module tt_um_crispy_vga (clk,
    ena,
    rst_n,
    ui_in,
    uio_in,
    uio_oe,
    uio_out,
    uo_out);
 input clk;
 input ena;
 input rst_n;
 input [7:0] ui_in;
 input [7:0] uio_in;
 output [7:0] uio_oe;
 output [7:0] uio_out;
 output [7:0] uo_out;

 wire _0000_;
 wire _0001_;
 wire _0002_;
 wire _0003_;
 wire _0004_;
 wire _0005_;
 wire _0006_;
 wire _0007_;
 wire _0008_;
 wire _0009_;
 wire _0010_;
 wire _0011_;
 wire _0012_;
 wire _0013_;
 wire _0014_;
 wire _0015_;
 wire _0016_;
 wire _0017_;
 wire _0018_;
 wire _0019_;
 wire _0020_;
 wire _0021_;
 wire _0022_;
 wire _0023_;
 wire _0024_;
 wire _0025_;
 wire _0026_;
 wire _0027_;
 wire _0028_;
 wire _0029_;
 wire _0030_;
 wire _0031_;
 wire _0032_;
 wire _0033_;
 wire _0034_;
 wire _0035_;
 wire _0036_;
 wire _0037_;
 wire _0038_;
 wire _0039_;
 wire _0040_;
 wire _0041_;
 wire _0042_;
 wire _0043_;
 wire _0044_;
 wire _0045_;
 wire _0046_;
 wire _0047_;
 wire _0048_;
 wire _0049_;
 wire _0050_;
 wire _0051_;
 wire _0052_;
 wire _0053_;
 wire _0054_;
 wire _0055_;
 wire _0056_;
 wire _0057_;
 wire _0058_;
 wire _0059_;
 wire _0060_;
 wire _0061_;
 wire _0062_;
 wire _0063_;
 wire _0064_;
 wire _0065_;
 wire _0066_;
 wire _0067_;
 wire _0068_;
 wire _0069_;
 wire _0070_;
 wire _0071_;
 wire _0072_;
 wire _0073_;
 wire _0074_;
 wire _0075_;
 wire _0076_;
 wire _0077_;
 wire _0078_;
 wire _0079_;
 wire _0080_;
 wire _0081_;
 wire _0082_;
 wire _0083_;
 wire _0084_;
 wire _0085_;
 wire _0086_;
 wire _0087_;
 wire _0088_;
 wire _0089_;
 wire _0090_;
 wire _0091_;
 wire _0092_;
 wire _0093_;
 wire _0094_;
 wire _0095_;
 wire _0096_;
 wire _0097_;
 wire _0098_;
 wire _0099_;
 wire _0100_;
 wire _0101_;
 wire _0102_;
 wire _0103_;
 wire _0104_;
 wire _0105_;
 wire _0106_;
 wire _0107_;
 wire _0108_;
 wire _0109_;
 wire _0110_;
 wire _0111_;
 wire _0112_;
 wire _0113_;
 wire _0114_;
 wire _0115_;
 wire _0116_;
 wire _0117_;
 wire _0118_;
 wire _0119_;
 wire _0120_;
 wire _0121_;
 wire _0122_;
 wire _0123_;
 wire _0124_;
 wire _0125_;
 wire _0126_;
 wire _0127_;
 wire _0128_;
 wire _0129_;
 wire _0130_;
 wire _0131_;
 wire _0132_;
 wire _0133_;
 wire _0134_;
 wire _0135_;
 wire _0136_;
 wire _0137_;
 wire _0138_;
 wire _0139_;
 wire _0140_;
 wire _0141_;
 wire _0142_;
 wire _0143_;
 wire _0144_;
 wire _0145_;
 wire _0146_;
 wire _0147_;
 wire _0148_;
 wire _0149_;
 wire _0150_;
 wire _0151_;
 wire _0152_;
 wire _0153_;
 wire _0154_;
 wire _0155_;
 wire _0156_;
 wire _0157_;
 wire _0158_;
 wire _0159_;
 wire _0160_;
 wire _0161_;
 wire _0162_;
 wire _0163_;
 wire _0164_;
 wire _0165_;
 wire _0166_;
 wire _0167_;
 wire _0168_;
 wire _0169_;
 wire _0170_;
 wire _0171_;
 wire _0172_;
 wire _0173_;
 wire _0174_;
 wire _0175_;
 wire _0176_;
 wire _0177_;
 wire _0178_;
 wire _0179_;
 wire _0180_;
 wire _0181_;
 wire _0182_;
 wire _0183_;
 wire _0184_;
 wire _0185_;
 wire _0186_;
 wire _0187_;
 wire _0188_;
 wire _0189_;
 wire _0190_;
 wire _0191_;
 wire _0192_;
 wire _0193_;
 wire _0194_;
 wire _0195_;
 wire _0196_;
 wire _0197_;
 wire _0198_;
 wire _0199_;
 wire _0200_;
 wire _0201_;
 wire _0202_;
 wire _0203_;
 wire _0204_;
 wire _0205_;
 wire _0206_;
 wire _0207_;
 wire _0208_;
 wire _0209_;
 wire _0210_;
 wire _0211_;
 wire _0212_;
 wire _0213_;
 wire _0214_;
 wire _0215_;
 wire _0216_;
 wire _0217_;
 wire _0218_;
 wire _0219_;
 wire _0220_;
 wire _0221_;
 wire _0222_;
 wire _0223_;
 wire _0224_;
 wire _0225_;
 wire _0226_;
 wire _0227_;
 wire _0228_;
 wire _0229_;
 wire _0230_;
 wire _0231_;
 wire _0232_;
 wire _0233_;
 wire _0234_;
 wire _0235_;
 wire _0236_;
 wire _0237_;
 wire _0238_;
 wire _0239_;
 wire _0240_;
 wire _0241_;
 wire _0242_;
 wire _0243_;
 wire _0244_;
 wire _0245_;
 wire _0246_;
 wire _0247_;
 wire _0248_;
 wire _0249_;
 wire _0250_;
 wire _0251_;
 wire _0252_;
 wire _0253_;
 wire _0254_;
 wire _0255_;
 wire _0256_;
 wire _0257_;
 wire _0258_;
 wire _0259_;
 wire _0260_;
 wire _0261_;
 wire _0262_;
 wire _0263_;
 wire _0264_;
 wire _0265_;
 wire _0266_;
 wire _0267_;
 wire _0268_;
 wire _0269_;
 wire _0270_;
 wire _0271_;
 wire _0272_;
 wire _0273_;
 wire _0274_;
 wire _0275_;
 wire _0276_;
 wire _0277_;
 wire _0278_;
 wire _0279_;
 wire _0280_;
 wire _0281_;
 wire _0282_;
 wire _0283_;
 wire _0284_;
 wire _0285_;
 wire _0286_;
 wire _0287_;
 wire _0288_;
 wire _0289_;
 wire _0290_;
 wire _0291_;
 wire _0292_;
 wire _0293_;
 wire _0294_;
 wire _0295_;
 wire _0296_;
 wire _0297_;
 wire _0298_;
 wire _0299_;
 wire _0300_;
 wire _0301_;
 wire _0302_;
 wire _0303_;
 wire _0304_;
 wire _0305_;
 wire _0306_;
 wire _0307_;
 wire _0308_;
 wire _0309_;
 wire _0310_;
 wire _0311_;
 wire _0312_;
 wire _0313_;
 wire _0314_;
 wire _0315_;
 wire _0316_;
 wire _0317_;
 wire _0318_;
 wire _0319_;
 wire _0320_;
 wire _0321_;
 wire _0322_;
 wire _0323_;
 wire _0324_;
 wire _0325_;
 wire _0326_;
 wire _0327_;
 wire _0328_;
 wire _0329_;
 wire _0330_;
 wire _0331_;
 wire _0332_;
 wire _0333_;
 wire _0334_;
 wire _0335_;
 wire _0336_;
 wire _0337_;
 wire _0338_;
 wire _0339_;
 wire _0340_;
 wire _0341_;
 wire _0342_;
 wire _0343_;
 wire _0344_;
 wire _0345_;
 wire _0346_;
 wire _0347_;
 wire _0348_;
 wire _0349_;
 wire _0350_;
 wire _0351_;
 wire _0352_;
 wire _0353_;
 wire _0354_;
 wire _0355_;
 wire _0356_;
 wire _0357_;
 wire _0358_;
 wire _0359_;
 wire _0360_;
 wire _0361_;
 wire _0362_;
 wire _0363_;
 wire _0364_;
 wire _0365_;
 wire _0366_;
 wire _0367_;
 wire _0368_;
 wire _0369_;
 wire _0370_;
 wire _0371_;
 wire _0372_;
 wire _0373_;
 wire _0374_;
 wire _0375_;
 wire _0376_;
 wire _0377_;
 wire _0378_;
 wire _0379_;
 wire _0380_;
 wire _0381_;
 wire _0382_;
 wire _0383_;
 wire _0384_;
 wire _0385_;
 wire _0386_;
 wire _0387_;
 wire _0388_;
 wire _0389_;
 wire _0390_;
 wire _0391_;
 wire _0392_;
 wire _0393_;
 wire _0394_;
 wire _0395_;
 wire _0396_;
 wire _0397_;
 wire _0398_;
 wire _0399_;
 wire _0400_;
 wire _0401_;
 wire _0402_;
 wire _0403_;
 wire _0404_;
 wire _0405_;
 wire _0406_;
 wire _0407_;
 wire _0408_;
 wire _0409_;
 wire _0410_;
 wire _0411_;
 wire _0412_;
 wire _0413_;
 wire _0414_;
 wire _0415_;
 wire _0416_;
 wire _0417_;
 wire _0418_;
 wire _0419_;
 wire _0420_;
 wire _0421_;
 wire _0422_;
 wire _0423_;
 wire _0424_;
 wire _0425_;
 wire _0426_;
 wire _0427_;
 wire _0428_;
 wire _0429_;
 wire _0430_;
 wire _0431_;
 wire _0432_;
 wire _0433_;
 wire _0434_;
 wire _0435_;
 wire _0436_;
 wire _0437_;
 wire _0438_;
 wire _0439_;
 wire _0440_;
 wire _0441_;
 wire _0442_;
 wire _0443_;
 wire _0444_;
 wire _0445_;
 wire _0446_;
 wire _0447_;
 wire _0448_;
 wire _0449_;
 wire _0450_;
 wire _0451_;
 wire _0452_;
 wire _0453_;
 wire _0454_;
 wire _0455_;
 wire _0456_;
 wire _0457_;
 wire _0458_;
 wire _0459_;
 wire _0460_;
 wire _0461_;
 wire _0462_;
 wire _0463_;
 wire _0464_;
 wire _0465_;
 wire _0466_;
 wire _0467_;
 wire _0468_;
 wire _0469_;
 wire _0470_;
 wire _0471_;
 wire _0472_;
 wire _0473_;
 wire _0474_;
 wire _0475_;
 wire _0476_;
 wire _0477_;
 wire _0478_;
 wire _0479_;
 wire _0480_;
 wire _0481_;
 wire _0482_;
 wire _0483_;
 wire _0484_;
 wire _0485_;
 wire _0486_;
 wire _0487_;
 wire _0488_;
 wire _0489_;
 wire _0490_;
 wire _0491_;
 wire _0492_;
 wire _0493_;
 wire _0494_;
 wire _0495_;
 wire _0496_;
 wire _0497_;
 wire _0498_;
 wire _0499_;
 wire _0500_;
 wire _0501_;
 wire _0502_;
 wire _0503_;
 wire _0504_;
 wire _0505_;
 wire _0506_;
 wire _0507_;
 wire _0508_;
 wire _0509_;
 wire _0510_;
 wire _0511_;
 wire _0512_;
 wire _0513_;
 wire _0514_;
 wire _0515_;
 wire _0516_;
 wire _0517_;
 wire _0518_;
 wire _0519_;
 wire _0520_;
 wire _0521_;
 wire _0522_;
 wire _0523_;
 wire _0524_;
 wire _0525_;
 wire _0526_;
 wire _0527_;
 wire _0528_;
 wire _0529_;
 wire _0530_;
 wire _0531_;
 wire _0532_;
 wire _0533_;
 wire _0534_;
 wire _0535_;
 wire _0536_;
 wire _0537_;
 wire _0538_;
 wire _0539_;
 wire _0540_;
 wire _0541_;
 wire _0542_;
 wire _0543_;
 wire _0544_;
 wire _0545_;
 wire _0546_;
 wire _0547_;
 wire _0548_;
 wire _0549_;
 wire _0550_;
 wire _0551_;
 wire _0552_;
 wire _0553_;
 wire _0554_;
 wire _0555_;
 wire _0556_;
 wire _0557_;
 wire _0558_;
 wire _0559_;
 wire _0560_;
 wire _0561_;
 wire _0562_;
 wire _0563_;
 wire _0564_;
 wire _0565_;
 wire _0566_;
 wire _0567_;
 wire _0568_;
 wire _0569_;
 wire _0570_;
 wire _0571_;
 wire _0572_;
 wire _0573_;
 wire _0574_;
 wire _0575_;
 wire _0576_;
 wire _0577_;
 wire _0578_;
 wire _0579_;
 wire _0580_;
 wire _0581_;
 wire _0582_;
 wire _0583_;
 wire _0584_;
 wire _0585_;
 wire _0586_;
 wire _0587_;
 wire _0588_;
 wire _0589_;
 wire _0590_;
 wire _0591_;
 wire _0592_;
 wire _0593_;
 wire _0594_;
 wire _0595_;
 wire _0596_;
 wire _0597_;
 wire _0598_;
 wire _0599_;
 wire _0600_;
 wire _0601_;
 wire _0602_;
 wire _0603_;
 wire _0604_;
 wire _0605_;
 wire _0606_;
 wire _0607_;
 wire _0608_;
 wire _0609_;
 wire _0610_;
 wire _0611_;
 wire _0612_;
 wire _0613_;
 wire _0614_;
 wire _0615_;
 wire _0616_;
 wire _0617_;
 wire _0618_;
 wire _0619_;
 wire _0620_;
 wire _0621_;
 wire _0622_;
 wire _0623_;
 wire _0624_;
 wire _0625_;
 wire _0626_;
 wire _0627_;
 wire _0628_;
 wire _0629_;
 wire _0630_;
 wire _0631_;
 wire _0632_;
 wire _0633_;
 wire _0634_;
 wire _0635_;
 wire _0636_;
 wire _0637_;
 wire _0638_;
 wire _0639_;
 wire _0640_;
 wire _0641_;
 wire _0642_;
 wire _0643_;
 wire _0644_;
 wire _0645_;
 wire _0646_;
 wire _0647_;
 wire _0648_;
 wire _0649_;
 wire _0650_;
 wire _0651_;
 wire _0652_;
 wire _0653_;
 wire _0654_;
 wire _0655_;
 wire _0656_;
 wire _0657_;
 wire _0658_;
 wire _0659_;
 wire _0660_;
 wire _0661_;
 wire _0662_;
 wire _0663_;
 wire _0664_;
 wire _0665_;
 wire _0666_;
 wire _0667_;
 wire _0668_;
 wire _0669_;
 wire _0670_;
 wire _0671_;
 wire _0672_;
 wire _0673_;
 wire _0674_;
 wire _0675_;
 wire _0676_;
 wire _0677_;
 wire _0678_;
 wire _0679_;
 wire _0680_;
 wire _0681_;
 wire _0682_;
 wire _0683_;
 wire _0684_;
 wire _0685_;
 wire _0686_;
 wire _0687_;
 wire _0688_;
 wire _0689_;
 wire _0690_;
 wire _0691_;
 wire _0692_;
 wire _0693_;
 wire _0694_;
 wire _0695_;
 wire _0696_;
 wire _0697_;
 wire _0698_;
 wire _0699_;
 wire _0700_;
 wire _0701_;
 wire _0702_;
 wire _0703_;
 wire _0704_;
 wire _0705_;
 wire _0706_;
 wire _0707_;
 wire _0708_;
 wire _0709_;
 wire _0710_;
 wire _0711_;
 wire _0712_;
 wire _0713_;
 wire _0714_;
 wire _0715_;
 wire _0716_;
 wire _0717_;
 wire _0718_;
 wire _0719_;
 wire _0720_;
 wire _0721_;
 wire _0722_;
 wire _0723_;
 wire _0724_;
 wire _0725_;
 wire _0726_;
 wire _0727_;
 wire _0728_;
 wire _0729_;
 wire _0730_;
 wire _0731_;
 wire _0732_;
 wire _0733_;
 wire _0734_;
 wire _0735_;
 wire _0736_;
 wire _0737_;
 wire _0738_;
 wire _0739_;
 wire _0740_;
 wire _0741_;
 wire _0742_;
 wire _0743_;
 wire _0744_;
 wire _0745_;
 wire _0746_;
 wire _0747_;
 wire _0748_;
 wire _0749_;
 wire _0750_;
 wire _0751_;
 wire _0752_;
 wire _0753_;
 wire _0754_;
 wire _0755_;
 wire _0756_;
 wire _0757_;
 wire _0758_;
 wire _0759_;
 wire _0760_;
 wire _0761_;
 wire _0762_;
 wire _0763_;
 wire _0764_;
 wire _0765_;
 wire _0766_;
 wire _0767_;
 wire _0768_;
 wire _0769_;
 wire _0770_;
 wire _0771_;
 wire _0772_;
 wire _0773_;
 wire _0774_;
 wire _0775_;
 wire _0776_;
 wire _0777_;
 wire _0778_;
 wire _0779_;
 wire _0780_;
 wire _0781_;
 wire _0782_;
 wire _0783_;
 wire _0784_;
 wire _0785_;
 wire _0786_;
 wire _0787_;
 wire _0788_;
 wire _0789_;
 wire _0790_;
 wire _0791_;
 wire _0792_;
 wire _0793_;
 wire _0794_;
 wire _0795_;
 wire _0796_;
 wire _0797_;
 wire _0798_;
 wire _0799_;
 wire _0800_;
 wire _0801_;
 wire _0802_;
 wire _0803_;
 wire _0804_;
 wire _0805_;
 wire _0806_;
 wire _0807_;
 wire _0808_;
 wire _0809_;
 wire _0810_;
 wire _0811_;
 wire _0812_;
 wire _0813_;
 wire _0814_;
 wire _0815_;
 wire _0816_;
 wire _0817_;
 wire _0818_;
 wire _0819_;
 wire _0820_;
 wire _0821_;
 wire _0822_;
 wire _0823_;
 wire _0824_;
 wire _0825_;
 wire _0826_;
 wire _0827_;
 wire _0828_;
 wire _0829_;
 wire _0830_;
 wire _0831_;
 wire _0832_;
 wire _0833_;
 wire _0834_;
 wire _0835_;
 wire _0836_;
 wire _0837_;
 wire _0838_;
 wire _0839_;
 wire _0840_;
 wire _0841_;
 wire _0842_;
 wire _0843_;
 wire _0844_;
 wire _0845_;
 wire _0846_;
 wire _0847_;
 wire _0848_;
 wire _0849_;
 wire _0850_;
 wire _0851_;
 wire _0852_;
 wire _0853_;
 wire _0854_;
 wire _0855_;
 wire _0856_;
 wire _0857_;
 wire _0858_;
 wire _0859_;
 wire _0860_;
 wire _0861_;
 wire _0862_;
 wire _0863_;
 wire _0864_;
 wire _0865_;
 wire _0866_;
 wire _0867_;
 wire _0868_;
 wire _0869_;
 wire _0870_;
 wire _0871_;
 wire _0872_;
 wire _0873_;
 wire _0874_;
 wire _0875_;
 wire _0876_;
 wire _0877_;
 wire _0878_;
 wire _0879_;
 wire _0880_;
 wire _0881_;
 wire _0882_;
 wire _0883_;
 wire _0884_;
 wire _0885_;
 wire _0886_;
 wire _0887_;
 wire _0888_;
 wire _0889_;
 wire _0890_;
 wire _0891_;
 wire _0892_;
 wire _0893_;
 wire _0894_;
 wire _0895_;
 wire _0896_;
 wire _0897_;
 wire _0898_;
 wire _0899_;
 wire _0900_;
 wire _0901_;
 wire _0902_;
 wire _0903_;
 wire _0904_;
 wire _0905_;
 wire _0906_;
 wire _0907_;
 wire _0908_;
 wire _0909_;
 wire _0910_;
 wire _0911_;
 wire _0912_;
 wire _0913_;
 wire _0914_;
 wire _0915_;
 wire _0916_;
 wire _0917_;
 wire _0918_;
 wire _0919_;
 wire _0920_;
 wire _0921_;
 wire _0922_;
 wire _0923_;
 wire _0924_;
 wire _0925_;
 wire _0926_;
 wire _0927_;
 wire _0928_;
 wire _0929_;
 wire _0930_;
 wire _0931_;
 wire _0932_;
 wire _0933_;
 wire _0934_;
 wire _0935_;
 wire _0936_;
 wire _0937_;
 wire _0938_;
 wire _0939_;
 wire _0940_;
 wire _0941_;
 wire _0942_;
 wire _0943_;
 wire _0944_;
 wire _0945_;
 wire _0946_;
 wire _0947_;
 wire _0948_;
 wire _0949_;
 wire _0950_;
 wire _0951_;
 wire _0952_;
 wire clknet_0_clk;
 wire net93;
 wire \pcg_out[0] ;
 wire \pcg_out[1] ;
 wire \pcg_out[2] ;
 wire \pcg_out[3] ;
 wire \pcg_out[4] ;
 wire \pcg_out[5] ;
 wire \pcg_out[6] ;
 wire \pcg_out[7] ;
 wire \state[0] ;
 wire \state[10] ;
 wire \state[11] ;
 wire \state[12] ;
 wire \state[13] ;
 wire \state[14] ;
 wire \state[15] ;
 wire \state[1] ;
 wire \state[2] ;
 wire \state[3] ;
 wire \state[4] ;
 wire \state[5] ;
 wire \state[6] ;
 wire \state[7] ;
 wire \state[8] ;
 wire \state[9] ;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire clknet_2_0__leaf_clk;
 wire clknet_2_1__leaf_clk;
 wire clknet_2_2__leaf_clk;
 wire clknet_2_3__leaf_clk;

 sg13g2_inv_1 _0955_ (.Y(_0706_),
    .A(net1));
 sg13g2_buf_1 _0956_ (.A(_0706_),
    .X(_0717_));
 sg13g2_buf_2 _0957_ (.A(\state[13] ),
    .X(_0728_));
 sg13g2_inv_2 _0958_ (.Y(_0738_),
    .A(_0728_));
 sg13g2_buf_2 _0959_ (.A(\state[15] ),
    .X(_0749_));
 sg13g2_buf_1 _0960_ (.A(_0749_),
    .X(_0760_));
 sg13g2_buf_1 _0961_ (.A(\state[5] ),
    .X(_0770_));
 sg13g2_buf_1 _0962_ (.A(\state[9] ),
    .X(_0781_));
 sg13g2_buf_1 _0963_ (.A(\state[11] ),
    .X(_0792_));
 sg13g2_buf_8 _0964_ (.A(\state[14] ),
    .X(_0802_));
 sg13g2_mux2_1 _0965_ (.A0(_0781_),
    .A1(net76),
    .S(_0802_),
    .X(_0813_));
 sg13g2_nor4_1 _0966_ (.A(_0738_),
    .B(_0760_),
    .C(_0770_),
    .D(_0813_),
    .Y(_0824_));
 sg13g2_nor2b_1 _0967_ (.A(_0749_),
    .B_N(_0728_),
    .Y(_0834_));
 sg13g2_and3_1 _0968_ (.X(_0845_),
    .A(_0770_),
    .B(_0834_),
    .C(_0813_));
 sg13g2_inv_1 _0969_ (.Y(_0856_),
    .A(_0749_));
 sg13g2_inv_1 _0970_ (.Y(_0866_),
    .A(_0770_));
 sg13g2_buf_1 _0971_ (.A(_0728_),
    .X(_0877_));
 sg13g2_buf_1 _0972_ (.A(\state[12] ),
    .X(_0888_));
 sg13g2_buf_8 _0973_ (.A(_0802_),
    .X(_0899_));
 sg13g2_nor3_1 _0974_ (.A(net67),
    .B(net75),
    .C(net66),
    .Y(_0907_));
 sg13g2_nor3_1 _0975_ (.A(_0856_),
    .B(net68),
    .C(_0907_),
    .Y(_0914_));
 sg13g2_buf_1 _0976_ (.A(_0728_),
    .X(_0922_));
 sg13g2_or2_1 _0977_ (.X(_0028_),
    .B(_0802_),
    .A(net75));
 sg13g2_buf_1 _0978_ (.A(_0028_),
    .X(_0035_));
 sg13g2_nor4_1 _0979_ (.A(net65),
    .B(_0856_),
    .C(_0770_),
    .D(_0035_),
    .Y(_0037_));
 sg13g2_nor4_2 _0980_ (.A(_0824_),
    .B(_0845_),
    .C(_0914_),
    .Y(_0038_),
    .D(_0037_));
 sg13g2_buf_2 _0981_ (.A(\state[8] ),
    .X(_0039_));
 sg13g2_mux2_1 _0982_ (.A0(_0039_),
    .A1(\state[10] ),
    .S(_0802_),
    .X(_0040_));
 sg13g2_buf_1 _0983_ (.A(_0040_),
    .X(_0041_));
 sg13g2_buf_1 _0984_ (.A(_0749_),
    .X(_0042_));
 sg13g2_nor3_1 _0985_ (.A(net65),
    .B(net64),
    .C(_0866_),
    .Y(_0043_));
 sg13g2_nor4_1 _0986_ (.A(net65),
    .B(net64),
    .C(_0770_),
    .D(_0041_),
    .Y(_0044_));
 sg13g2_a21oi_2 _0987_ (.B1(_0044_),
    .Y(_0045_),
    .A2(_0043_),
    .A1(_0041_));
 sg13g2_nand2_1 _0988_ (.Y(_0046_),
    .A(_0038_),
    .B(_0045_));
 sg13g2_buf_1 _0989_ (.A(_0046_),
    .X(_0047_));
 sg13g2_buf_1 _0990_ (.A(\state[6] ),
    .X(_0048_));
 sg13g2_buf_1 _0991_ (.A(\state[7] ),
    .X(_0049_));
 sg13g2_mux2_1 _0992_ (.A0(_0048_),
    .A1(net74),
    .S(_0728_),
    .X(_0050_));
 sg13g2_buf_1 _0993_ (.A(net66),
    .X(_0051_));
 sg13g2_nand2b_1 _0994_ (.Y(_0052_),
    .B(_0051_),
    .A_N(net69));
 sg13g2_nor2_1 _0995_ (.A(_0050_),
    .B(_0052_),
    .Y(_0053_));
 sg13g2_mux2_1 _0996_ (.A0(\state[4] ),
    .A1(_0770_),
    .S(_0877_),
    .X(_0054_));
 sg13g2_nor2_2 _0997_ (.A(net66),
    .B(_0749_),
    .Y(_0055_));
 sg13g2_nor2b_1 _0998_ (.A(_0054_),
    .B_N(_0055_),
    .Y(_0056_));
 sg13g2_nand2_1 _0999_ (.Y(_0057_),
    .A(net65),
    .B(net69));
 sg13g2_nor2_1 _1000_ (.A(_0813_),
    .B(_0057_),
    .Y(_0058_));
 sg13g2_nand2b_1 _1001_ (.Y(_0059_),
    .B(_0042_),
    .A_N(net65));
 sg13g2_nor2_1 _1002_ (.A(_0041_),
    .B(_0059_),
    .Y(_0060_));
 sg13g2_nor4_2 _1003_ (.A(_0053_),
    .B(_0056_),
    .C(_0058_),
    .Y(_0061_),
    .D(_0060_));
 sg13g2_xnor2_1 _1004_ (.Y(_0062_),
    .A(_0001_),
    .B(_0061_));
 sg13g2_buf_1 _1005_ (.A(\state[2] ),
    .X(_0063_));
 sg13g2_inv_1 _1006_ (.Y(_0064_),
    .A(_0063_));
 sg13g2_nor2b_1 _1007_ (.A(net67),
    .B_N(net69),
    .Y(_0065_));
 sg13g2_and2_1 _1008_ (.A(net67),
    .B(net69),
    .X(_0066_));
 sg13g2_mux2_1 _1009_ (.A0(\state[10] ),
    .A1(net75),
    .S(_0802_),
    .X(_0067_));
 sg13g2_a22oi_1 _1010_ (.Y(_0068_),
    .B1(_0066_),
    .B2(_0067_),
    .A2(_0813_),
    .A1(_0065_));
 sg13g2_mux2_1 _1011_ (.A0(_0770_),
    .A1(_0048_),
    .S(_0728_),
    .X(_0069_));
 sg13g2_mux2_1 _1012_ (.A0(_0049_),
    .A1(_0039_),
    .S(net67),
    .X(_0070_));
 sg13g2_nor2b_1 _1013_ (.A(_0749_),
    .B_N(net66),
    .Y(_0071_));
 sg13g2_a22oi_1 _1014_ (.Y(_0072_),
    .B1(_0070_),
    .B2(_0071_),
    .A2(_0069_),
    .A1(_0055_));
 sg13g2_nand2_1 _1015_ (.Y(_0073_),
    .A(_0068_),
    .B(_0072_));
 sg13g2_xnor2_1 _1016_ (.Y(_0074_),
    .A(_0064_),
    .B(_0073_));
 sg13g2_buf_2 _1017_ (.A(_0074_),
    .X(_0075_));
 sg13g2_xnor2_1 _1018_ (.Y(_0076_),
    .A(_0062_),
    .B(_0075_));
 sg13g2_xnor2_1 _1019_ (.Y(_0077_),
    .A(net46),
    .B(_0076_));
 sg13g2_buf_2 _1020_ (.A(_0077_),
    .X(_0078_));
 sg13g2_nor2_1 _1021_ (.A(net67),
    .B(_0067_),
    .Y(_0079_));
 sg13g2_or2_1 _1022_ (.X(_0080_),
    .B(\state[11] ),
    .A(_0899_));
 sg13g2_o21ai_1 _1023_ (.B1(net69),
    .Y(_0081_),
    .A1(_0738_),
    .A2(_0080_));
 sg13g2_mux2_1 _1024_ (.A0(_0039_),
    .A1(_0781_),
    .S(_0728_),
    .X(_0082_));
 sg13g2_a22oi_1 _1025_ (.Y(_0083_),
    .B1(_0071_),
    .B2(_0082_),
    .A2(_0055_),
    .A1(_0050_));
 sg13g2_o21ai_1 _1026_ (.B1(_0083_),
    .Y(_0084_),
    .A1(_0079_),
    .A2(_0081_));
 sg13g2_xnor2_1 _1027_ (.Y(_0085_),
    .A(_0002_),
    .B(_0084_));
 sg13g2_mux2_1 _1028_ (.A0(_0049_),
    .A1(_0781_),
    .S(net66),
    .X(_0086_));
 sg13g2_nor2b_1 _1029_ (.A(net49),
    .B_N(net76),
    .Y(_0087_));
 sg13g2_mux4_1 _1030_ (.S0(_0738_),
    .A0(_0041_),
    .A1(_0086_),
    .A2(_0035_),
    .A3(_0087_),
    .S1(_0042_),
    .X(_0088_));
 sg13g2_xor2_1 _1031_ (.B(_0088_),
    .A(\state[4] ),
    .X(_0089_));
 sg13g2_buf_1 _1032_ (.A(_0089_),
    .X(_0090_));
 sg13g2_nand2b_1 _1033_ (.Y(_0091_),
    .B(net45),
    .A_N(_0085_));
 sg13g2_nor2b_1 _1034_ (.A(net76),
    .B_N(net67),
    .Y(_0092_));
 sg13g2_nand3_1 _1035_ (.B(_0055_),
    .C(_0092_),
    .A(net74),
    .Y(_0093_));
 sg13g2_buf_1 _1036_ (.A(\state[10] ),
    .X(_0094_));
 sg13g2_nor2_1 _1037_ (.A(net66),
    .B(_0094_),
    .Y(_0095_));
 sg13g2_nor2b_1 _1038_ (.A(_0922_),
    .B_N(net74),
    .Y(_0096_));
 sg13g2_o21ai_1 _1039_ (.B1(_0096_),
    .Y(_0097_),
    .A1(net64),
    .A2(_0095_));
 sg13g2_nor2_1 _1040_ (.A(_0922_),
    .B(net75),
    .Y(_0098_));
 sg13g2_and2_1 _1041_ (.A(net49),
    .B(net74),
    .X(_0099_));
 sg13g2_o21ai_1 _1042_ (.B1(_0099_),
    .Y(_0100_),
    .A1(net64),
    .A2(_0098_));
 sg13g2_and3_1 _1043_ (.X(_0101_),
    .A(_0093_),
    .B(_0097_),
    .C(_0100_));
 sg13g2_buf_1 _1044_ (.A(_0101_),
    .X(_0102_));
 sg13g2_o21ai_1 _1045_ (.B1(_0738_),
    .Y(_0103_),
    .A1(net64),
    .A2(_0095_));
 sg13g2_o21ai_1 _1046_ (.B1(net49),
    .Y(_0104_),
    .A1(net64),
    .A2(_0098_));
 sg13g2_a21oi_1 _1047_ (.A1(_0055_),
    .A2(_0092_),
    .Y(_0105_),
    .B1(net74));
 sg13g2_nand3_1 _1048_ (.B(_0104_),
    .C(_0105_),
    .A(_0103_),
    .Y(_0106_));
 sg13g2_nand2_2 _1049_ (.Y(_0107_),
    .A(_0102_),
    .B(_0106_));
 sg13g2_buf_1 _1050_ (.A(_0107_),
    .X(_0108_));
 sg13g2_buf_1 _1051_ (.A(\state[4] ),
    .X(_0109_));
 sg13g2_xnor2_1 _1052_ (.Y(_0110_),
    .A(_0109_),
    .B(_0088_));
 sg13g2_buf_1 _1053_ (.A(_0110_),
    .X(_0111_));
 sg13g2_buf_1 _1054_ (.A(_0085_),
    .X(_0112_));
 sg13g2_nand3_1 _1055_ (.B(net43),
    .C(_0107_),
    .A(net44),
    .Y(_0113_));
 sg13g2_o21ai_1 _1056_ (.B1(_0113_),
    .Y(_0114_),
    .A1(_0091_),
    .A2(net32));
 sg13g2_buf_2 _1057_ (.A(_0003_),
    .X(_0115_));
 sg13g2_nor2_1 _1058_ (.A(_0052_),
    .B(_0069_),
    .Y(_0116_));
 sg13g2_mux2_1 _1059_ (.A0(\state[3] ),
    .A1(\state[4] ),
    .S(_0877_),
    .X(_0117_));
 sg13g2_nor2b_1 _1060_ (.A(_0117_),
    .B_N(_0055_),
    .Y(_0118_));
 sg13g2_nor2_1 _1061_ (.A(_0041_),
    .B(_0057_),
    .Y(_0119_));
 sg13g2_nor2_1 _1062_ (.A(_0086_),
    .B(_0059_),
    .Y(_0120_));
 sg13g2_nor4_2 _1063_ (.A(_0116_),
    .B(_0118_),
    .C(_0119_),
    .Y(_0121_),
    .D(_0120_));
 sg13g2_xor2_1 _1064_ (.B(_0121_),
    .A(_0115_),
    .X(_0122_));
 sg13g2_buf_1 _1065_ (.A(_0122_),
    .X(_0123_));
 sg13g2_buf_1 _1066_ (.A(\state[1] ),
    .X(_0124_));
 sg13g2_xnor2_1 _1067_ (.Y(_0125_),
    .A(_0124_),
    .B(_0061_));
 sg13g2_buf_2 _1068_ (.A(_0125_),
    .X(_0126_));
 sg13g2_nor2_1 _1069_ (.A(net39),
    .B(_0126_),
    .Y(_0127_));
 sg13g2_inv_2 _1070_ (.Y(_0128_),
    .A(_0039_));
 sg13g2_buf_1 _1071_ (.A(net65),
    .X(_0129_));
 sg13g2_nand3_1 _1072_ (.B(_0856_),
    .C(_0035_),
    .A(net48),
    .Y(_0130_));
 sg13g2_nor2_1 _1073_ (.A(_0749_),
    .B(net76),
    .Y(_0131_));
 sg13g2_nor2_1 _1074_ (.A(_0728_),
    .B(_0899_),
    .Y(_0132_));
 sg13g2_nand2b_1 _1075_ (.Y(_0133_),
    .B(_0132_),
    .A_N(_0131_));
 sg13g2_nand3_1 _1076_ (.B(_0130_),
    .C(_0133_),
    .A(_0128_),
    .Y(_0134_));
 sg13g2_a21o_1 _1077_ (.A2(_0133_),
    .A1(_0130_),
    .B1(_0128_),
    .X(_0135_));
 sg13g2_buf_1 _1078_ (.A(_0135_),
    .X(_0136_));
 sg13g2_nand2_1 _1079_ (.Y(_0137_),
    .A(_0134_),
    .B(_0136_));
 sg13g2_xnor2_1 _1080_ (.Y(_0138_),
    .A(_0127_),
    .B(_0137_));
 sg13g2_xnor2_1 _1081_ (.Y(_0139_),
    .A(_0114_),
    .B(_0138_));
 sg13g2_xnor2_1 _1082_ (.Y(_0140_),
    .A(_0078_),
    .B(_0139_));
 sg13g2_xor2_1 _1083_ (.B(_0084_),
    .A(\state[3] ),
    .X(_0141_));
 sg13g2_inv_1 _1084_ (.Y(_0142_),
    .A(_0000_));
 sg13g2_a21o_1 _1085_ (.A2(_0072_),
    .A1(_0068_),
    .B1(_0142_),
    .X(_0143_));
 sg13g2_nand3_1 _1086_ (.B(_0068_),
    .C(_0072_),
    .A(_0142_),
    .Y(_0144_));
 sg13g2_inv_2 _1087_ (.Y(_0145_),
    .A(\state[10] ));
 sg13g2_buf_1 _1088_ (.A(_0048_),
    .X(_0146_));
 sg13g2_nor4_1 _1089_ (.A(net49),
    .B(_0760_),
    .C(_0145_),
    .D(net62),
    .Y(_0147_));
 sg13g2_and2_1 _1090_ (.A(net65),
    .B(net49),
    .X(_0148_));
 sg13g2_nor2_1 _1091_ (.A(net69),
    .B(_0048_),
    .Y(_0149_));
 sg13g2_mux2_1 _1092_ (.A0(net62),
    .A1(_0149_),
    .S(_0888_),
    .X(_0150_));
 sg13g2_nand2b_1 _1093_ (.Y(_0151_),
    .B(net67),
    .A_N(net66));
 sg13g2_nand2b_1 _1094_ (.Y(_0152_),
    .B(net62),
    .A_N(net73));
 sg13g2_nand3_1 _1095_ (.B(net69),
    .C(net62),
    .A(net65),
    .Y(_0153_));
 sg13g2_o21ai_1 _1096_ (.B1(_0153_),
    .Y(_0154_),
    .A1(_0151_),
    .A2(_0152_));
 sg13g2_a221oi_1 _1097_ (.B2(_0150_),
    .C1(_0154_),
    .B1(_0148_),
    .A1(net48),
    .Y(_0155_),
    .A2(_0147_));
 sg13g2_buf_2 _1098_ (.A(_0155_),
    .X(_0156_));
 sg13g2_inv_1 _1099_ (.Y(_0157_),
    .A(_0048_));
 sg13g2_nand4_1 _1100_ (.B(_0781_),
    .C(_0157_),
    .A(_0856_),
    .Y(_0158_),
    .D(_0132_));
 sg13g2_nor2b_1 _1101_ (.A(net62),
    .B_N(_0749_),
    .Y(_0159_));
 sg13g2_nor2b_1 _1102_ (.A(net62),
    .B_N(net76),
    .Y(_0160_));
 sg13g2_nor2b_1 _1103_ (.A(net67),
    .B_N(net66),
    .Y(_0161_));
 sg13g2_o21ai_1 _1104_ (.B1(_0161_),
    .Y(_0162_),
    .A1(_0159_),
    .A2(_0160_));
 sg13g2_nand3_1 _1105_ (.B(_0131_),
    .C(_0161_),
    .A(net62),
    .Y(_0163_));
 sg13g2_nor2b_1 _1106_ (.A(_0781_),
    .B_N(_0048_),
    .Y(_0164_));
 sg13g2_nor2b_1 _1107_ (.A(_0051_),
    .B_N(net69),
    .Y(_0165_));
 sg13g2_a22oi_1 _1108_ (.Y(_0166_),
    .B1(_0165_),
    .B2(net62),
    .A2(_0164_),
    .A1(_0132_));
 sg13g2_and4_1 _1109_ (.A(_0158_),
    .B(_0162_),
    .C(_0163_),
    .D(_0166_),
    .X(_0167_));
 sg13g2_buf_2 _1110_ (.A(_0167_),
    .X(_0168_));
 sg13g2_nand4_1 _1111_ (.B(_0144_),
    .C(_0156_),
    .A(_0143_),
    .Y(_0169_),
    .D(_0168_));
 sg13g2_a22oi_1 _1112_ (.Y(_0170_),
    .B1(_0156_),
    .B2(_0168_),
    .A2(_0144_),
    .A1(_0143_));
 sg13g2_a21o_1 _1113_ (.A2(_0169_),
    .A1(_0141_),
    .B1(_0170_),
    .X(_0171_));
 sg13g2_buf_1 _1114_ (.A(_0171_),
    .X(_0172_));
 sg13g2_xnor2_1 _1115_ (.Y(_0173_),
    .A(_0115_),
    .B(_0121_));
 sg13g2_buf_1 _1116_ (.A(_0173_),
    .X(_0174_));
 sg13g2_xnor2_1 _1117_ (.Y(_0175_),
    .A(net38),
    .B(_0126_));
 sg13g2_xnor2_1 _1118_ (.Y(_0176_),
    .A(_0089_),
    .B(_0085_));
 sg13g2_xnor2_1 _1119_ (.Y(_0177_),
    .A(net32),
    .B(_0176_));
 sg13g2_a21o_1 _1120_ (.A2(_0175_),
    .A1(_0172_),
    .B1(_0177_),
    .X(_0178_));
 sg13g2_o21ai_1 _1121_ (.B1(_0178_),
    .Y(_0179_),
    .A1(_0172_),
    .A2(_0175_));
 sg13g2_xnor2_1 _1122_ (.Y(_0180_),
    .A(_0140_),
    .B(_0179_));
 sg13g2_buf_1 _1123_ (.A(net44),
    .X(_0181_));
 sg13g2_buf_1 _1124_ (.A(_0126_),
    .X(_0182_));
 sg13g2_nor4_1 _1125_ (.A(net37),
    .B(_0078_),
    .C(net38),
    .D(net31),
    .Y(_0183_));
 sg13g2_buf_1 _1126_ (.A(_0141_),
    .X(_0184_));
 sg13g2_nand2b_1 _1127_ (.Y(_0185_),
    .B(net42),
    .A_N(net31));
 sg13g2_buf_1 _1128_ (.A(\state[3] ),
    .X(_0186_));
 sg13g2_xnor2_1 _1129_ (.Y(_0187_),
    .A(_0186_),
    .B(_0084_));
 sg13g2_a21o_1 _1130_ (.A2(_0187_),
    .A1(net31),
    .B1(_0078_),
    .X(_0188_));
 sg13g2_a221oi_1 _1131_ (.B2(net37),
    .C1(net39),
    .B1(_0188_),
    .A1(_0078_),
    .Y(_0189_),
    .A2(_0185_));
 sg13g2_nand2_1 _1132_ (.Y(_0190_),
    .A(_0156_),
    .B(_0168_));
 sg13g2_buf_1 _1133_ (.A(_0190_),
    .X(_0191_));
 sg13g2_xnor2_1 _1134_ (.Y(_0192_),
    .A(_0191_),
    .B(_0141_));
 sg13g2_nand2_2 _1135_ (.Y(_0193_),
    .A(_0143_),
    .B(_0144_));
 sg13g2_buf_1 _1136_ (.A(_0047_),
    .X(_0194_));
 sg13g2_buf_1 _1137_ (.A(_0062_),
    .X(_0195_));
 sg13g2_xnor2_1 _1138_ (.Y(_0196_),
    .A(_0063_),
    .B(_0073_));
 sg13g2_nor2_1 _1139_ (.A(net46),
    .B(_0196_),
    .Y(_0197_));
 sg13g2_a21oi_1 _1140_ (.A1(net36),
    .A2(net35),
    .Y(_0198_),
    .B1(_0197_));
 sg13g2_nor4_1 _1141_ (.A(net46),
    .B(_0195_),
    .C(_0196_),
    .D(_0193_),
    .Y(_0199_));
 sg13g2_and2_1 _1142_ (.A(_0038_),
    .B(_0045_),
    .X(_0200_));
 sg13g2_buf_2 _1143_ (.A(_0200_),
    .X(_0201_));
 sg13g2_and3_1 _1144_ (.X(_0202_),
    .A(_0201_),
    .B(_0062_),
    .C(_0196_));
 sg13g2_or2_1 _1145_ (.X(_0203_),
    .B(_0202_),
    .A(_0199_));
 sg13g2_a21oi_1 _1146_ (.A1(_0193_),
    .A2(_0198_),
    .Y(_0204_),
    .B1(_0203_));
 sg13g2_xnor2_1 _1147_ (.Y(_0205_),
    .A(_0192_),
    .B(_0204_));
 sg13g2_mux2_1 _1148_ (.A0(_0183_),
    .A1(_0189_),
    .S(_0205_),
    .X(_0206_));
 sg13g2_buf_1 _1149_ (.A(_0201_),
    .X(_0207_));
 sg13g2_nand4_1 _1150_ (.B(_0075_),
    .C(_0193_),
    .A(_0207_),
    .Y(_0208_),
    .D(_0192_));
 sg13g2_and2_1 _1151_ (.A(_0156_),
    .B(_0168_),
    .X(_0209_));
 sg13g2_buf_1 _1152_ (.A(_0209_),
    .X(_0210_));
 sg13g2_xnor2_1 _1153_ (.Y(_0211_),
    .A(_0210_),
    .B(net42));
 sg13g2_nand2_1 _1154_ (.Y(_0212_),
    .A(_0211_),
    .B(_0202_));
 sg13g2_nor4_1 _1155_ (.A(_0047_),
    .B(_0195_),
    .C(_0196_),
    .D(net39),
    .Y(_0213_));
 sg13g2_a221oi_1 _1156_ (.B2(net38),
    .C1(_0213_),
    .B1(_0202_),
    .A1(_0211_),
    .Y(_0214_),
    .A2(_0199_));
 sg13g2_nand3_1 _1157_ (.B(_0212_),
    .C(_0214_),
    .A(_0208_),
    .Y(_0215_));
 sg13g2_and2_1 _1158_ (.A(_0143_),
    .B(_0144_),
    .X(_0216_));
 sg13g2_buf_2 _1159_ (.A(_0216_),
    .X(_0217_));
 sg13g2_nor2_2 _1160_ (.A(_0062_),
    .B(_0217_),
    .Y(_0218_));
 sg13g2_mux2_1 _1161_ (.A0(_0217_),
    .A1(_0218_),
    .S(_0211_),
    .X(_0219_));
 sg13g2_a21oi_1 _1162_ (.A1(net35),
    .A2(_0192_),
    .Y(_0220_),
    .B1(net38));
 sg13g2_nor2_1 _1163_ (.A(_0219_),
    .B(_0220_),
    .Y(_0221_));
 sg13g2_nor2_2 _1164_ (.A(_0215_),
    .B(_0221_),
    .Y(_0222_));
 sg13g2_xnor2_1 _1165_ (.Y(_0223_),
    .A(_0172_),
    .B(_0175_));
 sg13g2_xor2_1 _1166_ (.B(_0223_),
    .A(_0177_),
    .X(_0224_));
 sg13g2_and4_1 _1167_ (.A(_0174_),
    .B(_0193_),
    .C(_0192_),
    .D(_0202_),
    .X(_0225_));
 sg13g2_buf_1 _1168_ (.A(_0225_),
    .X(_0226_));
 sg13g2_inv_1 _1169_ (.Y(_0227_),
    .A(_0226_));
 sg13g2_nand2_1 _1170_ (.Y(_0228_),
    .A(_0224_),
    .B(_0227_));
 sg13g2_nor2b_1 _1171_ (.A(_0222_),
    .B_N(_0228_),
    .Y(_0229_));
 sg13g2_nand2_1 _1172_ (.Y(_0230_),
    .A(_0224_),
    .B(_0222_));
 sg13g2_o21ai_1 _1173_ (.B1(_0230_),
    .Y(_0231_),
    .A1(_0206_),
    .A2(_0229_));
 sg13g2_xnor2_1 _1174_ (.Y(_0232_),
    .A(_0180_),
    .B(_0231_));
 sg13g2_nor2_1 _1175_ (.A(net77),
    .B(_0232_),
    .Y(_0004_));
 sg13g2_buf_1 _1176_ (.A(net1),
    .X(_0233_));
 sg13g2_buf_1 _1177_ (.A(_0137_),
    .X(_0234_));
 sg13g2_nor2_1 _1178_ (.A(net44),
    .B(net33),
    .Y(_0235_));
 sg13g2_and2_1 _1179_ (.A(_0134_),
    .B(_0136_),
    .X(_0236_));
 sg13g2_buf_2 _1180_ (.A(_0236_),
    .X(_0237_));
 sg13g2_nand3_1 _1181_ (.B(_0038_),
    .C(_0045_),
    .A(net44),
    .Y(_0238_));
 sg13g2_nor2_1 _1182_ (.A(_0237_),
    .B(_0238_),
    .Y(_0239_));
 sg13g2_a21o_1 _1183_ (.A2(_0235_),
    .A1(net36),
    .B1(_0239_),
    .X(_0240_));
 sg13g2_buf_1 _1184_ (.A(_0781_),
    .X(_0241_));
 sg13g2_inv_2 _1185_ (.Y(_0242_),
    .A(net61));
 sg13g2_or3_1 _1186_ (.A(net64),
    .B(_0907_),
    .C(_0148_),
    .X(_0243_));
 sg13g2_xnor2_1 _1187_ (.Y(_0244_),
    .A(_0242_),
    .B(_0243_));
 sg13g2_buf_1 _1188_ (.A(_0244_),
    .X(_0245_));
 sg13g2_xnor2_1 _1189_ (.Y(_0246_),
    .A(_0218_),
    .B(_0245_));
 sg13g2_xnor2_1 _1190_ (.Y(_0247_),
    .A(_0192_),
    .B(_0246_));
 sg13g2_xnor2_1 _1191_ (.Y(_0248_),
    .A(_0240_),
    .B(_0247_));
 sg13g2_buf_1 _1192_ (.A(_0076_),
    .X(_0249_));
 sg13g2_xnor2_1 _1193_ (.Y(_0250_),
    .A(_0201_),
    .B(_0137_));
 sg13g2_buf_2 _1194_ (.A(_0250_),
    .X(_0251_));
 sg13g2_nand2b_1 _1195_ (.Y(_0252_),
    .B(_0251_),
    .A_N(_0113_));
 sg13g2_nor2_1 _1196_ (.A(net37),
    .B(_0251_),
    .Y(_0253_));
 sg13g2_o21ai_1 _1197_ (.B1(_0253_),
    .Y(_0254_),
    .A1(net43),
    .A2(_0108_));
 sg13g2_nand2_1 _1198_ (.Y(_0255_),
    .A(_0252_),
    .B(_0254_));
 sg13g2_nand3_1 _1199_ (.B(net39),
    .C(_0255_),
    .A(net29),
    .Y(_0256_));
 sg13g2_buf_1 _1200_ (.A(net38),
    .X(_0257_));
 sg13g2_nand2_1 _1201_ (.Y(_0258_),
    .A(net43),
    .B(_0108_));
 sg13g2_nand2_1 _1202_ (.Y(_0259_),
    .A(net37),
    .B(_0258_));
 sg13g2_nor2_1 _1203_ (.A(net44),
    .B(net43),
    .Y(_0260_));
 sg13g2_and2_1 _1204_ (.A(_0102_),
    .B(_0106_),
    .X(_0261_));
 sg13g2_buf_2 _1205_ (.A(_0261_),
    .X(_0262_));
 sg13g2_buf_1 _1206_ (.A(_0262_),
    .X(_0263_));
 sg13g2_nand3_1 _1207_ (.B(net27),
    .C(_0251_),
    .A(_0260_),
    .Y(_0264_));
 sg13g2_o21ai_1 _1208_ (.B1(_0264_),
    .Y(_0265_),
    .A1(_0251_),
    .A2(_0259_));
 sg13g2_nand3_1 _1209_ (.B(net28),
    .C(_0265_),
    .A(_0249_),
    .Y(_0266_));
 sg13g2_nor2_1 _1210_ (.A(net29),
    .B(_0126_),
    .Y(_0267_));
 sg13g2_nand3_1 _1211_ (.B(_0255_),
    .C(_0267_),
    .A(net28),
    .Y(_0268_));
 sg13g2_a22oi_1 _1212_ (.Y(_0269_),
    .B1(net29),
    .B2(_0112_),
    .A2(_0258_),
    .A1(net37));
 sg13g2_nand2_1 _1213_ (.Y(_0270_),
    .A(net44),
    .B(net43));
 sg13g2_a22oi_1 _1214_ (.Y(_0271_),
    .B1(_0270_),
    .B2(net29),
    .A2(net27),
    .A1(_0260_));
 sg13g2_mux2_1 _1215_ (.A0(_0269_),
    .A1(_0271_),
    .S(_0251_),
    .X(_0272_));
 sg13g2_a21oi_1 _1216_ (.A1(_0263_),
    .A2(net29),
    .Y(_0273_),
    .B1(net28));
 sg13g2_nand2_1 _1217_ (.Y(_0274_),
    .A(net45),
    .B(_0112_));
 sg13g2_nor2_1 _1218_ (.A(_0274_),
    .B(_0251_),
    .Y(_0275_));
 sg13g2_mux2_1 _1219_ (.A0(net45),
    .A1(net43),
    .S(_0107_),
    .X(_0276_));
 sg13g2_xnor2_1 _1220_ (.Y(_0277_),
    .A(_0251_),
    .B(_0276_));
 sg13g2_a21oi_1 _1221_ (.A1(_0274_),
    .A2(_0277_),
    .Y(_0278_),
    .B1(net29));
 sg13g2_mux2_1 _1222_ (.A0(_0091_),
    .A1(_0270_),
    .S(_0251_),
    .X(_0279_));
 sg13g2_nor2_1 _1223_ (.A(_0263_),
    .B(_0279_),
    .Y(_0280_));
 sg13g2_nand2_1 _1224_ (.Y(_0281_),
    .A(net38),
    .B(net31));
 sg13g2_nor4_1 _1225_ (.A(_0275_),
    .B(_0278_),
    .C(_0280_),
    .D(_0281_),
    .Y(_0282_));
 sg13g2_a21oi_1 _1226_ (.A1(_0272_),
    .A2(_0273_),
    .Y(_0283_),
    .B1(_0282_));
 sg13g2_nand4_1 _1227_ (.B(_0266_),
    .C(_0268_),
    .A(_0256_),
    .Y(_0284_),
    .D(_0283_));
 sg13g2_xnor2_1 _1228_ (.Y(_0285_),
    .A(_0248_),
    .B(_0284_));
 sg13g2_inv_1 _1229_ (.Y(_0286_),
    .A(_0206_));
 sg13g2_mux2_1 _1230_ (.A0(_0228_),
    .A1(_0224_),
    .S(_0222_),
    .X(_0287_));
 sg13g2_nand2b_1 _1231_ (.Y(_0288_),
    .B(_0226_),
    .A_N(_0224_));
 sg13g2_mux2_1 _1232_ (.A0(_0287_),
    .A1(_0288_),
    .S(_0180_),
    .X(_0289_));
 sg13g2_nand2_1 _1233_ (.Y(_0290_),
    .A(_0177_),
    .B(_0172_));
 sg13g2_nor2_1 _1234_ (.A(_0175_),
    .B(_0226_),
    .Y(_0291_));
 sg13g2_o21ai_1 _1235_ (.B1(_0291_),
    .Y(_0292_),
    .A1(_0140_),
    .A2(_0290_));
 sg13g2_and2_1 _1236_ (.A(_0177_),
    .B(_0172_),
    .X(_0293_));
 sg13g2_o21ai_1 _1237_ (.B1(_0293_),
    .Y(_0294_),
    .A1(_0215_),
    .A2(_0221_));
 sg13g2_nor2_1 _1238_ (.A(_0293_),
    .B(_0226_),
    .Y(_0295_));
 sg13g2_a22oi_1 _1239_ (.Y(_0296_),
    .B1(_0295_),
    .B2(_0222_),
    .A2(_0294_),
    .A1(_0140_));
 sg13g2_inv_1 _1240_ (.Y(_0297_),
    .A(_0175_));
 sg13g2_nand2_1 _1241_ (.Y(_0298_),
    .A(_0175_),
    .B(_0226_));
 sg13g2_nor2_1 _1242_ (.A(_0177_),
    .B(_0172_),
    .Y(_0299_));
 sg13g2_a221oi_1 _1243_ (.B2(_0140_),
    .C1(_0299_),
    .B1(_0298_),
    .A1(_0297_),
    .Y(_0300_),
    .A2(_0222_));
 sg13g2_a21oi_1 _1244_ (.A1(_0292_),
    .A2(_0296_),
    .Y(_0301_),
    .B1(_0300_));
 sg13g2_o21ai_1 _1245_ (.B1(_0301_),
    .Y(_0302_),
    .A1(_0286_),
    .A2(_0289_));
 sg13g2_nand2_1 _1246_ (.Y(_0303_),
    .A(_0285_),
    .B(_0302_));
 sg13g2_or2_1 _1247_ (.X(_0304_),
    .B(_0302_),
    .A(_0285_));
 sg13g2_and3_1 _1248_ (.X(_0005_),
    .A(net78),
    .B(_0303_),
    .C(_0304_));
 sg13g2_xnor2_1 _1249_ (.Y(_0305_),
    .A(net42),
    .B(_0218_));
 sg13g2_nand2_1 _1250_ (.Y(_0306_),
    .A(net45),
    .B(net34));
 sg13g2_or2_1 _1251_ (.X(_0307_),
    .B(_0306_),
    .A(_0305_));
 sg13g2_xnor2_1 _1252_ (.Y(_0308_),
    .A(_0241_),
    .B(_0243_));
 sg13g2_buf_1 _1253_ (.A(_0308_),
    .X(_0309_));
 sg13g2_a21oi_1 _1254_ (.A1(_0156_),
    .A2(_0168_),
    .Y(_0310_),
    .B1(net40));
 sg13g2_and3_1 _1255_ (.X(_0311_),
    .A(_0156_),
    .B(_0168_),
    .C(net40));
 sg13g2_or2_1 _1256_ (.X(_0312_),
    .B(_0311_),
    .A(_0310_));
 sg13g2_buf_1 _1257_ (.A(_0312_),
    .X(_0313_));
 sg13g2_nand3_1 _1258_ (.B(_0313_),
    .C(_0305_),
    .A(net34),
    .Y(_0314_));
 sg13g2_nor2_1 _1259_ (.A(net36),
    .B(_0237_),
    .Y(_0315_));
 sg13g2_a22oi_1 _1260_ (.Y(_0316_),
    .B1(_0305_),
    .B2(_0239_),
    .A2(_0313_),
    .A1(_0315_));
 sg13g2_nor2_1 _1261_ (.A(_0235_),
    .B(_0313_),
    .Y(_0317_));
 sg13g2_a21oi_1 _1262_ (.A1(_0235_),
    .A2(_0313_),
    .Y(_0318_),
    .B1(net34));
 sg13g2_o21ai_1 _1263_ (.B1(_0318_),
    .Y(_0319_),
    .A1(_0305_),
    .A2(_0317_));
 sg13g2_nand4_1 _1264_ (.B(_0314_),
    .C(_0316_),
    .A(_0307_),
    .Y(_0320_),
    .D(_0319_));
 sg13g2_nand2_1 _1265_ (.Y(_0321_),
    .A(_0193_),
    .B(_0141_));
 sg13g2_xnor2_1 _1266_ (.Y(_0322_),
    .A(_0176_),
    .B(_0321_));
 sg13g2_xnor2_1 _1267_ (.Y(_0323_),
    .A(_0145_),
    .B(_0262_));
 sg13g2_mux2_1 _1268_ (.A0(_0310_),
    .A1(_0311_),
    .S(net34),
    .X(_0324_));
 sg13g2_xnor2_1 _1269_ (.Y(_0325_),
    .A(_0323_),
    .B(_0324_));
 sg13g2_xnor2_1 _1270_ (.Y(_0326_),
    .A(_0322_),
    .B(_0325_));
 sg13g2_nand2_1 _1271_ (.Y(_0327_),
    .A(net35),
    .B(_0187_));
 sg13g2_nor2_1 _1272_ (.A(_0193_),
    .B(net42),
    .Y(_0328_));
 sg13g2_a221oi_1 _1273_ (.B2(_0327_),
    .C1(_0328_),
    .B1(_0306_),
    .A1(_0184_),
    .Y(_0329_),
    .A2(_0218_));
 sg13g2_xnor2_1 _1274_ (.Y(_0330_),
    .A(_0126_),
    .B(_0329_));
 sg13g2_xnor2_1 _1275_ (.Y(_0331_),
    .A(_0326_),
    .B(_0330_));
 sg13g2_xnor2_1 _1276_ (.Y(_0332_),
    .A(_0320_),
    .B(_0331_));
 sg13g2_nand2_1 _1277_ (.Y(_0333_),
    .A(net29),
    .B(_0126_));
 sg13g2_nor2b_1 _1278_ (.A(_0277_),
    .B_N(_0333_),
    .Y(_0334_));
 sg13g2_a21oi_1 _1279_ (.A1(net29),
    .A2(net31),
    .Y(_0335_),
    .B1(_0274_));
 sg13g2_nor3_1 _1280_ (.A(net39),
    .B(_0267_),
    .C(_0335_),
    .Y(_0336_));
 sg13g2_o21ai_1 _1281_ (.B1(_0336_),
    .Y(_0337_),
    .A1(_0280_),
    .A2(_0334_));
 sg13g2_or4_1 _1282_ (.A(_0123_),
    .B(_0274_),
    .C(_0277_),
    .D(_0333_),
    .X(_0338_));
 sg13g2_nand3_1 _1283_ (.B(_0337_),
    .C(_0338_),
    .A(_0248_),
    .Y(_0339_));
 sg13g2_or4_1 _1284_ (.A(net28),
    .B(_0275_),
    .C(_0278_),
    .D(_0280_),
    .X(_0340_));
 sg13g2_nor2_1 _1285_ (.A(_0267_),
    .B(_0335_),
    .Y(_0341_));
 sg13g2_nor2_1 _1286_ (.A(_0123_),
    .B(_0341_),
    .Y(_0342_));
 sg13g2_a21oi_1 _1287_ (.A1(_0339_),
    .A2(_0340_),
    .Y(_0343_),
    .B1(_0342_));
 sg13g2_nor2b_1 _1288_ (.A(_0268_),
    .B_N(_0339_),
    .Y(_0344_));
 sg13g2_nor2_1 _1289_ (.A(_0343_),
    .B(_0344_),
    .Y(_0345_));
 sg13g2_xor2_1 _1290_ (.B(_0345_),
    .A(_0332_),
    .X(_0346_));
 sg13g2_xnor2_1 _1291_ (.Y(_0347_),
    .A(_0303_),
    .B(_0346_));
 sg13g2_nor2_1 _1292_ (.A(net77),
    .B(_0347_),
    .Y(_0006_));
 sg13g2_nand3b_1 _1293_ (.B(_0339_),
    .C(_0340_),
    .Y(_0348_),
    .A_N(_0332_));
 sg13g2_nand2b_1 _1294_ (.Y(_0349_),
    .B(_0342_),
    .A_N(_0332_));
 sg13g2_nand3b_1 _1295_ (.B(_0348_),
    .C(_0349_),
    .Y(_0350_),
    .A_N(_0344_));
 sg13g2_a21o_1 _1296_ (.A2(_0302_),
    .A1(_0285_),
    .B1(_0350_),
    .X(_0351_));
 sg13g2_nand2_1 _1297_ (.Y(_0352_),
    .A(net34),
    .B(net40));
 sg13g2_a21oi_1 _1298_ (.A1(_0322_),
    .A2(_0352_),
    .Y(_0353_),
    .B1(_0323_));
 sg13g2_nor2_1 _1299_ (.A(_0322_),
    .B(_0352_),
    .Y(_0354_));
 sg13g2_buf_1 _1300_ (.A(_0210_),
    .X(_0355_));
 sg13g2_o21ai_1 _1301_ (.B1(_0355_),
    .Y(_0356_),
    .A1(_0353_),
    .A2(_0354_));
 sg13g2_nand2_1 _1302_ (.Y(_0357_),
    .A(net46),
    .B(_0245_));
 sg13g2_mux2_1 _1303_ (.A0(net36),
    .A1(_0357_),
    .S(_0322_),
    .X(_0358_));
 sg13g2_buf_1 _1304_ (.A(net73),
    .X(_0359_));
 sg13g2_xnor2_1 _1305_ (.Y(_0360_),
    .A(net60),
    .B(_0262_));
 sg13g2_nor2_1 _1306_ (.A(_0355_),
    .B(_0360_),
    .Y(_0361_));
 sg13g2_nor3_1 _1307_ (.A(net34),
    .B(net41),
    .C(_0322_),
    .Y(_0362_));
 sg13g2_a22oi_1 _1308_ (.Y(_0363_),
    .B1(_0362_),
    .B2(_0360_),
    .A2(_0361_),
    .A1(_0358_));
 sg13g2_and2_1 _1309_ (.A(_0356_),
    .B(_0363_),
    .X(_0364_));
 sg13g2_nand3_1 _1310_ (.B(_0262_),
    .C(net30),
    .A(_0094_),
    .Y(_0365_));
 sg13g2_nand3_1 _1311_ (.B(_0107_),
    .C(_0210_),
    .A(_0145_),
    .Y(_0366_));
 sg13g2_nand2_1 _1312_ (.Y(_0367_),
    .A(net49),
    .B(_0792_));
 sg13g2_o21ai_1 _1313_ (.B1(_0367_),
    .Y(_0368_),
    .A1(_0856_),
    .A2(_0080_));
 sg13g2_inv_1 _1314_ (.Y(_0369_),
    .A(_0792_));
 sg13g2_a21o_1 _1315_ (.A2(_0035_),
    .A1(_0856_),
    .B1(_0369_),
    .X(_0370_));
 sg13g2_nand2_1 _1316_ (.Y(_0371_),
    .A(_0035_),
    .B(_0131_));
 sg13g2_a21oi_1 _1317_ (.A1(_0370_),
    .A2(_0371_),
    .Y(_0372_),
    .B1(_0738_));
 sg13g2_a21oi_1 _1318_ (.A1(_0738_),
    .A2(_0368_),
    .Y(_0373_),
    .B1(_0372_));
 sg13g2_xnor2_1 _1319_ (.Y(_0374_),
    .A(_0039_),
    .B(_0373_));
 sg13g2_and3_1 _1320_ (.X(_0375_),
    .A(_0365_),
    .B(_0366_),
    .C(_0374_));
 sg13g2_a21oi_1 _1321_ (.A1(_0365_),
    .A2(_0366_),
    .Y(_0376_),
    .B1(_0374_));
 sg13g2_o21ai_1 _1322_ (.B1(_0046_),
    .Y(_0377_),
    .A1(net44),
    .A2(_0085_));
 sg13g2_nand3b_1 _1323_ (.B(_0201_),
    .C(net45),
    .Y(_0378_),
    .A_N(_0085_));
 sg13g2_buf_1 _1324_ (.A(_0378_),
    .X(_0379_));
 sg13g2_and2_1 _1325_ (.A(_0377_),
    .B(_0379_),
    .X(_0380_));
 sg13g2_o21ai_1 _1326_ (.B1(_0380_),
    .Y(_0381_),
    .A1(_0375_),
    .A2(_0376_));
 sg13g2_or3_1 _1327_ (.A(_0380_),
    .B(_0375_),
    .C(_0376_),
    .X(_0382_));
 sg13g2_nand2_2 _1328_ (.Y(_0383_),
    .A(_0381_),
    .B(_0382_));
 sg13g2_nand2_1 _1329_ (.Y(_0384_),
    .A(_0176_),
    .B(_0321_));
 sg13g2_nor2_1 _1330_ (.A(net46),
    .B(net26),
    .Y(_0385_));
 sg13g2_nor2_1 _1331_ (.A(_0176_),
    .B(_0321_),
    .Y(_0386_));
 sg13g2_a21oi_2 _1332_ (.B1(_0386_),
    .Y(_0387_),
    .A2(_0385_),
    .A1(_0384_));
 sg13g2_xnor2_1 _1333_ (.Y(_0388_),
    .A(_0075_),
    .B(_0387_));
 sg13g2_xnor2_1 _1334_ (.Y(_0389_),
    .A(_0383_),
    .B(_0388_));
 sg13g2_xnor2_1 _1335_ (.Y(_0390_),
    .A(_0364_),
    .B(_0389_));
 sg13g2_nor2_1 _1336_ (.A(_0326_),
    .B(_0330_),
    .Y(_0391_));
 sg13g2_nand2_1 _1337_ (.Y(_0392_),
    .A(_0326_),
    .B(_0330_));
 sg13g2_o21ai_1 _1338_ (.B1(_0392_),
    .Y(_0393_),
    .A1(_0320_),
    .A2(_0391_));
 sg13g2_a21oi_1 _1339_ (.A1(_0184_),
    .A2(_0306_),
    .Y(_0394_),
    .B1(_0328_));
 sg13g2_and2_1 _1340_ (.A(net35),
    .B(_0394_),
    .X(_0395_));
 sg13g2_xor2_1 _1341_ (.B(_0395_),
    .A(_0393_),
    .X(_0396_));
 sg13g2_xnor2_1 _1342_ (.Y(_0397_),
    .A(_0390_),
    .B(_0396_));
 sg13g2_and2_1 _1343_ (.A(_0332_),
    .B(_0343_),
    .X(_0398_));
 sg13g2_nor2_1 _1344_ (.A(_0397_),
    .B(_0398_),
    .Y(_0399_));
 sg13g2_nand2_1 _1345_ (.Y(_0400_),
    .A(_0351_),
    .B(_0399_));
 sg13g2_nand2b_1 _1346_ (.Y(_0401_),
    .B(_0351_),
    .A_N(_0398_));
 sg13g2_nand2_1 _1347_ (.Y(_0402_),
    .A(_0397_),
    .B(_0401_));
 sg13g2_and3_1 _1348_ (.X(_0007_),
    .A(net78),
    .B(_0400_),
    .C(_0402_));
 sg13g2_nand2_1 _1349_ (.Y(_0403_),
    .A(_0390_),
    .B(_0395_));
 sg13g2_o21ai_1 _1350_ (.B1(_0393_),
    .Y(_0404_),
    .A1(_0390_),
    .A2(_0395_));
 sg13g2_nand4_1 _1351_ (.B(_0363_),
    .C(_0383_),
    .A(_0356_),
    .Y(_0405_),
    .D(_0387_));
 sg13g2_a21o_1 _1352_ (.A2(_0385_),
    .A1(_0384_),
    .B1(_0386_),
    .X(_0406_));
 sg13g2_nand4_1 _1353_ (.B(_0381_),
    .C(_0382_),
    .A(_0075_),
    .Y(_0407_),
    .D(_0406_));
 sg13g2_a21o_1 _1354_ (.A2(_0363_),
    .A1(_0356_),
    .B1(_0407_),
    .X(_0408_));
 sg13g2_nand3_1 _1355_ (.B(_0382_),
    .C(_0406_),
    .A(_0381_),
    .Y(_0409_));
 sg13g2_nand4_1 _1356_ (.B(_0356_),
    .C(_0363_),
    .A(_0196_),
    .Y(_0410_),
    .D(_0409_));
 sg13g2_nand3_1 _1357_ (.B(_0383_),
    .C(_0387_),
    .A(_0196_),
    .Y(_0411_));
 sg13g2_nand4_1 _1358_ (.B(_0408_),
    .C(_0410_),
    .A(_0405_),
    .Y(_0412_),
    .D(_0411_));
 sg13g2_a21oi_1 _1359_ (.A1(_0377_),
    .A2(_0379_),
    .Y(_0413_),
    .B1(_0374_));
 sg13g2_nand2_1 _1360_ (.Y(_0414_),
    .A(net60),
    .B(net30));
 sg13g2_nand3_1 _1361_ (.B(_0379_),
    .C(_0374_),
    .A(_0377_),
    .Y(_0415_));
 sg13g2_o21ai_1 _1362_ (.B1(_0415_),
    .Y(_0416_),
    .A1(_0413_),
    .A2(_0414_));
 sg13g2_xnor2_1 _1363_ (.Y(_0417_),
    .A(_0128_),
    .B(_0373_));
 sg13g2_nand2_1 _1364_ (.Y(_0418_),
    .A(_0145_),
    .B(net26));
 sg13g2_a22oi_1 _1365_ (.Y(_0419_),
    .B1(_0417_),
    .B2(_0418_),
    .A2(_0379_),
    .A1(_0377_));
 sg13g2_and3_1 _1366_ (.X(_0420_),
    .A(net30),
    .B(_0377_),
    .C(_0379_));
 sg13g2_o21ai_1 _1367_ (.B1(net32),
    .Y(_0421_),
    .A1(net60),
    .A2(_0417_));
 sg13g2_nor3_1 _1368_ (.A(_0419_),
    .B(_0420_),
    .C(_0421_),
    .Y(_0422_));
 sg13g2_a21o_1 _1369_ (.A2(_0416_),
    .A1(net27),
    .B1(_0422_),
    .X(_0423_));
 sg13g2_buf_1 _1370_ (.A(net75),
    .X(_0424_));
 sg13g2_xnor2_1 _1371_ (.Y(_0425_),
    .A(net59),
    .B(net41));
 sg13g2_xnor2_1 _1372_ (.Y(_0426_),
    .A(_0210_),
    .B(_0238_));
 sg13g2_a22oi_1 _1373_ (.Y(_0427_),
    .B1(_0134_),
    .B2(_0136_),
    .A2(_0106_),
    .A1(_0102_));
 sg13g2_and4_1 _1374_ (.A(_0102_),
    .B(_0106_),
    .C(_0134_),
    .D(_0136_),
    .X(_0428_));
 sg13g2_mux2_1 _1375_ (.A0(_0427_),
    .A1(_0428_),
    .S(_0369_),
    .X(_0429_));
 sg13g2_xnor2_1 _1376_ (.Y(_0430_),
    .A(_0426_),
    .B(_0429_));
 sg13g2_xnor2_1 _1377_ (.Y(_0431_),
    .A(_0425_),
    .B(_0430_));
 sg13g2_xnor2_1 _1378_ (.Y(_0432_),
    .A(net38),
    .B(net42));
 sg13g2_nor3_1 _1379_ (.A(net44),
    .B(net43),
    .C(net46),
    .Y(_0433_));
 sg13g2_a22oi_1 _1380_ (.Y(_0434_),
    .B1(net30),
    .B2(net32),
    .A2(net46),
    .A1(net43));
 sg13g2_nor2_1 _1381_ (.A(net45),
    .B(net34),
    .Y(_0435_));
 sg13g2_nor3_1 _1382_ (.A(_0433_),
    .B(_0434_),
    .C(_0435_),
    .Y(_0436_));
 sg13g2_xor2_1 _1383_ (.B(_0436_),
    .A(_0432_),
    .X(_0437_));
 sg13g2_xor2_1 _1384_ (.B(_0437_),
    .A(_0431_),
    .X(_0438_));
 sg13g2_xnor2_1 _1385_ (.Y(_0439_),
    .A(_0423_),
    .B(_0438_));
 sg13g2_xnor2_1 _1386_ (.Y(_0440_),
    .A(_0412_),
    .B(_0439_));
 sg13g2_nand3_1 _1387_ (.B(_0404_),
    .C(_0440_),
    .A(_0403_),
    .Y(_0441_));
 sg13g2_nand2_1 _1388_ (.Y(_0442_),
    .A(_0403_),
    .B(_0404_));
 sg13g2_inv_1 _1389_ (.Y(_0443_),
    .A(_0440_));
 sg13g2_nand2_1 _1390_ (.Y(_0444_),
    .A(_0442_),
    .B(_0443_));
 sg13g2_nand2_1 _1391_ (.Y(_0445_),
    .A(_0441_),
    .B(_0444_));
 sg13g2_xnor2_1 _1392_ (.Y(_0446_),
    .A(_0400_),
    .B(_0445_));
 sg13g2_nor2_1 _1393_ (.A(_0717_),
    .B(_0446_),
    .Y(_0008_));
 sg13g2_inv_1 _1394_ (.Y(_0447_),
    .A(_0441_));
 sg13g2_a21oi_1 _1395_ (.A1(_0400_),
    .A2(_0444_),
    .Y(_0448_),
    .B1(_0447_));
 sg13g2_a21oi_1 _1396_ (.A1(_0409_),
    .A2(_0439_),
    .Y(_0449_),
    .B1(_0364_));
 sg13g2_and2_1 _1397_ (.A(_0364_),
    .B(_0409_),
    .X(_0450_));
 sg13g2_a221oi_1 _1398_ (.B2(_0196_),
    .C1(_0439_),
    .B1(_0450_),
    .A1(_0383_),
    .Y(_0451_),
    .A2(_0387_));
 sg13g2_a21o_1 _1399_ (.A2(_0449_),
    .A1(_0075_),
    .B1(_0451_),
    .X(_0452_));
 sg13g2_xnor2_1 _1400_ (.Y(_0453_),
    .A(net30),
    .B(_0238_));
 sg13g2_nor2_1 _1401_ (.A(_0369_),
    .B(net27),
    .Y(_0454_));
 sg13g2_o21ai_1 _1402_ (.B1(_0454_),
    .Y(_0455_),
    .A1(_0425_),
    .A2(_0453_));
 sg13g2_nand2_1 _1403_ (.Y(_0456_),
    .A(_0425_),
    .B(_0453_));
 sg13g2_and2_1 _1404_ (.A(_0455_),
    .B(_0456_),
    .X(_0457_));
 sg13g2_buf_1 _1405_ (.A(net76),
    .X(_0458_));
 sg13g2_nor2_1 _1406_ (.A(net58),
    .B(net32),
    .Y(_0459_));
 sg13g2_o21ai_1 _1407_ (.B1(_0426_),
    .Y(_0460_),
    .A1(_0425_),
    .A2(_0459_));
 sg13g2_a22oi_1 _1408_ (.Y(_0461_),
    .B1(_0453_),
    .B2(net32),
    .A2(_0425_),
    .A1(_0369_));
 sg13g2_a21oi_1 _1409_ (.A1(_0460_),
    .A2(_0461_),
    .Y(_0462_),
    .B1(net33));
 sg13g2_a21oi_1 _1410_ (.A1(net33),
    .A2(_0457_),
    .Y(_0463_),
    .B1(_0462_));
 sg13g2_nand2_1 _1411_ (.Y(_0464_),
    .A(net36),
    .B(net26));
 sg13g2_o21ai_1 _1412_ (.B1(net30),
    .Y(_0465_),
    .A1(_0262_),
    .A2(net33));
 sg13g2_a21oi_1 _1413_ (.A1(_0464_),
    .A2(_0465_),
    .Y(_0466_),
    .B1(net37));
 sg13g2_xnor2_1 _1414_ (.Y(_0467_),
    .A(net46),
    .B(net26));
 sg13g2_nor4_1 _1415_ (.A(net45),
    .B(net27),
    .C(net33),
    .D(_0467_),
    .Y(_0468_));
 sg13g2_nor2_1 _1416_ (.A(net39),
    .B(net42),
    .Y(_0469_));
 sg13g2_xnor2_1 _1417_ (.Y(_0470_),
    .A(net31),
    .B(_0469_));
 sg13g2_o21ai_1 _1418_ (.B1(_0470_),
    .Y(_0471_),
    .A1(_0466_),
    .A2(_0468_));
 sg13g2_or3_1 _1419_ (.A(_0466_),
    .B(_0468_),
    .C(_0470_),
    .X(_0472_));
 sg13g2_a22oi_1 _1420_ (.Y(_0473_),
    .B1(_0156_),
    .B2(_0168_),
    .A2(_0045_),
    .A1(_0038_));
 sg13g2_xnor2_1 _1421_ (.Y(_0474_),
    .A(_0262_),
    .B(_0473_));
 sg13g2_xnor2_1 _1422_ (.Y(_0475_),
    .A(net48),
    .B(net73));
 sg13g2_and2_1 _1423_ (.A(net75),
    .B(net41),
    .X(_0476_));
 sg13g2_nor2_1 _1424_ (.A(net59),
    .B(net41),
    .Y(_0477_));
 sg13g2_mux2_1 _1425_ (.A0(_0476_),
    .A1(_0477_),
    .S(net33),
    .X(_0478_));
 sg13g2_xnor2_1 _1426_ (.Y(_0479_),
    .A(_0475_),
    .B(_0478_));
 sg13g2_xnor2_1 _1427_ (.Y(_0480_),
    .A(_0474_),
    .B(_0479_));
 sg13g2_a21o_1 _1428_ (.A2(_0472_),
    .A1(_0471_),
    .B1(_0480_),
    .X(_0481_));
 sg13g2_nand3_1 _1429_ (.B(_0471_),
    .C(_0472_),
    .A(_0480_),
    .Y(_0482_));
 sg13g2_and3_1 _1430_ (.X(_0483_),
    .A(_0463_),
    .B(_0481_),
    .C(_0482_));
 sg13g2_a21oi_1 _1431_ (.A1(_0481_),
    .A2(_0482_),
    .Y(_0484_),
    .B1(_0463_));
 sg13g2_nor2_1 _1432_ (.A(_0483_),
    .B(_0484_),
    .Y(_0485_));
 sg13g2_nand2b_1 _1433_ (.Y(_0486_),
    .B(_0436_),
    .A_N(_0432_));
 sg13g2_nand2_1 _1434_ (.Y(_0487_),
    .A(_0431_),
    .B(_0437_));
 sg13g2_nor2_1 _1435_ (.A(_0431_),
    .B(_0437_),
    .Y(_0488_));
 sg13g2_a21o_1 _1436_ (.A2(_0487_),
    .A1(_0423_),
    .B1(_0488_),
    .X(_0489_));
 sg13g2_xnor2_1 _1437_ (.Y(_0490_),
    .A(_0486_),
    .B(_0489_));
 sg13g2_xnor2_1 _1438_ (.Y(_0491_),
    .A(_0485_),
    .B(_0490_));
 sg13g2_xor2_1 _1439_ (.B(_0491_),
    .A(_0452_),
    .X(_0492_));
 sg13g2_xnor2_1 _1440_ (.Y(_0493_),
    .A(_0448_),
    .B(_0492_));
 sg13g2_nor2_1 _1441_ (.A(_0717_),
    .B(_0493_),
    .Y(_0009_));
 sg13g2_o21ai_1 _1442_ (.B1(_0489_),
    .Y(_0494_),
    .A1(_0483_),
    .A2(_0484_));
 sg13g2_nor3_1 _1443_ (.A(_0489_),
    .B(_0483_),
    .C(_0484_),
    .Y(_0495_));
 sg13g2_a21oi_2 _1444_ (.B1(_0495_),
    .Y(_0496_),
    .A2(_0494_),
    .A1(_0486_));
 sg13g2_nand2_1 _1445_ (.Y(_0497_),
    .A(_0471_),
    .B(_0472_));
 sg13g2_nor2_1 _1446_ (.A(_0480_),
    .B(_0497_),
    .Y(_0498_));
 sg13g2_nand2_1 _1447_ (.Y(_0499_),
    .A(_0480_),
    .B(_0497_));
 sg13g2_o21ai_1 _1448_ (.B1(_0499_),
    .Y(_0500_),
    .A1(_0463_),
    .A2(_0498_));
 sg13g2_a22oi_1 _1449_ (.Y(_0501_),
    .B1(net26),
    .B2(net45),
    .A2(_0237_),
    .A1(net32));
 sg13g2_mux2_1 _1450_ (.A0(net34),
    .A1(_0238_),
    .S(net30),
    .X(_0502_));
 sg13g2_nand2b_1 _1451_ (.Y(_0503_),
    .B(_0502_),
    .A_N(_0501_));
 sg13g2_buf_1 _1452_ (.A(_0503_),
    .X(_0504_));
 sg13g2_a21o_1 _1453_ (.A2(net31),
    .A1(net37),
    .B1(_0504_),
    .X(_0505_));
 sg13g2_o21ai_1 _1454_ (.B1(net28),
    .Y(_0506_),
    .A1(_0185_),
    .A2(_0504_));
 sg13g2_o21ai_1 _1455_ (.B1(_0506_),
    .Y(_0507_),
    .A1(net28),
    .A2(_0505_));
 sg13g2_nor2_1 _1456_ (.A(_0181_),
    .B(net39),
    .Y(_0508_));
 sg13g2_mux2_1 _1457_ (.A0(_0508_),
    .A1(_0182_),
    .S(_0504_),
    .X(_0509_));
 sg13g2_nor2_1 _1458_ (.A(_0257_),
    .B(_0182_),
    .Y(_0510_));
 sg13g2_a21o_1 _1459_ (.A2(_0504_),
    .A1(net42),
    .B1(_0510_),
    .X(_0511_));
 sg13g2_a22oi_1 _1460_ (.Y(_0512_),
    .B1(_0511_),
    .B2(_0090_),
    .A2(_0509_),
    .A1(_0187_));
 sg13g2_and2_1 _1461_ (.A(_0507_),
    .B(_0512_),
    .X(_0513_));
 sg13g2_nor2_1 _1462_ (.A(_0234_),
    .B(net40),
    .Y(_0514_));
 sg13g2_a21oi_1 _1463_ (.A1(_0234_),
    .A2(_0474_),
    .Y(_0515_),
    .B1(_0514_));
 sg13g2_nand2_1 _1464_ (.Y(_0516_),
    .A(_0474_),
    .B(_0514_));
 sg13g2_o21ai_1 _1465_ (.B1(_0516_),
    .Y(_0517_),
    .A1(_0475_),
    .A2(_0515_));
 sg13g2_nor2_1 _1466_ (.A(_0424_),
    .B(_0237_),
    .Y(_0518_));
 sg13g2_mux2_1 _1467_ (.A0(_0518_),
    .A1(_0237_),
    .S(_0474_),
    .X(_0519_));
 sg13g2_nand2_1 _1468_ (.Y(_0520_),
    .A(_0309_),
    .B(_0475_));
 sg13g2_nand3b_1 _1469_ (.B(_0474_),
    .C(net41),
    .Y(_0521_),
    .A_N(_0475_));
 sg13g2_o21ai_1 _1470_ (.B1(_0521_),
    .Y(_0522_),
    .A1(_0519_),
    .A2(_0520_));
 sg13g2_a21o_1 _1471_ (.A2(_0517_),
    .A1(_0424_),
    .B1(_0522_),
    .X(_0523_));
 sg13g2_nor2_1 _1472_ (.A(net27),
    .B(net26),
    .Y(_0524_));
 sg13g2_a22oi_1 _1473_ (.Y(_0525_),
    .B1(_0237_),
    .B2(net40),
    .A2(_0207_),
    .A1(net27));
 sg13g2_a221oi_1 _1474_ (.B2(net36),
    .C1(_0525_),
    .B1(_0524_),
    .A1(net27),
    .Y(_0526_),
    .A2(net26));
 sg13g2_buf_1 _1475_ (.A(_0526_),
    .X(_0527_));
 sg13g2_nor2_1 _1476_ (.A(_0111_),
    .B(_0126_),
    .Y(_0528_));
 sg13g2_a21oi_1 _1477_ (.A1(_0181_),
    .A2(net38),
    .Y(_0529_),
    .B1(_0528_));
 sg13g2_xnor2_1 _1478_ (.Y(_0530_),
    .A(_0078_),
    .B(_0529_));
 sg13g2_xnor2_1 _1479_ (.Y(_0531_),
    .A(_0527_),
    .B(_0530_));
 sg13g2_nor2_1 _1480_ (.A(_0262_),
    .B(net30),
    .Y(_0532_));
 sg13g2_xnor2_1 _1481_ (.Y(_0533_),
    .A(_0237_),
    .B(_0532_));
 sg13g2_nor2b_1 _1482_ (.A(_0458_),
    .B_N(net49),
    .Y(_0534_));
 sg13g2_or2_1 _1483_ (.X(_0535_),
    .B(_0534_),
    .A(_0087_));
 sg13g2_buf_1 _1484_ (.A(_0535_),
    .X(_0536_));
 sg13g2_nor2_1 _1485_ (.A(net60),
    .B(net41),
    .Y(_0537_));
 sg13g2_nor3_1 _1486_ (.A(net48),
    .B(_0145_),
    .C(net40),
    .Y(_0538_));
 sg13g2_a21oi_1 _1487_ (.A1(net48),
    .A2(_0537_),
    .Y(_0539_),
    .B1(_0538_));
 sg13g2_xnor2_1 _1488_ (.Y(_0540_),
    .A(_0536_),
    .B(_0539_));
 sg13g2_xnor2_1 _1489_ (.Y(_0541_),
    .A(_0533_),
    .B(_0540_));
 sg13g2_xnor2_1 _1490_ (.Y(_0542_),
    .A(_0531_),
    .B(_0541_));
 sg13g2_xnor2_1 _1491_ (.Y(_0543_),
    .A(_0523_),
    .B(_0542_));
 sg13g2_xnor2_1 _1492_ (.Y(_0544_),
    .A(_0513_),
    .B(_0543_));
 sg13g2_xnor2_1 _1493_ (.Y(_0545_),
    .A(_0500_),
    .B(_0544_));
 sg13g2_xor2_1 _1494_ (.B(_0545_),
    .A(_0496_),
    .X(_0546_));
 sg13g2_a21oi_1 _1495_ (.A1(_0441_),
    .A2(_0452_),
    .Y(_0547_),
    .B1(_0491_));
 sg13g2_a221oi_1 _1496_ (.B2(_0443_),
    .C1(_0491_),
    .B1(_0442_),
    .A1(_0351_),
    .Y(_0548_),
    .A2(_0399_));
 sg13g2_nor2_1 _1497_ (.A(_0441_),
    .B(_0452_),
    .Y(_0549_));
 sg13g2_a221oi_1 _1498_ (.B2(_0443_),
    .C1(_0452_),
    .B1(_0442_),
    .A1(_0351_),
    .Y(_0550_),
    .A2(_0399_));
 sg13g2_or4_1 _1499_ (.A(_0547_),
    .B(_0548_),
    .C(_0549_),
    .D(_0550_),
    .X(_0551_));
 sg13g2_or2_1 _1500_ (.X(_0552_),
    .B(_0551_),
    .A(_0546_));
 sg13g2_nand2_1 _1501_ (.Y(_0553_),
    .A(_0546_),
    .B(_0551_));
 sg13g2_and3_1 _1502_ (.X(_0010_),
    .A(_0233_),
    .B(_0552_),
    .C(_0553_));
 sg13g2_inv_1 _1503_ (.Y(_0554_),
    .A(_0513_));
 sg13g2_xor2_1 _1504_ (.B(_0542_),
    .A(_0523_),
    .X(_0555_));
 sg13g2_nand2_1 _1505_ (.Y(_0556_),
    .A(_0554_),
    .B(_0555_));
 sg13g2_o21ai_1 _1506_ (.B1(_0500_),
    .Y(_0557_),
    .A1(_0554_),
    .A2(_0555_));
 sg13g2_a21o_1 _1507_ (.A2(_0557_),
    .A1(_0556_),
    .B1(_0496_),
    .X(_0558_));
 sg13g2_nor2_1 _1508_ (.A(_0513_),
    .B(_0543_),
    .Y(_0559_));
 sg13g2_nor3_1 _1509_ (.A(_0500_),
    .B(_0554_),
    .C(_0555_),
    .Y(_0560_));
 sg13g2_a22oi_1 _1510_ (.Y(_0561_),
    .B1(_0560_),
    .B2(_0496_),
    .A2(_0559_),
    .A1(_0500_));
 sg13g2_or2_1 _1511_ (.X(_0562_),
    .B(_0533_),
    .A(net60));
 sg13g2_nor2_1 _1512_ (.A(net40),
    .B(_0533_),
    .Y(_0563_));
 sg13g2_o21ai_1 _1513_ (.B1(_0536_),
    .Y(_0564_),
    .A1(_0537_),
    .A2(_0563_));
 sg13g2_o21ai_1 _1514_ (.B1(_0564_),
    .Y(_0565_),
    .A1(net41),
    .A2(_0562_));
 sg13g2_nand2_1 _1515_ (.Y(_0566_),
    .A(_0536_),
    .B(_0562_));
 sg13g2_o21ai_1 _1516_ (.B1(_0533_),
    .Y(_0567_),
    .A1(_0129_),
    .A2(net40));
 sg13g2_nand2b_1 _1517_ (.Y(_0568_),
    .B(_0567_),
    .A_N(_0563_));
 sg13g2_a21o_1 _1518_ (.A2(_0568_),
    .A1(_0359_),
    .B1(_0536_),
    .X(_0569_));
 sg13g2_a22oi_1 _1519_ (.Y(_0570_),
    .B1(_0566_),
    .B2(_0569_),
    .A2(_0565_),
    .A1(_0129_));
 sg13g2_nor3_1 _1520_ (.A(net35),
    .B(_0075_),
    .C(net39),
    .Y(_0571_));
 sg13g2_nor2_1 _1521_ (.A(net36),
    .B(net28),
    .Y(_0572_));
 sg13g2_a22oi_1 _1522_ (.Y(_0573_),
    .B1(_0572_),
    .B2(_0075_),
    .A2(_0571_),
    .A1(net36));
 sg13g2_o21ai_1 _1523_ (.B1(_0194_),
    .Y(_0574_),
    .A1(net35),
    .A2(_0217_));
 sg13g2_nand3b_1 _1524_ (.B(_0196_),
    .C(_0217_),
    .Y(_0575_),
    .A_N(net35));
 sg13g2_a21oi_1 _1525_ (.A1(_0574_),
    .A2(_0575_),
    .Y(_0576_),
    .B1(net28));
 sg13g2_nand2_1 _1526_ (.Y(_0577_),
    .A(_0174_),
    .B(_0217_));
 sg13g2_nand2_1 _1527_ (.Y(_0578_),
    .A(net35),
    .B(_0075_));
 sg13g2_a21oi_1 _1528_ (.A1(_0577_),
    .A2(_0578_),
    .Y(_0579_),
    .B1(_0194_));
 sg13g2_nor2_1 _1529_ (.A(_0249_),
    .B(_0577_),
    .Y(_0580_));
 sg13g2_nor3_1 _1530_ (.A(_0576_),
    .B(_0579_),
    .C(_0580_),
    .Y(_0581_));
 sg13g2_o21ai_1 _1531_ (.B1(_0581_),
    .Y(_0582_),
    .A1(_0217_),
    .A2(_0573_));
 sg13g2_a22oi_1 _1532_ (.Y(_0583_),
    .B1(_0534_),
    .B2(_0359_),
    .A2(_0095_),
    .A1(_0458_));
 sg13g2_xnor2_1 _1533_ (.Y(_0584_),
    .A(net64),
    .B(_0583_));
 sg13g2_xnor2_1 _1534_ (.Y(_0585_),
    .A(net31),
    .B(_0584_));
 sg13g2_xnor2_1 _1535_ (.Y(_0586_),
    .A(net42),
    .B(_0425_));
 sg13g2_xnor2_1 _1536_ (.Y(_0587_),
    .A(_0585_),
    .B(_0586_));
 sg13g2_nor2_1 _1537_ (.A(net32),
    .B(net26),
    .Y(_0588_));
 sg13g2_nor2_1 _1538_ (.A(_0145_),
    .B(net41),
    .Y(_0589_));
 sg13g2_a21o_1 _1539_ (.A2(_0589_),
    .A1(_0532_),
    .B1(_0588_),
    .X(_0590_));
 sg13g2_nor4_1 _1540_ (.A(net33),
    .B(_0588_),
    .C(_0532_),
    .D(_0589_),
    .Y(_0591_));
 sg13g2_a221oi_1 _1541_ (.B2(net33),
    .C1(_0591_),
    .B1(_0590_),
    .A1(_0588_),
    .Y(_0592_),
    .A2(_0589_));
 sg13g2_xnor2_1 _1542_ (.Y(_0593_),
    .A(_0587_),
    .B(_0592_));
 sg13g2_xnor2_1 _1543_ (.Y(_0594_),
    .A(_0582_),
    .B(_0593_));
 sg13g2_a21oi_1 _1544_ (.A1(_0187_),
    .A2(_0504_),
    .Y(_0595_),
    .B1(net37));
 sg13g2_nor2_1 _1545_ (.A(_0187_),
    .B(_0504_),
    .Y(_0596_));
 sg13g2_o21ai_1 _1546_ (.B1(_0127_),
    .Y(_0597_),
    .A1(_0595_),
    .A2(_0596_));
 sg13g2_xnor2_1 _1547_ (.Y(_0598_),
    .A(_0594_),
    .B(_0597_));
 sg13g2_xnor2_1 _1548_ (.Y(_0599_),
    .A(_0570_),
    .B(_0598_));
 sg13g2_a21o_1 _1549_ (.A2(_0541_),
    .A1(_0531_),
    .B1(_0523_),
    .X(_0600_));
 sg13g2_o21ai_1 _1550_ (.B1(_0600_),
    .Y(_0601_),
    .A1(_0531_),
    .A2(_0541_));
 sg13g2_nor2_1 _1551_ (.A(_0078_),
    .B(_0527_),
    .Y(_0602_));
 sg13g2_inv_1 _1552_ (.Y(_0603_),
    .A(_0078_));
 sg13g2_o21ai_1 _1553_ (.B1(_0510_),
    .Y(_0604_),
    .A1(_0603_),
    .A2(_0527_));
 sg13g2_o21ai_1 _1554_ (.B1(_0604_),
    .Y(_0605_),
    .A1(_0281_),
    .A2(_0602_));
 sg13g2_xnor2_1 _1555_ (.Y(_0606_),
    .A(_0078_),
    .B(_0257_));
 sg13g2_a22oi_1 _1556_ (.Y(_0607_),
    .B1(_0606_),
    .B2(_0527_),
    .A2(_0605_),
    .A1(_0090_));
 sg13g2_xor2_1 _1557_ (.B(_0607_),
    .A(_0601_),
    .X(_0608_));
 sg13g2_xnor2_1 _1558_ (.Y(_0609_),
    .A(_0599_),
    .B(_0608_));
 sg13g2_nand3_1 _1559_ (.B(_0561_),
    .C(_0609_),
    .A(_0558_),
    .Y(_0610_));
 sg13g2_a21o_1 _1560_ (.A2(_0561_),
    .A1(_0558_),
    .B1(_0609_),
    .X(_0611_));
 sg13g2_nand3_1 _1561_ (.B(_0610_),
    .C(_0611_),
    .A(_0233_),
    .Y(_0612_));
 sg13g2_a21oi_1 _1562_ (.A1(_0610_),
    .A2(_0611_),
    .Y(_0613_),
    .B1(_0706_));
 sg13g2_o21ai_1 _1563_ (.B1(_0613_),
    .Y(_0614_),
    .A1(_0546_),
    .A2(_0551_));
 sg13g2_o21ai_1 _1564_ (.B1(_0614_),
    .Y(_0011_),
    .A1(_0552_),
    .A2(_0612_));
 sg13g2_and2_1 _1565_ (.A(_0115_),
    .B(net78),
    .X(_0012_));
 sg13g2_buf_1 _1566_ (.A(_0146_),
    .X(_0615_));
 sg13g2_buf_1 _1567_ (.A(_0039_),
    .X(_0616_));
 sg13g2_xor2_1 _1568_ (.B(net57),
    .A(net47),
    .X(_0617_));
 sg13g2_nand2_1 _1569_ (.Y(_0618_),
    .A(net68),
    .B(net74));
 sg13g2_buf_1 _1570_ (.A(_0770_),
    .X(_0619_));
 sg13g2_nand2b_2 _1571_ (.Y(_0620_),
    .B(net56),
    .A_N(net74));
 sg13g2_nand2b_1 _1572_ (.Y(_0621_),
    .B(_0620_),
    .A_N(net72));
 sg13g2_nand2_1 _1573_ (.Y(_0622_),
    .A(_0618_),
    .B(_0621_));
 sg13g2_nand2b_1 _1574_ (.Y(_0623_),
    .B(_0622_),
    .A_N(_0617_));
 sg13g2_buf_1 _1575_ (.A(net72),
    .X(_0624_));
 sg13g2_o21ai_1 _1576_ (.B1(_0617_),
    .Y(_0625_),
    .A1(net56),
    .A2(net55));
 sg13g2_buf_1 _1577_ (.A(net71),
    .X(_0626_));
 sg13g2_a21oi_1 _1578_ (.A1(_0617_),
    .A2(_0620_),
    .Y(_0627_),
    .B1(net54));
 sg13g2_a21o_1 _1579_ (.A2(_0625_),
    .A1(_0623_),
    .B1(_0627_),
    .X(_0628_));
 sg13g2_buf_1 _1580_ (.A(net74),
    .X(_0629_));
 sg13g2_xnor2_1 _1581_ (.Y(_0630_),
    .A(net61),
    .B(net53));
 sg13g2_nand2_1 _1582_ (.Y(_0631_),
    .A(net57),
    .B(net68));
 sg13g2_nand2_1 _1583_ (.Y(_0632_),
    .A(net47),
    .B(_0128_));
 sg13g2_nor2_1 _1584_ (.A(_0157_),
    .B(net72),
    .Y(_0633_));
 sg13g2_nor2_1 _1585_ (.A(net57),
    .B(net68),
    .Y(_0634_));
 sg13g2_a22oi_1 _1586_ (.Y(_0635_),
    .B1(_0633_),
    .B2(_0634_),
    .A2(_0632_),
    .A1(net72));
 sg13g2_o21ai_1 _1587_ (.B1(_0635_),
    .Y(_0636_),
    .A1(net47),
    .A2(_0631_));
 sg13g2_xnor2_1 _1588_ (.Y(_0637_),
    .A(_0630_),
    .B(_0636_));
 sg13g2_nand2_1 _1589_ (.Y(_0638_),
    .A(_0628_),
    .B(_0637_));
 sg13g2_buf_1 _1590_ (.A(\state[0] ),
    .X(_0639_));
 sg13g2_inv_2 _1591_ (.Y(_0640_),
    .A(net70));
 sg13g2_o21ai_1 _1592_ (.B1(_0640_),
    .Y(_0641_),
    .A1(_0628_),
    .A2(_0637_));
 sg13g2_nand2_1 _1593_ (.Y(_0642_),
    .A(_0638_),
    .B(_0641_));
 sg13g2_nor2_1 _1594_ (.A(_0157_),
    .B(net68),
    .Y(_0643_));
 sg13g2_o21ai_1 _1595_ (.B1(_0643_),
    .Y(_0644_),
    .A1(_0616_),
    .A2(net55));
 sg13g2_nand2b_1 _1596_ (.Y(_0645_),
    .B(_0631_),
    .A_N(net55));
 sg13g2_a22oi_1 _1597_ (.Y(_0646_),
    .B1(_0645_),
    .B2(_0157_),
    .A2(net55),
    .A1(_0616_));
 sg13g2_mux2_1 _1598_ (.A0(_0644_),
    .A1(_0646_),
    .S(_0630_),
    .X(_0647_));
 sg13g2_inv_1 _1599_ (.Y(_0648_),
    .A(_0124_));
 sg13g2_xor2_1 _1600_ (.B(_0039_),
    .A(net73),
    .X(_0649_));
 sg13g2_nor2_1 _1601_ (.A(_0242_),
    .B(net53),
    .Y(_0650_));
 sg13g2_nor2_1 _1602_ (.A(net47),
    .B(net68),
    .Y(_0651_));
 sg13g2_nand2_1 _1603_ (.Y(_0652_),
    .A(net47),
    .B(net53));
 sg13g2_a21oi_1 _1604_ (.A1(net56),
    .A2(_0652_),
    .Y(_0653_),
    .B1(net61));
 sg13g2_a221oi_1 _1605_ (.B2(_0651_),
    .C1(_0653_),
    .B1(_0650_),
    .A1(net68),
    .Y(_0654_),
    .A2(net53));
 sg13g2_xnor2_1 _1606_ (.Y(_0655_),
    .A(_0649_),
    .B(_0654_));
 sg13g2_xnor2_1 _1607_ (.Y(_0656_),
    .A(net52),
    .B(_0655_));
 sg13g2_xnor2_1 _1608_ (.Y(_0657_),
    .A(_0647_),
    .B(_0656_));
 sg13g2_xnor2_1 _1609_ (.Y(_0658_),
    .A(_0642_),
    .B(_0657_));
 sg13g2_xor2_1 _1610_ (.B(net71),
    .A(net56),
    .X(_0659_));
 sg13g2_nor2_1 _1611_ (.A(_0063_),
    .B(_0124_),
    .Y(_0660_));
 sg13g2_o21ai_1 _1612_ (.B1(net72),
    .Y(_0661_),
    .A1(net70),
    .A2(_0660_));
 sg13g2_nand2_1 _1613_ (.Y(_0662_),
    .A(net63),
    .B(net70));
 sg13g2_buf_1 _1614_ (.A(_0063_),
    .X(_0663_));
 sg13g2_nor2_1 _1615_ (.A(net72),
    .B(\state[0] ),
    .Y(_0664_));
 sg13g2_nand3_1 _1616_ (.B(_0124_),
    .C(_0664_),
    .A(net51),
    .Y(_0665_));
 sg13g2_nand3_1 _1617_ (.B(_0662_),
    .C(_0665_),
    .A(_0661_),
    .Y(_0666_));
 sg13g2_xnor2_1 _1618_ (.Y(_0667_),
    .A(_0659_),
    .B(_0666_));
 sg13g2_nand2_1 _1619_ (.Y(_0668_),
    .A(net52),
    .B(net70));
 sg13g2_buf_1 _1620_ (.A(_0124_),
    .X(_0669_));
 sg13g2_nand2b_1 _1621_ (.Y(_0670_),
    .B(net50),
    .A_N(_0002_));
 sg13g2_o21ai_1 _1622_ (.B1(_0670_),
    .Y(_0671_),
    .A1(_0115_),
    .A2(_0668_));
 sg13g2_nor3_1 _1623_ (.A(net50),
    .B(_0115_),
    .C(net70),
    .Y(_0672_));
 sg13g2_xnor2_1 _1624_ (.Y(_0673_),
    .A(_0109_),
    .B(net51));
 sg13g2_mux2_1 _1625_ (.A0(_0671_),
    .A1(_0672_),
    .S(_0673_),
    .X(_0674_));
 sg13g2_xor2_1 _1626_ (.B(_0639_),
    .A(_0115_),
    .X(_0675_));
 sg13g2_nand2_1 _1627_ (.Y(_0676_),
    .A(_0002_),
    .B(_0669_));
 sg13g2_o21ai_1 _1628_ (.B1(_0676_),
    .Y(_0677_),
    .A1(net50),
    .A2(_0675_));
 sg13g2_xnor2_1 _1629_ (.Y(_0678_),
    .A(_0673_),
    .B(_0677_));
 sg13g2_nor2_1 _1630_ (.A(_0669_),
    .B(_0639_),
    .Y(_0679_));
 sg13g2_nand2_1 _1631_ (.Y(_0680_),
    .A(_0186_),
    .B(_0679_));
 sg13g2_o21ai_1 _1632_ (.B1(_0680_),
    .Y(_0681_),
    .A1(_0626_),
    .A2(net52));
 sg13g2_nand2_1 _1633_ (.Y(_0682_),
    .A(_0663_),
    .B(_0681_));
 sg13g2_nor2_1 _1634_ (.A(_0678_),
    .B(_0682_),
    .Y(_0683_));
 sg13g2_o21ai_1 _1635_ (.B1(_0683_),
    .Y(_0684_),
    .A1(_0667_),
    .A2(_0674_));
 sg13g2_nor3_1 _1636_ (.A(net63),
    .B(net52),
    .C(_0664_),
    .Y(_0685_));
 sg13g2_a21oi_1 _1637_ (.A1(_0661_),
    .A2(_0662_),
    .Y(_0686_),
    .B1(_0659_));
 sg13g2_a21o_1 _1638_ (.A2(_0685_),
    .A1(_0659_),
    .B1(_0686_),
    .X(_0687_));
 sg13g2_xnor2_1 _1639_ (.Y(_0688_),
    .A(_0146_),
    .B(net72));
 sg13g2_nor2_1 _1640_ (.A(net68),
    .B(net71),
    .Y(_0689_));
 sg13g2_nor2_1 _1641_ (.A(net51),
    .B(net52),
    .Y(_0690_));
 sg13g2_nand2_1 _1642_ (.Y(_0691_),
    .A(net71),
    .B(net51));
 sg13g2_a21oi_1 _1643_ (.A1(net50),
    .A2(_0691_),
    .Y(_0692_),
    .B1(net56));
 sg13g2_a221oi_1 _1644_ (.B2(_0690_),
    .C1(_0692_),
    .B1(_0689_),
    .A1(_0626_),
    .Y(_0693_),
    .A2(_0648_));
 sg13g2_xor2_1 _1645_ (.B(_0693_),
    .A(_0688_),
    .X(_0694_));
 sg13g2_nand2_1 _1646_ (.Y(_0695_),
    .A(_0667_),
    .B(_0674_));
 sg13g2_inv_1 _1647_ (.Y(_0696_),
    .A(_0695_));
 sg13g2_a21oi_1 _1648_ (.A1(_0687_),
    .A2(_0694_),
    .Y(_0697_),
    .B1(_0696_));
 sg13g2_nor2_1 _1649_ (.A(_0687_),
    .B(_0694_),
    .Y(_0698_));
 sg13g2_a21oi_2 _1650_ (.B1(_0698_),
    .Y(_0699_),
    .A2(_0697_),
    .A1(_0684_));
 sg13g2_nand2_2 _1651_ (.Y(_0700_),
    .A(_0620_),
    .B(_0618_));
 sg13g2_nor2_1 _1652_ (.A(net71),
    .B(net63),
    .Y(_0701_));
 sg13g2_nand2_1 _1653_ (.Y(_0702_),
    .A(net72),
    .B(net71));
 sg13g2_a21oi_1 _1654_ (.A1(net51),
    .A2(_0702_),
    .Y(_0703_),
    .B1(_0615_));
 sg13g2_a221oi_1 _1655_ (.B2(_0701_),
    .C1(_0703_),
    .B1(_0633_),
    .A1(net55),
    .Y(_0704_),
    .A2(net63));
 sg13g2_xnor2_1 _1656_ (.Y(_0705_),
    .A(_0700_),
    .B(_0704_));
 sg13g2_nor2_1 _1657_ (.A(net71),
    .B(net51),
    .Y(_0707_));
 sg13g2_o21ai_1 _1658_ (.B1(_0619_),
    .Y(_0708_),
    .A1(_0688_),
    .A2(_0707_));
 sg13g2_nand2_1 _1659_ (.Y(_0709_),
    .A(_0688_),
    .B(_0691_));
 sg13g2_nand2_1 _1660_ (.Y(_0710_),
    .A(_0708_),
    .B(_0709_));
 sg13g2_nor2_1 _1661_ (.A(_0688_),
    .B(_0691_),
    .Y(_0711_));
 sg13g2_a221oi_1 _1662_ (.B2(net50),
    .C1(_0711_),
    .B1(_0710_),
    .A1(_0689_),
    .Y(_0712_),
    .A2(_0688_));
 sg13g2_nand2_1 _1663_ (.Y(_0713_),
    .A(_0705_),
    .B(_0712_));
 sg13g2_inv_1 _1664_ (.Y(_0714_),
    .A(_0713_));
 sg13g2_nor2_1 _1665_ (.A(_0705_),
    .B(_0712_),
    .Y(_0715_));
 sg13g2_nor2_1 _1666_ (.A(_0714_),
    .B(_0715_),
    .Y(_0716_));
 sg13g2_xnor2_1 _1667_ (.Y(_0718_),
    .A(_0640_),
    .B(_0637_));
 sg13g2_xnor2_1 _1668_ (.Y(_0719_),
    .A(_0628_),
    .B(_0718_));
 sg13g2_nor2_1 _1669_ (.A(net54),
    .B(_0620_),
    .Y(_0720_));
 sg13g2_a21oi_1 _1670_ (.A1(net54),
    .A2(_0622_),
    .Y(_0721_),
    .B1(_0720_));
 sg13g2_xor2_1 _1671_ (.B(_0721_),
    .A(_0617_),
    .X(_0722_));
 sg13g2_nor2_1 _1672_ (.A(net55),
    .B(net71),
    .Y(_0723_));
 sg13g2_or2_1 _1673_ (.X(_0724_),
    .B(_0723_),
    .A(_0700_));
 sg13g2_a22oi_1 _1674_ (.Y(_0725_),
    .B1(_0724_),
    .B2(_0615_),
    .A2(_0702_),
    .A1(_0700_));
 sg13g2_nor2_1 _1675_ (.A(_0700_),
    .B(_0702_),
    .Y(_0726_));
 sg13g2_a21oi_1 _1676_ (.A1(_0633_),
    .A2(_0700_),
    .Y(_0727_),
    .B1(_0726_));
 sg13g2_o21ai_1 _1677_ (.B1(_0727_),
    .Y(_0729_),
    .A1(net63),
    .A2(_0725_));
 sg13g2_xnor2_1 _1678_ (.Y(_0730_),
    .A(_0722_),
    .B(_0729_));
 sg13g2_nor2_1 _1679_ (.A(_0719_),
    .B(_0730_),
    .Y(_0731_));
 sg13g2_nand3_1 _1680_ (.B(_0716_),
    .C(_0731_),
    .A(_0699_),
    .Y(_0732_));
 sg13g2_o21ai_1 _1681_ (.B1(_0729_),
    .Y(_0733_),
    .A1(_0715_),
    .A2(_0722_));
 sg13g2_nand2_1 _1682_ (.Y(_0734_),
    .A(_0715_),
    .B(_0722_));
 sg13g2_a21o_1 _1683_ (.A2(_0734_),
    .A1(_0733_),
    .B1(_0719_),
    .X(_0735_));
 sg13g2_nand2_1 _1684_ (.Y(_0736_),
    .A(_0732_),
    .B(_0735_));
 sg13g2_xor2_1 _1685_ (.B(_0736_),
    .A(_0658_),
    .X(_0737_));
 sg13g2_nor2_1 _1686_ (.A(net77),
    .B(_0737_),
    .Y(_0013_));
 sg13g2_nor2_1 _1687_ (.A(_0658_),
    .B(_0735_),
    .Y(_0739_));
 sg13g2_a21oi_1 _1688_ (.A1(_0658_),
    .A2(_0735_),
    .Y(_0740_),
    .B1(_0732_));
 sg13g2_nor2_1 _1689_ (.A(_0739_),
    .B(_0740_),
    .Y(_0741_));
 sg13g2_nor2_1 _1690_ (.A(_0642_),
    .B(_0657_),
    .Y(_0742_));
 sg13g2_nand2_1 _1691_ (.Y(_0743_),
    .A(_0647_),
    .B(_0655_));
 sg13g2_o21ai_1 _1692_ (.B1(net52),
    .Y(_0744_),
    .A1(_0647_),
    .A2(_0655_));
 sg13g2_nand2_1 _1693_ (.Y(_0745_),
    .A(_0743_),
    .B(_0744_));
 sg13g2_xnor2_1 _1694_ (.Y(_0746_),
    .A(net61),
    .B(net58));
 sg13g2_nand2_1 _1695_ (.Y(_0747_),
    .A(_0145_),
    .B(net57));
 sg13g2_nor2_1 _1696_ (.A(net47),
    .B(_0747_),
    .Y(_0748_));
 sg13g2_nor2_1 _1697_ (.A(net57),
    .B(net53),
    .Y(_0750_));
 sg13g2_a21oi_1 _1698_ (.A1(net57),
    .A2(net53),
    .Y(_0751_),
    .B1(_0157_));
 sg13g2_o21ai_1 _1699_ (.B1(_0751_),
    .Y(_0752_),
    .A1(net60),
    .A2(_0750_));
 sg13g2_nand2b_1 _1700_ (.Y(_0753_),
    .B(_0752_),
    .A_N(_0748_));
 sg13g2_xnor2_1 _1701_ (.Y(_0754_),
    .A(_0746_),
    .B(_0753_));
 sg13g2_nor2_1 _1702_ (.A(net47),
    .B(net53),
    .Y(_0755_));
 sg13g2_o21ai_1 _1703_ (.B1(net61),
    .Y(_0756_),
    .A1(_0649_),
    .A2(_0755_));
 sg13g2_nand2_1 _1704_ (.Y(_0757_),
    .A(_0649_),
    .B(_0652_));
 sg13g2_nand2_1 _1705_ (.Y(_0758_),
    .A(_0756_),
    .B(_0757_));
 sg13g2_nor2_1 _1706_ (.A(_0649_),
    .B(_0652_),
    .Y(_0759_));
 sg13g2_a221oi_1 _1707_ (.B2(net56),
    .C1(_0759_),
    .B1(_0758_),
    .A1(_0650_),
    .Y(_0761_),
    .A2(_0649_));
 sg13g2_xnor2_1 _1708_ (.Y(_0762_),
    .A(net63),
    .B(_0761_));
 sg13g2_xnor2_1 _1709_ (.Y(_0763_),
    .A(_0754_),
    .B(_0762_));
 sg13g2_xor2_1 _1710_ (.B(_0763_),
    .A(_0745_),
    .X(_0764_));
 sg13g2_xnor2_1 _1711_ (.Y(_0765_),
    .A(_0742_),
    .B(_0764_));
 sg13g2_nand2_1 _1712_ (.Y(_0766_),
    .A(_0741_),
    .B(_0765_));
 sg13g2_or2_1 _1713_ (.X(_0767_),
    .B(_0765_),
    .A(_0741_));
 sg13g2_buf_1 _1714_ (.A(_0767_),
    .X(_0768_));
 sg13g2_and3_1 _1715_ (.X(_0014_),
    .A(net78),
    .B(_0766_),
    .C(_0768_));
 sg13g2_nand2_1 _1716_ (.Y(_0769_),
    .A(_0742_),
    .B(_0764_));
 sg13g2_or2_1 _1717_ (.X(_0771_),
    .B(_0763_),
    .A(_0745_));
 sg13g2_buf_1 _1718_ (.A(_0771_),
    .X(_0772_));
 sg13g2_xnor2_1 _1719_ (.Y(_0773_),
    .A(net54),
    .B(net70));
 sg13g2_xnor2_1 _1720_ (.Y(_0774_),
    .A(net75),
    .B(net73));
 sg13g2_nor2_1 _1721_ (.A(net58),
    .B(_0128_),
    .Y(_0775_));
 sg13g2_a21oi_1 _1722_ (.A1(net76),
    .A2(_0128_),
    .Y(_0776_),
    .B1(net53));
 sg13g2_nand2_1 _1723_ (.Y(_0777_),
    .A(net58),
    .B(_0629_));
 sg13g2_o21ai_1 _1724_ (.B1(_0777_),
    .Y(_0778_),
    .A1(net61),
    .A2(_0776_));
 sg13g2_a21oi_1 _1725_ (.A1(_0650_),
    .A2(_0775_),
    .Y(_0779_),
    .B1(_0778_));
 sg13g2_xnor2_1 _1726_ (.Y(_0780_),
    .A(_0774_),
    .B(_0779_));
 sg13g2_mux2_1 _1727_ (.A0(_0750_),
    .A1(_0752_),
    .S(_0746_),
    .X(_0782_));
 sg13g2_nor2_1 _1728_ (.A(_0748_),
    .B(_0782_),
    .Y(_0783_));
 sg13g2_xnor2_1 _1729_ (.Y(_0784_),
    .A(_0780_),
    .B(_0783_));
 sg13g2_xnor2_1 _1730_ (.Y(_0785_),
    .A(_0773_),
    .B(_0784_));
 sg13g2_nand2_1 _1731_ (.Y(_0786_),
    .A(_0754_),
    .B(_0761_));
 sg13g2_o21ai_1 _1732_ (.B1(net63),
    .Y(_0787_),
    .A1(_0754_),
    .A2(_0761_));
 sg13g2_nand2_1 _1733_ (.Y(_0788_),
    .A(_0786_),
    .B(_0787_));
 sg13g2_or2_1 _1734_ (.X(_0789_),
    .B(_0788_),
    .A(_0785_));
 sg13g2_nand2_1 _1735_ (.Y(_0790_),
    .A(_0785_),
    .B(_0788_));
 sg13g2_nand2_1 _1736_ (.Y(_0791_),
    .A(_0789_),
    .B(_0790_));
 sg13g2_xnor2_1 _1737_ (.Y(_0793_),
    .A(_0772_),
    .B(_0791_));
 sg13g2_xnor2_1 _1738_ (.Y(_0794_),
    .A(_0769_),
    .B(_0793_));
 sg13g2_xnor2_1 _1739_ (.Y(_0795_),
    .A(_0768_),
    .B(_0794_));
 sg13g2_nand2_1 _1740_ (.Y(_0015_),
    .A(net78),
    .B(_0795_));
 sg13g2_nor2_1 _1741_ (.A(_0780_),
    .B(_0783_),
    .Y(_0796_));
 sg13g2_nand2_1 _1742_ (.Y(_0797_),
    .A(_0780_),
    .B(_0783_));
 sg13g2_o21ai_1 _1743_ (.B1(_0797_),
    .Y(_0798_),
    .A1(_0773_),
    .A2(_0796_));
 sg13g2_nor2_1 _1744_ (.A(net54),
    .B(_0640_),
    .Y(_0799_));
 sg13g2_xnor2_1 _1745_ (.Y(_0800_),
    .A(net55),
    .B(net50));
 sg13g2_xnor2_1 _1746_ (.Y(_0801_),
    .A(_0799_),
    .B(_0800_));
 sg13g2_nor2_1 _1747_ (.A(net58),
    .B(_0629_),
    .Y(_0803_));
 sg13g2_nor4_1 _1748_ (.A(_0242_),
    .B(_0128_),
    .C(_0774_),
    .D(_0803_),
    .Y(_0804_));
 sg13g2_a21oi_2 _1749_ (.B1(_0804_),
    .Y(_0805_),
    .A2(_0778_),
    .A1(_0774_));
 sg13g2_nand2_1 _1750_ (.Y(_0806_),
    .A(net61),
    .B(net73));
 sg13g2_nand2b_1 _1751_ (.Y(_0807_),
    .B(_0806_),
    .A_N(net59));
 sg13g2_o21ai_1 _1752_ (.B1(net59),
    .Y(_0808_),
    .A1(net61),
    .A2(_0747_));
 sg13g2_nor2b_1 _1753_ (.A(net73),
    .B_N(net75),
    .Y(_0809_));
 sg13g2_nor2_1 _1754_ (.A(net57),
    .B(_0809_),
    .Y(_0810_));
 sg13g2_a21oi_1 _1755_ (.A1(_0807_),
    .A2(_0808_),
    .Y(_0811_),
    .B1(_0810_));
 sg13g2_xnor2_1 _1756_ (.Y(_0812_),
    .A(net48),
    .B(net76));
 sg13g2_xnor2_1 _1757_ (.Y(_0814_),
    .A(_0811_),
    .B(_0812_));
 sg13g2_xnor2_1 _1758_ (.Y(_0815_),
    .A(_0805_),
    .B(_0814_));
 sg13g2_xnor2_1 _1759_ (.Y(_0816_),
    .A(_0801_),
    .B(_0815_));
 sg13g2_xor2_1 _1760_ (.B(_0816_),
    .A(_0798_),
    .X(_0817_));
 sg13g2_o21ai_1 _1761_ (.B1(_0788_),
    .Y(_0818_),
    .A1(_0772_),
    .A2(_0785_));
 sg13g2_nand2_1 _1762_ (.Y(_0819_),
    .A(_0772_),
    .B(_0785_));
 sg13g2_a22oi_1 _1763_ (.Y(_0820_),
    .B1(_0818_),
    .B2(_0819_),
    .A2(_0764_),
    .A1(_0742_));
 sg13g2_nor2b_1 _1764_ (.A(_0790_),
    .B_N(_0772_),
    .Y(_0821_));
 sg13g2_a21oi_1 _1765_ (.A1(_0768_),
    .A2(_0820_),
    .Y(_0822_),
    .B1(_0821_));
 sg13g2_xnor2_1 _1766_ (.Y(_0823_),
    .A(_0817_),
    .B(_0822_));
 sg13g2_nor2_1 _1767_ (.A(net77),
    .B(_0823_),
    .Y(_0016_));
 sg13g2_nand2b_1 _1768_ (.Y(_0825_),
    .B(_0790_),
    .A_N(_0772_));
 sg13g2_a21o_1 _1769_ (.A2(_0825_),
    .A1(_0768_),
    .B1(_0821_),
    .X(_0826_));
 sg13g2_nand2_1 _1770_ (.Y(_0827_),
    .A(_0789_),
    .B(_0817_));
 sg13g2_a221oi_1 _1771_ (.B2(_0769_),
    .C1(_0827_),
    .B1(_0826_),
    .A1(_0768_),
    .Y(_0828_),
    .A2(_0821_));
 sg13g2_and2_1 _1772_ (.A(_0798_),
    .B(_0816_),
    .X(_0829_));
 sg13g2_buf_1 _1773_ (.A(_0829_),
    .X(_0830_));
 sg13g2_nor2_1 _1774_ (.A(_0805_),
    .B(_0814_),
    .Y(_0831_));
 sg13g2_nor2_1 _1775_ (.A(_0801_),
    .B(_0831_),
    .Y(_0832_));
 sg13g2_a21oi_1 _1776_ (.A1(_0805_),
    .A2(_0814_),
    .Y(_0833_),
    .B1(_0832_));
 sg13g2_a21o_1 _1777_ (.A2(_0145_),
    .A1(_0242_),
    .B1(_0812_),
    .X(_0835_));
 sg13g2_a22oi_1 _1778_ (.Y(_0836_),
    .B1(_0835_),
    .B2(net59),
    .A2(_0812_),
    .A1(_0806_));
 sg13g2_inv_1 _1779_ (.Y(_0837_),
    .A(_0836_));
 sg13g2_nor2_1 _1780_ (.A(_0806_),
    .B(_0812_),
    .Y(_0838_));
 sg13g2_a221oi_1 _1781_ (.B2(net57),
    .C1(_0838_),
    .B1(_0837_),
    .A1(_0809_),
    .Y(_0839_),
    .A2(_0812_));
 sg13g2_xnor2_1 _1782_ (.Y(_0840_),
    .A(net56),
    .B(net51));
 sg13g2_nand2_1 _1783_ (.Y(_0841_),
    .A(_0624_),
    .B(net70));
 sg13g2_o21ai_1 _1784_ (.B1(_0841_),
    .Y(_0842_),
    .A1(net55),
    .A2(net52));
 sg13g2_xnor2_1 _1785_ (.Y(_0843_),
    .A(_0840_),
    .B(_0842_));
 sg13g2_xor2_1 _1786_ (.B(net49),
    .A(net59),
    .X(_0844_));
 sg13g2_nor2_1 _1787_ (.A(_0738_),
    .B(_0242_),
    .Y(_0846_));
 sg13g2_nor2_1 _1788_ (.A(net60),
    .B(net58),
    .Y(_0847_));
 sg13g2_nand2_1 _1789_ (.Y(_0848_),
    .A(net73),
    .B(net58));
 sg13g2_a21oi_1 _1790_ (.A1(_0241_),
    .A2(_0848_),
    .Y(_0849_),
    .B1(net48));
 sg13g2_a221oi_1 _1791_ (.B2(_0847_),
    .C1(_0849_),
    .B1(_0846_),
    .A1(_0242_),
    .Y(_0850_),
    .A2(net58));
 sg13g2_xor2_1 _1792_ (.B(_0850_),
    .A(_0844_),
    .X(_0851_));
 sg13g2_xor2_1 _1793_ (.B(_0851_),
    .A(_0843_),
    .X(_0852_));
 sg13g2_xnor2_1 _1794_ (.Y(_0853_),
    .A(_0839_),
    .B(_0852_));
 sg13g2_nand3_1 _1795_ (.B(net70),
    .C(_0800_),
    .A(net54),
    .Y(_0854_));
 sg13g2_nor2_1 _1796_ (.A(net52),
    .B(_0640_),
    .Y(_0855_));
 sg13g2_xnor2_1 _1797_ (.Y(_0857_),
    .A(_0854_),
    .B(_0855_));
 sg13g2_xnor2_1 _1798_ (.Y(_0858_),
    .A(_0853_),
    .B(_0857_));
 sg13g2_xnor2_1 _1799_ (.Y(_0859_),
    .A(_0833_),
    .B(_0858_));
 sg13g2_xor2_1 _1800_ (.B(_0859_),
    .A(_0830_),
    .X(_0860_));
 sg13g2_nand2b_1 _1801_ (.Y(_0861_),
    .B(_0817_),
    .A_N(_0789_));
 sg13g2_xnor2_1 _1802_ (.Y(_0862_),
    .A(_0860_),
    .B(_0861_));
 sg13g2_xnor2_1 _1803_ (.Y(_0863_),
    .A(_0828_),
    .B(_0862_));
 sg13g2_nor2_1 _1804_ (.A(net77),
    .B(_0863_),
    .Y(_0017_));
 sg13g2_or2_1 _1805_ (.X(_0864_),
    .B(_0853_),
    .A(_0833_));
 sg13g2_nor2_1 _1806_ (.A(_0830_),
    .B(_0864_),
    .Y(_0865_));
 sg13g2_and2_1 _1807_ (.A(_0833_),
    .B(_0853_),
    .X(_0867_));
 sg13g2_o21ai_1 _1808_ (.B1(_0864_),
    .Y(_0868_),
    .A1(_0830_),
    .A2(_0867_));
 sg13g2_nand2_1 _1809_ (.Y(_0869_),
    .A(_0830_),
    .B(_0867_));
 sg13g2_o21ai_1 _1810_ (.B1(_0869_),
    .Y(_0870_),
    .A1(_0854_),
    .A2(_0868_));
 sg13g2_a21oi_1 _1811_ (.A1(_0854_),
    .A2(_0868_),
    .Y(_0871_),
    .B1(_0865_));
 sg13g2_nor2_1 _1812_ (.A(_0855_),
    .B(_0871_),
    .Y(_0872_));
 sg13g2_a221oi_1 _1813_ (.B2(_0855_),
    .C1(_0872_),
    .B1(_0870_),
    .A1(_0854_),
    .Y(_0873_),
    .A2(_0865_));
 sg13g2_nor2_1 _1814_ (.A(net59),
    .B(_0087_),
    .Y(_0874_));
 sg13g2_or2_1 _1815_ (.X(_0875_),
    .B(_0874_),
    .A(_0534_));
 sg13g2_a22oi_1 _1816_ (.Y(_0876_),
    .B1(_0875_),
    .B2(net60),
    .A2(_0095_),
    .A1(net59));
 sg13g2_xnor2_1 _1817_ (.Y(_0878_),
    .A(net47),
    .B(net54));
 sg13g2_nor2_1 _1818_ (.A(_0834_),
    .B(_0065_),
    .Y(_0879_));
 sg13g2_xnor2_1 _1819_ (.Y(_0880_),
    .A(_0878_),
    .B(_0879_));
 sg13g2_xnor2_1 _1820_ (.Y(_0881_),
    .A(_0876_),
    .B(_0880_));
 sg13g2_nor3_1 _1821_ (.A(_0619_),
    .B(net63),
    .C(net50),
    .Y(_0882_));
 sg13g2_nand2_1 _1822_ (.Y(_0883_),
    .A(net50),
    .B(_0640_));
 sg13g2_a21oi_1 _1823_ (.A1(_0662_),
    .A2(_0883_),
    .Y(_0884_),
    .B1(_0866_));
 sg13g2_a21oi_1 _1824_ (.A1(_0640_),
    .A2(_0690_),
    .Y(_0885_),
    .B1(_0884_));
 sg13g2_nor2b_1 _1825_ (.A(_0885_),
    .B_N(_0624_),
    .Y(_0886_));
 sg13g2_a221oi_1 _1826_ (.B2(_0882_),
    .C1(_0886_),
    .B1(_0841_),
    .A1(net56),
    .Y(_0887_),
    .A2(_0690_));
 sg13g2_xnor2_1 _1827_ (.Y(_0889_),
    .A(_0881_),
    .B(_0887_));
 sg13g2_or2_1 _1828_ (.X(_0890_),
    .B(_0847_),
    .A(_0844_));
 sg13g2_a22oi_1 _1829_ (.Y(_0891_),
    .B1(_0890_),
    .B2(net48),
    .A2(_0848_),
    .A1(_0844_));
 sg13g2_nor2_1 _1830_ (.A(_0844_),
    .B(_0848_),
    .Y(_0892_));
 sg13g2_a21oi_1 _1831_ (.A1(_0092_),
    .A2(_0844_),
    .Y(_0893_),
    .B1(_0892_));
 sg13g2_o21ai_1 _1832_ (.B1(_0893_),
    .Y(_0894_),
    .A1(_0242_),
    .A2(_0891_));
 sg13g2_xnor2_1 _1833_ (.Y(_0895_),
    .A(_0889_),
    .B(_0894_));
 sg13g2_nor2_1 _1834_ (.A(_0843_),
    .B(_0851_),
    .Y(_0896_));
 sg13g2_nand2_1 _1835_ (.Y(_0897_),
    .A(_0843_),
    .B(_0851_));
 sg13g2_o21ai_1 _1836_ (.B1(_0897_),
    .Y(_0898_),
    .A1(_0839_),
    .A2(_0896_));
 sg13g2_xnor2_1 _1837_ (.Y(_0900_),
    .A(_0895_),
    .B(_0898_));
 sg13g2_xnor2_1 _1838_ (.Y(_0901_),
    .A(_0873_),
    .B(_0900_));
 sg13g2_nand3_1 _1839_ (.B(_0822_),
    .C(_0860_),
    .A(_0817_),
    .Y(_0902_));
 sg13g2_xnor2_1 _1840_ (.Y(_0903_),
    .A(_0901_),
    .B(_0902_));
 sg13g2_nor2_1 _1841_ (.A(net77),
    .B(_0903_),
    .Y(_0018_));
 sg13g2_a21oi_1 _1842_ (.A1(_0668_),
    .A2(_0883_),
    .Y(_0019_),
    .B1(_0706_));
 sg13g2_xnor2_1 _1843_ (.Y(_0904_),
    .A(net51),
    .B(_0668_));
 sg13g2_nand2_1 _1844_ (.Y(_0020_),
    .A(net78),
    .B(_0904_));
 sg13g2_a21oi_1 _1845_ (.A1(_0663_),
    .A2(_0679_),
    .Y(_0905_),
    .B1(_0690_));
 sg13g2_xor2_1 _1846_ (.B(_0905_),
    .A(net54),
    .X(_0906_));
 sg13g2_nor2_1 _1847_ (.A(net77),
    .B(_0906_),
    .Y(_0021_));
 sg13g2_xnor2_1 _1848_ (.Y(_0908_),
    .A(_0678_),
    .B(_0682_));
 sg13g2_nor2_1 _1849_ (.A(net77),
    .B(_0908_),
    .Y(_0022_));
 sg13g2_nor2_1 _1850_ (.A(_0683_),
    .B(_0674_),
    .Y(_0909_));
 sg13g2_xnor2_1 _1851_ (.Y(_0910_),
    .A(_0667_),
    .B(_0909_));
 sg13g2_and2_1 _1852_ (.A(net78),
    .B(_0910_),
    .X(_0023_));
 sg13g2_xnor2_1 _1853_ (.Y(_0911_),
    .A(_0687_),
    .B(_0684_));
 sg13g2_nor2_1 _1854_ (.A(_0696_),
    .B(_0911_),
    .Y(_0912_));
 sg13g2_xor2_1 _1855_ (.B(_0912_),
    .A(_0694_),
    .X(_0913_));
 sg13g2_nor2_1 _1856_ (.A(_0706_),
    .B(_0913_),
    .Y(_0024_));
 sg13g2_xnor2_1 _1857_ (.Y(_0915_),
    .A(_0699_),
    .B(_0716_));
 sg13g2_nor2_1 _1858_ (.A(_0706_),
    .B(_0915_),
    .Y(_0025_));
 sg13g2_o21ai_1 _1859_ (.B1(_0713_),
    .Y(_0916_),
    .A1(_0699_),
    .A2(_0715_));
 sg13g2_xnor2_1 _1860_ (.Y(_0917_),
    .A(_0730_),
    .B(_0916_));
 sg13g2_nand2_1 _1861_ (.Y(_0026_),
    .A(net78),
    .B(_0917_));
 sg13g2_nand2_1 _1862_ (.Y(_0918_),
    .A(_0722_),
    .B(_0729_));
 sg13g2_nor2_1 _1863_ (.A(_0722_),
    .B(_0729_),
    .Y(_0919_));
 sg13g2_a21oi_1 _1864_ (.A1(_0916_),
    .A2(_0918_),
    .Y(_0920_),
    .B1(_0919_));
 sg13g2_xor2_1 _1865_ (.B(_0920_),
    .A(_0719_),
    .X(_0921_));
 sg13g2_nor2_1 _1866_ (.A(_0706_),
    .B(_0921_),
    .Y(_0027_));
 sg13g2_xor2_1 _1867_ (.B(\pcg_out[6] ),
    .A(\pcg_out[7] ),
    .X(_0923_));
 sg13g2_nand2_1 _1868_ (.Y(_0924_),
    .A(net15),
    .B(_0923_));
 sg13g2_xor2_1 _1869_ (.B(\pcg_out[4] ),
    .A(\pcg_out[5] ),
    .X(_0925_));
 sg13g2_nand2_1 _1870_ (.Y(_0926_),
    .A(net14),
    .B(_0925_));
 sg13g2_nand2_1 _1871_ (.Y(_0927_),
    .A(net10),
    .B(\pcg_out[0] ));
 sg13g2_xnor2_1 _1872_ (.Y(_0928_),
    .A(net16),
    .B(_0927_));
 sg13g2_xnor2_1 _1873_ (.Y(_0929_),
    .A(_0926_),
    .B(_0928_));
 sg13g2_xnor2_1 _1874_ (.Y(_0930_),
    .A(_0924_),
    .B(_0929_));
 sg13g2_nand2_1 _1875_ (.Y(_0931_),
    .A(net11),
    .B(\pcg_out[1] ));
 sg13g2_nand2_1 _1876_ (.Y(_0932_),
    .A(net12),
    .B(\pcg_out[2] ));
 sg13g2_nand2_1 _1877_ (.Y(_0029_),
    .A(net13),
    .B(\pcg_out[3] ));
 sg13g2_xnor2_1 _1878_ (.Y(_0030_),
    .A(_0932_),
    .B(_0029_));
 sg13g2_xnor2_1 _1879_ (.Y(_0031_),
    .A(_0931_),
    .B(_0030_));
 sg13g2_xnor2_1 _1880_ (.Y(net17),
    .A(_0930_),
    .B(_0031_));
 sg13g2_nand3_1 _1881_ (.B(\pcg_out[7] ),
    .C(net15),
    .A(net13),
    .Y(_0032_));
 sg13g2_xnor2_1 _1882_ (.Y(net18),
    .A(net2),
    .B(_0032_));
 sg13g2_nand3_1 _1883_ (.B(net15),
    .C(\pcg_out[6] ),
    .A(net12),
    .Y(_0033_));
 sg13g2_xnor2_1 _1884_ (.Y(net19),
    .A(net3),
    .B(_0033_));
 sg13g2_nand3_1 _1885_ (.B(net15),
    .C(\pcg_out[5] ),
    .A(net11),
    .Y(_0034_));
 sg13g2_xnor2_1 _1886_ (.Y(net20),
    .A(net4),
    .B(_0034_));
 sg13g2_nand2_1 _1887_ (.Y(_0036_),
    .A(net14),
    .B(\pcg_out[4] ));
 sg13g2_xnor2_1 _1888_ (.Y(net21),
    .A(net5),
    .B(_0036_));
 sg13g2_xnor2_1 _1889_ (.Y(net22),
    .A(net6),
    .B(_0029_));
 sg13g2_xnor2_1 _1890_ (.Y(net23),
    .A(net7),
    .B(_0932_));
 sg13g2_xnor2_1 _1891_ (.Y(net24),
    .A(net8),
    .B(_0931_));
 sg13g2_xnor2_1 _1892_ (.Y(net25),
    .A(net9),
    .B(_0927_));
 sg13g2_buf_1 clkbuf_0_clk (.A(clk),
    .X(clknet_0_clk));
 sg13g2_tiehi _1902__93 (.L_HI(net93));
 sg13g2_buf_1 _1895_ (.A(net79),
    .X(uio_oe[0]));
 sg13g2_buf_1 _1896_ (.A(net80),
    .X(uio_oe[1]));
 sg13g2_buf_1 _1897_ (.A(net81),
    .X(uio_oe[2]));
 sg13g2_buf_1 _1898_ (.A(net82),
    .X(uio_oe[3]));
 sg13g2_buf_1 _1899_ (.A(net83),
    .X(uio_oe[4]));
 sg13g2_buf_1 _1900_ (.A(net84),
    .X(uio_oe[5]));
 sg13g2_buf_1 _1901_ (.A(net85),
    .X(uio_oe[6]));
 sg13g2_buf_1 _1902_ (.A(net93),
    .X(uio_oe[7]));
 sg13g2_buf_1 _1903_ (.A(net86),
    .X(uio_out[0]));
 sg13g2_buf_1 _1904_ (.A(net87),
    .X(uio_out[1]));
 sg13g2_buf_1 _1905_ (.A(net88),
    .X(uio_out[2]));
 sg13g2_buf_1 _1906_ (.A(net89),
    .X(uio_out[3]));
 sg13g2_buf_1 _1907_ (.A(net90),
    .X(uio_out[4]));
 sg13g2_buf_1 _1908_ (.A(net91),
    .X(uio_out[5]));
 sg13g2_buf_1 _1909_ (.A(net92),
    .X(uio_out[6]));
 sg13g2_dfrbp_1 \pcg_out[0]$_SDFF_PN0_  (.CLK(clknet_2_3__leaf_clk),
    .RESET_B(net94),
    .D(_0004_),
    .Q_N(_0952_),
    .Q(\pcg_out[0] ));
 sg13g2_dfrbp_1 \pcg_out[1]$_SDFF_PN0_  (.CLK(clknet_2_3__leaf_clk),
    .RESET_B(net95),
    .D(_0005_),
    .Q_N(_0951_),
    .Q(\pcg_out[1] ));
 sg13g2_dfrbp_1 \pcg_out[2]$_SDFF_PN0_  (.CLK(clknet_2_3__leaf_clk),
    .RESET_B(net96),
    .D(_0006_),
    .Q_N(_0950_),
    .Q(\pcg_out[2] ));
 sg13g2_dfrbp_1 \pcg_out[3]$_SDFF_PN0_  (.CLK(clknet_2_3__leaf_clk),
    .RESET_B(net97),
    .D(_0007_),
    .Q_N(_0949_),
    .Q(\pcg_out[3] ));
 sg13g2_dfrbp_1 \pcg_out[4]$_SDFF_PN0_  (.CLK(clknet_2_2__leaf_clk),
    .RESET_B(net98),
    .D(_0008_),
    .Q_N(_0948_),
    .Q(\pcg_out[4] ));
 sg13g2_dfrbp_1 \pcg_out[5]$_SDFF_PN0_  (.CLK(clknet_2_2__leaf_clk),
    .RESET_B(net99),
    .D(_0009_),
    .Q_N(_0947_),
    .Q(\pcg_out[5] ));
 sg13g2_dfrbp_1 \pcg_out[6]$_SDFF_PN0_  (.CLK(clknet_2_3__leaf_clk),
    .RESET_B(net100),
    .D(_0010_),
    .Q_N(_0946_),
    .Q(\pcg_out[6] ));
 sg13g2_dfrbp_1 \pcg_out[7]$_SDFF_PN0_  (.CLK(clknet_2_3__leaf_clk),
    .RESET_B(net101),
    .D(_0011_),
    .Q_N(_0945_),
    .Q(\pcg_out[7] ));
 sg13g2_dfrbp_1 \state[0]$_SDFF_PN0_  (.CLK(clknet_2_2__leaf_clk),
    .RESET_B(net102),
    .D(_0012_),
    .Q_N(_0003_),
    .Q(\state[0] ));
 sg13g2_dfrbp_1 \state[10]$_SDFF_PN0_  (.CLK(clknet_2_1__leaf_clk),
    .RESET_B(net103),
    .D(_0013_),
    .Q_N(_0944_),
    .Q(\state[10] ));
 sg13g2_dfrbp_1 \state[11]$_SDFF_PN0_  (.CLK(clknet_2_0__leaf_clk),
    .RESET_B(net104),
    .D(_0014_),
    .Q_N(_0943_),
    .Q(\state[11] ));
 sg13g2_dfrbp_1 \state[12]$_SDFF_PN1_  (.CLK(clknet_2_0__leaf_clk),
    .RESET_B(net105),
    .D(_0015_),
    .Q_N(_0942_),
    .Q(\state[12] ));
 sg13g2_dfrbp_1 \state[13]$_SDFF_PN0_  (.CLK(clknet_2_0__leaf_clk),
    .RESET_B(net106),
    .D(_0016_),
    .Q_N(_0941_),
    .Q(\state[13] ));
 sg13g2_dfrbp_1 \state[14]$_SDFF_PN0_  (.CLK(clknet_2_0__leaf_clk),
    .RESET_B(net107),
    .D(_0017_),
    .Q_N(_0940_),
    .Q(\state[14] ));
 sg13g2_dfrbp_1 \state[15]$_SDFF_PN0_  (.CLK(clknet_2_0__leaf_clk),
    .RESET_B(net108),
    .D(_0018_),
    .Q_N(_0939_),
    .Q(\state[15] ));
 sg13g2_dfrbp_1 \state[1]$_SDFF_PN0_  (.CLK(clknet_2_2__leaf_clk),
    .RESET_B(net109),
    .D(_0019_),
    .Q_N(_0001_),
    .Q(\state[1] ));
 sg13g2_dfrbp_1 \state[2]$_SDFF_PN1_  (.CLK(clknet_2_2__leaf_clk),
    .RESET_B(net110),
    .D(_0020_),
    .Q_N(_0000_),
    .Q(\state[2] ));
 sg13g2_dfrbp_1 \state[3]$_SDFF_PN0_  (.CLK(clknet_2_0__leaf_clk),
    .RESET_B(net111),
    .D(_0021_),
    .Q_N(_0002_),
    .Q(\state[3] ));
 sg13g2_dfrbp_1 \state[4]$_SDFF_PN0_  (.CLK(clknet_2_2__leaf_clk),
    .RESET_B(net112),
    .D(_0022_),
    .Q_N(_0938_),
    .Q(\state[4] ));
 sg13g2_dfrbp_1 \state[5]$_SDFF_PN0_  (.CLK(clknet_2_1__leaf_clk),
    .RESET_B(net113),
    .D(_0023_),
    .Q_N(_0937_),
    .Q(\state[5] ));
 sg13g2_dfrbp_1 \state[6]$_SDFF_PN0_  (.CLK(clknet_2_1__leaf_clk),
    .RESET_B(net114),
    .D(_0024_),
    .Q_N(_0936_),
    .Q(\state[6] ));
 sg13g2_dfrbp_1 \state[7]$_SDFF_PN0_  (.CLK(clknet_2_1__leaf_clk),
    .RESET_B(net115),
    .D(_0025_),
    .Q_N(_0935_),
    .Q(\state[7] ));
 sg13g2_dfrbp_1 \state[8]$_SDFF_PN1_  (.CLK(clknet_2_1__leaf_clk),
    .RESET_B(net116),
    .D(_0026_),
    .Q_N(_0934_),
    .Q(\state[8] ));
 sg13g2_dfrbp_1 \state[9]$_SDFF_PN0_  (.CLK(clknet_2_1__leaf_clk),
    .RESET_B(net117),
    .D(_0027_),
    .Q_N(_0933_),
    .Q(\state[9] ));
 sg13g2_buf_1 input1 (.A(rst_n),
    .X(net1));
 sg13g2_buf_1 input2 (.A(ui_in[0]),
    .X(net2));
 sg13g2_buf_1 input3 (.A(ui_in[1]),
    .X(net3));
 sg13g2_buf_1 input4 (.A(ui_in[2]),
    .X(net4));
 sg13g2_buf_1 input5 (.A(ui_in[3]),
    .X(net5));
 sg13g2_buf_1 input6 (.A(ui_in[4]),
    .X(net6));
 sg13g2_buf_1 input7 (.A(ui_in[5]),
    .X(net7));
 sg13g2_buf_1 input8 (.A(ui_in[6]),
    .X(net8));
 sg13g2_buf_1 input9 (.A(ui_in[7]),
    .X(net9));
 sg13g2_buf_1 input10 (.A(uio_in[0]),
    .X(net10));
 sg13g2_buf_1 input11 (.A(uio_in[1]),
    .X(net11));
 sg13g2_buf_1 input12 (.A(uio_in[2]),
    .X(net12));
 sg13g2_buf_1 input13 (.A(uio_in[3]),
    .X(net13));
 sg13g2_buf_1 input14 (.A(uio_in[4]),
    .X(net14));
 sg13g2_buf_1 input15 (.A(uio_in[5]),
    .X(net15));
 sg13g2_buf_1 input16 (.A(uio_in[6]),
    .X(net16));
 sg13g2_buf_1 output17 (.A(net17),
    .X(uio_out[7]));
 sg13g2_buf_1 output18 (.A(net18),
    .X(uo_out[0]));
 sg13g2_buf_1 output19 (.A(net19),
    .X(uo_out[1]));
 sg13g2_buf_1 output20 (.A(net20),
    .X(uo_out[2]));
 sg13g2_buf_1 output21 (.A(net21),
    .X(uo_out[3]));
 sg13g2_buf_1 output22 (.A(net22),
    .X(uo_out[4]));
 sg13g2_buf_1 output23 (.A(net23),
    .X(uo_out[5]));
 sg13g2_buf_1 output24 (.A(net24),
    .X(uo_out[6]));
 sg13g2_buf_1 output25 (.A(net25),
    .X(uo_out[7]));
 sg13g2_buf_2 fanout26 (.A(_0355_),
    .X(net26));
 sg13g2_buf_2 fanout27 (.A(_0263_),
    .X(net27));
 sg13g2_buf_2 fanout28 (.A(_0257_),
    .X(net28));
 sg13g2_buf_2 fanout29 (.A(_0249_),
    .X(net29));
 sg13g2_buf_2 fanout30 (.A(_0191_),
    .X(net30));
 sg13g2_buf_2 fanout31 (.A(_0182_),
    .X(net31));
 sg13g2_buf_2 fanout32 (.A(_0108_),
    .X(net32));
 sg13g2_buf_2 fanout33 (.A(_0234_),
    .X(net33));
 sg13g2_buf_2 fanout34 (.A(_0207_),
    .X(net34));
 sg13g2_buf_2 fanout35 (.A(_0195_),
    .X(net35));
 sg13g2_buf_2 fanout36 (.A(_0194_),
    .X(net36));
 sg13g2_buf_2 fanout37 (.A(_0181_),
    .X(net37));
 sg13g2_buf_2 fanout38 (.A(_0174_),
    .X(net38));
 sg13g2_buf_2 fanout39 (.A(_0123_),
    .X(net39));
 sg13g2_buf_2 fanout40 (.A(_0309_),
    .X(net40));
 sg13g2_buf_2 fanout41 (.A(_0245_),
    .X(net41));
 sg13g2_buf_2 fanout42 (.A(_0184_),
    .X(net42));
 sg13g2_buf_2 fanout43 (.A(_0112_),
    .X(net43));
 sg13g2_buf_2 fanout44 (.A(_0111_),
    .X(net44));
 sg13g2_buf_2 fanout45 (.A(_0090_),
    .X(net45));
 sg13g2_buf_2 fanout46 (.A(_0047_),
    .X(net46));
 sg13g2_buf_2 fanout47 (.A(_0615_),
    .X(net47));
 sg13g2_buf_2 fanout48 (.A(_0129_),
    .X(net48));
 sg13g2_buf_2 fanout49 (.A(_0051_),
    .X(net49));
 sg13g2_buf_2 fanout50 (.A(_0669_),
    .X(net50));
 sg13g2_buf_2 fanout51 (.A(_0663_),
    .X(net51));
 sg13g2_buf_2 fanout52 (.A(_0648_),
    .X(net52));
 sg13g2_buf_2 fanout53 (.A(_0629_),
    .X(net53));
 sg13g2_buf_2 fanout54 (.A(_0626_),
    .X(net54));
 sg13g2_buf_2 fanout55 (.A(_0624_),
    .X(net55));
 sg13g2_buf_2 fanout56 (.A(_0619_),
    .X(net56));
 sg13g2_buf_2 fanout57 (.A(_0616_),
    .X(net57));
 sg13g2_buf_2 fanout58 (.A(_0458_),
    .X(net58));
 sg13g2_buf_2 fanout59 (.A(_0424_),
    .X(net59));
 sg13g2_buf_2 fanout60 (.A(_0359_),
    .X(net60));
 sg13g2_buf_2 fanout61 (.A(_0241_),
    .X(net61));
 sg13g2_buf_2 fanout62 (.A(_0146_),
    .X(net62));
 sg13g2_buf_2 fanout63 (.A(_0064_),
    .X(net63));
 sg13g2_buf_2 fanout64 (.A(_0042_),
    .X(net64));
 sg13g2_buf_2 fanout65 (.A(_0922_),
    .X(net65));
 sg13g2_buf_2 fanout66 (.A(_0899_),
    .X(net66));
 sg13g2_buf_2 fanout67 (.A(_0877_),
    .X(net67));
 sg13g2_buf_2 fanout68 (.A(_0866_),
    .X(net68));
 sg13g2_buf_2 fanout69 (.A(_0760_),
    .X(net69));
 sg13g2_buf_2 fanout70 (.A(_0639_),
    .X(net70));
 sg13g2_buf_2 fanout71 (.A(_0186_),
    .X(net71));
 sg13g2_buf_2 fanout72 (.A(_0109_),
    .X(net72));
 sg13g2_buf_2 fanout73 (.A(_0094_),
    .X(net73));
 sg13g2_buf_2 fanout74 (.A(_0049_),
    .X(net74));
 sg13g2_buf_2 fanout75 (.A(_0888_),
    .X(net75));
 sg13g2_buf_2 fanout76 (.A(_0792_),
    .X(net76));
 sg13g2_buf_2 fanout77 (.A(_0717_),
    .X(net77));
 sg13g2_buf_2 fanout78 (.A(_0233_),
    .X(net78));
 sg13g2_tielo _1895__79 (.L_LO(net79));
 sg13g2_tielo _1896__80 (.L_LO(net80));
 sg13g2_tielo _1897__81 (.L_LO(net81));
 sg13g2_tielo _1898__82 (.L_LO(net82));
 sg13g2_tielo _1899__83 (.L_LO(net83));
 sg13g2_tielo _1900__84 (.L_LO(net84));
 sg13g2_tielo _1901__85 (.L_LO(net85));
 sg13g2_tielo _1903__86 (.L_LO(net86));
 sg13g2_tielo _1904__87 (.L_LO(net87));
 sg13g2_tielo _1905__88 (.L_LO(net88));
 sg13g2_tielo _1906__89 (.L_LO(net89));
 sg13g2_tielo _1907__90 (.L_LO(net90));
 sg13g2_tielo _1908__91 (.L_LO(net91));
 sg13g2_tielo _1909__92 (.L_LO(net92));
 sg13g2_tiehi \pcg_out[0]$_SDFF_PN0__94  (.L_HI(net94));
 sg13g2_tiehi \pcg_out[1]$_SDFF_PN0__95  (.L_HI(net95));
 sg13g2_tiehi \pcg_out[2]$_SDFF_PN0__96  (.L_HI(net96));
 sg13g2_tiehi \pcg_out[3]$_SDFF_PN0__97  (.L_HI(net97));
 sg13g2_tiehi \pcg_out[4]$_SDFF_PN0__98  (.L_HI(net98));
 sg13g2_tiehi \pcg_out[5]$_SDFF_PN0__99  (.L_HI(net99));
 sg13g2_tiehi \pcg_out[6]$_SDFF_PN0__100  (.L_HI(net100));
 sg13g2_tiehi \pcg_out[7]$_SDFF_PN0__101  (.L_HI(net101));
 sg13g2_tiehi \state[0]$_SDFF_PN0__102  (.L_HI(net102));
 sg13g2_tiehi \state[10]$_SDFF_PN0__103  (.L_HI(net103));
 sg13g2_tiehi \state[11]$_SDFF_PN0__104  (.L_HI(net104));
 sg13g2_tiehi \state[12]$_SDFF_PN1__105  (.L_HI(net105));
 sg13g2_tiehi \state[13]$_SDFF_PN0__106  (.L_HI(net106));
 sg13g2_tiehi \state[14]$_SDFF_PN0__107  (.L_HI(net107));
 sg13g2_tiehi \state[15]$_SDFF_PN0__108  (.L_HI(net108));
 sg13g2_tiehi \state[1]$_SDFF_PN0__109  (.L_HI(net109));
 sg13g2_tiehi \state[2]$_SDFF_PN1__110  (.L_HI(net110));
 sg13g2_tiehi \state[3]$_SDFF_PN0__111  (.L_HI(net111));
 sg13g2_tiehi \state[4]$_SDFF_PN0__112  (.L_HI(net112));
 sg13g2_tiehi \state[5]$_SDFF_PN0__113  (.L_HI(net113));
 sg13g2_tiehi \state[6]$_SDFF_PN0__114  (.L_HI(net114));
 sg13g2_tiehi \state[7]$_SDFF_PN0__115  (.L_HI(net115));
 sg13g2_tiehi \state[8]$_SDFF_PN1__116  (.L_HI(net116));
 sg13g2_tiehi \state[9]$_SDFF_PN0__117  (.L_HI(net117));
 sg13g2_buf_1 clkbuf_2_0__f_clk (.A(clknet_0_clk),
    .X(clknet_2_0__leaf_clk));
 sg13g2_buf_1 clkbuf_2_1__f_clk (.A(clknet_0_clk),
    .X(clknet_2_1__leaf_clk));
 sg13g2_buf_1 clkbuf_2_2__f_clk (.A(clknet_0_clk),
    .X(clknet_2_2__leaf_clk));
 sg13g2_buf_1 clkbuf_2_3__f_clk (.A(clknet_0_clk),
    .X(clknet_2_3__leaf_clk));
 sg13g2_decap_8 FILLER_0_0 ();
 sg13g2_decap_8 FILLER_0_7 ();
 sg13g2_decap_8 FILLER_0_14 ();
 sg13g2_decap_8 FILLER_0_21 ();
 sg13g2_decap_8 FILLER_0_28 ();
 sg13g2_decap_8 FILLER_0_35 ();
 sg13g2_decap_8 FILLER_0_42 ();
 sg13g2_decap_8 FILLER_0_49 ();
 sg13g2_decap_8 FILLER_0_56 ();
 sg13g2_decap_8 FILLER_0_63 ();
 sg13g2_decap_8 FILLER_0_70 ();
 sg13g2_decap_8 FILLER_0_77 ();
 sg13g2_decap_8 FILLER_0_84 ();
 sg13g2_decap_8 FILLER_0_91 ();
 sg13g2_decap_8 FILLER_0_98 ();
 sg13g2_decap_8 FILLER_0_105 ();
 sg13g2_decap_8 FILLER_0_112 ();
 sg13g2_decap_8 FILLER_0_119 ();
 sg13g2_decap_8 FILLER_0_126 ();
 sg13g2_decap_8 FILLER_0_133 ();
 sg13g2_decap_8 FILLER_0_140 ();
 sg13g2_decap_8 FILLER_0_147 ();
 sg13g2_decap_8 FILLER_0_154 ();
 sg13g2_decap_8 FILLER_0_161 ();
 sg13g2_decap_8 FILLER_0_168 ();
 sg13g2_decap_8 FILLER_0_175 ();
 sg13g2_decap_8 FILLER_0_182 ();
 sg13g2_decap_8 FILLER_0_189 ();
 sg13g2_decap_8 FILLER_0_196 ();
 sg13g2_decap_8 FILLER_0_203 ();
 sg13g2_decap_8 FILLER_0_210 ();
 sg13g2_decap_8 FILLER_0_217 ();
 sg13g2_decap_8 FILLER_0_224 ();
 sg13g2_decap_8 FILLER_0_231 ();
 sg13g2_decap_8 FILLER_0_238 ();
 sg13g2_decap_8 FILLER_0_245 ();
 sg13g2_decap_8 FILLER_0_252 ();
 sg13g2_decap_8 FILLER_0_259 ();
 sg13g2_decap_8 FILLER_0_266 ();
 sg13g2_decap_8 FILLER_0_273 ();
 sg13g2_decap_8 FILLER_0_280 ();
 sg13g2_decap_8 FILLER_0_287 ();
 sg13g2_decap_8 FILLER_0_294 ();
 sg13g2_decap_8 FILLER_0_301 ();
 sg13g2_decap_8 FILLER_0_308 ();
 sg13g2_decap_8 FILLER_0_315 ();
 sg13g2_decap_8 FILLER_0_322 ();
 sg13g2_decap_8 FILLER_0_329 ();
 sg13g2_decap_8 FILLER_0_336 ();
 sg13g2_decap_8 FILLER_0_343 ();
 sg13g2_decap_8 FILLER_0_350 ();
 sg13g2_decap_8 FILLER_0_357 ();
 sg13g2_decap_8 FILLER_0_364 ();
 sg13g2_decap_8 FILLER_0_371 ();
 sg13g2_decap_8 FILLER_0_378 ();
 sg13g2_decap_8 FILLER_0_385 ();
 sg13g2_decap_8 FILLER_0_392 ();
 sg13g2_decap_8 FILLER_0_399 ();
 sg13g2_decap_8 FILLER_0_406 ();
 sg13g2_decap_8 FILLER_0_413 ();
 sg13g2_decap_8 FILLER_0_420 ();
 sg13g2_fill_2 FILLER_0_427 ();
 sg13g2_fill_1 FILLER_0_429 ();
 sg13g2_decap_8 FILLER_1_0 ();
 sg13g2_decap_8 FILLER_1_7 ();
 sg13g2_decap_8 FILLER_1_14 ();
 sg13g2_decap_8 FILLER_1_21 ();
 sg13g2_decap_8 FILLER_1_28 ();
 sg13g2_decap_8 FILLER_1_35 ();
 sg13g2_decap_8 FILLER_1_42 ();
 sg13g2_decap_8 FILLER_1_49 ();
 sg13g2_decap_8 FILLER_1_56 ();
 sg13g2_decap_8 FILLER_1_63 ();
 sg13g2_decap_8 FILLER_1_70 ();
 sg13g2_decap_8 FILLER_1_77 ();
 sg13g2_decap_8 FILLER_1_84 ();
 sg13g2_decap_8 FILLER_1_91 ();
 sg13g2_decap_8 FILLER_1_98 ();
 sg13g2_decap_8 FILLER_1_105 ();
 sg13g2_decap_8 FILLER_1_112 ();
 sg13g2_decap_8 FILLER_1_119 ();
 sg13g2_decap_8 FILLER_1_126 ();
 sg13g2_decap_8 FILLER_1_133 ();
 sg13g2_decap_8 FILLER_1_140 ();
 sg13g2_decap_8 FILLER_1_147 ();
 sg13g2_decap_8 FILLER_1_154 ();
 sg13g2_decap_8 FILLER_1_161 ();
 sg13g2_decap_8 FILLER_1_168 ();
 sg13g2_decap_8 FILLER_1_175 ();
 sg13g2_decap_8 FILLER_1_182 ();
 sg13g2_decap_8 FILLER_1_189 ();
 sg13g2_decap_8 FILLER_1_196 ();
 sg13g2_decap_8 FILLER_1_203 ();
 sg13g2_decap_8 FILLER_1_210 ();
 sg13g2_decap_8 FILLER_1_217 ();
 sg13g2_decap_8 FILLER_1_224 ();
 sg13g2_decap_8 FILLER_1_231 ();
 sg13g2_decap_8 FILLER_1_238 ();
 sg13g2_decap_8 FILLER_1_245 ();
 sg13g2_decap_8 FILLER_1_252 ();
 sg13g2_decap_8 FILLER_1_259 ();
 sg13g2_decap_8 FILLER_1_266 ();
 sg13g2_decap_8 FILLER_1_273 ();
 sg13g2_decap_8 FILLER_1_280 ();
 sg13g2_decap_8 FILLER_1_287 ();
 sg13g2_decap_8 FILLER_1_294 ();
 sg13g2_decap_8 FILLER_1_301 ();
 sg13g2_decap_8 FILLER_1_308 ();
 sg13g2_decap_8 FILLER_1_315 ();
 sg13g2_decap_8 FILLER_1_322 ();
 sg13g2_decap_8 FILLER_1_329 ();
 sg13g2_decap_8 FILLER_1_336 ();
 sg13g2_decap_8 FILLER_1_343 ();
 sg13g2_decap_8 FILLER_1_350 ();
 sg13g2_decap_8 FILLER_1_357 ();
 sg13g2_decap_8 FILLER_1_364 ();
 sg13g2_decap_8 FILLER_1_371 ();
 sg13g2_decap_8 FILLER_1_378 ();
 sg13g2_decap_8 FILLER_1_385 ();
 sg13g2_decap_8 FILLER_1_392 ();
 sg13g2_decap_8 FILLER_1_399 ();
 sg13g2_decap_8 FILLER_1_406 ();
 sg13g2_decap_8 FILLER_1_413 ();
 sg13g2_decap_8 FILLER_1_420 ();
 sg13g2_fill_2 FILLER_1_427 ();
 sg13g2_fill_1 FILLER_1_429 ();
 sg13g2_decap_8 FILLER_2_0 ();
 sg13g2_decap_8 FILLER_2_7 ();
 sg13g2_decap_8 FILLER_2_14 ();
 sg13g2_decap_8 FILLER_2_21 ();
 sg13g2_decap_8 FILLER_2_28 ();
 sg13g2_decap_8 FILLER_2_35 ();
 sg13g2_decap_8 FILLER_2_42 ();
 sg13g2_decap_8 FILLER_2_49 ();
 sg13g2_decap_8 FILLER_2_56 ();
 sg13g2_decap_8 FILLER_2_63 ();
 sg13g2_decap_8 FILLER_2_70 ();
 sg13g2_decap_8 FILLER_2_77 ();
 sg13g2_decap_8 FILLER_2_84 ();
 sg13g2_decap_8 FILLER_2_91 ();
 sg13g2_decap_8 FILLER_2_98 ();
 sg13g2_decap_8 FILLER_2_105 ();
 sg13g2_decap_8 FILLER_2_112 ();
 sg13g2_decap_8 FILLER_2_119 ();
 sg13g2_decap_8 FILLER_2_126 ();
 sg13g2_decap_8 FILLER_2_133 ();
 sg13g2_decap_8 FILLER_2_140 ();
 sg13g2_decap_8 FILLER_2_147 ();
 sg13g2_decap_8 FILLER_2_154 ();
 sg13g2_decap_8 FILLER_2_161 ();
 sg13g2_decap_8 FILLER_2_168 ();
 sg13g2_decap_8 FILLER_2_175 ();
 sg13g2_decap_8 FILLER_2_182 ();
 sg13g2_decap_8 FILLER_2_189 ();
 sg13g2_decap_8 FILLER_2_196 ();
 sg13g2_decap_8 FILLER_2_203 ();
 sg13g2_decap_8 FILLER_2_210 ();
 sg13g2_decap_8 FILLER_2_217 ();
 sg13g2_decap_8 FILLER_2_224 ();
 sg13g2_decap_8 FILLER_2_231 ();
 sg13g2_decap_8 FILLER_2_238 ();
 sg13g2_decap_8 FILLER_2_245 ();
 sg13g2_decap_8 FILLER_2_252 ();
 sg13g2_decap_8 FILLER_2_259 ();
 sg13g2_decap_8 FILLER_2_266 ();
 sg13g2_decap_8 FILLER_2_273 ();
 sg13g2_decap_8 FILLER_2_280 ();
 sg13g2_decap_8 FILLER_2_287 ();
 sg13g2_decap_8 FILLER_2_294 ();
 sg13g2_decap_8 FILLER_2_301 ();
 sg13g2_decap_8 FILLER_2_308 ();
 sg13g2_decap_8 FILLER_2_315 ();
 sg13g2_decap_8 FILLER_2_322 ();
 sg13g2_decap_8 FILLER_2_329 ();
 sg13g2_decap_8 FILLER_2_336 ();
 sg13g2_decap_8 FILLER_2_343 ();
 sg13g2_decap_8 FILLER_2_350 ();
 sg13g2_decap_8 FILLER_2_357 ();
 sg13g2_decap_8 FILLER_2_364 ();
 sg13g2_decap_8 FILLER_2_371 ();
 sg13g2_decap_8 FILLER_2_378 ();
 sg13g2_decap_8 FILLER_2_385 ();
 sg13g2_decap_8 FILLER_2_392 ();
 sg13g2_decap_8 FILLER_2_399 ();
 sg13g2_decap_8 FILLER_2_406 ();
 sg13g2_decap_8 FILLER_2_413 ();
 sg13g2_decap_8 FILLER_2_420 ();
 sg13g2_fill_2 FILLER_2_427 ();
 sg13g2_fill_1 FILLER_2_429 ();
 sg13g2_decap_8 FILLER_3_0 ();
 sg13g2_decap_8 FILLER_3_7 ();
 sg13g2_decap_8 FILLER_3_14 ();
 sg13g2_decap_8 FILLER_3_21 ();
 sg13g2_decap_8 FILLER_3_28 ();
 sg13g2_decap_8 FILLER_3_35 ();
 sg13g2_decap_8 FILLER_3_42 ();
 sg13g2_decap_8 FILLER_3_49 ();
 sg13g2_decap_8 FILLER_3_56 ();
 sg13g2_decap_8 FILLER_3_63 ();
 sg13g2_decap_8 FILLER_3_70 ();
 sg13g2_decap_8 FILLER_3_77 ();
 sg13g2_decap_8 FILLER_3_84 ();
 sg13g2_decap_8 FILLER_3_91 ();
 sg13g2_decap_8 FILLER_3_98 ();
 sg13g2_decap_8 FILLER_3_105 ();
 sg13g2_decap_8 FILLER_3_112 ();
 sg13g2_decap_8 FILLER_3_119 ();
 sg13g2_decap_8 FILLER_3_126 ();
 sg13g2_decap_8 FILLER_3_133 ();
 sg13g2_decap_8 FILLER_3_140 ();
 sg13g2_decap_8 FILLER_3_147 ();
 sg13g2_decap_8 FILLER_3_154 ();
 sg13g2_decap_8 FILLER_3_161 ();
 sg13g2_decap_8 FILLER_3_168 ();
 sg13g2_decap_8 FILLER_3_175 ();
 sg13g2_decap_8 FILLER_3_182 ();
 sg13g2_decap_8 FILLER_3_189 ();
 sg13g2_decap_8 FILLER_3_196 ();
 sg13g2_decap_8 FILLER_3_203 ();
 sg13g2_decap_8 FILLER_3_210 ();
 sg13g2_decap_8 FILLER_3_217 ();
 sg13g2_decap_8 FILLER_3_224 ();
 sg13g2_decap_8 FILLER_3_231 ();
 sg13g2_decap_8 FILLER_3_238 ();
 sg13g2_decap_8 FILLER_3_245 ();
 sg13g2_decap_8 FILLER_3_252 ();
 sg13g2_decap_8 FILLER_3_259 ();
 sg13g2_decap_8 FILLER_3_266 ();
 sg13g2_decap_8 FILLER_3_273 ();
 sg13g2_decap_8 FILLER_3_280 ();
 sg13g2_decap_8 FILLER_3_287 ();
 sg13g2_decap_8 FILLER_3_294 ();
 sg13g2_decap_8 FILLER_3_301 ();
 sg13g2_decap_8 FILLER_3_308 ();
 sg13g2_decap_8 FILLER_3_315 ();
 sg13g2_decap_8 FILLER_3_322 ();
 sg13g2_decap_8 FILLER_3_329 ();
 sg13g2_decap_8 FILLER_3_336 ();
 sg13g2_decap_8 FILLER_3_343 ();
 sg13g2_decap_8 FILLER_3_350 ();
 sg13g2_decap_8 FILLER_3_357 ();
 sg13g2_decap_8 FILLER_3_364 ();
 sg13g2_decap_8 FILLER_3_371 ();
 sg13g2_decap_8 FILLER_3_378 ();
 sg13g2_decap_8 FILLER_3_385 ();
 sg13g2_decap_8 FILLER_3_392 ();
 sg13g2_decap_8 FILLER_3_399 ();
 sg13g2_decap_8 FILLER_3_406 ();
 sg13g2_decap_8 FILLER_3_413 ();
 sg13g2_decap_8 FILLER_3_420 ();
 sg13g2_fill_2 FILLER_3_427 ();
 sg13g2_fill_1 FILLER_3_429 ();
 sg13g2_decap_8 FILLER_4_0 ();
 sg13g2_decap_8 FILLER_4_7 ();
 sg13g2_decap_8 FILLER_4_14 ();
 sg13g2_decap_8 FILLER_4_21 ();
 sg13g2_decap_8 FILLER_4_28 ();
 sg13g2_decap_8 FILLER_4_35 ();
 sg13g2_decap_8 FILLER_4_42 ();
 sg13g2_decap_8 FILLER_4_49 ();
 sg13g2_decap_8 FILLER_4_56 ();
 sg13g2_decap_8 FILLER_4_63 ();
 sg13g2_decap_8 FILLER_4_70 ();
 sg13g2_decap_8 FILLER_4_77 ();
 sg13g2_decap_8 FILLER_4_84 ();
 sg13g2_decap_8 FILLER_4_91 ();
 sg13g2_decap_8 FILLER_4_98 ();
 sg13g2_decap_8 FILLER_4_105 ();
 sg13g2_decap_8 FILLER_4_112 ();
 sg13g2_decap_8 FILLER_4_119 ();
 sg13g2_decap_8 FILLER_4_126 ();
 sg13g2_decap_8 FILLER_4_133 ();
 sg13g2_decap_8 FILLER_4_140 ();
 sg13g2_decap_8 FILLER_4_147 ();
 sg13g2_decap_8 FILLER_4_154 ();
 sg13g2_decap_8 FILLER_4_161 ();
 sg13g2_decap_8 FILLER_4_168 ();
 sg13g2_decap_8 FILLER_4_175 ();
 sg13g2_decap_8 FILLER_4_182 ();
 sg13g2_decap_8 FILLER_4_189 ();
 sg13g2_decap_8 FILLER_4_196 ();
 sg13g2_decap_8 FILLER_4_203 ();
 sg13g2_decap_8 FILLER_4_210 ();
 sg13g2_decap_8 FILLER_4_217 ();
 sg13g2_decap_8 FILLER_4_224 ();
 sg13g2_decap_8 FILLER_4_231 ();
 sg13g2_decap_8 FILLER_4_238 ();
 sg13g2_decap_8 FILLER_4_245 ();
 sg13g2_decap_8 FILLER_4_252 ();
 sg13g2_decap_8 FILLER_4_259 ();
 sg13g2_decap_8 FILLER_4_266 ();
 sg13g2_decap_8 FILLER_4_273 ();
 sg13g2_decap_8 FILLER_4_280 ();
 sg13g2_decap_8 FILLER_4_287 ();
 sg13g2_decap_8 FILLER_4_294 ();
 sg13g2_decap_8 FILLER_4_301 ();
 sg13g2_decap_8 FILLER_4_308 ();
 sg13g2_decap_8 FILLER_4_315 ();
 sg13g2_decap_8 FILLER_4_322 ();
 sg13g2_decap_8 FILLER_4_329 ();
 sg13g2_decap_8 FILLER_4_336 ();
 sg13g2_decap_8 FILLER_4_343 ();
 sg13g2_decap_8 FILLER_4_350 ();
 sg13g2_decap_8 FILLER_4_357 ();
 sg13g2_decap_8 FILLER_4_364 ();
 sg13g2_decap_8 FILLER_4_371 ();
 sg13g2_decap_8 FILLER_4_378 ();
 sg13g2_decap_8 FILLER_4_385 ();
 sg13g2_decap_8 FILLER_4_392 ();
 sg13g2_decap_8 FILLER_4_399 ();
 sg13g2_decap_8 FILLER_4_406 ();
 sg13g2_decap_8 FILLER_4_413 ();
 sg13g2_decap_8 FILLER_4_420 ();
 sg13g2_fill_2 FILLER_4_427 ();
 sg13g2_fill_1 FILLER_4_429 ();
 sg13g2_decap_8 FILLER_5_0 ();
 sg13g2_decap_8 FILLER_5_7 ();
 sg13g2_decap_8 FILLER_5_14 ();
 sg13g2_decap_8 FILLER_5_21 ();
 sg13g2_decap_8 FILLER_5_28 ();
 sg13g2_decap_8 FILLER_5_35 ();
 sg13g2_decap_8 FILLER_5_42 ();
 sg13g2_decap_8 FILLER_5_49 ();
 sg13g2_decap_8 FILLER_5_56 ();
 sg13g2_decap_8 FILLER_5_63 ();
 sg13g2_decap_8 FILLER_5_70 ();
 sg13g2_decap_8 FILLER_5_77 ();
 sg13g2_decap_8 FILLER_5_84 ();
 sg13g2_decap_8 FILLER_5_91 ();
 sg13g2_decap_8 FILLER_5_98 ();
 sg13g2_decap_8 FILLER_5_105 ();
 sg13g2_decap_8 FILLER_5_112 ();
 sg13g2_decap_8 FILLER_5_119 ();
 sg13g2_decap_8 FILLER_5_126 ();
 sg13g2_decap_8 FILLER_5_133 ();
 sg13g2_decap_8 FILLER_5_140 ();
 sg13g2_decap_8 FILLER_5_147 ();
 sg13g2_decap_8 FILLER_5_154 ();
 sg13g2_decap_8 FILLER_5_161 ();
 sg13g2_decap_8 FILLER_5_168 ();
 sg13g2_decap_8 FILLER_5_175 ();
 sg13g2_decap_8 FILLER_5_182 ();
 sg13g2_decap_8 FILLER_5_189 ();
 sg13g2_decap_8 FILLER_5_196 ();
 sg13g2_decap_8 FILLER_5_203 ();
 sg13g2_decap_8 FILLER_5_210 ();
 sg13g2_decap_8 FILLER_5_217 ();
 sg13g2_decap_8 FILLER_5_224 ();
 sg13g2_decap_8 FILLER_5_231 ();
 sg13g2_decap_8 FILLER_5_238 ();
 sg13g2_decap_8 FILLER_5_245 ();
 sg13g2_decap_8 FILLER_5_252 ();
 sg13g2_decap_8 FILLER_5_259 ();
 sg13g2_decap_8 FILLER_5_266 ();
 sg13g2_decap_8 FILLER_5_273 ();
 sg13g2_decap_8 FILLER_5_280 ();
 sg13g2_decap_8 FILLER_5_287 ();
 sg13g2_decap_8 FILLER_5_294 ();
 sg13g2_decap_8 FILLER_5_301 ();
 sg13g2_decap_8 FILLER_5_308 ();
 sg13g2_decap_8 FILLER_5_315 ();
 sg13g2_decap_8 FILLER_5_322 ();
 sg13g2_decap_8 FILLER_5_329 ();
 sg13g2_decap_8 FILLER_5_336 ();
 sg13g2_decap_8 FILLER_5_343 ();
 sg13g2_decap_8 FILLER_5_350 ();
 sg13g2_decap_8 FILLER_5_357 ();
 sg13g2_decap_8 FILLER_5_364 ();
 sg13g2_decap_8 FILLER_5_371 ();
 sg13g2_decap_8 FILLER_5_378 ();
 sg13g2_decap_8 FILLER_5_385 ();
 sg13g2_decap_8 FILLER_5_392 ();
 sg13g2_decap_8 FILLER_5_399 ();
 sg13g2_decap_8 FILLER_5_406 ();
 sg13g2_decap_8 FILLER_5_413 ();
 sg13g2_decap_8 FILLER_5_420 ();
 sg13g2_fill_2 FILLER_5_427 ();
 sg13g2_fill_1 FILLER_5_429 ();
 sg13g2_decap_8 FILLER_6_0 ();
 sg13g2_decap_8 FILLER_6_7 ();
 sg13g2_decap_8 FILLER_6_14 ();
 sg13g2_decap_8 FILLER_6_21 ();
 sg13g2_decap_8 FILLER_6_28 ();
 sg13g2_decap_8 FILLER_6_35 ();
 sg13g2_decap_8 FILLER_6_42 ();
 sg13g2_decap_8 FILLER_6_49 ();
 sg13g2_decap_8 FILLER_6_56 ();
 sg13g2_decap_8 FILLER_6_63 ();
 sg13g2_decap_8 FILLER_6_70 ();
 sg13g2_decap_8 FILLER_6_77 ();
 sg13g2_decap_8 FILLER_6_84 ();
 sg13g2_decap_8 FILLER_6_91 ();
 sg13g2_decap_8 FILLER_6_98 ();
 sg13g2_decap_8 FILLER_6_105 ();
 sg13g2_decap_8 FILLER_6_112 ();
 sg13g2_decap_8 FILLER_6_119 ();
 sg13g2_decap_8 FILLER_6_126 ();
 sg13g2_decap_8 FILLER_6_133 ();
 sg13g2_decap_8 FILLER_6_140 ();
 sg13g2_decap_8 FILLER_6_147 ();
 sg13g2_decap_8 FILLER_6_154 ();
 sg13g2_decap_8 FILLER_6_161 ();
 sg13g2_decap_8 FILLER_6_168 ();
 sg13g2_decap_8 FILLER_6_175 ();
 sg13g2_decap_8 FILLER_6_182 ();
 sg13g2_decap_8 FILLER_6_189 ();
 sg13g2_decap_8 FILLER_6_196 ();
 sg13g2_decap_8 FILLER_6_203 ();
 sg13g2_decap_8 FILLER_6_210 ();
 sg13g2_decap_8 FILLER_6_217 ();
 sg13g2_decap_8 FILLER_6_224 ();
 sg13g2_decap_8 FILLER_6_231 ();
 sg13g2_decap_8 FILLER_6_238 ();
 sg13g2_decap_8 FILLER_6_245 ();
 sg13g2_decap_8 FILLER_6_252 ();
 sg13g2_decap_8 FILLER_6_259 ();
 sg13g2_decap_8 FILLER_6_266 ();
 sg13g2_decap_8 FILLER_6_273 ();
 sg13g2_decap_8 FILLER_6_280 ();
 sg13g2_decap_8 FILLER_6_287 ();
 sg13g2_decap_8 FILLER_6_294 ();
 sg13g2_decap_8 FILLER_6_301 ();
 sg13g2_decap_8 FILLER_6_308 ();
 sg13g2_decap_8 FILLER_6_315 ();
 sg13g2_decap_8 FILLER_6_322 ();
 sg13g2_decap_8 FILLER_6_329 ();
 sg13g2_decap_8 FILLER_6_336 ();
 sg13g2_decap_8 FILLER_6_343 ();
 sg13g2_decap_8 FILLER_6_350 ();
 sg13g2_decap_8 FILLER_6_357 ();
 sg13g2_decap_8 FILLER_6_364 ();
 sg13g2_decap_8 FILLER_6_371 ();
 sg13g2_decap_8 FILLER_6_378 ();
 sg13g2_decap_8 FILLER_6_385 ();
 sg13g2_decap_8 FILLER_6_392 ();
 sg13g2_decap_8 FILLER_6_399 ();
 sg13g2_decap_8 FILLER_6_406 ();
 sg13g2_decap_8 FILLER_6_413 ();
 sg13g2_decap_8 FILLER_6_420 ();
 sg13g2_fill_2 FILLER_6_427 ();
 sg13g2_fill_1 FILLER_6_429 ();
 sg13g2_decap_8 FILLER_7_0 ();
 sg13g2_decap_8 FILLER_7_7 ();
 sg13g2_decap_8 FILLER_7_14 ();
 sg13g2_decap_8 FILLER_7_21 ();
 sg13g2_decap_8 FILLER_7_28 ();
 sg13g2_decap_8 FILLER_7_35 ();
 sg13g2_decap_8 FILLER_7_42 ();
 sg13g2_decap_8 FILLER_7_49 ();
 sg13g2_decap_8 FILLER_7_56 ();
 sg13g2_decap_8 FILLER_7_63 ();
 sg13g2_decap_8 FILLER_7_70 ();
 sg13g2_decap_8 FILLER_7_77 ();
 sg13g2_decap_8 FILLER_7_84 ();
 sg13g2_decap_8 FILLER_7_91 ();
 sg13g2_decap_8 FILLER_7_98 ();
 sg13g2_decap_8 FILLER_7_105 ();
 sg13g2_decap_8 FILLER_7_112 ();
 sg13g2_decap_8 FILLER_7_119 ();
 sg13g2_decap_8 FILLER_7_126 ();
 sg13g2_decap_8 FILLER_7_133 ();
 sg13g2_decap_8 FILLER_7_140 ();
 sg13g2_decap_8 FILLER_7_147 ();
 sg13g2_decap_8 FILLER_7_154 ();
 sg13g2_decap_8 FILLER_7_161 ();
 sg13g2_decap_8 FILLER_7_168 ();
 sg13g2_decap_8 FILLER_7_175 ();
 sg13g2_decap_8 FILLER_7_182 ();
 sg13g2_decap_8 FILLER_7_189 ();
 sg13g2_decap_8 FILLER_7_196 ();
 sg13g2_decap_8 FILLER_7_203 ();
 sg13g2_decap_8 FILLER_7_210 ();
 sg13g2_decap_8 FILLER_7_217 ();
 sg13g2_decap_8 FILLER_7_224 ();
 sg13g2_decap_8 FILLER_7_231 ();
 sg13g2_decap_8 FILLER_7_238 ();
 sg13g2_decap_8 FILLER_7_245 ();
 sg13g2_decap_8 FILLER_7_252 ();
 sg13g2_decap_8 FILLER_7_259 ();
 sg13g2_decap_8 FILLER_7_266 ();
 sg13g2_decap_8 FILLER_7_273 ();
 sg13g2_decap_8 FILLER_7_280 ();
 sg13g2_decap_8 FILLER_7_287 ();
 sg13g2_decap_8 FILLER_7_294 ();
 sg13g2_decap_8 FILLER_7_301 ();
 sg13g2_decap_8 FILLER_7_308 ();
 sg13g2_decap_8 FILLER_7_315 ();
 sg13g2_decap_8 FILLER_7_322 ();
 sg13g2_decap_8 FILLER_7_329 ();
 sg13g2_decap_8 FILLER_7_336 ();
 sg13g2_decap_8 FILLER_7_343 ();
 sg13g2_decap_8 FILLER_7_350 ();
 sg13g2_decap_8 FILLER_7_357 ();
 sg13g2_decap_8 FILLER_7_364 ();
 sg13g2_decap_8 FILLER_7_371 ();
 sg13g2_decap_8 FILLER_7_378 ();
 sg13g2_decap_8 FILLER_7_385 ();
 sg13g2_decap_8 FILLER_7_392 ();
 sg13g2_decap_8 FILLER_7_399 ();
 sg13g2_decap_8 FILLER_7_406 ();
 sg13g2_decap_8 FILLER_7_413 ();
 sg13g2_decap_8 FILLER_7_420 ();
 sg13g2_fill_2 FILLER_7_427 ();
 sg13g2_fill_1 FILLER_7_429 ();
 sg13g2_decap_8 FILLER_8_0 ();
 sg13g2_decap_8 FILLER_8_7 ();
 sg13g2_decap_8 FILLER_8_14 ();
 sg13g2_decap_8 FILLER_8_21 ();
 sg13g2_decap_8 FILLER_8_28 ();
 sg13g2_decap_8 FILLER_8_35 ();
 sg13g2_decap_8 FILLER_8_42 ();
 sg13g2_decap_8 FILLER_8_49 ();
 sg13g2_decap_8 FILLER_8_56 ();
 sg13g2_decap_8 FILLER_8_63 ();
 sg13g2_decap_8 FILLER_8_70 ();
 sg13g2_decap_8 FILLER_8_77 ();
 sg13g2_decap_8 FILLER_8_84 ();
 sg13g2_decap_8 FILLER_8_91 ();
 sg13g2_decap_8 FILLER_8_98 ();
 sg13g2_decap_8 FILLER_8_105 ();
 sg13g2_decap_8 FILLER_8_112 ();
 sg13g2_decap_8 FILLER_8_119 ();
 sg13g2_decap_8 FILLER_8_126 ();
 sg13g2_decap_8 FILLER_8_133 ();
 sg13g2_decap_8 FILLER_8_140 ();
 sg13g2_decap_8 FILLER_8_147 ();
 sg13g2_decap_8 FILLER_8_154 ();
 sg13g2_decap_8 FILLER_8_161 ();
 sg13g2_decap_8 FILLER_8_168 ();
 sg13g2_decap_8 FILLER_8_175 ();
 sg13g2_decap_8 FILLER_8_182 ();
 sg13g2_decap_8 FILLER_8_189 ();
 sg13g2_decap_8 FILLER_8_196 ();
 sg13g2_decap_8 FILLER_8_203 ();
 sg13g2_decap_8 FILLER_8_210 ();
 sg13g2_decap_8 FILLER_8_217 ();
 sg13g2_decap_8 FILLER_8_224 ();
 sg13g2_decap_8 FILLER_8_231 ();
 sg13g2_decap_8 FILLER_8_238 ();
 sg13g2_decap_8 FILLER_8_245 ();
 sg13g2_decap_8 FILLER_8_252 ();
 sg13g2_decap_8 FILLER_8_259 ();
 sg13g2_decap_8 FILLER_8_266 ();
 sg13g2_decap_8 FILLER_8_273 ();
 sg13g2_decap_8 FILLER_8_280 ();
 sg13g2_decap_8 FILLER_8_287 ();
 sg13g2_decap_8 FILLER_8_294 ();
 sg13g2_decap_8 FILLER_8_301 ();
 sg13g2_decap_8 FILLER_8_308 ();
 sg13g2_decap_8 FILLER_8_315 ();
 sg13g2_decap_8 FILLER_8_322 ();
 sg13g2_decap_8 FILLER_8_329 ();
 sg13g2_decap_8 FILLER_8_336 ();
 sg13g2_decap_8 FILLER_8_343 ();
 sg13g2_decap_8 FILLER_8_350 ();
 sg13g2_decap_8 FILLER_8_357 ();
 sg13g2_decap_8 FILLER_8_364 ();
 sg13g2_decap_8 FILLER_8_371 ();
 sg13g2_decap_8 FILLER_8_378 ();
 sg13g2_decap_8 FILLER_8_385 ();
 sg13g2_decap_8 FILLER_8_392 ();
 sg13g2_decap_8 FILLER_8_399 ();
 sg13g2_decap_8 FILLER_8_406 ();
 sg13g2_decap_8 FILLER_8_413 ();
 sg13g2_decap_8 FILLER_8_420 ();
 sg13g2_fill_2 FILLER_8_427 ();
 sg13g2_fill_1 FILLER_8_429 ();
 sg13g2_decap_8 FILLER_9_0 ();
 sg13g2_decap_8 FILLER_9_7 ();
 sg13g2_decap_8 FILLER_9_14 ();
 sg13g2_decap_8 FILLER_9_21 ();
 sg13g2_decap_8 FILLER_9_28 ();
 sg13g2_decap_8 FILLER_9_35 ();
 sg13g2_decap_8 FILLER_9_42 ();
 sg13g2_decap_8 FILLER_9_49 ();
 sg13g2_decap_8 FILLER_9_56 ();
 sg13g2_decap_8 FILLER_9_63 ();
 sg13g2_decap_8 FILLER_9_70 ();
 sg13g2_decap_8 FILLER_9_77 ();
 sg13g2_decap_8 FILLER_9_84 ();
 sg13g2_decap_8 FILLER_9_91 ();
 sg13g2_decap_8 FILLER_9_98 ();
 sg13g2_decap_8 FILLER_9_105 ();
 sg13g2_decap_8 FILLER_9_112 ();
 sg13g2_decap_8 FILLER_9_119 ();
 sg13g2_decap_8 FILLER_9_126 ();
 sg13g2_decap_8 FILLER_9_133 ();
 sg13g2_decap_8 FILLER_9_140 ();
 sg13g2_decap_8 FILLER_9_147 ();
 sg13g2_decap_8 FILLER_9_154 ();
 sg13g2_decap_8 FILLER_9_161 ();
 sg13g2_decap_8 FILLER_9_168 ();
 sg13g2_decap_8 FILLER_9_175 ();
 sg13g2_decap_8 FILLER_9_182 ();
 sg13g2_decap_8 FILLER_9_189 ();
 sg13g2_decap_8 FILLER_9_196 ();
 sg13g2_decap_8 FILLER_9_203 ();
 sg13g2_decap_8 FILLER_9_210 ();
 sg13g2_decap_8 FILLER_9_217 ();
 sg13g2_decap_8 FILLER_9_224 ();
 sg13g2_decap_8 FILLER_9_231 ();
 sg13g2_decap_8 FILLER_9_238 ();
 sg13g2_decap_8 FILLER_9_245 ();
 sg13g2_decap_8 FILLER_9_252 ();
 sg13g2_decap_8 FILLER_9_259 ();
 sg13g2_decap_8 FILLER_9_266 ();
 sg13g2_decap_8 FILLER_9_273 ();
 sg13g2_decap_8 FILLER_9_280 ();
 sg13g2_decap_8 FILLER_9_287 ();
 sg13g2_decap_8 FILLER_9_294 ();
 sg13g2_decap_8 FILLER_9_301 ();
 sg13g2_decap_8 FILLER_9_308 ();
 sg13g2_decap_8 FILLER_9_315 ();
 sg13g2_decap_8 FILLER_9_322 ();
 sg13g2_decap_8 FILLER_9_329 ();
 sg13g2_decap_8 FILLER_9_336 ();
 sg13g2_decap_8 FILLER_9_343 ();
 sg13g2_decap_8 FILLER_9_350 ();
 sg13g2_decap_8 FILLER_9_357 ();
 sg13g2_decap_8 FILLER_9_364 ();
 sg13g2_decap_8 FILLER_9_371 ();
 sg13g2_decap_8 FILLER_9_378 ();
 sg13g2_decap_8 FILLER_9_385 ();
 sg13g2_decap_8 FILLER_9_392 ();
 sg13g2_decap_8 FILLER_9_399 ();
 sg13g2_decap_8 FILLER_9_406 ();
 sg13g2_decap_8 FILLER_9_413 ();
 sg13g2_decap_8 FILLER_9_420 ();
 sg13g2_fill_2 FILLER_9_427 ();
 sg13g2_fill_1 FILLER_9_429 ();
 sg13g2_decap_8 FILLER_10_0 ();
 sg13g2_decap_8 FILLER_10_7 ();
 sg13g2_decap_8 FILLER_10_14 ();
 sg13g2_decap_8 FILLER_10_21 ();
 sg13g2_decap_8 FILLER_10_28 ();
 sg13g2_decap_8 FILLER_10_35 ();
 sg13g2_decap_8 FILLER_10_42 ();
 sg13g2_decap_8 FILLER_10_49 ();
 sg13g2_decap_8 FILLER_10_56 ();
 sg13g2_decap_8 FILLER_10_63 ();
 sg13g2_decap_8 FILLER_10_70 ();
 sg13g2_decap_8 FILLER_10_77 ();
 sg13g2_decap_8 FILLER_10_84 ();
 sg13g2_decap_8 FILLER_10_91 ();
 sg13g2_decap_8 FILLER_10_98 ();
 sg13g2_decap_8 FILLER_10_105 ();
 sg13g2_decap_8 FILLER_10_112 ();
 sg13g2_decap_8 FILLER_10_119 ();
 sg13g2_decap_8 FILLER_10_126 ();
 sg13g2_decap_8 FILLER_10_133 ();
 sg13g2_decap_8 FILLER_10_140 ();
 sg13g2_decap_8 FILLER_10_147 ();
 sg13g2_decap_8 FILLER_10_154 ();
 sg13g2_decap_8 FILLER_10_161 ();
 sg13g2_decap_8 FILLER_10_168 ();
 sg13g2_decap_8 FILLER_10_175 ();
 sg13g2_decap_8 FILLER_10_182 ();
 sg13g2_decap_8 FILLER_10_189 ();
 sg13g2_decap_8 FILLER_10_196 ();
 sg13g2_decap_8 FILLER_10_203 ();
 sg13g2_decap_8 FILLER_10_210 ();
 sg13g2_decap_8 FILLER_10_217 ();
 sg13g2_decap_8 FILLER_10_224 ();
 sg13g2_decap_8 FILLER_10_231 ();
 sg13g2_decap_8 FILLER_10_238 ();
 sg13g2_decap_8 FILLER_10_245 ();
 sg13g2_decap_8 FILLER_10_252 ();
 sg13g2_decap_8 FILLER_10_259 ();
 sg13g2_decap_8 FILLER_10_266 ();
 sg13g2_decap_8 FILLER_10_273 ();
 sg13g2_decap_8 FILLER_10_280 ();
 sg13g2_decap_8 FILLER_10_287 ();
 sg13g2_decap_8 FILLER_10_294 ();
 sg13g2_decap_8 FILLER_10_301 ();
 sg13g2_decap_8 FILLER_10_308 ();
 sg13g2_decap_8 FILLER_10_315 ();
 sg13g2_decap_8 FILLER_10_322 ();
 sg13g2_decap_8 FILLER_10_329 ();
 sg13g2_decap_8 FILLER_10_336 ();
 sg13g2_decap_8 FILLER_10_343 ();
 sg13g2_decap_8 FILLER_10_350 ();
 sg13g2_decap_8 FILLER_10_357 ();
 sg13g2_decap_8 FILLER_10_364 ();
 sg13g2_decap_8 FILLER_10_371 ();
 sg13g2_decap_8 FILLER_10_378 ();
 sg13g2_decap_8 FILLER_10_385 ();
 sg13g2_decap_8 FILLER_10_392 ();
 sg13g2_decap_8 FILLER_10_399 ();
 sg13g2_decap_8 FILLER_10_406 ();
 sg13g2_decap_8 FILLER_10_413 ();
 sg13g2_decap_8 FILLER_10_420 ();
 sg13g2_fill_2 FILLER_10_427 ();
 sg13g2_fill_1 FILLER_10_429 ();
 sg13g2_decap_8 FILLER_11_0 ();
 sg13g2_decap_8 FILLER_11_7 ();
 sg13g2_decap_8 FILLER_11_14 ();
 sg13g2_decap_8 FILLER_11_21 ();
 sg13g2_decap_8 FILLER_11_28 ();
 sg13g2_decap_8 FILLER_11_35 ();
 sg13g2_decap_8 FILLER_11_42 ();
 sg13g2_decap_8 FILLER_11_49 ();
 sg13g2_decap_8 FILLER_11_56 ();
 sg13g2_decap_8 FILLER_11_63 ();
 sg13g2_decap_8 FILLER_11_70 ();
 sg13g2_decap_8 FILLER_11_77 ();
 sg13g2_decap_8 FILLER_11_84 ();
 sg13g2_decap_8 FILLER_11_91 ();
 sg13g2_decap_8 FILLER_11_98 ();
 sg13g2_decap_8 FILLER_11_105 ();
 sg13g2_decap_8 FILLER_11_112 ();
 sg13g2_decap_8 FILLER_11_119 ();
 sg13g2_decap_8 FILLER_11_126 ();
 sg13g2_decap_8 FILLER_11_133 ();
 sg13g2_decap_8 FILLER_11_140 ();
 sg13g2_decap_8 FILLER_11_147 ();
 sg13g2_decap_8 FILLER_11_154 ();
 sg13g2_decap_8 FILLER_11_161 ();
 sg13g2_decap_8 FILLER_11_168 ();
 sg13g2_decap_8 FILLER_11_175 ();
 sg13g2_decap_8 FILLER_11_182 ();
 sg13g2_decap_8 FILLER_11_189 ();
 sg13g2_decap_8 FILLER_11_196 ();
 sg13g2_decap_8 FILLER_11_203 ();
 sg13g2_decap_8 FILLER_11_210 ();
 sg13g2_decap_8 FILLER_11_217 ();
 sg13g2_decap_8 FILLER_11_224 ();
 sg13g2_decap_8 FILLER_11_231 ();
 sg13g2_decap_8 FILLER_11_238 ();
 sg13g2_decap_8 FILLER_11_245 ();
 sg13g2_decap_8 FILLER_11_252 ();
 sg13g2_decap_8 FILLER_11_259 ();
 sg13g2_decap_8 FILLER_11_266 ();
 sg13g2_decap_8 FILLER_11_273 ();
 sg13g2_decap_8 FILLER_11_280 ();
 sg13g2_decap_8 FILLER_11_287 ();
 sg13g2_decap_8 FILLER_11_294 ();
 sg13g2_decap_8 FILLER_11_301 ();
 sg13g2_decap_8 FILLER_11_308 ();
 sg13g2_decap_8 FILLER_11_315 ();
 sg13g2_decap_8 FILLER_11_322 ();
 sg13g2_decap_8 FILLER_11_329 ();
 sg13g2_decap_8 FILLER_11_336 ();
 sg13g2_decap_8 FILLER_11_343 ();
 sg13g2_decap_8 FILLER_11_350 ();
 sg13g2_decap_8 FILLER_11_357 ();
 sg13g2_decap_8 FILLER_11_364 ();
 sg13g2_decap_8 FILLER_11_371 ();
 sg13g2_decap_8 FILLER_11_378 ();
 sg13g2_decap_8 FILLER_11_385 ();
 sg13g2_decap_8 FILLER_11_392 ();
 sg13g2_decap_8 FILLER_11_399 ();
 sg13g2_decap_8 FILLER_11_406 ();
 sg13g2_decap_8 FILLER_11_413 ();
 sg13g2_decap_8 FILLER_11_420 ();
 sg13g2_fill_2 FILLER_11_427 ();
 sg13g2_fill_1 FILLER_11_429 ();
 sg13g2_decap_8 FILLER_12_0 ();
 sg13g2_decap_8 FILLER_12_7 ();
 sg13g2_decap_8 FILLER_12_14 ();
 sg13g2_decap_8 FILLER_12_21 ();
 sg13g2_decap_8 FILLER_12_28 ();
 sg13g2_decap_8 FILLER_12_35 ();
 sg13g2_decap_8 FILLER_12_42 ();
 sg13g2_decap_8 FILLER_12_49 ();
 sg13g2_decap_8 FILLER_12_56 ();
 sg13g2_decap_8 FILLER_12_63 ();
 sg13g2_decap_8 FILLER_12_70 ();
 sg13g2_decap_8 FILLER_12_77 ();
 sg13g2_decap_8 FILLER_12_84 ();
 sg13g2_decap_8 FILLER_12_91 ();
 sg13g2_decap_8 FILLER_12_98 ();
 sg13g2_decap_8 FILLER_12_105 ();
 sg13g2_decap_8 FILLER_12_112 ();
 sg13g2_decap_8 FILLER_12_119 ();
 sg13g2_decap_8 FILLER_12_126 ();
 sg13g2_decap_8 FILLER_12_133 ();
 sg13g2_decap_8 FILLER_12_140 ();
 sg13g2_decap_8 FILLER_12_147 ();
 sg13g2_decap_8 FILLER_12_154 ();
 sg13g2_decap_8 FILLER_12_161 ();
 sg13g2_decap_8 FILLER_12_168 ();
 sg13g2_decap_8 FILLER_12_175 ();
 sg13g2_decap_8 FILLER_12_182 ();
 sg13g2_decap_8 FILLER_12_189 ();
 sg13g2_decap_8 FILLER_12_196 ();
 sg13g2_decap_8 FILLER_12_203 ();
 sg13g2_decap_8 FILLER_12_210 ();
 sg13g2_decap_8 FILLER_12_217 ();
 sg13g2_decap_8 FILLER_12_224 ();
 sg13g2_decap_8 FILLER_12_231 ();
 sg13g2_decap_8 FILLER_12_238 ();
 sg13g2_decap_8 FILLER_12_245 ();
 sg13g2_decap_8 FILLER_12_252 ();
 sg13g2_decap_8 FILLER_12_259 ();
 sg13g2_decap_8 FILLER_12_266 ();
 sg13g2_decap_8 FILLER_12_281 ();
 sg13g2_fill_1 FILLER_12_288 ();
 sg13g2_decap_8 FILLER_12_297 ();
 sg13g2_fill_1 FILLER_12_304 ();
 sg13g2_decap_4 FILLER_12_309 ();
 sg13g2_decap_8 FILLER_12_323 ();
 sg13g2_fill_2 FILLER_12_330 ();
 sg13g2_decap_8 FILLER_12_336 ();
 sg13g2_decap_8 FILLER_12_343 ();
 sg13g2_fill_2 FILLER_12_350 ();
 sg13g2_fill_1 FILLER_12_352 ();
 sg13g2_decap_4 FILLER_12_361 ();
 sg13g2_fill_1 FILLER_12_378 ();
 sg13g2_decap_8 FILLER_12_387 ();
 sg13g2_decap_8 FILLER_12_394 ();
 sg13g2_decap_8 FILLER_12_401 ();
 sg13g2_decap_8 FILLER_12_408 ();
 sg13g2_decap_8 FILLER_12_415 ();
 sg13g2_decap_8 FILLER_12_422 ();
 sg13g2_fill_1 FILLER_12_429 ();
 sg13g2_decap_8 FILLER_13_0 ();
 sg13g2_decap_8 FILLER_13_7 ();
 sg13g2_decap_8 FILLER_13_14 ();
 sg13g2_decap_8 FILLER_13_21 ();
 sg13g2_decap_8 FILLER_13_28 ();
 sg13g2_decap_8 FILLER_13_35 ();
 sg13g2_decap_8 FILLER_13_42 ();
 sg13g2_decap_8 FILLER_13_49 ();
 sg13g2_decap_8 FILLER_13_56 ();
 sg13g2_decap_8 FILLER_13_63 ();
 sg13g2_decap_8 FILLER_13_70 ();
 sg13g2_decap_8 FILLER_13_77 ();
 sg13g2_decap_8 FILLER_13_84 ();
 sg13g2_decap_8 FILLER_13_91 ();
 sg13g2_decap_8 FILLER_13_98 ();
 sg13g2_decap_8 FILLER_13_105 ();
 sg13g2_decap_8 FILLER_13_112 ();
 sg13g2_decap_4 FILLER_13_119 ();
 sg13g2_fill_1 FILLER_13_123 ();
 sg13g2_decap_8 FILLER_13_128 ();
 sg13g2_decap_8 FILLER_13_135 ();
 sg13g2_decap_8 FILLER_13_142 ();
 sg13g2_decap_8 FILLER_13_149 ();
 sg13g2_decap_8 FILLER_13_156 ();
 sg13g2_decap_8 FILLER_13_163 ();
 sg13g2_decap_8 FILLER_13_170 ();
 sg13g2_decap_8 FILLER_13_177 ();
 sg13g2_fill_2 FILLER_13_184 ();
 sg13g2_decap_8 FILLER_13_190 ();
 sg13g2_decap_4 FILLER_13_202 ();
 sg13g2_fill_2 FILLER_13_206 ();
 sg13g2_decap_4 FILLER_13_262 ();
 sg13g2_fill_2 FILLER_13_273 ();
 sg13g2_fill_1 FILLER_13_275 ();
 sg13g2_fill_2 FILLER_13_291 ();
 sg13g2_fill_1 FILLER_13_297 ();
 sg13g2_fill_1 FILLER_13_325 ();
 sg13g2_fill_2 FILLER_13_331 ();
 sg13g2_fill_2 FILLER_13_338 ();
 sg13g2_fill_2 FILLER_13_348 ();
 sg13g2_fill_1 FILLER_13_350 ();
 sg13g2_fill_1 FILLER_13_376 ();
 sg13g2_decap_8 FILLER_13_389 ();
 sg13g2_decap_8 FILLER_13_396 ();
 sg13g2_decap_8 FILLER_13_403 ();
 sg13g2_decap_8 FILLER_13_410 ();
 sg13g2_decap_8 FILLER_13_417 ();
 sg13g2_decap_4 FILLER_13_424 ();
 sg13g2_fill_2 FILLER_13_428 ();
 sg13g2_decap_8 FILLER_14_0 ();
 sg13g2_decap_8 FILLER_14_7 ();
 sg13g2_decap_8 FILLER_14_14 ();
 sg13g2_decap_8 FILLER_14_21 ();
 sg13g2_decap_8 FILLER_14_28 ();
 sg13g2_decap_8 FILLER_14_35 ();
 sg13g2_decap_8 FILLER_14_42 ();
 sg13g2_decap_8 FILLER_14_49 ();
 sg13g2_decap_8 FILLER_14_56 ();
 sg13g2_decap_8 FILLER_14_63 ();
 sg13g2_decap_8 FILLER_14_70 ();
 sg13g2_decap_8 FILLER_14_77 ();
 sg13g2_fill_1 FILLER_14_84 ();
 sg13g2_fill_2 FILLER_14_93 ();
 sg13g2_decap_4 FILLER_14_112 ();
 sg13g2_fill_2 FILLER_14_116 ();
 sg13g2_fill_1 FILLER_14_123 ();
 sg13g2_fill_1 FILLER_14_128 ();
 sg13g2_fill_2 FILLER_14_153 ();
 sg13g2_fill_1 FILLER_14_155 ();
 sg13g2_fill_2 FILLER_14_160 ();
 sg13g2_fill_1 FILLER_14_162 ();
 sg13g2_decap_8 FILLER_14_176 ();
 sg13g2_decap_8 FILLER_14_183 ();
 sg13g2_decap_8 FILLER_14_190 ();
 sg13g2_decap_4 FILLER_14_197 ();
 sg13g2_fill_1 FILLER_14_206 ();
 sg13g2_fill_2 FILLER_14_216 ();
 sg13g2_fill_2 FILLER_14_225 ();
 sg13g2_fill_1 FILLER_14_227 ();
 sg13g2_fill_1 FILLER_14_233 ();
 sg13g2_fill_2 FILLER_14_259 ();
 sg13g2_fill_1 FILLER_14_261 ();
 sg13g2_fill_1 FILLER_14_266 ();
 sg13g2_decap_8 FILLER_14_284 ();
 sg13g2_decap_8 FILLER_14_291 ();
 sg13g2_decap_8 FILLER_14_298 ();
 sg13g2_decap_8 FILLER_14_305 ();
 sg13g2_decap_8 FILLER_14_316 ();
 sg13g2_decap_8 FILLER_14_323 ();
 sg13g2_fill_1 FILLER_14_330 ();
 sg13g2_decap_8 FILLER_14_347 ();
 sg13g2_decap_8 FILLER_14_354 ();
 sg13g2_fill_1 FILLER_14_361 ();
 sg13g2_decap_4 FILLER_14_374 ();
 sg13g2_fill_1 FILLER_14_378 ();
 sg13g2_decap_8 FILLER_14_395 ();
 sg13g2_decap_8 FILLER_14_402 ();
 sg13g2_decap_8 FILLER_14_409 ();
 sg13g2_decap_8 FILLER_14_416 ();
 sg13g2_decap_8 FILLER_14_423 ();
 sg13g2_decap_8 FILLER_15_0 ();
 sg13g2_decap_8 FILLER_15_7 ();
 sg13g2_decap_8 FILLER_15_14 ();
 sg13g2_decap_8 FILLER_15_21 ();
 sg13g2_decap_8 FILLER_15_28 ();
 sg13g2_decap_8 FILLER_15_35 ();
 sg13g2_decap_8 FILLER_15_42 ();
 sg13g2_decap_8 FILLER_15_49 ();
 sg13g2_decap_8 FILLER_15_56 ();
 sg13g2_decap_8 FILLER_15_63 ();
 sg13g2_decap_4 FILLER_15_70 ();
 sg13g2_fill_2 FILLER_15_82 ();
 sg13g2_fill_1 FILLER_15_84 ();
 sg13g2_fill_2 FILLER_15_97 ();
 sg13g2_decap_8 FILLER_15_108 ();
 sg13g2_fill_1 FILLER_15_115 ();
 sg13g2_fill_1 FILLER_15_128 ();
 sg13g2_fill_1 FILLER_15_137 ();
 sg13g2_decap_8 FILLER_15_143 ();
 sg13g2_fill_1 FILLER_15_150 ();
 sg13g2_decap_4 FILLER_15_164 ();
 sg13g2_fill_2 FILLER_15_168 ();
 sg13g2_fill_2 FILLER_15_178 ();
 sg13g2_fill_1 FILLER_15_189 ();
 sg13g2_fill_1 FILLER_15_201 ();
 sg13g2_fill_2 FILLER_15_211 ();
 sg13g2_decap_4 FILLER_15_217 ();
 sg13g2_decap_4 FILLER_15_231 ();
 sg13g2_fill_1 FILLER_15_235 ();
 sg13g2_decap_8 FILLER_15_241 ();
 sg13g2_decap_4 FILLER_15_248 ();
 sg13g2_decap_4 FILLER_15_258 ();
 sg13g2_decap_8 FILLER_15_266 ();
 sg13g2_decap_8 FILLER_15_273 ();
 sg13g2_decap_4 FILLER_15_280 ();
 sg13g2_fill_1 FILLER_15_284 ();
 sg13g2_fill_2 FILLER_15_316 ();
 sg13g2_decap_8 FILLER_15_325 ();
 sg13g2_fill_1 FILLER_15_332 ();
 sg13g2_decap_8 FILLER_15_346 ();
 sg13g2_fill_2 FILLER_15_353 ();
 sg13g2_fill_1 FILLER_15_355 ();
 sg13g2_decap_8 FILLER_15_372 ();
 sg13g2_decap_4 FILLER_15_379 ();
 sg13g2_decap_8 FILLER_15_395 ();
 sg13g2_decap_4 FILLER_15_402 ();
 sg13g2_fill_1 FILLER_15_406 ();
 sg13g2_decap_8 FILLER_15_415 ();
 sg13g2_decap_8 FILLER_15_422 ();
 sg13g2_fill_1 FILLER_15_429 ();
 sg13g2_decap_8 FILLER_16_0 ();
 sg13g2_decap_8 FILLER_16_7 ();
 sg13g2_decap_8 FILLER_16_14 ();
 sg13g2_decap_8 FILLER_16_21 ();
 sg13g2_decap_8 FILLER_16_28 ();
 sg13g2_decap_8 FILLER_16_35 ();
 sg13g2_decap_4 FILLER_16_42 ();
 sg13g2_fill_1 FILLER_16_46 ();
 sg13g2_decap_8 FILLER_16_51 ();
 sg13g2_fill_2 FILLER_16_58 ();
 sg13g2_decap_4 FILLER_16_81 ();
 sg13g2_fill_2 FILLER_16_85 ();
 sg13g2_fill_2 FILLER_16_95 ();
 sg13g2_fill_1 FILLER_16_102 ();
 sg13g2_decap_4 FILLER_16_112 ();
 sg13g2_decap_8 FILLER_16_124 ();
 sg13g2_fill_2 FILLER_16_135 ();
 sg13g2_fill_1 FILLER_16_137 ();
 sg13g2_fill_2 FILLER_16_146 ();
 sg13g2_decap_8 FILLER_16_152 ();
 sg13g2_decap_8 FILLER_16_159 ();
 sg13g2_decap_8 FILLER_16_166 ();
 sg13g2_fill_1 FILLER_16_183 ();
 sg13g2_fill_1 FILLER_16_208 ();
 sg13g2_decap_8 FILLER_16_217 ();
 sg13g2_decap_8 FILLER_16_224 ();
 sg13g2_decap_8 FILLER_16_231 ();
 sg13g2_decap_4 FILLER_16_238 ();
 sg13g2_fill_2 FILLER_16_242 ();
 sg13g2_fill_1 FILLER_16_259 ();
 sg13g2_decap_8 FILLER_16_268 ();
 sg13g2_fill_2 FILLER_16_275 ();
 sg13g2_fill_1 FILLER_16_277 ();
 sg13g2_fill_2 FILLER_16_286 ();
 sg13g2_decap_4 FILLER_16_300 ();
 sg13g2_fill_2 FILLER_16_325 ();
 sg13g2_decap_8 FILLER_16_335 ();
 sg13g2_decap_8 FILLER_16_342 ();
 sg13g2_fill_1 FILLER_16_349 ();
 sg13g2_decap_8 FILLER_16_366 ();
 sg13g2_fill_2 FILLER_16_373 ();
 sg13g2_fill_1 FILLER_16_390 ();
 sg13g2_decap_4 FILLER_16_399 ();
 sg13g2_fill_1 FILLER_16_403 ();
 sg13g2_fill_2 FILLER_16_412 ();
 sg13g2_decap_8 FILLER_16_421 ();
 sg13g2_fill_2 FILLER_16_428 ();
 sg13g2_decap_8 FILLER_17_0 ();
 sg13g2_fill_2 FILLER_17_7 ();
 sg13g2_fill_1 FILLER_17_9 ();
 sg13g2_decap_8 FILLER_17_23 ();
 sg13g2_decap_8 FILLER_17_30 ();
 sg13g2_decap_8 FILLER_17_37 ();
 sg13g2_fill_2 FILLER_17_44 ();
 sg13g2_fill_1 FILLER_17_55 ();
 sg13g2_decap_8 FILLER_17_72 ();
 sg13g2_fill_2 FILLER_17_79 ();
 sg13g2_decap_8 FILLER_17_108 ();
 sg13g2_decap_8 FILLER_17_115 ();
 sg13g2_decap_8 FILLER_17_122 ();
 sg13g2_fill_2 FILLER_17_129 ();
 sg13g2_fill_1 FILLER_17_152 ();
 sg13g2_decap_4 FILLER_17_158 ();
 sg13g2_fill_1 FILLER_17_171 ();
 sg13g2_fill_2 FILLER_17_177 ();
 sg13g2_fill_1 FILLER_17_179 ();
 sg13g2_fill_1 FILLER_17_190 ();
 sg13g2_fill_1 FILLER_17_217 ();
 sg13g2_decap_8 FILLER_17_222 ();
 sg13g2_decap_4 FILLER_17_229 ();
 sg13g2_fill_1 FILLER_17_243 ();
 sg13g2_fill_1 FILLER_17_266 ();
 sg13g2_fill_1 FILLER_17_302 ();
 sg13g2_decap_8 FILLER_17_311 ();
 sg13g2_fill_1 FILLER_17_318 ();
 sg13g2_decap_8 FILLER_17_323 ();
 sg13g2_decap_4 FILLER_17_330 ();
 sg13g2_fill_2 FILLER_17_334 ();
 sg13g2_fill_2 FILLER_17_340 ();
 sg13g2_fill_1 FILLER_17_342 ();
 sg13g2_decap_8 FILLER_17_351 ();
 sg13g2_decap_8 FILLER_17_358 ();
 sg13g2_decap_8 FILLER_17_365 ();
 sg13g2_fill_2 FILLER_17_372 ();
 sg13g2_decap_4 FILLER_17_387 ();
 sg13g2_fill_2 FILLER_17_391 ();
 sg13g2_decap_4 FILLER_17_425 ();
 sg13g2_fill_1 FILLER_17_429 ();
 sg13g2_decap_4 FILLER_18_0 ();
 sg13g2_fill_1 FILLER_18_4 ();
 sg13g2_decap_4 FILLER_18_26 ();
 sg13g2_fill_2 FILLER_18_34 ();
 sg13g2_fill_1 FILLER_18_36 ();
 sg13g2_decap_4 FILLER_18_42 ();
 sg13g2_decap_8 FILLER_18_54 ();
 sg13g2_decap_8 FILLER_18_61 ();
 sg13g2_fill_2 FILLER_18_68 ();
 sg13g2_fill_2 FILLER_18_78 ();
 sg13g2_fill_1 FILLER_18_80 ();
 sg13g2_fill_1 FILLER_18_98 ();
 sg13g2_decap_8 FILLER_18_120 ();
 sg13g2_decap_8 FILLER_18_127 ();
 sg13g2_decap_8 FILLER_18_134 ();
 sg13g2_fill_2 FILLER_18_156 ();
 sg13g2_fill_2 FILLER_18_183 ();
 sg13g2_fill_1 FILLER_18_185 ();
 sg13g2_decap_8 FILLER_18_191 ();
 sg13g2_fill_1 FILLER_18_198 ();
 sg13g2_decap_8 FILLER_18_202 ();
 sg13g2_decap_8 FILLER_18_209 ();
 sg13g2_decap_8 FILLER_18_216 ();
 sg13g2_decap_4 FILLER_18_223 ();
 sg13g2_fill_1 FILLER_18_227 ();
 sg13g2_decap_8 FILLER_18_265 ();
 sg13g2_decap_4 FILLER_18_272 ();
 sg13g2_fill_2 FILLER_18_276 ();
 sg13g2_fill_2 FILLER_18_286 ();
 sg13g2_decap_8 FILLER_18_292 ();
 sg13g2_fill_2 FILLER_18_299 ();
 sg13g2_fill_1 FILLER_18_301 ();
 sg13g2_fill_2 FILLER_18_330 ();
 sg13g2_fill_1 FILLER_18_332 ();
 sg13g2_decap_8 FILLER_18_338 ();
 sg13g2_fill_2 FILLER_18_345 ();
 sg13g2_decap_4 FILLER_18_351 ();
 sg13g2_decap_4 FILLER_18_369 ();
 sg13g2_fill_1 FILLER_18_373 ();
 sg13g2_fill_2 FILLER_18_408 ();
 sg13g2_decap_8 FILLER_18_414 ();
 sg13g2_decap_8 FILLER_18_421 ();
 sg13g2_fill_2 FILLER_18_428 ();
 sg13g2_decap_8 FILLER_19_0 ();
 sg13g2_decap_4 FILLER_19_7 ();
 sg13g2_decap_8 FILLER_19_29 ();
 sg13g2_decap_4 FILLER_19_65 ();
 sg13g2_fill_2 FILLER_19_69 ();
 sg13g2_decap_4 FILLER_19_85 ();
 sg13g2_fill_1 FILLER_19_102 ();
 sg13g2_decap_4 FILLER_19_107 ();
 sg13g2_decap_4 FILLER_19_116 ();
 sg13g2_fill_2 FILLER_19_120 ();
 sg13g2_decap_4 FILLER_19_126 ();
 sg13g2_fill_1 FILLER_19_130 ();
 sg13g2_fill_1 FILLER_19_175 ();
 sg13g2_fill_2 FILLER_19_182 ();
 sg13g2_fill_1 FILLER_19_184 ();
 sg13g2_fill_2 FILLER_19_195 ();
 sg13g2_fill_1 FILLER_19_204 ();
 sg13g2_fill_1 FILLER_19_210 ();
 sg13g2_decap_8 FILLER_19_227 ();
 sg13g2_decap_8 FILLER_19_243 ();
 sg13g2_fill_1 FILLER_19_250 ();
 sg13g2_decap_8 FILLER_19_256 ();
 sg13g2_fill_1 FILLER_19_263 ();
 sg13g2_fill_2 FILLER_19_269 ();
 sg13g2_fill_1 FILLER_19_275 ();
 sg13g2_fill_2 FILLER_19_286 ();
 sg13g2_fill_1 FILLER_19_288 ();
 sg13g2_decap_4 FILLER_19_300 ();
 sg13g2_decap_4 FILLER_19_310 ();
 sg13g2_fill_2 FILLER_19_314 ();
 sg13g2_decap_4 FILLER_19_322 ();
 sg13g2_fill_1 FILLER_19_326 ();
 sg13g2_decap_8 FILLER_19_337 ();
 sg13g2_decap_8 FILLER_19_344 ();
 sg13g2_decap_4 FILLER_19_351 ();
 sg13g2_fill_2 FILLER_19_367 ();
 sg13g2_fill_2 FILLER_19_373 ();
 sg13g2_fill_1 FILLER_19_375 ();
 sg13g2_decap_8 FILLER_19_399 ();
 sg13g2_decap_8 FILLER_19_406 ();
 sg13g2_decap_8 FILLER_19_413 ();
 sg13g2_decap_8 FILLER_19_420 ();
 sg13g2_fill_2 FILLER_19_427 ();
 sg13g2_fill_1 FILLER_19_429 ();
 sg13g2_decap_4 FILLER_20_0 ();
 sg13g2_fill_2 FILLER_20_4 ();
 sg13g2_fill_2 FILLER_20_27 ();
 sg13g2_fill_1 FILLER_20_29 ();
 sg13g2_decap_4 FILLER_20_38 ();
 sg13g2_fill_2 FILLER_20_42 ();
 sg13g2_decap_8 FILLER_20_52 ();
 sg13g2_decap_8 FILLER_20_59 ();
 sg13g2_fill_1 FILLER_20_66 ();
 sg13g2_fill_2 FILLER_20_80 ();
 sg13g2_fill_1 FILLER_20_82 ();
 sg13g2_fill_1 FILLER_20_97 ();
 sg13g2_fill_1 FILLER_20_107 ();
 sg13g2_decap_8 FILLER_20_112 ();
 sg13g2_decap_8 FILLER_20_119 ();
 sg13g2_decap_8 FILLER_20_126 ();
 sg13g2_fill_2 FILLER_20_133 ();
 sg13g2_fill_1 FILLER_20_140 ();
 sg13g2_fill_1 FILLER_20_146 ();
 sg13g2_fill_2 FILLER_20_152 ();
 sg13g2_fill_2 FILLER_20_159 ();
 sg13g2_fill_2 FILLER_20_167 ();
 sg13g2_fill_1 FILLER_20_169 ();
 sg13g2_fill_1 FILLER_20_174 ();
 sg13g2_fill_2 FILLER_20_183 ();
 sg13g2_fill_1 FILLER_20_189 ();
 sg13g2_fill_1 FILLER_20_199 ();
 sg13g2_decap_8 FILLER_20_204 ();
 sg13g2_decap_8 FILLER_20_224 ();
 sg13g2_decap_8 FILLER_20_231 ();
 sg13g2_decap_8 FILLER_20_238 ();
 sg13g2_decap_4 FILLER_20_245 ();
 sg13g2_fill_1 FILLER_20_249 ();
 sg13g2_decap_8 FILLER_20_258 ();
 sg13g2_fill_1 FILLER_20_269 ();
 sg13g2_fill_1 FILLER_20_283 ();
 sg13g2_fill_1 FILLER_20_289 ();
 sg13g2_fill_1 FILLER_20_295 ();
 sg13g2_decap_8 FILLER_20_301 ();
 sg13g2_decap_8 FILLER_20_308 ();
 sg13g2_fill_1 FILLER_20_323 ();
 sg13g2_fill_1 FILLER_20_328 ();
 sg13g2_fill_2 FILLER_20_357 ();
 sg13g2_fill_1 FILLER_20_359 ();
 sg13g2_fill_1 FILLER_20_407 ();
 sg13g2_fill_2 FILLER_20_413 ();
 sg13g2_decap_8 FILLER_20_420 ();
 sg13g2_fill_2 FILLER_20_427 ();
 sg13g2_fill_1 FILLER_20_429 ();
 sg13g2_decap_8 FILLER_21_0 ();
 sg13g2_fill_1 FILLER_21_7 ();
 sg13g2_fill_2 FILLER_21_13 ();
 sg13g2_fill_1 FILLER_21_15 ();
 sg13g2_decap_8 FILLER_21_20 ();
 sg13g2_fill_2 FILLER_21_27 ();
 sg13g2_fill_1 FILLER_21_42 ();
 sg13g2_fill_2 FILLER_21_51 ();
 sg13g2_fill_1 FILLER_21_53 ();
 sg13g2_decap_8 FILLER_21_67 ();
 sg13g2_decap_8 FILLER_21_74 ();
 sg13g2_decap_8 FILLER_21_81 ();
 sg13g2_fill_2 FILLER_21_88 ();
 sg13g2_decap_4 FILLER_21_110 ();
 sg13g2_fill_2 FILLER_21_114 ();
 sg13g2_decap_8 FILLER_21_124 ();
 sg13g2_fill_2 FILLER_21_140 ();
 sg13g2_fill_1 FILLER_21_154 ();
 sg13g2_fill_2 FILLER_21_174 ();
 sg13g2_fill_1 FILLER_21_176 ();
 sg13g2_decap_8 FILLER_21_182 ();
 sg13g2_decap_4 FILLER_21_210 ();
 sg13g2_fill_1 FILLER_21_214 ();
 sg13g2_decap_8 FILLER_21_223 ();
 sg13g2_decap_8 FILLER_21_230 ();
 sg13g2_fill_1 FILLER_21_237 ();
 sg13g2_fill_2 FILLER_21_249 ();
 sg13g2_fill_1 FILLER_21_251 ();
 sg13g2_decap_4 FILLER_21_272 ();
 sg13g2_fill_2 FILLER_21_276 ();
 sg13g2_fill_2 FILLER_21_283 ();
 sg13g2_fill_2 FILLER_21_298 ();
 sg13g2_decap_8 FILLER_21_305 ();
 sg13g2_decap_4 FILLER_21_312 ();
 sg13g2_fill_1 FILLER_21_324 ();
 sg13g2_decap_8 FILLER_21_329 ();
 sg13g2_decap_8 FILLER_21_336 ();
 sg13g2_fill_2 FILLER_21_352 ();
 sg13g2_fill_2 FILLER_21_359 ();
 sg13g2_fill_1 FILLER_21_361 ();
 sg13g2_fill_2 FILLER_21_372 ();
 sg13g2_fill_1 FILLER_21_415 ();
 sg13g2_decap_4 FILLER_21_426 ();
 sg13g2_decap_4 FILLER_22_0 ();
 sg13g2_fill_2 FILLER_22_4 ();
 sg13g2_fill_2 FILLER_22_11 ();
 sg13g2_fill_1 FILLER_22_13 ();
 sg13g2_decap_8 FILLER_22_22 ();
 sg13g2_decap_8 FILLER_22_29 ();
 sg13g2_decap_8 FILLER_22_36 ();
 sg13g2_fill_2 FILLER_22_43 ();
 sg13g2_fill_2 FILLER_22_49 ();
 sg13g2_fill_1 FILLER_22_51 ();
 sg13g2_decap_8 FILLER_22_56 ();
 sg13g2_fill_2 FILLER_22_63 ();
 sg13g2_fill_1 FILLER_22_65 ();
 sg13g2_decap_4 FILLER_22_79 ();
 sg13g2_fill_1 FILLER_22_83 ();
 sg13g2_decap_8 FILLER_22_113 ();
 sg13g2_decap_4 FILLER_22_120 ();
 sg13g2_decap_8 FILLER_22_128 ();
 sg13g2_decap_4 FILLER_22_135 ();
 sg13g2_fill_1 FILLER_22_174 ();
 sg13g2_fill_2 FILLER_22_179 ();
 sg13g2_decap_8 FILLER_22_193 ();
 sg13g2_fill_2 FILLER_22_200 ();
 sg13g2_decap_8 FILLER_22_221 ();
 sg13g2_decap_8 FILLER_22_228 ();
 sg13g2_fill_2 FILLER_22_240 ();
 sg13g2_fill_1 FILLER_22_242 ();
 sg13g2_fill_1 FILLER_22_256 ();
 sg13g2_fill_2 FILLER_22_262 ();
 sg13g2_fill_1 FILLER_22_278 ();
 sg13g2_decap_4 FILLER_22_288 ();
 sg13g2_fill_2 FILLER_22_296 ();
 sg13g2_fill_1 FILLER_22_298 ();
 sg13g2_fill_2 FILLER_22_306 ();
 sg13g2_decap_4 FILLER_22_317 ();
 sg13g2_fill_1 FILLER_22_321 ();
 sg13g2_fill_1 FILLER_22_328 ();
 sg13g2_decap_8 FILLER_22_345 ();
 sg13g2_fill_2 FILLER_22_352 ();
 sg13g2_fill_1 FILLER_22_354 ();
 sg13g2_fill_2 FILLER_22_379 ();
 sg13g2_fill_2 FILLER_22_386 ();
 sg13g2_fill_1 FILLER_22_388 ();
 sg13g2_fill_2 FILLER_22_397 ();
 sg13g2_fill_1 FILLER_22_399 ();
 sg13g2_fill_2 FILLER_22_405 ();
 sg13g2_decap_4 FILLER_22_413 ();
 sg13g2_decap_8 FILLER_22_422 ();
 sg13g2_fill_1 FILLER_22_429 ();
 sg13g2_decap_4 FILLER_23_0 ();
 sg13g2_fill_1 FILLER_23_4 ();
 sg13g2_fill_1 FILLER_23_18 ();
 sg13g2_fill_2 FILLER_23_24 ();
 sg13g2_decap_4 FILLER_23_30 ();
 sg13g2_decap_4 FILLER_23_43 ();
 sg13g2_decap_4 FILLER_23_55 ();
 sg13g2_fill_1 FILLER_23_59 ();
 sg13g2_decap_8 FILLER_23_76 ();
 sg13g2_fill_1 FILLER_23_88 ();
 sg13g2_fill_2 FILLER_23_93 ();
 sg13g2_fill_1 FILLER_23_95 ();
 sg13g2_decap_4 FILLER_23_108 ();
 sg13g2_decap_8 FILLER_23_117 ();
 sg13g2_decap_8 FILLER_23_124 ();
 sg13g2_decap_8 FILLER_23_131 ();
 sg13g2_fill_1 FILLER_23_152 ();
 sg13g2_fill_2 FILLER_23_173 ();
 sg13g2_fill_2 FILLER_23_179 ();
 sg13g2_fill_1 FILLER_23_181 ();
 sg13g2_fill_1 FILLER_23_187 ();
 sg13g2_fill_1 FILLER_23_192 ();
 sg13g2_fill_1 FILLER_23_214 ();
 sg13g2_fill_2 FILLER_23_220 ();
 sg13g2_decap_8 FILLER_23_230 ();
 sg13g2_decap_4 FILLER_23_237 ();
 sg13g2_fill_2 FILLER_23_241 ();
 sg13g2_fill_2 FILLER_23_260 ();
 sg13g2_decap_4 FILLER_23_270 ();
 sg13g2_fill_1 FILLER_23_274 ();
 sg13g2_decap_8 FILLER_23_279 ();
 sg13g2_decap_8 FILLER_23_286 ();
 sg13g2_decap_8 FILLER_23_293 ();
 sg13g2_decap_8 FILLER_23_308 ();
 sg13g2_fill_1 FILLER_23_315 ();
 sg13g2_decap_8 FILLER_23_340 ();
 sg13g2_decap_4 FILLER_23_347 ();
 sg13g2_fill_1 FILLER_23_372 ();
 sg13g2_fill_1 FILLER_23_382 ();
 sg13g2_decap_4 FILLER_23_393 ();
 sg13g2_fill_2 FILLER_23_414 ();
 sg13g2_decap_8 FILLER_23_421 ();
 sg13g2_fill_2 FILLER_23_428 ();
 sg13g2_decap_4 FILLER_24_0 ();
 sg13g2_fill_2 FILLER_24_4 ();
 sg13g2_fill_2 FILLER_24_19 ();
 sg13g2_fill_1 FILLER_24_21 ();
 sg13g2_decap_4 FILLER_24_28 ();
 sg13g2_decap_8 FILLER_24_61 ();
 sg13g2_decap_8 FILLER_24_68 ();
 sg13g2_fill_1 FILLER_24_101 ();
 sg13g2_fill_2 FILLER_24_108 ();
 sg13g2_decap_8 FILLER_24_114 ();
 sg13g2_decap_8 FILLER_24_121 ();
 sg13g2_fill_2 FILLER_24_128 ();
 sg13g2_decap_4 FILLER_24_186 ();
 sg13g2_fill_1 FILLER_24_190 ();
 sg13g2_fill_1 FILLER_24_195 ();
 sg13g2_fill_2 FILLER_24_200 ();
 sg13g2_fill_2 FILLER_24_215 ();
 sg13g2_decap_4 FILLER_24_221 ();
 sg13g2_fill_1 FILLER_24_225 ();
 sg13g2_decap_8 FILLER_24_234 ();
 sg13g2_decap_8 FILLER_24_241 ();
 sg13g2_fill_2 FILLER_24_248 ();
 sg13g2_fill_1 FILLER_24_260 ();
 sg13g2_fill_2 FILLER_24_269 ();
 sg13g2_fill_1 FILLER_24_271 ();
 sg13g2_fill_1 FILLER_24_286 ();
 sg13g2_fill_1 FILLER_24_292 ();
 sg13g2_fill_1 FILLER_24_297 ();
 sg13g2_fill_2 FILLER_24_304 ();
 sg13g2_fill_1 FILLER_24_310 ();
 sg13g2_decap_4 FILLER_24_316 ();
 sg13g2_decap_8 FILLER_24_333 ();
 sg13g2_decap_8 FILLER_24_340 ();
 sg13g2_decap_8 FILLER_24_347 ();
 sg13g2_fill_2 FILLER_24_354 ();
 sg13g2_fill_1 FILLER_24_356 ();
 sg13g2_decap_8 FILLER_24_384 ();
 sg13g2_decap_8 FILLER_24_391 ();
 sg13g2_fill_1 FILLER_24_402 ();
 sg13g2_decap_4 FILLER_24_424 ();
 sg13g2_fill_2 FILLER_24_428 ();
 sg13g2_decap_8 FILLER_25_0 ();
 sg13g2_fill_2 FILLER_25_7 ();
 sg13g2_fill_2 FILLER_25_20 ();
 sg13g2_decap_4 FILLER_25_27 ();
 sg13g2_decap_8 FILLER_25_39 ();
 sg13g2_decap_8 FILLER_25_46 ();
 sg13g2_decap_8 FILLER_25_53 ();
 sg13g2_decap_8 FILLER_25_60 ();
 sg13g2_decap_4 FILLER_25_67 ();
 sg13g2_fill_2 FILLER_25_71 ();
 sg13g2_decap_4 FILLER_25_81 ();
 sg13g2_fill_2 FILLER_25_85 ();
 sg13g2_decap_4 FILLER_25_99 ();
 sg13g2_fill_1 FILLER_25_103 ();
 sg13g2_fill_2 FILLER_25_108 ();
 sg13g2_fill_1 FILLER_25_110 ();
 sg13g2_decap_8 FILLER_25_119 ();
 sg13g2_fill_2 FILLER_25_126 ();
 sg13g2_fill_2 FILLER_25_138 ();
 sg13g2_decap_4 FILLER_25_160 ();
 sg13g2_fill_2 FILLER_25_188 ();
 sg13g2_decap_8 FILLER_25_194 ();
 sg13g2_fill_1 FILLER_25_201 ();
 sg13g2_decap_8 FILLER_25_224 ();
 sg13g2_decap_8 FILLER_25_231 ();
 sg13g2_decap_4 FILLER_25_238 ();
 sg13g2_fill_2 FILLER_25_242 ();
 sg13g2_decap_4 FILLER_25_257 ();
 sg13g2_fill_1 FILLER_25_261 ();
 sg13g2_decap_8 FILLER_25_266 ();
 sg13g2_decap_4 FILLER_25_273 ();
 sg13g2_fill_1 FILLER_25_277 ();
 sg13g2_decap_8 FILLER_25_304 ();
 sg13g2_decap_8 FILLER_25_311 ();
 sg13g2_fill_1 FILLER_25_318 ();
 sg13g2_decap_4 FILLER_25_343 ();
 sg13g2_fill_1 FILLER_25_361 ();
 sg13g2_fill_1 FILLER_25_376 ();
 sg13g2_decap_8 FILLER_25_382 ();
 sg13g2_decap_8 FILLER_25_389 ();
 sg13g2_decap_8 FILLER_25_418 ();
 sg13g2_decap_4 FILLER_25_425 ();
 sg13g2_fill_1 FILLER_25_429 ();
 sg13g2_decap_8 FILLER_26_0 ();
 sg13g2_fill_2 FILLER_26_7 ();
 sg13g2_fill_1 FILLER_26_9 ();
 sg13g2_decap_8 FILLER_26_26 ();
 sg13g2_decap_4 FILLER_26_33 ();
 sg13g2_fill_1 FILLER_26_45 ();
 sg13g2_fill_1 FILLER_26_72 ();
 sg13g2_decap_8 FILLER_26_99 ();
 sg13g2_fill_2 FILLER_26_114 ();
 sg13g2_fill_1 FILLER_26_116 ();
 sg13g2_decap_4 FILLER_26_122 ();
 sg13g2_fill_1 FILLER_26_126 ();
 sg13g2_decap_8 FILLER_26_132 ();
 sg13g2_decap_8 FILLER_26_139 ();
 sg13g2_fill_1 FILLER_26_146 ();
 sg13g2_decap_4 FILLER_26_171 ();
 sg13g2_decap_4 FILLER_26_186 ();
 sg13g2_fill_1 FILLER_26_190 ();
 sg13g2_fill_1 FILLER_26_197 ();
 sg13g2_fill_1 FILLER_26_202 ();
 sg13g2_decap_8 FILLER_26_215 ();
 sg13g2_fill_1 FILLER_26_222 ();
 sg13g2_decap_8 FILLER_26_231 ();
 sg13g2_decap_8 FILLER_26_238 ();
 sg13g2_fill_2 FILLER_26_245 ();
 sg13g2_decap_8 FILLER_26_259 ();
 sg13g2_fill_2 FILLER_26_266 ();
 sg13g2_fill_1 FILLER_26_268 ();
 sg13g2_decap_8 FILLER_26_277 ();
 sg13g2_fill_1 FILLER_26_284 ();
 sg13g2_decap_8 FILLER_26_297 ();
 sg13g2_decap_4 FILLER_26_304 ();
 sg13g2_decap_8 FILLER_26_316 ();
 sg13g2_fill_2 FILLER_26_323 ();
 sg13g2_fill_1 FILLER_26_325 ();
 sg13g2_decap_8 FILLER_26_332 ();
 sg13g2_decap_8 FILLER_26_339 ();
 sg13g2_fill_2 FILLER_26_370 ();
 sg13g2_fill_2 FILLER_26_379 ();
 sg13g2_fill_1 FILLER_26_381 ();
 sg13g2_decap_4 FILLER_26_392 ();
 sg13g2_fill_1 FILLER_26_396 ();
 sg13g2_fill_1 FILLER_26_416 ();
 sg13g2_decap_4 FILLER_26_425 ();
 sg13g2_fill_1 FILLER_26_429 ();
 sg13g2_decap_4 FILLER_27_0 ();
 sg13g2_fill_2 FILLER_27_4 ();
 sg13g2_fill_1 FILLER_27_14 ();
 sg13g2_fill_2 FILLER_27_19 ();
 sg13g2_fill_2 FILLER_27_51 ();
 sg13g2_fill_1 FILLER_27_57 ();
 sg13g2_decap_8 FILLER_27_62 ();
 sg13g2_decap_8 FILLER_27_69 ();
 sg13g2_decap_4 FILLER_27_76 ();
 sg13g2_fill_1 FILLER_27_80 ();
 sg13g2_decap_8 FILLER_27_98 ();
 sg13g2_fill_1 FILLER_27_113 ();
 sg13g2_fill_1 FILLER_27_123 ();
 sg13g2_fill_2 FILLER_27_128 ();
 sg13g2_decap_8 FILLER_27_134 ();
 sg13g2_decap_8 FILLER_27_141 ();
 sg13g2_decap_8 FILLER_27_148 ();
 sg13g2_decap_8 FILLER_27_155 ();
 sg13g2_decap_8 FILLER_27_162 ();
 sg13g2_decap_8 FILLER_27_169 ();
 sg13g2_decap_4 FILLER_27_176 ();
 sg13g2_decap_8 FILLER_27_190 ();
 sg13g2_decap_4 FILLER_27_197 ();
 sg13g2_fill_1 FILLER_27_201 ();
 sg13g2_decap_8 FILLER_27_233 ();
 sg13g2_fill_1 FILLER_27_240 ();
 sg13g2_decap_4 FILLER_27_302 ();
 sg13g2_fill_1 FILLER_27_306 ();
 sg13g2_fill_1 FILLER_27_312 ();
 sg13g2_fill_2 FILLER_27_318 ();
 sg13g2_fill_1 FILLER_27_320 ();
 sg13g2_fill_1 FILLER_27_325 ();
 sg13g2_decap_4 FILLER_27_330 ();
 sg13g2_decap_4 FILLER_27_338 ();
 sg13g2_fill_1 FILLER_27_342 ();
 sg13g2_fill_2 FILLER_27_349 ();
 sg13g2_fill_2 FILLER_27_359 ();
 sg13g2_fill_2 FILLER_27_367 ();
 sg13g2_fill_1 FILLER_27_369 ();
 sg13g2_fill_1 FILLER_27_375 ();
 sg13g2_decap_8 FILLER_27_384 ();
 sg13g2_decap_8 FILLER_27_391 ();
 sg13g2_decap_4 FILLER_27_398 ();
 sg13g2_decap_8 FILLER_27_406 ();
 sg13g2_fill_2 FILLER_27_413 ();
 sg13g2_decap_8 FILLER_27_420 ();
 sg13g2_fill_2 FILLER_27_427 ();
 sg13g2_fill_1 FILLER_27_429 ();
 sg13g2_decap_8 FILLER_28_0 ();
 sg13g2_decap_4 FILLER_28_7 ();
 sg13g2_fill_1 FILLER_28_11 ();
 sg13g2_decap_8 FILLER_28_20 ();
 sg13g2_decap_4 FILLER_28_27 ();
 sg13g2_fill_2 FILLER_28_31 ();
 sg13g2_decap_4 FILLER_28_37 ();
 sg13g2_fill_2 FILLER_28_41 ();
 sg13g2_decap_8 FILLER_28_76 ();
 sg13g2_fill_2 FILLER_28_83 ();
 sg13g2_fill_1 FILLER_28_85 ();
 sg13g2_fill_1 FILLER_28_106 ();
 sg13g2_decap_8 FILLER_28_116 ();
 sg13g2_decap_8 FILLER_28_123 ();
 sg13g2_fill_1 FILLER_28_130 ();
 sg13g2_fill_2 FILLER_28_148 ();
 sg13g2_fill_1 FILLER_28_150 ();
 sg13g2_decap_4 FILLER_28_169 ();
 sg13g2_fill_1 FILLER_28_173 ();
 sg13g2_fill_2 FILLER_28_182 ();
 sg13g2_fill_2 FILLER_28_188 ();
 sg13g2_decap_8 FILLER_28_220 ();
 sg13g2_decap_4 FILLER_28_227 ();
 sg13g2_fill_2 FILLER_28_231 ();
 sg13g2_fill_1 FILLER_28_241 ();
 sg13g2_fill_1 FILLER_28_246 ();
 sg13g2_fill_1 FILLER_28_255 ();
 sg13g2_fill_2 FILLER_28_264 ();
 sg13g2_decap_4 FILLER_28_270 ();
 sg13g2_fill_2 FILLER_28_301 ();
 sg13g2_decap_8 FILLER_28_307 ();
 sg13g2_fill_2 FILLER_28_314 ();
 sg13g2_fill_1 FILLER_28_316 ();
 sg13g2_fill_2 FILLER_28_344 ();
 sg13g2_fill_1 FILLER_28_346 ();
 sg13g2_fill_1 FILLER_28_357 ();
 sg13g2_decap_4 FILLER_28_376 ();
 sg13g2_decap_8 FILLER_28_385 ();
 sg13g2_decap_8 FILLER_28_392 ();
 sg13g2_decap_8 FILLER_28_399 ();
 sg13g2_decap_8 FILLER_28_423 ();
 sg13g2_decap_8 FILLER_29_0 ();
 sg13g2_fill_1 FILLER_29_7 ();
 sg13g2_fill_1 FILLER_29_16 ();
 sg13g2_fill_2 FILLER_29_21 ();
 sg13g2_fill_2 FILLER_29_49 ();
 sg13g2_fill_1 FILLER_29_51 ();
 sg13g2_decap_8 FILLER_29_56 ();
 sg13g2_fill_1 FILLER_29_63 ();
 sg13g2_decap_4 FILLER_29_84 ();
 sg13g2_fill_1 FILLER_29_88 ();
 sg13g2_fill_1 FILLER_29_99 ();
 sg13g2_decap_8 FILLER_29_116 ();
 sg13g2_fill_2 FILLER_29_140 ();
 sg13g2_decap_8 FILLER_29_155 ();
 sg13g2_decap_4 FILLER_29_162 ();
 sg13g2_fill_1 FILLER_29_166 ();
 sg13g2_fill_2 FILLER_29_177 ();
 sg13g2_fill_1 FILLER_29_188 ();
 sg13g2_fill_1 FILLER_29_198 ();
 sg13g2_fill_2 FILLER_29_203 ();
 sg13g2_decap_8 FILLER_29_251 ();
 sg13g2_decap_4 FILLER_29_258 ();
 sg13g2_fill_1 FILLER_29_262 ();
 sg13g2_decap_8 FILLER_29_268 ();
 sg13g2_fill_2 FILLER_29_275 ();
 sg13g2_fill_1 FILLER_29_277 ();
 sg13g2_fill_2 FILLER_29_284 ();
 sg13g2_decap_4 FILLER_29_304 ();
 sg13g2_fill_1 FILLER_29_308 ();
 sg13g2_fill_2 FILLER_29_327 ();
 sg13g2_fill_1 FILLER_29_329 ();
 sg13g2_decap_4 FILLER_29_346 ();
 sg13g2_fill_1 FILLER_29_350 ();
 sg13g2_decap_4 FILLER_29_365 ();
 sg13g2_fill_2 FILLER_29_369 ();
 sg13g2_decap_8 FILLER_29_375 ();
 sg13g2_decap_8 FILLER_29_382 ();
 sg13g2_decap_4 FILLER_29_401 ();
 sg13g2_fill_1 FILLER_29_412 ();
 sg13g2_decap_4 FILLER_29_424 ();
 sg13g2_fill_2 FILLER_29_428 ();
 sg13g2_decap_8 FILLER_30_0 ();
 sg13g2_decap_8 FILLER_30_7 ();
 sg13g2_decap_8 FILLER_30_23 ();
 sg13g2_fill_2 FILLER_30_34 ();
 sg13g2_fill_1 FILLER_30_36 ();
 sg13g2_decap_8 FILLER_30_41 ();
 sg13g2_decap_8 FILLER_30_48 ();
 sg13g2_decap_8 FILLER_30_55 ();
 sg13g2_decap_8 FILLER_30_62 ();
 sg13g2_decap_4 FILLER_30_69 ();
 sg13g2_fill_2 FILLER_30_73 ();
 sg13g2_fill_2 FILLER_30_98 ();
 sg13g2_fill_1 FILLER_30_100 ();
 sg13g2_decap_4 FILLER_30_109 ();
 sg13g2_decap_4 FILLER_30_117 ();
 sg13g2_fill_1 FILLER_30_121 ();
 sg13g2_decap_8 FILLER_30_149 ();
 sg13g2_decap_8 FILLER_30_156 ();
 sg13g2_fill_2 FILLER_30_163 ();
 sg13g2_fill_1 FILLER_30_187 ();
 sg13g2_fill_1 FILLER_30_201 ();
 sg13g2_decap_8 FILLER_30_211 ();
 sg13g2_fill_2 FILLER_30_218 ();
 sg13g2_decap_8 FILLER_30_224 ();
 sg13g2_decap_8 FILLER_30_231 ();
 sg13g2_decap_8 FILLER_30_238 ();
 sg13g2_decap_4 FILLER_30_245 ();
 sg13g2_decap_4 FILLER_30_252 ();
 sg13g2_fill_1 FILLER_30_256 ();
 sg13g2_decap_8 FILLER_30_270 ();
 sg13g2_decap_4 FILLER_30_277 ();
 sg13g2_fill_1 FILLER_30_281 ();
 sg13g2_fill_2 FILLER_30_287 ();
 sg13g2_fill_1 FILLER_30_289 ();
 sg13g2_fill_2 FILLER_30_300 ();
 sg13g2_fill_1 FILLER_30_302 ();
 sg13g2_decap_8 FILLER_30_311 ();
 sg13g2_decap_4 FILLER_30_318 ();
 sg13g2_fill_1 FILLER_30_322 ();
 sg13g2_decap_8 FILLER_30_336 ();
 sg13g2_fill_2 FILLER_30_343 ();
 sg13g2_fill_1 FILLER_30_345 ();
 sg13g2_decap_8 FILLER_30_351 ();
 sg13g2_fill_1 FILLER_30_358 ();
 sg13g2_fill_2 FILLER_30_375 ();
 sg13g2_fill_1 FILLER_30_377 ();
 sg13g2_fill_1 FILLER_30_387 ();
 sg13g2_fill_1 FILLER_30_395 ();
 sg13g2_fill_2 FILLER_30_404 ();
 sg13g2_fill_2 FILLER_30_419 ();
 sg13g2_fill_1 FILLER_30_421 ();
 sg13g2_decap_8 FILLER_31_0 ();
 sg13g2_decap_8 FILLER_31_7 ();
 sg13g2_fill_2 FILLER_31_14 ();
 sg13g2_fill_1 FILLER_31_16 ();
 sg13g2_fill_2 FILLER_31_28 ();
 sg13g2_decap_8 FILLER_31_56 ();
 sg13g2_decap_8 FILLER_31_63 ();
 sg13g2_decap_8 FILLER_31_70 ();
 sg13g2_fill_1 FILLER_31_77 ();
 sg13g2_fill_2 FILLER_31_83 ();
 sg13g2_decap_8 FILLER_31_106 ();
 sg13g2_decap_8 FILLER_31_113 ();
 sg13g2_decap_4 FILLER_31_120 ();
 sg13g2_fill_1 FILLER_31_128 ();
 sg13g2_fill_1 FILLER_31_137 ();
 sg13g2_decap_8 FILLER_31_143 ();
 sg13g2_fill_1 FILLER_31_158 ();
 sg13g2_fill_1 FILLER_31_184 ();
 sg13g2_fill_1 FILLER_31_193 ();
 sg13g2_fill_2 FILLER_31_198 ();
 sg13g2_fill_1 FILLER_31_208 ();
 sg13g2_fill_1 FILLER_31_217 ();
 sg13g2_fill_1 FILLER_31_223 ();
 sg13g2_fill_2 FILLER_31_228 ();
 sg13g2_fill_1 FILLER_31_256 ();
 sg13g2_decap_8 FILLER_31_265 ();
 sg13g2_fill_1 FILLER_31_272 ();
 sg13g2_fill_2 FILLER_31_297 ();
 sg13g2_decap_8 FILLER_31_307 ();
 sg13g2_fill_2 FILLER_31_314 ();
 sg13g2_fill_1 FILLER_31_325 ();
 sg13g2_decap_8 FILLER_31_342 ();
 sg13g2_decap_8 FILLER_31_349 ();
 sg13g2_decap_8 FILLER_31_356 ();
 sg13g2_fill_1 FILLER_31_363 ();
 sg13g2_fill_1 FILLER_31_374 ();
 sg13g2_fill_1 FILLER_31_378 ();
 sg13g2_fill_1 FILLER_31_404 ();
 sg13g2_decap_4 FILLER_31_410 ();
 sg13g2_fill_1 FILLER_31_414 ();
 sg13g2_decap_8 FILLER_31_423 ();
 sg13g2_decap_8 FILLER_32_0 ();
 sg13g2_decap_8 FILLER_32_7 ();
 sg13g2_decap_8 FILLER_32_14 ();
 sg13g2_decap_8 FILLER_32_21 ();
 sg13g2_decap_8 FILLER_32_28 ();
 sg13g2_decap_4 FILLER_32_35 ();
 sg13g2_fill_2 FILLER_32_39 ();
 sg13g2_fill_1 FILLER_32_49 ();
 sg13g2_decap_8 FILLER_32_55 ();
 sg13g2_decap_4 FILLER_32_62 ();
 sg13g2_fill_1 FILLER_32_66 ();
 sg13g2_fill_1 FILLER_32_71 ();
 sg13g2_fill_1 FILLER_32_81 ();
 sg13g2_decap_8 FILLER_32_86 ();
 sg13g2_decap_8 FILLER_32_93 ();
 sg13g2_fill_2 FILLER_32_100 ();
 sg13g2_decap_8 FILLER_32_110 ();
 sg13g2_decap_8 FILLER_32_117 ();
 sg13g2_decap_4 FILLER_32_136 ();
 sg13g2_decap_8 FILLER_32_152 ();
 sg13g2_decap_8 FILLER_32_174 ();
 sg13g2_decap_8 FILLER_32_181 ();
 sg13g2_decap_8 FILLER_32_188 ();
 sg13g2_fill_2 FILLER_32_195 ();
 sg13g2_decap_4 FILLER_32_201 ();
 sg13g2_fill_1 FILLER_32_205 ();
 sg13g2_fill_1 FILLER_32_211 ();
 sg13g2_fill_1 FILLER_32_222 ();
 sg13g2_decap_4 FILLER_32_231 ();
 sg13g2_fill_2 FILLER_32_235 ();
 sg13g2_decap_8 FILLER_32_241 ();
 sg13g2_fill_2 FILLER_32_251 ();
 sg13g2_fill_1 FILLER_32_253 ();
 sg13g2_decap_8 FILLER_32_258 ();
 sg13g2_decap_8 FILLER_32_265 ();
 sg13g2_decap_8 FILLER_32_272 ();
 sg13g2_decap_8 FILLER_32_279 ();
 sg13g2_decap_4 FILLER_32_286 ();
 sg13g2_decap_8 FILLER_32_297 ();
 sg13g2_decap_8 FILLER_32_304 ();
 sg13g2_fill_2 FILLER_32_323 ();
 sg13g2_decap_4 FILLER_32_333 ();
 sg13g2_fill_1 FILLER_32_337 ();
 sg13g2_decap_8 FILLER_32_351 ();
 sg13g2_fill_2 FILLER_32_358 ();
 sg13g2_decap_8 FILLER_32_370 ();
 sg13g2_decap_4 FILLER_32_410 ();
 sg13g2_fill_2 FILLER_32_414 ();
 sg13g2_decap_8 FILLER_32_423 ();
 sg13g2_decap_8 FILLER_33_0 ();
 sg13g2_decap_8 FILLER_33_7 ();
 sg13g2_decap_8 FILLER_33_14 ();
 sg13g2_decap_8 FILLER_33_21 ();
 sg13g2_decap_8 FILLER_33_28 ();
 sg13g2_decap_8 FILLER_33_35 ();
 sg13g2_decap_8 FILLER_33_54 ();
 sg13g2_fill_2 FILLER_33_61 ();
 sg13g2_fill_2 FILLER_33_78 ();
 sg13g2_fill_2 FILLER_33_85 ();
 sg13g2_fill_1 FILLER_33_87 ();
 sg13g2_fill_1 FILLER_33_96 ();
 sg13g2_fill_2 FILLER_33_105 ();
 sg13g2_fill_2 FILLER_33_154 ();
 sg13g2_fill_2 FILLER_33_164 ();
 sg13g2_decap_4 FILLER_33_182 ();
 sg13g2_fill_2 FILLER_33_190 ();
 sg13g2_fill_1 FILLER_33_192 ();
 sg13g2_fill_1 FILLER_33_201 ();
 sg13g2_decap_4 FILLER_33_225 ();
 sg13g2_decap_4 FILLER_33_234 ();
 sg13g2_decap_4 FILLER_33_242 ();
 sg13g2_decap_8 FILLER_33_251 ();
 sg13g2_decap_8 FILLER_33_258 ();
 sg13g2_decap_8 FILLER_33_265 ();
 sg13g2_decap_8 FILLER_33_272 ();
 sg13g2_decap_8 FILLER_33_279 ();
 sg13g2_decap_8 FILLER_33_286 ();
 sg13g2_fill_1 FILLER_33_293 ();
 sg13g2_fill_2 FILLER_33_302 ();
 sg13g2_fill_1 FILLER_33_304 ();
 sg13g2_decap_4 FILLER_33_345 ();
 sg13g2_fill_1 FILLER_33_349 ();
 sg13g2_decap_8 FILLER_33_369 ();
 sg13g2_fill_2 FILLER_33_376 ();
 sg13g2_decap_8 FILLER_33_383 ();
 sg13g2_decap_4 FILLER_33_390 ();
 sg13g2_fill_2 FILLER_33_394 ();
 sg13g2_decap_8 FILLER_33_401 ();
 sg13g2_fill_2 FILLER_33_408 ();
 sg13g2_decap_8 FILLER_33_419 ();
 sg13g2_decap_4 FILLER_33_426 ();
 sg13g2_decap_8 FILLER_34_0 ();
 sg13g2_decap_8 FILLER_34_7 ();
 sg13g2_decap_8 FILLER_34_14 ();
 sg13g2_decap_8 FILLER_34_21 ();
 sg13g2_decap_8 FILLER_34_28 ();
 sg13g2_decap_4 FILLER_34_35 ();
 sg13g2_fill_1 FILLER_34_39 ();
 sg13g2_fill_2 FILLER_34_44 ();
 sg13g2_fill_2 FILLER_34_72 ();
 sg13g2_fill_1 FILLER_34_74 ();
 sg13g2_fill_1 FILLER_34_83 ();
 sg13g2_fill_2 FILLER_34_88 ();
 sg13g2_fill_1 FILLER_34_90 ();
 sg13g2_decap_8 FILLER_34_96 ();
 sg13g2_decap_4 FILLER_34_103 ();
 sg13g2_fill_1 FILLER_34_107 ();
 sg13g2_decap_4 FILLER_34_116 ();
 sg13g2_fill_2 FILLER_34_120 ();
 sg13g2_decap_8 FILLER_34_130 ();
 sg13g2_decap_4 FILLER_34_137 ();
 sg13g2_decap_4 FILLER_34_153 ();
 sg13g2_decap_4 FILLER_34_161 ();
 sg13g2_fill_1 FILLER_34_165 ();
 sg13g2_fill_2 FILLER_34_170 ();
 sg13g2_decap_4 FILLER_34_180 ();
 sg13g2_fill_2 FILLER_34_184 ();
 sg13g2_fill_2 FILLER_34_194 ();
 sg13g2_fill_1 FILLER_34_196 ();
 sg13g2_fill_1 FILLER_34_201 ();
 sg13g2_fill_2 FILLER_34_228 ();
 sg13g2_fill_1 FILLER_34_230 ();
 sg13g2_decap_8 FILLER_34_257 ();
 sg13g2_decap_8 FILLER_34_264 ();
 sg13g2_decap_8 FILLER_34_271 ();
 sg13g2_decap_8 FILLER_34_278 ();
 sg13g2_decap_8 FILLER_34_285 ();
 sg13g2_decap_4 FILLER_34_292 ();
 sg13g2_decap_8 FILLER_34_321 ();
 sg13g2_fill_2 FILLER_34_328 ();
 sg13g2_decap_8 FILLER_34_337 ();
 sg13g2_decap_8 FILLER_34_344 ();
 sg13g2_fill_2 FILLER_34_351 ();
 sg13g2_fill_2 FILLER_34_360 ();
 sg13g2_fill_2 FILLER_34_366 ();
 sg13g2_fill_2 FILLER_34_402 ();
 sg13g2_fill_2 FILLER_34_411 ();
 sg13g2_fill_1 FILLER_34_413 ();
 sg13g2_decap_8 FILLER_34_422 ();
 sg13g2_fill_1 FILLER_34_429 ();
 sg13g2_decap_8 FILLER_35_0 ();
 sg13g2_decap_8 FILLER_35_7 ();
 sg13g2_decap_8 FILLER_35_14 ();
 sg13g2_decap_8 FILLER_35_21 ();
 sg13g2_decap_8 FILLER_35_28 ();
 sg13g2_decap_8 FILLER_35_35 ();
 sg13g2_decap_8 FILLER_35_42 ();
 sg13g2_decap_4 FILLER_35_49 ();
 sg13g2_fill_2 FILLER_35_53 ();
 sg13g2_decap_8 FILLER_35_59 ();
 sg13g2_decap_8 FILLER_35_66 ();
 sg13g2_decap_4 FILLER_35_73 ();
 sg13g2_fill_2 FILLER_35_77 ();
 sg13g2_fill_2 FILLER_35_109 ();
 sg13g2_fill_1 FILLER_35_111 ();
 sg13g2_fill_1 FILLER_35_142 ();
 sg13g2_decap_4 FILLER_35_169 ();
 sg13g2_decap_8 FILLER_35_212 ();
 sg13g2_decap_8 FILLER_35_219 ();
 sg13g2_decap_8 FILLER_35_226 ();
 sg13g2_decap_8 FILLER_35_233 ();
 sg13g2_decap_4 FILLER_35_240 ();
 sg13g2_fill_1 FILLER_35_244 ();
 sg13g2_decap_8 FILLER_35_249 ();
 sg13g2_decap_8 FILLER_35_256 ();
 sg13g2_decap_8 FILLER_35_263 ();
 sg13g2_fill_1 FILLER_35_270 ();
 sg13g2_decap_8 FILLER_35_275 ();
 sg13g2_decap_8 FILLER_35_282 ();
 sg13g2_decap_4 FILLER_35_289 ();
 sg13g2_decap_4 FILLER_35_327 ();
 sg13g2_decap_4 FILLER_35_357 ();
 sg13g2_decap_8 FILLER_35_369 ();
 sg13g2_fill_1 FILLER_35_380 ();
 sg13g2_decap_8 FILLER_35_385 ();
 sg13g2_fill_2 FILLER_35_392 ();
 sg13g2_fill_1 FILLER_35_394 ();
 sg13g2_fill_1 FILLER_35_403 ();
 sg13g2_decap_8 FILLER_36_0 ();
 sg13g2_decap_8 FILLER_36_7 ();
 sg13g2_decap_8 FILLER_36_14 ();
 sg13g2_decap_8 FILLER_36_21 ();
 sg13g2_decap_8 FILLER_36_28 ();
 sg13g2_decap_8 FILLER_36_35 ();
 sg13g2_decap_8 FILLER_36_42 ();
 sg13g2_decap_8 FILLER_36_49 ();
 sg13g2_decap_8 FILLER_36_56 ();
 sg13g2_decap_8 FILLER_36_63 ();
 sg13g2_decap_8 FILLER_36_70 ();
 sg13g2_decap_8 FILLER_36_77 ();
 sg13g2_decap_4 FILLER_36_84 ();
 sg13g2_fill_2 FILLER_36_88 ();
 sg13g2_decap_8 FILLER_36_94 ();
 sg13g2_decap_4 FILLER_36_101 ();
 sg13g2_fill_1 FILLER_36_110 ();
 sg13g2_decap_4 FILLER_36_115 ();
 sg13g2_decap_8 FILLER_36_123 ();
 sg13g2_decap_8 FILLER_36_130 ();
 sg13g2_decap_8 FILLER_36_137 ();
 sg13g2_decap_4 FILLER_36_144 ();
 sg13g2_fill_2 FILLER_36_148 ();
 sg13g2_decap_8 FILLER_36_154 ();
 sg13g2_decap_8 FILLER_36_161 ();
 sg13g2_decap_8 FILLER_36_168 ();
 sg13g2_decap_8 FILLER_36_175 ();
 sg13g2_fill_2 FILLER_36_182 ();
 sg13g2_fill_1 FILLER_36_184 ();
 sg13g2_decap_8 FILLER_36_189 ();
 sg13g2_decap_8 FILLER_36_196 ();
 sg13g2_decap_8 FILLER_36_203 ();
 sg13g2_decap_8 FILLER_36_210 ();
 sg13g2_decap_8 FILLER_36_217 ();
 sg13g2_decap_8 FILLER_36_224 ();
 sg13g2_decap_8 FILLER_36_231 ();
 sg13g2_decap_8 FILLER_36_238 ();
 sg13g2_decap_8 FILLER_36_245 ();
 sg13g2_decap_8 FILLER_36_252 ();
 sg13g2_decap_4 FILLER_36_259 ();
 sg13g2_fill_1 FILLER_36_263 ();
 sg13g2_decap_8 FILLER_36_298 ();
 sg13g2_fill_2 FILLER_36_305 ();
 sg13g2_decap_8 FILLER_36_311 ();
 sg13g2_decap_8 FILLER_36_318 ();
 sg13g2_decap_8 FILLER_36_325 ();
 sg13g2_fill_2 FILLER_36_336 ();
 sg13g2_decap_8 FILLER_36_342 ();
 sg13g2_fill_2 FILLER_36_349 ();
 sg13g2_decap_4 FILLER_36_355 ();
 sg13g2_decap_8 FILLER_36_385 ();
 sg13g2_decap_8 FILLER_36_392 ();
 sg13g2_fill_1 FILLER_36_399 ();
 sg13g2_decap_8 FILLER_37_0 ();
 sg13g2_decap_8 FILLER_37_7 ();
 sg13g2_decap_8 FILLER_37_14 ();
 sg13g2_decap_8 FILLER_37_21 ();
 sg13g2_decap_8 FILLER_37_28 ();
 sg13g2_decap_8 FILLER_37_35 ();
 sg13g2_decap_8 FILLER_37_42 ();
 sg13g2_decap_8 FILLER_37_49 ();
 sg13g2_decap_8 FILLER_37_56 ();
 sg13g2_decap_8 FILLER_37_63 ();
 sg13g2_decap_8 FILLER_37_70 ();
 sg13g2_decap_8 FILLER_37_77 ();
 sg13g2_decap_8 FILLER_37_84 ();
 sg13g2_decap_8 FILLER_37_95 ();
 sg13g2_decap_8 FILLER_37_102 ();
 sg13g2_decap_8 FILLER_37_109 ();
 sg13g2_decap_8 FILLER_37_116 ();
 sg13g2_decap_8 FILLER_37_123 ();
 sg13g2_decap_8 FILLER_37_130 ();
 sg13g2_decap_8 FILLER_37_137 ();
 sg13g2_decap_8 FILLER_37_144 ();
 sg13g2_decap_8 FILLER_37_151 ();
 sg13g2_decap_8 FILLER_37_158 ();
 sg13g2_decap_8 FILLER_37_165 ();
 sg13g2_decap_8 FILLER_37_172 ();
 sg13g2_decap_8 FILLER_37_179 ();
 sg13g2_decap_8 FILLER_37_186 ();
 sg13g2_decap_8 FILLER_37_193 ();
 sg13g2_decap_8 FILLER_37_200 ();
 sg13g2_decap_8 FILLER_37_207 ();
 sg13g2_decap_8 FILLER_37_214 ();
 sg13g2_decap_8 FILLER_37_221 ();
 sg13g2_decap_8 FILLER_37_228 ();
 sg13g2_decap_8 FILLER_37_235 ();
 sg13g2_decap_8 FILLER_37_242 ();
 sg13g2_decap_8 FILLER_37_249 ();
 sg13g2_decap_8 FILLER_37_256 ();
 sg13g2_decap_8 FILLER_37_263 ();
 sg13g2_decap_4 FILLER_37_270 ();
 sg13g2_fill_2 FILLER_37_274 ();
 sg13g2_fill_2 FILLER_37_300 ();
 sg13g2_decap_4 FILLER_37_310 ();
 sg13g2_fill_2 FILLER_37_314 ();
 sg13g2_fill_1 FILLER_37_324 ();
 sg13g2_fill_1 FILLER_37_330 ();
 sg13g2_fill_1 FILLER_37_363 ();
 sg13g2_fill_1 FILLER_37_372 ();
 sg13g2_fill_2 FILLER_37_378 ();
 sg13g2_fill_1 FILLER_37_388 ();
 sg13g2_fill_2 FILLER_37_415 ();
 sg13g2_decap_8 FILLER_37_421 ();
 sg13g2_fill_2 FILLER_37_428 ();
 sg13g2_decap_8 FILLER_38_0 ();
 sg13g2_decap_8 FILLER_38_7 ();
 sg13g2_decap_8 FILLER_38_14 ();
 sg13g2_decap_8 FILLER_38_21 ();
 sg13g2_decap_8 FILLER_38_28 ();
 sg13g2_decap_8 FILLER_38_35 ();
 sg13g2_decap_8 FILLER_38_42 ();
 sg13g2_decap_8 FILLER_38_49 ();
 sg13g2_decap_8 FILLER_38_56 ();
 sg13g2_decap_8 FILLER_38_63 ();
 sg13g2_fill_2 FILLER_38_70 ();
 sg13g2_fill_1 FILLER_38_72 ();
 sg13g2_fill_2 FILLER_38_81 ();
 sg13g2_fill_1 FILLER_38_83 ();
 sg13g2_fill_1 FILLER_38_112 ();
 sg13g2_fill_2 FILLER_38_137 ();
 sg13g2_fill_1 FILLER_38_139 ();
 sg13g2_decap_8 FILLER_38_200 ();
 sg13g2_decap_8 FILLER_38_207 ();
 sg13g2_fill_2 FILLER_38_214 ();
 sg13g2_fill_1 FILLER_38_216 ();
 sg13g2_decap_8 FILLER_38_221 ();
 sg13g2_decap_4 FILLER_38_228 ();
 sg13g2_fill_1 FILLER_38_232 ();
 sg13g2_fill_2 FILLER_38_241 ();
 sg13g2_decap_4 FILLER_38_247 ();
 sg13g2_decap_8 FILLER_38_263 ();
 sg13g2_fill_1 FILLER_38_278 ();
 sg13g2_fill_1 FILLER_38_303 ();
 sg13g2_fill_2 FILLER_38_340 ();
 sg13g2_fill_1 FILLER_38_346 ();
 sg13g2_fill_1 FILLER_38_355 ();
 sg13g2_fill_1 FILLER_38_401 ();
 sg13g2_fill_1 FILLER_38_406 ();
 sg13g2_decap_8 FILLER_38_411 ();
 sg13g2_decap_8 FILLER_38_418 ();
 sg13g2_decap_4 FILLER_38_425 ();
 sg13g2_fill_1 FILLER_38_429 ();
endmodule
