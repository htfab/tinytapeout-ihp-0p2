module tt_um_toivoh_demo_deluxe (clk,
    ena,
    rst_n,
    ui_in,
    uio_in,
    uio_oe,
    uio_out,
    uo_out);
 input clk;
 input ena;
 input rst_n;
 input [7:0] ui_in;
 input [7:0] uio_in;
 output [7:0] uio_oe;
 output [7:0] uio_out;
 output [7:0] uo_out;

 wire _00000_;
 wire _00001_;
 wire _00002_;
 wire _00003_;
 wire _00004_;
 wire _00005_;
 wire _00006_;
 wire _00007_;
 wire _00008_;
 wire _00009_;
 wire _00010_;
 wire _00011_;
 wire _00012_;
 wire _00013_;
 wire _00014_;
 wire _00015_;
 wire _00016_;
 wire _00017_;
 wire _00018_;
 wire _00019_;
 wire _00020_;
 wire _00021_;
 wire _00022_;
 wire _00023_;
 wire _00024_;
 wire _00025_;
 wire _00026_;
 wire _00027_;
 wire _00028_;
 wire _00029_;
 wire _00030_;
 wire _00031_;
 wire _00032_;
 wire _00033_;
 wire _00034_;
 wire _00035_;
 wire _00036_;
 wire _00037_;
 wire _00038_;
 wire _00039_;
 wire _00040_;
 wire _00041_;
 wire _00042_;
 wire _00043_;
 wire _00044_;
 wire _00045_;
 wire _00046_;
 wire _00047_;
 wire _00048_;
 wire _00049_;
 wire _00050_;
 wire _00051_;
 wire _00052_;
 wire _00053_;
 wire _00054_;
 wire _00055_;
 wire _00056_;
 wire _00057_;
 wire _00058_;
 wire _00059_;
 wire _00060_;
 wire _00061_;
 wire _00062_;
 wire _00063_;
 wire _00064_;
 wire _00065_;
 wire _00066_;
 wire _00067_;
 wire _00068_;
 wire _00069_;
 wire _00070_;
 wire _00071_;
 wire _00072_;
 wire _00073_;
 wire _00074_;
 wire _00075_;
 wire _00076_;
 wire _00077_;
 wire _00078_;
 wire _00079_;
 wire _00080_;
 wire _00081_;
 wire _00082_;
 wire _00083_;
 wire _00084_;
 wire _00085_;
 wire _00086_;
 wire _00087_;
 wire _00088_;
 wire _00089_;
 wire _00090_;
 wire _00091_;
 wire _00092_;
 wire _00093_;
 wire _00094_;
 wire _00095_;
 wire _00096_;
 wire _00097_;
 wire _00098_;
 wire _00099_;
 wire _00100_;
 wire _00101_;
 wire _00102_;
 wire _00103_;
 wire _00104_;
 wire _00105_;
 wire _00106_;
 wire _00107_;
 wire _00108_;
 wire _00109_;
 wire _00110_;
 wire _00111_;
 wire _00112_;
 wire _00113_;
 wire _00114_;
 wire _00115_;
 wire _00116_;
 wire _00117_;
 wire _00118_;
 wire _00119_;
 wire _00120_;
 wire _00121_;
 wire _00122_;
 wire _00123_;
 wire _00124_;
 wire _00125_;
 wire _00126_;
 wire _00127_;
 wire _00128_;
 wire _00129_;
 wire _00130_;
 wire _00131_;
 wire _00132_;
 wire _00133_;
 wire _00134_;
 wire _00135_;
 wire _00136_;
 wire _00137_;
 wire _00138_;
 wire _00139_;
 wire _00140_;
 wire _00141_;
 wire _00142_;
 wire _00143_;
 wire _00144_;
 wire _00145_;
 wire _00146_;
 wire _00147_;
 wire _00148_;
 wire _00149_;
 wire _00150_;
 wire _00151_;
 wire _00152_;
 wire _00153_;
 wire _00154_;
 wire _00155_;
 wire _00156_;
 wire _00157_;
 wire _00158_;
 wire _00159_;
 wire _00160_;
 wire _00161_;
 wire _00162_;
 wire _00163_;
 wire _00164_;
 wire _00165_;
 wire _00166_;
 wire _00167_;
 wire _00168_;
 wire _00169_;
 wire _00170_;
 wire _00171_;
 wire _00172_;
 wire _00173_;
 wire _00174_;
 wire _00175_;
 wire _00176_;
 wire _00177_;
 wire _00178_;
 wire _00179_;
 wire _00180_;
 wire _00181_;
 wire _00182_;
 wire _00183_;
 wire _00184_;
 wire _00185_;
 wire _00186_;
 wire _00187_;
 wire _00188_;
 wire _00189_;
 wire _00190_;
 wire _00191_;
 wire _00192_;
 wire _00193_;
 wire _00194_;
 wire _00195_;
 wire _00196_;
 wire _00197_;
 wire _00198_;
 wire _00199_;
 wire _00200_;
 wire _00201_;
 wire _00202_;
 wire _00203_;
 wire _00204_;
 wire _00205_;
 wire _00206_;
 wire _00207_;
 wire _00208_;
 wire _00209_;
 wire _00210_;
 wire _00211_;
 wire _00212_;
 wire _00213_;
 wire _00214_;
 wire _00215_;
 wire _00216_;
 wire _00217_;
 wire _00218_;
 wire _00219_;
 wire _00220_;
 wire _00221_;
 wire _00222_;
 wire _00223_;
 wire _00224_;
 wire _00225_;
 wire _00226_;
 wire _00227_;
 wire _00228_;
 wire _00229_;
 wire _00230_;
 wire _00231_;
 wire _00232_;
 wire _00233_;
 wire _00234_;
 wire _00235_;
 wire _00236_;
 wire _00237_;
 wire _00238_;
 wire _00239_;
 wire _00240_;
 wire _00241_;
 wire _00242_;
 wire _00243_;
 wire _00244_;
 wire _00245_;
 wire _00246_;
 wire _00247_;
 wire _00248_;
 wire _00249_;
 wire _00250_;
 wire _00251_;
 wire _00252_;
 wire _00253_;
 wire _00254_;
 wire _00255_;
 wire _00256_;
 wire _00257_;
 wire _00258_;
 wire _00259_;
 wire _00260_;
 wire _00261_;
 wire _00262_;
 wire _00263_;
 wire _00264_;
 wire _00265_;
 wire _00266_;
 wire _00267_;
 wire _00268_;
 wire _00269_;
 wire _00270_;
 wire _00271_;
 wire _00272_;
 wire _00273_;
 wire _00274_;
 wire _00275_;
 wire _00276_;
 wire _00277_;
 wire _00278_;
 wire _00279_;
 wire _00280_;
 wire _00281_;
 wire _00282_;
 wire _00283_;
 wire _00284_;
 wire _00285_;
 wire _00286_;
 wire _00287_;
 wire _00288_;
 wire _00289_;
 wire _00290_;
 wire _00291_;
 wire _00292_;
 wire _00293_;
 wire _00294_;
 wire _00295_;
 wire _00296_;
 wire _00297_;
 wire _00298_;
 wire _00299_;
 wire _00300_;
 wire _00301_;
 wire _00302_;
 wire _00303_;
 wire _00304_;
 wire _00305_;
 wire _00306_;
 wire _00307_;
 wire _00308_;
 wire _00309_;
 wire _00310_;
 wire _00311_;
 wire _00312_;
 wire _00313_;
 wire _00314_;
 wire _00315_;
 wire _00316_;
 wire _00317_;
 wire _00318_;
 wire _00319_;
 wire _00320_;
 wire _00321_;
 wire _00322_;
 wire _00323_;
 wire _00324_;
 wire _00325_;
 wire _00326_;
 wire _00327_;
 wire _00328_;
 wire _00329_;
 wire _00330_;
 wire _00331_;
 wire _00332_;
 wire _00333_;
 wire _00334_;
 wire _00335_;
 wire _00336_;
 wire _00337_;
 wire _00338_;
 wire _00339_;
 wire _00340_;
 wire _00341_;
 wire _00342_;
 wire _00343_;
 wire _00344_;
 wire _00345_;
 wire _00346_;
 wire _00347_;
 wire _00348_;
 wire _00349_;
 wire _00350_;
 wire _00351_;
 wire _00352_;
 wire _00353_;
 wire _00354_;
 wire _00355_;
 wire _00356_;
 wire _00357_;
 wire _00358_;
 wire _00359_;
 wire _00360_;
 wire _00361_;
 wire _00362_;
 wire _00363_;
 wire _00364_;
 wire _00365_;
 wire _00366_;
 wire _00367_;
 wire _00368_;
 wire _00369_;
 wire _00370_;
 wire _00371_;
 wire _00372_;
 wire _00373_;
 wire _00374_;
 wire _00375_;
 wire _00376_;
 wire _00377_;
 wire _00378_;
 wire _00379_;
 wire _00380_;
 wire _00381_;
 wire _00382_;
 wire _00383_;
 wire _00384_;
 wire _00385_;
 wire _00386_;
 wire _00387_;
 wire _00388_;
 wire _00389_;
 wire _00390_;
 wire _00391_;
 wire _00392_;
 wire _00393_;
 wire _00394_;
 wire _00395_;
 wire _00396_;
 wire _00397_;
 wire _00398_;
 wire _00399_;
 wire _00400_;
 wire _00401_;
 wire _00402_;
 wire _00403_;
 wire _00404_;
 wire _00405_;
 wire _00406_;
 wire _00407_;
 wire _00408_;
 wire _00409_;
 wire _00410_;
 wire _00411_;
 wire _00412_;
 wire _00413_;
 wire _00414_;
 wire _00415_;
 wire _00416_;
 wire _00417_;
 wire _00418_;
 wire _00419_;
 wire _00420_;
 wire _00421_;
 wire _00422_;
 wire _00423_;
 wire _00424_;
 wire _00425_;
 wire _00426_;
 wire _00427_;
 wire _00428_;
 wire _00429_;
 wire _00430_;
 wire _00431_;
 wire _00432_;
 wire _00433_;
 wire _00434_;
 wire _00435_;
 wire _00436_;
 wire _00437_;
 wire _00438_;
 wire _00439_;
 wire _00440_;
 wire _00441_;
 wire _00442_;
 wire _00443_;
 wire _00444_;
 wire _00445_;
 wire _00446_;
 wire _00447_;
 wire _00448_;
 wire _00449_;
 wire _00450_;
 wire _00451_;
 wire _00452_;
 wire _00453_;
 wire _00454_;
 wire _00455_;
 wire _00456_;
 wire _00457_;
 wire _00458_;
 wire _00459_;
 wire _00460_;
 wire _00461_;
 wire _00462_;
 wire _00463_;
 wire _00464_;
 wire _00465_;
 wire _00466_;
 wire _00467_;
 wire _00468_;
 wire _00469_;
 wire _00470_;
 wire _00471_;
 wire _00472_;
 wire _00473_;
 wire _00474_;
 wire _00475_;
 wire _00476_;
 wire _00477_;
 wire _00478_;
 wire _00479_;
 wire _00480_;
 wire _00481_;
 wire _00482_;
 wire _00483_;
 wire _00484_;
 wire _00485_;
 wire _00486_;
 wire _00487_;
 wire _00488_;
 wire _00489_;
 wire _00490_;
 wire _00491_;
 wire _00492_;
 wire _00493_;
 wire _00494_;
 wire _00495_;
 wire _00496_;
 wire _00497_;
 wire _00498_;
 wire _00499_;
 wire _00500_;
 wire _00501_;
 wire _00502_;
 wire _00503_;
 wire _00504_;
 wire _00505_;
 wire _00506_;
 wire _00507_;
 wire _00508_;
 wire _00509_;
 wire _00510_;
 wire _00511_;
 wire _00512_;
 wire _00513_;
 wire _00514_;
 wire _00515_;
 wire _00516_;
 wire _00517_;
 wire _00518_;
 wire _00519_;
 wire _00520_;
 wire _00521_;
 wire _00522_;
 wire _00523_;
 wire _00524_;
 wire _00525_;
 wire _00526_;
 wire _00527_;
 wire _00528_;
 wire _00529_;
 wire _00530_;
 wire _00531_;
 wire _00532_;
 wire _00533_;
 wire _00534_;
 wire _00535_;
 wire _00536_;
 wire _00537_;
 wire _00538_;
 wire _00539_;
 wire _00540_;
 wire _00541_;
 wire _00542_;
 wire _00543_;
 wire _00544_;
 wire _00545_;
 wire _00546_;
 wire _00547_;
 wire _00548_;
 wire _00549_;
 wire _00550_;
 wire _00551_;
 wire _00552_;
 wire _00553_;
 wire _00554_;
 wire _00555_;
 wire _00556_;
 wire _00557_;
 wire _00558_;
 wire _00559_;
 wire _00560_;
 wire _00561_;
 wire _00562_;
 wire _00563_;
 wire _00564_;
 wire _00565_;
 wire _00566_;
 wire _00567_;
 wire _00568_;
 wire _00569_;
 wire _00570_;
 wire _00571_;
 wire _00572_;
 wire _00573_;
 wire _00574_;
 wire _00575_;
 wire _00576_;
 wire _00577_;
 wire _00578_;
 wire _00579_;
 wire _00580_;
 wire _00581_;
 wire _00582_;
 wire _00583_;
 wire _00584_;
 wire _00585_;
 wire _00586_;
 wire _00587_;
 wire _00588_;
 wire _00589_;
 wire _00590_;
 wire _00591_;
 wire _00592_;
 wire _00593_;
 wire _00594_;
 wire _00595_;
 wire _00596_;
 wire _00597_;
 wire _00598_;
 wire _00599_;
 wire _00600_;
 wire _00601_;
 wire _00602_;
 wire _00603_;
 wire _00604_;
 wire _00605_;
 wire _00606_;
 wire _00607_;
 wire _00608_;
 wire _00609_;
 wire _00610_;
 wire _00611_;
 wire _00612_;
 wire _00613_;
 wire _00614_;
 wire _00615_;
 wire _00616_;
 wire _00617_;
 wire _00618_;
 wire _00619_;
 wire _00620_;
 wire _00621_;
 wire _00622_;
 wire _00623_;
 wire _00624_;
 wire _00625_;
 wire _00626_;
 wire _00627_;
 wire _00628_;
 wire _00629_;
 wire _00630_;
 wire _00631_;
 wire _00632_;
 wire _00633_;
 wire _00634_;
 wire _00635_;
 wire _00636_;
 wire _00637_;
 wire _00638_;
 wire _00639_;
 wire _00640_;
 wire _00641_;
 wire _00642_;
 wire _00643_;
 wire _00644_;
 wire _00645_;
 wire _00646_;
 wire _00647_;
 wire _00648_;
 wire _00649_;
 wire _00650_;
 wire _00651_;
 wire _00652_;
 wire _00653_;
 wire _00654_;
 wire _00655_;
 wire _00656_;
 wire _00657_;
 wire _00658_;
 wire _00659_;
 wire _00660_;
 wire _00661_;
 wire _00662_;
 wire _00663_;
 wire _00664_;
 wire _00665_;
 wire _00666_;
 wire _00667_;
 wire _00668_;
 wire _00669_;
 wire _00670_;
 wire _00671_;
 wire _00672_;
 wire _00673_;
 wire _00674_;
 wire _00675_;
 wire _00676_;
 wire _00677_;
 wire _00678_;
 wire _00679_;
 wire _00680_;
 wire _00681_;
 wire _00682_;
 wire _00683_;
 wire _00684_;
 wire _00685_;
 wire _00686_;
 wire _00687_;
 wire _00688_;
 wire _00689_;
 wire _00690_;
 wire _00691_;
 wire _00692_;
 wire _00693_;
 wire _00694_;
 wire _00695_;
 wire _00696_;
 wire _00697_;
 wire _00698_;
 wire _00699_;
 wire _00700_;
 wire _00701_;
 wire _00702_;
 wire _00703_;
 wire _00704_;
 wire _00705_;
 wire _00706_;
 wire _00707_;
 wire _00708_;
 wire _00709_;
 wire _00710_;
 wire _00711_;
 wire _00712_;
 wire _00713_;
 wire _00714_;
 wire _00715_;
 wire _00716_;
 wire _00717_;
 wire _00718_;
 wire _00719_;
 wire _00720_;
 wire _00721_;
 wire _00722_;
 wire _00723_;
 wire _00724_;
 wire _00725_;
 wire _00726_;
 wire _00727_;
 wire _00728_;
 wire _00729_;
 wire _00730_;
 wire _00731_;
 wire _00732_;
 wire _00733_;
 wire _00734_;
 wire _00735_;
 wire _00736_;
 wire _00737_;
 wire _00738_;
 wire _00739_;
 wire _00740_;
 wire _00741_;
 wire _00742_;
 wire _00743_;
 wire _00744_;
 wire _00745_;
 wire _00746_;
 wire _00747_;
 wire _00748_;
 wire _00749_;
 wire _00750_;
 wire _00751_;
 wire _00752_;
 wire _00753_;
 wire _00754_;
 wire _00755_;
 wire _00756_;
 wire _00757_;
 wire _00758_;
 wire _00759_;
 wire _00760_;
 wire _00761_;
 wire _00762_;
 wire _00763_;
 wire _00764_;
 wire _00765_;
 wire _00766_;
 wire _00767_;
 wire _00768_;
 wire _00769_;
 wire _00770_;
 wire _00771_;
 wire _00772_;
 wire _00773_;
 wire _00774_;
 wire _00775_;
 wire _00776_;
 wire _00777_;
 wire _00778_;
 wire _00779_;
 wire _00780_;
 wire _00781_;
 wire _00782_;
 wire _00783_;
 wire _00784_;
 wire _00785_;
 wire _00786_;
 wire _00787_;
 wire _00788_;
 wire _00789_;
 wire _00790_;
 wire _00791_;
 wire _00792_;
 wire _00793_;
 wire _00794_;
 wire _00795_;
 wire _00796_;
 wire _00797_;
 wire _00798_;
 wire _00799_;
 wire _00800_;
 wire _00801_;
 wire _00802_;
 wire _00803_;
 wire _00804_;
 wire _00805_;
 wire _00806_;
 wire _00807_;
 wire _00808_;
 wire _00809_;
 wire _00810_;
 wire _00811_;
 wire _00812_;
 wire _00813_;
 wire _00814_;
 wire _00815_;
 wire _00816_;
 wire _00817_;
 wire _00818_;
 wire _00819_;
 wire _00820_;
 wire _00821_;
 wire _00822_;
 wire _00823_;
 wire _00824_;
 wire _00825_;
 wire _00826_;
 wire _00827_;
 wire _00828_;
 wire _00829_;
 wire _00830_;
 wire _00831_;
 wire _00832_;
 wire _00833_;
 wire _00834_;
 wire _00835_;
 wire _00836_;
 wire _00837_;
 wire _00838_;
 wire _00839_;
 wire _00840_;
 wire _00841_;
 wire _00842_;
 wire _00843_;
 wire _00844_;
 wire _00845_;
 wire _00846_;
 wire _00847_;
 wire _00848_;
 wire _00849_;
 wire _00850_;
 wire _00851_;
 wire _00852_;
 wire _00853_;
 wire _00854_;
 wire _00855_;
 wire _00856_;
 wire _00857_;
 wire _00858_;
 wire _00859_;
 wire _00860_;
 wire _00861_;
 wire _00862_;
 wire _00863_;
 wire _00864_;
 wire _00865_;
 wire _00866_;
 wire _00867_;
 wire _00868_;
 wire _00869_;
 wire _00870_;
 wire _00871_;
 wire _00872_;
 wire _00873_;
 wire _00874_;
 wire _00875_;
 wire _00876_;
 wire _00877_;
 wire _00878_;
 wire _00879_;
 wire _00880_;
 wire _00881_;
 wire _00882_;
 wire _00883_;
 wire _00884_;
 wire _00885_;
 wire _00886_;
 wire _00887_;
 wire _00888_;
 wire _00889_;
 wire _00890_;
 wire _00891_;
 wire _00892_;
 wire _00893_;
 wire _00894_;
 wire _00895_;
 wire _00896_;
 wire _00897_;
 wire _00898_;
 wire _00899_;
 wire _00900_;
 wire _00901_;
 wire _00902_;
 wire _00903_;
 wire _00904_;
 wire _00905_;
 wire _00906_;
 wire _00907_;
 wire _00908_;
 wire _00909_;
 wire _00910_;
 wire _00911_;
 wire _00912_;
 wire _00913_;
 wire _00914_;
 wire _00915_;
 wire _00916_;
 wire _00917_;
 wire _00918_;
 wire _00919_;
 wire _00920_;
 wire _00921_;
 wire _00922_;
 wire _00923_;
 wire _00924_;
 wire _00925_;
 wire _00926_;
 wire _00927_;
 wire _00928_;
 wire _00929_;
 wire _00930_;
 wire _00931_;
 wire _00932_;
 wire _00933_;
 wire _00934_;
 wire _00935_;
 wire _00936_;
 wire _00937_;
 wire _00938_;
 wire _00939_;
 wire _00940_;
 wire _00941_;
 wire _00942_;
 wire _00943_;
 wire _00944_;
 wire _00945_;
 wire _00946_;
 wire _00947_;
 wire _00948_;
 wire _00949_;
 wire _00950_;
 wire _00951_;
 wire _00952_;
 wire _00953_;
 wire _00954_;
 wire _00955_;
 wire _00956_;
 wire _00957_;
 wire _00958_;
 wire _00959_;
 wire _00960_;
 wire _00961_;
 wire _00962_;
 wire _00963_;
 wire _00964_;
 wire _00965_;
 wire _00966_;
 wire _00967_;
 wire _00968_;
 wire _00969_;
 wire _00970_;
 wire _00971_;
 wire _00972_;
 wire _00973_;
 wire _00974_;
 wire _00975_;
 wire _00976_;
 wire _00977_;
 wire _00978_;
 wire _00979_;
 wire _00980_;
 wire _00981_;
 wire _00982_;
 wire _00983_;
 wire _00984_;
 wire _00985_;
 wire _00986_;
 wire _00987_;
 wire _00988_;
 wire _00989_;
 wire _00990_;
 wire _00991_;
 wire _00992_;
 wire _00993_;
 wire _00994_;
 wire _00995_;
 wire _00996_;
 wire _00997_;
 wire _00998_;
 wire _00999_;
 wire _01000_;
 wire _01001_;
 wire _01002_;
 wire _01003_;
 wire _01004_;
 wire _01005_;
 wire _01006_;
 wire _01007_;
 wire _01008_;
 wire _01009_;
 wire _01010_;
 wire _01011_;
 wire _01012_;
 wire _01013_;
 wire _01014_;
 wire _01015_;
 wire _01016_;
 wire _01017_;
 wire _01018_;
 wire _01019_;
 wire _01020_;
 wire _01021_;
 wire _01022_;
 wire _01023_;
 wire _01024_;
 wire _01025_;
 wire _01026_;
 wire _01027_;
 wire _01028_;
 wire _01029_;
 wire _01030_;
 wire _01031_;
 wire _01032_;
 wire _01033_;
 wire _01034_;
 wire _01035_;
 wire _01036_;
 wire _01037_;
 wire _01038_;
 wire _01039_;
 wire _01040_;
 wire _01041_;
 wire _01042_;
 wire _01043_;
 wire _01044_;
 wire _01045_;
 wire _01046_;
 wire _01047_;
 wire _01048_;
 wire _01049_;
 wire _01050_;
 wire _01051_;
 wire _01052_;
 wire _01053_;
 wire _01054_;
 wire _01055_;
 wire _01056_;
 wire _01057_;
 wire _01058_;
 wire _01059_;
 wire _01060_;
 wire _01061_;
 wire _01062_;
 wire _01063_;
 wire _01064_;
 wire _01065_;
 wire _01066_;
 wire _01067_;
 wire _01068_;
 wire _01069_;
 wire _01070_;
 wire _01071_;
 wire _01072_;
 wire _01073_;
 wire _01074_;
 wire _01075_;
 wire _01076_;
 wire _01077_;
 wire _01078_;
 wire _01079_;
 wire _01080_;
 wire _01081_;
 wire _01082_;
 wire _01083_;
 wire _01084_;
 wire _01085_;
 wire _01086_;
 wire _01087_;
 wire _01088_;
 wire _01089_;
 wire _01090_;
 wire _01091_;
 wire _01092_;
 wire _01093_;
 wire _01094_;
 wire _01095_;
 wire _01096_;
 wire _01097_;
 wire _01098_;
 wire _01099_;
 wire _01100_;
 wire _01101_;
 wire _01102_;
 wire _01103_;
 wire _01104_;
 wire _01105_;
 wire _01106_;
 wire _01107_;
 wire _01108_;
 wire _01109_;
 wire _01110_;
 wire _01111_;
 wire _01112_;
 wire _01113_;
 wire _01114_;
 wire _01115_;
 wire _01116_;
 wire _01117_;
 wire _01118_;
 wire _01119_;
 wire _01120_;
 wire _01121_;
 wire _01122_;
 wire _01123_;
 wire _01124_;
 wire _01125_;
 wire _01126_;
 wire _01127_;
 wire _01128_;
 wire _01129_;
 wire _01130_;
 wire _01131_;
 wire _01132_;
 wire _01133_;
 wire _01134_;
 wire _01135_;
 wire _01136_;
 wire _01137_;
 wire _01138_;
 wire _01139_;
 wire _01140_;
 wire _01141_;
 wire _01142_;
 wire _01143_;
 wire _01144_;
 wire _01145_;
 wire _01146_;
 wire _01147_;
 wire _01148_;
 wire _01149_;
 wire _01150_;
 wire _01151_;
 wire _01152_;
 wire _01153_;
 wire _01154_;
 wire _01155_;
 wire _01156_;
 wire _01157_;
 wire _01158_;
 wire _01159_;
 wire _01160_;
 wire _01161_;
 wire _01162_;
 wire _01163_;
 wire _01164_;
 wire _01165_;
 wire _01166_;
 wire _01167_;
 wire _01168_;
 wire _01169_;
 wire _01170_;
 wire _01171_;
 wire _01172_;
 wire _01173_;
 wire _01174_;
 wire _01175_;
 wire _01176_;
 wire _01177_;
 wire _01178_;
 wire _01179_;
 wire _01180_;
 wire _01181_;
 wire _01182_;
 wire _01183_;
 wire _01184_;
 wire _01185_;
 wire _01186_;
 wire _01187_;
 wire _01188_;
 wire _01189_;
 wire _01190_;
 wire _01191_;
 wire _01192_;
 wire _01193_;
 wire _01194_;
 wire _01195_;
 wire _01196_;
 wire _01197_;
 wire _01198_;
 wire _01199_;
 wire _01200_;
 wire _01201_;
 wire _01202_;
 wire _01203_;
 wire _01204_;
 wire _01205_;
 wire _01206_;
 wire _01207_;
 wire _01208_;
 wire _01209_;
 wire _01210_;
 wire _01211_;
 wire _01212_;
 wire _01213_;
 wire _01214_;
 wire _01215_;
 wire _01216_;
 wire _01217_;
 wire _01218_;
 wire _01219_;
 wire _01220_;
 wire _01221_;
 wire _01222_;
 wire _01223_;
 wire _01224_;
 wire _01225_;
 wire _01226_;
 wire _01227_;
 wire _01228_;
 wire _01229_;
 wire _01230_;
 wire _01231_;
 wire _01232_;
 wire _01233_;
 wire _01234_;
 wire _01235_;
 wire _01236_;
 wire _01237_;
 wire _01238_;
 wire _01239_;
 wire _01240_;
 wire _01241_;
 wire _01242_;
 wire _01243_;
 wire _01244_;
 wire _01245_;
 wire _01246_;
 wire _01247_;
 wire _01248_;
 wire _01249_;
 wire _01250_;
 wire _01251_;
 wire _01252_;
 wire _01253_;
 wire _01254_;
 wire _01255_;
 wire _01256_;
 wire _01257_;
 wire _01258_;
 wire _01259_;
 wire _01260_;
 wire _01261_;
 wire _01262_;
 wire _01263_;
 wire _01264_;
 wire _01265_;
 wire _01266_;
 wire _01267_;
 wire _01268_;
 wire _01269_;
 wire _01270_;
 wire _01271_;
 wire _01272_;
 wire _01273_;
 wire _01274_;
 wire _01275_;
 wire _01276_;
 wire _01277_;
 wire _01278_;
 wire _01279_;
 wire _01280_;
 wire _01281_;
 wire _01282_;
 wire _01283_;
 wire _01284_;
 wire _01285_;
 wire _01286_;
 wire _01287_;
 wire _01288_;
 wire _01289_;
 wire _01290_;
 wire _01291_;
 wire _01292_;
 wire _01293_;
 wire _01294_;
 wire _01295_;
 wire _01296_;
 wire _01297_;
 wire _01298_;
 wire _01299_;
 wire _01300_;
 wire _01301_;
 wire _01302_;
 wire _01303_;
 wire _01304_;
 wire _01305_;
 wire _01306_;
 wire _01307_;
 wire _01308_;
 wire _01309_;
 wire _01310_;
 wire _01311_;
 wire _01312_;
 wire _01313_;
 wire _01314_;
 wire _01315_;
 wire _01316_;
 wire _01317_;
 wire _01318_;
 wire _01319_;
 wire _01320_;
 wire _01321_;
 wire _01322_;
 wire _01323_;
 wire _01324_;
 wire _01325_;
 wire _01326_;
 wire _01327_;
 wire _01328_;
 wire _01329_;
 wire _01330_;
 wire _01331_;
 wire _01332_;
 wire _01333_;
 wire _01334_;
 wire _01335_;
 wire _01336_;
 wire _01337_;
 wire _01338_;
 wire _01339_;
 wire _01340_;
 wire _01341_;
 wire _01342_;
 wire _01343_;
 wire _01344_;
 wire _01345_;
 wire _01346_;
 wire _01347_;
 wire _01348_;
 wire _01349_;
 wire _01350_;
 wire _01351_;
 wire _01352_;
 wire _01353_;
 wire _01354_;
 wire _01355_;
 wire _01356_;
 wire _01357_;
 wire _01358_;
 wire _01359_;
 wire _01360_;
 wire _01361_;
 wire _01362_;
 wire _01363_;
 wire _01364_;
 wire _01365_;
 wire _01366_;
 wire _01367_;
 wire _01368_;
 wire _01369_;
 wire _01370_;
 wire _01371_;
 wire _01372_;
 wire _01373_;
 wire _01374_;
 wire _01375_;
 wire _01376_;
 wire _01377_;
 wire _01378_;
 wire _01379_;
 wire _01380_;
 wire _01381_;
 wire _01382_;
 wire _01383_;
 wire _01384_;
 wire _01385_;
 wire _01386_;
 wire _01387_;
 wire _01388_;
 wire _01389_;
 wire _01390_;
 wire _01391_;
 wire _01392_;
 wire _01393_;
 wire _01394_;
 wire _01395_;
 wire _01396_;
 wire _01397_;
 wire _01398_;
 wire _01399_;
 wire _01400_;
 wire _01401_;
 wire _01402_;
 wire _01403_;
 wire _01404_;
 wire _01405_;
 wire _01406_;
 wire _01407_;
 wire _01408_;
 wire _01409_;
 wire _01410_;
 wire _01411_;
 wire _01412_;
 wire _01413_;
 wire _01414_;
 wire _01415_;
 wire _01416_;
 wire _01417_;
 wire _01418_;
 wire _01419_;
 wire _01420_;
 wire _01421_;
 wire _01422_;
 wire _01423_;
 wire _01424_;
 wire _01425_;
 wire _01426_;
 wire _01427_;
 wire _01428_;
 wire _01429_;
 wire _01430_;
 wire _01431_;
 wire _01432_;
 wire _01433_;
 wire _01434_;
 wire _01435_;
 wire _01436_;
 wire _01437_;
 wire _01438_;
 wire _01439_;
 wire _01440_;
 wire _01441_;
 wire _01442_;
 wire _01443_;
 wire _01444_;
 wire _01445_;
 wire _01446_;
 wire _01447_;
 wire _01448_;
 wire _01449_;
 wire _01450_;
 wire _01451_;
 wire _01452_;
 wire _01453_;
 wire _01454_;
 wire _01455_;
 wire _01456_;
 wire _01457_;
 wire _01458_;
 wire _01459_;
 wire _01460_;
 wire _01461_;
 wire _01462_;
 wire _01463_;
 wire _01464_;
 wire _01465_;
 wire _01466_;
 wire _01467_;
 wire _01468_;
 wire _01469_;
 wire _01470_;
 wire _01471_;
 wire _01472_;
 wire _01473_;
 wire _01474_;
 wire _01475_;
 wire _01476_;
 wire _01477_;
 wire _01478_;
 wire _01479_;
 wire _01480_;
 wire _01481_;
 wire _01482_;
 wire _01483_;
 wire _01484_;
 wire _01485_;
 wire _01486_;
 wire _01487_;
 wire _01488_;
 wire _01489_;
 wire _01490_;
 wire _01491_;
 wire _01492_;
 wire _01493_;
 wire _01494_;
 wire _01495_;
 wire _01496_;
 wire _01497_;
 wire _01498_;
 wire _01499_;
 wire _01500_;
 wire _01501_;
 wire _01502_;
 wire _01503_;
 wire _01504_;
 wire _01505_;
 wire _01506_;
 wire _01507_;
 wire _01508_;
 wire _01509_;
 wire _01510_;
 wire _01511_;
 wire _01512_;
 wire _01513_;
 wire _01514_;
 wire _01515_;
 wire _01516_;
 wire _01517_;
 wire _01518_;
 wire _01519_;
 wire _01520_;
 wire _01521_;
 wire _01522_;
 wire _01523_;
 wire _01524_;
 wire _01525_;
 wire _01526_;
 wire _01527_;
 wire _01528_;
 wire _01529_;
 wire _01530_;
 wire _01531_;
 wire _01532_;
 wire _01533_;
 wire _01534_;
 wire _01535_;
 wire _01536_;
 wire _01537_;
 wire _01538_;
 wire _01539_;
 wire _01540_;
 wire _01541_;
 wire _01542_;
 wire _01543_;
 wire _01544_;
 wire _01545_;
 wire _01546_;
 wire _01547_;
 wire _01548_;
 wire _01549_;
 wire _01550_;
 wire _01551_;
 wire _01552_;
 wire _01553_;
 wire _01554_;
 wire _01555_;
 wire _01556_;
 wire _01557_;
 wire _01558_;
 wire _01559_;
 wire _01560_;
 wire _01561_;
 wire _01562_;
 wire _01563_;
 wire _01564_;
 wire _01565_;
 wire _01566_;
 wire _01567_;
 wire _01568_;
 wire _01569_;
 wire _01570_;
 wire _01571_;
 wire _01572_;
 wire _01573_;
 wire _01574_;
 wire _01575_;
 wire _01576_;
 wire _01577_;
 wire _01578_;
 wire _01579_;
 wire _01580_;
 wire _01581_;
 wire _01582_;
 wire _01583_;
 wire _01584_;
 wire _01585_;
 wire _01586_;
 wire _01587_;
 wire _01588_;
 wire _01589_;
 wire _01590_;
 wire _01591_;
 wire _01592_;
 wire _01593_;
 wire _01594_;
 wire _01595_;
 wire _01596_;
 wire _01597_;
 wire _01598_;
 wire _01599_;
 wire _01600_;
 wire _01601_;
 wire _01602_;
 wire _01603_;
 wire _01604_;
 wire _01605_;
 wire _01606_;
 wire _01607_;
 wire _01608_;
 wire _01609_;
 wire _01610_;
 wire _01611_;
 wire _01612_;
 wire _01613_;
 wire _01614_;
 wire _01615_;
 wire _01616_;
 wire _01617_;
 wire _01618_;
 wire _01619_;
 wire _01620_;
 wire _01621_;
 wire _01622_;
 wire _01623_;
 wire _01624_;
 wire _01625_;
 wire _01626_;
 wire _01627_;
 wire _01628_;
 wire _01629_;
 wire _01630_;
 wire _01631_;
 wire _01632_;
 wire _01633_;
 wire _01634_;
 wire _01635_;
 wire _01636_;
 wire _01637_;
 wire _01638_;
 wire _01639_;
 wire _01640_;
 wire _01641_;
 wire _01642_;
 wire _01643_;
 wire _01644_;
 wire _01645_;
 wire _01646_;
 wire _01647_;
 wire _01648_;
 wire _01649_;
 wire _01650_;
 wire _01651_;
 wire _01652_;
 wire _01653_;
 wire _01654_;
 wire _01655_;
 wire _01656_;
 wire _01657_;
 wire _01658_;
 wire _01659_;
 wire _01660_;
 wire _01661_;
 wire _01662_;
 wire _01663_;
 wire _01664_;
 wire _01665_;
 wire _01666_;
 wire _01667_;
 wire _01668_;
 wire _01669_;
 wire _01670_;
 wire _01671_;
 wire _01672_;
 wire _01673_;
 wire _01674_;
 wire _01675_;
 wire _01676_;
 wire _01677_;
 wire _01678_;
 wire _01679_;
 wire _01680_;
 wire _01681_;
 wire _01682_;
 wire _01683_;
 wire _01684_;
 wire _01685_;
 wire _01686_;
 wire _01687_;
 wire _01688_;
 wire _01689_;
 wire _01690_;
 wire _01691_;
 wire _01692_;
 wire _01693_;
 wire _01694_;
 wire _01695_;
 wire _01696_;
 wire _01697_;
 wire _01698_;
 wire _01699_;
 wire _01700_;
 wire _01701_;
 wire _01702_;
 wire _01703_;
 wire _01704_;
 wire _01705_;
 wire _01706_;
 wire _01707_;
 wire _01708_;
 wire _01709_;
 wire _01710_;
 wire _01711_;
 wire _01712_;
 wire _01713_;
 wire _01714_;
 wire _01715_;
 wire _01716_;
 wire _01717_;
 wire _01718_;
 wire _01719_;
 wire _01720_;
 wire _01721_;
 wire _01722_;
 wire _01723_;
 wire _01724_;
 wire _01725_;
 wire _01726_;
 wire _01727_;
 wire _01728_;
 wire _01729_;
 wire _01730_;
 wire _01731_;
 wire _01732_;
 wire _01733_;
 wire _01734_;
 wire _01735_;
 wire _01736_;
 wire _01737_;
 wire _01738_;
 wire _01739_;
 wire _01740_;
 wire _01741_;
 wire _01742_;
 wire _01743_;
 wire _01744_;
 wire _01745_;
 wire _01746_;
 wire _01747_;
 wire _01748_;
 wire _01749_;
 wire _01750_;
 wire _01751_;
 wire _01752_;
 wire _01753_;
 wire _01754_;
 wire _01755_;
 wire _01756_;
 wire _01757_;
 wire _01758_;
 wire _01759_;
 wire _01760_;
 wire _01761_;
 wire _01762_;
 wire _01763_;
 wire _01764_;
 wire _01765_;
 wire _01766_;
 wire _01767_;
 wire _01768_;
 wire _01769_;
 wire _01770_;
 wire _01771_;
 wire _01772_;
 wire _01773_;
 wire _01774_;
 wire _01775_;
 wire _01776_;
 wire _01777_;
 wire _01778_;
 wire _01779_;
 wire _01780_;
 wire _01781_;
 wire _01782_;
 wire _01783_;
 wire _01784_;
 wire _01785_;
 wire _01786_;
 wire _01787_;
 wire _01788_;
 wire _01789_;
 wire _01790_;
 wire _01791_;
 wire _01792_;
 wire _01793_;
 wire _01794_;
 wire _01795_;
 wire _01796_;
 wire _01797_;
 wire _01798_;
 wire _01799_;
 wire _01800_;
 wire _01801_;
 wire _01802_;
 wire _01803_;
 wire _01804_;
 wire _01805_;
 wire _01806_;
 wire _01807_;
 wire _01808_;
 wire _01809_;
 wire _01810_;
 wire _01811_;
 wire _01812_;
 wire _01813_;
 wire _01814_;
 wire _01815_;
 wire _01816_;
 wire _01817_;
 wire _01818_;
 wire _01819_;
 wire _01820_;
 wire _01821_;
 wire _01822_;
 wire _01823_;
 wire _01824_;
 wire _01825_;
 wire _01826_;
 wire _01827_;
 wire _01828_;
 wire _01829_;
 wire _01830_;
 wire _01831_;
 wire _01832_;
 wire _01833_;
 wire _01834_;
 wire _01835_;
 wire _01836_;
 wire _01837_;
 wire _01838_;
 wire _01839_;
 wire _01840_;
 wire _01841_;
 wire _01842_;
 wire _01843_;
 wire _01844_;
 wire _01845_;
 wire _01846_;
 wire _01847_;
 wire _01848_;
 wire _01849_;
 wire _01850_;
 wire _01851_;
 wire _01852_;
 wire _01853_;
 wire _01854_;
 wire _01855_;
 wire _01856_;
 wire _01857_;
 wire _01858_;
 wire _01859_;
 wire _01860_;
 wire _01861_;
 wire _01862_;
 wire _01863_;
 wire _01864_;
 wire _01865_;
 wire _01866_;
 wire _01867_;
 wire _01868_;
 wire _01869_;
 wire _01870_;
 wire _01871_;
 wire _01872_;
 wire _01873_;
 wire _01874_;
 wire _01875_;
 wire _01876_;
 wire _01877_;
 wire _01878_;
 wire _01879_;
 wire _01880_;
 wire _01881_;
 wire _01882_;
 wire _01883_;
 wire _01884_;
 wire _01885_;
 wire _01886_;
 wire _01887_;
 wire _01888_;
 wire _01889_;
 wire _01890_;
 wire _01891_;
 wire _01892_;
 wire _01893_;
 wire _01894_;
 wire _01895_;
 wire _01896_;
 wire _01897_;
 wire _01898_;
 wire _01899_;
 wire _01900_;
 wire _01901_;
 wire _01902_;
 wire _01903_;
 wire _01904_;
 wire _01905_;
 wire _01906_;
 wire _01907_;
 wire _01908_;
 wire _01909_;
 wire _01910_;
 wire _01911_;
 wire _01912_;
 wire _01913_;
 wire _01914_;
 wire _01915_;
 wire _01916_;
 wire _01917_;
 wire _01918_;
 wire _01919_;
 wire _01920_;
 wire _01921_;
 wire _01922_;
 wire _01923_;
 wire _01924_;
 wire _01925_;
 wire _01926_;
 wire _01927_;
 wire _01928_;
 wire _01929_;
 wire _01930_;
 wire _01931_;
 wire _01932_;
 wire _01933_;
 wire _01934_;
 wire _01935_;
 wire _01936_;
 wire _01937_;
 wire _01938_;
 wire _01939_;
 wire _01940_;
 wire _01941_;
 wire _01942_;
 wire _01943_;
 wire _01944_;
 wire _01945_;
 wire _01946_;
 wire _01947_;
 wire _01948_;
 wire _01949_;
 wire _01950_;
 wire _01951_;
 wire _01952_;
 wire _01953_;
 wire _01954_;
 wire _01955_;
 wire _01956_;
 wire _01957_;
 wire _01958_;
 wire _01959_;
 wire _01960_;
 wire _01961_;
 wire _01962_;
 wire _01963_;
 wire _01964_;
 wire _01965_;
 wire _01966_;
 wire _01967_;
 wire _01968_;
 wire _01969_;
 wire _01970_;
 wire _01971_;
 wire _01972_;
 wire _01973_;
 wire _01974_;
 wire _01975_;
 wire _01976_;
 wire _01977_;
 wire _01978_;
 wire _01979_;
 wire _01980_;
 wire _01981_;
 wire _01982_;
 wire _01983_;
 wire _01984_;
 wire _01985_;
 wire _01986_;
 wire _01987_;
 wire _01988_;
 wire _01989_;
 wire _01990_;
 wire _01991_;
 wire _01992_;
 wire _01993_;
 wire _01994_;
 wire _01995_;
 wire _01996_;
 wire _01997_;
 wire _01998_;
 wire _01999_;
 wire _02000_;
 wire _02001_;
 wire _02002_;
 wire _02003_;
 wire _02004_;
 wire _02005_;
 wire _02006_;
 wire _02007_;
 wire _02008_;
 wire _02009_;
 wire _02010_;
 wire _02011_;
 wire _02012_;
 wire _02013_;
 wire _02014_;
 wire _02015_;
 wire _02016_;
 wire _02017_;
 wire _02018_;
 wire _02019_;
 wire _02020_;
 wire _02021_;
 wire _02022_;
 wire _02023_;
 wire _02024_;
 wire _02025_;
 wire _02026_;
 wire _02027_;
 wire _02028_;
 wire _02029_;
 wire _02030_;
 wire _02031_;
 wire _02032_;
 wire _02033_;
 wire _02034_;
 wire _02035_;
 wire _02036_;
 wire _02037_;
 wire _02038_;
 wire _02039_;
 wire _02040_;
 wire _02041_;
 wire _02042_;
 wire _02043_;
 wire _02044_;
 wire _02045_;
 wire _02046_;
 wire _02047_;
 wire _02048_;
 wire _02049_;
 wire _02050_;
 wire _02051_;
 wire _02052_;
 wire _02053_;
 wire _02054_;
 wire _02055_;
 wire _02056_;
 wire _02057_;
 wire _02058_;
 wire _02059_;
 wire _02060_;
 wire _02061_;
 wire _02062_;
 wire _02063_;
 wire _02064_;
 wire _02065_;
 wire _02066_;
 wire _02067_;
 wire _02068_;
 wire _02069_;
 wire _02070_;
 wire _02071_;
 wire _02072_;
 wire _02073_;
 wire _02074_;
 wire _02075_;
 wire _02076_;
 wire _02077_;
 wire _02078_;
 wire _02079_;
 wire _02080_;
 wire _02081_;
 wire _02082_;
 wire _02083_;
 wire _02084_;
 wire _02085_;
 wire _02086_;
 wire _02087_;
 wire _02088_;
 wire _02089_;
 wire _02090_;
 wire _02091_;
 wire _02092_;
 wire _02093_;
 wire _02094_;
 wire _02095_;
 wire _02096_;
 wire _02097_;
 wire _02098_;
 wire _02099_;
 wire _02100_;
 wire _02101_;
 wire _02102_;
 wire _02103_;
 wire _02104_;
 wire _02105_;
 wire _02106_;
 wire _02107_;
 wire _02108_;
 wire _02109_;
 wire _02110_;
 wire _02111_;
 wire _02112_;
 wire _02113_;
 wire _02114_;
 wire _02115_;
 wire _02116_;
 wire _02117_;
 wire _02118_;
 wire _02119_;
 wire _02120_;
 wire _02121_;
 wire _02122_;
 wire _02123_;
 wire _02124_;
 wire _02125_;
 wire _02126_;
 wire _02127_;
 wire _02128_;
 wire _02129_;
 wire _02130_;
 wire _02131_;
 wire _02132_;
 wire _02133_;
 wire _02134_;
 wire _02135_;
 wire _02136_;
 wire _02137_;
 wire _02138_;
 wire _02139_;
 wire _02140_;
 wire _02141_;
 wire _02142_;
 wire _02143_;
 wire _02144_;
 wire _02145_;
 wire _02146_;
 wire _02147_;
 wire _02148_;
 wire _02149_;
 wire _02150_;
 wire _02151_;
 wire _02152_;
 wire _02153_;
 wire _02154_;
 wire _02155_;
 wire _02156_;
 wire _02157_;
 wire _02158_;
 wire _02159_;
 wire _02160_;
 wire _02161_;
 wire _02162_;
 wire _02163_;
 wire _02164_;
 wire _02165_;
 wire _02166_;
 wire _02167_;
 wire _02168_;
 wire _02169_;
 wire _02170_;
 wire _02171_;
 wire _02172_;
 wire _02173_;
 wire _02174_;
 wire _02175_;
 wire _02176_;
 wire _02177_;
 wire _02178_;
 wire _02179_;
 wire _02180_;
 wire _02181_;
 wire _02182_;
 wire _02183_;
 wire _02184_;
 wire _02185_;
 wire _02186_;
 wire _02187_;
 wire _02188_;
 wire _02189_;
 wire _02190_;
 wire _02191_;
 wire _02192_;
 wire _02193_;
 wire _02194_;
 wire _02195_;
 wire _02196_;
 wire _02197_;
 wire _02198_;
 wire _02199_;
 wire _02200_;
 wire _02201_;
 wire _02202_;
 wire _02203_;
 wire _02204_;
 wire _02205_;
 wire _02206_;
 wire _02207_;
 wire _02208_;
 wire _02209_;
 wire _02210_;
 wire _02211_;
 wire _02212_;
 wire _02213_;
 wire _02214_;
 wire _02215_;
 wire _02216_;
 wire _02217_;
 wire _02218_;
 wire _02219_;
 wire _02220_;
 wire _02221_;
 wire _02222_;
 wire _02223_;
 wire _02224_;
 wire _02225_;
 wire _02226_;
 wire _02227_;
 wire _02228_;
 wire _02229_;
 wire _02230_;
 wire _02231_;
 wire _02232_;
 wire _02233_;
 wire _02234_;
 wire _02235_;
 wire _02236_;
 wire _02237_;
 wire _02238_;
 wire _02239_;
 wire _02240_;
 wire _02241_;
 wire _02242_;
 wire _02243_;
 wire _02244_;
 wire _02245_;
 wire _02246_;
 wire _02247_;
 wire _02248_;
 wire _02249_;
 wire _02250_;
 wire _02251_;
 wire _02252_;
 wire _02253_;
 wire _02254_;
 wire _02255_;
 wire _02256_;
 wire _02257_;
 wire _02258_;
 wire _02259_;
 wire _02260_;
 wire _02261_;
 wire _02262_;
 wire _02263_;
 wire _02264_;
 wire _02265_;
 wire _02266_;
 wire _02267_;
 wire _02268_;
 wire _02269_;
 wire _02270_;
 wire _02271_;
 wire _02272_;
 wire _02273_;
 wire _02274_;
 wire _02275_;
 wire _02276_;
 wire _02277_;
 wire _02278_;
 wire _02279_;
 wire _02280_;
 wire _02281_;
 wire _02282_;
 wire _02283_;
 wire _02284_;
 wire _02285_;
 wire _02286_;
 wire _02287_;
 wire _02288_;
 wire _02289_;
 wire _02290_;
 wire _02291_;
 wire _02292_;
 wire _02293_;
 wire _02294_;
 wire _02295_;
 wire _02296_;
 wire _02297_;
 wire _02298_;
 wire _02299_;
 wire _02300_;
 wire _02301_;
 wire _02302_;
 wire _02303_;
 wire _02304_;
 wire _02305_;
 wire _02306_;
 wire _02307_;
 wire _02308_;
 wire _02309_;
 wire _02310_;
 wire _02311_;
 wire _02312_;
 wire _02313_;
 wire _02314_;
 wire _02315_;
 wire _02316_;
 wire _02317_;
 wire _02318_;
 wire _02319_;
 wire _02320_;
 wire _02321_;
 wire _02322_;
 wire _02323_;
 wire _02324_;
 wire _02325_;
 wire _02326_;
 wire _02327_;
 wire _02328_;
 wire _02329_;
 wire _02330_;
 wire _02331_;
 wire _02332_;
 wire _02333_;
 wire _02334_;
 wire _02335_;
 wire _02336_;
 wire _02337_;
 wire _02338_;
 wire _02339_;
 wire _02340_;
 wire _02341_;
 wire _02342_;
 wire _02343_;
 wire _02344_;
 wire _02345_;
 wire _02346_;
 wire _02347_;
 wire _02348_;
 wire _02349_;
 wire _02350_;
 wire _02351_;
 wire _02352_;
 wire _02353_;
 wire _02354_;
 wire _02355_;
 wire _02356_;
 wire _02357_;
 wire _02358_;
 wire _02359_;
 wire _02360_;
 wire _02361_;
 wire _02362_;
 wire _02363_;
 wire _02364_;
 wire _02365_;
 wire _02366_;
 wire _02367_;
 wire _02368_;
 wire _02369_;
 wire _02370_;
 wire _02371_;
 wire _02372_;
 wire _02373_;
 wire _02374_;
 wire _02375_;
 wire _02376_;
 wire _02377_;
 wire _02378_;
 wire _02379_;
 wire _02380_;
 wire _02381_;
 wire _02382_;
 wire _02383_;
 wire _02384_;
 wire _02385_;
 wire _02386_;
 wire _02387_;
 wire _02388_;
 wire _02389_;
 wire _02390_;
 wire _02391_;
 wire _02392_;
 wire _02393_;
 wire _02394_;
 wire _02395_;
 wire _02396_;
 wire _02397_;
 wire _02398_;
 wire _02399_;
 wire _02400_;
 wire _02401_;
 wire _02402_;
 wire _02403_;
 wire _02404_;
 wire _02405_;
 wire _02406_;
 wire _02407_;
 wire _02408_;
 wire _02409_;
 wire _02410_;
 wire _02411_;
 wire _02412_;
 wire _02413_;
 wire _02414_;
 wire _02415_;
 wire _02416_;
 wire _02417_;
 wire _02418_;
 wire _02419_;
 wire _02420_;
 wire _02421_;
 wire _02422_;
 wire _02423_;
 wire _02424_;
 wire _02425_;
 wire _02426_;
 wire _02427_;
 wire _02428_;
 wire _02429_;
 wire _02430_;
 wire _02431_;
 wire _02432_;
 wire _02433_;
 wire _02434_;
 wire _02435_;
 wire _02436_;
 wire _02437_;
 wire _02438_;
 wire _02439_;
 wire _02440_;
 wire _02441_;
 wire _02442_;
 wire _02443_;
 wire _02444_;
 wire _02445_;
 wire _02446_;
 wire _02447_;
 wire _02448_;
 wire _02449_;
 wire _02450_;
 wire _02451_;
 wire _02452_;
 wire _02453_;
 wire _02454_;
 wire _02455_;
 wire _02456_;
 wire _02457_;
 wire _02458_;
 wire _02459_;
 wire _02460_;
 wire _02461_;
 wire _02462_;
 wire _02463_;
 wire _02464_;
 wire _02465_;
 wire _02466_;
 wire _02467_;
 wire _02468_;
 wire _02469_;
 wire _02470_;
 wire _02471_;
 wire _02472_;
 wire _02473_;
 wire _02474_;
 wire _02475_;
 wire _02476_;
 wire _02477_;
 wire _02478_;
 wire _02479_;
 wire _02480_;
 wire _02481_;
 wire _02482_;
 wire _02483_;
 wire _02484_;
 wire _02485_;
 wire _02486_;
 wire _02487_;
 wire _02488_;
 wire _02489_;
 wire _02490_;
 wire _02491_;
 wire _02492_;
 wire _02493_;
 wire _02494_;
 wire _02495_;
 wire _02496_;
 wire _02497_;
 wire _02498_;
 wire _02499_;
 wire _02500_;
 wire _02501_;
 wire _02502_;
 wire _02503_;
 wire _02504_;
 wire _02505_;
 wire _02506_;
 wire _02507_;
 wire _02508_;
 wire _02509_;
 wire _02510_;
 wire _02511_;
 wire _02512_;
 wire _02513_;
 wire _02514_;
 wire _02515_;
 wire _02516_;
 wire _02517_;
 wire _02518_;
 wire _02519_;
 wire _02520_;
 wire _02521_;
 wire _02522_;
 wire _02523_;
 wire _02524_;
 wire _02525_;
 wire _02526_;
 wire _02527_;
 wire _02528_;
 wire _02529_;
 wire _02530_;
 wire _02531_;
 wire _02532_;
 wire _02533_;
 wire _02534_;
 wire _02535_;
 wire _02536_;
 wire _02537_;
 wire _02538_;
 wire _02539_;
 wire _02540_;
 wire _02541_;
 wire _02542_;
 wire _02543_;
 wire _02544_;
 wire _02545_;
 wire _02546_;
 wire _02547_;
 wire _02548_;
 wire _02549_;
 wire _02550_;
 wire _02551_;
 wire _02552_;
 wire _02553_;
 wire _02554_;
 wire _02555_;
 wire _02556_;
 wire _02557_;
 wire _02558_;
 wire _02559_;
 wire _02560_;
 wire _02561_;
 wire _02562_;
 wire _02563_;
 wire _02564_;
 wire _02565_;
 wire _02566_;
 wire _02567_;
 wire _02568_;
 wire _02569_;
 wire _02570_;
 wire _02571_;
 wire _02572_;
 wire _02573_;
 wire _02574_;
 wire _02575_;
 wire _02576_;
 wire _02577_;
 wire _02578_;
 wire _02579_;
 wire _02580_;
 wire _02581_;
 wire _02582_;
 wire _02583_;
 wire _02584_;
 wire _02585_;
 wire _02586_;
 wire _02587_;
 wire _02588_;
 wire _02589_;
 wire _02590_;
 wire _02591_;
 wire _02592_;
 wire _02593_;
 wire _02594_;
 wire _02595_;
 wire _02596_;
 wire _02597_;
 wire _02598_;
 wire _02599_;
 wire _02600_;
 wire _02601_;
 wire _02602_;
 wire _02603_;
 wire _02604_;
 wire _02605_;
 wire _02606_;
 wire _02607_;
 wire _02608_;
 wire _02609_;
 wire _02610_;
 wire _02611_;
 wire _02612_;
 wire _02613_;
 wire _02614_;
 wire _02615_;
 wire _02616_;
 wire _02617_;
 wire _02618_;
 wire _02619_;
 wire _02620_;
 wire _02621_;
 wire _02622_;
 wire _02623_;
 wire _02624_;
 wire _02625_;
 wire _02626_;
 wire _02627_;
 wire _02628_;
 wire _02629_;
 wire _02630_;
 wire _02631_;
 wire _02632_;
 wire _02633_;
 wire _02634_;
 wire _02635_;
 wire _02636_;
 wire _02637_;
 wire _02638_;
 wire _02639_;
 wire _02640_;
 wire _02641_;
 wire _02642_;
 wire _02643_;
 wire _02644_;
 wire _02645_;
 wire _02646_;
 wire _02647_;
 wire _02648_;
 wire _02649_;
 wire _02650_;
 wire _02651_;
 wire _02652_;
 wire _02653_;
 wire _02654_;
 wire _02655_;
 wire _02656_;
 wire _02657_;
 wire _02658_;
 wire _02659_;
 wire _02660_;
 wire _02661_;
 wire _02662_;
 wire _02663_;
 wire _02664_;
 wire _02665_;
 wire _02666_;
 wire _02667_;
 wire _02668_;
 wire _02669_;
 wire _02670_;
 wire _02671_;
 wire _02672_;
 wire _02673_;
 wire _02674_;
 wire _02675_;
 wire _02676_;
 wire _02677_;
 wire _02678_;
 wire _02679_;
 wire _02680_;
 wire _02681_;
 wire _02682_;
 wire _02683_;
 wire _02684_;
 wire _02685_;
 wire _02686_;
 wire _02687_;
 wire _02688_;
 wire _02689_;
 wire _02690_;
 wire _02691_;
 wire _02692_;
 wire _02693_;
 wire _02694_;
 wire _02695_;
 wire _02696_;
 wire _02697_;
 wire _02698_;
 wire _02699_;
 wire _02700_;
 wire _02701_;
 wire _02702_;
 wire _02703_;
 wire _02704_;
 wire _02705_;
 wire _02706_;
 wire _02707_;
 wire _02708_;
 wire _02709_;
 wire _02710_;
 wire _02711_;
 wire _02712_;
 wire _02713_;
 wire _02714_;
 wire _02715_;
 wire _02716_;
 wire _02717_;
 wire _02718_;
 wire _02719_;
 wire _02720_;
 wire _02721_;
 wire _02722_;
 wire _02723_;
 wire _02724_;
 wire _02725_;
 wire _02726_;
 wire _02727_;
 wire _02728_;
 wire _02729_;
 wire _02730_;
 wire _02731_;
 wire _02732_;
 wire _02733_;
 wire _02734_;
 wire _02735_;
 wire _02736_;
 wire _02737_;
 wire _02738_;
 wire _02739_;
 wire _02740_;
 wire _02741_;
 wire _02742_;
 wire _02743_;
 wire _02744_;
 wire _02745_;
 wire _02746_;
 wire _02747_;
 wire _02748_;
 wire _02749_;
 wire _02750_;
 wire _02751_;
 wire _02752_;
 wire _02753_;
 wire _02754_;
 wire _02755_;
 wire _02756_;
 wire _02757_;
 wire _02758_;
 wire _02759_;
 wire _02760_;
 wire _02761_;
 wire _02762_;
 wire _02763_;
 wire _02764_;
 wire _02765_;
 wire _02766_;
 wire _02767_;
 wire _02768_;
 wire _02769_;
 wire _02770_;
 wire _02771_;
 wire _02772_;
 wire _02773_;
 wire _02774_;
 wire _02775_;
 wire _02776_;
 wire _02777_;
 wire _02778_;
 wire _02779_;
 wire _02780_;
 wire _02781_;
 wire _02782_;
 wire _02783_;
 wire _02784_;
 wire _02785_;
 wire _02786_;
 wire _02787_;
 wire _02788_;
 wire _02789_;
 wire _02790_;
 wire _02791_;
 wire _02792_;
 wire _02793_;
 wire _02794_;
 wire _02795_;
 wire _02796_;
 wire _02797_;
 wire _02798_;
 wire _02799_;
 wire _02800_;
 wire _02801_;
 wire _02802_;
 wire _02803_;
 wire _02804_;
 wire _02805_;
 wire _02806_;
 wire _02807_;
 wire _02808_;
 wire _02809_;
 wire _02810_;
 wire _02811_;
 wire _02812_;
 wire _02813_;
 wire _02814_;
 wire _02815_;
 wire _02816_;
 wire _02817_;
 wire _02818_;
 wire _02819_;
 wire _02820_;
 wire _02821_;
 wire _02822_;
 wire _02823_;
 wire _02824_;
 wire _02825_;
 wire _02826_;
 wire _02827_;
 wire _02828_;
 wire _02829_;
 wire _02830_;
 wire _02831_;
 wire _02832_;
 wire _02833_;
 wire _02834_;
 wire _02835_;
 wire _02836_;
 wire _02837_;
 wire _02838_;
 wire _02839_;
 wire _02840_;
 wire _02841_;
 wire _02842_;
 wire _02843_;
 wire _02844_;
 wire _02845_;
 wire _02846_;
 wire _02847_;
 wire _02848_;
 wire _02849_;
 wire _02850_;
 wire _02851_;
 wire _02852_;
 wire _02853_;
 wire _02854_;
 wire _02855_;
 wire _02856_;
 wire _02857_;
 wire _02858_;
 wire _02859_;
 wire _02860_;
 wire _02861_;
 wire _02862_;
 wire _02863_;
 wire _02864_;
 wire _02865_;
 wire _02866_;
 wire _02867_;
 wire _02868_;
 wire _02869_;
 wire _02870_;
 wire _02871_;
 wire _02872_;
 wire _02873_;
 wire _02874_;
 wire _02875_;
 wire _02876_;
 wire _02877_;
 wire _02878_;
 wire _02879_;
 wire _02880_;
 wire _02881_;
 wire _02882_;
 wire _02883_;
 wire _02884_;
 wire _02885_;
 wire _02886_;
 wire _02887_;
 wire _02888_;
 wire _02889_;
 wire _02890_;
 wire _02891_;
 wire _02892_;
 wire _02893_;
 wire _02894_;
 wire _02895_;
 wire _02896_;
 wire _02897_;
 wire _02898_;
 wire _02899_;
 wire _02900_;
 wire _02901_;
 wire _02902_;
 wire _02903_;
 wire _02904_;
 wire _02905_;
 wire _02906_;
 wire _02907_;
 wire _02908_;
 wire _02909_;
 wire _02910_;
 wire _02911_;
 wire _02912_;
 wire _02913_;
 wire _02914_;
 wire _02915_;
 wire _02916_;
 wire _02917_;
 wire _02918_;
 wire _02919_;
 wire _02920_;
 wire _02921_;
 wire _02922_;
 wire _02923_;
 wire _02924_;
 wire _02925_;
 wire _02926_;
 wire _02927_;
 wire _02928_;
 wire _02929_;
 wire _02930_;
 wire _02931_;
 wire _02932_;
 wire _02933_;
 wire _02934_;
 wire _02935_;
 wire _02936_;
 wire _02937_;
 wire _02938_;
 wire _02939_;
 wire _02940_;
 wire _02941_;
 wire _02942_;
 wire _02943_;
 wire _02944_;
 wire _02945_;
 wire _02946_;
 wire _02947_;
 wire _02948_;
 wire _02949_;
 wire _02950_;
 wire _02951_;
 wire _02952_;
 wire _02953_;
 wire _02954_;
 wire _02955_;
 wire _02956_;
 wire _02957_;
 wire _02958_;
 wire _02959_;
 wire _02960_;
 wire _02961_;
 wire _02962_;
 wire _02963_;
 wire _02964_;
 wire _02965_;
 wire _02966_;
 wire _02967_;
 wire _02968_;
 wire _02969_;
 wire _02970_;
 wire _02971_;
 wire _02972_;
 wire _02973_;
 wire _02974_;
 wire _02975_;
 wire _02976_;
 wire _02977_;
 wire _02978_;
 wire _02979_;
 wire _02980_;
 wire _02981_;
 wire _02982_;
 wire _02983_;
 wire _02984_;
 wire _02985_;
 wire _02986_;
 wire _02987_;
 wire _02988_;
 wire _02989_;
 wire _02990_;
 wire _02991_;
 wire _02992_;
 wire _02993_;
 wire _02994_;
 wire _02995_;
 wire _02996_;
 wire _02997_;
 wire _02998_;
 wire _02999_;
 wire _03000_;
 wire _03001_;
 wire _03002_;
 wire _03003_;
 wire _03004_;
 wire _03005_;
 wire _03006_;
 wire _03007_;
 wire _03008_;
 wire _03009_;
 wire _03010_;
 wire _03011_;
 wire _03012_;
 wire _03013_;
 wire _03014_;
 wire _03015_;
 wire _03016_;
 wire _03017_;
 wire _03018_;
 wire _03019_;
 wire _03020_;
 wire _03021_;
 wire _03022_;
 wire _03023_;
 wire _03024_;
 wire _03025_;
 wire _03026_;
 wire _03027_;
 wire _03028_;
 wire _03029_;
 wire _03030_;
 wire _03031_;
 wire _03032_;
 wire _03033_;
 wire _03034_;
 wire _03035_;
 wire _03036_;
 wire _03037_;
 wire _03038_;
 wire _03039_;
 wire _03040_;
 wire _03041_;
 wire _03042_;
 wire _03043_;
 wire _03044_;
 wire _03045_;
 wire _03046_;
 wire _03047_;
 wire _03048_;
 wire _03049_;
 wire _03050_;
 wire _03051_;
 wire _03052_;
 wire _03053_;
 wire _03054_;
 wire _03055_;
 wire _03056_;
 wire _03057_;
 wire _03058_;
 wire _03059_;
 wire _03060_;
 wire _03061_;
 wire _03062_;
 wire _03063_;
 wire _03064_;
 wire _03065_;
 wire _03066_;
 wire _03067_;
 wire _03068_;
 wire _03069_;
 wire _03070_;
 wire _03071_;
 wire _03072_;
 wire _03073_;
 wire _03074_;
 wire _03075_;
 wire _03076_;
 wire _03077_;
 wire _03078_;
 wire _03079_;
 wire _03080_;
 wire _03081_;
 wire _03082_;
 wire _03083_;
 wire _03084_;
 wire _03085_;
 wire _03086_;
 wire _03087_;
 wire _03088_;
 wire _03089_;
 wire _03090_;
 wire _03091_;
 wire _03092_;
 wire _03093_;
 wire _03094_;
 wire _03095_;
 wire _03096_;
 wire _03097_;
 wire _03098_;
 wire _03099_;
 wire _03100_;
 wire _03101_;
 wire _03102_;
 wire _03103_;
 wire _03104_;
 wire _03105_;
 wire _03106_;
 wire _03107_;
 wire _03108_;
 wire _03109_;
 wire _03110_;
 wire _03111_;
 wire _03112_;
 wire _03113_;
 wire _03114_;
 wire _03115_;
 wire _03116_;
 wire _03117_;
 wire _03118_;
 wire _03119_;
 wire _03120_;
 wire _03121_;
 wire _03122_;
 wire _03123_;
 wire _03124_;
 wire _03125_;
 wire _03126_;
 wire _03127_;
 wire _03128_;
 wire _03129_;
 wire _03130_;
 wire _03131_;
 wire _03132_;
 wire _03133_;
 wire _03134_;
 wire _03135_;
 wire _03136_;
 wire _03137_;
 wire _03138_;
 wire _03139_;
 wire _03140_;
 wire _03141_;
 wire _03142_;
 wire _03143_;
 wire _03144_;
 wire _03145_;
 wire _03146_;
 wire _03147_;
 wire _03148_;
 wire _03149_;
 wire _03150_;
 wire _03151_;
 wire _03152_;
 wire _03153_;
 wire _03154_;
 wire _03155_;
 wire _03156_;
 wire _03157_;
 wire _03158_;
 wire _03159_;
 wire _03160_;
 wire _03161_;
 wire _03162_;
 wire _03163_;
 wire _03164_;
 wire _03165_;
 wire _03166_;
 wire _03167_;
 wire _03168_;
 wire _03169_;
 wire _03170_;
 wire _03171_;
 wire _03172_;
 wire _03173_;
 wire _03174_;
 wire _03175_;
 wire _03176_;
 wire _03177_;
 wire _03178_;
 wire _03179_;
 wire _03180_;
 wire _03181_;
 wire _03182_;
 wire _03183_;
 wire _03184_;
 wire _03185_;
 wire _03186_;
 wire _03187_;
 wire _03188_;
 wire _03189_;
 wire _03190_;
 wire _03191_;
 wire _03192_;
 wire _03193_;
 wire _03194_;
 wire _03195_;
 wire _03196_;
 wire _03197_;
 wire _03198_;
 wire _03199_;
 wire _03200_;
 wire _03201_;
 wire _03202_;
 wire _03203_;
 wire _03204_;
 wire _03205_;
 wire _03206_;
 wire _03207_;
 wire _03208_;
 wire _03209_;
 wire _03210_;
 wire _03211_;
 wire _03212_;
 wire _03213_;
 wire _03214_;
 wire _03215_;
 wire _03216_;
 wire _03217_;
 wire _03218_;
 wire _03219_;
 wire _03220_;
 wire _03221_;
 wire _03222_;
 wire _03223_;
 wire _03224_;
 wire _03225_;
 wire _03226_;
 wire _03227_;
 wire _03228_;
 wire _03229_;
 wire _03230_;
 wire _03231_;
 wire _03232_;
 wire _03233_;
 wire _03234_;
 wire _03235_;
 wire _03236_;
 wire _03237_;
 wire _03238_;
 wire _03239_;
 wire _03240_;
 wire _03241_;
 wire _03242_;
 wire _03243_;
 wire _03244_;
 wire _03245_;
 wire _03246_;
 wire _03247_;
 wire _03248_;
 wire _03249_;
 wire _03250_;
 wire _03251_;
 wire _03252_;
 wire _03253_;
 wire _03254_;
 wire _03255_;
 wire _03256_;
 wire _03257_;
 wire _03258_;
 wire _03259_;
 wire _03260_;
 wire _03261_;
 wire _03262_;
 wire _03263_;
 wire _03264_;
 wire _03265_;
 wire _03266_;
 wire _03267_;
 wire _03268_;
 wire _03269_;
 wire _03270_;
 wire _03271_;
 wire _03272_;
 wire _03273_;
 wire _03274_;
 wire _03275_;
 wire _03276_;
 wire _03277_;
 wire _03278_;
 wire _03279_;
 wire _03280_;
 wire _03281_;
 wire _03282_;
 wire _03283_;
 wire _03284_;
 wire _03285_;
 wire _03286_;
 wire _03287_;
 wire _03288_;
 wire _03289_;
 wire _03290_;
 wire _03291_;
 wire _03292_;
 wire _03293_;
 wire _03294_;
 wire _03295_;
 wire _03296_;
 wire _03297_;
 wire _03298_;
 wire _03299_;
 wire _03300_;
 wire _03301_;
 wire _03302_;
 wire _03303_;
 wire _03304_;
 wire _03305_;
 wire _03306_;
 wire _03307_;
 wire _03308_;
 wire _03309_;
 wire _03310_;
 wire _03311_;
 wire _03312_;
 wire _03313_;
 wire _03314_;
 wire _03315_;
 wire _03316_;
 wire _03317_;
 wire _03318_;
 wire _03319_;
 wire _03320_;
 wire _03321_;
 wire _03322_;
 wire _03323_;
 wire _03324_;
 wire _03325_;
 wire _03326_;
 wire _03327_;
 wire _03328_;
 wire _03329_;
 wire _03330_;
 wire _03331_;
 wire _03332_;
 wire _03333_;
 wire _03334_;
 wire _03335_;
 wire _03336_;
 wire _03337_;
 wire _03338_;
 wire _03339_;
 wire _03340_;
 wire _03341_;
 wire _03342_;
 wire _03343_;
 wire _03344_;
 wire _03345_;
 wire _03346_;
 wire _03347_;
 wire _03348_;
 wire _03349_;
 wire _03350_;
 wire _03351_;
 wire _03352_;
 wire _03353_;
 wire _03354_;
 wire _03355_;
 wire _03356_;
 wire _03357_;
 wire _03358_;
 wire _03359_;
 wire _03360_;
 wire _03361_;
 wire _03362_;
 wire _03363_;
 wire _03364_;
 wire _03365_;
 wire _03366_;
 wire _03367_;
 wire _03368_;
 wire _03369_;
 wire _03370_;
 wire _03371_;
 wire _03372_;
 wire _03373_;
 wire _03374_;
 wire _03375_;
 wire _03376_;
 wire _03377_;
 wire _03378_;
 wire _03379_;
 wire _03380_;
 wire _03381_;
 wire _03382_;
 wire _03383_;
 wire _03384_;
 wire _03385_;
 wire _03386_;
 wire _03387_;
 wire _03388_;
 wire _03389_;
 wire _03390_;
 wire _03391_;
 wire _03392_;
 wire _03393_;
 wire _03394_;
 wire _03395_;
 wire _03396_;
 wire _03397_;
 wire _03398_;
 wire _03399_;
 wire _03400_;
 wire _03401_;
 wire _03402_;
 wire _03403_;
 wire _03404_;
 wire _03405_;
 wire _03406_;
 wire _03407_;
 wire _03408_;
 wire _03409_;
 wire _03410_;
 wire _03411_;
 wire _03412_;
 wire _03413_;
 wire _03414_;
 wire _03415_;
 wire _03416_;
 wire _03417_;
 wire _03418_;
 wire _03419_;
 wire _03420_;
 wire _03421_;
 wire _03422_;
 wire _03423_;
 wire _03424_;
 wire _03425_;
 wire _03426_;
 wire _03427_;
 wire _03428_;
 wire _03429_;
 wire _03430_;
 wire _03431_;
 wire _03432_;
 wire _03433_;
 wire _03434_;
 wire _03435_;
 wire _03436_;
 wire _03437_;
 wire _03438_;
 wire _03439_;
 wire _03440_;
 wire _03441_;
 wire _03442_;
 wire _03443_;
 wire _03444_;
 wire _03445_;
 wire _03446_;
 wire _03447_;
 wire _03448_;
 wire _03449_;
 wire _03450_;
 wire _03451_;
 wire _03452_;
 wire _03453_;
 wire _03454_;
 wire _03455_;
 wire _03456_;
 wire _03457_;
 wire _03458_;
 wire _03459_;
 wire _03460_;
 wire _03461_;
 wire _03462_;
 wire _03463_;
 wire _03464_;
 wire _03465_;
 wire _03466_;
 wire _03467_;
 wire _03468_;
 wire _03469_;
 wire _03470_;
 wire _03471_;
 wire _03472_;
 wire _03473_;
 wire _03474_;
 wire _03475_;
 wire _03476_;
 wire _03477_;
 wire _03478_;
 wire _03479_;
 wire _03480_;
 wire _03481_;
 wire _03482_;
 wire _03483_;
 wire _03484_;
 wire _03485_;
 wire _03486_;
 wire _03487_;
 wire _03488_;
 wire _03489_;
 wire _03490_;
 wire _03491_;
 wire _03492_;
 wire _03493_;
 wire _03494_;
 wire _03495_;
 wire _03496_;
 wire _03497_;
 wire _03498_;
 wire _03499_;
 wire _03500_;
 wire _03501_;
 wire _03502_;
 wire _03503_;
 wire _03504_;
 wire _03505_;
 wire _03506_;
 wire _03507_;
 wire _03508_;
 wire _03509_;
 wire _03510_;
 wire _03511_;
 wire _03512_;
 wire _03513_;
 wire _03514_;
 wire _03515_;
 wire _03516_;
 wire _03517_;
 wire _03518_;
 wire _03519_;
 wire _03520_;
 wire _03521_;
 wire _03522_;
 wire _03523_;
 wire _03524_;
 wire _03525_;
 wire _03526_;
 wire _03527_;
 wire _03528_;
 wire _03529_;
 wire _03530_;
 wire _03531_;
 wire _03532_;
 wire _03533_;
 wire _03534_;
 wire _03535_;
 wire _03536_;
 wire _03537_;
 wire _03538_;
 wire _03539_;
 wire _03540_;
 wire _03541_;
 wire _03542_;
 wire _03543_;
 wire _03544_;
 wire _03545_;
 wire _03546_;
 wire _03547_;
 wire _03548_;
 wire _03549_;
 wire _03550_;
 wire _03551_;
 wire _03552_;
 wire _03553_;
 wire _03554_;
 wire _03555_;
 wire _03556_;
 wire _03557_;
 wire _03558_;
 wire _03559_;
 wire _03560_;
 wire _03561_;
 wire _03562_;
 wire _03563_;
 wire _03564_;
 wire _03565_;
 wire _03566_;
 wire _03567_;
 wire _03568_;
 wire _03569_;
 wire _03570_;
 wire _03571_;
 wire _03572_;
 wire _03573_;
 wire _03574_;
 wire _03575_;
 wire _03576_;
 wire _03577_;
 wire _03578_;
 wire _03579_;
 wire _03580_;
 wire _03581_;
 wire _03582_;
 wire _03583_;
 wire _03584_;
 wire _03585_;
 wire _03586_;
 wire _03587_;
 wire _03588_;
 wire _03589_;
 wire _03590_;
 wire _03591_;
 wire _03592_;
 wire _03593_;
 wire _03594_;
 wire _03595_;
 wire _03596_;
 wire _03597_;
 wire _03598_;
 wire _03599_;
 wire _03600_;
 wire _03601_;
 wire _03602_;
 wire _03603_;
 wire _03604_;
 wire _03605_;
 wire _03606_;
 wire _03607_;
 wire _03608_;
 wire _03609_;
 wire _03610_;
 wire _03611_;
 wire _03612_;
 wire _03613_;
 wire _03614_;
 wire _03615_;
 wire _03616_;
 wire _03617_;
 wire _03618_;
 wire _03619_;
 wire _03620_;
 wire _03621_;
 wire _03622_;
 wire _03623_;
 wire _03624_;
 wire _03625_;
 wire _03626_;
 wire _03627_;
 wire _03628_;
 wire _03629_;
 wire _03630_;
 wire _03631_;
 wire _03632_;
 wire _03633_;
 wire _03634_;
 wire _03635_;
 wire _03636_;
 wire _03637_;
 wire _03638_;
 wire _03639_;
 wire _03640_;
 wire _03641_;
 wire _03642_;
 wire _03643_;
 wire _03644_;
 wire _03645_;
 wire _03646_;
 wire _03647_;
 wire _03648_;
 wire _03649_;
 wire _03650_;
 wire _03651_;
 wire _03652_;
 wire _03653_;
 wire _03654_;
 wire _03655_;
 wire _03656_;
 wire _03657_;
 wire _03658_;
 wire _03659_;
 wire _03660_;
 wire _03661_;
 wire _03662_;
 wire _03663_;
 wire _03664_;
 wire _03665_;
 wire _03666_;
 wire _03667_;
 wire _03668_;
 wire _03669_;
 wire _03670_;
 wire _03671_;
 wire _03672_;
 wire _03673_;
 wire _03674_;
 wire _03675_;
 wire _03676_;
 wire _03677_;
 wire _03678_;
 wire _03679_;
 wire _03680_;
 wire _03681_;
 wire _03682_;
 wire _03683_;
 wire _03684_;
 wire _03685_;
 wire _03686_;
 wire _03687_;
 wire _03688_;
 wire _03689_;
 wire _03690_;
 wire _03691_;
 wire _03692_;
 wire _03693_;
 wire _03694_;
 wire _03695_;
 wire _03696_;
 wire _03697_;
 wire _03698_;
 wire _03699_;
 wire _03700_;
 wire _03701_;
 wire _03702_;
 wire _03703_;
 wire _03704_;
 wire _03705_;
 wire _03706_;
 wire _03707_;
 wire _03708_;
 wire _03709_;
 wire _03710_;
 wire _03711_;
 wire _03712_;
 wire _03713_;
 wire _03714_;
 wire _03715_;
 wire _03716_;
 wire _03717_;
 wire _03718_;
 wire _03719_;
 wire _03720_;
 wire _03721_;
 wire _03722_;
 wire _03723_;
 wire _03724_;
 wire _03725_;
 wire _03726_;
 wire _03727_;
 wire _03728_;
 wire _03729_;
 wire _03730_;
 wire _03731_;
 wire _03732_;
 wire _03733_;
 wire _03734_;
 wire _03735_;
 wire _03736_;
 wire _03737_;
 wire _03738_;
 wire _03739_;
 wire _03740_;
 wire _03741_;
 wire _03742_;
 wire _03743_;
 wire _03744_;
 wire _03745_;
 wire _03746_;
 wire _03747_;
 wire _03748_;
 wire _03749_;
 wire _03750_;
 wire _03751_;
 wire _03752_;
 wire _03753_;
 wire _03754_;
 wire _03755_;
 wire _03756_;
 wire _03757_;
 wire _03758_;
 wire _03759_;
 wire _03760_;
 wire _03761_;
 wire _03762_;
 wire _03763_;
 wire _03764_;
 wire _03765_;
 wire _03766_;
 wire _03767_;
 wire _03768_;
 wire _03769_;
 wire _03770_;
 wire _03771_;
 wire _03772_;
 wire _03773_;
 wire _03774_;
 wire _03775_;
 wire _03776_;
 wire _03777_;
 wire _03778_;
 wire _03779_;
 wire _03780_;
 wire _03781_;
 wire _03782_;
 wire _03783_;
 wire _03784_;
 wire _03785_;
 wire _03786_;
 wire _03787_;
 wire _03788_;
 wire _03789_;
 wire _03790_;
 wire _03791_;
 wire _03792_;
 wire _03793_;
 wire _03794_;
 wire _03795_;
 wire _03796_;
 wire _03797_;
 wire _03798_;
 wire _03799_;
 wire _03800_;
 wire _03801_;
 wire _03802_;
 wire _03803_;
 wire _03804_;
 wire _03805_;
 wire _03806_;
 wire _03807_;
 wire _03808_;
 wire _03809_;
 wire _03810_;
 wire _03811_;
 wire _03812_;
 wire _03813_;
 wire _03814_;
 wire _03815_;
 wire _03816_;
 wire _03817_;
 wire _03818_;
 wire _03819_;
 wire _03820_;
 wire _03821_;
 wire _03822_;
 wire _03823_;
 wire _03824_;
 wire _03825_;
 wire _03826_;
 wire _03827_;
 wire _03828_;
 wire _03829_;
 wire _03830_;
 wire _03831_;
 wire _03832_;
 wire _03833_;
 wire _03834_;
 wire _03835_;
 wire _03836_;
 wire _03837_;
 wire _03838_;
 wire _03839_;
 wire _03840_;
 wire _03841_;
 wire _03842_;
 wire _03843_;
 wire _03844_;
 wire _03845_;
 wire _03846_;
 wire _03847_;
 wire _03848_;
 wire _03849_;
 wire _03850_;
 wire _03851_;
 wire _03852_;
 wire _03853_;
 wire _03854_;
 wire _03855_;
 wire _03856_;
 wire _03857_;
 wire _03858_;
 wire _03859_;
 wire _03860_;
 wire _03861_;
 wire _03862_;
 wire _03863_;
 wire _03864_;
 wire _03865_;
 wire _03866_;
 wire _03867_;
 wire _03868_;
 wire _03869_;
 wire _03870_;
 wire _03871_;
 wire _03872_;
 wire _03873_;
 wire _03874_;
 wire _03875_;
 wire _03876_;
 wire _03877_;
 wire _03878_;
 wire _03879_;
 wire _03880_;
 wire _03881_;
 wire _03882_;
 wire _03883_;
 wire _03884_;
 wire _03885_;
 wire _03886_;
 wire _03887_;
 wire _03888_;
 wire _03889_;
 wire _03890_;
 wire _03891_;
 wire _03892_;
 wire _03893_;
 wire _03894_;
 wire _03895_;
 wire _03896_;
 wire _03897_;
 wire _03898_;
 wire _03899_;
 wire _03900_;
 wire _03901_;
 wire _03902_;
 wire _03903_;
 wire _03904_;
 wire _03905_;
 wire _03906_;
 wire _03907_;
 wire _03908_;
 wire _03909_;
 wire _03910_;
 wire _03911_;
 wire _03912_;
 wire _03913_;
 wire _03914_;
 wire _03915_;
 wire _03916_;
 wire _03917_;
 wire _03918_;
 wire _03919_;
 wire _03920_;
 wire _03921_;
 wire _03922_;
 wire _03923_;
 wire _03924_;
 wire _03925_;
 wire _03926_;
 wire _03927_;
 wire _03928_;
 wire _03929_;
 wire _03930_;
 wire _03931_;
 wire _03932_;
 wire _03933_;
 wire _03934_;
 wire _03935_;
 wire _03936_;
 wire _03937_;
 wire _03938_;
 wire _03939_;
 wire _03940_;
 wire _03941_;
 wire _03942_;
 wire _03943_;
 wire _03944_;
 wire _03945_;
 wire _03946_;
 wire _03947_;
 wire _03948_;
 wire _03949_;
 wire _03950_;
 wire _03951_;
 wire _03952_;
 wire _03953_;
 wire _03954_;
 wire _03955_;
 wire _03956_;
 wire _03957_;
 wire _03958_;
 wire _03959_;
 wire _03960_;
 wire _03961_;
 wire _03962_;
 wire _03963_;
 wire _03964_;
 wire _03965_;
 wire _03966_;
 wire _03967_;
 wire _03968_;
 wire _03969_;
 wire _03970_;
 wire _03971_;
 wire _03972_;
 wire _03973_;
 wire _03974_;
 wire _03975_;
 wire _03976_;
 wire _03977_;
 wire _03978_;
 wire _03979_;
 wire _03980_;
 wire _03981_;
 wire _03982_;
 wire _03983_;
 wire _03984_;
 wire _03985_;
 wire _03986_;
 wire _03987_;
 wire _03988_;
 wire _03989_;
 wire _03990_;
 wire _03991_;
 wire _03992_;
 wire _03993_;
 wire _03994_;
 wire _03995_;
 wire _03996_;
 wire _03997_;
 wire _03998_;
 wire _03999_;
 wire _04000_;
 wire _04001_;
 wire _04002_;
 wire _04003_;
 wire _04004_;
 wire _04005_;
 wire _04006_;
 wire _04007_;
 wire _04008_;
 wire _04009_;
 wire _04010_;
 wire _04011_;
 wire _04012_;
 wire _04013_;
 wire _04014_;
 wire _04015_;
 wire _04016_;
 wire _04017_;
 wire _04018_;
 wire _04019_;
 wire _04020_;
 wire _04021_;
 wire _04022_;
 wire _04023_;
 wire _04024_;
 wire _04025_;
 wire _04026_;
 wire _04027_;
 wire _04028_;
 wire _04029_;
 wire _04030_;
 wire _04031_;
 wire _04032_;
 wire _04033_;
 wire _04034_;
 wire _04035_;
 wire _04036_;
 wire _04037_;
 wire _04038_;
 wire _04039_;
 wire _04040_;
 wire _04041_;
 wire _04042_;
 wire _04043_;
 wire _04044_;
 wire _04045_;
 wire _04046_;
 wire _04047_;
 wire _04048_;
 wire _04049_;
 wire _04050_;
 wire _04051_;
 wire _04052_;
 wire _04053_;
 wire _04054_;
 wire _04055_;
 wire _04056_;
 wire _04057_;
 wire _04058_;
 wire _04059_;
 wire _04060_;
 wire _04061_;
 wire _04062_;
 wire _04063_;
 wire _04064_;
 wire _04065_;
 wire _04066_;
 wire _04067_;
 wire _04068_;
 wire _04069_;
 wire _04070_;
 wire _04071_;
 wire _04072_;
 wire _04073_;
 wire _04074_;
 wire _04075_;
 wire _04076_;
 wire _04077_;
 wire _04078_;
 wire _04079_;
 wire _04080_;
 wire _04081_;
 wire _04082_;
 wire _04083_;
 wire _04084_;
 wire _04085_;
 wire _04086_;
 wire _04087_;
 wire _04088_;
 wire _04089_;
 wire _04090_;
 wire _04091_;
 wire _04092_;
 wire _04093_;
 wire _04094_;
 wire _04095_;
 wire _04096_;
 wire _04097_;
 wire _04098_;
 wire _04099_;
 wire _04100_;
 wire _04101_;
 wire _04102_;
 wire _04103_;
 wire _04104_;
 wire _04105_;
 wire _04106_;
 wire _04107_;
 wire _04108_;
 wire _04109_;
 wire _04110_;
 wire _04111_;
 wire _04112_;
 wire _04113_;
 wire _04114_;
 wire _04115_;
 wire _04116_;
 wire _04117_;
 wire _04118_;
 wire _04119_;
 wire _04120_;
 wire _04121_;
 wire _04122_;
 wire _04123_;
 wire _04124_;
 wire _04125_;
 wire _04126_;
 wire _04127_;
 wire _04128_;
 wire _04129_;
 wire _04130_;
 wire _04131_;
 wire _04132_;
 wire _04133_;
 wire _04134_;
 wire _04135_;
 wire _04136_;
 wire _04137_;
 wire _04138_;
 wire _04139_;
 wire _04140_;
 wire _04141_;
 wire _04142_;
 wire _04143_;
 wire _04144_;
 wire _04145_;
 wire _04146_;
 wire _04147_;
 wire _04148_;
 wire _04149_;
 wire _04150_;
 wire _04151_;
 wire _04152_;
 wire _04153_;
 wire _04154_;
 wire _04155_;
 wire _04156_;
 wire _04157_;
 wire _04158_;
 wire _04159_;
 wire _04160_;
 wire _04161_;
 wire _04162_;
 wire _04163_;
 wire _04164_;
 wire _04165_;
 wire _04166_;
 wire _04167_;
 wire _04168_;
 wire _04169_;
 wire _04170_;
 wire _04171_;
 wire _04172_;
 wire _04173_;
 wire _04174_;
 wire _04175_;
 wire _04176_;
 wire _04177_;
 wire _04178_;
 wire _04179_;
 wire _04180_;
 wire _04181_;
 wire _04182_;
 wire _04183_;
 wire _04184_;
 wire _04185_;
 wire _04186_;
 wire _04187_;
 wire _04188_;
 wire _04189_;
 wire _04190_;
 wire _04191_;
 wire _04192_;
 wire _04193_;
 wire _04194_;
 wire _04195_;
 wire _04196_;
 wire _04197_;
 wire _04198_;
 wire _04199_;
 wire _04200_;
 wire _04201_;
 wire _04202_;
 wire _04203_;
 wire _04204_;
 wire _04205_;
 wire _04206_;
 wire _04207_;
 wire _04208_;
 wire _04209_;
 wire _04210_;
 wire _04211_;
 wire _04212_;
 wire _04213_;
 wire _04214_;
 wire _04215_;
 wire _04216_;
 wire _04217_;
 wire _04218_;
 wire _04219_;
 wire _04220_;
 wire _04221_;
 wire _04222_;
 wire _04223_;
 wire _04224_;
 wire _04225_;
 wire _04226_;
 wire _04227_;
 wire _04228_;
 wire _04229_;
 wire _04230_;
 wire _04231_;
 wire _04232_;
 wire _04233_;
 wire _04234_;
 wire _04235_;
 wire _04236_;
 wire _04237_;
 wire _04238_;
 wire _04239_;
 wire _04240_;
 wire _04241_;
 wire _04242_;
 wire _04243_;
 wire _04244_;
 wire _04245_;
 wire _04246_;
 wire _04247_;
 wire _04248_;
 wire _04249_;
 wire _04250_;
 wire _04251_;
 wire _04252_;
 wire _04253_;
 wire _04254_;
 wire _04255_;
 wire _04256_;
 wire _04257_;
 wire _04258_;
 wire _04259_;
 wire _04260_;
 wire _04261_;
 wire _04262_;
 wire _04263_;
 wire _04264_;
 wire _04265_;
 wire _04266_;
 wire _04267_;
 wire _04268_;
 wire _04269_;
 wire _04270_;
 wire _04271_;
 wire _04272_;
 wire _04273_;
 wire _04274_;
 wire _04275_;
 wire _04276_;
 wire _04277_;
 wire _04278_;
 wire _04279_;
 wire _04280_;
 wire _04281_;
 wire _04282_;
 wire _04283_;
 wire _04284_;
 wire _04285_;
 wire _04286_;
 wire _04287_;
 wire _04288_;
 wire _04289_;
 wire _04290_;
 wire _04291_;
 wire _04292_;
 wire _04293_;
 wire _04294_;
 wire _04295_;
 wire _04296_;
 wire _04297_;
 wire _04298_;
 wire _04299_;
 wire _04300_;
 wire _04301_;
 wire _04302_;
 wire _04303_;
 wire _04304_;
 wire _04305_;
 wire _04306_;
 wire _04307_;
 wire _04308_;
 wire _04309_;
 wire _04310_;
 wire _04311_;
 wire _04312_;
 wire _04313_;
 wire _04314_;
 wire _04315_;
 wire _04316_;
 wire _04317_;
 wire _04318_;
 wire _04319_;
 wire _04320_;
 wire _04321_;
 wire _04322_;
 wire _04323_;
 wire _04324_;
 wire _04325_;
 wire _04326_;
 wire _04327_;
 wire _04328_;
 wire _04329_;
 wire _04330_;
 wire _04331_;
 wire _04332_;
 wire _04333_;
 wire _04334_;
 wire _04335_;
 wire _04336_;
 wire _04337_;
 wire _04338_;
 wire _04339_;
 wire _04340_;
 wire _04341_;
 wire _04342_;
 wire _04343_;
 wire _04344_;
 wire _04345_;
 wire _04346_;
 wire _04347_;
 wire _04348_;
 wire _04349_;
 wire _04350_;
 wire _04351_;
 wire _04352_;
 wire _04353_;
 wire _04354_;
 wire _04355_;
 wire _04356_;
 wire _04357_;
 wire _04358_;
 wire _04359_;
 wire _04360_;
 wire _04361_;
 wire _04362_;
 wire _04363_;
 wire _04364_;
 wire _04365_;
 wire _04366_;
 wire _04367_;
 wire _04368_;
 wire _04369_;
 wire _04370_;
 wire _04371_;
 wire _04372_;
 wire _04373_;
 wire _04374_;
 wire _04375_;
 wire _04376_;
 wire _04377_;
 wire _04378_;
 wire _04379_;
 wire _04380_;
 wire _04381_;
 wire _04382_;
 wire _04383_;
 wire _04384_;
 wire _04385_;
 wire _04386_;
 wire _04387_;
 wire _04388_;
 wire _04389_;
 wire _04390_;
 wire _04391_;
 wire _04392_;
 wire _04393_;
 wire _04394_;
 wire _04395_;
 wire _04396_;
 wire _04397_;
 wire _04398_;
 wire _04399_;
 wire _04400_;
 wire _04401_;
 wire _04402_;
 wire _04403_;
 wire _04404_;
 wire _04405_;
 wire _04406_;
 wire _04407_;
 wire _04408_;
 wire _04409_;
 wire _04410_;
 wire _04411_;
 wire _04412_;
 wire _04413_;
 wire _04414_;
 wire _04415_;
 wire _04416_;
 wire _04417_;
 wire _04418_;
 wire _04419_;
 wire _04420_;
 wire _04421_;
 wire _04422_;
 wire _04423_;
 wire _04424_;
 wire _04425_;
 wire _04426_;
 wire _04427_;
 wire _04428_;
 wire _04429_;
 wire _04430_;
 wire _04431_;
 wire _04432_;
 wire _04433_;
 wire _04434_;
 wire _04435_;
 wire _04436_;
 wire _04437_;
 wire _04438_;
 wire _04439_;
 wire _04440_;
 wire _04441_;
 wire _04442_;
 wire _04443_;
 wire _04444_;
 wire _04445_;
 wire _04446_;
 wire _04447_;
 wire _04448_;
 wire _04449_;
 wire _04450_;
 wire _04451_;
 wire _04452_;
 wire _04453_;
 wire _04454_;
 wire _04455_;
 wire _04456_;
 wire _04457_;
 wire _04458_;
 wire _04459_;
 wire _04460_;
 wire _04461_;
 wire _04462_;
 wire _04463_;
 wire _04464_;
 wire _04465_;
 wire _04466_;
 wire _04467_;
 wire _04468_;
 wire _04469_;
 wire _04470_;
 wire _04471_;
 wire _04472_;
 wire _04473_;
 wire _04474_;
 wire _04475_;
 wire _04476_;
 wire _04477_;
 wire _04478_;
 wire _04479_;
 wire _04480_;
 wire _04481_;
 wire _04482_;
 wire _04483_;
 wire _04484_;
 wire _04485_;
 wire _04486_;
 wire _04487_;
 wire _04488_;
 wire _04489_;
 wire _04490_;
 wire _04491_;
 wire _04492_;
 wire _04493_;
 wire _04494_;
 wire _04495_;
 wire _04496_;
 wire _04497_;
 wire _04498_;
 wire _04499_;
 wire _04500_;
 wire _04501_;
 wire _04502_;
 wire _04503_;
 wire _04504_;
 wire _04505_;
 wire _04506_;
 wire _04507_;
 wire _04508_;
 wire _04509_;
 wire _04510_;
 wire _04511_;
 wire _04512_;
 wire _04513_;
 wire _04514_;
 wire _04515_;
 wire _04516_;
 wire _04517_;
 wire _04518_;
 wire _04519_;
 wire _04520_;
 wire _04521_;
 wire _04522_;
 wire _04523_;
 wire _04524_;
 wire _04525_;
 wire _04526_;
 wire _04527_;
 wire _04528_;
 wire _04529_;
 wire _04530_;
 wire _04531_;
 wire _04532_;
 wire _04533_;
 wire _04534_;
 wire _04535_;
 wire _04536_;
 wire _04537_;
 wire _04538_;
 wire _04539_;
 wire _04540_;
 wire _04541_;
 wire _04542_;
 wire _04543_;
 wire _04544_;
 wire _04545_;
 wire _04546_;
 wire _04547_;
 wire _04548_;
 wire _04549_;
 wire _04550_;
 wire _04551_;
 wire _04552_;
 wire _04553_;
 wire _04554_;
 wire _04555_;
 wire _04556_;
 wire _04557_;
 wire _04558_;
 wire _04559_;
 wire _04560_;
 wire _04561_;
 wire _04562_;
 wire _04563_;
 wire _04564_;
 wire _04565_;
 wire _04566_;
 wire _04567_;
 wire _04568_;
 wire _04569_;
 wire _04570_;
 wire _04571_;
 wire _04572_;
 wire _04573_;
 wire _04574_;
 wire _04575_;
 wire _04576_;
 wire _04577_;
 wire _04578_;
 wire _04579_;
 wire _04580_;
 wire _04581_;
 wire _04582_;
 wire _04583_;
 wire _04584_;
 wire _04585_;
 wire _04586_;
 wire _04587_;
 wire _04588_;
 wire _04589_;
 wire _04590_;
 wire _04591_;
 wire _04592_;
 wire _04593_;
 wire _04594_;
 wire _04595_;
 wire _04596_;
 wire _04597_;
 wire _04598_;
 wire _04599_;
 wire _04600_;
 wire _04601_;
 wire _04602_;
 wire _04603_;
 wire _04604_;
 wire _04605_;
 wire _04606_;
 wire _04607_;
 wire _04608_;
 wire _04609_;
 wire _04610_;
 wire _04611_;
 wire _04612_;
 wire _04613_;
 wire _04614_;
 wire _04615_;
 wire _04616_;
 wire _04617_;
 wire _04618_;
 wire _04619_;
 wire _04620_;
 wire _04621_;
 wire _04622_;
 wire _04623_;
 wire _04624_;
 wire _04625_;
 wire _04626_;
 wire _04627_;
 wire _04628_;
 wire _04629_;
 wire _04630_;
 wire _04631_;
 wire _04632_;
 wire _04633_;
 wire _04634_;
 wire _04635_;
 wire _04636_;
 wire _04637_;
 wire _04638_;
 wire _04639_;
 wire _04640_;
 wire _04641_;
 wire _04642_;
 wire _04643_;
 wire _04644_;
 wire _04645_;
 wire _04646_;
 wire _04647_;
 wire _04648_;
 wire _04649_;
 wire _04650_;
 wire _04651_;
 wire _04652_;
 wire _04653_;
 wire _04654_;
 wire _04655_;
 wire _04656_;
 wire _04657_;
 wire _04658_;
 wire _04659_;
 wire _04660_;
 wire _04661_;
 wire _04662_;
 wire _04663_;
 wire _04664_;
 wire _04665_;
 wire _04666_;
 wire _04667_;
 wire _04668_;
 wire _04669_;
 wire _04670_;
 wire _04671_;
 wire _04672_;
 wire _04673_;
 wire _04674_;
 wire _04675_;
 wire _04676_;
 wire _04677_;
 wire _04678_;
 wire _04679_;
 wire _04680_;
 wire _04681_;
 wire _04682_;
 wire _04683_;
 wire _04684_;
 wire _04685_;
 wire _04686_;
 wire _04687_;
 wire _04688_;
 wire _04689_;
 wire _04690_;
 wire _04691_;
 wire _04692_;
 wire _04693_;
 wire _04694_;
 wire _04695_;
 wire _04696_;
 wire _04697_;
 wire _04698_;
 wire _04699_;
 wire _04700_;
 wire _04701_;
 wire _04702_;
 wire _04703_;
 wire _04704_;
 wire _04705_;
 wire _04706_;
 wire _04707_;
 wire _04708_;
 wire _04709_;
 wire _04710_;
 wire _04711_;
 wire _04712_;
 wire _04713_;
 wire _04714_;
 wire _04715_;
 wire _04716_;
 wire _04717_;
 wire _04718_;
 wire _04719_;
 wire _04720_;
 wire _04721_;
 wire _04722_;
 wire _04723_;
 wire _04724_;
 wire _04725_;
 wire _04726_;
 wire _04727_;
 wire _04728_;
 wire _04729_;
 wire _04730_;
 wire _04731_;
 wire _04732_;
 wire _04733_;
 wire _04734_;
 wire _04735_;
 wire _04736_;
 wire _04737_;
 wire _04738_;
 wire _04739_;
 wire _04740_;
 wire _04741_;
 wire _04742_;
 wire _04743_;
 wire _04744_;
 wire _04745_;
 wire _04746_;
 wire _04747_;
 wire _04748_;
 wire _04749_;
 wire _04750_;
 wire _04751_;
 wire _04752_;
 wire _04753_;
 wire _04754_;
 wire _04755_;
 wire _04756_;
 wire _04757_;
 wire _04758_;
 wire _04759_;
 wire _04760_;
 wire _04761_;
 wire _04762_;
 wire _04763_;
 wire _04764_;
 wire _04765_;
 wire _04766_;
 wire _04767_;
 wire _04768_;
 wire _04769_;
 wire _04770_;
 wire _04771_;
 wire _04772_;
 wire _04773_;
 wire _04774_;
 wire _04775_;
 wire _04776_;
 wire _04777_;
 wire _04778_;
 wire _04779_;
 wire _04780_;
 wire _04781_;
 wire _04782_;
 wire _04783_;
 wire _04784_;
 wire _04785_;
 wire _04786_;
 wire _04787_;
 wire _04788_;
 wire _04789_;
 wire _04790_;
 wire _04791_;
 wire _04792_;
 wire _04793_;
 wire _04794_;
 wire _04795_;
 wire _04796_;
 wire _04797_;
 wire _04798_;
 wire _04799_;
 wire _04800_;
 wire _04801_;
 wire _04802_;
 wire _04803_;
 wire _04804_;
 wire _04805_;
 wire _04806_;
 wire _04807_;
 wire _04808_;
 wire _04809_;
 wire _04810_;
 wire _04811_;
 wire _04812_;
 wire _04813_;
 wire _04814_;
 wire _04815_;
 wire _04816_;
 wire _04817_;
 wire _04818_;
 wire _04819_;
 wire _04820_;
 wire _04821_;
 wire _04822_;
 wire _04823_;
 wire _04824_;
 wire _04825_;
 wire _04826_;
 wire _04827_;
 wire _04828_;
 wire _04829_;
 wire _04830_;
 wire _04831_;
 wire _04832_;
 wire _04833_;
 wire _04834_;
 wire _04835_;
 wire _04836_;
 wire _04837_;
 wire _04838_;
 wire _04839_;
 wire _04840_;
 wire _04841_;
 wire _04842_;
 wire _04843_;
 wire _04844_;
 wire _04845_;
 wire _04846_;
 wire _04847_;
 wire _04848_;
 wire _04849_;
 wire _04850_;
 wire _04851_;
 wire _04852_;
 wire _04853_;
 wire _04854_;
 wire _04855_;
 wire _04856_;
 wire _04857_;
 wire _04858_;
 wire _04859_;
 wire _04860_;
 wire _04861_;
 wire _04862_;
 wire _04863_;
 wire _04864_;
 wire _04865_;
 wire _04866_;
 wire _04867_;
 wire _04868_;
 wire _04869_;
 wire _04870_;
 wire _04871_;
 wire _04872_;
 wire _04873_;
 wire _04874_;
 wire _04875_;
 wire _04876_;
 wire _04877_;
 wire _04878_;
 wire _04879_;
 wire _04880_;
 wire _04881_;
 wire _04882_;
 wire _04883_;
 wire _04884_;
 wire _04885_;
 wire _04886_;
 wire _04887_;
 wire _04888_;
 wire _04889_;
 wire _04890_;
 wire _04891_;
 wire _04892_;
 wire _04893_;
 wire _04894_;
 wire _04895_;
 wire _04896_;
 wire _04897_;
 wire _04898_;
 wire _04899_;
 wire _04900_;
 wire _04901_;
 wire _04902_;
 wire _04903_;
 wire _04904_;
 wire _04905_;
 wire _04906_;
 wire _04907_;
 wire _04908_;
 wire _04909_;
 wire _04910_;
 wire _04911_;
 wire _04912_;
 wire _04913_;
 wire _04914_;
 wire _04915_;
 wire _04916_;
 wire _04917_;
 wire _04918_;
 wire _04919_;
 wire _04920_;
 wire _04921_;
 wire _04922_;
 wire _04923_;
 wire _04924_;
 wire _04925_;
 wire _04926_;
 wire _04927_;
 wire _04928_;
 wire _04929_;
 wire _04930_;
 wire _04931_;
 wire _04932_;
 wire _04933_;
 wire _04934_;
 wire _04935_;
 wire _04936_;
 wire _04937_;
 wire _04938_;
 wire _04939_;
 wire _04940_;
 wire _04941_;
 wire _04942_;
 wire _04943_;
 wire _04944_;
 wire _04945_;
 wire _04946_;
 wire _04947_;
 wire _04948_;
 wire _04949_;
 wire _04950_;
 wire _04951_;
 wire _04952_;
 wire _04953_;
 wire _04954_;
 wire _04955_;
 wire _04956_;
 wire _04957_;
 wire _04958_;
 wire _04959_;
 wire _04960_;
 wire _04961_;
 wire _04962_;
 wire _04963_;
 wire _04964_;
 wire _04965_;
 wire _04966_;
 wire _04967_;
 wire _04968_;
 wire _04969_;
 wire _04970_;
 wire _04971_;
 wire _04972_;
 wire _04973_;
 wire _04974_;
 wire _04975_;
 wire _04976_;
 wire _04977_;
 wire _04978_;
 wire _04979_;
 wire _04980_;
 wire _04981_;
 wire _04982_;
 wire _04983_;
 wire _04984_;
 wire _04985_;
 wire _04986_;
 wire _04987_;
 wire _04988_;
 wire _04989_;
 wire _04990_;
 wire _04991_;
 wire _04992_;
 wire _04993_;
 wire _04994_;
 wire _04995_;
 wire _04996_;
 wire _04997_;
 wire _04998_;
 wire _04999_;
 wire _05000_;
 wire _05001_;
 wire _05002_;
 wire _05003_;
 wire _05004_;
 wire _05005_;
 wire _05006_;
 wire _05007_;
 wire _05008_;
 wire _05009_;
 wire _05010_;
 wire _05011_;
 wire _05012_;
 wire _05013_;
 wire _05014_;
 wire _05015_;
 wire _05016_;
 wire _05017_;
 wire _05018_;
 wire _05019_;
 wire _05020_;
 wire _05021_;
 wire _05022_;
 wire _05023_;
 wire _05024_;
 wire _05025_;
 wire _05026_;
 wire _05027_;
 wire _05028_;
 wire _05029_;
 wire _05030_;
 wire _05031_;
 wire _05032_;
 wire _05033_;
 wire _05034_;
 wire _05035_;
 wire _05036_;
 wire _05037_;
 wire _05038_;
 wire _05039_;
 wire _05040_;
 wire _05041_;
 wire _05042_;
 wire _05043_;
 wire _05044_;
 wire _05045_;
 wire _05046_;
 wire _05047_;
 wire _05048_;
 wire _05049_;
 wire _05050_;
 wire _05051_;
 wire _05052_;
 wire _05053_;
 wire _05054_;
 wire _05055_;
 wire _05056_;
 wire _05057_;
 wire _05058_;
 wire _05059_;
 wire _05060_;
 wire _05061_;
 wire _05062_;
 wire _05063_;
 wire _05064_;
 wire _05065_;
 wire _05066_;
 wire _05067_;
 wire _05068_;
 wire _05069_;
 wire _05070_;
 wire _05071_;
 wire _05072_;
 wire _05073_;
 wire _05074_;
 wire _05075_;
 wire _05076_;
 wire _05077_;
 wire _05078_;
 wire _05079_;
 wire _05080_;
 wire _05081_;
 wire _05082_;
 wire _05083_;
 wire _05084_;
 wire _05085_;
 wire _05086_;
 wire _05087_;
 wire _05088_;
 wire _05089_;
 wire _05090_;
 wire _05091_;
 wire _05092_;
 wire _05093_;
 wire _05094_;
 wire _05095_;
 wire _05096_;
 wire _05097_;
 wire _05098_;
 wire _05099_;
 wire _05100_;
 wire _05101_;
 wire _05102_;
 wire _05103_;
 wire _05104_;
 wire _05105_;
 wire _05106_;
 wire _05107_;
 wire _05108_;
 wire _05109_;
 wire _05110_;
 wire _05111_;
 wire _05112_;
 wire _05113_;
 wire _05114_;
 wire _05115_;
 wire _05116_;
 wire _05117_;
 wire _05118_;
 wire _05119_;
 wire _05120_;
 wire _05121_;
 wire _05122_;
 wire _05123_;
 wire _05124_;
 wire _05125_;
 wire _05126_;
 wire _05127_;
 wire _05128_;
 wire _05129_;
 wire _05130_;
 wire _05131_;
 wire _05132_;
 wire _05133_;
 wire _05134_;
 wire _05135_;
 wire _05136_;
 wire _05137_;
 wire _05138_;
 wire _05139_;
 wire _05140_;
 wire _05141_;
 wire _05142_;
 wire _05143_;
 wire _05144_;
 wire _05145_;
 wire _05146_;
 wire _05147_;
 wire _05148_;
 wire _05149_;
 wire _05150_;
 wire _05151_;
 wire _05152_;
 wire _05153_;
 wire _05154_;
 wire _05155_;
 wire _05156_;
 wire _05157_;
 wire _05158_;
 wire _05159_;
 wire _05160_;
 wire _05161_;
 wire _05162_;
 wire _05163_;
 wire _05164_;
 wire _05165_;
 wire _05166_;
 wire _05167_;
 wire _05168_;
 wire _05169_;
 wire _05170_;
 wire _05171_;
 wire _05172_;
 wire _05173_;
 wire _05174_;
 wire _05175_;
 wire _05176_;
 wire _05177_;
 wire _05178_;
 wire _05179_;
 wire _05180_;
 wire _05181_;
 wire _05182_;
 wire _05183_;
 wire _05184_;
 wire _05185_;
 wire _05186_;
 wire _05187_;
 wire _05188_;
 wire _05189_;
 wire _05190_;
 wire _05191_;
 wire _05192_;
 wire _05193_;
 wire _05194_;
 wire _05195_;
 wire _05196_;
 wire _05197_;
 wire _05198_;
 wire _05199_;
 wire _05200_;
 wire _05201_;
 wire _05202_;
 wire _05203_;
 wire _05204_;
 wire _05205_;
 wire _05206_;
 wire _05207_;
 wire _05208_;
 wire _05209_;
 wire _05210_;
 wire _05211_;
 wire _05212_;
 wire _05213_;
 wire _05214_;
 wire _05215_;
 wire _05216_;
 wire _05217_;
 wire _05218_;
 wire _05219_;
 wire _05220_;
 wire _05221_;
 wire _05222_;
 wire _05223_;
 wire _05224_;
 wire _05225_;
 wire _05226_;
 wire _05227_;
 wire _05228_;
 wire _05229_;
 wire _05230_;
 wire _05231_;
 wire _05232_;
 wire _05233_;
 wire _05234_;
 wire _05235_;
 wire _05236_;
 wire _05237_;
 wire _05238_;
 wire _05239_;
 wire _05240_;
 wire _05241_;
 wire _05242_;
 wire _05243_;
 wire _05244_;
 wire _05245_;
 wire _05246_;
 wire _05247_;
 wire _05248_;
 wire _05249_;
 wire _05250_;
 wire _05251_;
 wire _05252_;
 wire _05253_;
 wire _05254_;
 wire _05255_;
 wire _05256_;
 wire _05257_;
 wire _05258_;
 wire _05259_;
 wire _05260_;
 wire _05261_;
 wire _05262_;
 wire _05263_;
 wire _05264_;
 wire _05265_;
 wire _05266_;
 wire _05267_;
 wire _05268_;
 wire _05269_;
 wire _05270_;
 wire _05271_;
 wire _05272_;
 wire _05273_;
 wire _05274_;
 wire _05275_;
 wire _05276_;
 wire _05277_;
 wire _05278_;
 wire _05279_;
 wire _05280_;
 wire _05281_;
 wire _05282_;
 wire _05283_;
 wire _05284_;
 wire _05285_;
 wire _05286_;
 wire _05287_;
 wire _05288_;
 wire _05289_;
 wire _05290_;
 wire _05291_;
 wire _05292_;
 wire _05293_;
 wire _05294_;
 wire _05295_;
 wire _05296_;
 wire _05297_;
 wire _05298_;
 wire _05299_;
 wire _05300_;
 wire _05301_;
 wire _05302_;
 wire _05303_;
 wire _05304_;
 wire _05305_;
 wire _05306_;
 wire _05307_;
 wire _05308_;
 wire _05309_;
 wire _05310_;
 wire _05311_;
 wire _05312_;
 wire _05313_;
 wire _05314_;
 wire _05315_;
 wire _05316_;
 wire _05317_;
 wire _05318_;
 wire _05319_;
 wire _05320_;
 wire _05321_;
 wire _05322_;
 wire _05323_;
 wire _05324_;
 wire _05325_;
 wire _05326_;
 wire _05327_;
 wire _05328_;
 wire _05329_;
 wire _05330_;
 wire _05331_;
 wire _05332_;
 wire _05333_;
 wire _05334_;
 wire _05335_;
 wire _05336_;
 wire _05337_;
 wire _05338_;
 wire _05339_;
 wire _05340_;
 wire _05341_;
 wire _05342_;
 wire _05343_;
 wire _05344_;
 wire _05345_;
 wire _05346_;
 wire _05347_;
 wire _05348_;
 wire _05349_;
 wire _05350_;
 wire _05351_;
 wire _05352_;
 wire _05353_;
 wire _05354_;
 wire _05355_;
 wire _05356_;
 wire _05357_;
 wire _05358_;
 wire _05359_;
 wire _05360_;
 wire _05361_;
 wire _05362_;
 wire _05363_;
 wire _05364_;
 wire _05365_;
 wire _05366_;
 wire _05367_;
 wire _05368_;
 wire _05369_;
 wire _05370_;
 wire _05371_;
 wire _05372_;
 wire _05373_;
 wire _05374_;
 wire _05375_;
 wire _05376_;
 wire _05377_;
 wire _05378_;
 wire _05379_;
 wire _05380_;
 wire _05381_;
 wire _05382_;
 wire _05383_;
 wire _05384_;
 wire _05385_;
 wire _05386_;
 wire _05387_;
 wire _05388_;
 wire _05389_;
 wire _05390_;
 wire _05391_;
 wire _05392_;
 wire _05393_;
 wire _05394_;
 wire _05395_;
 wire _05396_;
 wire _05397_;
 wire _05398_;
 wire _05399_;
 wire _05400_;
 wire _05401_;
 wire _05402_;
 wire _05403_;
 wire _05404_;
 wire _05405_;
 wire _05406_;
 wire _05407_;
 wire _05408_;
 wire _05409_;
 wire _05410_;
 wire _05411_;
 wire _05412_;
 wire _05413_;
 wire _05414_;
 wire _05415_;
 wire _05416_;
 wire _05417_;
 wire _05418_;
 wire _05419_;
 wire _05420_;
 wire _05421_;
 wire _05422_;
 wire _05423_;
 wire _05424_;
 wire _05425_;
 wire _05426_;
 wire _05427_;
 wire _05428_;
 wire _05429_;
 wire _05430_;
 wire _05431_;
 wire _05432_;
 wire _05433_;
 wire _05434_;
 wire _05435_;
 wire _05436_;
 wire _05437_;
 wire _05438_;
 wire _05439_;
 wire _05440_;
 wire _05441_;
 wire _05442_;
 wire _05443_;
 wire _05444_;
 wire _05445_;
 wire _05446_;
 wire _05447_;
 wire _05448_;
 wire _05449_;
 wire _05450_;
 wire _05451_;
 wire _05452_;
 wire _05453_;
 wire _05454_;
 wire _05455_;
 wire _05456_;
 wire _05457_;
 wire _05458_;
 wire _05459_;
 wire _05460_;
 wire _05461_;
 wire _05462_;
 wire _05463_;
 wire _05464_;
 wire _05465_;
 wire _05466_;
 wire _05467_;
 wire _05468_;
 wire _05469_;
 wire _05470_;
 wire _05471_;
 wire _05472_;
 wire _05473_;
 wire _05474_;
 wire _05475_;
 wire _05476_;
 wire _05477_;
 wire _05478_;
 wire _05479_;
 wire _05480_;
 wire _05481_;
 wire _05482_;
 wire _05483_;
 wire _05484_;
 wire _05485_;
 wire _05486_;
 wire _05487_;
 wire _05488_;
 wire _05489_;
 wire _05490_;
 wire _05491_;
 wire _05492_;
 wire _05493_;
 wire _05494_;
 wire _05495_;
 wire _05496_;
 wire _05497_;
 wire _05498_;
 wire _05499_;
 wire _05500_;
 wire _05501_;
 wire _05502_;
 wire _05503_;
 wire _05504_;
 wire _05505_;
 wire _05506_;
 wire _05507_;
 wire _05508_;
 wire _05509_;
 wire _05510_;
 wire _05511_;
 wire _05512_;
 wire _05513_;
 wire _05514_;
 wire _05515_;
 wire _05516_;
 wire _05517_;
 wire _05518_;
 wire _05519_;
 wire _05520_;
 wire _05521_;
 wire _05522_;
 wire _05523_;
 wire _05524_;
 wire _05525_;
 wire _05526_;
 wire _05527_;
 wire _05528_;
 wire _05529_;
 wire _05530_;
 wire _05531_;
 wire _05532_;
 wire _05533_;
 wire _05534_;
 wire _05535_;
 wire _05536_;
 wire _05537_;
 wire _05538_;
 wire _05539_;
 wire _05540_;
 wire _05541_;
 wire _05542_;
 wire _05543_;
 wire _05544_;
 wire _05545_;
 wire _05546_;
 wire _05547_;
 wire _05548_;
 wire _05549_;
 wire _05550_;
 wire _05551_;
 wire _05552_;
 wire _05553_;
 wire _05554_;
 wire _05555_;
 wire _05556_;
 wire _05557_;
 wire _05558_;
 wire _05559_;
 wire _05560_;
 wire _05561_;
 wire _05562_;
 wire _05563_;
 wire _05564_;
 wire _05565_;
 wire _05566_;
 wire _05567_;
 wire _05568_;
 wire _05569_;
 wire _05570_;
 wire _05571_;
 wire _05572_;
 wire _05573_;
 wire _05574_;
 wire _05575_;
 wire _05576_;
 wire _05577_;
 wire _05578_;
 wire _05579_;
 wire _05580_;
 wire _05581_;
 wire _05582_;
 wire _05583_;
 wire _05584_;
 wire _05585_;
 wire _05586_;
 wire _05587_;
 wire _05588_;
 wire _05589_;
 wire _05590_;
 wire _05591_;
 wire _05592_;
 wire _05593_;
 wire _05594_;
 wire _05595_;
 wire _05596_;
 wire _05597_;
 wire _05598_;
 wire _05599_;
 wire _05600_;
 wire _05601_;
 wire _05602_;
 wire _05603_;
 wire _05604_;
 wire _05605_;
 wire _05606_;
 wire _05607_;
 wire _05608_;
 wire _05609_;
 wire _05610_;
 wire _05611_;
 wire _05612_;
 wire _05613_;
 wire _05614_;
 wire _05615_;
 wire _05616_;
 wire _05617_;
 wire _05618_;
 wire _05619_;
 wire _05620_;
 wire _05621_;
 wire _05622_;
 wire _05623_;
 wire _05624_;
 wire _05625_;
 wire _05626_;
 wire _05627_;
 wire _05628_;
 wire _05629_;
 wire _05630_;
 wire _05631_;
 wire _05632_;
 wire _05633_;
 wire _05634_;
 wire _05635_;
 wire clknet_leaf_0_clk;
 wire advance_frame;
 wire \dtop.detune_counter[10] ;
 wire \dtop.detune_counter[11] ;
 wire \dtop.detune_counter[12] ;
 wire \dtop.detune_counter[13] ;
 wire \dtop.detune_counter[14] ;
 wire \dtop.detune_counter[15] ;
 wire \dtop.detune_counter[16] ;
 wire \dtop.detune_counter[17] ;
 wire \dtop.detune_counter[4] ;
 wire \dtop.detune_counter[5] ;
 wire \dtop.detune_counter[6] ;
 wire \dtop.detune_counter[7] ;
 wire \dtop.detune_counter[8] ;
 wire \dtop.detune_counter[9] ;
 wire \dtop.enable ;
 wire \dtop.ext_control[0] ;
 wire \dtop.ext_control[1] ;
 wire \dtop.ext_control[2] ;
 wire \dtop.ext_control[3] ;
 wire \dtop.ext_control[4] ;
 wire \dtop.ext_control[5] ;
 wire \dtop.ext_control[6] ;
 wire \dtop.out_sample[0] ;
 wire \dtop.out_sample[1] ;
 wire \dtop.out_sample[2] ;
 wire \dtop.out_sample[3] ;
 wire \dtop.out_sample[4] ;
 wire \dtop.out_sample[5] ;
 wire \dtop.out_sample[6] ;
 wire \dtop.player_inst.oct_counter[0] ;
 wire \dtop.player_inst.oct_counter[1] ;
 wire \dtop.player_inst.oct_counter[2] ;
 wire \dtop.player_inst.oct_counter[3] ;
 wire \dtop.player_inst.oct_counter[4] ;
 wire \dtop.player_inst.oct_counter[5] ;
 wire \dtop.player_inst.oct_counter[6] ;
 wire \dtop.player_inst.program_addr[0] ;
 wire \dtop.player_inst.program_addr[1] ;
 wire \dtop.player_inst.program_addr[2] ;
 wire \dtop.player_inst.program_addr[3] ;
 wire \dtop.player_inst.program_addr[4] ;
 wire \dtop.player_inst.program_addr[5] ;
 wire \dtop.player_inst.program_addr[6] ;
 wire \dtop.player_inst.synth.alu.acc[0] ;
 wire \dtop.player_inst.synth.alu.acc[10] ;
 wire \dtop.player_inst.synth.alu.acc[1] ;
 wire \dtop.player_inst.synth.alu.acc[2] ;
 wire \dtop.player_inst.synth.alu.acc[3] ;
 wire \dtop.player_inst.synth.alu.acc[4] ;
 wire \dtop.player_inst.synth.alu.acc[5] ;
 wire \dtop.player_inst.synth.alu.acc[6] ;
 wire \dtop.player_inst.synth.alu.acc[7] ;
 wire \dtop.player_inst.synth.alu.acc[8] ;
 wire \dtop.player_inst.synth.alu.acc[9] ;
 wire \dtop.player_inst.synth.alu.carry ;
 wire \dtop.player_inst.synth.alu.oct_en ;
 wire \dtop.player_inst.synth.alu.registers[0][0] ;
 wire \dtop.player_inst.synth.alu.registers[0][10] ;
 wire \dtop.player_inst.synth.alu.registers[0][1] ;
 wire \dtop.player_inst.synth.alu.registers[0][2] ;
 wire \dtop.player_inst.synth.alu.registers[0][3] ;
 wire \dtop.player_inst.synth.alu.registers[0][4] ;
 wire \dtop.player_inst.synth.alu.registers[0][5] ;
 wire \dtop.player_inst.synth.alu.registers[0][6] ;
 wire \dtop.player_inst.synth.alu.registers[0][7] ;
 wire \dtop.player_inst.synth.alu.registers[0][8] ;
 wire \dtop.player_inst.synth.alu.registers[0][9] ;
 wire \dtop.player_inst.synth.alu.registers[1][0] ;
 wire \dtop.player_inst.synth.alu.registers[1][10] ;
 wire \dtop.player_inst.synth.alu.registers[1][1] ;
 wire \dtop.player_inst.synth.alu.registers[1][2] ;
 wire \dtop.player_inst.synth.alu.registers[1][3] ;
 wire \dtop.player_inst.synth.alu.registers[1][4] ;
 wire \dtop.player_inst.synth.alu.registers[1][5] ;
 wire \dtop.player_inst.synth.alu.registers[1][6] ;
 wire \dtop.player_inst.synth.alu.registers[1][7] ;
 wire \dtop.player_inst.synth.alu.registers[1][8] ;
 wire \dtop.player_inst.synth.alu.registers[1][9] ;
 wire \dtop.player_inst.synth.alu.registers[2][0] ;
 wire \dtop.player_inst.synth.alu.registers[2][1] ;
 wire \dtop.player_inst.synth.alu.registers[2][2] ;
 wire \dtop.player_inst.synth.alu.registers[2][3] ;
 wire \dtop.player_inst.synth.alu.registers[2][4] ;
 wire \dtop.player_inst.synth.alu.registers[2][5] ;
 wire \dtop.player_inst.synth.alu.registers[2][6] ;
 wire \dtop.player_inst.synth.alu.registers[2][7] ;
 wire \dtop.player_inst.synth.alu.registers[3][0] ;
 wire \dtop.player_inst.synth.alu.registers[3][1] ;
 wire \dtop.player_inst.synth.alu.registers[3][2] ;
 wire \dtop.player_inst.synth.alu.registers[3][3] ;
 wire \dtop.player_inst.synth.alu.registers[3][4] ;
 wire \dtop.player_inst.synth.alu.registers[3][5] ;
 wire \dtop.player_inst.synth.alu.registers[3][6] ;
 wire \dtop.player_inst.synth.alu.registers[3][7] ;
 wire \dtop.player_inst.synth.alu.registers[4][0] ;
 wire \dtop.player_inst.synth.alu.registers[4][10] ;
 wire \dtop.player_inst.synth.alu.registers[4][1] ;
 wire \dtop.player_inst.synth.alu.registers[4][2] ;
 wire \dtop.player_inst.synth.alu.registers[4][3] ;
 wire \dtop.player_inst.synth.alu.registers[4][4] ;
 wire \dtop.player_inst.synth.alu.registers[4][5] ;
 wire \dtop.player_inst.synth.alu.registers[4][6] ;
 wire \dtop.player_inst.synth.alu.registers[4][7] ;
 wire \dtop.player_inst.synth.alu.registers[4][8] ;
 wire \dtop.player_inst.synth.alu.registers[4][9] ;
 wire \dtop.player_inst.synth.alu.registers[5][0] ;
 wire \dtop.player_inst.synth.alu.registers[5][1] ;
 wire \dtop.player_inst.synth.alu.registers[5][2] ;
 wire \dtop.player_inst.synth.alu.registers[5][3] ;
 wire \dtop.player_inst.synth.alu.registers[5][4] ;
 wire \dtop.player_inst.synth.alu.registers[5][5] ;
 wire \dtop.player_inst.synth.alu.registers[5][6] ;
 wire \dtop.vsync ;
 wire \dtop.vtop.color[10] ;
 wire \dtop.vtop.color[11] ;
 wire \dtop.vtop.color[6] ;
 wire \dtop.vtop.color[7] ;
 wire \dtop.vtop.color[8] ;
 wire \dtop.vtop.color[9] ;
 wire \dtop.vtop.dphases[0][0] ;
 wire \dtop.vtop.dphases[0][10] ;
 wire \dtop.vtop.dphases[0][1] ;
 wire \dtop.vtop.dphases[0][2] ;
 wire \dtop.vtop.dphases[0][3] ;
 wire \dtop.vtop.dphases[0][4] ;
 wire \dtop.vtop.dphases[0][5] ;
 wire \dtop.vtop.dphases[0][6] ;
 wire \dtop.vtop.dphases[0][7] ;
 wire \dtop.vtop.dphases[0][8] ;
 wire \dtop.vtop.dphases[0][9] ;
 wire \dtop.vtop.dphases[1][0] ;
 wire \dtop.vtop.dphases[1][10] ;
 wire \dtop.vtop.dphases[1][1] ;
 wire \dtop.vtop.dphases[1][2] ;
 wire \dtop.vtop.dphases[1][3] ;
 wire \dtop.vtop.dphases[1][4] ;
 wire \dtop.vtop.dphases[1][5] ;
 wire \dtop.vtop.dphases[1][6] ;
 wire \dtop.vtop.dphases[1][7] ;
 wire \dtop.vtop.dphases[1][8] ;
 wire \dtop.vtop.dphases[1][9] ;
 wire \dtop.vtop.dphases[2][0] ;
 wire \dtop.vtop.dphases[2][10] ;
 wire \dtop.vtop.dphases[2][1] ;
 wire \dtop.vtop.dphases[2][2] ;
 wire \dtop.vtop.dphases[2][3] ;
 wire \dtop.vtop.dphases[2][4] ;
 wire \dtop.vtop.dphases[2][5] ;
 wire \dtop.vtop.dphases[2][6] ;
 wire \dtop.vtop.dphases[2][7] ;
 wire \dtop.vtop.dphases[2][8] ;
 wire \dtop.vtop.dphases[2][9] ;
 wire \dtop.vtop.force_sat0 ;
 wire \dtop.vtop.logo.addr[10] ;
 wire \dtop.vtop.logo.addr[11] ;
 wire \dtop.vtop.logo.addr[7] ;
 wire \dtop.vtop.logo.addr[8] ;
 wire \dtop.vtop.logo.addr[9] ;
 wire \dtop.vtop.logo_d[1] ;
 wire \dtop.vtop.pipeline.cosappr_acc[0] ;
 wire \dtop.vtop.pipeline.cosappr_acc[1] ;
 wire \dtop.vtop.pipeline.cosappr_acc[2] ;
 wire \dtop.vtop.pipeline.cosappr_acc[3] ;
 wire \dtop.vtop.pipeline.cosappr_acc[4] ;
 wire \dtop.vtop.pipeline.cosappr_acc[5] ;
 wire \dtop.vtop.pipeline.cosappr_acc[6] ;
 wire \dtop.vtop.pipeline.cosappr_acc[7] ;
 wire \dtop.vtop.pipeline.cosappr_acc[8] ;
 wire \dtop.vtop.pipeline.dz[0] ;
 wire \dtop.vtop.pipeline.dz[1] ;
 wire \dtop.vtop.pipeline.dz[2] ;
 wire \dtop.vtop.pipeline.dz[3] ;
 wire \dtop.vtop.pipeline.dz[4] ;
 wire \dtop.vtop.pipeline.dz[5] ;
 wire \dtop.vtop.pipeline.dz[6] ;
 wire \dtop.vtop.pipeline.dz[7] ;
 wire \dtop.vtop.pipeline.dz[8] ;
 wire \dtop.vtop.pipeline.neg_t[0] ;
 wire \dtop.vtop.pipeline.neg_t[1] ;
 wire \dtop.vtop.pipeline.neg_t[2] ;
 wire \dtop.vtop.pipeline.neg_t[3] ;
 wire \dtop.vtop.pipeline.neg_t[4] ;
 wire \dtop.vtop.pipeline.neg_t[5] ;
 wire \dtop.vtop.pipeline.neg_t[6] ;
 wire \dtop.vtop.pipeline.neg_t[7] ;
 wire \dtop.vtop.pipeline.neg_t[8] ;
 wire \dtop.vtop.pipeline.neg_t[9] ;
 wire \dtop.vtop.pipeline.next_nstep_counter[0] ;
 wire \dtop.vtop.pipeline.nstep[0] ;
 wire \dtop.vtop.pipeline.nstep[1] ;
 wire \dtop.vtop.pipeline.nstep_counter[0] ;
 wire \dtop.vtop.pipeline.nstep_counter[1] ;
 wire \dtop.vtop.pipeline.nstep_counter[2] ;
 wire \dtop.vtop.pipeline.nstep_counter[3] ;
 wire \dtop.vtop.pipeline.nstep_counter[4] ;
 wire \dtop.vtop.pipeline.nstep_zg[0] ;
 wire \dtop.vtop.pipeline.nstep_zg[1] ;
 wire \dtop.vtop.pipeline.phases[0][0] ;
 wire \dtop.vtop.pipeline.phases[0][10] ;
 wire \dtop.vtop.pipeline.phases[0][11] ;
 wire \dtop.vtop.pipeline.phases[0][12] ;
 wire \dtop.vtop.pipeline.phases[0][13] ;
 wire \dtop.vtop.pipeline.phases[0][14] ;
 wire \dtop.vtop.pipeline.phases[0][15] ;
 wire \dtop.vtop.pipeline.phases[0][1] ;
 wire \dtop.vtop.pipeline.phases[0][2] ;
 wire \dtop.vtop.pipeline.phases[0][3] ;
 wire \dtop.vtop.pipeline.phases[0][4] ;
 wire \dtop.vtop.pipeline.phases[0][5] ;
 wire \dtop.vtop.pipeline.phases[0][6] ;
 wire \dtop.vtop.pipeline.phases[0][7] ;
 wire \dtop.vtop.pipeline.phases[0][8] ;
 wire \dtop.vtop.pipeline.phases[0][9] ;
 wire \dtop.vtop.pipeline.phases[1][0] ;
 wire \dtop.vtop.pipeline.phases[1][10] ;
 wire \dtop.vtop.pipeline.phases[1][11] ;
 wire \dtop.vtop.pipeline.phases[1][12] ;
 wire \dtop.vtop.pipeline.phases[1][13] ;
 wire \dtop.vtop.pipeline.phases[1][14] ;
 wire \dtop.vtop.pipeline.phases[1][15] ;
 wire \dtop.vtop.pipeline.phases[1][1] ;
 wire \dtop.vtop.pipeline.phases[1][2] ;
 wire \dtop.vtop.pipeline.phases[1][3] ;
 wire \dtop.vtop.pipeline.phases[1][4] ;
 wire \dtop.vtop.pipeline.phases[1][5] ;
 wire \dtop.vtop.pipeline.phases[1][6] ;
 wire \dtop.vtop.pipeline.phases[1][7] ;
 wire \dtop.vtop.pipeline.phases[1][8] ;
 wire \dtop.vtop.pipeline.phases[1][9] ;
 wire \dtop.vtop.pipeline.phases[2][0] ;
 wire \dtop.vtop.pipeline.phases[2][10] ;
 wire \dtop.vtop.pipeline.phases[2][11] ;
 wire \dtop.vtop.pipeline.phases[2][12] ;
 wire \dtop.vtop.pipeline.phases[2][13] ;
 wire \dtop.vtop.pipeline.phases[2][14] ;
 wire \dtop.vtop.pipeline.phases[2][15] ;
 wire \dtop.vtop.pipeline.phases[2][1] ;
 wire \dtop.vtop.pipeline.phases[2][2] ;
 wire \dtop.vtop.pipeline.phases[2][3] ;
 wire \dtop.vtop.pipeline.phases[2][4] ;
 wire \dtop.vtop.pipeline.phases[2][5] ;
 wire \dtop.vtop.pipeline.phases[2][6] ;
 wire \dtop.vtop.pipeline.phases[2][7] ;
 wire \dtop.vtop.pipeline.phases[2][8] ;
 wire \dtop.vtop.pipeline.phases[2][9] ;
 wire \dtop.vtop.pipeline.wave_index[0] ;
 wire \dtop.vtop.pipeline.wave_index[1] ;
 wire \dtop.vtop.pipeline.z[0] ;
 wire \dtop.vtop.pipeline.z[10] ;
 wire \dtop.vtop.pipeline.z[11] ;
 wire \dtop.vtop.pipeline.z[12] ;
 wire \dtop.vtop.pipeline.z[13] ;
 wire \dtop.vtop.pipeline.z[14] ;
 wire \dtop.vtop.pipeline.z[1] ;
 wire \dtop.vtop.pipeline.z[2] ;
 wire \dtop.vtop.pipeline.z[3] ;
 wire \dtop.vtop.pipeline.z[4] ;
 wire \dtop.vtop.pipeline.z[5] ;
 wire \dtop.vtop.pipeline.z[6] ;
 wire \dtop.vtop.pipeline.z[7] ;
 wire \dtop.vtop.pipeline.z[8] ;
 wire \dtop.vtop.pipeline.z[9] ;
 wire \dtop.vtop.pipeline.zg[0] ;
 wire \dtop.vtop.pipeline.zg[1] ;
 wire \dtop.vtop.pipeline.zg[2] ;
 wire \dtop.vtop.pipeline.zg[3] ;
 wire \dtop.vtop.pipeline.zg[4] ;
 wire \dtop.vtop.pipeline.zg[5] ;
 wire \dtop.vtop.pipeline.zg[6] ;
 wire \dtop.vtop.pipeline.zg[7] ;
 wire \dtop.vtop.pipeline.zg[8] ;
 wire \dtop.vtop.pipeline.zg[9] ;
 wire \dtop.vtop.pipeline.zg_acc[0] ;
 wire \dtop.vtop.pipeline.zg_acc[1] ;
 wire \dtop.vtop.pipeline.zg_acc[2] ;
 wire \dtop.vtop.pipeline.zg_acc[3] ;
 wire \dtop.vtop.pipeline.zg_acc[4] ;
 wire \dtop.vtop.pipeline.zg_acc[5] ;
 wire \dtop.vtop.pipeline.zg_acc[6] ;
 wire \dtop.vtop.pipeline.zg_acc[7] ;
 wire \dtop.vtop.pipeline.zg_acc[8] ;
 wire \dtop.vtop.pipeline.zg_acc[9] ;
 wire \dtop.vtop.pipeline.zg_valid ;
 wire \dtop.vtop.rs.saturated ;
 wire \dtop.vtop.rs.scan_y.phase[0] ;
 wire \dtop.vtop.rs.scan_y.phase[1] ;
 wire \dtop.vtop.rs.x_scan.phase[0] ;
 wire \dtop.vtop.rs.x_scan.phase[1] ;
 wire rst_n_reg;
 wire \uio_out0b[5] ;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net180;
 wire net181;
 wire net182;
 wire net183;
 wire net184;
 wire net185;
 wire net186;
 wire net187;
 wire net188;
 wire net189;
 wire net190;
 wire net191;
 wire net192;
 wire net193;
 wire net194;
 wire net195;
 wire net196;
 wire net197;
 wire net198;
 wire net199;
 wire net200;
 wire net201;
 wire net202;
 wire net203;
 wire net204;
 wire net205;
 wire net206;
 wire net207;
 wire net208;
 wire net209;
 wire net210;
 wire net211;
 wire net212;
 wire net213;
 wire net214;
 wire net215;
 wire net216;
 wire net217;
 wire net218;
 wire net219;
 wire net220;
 wire net221;
 wire net222;
 wire net223;
 wire net224;
 wire net225;
 wire net226;
 wire net227;
 wire net228;
 wire net229;
 wire net230;
 wire net231;
 wire net232;
 wire net233;
 wire net234;
 wire net235;
 wire net236;
 wire net237;
 wire net238;
 wire net239;
 wire net240;
 wire net241;
 wire net242;
 wire net243;
 wire net244;
 wire net245;
 wire net246;
 wire net247;
 wire net248;
 wire net249;
 wire net250;
 wire net251;
 wire net252;
 wire net253;
 wire net254;
 wire net255;
 wire net256;
 wire net257;
 wire net258;
 wire net259;
 wire net260;
 wire net261;
 wire net262;
 wire net263;
 wire net264;
 wire net265;
 wire net266;
 wire net267;
 wire net268;
 wire net269;
 wire net270;
 wire net271;
 wire net272;
 wire net273;
 wire net274;
 wire net275;
 wire net276;
 wire net277;
 wire net278;
 wire net279;
 wire net280;
 wire net281;
 wire net282;
 wire net283;
 wire net284;
 wire net285;
 wire net286;
 wire net287;
 wire net288;
 wire net289;
 wire net290;
 wire net291;
 wire net292;
 wire net293;
 wire net294;
 wire net295;
 wire net296;
 wire net297;
 wire net298;
 wire net299;
 wire net300;
 wire net301;
 wire net302;
 wire net303;
 wire net304;
 wire net305;
 wire net306;
 wire net307;
 wire net308;
 wire net309;
 wire net310;
 wire net311;
 wire net312;
 wire net313;
 wire net314;
 wire net315;
 wire net316;
 wire net317;
 wire net318;
 wire net319;
 wire net320;
 wire net321;
 wire net322;
 wire net323;
 wire net324;
 wire net325;
 wire net326;
 wire net327;
 wire net328;
 wire net329;
 wire net330;
 wire net331;
 wire net332;
 wire net333;
 wire net334;
 wire net335;
 wire net336;
 wire net337;
 wire net338;
 wire net339;
 wire net340;
 wire net341;
 wire net342;
 wire net343;
 wire net344;
 wire net345;
 wire net346;
 wire net347;
 wire net348;
 wire net349;
 wire net350;
 wire net351;
 wire net352;
 wire net353;
 wire net354;
 wire net355;
 wire net356;
 wire net357;
 wire net358;
 wire net359;
 wire net360;
 wire net361;
 wire net362;
 wire net363;
 wire net364;
 wire net365;
 wire net366;
 wire net367;
 wire net368;
 wire net369;
 wire net370;
 wire net371;
 wire net372;
 wire net373;
 wire net374;
 wire net375;
 wire net376;
 wire net377;
 wire net378;
 wire net379;
 wire net380;
 wire net381;
 wire net382;
 wire net383;
 wire net384;
 wire net385;
 wire net386;
 wire net387;
 wire net388;
 wire net389;
 wire net390;
 wire net391;
 wire net392;
 wire net393;
 wire net394;
 wire net395;
 wire net396;
 wire net397;
 wire net398;
 wire net399;
 wire net400;
 wire net401;
 wire net402;
 wire net403;
 wire net404;
 wire net405;
 wire net406;
 wire net407;
 wire net408;
 wire net409;
 wire net410;
 wire net411;
 wire net412;
 wire net413;
 wire net414;
 wire net415;
 wire net416;
 wire net417;
 wire net418;
 wire net419;
 wire net420;
 wire net421;
 wire net422;
 wire net423;
 wire net424;
 wire net425;
 wire net426;
 wire net427;
 wire net428;
 wire net429;
 wire net430;
 wire net431;
 wire net432;
 wire net433;
 wire net434;
 wire net435;
 wire net436;
 wire net437;
 wire net438;
 wire net439;
 wire net440;
 wire net441;
 wire net442;
 wire net443;
 wire net444;
 wire net445;
 wire net446;
 wire net447;
 wire net448;
 wire net449;
 wire net450;
 wire net451;
 wire net452;
 wire net453;
 wire net454;
 wire net455;
 wire net456;
 wire net457;
 wire net458;
 wire net459;
 wire net460;
 wire net461;
 wire net462;
 wire net463;
 wire net464;
 wire net465;
 wire net466;
 wire net467;
 wire net468;
 wire net469;
 wire net470;
 wire net471;
 wire net472;
 wire net473;
 wire net474;
 wire net475;
 wire net476;
 wire net477;
 wire net478;
 wire net479;
 wire net480;
 wire net481;
 wire net482;
 wire net483;
 wire net484;
 wire net485;
 wire net486;
 wire net487;
 wire net488;
 wire net489;
 wire net490;
 wire net491;
 wire net492;
 wire net493;
 wire net494;
 wire net495;
 wire net496;
 wire net497;
 wire net498;
 wire net499;
 wire net500;
 wire net501;
 wire net502;
 wire net503;
 wire net504;
 wire net505;
 wire net506;
 wire net507;
 wire net508;
 wire net509;
 wire net510;
 wire net511;
 wire net512;
 wire net513;
 wire net514;
 wire net515;
 wire net516;
 wire net517;
 wire net518;
 wire net519;
 wire net520;
 wire net521;
 wire net522;
 wire net523;
 wire net524;
 wire net525;
 wire net526;
 wire net527;
 wire net528;
 wire net529;
 wire net530;
 wire net531;
 wire net532;
 wire net533;
 wire net534;
 wire net535;
 wire net536;
 wire net537;
 wire net538;
 wire net539;
 wire net540;
 wire net541;
 wire net542;
 wire net543;
 wire net544;
 wire net545;
 wire net546;
 wire net547;
 wire net548;
 wire net549;
 wire net550;
 wire net551;
 wire net552;
 wire net553;
 wire net554;
 wire net555;
 wire net556;
 wire net557;
 wire net558;
 wire net559;
 wire net560;
 wire net561;
 wire net562;
 wire net563;
 wire net564;
 wire net565;
 wire net566;
 wire net567;
 wire net568;
 wire net569;
 wire net570;
 wire net571;
 wire net572;
 wire net573;
 wire net574;
 wire net575;
 wire net576;
 wire net577;
 wire net578;
 wire net579;
 wire net580;
 wire net581;
 wire net582;
 wire net583;
 wire net584;
 wire net585;
 wire net586;
 wire net587;
 wire net588;
 wire net589;
 wire net590;
 wire net591;
 wire net592;
 wire net593;
 wire net594;
 wire net595;
 wire net596;
 wire net597;
 wire net598;
 wire net599;
 wire net600;
 wire net601;
 wire net602;
 wire net603;
 wire net604;
 wire net605;
 wire net606;
 wire net607;
 wire net608;
 wire net609;
 wire net610;
 wire net611;
 wire net612;
 wire net613;
 wire net614;
 wire net615;
 wire net616;
 wire net617;
 wire net618;
 wire net619;
 wire net620;
 wire net621;
 wire net622;
 wire net623;
 wire net624;
 wire net625;
 wire net626;
 wire net627;
 wire net628;
 wire net629;
 wire net630;
 wire net631;
 wire net632;
 wire net633;
 wire net634;
 wire net635;
 wire net636;
 wire net637;
 wire net638;
 wire net639;
 wire net640;
 wire net641;
 wire net642;
 wire net643;
 wire net644;
 wire net645;
 wire net646;
 wire net647;
 wire net648;
 wire net649;
 wire net650;
 wire net651;
 wire net652;
 wire net653;
 wire net654;
 wire net655;
 wire net656;
 wire net657;
 wire net658;
 wire net659;
 wire net660;
 wire net661;
 wire net662;
 wire net663;
 wire net664;
 wire net665;
 wire net666;
 wire net667;
 wire net668;
 wire net669;
 wire net670;
 wire net671;
 wire net672;
 wire net673;
 wire net674;
 wire net675;
 wire net676;
 wire net677;
 wire net678;
 wire net679;
 wire net680;
 wire net681;
 wire net682;
 wire net683;
 wire net684;
 wire net685;
 wire net686;
 wire net687;
 wire net688;
 wire net689;
 wire net690;
 wire net691;
 wire net692;
 wire net693;
 wire net694;
 wire net695;
 wire net696;
 wire net697;
 wire net698;
 wire net699;
 wire net700;
 wire net701;
 wire net702;
 wire net703;
 wire net704;
 wire net705;
 wire net706;
 wire net707;
 wire net708;
 wire net709;
 wire net710;
 wire net711;
 wire net712;
 wire net713;
 wire net714;
 wire net715;
 wire net716;
 wire net717;
 wire net718;
 wire net719;
 wire net720;
 wire net721;
 wire net722;
 wire net723;
 wire net724;
 wire net725;
 wire net726;
 wire net727;
 wire net728;
 wire net729;
 wire net730;
 wire net731;
 wire net732;
 wire net733;
 wire net734;
 wire net735;
 wire net736;
 wire net737;
 wire clknet_leaf_1_clk;
 wire clknet_leaf_2_clk;
 wire clknet_leaf_3_clk;
 wire clknet_leaf_4_clk;
 wire clknet_leaf_5_clk;
 wire clknet_leaf_6_clk;
 wire clknet_leaf_7_clk;
 wire clknet_leaf_8_clk;
 wire clknet_leaf_10_clk;
 wire clknet_leaf_11_clk;
 wire clknet_leaf_12_clk;
 wire clknet_leaf_13_clk;
 wire clknet_leaf_14_clk;
 wire clknet_leaf_15_clk;
 wire clknet_leaf_16_clk;
 wire clknet_leaf_17_clk;
 wire clknet_leaf_18_clk;
 wire clknet_leaf_19_clk;
 wire clknet_leaf_20_clk;
 wire clknet_leaf_21_clk;
 wire clknet_leaf_22_clk;
 wire clknet_leaf_23_clk;
 wire clknet_leaf_24_clk;
 wire clknet_leaf_26_clk;
 wire clknet_leaf_27_clk;
 wire clknet_leaf_28_clk;
 wire clknet_leaf_29_clk;
 wire clknet_leaf_30_clk;
 wire clknet_leaf_31_clk;
 wire clknet_leaf_33_clk;
 wire clknet_leaf_34_clk;
 wire clknet_leaf_36_clk;
 wire clknet_leaf_37_clk;
 wire clknet_leaf_38_clk;
 wire clknet_leaf_39_clk;
 wire clknet_leaf_40_clk;
 wire clknet_leaf_41_clk;
 wire clknet_leaf_42_clk;
 wire clknet_leaf_44_clk;
 wire clknet_leaf_45_clk;
 wire clknet_leaf_46_clk;
 wire clknet_leaf_47_clk;
 wire clknet_leaf_48_clk;
 wire clknet_leaf_49_clk;
 wire clknet_leaf_50_clk;
 wire clknet_leaf_51_clk;
 wire clknet_leaf_52_clk;
 wire clknet_leaf_53_clk;
 wire clknet_leaf_55_clk;
 wire clknet_leaf_56_clk;
 wire clknet_leaf_57_clk;
 wire clknet_0_clk;
 wire clknet_4_0_0_clk;
 wire clknet_4_1_0_clk;
 wire clknet_4_2_0_clk;
 wire clknet_4_3_0_clk;
 wire clknet_4_4_0_clk;
 wire clknet_4_5_0_clk;
 wire clknet_4_6_0_clk;
 wire clknet_4_7_0_clk;
 wire clknet_4_8_0_clk;
 wire clknet_4_9_0_clk;
 wire clknet_4_10_0_clk;
 wire clknet_4_11_0_clk;
 wire clknet_4_12_0_clk;
 wire clknet_4_13_0_clk;
 wire clknet_4_14_0_clk;
 wire clknet_4_15_0_clk;

 sg13g2_buf_1 _05637_ (.A(\dtop.detune_counter[16] ),
    .X(_05129_));
 sg13g2_buf_2 _05638_ (.A(\dtop.detune_counter[17] ),
    .X(_05130_));
 sg13g2_buf_1 _05639_ (.A(\dtop.detune_counter[15] ),
    .X(_05131_));
 sg13g2_buf_1 _05640_ (.A(_05131_),
    .X(_05132_));
 sg13g2_nand3b_1 _05641_ (.B(_05130_),
    .C(net402),
    .Y(_05133_),
    .A_N(_05129_));
 sg13g2_buf_2 _05642_ (.A(_05133_),
    .X(_05134_));
 sg13g2_buf_1 _05643_ (.A(_05134_),
    .X(_05135_));
 sg13g2_buf_2 _05644_ (.A(\dtop.detune_counter[13] ),
    .X(_05136_));
 sg13g2_buf_1 _05645_ (.A(_05136_),
    .X(_05137_));
 sg13g2_buf_8 _05646_ (.A(\dtop.player_inst.program_addr[3] ),
    .X(_05138_));
 sg13g2_buf_8 _05647_ (.A(_05138_),
    .X(_05139_));
 sg13g2_buf_8 _05648_ (.A(net400),
    .X(_05140_));
 sg13g2_buf_1 _05649_ (.A(net358),
    .X(_05141_));
 sg13g2_buf_1 _05650_ (.A(net329),
    .X(_05142_));
 sg13g2_buf_1 _05651_ (.A(net304),
    .X(_05143_));
 sg13g2_buf_1 _05652_ (.A(net402),
    .X(_05144_));
 sg13g2_nand2b_1 _05653_ (.Y(_05145_),
    .B(_05130_),
    .A_N(_05129_));
 sg13g2_buf_1 _05654_ (.A(_05145_),
    .X(_05146_));
 sg13g2_buf_1 _05655_ (.A(_05146_),
    .X(_05147_));
 sg13g2_nor2_2 _05656_ (.A(net357),
    .B(net328),
    .Y(_05148_));
 sg13g2_buf_1 _05657_ (.A(\dtop.detune_counter[12] ),
    .X(_05149_));
 sg13g2_buf_1 _05658_ (.A(_05149_),
    .X(_05150_));
 sg13g2_buf_2 _05659_ (.A(\dtop.detune_counter[11] ),
    .X(_05151_));
 sg13g2_buf_1 _05660_ (.A(_05151_),
    .X(_05152_));
 sg13g2_and2_1 _05661_ (.A(net399),
    .B(net398),
    .X(_05153_));
 sg13g2_buf_2 _05662_ (.A(_05153_),
    .X(_05154_));
 sg13g2_buf_1 _05663_ (.A(\dtop.player_inst.program_addr[1] ),
    .X(_05155_));
 sg13g2_buf_8 _05664_ (.A(net429),
    .X(_05156_));
 sg13g2_buf_8 _05665_ (.A(net397),
    .X(_05157_));
 sg13g2_buf_8 _05666_ (.A(\dtop.player_inst.program_addr[2] ),
    .X(_05158_));
 sg13g2_buf_8 _05667_ (.A(_05158_),
    .X(_05159_));
 sg13g2_buf_1 _05668_ (.A(net396),
    .X(_05160_));
 sg13g2_buf_1 _05669_ (.A(net355),
    .X(_05161_));
 sg13g2_nor2b_1 _05670_ (.A(net356),
    .B_N(_05161_),
    .Y(_05162_));
 sg13g2_buf_2 _05671_ (.A(_05162_),
    .X(_05163_));
 sg13g2_nand4_1 _05672_ (.B(_05148_),
    .C(_05154_),
    .A(net291),
    .Y(_05164_),
    .D(_05163_));
 sg13g2_buf_2 _05673_ (.A(_00020_),
    .X(_05165_));
 sg13g2_inv_1 _05674_ (.Y(_05166_),
    .A(_05165_));
 sg13g2_buf_1 _05675_ (.A(\dtop.player_inst.oct_counter[0] ),
    .X(_05167_));
 sg13g2_buf_8 _05676_ (.A(\dtop.player_inst.oct_counter[1] ),
    .X(_05168_));
 sg13g2_or2_1 _05677_ (.X(_05169_),
    .B(_05168_),
    .A(_05167_));
 sg13g2_buf_2 _05678_ (.A(_05169_),
    .X(_05170_));
 sg13g2_buf_8 _05679_ (.A(\dtop.player_inst.program_addr[4] ),
    .X(_05171_));
 sg13g2_nand2b_1 _05680_ (.Y(_05172_),
    .B(_00078_),
    .A_N(_05171_));
 sg13g2_buf_2 _05681_ (.A(_05172_),
    .X(_05173_));
 sg13g2_buf_2 _05682_ (.A(_00077_),
    .X(_05174_));
 sg13g2_nand2b_1 _05683_ (.Y(_05175_),
    .B(_05174_),
    .A_N(\dtop.player_inst.program_addr[5] ));
 sg13g2_or3_1 _05684_ (.A(_05170_),
    .B(_05173_),
    .C(_05175_),
    .X(_05176_));
 sg13g2_buf_1 _05685_ (.A(_05176_),
    .X(_05177_));
 sg13g2_buf_8 _05686_ (.A(net303),
    .X(_05178_));
 sg13g2_buf_1 _05687_ (.A(net290),
    .X(_05179_));
 sg13g2_inv_2 _05688_ (.Y(_05180_),
    .A(net400));
 sg13g2_buf_1 _05689_ (.A(_05180_),
    .X(_05181_));
 sg13g2_buf_2 _05690_ (.A(_05167_),
    .X(_05182_));
 sg13g2_buf_1 _05691_ (.A(\dtop.player_inst.oct_counter[2] ),
    .X(_05183_));
 sg13g2_nor2_1 _05692_ (.A(_05174_),
    .B(_05183_),
    .Y(_05184_));
 sg13g2_buf_1 _05693_ (.A(_00090_),
    .X(_05185_));
 sg13g2_inv_2 _05694_ (.Y(_05186_),
    .A(net428));
 sg13g2_o21ai_1 _05695_ (.B1(_05186_),
    .Y(_05187_),
    .A1(net395),
    .A2(_05184_));
 sg13g2_buf_1 _05696_ (.A(net428),
    .X(_05188_));
 sg13g2_nor2b_1 _05697_ (.A(net395),
    .B_N(_05183_),
    .Y(_05189_));
 sg13g2_nor3_1 _05698_ (.A(_05168_),
    .B(_05188_),
    .C(_05189_),
    .Y(_05190_));
 sg13g2_a21o_1 _05699_ (.A2(_05187_),
    .A1(_05168_),
    .B1(_05190_),
    .X(_05191_));
 sg13g2_xnor2_1 _05700_ (.Y(_05192_),
    .A(net326),
    .B(_05191_));
 sg13g2_buf_2 _05701_ (.A(_05192_),
    .X(_05193_));
 sg13g2_buf_2 _05702_ (.A(_00005_),
    .X(_05194_));
 sg13g2_inv_1 _05703_ (.Y(_05195_),
    .A(_05194_));
 sg13g2_inv_1 _05704_ (.Y(_05196_),
    .A(_05132_));
 sg13g2_buf_1 _05705_ (.A(_05129_),
    .X(_05197_));
 sg13g2_nor2b_1 _05706_ (.A(_05197_),
    .B_N(_05130_),
    .Y(_05198_));
 sg13g2_buf_1 _05707_ (.A(_05198_),
    .X(_05199_));
 sg13g2_nand3_1 _05708_ (.B(net304),
    .C(_05199_),
    .A(_05196_),
    .Y(_05200_));
 sg13g2_and2_1 _05709_ (.A(_05195_),
    .B(_05200_),
    .X(_05201_));
 sg13g2_inv_2 _05710_ (.Y(_05202_),
    .A(net397));
 sg13g2_nor2_1 _05711_ (.A(net398),
    .B(net354),
    .Y(_05203_));
 sg13g2_buf_1 _05712_ (.A(net327),
    .X(_05204_));
 sg13g2_buf_1 _05713_ (.A(net356),
    .X(_05205_));
 sg13g2_nand2b_1 _05714_ (.Y(_05206_),
    .B(net398),
    .A_N(net325));
 sg13g2_a21oi_1 _05715_ (.A1(net399),
    .A2(net302),
    .Y(_05207_),
    .B1(_05206_));
 sg13g2_nor3_1 _05716_ (.A(_05200_),
    .B(_05203_),
    .C(_05207_),
    .Y(_05208_));
 sg13g2_nor3_1 _05717_ (.A(net290),
    .B(_05201_),
    .C(_05208_),
    .Y(_05209_));
 sg13g2_buf_2 _05718_ (.A(_05209_),
    .X(_05210_));
 sg13g2_a21oi_1 _05719_ (.A1(net278),
    .A2(_05193_),
    .Y(_05211_),
    .B1(_05210_));
 sg13g2_buf_2 _05720_ (.A(_05211_),
    .X(_05212_));
 sg13g2_buf_1 _05721_ (.A(_05212_),
    .X(_05213_));
 sg13g2_buf_1 _05722_ (.A(\dtop.detune_counter[8] ),
    .X(_05214_));
 sg13g2_buf_1 _05723_ (.A(_05214_),
    .X(_05215_));
 sg13g2_buf_1 _05724_ (.A(net392),
    .X(_05216_));
 sg13g2_nand2_1 _05725_ (.Y(_05217_),
    .A(net353),
    .B(_05212_));
 sg13g2_o21ai_1 _05726_ (.B1(_05217_),
    .Y(_05218_),
    .A1(_05166_),
    .A2(net208));
 sg13g2_buf_1 _05727_ (.A(\dtop.detune_counter[10] ),
    .X(_05219_));
 sg13g2_buf_1 _05728_ (.A(_05219_),
    .X(_05220_));
 sg13g2_inv_2 _05729_ (.Y(_05221_),
    .A(net391));
 sg13g2_a21o_1 _05730_ (.A2(_05193_),
    .A1(net290),
    .B1(_05210_),
    .X(_05222_));
 sg13g2_buf_1 _05731_ (.A(_05222_),
    .X(_05223_));
 sg13g2_buf_1 _05732_ (.A(_05223_),
    .X(_05224_));
 sg13g2_buf_1 _05733_ (.A(_00001_),
    .X(_05225_));
 sg13g2_nand2_1 _05734_ (.Y(_05226_),
    .A(net427),
    .B(_05224_));
 sg13g2_o21ai_1 _05735_ (.B1(_05226_),
    .Y(_05227_),
    .A1(_05221_),
    .A2(_05224_));
 sg13g2_xnor2_1 _05736_ (.Y(_05228_),
    .A(net291),
    .B(_05191_));
 sg13g2_inv_1 _05737_ (.Y(_05229_),
    .A(_05149_));
 sg13g2_xor2_1 _05738_ (.B(net325),
    .A(net398),
    .X(_05230_));
 sg13g2_xnor2_1 _05739_ (.Y(_05231_),
    .A(_05229_),
    .B(_05230_));
 sg13g2_nor2_1 _05740_ (.A(_05200_),
    .B(_05231_),
    .Y(_05232_));
 sg13g2_xnor2_1 _05741_ (.Y(_05233_),
    .A(net302),
    .B(_05232_));
 sg13g2_nor3_1 _05742_ (.A(_05170_),
    .B(_05173_),
    .C(_05175_),
    .Y(_05234_));
 sg13g2_buf_8 _05743_ (.A(_05234_),
    .X(_05235_));
 sg13g2_buf_8 _05744_ (.A(_05235_),
    .X(_05236_));
 sg13g2_mux2_1 _05745_ (.A0(_05228_),
    .A1(_05233_),
    .S(net289),
    .X(_05237_));
 sg13g2_buf_1 _05746_ (.A(_05237_),
    .X(_05238_));
 sg13g2_buf_1 _05747_ (.A(_05238_),
    .X(_05239_));
 sg13g2_buf_1 _05748_ (.A(net232),
    .X(_05240_));
 sg13g2_mux2_1 _05749_ (.A0(_05218_),
    .A1(_05227_),
    .S(net206),
    .X(_05241_));
 sg13g2_buf_1 _05750_ (.A(_00002_),
    .X(_05242_));
 sg13g2_nand2_1 _05751_ (.Y(_05243_),
    .A(_05196_),
    .B(_05199_));
 sg13g2_buf_1 _05752_ (.A(_05243_),
    .X(_05244_));
 sg13g2_xor2_1 _05753_ (.B(net302),
    .A(net399),
    .X(_05245_));
 sg13g2_nor3_1 _05754_ (.A(net288),
    .B(_05230_),
    .C(_05245_),
    .Y(_05246_));
 sg13g2_nor3_2 _05755_ (.A(net426),
    .B(net278),
    .C(_05246_),
    .Y(_05247_));
 sg13g2_buf_1 _05756_ (.A(_05247_),
    .X(_05248_));
 sg13g2_buf_2 _05757_ (.A(_00000_),
    .X(_05249_));
 sg13g2_inv_2 _05758_ (.Y(_05250_),
    .A(_05249_));
 sg13g2_nand2_1 _05759_ (.Y(_05251_),
    .A(net399),
    .B(net208));
 sg13g2_o21ai_1 _05760_ (.B1(_05251_),
    .Y(_05252_),
    .A1(_05250_),
    .A2(net208));
 sg13g2_buf_1 _05761_ (.A(\dtop.detune_counter[14] ),
    .X(_05253_));
 sg13g2_buf_1 _05762_ (.A(_05253_),
    .X(_05254_));
 sg13g2_a22oi_1 _05763_ (.Y(_05255_),
    .B1(net208),
    .B2(net390),
    .A2(_05210_),
    .A1(_00059_));
 sg13g2_nand2_1 _05764_ (.Y(_05256_),
    .A(net206),
    .B(_05255_));
 sg13g2_o21ai_1 _05765_ (.B1(_05256_),
    .Y(_05257_),
    .A1(net206),
    .A2(_05252_));
 sg13g2_nor2_1 _05766_ (.A(net263),
    .B(_05257_),
    .Y(_05258_));
 sg13g2_a21oi_1 _05767_ (.A1(_05241_),
    .A2(net263),
    .Y(_05259_),
    .B1(_05258_));
 sg13g2_nand2_1 _05768_ (.Y(_05260_),
    .A(_05164_),
    .B(_05259_));
 sg13g2_inv_1 _05769_ (.Y(_05261_),
    .A(net426));
 sg13g2_buf_2 _05770_ (.A(_00086_),
    .X(_05262_));
 sg13g2_nand3b_1 _05771_ (.B(_05262_),
    .C(_05131_),
    .Y(_05263_),
    .A_N(_05129_));
 sg13g2_buf_1 _05772_ (.A(_05263_),
    .X(_05264_));
 sg13g2_inv_1 _05773_ (.Y(_05265_),
    .A(_05264_));
 sg13g2_nand3_1 _05774_ (.B(net426),
    .C(_05265_),
    .A(net401),
    .Y(_05266_));
 sg13g2_o21ai_1 _05775_ (.B1(_05266_),
    .Y(_05267_),
    .A1(net401),
    .A2(net426));
 sg13g2_inv_1 _05776_ (.Y(_05268_),
    .A(_05254_));
 sg13g2_a22oi_1 _05777_ (.Y(_05269_),
    .B1(_05267_),
    .B2(_05268_),
    .A2(_05264_),
    .A1(_05261_));
 sg13g2_nor2_1 _05778_ (.A(net278),
    .B(_05269_),
    .Y(_05270_));
 sg13g2_buf_1 _05779_ (.A(_05270_),
    .X(_05271_));
 sg13g2_buf_2 _05780_ (.A(\dtop.detune_counter[6] ),
    .X(_05272_));
 sg13g2_buf_2 _05781_ (.A(_00017_),
    .X(_05273_));
 sg13g2_mux4_1 _05782_ (.S0(_05223_),
    .A0(_05272_),
    .A1(_05273_),
    .A2(net353),
    .A3(_05165_),
    .S1(_05239_),
    .X(_05274_));
 sg13g2_mux2_1 _05783_ (.A0(_05227_),
    .A1(_05252_),
    .S(net206),
    .X(_05275_));
 sg13g2_or3_1 _05784_ (.A(net426),
    .B(_05179_),
    .C(_05246_),
    .X(_05276_));
 sg13g2_buf_1 _05785_ (.A(_05276_),
    .X(_05277_));
 sg13g2_mux2_1 _05786_ (.A0(_05274_),
    .A1(_05275_),
    .S(_05277_),
    .X(_05278_));
 sg13g2_buf_1 _05787_ (.A(_05278_),
    .X(_05279_));
 sg13g2_buf_1 _05788_ (.A(\dtop.vtop.logo.addr[11] ),
    .X(_05280_));
 sg13g2_buf_1 _05789_ (.A(_05280_),
    .X(_05281_));
 sg13g2_buf_1 _05790_ (.A(net289),
    .X(_05282_));
 sg13g2_nand2b_1 _05791_ (.Y(_05283_),
    .B(net277),
    .A_N(_05269_));
 sg13g2_buf_1 _05792_ (.A(_05283_),
    .X(_05284_));
 sg13g2_nand2_1 _05793_ (.Y(_05285_),
    .A(net389),
    .B(net260));
 sg13g2_and2_1 _05794_ (.A(_05279_),
    .B(_05285_),
    .X(_05286_));
 sg13g2_buf_1 _05795_ (.A(_05286_),
    .X(_05287_));
 sg13g2_inv_1 _05796_ (.Y(_05288_),
    .A(_05279_));
 sg13g2_nor2_1 _05797_ (.A(_05210_),
    .B(net261),
    .Y(_05289_));
 sg13g2_buf_1 _05798_ (.A(_00080_),
    .X(_05290_));
 sg13g2_nor3_1 _05799_ (.A(net425),
    .B(_05212_),
    .C(_05247_),
    .Y(_05291_));
 sg13g2_o21ai_1 _05800_ (.B1(net232),
    .Y(_05292_),
    .A1(_05289_),
    .A2(_05291_));
 sg13g2_buf_2 _05801_ (.A(\dtop.detune_counter[4] ),
    .X(_05293_));
 sg13g2_nand2_1 _05802_ (.Y(_05294_),
    .A(_05293_),
    .B(_05238_));
 sg13g2_nand2b_1 _05803_ (.Y(_05295_),
    .B(_05247_),
    .A_N(net232));
 sg13g2_nand3_1 _05804_ (.B(_05294_),
    .C(_05295_),
    .A(_05212_),
    .Y(_05296_));
 sg13g2_buf_1 _05805_ (.A(_05296_),
    .X(_05297_));
 sg13g2_buf_2 _05806_ (.A(\dtop.player_inst.oct_counter[3] ),
    .X(_05298_));
 sg13g2_nand2_1 _05807_ (.Y(_05299_),
    .A(_05298_),
    .B(net260));
 sg13g2_a21oi_1 _05808_ (.A1(_05292_),
    .A2(_05297_),
    .Y(_05300_),
    .B1(_05299_));
 sg13g2_inv_1 _05809_ (.Y(_05301_),
    .A(\dtop.player_inst.oct_counter[4] ));
 sg13g2_nor2_1 _05810_ (.A(_05301_),
    .B(net262),
    .Y(_05302_));
 sg13g2_buf_2 _05811_ (.A(_00019_),
    .X(_05303_));
 sg13g2_inv_1 _05812_ (.Y(_05304_),
    .A(_05303_));
 sg13g2_mux2_1 _05813_ (.A0(_05293_),
    .A1(_05304_),
    .S(_05238_),
    .X(_05305_));
 sg13g2_buf_2 _05814_ (.A(\dtop.detune_counter[5] ),
    .X(_05306_));
 sg13g2_nand3_1 _05815_ (.B(_05239_),
    .C(_05212_),
    .A(_05306_),
    .Y(_05307_));
 sg13g2_o21ai_1 _05816_ (.B1(_05307_),
    .Y(_05308_),
    .A1(_05212_),
    .A2(_05305_));
 sg13g2_nand3_1 _05817_ (.B(net208),
    .C(_05247_),
    .A(_05240_),
    .Y(_05309_));
 sg13g2_o21ai_1 _05818_ (.B1(_05309_),
    .Y(_05310_),
    .A1(_05248_),
    .A2(_05308_));
 sg13g2_buf_1 _05819_ (.A(_05310_),
    .X(_05311_));
 sg13g2_o21ai_1 _05820_ (.B1(_05311_),
    .Y(_05312_),
    .A1(_05300_),
    .A2(_05302_));
 sg13g2_nand2_1 _05821_ (.Y(_05313_),
    .A(_05292_),
    .B(_05297_));
 sg13g2_inv_1 _05822_ (.Y(_05314_),
    .A(_05298_));
 sg13g2_nor3_1 _05823_ (.A(_05301_),
    .B(_05314_),
    .C(_05270_),
    .Y(_05315_));
 sg13g2_mux2_1 _05824_ (.A0(_05290_),
    .A1(_05273_),
    .S(net232),
    .X(_05316_));
 sg13g2_nand2b_1 _05825_ (.Y(_05317_),
    .B(net261),
    .A_N(_05316_));
 sg13g2_nor2_1 _05826_ (.A(net207),
    .B(net263),
    .Y(_05318_));
 sg13g2_mux2_1 _05827_ (.A0(_05293_),
    .A1(_05272_),
    .S(net232),
    .X(_05319_));
 sg13g2_a22oi_1 _05828_ (.Y(_05320_),
    .B1(_05318_),
    .B2(_05319_),
    .A2(_05317_),
    .A1(net207));
 sg13g2_a21oi_1 _05829_ (.A1(_05313_),
    .A2(_05315_),
    .Y(_05321_),
    .B1(_05320_));
 sg13g2_buf_2 _05830_ (.A(\dtop.vtop.logo.addr[7] ),
    .X(_05322_));
 sg13g2_nand2_1 _05831_ (.Y(_05323_),
    .A(net261),
    .B(_05274_));
 sg13g2_inv_2 _05832_ (.Y(_05324_),
    .A(net425));
 sg13g2_nand3_1 _05833_ (.B(net232),
    .C(net207),
    .A(_05324_),
    .Y(_05325_));
 sg13g2_a21o_1 _05834_ (.A2(net232),
    .A1(_05293_),
    .B1(net207),
    .X(_05326_));
 sg13g2_nand3_1 _05835_ (.B(_05325_),
    .C(_05326_),
    .A(net263),
    .Y(_05327_));
 sg13g2_and2_1 _05836_ (.A(_05323_),
    .B(_05327_),
    .X(_05328_));
 sg13g2_buf_1 _05837_ (.A(_05328_),
    .X(_05329_));
 sg13g2_mux2_1 _05838_ (.A0(_05306_),
    .A1(_05303_),
    .S(net207),
    .X(_05330_));
 sg13g2_buf_1 _05839_ (.A(\dtop.detune_counter[7] ),
    .X(_05331_));
 sg13g2_buf_1 _05840_ (.A(_05331_),
    .X(_05332_));
 sg13g2_buf_1 _05841_ (.A(net388),
    .X(_05333_));
 sg13g2_buf_1 _05842_ (.A(_00022_),
    .X(_05334_));
 sg13g2_mux2_1 _05843_ (.A0(_05333_),
    .A1(net424),
    .S(net207),
    .X(_05335_));
 sg13g2_mux2_1 _05844_ (.A0(_05330_),
    .A1(_05335_),
    .S(net232),
    .X(_05336_));
 sg13g2_nor2_1 _05845_ (.A(net208),
    .B(net261),
    .Y(_05337_));
 sg13g2_a22oi_1 _05846_ (.Y(_05338_),
    .B1(_05294_),
    .B2(_05337_),
    .A2(_05336_),
    .A1(net261));
 sg13g2_buf_1 _05847_ (.A(_05338_),
    .X(_05339_));
 sg13g2_o21ai_1 _05848_ (.B1(_05339_),
    .Y(_05340_),
    .A1(_05322_),
    .A2(_05329_));
 sg13g2_a21oi_1 _05849_ (.A1(_05312_),
    .A2(_05321_),
    .Y(_05341_),
    .B1(_05340_));
 sg13g2_buf_1 _05850_ (.A(\dtop.player_inst.oct_counter[6] ),
    .X(_05342_));
 sg13g2_o21ai_1 _05851_ (.B1(net423),
    .Y(_05343_),
    .A1(_05322_),
    .A2(_05329_));
 sg13g2_a21oi_1 _05852_ (.A1(_05312_),
    .A2(_05321_),
    .Y(_05344_),
    .B1(_05343_));
 sg13g2_a21oi_2 _05853_ (.B1(_05314_),
    .Y(_05345_),
    .A2(_05297_),
    .A1(_05292_));
 sg13g2_buf_1 _05854_ (.A(\dtop.player_inst.oct_counter[4] ),
    .X(_05346_));
 sg13g2_a21oi_1 _05855_ (.A1(_05311_),
    .A2(_05345_),
    .Y(_05347_),
    .B1(net422));
 sg13g2_a221oi_1 _05856_ (.B2(_05319_),
    .C1(net262),
    .B1(_05318_),
    .A1(net207),
    .Y(_05348_),
    .A2(_05317_));
 sg13g2_o21ai_1 _05857_ (.B1(_05348_),
    .Y(_05349_),
    .A1(_05311_),
    .A2(_05345_));
 sg13g2_buf_1 _05858_ (.A(\dtop.player_inst.oct_counter[5] ),
    .X(_05350_));
 sg13g2_inv_1 _05859_ (.Y(_05351_),
    .A(net421));
 sg13g2_o21ai_1 _05860_ (.B1(_05351_),
    .Y(_05352_),
    .A1(_05347_),
    .A2(_05349_));
 sg13g2_o21ai_1 _05861_ (.B1(_05352_),
    .Y(_05353_),
    .A1(_05341_),
    .A2(_05344_));
 sg13g2_buf_1 _05862_ (.A(_05322_),
    .X(_05354_));
 sg13g2_nor2_1 _05863_ (.A(net387),
    .B(_05329_),
    .Y(_05355_));
 sg13g2_nand2_1 _05864_ (.Y(_05356_),
    .A(net423),
    .B(_05339_));
 sg13g2_nor2_1 _05865_ (.A(_05355_),
    .B(_05356_),
    .Y(_05357_));
 sg13g2_a21oi_1 _05866_ (.A1(net387),
    .A2(_05329_),
    .Y(_05358_),
    .B1(_05357_));
 sg13g2_buf_1 _05867_ (.A(\dtop.vtop.logo.addr[9] ),
    .X(_05359_));
 sg13g2_inv_2 _05868_ (.Y(_05360_),
    .A(_05359_));
 sg13g2_mux2_1 _05869_ (.A0(_05319_),
    .A1(_05316_),
    .S(net207),
    .X(_05361_));
 sg13g2_mux2_1 _05870_ (.A0(_05241_),
    .A1(_05361_),
    .S(net263),
    .X(_05362_));
 sg13g2_buf_1 _05871_ (.A(_05362_),
    .X(_05363_));
 sg13g2_nand2_2 _05872_ (.Y(_05364_),
    .A(_05360_),
    .B(_05363_));
 sg13g2_buf_2 _05873_ (.A(_00024_),
    .X(_05365_));
 sg13g2_inv_1 _05874_ (.Y(_05366_),
    .A(_05365_));
 sg13g2_buf_1 _05875_ (.A(\dtop.detune_counter[9] ),
    .X(_05367_));
 sg13g2_buf_1 _05876_ (.A(net420),
    .X(_05368_));
 sg13g2_nand2_1 _05877_ (.Y(_05369_),
    .A(net386),
    .B(_05212_));
 sg13g2_o21ai_1 _05878_ (.B1(_05369_),
    .Y(_05370_),
    .A1(_05366_),
    .A2(net208));
 sg13g2_mux2_1 _05879_ (.A0(_05335_),
    .A1(_05370_),
    .S(net206),
    .X(_05371_));
 sg13g2_and2_1 _05880_ (.A(net261),
    .B(_05371_),
    .X(_05372_));
 sg13g2_a21oi_1 _05881_ (.A1(_05248_),
    .A2(_05308_),
    .Y(_05373_),
    .B1(_05372_));
 sg13g2_buf_2 _05882_ (.A(_05373_),
    .X(_05374_));
 sg13g2_nand3_1 _05883_ (.B(_05364_),
    .C(_05374_),
    .A(net260),
    .Y(_05375_));
 sg13g2_buf_2 _05884_ (.A(\dtop.vtop.logo.addr[8] ),
    .X(_05376_));
 sg13g2_nand3_1 _05885_ (.B(net260),
    .C(_05364_),
    .A(_05376_),
    .Y(_05377_));
 sg13g2_a22oi_1 _05886_ (.Y(_05378_),
    .B1(_05375_),
    .B2(_05377_),
    .A2(_05358_),
    .A1(_05353_));
 sg13g2_nand3_1 _05887_ (.B(_05364_),
    .C(_05374_),
    .A(_05376_),
    .Y(_05379_));
 sg13g2_o21ai_1 _05888_ (.B1(_05379_),
    .Y(_05380_),
    .A1(_05360_),
    .A2(_05363_));
 sg13g2_or2_1 _05889_ (.X(_05381_),
    .B(_05380_),
    .A(_05378_));
 sg13g2_buf_1 _05890_ (.A(_05381_),
    .X(_05382_));
 sg13g2_buf_2 _05891_ (.A(\dtop.vtop.logo.addr[10] ),
    .X(_05383_));
 sg13g2_inv_1 _05892_ (.Y(_05384_),
    .A(_05383_));
 sg13g2_buf_2 _05893_ (.A(_00028_),
    .X(_05385_));
 sg13g2_inv_1 _05894_ (.Y(_05386_),
    .A(_05385_));
 sg13g2_buf_1 _05895_ (.A(net398),
    .X(_05387_));
 sg13g2_nand2_1 _05896_ (.Y(_05388_),
    .A(net351),
    .B(net208));
 sg13g2_o21ai_1 _05897_ (.B1(_05388_),
    .Y(_05389_),
    .A1(_05386_),
    .A2(_05213_));
 sg13g2_mux2_1 _05898_ (.A0(_05370_),
    .A1(_05389_),
    .S(net206),
    .X(_05390_));
 sg13g2_mux2_1 _05899_ (.A0(_05336_),
    .A1(_05390_),
    .S(net261),
    .X(_05391_));
 sg13g2_buf_1 _05900_ (.A(_05391_),
    .X(_05392_));
 sg13g2_nand2_1 _05901_ (.Y(_05393_),
    .A(net385),
    .B(_05392_));
 sg13g2_nor2_1 _05902_ (.A(_05384_),
    .B(_05392_),
    .Y(_05394_));
 sg13g2_a221oi_1 _05903_ (.B2(_05393_),
    .C1(_05394_),
    .B1(_05382_),
    .A1(net389),
    .Y(_05395_),
    .A2(_05288_));
 sg13g2_nor3_1 _05904_ (.A(net262),
    .B(_05287_),
    .C(_05395_),
    .Y(_05396_));
 sg13g2_buf_1 _05905_ (.A(_00029_),
    .X(_05397_));
 sg13g2_a22oi_1 _05906_ (.Y(_05398_),
    .B1(_05213_),
    .B2(net401),
    .A2(_05210_),
    .A1(_05397_));
 sg13g2_nand2_1 _05907_ (.Y(_05399_),
    .A(net206),
    .B(_05398_));
 sg13g2_o21ai_1 _05908_ (.B1(_05399_),
    .Y(_05400_),
    .A1(net206),
    .A2(_05389_));
 sg13g2_nor2_1 _05909_ (.A(net263),
    .B(_05400_),
    .Y(_05401_));
 sg13g2_a21oi_1 _05910_ (.A1(net263),
    .A2(_05371_),
    .Y(_05402_),
    .B1(_05401_));
 sg13g2_and2_1 _05911_ (.A(_05164_),
    .B(_05402_),
    .X(_05403_));
 sg13g2_buf_1 _05912_ (.A(_05403_),
    .X(_05404_));
 sg13g2_nand2_1 _05913_ (.Y(_05405_),
    .A(net426),
    .B(_05282_));
 sg13g2_inv_1 _05914_ (.Y(_05406_),
    .A(_05137_));
 sg13g2_nor3_1 _05915_ (.A(net390),
    .B(_05406_),
    .C(_05264_),
    .Y(_05407_));
 sg13g2_nor3_1 _05916_ (.A(_05194_),
    .B(_05405_),
    .C(_05407_),
    .Y(_05408_));
 sg13g2_and2_1 _05917_ (.A(_05404_),
    .B(_05408_),
    .X(_05409_));
 sg13g2_or2_1 _05918_ (.X(_05410_),
    .B(_05408_),
    .A(_05404_));
 sg13g2_o21ai_1 _05919_ (.B1(_05410_),
    .Y(_05411_),
    .A1(_05396_),
    .A2(_05409_));
 sg13g2_xnor2_1 _05920_ (.Y(_05412_),
    .A(_05260_),
    .B(_05411_));
 sg13g2_xnor2_1 _05921_ (.Y(_05413_),
    .A(_05404_),
    .B(_05408_));
 sg13g2_inv_1 _05922_ (.Y(_05414_),
    .A(_05413_));
 sg13g2_xnor2_1 _05923_ (.Y(_05415_),
    .A(_05396_),
    .B(_05414_));
 sg13g2_nand3_1 _05924_ (.B(_05382_),
    .C(_05394_),
    .A(net260),
    .Y(_05416_));
 sg13g2_a21o_1 _05925_ (.A2(_05285_),
    .A1(_05279_),
    .B1(_05416_),
    .X(_05417_));
 sg13g2_nor2_1 _05926_ (.A(_05279_),
    .B(_05285_),
    .Y(_05418_));
 sg13g2_inv_1 _05927_ (.Y(_05419_),
    .A(_05393_));
 sg13g2_nand2_1 _05928_ (.Y(_05420_),
    .A(_05364_),
    .B(_05374_));
 sg13g2_buf_1 _05929_ (.A(_05376_),
    .X(_05421_));
 sg13g2_nand2_1 _05930_ (.Y(_05422_),
    .A(net384),
    .B(_05364_));
 sg13g2_a22oi_1 _05931_ (.Y(_05423_),
    .B1(_05420_),
    .B2(_05422_),
    .A2(_05358_),
    .A1(_05353_));
 sg13g2_nor2_1 _05932_ (.A(_05380_),
    .B(_05423_),
    .Y(_05424_));
 sg13g2_a22oi_1 _05933_ (.Y(_05425_),
    .B1(_05419_),
    .B2(_05424_),
    .A2(_05392_),
    .A1(net262));
 sg13g2_a21oi_1 _05934_ (.A1(_05418_),
    .A2(_05425_),
    .Y(_05426_),
    .B1(_05414_));
 sg13g2_inv_1 _05935_ (.Y(_05427_),
    .A(_05287_));
 sg13g2_o21ai_1 _05936_ (.B1(_05427_),
    .Y(_00393_),
    .A1(_05271_),
    .A2(_05395_));
 sg13g2_a21oi_1 _05937_ (.A1(_05287_),
    .A2(_05425_),
    .Y(_00394_),
    .B1(_05413_));
 sg13g2_a221oi_1 _05938_ (.B2(_00394_),
    .C1(_05228_),
    .B1(_00393_),
    .A1(_05417_),
    .Y(_00395_),
    .A2(_05426_));
 sg13g2_a21oi_1 _05939_ (.A1(_05228_),
    .A2(_05415_),
    .Y(_00396_),
    .B1(_00395_));
 sg13g2_xnor2_1 _05940_ (.Y(_00397_),
    .A(_05412_),
    .B(_00396_));
 sg13g2_a21oi_1 _05941_ (.A1(net401),
    .A2(_00397_),
    .Y(_00398_),
    .B1(net390));
 sg13g2_nor2_1 _05942_ (.A(net305),
    .B(_00398_),
    .Y(_00399_));
 sg13g2_or4_1 _05943_ (.A(net402),
    .B(net390),
    .C(net393),
    .D(_05130_),
    .X(_00400_));
 sg13g2_buf_1 _05944_ (.A(_00400_),
    .X(_00401_));
 sg13g2_a21oi_1 _05945_ (.A1(net401),
    .A2(_00397_),
    .Y(_00402_),
    .B1(_00401_));
 sg13g2_inv_2 _05946_ (.Y(_00403_),
    .A(_05397_));
 sg13g2_o21ai_1 _05947_ (.B1(_05154_),
    .Y(_00404_),
    .A1(_05250_),
    .A2(_05148_));
 sg13g2_nor2_1 _05948_ (.A(net424),
    .B(_00404_),
    .Y(_00405_));
 sg13g2_inv_1 _05949_ (.Y(_00406_),
    .A(_05214_));
 sg13g2_buf_1 _05950_ (.A(_00406_),
    .X(_00407_));
 sg13g2_nand2b_1 _05951_ (.Y(_00408_),
    .B(_00407_),
    .A_N(_00404_));
 sg13g2_buf_1 _05952_ (.A(_00408_),
    .X(_00409_));
 sg13g2_nand2_1 _05953_ (.Y(_00410_),
    .A(\dtop.enable ),
    .B(_05193_));
 sg13g2_buf_2 _05954_ (.A(_05428_),
    .X(_00411_));
 sg13g2_inv_1 _05955_ (.Y(_00412_),
    .A(_05167_));
 sg13g2_nor2b_1 _05956_ (.A(net395),
    .B_N(_05174_),
    .Y(_00413_));
 sg13g2_nor2_1 _05957_ (.A(_05168_),
    .B(net329),
    .Y(_00414_));
 sg13g2_a221oi_1 _05958_ (.B2(_00413_),
    .C1(_00414_),
    .B1(_05180_),
    .A1(_00412_),
    .Y(_00415_),
    .A2(_05183_));
 sg13g2_a22oi_1 _05959_ (.Y(_00416_),
    .B1(_05186_),
    .B2(_00415_),
    .A2(net304),
    .A1(_05168_));
 sg13g2_buf_2 _05960_ (.A(_00416_),
    .X(_00417_));
 sg13g2_buf_8 _05961_ (.A(_05171_),
    .X(_00418_));
 sg13g2_buf_1 _05962_ (.A(net383),
    .X(_00419_));
 sg13g2_buf_1 _05963_ (.A(net349),
    .X(_00420_));
 sg13g2_buf_1 _05964_ (.A(_05183_),
    .X(_00421_));
 sg13g2_xnor2_1 _05965_ (.Y(_00422_),
    .A(net324),
    .B(net382));
 sg13g2_xor2_1 _05966_ (.B(_00422_),
    .A(_00417_),
    .X(_00423_));
 sg13g2_xnor2_1 _05967_ (.Y(_00424_),
    .A(_00411_),
    .B(_00423_));
 sg13g2_xor2_1 _05968_ (.B(_00424_),
    .A(_00410_),
    .X(_00425_));
 sg13g2_nor2_2 _05969_ (.A(_05221_),
    .B(net420),
    .Y(_00426_));
 sg13g2_nand2_1 _05970_ (.Y(_00427_),
    .A(net391),
    .B(_00064_));
 sg13g2_a22oi_1 _05971_ (.Y(_00428_),
    .B1(_00427_),
    .B2(net386),
    .A2(_00426_),
    .A1(_00425_));
 sg13g2_xnor2_1 _05972_ (.Y(_00429_),
    .A(_05303_),
    .B(_00428_));
 sg13g2_nor2_1 _05973_ (.A(_00409_),
    .B(_00429_),
    .Y(_00430_));
 sg13g2_or2_1 _05974_ (.X(_00431_),
    .B(_00430_),
    .A(_00405_));
 sg13g2_buf_2 _05975_ (.A(\dtop.player_inst.program_addr[0] ),
    .X(_00432_));
 sg13g2_buf_8 _05976_ (.A(_00432_),
    .X(_00433_));
 sg13g2_inv_1 _05977_ (.Y(_00434_),
    .A(net381));
 sg13g2_buf_1 _05978_ (.A(_00434_),
    .X(_00435_));
 sg13g2_o21ai_1 _05979_ (.B1(net354),
    .Y(_00436_),
    .A1(net323),
    .A2(_05298_));
 sg13g2_and2_1 _05980_ (.A(net429),
    .B(_00432_),
    .X(_00437_));
 sg13g2_buf_1 _05981_ (.A(_00437_),
    .X(_00438_));
 sg13g2_a22oi_1 _05982_ (.Y(_00439_),
    .B1(_00438_),
    .B2(_05314_),
    .A2(_00436_),
    .A1(_05301_));
 sg13g2_inv_1 _05983_ (.Y(_00440_),
    .A(_00439_));
 sg13g2_inv_2 _05984_ (.Y(_00441_),
    .A(net355));
 sg13g2_buf_1 _05985_ (.A(_00441_),
    .X(_00442_));
 sg13g2_a21oi_1 _05986_ (.A1(_05168_),
    .A2(_05174_),
    .Y(_00443_),
    .B1(_05183_));
 sg13g2_nor2_2 _05987_ (.A(net395),
    .B(_00443_),
    .Y(_00444_));
 sg13g2_xnor2_1 _05988_ (.Y(_00445_),
    .A(net300),
    .B(_00444_));
 sg13g2_xor2_1 _05989_ (.B(_00445_),
    .A(_00066_),
    .X(_00446_));
 sg13g2_nand2_1 _05990_ (.Y(_00447_),
    .A(net421),
    .B(_00445_));
 sg13g2_o21ai_1 _05991_ (.B1(_00447_),
    .Y(_00448_),
    .A1(_00440_),
    .A2(_00446_));
 sg13g2_buf_1 _05992_ (.A(_00065_),
    .X(_00449_));
 sg13g2_buf_1 _05993_ (.A(\dtop.enable ),
    .X(_00450_));
 sg13g2_xnor2_1 _05994_ (.Y(_00451_),
    .A(net419),
    .B(_05228_));
 sg13g2_nand2_1 _05995_ (.Y(_00452_),
    .A(_00449_),
    .B(_00451_));
 sg13g2_nor2_1 _05996_ (.A(_00449_),
    .B(_00451_),
    .Y(_00453_));
 sg13g2_a21oi_1 _05997_ (.A1(_00448_),
    .A2(_00452_),
    .Y(_00454_),
    .B1(_00453_));
 sg13g2_buf_1 _05998_ (.A(_00454_),
    .X(_00455_));
 sg13g2_nand2b_1 _05999_ (.Y(_00456_),
    .B(_00455_),
    .A_N(_00405_));
 sg13g2_xnor2_1 _06000_ (.Y(_00457_),
    .A(_00451_),
    .B(_00448_));
 sg13g2_xnor2_1 _06001_ (.Y(_00458_),
    .A(_00449_),
    .B(_00457_));
 sg13g2_buf_1 _06002_ (.A(net381),
    .X(_00459_));
 sg13g2_buf_1 _06003_ (.A(_00459_),
    .X(_00460_));
 sg13g2_buf_1 _06004_ (.A(net322),
    .X(_00461_));
 sg13g2_buf_1 _06005_ (.A(net299),
    .X(_00462_));
 sg13g2_xnor2_1 _06006_ (.Y(_00463_),
    .A(net287),
    .B(_05298_));
 sg13g2_buf_1 _06007_ (.A(net325),
    .X(_00464_));
 sg13g2_buf_1 _06008_ (.A(net298),
    .X(_00465_));
 sg13g2_xnor2_1 _06009_ (.Y(_00466_),
    .A(net422),
    .B(net286));
 sg13g2_buf_2 _06010_ (.A(_00014_),
    .X(_00467_));
 sg13g2_inv_1 _06011_ (.Y(_00468_),
    .A(_00467_));
 sg13g2_a21oi_1 _06012_ (.A1(_00463_),
    .A2(_00466_),
    .Y(_00469_),
    .B1(_00468_));
 sg13g2_xnor2_1 _06013_ (.Y(_00470_),
    .A(_00410_),
    .B(_00424_));
 sg13g2_inv_2 _06014_ (.Y(_00471_),
    .A(net420));
 sg13g2_nand2_1 _06015_ (.Y(_00472_),
    .A(net391),
    .B(_00471_));
 sg13g2_nand2_1 _06016_ (.Y(_00473_),
    .A(net386),
    .B(_00427_));
 sg13g2_o21ai_1 _06017_ (.B1(_00473_),
    .Y(_00474_),
    .A1(_00470_),
    .A2(_00472_));
 sg13g2_o21ai_1 _06018_ (.B1(_00474_),
    .Y(_00475_),
    .A1(_00458_),
    .A2(_00469_));
 sg13g2_o21ai_1 _06019_ (.B1(_00458_),
    .Y(_00476_),
    .A1(_00428_),
    .A2(_00469_));
 sg13g2_mux2_1 _06020_ (.A0(_00475_),
    .A1(_00476_),
    .S(_05324_),
    .X(_00477_));
 sg13g2_and3_1 _06021_ (.X(_00478_),
    .A(_00468_),
    .B(_00463_),
    .C(_00466_));
 sg13g2_nor2_1 _06022_ (.A(_05324_),
    .B(_00478_),
    .Y(_00479_));
 sg13g2_nor2_1 _06023_ (.A(net425),
    .B(_00478_),
    .Y(_00480_));
 sg13g2_a22oi_1 _06024_ (.Y(_00481_),
    .B1(_00480_),
    .B2(_00458_),
    .A2(_00479_),
    .A1(_00474_));
 sg13g2_nor2_1 _06025_ (.A(net425),
    .B(_00467_),
    .Y(_00482_));
 sg13g2_nor2_1 _06026_ (.A(_05324_),
    .B(_00467_),
    .Y(_00483_));
 sg13g2_a22oi_1 _06027_ (.Y(_00484_),
    .B1(_00483_),
    .B2(_00458_),
    .A2(_00482_),
    .A1(_00428_));
 sg13g2_xnor2_1 _06028_ (.Y(_00485_),
    .A(_00440_),
    .B(_00446_));
 sg13g2_a21o_1 _06029_ (.A2(_00484_),
    .A1(_00481_),
    .B1(_00485_),
    .X(_00486_));
 sg13g2_a21oi_1 _06030_ (.A1(_00477_),
    .A2(_00486_),
    .Y(_00487_),
    .B1(_00409_));
 sg13g2_a21oi_2 _06031_ (.B1(_00487_),
    .Y(_00488_),
    .A2(_00456_),
    .A1(_00431_));
 sg13g2_nor2_2 _06032_ (.A(_05221_),
    .B(_00471_),
    .Y(_00489_));
 sg13g2_o21ai_1 _06033_ (.B1(_00489_),
    .Y(_00490_),
    .A1(_00430_),
    .A2(_00456_));
 sg13g2_buf_1 _06034_ (.A(_00490_),
    .X(_00491_));
 sg13g2_nor3_2 _06035_ (.A(_05249_),
    .B(_00488_),
    .C(_00491_),
    .Y(_00492_));
 sg13g2_nor2_1 _06036_ (.A(_05250_),
    .B(_00403_),
    .Y(_00493_));
 sg13g2_buf_1 _06037_ (.A(_00487_),
    .X(_00494_));
 sg13g2_a21o_1 _06038_ (.A2(_00456_),
    .A1(_00431_),
    .B1(_00494_),
    .X(_00495_));
 sg13g2_inv_1 _06039_ (.Y(_00496_),
    .A(_00491_));
 sg13g2_nand2_1 _06040_ (.Y(_00497_),
    .A(_00495_),
    .B(_00496_));
 sg13g2_a221oi_1 _06041_ (.B2(_00497_),
    .C1(net288),
    .B1(_00493_),
    .A1(_00403_),
    .Y(_00498_),
    .A2(_00492_));
 sg13g2_buf_1 _06042_ (.A(_00498_),
    .X(_00499_));
 sg13g2_buf_1 _06043_ (.A(net60),
    .X(_00500_));
 sg13g2_buf_8 _06044_ (.A(\dtop.player_inst.program_addr[5] ),
    .X(_00501_));
 sg13g2_buf_1 _06045_ (.A(net418),
    .X(_00502_));
 sg13g2_inv_1 _06046_ (.Y(_00503_),
    .A(net380));
 sg13g2_buf_1 _06047_ (.A(_00503_),
    .X(_00504_));
 sg13g2_nand2_1 _06048_ (.Y(_00505_),
    .A(net321),
    .B(_00444_));
 sg13g2_nand2_1 _06049_ (.Y(_00506_),
    .A(net324),
    .B(_00421_));
 sg13g2_buf_1 _06050_ (.A(net324),
    .X(_00507_));
 sg13g2_nor2_1 _06051_ (.A(net297),
    .B(net382),
    .Y(_00508_));
 sg13g2_a21oi_2 _06052_ (.B1(_00508_),
    .Y(_00509_),
    .A2(_00506_),
    .A1(_00417_));
 sg13g2_nor2_1 _06053_ (.A(net321),
    .B(_00444_),
    .Y(_00510_));
 sg13g2_a21oi_2 _06054_ (.B1(_00510_),
    .Y(_00511_),
    .A2(_00509_),
    .A1(_00505_));
 sg13g2_buf_8 _06055_ (.A(\dtop.player_inst.program_addr[6] ),
    .X(_00512_));
 sg13g2_inv_2 _06056_ (.Y(_00513_),
    .A(net417));
 sg13g2_buf_1 _06057_ (.A(net379),
    .X(_00514_));
 sg13g2_inv_1 _06058_ (.Y(_00515_),
    .A(net382));
 sg13g2_buf_1 _06059_ (.A(_05168_),
    .X(_00516_));
 sg13g2_nand3b_1 _06060_ (.B(net378),
    .C(net395),
    .Y(_00517_),
    .A_N(_05184_));
 sg13g2_o21ai_1 _06061_ (.B1(_00517_),
    .Y(_00518_),
    .A1(_00515_),
    .A2(_05170_));
 sg13g2_xnor2_1 _06062_ (.Y(_00519_),
    .A(net346),
    .B(_00518_));
 sg13g2_nor2_1 _06063_ (.A(_00511_),
    .B(_00519_),
    .Y(_00520_));
 sg13g2_buf_1 _06064_ (.A(_00078_),
    .X(_00521_));
 sg13g2_buf_1 _06065_ (.A(net416),
    .X(_00522_));
 sg13g2_nor2_1 _06066_ (.A(net377),
    .B(_00518_),
    .Y(_00523_));
 sg13g2_nor2_2 _06067_ (.A(_00520_),
    .B(_00523_),
    .Y(_00524_));
 sg13g2_o21ai_1 _06068_ (.B1(net378),
    .Y(_00525_),
    .A1(_00412_),
    .A2(_05174_));
 sg13g2_and4_1 _06069_ (.A(_00412_),
    .B(net378),
    .C(_05174_),
    .D(_00515_),
    .X(_00526_));
 sg13g2_a21oi_2 _06070_ (.B1(_00526_),
    .Y(_00527_),
    .A2(_00525_),
    .A1(net382));
 sg13g2_xor2_1 _06071_ (.B(_00527_),
    .A(_00524_),
    .X(_00528_));
 sg13g2_buf_1 _06072_ (.A(_00528_),
    .X(_00529_));
 sg13g2_buf_1 _06073_ (.A(net137),
    .X(_00530_));
 sg13g2_buf_1 _06074_ (.A(net110),
    .X(_00531_));
 sg13g2_buf_1 _06075_ (.A(_00531_),
    .X(_00532_));
 sg13g2_xnor2_1 _06076_ (.Y(_00533_),
    .A(_00430_),
    .B(_00455_));
 sg13g2_buf_2 _06077_ (.A(_00533_),
    .X(_00534_));
 sg13g2_xor2_1 _06078_ (.B(_00534_),
    .A(net94),
    .X(_00535_));
 sg13g2_buf_1 _06079_ (.A(_00535_),
    .X(_00536_));
 sg13g2_xor2_1 _06080_ (.B(_00519_),
    .A(_00511_),
    .X(_00537_));
 sg13g2_buf_2 _06081_ (.A(_00537_),
    .X(_00538_));
 sg13g2_buf_1 _06082_ (.A(net380),
    .X(_00539_));
 sg13g2_xnor2_1 _06083_ (.Y(_00540_),
    .A(net345),
    .B(_00444_));
 sg13g2_xnor2_1 _06084_ (.Y(_00541_),
    .A(_00509_),
    .B(_00540_));
 sg13g2_nand3_1 _06085_ (.B(_05193_),
    .C(_00423_),
    .A(net419),
    .Y(_00542_));
 sg13g2_a21oi_1 _06086_ (.A1(net419),
    .A2(_05193_),
    .Y(_00543_),
    .B1(_00423_));
 sg13g2_a21o_1 _06087_ (.A2(_00542_),
    .A1(_00411_),
    .B1(_00543_),
    .X(_00544_));
 sg13g2_buf_2 _06088_ (.A(_00544_),
    .X(_00545_));
 sg13g2_nor2_1 _06089_ (.A(_00541_),
    .B(_00545_),
    .Y(_00546_));
 sg13g2_buf_1 _06090_ (.A(_00546_),
    .X(_00547_));
 sg13g2_nand2_1 _06091_ (.Y(_00548_),
    .A(_00538_),
    .B(net136));
 sg13g2_xnor2_1 _06092_ (.Y(_00549_),
    .A(_00511_),
    .B(_00519_));
 sg13g2_xor2_1 _06093_ (.B(_00540_),
    .A(_00509_),
    .X(_00550_));
 sg13g2_buf_1 _06094_ (.A(_00550_),
    .X(_00551_));
 sg13g2_a21oi_1 _06095_ (.A1(_00411_),
    .A2(_00542_),
    .Y(_00552_),
    .B1(_00543_));
 sg13g2_nand2_1 _06096_ (.Y(_00553_),
    .A(_00551_),
    .B(_00552_));
 sg13g2_nand2_1 _06097_ (.Y(_00554_),
    .A(_00549_),
    .B(_00553_));
 sg13g2_buf_2 _06098_ (.A(_00554_),
    .X(_00555_));
 sg13g2_nand2_1 _06099_ (.Y(_00556_),
    .A(_00548_),
    .B(_00555_));
 sg13g2_buf_2 _06100_ (.A(_00556_),
    .X(_00557_));
 sg13g2_nor2_1 _06101_ (.A(_00536_),
    .B(_00557_),
    .Y(_00558_));
 sg13g2_buf_1 _06102_ (.A(_00552_),
    .X(_00559_));
 sg13g2_nor2_1 _06103_ (.A(_00551_),
    .B(net205),
    .Y(_00560_));
 sg13g2_buf_1 _06104_ (.A(_00560_),
    .X(_00561_));
 sg13g2_nor2_1 _06105_ (.A(net135),
    .B(_00546_),
    .Y(_00562_));
 sg13g2_buf_1 _06106_ (.A(_00562_),
    .X(_00563_));
 sg13g2_nor2_2 _06107_ (.A(net92),
    .B(_00557_),
    .Y(_00564_));
 sg13g2_xnor2_1 _06108_ (.Y(_00565_),
    .A(net94),
    .B(_00534_));
 sg13g2_buf_1 _06109_ (.A(_00565_),
    .X(_00566_));
 sg13g2_buf_8 _06110_ (.A(net72),
    .X(_00567_));
 sg13g2_xnor2_1 _06111_ (.Y(_00568_),
    .A(_00524_),
    .B(_00527_));
 sg13g2_buf_1 _06112_ (.A(_00568_),
    .X(_00569_));
 sg13g2_buf_1 _06113_ (.A(_00549_),
    .X(_00570_));
 sg13g2_buf_1 _06114_ (.A(_00553_),
    .X(_00571_));
 sg13g2_nor2_2 _06115_ (.A(net204),
    .B(net172),
    .Y(_00572_));
 sg13g2_xnor2_1 _06116_ (.Y(_00573_),
    .A(_00569_),
    .B(_00572_));
 sg13g2_buf_1 _06117_ (.A(_00573_),
    .X(_00574_));
 sg13g2_nor2_1 _06118_ (.A(_00567_),
    .B(net91),
    .Y(_00575_));
 sg13g2_buf_1 _06119_ (.A(_00425_),
    .X(_00576_));
 sg13g2_buf_1 _06120_ (.A(net203),
    .X(_00577_));
 sg13g2_buf_1 _06121_ (.A(net171),
    .X(_00578_));
 sg13g2_buf_1 _06122_ (.A(net134),
    .X(_00579_));
 sg13g2_buf_1 _06123_ (.A(net109),
    .X(_00580_));
 sg13g2_buf_1 _06124_ (.A(net67),
    .X(_00581_));
 sg13g2_xnor2_1 _06125_ (.Y(_00582_),
    .A(net137),
    .B(_00572_));
 sg13g2_buf_1 _06126_ (.A(_00582_),
    .X(_00583_));
 sg13g2_buf_1 _06127_ (.A(net89),
    .X(_00584_));
 sg13g2_buf_1 _06128_ (.A(_00538_),
    .X(_00585_));
 sg13g2_nand2_1 _06129_ (.Y(_00586_),
    .A(_00541_),
    .B(_00545_));
 sg13g2_buf_1 _06130_ (.A(_00586_),
    .X(_00587_));
 sg13g2_nand2_1 _06131_ (.Y(_00588_),
    .A(net133),
    .B(net172));
 sg13g2_buf_1 _06132_ (.A(_00588_),
    .X(_00589_));
 sg13g2_nor2_1 _06133_ (.A(_00585_),
    .B(_00589_),
    .Y(_00590_));
 sg13g2_buf_1 _06134_ (.A(_00590_),
    .X(_00591_));
 sg13g2_o21ai_1 _06135_ (.B1(net71),
    .Y(_00592_),
    .A1(net59),
    .A2(net79));
 sg13g2_nand2_1 _06136_ (.Y(_00593_),
    .A(net90),
    .B(_00592_));
 sg13g2_a221oi_1 _06137_ (.B2(_00575_),
    .C1(_00593_),
    .B1(_00564_),
    .A1(net80),
    .Y(_00594_),
    .A2(_00558_));
 sg13g2_buf_1 _06138_ (.A(_00589_),
    .X(_00595_));
 sg13g2_buf_1 _06139_ (.A(net78),
    .X(_00596_));
 sg13g2_buf_1 _06140_ (.A(net70),
    .X(_00597_));
 sg13g2_nor2_2 _06141_ (.A(_00536_),
    .B(net91),
    .Y(_00598_));
 sg13g2_nor2_1 _06142_ (.A(_00538_),
    .B(_00546_),
    .Y(_00599_));
 sg13g2_buf_2 _06143_ (.A(_00599_),
    .X(_00600_));
 sg13g2_nor2_1 _06144_ (.A(_00572_),
    .B(_00600_),
    .Y(_00601_));
 sg13g2_buf_1 _06145_ (.A(_00601_),
    .X(_00602_));
 sg13g2_nor2_2 _06146_ (.A(net77),
    .B(net89),
    .Y(_00603_));
 sg13g2_o21ai_1 _06147_ (.B1(net78),
    .Y(_00604_),
    .A1(_00557_),
    .A2(net91));
 sg13g2_nand2b_1 _06148_ (.Y(_00605_),
    .B(_00604_),
    .A_N(_00603_));
 sg13g2_buf_1 _06149_ (.A(net73),
    .X(_00606_));
 sg13g2_buf_1 _06150_ (.A(net65),
    .X(_00607_));
 sg13g2_nand2_1 _06151_ (.Y(_00608_),
    .A(net204),
    .B(_00562_));
 sg13g2_buf_2 _06152_ (.A(_00608_),
    .X(_00609_));
 sg13g2_buf_1 _06153_ (.A(_00470_),
    .X(_00610_));
 sg13g2_buf_1 _06154_ (.A(net202),
    .X(_00611_));
 sg13g2_buf_1 _06155_ (.A(net169),
    .X(_00612_));
 sg13g2_buf_1 _06156_ (.A(net132),
    .X(_00613_));
 sg13g2_o21ai_1 _06157_ (.B1(net108),
    .Y(_00614_),
    .A1(net58),
    .A2(_00609_));
 sg13g2_a221oi_1 _06158_ (.B2(net58),
    .C1(_00614_),
    .B1(_00605_),
    .A1(net66),
    .Y(_00615_),
    .A2(_00598_));
 sg13g2_nor3_1 _06159_ (.A(net51),
    .B(_00594_),
    .C(_00615_),
    .Y(_00616_));
 sg13g2_nor2_2 _06160_ (.A(net203),
    .B(_00589_),
    .Y(_00617_));
 sg13g2_nand3_1 _06161_ (.B(_00495_),
    .C(_00496_),
    .A(_05249_),
    .Y(_00618_));
 sg13g2_buf_1 _06162_ (.A(_00618_),
    .X(_00619_));
 sg13g2_nor2_1 _06163_ (.A(_05249_),
    .B(net288),
    .Y(_00620_));
 sg13g2_o21ai_1 _06164_ (.B1(_00620_),
    .Y(_00621_),
    .A1(_00488_),
    .A2(_00491_));
 sg13g2_buf_1 _06165_ (.A(_00621_),
    .X(_00622_));
 sg13g2_and2_1 _06166_ (.A(_00619_),
    .B(_00622_),
    .X(_00623_));
 sg13g2_buf_2 _06167_ (.A(_00623_),
    .X(_00624_));
 sg13g2_nand2_2 _06168_ (.Y(_00625_),
    .A(_00557_),
    .B(_00583_));
 sg13g2_nor3_2 _06169_ (.A(_00403_),
    .B(_00624_),
    .C(_00625_),
    .Y(_00626_));
 sg13g2_and2_1 _06170_ (.A(_00617_),
    .B(_00626_),
    .X(_00627_));
 sg13g2_nand4_1 _06171_ (.B(_00602_),
    .C(_00574_),
    .A(_05148_),
    .Y(_00628_),
    .D(_00617_));
 sg13g2_buf_1 _06172_ (.A(_05397_),
    .X(_00629_));
 sg13g2_nor2_1 _06173_ (.A(_05250_),
    .B(net376),
    .Y(_00630_));
 sg13g2_a22oi_1 _06174_ (.Y(_00631_),
    .B1(_00630_),
    .B2(_00497_),
    .A2(_00492_),
    .A1(net376));
 sg13g2_or2_1 _06175_ (.X(_00632_),
    .B(_00631_),
    .A(_00628_));
 sg13g2_buf_1 _06176_ (.A(_00632_),
    .X(_00633_));
 sg13g2_nor2_1 _06177_ (.A(net77),
    .B(_00573_),
    .Y(_00634_));
 sg13g2_a21oi_2 _06178_ (.B1(net376),
    .Y(_00635_),
    .A2(_00622_),
    .A1(_00619_));
 sg13g2_and2_1 _06179_ (.A(_00634_),
    .B(_00635_),
    .X(_00636_));
 sg13g2_buf_2 _06180_ (.A(_00636_),
    .X(_00637_));
 sg13g2_buf_1 _06181_ (.A(net92),
    .X(_00638_));
 sg13g2_nor2_1 _06182_ (.A(net203),
    .B(net73),
    .Y(_00639_));
 sg13g2_buf_1 _06183_ (.A(_00639_),
    .X(_00640_));
 sg13g2_nor2_1 _06184_ (.A(_00638_),
    .B(_00640_),
    .Y(_00641_));
 sg13g2_buf_1 _06185_ (.A(net387),
    .X(_00642_));
 sg13g2_a21oi_1 _06186_ (.A1(_00637_),
    .A2(_00641_),
    .Y(_00643_),
    .B1(net344));
 sg13g2_nand3b_1 _06187_ (.B(_00633_),
    .C(_00643_),
    .Y(_00644_),
    .A_N(_00627_));
 sg13g2_nor2_1 _06188_ (.A(_05359_),
    .B(_05376_),
    .Y(_00645_));
 sg13g2_o21ai_1 _06189_ (.B1(_00645_),
    .Y(_00646_),
    .A1(_00616_),
    .A2(_00644_));
 sg13g2_nor4_1 _06190_ (.A(_05249_),
    .B(net376),
    .C(_00488_),
    .D(_00491_),
    .Y(_00647_));
 sg13g2_o21ai_1 _06191_ (.B1(_00493_),
    .Y(_00648_),
    .A1(_00488_),
    .A2(_00491_));
 sg13g2_nand3b_1 _06192_ (.B(_00648_),
    .C(_05148_),
    .Y(_00649_),
    .A_N(_00647_));
 sg13g2_buf_1 _06193_ (.A(_00649_),
    .X(_00650_));
 sg13g2_buf_1 _06194_ (.A(_00650_),
    .X(_00651_));
 sg13g2_buf_1 _06195_ (.A(net56),
    .X(_00652_));
 sg13g2_nand2_1 _06196_ (.Y(_00653_),
    .A(_00610_),
    .B(net72));
 sg13g2_buf_1 _06197_ (.A(_00653_),
    .X(_00654_));
 sg13g2_nor2_2 _06198_ (.A(_00538_),
    .B(_00587_),
    .Y(_00655_));
 sg13g2_nor2_1 _06199_ (.A(net73),
    .B(net89),
    .Y(_00656_));
 sg13g2_nand2_1 _06200_ (.Y(_00657_),
    .A(net73),
    .B(net89));
 sg13g2_nand2b_1 _06201_ (.Y(_00658_),
    .B(_00657_),
    .A_N(_00656_));
 sg13g2_buf_1 _06202_ (.A(net109),
    .X(_00659_));
 sg13g2_nor2_2 _06203_ (.A(net204),
    .B(net135),
    .Y(_00660_));
 sg13g2_o21ai_1 _06204_ (.B1(_00660_),
    .Y(_00661_),
    .A1(_00571_),
    .A2(net55));
 sg13g2_o21ai_1 _06205_ (.B1(_00661_),
    .Y(_00662_),
    .A1(net88),
    .A2(_00658_));
 sg13g2_a221oi_1 _06206_ (.B2(net88),
    .C1(_00662_),
    .B1(_00658_),
    .A1(net55),
    .Y(_00663_),
    .A2(_00655_));
 sg13g2_nand2_1 _06207_ (.Y(_00664_),
    .A(_00619_),
    .B(_00622_));
 sg13g2_buf_1 _06208_ (.A(_00664_),
    .X(_00665_));
 sg13g2_buf_1 _06209_ (.A(_00634_),
    .X(_00666_));
 sg13g2_nor2_1 _06210_ (.A(net202),
    .B(_00565_),
    .Y(_00667_));
 sg13g2_buf_1 _06211_ (.A(_00667_),
    .X(_00668_));
 sg13g2_nand3_1 _06212_ (.B(net64),
    .C(_00668_),
    .A(net49),
    .Y(_00669_));
 sg13g2_buf_1 _06213_ (.A(net72),
    .X(_00670_));
 sg13g2_buf_1 _06214_ (.A(net62),
    .X(_00671_));
 sg13g2_nor2_1 _06215_ (.A(net54),
    .B(_00609_),
    .Y(_00672_));
 sg13g2_buf_1 _06216_ (.A(net65),
    .X(_00673_));
 sg13g2_buf_1 _06217_ (.A(net204),
    .X(_00674_));
 sg13g2_nor4_1 _06218_ (.A(_00673_),
    .B(_00674_),
    .C(_00571_),
    .D(_00624_),
    .Y(_00675_));
 sg13g2_o21ai_1 _06219_ (.B1(net80),
    .Y(_00676_),
    .A1(_00672_),
    .A2(_00675_));
 sg13g2_nor2_1 _06220_ (.A(_00569_),
    .B(_00609_),
    .Y(_00677_));
 sg13g2_nand2_1 _06221_ (.Y(_00678_),
    .A(net88),
    .B(_00677_));
 sg13g2_nor2_1 _06222_ (.A(net137),
    .B(net73),
    .Y(_00679_));
 sg13g2_buf_2 _06223_ (.A(_00679_),
    .X(_00680_));
 sg13g2_nand3_1 _06224_ (.B(net49),
    .C(_00655_),
    .A(_00680_),
    .Y(_00681_));
 sg13g2_nand4_1 _06225_ (.B(_00676_),
    .C(_00678_),
    .A(_00669_),
    .Y(_00682_),
    .D(_00681_));
 sg13g2_nor2_1 _06226_ (.A(net376),
    .B(net288),
    .Y(_00683_));
 sg13g2_nor2_1 _06227_ (.A(_00403_),
    .B(net288),
    .Y(_00684_));
 sg13g2_mux2_1 _06228_ (.A0(_00683_),
    .A1(_00684_),
    .S(_00492_),
    .X(_00685_));
 sg13g2_buf_1 _06229_ (.A(_00685_),
    .X(_00686_));
 sg13g2_buf_1 _06230_ (.A(_00686_),
    .X(_00687_));
 sg13g2_buf_1 _06231_ (.A(net344),
    .X(_00688_));
 sg13g2_nand2_1 _06232_ (.Y(_00689_),
    .A(_00629_),
    .B(_00664_));
 sg13g2_nand2_2 _06233_ (.Y(_00690_),
    .A(net73),
    .B(net92));
 sg13g2_nor2_1 _06234_ (.A(net109),
    .B(_00625_),
    .Y(_00691_));
 sg13g2_nand2_1 _06235_ (.Y(_00692_),
    .A(net65),
    .B(net91));
 sg13g2_o21ai_1 _06236_ (.B1(_00692_),
    .Y(_00693_),
    .A1(net132),
    .A2(_00598_));
 sg13g2_a22oi_1 _06237_ (.Y(_00694_),
    .B1(_00693_),
    .B2(net71),
    .A2(_00691_),
    .A1(_00690_));
 sg13g2_or2_1 _06238_ (.X(_00695_),
    .B(_00694_),
    .A(_00689_));
 sg13g2_nand3_1 _06239_ (.B(_00633_),
    .C(_00695_),
    .A(net320),
    .Y(_00696_));
 sg13g2_a221oi_1 _06240_ (.B2(net52),
    .C1(_00696_),
    .B1(_00682_),
    .A1(net50),
    .Y(_00697_),
    .A2(_00663_));
 sg13g2_nor2_1 _06241_ (.A(_00646_),
    .B(_00697_),
    .Y(_00698_));
 sg13g2_buf_1 _06242_ (.A(_00624_),
    .X(_00699_));
 sg13g2_and2_1 _06243_ (.A(_00634_),
    .B(_00686_),
    .X(_00700_));
 sg13g2_buf_2 _06244_ (.A(_00700_),
    .X(_00701_));
 sg13g2_nand2_1 _06245_ (.Y(_00702_),
    .A(net41),
    .B(_00701_));
 sg13g2_nand2_1 _06246_ (.Y(_00703_),
    .A(net72),
    .B(net78));
 sg13g2_nand3_1 _06247_ (.B(_00701_),
    .C(_00703_),
    .A(net41),
    .Y(_00704_));
 sg13g2_nand2_1 _06248_ (.Y(_00705_),
    .A(net64),
    .B(_00635_));
 sg13g2_a221oi_1 _06249_ (.B2(_00705_),
    .C1(net63),
    .B1(_00704_),
    .A1(_00638_),
    .Y(_00706_),
    .A2(_00702_));
 sg13g2_a21oi_1 _06250_ (.A1(net169),
    .A2(_00680_),
    .Y(_00707_),
    .B1(_00667_));
 sg13g2_o21ai_1 _06251_ (.B1(net76),
    .Y(_00708_),
    .A1(net170),
    .A2(net57));
 sg13g2_nand2_2 _06252_ (.Y(_00709_),
    .A(net110),
    .B(net73));
 sg13g2_buf_1 _06253_ (.A(_00572_),
    .X(_00710_));
 sg13g2_nand2_1 _06254_ (.Y(_00711_),
    .A(net110),
    .B(_00600_));
 sg13g2_o21ai_1 _06255_ (.B1(net134),
    .Y(_00712_),
    .A1(net93),
    .A2(_00600_));
 sg13g2_nand2_1 _06256_ (.Y(_00713_),
    .A(_00711_),
    .B(_00712_));
 sg13g2_a22oi_1 _06257_ (.Y(_00714_),
    .B1(_00713_),
    .B2(net66),
    .A2(net107),
    .A1(_00709_));
 sg13g2_nand3_1 _06258_ (.B(_00708_),
    .C(_00714_),
    .A(_00707_),
    .Y(_00715_));
 sg13g2_buf_1 _06259_ (.A(_00557_),
    .X(_00716_));
 sg13g2_nand2_1 _06260_ (.Y(_00717_),
    .A(_00576_),
    .B(_00589_));
 sg13g2_nor3_2 _06261_ (.A(net69),
    .B(net89),
    .C(_00717_),
    .Y(_00718_));
 sg13g2_buf_8 _06262_ (.A(net73),
    .X(_00719_));
 sg13g2_nand2_1 _06263_ (.Y(_00720_),
    .A(net169),
    .B(net61));
 sg13g2_nor2_1 _06264_ (.A(net203),
    .B(_00562_),
    .Y(_00721_));
 sg13g2_nand2_1 _06265_ (.Y(_00722_),
    .A(_00576_),
    .B(net92));
 sg13g2_nor2_1 _06266_ (.A(_00566_),
    .B(_00722_),
    .Y(_00723_));
 sg13g2_o21ai_1 _06267_ (.B1(_00666_),
    .Y(_00724_),
    .A1(_00721_),
    .A2(_00723_));
 sg13g2_a21oi_1 _06268_ (.A1(_00664_),
    .A2(_00724_),
    .Y(_00725_),
    .B1(net52));
 sg13g2_a221oi_1 _06269_ (.B2(_00677_),
    .C1(_00725_),
    .B1(_00720_),
    .A1(net58),
    .Y(_00726_),
    .A2(_00718_));
 sg13g2_a21oi_1 _06270_ (.A1(net50),
    .A2(_00715_),
    .Y(_00727_),
    .B1(_00726_));
 sg13g2_nor2_1 _06271_ (.A(_00610_),
    .B(_00595_),
    .Y(_00728_));
 sg13g2_nand2_2 _06272_ (.Y(_00729_),
    .A(net61),
    .B(_00728_));
 sg13g2_inv_2 _06273_ (.Y(_00730_),
    .A(_05354_));
 sg13g2_nor2_1 _06274_ (.A(net384),
    .B(_00730_),
    .Y(_00731_));
 sg13g2_o21ai_1 _06275_ (.B1(_00731_),
    .Y(_00732_),
    .A1(_00705_),
    .A2(_00729_));
 sg13g2_nor3_1 _06276_ (.A(_00706_),
    .B(_00727_),
    .C(_00732_),
    .Y(_00733_));
 sg13g2_buf_1 _06277_ (.A(net77),
    .X(_00734_));
 sg13g2_nor2_1 _06278_ (.A(net169),
    .B(net61),
    .Y(_00735_));
 sg13g2_o21ai_1 _06279_ (.B1(net76),
    .Y(_00736_),
    .A1(net68),
    .A2(_00735_));
 sg13g2_buf_1 _06280_ (.A(net169),
    .X(_00737_));
 sg13g2_nand3_1 _06281_ (.B(net53),
    .C(_00604_),
    .A(net131),
    .Y(_00738_));
 sg13g2_nor2_2 _06282_ (.A(net92),
    .B(net77),
    .Y(_00739_));
 sg13g2_o21ai_1 _06283_ (.B1(net109),
    .Y(_00740_),
    .A1(_00598_),
    .A2(_00739_));
 sg13g2_nand3_1 _06284_ (.B(_00738_),
    .C(_00740_),
    .A(_00736_),
    .Y(_00741_));
 sg13g2_nor2_1 _06285_ (.A(net171),
    .B(_00583_),
    .Y(_00742_));
 sg13g2_nand3_1 _06286_ (.B(net71),
    .C(_00742_),
    .A(net61),
    .Y(_00743_));
 sg13g2_buf_1 _06287_ (.A(_00569_),
    .X(_00744_));
 sg13g2_nor3_2 _06288_ (.A(_00744_),
    .B(_00660_),
    .C(_00655_),
    .Y(_00745_));
 sg13g2_nand3_1 _06289_ (.B(_00566_),
    .C(_00745_),
    .A(net134),
    .Y(_00746_));
 sg13g2_nand2_1 _06290_ (.Y(_00747_),
    .A(_00743_),
    .B(_00746_));
 sg13g2_nand2_1 _06291_ (.Y(_00748_),
    .A(net60),
    .B(_00747_));
 sg13g2_o21ai_1 _06292_ (.B1(_00748_),
    .Y(_00749_),
    .A1(net51),
    .A2(_00741_));
 sg13g2_nand2_2 _06293_ (.Y(_00750_),
    .A(net67),
    .B(net92));
 sg13g2_xnor2_1 _06294_ (.Y(_00751_),
    .A(net131),
    .B(_00750_));
 sg13g2_and2_1 _06295_ (.A(_00626_),
    .B(_00751_),
    .X(_00752_));
 sg13g2_a21oi_2 _06296_ (.B1(net169),
    .Y(_00753_),
    .A2(_00595_),
    .A1(net67));
 sg13g2_and2_1 _06297_ (.A(_00637_),
    .B(_00753_),
    .X(_00754_));
 sg13g2_buf_1 _06298_ (.A(net384),
    .X(_00755_));
 sg13g2_buf_1 _06299_ (.A(_00730_),
    .X(_00756_));
 sg13g2_nand2_1 _06300_ (.Y(_00757_),
    .A(net67),
    .B(_00721_));
 sg13g2_nand2_1 _06301_ (.Y(_00758_),
    .A(_00729_),
    .B(_00757_));
 sg13g2_nand3_1 _06302_ (.B(_00701_),
    .C(_00758_),
    .A(_00699_),
    .Y(_00759_));
 sg13g2_nand3_1 _06303_ (.B(net319),
    .C(_00759_),
    .A(net343),
    .Y(_00760_));
 sg13g2_nor4_1 _06304_ (.A(_00749_),
    .B(_00752_),
    .C(_00754_),
    .D(_00760_),
    .Y(_00761_));
 sg13g2_buf_1 _06305_ (.A(net91),
    .X(_00762_));
 sg13g2_a22oi_1 _06306_ (.Y(_00763_),
    .B1(_00739_),
    .B2(net53),
    .A2(_00558_),
    .A1(net131));
 sg13g2_nor2_1 _06307_ (.A(net75),
    .B(_00763_),
    .Y(_00764_));
 sg13g2_o21ai_1 _06308_ (.B1(_00579_),
    .Y(_00765_),
    .A1(net53),
    .A2(_00739_));
 sg13g2_nand3_1 _06309_ (.B(_00708_),
    .C(_00765_),
    .A(net344),
    .Y(_00766_));
 sg13g2_o21ai_1 _06310_ (.B1(net50),
    .Y(_00767_),
    .A1(_00764_),
    .A2(_00766_));
 sg13g2_nand2_1 _06311_ (.Y(_00768_),
    .A(_00690_),
    .B(net55));
 sg13g2_nand2_1 _06312_ (.Y(_00769_),
    .A(_00626_),
    .B(_00768_));
 sg13g2_nand2_1 _06313_ (.Y(_00770_),
    .A(_00611_),
    .B(net71));
 sg13g2_nand3_1 _06314_ (.B(_00719_),
    .C(_00564_),
    .A(net134),
    .Y(_00771_));
 sg13g2_o21ai_1 _06315_ (.B1(_00771_),
    .Y(_00772_),
    .A1(net65),
    .A2(_00770_));
 sg13g2_nand2_1 _06316_ (.Y(_00773_),
    .A(net75),
    .B(_00772_));
 sg13g2_nand3_1 _06317_ (.B(_00769_),
    .C(_00773_),
    .A(net51),
    .Y(_00774_));
 sg13g2_nand2_1 _06318_ (.Y(_00775_),
    .A(net49),
    .B(net55));
 sg13g2_a221oi_1 _06319_ (.B2(net66),
    .C1(net63),
    .B1(_00775_),
    .A1(_00617_),
    .Y(_00776_),
    .A2(net49));
 sg13g2_nand2_1 _06320_ (.Y(_00777_),
    .A(net343),
    .B(_00688_));
 sg13g2_a221oi_1 _06321_ (.B2(_00701_),
    .C1(_00777_),
    .B1(_00776_),
    .A1(_00767_),
    .Y(_00778_),
    .A2(_00774_));
 sg13g2_buf_1 _06322_ (.A(_05359_),
    .X(_00779_));
 sg13g2_nand3_1 _06323_ (.B(_00690_),
    .C(_00637_),
    .A(net88),
    .Y(_00780_));
 sg13g2_nand3_1 _06324_ (.B(_00701_),
    .C(_00768_),
    .A(net41),
    .Y(_00781_));
 sg13g2_nor2_1 _06325_ (.A(_00577_),
    .B(net77),
    .Y(_00782_));
 sg13g2_nor2_1 _06326_ (.A(_00564_),
    .B(net71),
    .Y(_00783_));
 sg13g2_nand2_1 _06327_ (.Y(_00784_),
    .A(net134),
    .B(_00719_));
 sg13g2_nor2_1 _06328_ (.A(_00783_),
    .B(_00784_),
    .Y(_00785_));
 sg13g2_a221oi_1 _06329_ (.B2(net55),
    .C1(_00785_),
    .B1(_00745_),
    .A1(net59),
    .Y(_00786_),
    .A2(_00782_));
 sg13g2_a21oi_1 _06330_ (.A1(_00567_),
    .A2(_00564_),
    .Y(_00787_),
    .B1(_00591_));
 sg13g2_nor2_1 _06331_ (.A(net57),
    .B(_00787_),
    .Y(_00788_));
 sg13g2_a21oi_1 _06332_ (.A1(net75),
    .A2(_00788_),
    .Y(_00789_),
    .B1(net56));
 sg13g2_a21o_1 _06333_ (.A2(_00786_),
    .A1(net56),
    .B1(_00789_),
    .X(_00790_));
 sg13g2_nor2_1 _06334_ (.A(_00597_),
    .B(net63),
    .Y(_00791_));
 sg13g2_or2_1 _06335_ (.X(_00792_),
    .B(net387),
    .A(_05421_));
 sg13g2_a21oi_1 _06336_ (.A1(_00626_),
    .A2(_00791_),
    .Y(_00793_),
    .B1(_00792_));
 sg13g2_nand4_1 _06337_ (.B(_00781_),
    .C(_00790_),
    .A(_00780_),
    .Y(_00794_),
    .D(_00793_));
 sg13g2_nand2_1 _06338_ (.Y(_00795_),
    .A(net375),
    .B(_00794_));
 sg13g2_nor4_1 _06339_ (.A(_00733_),
    .B(_00761_),
    .C(_00778_),
    .D(_00795_),
    .Y(_00796_));
 sg13g2_a21oi_1 _06340_ (.A1(net91),
    .A2(_00639_),
    .Y(_00797_),
    .B1(net68));
 sg13g2_nor2_1 _06341_ (.A(net70),
    .B(_00797_),
    .Y(_00798_));
 sg13g2_buf_1 _06342_ (.A(net106),
    .X(_00799_));
 sg13g2_buf_1 _06343_ (.A(net87),
    .X(_00800_));
 sg13g2_nor2_1 _06344_ (.A(_00670_),
    .B(net78),
    .Y(_00801_));
 sg13g2_a22oi_1 _06345_ (.Y(_00802_),
    .B1(_00656_),
    .B2(net68),
    .A2(_00801_),
    .A1(_00800_));
 sg13g2_nand3_1 _06346_ (.B(net68),
    .C(net75),
    .A(net58),
    .Y(_00803_));
 sg13g2_a221oi_1 _06347_ (.B2(net59),
    .C1(net131),
    .B1(net64),
    .A1(_00596_),
    .Y(_00804_),
    .A2(net69));
 sg13g2_a22oi_1 _06348_ (.Y(_00805_),
    .B1(_00803_),
    .B2(_00804_),
    .A2(_00802_),
    .A1(net108));
 sg13g2_nor3_1 _06349_ (.A(_00500_),
    .B(_00798_),
    .C(_00805_),
    .Y(_00806_));
 sg13g2_nor2_1 _06350_ (.A(_00744_),
    .B(net78),
    .Y(_00807_));
 sg13g2_nor2_1 _06351_ (.A(net93),
    .B(net92),
    .Y(_00808_));
 sg13g2_a22oi_1 _06352_ (.Y(_00809_),
    .B1(_00808_),
    .B2(_00600_),
    .A2(_00807_),
    .A1(net62));
 sg13g2_nand2_1 _06353_ (.Y(_00810_),
    .A(net110),
    .B(net136));
 sg13g2_o21ai_1 _06354_ (.B1(_00810_),
    .Y(_00811_),
    .A1(net110),
    .A2(_00555_));
 sg13g2_nor2_2 _06355_ (.A(net202),
    .B(_00563_),
    .Y(_00812_));
 sg13g2_nor2_1 _06356_ (.A(net171),
    .B(net172),
    .Y(_00813_));
 sg13g2_a21o_1 _06357_ (.A2(_00812_),
    .A1(net61),
    .B1(_00813_),
    .X(_00814_));
 sg13g2_nor2_1 _06358_ (.A(_00569_),
    .B(net204),
    .Y(_00815_));
 sg13g2_and2_1 _06359_ (.A(net72),
    .B(_00677_),
    .X(_00816_));
 sg13g2_buf_1 _06360_ (.A(_00816_),
    .X(_00817_));
 sg13g2_a221oi_1 _06361_ (.B2(_00815_),
    .C1(_00817_),
    .B1(_00814_),
    .A1(net63),
    .Y(_00818_),
    .A2(_00811_));
 sg13g2_o21ai_1 _06362_ (.B1(_00818_),
    .Y(_00819_),
    .A1(net90),
    .A2(_00809_));
 sg13g2_nor2_1 _06363_ (.A(net67),
    .B(net92),
    .Y(_00820_));
 sg13g2_a21oi_1 _06364_ (.A1(_00612_),
    .A2(_00820_),
    .Y(_00821_),
    .B1(_00735_));
 sg13g2_nor2_1 _06365_ (.A(_00624_),
    .B(_00821_),
    .Y(_00822_));
 sg13g2_a22oi_1 _06366_ (.Y(_00823_),
    .B1(_00822_),
    .B2(net64),
    .A2(_00819_),
    .A1(net41));
 sg13g2_nor2b_1 _06367_ (.A(_00823_),
    .B_N(net52),
    .Y(_00824_));
 sg13g2_a21oi_1 _06368_ (.A1(net58),
    .A2(_00718_),
    .Y(_00825_),
    .B1(_00817_));
 sg13g2_o21ai_1 _06369_ (.B1(net319),
    .Y(_00826_),
    .A1(_00699_),
    .A2(_00825_));
 sg13g2_nor4_1 _06370_ (.A(_00752_),
    .B(_00806_),
    .C(_00824_),
    .D(_00826_),
    .Y(_00827_));
 sg13g2_nor2_2 _06371_ (.A(net57),
    .B(net63),
    .Y(_00828_));
 sg13g2_nor2_1 _06372_ (.A(net76),
    .B(_00653_),
    .Y(_00829_));
 sg13g2_a21oi_1 _06373_ (.A1(_00624_),
    .A2(_00828_),
    .Y(_00830_),
    .B1(_00829_));
 sg13g2_o21ai_1 _06374_ (.B1(_00830_),
    .Y(_00831_),
    .A1(net41),
    .A2(_00784_));
 sg13g2_a21o_1 _06375_ (.A2(_00831_),
    .A1(_00701_),
    .B1(_00756_),
    .X(_00832_));
 sg13g2_a21oi_1 _06376_ (.A1(_00626_),
    .A2(_00768_),
    .Y(_00833_),
    .B1(_00718_));
 sg13g2_nor2_2 _06377_ (.A(net137),
    .B(_00538_),
    .Y(_00834_));
 sg13g2_o21ai_1 _06378_ (.B1(_00720_),
    .Y(_00835_),
    .A1(net131),
    .A2(_00750_));
 sg13g2_nor2_1 _06379_ (.A(_00558_),
    .B(net89),
    .Y(_00836_));
 sg13g2_nand2_1 _06380_ (.Y(_00837_),
    .A(_00558_),
    .B(net79));
 sg13g2_o21ai_1 _06381_ (.B1(_00837_),
    .Y(_00838_),
    .A1(net90),
    .A2(_00836_));
 sg13g2_a221oi_1 _06382_ (.B2(net66),
    .C1(net60),
    .B1(_00838_),
    .A1(_00834_),
    .Y(_00839_),
    .A2(_00835_));
 sg13g2_a21oi_1 _06383_ (.A1(net51),
    .A2(_00833_),
    .Y(_00840_),
    .B1(_00839_));
 sg13g2_nor2b_1 _06384_ (.A(net375),
    .B_N(net384),
    .Y(_00841_));
 sg13g2_o21ai_1 _06385_ (.B1(_00841_),
    .Y(_00842_),
    .A1(_00832_),
    .A2(_00840_));
 sg13g2_o21ai_1 _06386_ (.B1(_05383_),
    .Y(_00843_),
    .A1(_00827_),
    .A2(_00842_));
 sg13g2_or3_1 _06387_ (.A(_00698_),
    .B(_00796_),
    .C(_00843_),
    .X(_00844_));
 sg13g2_nand2_2 _06388_ (.Y(_00845_),
    .A(net106),
    .B(net72));
 sg13g2_o21ai_1 _06389_ (.B1(_00709_),
    .Y(_00846_),
    .A1(_00845_),
    .A2(net136));
 sg13g2_nand2_1 _06390_ (.Y(_00847_),
    .A(net87),
    .B(net61));
 sg13g2_a21oi_1 _06391_ (.A1(_00847_),
    .A2(net172),
    .Y(_00848_),
    .B1(net168));
 sg13g2_a221oi_1 _06392_ (.B2(net168),
    .C1(_00848_),
    .B1(_00846_),
    .A1(_00845_),
    .Y(_00849_),
    .A2(net70));
 sg13g2_nand2_1 _06393_ (.Y(_00850_),
    .A(net137),
    .B(net170));
 sg13g2_a21o_1 _06394_ (.A2(_00850_),
    .A1(_00847_),
    .B1(net172),
    .X(_00851_));
 sg13g2_o21ai_1 _06395_ (.B1(_00711_),
    .Y(_00852_),
    .A1(net93),
    .A2(net133));
 sg13g2_a22oi_1 _06396_ (.Y(_00853_),
    .B1(_00852_),
    .B2(net65),
    .A2(_00600_),
    .A1(_00680_));
 sg13g2_a21oi_1 _06397_ (.A1(_00851_),
    .A2(_00853_),
    .Y(_00854_),
    .B1(net90));
 sg13g2_a21o_1 _06398_ (.A2(_00849_),
    .A1(net88),
    .B1(_00854_),
    .X(_00855_));
 sg13g2_o21ai_1 _06399_ (.B1(_00725_),
    .Y(_00856_),
    .A1(net49),
    .A2(_00855_));
 sg13g2_nand2_1 _06400_ (.Y(_00857_),
    .A(net319),
    .B(_00856_));
 sg13g2_nor3_1 _06401_ (.A(net70),
    .B(_00640_),
    .C(net63),
    .Y(_00858_));
 sg13g2_o21ai_1 _06402_ (.B1(_00626_),
    .Y(_00859_),
    .A1(_00829_),
    .A2(_00858_));
 sg13g2_nand2b_1 _06403_ (.Y(_00860_),
    .B(net58),
    .A_N(_00633_));
 sg13g2_o21ai_1 _06404_ (.B1(net70),
    .Y(_00861_),
    .A1(net62),
    .A2(_00834_));
 sg13g2_a22oi_1 _06405_ (.Y(_00862_),
    .B1(net71),
    .B2(_00845_),
    .A2(net135),
    .A1(net87));
 sg13g2_nor2_1 _06406_ (.A(net106),
    .B(net72),
    .Y(_00863_));
 sg13g2_o21ai_1 _06407_ (.B1(net107),
    .Y(_00864_),
    .A1(_00680_),
    .A2(_00863_));
 sg13g2_nand4_1 _06408_ (.B(_00861_),
    .C(_00862_),
    .A(net131),
    .Y(_00865_),
    .D(_00864_));
 sg13g2_buf_1 _06409_ (.A(net170),
    .X(_00866_));
 sg13g2_a22oi_1 _06410_ (.Y(_00867_),
    .B1(net76),
    .B2(_00680_),
    .A2(net136),
    .A1(_00863_));
 sg13g2_nor2_1 _06411_ (.A(_00570_),
    .B(net136),
    .Y(_00868_));
 sg13g2_nand2_1 _06412_ (.Y(_00869_),
    .A(net72),
    .B(_00570_));
 sg13g2_a221oi_1 _06413_ (.B2(_00807_),
    .C1(net132),
    .B1(_00869_),
    .A1(_00863_),
    .Y(_00870_),
    .A2(_00868_));
 sg13g2_o21ai_1 _06414_ (.B1(_00870_),
    .Y(_00871_),
    .A1(net130),
    .A2(_00867_));
 sg13g2_nand3_1 _06415_ (.B(_00865_),
    .C(_00871_),
    .A(net56),
    .Y(_00872_));
 sg13g2_nand4_1 _06416_ (.B(_00859_),
    .C(_00860_),
    .A(net344),
    .Y(_00873_),
    .D(_00872_));
 sg13g2_and2_1 _06417_ (.A(net343),
    .B(_00873_),
    .X(_00874_));
 sg13g2_nor2_1 _06418_ (.A(net384),
    .B(net60),
    .Y(_00875_));
 sg13g2_o21ai_1 _06419_ (.B1(_00555_),
    .Y(_00876_),
    .A1(net107),
    .A2(_00703_));
 sg13g2_nor2_1 _06420_ (.A(net108),
    .B(_00532_),
    .Y(_00877_));
 sg13g2_nand2_1 _06421_ (.Y(_00878_),
    .A(net202),
    .B(net137));
 sg13g2_nand2_1 _06422_ (.Y(_00879_),
    .A(net87),
    .B(net107));
 sg13g2_o21ai_1 _06423_ (.B1(_00879_),
    .Y(_00880_),
    .A1(_00878_),
    .A2(_00660_));
 sg13g2_a221oi_1 _06424_ (.B2(_00673_),
    .C1(_00730_),
    .B1(_00880_),
    .A1(_00603_),
    .Y(_00881_),
    .A2(_00812_));
 sg13g2_o21ai_1 _06425_ (.B1(_00881_),
    .Y(_00882_),
    .A1(_00869_),
    .A2(_00722_));
 sg13g2_a21o_1 _06426_ (.A2(_00877_),
    .A1(_00876_),
    .B1(_00882_),
    .X(_00883_));
 sg13g2_o21ai_1 _06427_ (.B1(net133),
    .Y(_00884_),
    .A1(net130),
    .A2(net172));
 sg13g2_a221oi_1 _06428_ (.B2(_00884_),
    .C1(_00655_),
    .B1(_00828_),
    .A1(_00866_),
    .Y(_00885_),
    .A2(_00617_));
 sg13g2_a21oi_1 _06429_ (.A1(_00750_),
    .A2(_00720_),
    .Y(_00886_),
    .B1(_00600_));
 sg13g2_nor3_1 _06430_ (.A(net74),
    .B(net107),
    .C(_00886_),
    .Y(_00887_));
 sg13g2_a21oi_1 _06431_ (.A1(_00800_),
    .A2(_00885_),
    .Y(_00888_),
    .B1(_00887_));
 sg13g2_a22oi_1 _06432_ (.Y(_00889_),
    .B1(net76),
    .B2(net54),
    .A2(net136),
    .A1(net80));
 sg13g2_nand2_1 _06433_ (.Y(_00890_),
    .A(net74),
    .B(net70));
 sg13g2_a221oi_1 _06434_ (.B2(net58),
    .C1(net90),
    .B1(_00890_),
    .A1(_00680_),
    .Y(_00891_),
    .A2(net135));
 sg13g2_a21oi_1 _06435_ (.A1(net88),
    .A2(_00889_),
    .Y(_00892_),
    .B1(_00891_));
 sg13g2_nand3_1 _06436_ (.B(_00709_),
    .C(_00813_),
    .A(_00845_),
    .Y(_00893_));
 sg13g2_nand2_1 _06437_ (.Y(_00894_),
    .A(net87),
    .B(net76));
 sg13g2_o21ai_1 _06438_ (.B1(_00894_),
    .Y(_00895_),
    .A1(net87),
    .A2(net133));
 sg13g2_a221oi_1 _06439_ (.B2(net90),
    .C1(net168),
    .B1(_00895_),
    .A1(net135),
    .Y(_00896_),
    .A2(_00863_));
 sg13g2_a21oi_1 _06440_ (.A1(_00893_),
    .A2(_00896_),
    .Y(_00897_),
    .B1(net344));
 sg13g2_o21ai_1 _06441_ (.B1(_00897_),
    .Y(_00898_),
    .A1(_00866_),
    .A2(_00892_));
 sg13g2_o21ai_1 _06442_ (.B1(_00898_),
    .Y(_00899_),
    .A1(_00883_),
    .A2(_00888_));
 sg13g2_a21oi_1 _06443_ (.A1(_00642_),
    .A2(_00829_),
    .Y(_00900_),
    .B1(_00728_));
 sg13g2_o21ai_1 _06444_ (.B1(_00900_),
    .Y(_00901_),
    .A1(_00642_),
    .A2(_00821_));
 sg13g2_nand2_1 _06445_ (.Y(_00902_),
    .A(_00637_),
    .B(_00901_));
 sg13g2_nand3_1 _06446_ (.B(net375),
    .C(_00902_),
    .A(net385),
    .Y(_00903_));
 sg13g2_a221oi_1 _06447_ (.B2(_00899_),
    .C1(_00903_),
    .B1(_00875_),
    .A1(_00857_),
    .Y(_00904_),
    .A2(_00874_));
 sg13g2_o21ai_1 _06448_ (.B1(net205),
    .Y(_00905_),
    .A1(net130),
    .A2(net57));
 sg13g2_buf_1 _06449_ (.A(_00541_),
    .X(_00906_));
 sg13g2_a22oi_1 _06450_ (.Y(_00907_),
    .B1(_00905_),
    .B2(net231),
    .A2(net55),
    .A1(_00710_));
 sg13g2_nor2_1 _06451_ (.A(net170),
    .B(net205),
    .Y(_00908_));
 sg13g2_a22oi_1 _06452_ (.Y(_00909_),
    .B1(net55),
    .B2(_00908_),
    .A2(net136),
    .A1(net74));
 sg13g2_a21oi_1 _06453_ (.A1(_00907_),
    .A2(_00909_),
    .Y(_00910_),
    .B1(net51));
 sg13g2_a21o_1 _06454_ (.A2(net130),
    .A1(net231),
    .B1(_00834_),
    .X(_00911_));
 sg13g2_a22oi_1 _06455_ (.Y(_00912_),
    .B1(net57),
    .B2(_00911_),
    .A2(_00815_),
    .A1(net231));
 sg13g2_buf_1 _06456_ (.A(_00551_),
    .X(_00913_));
 sg13g2_nand2_1 _06457_ (.Y(_00914_),
    .A(net201),
    .B(net170));
 sg13g2_nand2_1 _06458_ (.Y(_00915_),
    .A(net168),
    .B(net135));
 sg13g2_nand3_1 _06459_ (.B(net53),
    .C(_00908_),
    .A(net74),
    .Y(_00916_));
 sg13g2_nand4_1 _06460_ (.B(net53),
    .C(net231),
    .A(net74),
    .Y(_00917_),
    .D(net168));
 sg13g2_nand4_1 _06461_ (.B(_00915_),
    .C(_00916_),
    .A(_00914_),
    .Y(_00918_),
    .D(_00917_));
 sg13g2_nand2_1 _06462_ (.Y(_00919_),
    .A(net88),
    .B(_00918_));
 sg13g2_nand3_1 _06463_ (.B(_00912_),
    .C(_00919_),
    .A(_00910_),
    .Y(_00920_));
 sg13g2_a22oi_1 _06464_ (.Y(_00921_),
    .B1(_00729_),
    .B2(_00757_),
    .A2(net68),
    .A1(_00532_));
 sg13g2_xnor2_1 _06465_ (.Y(_00922_),
    .A(net132),
    .B(net69));
 sg13g2_a22oi_1 _06466_ (.Y(_00923_),
    .B1(_00922_),
    .B2(net66),
    .A2(_00782_),
    .A1(_00671_));
 sg13g2_o21ai_1 _06467_ (.B1(_00771_),
    .Y(_00924_),
    .A1(net75),
    .A2(_00923_));
 sg13g2_o21ai_1 _06468_ (.B1(net50),
    .Y(_00925_),
    .A1(_00921_),
    .A2(_00924_));
 sg13g2_a22oi_1 _06469_ (.Y(_00926_),
    .B1(_00925_),
    .B2(net320),
    .A2(_00920_),
    .A1(_00643_));
 sg13g2_and2_1 _06470_ (.A(_05376_),
    .B(_05322_),
    .X(_00927_));
 sg13g2_buf_1 _06471_ (.A(_00927_),
    .X(_00928_));
 sg13g2_nand3_1 _06472_ (.B(_00758_),
    .C(_00928_),
    .A(_00637_),
    .Y(_00929_));
 sg13g2_nand2_1 _06473_ (.Y(_00930_),
    .A(net78),
    .B(net77));
 sg13g2_nor4_1 _06474_ (.A(_00730_),
    .B(net108),
    .C(_00930_),
    .D(_00657_),
    .Y(_00931_));
 sg13g2_o21ai_1 _06475_ (.B1(net387),
    .Y(_00932_),
    .A1(net76),
    .A2(_00575_));
 sg13g2_nand3_1 _06476_ (.B(_00750_),
    .C(_00932_),
    .A(net108),
    .Y(_00933_));
 sg13g2_a21oi_1 _06477_ (.A1(net387),
    .A2(net59),
    .Y(_00934_),
    .B1(net70));
 sg13g2_nand2_1 _06478_ (.Y(_00935_),
    .A(net90),
    .B(_00934_));
 sg13g2_nor2_1 _06479_ (.A(net344),
    .B(net79),
    .Y(_00936_));
 sg13g2_nand2_1 _06480_ (.Y(_00937_),
    .A(net65),
    .B(net78));
 sg13g2_a221oi_1 _06481_ (.B2(_00937_),
    .C1(_00734_),
    .B1(_00936_),
    .A1(_00933_),
    .Y(_00938_),
    .A2(_00935_));
 sg13g2_o21ai_1 _06482_ (.B1(_00875_),
    .Y(_00939_),
    .A1(_00931_),
    .A2(_00938_));
 sg13g2_nand4_1 _06483_ (.B(_05360_),
    .C(_00929_),
    .A(net385),
    .Y(_00940_),
    .D(_00939_));
 sg13g2_a21oi_1 _06484_ (.A1(net343),
    .A2(_00926_),
    .Y(_00941_),
    .B1(_00940_));
 sg13g2_o21ai_1 _06485_ (.B1(_00524_),
    .Y(_00942_),
    .A1(_05184_),
    .A2(_05189_));
 sg13g2_nand4_1 _06486_ (.B(net378),
    .C(_05174_),
    .A(net395),
    .Y(_00943_),
    .D(_00520_));
 sg13g2_inv_1 _06487_ (.Y(_00944_),
    .A(net378));
 sg13g2_o21ai_1 _06488_ (.B1(_00944_),
    .Y(_00945_),
    .A1(net382),
    .A2(_00524_));
 sg13g2_nand3_1 _06489_ (.B(_00943_),
    .C(_00945_),
    .A(_00942_),
    .Y(_00946_));
 sg13g2_buf_1 _06490_ (.A(_00946_),
    .X(_00947_));
 sg13g2_xor2_1 _06491_ (.B(_00947_),
    .A(_00879_),
    .X(_00948_));
 sg13g2_nor4_1 _06492_ (.A(net389),
    .B(_00904_),
    .C(_00941_),
    .D(_00948_),
    .Y(_00949_));
 sg13g2_inv_1 _06493_ (.Y(_00950_),
    .A(net389));
 sg13g2_xnor2_1 _06494_ (.Y(_00951_),
    .A(_00737_),
    .B(_00635_));
 sg13g2_nand2_1 _06495_ (.Y(_00952_),
    .A(_00575_),
    .B(net71));
 sg13g2_nand2_1 _06496_ (.Y(_00953_),
    .A(net77),
    .B(_00721_));
 sg13g2_nand2_1 _06497_ (.Y(_00954_),
    .A(_00578_),
    .B(net71));
 sg13g2_o21ai_1 _06498_ (.B1(_00954_),
    .Y(_00955_),
    .A1(_00606_),
    .A2(_00953_));
 sg13g2_a22oi_1 _06499_ (.Y(_00956_),
    .B1(_00955_),
    .B2(net80),
    .A2(_00828_),
    .A1(_00603_));
 sg13g2_o21ai_1 _06500_ (.B1(_00956_),
    .Y(_00957_),
    .A1(_00951_),
    .A2(_00952_));
 sg13g2_o21ai_1 _06501_ (.B1(_00906_),
    .Y(_00958_),
    .A1(net171),
    .A2(_00834_));
 sg13g2_o21ai_1 _06502_ (.B1(_00958_),
    .Y(_00959_),
    .A1(net110),
    .A2(_00914_));
 sg13g2_a21oi_1 _06503_ (.A1(net169),
    .A2(_00850_),
    .Y(_00960_),
    .B1(net172));
 sg13g2_a221oi_1 _06504_ (.B2(_00959_),
    .C1(_00960_),
    .B1(_00545_),
    .A1(net134),
    .Y(_00961_),
    .A2(net93));
 sg13g2_nand2_1 _06505_ (.Y(_00962_),
    .A(_00578_),
    .B(net91));
 sg13g2_nand2_1 _06506_ (.Y(_00963_),
    .A(_00611_),
    .B(net89));
 sg13g2_nand3_1 _06507_ (.B(_00962_),
    .C(_00963_),
    .A(net53),
    .Y(_00964_));
 sg13g2_o21ai_1 _06508_ (.B1(_00964_),
    .Y(_00965_),
    .A1(net53),
    .A2(_00961_));
 sg13g2_a21oi_1 _06509_ (.A1(net132),
    .A2(_00598_),
    .Y(_00966_),
    .B1(net170));
 sg13g2_nor2_1 _06510_ (.A(net70),
    .B(_00966_),
    .Y(_00967_));
 sg13g2_o21ai_1 _06511_ (.B1(net56),
    .Y(_00968_),
    .A1(_00965_),
    .A2(_00967_));
 sg13g2_o21ai_1 _06512_ (.B1(_00968_),
    .Y(_00969_),
    .A1(net50),
    .A2(_00957_));
 sg13g2_a21oi_1 _06513_ (.A1(_00812_),
    .A2(_00836_),
    .Y(_00970_),
    .B1(_00817_));
 sg13g2_nand4_1 _06514_ (.B(_00690_),
    .C(_00634_),
    .A(net132),
    .Y(_00971_),
    .D(_00703_));
 sg13g2_a21o_1 _06515_ (.A2(_00937_),
    .A1(_00686_),
    .B1(_00971_),
    .X(_00972_));
 sg13g2_a21oi_1 _06516_ (.A1(_00970_),
    .A2(_00972_),
    .Y(_00973_),
    .B1(_00635_));
 sg13g2_nor2_1 _06517_ (.A(net87),
    .B(net61),
    .Y(_00974_));
 sg13g2_a21oi_1 _06518_ (.A1(net67),
    .A2(_00561_),
    .Y(_00975_),
    .B1(_00547_));
 sg13g2_nor4_1 _06519_ (.A(net109),
    .B(_00674_),
    .C(_00974_),
    .D(_00975_),
    .Y(_00976_));
 sg13g2_a21oi_1 _06520_ (.A1(_00668_),
    .A2(_00745_),
    .Y(_00977_),
    .B1(_00976_));
 sg13g2_and2_1 _06521_ (.A(_00477_),
    .B(_00486_),
    .X(_00978_));
 sg13g2_nand3_1 _06522_ (.B(_00534_),
    .C(net133),
    .A(_00530_),
    .Y(_00979_));
 sg13g2_o21ai_1 _06523_ (.B1(_00979_),
    .Y(_00980_),
    .A1(net93),
    .A2(_00534_));
 sg13g2_nor3_1 _06524_ (.A(net106),
    .B(_00534_),
    .C(net135),
    .Y(_00981_));
 sg13g2_a21o_1 _06525_ (.A2(_00534_),
    .A1(_00799_),
    .B1(_00981_),
    .X(_00982_));
 sg13g2_nor3_1 _06526_ (.A(_00455_),
    .B(net106),
    .C(net135),
    .Y(_00983_));
 sg13g2_and2_1 _06527_ (.A(_00455_),
    .B(net106),
    .X(_00984_));
 sg13g2_o21ai_1 _06528_ (.B1(_00409_),
    .Y(_00985_),
    .A1(_00983_),
    .A2(_00984_));
 sg13g2_nand3_1 _06529_ (.B(_00600_),
    .C(_00985_),
    .A(_00612_),
    .Y(_00986_));
 sg13g2_a221oi_1 _06530_ (.B2(_00494_),
    .C1(_00986_),
    .B1(_00982_),
    .A1(_00978_),
    .Y(_00987_),
    .A2(_00980_));
 sg13g2_xnor2_1 _06531_ (.Y(_00988_),
    .A(net202),
    .B(net205));
 sg13g2_nand2_1 _06532_ (.Y(_00989_),
    .A(net203),
    .B(net205));
 sg13g2_nor2_1 _06533_ (.A(net201),
    .B(_00989_),
    .Y(_00990_));
 sg13g2_a21oi_1 _06534_ (.A1(net201),
    .A2(_00988_),
    .Y(_00991_),
    .B1(_00990_));
 sg13g2_nor3_1 _06535_ (.A(_00845_),
    .B(net130),
    .C(_00991_),
    .Y(_00992_));
 sg13g2_nor2_1 _06536_ (.A(_00987_),
    .B(_00992_),
    .Y(_00993_));
 sg13g2_nand3_1 _06537_ (.B(_00977_),
    .C(_00993_),
    .A(net56),
    .Y(_00994_));
 sg13g2_o21ai_1 _06538_ (.B1(_00994_),
    .Y(_00995_),
    .A1(net50),
    .A2(_00973_));
 sg13g2_nand3_1 _06539_ (.B(net64),
    .C(_00703_),
    .A(_00690_),
    .Y(_00996_));
 sg13g2_o21ai_1 _06540_ (.B1(_00970_),
    .Y(_00997_),
    .A1(_00613_),
    .A2(_00996_));
 sg13g2_a21oi_1 _06541_ (.A1(_00635_),
    .A2(_00997_),
    .Y(_00998_),
    .B1(net343));
 sg13g2_nand2_1 _06542_ (.Y(_00999_),
    .A(net375),
    .B(net319));
 sg13g2_a221oi_1 _06543_ (.B2(_00998_),
    .C1(_00999_),
    .B1(_00995_),
    .A1(net343),
    .Y(_01000_),
    .A2(_00969_));
 sg13g2_nand2_1 _06544_ (.Y(_01001_),
    .A(_00745_),
    .B(_00828_));
 sg13g2_nand2_1 _06545_ (.Y(_01002_),
    .A(net50),
    .B(_01001_));
 sg13g2_nand4_1 _06546_ (.B(net64),
    .C(net55),
    .A(net49),
    .Y(_01003_),
    .D(_00722_));
 sg13g2_nand3_1 _06547_ (.B(_00773_),
    .C(_01003_),
    .A(net52),
    .Y(_01004_));
 sg13g2_nand2_1 _06548_ (.Y(_01005_),
    .A(_00425_),
    .B(net204));
 sg13g2_or2_1 _06549_ (.X(_01006_),
    .B(_01005_),
    .A(_00657_));
 sg13g2_a21oi_1 _06550_ (.A1(_00670_),
    .A2(_00782_),
    .Y(_01007_),
    .B1(_00596_));
 sg13g2_nand3_1 _06551_ (.B(net65),
    .C(_00734_),
    .A(net109),
    .Y(_01008_));
 sg13g2_a21oi_1 _06552_ (.A1(net132),
    .A2(net64),
    .Y(_01009_),
    .B1(net76));
 sg13g2_a22oi_1 _06553_ (.Y(_01010_),
    .B1(_01008_),
    .B2(_01009_),
    .A2(_01007_),
    .A1(_01006_));
 sg13g2_or2_1 _06554_ (.X(_01011_),
    .B(_01010_),
    .A(_00689_));
 sg13g2_nand3_1 _06555_ (.B(_01004_),
    .C(_01011_),
    .A(_01002_),
    .Y(_01012_));
 sg13g2_nor2_1 _06556_ (.A(_00557_),
    .B(_00717_),
    .Y(_01013_));
 sg13g2_nand2_1 _06557_ (.Y(_01014_),
    .A(net67),
    .B(_01013_));
 sg13g2_o21ai_1 _06558_ (.B1(_01014_),
    .Y(_01015_),
    .A1(net62),
    .A2(_00953_));
 sg13g2_nor3_1 _06559_ (.A(_00579_),
    .B(_00606_),
    .C(_00555_),
    .Y(_01016_));
 sg13g2_nor3_1 _06560_ (.A(net62),
    .B(_00555_),
    .C(_00989_),
    .Y(_01017_));
 sg13g2_nor3_1 _06561_ (.A(_01015_),
    .B(_01016_),
    .C(_01017_),
    .Y(_01018_));
 sg13g2_nor4_1 _06562_ (.A(net134),
    .B(net65),
    .C(net168),
    .D(_00545_),
    .Y(_01019_));
 sg13g2_nand3_1 _06563_ (.B(net201),
    .C(_00545_),
    .A(net171),
    .Y(_01020_));
 sg13g2_nor3_1 _06564_ (.A(net62),
    .B(net130),
    .C(_01020_),
    .Y(_01021_));
 sg13g2_a21oi_1 _06565_ (.A1(_00913_),
    .A2(_01019_),
    .Y(_01022_),
    .B1(_01021_));
 sg13g2_nand2_1 _06566_ (.Y(_01023_),
    .A(net79),
    .B(_00624_));
 sg13g2_a21oi_1 _06567_ (.A1(_01018_),
    .A2(_01022_),
    .Y(_01024_),
    .B1(_01023_));
 sg13g2_nor3_1 _06568_ (.A(_05383_),
    .B(net319),
    .C(_01024_),
    .Y(_01025_));
 sg13g2_o21ai_1 _06569_ (.B1(net58),
    .Y(_01026_),
    .A1(_00782_),
    .A2(_01013_));
 sg13g2_a21oi_1 _06570_ (.A1(_00770_),
    .A2(_01026_),
    .Y(_01027_),
    .B1(_01023_));
 sg13g2_o21ai_1 _06571_ (.B1(net52),
    .Y(_01028_),
    .A1(_00747_),
    .A2(_01027_));
 sg13g2_nand2_1 _06572_ (.Y(_01029_),
    .A(_00730_),
    .B(net60));
 sg13g2_nand2_1 _06573_ (.Y(_01030_),
    .A(net62),
    .B(_00906_));
 sg13g2_nand4_1 _06574_ (.B(_00709_),
    .C(_00908_),
    .A(net131),
    .Y(_01031_),
    .D(_01030_));
 sg13g2_nor4_1 _06575_ (.A(_00530_),
    .B(net201),
    .C(net170),
    .D(_00545_),
    .Y(_01032_));
 sg13g2_and3_1 _06576_ (.X(_01033_),
    .A(net169),
    .B(_00534_),
    .C(_00710_));
 sg13g2_xnor2_1 _06577_ (.Y(_01034_),
    .A(net94),
    .B(_00799_));
 sg13g2_a221oi_1 _06578_ (.B2(_01034_),
    .C1(net387),
    .B1(_01033_),
    .A1(net131),
    .Y(_01035_),
    .A2(_01032_));
 sg13g2_nor2_1 _06579_ (.A(net168),
    .B(net133),
    .Y(_01036_));
 sg13g2_nand2b_1 _06580_ (.Y(_01037_),
    .B(_01036_),
    .A_N(_00707_));
 sg13g2_nor2_1 _06581_ (.A(_00529_),
    .B(net205),
    .Y(_01038_));
 sg13g2_nand3_1 _06582_ (.B(net205),
    .C(_00815_),
    .A(_00470_),
    .Y(_01039_));
 sg13g2_o21ai_1 _06583_ (.B1(_01039_),
    .Y(_01040_),
    .A1(_01005_),
    .A2(_01038_));
 sg13g2_o21ai_1 _06584_ (.B1(_00569_),
    .Y(_01041_),
    .A1(net204),
    .A2(_00559_));
 sg13g2_nor3_1 _06585_ (.A(net203),
    .B(net94),
    .C(_01041_),
    .Y(_01042_));
 sg13g2_a21o_1 _06586_ (.A2(_01040_),
    .A1(net94),
    .B1(_01042_),
    .X(_01043_));
 sg13g2_nand2_1 _06587_ (.Y(_01044_),
    .A(net202),
    .B(net231));
 sg13g2_mux2_1 _06588_ (.A0(_01044_),
    .A1(_00989_),
    .S(net94),
    .X(_01045_));
 sg13g2_nor3_1 _06589_ (.A(net106),
    .B(net170),
    .C(_01045_),
    .Y(_01046_));
 sg13g2_a21oi_1 _06590_ (.A1(net201),
    .A2(_01043_),
    .Y(_01047_),
    .B1(_01046_));
 sg13g2_xnor2_1 _06591_ (.Y(_01048_),
    .A(_00529_),
    .B(_00551_));
 sg13g2_nor4_1 _06592_ (.A(_00409_),
    .B(net171),
    .C(_00978_),
    .D(_01048_),
    .Y(_01049_));
 sg13g2_nor2_1 _06593_ (.A(net231),
    .B(_01038_),
    .Y(_01050_));
 sg13g2_a21oi_1 _06594_ (.A1(net137),
    .A2(_00559_),
    .Y(_01051_),
    .B1(_01050_));
 sg13g2_nor3_1 _06595_ (.A(net202),
    .B(net94),
    .C(_01051_),
    .Y(_01052_));
 sg13g2_o21ai_1 _06596_ (.B1(net204),
    .Y(_01053_),
    .A1(_01049_),
    .A2(_01052_));
 sg13g2_mux2_1 _06597_ (.A0(_01047_),
    .A1(_01053_),
    .S(_00534_),
    .X(_01054_));
 sg13g2_nand4_1 _06598_ (.B(_01035_),
    .C(_01037_),
    .A(_01031_),
    .Y(_01055_),
    .D(_01054_));
 sg13g2_a21oi_1 _06599_ (.A1(_00750_),
    .A2(_00720_),
    .Y(_01056_),
    .B1(_00625_));
 sg13g2_nor2_1 _06600_ (.A(_00747_),
    .B(_01056_),
    .Y(_01057_));
 sg13g2_o21ai_1 _06601_ (.B1(net385),
    .Y(_01058_),
    .A1(_00689_),
    .A2(_01057_));
 sg13g2_a221oi_1 _06602_ (.B2(_01055_),
    .C1(_01058_),
    .B1(_01029_),
    .A1(_00637_),
    .Y(_01059_),
    .A2(_00829_));
 sg13g2_nor2_1 _06603_ (.A(_05383_),
    .B(_00645_),
    .Y(_01060_));
 sg13g2_a221oi_1 _06604_ (.B2(_01059_),
    .C1(_01060_),
    .B1(_01028_),
    .A1(_01012_),
    .Y(_01061_),
    .A2(_01025_));
 sg13g2_o21ai_1 _06605_ (.B1(net69),
    .Y(_01062_),
    .A1(_00801_),
    .A2(_00753_));
 sg13g2_a21oi_1 _06606_ (.A1(_01014_),
    .A2(_01062_),
    .Y(_01063_),
    .B1(net79));
 sg13g2_nor3_1 _06607_ (.A(_00629_),
    .B(net41),
    .C(_00954_),
    .Y(_01064_));
 sg13g2_o21ai_1 _06608_ (.B1(net51),
    .Y(_01065_),
    .A1(_01063_),
    .A2(_01064_));
 sg13g2_nand3_1 _06609_ (.B(_00624_),
    .C(_00687_),
    .A(net79),
    .Y(_01066_));
 sg13g2_nor4_1 _06610_ (.A(net56),
    .B(_00654_),
    .C(_00783_),
    .D(_01066_),
    .Y(_01067_));
 sg13g2_nand2_1 _06611_ (.Y(_01068_),
    .A(net79),
    .B(_00739_));
 sg13g2_a21oi_1 _06612_ (.A1(_00962_),
    .A2(_01068_),
    .Y(_01069_),
    .B1(_00581_));
 sg13g2_nor2_1 _06613_ (.A(net69),
    .B(_00598_),
    .Y(_01070_));
 sg13g2_nor2_1 _06614_ (.A(_00717_),
    .B(_01070_),
    .Y(_01071_));
 sg13g2_nor4_1 _06615_ (.A(net60),
    .B(_00798_),
    .C(_01069_),
    .D(_01071_),
    .Y(_01072_));
 sg13g2_nor4_1 _06616_ (.A(_00730_),
    .B(_00627_),
    .C(_01067_),
    .D(_01072_),
    .Y(_01073_));
 sg13g2_nor3_1 _06617_ (.A(net387),
    .B(net56),
    .C(_00718_),
    .Y(_01074_));
 sg13g2_nand3_1 _06618_ (.B(net69),
    .C(_00664_),
    .A(net54),
    .Y(_01075_));
 sg13g2_o21ai_1 _06619_ (.B1(_01075_),
    .Y(_01076_),
    .A1(_00659_),
    .A2(net49));
 sg13g2_nand2_1 _06620_ (.Y(_01077_),
    .A(_00653_),
    .B(_00729_));
 sg13g2_o21ai_1 _06621_ (.B1(net52),
    .Y(_01078_),
    .A1(_00609_),
    .A2(net49));
 sg13g2_a221oi_1 _06622_ (.B2(net69),
    .C1(_01078_),
    .B1(_01077_),
    .A1(_00597_),
    .Y(_01079_),
    .A2(_01076_));
 sg13g2_nand4_1 _06623_ (.B(_00680_),
    .C(net168),
    .A(net109),
    .Y(_01080_),
    .D(net205));
 sg13g2_o21ai_1 _06624_ (.B1(_00850_),
    .Y(_01081_),
    .A1(net134),
    .A2(_00834_));
 sg13g2_nand2_1 _06625_ (.Y(_01082_),
    .A(_00545_),
    .B(_01081_));
 sg13g2_a21oi_1 _06626_ (.A1(_01080_),
    .A2(_01082_),
    .Y(_01083_),
    .B1(_00913_));
 sg13g2_o21ai_1 _06627_ (.B1(_00878_),
    .Y(_01084_),
    .A1(net110),
    .A2(_01020_));
 sg13g2_nand2_1 _06628_ (.Y(_01085_),
    .A(net171),
    .B(net106));
 sg13g2_and4_1 _06629_ (.A(net61),
    .B(net133),
    .C(_00878_),
    .D(_01085_),
    .X(_01086_));
 sg13g2_a221oi_1 _06630_ (.B2(net62),
    .C1(_01086_),
    .B1(_01084_),
    .A1(net93),
    .Y(_01087_),
    .A2(net136));
 sg13g2_a21oi_1 _06631_ (.A1(net74),
    .A2(_00813_),
    .Y(_01088_),
    .B1(_05354_));
 sg13g2_o21ai_1 _06632_ (.B1(_01088_),
    .Y(_01089_),
    .A1(net130),
    .A2(_01087_));
 sg13g2_or3_1 _06633_ (.A(net60),
    .B(_01083_),
    .C(_01089_),
    .X(_01090_));
 sg13g2_o21ai_1 _06634_ (.B1(net79),
    .Y(_01091_),
    .A1(_00687_),
    .A2(_00788_));
 sg13g2_nand2_1 _06635_ (.Y(_01092_),
    .A(_01074_),
    .B(_01091_));
 sg13g2_nand3_1 _06636_ (.B(_01090_),
    .C(_01092_),
    .A(_00841_),
    .Y(_01093_));
 sg13g2_a221oi_1 _06637_ (.B2(_01079_),
    .C1(_01093_),
    .B1(_01074_),
    .A1(_01065_),
    .Y(_01094_),
    .A2(_01073_));
 sg13g2_a21oi_1 _06638_ (.A1(_00531_),
    .A2(net68),
    .Y(_01095_),
    .B1(net64));
 sg13g2_nor3_1 _06639_ (.A(net202),
    .B(net77),
    .C(net89),
    .Y(_01096_));
 sg13g2_nor3_1 _06640_ (.A(_00577_),
    .B(_00557_),
    .C(net91),
    .Y(_01097_));
 sg13g2_o21ai_1 _06641_ (.B1(net78),
    .Y(_01098_),
    .A1(_01096_),
    .A2(_01097_));
 sg13g2_nand2_1 _06642_ (.Y(_01099_),
    .A(net384),
    .B(_01098_));
 sg13g2_a221oi_1 _06643_ (.B2(_00820_),
    .C1(_01099_),
    .B1(_01095_),
    .A1(_00666_),
    .Y(_01100_),
    .A2(_01077_));
 sg13g2_nand3_1 _06644_ (.B(_01001_),
    .C(_01100_),
    .A(_00652_),
    .Y(_01101_));
 sg13g2_nand3_1 _06645_ (.B(net320),
    .C(_01101_),
    .A(net375),
    .Y(_01102_));
 sg13g2_o21ai_1 _06646_ (.B1(_00737_),
    .Y(_01103_),
    .A1(_00581_),
    .A2(_00716_));
 sg13g2_and4_1 _06647_ (.A(net66),
    .B(_00762_),
    .C(_01008_),
    .D(_01103_),
    .X(_01104_));
 sg13g2_nand3_1 _06648_ (.B(_00716_),
    .C(_00812_),
    .A(net54),
    .Y(_01105_));
 sg13g2_o21ai_1 _06649_ (.B1(net52),
    .Y(_01106_),
    .A1(net41),
    .A2(_01105_));
 sg13g2_nor2_1 _06650_ (.A(_00625_),
    .B(_00757_),
    .Y(_01107_));
 sg13g2_and2_1 _06651_ (.A(net41),
    .B(_01107_),
    .X(_01108_));
 sg13g2_nor4_1 _06652_ (.A(net343),
    .B(_01104_),
    .C(_01106_),
    .D(_01108_),
    .Y(_01109_));
 sg13g2_a21oi_1 _06653_ (.A1(net59),
    .A2(_00807_),
    .Y(_01110_),
    .B1(_00575_));
 sg13g2_a22oi_1 _06654_ (.Y(_01111_),
    .B1(_01110_),
    .B2(_00613_),
    .A2(_00728_),
    .A1(_00658_));
 sg13g2_nand3_1 _06655_ (.B(_00665_),
    .C(_00812_),
    .A(_00762_),
    .Y(_01112_));
 sg13g2_o21ai_1 _06656_ (.B1(_01112_),
    .Y(_01113_),
    .A1(_00665_),
    .A2(_01111_));
 sg13g2_nand2_1 _06657_ (.Y(_01114_),
    .A(_00607_),
    .B(_00564_));
 sg13g2_nor4_1 _06658_ (.A(_00584_),
    .B(_00930_),
    .C(net57),
    .D(net63),
    .Y(_01115_));
 sg13g2_nor4_1 _06659_ (.A(_05421_),
    .B(net52),
    .C(_01107_),
    .D(_01115_),
    .Y(_01116_));
 sg13g2_o21ai_1 _06660_ (.B1(_01116_),
    .Y(_01117_),
    .A1(_01114_),
    .A2(_01023_));
 sg13g2_a21oi_1 _06661_ (.A1(net69),
    .A2(_01113_),
    .Y(_01118_),
    .B1(_01117_));
 sg13g2_nor3_1 _06662_ (.A(_00409_),
    .B(_00429_),
    .C(_00455_),
    .Y(_01119_));
 sg13g2_o21ai_1 _06663_ (.B1(_00455_),
    .Y(_01120_),
    .A1(_00409_),
    .A2(_00429_));
 sg13g2_o21ai_1 _06664_ (.B1(_01120_),
    .Y(_01121_),
    .A1(net94),
    .A2(_01119_));
 sg13g2_xnor2_1 _06665_ (.Y(_01122_),
    .A(_05250_),
    .B(net171));
 sg13g2_nor4_1 _06666_ (.A(net376),
    .B(net288),
    .C(_00405_),
    .D(_01122_),
    .Y(_01123_));
 sg13g2_nor3_1 _06667_ (.A(net376),
    .B(_00489_),
    .C(_00425_),
    .Y(_01124_));
 sg13g2_a21oi_1 _06668_ (.A1(net376),
    .A2(net203),
    .Y(_01125_),
    .B1(_01124_));
 sg13g2_nand2_2 _06669_ (.Y(_01126_),
    .A(_05219_),
    .B(net420));
 sg13g2_nand3_1 _06670_ (.B(net203),
    .C(_00630_),
    .A(_01126_),
    .Y(_01127_));
 sg13g2_o21ai_1 _06671_ (.B1(_01127_),
    .Y(_01128_),
    .A1(_05249_),
    .A2(_01125_));
 sg13g2_a21oi_1 _06672_ (.A1(_05148_),
    .A2(_01128_),
    .Y(_01129_),
    .B1(_00625_));
 sg13g2_nand3_1 _06673_ (.B(_00563_),
    .C(_01129_),
    .A(net67),
    .Y(_01130_));
 sg13g2_a21oi_1 _06674_ (.A1(_01121_),
    .A2(_01123_),
    .Y(_01131_),
    .B1(_01130_));
 sg13g2_a21oi_1 _06675_ (.A1(_00497_),
    .A2(_01131_),
    .Y(_01132_),
    .B1(net288));
 sg13g2_a22oi_1 _06676_ (.Y(_01133_),
    .B1(_00745_),
    .B2(_00753_),
    .A2(net57),
    .A1(_00603_));
 sg13g2_nand3_1 _06677_ (.B(_01132_),
    .C(_01133_),
    .A(net384),
    .Y(_01134_));
 sg13g2_a21oi_1 _06678_ (.A1(_00659_),
    .A2(_01131_),
    .Y(_01135_),
    .B1(_00492_));
 sg13g2_a221oi_1 _06679_ (.B2(net108),
    .C1(_00403_),
    .B1(_01131_),
    .A1(_05249_),
    .Y(_01136_),
    .A2(_00497_));
 sg13g2_a21oi_1 _06680_ (.A1(_00403_),
    .A2(_01135_),
    .Y(_01137_),
    .B1(_01136_));
 sg13g2_nor2_1 _06681_ (.A(_01134_),
    .B(_01137_),
    .Y(_01138_));
 sg13g2_nor4_1 _06682_ (.A(_01102_),
    .B(_01109_),
    .C(_01118_),
    .D(_01138_),
    .Y(_01139_));
 sg13g2_nor4_1 _06683_ (.A(_01000_),
    .B(_01061_),
    .C(_01094_),
    .D(_01139_),
    .Y(_01140_));
 sg13g2_nor4_1 _06684_ (.A(net60),
    .B(_00574_),
    .C(_00609_),
    .D(_00784_),
    .Y(_01141_));
 sg13g2_nor4_1 _06685_ (.A(_00650_),
    .B(_00584_),
    .C(_00609_),
    .D(_00654_),
    .Y(_01142_));
 sg13g2_nor4_1 _06686_ (.A(_00580_),
    .B(_00499_),
    .C(net68),
    .D(_00658_),
    .Y(_01143_));
 sg13g2_nor3_1 _06687_ (.A(_01141_),
    .B(_01142_),
    .C(_01143_),
    .Y(_01144_));
 sg13g2_o21ai_1 _06688_ (.B1(_00657_),
    .Y(_01145_),
    .A1(_00580_),
    .A2(_00656_));
 sg13g2_nand4_1 _06689_ (.B(net66),
    .C(net68),
    .A(_00651_),
    .Y(_01146_),
    .D(_01145_));
 sg13g2_nand3_1 _06690_ (.B(_00607_),
    .C(_00718_),
    .A(_00499_),
    .Y(_01147_));
 sg13g2_nand4_1 _06691_ (.B(net54),
    .C(net75),
    .A(_00651_),
    .Y(_01148_),
    .D(_00812_));
 sg13g2_nand4_1 _06692_ (.B(_01146_),
    .C(_01147_),
    .A(_01144_),
    .Y(_01149_),
    .D(_01148_));
 sg13g2_a221oi_1 _06693_ (.B2(_00914_),
    .C1(net93),
    .B1(net63),
    .A1(net59),
    .Y(_01150_),
    .A2(_00655_));
 sg13g2_nand2_1 _06694_ (.Y(_01151_),
    .A(net132),
    .B(net107));
 sg13g2_o21ai_1 _06695_ (.B1(_00915_),
    .Y(_01152_),
    .A1(net59),
    .A2(_01151_));
 sg13g2_nor3_1 _06696_ (.A(net74),
    .B(_00660_),
    .C(_00828_),
    .Y(_01153_));
 sg13g2_a221oi_1 _06697_ (.B2(net80),
    .C1(_01153_),
    .B1(_01152_),
    .A1(_00708_),
    .Y(_01154_),
    .A2(_01150_));
 sg13g2_o21ai_1 _06698_ (.B1(_00748_),
    .Y(_01155_),
    .A1(_00500_),
    .A2(_01154_));
 sg13g2_mux2_1 _06699_ (.A0(_01149_),
    .A1(_01155_),
    .S(net319),
    .X(_01156_));
 sg13g2_o21ai_1 _06700_ (.B1(_00609_),
    .Y(_01157_),
    .A1(net54),
    .A2(_00930_));
 sg13g2_o21ai_1 _06701_ (.B1(net75),
    .Y(_01158_),
    .A1(_00591_),
    .A2(_01013_));
 sg13g2_o21ai_1 _06702_ (.B1(_01158_),
    .Y(_01159_),
    .A1(net75),
    .A2(_00953_));
 sg13g2_a22oi_1 _06703_ (.Y(_01160_),
    .B1(_01159_),
    .B2(_00671_),
    .A2(_01157_),
    .A1(_00742_));
 sg13g2_nand3b_1 _06704_ (.B(net320),
    .C(_00652_),
    .Y(_01161_),
    .A_N(_01160_));
 sg13g2_nand4_1 _06705_ (.B(net51),
    .C(net54),
    .A(net319),
    .Y(_01162_),
    .D(_00718_));
 sg13g2_o21ai_1 _06706_ (.B1(net108),
    .Y(_01163_),
    .A1(_00709_),
    .A2(net107));
 sg13g2_nand3_1 _06707_ (.B(net80),
    .C(_00555_),
    .A(net88),
    .Y(_01164_));
 sg13g2_nand3_1 _06708_ (.B(_01163_),
    .C(_01164_),
    .A(net66),
    .Y(_01165_));
 sg13g2_nor2_1 _06709_ (.A(net108),
    .B(_00548_),
    .Y(_01166_));
 sg13g2_nand3_1 _06710_ (.B(net80),
    .C(net59),
    .A(net109),
    .Y(_01167_));
 sg13g2_o21ai_1 _06711_ (.B1(_01167_),
    .Y(_01168_),
    .A1(net54),
    .A2(_00879_));
 sg13g2_nor4_1 _06712_ (.A(net344),
    .B(_00967_),
    .C(_01166_),
    .D(_01168_),
    .Y(_01169_));
 sg13g2_nand3_1 _06713_ (.B(_01165_),
    .C(_01169_),
    .A(net50),
    .Y(_01170_));
 sg13g2_nand3_1 _06714_ (.B(_01162_),
    .C(_01170_),
    .A(_01161_),
    .Y(_01171_));
 sg13g2_a21oi_1 _06715_ (.A1(net53),
    .A2(_00555_),
    .Y(_01172_),
    .B1(net107));
 sg13g2_o21ai_1 _06716_ (.B1(_00561_),
    .Y(_01173_),
    .A1(net87),
    .A2(_00585_));
 sg13g2_a21oi_1 _06717_ (.A1(net172),
    .A2(_01173_),
    .Y(_01174_),
    .B1(net90));
 sg13g2_o21ai_1 _06718_ (.B1(_01174_),
    .Y(_01175_),
    .A1(net80),
    .A2(_01172_));
 sg13g2_nand2_1 _06719_ (.Y(_01176_),
    .A(_00974_),
    .B(_00564_));
 sg13g2_nand3_1 _06720_ (.B(_01175_),
    .C(_01176_),
    .A(net320),
    .Y(_01177_));
 sg13g2_o21ai_1 _06721_ (.B1(net74),
    .Y(_01178_),
    .A1(net201),
    .A2(_01005_));
 sg13g2_a221oi_1 _06722_ (.B2(net57),
    .C1(_01178_),
    .B1(_00555_),
    .A1(net130),
    .Y(_01179_),
    .A2(net133));
 sg13g2_nor2_1 _06723_ (.A(_00547_),
    .B(_01036_),
    .Y(_01180_));
 sg13g2_nor2_1 _06724_ (.A(_00878_),
    .B(_01180_),
    .Y(_01181_));
 sg13g2_or4_1 _06725_ (.A(net344),
    .B(_01032_),
    .C(_01179_),
    .D(_01181_),
    .X(_01182_));
 sg13g2_nand3_1 _06726_ (.B(_01177_),
    .C(_01182_),
    .A(net375),
    .Y(_01183_));
 sg13g2_o21ai_1 _06727_ (.B1(_05383_),
    .Y(_01184_),
    .A1(net51),
    .A2(_01183_));
 sg13g2_a221oi_1 _06728_ (.B2(_00841_),
    .C1(_01184_),
    .B1(_01171_),
    .A1(_00645_),
    .Y(_01185_),
    .A2(_01156_));
 sg13g2_nor4_1 _06729_ (.A(_00950_),
    .B(_00948_),
    .C(_01140_),
    .D(_01185_),
    .Y(_01186_));
 sg13g2_a21oi_1 _06730_ (.A1(_00844_),
    .A2(_00949_),
    .Y(_01187_),
    .B1(_01186_));
 sg13g2_nor3_1 _06731_ (.A(_00399_),
    .B(_00402_),
    .C(_01187_),
    .Y(_01188_));
 sg13g2_buf_1 _06732_ (.A(net419),
    .X(_01189_));
 sg13g2_mux2_1 _06733_ (.A0(\dtop.vtop.logo_d[1] ),
    .A1(_01188_),
    .S(net374),
    .X(_00096_));
 sg13g2_o21ai_1 _06734_ (.B1(_05134_),
    .Y(_01190_),
    .A1(_05151_),
    .A2(_05386_));
 sg13g2_buf_2 _06735_ (.A(_01190_),
    .X(_01191_));
 sg13g2_nand3b_1 _06736_ (.B(_05129_),
    .C(_05131_),
    .Y(_01192_),
    .A_N(_05130_));
 sg13g2_buf_2 _06737_ (.A(_01192_),
    .X(_01193_));
 sg13g2_nand4_1 _06738_ (.B(_05149_),
    .C(_05136_),
    .A(_05253_),
    .Y(_01194_),
    .D(_05151_));
 sg13g2_buf_1 _06739_ (.A(_01194_),
    .X(_01195_));
 sg13g2_o21ai_1 _06740_ (.B1(_05146_),
    .Y(_01196_),
    .A1(_01193_),
    .A2(_01195_));
 sg13g2_buf_1 _06741_ (.A(_01196_),
    .X(_01197_));
 sg13g2_nand2_1 _06742_ (.Y(_01198_),
    .A(_01191_),
    .B(net296));
 sg13g2_nand2b_1 _06743_ (.Y(_01199_),
    .B(_05197_),
    .A_N(_05130_));
 sg13g2_nor2_1 _06744_ (.A(net402),
    .B(_01199_),
    .Y(_01200_));
 sg13g2_buf_1 _06745_ (.A(_01200_),
    .X(_01201_));
 sg13g2_nand2b_1 _06746_ (.Y(_01202_),
    .B(_00501_),
    .A_N(net383));
 sg13g2_buf_1 _06747_ (.A(_01202_),
    .X(_01203_));
 sg13g2_nor2_1 _06748_ (.A(net417),
    .B(net318),
    .Y(_01204_));
 sg13g2_buf_2 _06749_ (.A(_01204_),
    .X(_01205_));
 sg13g2_nand2_1 _06750_ (.Y(_01206_),
    .A(_05158_),
    .B(_05138_));
 sg13g2_buf_1 _06751_ (.A(_01206_),
    .X(_01207_));
 sg13g2_nand2b_1 _06752_ (.Y(_01208_),
    .B(net429),
    .A_N(net381));
 sg13g2_buf_2 _06753_ (.A(_01208_),
    .X(_01209_));
 sg13g2_nor2_2 _06754_ (.A(net342),
    .B(_01209_),
    .Y(_01210_));
 sg13g2_nand2b_1 _06755_ (.Y(_01211_),
    .B(_05158_),
    .A_N(_05138_));
 sg13g2_buf_2 _06756_ (.A(_01211_),
    .X(_01212_));
 sg13g2_nor2_1 _06757_ (.A(_01212_),
    .B(_01209_),
    .Y(_01213_));
 sg13g2_buf_1 _06758_ (.A(net417),
    .X(_01214_));
 sg13g2_nand2b_1 _06759_ (.Y(_01215_),
    .B(net383),
    .A_N(net418));
 sg13g2_buf_1 _06760_ (.A(_01215_),
    .X(_01216_));
 sg13g2_nor2_1 _06761_ (.A(net373),
    .B(_01216_),
    .Y(_01217_));
 sg13g2_buf_1 _06762_ (.A(_01217_),
    .X(_01218_));
 sg13g2_a22oi_1 _06763_ (.Y(_01219_),
    .B1(_01213_),
    .B2(net285),
    .A2(_01210_),
    .A1(_01205_));
 sg13g2_buf_1 _06764_ (.A(_01219_),
    .X(_01220_));
 sg13g2_nand2_1 _06765_ (.Y(_01221_),
    .A(_05151_),
    .B(_05386_));
 sg13g2_a22oi_1 _06766_ (.Y(_01222_),
    .B1(_01195_),
    .B2(_05134_),
    .A2(_01193_),
    .A1(_05146_));
 sg13g2_buf_1 _06767_ (.A(_01222_),
    .X(_01223_));
 sg13g2_nor2_1 _06768_ (.A(_01221_),
    .B(_01223_),
    .Y(_01224_));
 sg13g2_buf_1 _06769_ (.A(_01224_),
    .X(_01225_));
 sg13g2_nand2_1 _06770_ (.Y(_01226_),
    .A(_01220_),
    .B(net274));
 sg13g2_nor2b_1 _06771_ (.A(_05385_),
    .B_N(_05152_),
    .Y(_01227_));
 sg13g2_nand2b_1 _06772_ (.Y(_01228_),
    .B(_01227_),
    .A_N(_01223_));
 sg13g2_buf_1 _06773_ (.A(_01195_),
    .X(_01229_));
 sg13g2_o21ai_1 _06774_ (.B1(net328),
    .Y(_01230_),
    .A1(_01199_),
    .A2(net317));
 sg13g2_o21ai_1 _06775_ (.B1(_05386_),
    .Y(_01231_),
    .A1(_05146_),
    .A2(_01195_));
 sg13g2_a21oi_1 _06776_ (.A1(net402),
    .A2(_01230_),
    .Y(_01232_),
    .B1(_01231_));
 sg13g2_buf_2 _06777_ (.A(_01232_),
    .X(_01233_));
 sg13g2_nor2_1 _06778_ (.A(net418),
    .B(net383),
    .Y(_01234_));
 sg13g2_buf_1 _06779_ (.A(_01234_),
    .X(_01235_));
 sg13g2_nand2_2 _06780_ (.Y(_01236_),
    .A(net377),
    .B(net316));
 sg13g2_nand3_1 _06781_ (.B(_05160_),
    .C(net358),
    .A(net397),
    .Y(_01237_));
 sg13g2_nor2b_1 _06782_ (.A(net383),
    .B_N(net418),
    .Y(_01238_));
 sg13g2_buf_1 _06783_ (.A(_01238_),
    .X(_01239_));
 sg13g2_nor2_1 _06784_ (.A(_05138_),
    .B(\dtop.player_inst.program_addr[6] ),
    .Y(_01240_));
 sg13g2_and2_1 _06785_ (.A(_05155_),
    .B(_05158_),
    .X(_01241_));
 sg13g2_buf_1 _06786_ (.A(_01241_),
    .X(_01242_));
 sg13g2_nand3_1 _06787_ (.B(_01240_),
    .C(_01242_),
    .A(_01239_),
    .Y(_01243_));
 sg13g2_buf_1 _06788_ (.A(_01243_),
    .X(_01244_));
 sg13g2_o21ai_1 _06789_ (.B1(_01244_),
    .Y(_01245_),
    .A1(_01236_),
    .A2(_01237_));
 sg13g2_nand3_1 _06790_ (.B(_01233_),
    .C(_01245_),
    .A(_01228_),
    .Y(_01246_));
 sg13g2_nand2_1 _06791_ (.Y(_01247_),
    .A(net429),
    .B(net381));
 sg13g2_nor2_1 _06792_ (.A(_01247_),
    .B(net342),
    .Y(_01248_));
 sg13g2_buf_2 _06793_ (.A(_01248_),
    .X(_01249_));
 sg13g2_and2_1 _06794_ (.A(net416),
    .B(net316),
    .X(_01250_));
 sg13g2_buf_2 _06795_ (.A(_01250_),
    .X(_01251_));
 sg13g2_or2_1 _06796_ (.X(_01252_),
    .B(net417),
    .A(net358));
 sg13g2_buf_2 _06797_ (.A(_01252_),
    .X(_01253_));
 sg13g2_nor4_1 _06798_ (.A(net354),
    .B(_00441_),
    .C(net318),
    .D(_01253_),
    .Y(_01254_));
 sg13g2_a22oi_1 _06799_ (.Y(_01255_),
    .B1(_01254_),
    .B2(net322),
    .A2(_01251_),
    .A1(_01249_));
 sg13g2_buf_1 _06800_ (.A(_01255_),
    .X(_01256_));
 sg13g2_inv_1 _06801_ (.Y(_01257_),
    .A(_01256_));
 sg13g2_a21oi_1 _06802_ (.A1(_01226_),
    .A2(_01246_),
    .Y(_01258_),
    .B1(_01257_));
 sg13g2_and2_1 _06803_ (.A(net329),
    .B(_01242_),
    .X(_01259_));
 sg13g2_a21oi_1 _06804_ (.A1(_01251_),
    .A2(_01259_),
    .Y(_01260_),
    .B1(_01254_));
 sg13g2_or3_1 _06805_ (.A(net397),
    .B(net381),
    .C(net396),
    .X(_01261_));
 sg13g2_buf_1 _06806_ (.A(_01261_),
    .X(_01262_));
 sg13g2_nor2b_1 _06807_ (.A(net418),
    .B_N(net416),
    .Y(_01263_));
 sg13g2_a22oi_1 _06808_ (.Y(_01264_),
    .B1(_01263_),
    .B2(net400),
    .A2(_01240_),
    .A1(net380));
 sg13g2_buf_1 _06809_ (.A(_01264_),
    .X(_01265_));
 sg13g2_nor3_2 _06810_ (.A(net349),
    .B(_01262_),
    .C(_01265_),
    .Y(_01266_));
 sg13g2_nor2b_1 _06811_ (.A(_01266_),
    .B_N(_01256_),
    .Y(_01267_));
 sg13g2_nor4_1 _06812_ (.A(net274),
    .B(_01233_),
    .C(_01260_),
    .D(_01267_),
    .Y(_01268_));
 sg13g2_nor3_1 _06813_ (.A(_01201_),
    .B(_01258_),
    .C(_01268_),
    .Y(_01269_));
 sg13g2_and3_1 _06814_ (.X(_01270_),
    .A(net418),
    .B(_05171_),
    .C(net416));
 sg13g2_buf_1 _06815_ (.A(_01270_),
    .X(_01271_));
 sg13g2_buf_1 _06816_ (.A(_01271_),
    .X(_01272_));
 sg13g2_buf_1 _06817_ (.A(net315),
    .X(_01273_));
 sg13g2_or2_1 _06818_ (.X(_01274_),
    .B(net400),
    .A(net396));
 sg13g2_buf_2 _06819_ (.A(_01274_),
    .X(_01275_));
 sg13g2_mux2_1 _06820_ (.A0(_01207_),
    .A1(_01275_),
    .S(net322),
    .X(_01276_));
 sg13g2_and2_1 _06821_ (.A(net396),
    .B(_05138_),
    .X(_01277_));
 sg13g2_buf_1 _06822_ (.A(_01277_),
    .X(_01278_));
 sg13g2_a21oi_1 _06823_ (.A1(net322),
    .A2(net314),
    .Y(_01279_),
    .B1(net325));
 sg13g2_xnor2_1 _06824_ (.Y(_01280_),
    .A(_05159_),
    .B(net400));
 sg13g2_or2_1 _06825_ (.X(_01281_),
    .B(_01280_),
    .A(net322));
 sg13g2_a22oi_1 _06826_ (.Y(_01282_),
    .B1(_01279_),
    .B2(_01281_),
    .A2(_01276_),
    .A1(net325));
 sg13g2_nand2_1 _06827_ (.Y(_01283_),
    .A(net295),
    .B(_01282_));
 sg13g2_nor2b_1 _06828_ (.A(net417),
    .B_N(_05138_),
    .Y(_01284_));
 sg13g2_buf_1 _06829_ (.A(_01284_),
    .X(_01285_));
 sg13g2_nor2b_1 _06830_ (.A(net322),
    .B_N(net355),
    .Y(_01286_));
 sg13g2_buf_1 _06831_ (.A(_01216_),
    .X(_01287_));
 sg13g2_o21ai_1 _06832_ (.B1(net294),
    .Y(_01288_),
    .A1(net356),
    .A2(net318));
 sg13g2_nor2_1 _06833_ (.A(net429),
    .B(net381),
    .Y(_01289_));
 sg13g2_buf_1 _06834_ (.A(_01289_),
    .X(_01290_));
 sg13g2_nor3_1 _06835_ (.A(net327),
    .B(net318),
    .C(net313),
    .Y(_01291_));
 sg13g2_a21o_1 _06836_ (.A2(_01288_),
    .A1(_01286_),
    .B1(_01291_),
    .X(_01292_));
 sg13g2_buf_1 _06837_ (.A(net373),
    .X(_01293_));
 sg13g2_nand2_1 _06838_ (.Y(_01294_),
    .A(net341),
    .B(net316));
 sg13g2_nand2_1 _06839_ (.Y(_01295_),
    .A(net315),
    .B(_01242_));
 sg13g2_o21ai_1 _06840_ (.B1(_01295_),
    .Y(_01296_),
    .A1(_01294_),
    .A2(_01262_));
 sg13g2_nand3b_1 _06841_ (.B(_00418_),
    .C(net417),
    .Y(_01297_),
    .A_N(net380));
 sg13g2_buf_2 _06842_ (.A(_01297_),
    .X(_01298_));
 sg13g2_nor2b_1 _06843_ (.A(_05138_),
    .B_N(_05158_),
    .Y(_01299_));
 sg13g2_buf_2 _06844_ (.A(_01299_),
    .X(_01300_));
 sg13g2_nor2b_1 _06845_ (.A(_05158_),
    .B_N(_05138_),
    .Y(_01301_));
 sg13g2_buf_1 _06846_ (.A(_01301_),
    .X(_01302_));
 sg13g2_buf_1 _06847_ (.A(_01302_),
    .X(_01303_));
 sg13g2_a22oi_1 _06848_ (.Y(_01304_),
    .B1(net313),
    .B2(_01303_),
    .A2(_01300_),
    .A1(net356));
 sg13g2_and3_1 _06849_ (.X(_01305_),
    .A(net380),
    .B(_00419_),
    .C(net356));
 sg13g2_nor3_1 _06850_ (.A(_00502_),
    .B(_00419_),
    .C(_05157_),
    .Y(_01306_));
 sg13g2_and4_1 _06851_ (.A(net416),
    .B(net347),
    .C(_05160_),
    .D(net329),
    .X(_01307_));
 sg13g2_o21ai_1 _06852_ (.B1(_01307_),
    .Y(_01308_),
    .A1(_01305_),
    .A2(_01306_));
 sg13g2_o21ai_1 _06853_ (.B1(_01308_),
    .Y(_01309_),
    .A1(_01298_),
    .A2(_01304_));
 sg13g2_a221oi_1 _06854_ (.B2(_05181_),
    .C1(_01309_),
    .B1(_01296_),
    .A1(_01285_),
    .Y(_01310_),
    .A2(_01292_));
 sg13g2_or2_1 _06855_ (.X(_01311_),
    .B(_05171_),
    .A(net418));
 sg13g2_buf_2 _06856_ (.A(_01311_),
    .X(_01312_));
 sg13g2_nand2b_1 _06857_ (.Y(_01313_),
    .B(net417),
    .A_N(net400));
 sg13g2_nand2b_1 _06858_ (.Y(_01314_),
    .B(net429),
    .A_N(_05158_));
 sg13g2_buf_1 _06859_ (.A(_01314_),
    .X(_01315_));
 sg13g2_nor3_2 _06860_ (.A(_01312_),
    .B(_01313_),
    .C(_01315_),
    .Y(_01316_));
 sg13g2_nand2_1 _06861_ (.Y(_01317_),
    .A(net323),
    .B(_01316_));
 sg13g2_and3_1 _06862_ (.X(_01318_),
    .A(_01256_),
    .B(_01220_),
    .C(_01317_));
 sg13g2_buf_1 _06863_ (.A(_01318_),
    .X(_01319_));
 sg13g2_nor2_1 _06864_ (.A(_05159_),
    .B(_05139_),
    .Y(_01320_));
 sg13g2_nor2b_1 _06865_ (.A(net418),
    .B_N(_05171_),
    .Y(_01321_));
 sg13g2_buf_1 _06866_ (.A(_01321_),
    .X(_01322_));
 sg13g2_nor2b_1 _06867_ (.A(_00432_),
    .B_N(_05155_),
    .Y(_01323_));
 sg13g2_buf_2 _06868_ (.A(_01323_),
    .X(_01324_));
 sg13g2_nand4_1 _06869_ (.B(_01320_),
    .C(net340),
    .A(_00512_),
    .Y(_01325_),
    .D(_01324_));
 sg13g2_nand3_1 _06870_ (.B(_01271_),
    .C(_01302_),
    .A(net348),
    .Y(_01326_));
 sg13g2_nand4_1 _06871_ (.B(_01234_),
    .C(_01289_),
    .A(_00512_),
    .Y(_01327_),
    .D(_01302_));
 sg13g2_nand3_1 _06872_ (.B(_01326_),
    .C(_01327_),
    .A(_01325_),
    .Y(_01328_));
 sg13g2_buf_1 _06873_ (.A(_01328_),
    .X(_01329_));
 sg13g2_nand4_1 _06874_ (.B(net314),
    .C(net316),
    .A(net377),
    .Y(_01330_),
    .D(_01324_));
 sg13g2_o21ai_1 _06875_ (.B1(_01330_),
    .Y(_01331_),
    .A1(net299),
    .A2(_01244_));
 sg13g2_nor2_1 _06876_ (.A(net379),
    .B(_01216_),
    .Y(_01332_));
 sg13g2_buf_1 _06877_ (.A(_01332_),
    .X(_01333_));
 sg13g2_xor2_1 _06878_ (.B(net358),
    .A(net347),
    .X(_01334_));
 sg13g2_nor3_1 _06879_ (.A(net298),
    .B(net302),
    .C(_01334_),
    .Y(_01335_));
 sg13g2_and2_1 _06880_ (.A(net284),
    .B(_01335_),
    .X(_01336_));
 sg13g2_nor3_1 _06881_ (.A(_01329_),
    .B(_01331_),
    .C(_01336_),
    .Y(_01337_));
 sg13g2_and4_1 _06882_ (.A(_01283_),
    .B(_01310_),
    .C(_01319_),
    .D(_01337_),
    .X(_01338_));
 sg13g2_nor2b_1 _06883_ (.A(net304),
    .B_N(net325),
    .Y(_01339_));
 sg13g2_buf_1 _06884_ (.A(net341),
    .X(_01340_));
 sg13g2_nor2b_1 _06885_ (.A(net298),
    .B_N(net311),
    .Y(_01341_));
 sg13g2_nor3_1 _06886_ (.A(net294),
    .B(_01339_),
    .C(_01341_),
    .Y(_01342_));
 sg13g2_nor3_1 _06887_ (.A(net298),
    .B(net318),
    .C(_01313_),
    .Y(_01343_));
 sg13g2_o21ai_1 _06888_ (.B1(net300),
    .Y(_01344_),
    .A1(_01342_),
    .A2(_01343_));
 sg13g2_nor2_1 _06889_ (.A(net318),
    .B(_01253_),
    .Y(_01345_));
 sg13g2_or2_1 _06890_ (.X(_01346_),
    .B(_00432_),
    .A(\dtop.player_inst.program_addr[1] ));
 sg13g2_buf_1 _06891_ (.A(_01346_),
    .X(_01347_));
 sg13g2_nor2_1 _06892_ (.A(_01212_),
    .B(_01347_),
    .Y(_01348_));
 sg13g2_buf_1 _06893_ (.A(_01348_),
    .X(_01349_));
 sg13g2_a22oi_1 _06894_ (.Y(_01350_),
    .B1(net293),
    .B2(net284),
    .A2(_01345_),
    .A1(_05163_));
 sg13g2_nor2_1 _06895_ (.A(_00502_),
    .B(net323),
    .Y(_01351_));
 sg13g2_nand2b_1 _06896_ (.Y(_01352_),
    .B(net349),
    .A_N(net358));
 sg13g2_nand3b_1 _06897_ (.B(net355),
    .C(net358),
    .Y(_01353_),
    .A_N(net349));
 sg13g2_o21ai_1 _06898_ (.B1(_01353_),
    .Y(_01354_),
    .A1(net327),
    .A2(_01352_));
 sg13g2_nand4_1 _06899_ (.B(net311),
    .C(_01351_),
    .A(net298),
    .Y(_01355_),
    .D(_01354_));
 sg13g2_nand3_1 _06900_ (.B(_01350_),
    .C(_01355_),
    .A(_01344_),
    .Y(_01356_));
 sg13g2_nand3_1 _06901_ (.B(net312),
    .C(_01324_),
    .A(net315),
    .Y(_01357_));
 sg13g2_buf_1 _06902_ (.A(_01320_),
    .X(_01358_));
 sg13g2_nor2b_1 _06903_ (.A(net429),
    .B_N(_00432_),
    .Y(_01359_));
 sg13g2_buf_2 _06904_ (.A(_01359_),
    .X(_01360_));
 sg13g2_nand4_1 _06905_ (.B(net310),
    .C(net340),
    .A(net311),
    .Y(_01361_),
    .D(_01360_));
 sg13g2_nand4_1 _06906_ (.B(net316),
    .C(_01300_),
    .A(_00522_),
    .Y(_01362_),
    .D(_01324_));
 sg13g2_nand3_1 _06907_ (.B(_01361_),
    .C(_01362_),
    .A(_01357_),
    .Y(_01363_));
 sg13g2_nand3_1 _06908_ (.B(_05140_),
    .C(net417),
    .A(net383),
    .Y(_01364_));
 sg13g2_o21ai_1 _06909_ (.B1(_01364_),
    .Y(_01365_),
    .A1(net358),
    .A2(_05173_));
 sg13g2_nand3_1 _06910_ (.B(_05163_),
    .C(_01365_),
    .A(net321),
    .Y(_01366_));
 sg13g2_nand2b_1 _06911_ (.Y(_01367_),
    .B(_01366_),
    .A_N(_01363_));
 sg13g2_buf_1 _06912_ (.A(_01347_),
    .X(_01368_));
 sg13g2_nand3_1 _06913_ (.B(net291),
    .C(net311),
    .A(_00464_),
    .Y(_01369_));
 sg13g2_o21ai_1 _06914_ (.B1(_01369_),
    .Y(_01370_),
    .A1(_01253_),
    .A2(net309));
 sg13g2_nor2b_1 _06915_ (.A(net341),
    .B_N(net356),
    .Y(_01371_));
 sg13g2_nor2b_1 _06916_ (.A(_01286_),
    .B_N(_01371_),
    .Y(_01372_));
 sg13g2_a22oi_1 _06917_ (.Y(_01373_),
    .B1(_01372_),
    .B2(net326),
    .A2(_01370_),
    .A1(net302));
 sg13g2_nor2_1 _06918_ (.A(_00513_),
    .B(_01312_),
    .Y(_01374_));
 sg13g2_buf_2 _06919_ (.A(_01374_),
    .X(_01375_));
 sg13g2_o21ai_1 _06920_ (.B1(net327),
    .Y(_01376_),
    .A1(net356),
    .A2(net322));
 sg13g2_and3_1 _06921_ (.X(_01377_),
    .A(net329),
    .B(_01262_),
    .C(_01376_));
 sg13g2_nand3_1 _06922_ (.B(_00418_),
    .C(net416),
    .A(_00501_),
    .Y(_01378_));
 sg13g2_buf_2 _06923_ (.A(_01378_),
    .X(_01379_));
 sg13g2_nor3_1 _06924_ (.A(net348),
    .B(_01379_),
    .C(_01275_),
    .Y(_01380_));
 sg13g2_a221oi_1 _06925_ (.B2(_01377_),
    .C1(_01380_),
    .B1(_01375_),
    .A1(_01249_),
    .Y(_01381_),
    .A2(_01205_));
 sg13g2_o21ai_1 _06926_ (.B1(_01381_),
    .Y(_01382_),
    .A1(net294),
    .A2(_01373_));
 sg13g2_xor2_1 _06927_ (.B(_00433_),
    .A(_05156_),
    .X(_01383_));
 sg13g2_buf_2 _06928_ (.A(_01383_),
    .X(_01384_));
 sg13g2_or2_1 _06929_ (.X(_01385_),
    .B(_01384_),
    .A(net326));
 sg13g2_nor3_1 _06930_ (.A(_00441_),
    .B(net346),
    .C(_01312_),
    .Y(_01386_));
 sg13g2_nor4_2 _06931_ (.A(net346),
    .B(_01203_),
    .C(_01275_),
    .Y(_01387_),
    .D(_01209_));
 sg13g2_a21oi_1 _06932_ (.A1(_01385_),
    .A2(_01386_),
    .Y(_01388_),
    .B1(_01387_));
 sg13g2_nor2_1 _06933_ (.A(net329),
    .B(net379),
    .Y(_01389_));
 sg13g2_mux2_1 _06934_ (.A0(_00441_),
    .A1(_05163_),
    .S(net324),
    .X(_01390_));
 sg13g2_nand3_1 _06935_ (.B(_01351_),
    .C(_01390_),
    .A(_01389_),
    .Y(_01391_));
 sg13g2_nand4_1 _06936_ (.B(_01239_),
    .C(_01289_),
    .A(net379),
    .Y(_01392_),
    .D(_01302_));
 sg13g2_nand4_1 _06937_ (.B(net314),
    .C(net316),
    .A(net416),
    .Y(_01393_),
    .D(net313));
 sg13g2_nand4_1 _06938_ (.B(_01239_),
    .C(_01358_),
    .A(net379),
    .Y(_01394_),
    .D(net309));
 sg13g2_nand4_1 _06939_ (.B(_01235_),
    .C(net309),
    .A(_00521_),
    .Y(_01395_),
    .D(net312));
 sg13g2_and4_1 _06940_ (.A(_01392_),
    .B(_01393_),
    .C(_01394_),
    .D(_01395_),
    .X(_01396_));
 sg13g2_buf_1 _06941_ (.A(_01396_),
    .X(_01397_));
 sg13g2_buf_8 _06942_ (.A(_01247_),
    .X(_01398_));
 sg13g2_nor2_1 _06943_ (.A(net308),
    .B(_01275_),
    .Y(_01399_));
 sg13g2_nor2_1 _06944_ (.A(net346),
    .B(net318),
    .Y(_01400_));
 sg13g2_nand4_1 _06945_ (.B(net324),
    .C(net377),
    .A(net345),
    .Y(_01401_),
    .D(net329));
 sg13g2_buf_1 _06946_ (.A(_01401_),
    .X(_01402_));
 sg13g2_xnor2_1 _06947_ (.Y(_01403_),
    .A(net347),
    .B(net355));
 sg13g2_nor3_1 _06948_ (.A(_00464_),
    .B(_01402_),
    .C(_01403_),
    .Y(_01404_));
 sg13g2_a221oi_1 _06949_ (.B2(_01400_),
    .C1(_01404_),
    .B1(_01399_),
    .A1(_01251_),
    .Y(_01405_),
    .A2(net310));
 sg13g2_nand4_1 _06950_ (.B(_01391_),
    .C(_01397_),
    .A(_01388_),
    .Y(_01406_),
    .D(_01405_));
 sg13g2_nor4_2 _06951_ (.A(_01356_),
    .B(_01367_),
    .C(_01382_),
    .Y(_01407_),
    .D(_01406_));
 sg13g2_nand2b_1 _06952_ (.Y(_01408_),
    .B(_00433_),
    .A_N(net429));
 sg13g2_buf_2 _06953_ (.A(_01408_),
    .X(_01409_));
 sg13g2_nor2_1 _06954_ (.A(_01212_),
    .B(_01409_),
    .Y(_01410_));
 sg13g2_o21ai_1 _06955_ (.B1(_01410_),
    .Y(_01411_),
    .A1(_01273_),
    .A2(net285));
 sg13g2_nand2_1 _06956_ (.Y(_01412_),
    .A(net381),
    .B(net396));
 sg13g2_nand2_1 _06957_ (.Y(_01413_),
    .A(_00503_),
    .B(net397));
 sg13g2_nor2b_1 _06958_ (.A(net383),
    .B_N(net416),
    .Y(_01414_));
 sg13g2_a22oi_1 _06959_ (.Y(_01415_),
    .B1(_01285_),
    .B2(net349),
    .A2(_01414_),
    .A1(_05180_));
 sg13g2_nor3_2 _06960_ (.A(_01412_),
    .B(_01413_),
    .C(_01415_),
    .Y(_01416_));
 sg13g2_nor2_1 _06961_ (.A(net342),
    .B(_01409_),
    .Y(_01417_));
 sg13g2_and2_1 _06962_ (.A(_01205_),
    .B(_01417_),
    .X(_01418_));
 sg13g2_nor4_2 _06963_ (.A(_01266_),
    .B(_01416_),
    .C(_01329_),
    .Y(_01419_),
    .D(_01418_));
 sg13g2_nand3_1 _06964_ (.B(_01419_),
    .C(_01319_),
    .A(_01411_),
    .Y(_01420_));
 sg13g2_a21o_1 _06965_ (.A2(_01407_),
    .A1(_01338_),
    .B1(_01420_),
    .X(_01421_));
 sg13g2_nor3_1 _06966_ (.A(net324),
    .B(net323),
    .C(_01265_),
    .Y(_01422_));
 sg13g2_nand3_1 _06967_ (.B(net340),
    .C(_01285_),
    .A(net323),
    .Y(_01423_));
 sg13g2_nand2b_1 _06968_ (.Y(_01424_),
    .B(_01423_),
    .A_N(_01422_));
 sg13g2_nand3b_1 _06969_ (.B(net377),
    .C(net329),
    .Y(_01425_),
    .A_N(net345));
 sg13g2_o21ai_1 _06970_ (.B1(_01425_),
    .Y(_01426_),
    .A1(net321),
    .A2(_01253_));
 sg13g2_nor2b_1 _06971_ (.A(net345),
    .B_N(net341),
    .Y(_01427_));
 sg13g2_nand2b_1 _06972_ (.Y(_01428_),
    .B(net400),
    .A_N(_05158_));
 sg13g2_buf_2 _06973_ (.A(_01428_),
    .X(_01429_));
 sg13g2_nand2_1 _06974_ (.Y(_01430_),
    .A(_01429_),
    .B(_01352_));
 sg13g2_a22oi_1 _06975_ (.Y(_01431_),
    .B1(_01427_),
    .B2(_01430_),
    .A2(_01426_),
    .A1(net302));
 sg13g2_nand2_1 _06976_ (.Y(_01432_),
    .A(_05180_),
    .B(_01427_));
 sg13g2_a21o_1 _06977_ (.A2(_01432_),
    .A1(net324),
    .B1(net299),
    .X(_01433_));
 sg13g2_nor3_1 _06978_ (.A(_01312_),
    .B(_01412_),
    .C(_01313_),
    .Y(_01434_));
 sg13g2_nor3_1 _06979_ (.A(net341),
    .B(net294),
    .C(_01429_),
    .Y(_01435_));
 sg13g2_nor3_1 _06980_ (.A(net298),
    .B(_01434_),
    .C(_01435_),
    .Y(_01436_));
 sg13g2_o21ai_1 _06981_ (.B1(_01436_),
    .Y(_01437_),
    .A1(_01431_),
    .A2(_01433_));
 sg13g2_nor3_1 _06982_ (.A(net324),
    .B(net327),
    .C(_01265_),
    .Y(_01438_));
 sg13g2_and2_1 _06983_ (.A(_05141_),
    .B(net373),
    .X(_01439_));
 sg13g2_a21oi_1 _06984_ (.A1(_00460_),
    .A2(_01240_),
    .Y(_01440_),
    .B1(_01439_));
 sg13g2_nor3_1 _06985_ (.A(_00441_),
    .B(net294),
    .C(_01440_),
    .Y(_01441_));
 sg13g2_and3_1 _06986_ (.X(_01442_),
    .A(net311),
    .B(_01351_),
    .C(_01354_));
 sg13g2_or4_1 _06987_ (.A(net354),
    .B(_01438_),
    .C(_01441_),
    .D(_01442_),
    .X(_01443_));
 sg13g2_inv_1 _06988_ (.Y(_01444_),
    .A(_01381_));
 sg13g2_a221oi_1 _06989_ (.B2(_01443_),
    .C1(_01444_),
    .B1(_01437_),
    .A1(net300),
    .Y(_01445_),
    .A2(_01424_));
 sg13g2_buf_1 _06990_ (.A(_01445_),
    .X(_01446_));
 sg13g2_a22oi_1 _06991_ (.Y(_01447_),
    .B1(_01410_),
    .B2(net295),
    .A2(_01377_),
    .A1(_01332_));
 sg13g2_nor2_1 _06992_ (.A(net323),
    .B(net304),
    .Y(_01448_));
 sg13g2_o21ai_1 _06993_ (.B1(net302),
    .Y(_01449_),
    .A1(net298),
    .A2(_01448_));
 sg13g2_nor2_2 _06994_ (.A(net397),
    .B(net396),
    .Y(_01450_));
 sg13g2_o21ai_1 _06995_ (.B1(net291),
    .Y(_01451_),
    .A1(_00435_),
    .A2(_01450_));
 sg13g2_nand3_1 _06996_ (.B(_01449_),
    .C(_01451_),
    .A(net285),
    .Y(_01452_));
 sg13g2_nand2b_1 _06997_ (.Y(_01453_),
    .B(net396),
    .A_N(net397));
 sg13g2_xnor2_1 _06998_ (.Y(_01454_),
    .A(net383),
    .B(net400));
 sg13g2_nor4_1 _06999_ (.A(net380),
    .B(_00434_),
    .C(_01453_),
    .D(_01454_),
    .Y(_01455_));
 sg13g2_buf_1 _07000_ (.A(_01239_),
    .X(_01456_));
 sg13g2_nor3_2 _07001_ (.A(net381),
    .B(net396),
    .C(_05139_),
    .Y(_01457_));
 sg13g2_nand3_1 _07002_ (.B(net292),
    .C(_01457_),
    .A(net325),
    .Y(_01458_));
 sg13g2_nand2b_1 _07003_ (.Y(_01459_),
    .B(_01458_),
    .A_N(_01455_));
 sg13g2_o21ai_1 _07004_ (.B1(_05205_),
    .Y(_01460_),
    .A1(_05180_),
    .A2(_01286_));
 sg13g2_o21ai_1 _07005_ (.B1(_01460_),
    .Y(_01461_),
    .A1(net291),
    .A2(_01403_));
 sg13g2_buf_1 _07006_ (.A(_01375_),
    .X(_01462_));
 sg13g2_a22oi_1 _07007_ (.Y(_01463_),
    .B1(_01461_),
    .B2(net283),
    .A2(_01459_),
    .A1(_01340_));
 sg13g2_and3_1 _07008_ (.X(_01464_),
    .A(_01447_),
    .B(_01452_),
    .C(_01463_));
 sg13g2_buf_1 _07009_ (.A(_01464_),
    .X(_01465_));
 sg13g2_nand3_1 _07010_ (.B(_01360_),
    .C(_01365_),
    .A(net321),
    .Y(_01466_));
 sg13g2_nand3_1 _07011_ (.B(_01251_),
    .C(_01324_),
    .A(_05180_),
    .Y(_01467_));
 sg13g2_a21o_1 _07012_ (.A2(_01467_),
    .A1(_01466_),
    .B1(_00441_),
    .X(_01468_));
 sg13g2_nor2_1 _07013_ (.A(net325),
    .B(net318),
    .Y(_01469_));
 sg13g2_mux2_1 _07014_ (.A0(_01212_),
    .A1(_01429_),
    .S(_00434_),
    .X(_01470_));
 sg13g2_nand2_1 _07015_ (.Y(_01471_),
    .A(net341),
    .B(net310));
 sg13g2_o21ai_1 _07016_ (.B1(_01471_),
    .Y(_01472_),
    .A1(net341),
    .A2(_01470_));
 sg13g2_a22oi_1 _07017_ (.Y(_01473_),
    .B1(net309),
    .B2(net327),
    .A2(_01236_),
    .A1(_05180_));
 sg13g2_nor2_1 _07018_ (.A(net327),
    .B(net309),
    .Y(_01474_));
 sg13g2_o21ai_1 _07019_ (.B1(net304),
    .Y(_01475_),
    .A1(_01379_),
    .A2(_01474_));
 sg13g2_a22oi_1 _07020_ (.Y(_01476_),
    .B1(net340),
    .B2(_01384_),
    .A2(net292),
    .A1(net348));
 sg13g2_nor2_1 _07021_ (.A(_01471_),
    .B(_01476_),
    .Y(_01477_));
 sg13g2_a221oi_1 _07022_ (.B2(_01475_),
    .C1(_01477_),
    .B1(_01473_),
    .A1(_01469_),
    .Y(_01478_),
    .A2(_01472_));
 sg13g2_and4_1 _07023_ (.A(_01468_),
    .B(_01478_),
    .C(_01283_),
    .D(_01310_),
    .X(_01479_));
 sg13g2_buf_1 _07024_ (.A(_01479_),
    .X(_01480_));
 sg13g2_nand3_1 _07025_ (.B(_01465_),
    .C(_01480_),
    .A(_01446_),
    .Y(_01481_));
 sg13g2_buf_2 _07026_ (.A(_01481_),
    .X(_01482_));
 sg13g2_mux2_1 _07027_ (.A0(_01269_),
    .A1(_01421_),
    .S(_01482_),
    .X(_01483_));
 sg13g2_buf_1 _07028_ (.A(_01483_),
    .X(_01484_));
 sg13g2_buf_1 _07029_ (.A(_01484_),
    .X(_01485_));
 sg13g2_nor2_1 _07030_ (.A(_05253_),
    .B(_05136_),
    .Y(_01486_));
 sg13g2_or2_1 _07031_ (.X(_01487_),
    .B(_01486_),
    .A(net305));
 sg13g2_nor2_1 _07032_ (.A(_05150_),
    .B(net398),
    .Y(_01488_));
 sg13g2_nor3_1 _07033_ (.A(net391),
    .B(net392),
    .C(net420),
    .Y(_01489_));
 sg13g2_o21ai_1 _07034_ (.B1(_01489_),
    .Y(_01490_),
    .A1(net305),
    .A2(_01488_));
 sg13g2_nand2_2 _07035_ (.Y(_01491_),
    .A(_01487_),
    .B(_01490_));
 sg13g2_and2_1 _07036_ (.A(_01319_),
    .B(_01337_),
    .X(_01492_));
 sg13g2_buf_1 _07037_ (.A(_01492_),
    .X(_01493_));
 sg13g2_nor2b_1 _07038_ (.A(net373),
    .B_N(net355),
    .Y(_01494_));
 sg13g2_nand3b_1 _07039_ (.B(_05140_),
    .C(net380),
    .Y(_01495_),
    .A_N(net349));
 sg13g2_o21ai_1 _07040_ (.B1(_01495_),
    .Y(_01496_),
    .A1(net345),
    .A2(_01352_));
 sg13g2_and3_1 _07041_ (.X(_01497_),
    .A(_01360_),
    .B(_01494_),
    .C(_01496_));
 sg13g2_nand2_1 _07042_ (.Y(_01498_),
    .A(_05151_),
    .B(_05134_));
 sg13g2_buf_2 _07043_ (.A(_01498_),
    .X(_01499_));
 sg13g2_a221oi_1 _07044_ (.B2(_01245_),
    .C1(_01201_),
    .B1(_01191_),
    .A1(_01497_),
    .Y(_01500_),
    .A2(_01499_));
 sg13g2_nor2_2 _07045_ (.A(_05151_),
    .B(_05385_),
    .Y(_01501_));
 sg13g2_and2_1 _07046_ (.A(_05134_),
    .B(_01501_),
    .X(_01502_));
 sg13g2_buf_1 _07047_ (.A(_01502_),
    .X(_01503_));
 sg13g2_nand3_1 _07048_ (.B(_01260_),
    .C(_01503_),
    .A(_01220_),
    .Y(_01504_));
 sg13g2_nand2b_1 _07049_ (.Y(_01505_),
    .B(net274),
    .A_N(_01220_));
 sg13g2_a21o_1 _07050_ (.A2(_01230_),
    .A1(net402),
    .B1(_01231_),
    .X(_01506_));
 sg13g2_buf_1 _07051_ (.A(_01506_),
    .X(_01507_));
 sg13g2_inv_1 _07052_ (.Y(_01508_),
    .A(_05151_));
 sg13g2_nor2_2 _07053_ (.A(_05196_),
    .B(_05147_),
    .Y(_01509_));
 sg13g2_nor2_1 _07054_ (.A(net372),
    .B(_01509_),
    .Y(_01510_));
 sg13g2_nand4_1 _07055_ (.B(_01220_),
    .C(_01507_),
    .A(_01256_),
    .Y(_01511_),
    .D(_01510_));
 sg13g2_and4_1 _07056_ (.A(_01500_),
    .B(_01504_),
    .C(_01505_),
    .D(_01511_),
    .X(_01512_));
 sg13g2_and4_1 _07057_ (.A(_01446_),
    .B(_01465_),
    .C(_01480_),
    .D(_01512_),
    .X(_01513_));
 sg13g2_buf_1 _07058_ (.A(_01513_),
    .X(_01514_));
 sg13g2_a21o_1 _07059_ (.A2(_01493_),
    .A1(_01482_),
    .B1(_01514_),
    .X(_01515_));
 sg13g2_buf_2 _07060_ (.A(_01515_),
    .X(_01516_));
 sg13g2_buf_1 _07061_ (.A(_01516_),
    .X(_01517_));
 sg13g2_nand2b_1 _07062_ (.Y(_01518_),
    .B(net104),
    .A_N(_01491_));
 sg13g2_nor2_1 _07063_ (.A(net105),
    .B(_01518_),
    .Y(_01519_));
 sg13g2_or3_1 _07064_ (.A(_01201_),
    .B(_01258_),
    .C(_01268_),
    .X(_01520_));
 sg13g2_buf_1 _07065_ (.A(_01520_),
    .X(_01521_));
 sg13g2_a21oi_2 _07066_ (.B1(_01420_),
    .Y(_01522_),
    .A2(_01407_),
    .A1(_01338_));
 sg13g2_mux2_1 _07067_ (.A0(_01521_),
    .A1(_01522_),
    .S(_01482_),
    .X(_01523_));
 sg13g2_buf_1 _07068_ (.A(_01523_),
    .X(_01524_));
 sg13g2_buf_1 _07069_ (.A(net129),
    .X(_01525_));
 sg13g2_nor2_1 _07070_ (.A(net402),
    .B(net317),
    .Y(_01526_));
 sg13g2_nor3_1 _07071_ (.A(net328),
    .B(_01126_),
    .C(_01526_),
    .Y(_01527_));
 sg13g2_buf_2 _07072_ (.A(_01527_),
    .X(_01528_));
 sg13g2_inv_1 _07073_ (.Y(_01529_),
    .A(_05331_));
 sg13g2_nand2_1 _07074_ (.Y(_01530_),
    .A(_00406_),
    .B(_01529_));
 sg13g2_o21ai_1 _07075_ (.B1(_01530_),
    .Y(_01531_),
    .A1(_01221_),
    .A2(_01223_));
 sg13g2_nand2_1 _07076_ (.Y(_01532_),
    .A(_05152_),
    .B(_05166_));
 sg13g2_nor2_1 _07077_ (.A(_00022_),
    .B(_05365_),
    .Y(_01533_));
 sg13g2_o21ai_1 _07078_ (.B1(_01533_),
    .Y(_01534_),
    .A1(net296),
    .A2(_01532_));
 sg13g2_buf_1 _07079_ (.A(_01534_),
    .X(_01535_));
 sg13g2_a21o_1 _07080_ (.A2(_01229_),
    .A1(_05199_),
    .B1(_05365_),
    .X(_01536_));
 sg13g2_nand3_1 _07081_ (.B(net424),
    .C(_01536_),
    .A(_05166_),
    .Y(_01537_));
 sg13g2_xor2_1 _07082_ (.B(net424),
    .A(_05165_),
    .X(_01538_));
 sg13g2_o21ai_1 _07083_ (.B1(_05135_),
    .Y(_01539_),
    .A1(_05366_),
    .A2(_01538_));
 sg13g2_a221oi_1 _07084_ (.B2(_01537_),
    .C1(_01539_),
    .B1(_01535_),
    .A1(_01528_),
    .Y(_01540_),
    .A2(_01531_));
 sg13g2_nand3b_1 _07085_ (.B(net274),
    .C(_01528_),
    .Y(_01541_),
    .A_N(net424));
 sg13g2_nand2b_1 _07086_ (.Y(_01542_),
    .B(_01541_),
    .A_N(_01540_));
 sg13g2_buf_2 _07087_ (.A(_01542_),
    .X(_01543_));
 sg13g2_nor2_1 _07088_ (.A(_01233_),
    .B(_01499_),
    .Y(_01544_));
 sg13g2_nor2_1 _07089_ (.A(_01193_),
    .B(net317),
    .Y(_01545_));
 sg13g2_nor2_1 _07090_ (.A(_05199_),
    .B(_01545_),
    .Y(_01546_));
 sg13g2_nor2_1 _07091_ (.A(_01191_),
    .B(_01530_),
    .Y(_01547_));
 sg13g2_or2_1 _07092_ (.X(_01548_),
    .B(_01547_),
    .A(_01225_));
 sg13g2_buf_1 _07093_ (.A(_01548_),
    .X(_01549_));
 sg13g2_nand2_1 _07094_ (.Y(_01550_),
    .A(net424),
    .B(_01227_));
 sg13g2_o21ai_1 _07095_ (.B1(_05366_),
    .Y(_01551_),
    .A1(net296),
    .A2(_01550_));
 sg13g2_nand2_1 _07096_ (.Y(_01552_),
    .A(_05166_),
    .B(_01551_));
 sg13g2_or4_1 _07097_ (.A(net328),
    .B(_01126_),
    .C(_01526_),
    .D(_01530_),
    .X(_01553_));
 sg13g2_nand2b_1 _07098_ (.Y(_01554_),
    .B(_05165_),
    .A_N(_05334_));
 sg13g2_a21oi_1 _07099_ (.A1(_05365_),
    .A2(_01554_),
    .Y(_01555_),
    .B1(_01509_));
 sg13g2_and3_1 _07100_ (.X(_01556_),
    .A(_01535_),
    .B(_01553_),
    .C(_01555_));
 sg13g2_buf_1 _07101_ (.A(_01556_),
    .X(_01557_));
 sg13g2_a22oi_1 _07102_ (.Y(_01558_),
    .B1(_01552_),
    .B2(_01557_),
    .A2(_01549_),
    .A1(_01528_));
 sg13g2_buf_1 _07103_ (.A(_01558_),
    .X(_01559_));
 sg13g2_o21ai_1 _07104_ (.B1(_01559_),
    .Y(_01560_),
    .A1(_01544_),
    .A2(_01546_));
 sg13g2_nor3_1 _07105_ (.A(net103),
    .B(_01543_),
    .C(_01560_),
    .Y(_01561_));
 sg13g2_a21oi_1 _07106_ (.A1(_05273_),
    .A2(_01525_),
    .Y(_01562_),
    .B1(_01561_));
 sg13g2_nor4_2 _07107_ (.A(net357),
    .B(net390),
    .C(net393),
    .Y(_01563_),
    .D(_05130_));
 sg13g2_nor2_1 _07108_ (.A(net398),
    .B(_05199_),
    .Y(_01564_));
 sg13g2_buf_1 _07109_ (.A(_01529_),
    .X(_01565_));
 sg13g2_xnor2_1 _07110_ (.Y(_01566_),
    .A(_05219_),
    .B(net420));
 sg13g2_buf_1 _07111_ (.A(_01566_),
    .X(_01567_));
 sg13g2_a21oi_1 _07112_ (.A1(net339),
    .A2(_01567_),
    .Y(_01568_),
    .B1(net350));
 sg13g2_nor2_2 _07113_ (.A(_05220_),
    .B(net420),
    .Y(_01569_));
 sg13g2_a21oi_1 _07114_ (.A1(net351),
    .A2(_00489_),
    .Y(_01570_),
    .B1(_01569_));
 sg13g2_o21ai_1 _07115_ (.B1(net350),
    .Y(_01571_),
    .A1(net386),
    .A2(_01529_));
 sg13g2_o21ai_1 _07116_ (.B1(_01571_),
    .Y(_01572_),
    .A1(net352),
    .A2(_01570_));
 sg13g2_o21ai_1 _07117_ (.B1(_01572_),
    .Y(_01573_),
    .A1(_01564_),
    .A2(_01568_));
 sg13g2_nor2_1 _07118_ (.A(_00406_),
    .B(_01567_),
    .Y(_01574_));
 sg13g2_nor2b_1 _07119_ (.A(_01574_),
    .B_N(_01564_),
    .Y(_01575_));
 sg13g2_nand3_1 _07120_ (.B(_01563_),
    .C(_01575_),
    .A(net339),
    .Y(_01576_));
 sg13g2_o21ai_1 _07121_ (.B1(_01576_),
    .Y(_01577_),
    .A1(_01563_),
    .A2(_01573_));
 sg13g2_buf_1 _07122_ (.A(_01577_),
    .X(_01578_));
 sg13g2_nand2_1 _07123_ (.Y(_01579_),
    .A(net399),
    .B(net398));
 sg13g2_buf_1 _07124_ (.A(_01579_),
    .X(_01580_));
 sg13g2_o21ai_1 _07125_ (.B1(net350),
    .Y(_01581_),
    .A1(net307),
    .A2(_00426_));
 sg13g2_o21ai_1 _07126_ (.B1(_01573_),
    .Y(_01582_),
    .A1(net339),
    .A2(_00472_));
 sg13g2_a22oi_1 _07127_ (.Y(_01583_),
    .B1(_01582_),
    .B2(net307),
    .A2(_01581_),
    .A1(net352));
 sg13g2_nand3_1 _07128_ (.B(net388),
    .C(_01567_),
    .A(net350),
    .Y(_01584_));
 sg13g2_o21ai_1 _07129_ (.B1(_01584_),
    .Y(_01585_),
    .A1(net352),
    .A2(_01575_));
 sg13g2_mux2_1 _07130_ (.A0(_01583_),
    .A1(_01585_),
    .S(_01563_),
    .X(_01586_));
 sg13g2_nand3_1 _07131_ (.B(_05221_),
    .C(_01229_),
    .A(_05254_),
    .Y(_01587_));
 sg13g2_nand2b_1 _07132_ (.Y(_01588_),
    .B(_01587_),
    .A_N(_01193_));
 sg13g2_buf_1 _07133_ (.A(_01588_),
    .X(_01589_));
 sg13g2_nor2_1 _07134_ (.A(\dtop.ext_control[2] ),
    .B(net276),
    .Y(_01590_));
 sg13g2_a22oi_1 _07135_ (.Y(_01591_),
    .B1(_01586_),
    .B2(_01590_),
    .A2(_01578_),
    .A1(\dtop.ext_control[2] ));
 sg13g2_a21oi_1 _07136_ (.A1(net276),
    .A2(_01578_),
    .Y(_01592_),
    .B1(net103));
 sg13g2_o21ai_1 _07137_ (.B1(_01592_),
    .Y(_01593_),
    .A1(\dtop.ext_control[0] ),
    .A2(_01591_));
 sg13g2_nand2_1 _07138_ (.Y(_01594_),
    .A(net104),
    .B(_01593_));
 sg13g2_o21ai_1 _07139_ (.B1(_01594_),
    .Y(_01595_),
    .A1(net104),
    .A2(_01562_));
 sg13g2_a21oi_1 _07140_ (.A1(_01482_),
    .A2(_01493_),
    .Y(_01596_),
    .B1(_01514_));
 sg13g2_buf_4 _07141_ (.X(_01597_),
    .A(_01596_));
 sg13g2_buf_1 _07142_ (.A(_01597_),
    .X(_01598_));
 sg13g2_nor2b_1 _07143_ (.A(_01193_),
    .B_N(_01587_),
    .Y(_01599_));
 sg13g2_buf_2 _07144_ (.A(_01599_),
    .X(_01600_));
 sg13g2_o21ai_1 _07145_ (.B1(_01600_),
    .Y(_01601_),
    .A1(_05216_),
    .A2(\dtop.ext_control[1] ));
 sg13g2_nand3_1 _07146_ (.B(_01598_),
    .C(_01601_),
    .A(net305),
    .Y(_01602_));
 sg13g2_nor2_1 _07147_ (.A(net103),
    .B(net104),
    .Y(_01603_));
 sg13g2_a21oi_1 _07148_ (.A1(_05385_),
    .A2(_01486_),
    .Y(_01604_),
    .B1(_05196_));
 sg13g2_nor2_1 _07149_ (.A(net328),
    .B(_01604_),
    .Y(_01605_));
 sg13g2_a21oi_2 _07150_ (.B1(_01605_),
    .Y(_01606_),
    .A2(net328),
    .A1(net390));
 sg13g2_a22oi_1 _07151_ (.Y(_01607_),
    .B1(_01603_),
    .B2(_01606_),
    .A2(_01602_),
    .A1(net103));
 sg13g2_a22oi_1 _07152_ (.Y(_01608_),
    .B1(_01595_),
    .B2(_01607_),
    .A2(_01519_),
    .A1(_01198_));
 sg13g2_buf_1 _07153_ (.A(_01608_),
    .X(_01609_));
 sg13g2_and3_1 _07154_ (.X(_01610_),
    .A(_01446_),
    .B(_01465_),
    .C(_01480_));
 sg13g2_buf_2 _07155_ (.A(_01610_),
    .X(_01611_));
 sg13g2_nand3b_1 _07156_ (.B(_01256_),
    .C(_01220_),
    .Y(_01612_),
    .A_N(_01266_));
 sg13g2_a21oi_1 _07157_ (.A1(_05196_),
    .A2(net317),
    .Y(_01613_),
    .B1(_05147_));
 sg13g2_a21oi_1 _07158_ (.A1(_05144_),
    .A2(net317),
    .Y(_01614_),
    .B1(_01199_));
 sg13g2_nor3_2 _07159_ (.A(_05385_),
    .B(_01613_),
    .C(_01614_),
    .Y(_01615_));
 sg13g2_o21ai_1 _07160_ (.B1(_01615_),
    .Y(_01616_),
    .A1(_01245_),
    .A2(_01510_));
 sg13g2_nor2_1 _07161_ (.A(_01612_),
    .B(_01616_),
    .Y(_01617_));
 sg13g2_nand2_1 _07162_ (.Y(_01618_),
    .A(net285),
    .B(_01417_));
 sg13g2_nand4_1 _07163_ (.B(net310),
    .C(_01322_),
    .A(_01214_),
    .Y(_01619_),
    .D(_01290_));
 sg13g2_nand2_1 _07164_ (.Y(_01620_),
    .A(_01618_),
    .B(_01619_));
 sg13g2_a21oi_2 _07165_ (.B1(_01620_),
    .Y(_01621_),
    .A2(_01617_),
    .A1(_01611_));
 sg13g2_buf_1 _07166_ (.A(_01621_),
    .X(_01622_));
 sg13g2_nor2_1 _07167_ (.A(net308),
    .B(_01429_),
    .Y(_01623_));
 sg13g2_nor3_1 _07168_ (.A(net308),
    .B(_01275_),
    .C(_01298_),
    .Y(_01624_));
 sg13g2_a21o_1 _07169_ (.A2(_01623_),
    .A1(_01375_),
    .B1(_01624_),
    .X(_01625_));
 sg13g2_nand4_1 _07170_ (.B(net292),
    .C(_01371_),
    .A(net304),
    .Y(_01626_),
    .D(_01403_));
 sg13g2_nand3_1 _07171_ (.B(net315),
    .C(net310),
    .A(net354),
    .Y(_01627_));
 sg13g2_nand3b_1 _07172_ (.B(_01626_),
    .C(_01627_),
    .Y(_01628_),
    .A_N(_01625_));
 sg13g2_buf_1 _07173_ (.A(_01628_),
    .X(_01629_));
 sg13g2_nor2_1 _07174_ (.A(_01429_),
    .B(_01209_),
    .Y(_01630_));
 sg13g2_nor3_1 _07175_ (.A(net342),
    .B(_01379_),
    .C(net309),
    .Y(_01631_));
 sg13g2_a221oi_1 _07176_ (.B2(_01630_),
    .C1(_01631_),
    .B1(_01375_),
    .A1(_01249_),
    .Y(_01632_),
    .A2(_01332_));
 sg13g2_buf_1 _07177_ (.A(_01632_),
    .X(_01633_));
 sg13g2_nor2_1 _07178_ (.A(net342),
    .B(net309),
    .Y(_01634_));
 sg13g2_and3_1 _07179_ (.X(_01635_),
    .A(_01278_),
    .B(net315),
    .C(_01384_));
 sg13g2_a221oi_1 _07180_ (.B2(_01375_),
    .C1(_01635_),
    .B1(_01634_),
    .A1(_01332_),
    .Y(_01636_),
    .A2(net293));
 sg13g2_nor2_1 _07181_ (.A(_01398_),
    .B(_01212_),
    .Y(_01637_));
 sg13g2_o21ai_1 _07182_ (.B1(net397),
    .Y(_01638_),
    .A1(net347),
    .A2(net358));
 sg13g2_and3_1 _07183_ (.X(_01639_),
    .A(net379),
    .B(net340),
    .C(_01638_));
 sg13g2_and4_1 _07184_ (.A(net347),
    .B(_01456_),
    .C(_01285_),
    .D(_01450_),
    .X(_01640_));
 sg13g2_a221oi_1 _07185_ (.B2(_00441_),
    .C1(_01640_),
    .B1(_01639_),
    .A1(net285),
    .Y(_01641_),
    .A2(_01637_));
 sg13g2_nand4_1 _07186_ (.B(_01633_),
    .C(_01636_),
    .A(_01397_),
    .Y(_01642_),
    .D(_01641_));
 sg13g2_buf_2 _07187_ (.A(_01642_),
    .X(_01643_));
 sg13g2_nand4_1 _07188_ (.B(_01235_),
    .C(_01300_),
    .A(_00521_),
    .Y(_01644_),
    .D(_01289_));
 sg13g2_nand4_1 _07189_ (.B(net314),
    .C(net340),
    .A(net373),
    .Y(_01645_),
    .D(net313));
 sg13g2_nand4_1 _07190_ (.B(_01234_),
    .C(_01300_),
    .A(net373),
    .Y(_01646_),
    .D(_01360_));
 sg13g2_nand3_1 _07191_ (.B(_01290_),
    .C(net312),
    .A(_01272_),
    .Y(_01647_));
 sg13g2_nand4_1 _07192_ (.B(_01645_),
    .C(_01646_),
    .A(_01644_),
    .Y(_01648_),
    .D(_01647_));
 sg13g2_buf_2 _07193_ (.A(_01648_),
    .X(_01649_));
 sg13g2_nor3_2 _07194_ (.A(_01629_),
    .B(_01643_),
    .C(_01649_),
    .Y(_01650_));
 sg13g2_nor3_2 _07195_ (.A(_05181_),
    .B(_01298_),
    .C(_01209_),
    .Y(_01651_));
 sg13g2_nand3_1 _07196_ (.B(_01365_),
    .C(_01450_),
    .A(net321),
    .Y(_01652_));
 sg13g2_nor2_1 _07197_ (.A(_01379_),
    .B(_01212_),
    .Y(_01653_));
 sg13g2_nor4_1 _07198_ (.A(net379),
    .B(_01312_),
    .C(_01275_),
    .D(_01409_),
    .Y(_01654_));
 sg13g2_a221oi_1 _07199_ (.B2(net354),
    .C1(_01654_),
    .B1(_01653_),
    .A1(_00434_),
    .Y(_01655_),
    .A2(_01316_));
 sg13g2_nand2_1 _07200_ (.Y(_01656_),
    .A(_01652_),
    .B(_01655_));
 sg13g2_buf_1 _07201_ (.A(_01656_),
    .X(_01657_));
 sg13g2_and2_1 _07202_ (.A(net292),
    .B(_01457_),
    .X(_01658_));
 sg13g2_o21ai_1 _07203_ (.B1(_01293_),
    .Y(_01659_),
    .A1(_01455_),
    .A2(_01658_));
 sg13g2_a21o_1 _07204_ (.A2(net314),
    .A1(net347),
    .B1(_01457_),
    .X(_01660_));
 sg13g2_nand3_1 _07205_ (.B(net315),
    .C(_01660_),
    .A(_05157_),
    .Y(_01661_));
 sg13g2_nand2_1 _07206_ (.Y(_01662_),
    .A(_01205_),
    .B(net293));
 sg13g2_and2_1 _07207_ (.A(net340),
    .B(_01334_),
    .X(_01663_));
 sg13g2_nor2_1 _07208_ (.A(_00434_),
    .B(_01495_),
    .Y(_01664_));
 sg13g2_nor2_1 _07209_ (.A(_01293_),
    .B(_01315_),
    .Y(_01665_));
 sg13g2_o21ai_1 _07210_ (.B1(_01665_),
    .Y(_01666_),
    .A1(_01663_),
    .A2(_01664_));
 sg13g2_nand4_1 _07211_ (.B(_01661_),
    .C(_01662_),
    .A(_01659_),
    .Y(_01667_),
    .D(_01666_));
 sg13g2_buf_1 _07212_ (.A(_01667_),
    .X(_01668_));
 sg13g2_nand3_1 _07213_ (.B(net316),
    .C(net310),
    .A(net341),
    .Y(_01669_));
 sg13g2_nor2_1 _07214_ (.A(net304),
    .B(_01379_),
    .Y(_01670_));
 sg13g2_nor3_1 _07215_ (.A(net326),
    .B(net346),
    .C(_01312_),
    .Y(_01671_));
 sg13g2_o21ai_1 _07216_ (.B1(net302),
    .Y(_01672_),
    .A1(_01670_),
    .A2(_01671_));
 sg13g2_a21oi_1 _07217_ (.A1(_01669_),
    .A2(_01672_),
    .Y(_01673_),
    .B1(net308));
 sg13g2_nor4_2 _07218_ (.A(_01651_),
    .B(net273),
    .C(net259),
    .Y(_01674_),
    .D(_01673_));
 sg13g2_nand2_1 _07219_ (.Y(_01675_),
    .A(_01650_),
    .B(_01674_));
 sg13g2_a21oi_1 _07220_ (.A1(_01466_),
    .A2(_01467_),
    .Y(_01676_),
    .B1(net300));
 sg13g2_nand2_1 _07221_ (.Y(_01677_),
    .A(_01375_),
    .B(_01259_));
 sg13g2_nand3_1 _07222_ (.B(net314),
    .C(net292),
    .A(net379),
    .Y(_01678_));
 sg13g2_a21o_1 _07223_ (.A2(_01678_),
    .A1(_01669_),
    .B1(_05205_),
    .X(_01679_));
 sg13g2_a21oi_2 _07224_ (.B1(net299),
    .Y(_01680_),
    .A2(_01679_),
    .A1(_01677_));
 sg13g2_nor2_1 _07225_ (.A(_01429_),
    .B(_01409_),
    .Y(_01681_));
 sg13g2_nand2_1 _07226_ (.Y(_01682_),
    .A(net315),
    .B(_01681_));
 sg13g2_nor2b_1 _07227_ (.A(net327),
    .B_N(net347),
    .Y(_01683_));
 sg13g2_a22oi_1 _07228_ (.Y(_01684_),
    .B1(_01683_),
    .B2(net292),
    .A2(_01242_),
    .A1(_00504_));
 sg13g2_nand2b_1 _07229_ (.Y(_01685_),
    .B(_01389_),
    .A_N(_01684_));
 sg13g2_a22oi_1 _07230_ (.Y(_01686_),
    .B1(_01410_),
    .B2(_01205_),
    .A2(_01399_),
    .A1(net315));
 sg13g2_o21ai_1 _07231_ (.B1(net285),
    .Y(_01687_),
    .A1(_01623_),
    .A2(net293));
 sg13g2_nand4_1 _07232_ (.B(_01685_),
    .C(_01686_),
    .A(_01682_),
    .Y(_01688_),
    .D(_01687_));
 sg13g2_nor2b_1 _07233_ (.A(net322),
    .B_N(net349),
    .Y(_01689_));
 sg13g2_a22oi_1 _07234_ (.Y(_01690_),
    .B1(_01371_),
    .B2(_01689_),
    .A2(_01360_),
    .A1(_01414_));
 sg13g2_or3_1 _07235_ (.A(net345),
    .B(net342),
    .C(_01690_),
    .X(_01691_));
 sg13g2_nand3_1 _07236_ (.B(_01691_),
    .C(_01361_),
    .A(_01357_),
    .Y(_01692_));
 sg13g2_nor4_2 _07237_ (.A(_01676_),
    .B(_01680_),
    .C(_01688_),
    .Y(_01693_),
    .D(_01692_));
 sg13g2_and2_1 _07238_ (.A(_01244_),
    .B(_01619_),
    .X(_01694_));
 sg13g2_o21ai_1 _07239_ (.B1(_01409_),
    .Y(_01695_),
    .A1(_05141_),
    .A2(_01209_));
 sg13g2_nor3_1 _07240_ (.A(_00441_),
    .B(_01214_),
    .C(_01287_),
    .Y(_01696_));
 sg13g2_nor2_1 _07241_ (.A(net349),
    .B(_01237_),
    .Y(_01697_));
 sg13g2_nor2_1 _07242_ (.A(_00459_),
    .B(net373),
    .Y(_01698_));
 sg13g2_a21o_1 _07243_ (.A2(_01698_),
    .A1(net380),
    .B1(_01263_),
    .X(_01699_));
 sg13g2_a22oi_1 _07244_ (.Y(_01700_),
    .B1(_01697_),
    .B2(_01699_),
    .A2(_01696_),
    .A1(_01695_));
 sg13g2_and4_1 _07245_ (.A(_01652_),
    .B(_01655_),
    .C(_01694_),
    .D(_01700_),
    .X(_01701_));
 sg13g2_nor2_1 _07246_ (.A(net347),
    .B(net355),
    .Y(_01702_));
 sg13g2_nand2_1 _07247_ (.Y(_01703_),
    .A(net316),
    .B(_01702_));
 sg13g2_nand3_1 _07248_ (.B(_00420_),
    .C(_05161_),
    .A(net345),
    .Y(_01704_));
 sg13g2_nand2_1 _07249_ (.Y(_01705_),
    .A(_00522_),
    .B(net356));
 sg13g2_a21oi_1 _07250_ (.A1(_01703_),
    .A2(_01704_),
    .Y(_01706_),
    .B1(_01705_));
 sg13g2_nor2b_1 _07251_ (.A(net355),
    .B_N(net373),
    .Y(_01707_));
 sg13g2_a22oi_1 _07252_ (.Y(_01708_),
    .B1(_01494_),
    .B2(net313),
    .A2(_01707_),
    .A1(net348));
 sg13g2_o21ai_1 _07253_ (.B1(_05142_),
    .Y(_01709_),
    .A1(_01287_),
    .A2(_01708_));
 sg13g2_o21ai_1 _07254_ (.B1(_01709_),
    .Y(_01710_),
    .A1(_05142_),
    .A2(_01706_));
 sg13g2_mux2_1 _07255_ (.A0(net312),
    .A1(_01280_),
    .S(_05156_),
    .X(_01711_));
 sg13g2_a21o_1 _07256_ (.A2(_01711_),
    .A1(_00460_),
    .B1(net293),
    .X(_01712_));
 sg13g2_a21oi_1 _07257_ (.A1(_01375_),
    .A2(_01712_),
    .Y(_01713_),
    .B1(_01649_));
 sg13g2_and4_1 _07258_ (.A(_01419_),
    .B(_01701_),
    .C(_01710_),
    .D(_01713_),
    .X(_01714_));
 sg13g2_buf_1 _07259_ (.A(_01714_),
    .X(_01715_));
 sg13g2_and2_1 _07260_ (.A(_01693_),
    .B(_01715_),
    .X(_01716_));
 sg13g2_buf_2 _07261_ (.A(_01716_),
    .X(_01717_));
 sg13g2_nor2_1 _07262_ (.A(_01629_),
    .B(_01643_),
    .Y(_01718_));
 sg13g2_and2_1 _07263_ (.A(_01419_),
    .B(_01701_),
    .X(_01719_));
 sg13g2_a21oi_1 _07264_ (.A1(_01462_),
    .A2(_01681_),
    .Y(_01720_),
    .B1(net259));
 sg13g2_and3_1 _07265_ (.X(_01721_),
    .A(_01718_),
    .B(_01719_),
    .C(_01720_));
 sg13g2_buf_1 _07266_ (.A(_01721_),
    .X(_01722_));
 sg13g2_o21ai_1 _07267_ (.B1(_01375_),
    .Y(_01723_),
    .A1(net293),
    .A2(_01681_));
 sg13g2_nand2b_1 _07268_ (.Y(_01724_),
    .B(_01723_),
    .A_N(_01649_));
 sg13g2_nor3_1 _07269_ (.A(_01629_),
    .B(_01643_),
    .C(_01724_),
    .Y(_01725_));
 sg13g2_buf_2 _07270_ (.A(_01725_),
    .X(_01726_));
 sg13g2_nor3_1 _07271_ (.A(_01379_),
    .B(_01212_),
    .C(_01209_),
    .Y(_01727_));
 sg13g2_buf_1 _07272_ (.A(_01727_),
    .X(_01728_));
 sg13g2_a21oi_1 _07273_ (.A1(net283),
    .A2(_01712_),
    .Y(_01729_),
    .B1(net282));
 sg13g2_nand2_1 _07274_ (.Y(_01730_),
    .A(_01272_),
    .B(_01300_));
 sg13g2_nand2b_1 _07275_ (.Y(_01731_),
    .B(_01303_),
    .A_N(_01298_));
 sg13g2_a21oi_1 _07276_ (.A1(_01730_),
    .A2(_01731_),
    .Y(_01732_),
    .B1(net308));
 sg13g2_nor3_1 _07277_ (.A(_01732_),
    .B(_01620_),
    .C(net273),
    .Y(_01733_));
 sg13g2_nand3_1 _07278_ (.B(_01729_),
    .C(_01733_),
    .A(_01726_),
    .Y(_01734_));
 sg13g2_nor4_1 _07279_ (.A(_01675_),
    .B(_01717_),
    .C(_01722_),
    .D(_01734_),
    .Y(_01735_));
 sg13g2_buf_2 _07280_ (.A(_01735_),
    .X(_01736_));
 sg13g2_mux2_1 _07281_ (.A0(net353),
    .A1(\dtop.player_inst.synth.alu.registers[4][1] ),
    .S(_01736_),
    .X(_01737_));
 sg13g2_buf_1 _07282_ (.A(_01737_),
    .X(_01738_));
 sg13g2_buf_8 _07283_ (.A(_01736_),
    .X(_01739_));
 sg13g2_mux2_1 _07284_ (.A0(net386),
    .A1(\dtop.player_inst.synth.alu.registers[4][2] ),
    .S(net101),
    .X(_01740_));
 sg13g2_nor2_1 _07285_ (.A(_05303_),
    .B(net101),
    .Y(_01741_));
 sg13g2_mux2_1 _07286_ (.A0(net352),
    .A1(\dtop.player_inst.synth.alu.registers[4][0] ),
    .S(_01736_),
    .X(_01742_));
 sg13g2_buf_1 _07287_ (.A(_01742_),
    .X(_01743_));
 sg13g2_mux4_1 _07288_ (.S0(net104),
    .A0(_01738_),
    .A1(_01740_),
    .A2(_01741_),
    .A3(_01743_),
    .S1(_01485_),
    .X(_01744_));
 sg13g2_nand2_1 _07289_ (.Y(_01745_),
    .A(net128),
    .B(_01744_));
 sg13g2_buf_1 _07290_ (.A(_01675_),
    .X(_01746_));
 sg13g2_nor3_2 _07291_ (.A(net200),
    .B(_01717_),
    .C(_01722_),
    .Y(_01747_));
 sg13g2_nand2_1 _07292_ (.Y(_01748_),
    .A(_01726_),
    .B(_01747_));
 sg13g2_buf_1 _07293_ (.A(_01748_),
    .X(_01749_));
 sg13g2_buf_1 _07294_ (.A(_01749_),
    .X(_01750_));
 sg13g2_mux2_1 _07295_ (.A0(_05324_),
    .A1(_00468_),
    .S(_01597_),
    .X(_01751_));
 sg13g2_mux2_1 _07296_ (.A0(_05281_),
    .A1(_05383_),
    .S(net102),
    .X(_01752_));
 sg13g2_buf_2 _07297_ (.A(\dtop.vtop.rs.saturated ),
    .X(_01753_));
 sg13g2_nor2_1 _07298_ (.A(_01753_),
    .B(net129),
    .Y(_01754_));
 sg13g2_a22oi_1 _07299_ (.Y(_01755_),
    .B1(_01752_),
    .B2(_01754_),
    .A2(_01751_),
    .A1(_01524_));
 sg13g2_or2_1 _07300_ (.X(_01756_),
    .B(net101),
    .A(net128));
 sg13g2_nor2_1 _07301_ (.A(_01755_),
    .B(_01756_),
    .Y(_01757_));
 sg13g2_nor2_1 _07302_ (.A(net86),
    .B(_01757_),
    .Y(_01758_));
 sg13g2_nand3_1 _07303_ (.B(_01719_),
    .C(_01720_),
    .A(_01718_),
    .Y(_01759_));
 sg13g2_nor4_1 _07304_ (.A(net200),
    .B(_01717_),
    .C(_01759_),
    .D(_01734_),
    .Y(_01760_));
 sg13g2_buf_1 _07305_ (.A(_01760_),
    .X(_01761_));
 sg13g2_nand2_1 _07306_ (.Y(_01762_),
    .A(\dtop.player_inst.synth.alu.registers[0][2] ),
    .B(net127));
 sg13g2_a21o_1 _07307_ (.A2(_01712_),
    .A1(_01462_),
    .B1(net282),
    .X(_01763_));
 sg13g2_nor4_1 _07308_ (.A(_01629_),
    .B(_01643_),
    .C(_01649_),
    .D(_01763_),
    .Y(_01764_));
 sg13g2_buf_2 _07309_ (.A(_01764_),
    .X(_01765_));
 sg13g2_a21oi_1 _07310_ (.A1(_01650_),
    .A2(_01674_),
    .Y(_01766_),
    .B1(_01765_));
 sg13g2_and4_1 _07311_ (.A(_01722_),
    .B(_01726_),
    .C(_01733_),
    .D(_01766_),
    .X(_01767_));
 sg13g2_buf_2 _07312_ (.A(_01767_),
    .X(_01768_));
 sg13g2_inv_2 _07313_ (.Y(_01769_),
    .A(_01753_));
 sg13g2_nor3_2 _07314_ (.A(net308),
    .B(_01298_),
    .C(_01429_),
    .Y(_01770_));
 sg13g2_and2_1 _07315_ (.A(_01769_),
    .B(_01770_),
    .X(_01771_));
 sg13g2_buf_1 _07316_ (.A(_01771_),
    .X(_01772_));
 sg13g2_nand2_1 _07317_ (.Y(_01773_),
    .A(_05322_),
    .B(_01772_));
 sg13g2_buf_1 _07318_ (.A(_01651_),
    .X(_01774_));
 sg13g2_a22oi_1 _07319_ (.Y(_01775_),
    .B1(net282),
    .B2(\dtop.player_inst.synth.alu.registers[2][2] ),
    .A2(net281),
    .A1(\dtop.player_inst.synth.alu.registers[1][2] ));
 sg13g2_a22oi_1 _07320_ (.Y(_01776_),
    .B1(net259),
    .B2(\dtop.player_inst.synth.alu.registers[5][2] ),
    .A2(_01657_),
    .A1(_00421_));
 sg13g2_nand3_1 _07321_ (.B(_01775_),
    .C(_01776_),
    .A(_01773_),
    .Y(_01777_));
 sg13g2_a221oi_1 _07322_ (.B2(\dtop.player_inst.synth.alu.registers[3][2] ),
    .C1(_01777_),
    .B1(_01768_),
    .A1(_01726_),
    .Y(_01778_),
    .A2(_01747_));
 sg13g2_and2_1 _07323_ (.A(_01762_),
    .B(_01778_),
    .X(_01779_));
 sg13g2_buf_1 _07324_ (.A(_01779_),
    .X(_01780_));
 sg13g2_a21oi_1 _07325_ (.A1(_01745_),
    .A2(_01758_),
    .Y(_01781_),
    .B1(_01780_));
 sg13g2_buf_1 _07326_ (.A(\dtop.player_inst.synth.alu.acc[3] ),
    .X(_01782_));
 sg13g2_inv_2 _07327_ (.Y(_01783_),
    .A(_01782_));
 sg13g2_nor2_1 _07328_ (.A(_01680_),
    .B(_01688_),
    .Y(_01784_));
 sg13g2_a22oi_1 _07329_ (.Y(_01785_),
    .B1(net283),
    .B2(net293),
    .A2(_01399_),
    .A1(_01251_));
 sg13g2_nand2b_1 _07330_ (.Y(_01786_),
    .B(_01785_),
    .A_N(_01732_));
 sg13g2_buf_1 _07331_ (.A(_01786_),
    .X(_01787_));
 sg13g2_nand2_1 _07332_ (.Y(_01788_),
    .A(_01251_),
    .B(_01417_));
 sg13g2_nor3_1 _07333_ (.A(net311),
    .B(net294),
    .C(_01237_),
    .Y(_01789_));
 sg13g2_o21ai_1 _07334_ (.B1(_00435_),
    .Y(_01790_),
    .A1(_01316_),
    .A2(_01789_));
 sg13g2_and2_1 _07335_ (.A(_01646_),
    .B(_01647_),
    .X(_01791_));
 sg13g2_o21ai_1 _07336_ (.B1(net284),
    .Y(_01792_),
    .A1(_01210_),
    .A2(_01335_));
 sg13g2_nand4_1 _07337_ (.B(_01790_),
    .C(_01791_),
    .A(_01788_),
    .Y(_01793_),
    .D(_01792_));
 sg13g2_nor4_1 _07338_ (.A(_01787_),
    .B(_01367_),
    .C(_01612_),
    .D(_01793_),
    .Y(_01794_));
 sg13g2_nand3_1 _07339_ (.B(_05204_),
    .C(_01285_),
    .A(_00420_),
    .Y(_01795_));
 sg13g2_o21ai_1 _07340_ (.B1(_01795_),
    .Y(_01796_),
    .A1(_05173_),
    .A2(_01275_));
 sg13g2_a221oi_1 _07341_ (.B2(net321),
    .C1(net298),
    .B1(_01796_),
    .A1(net295),
    .Y(_01797_),
    .A2(_01300_));
 sg13g2_o21ai_1 _07342_ (.B1(net286),
    .Y(_01798_),
    .A1(net342),
    .A2(_01379_));
 sg13g2_nand3b_1 _07343_ (.B(net299),
    .C(_01798_),
    .Y(_01799_),
    .A_N(_01797_));
 sg13g2_and3_1 _07344_ (.X(_01800_),
    .A(_01784_),
    .B(_01794_),
    .C(_01799_));
 sg13g2_buf_1 _07345_ (.A(_01800_),
    .X(_01801_));
 sg13g2_a21oi_1 _07346_ (.A1(_01273_),
    .A2(net293),
    .Y(_01802_),
    .B1(_01654_));
 sg13g2_nor2_1 _07347_ (.A(_01368_),
    .B(_01429_),
    .Y(_01803_));
 sg13g2_nor2_1 _07348_ (.A(_01275_),
    .B(_01368_),
    .Y(_01804_));
 sg13g2_a22oi_1 _07349_ (.Y(_01805_),
    .B1(_01804_),
    .B2(_01251_),
    .A2(_01803_),
    .A1(net284));
 sg13g2_nand2_1 _07350_ (.Y(_01806_),
    .A(_01802_),
    .B(_01805_));
 sg13g2_buf_1 _07351_ (.A(_05204_),
    .X(_01807_));
 sg13g2_nand2_1 _07352_ (.Y(_01808_),
    .A(net280),
    .B(net348));
 sg13g2_nor2_1 _07353_ (.A(net294),
    .B(_01253_),
    .Y(_01809_));
 sg13g2_a21oi_1 _07354_ (.A1(net291),
    .A2(_01205_),
    .Y(_01810_),
    .B1(_01809_));
 sg13g2_or2_1 _07355_ (.X(_01811_),
    .B(_01400_),
    .A(net285));
 sg13g2_a21oi_1 _07356_ (.A1(_01804_),
    .A2(_01811_),
    .Y(_01812_),
    .B1(_01625_));
 sg13g2_o21ai_1 _07357_ (.B1(_01812_),
    .Y(_01813_),
    .A1(_01808_),
    .A2(_01810_));
 sg13g2_or2_1 _07358_ (.X(_01814_),
    .B(_01412_),
    .A(_01402_));
 sg13g2_nand2_1 _07359_ (.Y(_01815_),
    .A(net346),
    .B(net292));
 sg13g2_nor3_1 _07360_ (.A(net299),
    .B(net326),
    .C(_01815_),
    .Y(_01816_));
 sg13g2_o21ai_1 _07361_ (.B1(net300),
    .Y(_01817_),
    .A1(_01422_),
    .A2(_01816_));
 sg13g2_a21oi_1 _07362_ (.A1(_01814_),
    .A2(_01817_),
    .Y(_01818_),
    .B1(net286));
 sg13g2_nor3_1 _07363_ (.A(_01806_),
    .B(_01813_),
    .C(_01818_),
    .Y(_01819_));
 sg13g2_and2_1 _07364_ (.A(_01801_),
    .B(_01819_),
    .X(_01820_));
 sg13g2_buf_1 _07365_ (.A(_01820_),
    .X(_01821_));
 sg13g2_nand2_1 _07366_ (.Y(_01822_),
    .A(net280),
    .B(net295));
 sg13g2_o21ai_1 _07367_ (.B1(_01822_),
    .Y(_01823_),
    .A1(net280),
    .A2(_01236_));
 sg13g2_nor4_1 _07368_ (.A(net300),
    .B(net326),
    .C(net311),
    .D(net294),
    .Y(_01824_));
 sg13g2_a22oi_1 _07369_ (.Y(_01825_),
    .B1(_01824_),
    .B2(net354),
    .A2(_01339_),
    .A1(_01823_));
 sg13g2_a22oi_1 _07370_ (.Y(_01826_),
    .B1(_01630_),
    .B2(net284),
    .A2(_01316_),
    .A1(_00461_));
 sg13g2_o21ai_1 _07371_ (.B1(_01826_),
    .Y(_01827_),
    .A1(_00461_),
    .A2(_01825_));
 sg13g2_nor2_1 _07372_ (.A(_01329_),
    .B(_01331_),
    .Y(_01828_));
 sg13g2_nand2_1 _07373_ (.Y(_01829_),
    .A(_00438_),
    .B(net314));
 sg13g2_nand2_1 _07374_ (.Y(_01830_),
    .A(net312),
    .B(_01360_));
 sg13g2_a21oi_1 _07375_ (.A1(_01829_),
    .A2(_01830_),
    .Y(_01831_),
    .B1(_01294_));
 sg13g2_nor4_1 _07376_ (.A(_01416_),
    .B(_01387_),
    .C(_01497_),
    .D(_01831_),
    .Y(_01832_));
 sg13g2_nand3_1 _07377_ (.B(_01633_),
    .C(_01832_),
    .A(_01828_),
    .Y(_01833_));
 sg13g2_nor2_1 _07378_ (.A(_01827_),
    .B(_01833_),
    .Y(_01834_));
 sg13g2_nand2_1 _07379_ (.Y(_01835_),
    .A(_01821_),
    .B(_01834_));
 sg13g2_buf_1 _07380_ (.A(_01835_),
    .X(_01836_));
 sg13g2_buf_1 _07381_ (.A(\dtop.player_inst.synth.alu.acc[8] ),
    .X(_01837_));
 sg13g2_buf_1 _07382_ (.A(_01787_),
    .X(_01838_));
 sg13g2_or2_1 _07383_ (.X(_01839_),
    .B(_01818_),
    .A(_01813_));
 sg13g2_buf_1 _07384_ (.A(_01839_),
    .X(_01840_));
 sg13g2_or2_1 _07385_ (.X(_01841_),
    .B(_01840_),
    .A(net249));
 sg13g2_nand3_1 _07386_ (.B(_01794_),
    .C(_01799_),
    .A(_01784_),
    .Y(_01842_));
 sg13g2_nor3_1 _07387_ (.A(_01787_),
    .B(_01813_),
    .C(_01818_),
    .Y(_01843_));
 sg13g2_and2_1 _07388_ (.A(_01842_),
    .B(_01843_),
    .X(_01844_));
 sg13g2_buf_1 _07389_ (.A(_01844_),
    .X(_01845_));
 sg13g2_buf_1 _07390_ (.A(\dtop.player_inst.synth.alu.acc[2] ),
    .X(_01846_));
 sg13g2_a22oi_1 _07391_ (.Y(_01847_),
    .B1(net167),
    .B2(net415),
    .A2(_01841_),
    .A1(_01837_));
 sg13g2_o21ai_1 _07392_ (.B1(_01847_),
    .Y(_01848_),
    .A1(_01783_),
    .A2(_01836_));
 sg13g2_buf_2 _07393_ (.A(\dtop.player_inst.synth.alu.acc[10] ),
    .X(_01849_));
 sg13g2_buf_1 _07394_ (.A(\dtop.player_inst.synth.alu.acc[1] ),
    .X(_01850_));
 sg13g2_xor2_1 _07395_ (.B(net414),
    .A(_01849_),
    .X(_01851_));
 sg13g2_and3_1 _07396_ (.X(_01852_),
    .A(_01801_),
    .B(_01819_),
    .C(_01834_));
 sg13g2_buf_1 _07397_ (.A(_01852_),
    .X(_01853_));
 sg13g2_nor2_1 _07398_ (.A(_01387_),
    .B(net249),
    .Y(_01854_));
 sg13g2_nor2b_1 _07399_ (.A(_01853_),
    .B_N(_01854_),
    .Y(_01855_));
 sg13g2_and3_1 _07400_ (.X(_01856_),
    .A(_01821_),
    .B(_01851_),
    .C(_01855_));
 sg13g2_buf_1 _07401_ (.A(_01633_),
    .X(_01857_));
 sg13g2_nand3_1 _07402_ (.B(_01821_),
    .C(_01855_),
    .A(net272),
    .Y(_01858_));
 sg13g2_o21ai_1 _07403_ (.B1(_01858_),
    .Y(_01859_),
    .A1(_01848_),
    .A2(_01856_));
 sg13g2_buf_1 _07404_ (.A(_01859_),
    .X(_01860_));
 sg13g2_nor2_1 _07405_ (.A(_01781_),
    .B(_01860_),
    .Y(_01861_));
 sg13g2_and2_1 _07406_ (.A(_01726_),
    .B(_01747_),
    .X(_01862_));
 sg13g2_buf_1 _07407_ (.A(_01862_),
    .X(_01863_));
 sg13g2_mux2_1 _07408_ (.A0(_05324_),
    .A1(_05304_),
    .S(_01516_),
    .X(_01864_));
 sg13g2_nor2_1 _07409_ (.A(net129),
    .B(_01736_),
    .Y(_01865_));
 sg13g2_nand3_1 _07410_ (.B(_01864_),
    .C(_01865_),
    .A(_01621_),
    .Y(_01866_));
 sg13g2_a21o_1 _07411_ (.A2(_01617_),
    .A1(_01611_),
    .B1(_01620_),
    .X(_01867_));
 sg13g2_buf_1 _07412_ (.A(_01867_),
    .X(_01868_));
 sg13g2_nor3_1 _07413_ (.A(_01484_),
    .B(_01598_),
    .C(_01868_),
    .Y(_01869_));
 sg13g2_buf_1 _07414_ (.A(_01868_),
    .X(_01870_));
 sg13g2_nor3_1 _07415_ (.A(net105),
    .B(_01516_),
    .C(net99),
    .Y(_01871_));
 sg13g2_a22oi_1 _07416_ (.Y(_01872_),
    .B1(_01871_),
    .B2(_01743_),
    .A2(_01869_),
    .A1(_01738_));
 sg13g2_nand2_1 _07417_ (.Y(_01873_),
    .A(_01521_),
    .B(_01611_));
 sg13g2_nand2_1 _07418_ (.Y(_01874_),
    .A(_01482_),
    .B(_01522_));
 sg13g2_a221oi_1 _07419_ (.B2(_01493_),
    .C1(_01514_),
    .B1(_01482_),
    .A1(net389),
    .Y(_01875_),
    .A2(_01769_));
 sg13g2_a221oi_1 _07420_ (.B2(_00467_),
    .C1(_01875_),
    .B1(_01516_),
    .A1(_01873_),
    .Y(_01876_),
    .A2(_01874_));
 sg13g2_nor4_1 _07421_ (.A(net385),
    .B(_01753_),
    .C(net129),
    .D(_01597_),
    .Y(_01877_));
 sg13g2_nor2_1 _07422_ (.A(_01621_),
    .B(_01739_),
    .Y(_01878_));
 sg13g2_o21ai_1 _07423_ (.B1(_01878_),
    .Y(_01879_),
    .A1(_01876_),
    .A2(_01877_));
 sg13g2_nand4_1 _07424_ (.B(_01866_),
    .C(_01872_),
    .A(_01863_),
    .Y(_01880_),
    .D(_01879_));
 sg13g2_buf_2 _07425_ (.A(_01880_),
    .X(_01881_));
 sg13g2_nand2_1 _07426_ (.Y(_01882_),
    .A(\dtop.player_inst.synth.alu.registers[3][1] ),
    .B(_01768_));
 sg13g2_nand2_1 _07427_ (.Y(_01883_),
    .A(net423),
    .B(_01772_));
 sg13g2_a22oi_1 _07428_ (.Y(_01884_),
    .B1(net282),
    .B2(\dtop.player_inst.synth.alu.registers[2][1] ),
    .A2(_01651_),
    .A1(\dtop.player_inst.synth.alu.registers[1][1] ));
 sg13g2_buf_2 _07429_ (.A(\dtop.player_inst.synth.alu.acc[0] ),
    .X(_01885_));
 sg13g2_inv_2 _07430_ (.Y(_01886_),
    .A(_01885_));
 sg13g2_nand4_1 _07431_ (.B(\dtop.player_inst.synth.alu.carry ),
    .C(\dtop.player_inst.synth.alu.oct_en ),
    .A(_01886_),
    .Y(_01887_),
    .D(_01649_));
 sg13g2_nand3_1 _07432_ (.B(_01884_),
    .C(_01887_),
    .A(_01883_),
    .Y(_01888_));
 sg13g2_a221oi_1 _07433_ (.B2(\dtop.player_inst.synth.alu.registers[5][1] ),
    .C1(_01888_),
    .B1(net259),
    .A1(_00516_),
    .Y(_01889_),
    .A2(net273));
 sg13g2_nand2_1 _07434_ (.Y(_01890_),
    .A(\dtop.player_inst.synth.alu.registers[0][1] ),
    .B(net127));
 sg13g2_nand4_1 _07435_ (.B(_01882_),
    .C(_01889_),
    .A(net100),
    .Y(_01891_),
    .D(_01890_));
 sg13g2_buf_2 _07436_ (.A(_01891_),
    .X(_01892_));
 sg13g2_and2_1 _07437_ (.A(_01881_),
    .B(_01892_),
    .X(_01893_));
 sg13g2_nand3_1 _07438_ (.B(_01842_),
    .C(_01843_),
    .A(net414),
    .Y(_01894_));
 sg13g2_buf_1 _07439_ (.A(\dtop.player_inst.synth.alu.acc[9] ),
    .X(_01895_));
 sg13g2_buf_2 _07440_ (.A(\dtop.player_inst.synth.alu.acc[7] ),
    .X(_01896_));
 sg13g2_xnor2_1 _07441_ (.Y(_01897_),
    .A(_01849_),
    .B(_01885_));
 sg13g2_nor2_1 _07442_ (.A(_01633_),
    .B(_01897_),
    .Y(_01898_));
 sg13g2_a221oi_1 _07443_ (.B2(_01896_),
    .C1(_01898_),
    .B1(_01840_),
    .A1(net413),
    .Y(_01899_),
    .A2(_01787_));
 sg13g2_nand4_1 _07444_ (.B(_01801_),
    .C(_01819_),
    .A(net415),
    .Y(_01900_),
    .D(_01834_));
 sg13g2_and3_1 _07445_ (.X(_01901_),
    .A(_01894_),
    .B(_01899_),
    .C(_01900_));
 sg13g2_buf_1 _07446_ (.A(_01901_),
    .X(_01902_));
 sg13g2_nor3_1 _07447_ (.A(_01609_),
    .B(_01893_),
    .C(_01902_),
    .Y(_01903_));
 sg13g2_a21o_1 _07448_ (.A2(_01861_),
    .A1(_01609_),
    .B1(_01903_),
    .X(_01904_));
 sg13g2_nand2_1 _07449_ (.Y(_01905_),
    .A(\dtop.player_inst.synth.alu.registers[5][0] ),
    .B(net259));
 sg13g2_nand2_1 _07450_ (.Y(_01906_),
    .A(net421),
    .B(_01772_));
 sg13g2_a22oi_1 _07451_ (.Y(_01907_),
    .B1(net282),
    .B2(\dtop.player_inst.synth.alu.registers[2][0] ),
    .A2(net281),
    .A1(\dtop.player_inst.synth.alu.registers[1][0] ));
 sg13g2_nand2_1 _07452_ (.Y(_01908_),
    .A(_01886_),
    .B(\dtop.player_inst.synth.alu.carry ));
 sg13g2_nand3_1 _07453_ (.B(_01649_),
    .C(_01908_),
    .A(\dtop.player_inst.synth.alu.oct_en ),
    .Y(_01909_));
 sg13g2_nand4_1 _07454_ (.B(_01906_),
    .C(_01907_),
    .A(_01905_),
    .Y(_01910_),
    .D(_01909_));
 sg13g2_a221oi_1 _07455_ (.B2(\dtop.player_inst.synth.alu.registers[3][0] ),
    .C1(_01910_),
    .B1(_01768_),
    .A1(_05182_),
    .Y(_01911_),
    .A2(net273));
 sg13g2_nand2_1 _07456_ (.Y(_01912_),
    .A(\dtop.player_inst.synth.alu.registers[0][0] ),
    .B(net127));
 sg13g2_nand3_1 _07457_ (.B(_01911_),
    .C(_01912_),
    .A(net100),
    .Y(_01913_));
 sg13g2_buf_2 _07458_ (.A(_01913_),
    .X(_01914_));
 sg13g2_nor2_1 _07459_ (.A(_01621_),
    .B(net100),
    .Y(_01915_));
 sg13g2_nor2_1 _07460_ (.A(net385),
    .B(_01516_),
    .Y(_01916_));
 sg13g2_and2_1 _07461_ (.A(_05280_),
    .B(_01493_),
    .X(_01917_));
 sg13g2_mux2_1 _07462_ (.A0(net375),
    .A1(_01917_),
    .S(_01522_),
    .X(_01918_));
 sg13g2_and2_1 _07463_ (.A(_05280_),
    .B(_01512_),
    .X(_01919_));
 sg13g2_mux2_1 _07464_ (.A0(_00779_),
    .A1(_01919_),
    .S(_01521_),
    .X(_01920_));
 sg13g2_mux2_1 _07465_ (.A0(_01918_),
    .A1(_01920_),
    .S(_01611_),
    .X(_01921_));
 sg13g2_nor2_1 _07466_ (.A(_01753_),
    .B(_01739_),
    .Y(_01922_));
 sg13g2_o21ai_1 _07467_ (.B1(_01922_),
    .Y(_01923_),
    .A1(_01916_),
    .A2(_01921_));
 sg13g2_nor2_1 _07468_ (.A(_01484_),
    .B(_01597_),
    .Y(_01924_));
 sg13g2_nor4_1 _07469_ (.A(_05303_),
    .B(_01484_),
    .C(_01516_),
    .D(_01736_),
    .Y(_01925_));
 sg13g2_a221oi_1 _07470_ (.B2(_01743_),
    .C1(_01925_),
    .B1(_01924_),
    .A1(_01751_),
    .Y(_01926_),
    .A2(_01865_));
 sg13g2_nor2_1 _07471_ (.A(net99),
    .B(net100),
    .Y(_01927_));
 sg13g2_a22oi_1 _07472_ (.Y(_01928_),
    .B1(_01926_),
    .B2(_01927_),
    .A2(_01923_),
    .A1(_01915_));
 sg13g2_buf_1 _07473_ (.A(_01928_),
    .X(_01929_));
 sg13g2_nand2_1 _07474_ (.Y(_01930_),
    .A(_01914_),
    .B(_01929_));
 sg13g2_nand2_1 _07475_ (.Y(_01931_),
    .A(net414),
    .B(_01853_));
 sg13g2_a22oi_1 _07476_ (.Y(_01932_),
    .B1(_01845_),
    .B2(_01885_),
    .A2(_01838_),
    .A1(_01849_));
 sg13g2_buf_1 _07477_ (.A(\dtop.player_inst.synth.alu.acc[6] ),
    .X(_01933_));
 sg13g2_a22oi_1 _07478_ (.Y(_01934_),
    .B1(_01840_),
    .B2(net412),
    .A2(_01801_),
    .A1(_01806_));
 sg13g2_nand3_1 _07479_ (.B(_01932_),
    .C(_01934_),
    .A(_01931_),
    .Y(_01935_));
 sg13g2_buf_1 _07480_ (.A(_01935_),
    .X(_01936_));
 sg13g2_nand2_1 _07481_ (.Y(_01937_),
    .A(_01930_),
    .B(_01936_));
 sg13g2_nand2_1 _07482_ (.Y(_01938_),
    .A(_01609_),
    .B(_01937_));
 sg13g2_nand2b_1 _07483_ (.Y(_01939_),
    .B(net103),
    .A_N(_01518_));
 sg13g2_nor2_1 _07484_ (.A(_05334_),
    .B(_01485_),
    .Y(_01940_));
 sg13g2_o21ai_1 _07485_ (.B1(net102),
    .Y(_01941_),
    .A1(_01561_),
    .A2(_01940_));
 sg13g2_nor2b_1 _07486_ (.A(\dtop.ext_control[0] ),
    .B_N(\dtop.ext_control[2] ),
    .Y(_01942_));
 sg13g2_o21ai_1 _07487_ (.B1(_01578_),
    .Y(_01943_),
    .A1(_01589_),
    .A2(_01942_));
 sg13g2_nand3_1 _07488_ (.B(_01517_),
    .C(_01943_),
    .A(net105),
    .Y(_01944_));
 sg13g2_nand3_1 _07489_ (.B(_01941_),
    .C(_01944_),
    .A(_01607_),
    .Y(_01945_));
 sg13g2_o21ai_1 _07490_ (.B1(_01945_),
    .Y(_01946_),
    .A1(_01198_),
    .A2(_01939_));
 sg13g2_mux2_1 _07491_ (.A0(_01904_),
    .A1(_01938_),
    .S(_01946_),
    .X(_01947_));
 sg13g2_and2_1 _07492_ (.A(_00779_),
    .B(_01772_),
    .X(_01948_));
 sg13g2_a221oi_1 _07493_ (.B2(\dtop.player_inst.synth.alu.registers[2][4] ),
    .C1(_01948_),
    .B1(net282),
    .A1(\dtop.player_inst.synth.alu.registers[1][4] ),
    .Y(_01949_),
    .A2(net281));
 sg13g2_a22oi_1 _07494_ (.Y(_01950_),
    .B1(net259),
    .B2(\dtop.player_inst.synth.alu.registers[5][4] ),
    .A2(net273),
    .A1(_05346_));
 sg13g2_a22oi_1 _07495_ (.Y(_01951_),
    .B1(_01768_),
    .B2(\dtop.player_inst.synth.alu.registers[3][4] ),
    .A2(net127),
    .A1(\dtop.player_inst.synth.alu.registers[0][4] ));
 sg13g2_nand4_1 _07496_ (.B(_01949_),
    .C(_01950_),
    .A(_01749_),
    .Y(_01952_),
    .D(_01951_));
 sg13g2_nand2_1 _07497_ (.Y(_01953_),
    .A(_01535_),
    .B(_01537_));
 sg13g2_a21oi_1 _07498_ (.A1(_01528_),
    .A2(_01531_),
    .Y(_01954_),
    .B1(_01539_));
 sg13g2_and2_1 _07499_ (.A(_05166_),
    .B(_01551_),
    .X(_01955_));
 sg13g2_nand3_1 _07500_ (.B(_01553_),
    .C(_01555_),
    .A(_01535_),
    .Y(_01956_));
 sg13g2_o21ai_1 _07501_ (.B1(_01528_),
    .Y(_01957_),
    .A1(_01225_),
    .A2(_01547_));
 sg13g2_o21ai_1 _07502_ (.B1(_01957_),
    .Y(_01958_),
    .A1(_01955_),
    .A2(_01956_));
 sg13g2_buf_2 _07503_ (.A(_01958_),
    .X(_01959_));
 sg13g2_a221oi_1 _07504_ (.B2(_01557_),
    .C1(_01499_),
    .B1(_01552_),
    .A1(_01528_),
    .Y(_01960_),
    .A2(_01549_));
 sg13g2_a221oi_1 _07505_ (.B2(_01233_),
    .C1(_01960_),
    .B1(_01959_),
    .A1(_01953_),
    .Y(_01961_),
    .A2(_01954_));
 sg13g2_nor2_1 _07506_ (.A(_01228_),
    .B(_01959_),
    .Y(_01962_));
 sg13g2_a221oi_1 _07507_ (.B2(_01650_),
    .C1(_01606_),
    .B1(_01729_),
    .A1(_01693_),
    .Y(_01963_),
    .A2(_01715_));
 sg13g2_o21ai_1 _07508_ (.B1(_01963_),
    .Y(_01964_),
    .A1(_01961_),
    .A2(_01962_));
 sg13g2_buf_1 _07509_ (.A(_01765_),
    .X(_01965_));
 sg13g2_a21oi_1 _07510_ (.A1(_01201_),
    .A2(_01227_),
    .Y(_01966_),
    .B1(_01191_));
 sg13g2_or2_1 _07511_ (.X(_01967_),
    .B(_01966_),
    .A(_01491_));
 sg13g2_inv_1 _07512_ (.Y(_01968_),
    .A(_01967_));
 sg13g2_a21oi_1 _07513_ (.A1(net199),
    .A2(_01968_),
    .Y(_01969_),
    .B1(net200));
 sg13g2_and2_1 _07514_ (.A(_01650_),
    .B(_01674_),
    .X(_01970_));
 sg13g2_buf_1 _07515_ (.A(_01970_),
    .X(_01971_));
 sg13g2_nor2_1 _07516_ (.A(_01765_),
    .B(_01967_),
    .Y(_01972_));
 sg13g2_nor2_1 _07517_ (.A(_01971_),
    .B(_01972_),
    .Y(_01973_));
 sg13g2_nor2b_1 _07518_ (.A(_05367_),
    .B_N(_05214_),
    .Y(_01974_));
 sg13g2_mux2_1 _07519_ (.A0(_05368_),
    .A1(_01974_),
    .S(_01233_),
    .X(_01975_));
 sg13g2_nand2_1 _07520_ (.Y(_01976_),
    .A(net391),
    .B(_01975_));
 sg13g2_nand2_1 _07521_ (.Y(_01977_),
    .A(net388),
    .B(_01569_));
 sg13g2_nand2_1 _07522_ (.Y(_01978_),
    .A(net274),
    .B(_01977_));
 sg13g2_nand2_1 _07523_ (.Y(_01979_),
    .A(net392),
    .B(net420));
 sg13g2_o21ai_1 _07524_ (.B1(_00471_),
    .Y(_01980_),
    .A1(_01221_),
    .A2(_01223_));
 sg13g2_o21ai_1 _07525_ (.B1(_01980_),
    .Y(_01981_),
    .A1(_01507_),
    .A2(_01979_));
 sg13g2_a22oi_1 _07526_ (.Y(_01982_),
    .B1(_01981_),
    .B2(_05221_),
    .A2(_01978_),
    .A1(net350));
 sg13g2_o21ai_1 _07527_ (.B1(_01980_),
    .Y(_01983_),
    .A1(_01228_),
    .A2(_01569_));
 sg13g2_a21oi_1 _07528_ (.A1(net388),
    .A2(_00426_),
    .Y(_01984_),
    .B1(_05154_));
 sg13g2_o21ai_1 _07529_ (.B1(net339),
    .Y(_01985_),
    .A1(net351),
    .A2(_01569_));
 sg13g2_nand2_1 _07530_ (.Y(_01986_),
    .A(net353),
    .B(_01985_));
 sg13g2_nand2_1 _07531_ (.Y(_01987_),
    .A(_01984_),
    .B(_01986_));
 sg13g2_a221oi_1 _07532_ (.B2(net352),
    .C1(_01987_),
    .B1(_01983_),
    .A1(_01976_),
    .Y(_01988_),
    .A2(_01982_));
 sg13g2_nor2_1 _07533_ (.A(net339),
    .B(_00426_),
    .Y(_01989_));
 sg13g2_nor3_1 _07534_ (.A(net392),
    .B(net274),
    .C(_01989_),
    .Y(_01990_));
 sg13g2_nor3_1 _07535_ (.A(net350),
    .B(net388),
    .C(_01507_),
    .Y(_01991_));
 sg13g2_o21ai_1 _07536_ (.B1(_05154_),
    .Y(_01992_),
    .A1(_01990_),
    .A2(_01991_));
 sg13g2_nand2_1 _07537_ (.Y(_01993_),
    .A(_00401_),
    .B(_01992_));
 sg13g2_and2_1 _07538_ (.A(_05332_),
    .B(_01567_),
    .X(_01994_));
 sg13g2_mux2_1 _07539_ (.A0(_01565_),
    .A1(_01994_),
    .S(net274),
    .X(_01995_));
 sg13g2_mux2_1 _07540_ (.A0(_01567_),
    .A1(_01574_),
    .S(net274),
    .X(_01996_));
 sg13g2_a221oi_1 _07541_ (.B2(_01565_),
    .C1(_00401_),
    .B1(_01996_),
    .A1(net350),
    .Y(_01997_),
    .A2(_01995_));
 sg13g2_nor2b_1 _07542_ (.A(_01997_),
    .B_N(_01765_),
    .Y(_01998_));
 sg13g2_o21ai_1 _07543_ (.B1(_01998_),
    .Y(_01999_),
    .A1(_01988_),
    .A2(_01993_));
 sg13g2_a22oi_1 _07544_ (.Y(_02000_),
    .B1(_01973_),
    .B2(_01999_),
    .A2(_01969_),
    .A1(_01964_));
 sg13g2_buf_1 _07545_ (.A(_02000_),
    .X(_02001_));
 sg13g2_nor2_1 _07546_ (.A(net296),
    .B(_02001_),
    .Y(_02002_));
 sg13g2_a221oi_1 _07547_ (.B2(_01999_),
    .C1(_01546_),
    .B1(_01973_),
    .A1(_01964_),
    .Y(_02003_),
    .A2(_01969_));
 sg13g2_buf_1 _07548_ (.A(_02003_),
    .X(_02004_));
 sg13g2_nor2_1 _07549_ (.A(_02002_),
    .B(_02004_),
    .Y(_02005_));
 sg13g2_or2_1 _07550_ (.X(_02006_),
    .B(_01765_),
    .A(_01606_));
 sg13g2_nor3_2 _07551_ (.A(_01675_),
    .B(_01717_),
    .C(_02006_),
    .Y(_02007_));
 sg13g2_a21oi_1 _07552_ (.A1(net288),
    .A2(_01193_),
    .Y(_02008_),
    .B1(net317));
 sg13g2_nand2_1 _07553_ (.Y(_02009_),
    .A(_00426_),
    .B(_02008_));
 sg13g2_a21oi_1 _07554_ (.A1(_01959_),
    .A2(_02009_),
    .Y(_02010_),
    .B1(_01543_));
 sg13g2_a21o_1 _07555_ (.A2(_01559_),
    .A1(_01503_),
    .B1(_02010_),
    .X(_02011_));
 sg13g2_a21oi_1 _07556_ (.A1(net372),
    .A2(_05385_),
    .Y(_02012_),
    .B1(_01509_));
 sg13g2_nor2_1 _07557_ (.A(_02012_),
    .B(_01491_),
    .Y(_02013_));
 sg13g2_a21oi_1 _07558_ (.A1(net386),
    .A2(net307),
    .Y(_02014_),
    .B1(_01529_));
 sg13g2_nand3_1 _07559_ (.B(net307),
    .C(_01569_),
    .A(net339),
    .Y(_02015_));
 sg13g2_o21ai_1 _07560_ (.B1(_02015_),
    .Y(_02016_),
    .A1(net392),
    .A2(_02014_));
 sg13g2_nor4_1 _07561_ (.A(_00471_),
    .B(_05331_),
    .C(net427),
    .D(_05154_),
    .Y(_02017_));
 sg13g2_nor3_1 _07562_ (.A(net392),
    .B(net386),
    .C(net307),
    .Y(_02018_));
 sg13g2_o21ai_1 _07563_ (.B1(net391),
    .Y(_02019_),
    .A1(_02017_),
    .A2(_02018_));
 sg13g2_nor2b_1 _07564_ (.A(_02016_),
    .B_N(_02019_),
    .Y(_02020_));
 sg13g2_nand2_1 _07565_ (.Y(_02021_),
    .A(_00401_),
    .B(_01499_));
 sg13g2_o21ai_1 _07566_ (.B1(_01576_),
    .Y(_02022_),
    .A1(_02020_),
    .A2(_02021_));
 sg13g2_mux2_1 _07567_ (.A0(_02013_),
    .A1(_02022_),
    .S(_01765_),
    .X(_02023_));
 sg13g2_and2_1 _07568_ (.A(_01765_),
    .B(_02013_),
    .X(_02024_));
 sg13g2_mux2_1 _07569_ (.A0(_02023_),
    .A1(_02024_),
    .S(_01971_),
    .X(_02025_));
 sg13g2_a21o_1 _07570_ (.A2(_02011_),
    .A1(_02007_),
    .B1(_02025_),
    .X(_02026_));
 sg13g2_buf_1 _07571_ (.A(_02026_),
    .X(_02027_));
 sg13g2_and2_1 _07572_ (.A(_00426_),
    .B(_02008_),
    .X(_02028_));
 sg13g2_a21oi_1 _07573_ (.A1(_01959_),
    .A2(_02028_),
    .Y(_02029_),
    .B1(_01543_));
 sg13g2_xnor2_1 _07574_ (.Y(_02030_),
    .A(net372),
    .B(_01559_));
 sg13g2_and2_1 _07575_ (.A(_01233_),
    .B(_01543_),
    .X(_02031_));
 sg13g2_a22oi_1 _07576_ (.Y(_02032_),
    .B1(_02030_),
    .B2(_02031_),
    .A2(_02029_),
    .A1(_01507_));
 sg13g2_nand2b_1 _07577_ (.Y(_02033_),
    .B(_02012_),
    .A_N(_02032_));
 sg13g2_nor2_1 _07578_ (.A(_01191_),
    .B(_01559_),
    .Y(_02034_));
 sg13g2_nor2_1 _07579_ (.A(_01546_),
    .B(_01959_),
    .Y(_02035_));
 sg13g2_nor3_1 _07580_ (.A(_01543_),
    .B(_02034_),
    .C(_02035_),
    .Y(_02036_));
 sg13g2_nor4_2 _07581_ (.A(net200),
    .B(net199),
    .C(_02006_),
    .Y(_02037_),
    .D(_02036_));
 sg13g2_nor3_1 _07582_ (.A(_01503_),
    .B(_01491_),
    .C(_01615_),
    .Y(_02038_));
 sg13g2_nand3_1 _07583_ (.B(net199),
    .C(_02038_),
    .A(_01971_),
    .Y(_02039_));
 sg13g2_nand2_1 _07584_ (.Y(_02040_),
    .A(_01766_),
    .B(_02038_));
 sg13g2_nand2_2 _07585_ (.Y(_02041_),
    .A(net305),
    .B(_01501_));
 sg13g2_nand2_1 _07586_ (.Y(_02042_),
    .A(_02041_),
    .B(_01994_));
 sg13g2_o21ai_1 _07587_ (.B1(_02042_),
    .Y(_02043_),
    .A1(net388),
    .A2(_01510_));
 sg13g2_a22oi_1 _07588_ (.Y(_02044_),
    .B1(_01574_),
    .B2(_02041_),
    .A2(_01567_),
    .A1(_01499_));
 sg13g2_nor2_1 _07589_ (.A(net388),
    .B(_02044_),
    .Y(_02045_));
 sg13g2_a21oi_1 _07590_ (.A1(_00407_),
    .A2(_02043_),
    .Y(_02046_),
    .B1(_02045_));
 sg13g2_nand2_1 _07591_ (.Y(_02047_),
    .A(_01563_),
    .B(_02046_));
 sg13g2_a21oi_1 _07592_ (.A1(net305),
    .A2(_01501_),
    .Y(_02048_),
    .B1(_01979_));
 sg13g2_a21oi_1 _07593_ (.A1(net351),
    .A2(net305),
    .Y(_02049_),
    .B1(_05368_));
 sg13g2_o21ai_1 _07594_ (.B1(_05221_),
    .Y(_02050_),
    .A1(_02048_),
    .A2(_02049_));
 sg13g2_nand3_1 _07595_ (.B(net305),
    .C(_01501_),
    .A(net392),
    .Y(_02051_));
 sg13g2_and2_1 _07596_ (.A(_05220_),
    .B(_01974_),
    .X(_02052_));
 sg13g2_a22oi_1 _07597_ (.Y(_02053_),
    .B1(_02052_),
    .B2(_02041_),
    .A2(_02051_),
    .A1(_01499_));
 sg13g2_a21oi_1 _07598_ (.A1(_02050_),
    .A2(_02053_),
    .Y(_02054_),
    .B1(_05332_));
 sg13g2_nand2_1 _07599_ (.Y(_02055_),
    .A(net386),
    .B(_01499_));
 sg13g2_nand2b_1 _07600_ (.Y(_02056_),
    .B(_02041_),
    .A_N(_01977_));
 sg13g2_a21oi_1 _07601_ (.A1(_02055_),
    .A2(_02056_),
    .Y(_02057_),
    .B1(_05215_));
 sg13g2_o21ai_1 _07602_ (.B1(net307),
    .Y(_02058_),
    .A1(_02054_),
    .A2(_02057_));
 sg13g2_o21ai_1 _07603_ (.B1(net388),
    .Y(_02059_),
    .A1(net392),
    .A2(_00472_));
 sg13g2_nand2_1 _07604_ (.Y(_02060_),
    .A(net350),
    .B(_05135_));
 sg13g2_nand3_1 _07605_ (.B(_02059_),
    .C(_02060_),
    .A(_05154_),
    .Y(_02061_));
 sg13g2_nand3_1 _07606_ (.B(_02058_),
    .C(_02061_),
    .A(_00401_),
    .Y(_02062_));
 sg13g2_nand4_1 _07607_ (.B(net199),
    .C(_02047_),
    .A(net200),
    .Y(_02063_),
    .D(_02062_));
 sg13g2_and3_1 _07608_ (.X(_02064_),
    .A(_02039_),
    .B(_02040_),
    .C(_02063_));
 sg13g2_a21oi_1 _07609_ (.A1(_01543_),
    .A2(_01959_),
    .Y(_02065_),
    .B1(_02012_));
 sg13g2_nor2_1 _07610_ (.A(_01233_),
    .B(_02028_),
    .Y(_02066_));
 sg13g2_nor3_1 _07611_ (.A(_01233_),
    .B(_01499_),
    .C(_02008_),
    .Y(_02067_));
 sg13g2_a221oi_1 _07612_ (.B2(_01557_),
    .C1(_02067_),
    .B1(_01552_),
    .A1(_01528_),
    .Y(_02068_),
    .A2(_01549_));
 sg13g2_a22oi_1 _07613_ (.Y(_02069_),
    .B1(_02068_),
    .B2(_01543_),
    .A2(_02066_),
    .A1(_01959_));
 sg13g2_or3_1 _07614_ (.A(net351),
    .B(_02065_),
    .C(_02069_),
    .X(_02070_));
 sg13g2_a22oi_1 _07615_ (.Y(_02071_),
    .B1(_02068_),
    .B2(_01507_),
    .A2(_02009_),
    .A1(_01959_));
 sg13g2_or3_1 _07616_ (.A(_01191_),
    .B(_01543_),
    .C(_02071_),
    .X(_02072_));
 sg13g2_nand3_1 _07617_ (.B(_02070_),
    .C(_02072_),
    .A(_02007_),
    .Y(_02073_));
 sg13g2_a221oi_1 _07618_ (.B2(net351),
    .C1(_01491_),
    .B1(_01615_),
    .A1(_01191_),
    .Y(_02074_),
    .A2(_01546_));
 sg13g2_inv_1 _07619_ (.Y(_02075_),
    .A(_02074_));
 sg13g2_xnor2_1 _07620_ (.Y(_02076_),
    .A(net200),
    .B(net199));
 sg13g2_inv_1 _07621_ (.Y(_02077_),
    .A(_01569_));
 sg13g2_nor2_1 _07622_ (.A(_05132_),
    .B(net372),
    .Y(_02078_));
 sg13g2_a221oi_1 _07623_ (.B2(_02078_),
    .C1(_01545_),
    .B1(_01231_),
    .A1(net328),
    .Y(_02079_),
    .A2(_01221_));
 sg13g2_buf_1 _07624_ (.A(_02079_),
    .X(_02080_));
 sg13g2_o21ai_1 _07625_ (.B1(net339),
    .Y(_02081_),
    .A1(_02077_),
    .A2(_02080_));
 sg13g2_o21ai_1 _07626_ (.B1(_01984_),
    .Y(_02082_),
    .A1(_01571_),
    .A2(_02080_));
 sg13g2_a221oi_1 _07627_ (.B2(net353),
    .C1(_02082_),
    .B1(_02081_),
    .A1(_00489_),
    .Y(_02083_),
    .A2(_01544_));
 sg13g2_nor2_1 _07628_ (.A(_05215_),
    .B(_02080_),
    .Y(_02084_));
 sg13g2_nand2_1 _07629_ (.Y(_02085_),
    .A(_05154_),
    .B(_02059_));
 sg13g2_o21ai_1 _07630_ (.B1(_00401_),
    .Y(_02086_),
    .A1(_02084_),
    .A2(_02085_));
 sg13g2_o21ai_1 _07631_ (.B1(net339),
    .Y(_02087_),
    .A1(_01574_),
    .A2(_02080_));
 sg13g2_nand3_1 _07632_ (.B(_01584_),
    .C(_02087_),
    .A(_01563_),
    .Y(_02088_));
 sg13g2_o21ai_1 _07633_ (.B1(_02088_),
    .Y(_02089_),
    .A1(_02083_),
    .A2(_02086_));
 sg13g2_nand3b_1 _07634_ (.B(net200),
    .C(net199),
    .Y(_02090_),
    .A_N(_02089_));
 sg13g2_o21ai_1 _07635_ (.B1(_02090_),
    .Y(_02091_),
    .A1(_02075_),
    .A2(_02076_));
 sg13g2_a221oi_1 _07636_ (.B2(_02073_),
    .C1(_02091_),
    .B1(_02064_),
    .A1(_02033_),
    .Y(_02092_),
    .A2(_02037_));
 sg13g2_buf_2 _07637_ (.A(_02092_),
    .X(_02093_));
 sg13g2_nor2_1 _07638_ (.A(_02027_),
    .B(_02093_),
    .Y(_02094_));
 sg13g2_nand2b_1 _07639_ (.Y(_02095_),
    .B(_01746_),
    .A_N(_01732_));
 sg13g2_nor2_1 _07640_ (.A(_01746_),
    .B(_01717_),
    .Y(_02096_));
 sg13g2_o21ai_1 _07641_ (.B1(_02096_),
    .Y(_02097_),
    .A1(_01759_),
    .A2(_01726_));
 sg13g2_nand2_1 _07642_ (.Y(_02098_),
    .A(_01650_),
    .B(_01723_));
 sg13g2_nor3_1 _07643_ (.A(_01722_),
    .B(_02098_),
    .C(_01965_),
    .Y(_02099_));
 sg13g2_a21oi_1 _07644_ (.A1(_02095_),
    .A2(_02097_),
    .Y(_02100_),
    .B1(_02099_));
 sg13g2_buf_1 _07645_ (.A(_02100_),
    .X(_02101_));
 sg13g2_a21oi_1 _07646_ (.A1(_02005_),
    .A2(_02094_),
    .Y(_02102_),
    .B1(_02101_));
 sg13g2_mux2_1 _07647_ (.A0(net391),
    .A1(\dtop.player_inst.synth.alu.registers[4][3] ),
    .S(net101),
    .X(_02103_));
 sg13g2_mux2_1 _07648_ (.A0(_05387_),
    .A1(\dtop.player_inst.synth.alu.registers[4][4] ),
    .S(net101),
    .X(_02104_));
 sg13g2_mux4_1 _07649_ (.S0(net104),
    .A0(_01738_),
    .A1(_01740_),
    .A2(_02103_),
    .A3(_02104_),
    .S1(net129),
    .X(_02105_));
 sg13g2_nor2_1 _07650_ (.A(net99),
    .B(_02105_),
    .Y(_02106_));
 sg13g2_and2_1 _07651_ (.A(_01870_),
    .B(_01926_),
    .X(_02107_));
 sg13g2_o21ai_1 _07652_ (.B1(_01863_),
    .Y(_02108_),
    .A1(_02106_),
    .A2(_02107_));
 sg13g2_o21ai_1 _07653_ (.B1(_02108_),
    .Y(_02109_),
    .A1(_01952_),
    .A2(_02102_));
 sg13g2_buf_1 _07654_ (.A(_02109_),
    .X(_02110_));
 sg13g2_buf_2 _07655_ (.A(\dtop.player_inst.synth.alu.acc[5] ),
    .X(_02111_));
 sg13g2_inv_1 _07656_ (.Y(_02112_),
    .A(_02111_));
 sg13g2_buf_1 _07657_ (.A(\dtop.player_inst.synth.alu.acc[4] ),
    .X(_02113_));
 sg13g2_buf_1 _07658_ (.A(_01849_),
    .X(_02114_));
 sg13g2_xnor2_1 _07659_ (.Y(_02115_),
    .A(net371),
    .B(_01782_));
 sg13g2_nand2_1 _07660_ (.Y(_02116_),
    .A(_01933_),
    .B(net249));
 sg13g2_o21ai_1 _07661_ (.B1(_02116_),
    .Y(_02117_),
    .A1(net272),
    .A2(_02115_));
 sg13g2_a221oi_1 _07662_ (.B2(_02113_),
    .C1(_02117_),
    .B1(net167),
    .A1(_00060_),
    .Y(_02118_),
    .A2(_01840_));
 sg13g2_o21ai_1 _07663_ (.B1(_02118_),
    .Y(_02119_),
    .A1(_02112_),
    .A2(_01836_));
 sg13g2_buf_1 _07664_ (.A(_02119_),
    .X(_02120_));
 sg13g2_nand4_1 _07665_ (.B(_01609_),
    .C(_02110_),
    .A(_01946_),
    .Y(_02121_),
    .D(_02120_));
 sg13g2_inv_2 _07666_ (.Y(_02122_),
    .A(_02113_));
 sg13g2_xnor2_1 _07667_ (.Y(_02123_),
    .A(_01849_),
    .B(net415));
 sg13g2_nand2_1 _07668_ (.Y(_02124_),
    .A(_01896_),
    .B(net249));
 sg13g2_o21ai_1 _07669_ (.B1(_02124_),
    .Y(_02125_),
    .A1(net272),
    .A2(_02123_));
 sg13g2_a221oi_1 _07670_ (.B2(_01782_),
    .C1(_02125_),
    .B1(net167),
    .A1(net413),
    .Y(_02126_),
    .A2(_01840_));
 sg13g2_o21ai_1 _07671_ (.B1(_02126_),
    .Y(_02127_),
    .A1(_02122_),
    .A2(_01836_));
 sg13g2_buf_1 _07672_ (.A(_02127_),
    .X(_02128_));
 sg13g2_nand2_1 _07673_ (.Y(_02129_),
    .A(net199),
    .B(_02074_));
 sg13g2_nand2_1 _07674_ (.Y(_02130_),
    .A(_01693_),
    .B(_01715_));
 sg13g2_or3_1 _07675_ (.A(_02130_),
    .B(net199),
    .C(_02089_),
    .X(_02131_));
 sg13g2_nand3_1 _07676_ (.B(_02129_),
    .C(_02131_),
    .A(_01971_),
    .Y(_02132_));
 sg13g2_mux2_1 _07677_ (.A0(_02075_),
    .A1(_02089_),
    .S(_01965_),
    .X(_02133_));
 sg13g2_nand2_1 _07678_ (.Y(_02134_),
    .A(net200),
    .B(_02133_));
 sg13g2_a221oi_1 _07679_ (.B2(_02037_),
    .C1(_02027_),
    .B1(_02033_),
    .A1(_02132_),
    .Y(_02135_),
    .A2(_02134_));
 sg13g2_nand3_1 _07680_ (.B(_02040_),
    .C(_02063_),
    .A(_02039_),
    .Y(_02136_));
 sg13g2_buf_1 _07681_ (.A(_02136_),
    .X(_02137_));
 sg13g2_and3_1 _07682_ (.X(_02138_),
    .A(_02007_),
    .B(_02070_),
    .C(_02072_));
 sg13g2_buf_1 _07683_ (.A(_02138_),
    .X(_02139_));
 sg13g2_nor4_2 _07684_ (.A(net296),
    .B(_02001_),
    .C(_02137_),
    .Y(_02140_),
    .D(_02139_));
 sg13g2_nand2b_1 _07685_ (.Y(_02141_),
    .B(_02140_),
    .A_N(_02135_));
 sg13g2_nand2_1 _07686_ (.Y(_02142_),
    .A(_05376_),
    .B(_01772_));
 sg13g2_a22oi_1 _07687_ (.Y(_02143_),
    .B1(net282),
    .B2(\dtop.player_inst.synth.alu.registers[2][3] ),
    .A2(net281),
    .A1(\dtop.player_inst.synth.alu.registers[1][3] ));
 sg13g2_a22oi_1 _07688_ (.Y(_02144_),
    .B1(net259),
    .B2(\dtop.player_inst.synth.alu.registers[5][3] ),
    .A2(net273),
    .A1(_05298_));
 sg13g2_nand4_1 _07689_ (.B(_02142_),
    .C(_02143_),
    .A(net100),
    .Y(_02145_),
    .D(_02144_));
 sg13g2_a221oi_1 _07690_ (.B2(\dtop.player_inst.synth.alu.registers[3][3] ),
    .C1(_02145_),
    .B1(_01768_),
    .A1(\dtop.player_inst.synth.alu.registers[0][3] ),
    .Y(_02146_),
    .A2(_01761_));
 sg13g2_a21oi_1 _07691_ (.A1(_02007_),
    .A2(_02011_),
    .Y(_02147_),
    .B1(_02025_));
 sg13g2_buf_2 _07692_ (.A(_02147_),
    .X(_02148_));
 sg13g2_nand2_1 _07693_ (.Y(_02149_),
    .A(_02148_),
    .B(_02093_));
 sg13g2_o21ai_1 _07694_ (.B1(_02004_),
    .Y(_02150_),
    .A1(_02148_),
    .A2(_02093_));
 sg13g2_nand4_1 _07695_ (.B(_02146_),
    .C(_02149_),
    .A(_02141_),
    .Y(_02151_),
    .D(_02150_));
 sg13g2_mux4_1 _07696_ (.S0(net102),
    .A0(_01738_),
    .A1(_01743_),
    .A2(_02103_),
    .A3(_01740_),
    .S1(net129),
    .X(_02152_));
 sg13g2_buf_1 _07697_ (.A(net101),
    .X(_02153_));
 sg13g2_nand2_1 _07698_ (.Y(_02154_),
    .A(net389),
    .B(_01769_));
 sg13g2_mux4_1 _07699_ (.S0(_01516_),
    .A0(net425),
    .A1(_05303_),
    .A2(_02154_),
    .A3(_00467_),
    .S1(net105),
    .X(_02155_));
 sg13g2_nor3_1 _07700_ (.A(net128),
    .B(net85),
    .C(_02155_),
    .Y(_02156_));
 sg13g2_a21oi_1 _07701_ (.A1(net128),
    .A2(_02152_),
    .Y(_02157_),
    .B1(_02156_));
 sg13g2_a22oi_1 _07702_ (.Y(_02158_),
    .B1(_02157_),
    .B2(_01863_),
    .A2(_02101_),
    .A1(_02146_));
 sg13g2_nand2_1 _07703_ (.Y(_02159_),
    .A(_02151_),
    .B(_02158_));
 sg13g2_nand2_1 _07704_ (.Y(_02160_),
    .A(_02128_),
    .B(_02159_));
 sg13g2_a21o_1 _07705_ (.A2(_02160_),
    .A1(_01946_),
    .B1(_01609_),
    .X(_02161_));
 sg13g2_nand2_1 _07706_ (.Y(_02162_),
    .A(_02121_),
    .B(_02161_));
 sg13g2_and2_1 _07707_ (.A(_01578_),
    .B(_01590_),
    .X(_02163_));
 sg13g2_nand2_1 _07708_ (.Y(_02164_),
    .A(\dtop.ext_control[0] ),
    .B(_01600_));
 sg13g2_o21ai_1 _07709_ (.B1(_02164_),
    .Y(_02165_),
    .A1(_01586_),
    .A2(_02163_));
 sg13g2_nand2_1 _07710_ (.Y(_02166_),
    .A(_01517_),
    .B(_02165_));
 sg13g2_a21oi_1 _07711_ (.A1(_01602_),
    .A2(_01518_),
    .Y(_02167_),
    .B1(net105));
 sg13g2_a21oi_1 _07712_ (.A1(_01607_),
    .A2(_02166_),
    .Y(_02168_),
    .B1(_02167_));
 sg13g2_mux2_1 _07713_ (.A0(_01947_),
    .A1(_02162_),
    .S(_02168_),
    .X(_02169_));
 sg13g2_buf_1 _07714_ (.A(rst_n_reg),
    .X(_02170_));
 sg13g2_buf_1 _07715_ (.A(net411),
    .X(_02171_));
 sg13g2_nand3_1 _07716_ (.B(_01324_),
    .C(_01400_),
    .A(net310),
    .Y(_02172_));
 sg13g2_nand3_1 _07717_ (.B(net283),
    .C(_01384_),
    .A(net312),
    .Y(_02173_));
 sg13g2_nand2_1 _07718_ (.Y(_02174_),
    .A(net284),
    .B(_01213_));
 sg13g2_o21ai_1 _07719_ (.B1(_01249_),
    .Y(_02175_),
    .A1(_01251_),
    .A2(_01205_));
 sg13g2_a22oi_1 _07720_ (.Y(_02176_),
    .B1(net284),
    .B2(_01803_),
    .A2(_01457_),
    .A1(net285));
 sg13g2_a21oi_1 _07721_ (.A1(net300),
    .A2(net348),
    .Y(_02177_),
    .B1(_05163_));
 sg13g2_a21oi_1 _07722_ (.A1(_01670_),
    .A2(_02177_),
    .Y(_02178_),
    .B1(_01625_));
 sg13g2_and4_1 _07723_ (.A(_02175_),
    .B(_02176_),
    .C(_02178_),
    .D(_01447_),
    .X(_02179_));
 sg13g2_a22oi_1 _07724_ (.Y(_02180_),
    .B1(_01384_),
    .B2(net314),
    .A2(net312),
    .A1(net309));
 sg13g2_nor2_1 _07725_ (.A(_01815_),
    .B(_02180_),
    .Y(_02181_));
 sg13g2_nand2_1 _07726_ (.Y(_02182_),
    .A(_01330_),
    .B(_01618_));
 sg13g2_nor4_1 _07727_ (.A(_01266_),
    .B(_01416_),
    .C(_02181_),
    .D(_02182_),
    .Y(_02183_));
 sg13g2_nand2_1 _07728_ (.Y(_02184_),
    .A(net287),
    .B(_01809_));
 sg13g2_nand3_1 _07729_ (.B(net295),
    .C(_01702_),
    .A(net291),
    .Y(_02185_));
 sg13g2_nand2_1 _07730_ (.Y(_02186_),
    .A(_02184_),
    .B(_02185_));
 sg13g2_nor2_1 _07731_ (.A(_01707_),
    .B(_01494_),
    .Y(_02187_));
 sg13g2_a22oi_1 _07732_ (.Y(_02188_),
    .B1(_02187_),
    .B2(net348),
    .A2(_01474_),
    .A1(_01340_));
 sg13g2_a21oi_1 _07733_ (.A1(net287),
    .A2(net280),
    .Y(_02189_),
    .B1(net286));
 sg13g2_o21ai_1 _07734_ (.B1(_01285_),
    .Y(_02190_),
    .A1(_01702_),
    .A2(_02189_));
 sg13g2_o21ai_1 _07735_ (.B1(_02190_),
    .Y(_02191_),
    .A1(net291),
    .A2(_02188_));
 sg13g2_a22oi_1 _07736_ (.Y(_02192_),
    .B1(_02191_),
    .B2(net340),
    .A2(_02186_),
    .A1(_05202_));
 sg13g2_o21ai_1 _07737_ (.B1(_05143_),
    .Y(_02193_),
    .A1(net297),
    .A2(_01249_));
 sg13g2_mux2_1 _07738_ (.A0(_02193_),
    .A1(_01352_),
    .S(net346),
    .X(_02194_));
 sg13g2_o21ai_1 _07739_ (.B1(_02184_),
    .Y(_02195_),
    .A1(_01413_),
    .A2(_02194_));
 sg13g2_nand2_1 _07740_ (.Y(_02196_),
    .A(net280),
    .B(_02195_));
 sg13g2_nand4_1 _07741_ (.B(_02183_),
    .C(_02192_),
    .A(_02179_),
    .Y(_02197_),
    .D(_02196_));
 sg13g2_nand4_1 _07742_ (.B(_01391_),
    .C(_01788_),
    .A(_01388_),
    .Y(_02198_),
    .D(_01790_));
 sg13g2_a22oi_1 _07743_ (.Y(_02199_),
    .B1(_01634_),
    .B2(net283),
    .A2(_01349_),
    .A1(_01333_));
 sg13g2_nand2_1 _07744_ (.Y(_02200_),
    .A(net295),
    .B(_01210_));
 sg13g2_nand3_1 _07745_ (.B(_02173_),
    .C(_02200_),
    .A(_02199_),
    .Y(_02201_));
 sg13g2_nand3_1 _07746_ (.B(_01244_),
    .C(_02174_),
    .A(_01814_),
    .Y(_02202_));
 sg13g2_nor3_1 _07747_ (.A(_02198_),
    .B(_02201_),
    .C(_02202_),
    .Y(_02203_));
 sg13g2_nor2_1 _07748_ (.A(net297),
    .B(_01265_),
    .Y(_02204_));
 sg13g2_o21ai_1 _07749_ (.B1(net313),
    .Y(_02205_),
    .A1(_01670_),
    .A2(_02204_));
 sg13g2_nand2_1 _07750_ (.Y(_02206_),
    .A(_01294_),
    .B(_01474_));
 sg13g2_o21ai_1 _07751_ (.B1(_02206_),
    .Y(_02207_),
    .A1(net313),
    .A2(_02204_));
 sg13g2_a21o_1 _07752_ (.A2(_02205_),
    .A1(net280),
    .B1(_02207_),
    .X(_02208_));
 sg13g2_nand4_1 _07753_ (.B(_01478_),
    .C(_02203_),
    .A(_01468_),
    .Y(_02209_),
    .D(_02208_));
 sg13g2_or2_1 _07754_ (.X(_02210_),
    .B(_02209_),
    .A(_02197_));
 sg13g2_nand4_1 _07755_ (.B(_02173_),
    .C(_02174_),
    .A(_02172_),
    .Y(_02211_),
    .D(_02210_));
 sg13g2_o21ai_1 _07756_ (.B1(_01210_),
    .Y(_02212_),
    .A1(net295),
    .A2(net284));
 sg13g2_and2_1 _07757_ (.A(_02173_),
    .B(_02212_),
    .X(_02213_));
 sg13g2_buf_1 _07758_ (.A(_02213_),
    .X(_02214_));
 sg13g2_nand2_1 _07759_ (.Y(_02215_),
    .A(_02210_),
    .B(_02214_));
 sg13g2_xnor2_1 _07760_ (.Y(_02216_),
    .A(_02215_),
    .B(_01201_));
 sg13g2_and2_1 _07761_ (.A(_02211_),
    .B(_02216_),
    .X(_02217_));
 sg13g2_nand2b_1 _07762_ (.Y(_02218_),
    .B(_02172_),
    .A_N(_02201_));
 sg13g2_nand2b_1 _07763_ (.Y(_02219_),
    .B(_00404_),
    .A_N(_02218_));
 sg13g2_nand3b_1 _07764_ (.B(_05199_),
    .C(_05144_),
    .Y(_02220_),
    .A_N(_05225_));
 sg13g2_nand3_1 _07765_ (.B(_01580_),
    .C(_00489_),
    .A(net328),
    .Y(_02221_));
 sg13g2_nand3_1 _07766_ (.B(_02220_),
    .C(_02221_),
    .A(_02214_),
    .Y(_02222_));
 sg13g2_o21ai_1 _07767_ (.B1(_02222_),
    .Y(_02223_),
    .A1(_02214_),
    .A2(_01600_));
 sg13g2_o21ai_1 _07768_ (.B1(_02218_),
    .Y(_02224_),
    .A1(_02211_),
    .A2(_02223_));
 sg13g2_o21ai_1 _07769_ (.B1(_02224_),
    .Y(_02225_),
    .A1(_02212_),
    .A2(_02219_));
 sg13g2_nand2_1 _07770_ (.Y(_02226_),
    .A(_00412_),
    .B(_02214_));
 sg13g2_xnor2_1 _07771_ (.Y(_02227_),
    .A(_05268_),
    .B(_01126_));
 sg13g2_o21ai_1 _07772_ (.B1(_02215_),
    .Y(_02228_),
    .A1(_05244_),
    .A2(_02227_));
 sg13g2_nand4_1 _07773_ (.B(_02218_),
    .C(_02226_),
    .A(_02211_),
    .Y(_02229_),
    .D(_02228_));
 sg13g2_o21ai_1 _07774_ (.B1(_02229_),
    .Y(_02230_),
    .A1(_02217_),
    .A2(_02225_));
 sg13g2_and2_1 _07775_ (.A(net419),
    .B(_02230_),
    .X(_02231_));
 sg13g2_buf_1 _07776_ (.A(_02231_),
    .X(_02232_));
 sg13g2_o21ai_1 _07777_ (.B1(_01402_),
    .Y(_02233_),
    .A1(_05143_),
    .A2(_01236_));
 sg13g2_nor2_1 _07778_ (.A(net308),
    .B(_01402_),
    .Y(_02234_));
 sg13g2_a21oi_1 _07779_ (.A1(net313),
    .A2(_02233_),
    .Y(_02235_),
    .B1(_02234_));
 sg13g2_o21ai_1 _07780_ (.B1(_02183_),
    .Y(_02236_),
    .A1(net280),
    .A2(_02235_));
 sg13g2_nand2_1 _07781_ (.Y(_02237_),
    .A(_01659_),
    .B(_01802_));
 sg13g2_o21ai_1 _07782_ (.B1(_01379_),
    .Y(_02238_),
    .A1(_01398_),
    .A2(_01236_));
 sg13g2_a21oi_1 _07783_ (.A1(_01358_),
    .A2(_01324_),
    .Y(_02239_),
    .B1(_01803_));
 sg13g2_a21oi_1 _07784_ (.A1(_01298_),
    .A2(_01392_),
    .Y(_02240_),
    .B1(_02239_));
 sg13g2_a21oi_1 _07785_ (.A1(_01278_),
    .A2(_02238_),
    .Y(_02241_),
    .B1(_02240_));
 sg13g2_o21ai_1 _07786_ (.B1(_01809_),
    .Y(_02242_),
    .A1(_00442_),
    .A2(_01384_));
 sg13g2_and2_1 _07787_ (.A(_01644_),
    .B(_01645_),
    .X(_02243_));
 sg13g2_nand4_1 _07788_ (.B(_02241_),
    .C(_02242_),
    .A(_01244_),
    .Y(_02244_),
    .D(_02243_));
 sg13g2_nor3_1 _07789_ (.A(_02236_),
    .B(_02237_),
    .C(_02244_),
    .Y(_02245_));
 sg13g2_nand3b_1 _07790_ (.B(_01446_),
    .C(_02245_),
    .Y(_02246_),
    .A_N(_01827_));
 sg13g2_nor2_1 _07791_ (.A(net249),
    .B(_02246_),
    .Y(_02247_));
 sg13g2_nand4_1 _07792_ (.B(_02232_),
    .C(_01693_),
    .A(net370),
    .Y(_02248_),
    .D(_02247_));
 sg13g2_mux2_1 _07793_ (.A0(_02169_),
    .A1(\dtop.player_inst.synth.alu.oct_en ),
    .S(_02248_),
    .X(_00110_));
 sg13g2_buf_1 _07794_ (.A(\dtop.vtop.pipeline.wave_index[0] ),
    .X(_02249_));
 sg13g2_buf_2 _07795_ (.A(\dtop.vtop.pipeline.wave_index[1] ),
    .X(_02250_));
 sg13g2_inv_1 _07796_ (.Y(_02251_),
    .A(_02250_));
 sg13g2_nor3_2 _07797_ (.A(_02249_),
    .B(_02251_),
    .C(net277),
    .Y(_02252_));
 sg13g2_a21oi_1 _07798_ (.A1(net394),
    .A2(net277),
    .Y(_02253_),
    .B1(_02252_));
 sg13g2_buf_1 _07799_ (.A(_02253_),
    .X(_02254_));
 sg13g2_and2_1 _07800_ (.A(net428),
    .B(_05194_),
    .X(_02255_));
 sg13g2_buf_1 _07801_ (.A(_02255_),
    .X(_02256_));
 sg13g2_buf_1 _07802_ (.A(_00004_),
    .X(_02257_));
 sg13g2_buf_2 _07803_ (.A(_00006_),
    .X(_02258_));
 sg13g2_and2_1 _07804_ (.A(_02257_),
    .B(_02258_),
    .X(_02259_));
 sg13g2_buf_1 _07805_ (.A(_02259_),
    .X(_02260_));
 sg13g2_mux2_1 _07806_ (.A0(_02256_),
    .A1(_02260_),
    .S(net303),
    .X(_02261_));
 sg13g2_buf_2 _07807_ (.A(_02261_),
    .X(_02262_));
 sg13g2_nand2_1 _07808_ (.Y(_02263_),
    .A(_00003_),
    .B(_02262_));
 sg13g2_inv_1 _07809_ (.Y(_02264_),
    .A(_02257_));
 sg13g2_mux2_1 _07810_ (.A0(_02264_),
    .A1(_05195_),
    .S(net301),
    .X(_02265_));
 sg13g2_buf_8 _07811_ (.A(_02265_),
    .X(_02266_));
 sg13g2_nor2_1 _07812_ (.A(_02258_),
    .B(\dtop.vtop.pipeline.phases[2][15] ),
    .Y(_02267_));
 sg13g2_nor2_1 _07813_ (.A(net428),
    .B(\dtop.vtop.pipeline.phases[2][15] ),
    .Y(_02268_));
 sg13g2_mux2_1 _07814_ (.A0(_02267_),
    .A1(_02268_),
    .S(net301),
    .X(_02269_));
 sg13g2_mux2_1 _07815_ (.A0(\dtop.vtop.pipeline.zg_acc[8] ),
    .A1(\dtop.vtop.pipeline.phases[1][15] ),
    .S(_02258_),
    .X(_02270_));
 sg13g2_nand2_1 _07816_ (.Y(_02271_),
    .A(_02264_),
    .B(_02270_));
 sg13g2_mux2_1 _07817_ (.A0(\dtop.vtop.pipeline.zg_acc[8] ),
    .A1(\dtop.vtop.pipeline.phases[1][15] ),
    .S(net428),
    .X(_02272_));
 sg13g2_nand2_1 _07818_ (.Y(_02273_),
    .A(_05195_),
    .B(_02272_));
 sg13g2_mux2_1 _07819_ (.A0(_02271_),
    .A1(_02273_),
    .S(net301),
    .X(_02274_));
 sg13g2_o21ai_1 _07820_ (.B1(_02274_),
    .Y(_02275_),
    .A1(_02266_),
    .A2(_02269_));
 sg13g2_nand2_1 _07821_ (.Y(_02276_),
    .A(_02263_),
    .B(_02275_));
 sg13g2_buf_1 _07822_ (.A(_02276_),
    .X(_02277_));
 sg13g2_nand2b_1 _07823_ (.Y(_02278_),
    .B(_05397_),
    .A_N(_05131_));
 sg13g2_nand3b_1 _07824_ (.B(_05149_),
    .C(net402),
    .Y(_02279_),
    .A_N(_05136_));
 sg13g2_a21oi_1 _07825_ (.A1(_02278_),
    .A2(_02279_),
    .Y(_02280_),
    .B1(_01199_));
 sg13g2_nand2_1 _07826_ (.Y(_02281_),
    .A(_05253_),
    .B(_05136_));
 sg13g2_nor2_1 _07827_ (.A(_05264_),
    .B(_02281_),
    .Y(_02282_));
 sg13g2_a21oi_1 _07828_ (.A1(net303),
    .A2(_02280_),
    .Y(_02283_),
    .B1(_02282_));
 sg13g2_inv_1 _07829_ (.Y(_02284_),
    .A(_02283_));
 sg13g2_nor2_1 _07830_ (.A(net247),
    .B(_02284_),
    .Y(_02285_));
 sg13g2_buf_1 _07831_ (.A(_02285_),
    .X(_02286_));
 sg13g2_buf_2 _07832_ (.A(_02286_),
    .X(_02287_));
 sg13g2_nor2b_1 _07833_ (.A(_02258_),
    .B_N(_02257_),
    .Y(_02288_));
 sg13g2_nand2b_1 _07834_ (.Y(_02289_),
    .B(_05194_),
    .A_N(_00090_));
 sg13g2_nor4_2 _07835_ (.A(_05170_),
    .B(_05173_),
    .C(_05175_),
    .Y(_02290_),
    .D(_02289_));
 sg13g2_a21o_1 _07836_ (.A2(_02288_),
    .A1(net303),
    .B1(_02290_),
    .X(_02291_));
 sg13g2_buf_1 _07837_ (.A(_02291_),
    .X(_02292_));
 sg13g2_inv_1 _07838_ (.Y(_02293_),
    .A(\dtop.vtop.pipeline.phases[2][9] ));
 sg13g2_a22oi_1 _07839_ (.Y(_02294_),
    .B1(net275),
    .B2(_02293_),
    .A2(_02262_),
    .A1(_00049_));
 sg13g2_buf_1 _07840_ (.A(_02294_),
    .X(_02295_));
 sg13g2_buf_1 _07841_ (.A(_02258_),
    .X(_02296_));
 sg13g2_and2_1 _07842_ (.A(_02296_),
    .B(\dtop.vtop.pipeline.phases[1][9] ),
    .X(_02297_));
 sg13g2_buf_1 _07843_ (.A(\dtop.vtop.pipeline.zg_acc[2] ),
    .X(_02298_));
 sg13g2_inv_2 _07844_ (.Y(_02299_),
    .A(_02298_));
 sg13g2_nor2_1 _07845_ (.A(net369),
    .B(_02299_),
    .Y(_02300_));
 sg13g2_o21ai_1 _07846_ (.B1(net303),
    .Y(_02301_),
    .A1(_02297_),
    .A2(_02300_));
 sg13g2_and2_1 _07847_ (.A(net428),
    .B(\dtop.vtop.pipeline.phases[1][9] ),
    .X(_02302_));
 sg13g2_nor2_1 _07848_ (.A(net394),
    .B(_02299_),
    .Y(_02303_));
 sg13g2_o21ai_1 _07849_ (.B1(net301),
    .Y(_02304_),
    .A1(_02302_),
    .A2(_02303_));
 sg13g2_nand3_1 _07850_ (.B(_02301_),
    .C(_02304_),
    .A(_02266_),
    .Y(_02305_));
 sg13g2_buf_1 _07851_ (.A(_02305_),
    .X(_02306_));
 sg13g2_nand2_1 _07852_ (.Y(_02307_),
    .A(_02295_),
    .B(_02306_));
 sg13g2_buf_1 _07853_ (.A(_02307_),
    .X(_02308_));
 sg13g2_buf_1 _07854_ (.A(_02308_),
    .X(_02309_));
 sg13g2_mux2_1 _07855_ (.A0(_05185_),
    .A1(_02258_),
    .S(net303),
    .X(_02310_));
 sg13g2_buf_2 _07856_ (.A(_02310_),
    .X(_02311_));
 sg13g2_mux2_1 _07857_ (.A0(_02257_),
    .A1(_05194_),
    .S(net301),
    .X(_02312_));
 sg13g2_buf_2 _07858_ (.A(_02312_),
    .X(_02313_));
 sg13g2_a21o_1 _07859_ (.A2(_02311_),
    .A1(\dtop.vtop.pipeline.phases[1][6] ),
    .B1(_02313_),
    .X(_02314_));
 sg13g2_buf_1 _07860_ (.A(_02314_),
    .X(_02315_));
 sg13g2_and2_1 _07861_ (.A(net369),
    .B(\dtop.vtop.pipeline.phases[0][6] ),
    .X(_02316_));
 sg13g2_nor2b_1 _07862_ (.A(_02296_),
    .B_N(\dtop.vtop.pipeline.phases[2][6] ),
    .Y(_02317_));
 sg13g2_o21ai_1 _07863_ (.B1(net290),
    .Y(_02318_),
    .A1(_02316_),
    .A2(_02317_));
 sg13g2_and2_1 _07864_ (.A(net428),
    .B(\dtop.vtop.pipeline.phases[0][6] ),
    .X(_02319_));
 sg13g2_nor2b_1 _07865_ (.A(net394),
    .B_N(\dtop.vtop.pipeline.phases[2][6] ),
    .Y(_02320_));
 sg13g2_o21ai_1 _07866_ (.B1(net289),
    .Y(_02321_),
    .A1(_02319_),
    .A2(_02320_));
 sg13g2_nand3_1 _07867_ (.B(_02318_),
    .C(_02321_),
    .A(_02313_),
    .Y(_02322_));
 sg13g2_buf_1 _07868_ (.A(_02322_),
    .X(_02323_));
 sg13g2_nand2_1 _07869_ (.Y(_02324_),
    .A(_02315_),
    .B(net258));
 sg13g2_buf_1 _07870_ (.A(_02324_),
    .X(_02325_));
 sg13g2_nand2_1 _07871_ (.Y(_02326_),
    .A(net198),
    .B(_02325_));
 sg13g2_buf_1 _07872_ (.A(_02306_),
    .X(_02327_));
 sg13g2_and2_1 _07873_ (.A(_02295_),
    .B(net246),
    .X(_02328_));
 sg13g2_buf_1 _07874_ (.A(_02328_),
    .X(_02329_));
 sg13g2_buf_1 _07875_ (.A(_02315_),
    .X(_02330_));
 sg13g2_and2_1 _07876_ (.A(net245),
    .B(net258),
    .X(_02331_));
 sg13g2_buf_2 _07877_ (.A(_02331_),
    .X(_02332_));
 sg13g2_inv_1 _07878_ (.Y(_02333_),
    .A(\dtop.vtop.pipeline.phases[2][8] ));
 sg13g2_and2_1 _07879_ (.A(_02333_),
    .B(_02288_),
    .X(_02334_));
 sg13g2_a22oi_1 _07880_ (.Y(_02335_),
    .B1(_02334_),
    .B2(net303),
    .A2(_02290_),
    .A1(_02333_));
 sg13g2_nand2_1 _07881_ (.Y(_02336_),
    .A(_00046_),
    .B(_02260_));
 sg13g2_nand2_1 _07882_ (.Y(_02337_),
    .A(_00046_),
    .B(_02256_));
 sg13g2_mux2_1 _07883_ (.A0(_02336_),
    .A1(_02337_),
    .S(net301),
    .X(_02338_));
 sg13g2_nand2_1 _07884_ (.Y(_02339_),
    .A(_02335_),
    .B(_02338_));
 sg13g2_inv_1 _07885_ (.Y(_02340_),
    .A(_02258_));
 sg13g2_nor2_1 _07886_ (.A(_02340_),
    .B(\dtop.vtop.pipeline.phases[1][8] ),
    .Y(_02341_));
 sg13g2_buf_2 _07887_ (.A(_00047_),
    .X(_02342_));
 sg13g2_nor2b_1 _07888_ (.A(net369),
    .B_N(_02342_),
    .Y(_02343_));
 sg13g2_o21ai_1 _07889_ (.B1(net303),
    .Y(_02344_),
    .A1(_02341_),
    .A2(_02343_));
 sg13g2_nor2_1 _07890_ (.A(_05186_),
    .B(\dtop.vtop.pipeline.phases[1][8] ),
    .Y(_02345_));
 sg13g2_nor2b_1 _07891_ (.A(net394),
    .B_N(_02342_),
    .Y(_02346_));
 sg13g2_o21ai_1 _07892_ (.B1(net301),
    .Y(_02347_),
    .A1(_02345_),
    .A2(_02346_));
 sg13g2_a21oi_1 _07893_ (.A1(_02344_),
    .A2(_02347_),
    .Y(_02348_),
    .B1(_02313_));
 sg13g2_nor2_1 _07894_ (.A(_02339_),
    .B(_02348_),
    .Y(_02349_));
 sg13g2_buf_2 _07895_ (.A(_02349_),
    .X(_02350_));
 sg13g2_nand3_1 _07896_ (.B(_02332_),
    .C(_02350_),
    .A(net197),
    .Y(_02351_));
 sg13g2_inv_1 _07897_ (.Y(_02352_),
    .A(\dtop.vtop.pipeline.phases[2][7] ));
 sg13g2_a22oi_1 _07898_ (.Y(_02353_),
    .B1(net275),
    .B2(_02352_),
    .A2(_02262_),
    .A1(_00044_));
 sg13g2_buf_1 _07899_ (.A(_02353_),
    .X(_02354_));
 sg13g2_and2_1 _07900_ (.A(net369),
    .B(\dtop.vtop.pipeline.phases[1][7] ),
    .X(_02355_));
 sg13g2_buf_1 _07901_ (.A(\dtop.vtop.pipeline.zg_acc[0] ),
    .X(_02356_));
 sg13g2_inv_1 _07902_ (.Y(_02357_),
    .A(_02356_));
 sg13g2_nor2_1 _07903_ (.A(net369),
    .B(_02357_),
    .Y(_02358_));
 sg13g2_o21ai_1 _07904_ (.B1(net290),
    .Y(_02359_),
    .A1(_02355_),
    .A2(_02358_));
 sg13g2_and2_1 _07905_ (.A(net428),
    .B(\dtop.vtop.pipeline.phases[1][7] ),
    .X(_02360_));
 sg13g2_nor2_1 _07906_ (.A(net394),
    .B(_02357_),
    .Y(_02361_));
 sg13g2_o21ai_1 _07907_ (.B1(net289),
    .Y(_02362_),
    .A1(_02360_),
    .A2(_02361_));
 sg13g2_nand3_1 _07908_ (.B(_02359_),
    .C(_02362_),
    .A(_02266_),
    .Y(_02363_));
 sg13g2_buf_1 _07909_ (.A(_02363_),
    .X(_02364_));
 sg13g2_nand2_1 _07910_ (.Y(_02365_),
    .A(net257),
    .B(net256));
 sg13g2_buf_1 _07911_ (.A(_02365_),
    .X(_02366_));
 sg13g2_buf_1 _07912_ (.A(net229),
    .X(_02367_));
 sg13g2_a21oi_1 _07913_ (.A1(_02326_),
    .A2(_02351_),
    .Y(_02368_),
    .B1(net196));
 sg13g2_and2_1 _07914_ (.A(net257),
    .B(net256),
    .X(_02369_));
 sg13g2_buf_1 _07915_ (.A(_02369_),
    .X(_02370_));
 sg13g2_buf_1 _07916_ (.A(net228),
    .X(_02371_));
 sg13g2_buf_1 _07917_ (.A(net195),
    .X(_02372_));
 sg13g2_buf_1 _07918_ (.A(_02332_),
    .X(_02373_));
 sg13g2_buf_1 _07919_ (.A(net164),
    .X(_02374_));
 sg13g2_buf_1 _07920_ (.A(_02350_),
    .X(_02375_));
 sg13g2_buf_1 _07921_ (.A(_02375_),
    .X(_02376_));
 sg13g2_buf_1 _07922_ (.A(_02329_),
    .X(_02377_));
 sg13g2_buf_1 _07923_ (.A(net163),
    .X(_02378_));
 sg13g2_a21oi_1 _07924_ (.A1(_02374_),
    .A2(net194),
    .Y(_02379_),
    .B1(net125));
 sg13g2_nor2_1 _07925_ (.A(_02372_),
    .B(_02379_),
    .Y(_02380_));
 sg13g2_buf_1 _07926_ (.A(_00058_),
    .X(_02381_));
 sg13g2_nor2_1 _07927_ (.A(_02381_),
    .B(_02311_),
    .Y(_02382_));
 sg13g2_a21o_1 _07928_ (.A2(_02311_),
    .A1(\dtop.vtop.pipeline.phases[1][14] ),
    .B1(_02313_),
    .X(_02383_));
 sg13g2_inv_1 _07929_ (.Y(_02384_),
    .A(\dtop.vtop.pipeline.phases[2][14] ));
 sg13g2_a22oi_1 _07930_ (.Y(_02385_),
    .B1(net275),
    .B2(_02384_),
    .A2(_02262_),
    .A1(_00057_));
 sg13g2_o21ai_1 _07931_ (.B1(_02385_),
    .Y(_02386_),
    .A1(_02382_),
    .A2(_02383_));
 sg13g2_buf_8 _07932_ (.A(_02386_),
    .X(_02387_));
 sg13g2_nand3_1 _07933_ (.B(_02275_),
    .C(_02284_),
    .A(_02263_),
    .Y(_02388_));
 sg13g2_buf_2 _07934_ (.A(_02388_),
    .X(_02389_));
 sg13g2_xor2_1 _07935_ (.B(_02389_),
    .A(_02387_),
    .X(_02390_));
 sg13g2_buf_8 _07936_ (.A(_02390_),
    .X(_02391_));
 sg13g2_buf_8 _07937_ (.A(_02391_),
    .X(_02392_));
 sg13g2_buf_8 _07938_ (.A(_02392_),
    .X(_02393_));
 sg13g2_inv_1 _07939_ (.Y(_02394_),
    .A(\dtop.vtop.pipeline.phases[2][10] ));
 sg13g2_a22oi_1 _07940_ (.Y(_02395_),
    .B1(_02292_),
    .B2(_02394_),
    .A2(_02262_),
    .A1(_00051_));
 sg13g2_buf_2 _07941_ (.A(_02395_),
    .X(_02396_));
 sg13g2_inv_1 _07942_ (.Y(_02397_),
    .A(\dtop.vtop.pipeline.phases[1][10] ));
 sg13g2_nor2_1 _07943_ (.A(_02340_),
    .B(_02397_),
    .Y(_02398_));
 sg13g2_buf_1 _07944_ (.A(\dtop.vtop.pipeline.zg_acc[3] ),
    .X(_02399_));
 sg13g2_inv_1 _07945_ (.Y(_02400_),
    .A(_02399_));
 sg13g2_nor2_1 _07946_ (.A(net369),
    .B(_02400_),
    .Y(_02401_));
 sg13g2_o21ai_1 _07947_ (.B1(_05177_),
    .Y(_02402_),
    .A1(_02398_),
    .A2(_02401_));
 sg13g2_nor2_1 _07948_ (.A(_05186_),
    .B(_02397_),
    .Y(_02403_));
 sg13g2_nor2_1 _07949_ (.A(net394),
    .B(_02400_),
    .Y(_02404_));
 sg13g2_o21ai_1 _07950_ (.B1(net301),
    .Y(_02405_),
    .A1(_02403_),
    .A2(_02404_));
 sg13g2_nand3_1 _07951_ (.B(_02402_),
    .C(_02405_),
    .A(_02266_),
    .Y(_02406_));
 sg13g2_buf_1 _07952_ (.A(_02406_),
    .X(_02407_));
 sg13g2_nand2_1 _07953_ (.Y(_02408_),
    .A(_02396_),
    .B(_02407_));
 sg13g2_buf_2 _07954_ (.A(_02408_),
    .X(_02409_));
 sg13g2_buf_1 _07955_ (.A(_02409_),
    .X(_02410_));
 sg13g2_buf_1 _07956_ (.A(net193),
    .X(_02411_));
 sg13g2_nor2_1 _07957_ (.A(net124),
    .B(net161),
    .Y(_02412_));
 sg13g2_o21ai_1 _07958_ (.B1(_02412_),
    .Y(_02413_),
    .A1(_02368_),
    .A2(_02380_));
 sg13g2_nor2_1 _07959_ (.A(net228),
    .B(net230),
    .Y(_02414_));
 sg13g2_o21ai_1 _07960_ (.B1(net229),
    .Y(_02415_),
    .A1(net198),
    .A2(_02332_));
 sg13g2_xnor2_1 _07961_ (.Y(_02416_),
    .A(_02387_),
    .B(_02389_));
 sg13g2_buf_8 _07962_ (.A(_02416_),
    .X(_02417_));
 sg13g2_mux2_1 _07963_ (.A0(_02414_),
    .A1(_02415_),
    .S(_02417_),
    .X(_02418_));
 sg13g2_buf_1 _07964_ (.A(_02308_),
    .X(_02419_));
 sg13g2_and4_1 _07965_ (.A(net257),
    .B(net256),
    .C(net245),
    .D(net258),
    .X(_02420_));
 sg13g2_buf_1 _07966_ (.A(_02420_),
    .X(_02421_));
 sg13g2_buf_1 _07967_ (.A(_02421_),
    .X(_02422_));
 sg13g2_buf_1 _07968_ (.A(_02350_),
    .X(_02423_));
 sg13g2_o21ai_1 _07969_ (.B1(net226),
    .Y(_02424_),
    .A1(net192),
    .A2(net160));
 sg13g2_buf_1 _07970_ (.A(net229),
    .X(_02425_));
 sg13g2_nor2_1 _07971_ (.A(_02417_),
    .B(net191),
    .Y(_02426_));
 sg13g2_buf_8 _07972_ (.A(_02417_),
    .X(_02427_));
 sg13g2_and2_1 _07973_ (.A(_02335_),
    .B(_02338_),
    .X(_02428_));
 sg13g2_buf_2 _07974_ (.A(_02428_),
    .X(_02429_));
 sg13g2_a21o_1 _07975_ (.A2(_02347_),
    .A1(_02344_),
    .B1(_02313_),
    .X(_02430_));
 sg13g2_buf_2 _07976_ (.A(_02430_),
    .X(_02431_));
 sg13g2_nand2_1 _07977_ (.Y(_02432_),
    .A(_02429_),
    .B(_02431_));
 sg13g2_buf_2 _07978_ (.A(_02432_),
    .X(_02433_));
 sg13g2_nand2_1 _07979_ (.Y(_02434_),
    .A(net230),
    .B(_02433_));
 sg13g2_a22oi_1 _07980_ (.Y(_02435_),
    .B1(_02429_),
    .B2(_02431_),
    .A2(net256),
    .A1(net257));
 sg13g2_buf_1 _07981_ (.A(_02435_),
    .X(_02436_));
 sg13g2_nand2_1 _07982_ (.Y(_02437_),
    .A(_02308_),
    .B(_02436_));
 sg13g2_o21ai_1 _07983_ (.B1(_02437_),
    .Y(_02438_),
    .A1(net159),
    .A2(_02434_));
 sg13g2_a221oi_1 _07984_ (.B2(_02426_),
    .C1(_02438_),
    .B1(_02424_),
    .A1(net194),
    .Y(_02439_),
    .A2(_02418_));
 sg13g2_buf_8 _07985_ (.A(_02391_),
    .X(_02440_));
 sg13g2_a22oi_1 _07986_ (.Y(_02441_),
    .B1(net245),
    .B2(net258),
    .A2(net256),
    .A1(net257));
 sg13g2_buf_2 _07987_ (.A(_02441_),
    .X(_02442_));
 sg13g2_buf_1 _07988_ (.A(_02442_),
    .X(_02443_));
 sg13g2_a21oi_1 _07989_ (.A1(net158),
    .A2(net157),
    .Y(_02444_),
    .B1(net160));
 sg13g2_nor2_1 _07990_ (.A(net125),
    .B(_02444_),
    .Y(_02445_));
 sg13g2_buf_8 _07991_ (.A(net159),
    .X(_02446_));
 sg13g2_and2_1 _07992_ (.A(_02396_),
    .B(_02407_),
    .X(_02447_));
 sg13g2_buf_2 _07993_ (.A(_02447_),
    .X(_02448_));
 sg13g2_buf_8 _07994_ (.A(_02448_),
    .X(_02449_));
 sg13g2_buf_1 _07995_ (.A(net190),
    .X(_02450_));
 sg13g2_buf_1 _07996_ (.A(net156),
    .X(_02451_));
 sg13g2_nor2_1 _07997_ (.A(net123),
    .B(net122),
    .Y(_02452_));
 sg13g2_o21ai_1 _07998_ (.B1(_02452_),
    .Y(_02453_),
    .A1(_02439_),
    .A2(_02445_));
 sg13g2_buf_2 _07999_ (.A(_02313_),
    .X(_02454_));
 sg13g2_buf_2 _08000_ (.A(\dtop.vtop.pipeline.zg_acc[4] ),
    .X(_02455_));
 sg13g2_mux2_1 _08001_ (.A0(_02455_),
    .A1(\dtop.vtop.pipeline.phases[1][11] ),
    .S(_02311_),
    .X(_02456_));
 sg13g2_inv_1 _08002_ (.Y(_02457_),
    .A(\dtop.vtop.pipeline.phases[2][11] ));
 sg13g2_a22oi_1 _08003_ (.Y(_02458_),
    .B1(net275),
    .B2(_02457_),
    .A2(_02262_),
    .A1(_00053_));
 sg13g2_o21ai_1 _08004_ (.B1(_02458_),
    .Y(_02459_),
    .A1(net271),
    .A2(_02456_));
 sg13g2_buf_1 _08005_ (.A(_02459_),
    .X(_02460_));
 sg13g2_buf_1 _08006_ (.A(net244),
    .X(_02461_));
 sg13g2_buf_1 _08007_ (.A(net225),
    .X(_02462_));
 sg13g2_a21oi_1 _08008_ (.A1(_02413_),
    .A2(_02453_),
    .Y(_02463_),
    .B1(_02462_));
 sg13g2_mux2_1 _08009_ (.A0(_05186_),
    .A1(_02340_),
    .S(net290),
    .X(_02464_));
 sg13g2_buf_1 _08010_ (.A(_02464_),
    .X(_02465_));
 sg13g2_nand2_1 _08011_ (.Y(_02466_),
    .A(_02455_),
    .B(_02465_));
 sg13g2_a21oi_1 _08012_ (.A1(\dtop.vtop.pipeline.phases[1][11] ),
    .A2(_02311_),
    .Y(_02467_),
    .B1(_02313_));
 sg13g2_a21oi_1 _08013_ (.A1(net290),
    .A2(_02288_),
    .Y(_02468_),
    .B1(_02290_));
 sg13g2_buf_2 _08014_ (.A(_02468_),
    .X(_02469_));
 sg13g2_nor2_1 _08015_ (.A(\dtop.vtop.pipeline.phases[2][11] ),
    .B(_02469_),
    .Y(_02470_));
 sg13g2_a221oi_1 _08016_ (.B2(_02467_),
    .C1(_02470_),
    .B1(_02466_),
    .A1(_00053_),
    .Y(_02471_),
    .A2(_02262_));
 sg13g2_buf_1 _08017_ (.A(_02471_),
    .X(_02472_));
 sg13g2_buf_1 _08018_ (.A(_02472_),
    .X(_02473_));
 sg13g2_buf_1 _08019_ (.A(net188),
    .X(_02474_));
 sg13g2_buf_1 _08020_ (.A(net155),
    .X(_02475_));
 sg13g2_xnor2_1 _08021_ (.Y(_02476_),
    .A(_02391_),
    .B(_02350_));
 sg13g2_buf_2 _08022_ (.A(_02476_),
    .X(_02477_));
 sg13g2_buf_1 _08023_ (.A(net230),
    .X(_02478_));
 sg13g2_buf_1 _08024_ (.A(_02478_),
    .X(_02479_));
 sg13g2_nor2_2 _08025_ (.A(net191),
    .B(_02309_),
    .Y(_02480_));
 sg13g2_nand2_1 _08026_ (.Y(_02481_),
    .A(net229),
    .B(net198));
 sg13g2_o21ai_1 _08027_ (.B1(_02481_),
    .Y(_02482_),
    .A1(net154),
    .A2(_02480_));
 sg13g2_nand2b_1 _08028_ (.Y(_02483_),
    .B(_02482_),
    .A_N(_02477_));
 sg13g2_buf_1 _08029_ (.A(net161),
    .X(_02484_));
 sg13g2_buf_1 _08030_ (.A(_02417_),
    .X(_02485_));
 sg13g2_nand2_1 _08031_ (.Y(_02486_),
    .A(net230),
    .B(_02350_));
 sg13g2_nor2_1 _08032_ (.A(_02485_),
    .B(_02486_),
    .Y(_02487_));
 sg13g2_buf_8 _08033_ (.A(_02391_),
    .X(_02488_));
 sg13g2_nor3_1 _08034_ (.A(_02488_),
    .B(net154),
    .C(_02481_),
    .Y(_02489_));
 sg13g2_nor3_1 _08035_ (.A(net120),
    .B(_02487_),
    .C(_02489_),
    .Y(_02490_));
 sg13g2_buf_1 _08036_ (.A(_02295_),
    .X(_02491_));
 sg13g2_and4_1 _08037_ (.A(net243),
    .B(net246),
    .C(_02429_),
    .D(_02431_),
    .X(_02492_));
 sg13g2_buf_1 _08038_ (.A(_02492_),
    .X(_02493_));
 sg13g2_and2_1 _08039_ (.A(net162),
    .B(_02493_),
    .X(_02494_));
 sg13g2_nor2_1 _08040_ (.A(net197),
    .B(_02433_),
    .Y(_02495_));
 sg13g2_nor3_1 _08041_ (.A(net162),
    .B(net164),
    .C(_02495_),
    .Y(_02496_));
 sg13g2_o21ai_1 _08042_ (.B1(net165),
    .Y(_02497_),
    .A1(_02494_),
    .A2(_02496_));
 sg13g2_nand3_1 _08043_ (.B(_02490_),
    .C(_02497_),
    .A(_02483_),
    .Y(_02498_));
 sg13g2_and2_1 _08044_ (.A(_02301_),
    .B(_02304_),
    .X(_02499_));
 sg13g2_buf_1 _08045_ (.A(_02266_),
    .X(_02500_));
 sg13g2_nand2_1 _08046_ (.Y(_02501_),
    .A(_00049_),
    .B(_02260_));
 sg13g2_nand2_1 _08047_ (.Y(_02502_),
    .A(_00049_),
    .B(_02256_));
 sg13g2_mux2_1 _08048_ (.A0(_02501_),
    .A1(_02502_),
    .S(net289),
    .X(_02503_));
 sg13g2_o21ai_1 _08049_ (.B1(_02503_),
    .Y(_02504_),
    .A1(\dtop.vtop.pipeline.phases[2][9] ),
    .A2(_02469_));
 sg13g2_a221oi_1 _08050_ (.B2(net270),
    .C1(_02504_),
    .B1(_02499_),
    .A1(net257),
    .Y(_02505_),
    .A2(net256));
 sg13g2_buf_2 _08051_ (.A(_02505_),
    .X(_02506_));
 sg13g2_and2_1 _08052_ (.A(_02359_),
    .B(_02362_),
    .X(_02507_));
 sg13g2_buf_8 _08053_ (.A(_02469_),
    .X(_02508_));
 sg13g2_nand2_1 _08054_ (.Y(_02509_),
    .A(_00044_),
    .B(_02260_));
 sg13g2_nand2_1 _08055_ (.Y(_02510_),
    .A(_00044_),
    .B(_02256_));
 sg13g2_mux2_1 _08056_ (.A0(_02509_),
    .A1(_02510_),
    .S(_05236_),
    .X(_02511_));
 sg13g2_o21ai_1 _08057_ (.B1(_02511_),
    .Y(_02512_),
    .A1(\dtop.vtop.pipeline.phases[2][7] ),
    .A2(_02508_));
 sg13g2_a221oi_1 _08058_ (.B2(net246),
    .C1(_02512_),
    .B1(net243),
    .A1(net270),
    .Y(_02513_),
    .A2(_02507_));
 sg13g2_buf_2 _08059_ (.A(_02513_),
    .X(_02514_));
 sg13g2_nor3_1 _08060_ (.A(net152),
    .B(net156),
    .C(_02514_),
    .Y(_02515_));
 sg13g2_buf_1 _08061_ (.A(net227),
    .X(_02516_));
 sg13g2_buf_1 _08062_ (.A(net186),
    .X(_02517_));
 sg13g2_o21ai_1 _08063_ (.B1(net151),
    .Y(_02518_),
    .A1(_02506_),
    .A2(_02515_));
 sg13g2_nand2_1 _08064_ (.Y(_02519_),
    .A(net196),
    .B(net186));
 sg13g2_and2_1 _08065_ (.A(_02402_),
    .B(_02405_),
    .X(_02520_));
 sg13g2_nand2_1 _08066_ (.Y(_02521_),
    .A(_00051_),
    .B(_02260_));
 sg13g2_nand2_1 _08067_ (.Y(_02522_),
    .A(_00051_),
    .B(_02256_));
 sg13g2_mux2_1 _08068_ (.A0(_02521_),
    .A1(_02522_),
    .S(_05236_),
    .X(_02523_));
 sg13g2_o21ai_1 _08069_ (.B1(_02523_),
    .Y(_02524_),
    .A1(\dtop.vtop.pipeline.phases[2][10] ),
    .A2(_02469_));
 sg13g2_a221oi_1 _08070_ (.B2(_02306_),
    .C1(_02524_),
    .B1(net243),
    .A1(_02266_),
    .Y(_02525_),
    .A2(_02520_));
 sg13g2_buf_1 _08071_ (.A(_02525_),
    .X(_02526_));
 sg13g2_a221oi_1 _08072_ (.B2(_02266_),
    .C1(_02504_),
    .B1(_02499_),
    .A1(_02396_),
    .Y(_02527_),
    .A2(_02407_));
 sg13g2_buf_1 _08073_ (.A(_02527_),
    .X(_02528_));
 sg13g2_buf_1 _08074_ (.A(_02528_),
    .X(_02529_));
 sg13g2_and2_1 _08075_ (.A(_02366_),
    .B(net184),
    .X(_02530_));
 sg13g2_buf_1 _08076_ (.A(_02530_),
    .X(_02531_));
 sg13g2_a221oi_1 _08077_ (.B2(_02526_),
    .C1(_02531_),
    .B1(_02519_),
    .A1(net124),
    .Y(_02532_),
    .A2(_02514_));
 sg13g2_buf_1 _08078_ (.A(net154),
    .X(_02533_));
 sg13g2_a21o_1 _08079_ (.A2(_02532_),
    .A1(_02518_),
    .B1(net119),
    .X(_02534_));
 sg13g2_xnor2_1 _08080_ (.Y(_02535_),
    .A(_02449_),
    .B(net228));
 sg13g2_buf_1 _08081_ (.A(_02449_),
    .X(_02536_));
 sg13g2_buf_1 _08082_ (.A(_02370_),
    .X(_02537_));
 sg13g2_buf_1 _08083_ (.A(net197),
    .X(_02538_));
 sg13g2_buf_1 _08084_ (.A(_02433_),
    .X(_02539_));
 sg13g2_buf_1 _08085_ (.A(_02539_),
    .X(_02540_));
 sg13g2_nand4_1 _08086_ (.B(net183),
    .C(_02538_),
    .A(_02536_),
    .Y(_02541_),
    .D(net148));
 sg13g2_o21ai_1 _08087_ (.B1(_02541_),
    .Y(_02542_),
    .A1(net125),
    .A2(_02535_));
 sg13g2_or2_1 _08088_ (.X(_02543_),
    .B(_02514_),
    .A(_02506_));
 sg13g2_o21ai_1 _08089_ (.B1(_02462_),
    .Y(_02544_),
    .A1(_02434_),
    .A2(_02543_));
 sg13g2_a21oi_1 _08090_ (.A1(net119),
    .A2(_02542_),
    .Y(_02545_),
    .B1(_02544_));
 sg13g2_buf_1 _08091_ (.A(net123),
    .X(_02546_));
 sg13g2_a221oi_1 _08092_ (.B2(_02545_),
    .C1(_02546_),
    .B1(_02534_),
    .A1(_02475_),
    .Y(_02547_),
    .A2(_02498_));
 sg13g2_buf_8 _08093_ (.A(_02392_),
    .X(_02548_));
 sg13g2_buf_8 _08094_ (.A(net118),
    .X(_02549_));
 sg13g2_inv_1 _08095_ (.Y(_02550_),
    .A(\dtop.vtop.pipeline.phases[2][12] ));
 sg13g2_a22oi_1 _08096_ (.Y(_02551_),
    .B1(_02292_),
    .B2(_02550_),
    .A2(_02262_),
    .A1(_00054_));
 sg13g2_and2_1 _08097_ (.A(net369),
    .B(\dtop.vtop.pipeline.phases[1][12] ),
    .X(_02552_));
 sg13g2_buf_1 _08098_ (.A(\dtop.vtop.pipeline.zg_acc[5] ),
    .X(_02553_));
 sg13g2_nor2b_1 _08099_ (.A(net369),
    .B_N(_02553_),
    .Y(_02554_));
 sg13g2_o21ai_1 _08100_ (.B1(net290),
    .Y(_02555_),
    .A1(_02552_),
    .A2(_02554_));
 sg13g2_nand3_1 _08101_ (.B(\dtop.vtop.pipeline.phases[1][12] ),
    .C(net289),
    .A(net394),
    .Y(_02556_));
 sg13g2_nand3_1 _08102_ (.B(_02553_),
    .C(net289),
    .A(_05186_),
    .Y(_02557_));
 sg13g2_nand4_1 _08103_ (.B(_02555_),
    .C(_02556_),
    .A(_02266_),
    .Y(_02558_),
    .D(_02557_));
 sg13g2_nand2_1 _08104_ (.Y(_02559_),
    .A(_02551_),
    .B(_02558_));
 sg13g2_buf_2 _08105_ (.A(_02559_),
    .X(_02560_));
 sg13g2_buf_1 _08106_ (.A(_02560_),
    .X(_02561_));
 sg13g2_nor2_1 _08107_ (.A(net97),
    .B(net224),
    .Y(_02562_));
 sg13g2_buf_1 _08108_ (.A(net198),
    .X(_02563_));
 sg13g2_buf_1 _08109_ (.A(net147),
    .X(_02564_));
 sg13g2_nand2_2 _08110_ (.Y(_02565_),
    .A(net229),
    .B(net230));
 sg13g2_nor2_1 _08111_ (.A(net117),
    .B(_02565_),
    .Y(_02566_));
 sg13g2_buf_1 _08112_ (.A(_02433_),
    .X(_02567_));
 sg13g2_buf_1 _08113_ (.A(net181),
    .X(_02568_));
 sg13g2_a22oi_1 _08114_ (.Y(_02569_),
    .B1(net243),
    .B2(net246),
    .A2(net256),
    .A1(net257));
 sg13g2_buf_1 _08115_ (.A(_02569_),
    .X(_02570_));
 sg13g2_a21oi_1 _08116_ (.A1(net126),
    .A2(_02570_),
    .Y(_02571_),
    .B1(_02480_));
 sg13g2_a22oi_1 _08117_ (.Y(_02572_),
    .B1(_02429_),
    .B2(_02431_),
    .A2(net246),
    .A1(net243));
 sg13g2_buf_1 _08118_ (.A(_02572_),
    .X(_02573_));
 sg13g2_mux2_1 _08119_ (.A0(net163),
    .A1(_02573_),
    .S(net187),
    .X(_02574_));
 sg13g2_nand2_1 _08120_ (.Y(_02575_),
    .A(net165),
    .B(_02574_));
 sg13g2_o21ai_1 _08121_ (.B1(_02575_),
    .Y(_02576_),
    .A1(net146),
    .A2(_02571_));
 sg13g2_nor2_1 _08122_ (.A(net189),
    .B(net122),
    .Y(_02577_));
 sg13g2_o21ai_1 _08123_ (.B1(_02577_),
    .Y(_02578_),
    .A1(_02566_),
    .A2(_02576_));
 sg13g2_and2_1 _08124_ (.A(_02551_),
    .B(_02558_),
    .X(_02579_));
 sg13g2_buf_1 _08125_ (.A(_02579_),
    .X(_02580_));
 sg13g2_buf_1 _08126_ (.A(_02580_),
    .X(_02581_));
 sg13g2_nor2_1 _08127_ (.A(net123),
    .B(_02581_),
    .Y(_02582_));
 sg13g2_a21oi_1 _08128_ (.A1(_02562_),
    .A2(_02578_),
    .Y(_02583_),
    .B1(_02582_));
 sg13g2_a22oi_1 _08129_ (.Y(_02584_),
    .B1(_02335_),
    .B2(_02338_),
    .A2(_02321_),
    .A1(_02318_));
 sg13g2_o21ai_1 _08130_ (.B1(net245),
    .Y(_02585_),
    .A1(_02348_),
    .A2(_02584_));
 sg13g2_buf_2 _08131_ (.A(_02585_),
    .X(_02586_));
 sg13g2_and2_1 _08132_ (.A(net120),
    .B(_02586_),
    .X(_02587_));
 sg13g2_o21ai_1 _08133_ (.B1(_02587_),
    .Y(_02588_),
    .A1(_02439_),
    .A2(_02445_));
 sg13g2_nand2_1 _08134_ (.Y(_02589_),
    .A(net225),
    .B(net123));
 sg13g2_a21oi_1 _08135_ (.A1(_02498_),
    .A2(_02588_),
    .Y(_02590_),
    .B1(_02589_));
 sg13g2_or4_1 _08136_ (.A(_02463_),
    .B(_02547_),
    .C(_02583_),
    .D(_02590_),
    .X(_02591_));
 sg13g2_nor2_2 _08137_ (.A(_02409_),
    .B(_02350_),
    .Y(_02592_));
 sg13g2_buf_8 _08138_ (.A(_02396_),
    .X(_02593_));
 sg13g2_buf_1 _08139_ (.A(_02407_),
    .X(_02594_));
 sg13g2_nand4_1 _08140_ (.B(net241),
    .C(net243),
    .A(net242),
    .Y(_02595_),
    .D(net246));
 sg13g2_buf_1 _08141_ (.A(_02595_),
    .X(_02596_));
 sg13g2_and4_1 _08142_ (.A(_02396_),
    .B(_02407_),
    .C(_02295_),
    .D(_02306_),
    .X(_02597_));
 sg13g2_buf_1 _08143_ (.A(_02597_),
    .X(_02598_));
 sg13g2_buf_1 _08144_ (.A(_02598_),
    .X(_02599_));
 sg13g2_o21ai_1 _08145_ (.B1(net126),
    .Y(_02600_),
    .A1(net148),
    .A2(net180));
 sg13g2_o21ai_1 _08146_ (.B1(_02600_),
    .Y(_02601_),
    .A1(net151),
    .A2(_02596_));
 sg13g2_buf_1 _08147_ (.A(net191),
    .X(_02602_));
 sg13g2_nand2_1 _08148_ (.Y(_02603_),
    .A(net187),
    .B(_02596_));
 sg13g2_a22oi_1 _08149_ (.Y(_02604_),
    .B1(net243),
    .B2(net246),
    .A2(net241),
    .A1(_02593_));
 sg13g2_buf_1 _08150_ (.A(_02604_),
    .X(_02605_));
 sg13g2_buf_1 _08151_ (.A(_02605_),
    .X(_02606_));
 sg13g2_o21ai_1 _08152_ (.B1(net183),
    .Y(_02607_),
    .A1(net154),
    .A2(net144));
 sg13g2_a21oi_1 _08153_ (.A1(_02603_),
    .A2(_02607_),
    .Y(_02608_),
    .B1(_02568_));
 sg13g2_a221oi_1 _08154_ (.B2(net145),
    .C1(_02608_),
    .B1(_02601_),
    .A1(net126),
    .Y(_02609_),
    .A2(_02592_));
 sg13g2_nand2_1 _08155_ (.Y(_02610_),
    .A(net152),
    .B(net223));
 sg13g2_nand4_1 _08156_ (.B(_02364_),
    .C(net245),
    .A(_02354_),
    .Y(_02611_),
    .D(net258));
 sg13g2_buf_1 _08157_ (.A(_02611_),
    .X(_02612_));
 sg13g2_buf_1 _08158_ (.A(_02612_),
    .X(_02613_));
 sg13g2_nand2_1 _08159_ (.Y(_02614_),
    .A(net143),
    .B(_02565_));
 sg13g2_xnor2_1 _08160_ (.Y(_02615_),
    .A(net146),
    .B(_02614_));
 sg13g2_nand3_1 _08161_ (.B(net224),
    .C(_02615_),
    .A(net98),
    .Y(_02616_));
 sg13g2_o21ai_1 _08162_ (.B1(_02616_),
    .Y(_02617_),
    .A1(_02609_),
    .A2(_02610_));
 sg13g2_buf_1 _08163_ (.A(net223),
    .X(_02618_));
 sg13g2_nand2_1 _08164_ (.Y(_02619_),
    .A(net189),
    .B(net179));
 sg13g2_buf_1 _08165_ (.A(_00056_),
    .X(_02620_));
 sg13g2_inv_1 _08166_ (.Y(_02621_),
    .A(\dtop.vtop.pipeline.phases[2][13] ));
 sg13g2_inv_1 _08167_ (.Y(_02622_),
    .A(\dtop.vtop.pipeline.phases[1][13] ));
 sg13g2_buf_1 _08168_ (.A(_02311_),
    .X(_02623_));
 sg13g2_mux4_1 _08169_ (.S0(net271),
    .A0(_02620_),
    .A1(_02621_),
    .A2(_02622_),
    .A3(_00055_),
    .S1(net269),
    .X(_02624_));
 sg13g2_buf_2 _08170_ (.A(_02624_),
    .X(_02625_));
 sg13g2_nor2_1 _08171_ (.A(net159),
    .B(_02625_),
    .Y(_02626_));
 sg13g2_o21ai_1 _08172_ (.B1(_02626_),
    .Y(_02627_),
    .A1(_02615_),
    .A2(_02619_));
 sg13g2_buf_1 _08173_ (.A(_02625_),
    .X(_02628_));
 sg13g2_nand2_1 _08174_ (.Y(_02629_),
    .A(net98),
    .B(net222));
 sg13g2_nand3_1 _08175_ (.B(_02603_),
    .C(_02607_),
    .A(net146),
    .Y(_02630_));
 sg13g2_nand2_1 _08176_ (.Y(_02631_),
    .A(_02344_),
    .B(_02347_));
 sg13g2_a221oi_1 _08177_ (.B2(net270),
    .C1(_02339_),
    .B1(_02631_),
    .A1(net242),
    .Y(_02632_),
    .A2(net241));
 sg13g2_buf_1 _08178_ (.A(_02632_),
    .X(_02633_));
 sg13g2_and2_1 _08179_ (.A(net227),
    .B(_02605_),
    .X(_02634_));
 sg13g2_o21ai_1 _08180_ (.B1(net119),
    .Y(_02635_),
    .A1(net151),
    .A2(net144));
 sg13g2_nand2b_1 _08181_ (.Y(_02636_),
    .B(_02635_),
    .A_N(_02634_));
 sg13g2_a22oi_1 _08182_ (.Y(_02637_),
    .B1(_02636_),
    .B2(net165),
    .A2(_02633_),
    .A1(net119));
 sg13g2_nor2_1 _08183_ (.A(_02472_),
    .B(_02580_),
    .Y(_02638_));
 sg13g2_buf_2 _08184_ (.A(_02638_),
    .X(_02639_));
 sg13g2_nand2_1 _08185_ (.Y(_02640_),
    .A(net153),
    .B(_02639_));
 sg13g2_a21oi_1 _08186_ (.A1(_02630_),
    .A2(_02637_),
    .Y(_02641_),
    .B1(_02640_));
 sg13g2_a221oi_1 _08187_ (.B2(_02629_),
    .C1(_02641_),
    .B1(_02627_),
    .A1(net121),
    .Y(_02642_),
    .A2(_02617_));
 sg13g2_nand2_1 _08188_ (.Y(_02643_),
    .A(net125),
    .B(_02535_));
 sg13g2_o21ai_1 _08189_ (.B1(_02486_),
    .Y(_02644_),
    .A1(net150),
    .A2(_02514_));
 sg13g2_nand2_2 _08190_ (.Y(_02645_),
    .A(net188),
    .B(net159));
 sg13g2_a221oi_1 _08191_ (.B2(_02644_),
    .C1(_02645_),
    .B1(_02643_),
    .A1(net117),
    .Y(_02646_),
    .A2(net157));
 sg13g2_nand2b_1 _08192_ (.Y(_02647_),
    .B(_02389_),
    .A_N(_02387_));
 sg13g2_nand2b_1 _08193_ (.Y(_02648_),
    .B(_02387_),
    .A_N(_02389_));
 sg13g2_a221oi_1 _08194_ (.B2(_02570_),
    .C1(_02474_),
    .B1(net122),
    .A1(_02647_),
    .Y(_02649_),
    .A2(_02648_));
 sg13g2_nand2_1 _08195_ (.Y(_02650_),
    .A(net123),
    .B(net125));
 sg13g2_nor2_1 _08196_ (.A(_02573_),
    .B(_02506_),
    .Y(_02651_));
 sg13g2_o21ai_1 _08197_ (.B1(net195),
    .Y(_02652_),
    .A1(net193),
    .A2(net164));
 sg13g2_a21oi_1 _08198_ (.A1(_02612_),
    .A2(_02586_),
    .Y(_02653_),
    .B1(net192));
 sg13g2_a21o_1 _08199_ (.A2(_02652_),
    .A1(_02651_),
    .B1(_02653_),
    .X(_02654_));
 sg13g2_nand2_1 _08200_ (.Y(_02655_),
    .A(net228),
    .B(net182));
 sg13g2_o21ai_1 _08201_ (.B1(_02655_),
    .Y(_02656_),
    .A1(net150),
    .A2(_02586_));
 sg13g2_buf_1 _08202_ (.A(net149),
    .X(_02657_));
 sg13g2_buf_1 _08203_ (.A(_02417_),
    .X(_02658_));
 sg13g2_nor4_1 _08204_ (.A(net142),
    .B(net150),
    .C(net194),
    .D(net143),
    .Y(_02659_));
 sg13g2_a221oi_1 _08205_ (.B2(net116),
    .C1(_02659_),
    .B1(_02656_),
    .A1(_02650_),
    .Y(_02660_),
    .A2(_02654_));
 sg13g2_o21ai_1 _08206_ (.B1(_02660_),
    .Y(_02661_),
    .A1(_02646_),
    .A2(_02649_));
 sg13g2_nand2_1 _08207_ (.Y(_02662_),
    .A(net151),
    .B(net184));
 sg13g2_nand2_1 _08208_ (.Y(_02663_),
    .A(net182),
    .B(net185));
 sg13g2_a22oi_1 _08209_ (.Y(_02664_),
    .B1(_02663_),
    .B2(net157),
    .A2(_02662_),
    .A1(net160));
 sg13g2_a221oi_1 _08210_ (.B2(_02500_),
    .C1(_02339_),
    .B1(_02631_),
    .A1(net245),
    .Y(_02665_),
    .A2(net258));
 sg13g2_buf_1 _08211_ (.A(_02665_),
    .X(_02666_));
 sg13g2_nand2_1 _08212_ (.Y(_02667_),
    .A(net244),
    .B(_02560_));
 sg13g2_a221oi_1 _08213_ (.B2(net184),
    .C1(_02667_),
    .B1(_02666_),
    .A1(net165),
    .Y(_02668_),
    .A2(_02374_));
 sg13g2_and2_1 _08214_ (.A(_02318_),
    .B(_02321_),
    .X(_02669_));
 sg13g2_nand4_1 _08215_ (.B(_02397_),
    .C(_02500_),
    .A(\dtop.vtop.pipeline.phases[1][6] ),
    .Y(_02670_),
    .D(_02623_));
 sg13g2_a21oi_1 _08216_ (.A1(\dtop.vtop.pipeline.phases[1][6] ),
    .A2(_02623_),
    .Y(_02671_),
    .B1(net271));
 sg13g2_a221oi_1 _08217_ (.B2(net242),
    .C1(_02671_),
    .B1(_02670_),
    .A1(net271),
    .Y(_02672_),
    .A2(_02669_));
 sg13g2_a221oi_1 _08218_ (.B2(net183),
    .C1(net148),
    .B1(_02672_),
    .A1(_02536_),
    .Y(_02673_),
    .A2(_02506_));
 sg13g2_nor3_1 _08219_ (.A(net194),
    .B(net143),
    .C(net180),
    .Y(_02674_));
 sg13g2_nor3_1 _08220_ (.A(net155),
    .B(_02673_),
    .C(_02674_),
    .Y(_02675_));
 sg13g2_nor2_1 _08221_ (.A(_02561_),
    .B(_02675_),
    .Y(_02676_));
 sg13g2_a21oi_2 _08222_ (.B1(net192),
    .Y(_02677_),
    .A2(_02612_),
    .A1(net182));
 sg13g2_o21ai_1 _08223_ (.B1(net198),
    .Y(_02678_),
    .A1(_02433_),
    .A2(_02442_));
 sg13g2_nor2_1 _08224_ (.A(net158),
    .B(_02678_),
    .Y(_02679_));
 sg13g2_a21oi_1 _08225_ (.A1(net118),
    .A2(_02677_),
    .Y(_02680_),
    .B1(_02679_));
 sg13g2_nor2_2 _08226_ (.A(_02391_),
    .B(net192),
    .Y(_02681_));
 sg13g2_nor2_2 _08227_ (.A(_02366_),
    .B(net182),
    .Y(_02682_));
 sg13g2_nor2_1 _08228_ (.A(_02417_),
    .B(_02437_),
    .Y(_02683_));
 sg13g2_a21oi_2 _08229_ (.B1(_02683_),
    .Y(_02684_),
    .A2(_02682_),
    .A1(_02681_));
 sg13g2_nand3_1 _08230_ (.B(_02680_),
    .C(_02684_),
    .A(_02577_),
    .Y(_02685_));
 sg13g2_inv_1 _08231_ (.Y(_02686_),
    .A(_02620_));
 sg13g2_inv_1 _08232_ (.Y(_02687_),
    .A(_00055_));
 sg13g2_mux4_1 _08233_ (.S0(net271),
    .A0(_02686_),
    .A1(\dtop.vtop.pipeline.phases[2][13] ),
    .A2(\dtop.vtop.pipeline.phases[1][13] ),
    .A3(_02687_),
    .S1(net269),
    .X(_02688_));
 sg13g2_buf_2 _08234_ (.A(_02688_),
    .X(_02689_));
 sg13g2_buf_1 _08235_ (.A(_02689_),
    .X(_02690_));
 sg13g2_nand2_1 _08236_ (.Y(_02691_),
    .A(net142),
    .B(net221));
 sg13g2_a221oi_1 _08237_ (.B2(_02685_),
    .C1(_02691_),
    .B1(_02676_),
    .A1(_02664_),
    .Y(_02692_),
    .A2(_02668_));
 sg13g2_or3_1 _08238_ (.A(net224),
    .B(_02661_),
    .C(_02692_),
    .X(_02693_));
 sg13g2_nand2b_1 _08239_ (.Y(_02694_),
    .B(net224),
    .A_N(_02661_));
 sg13g2_buf_1 _08240_ (.A(net150),
    .X(_02695_));
 sg13g2_nand4_1 _08241_ (.B(net115),
    .C(_02680_),
    .A(net189),
    .Y(_02696_),
    .D(_02684_));
 sg13g2_buf_1 _08242_ (.A(_02436_),
    .X(_02697_));
 sg13g2_or2_1 _08243_ (.X(_02698_),
    .B(_02697_),
    .A(_02448_));
 sg13g2_buf_1 _08244_ (.A(_02698_),
    .X(_02699_));
 sg13g2_nand2b_1 _08245_ (.Y(_02700_),
    .B(net227),
    .A_N(_02442_));
 sg13g2_nand4_1 _08246_ (.B(net229),
    .C(net230),
    .A(net190),
    .Y(_02701_),
    .D(_02539_));
 sg13g2_and2_1 _08247_ (.A(_02700_),
    .B(_02701_),
    .X(_02702_));
 sg13g2_o21ai_1 _08248_ (.B1(_02702_),
    .Y(_02703_),
    .A1(net116),
    .A2(_02699_));
 sg13g2_a21oi_1 _08249_ (.A1(_02475_),
    .A2(_02703_),
    .Y(_02704_),
    .B1(net179));
 sg13g2_o21ai_1 _08250_ (.B1(net246),
    .Y(_02705_),
    .A1(net243),
    .A2(_02669_));
 sg13g2_and2_1 _08251_ (.A(net245),
    .B(_02705_),
    .X(_02706_));
 sg13g2_buf_1 _08252_ (.A(_02706_),
    .X(_02707_));
 sg13g2_nand2_1 _08253_ (.Y(_02708_),
    .A(_02472_),
    .B(_02580_));
 sg13g2_a221oi_1 _08254_ (.B2(_02707_),
    .C1(_02708_),
    .B1(_02592_),
    .A1(net145),
    .Y(_02709_),
    .A2(net119));
 sg13g2_nor2_1 _08255_ (.A(net153),
    .B(_02689_),
    .Y(_02710_));
 sg13g2_inv_1 _08256_ (.Y(_02711_),
    .A(_02710_));
 sg13g2_a221oi_1 _08257_ (.B2(_02709_),
    .C1(_02711_),
    .B1(_02664_),
    .A1(_02696_),
    .Y(_02712_),
    .A2(_02704_));
 sg13g2_a21o_1 _08258_ (.A2(_02694_),
    .A1(_02692_),
    .B1(_02712_),
    .X(_02713_));
 sg13g2_a22oi_1 _08259_ (.Y(_02714_),
    .B1(_02693_),
    .B2(_02713_),
    .A2(_02642_),
    .A1(_02591_));
 sg13g2_buf_2 _08260_ (.A(_02714_),
    .X(_02715_));
 sg13g2_nand3_1 _08261_ (.B(net164),
    .C(net227),
    .A(net196),
    .Y(_02716_));
 sg13g2_buf_1 _08262_ (.A(net152),
    .X(_02717_));
 sg13g2_a21oi_1 _08263_ (.A1(_02434_),
    .A2(_02716_),
    .Y(_02718_),
    .B1(_02717_));
 sg13g2_a221oi_1 _08264_ (.B2(_02568_),
    .C1(_02718_),
    .B1(_02614_),
    .A1(_02426_),
    .Y(_02719_),
    .A2(_02666_));
 sg13g2_nor2_1 _08265_ (.A(net117),
    .B(_02719_),
    .Y(_02720_));
 sg13g2_buf_1 _08266_ (.A(net159),
    .X(_02721_));
 sg13g2_nor2_1 _08267_ (.A(net191),
    .B(_02373_),
    .Y(_02722_));
 sg13g2_nor2_1 _08268_ (.A(net195),
    .B(_02567_),
    .Y(_02723_));
 sg13g2_a21oi_1 _08269_ (.A1(net148),
    .A2(_02722_),
    .Y(_02724_),
    .B1(_02723_));
 sg13g2_nand2_1 _08270_ (.Y(_02725_),
    .A(net194),
    .B(_02614_));
 sg13g2_o21ai_1 _08271_ (.B1(_02725_),
    .Y(_02726_),
    .A1(net113),
    .A2(_02724_));
 sg13g2_nand2_1 _08272_ (.Y(_02727_),
    .A(net178),
    .B(_02707_));
 sg13g2_a21oi_1 _08273_ (.A1(_02412_),
    .A2(_02727_),
    .Y(_02728_),
    .B1(_02452_));
 sg13g2_a21o_1 _08274_ (.A2(_02726_),
    .A1(net117),
    .B1(_02728_),
    .X(_02729_));
 sg13g2_and3_1 _08275_ (.X(_02730_),
    .A(net196),
    .B(_02326_),
    .C(_02351_));
 sg13g2_o21ai_1 _08276_ (.B1(_02484_),
    .Y(_02731_),
    .A1(_02368_),
    .A2(_02730_));
 sg13g2_nor2_2 _08277_ (.A(_02560_),
    .B(_02689_),
    .Y(_02732_));
 sg13g2_nand2_1 _08278_ (.Y(_02733_),
    .A(_02731_),
    .B(_02732_));
 sg13g2_xnor2_1 _08279_ (.Y(_02734_),
    .A(net165),
    .B(_02574_));
 sg13g2_nand2_1 _08280_ (.Y(_02735_),
    .A(net188),
    .B(net162));
 sg13g2_nand2_1 _08281_ (.Y(_02736_),
    .A(_02560_),
    .B(_02689_));
 sg13g2_nor2_1 _08282_ (.A(_02735_),
    .B(_02736_),
    .Y(_02737_));
 sg13g2_o21ai_1 _08283_ (.B1(_02737_),
    .Y(_02738_),
    .A1(_02484_),
    .A2(_02734_));
 sg13g2_o21ai_1 _08284_ (.B1(_02738_),
    .Y(_02739_),
    .A1(_02589_),
    .A2(_02733_));
 sg13g2_o21ai_1 _08285_ (.B1(_02739_),
    .Y(_02740_),
    .A1(_02720_),
    .A2(_02729_));
 sg13g2_nand2_1 _08286_ (.Y(_02741_),
    .A(net223),
    .B(_02625_));
 sg13g2_mux2_1 _08287_ (.A0(_02741_),
    .A1(_02736_),
    .S(net159),
    .X(_02742_));
 sg13g2_nor2_1 _08288_ (.A(_02473_),
    .B(net162),
    .Y(_02743_));
 sg13g2_a21o_1 _08289_ (.A2(_02570_),
    .A1(_02448_),
    .B1(_02332_),
    .X(_02744_));
 sg13g2_nand2_1 _08290_ (.Y(_02745_),
    .A(net228),
    .B(_02528_));
 sg13g2_a22oi_1 _08291_ (.Y(_02746_),
    .B1(_02745_),
    .B2(_02373_),
    .A2(_02744_),
    .A1(net182));
 sg13g2_nor2_1 _08292_ (.A(_02735_),
    .B(_02746_),
    .Y(_02747_));
 sg13g2_a21oi_1 _08293_ (.A1(_02743_),
    .A2(_02746_),
    .Y(_02748_),
    .B1(_02747_));
 sg13g2_nor2_1 _08294_ (.A(net193),
    .B(net187),
    .Y(_02749_));
 sg13g2_nand2_1 _08295_ (.Y(_02750_),
    .A(net124),
    .B(_02749_));
 sg13g2_a22oi_1 _08296_ (.Y(_02751_),
    .B1(net245),
    .B2(net258),
    .A2(_02594_),
    .A1(_02593_));
 sg13g2_buf_1 _08297_ (.A(_02751_),
    .X(_02752_));
 sg13g2_nand2_1 _08298_ (.Y(_02753_),
    .A(net142),
    .B(_02752_));
 sg13g2_a21oi_1 _08299_ (.A1(_02750_),
    .A2(_02753_),
    .Y(_02754_),
    .B1(_02684_));
 sg13g2_nor2_1 _08300_ (.A(_02748_),
    .B(_02754_),
    .Y(_02755_));
 sg13g2_xnor2_1 _08301_ (.Y(_02756_),
    .A(net191),
    .B(net180));
 sg13g2_nand2_1 _08302_ (.Y(_02757_),
    .A(_02409_),
    .B(net197));
 sg13g2_nand3_1 _08303_ (.B(_02481_),
    .C(_02757_),
    .A(net187),
    .Y(_02758_));
 sg13g2_o21ai_1 _08304_ (.B1(_02758_),
    .Y(_02759_),
    .A1(_02479_),
    .A2(_02756_));
 sg13g2_a21o_1 _08305_ (.A2(_02598_),
    .A1(_02370_),
    .B1(_02605_),
    .X(_02760_));
 sg13g2_nand2_1 _08306_ (.Y(_02761_),
    .A(net190),
    .B(net198));
 sg13g2_nand2_1 _08307_ (.Y(_02762_),
    .A(_02757_),
    .B(_02761_));
 sg13g2_a221oi_1 _08308_ (.B2(_02414_),
    .C1(net194),
    .B1(_02762_),
    .A1(_02479_),
    .Y(_02763_),
    .A2(_02760_));
 sg13g2_a21oi_1 _08309_ (.A1(net151),
    .A2(_02759_),
    .Y(_02764_),
    .B1(_02763_));
 sg13g2_nor2_1 _08310_ (.A(_02645_),
    .B(_02764_),
    .Y(_02765_));
 sg13g2_nand2_2 _08311_ (.Y(_02766_),
    .A(_02409_),
    .B(net198));
 sg13g2_a221oi_1 _08312_ (.B2(net196),
    .C1(net164),
    .B1(_02766_),
    .A1(net193),
    .Y(_02767_),
    .A2(_02514_));
 sg13g2_nor3_1 _08313_ (.A(net154),
    .B(_02480_),
    .C(_02526_),
    .Y(_02768_));
 sg13g2_nor3_1 _08314_ (.A(_02517_),
    .B(_02767_),
    .C(_02768_),
    .Y(_02769_));
 sg13g2_a21o_1 _08315_ (.A2(_02605_),
    .A1(_02425_),
    .B1(_02599_),
    .X(_02770_));
 sg13g2_a22oi_1 _08316_ (.Y(_02771_),
    .B1(_02770_),
    .B2(net126),
    .A2(_02762_),
    .A1(_02722_));
 sg13g2_nor2_1 _08317_ (.A(net146),
    .B(_02771_),
    .Y(_02772_));
 sg13g2_nor4_1 _08318_ (.A(net121),
    .B(net98),
    .C(_02769_),
    .D(_02772_),
    .Y(_02773_));
 sg13g2_or4_1 _08319_ (.A(_02742_),
    .B(_02755_),
    .C(_02765_),
    .D(_02773_),
    .X(_02774_));
 sg13g2_nand4_1 _08320_ (.B(net241),
    .C(_02429_),
    .A(net242),
    .Y(_02775_),
    .D(_02431_));
 sg13g2_buf_1 _08321_ (.A(_02775_),
    .X(_02776_));
 sg13g2_a22oi_1 _08322_ (.Y(_02777_),
    .B1(_02429_),
    .B2(_02431_),
    .A2(_02594_),
    .A1(_02396_));
 sg13g2_buf_2 _08323_ (.A(_02777_),
    .X(_02778_));
 sg13g2_a221oi_1 _08324_ (.B2(_02538_),
    .C1(net154),
    .B1(_02778_),
    .A1(net148),
    .Y(_02779_),
    .A2(_02514_));
 sg13g2_o21ai_1 _08325_ (.B1(_02779_),
    .Y(_02780_),
    .A1(_02543_),
    .A2(_02776_));
 sg13g2_nand4_1 _08326_ (.B(net256),
    .C(_02429_),
    .A(net257),
    .Y(_02781_),
    .D(_02431_));
 sg13g2_buf_1 _08327_ (.A(_02781_),
    .X(_02782_));
 sg13g2_nor2_1 _08328_ (.A(net178),
    .B(_02603_),
    .Y(_02783_));
 sg13g2_o21ai_1 _08329_ (.B1(_02783_),
    .Y(_02784_),
    .A1(net122),
    .A2(_02782_));
 sg13g2_nor2_1 _08330_ (.A(net124),
    .B(_02708_),
    .Y(_02785_));
 sg13g2_nand3_1 _08331_ (.B(_02784_),
    .C(_02785_),
    .A(_02780_),
    .Y(_02786_));
 sg13g2_nand2_1 _08332_ (.Y(_02787_),
    .A(net222),
    .B(_02786_));
 sg13g2_o21ai_1 _08333_ (.B1(net186),
    .Y(_02788_),
    .A1(_02506_),
    .A2(net185));
 sg13g2_a22oi_1 _08334_ (.Y(_02789_),
    .B1(_02778_),
    .B2(_02480_),
    .A2(net144),
    .A1(net178));
 sg13g2_nand3_1 _08335_ (.B(_02788_),
    .C(_02789_),
    .A(_02533_),
    .Y(_02790_));
 sg13g2_nand3_1 _08336_ (.B(net196),
    .C(net181),
    .A(net156),
    .Y(_02791_));
 sg13g2_nand4_1 _08337_ (.B(_02766_),
    .C(_02782_),
    .A(net126),
    .Y(_02792_),
    .D(_02791_));
 sg13g2_nand4_1 _08338_ (.B(_02639_),
    .C(_02790_),
    .A(net97),
    .Y(_02793_),
    .D(_02792_));
 sg13g2_nand2_1 _08339_ (.Y(_02794_),
    .A(net221),
    .B(_02793_));
 sg13g2_xnor2_1 _08340_ (.Y(_02795_),
    .A(net188),
    .B(_02417_));
 sg13g2_buf_2 _08341_ (.A(_02795_),
    .X(_02796_));
 sg13g2_o21ai_1 _08342_ (.B1(_02586_),
    .Y(_02797_),
    .A1(net163),
    .A2(_02666_));
 sg13g2_xnor2_1 _08343_ (.Y(_02798_),
    .A(net183),
    .B(_02797_));
 sg13g2_o21ai_1 _08344_ (.B1(net150),
    .Y(_02799_),
    .A1(net195),
    .A2(net154));
 sg13g2_a21oi_1 _08345_ (.A1(net195),
    .A2(net187),
    .Y(_02800_),
    .B1(net156));
 sg13g2_nor2_1 _08346_ (.A(net225),
    .B(_02800_),
    .Y(_02801_));
 sg13g2_a22oi_1 _08347_ (.Y(_02802_),
    .B1(_02801_),
    .B2(_02717_),
    .A2(_02799_),
    .A1(_02743_));
 sg13g2_o21ai_1 _08348_ (.B1(_02802_),
    .Y(_02803_),
    .A1(_02796_),
    .A2(_02798_));
 sg13g2_a221oi_1 _08349_ (.B2(net160),
    .C1(net161),
    .B1(net148),
    .A1(_02647_),
    .Y(_02804_),
    .A2(_02648_));
 sg13g2_a221oi_1 _08350_ (.B2(net157),
    .C1(net124),
    .B1(net194),
    .A1(net242),
    .Y(_02805_),
    .A2(net241));
 sg13g2_a22oi_1 _08351_ (.Y(_02806_),
    .B1(_02514_),
    .B2(_02486_),
    .A2(_02506_),
    .A1(_02586_));
 sg13g2_o21ai_1 _08352_ (.B1(_02806_),
    .Y(_02807_),
    .A1(_02804_),
    .A2(_02805_));
 sg13g2_a21oi_1 _08353_ (.A1(net155),
    .A2(net165),
    .Y(_02808_),
    .B1(_02618_));
 sg13g2_nand3_1 _08354_ (.B(_02628_),
    .C(_02808_),
    .A(_02546_),
    .Y(_02809_));
 sg13g2_nand2_1 _08355_ (.Y(_02810_),
    .A(net189),
    .B(net145));
 sg13g2_nand4_1 _08356_ (.B(_02618_),
    .C(_02690_),
    .A(_02549_),
    .Y(_02811_),
    .D(_02810_));
 sg13g2_a22oi_1 _08357_ (.Y(_02812_),
    .B1(_02809_),
    .B2(_02811_),
    .A2(_02807_),
    .A1(_02803_));
 sg13g2_a21oi_1 _08358_ (.A1(_02787_),
    .A2(_02794_),
    .Y(_02813_),
    .B1(_02812_));
 sg13g2_a22oi_1 _08359_ (.Y(_02814_),
    .B1(_02495_),
    .B2(net195),
    .A2(_02570_),
    .A1(net164));
 sg13g2_nor2_1 _08360_ (.A(net123),
    .B(_02814_),
    .Y(_02815_));
 sg13g2_a221oi_1 _08361_ (.B2(net113),
    .C1(_02815_),
    .B1(_02614_),
    .A1(net117),
    .Y(_02816_),
    .A2(net178));
 sg13g2_nand2_1 _08362_ (.Y(_02817_),
    .A(_02589_),
    .B(_02735_));
 sg13g2_o21ai_1 _08363_ (.B1(_02817_),
    .Y(_02818_),
    .A1(_02695_),
    .A2(_02816_));
 sg13g2_a21oi_1 _08364_ (.A1(net153),
    .A2(_02480_),
    .Y(_02819_),
    .B1(_02570_));
 sg13g2_nand2_1 _08365_ (.Y(_02820_),
    .A(net193),
    .B(net191));
 sg13g2_o21ai_1 _08366_ (.B1(_02820_),
    .Y(_02821_),
    .A1(_02533_),
    .A2(_02819_));
 sg13g2_nand2_1 _08367_ (.Y(_02822_),
    .A(net113),
    .B(net147));
 sg13g2_a22oi_1 _08368_ (.Y(_02823_),
    .B1(_02603_),
    .B2(_02822_),
    .A2(net146),
    .A1(_02326_));
 sg13g2_a21oi_1 _08369_ (.A1(net227),
    .A2(_02506_),
    .Y(_02824_),
    .B1(net193));
 sg13g2_and2_1 _08370_ (.A(net142),
    .B(_02824_),
    .X(_02825_));
 sg13g2_a221oi_1 _08371_ (.B2(_02722_),
    .C1(net123),
    .B1(_02592_),
    .A1(net126),
    .Y(_02826_),
    .A2(net143));
 sg13g2_o21ai_1 _08372_ (.B1(_02766_),
    .Y(_02827_),
    .A1(_02825_),
    .A2(_02826_));
 sg13g2_a221oi_1 _08373_ (.B2(_02372_),
    .C1(_02827_),
    .B1(_02823_),
    .A1(net146),
    .Y(_02828_),
    .A2(_02821_));
 sg13g2_nor3_1 _08374_ (.A(net118),
    .B(net224),
    .C(net222),
    .Y(_02829_));
 sg13g2_a21oi_1 _08375_ (.A1(_02582_),
    .A2(_02628_),
    .Y(_02830_),
    .B1(_02829_));
 sg13g2_nand2b_1 _08376_ (.Y(_02831_),
    .B(_02716_),
    .A_N(_02592_));
 sg13g2_nand2_1 _08377_ (.Y(_02832_),
    .A(net122),
    .B(_02481_));
 sg13g2_nand2_1 _08378_ (.Y(_02833_),
    .A(_02433_),
    .B(_02442_));
 sg13g2_nand3_1 _08379_ (.B(_02782_),
    .C(_02833_),
    .A(net161),
    .Y(_02834_));
 sg13g2_a221oi_1 _08380_ (.B2(_02834_),
    .C1(_02645_),
    .B1(_02832_),
    .A1(_02564_),
    .Y(_02835_),
    .A2(_02831_));
 sg13g2_nor3_1 _08381_ (.A(_02409_),
    .B(net229),
    .C(_02325_),
    .Y(_02836_));
 sg13g2_o21ai_1 _08382_ (.B1(_02376_),
    .Y(_02837_),
    .A1(_02529_),
    .A2(_02836_));
 sg13g2_nand2_1 _08383_ (.Y(_02838_),
    .A(net197),
    .B(net230));
 sg13g2_nand2_1 _08384_ (.Y(_02839_),
    .A(net195),
    .B(_02838_));
 sg13g2_a221oi_1 _08385_ (.B2(_02592_),
    .C1(net123),
    .B1(_02839_),
    .A1(net183),
    .Y(_02840_),
    .A2(_02529_));
 sg13g2_and3_1 _08386_ (.X(_02841_),
    .A(net189),
    .B(_02837_),
    .C(_02840_));
 sg13g2_nor3_1 _08387_ (.A(_02830_),
    .B(_02835_),
    .C(_02841_),
    .Y(_02842_));
 sg13g2_o21ai_1 _08388_ (.B1(_02842_),
    .Y(_02843_),
    .A1(_02818_),
    .A2(_02828_));
 sg13g2_and4_1 _08389_ (.A(_02740_),
    .B(_02774_),
    .C(_02813_),
    .D(_02843_),
    .X(_02844_));
 sg13g2_buf_1 _08390_ (.A(_02844_),
    .X(_02845_));
 sg13g2_inv_1 _08391_ (.Y(_02846_),
    .A(_02249_));
 sg13g2_nor2_1 _08392_ (.A(_02846_),
    .B(_02251_),
    .Y(_02847_));
 sg13g2_nor3_1 _08393_ (.A(net399),
    .B(_05136_),
    .C(_01193_),
    .Y(_02848_));
 sg13g2_or2_1 _08394_ (.X(_02849_),
    .B(_02848_),
    .A(_05265_));
 sg13g2_buf_1 _08395_ (.A(_02849_),
    .X(_02850_));
 sg13g2_nor2_1 _08396_ (.A(_02264_),
    .B(_02847_),
    .Y(_02851_));
 sg13g2_a21oi_1 _08397_ (.A1(_02847_),
    .A2(_02850_),
    .Y(_02852_),
    .B1(_02851_));
 sg13g2_nor2_1 _08398_ (.A(net289),
    .B(_02852_),
    .Y(_02853_));
 sg13g2_a21o_1 _08399_ (.A2(net277),
    .A1(net286),
    .B1(_02853_),
    .X(_02854_));
 sg13g2_buf_1 _08400_ (.A(_02854_),
    .X(_02855_));
 sg13g2_buf_1 _08401_ (.A(net240),
    .X(_02856_));
 sg13g2_mux2_1 _08402_ (.A0(_02715_),
    .A1(_02845_),
    .S(net220),
    .X(_02857_));
 sg13g2_xnor2_1 _08403_ (.Y(_02858_),
    .A(net166),
    .B(_02857_));
 sg13g2_nor2_1 _08404_ (.A(net248),
    .B(_02858_),
    .Y(_02859_));
 sg13g2_nor2b_1 _08405_ (.A(_05405_),
    .B_N(_01450_),
    .Y(_02860_));
 sg13g2_buf_2 _08406_ (.A(_02860_),
    .X(_02861_));
 sg13g2_mux2_1 _08407_ (.A0(\dtop.vtop.dphases[0][0] ),
    .A1(_02859_),
    .S(_02861_),
    .X(_00174_));
 sg13g2_buf_1 _08408_ (.A(net277),
    .X(_02862_));
 sg13g2_nand3_1 _08409_ (.B(_02862_),
    .C(_01450_),
    .A(net426),
    .Y(_02863_));
 sg13g2_buf_1 _08410_ (.A(_02863_),
    .X(_02864_));
 sg13g2_nand2_1 _08411_ (.Y(_02865_),
    .A(\dtop.vtop.dphases[0][10] ),
    .B(net239));
 sg13g2_o21ai_1 _08412_ (.B1(_02865_),
    .Y(_00175_),
    .A1(net247),
    .A2(net239));
 sg13g2_a21oi_1 _08413_ (.A1(net286),
    .A2(net277),
    .Y(_02866_),
    .B1(_02853_));
 sg13g2_buf_2 _08414_ (.A(_02866_),
    .X(_02867_));
 sg13g2_a21o_1 _08415_ (.A2(net277),
    .A1(net394),
    .B1(_02252_),
    .X(_02868_));
 sg13g2_buf_1 _08416_ (.A(_02868_),
    .X(_02869_));
 sg13g2_buf_1 _08417_ (.A(_02869_),
    .X(_02870_));
 sg13g2_buf_1 _08418_ (.A(net219),
    .X(_02871_));
 sg13g2_nor2_1 _08419_ (.A(net158),
    .B(net183),
    .Y(_02872_));
 sg13g2_nor2_2 _08420_ (.A(_02410_),
    .B(net182),
    .Y(_02873_));
 sg13g2_and2_1 _08421_ (.A(_02442_),
    .B(_02778_),
    .X(_02874_));
 sg13g2_buf_1 _08422_ (.A(_02874_),
    .X(_02875_));
 sg13g2_nor2_1 _08423_ (.A(_02873_),
    .B(_02875_),
    .Y(_02876_));
 sg13g2_o21ai_1 _08424_ (.B1(net142),
    .Y(_02877_),
    .A1(_02873_),
    .A2(_02875_));
 sg13g2_nor2_1 _08425_ (.A(_02592_),
    .B(_02633_),
    .Y(_02878_));
 sg13g2_a221oi_1 _08426_ (.B2(_02878_),
    .C1(_02564_),
    .B1(_02877_),
    .A1(_02872_),
    .Y(_02879_),
    .A2(_02876_));
 sg13g2_nor2_1 _08427_ (.A(net230),
    .B(_02776_),
    .Y(_02880_));
 sg13g2_nor2_1 _08428_ (.A(_02778_),
    .B(_02880_),
    .Y(_02881_));
 sg13g2_a221oi_1 _08429_ (.B2(_02426_),
    .C1(net116),
    .B1(_02881_),
    .A1(net113),
    .Y(_02882_),
    .A2(_02878_));
 sg13g2_nand3_1 _08430_ (.B(net186),
    .C(net185),
    .A(net145),
    .Y(_02883_));
 sg13g2_nand4_1 _08431_ (.B(net114),
    .C(net179),
    .A(net189),
    .Y(_02884_),
    .D(_02883_));
 sg13g2_o21ai_1 _08432_ (.B1(_02884_),
    .Y(_02885_),
    .A1(net179),
    .A2(_02645_));
 sg13g2_o21ai_1 _08433_ (.B1(_02885_),
    .Y(_02886_),
    .A1(_02879_),
    .A2(_02882_));
 sg13g2_a21oi_1 _08434_ (.A1(_02376_),
    .A2(_02745_),
    .Y(_02887_),
    .B1(net160));
 sg13g2_nor2_1 _08435_ (.A(_02460_),
    .B(_02560_),
    .Y(_02888_));
 sg13g2_buf_2 _08436_ (.A(_02888_),
    .X(_02889_));
 sg13g2_nand2_1 _08437_ (.Y(_02890_),
    .A(net124),
    .B(_02889_));
 sg13g2_o21ai_1 _08438_ (.B1(_02890_),
    .Y(_02891_),
    .A1(_02640_),
    .A2(_02887_));
 sg13g2_nand2_1 _08439_ (.Y(_02892_),
    .A(net190),
    .B(_02367_));
 sg13g2_nor2b_1 _08440_ (.A(_02892_),
    .B_N(_02707_),
    .Y(_02893_));
 sg13g2_nand2_1 _08441_ (.Y(_02894_),
    .A(net227),
    .B(_02421_));
 sg13g2_o21ai_1 _08442_ (.B1(_02894_),
    .Y(_02895_),
    .A1(net153),
    .A2(_02700_));
 sg13g2_a221oi_1 _08443_ (.B2(net118),
    .C1(_02895_),
    .B1(_02893_),
    .A1(net146),
    .Y(_02896_),
    .A2(net157));
 sg13g2_nor2_1 _08444_ (.A(_02472_),
    .B(_02560_),
    .Y(_02897_));
 sg13g2_nor2_1 _08445_ (.A(net244),
    .B(_02580_),
    .Y(_02898_));
 sg13g2_mux2_1 _08446_ (.A0(_02897_),
    .A1(_02898_),
    .S(_02391_),
    .X(_02899_));
 sg13g2_buf_2 _08447_ (.A(_02899_),
    .X(_02900_));
 sg13g2_a22oi_1 _08448_ (.Y(_02901_),
    .B1(_02672_),
    .B2(_02682_),
    .A2(_02701_),
    .A1(net152));
 sg13g2_xnor2_1 _08449_ (.Y(_02902_),
    .A(net125),
    .B(_02901_));
 sg13g2_nand3_1 _08450_ (.B(_02639_),
    .C(_02677_),
    .A(net122),
    .Y(_02903_));
 sg13g2_nand3_1 _08451_ (.B(_02700_),
    .C(_02889_),
    .A(net144),
    .Y(_02904_));
 sg13g2_nor2_1 _08452_ (.A(net158),
    .B(net222),
    .Y(_02905_));
 sg13g2_a22oi_1 _08453_ (.Y(_02906_),
    .B1(_02904_),
    .B2(_02905_),
    .A2(_02903_),
    .A1(_02710_));
 sg13g2_a221oi_1 _08454_ (.B2(_02902_),
    .C1(_02906_),
    .B1(_02900_),
    .A1(_02891_),
    .Y(_02907_),
    .A2(_02896_));
 sg13g2_nand2_1 _08455_ (.Y(_02908_),
    .A(_02886_),
    .B(_02907_));
 sg13g2_a22oi_1 _08456_ (.Y(_02909_),
    .B1(_02330_),
    .B2(net258),
    .A2(_02327_),
    .A1(_02491_));
 sg13g2_o21ai_1 _08457_ (.B1(_02371_),
    .Y(_02910_),
    .A1(net163),
    .A2(_02752_));
 sg13g2_o21ai_1 _08458_ (.B1(_02672_),
    .Y(_02911_),
    .A1(net163),
    .A2(net182));
 sg13g2_nand3_1 _08459_ (.B(_02910_),
    .C(_02911_),
    .A(_02440_),
    .Y(_02912_));
 sg13g2_o21ai_1 _08460_ (.B1(_02367_),
    .Y(_02913_),
    .A1(net192),
    .A2(_02752_));
 sg13g2_nand2_1 _08461_ (.Y(_02914_),
    .A(net142),
    .B(_02913_));
 sg13g2_nand2_1 _08462_ (.Y(_02915_),
    .A(_02377_),
    .B(net182));
 sg13g2_a21oi_1 _08463_ (.A1(net150),
    .A2(net154),
    .Y(_02916_),
    .B1(_02915_));
 sg13g2_a221oi_1 _08464_ (.B2(_02914_),
    .C1(_02916_),
    .B1(_02912_),
    .A1(_02909_),
    .Y(_02917_),
    .A2(_02517_));
 sg13g2_nand3b_1 _08465_ (.B(net142),
    .C(_02326_),
    .Y(_02918_),
    .A_N(_02414_));
 sg13g2_a21oi_1 _08466_ (.A1(_02440_),
    .A2(net143),
    .Y(_02919_),
    .B1(net161));
 sg13g2_o21ai_1 _08467_ (.B1(_02378_),
    .Y(_02920_),
    .A1(net158),
    .A2(net126));
 sg13g2_a22oi_1 _08468_ (.Y(_02921_),
    .B1(_02920_),
    .B2(_02873_),
    .A2(_02919_),
    .A1(_02918_));
 sg13g2_mux2_1 _08469_ (.A0(net149),
    .A1(net185),
    .S(_02375_),
    .X(_02922_));
 sg13g2_nand3_1 _08470_ (.B(net145),
    .C(_02922_),
    .A(_02721_),
    .Y(_02923_));
 sg13g2_mux2_1 _08471_ (.A0(_02423_),
    .A1(_02778_),
    .S(_02377_),
    .X(_02924_));
 sg13g2_nand3_1 _08472_ (.B(net183),
    .C(_02924_),
    .A(_02548_),
    .Y(_02925_));
 sg13g2_nand3_1 _08473_ (.B(_02923_),
    .C(_02925_),
    .A(_02900_),
    .Y(_02926_));
 sg13g2_a21o_1 _08474_ (.A2(_02921_),
    .A1(_02917_),
    .B1(_02926_),
    .X(_02927_));
 sg13g2_nor2_1 _08475_ (.A(net162),
    .B(_02689_),
    .Y(_02928_));
 sg13g2_xnor2_1 _08476_ (.Y(_02929_),
    .A(net190),
    .B(_02909_));
 sg13g2_a22oi_1 _08477_ (.Y(_02930_),
    .B1(_02929_),
    .B2(_02723_),
    .A2(_02770_),
    .A1(_02540_));
 sg13g2_nor2_1 _08478_ (.A(net187),
    .B(_02596_),
    .Y(_02931_));
 sg13g2_o21ai_1 _08479_ (.B1(_02537_),
    .Y(_02932_),
    .A1(_02634_),
    .A2(_02931_));
 sg13g2_nand4_1 _08480_ (.B(_02327_),
    .C(_02330_),
    .A(_02491_),
    .Y(_02933_),
    .D(_02323_));
 sg13g2_a21o_1 _08481_ (.A2(_02933_),
    .A1(_02411_),
    .B1(_02655_),
    .X(_02934_));
 sg13g2_nand4_1 _08482_ (.B(_02930_),
    .C(_02932_),
    .A(_02889_),
    .Y(_02935_),
    .D(_02934_));
 sg13g2_o21ai_1 _08483_ (.B1(_02423_),
    .Y(_02936_),
    .A1(_02410_),
    .A2(_02909_));
 sg13g2_a22oi_1 _08484_ (.Y(_02937_),
    .B1(_02605_),
    .B2(_02478_),
    .A2(_02599_),
    .A1(net181));
 sg13g2_a21o_1 _08485_ (.A2(_02937_),
    .A1(_02936_),
    .B1(_02537_),
    .X(_02938_));
 sg13g2_xnor2_1 _08486_ (.Y(_02939_),
    .A(net190),
    .B(_02933_));
 sg13g2_nor2_1 _08487_ (.A(net196),
    .B(net226),
    .Y(_02940_));
 sg13g2_a221oi_1 _08488_ (.B2(_02940_),
    .C1(_02667_),
    .B1(_02939_),
    .A1(net186),
    .Y(_02941_),
    .A2(_02760_));
 sg13g2_nand2_1 _08489_ (.Y(_02942_),
    .A(net124),
    .B(_02690_));
 sg13g2_a21oi_1 _08490_ (.A1(_02938_),
    .A2(_02941_),
    .Y(_02943_),
    .B1(_02942_));
 sg13g2_a21o_1 _08491_ (.A2(_02935_),
    .A1(_02928_),
    .B1(_02943_),
    .X(_02944_));
 sg13g2_mux2_1 _08492_ (.A0(_02378_),
    .A1(_02915_),
    .S(net152),
    .X(_02945_));
 sg13g2_a22oi_1 _08493_ (.Y(_02946_),
    .B1(net180),
    .B2(net164),
    .A2(_02586_),
    .A1(_02419_));
 sg13g2_a21oi_1 _08494_ (.A1(_02666_),
    .A2(net184),
    .Y(_02947_),
    .B1(_02573_));
 sg13g2_mux2_1 _08495_ (.A0(_02946_),
    .A1(_02947_),
    .S(_02658_),
    .X(_02948_));
 sg13g2_o21ai_1 _08496_ (.B1(_02948_),
    .Y(_02949_),
    .A1(_02752_),
    .A2(_02945_));
 sg13g2_xnor2_1 _08497_ (.Y(_02950_),
    .A(net159),
    .B(net223));
 sg13g2_nor3_1 _08498_ (.A(net165),
    .B(_02796_),
    .C(_02950_),
    .Y(_02951_));
 sg13g2_nor2_1 _08499_ (.A(net153),
    .B(_02516_),
    .Y(_02952_));
 sg13g2_a21oi_1 _08500_ (.A1(net156),
    .A2(net181),
    .Y(_02953_),
    .B1(net164));
 sg13g2_o21ai_1 _08501_ (.B1(_02446_),
    .Y(_02954_),
    .A1(_02633_),
    .A2(_02953_));
 sg13g2_a21oi_1 _08502_ (.A1(net158),
    .A2(_02749_),
    .Y(_02955_),
    .B1(net125));
 sg13g2_and2_1 _08503_ (.A(net187),
    .B(_02493_),
    .X(_02956_));
 sg13g2_mux2_1 _08504_ (.A0(_02495_),
    .A1(_02956_),
    .S(_02485_),
    .X(_02957_));
 sg13g2_a221oi_1 _08505_ (.B2(_02955_),
    .C1(_02957_),
    .B1(_02954_),
    .A1(_02952_),
    .Y(_02958_),
    .A2(_02931_));
 sg13g2_nor3_1 _08506_ (.A(_02602_),
    .B(_02796_),
    .C(_02950_),
    .Y(_02959_));
 sg13g2_a22oi_1 _08507_ (.Y(_02960_),
    .B1(_02958_),
    .B2(_02959_),
    .A2(_02951_),
    .A1(_02949_));
 sg13g2_xnor2_1 _08508_ (.Y(_02961_),
    .A(_02391_),
    .B(_02580_));
 sg13g2_buf_2 _08509_ (.A(_02961_),
    .X(_02962_));
 sg13g2_a21oi_1 _08510_ (.A1(_02602_),
    .A2(_02586_),
    .Y(_02963_),
    .B1(_02666_));
 sg13g2_xnor2_1 _08511_ (.Y(_02964_),
    .A(_02657_),
    .B(_02963_));
 sg13g2_nand3_1 _08512_ (.B(_02962_),
    .C(_02964_),
    .A(_02796_),
    .Y(_02965_));
 sg13g2_nand4_1 _08513_ (.B(_02944_),
    .C(_02960_),
    .A(_02927_),
    .Y(_02966_),
    .D(_02965_));
 sg13g2_and2_1 _08514_ (.A(_02908_),
    .B(_02966_),
    .X(_02967_));
 sg13g2_buf_1 _08515_ (.A(_02967_),
    .X(_02968_));
 sg13g2_nand2_1 _08516_ (.Y(_02969_),
    .A(net177),
    .B(_02968_));
 sg13g2_o21ai_1 _08517_ (.B1(_02969_),
    .Y(_02970_),
    .A1(net177),
    .A2(_02845_));
 sg13g2_xnor2_1 _08518_ (.Y(_02971_),
    .A(_02287_),
    .B(_02970_));
 sg13g2_xnor2_1 _08519_ (.Y(_02972_),
    .A(net166),
    .B(_02715_));
 sg13g2_nor3_1 _08520_ (.A(_02254_),
    .B(_02867_),
    .C(_02972_),
    .Y(_02973_));
 sg13g2_a21o_1 _08521_ (.A2(_02971_),
    .A1(_02867_),
    .B1(_02973_),
    .X(_02974_));
 sg13g2_mux2_1 _08522_ (.A0(\dtop.vtop.dphases[0][1] ),
    .A1(_02974_),
    .S(_02861_),
    .X(_00176_));
 sg13g2_nand3_1 _08523_ (.B(_02796_),
    .C(_02962_),
    .A(net120),
    .Y(_02975_));
 sg13g2_nand3_1 _08524_ (.B(_02796_),
    .C(_02962_),
    .A(net122),
    .Y(_02976_));
 sg13g2_or2_1 _08525_ (.X(_02977_),
    .B(_02442_),
    .A(net197));
 sg13g2_mux2_1 _08526_ (.A0(_02838_),
    .A1(_02977_),
    .S(_02391_),
    .X(_02978_));
 sg13g2_nor4_1 _08527_ (.A(net196),
    .B(net163),
    .C(net187),
    .D(net181),
    .Y(_02979_));
 sg13g2_nor4_1 _08528_ (.A(net162),
    .B(net147),
    .C(_02422_),
    .D(_02697_),
    .Y(_02980_));
 sg13g2_a221oi_1 _08529_ (.B2(_02393_),
    .C1(_02980_),
    .B1(_02979_),
    .A1(net146),
    .Y(_02981_),
    .A2(_02978_));
 sg13g2_mux2_1 _08530_ (.A0(_02975_),
    .A1(_02976_),
    .S(_02981_),
    .X(_02982_));
 sg13g2_and2_1 _08531_ (.A(net191),
    .B(_02778_),
    .X(_02983_));
 sg13g2_o21ai_1 _08532_ (.B1(net149),
    .Y(_02984_),
    .A1(_02836_),
    .A2(_02983_));
 sg13g2_and2_1 _08533_ (.A(net153),
    .B(_02663_),
    .X(_02985_));
 sg13g2_a21o_1 _08534_ (.A2(net185),
    .A1(net228),
    .B1(net184),
    .X(_02986_));
 sg13g2_a221oi_1 _08535_ (.B2(_02516_),
    .C1(net153),
    .B1(_02986_),
    .A1(net157),
    .Y(_02987_),
    .A2(_02606_));
 sg13g2_a21o_1 _08536_ (.A2(_02985_),
    .A1(_02984_),
    .B1(_02987_),
    .X(_02988_));
 sg13g2_nand2_1 _08537_ (.Y(_02989_),
    .A(_02658_),
    .B(_02897_));
 sg13g2_nand2_1 _08538_ (.Y(_02990_),
    .A(_02393_),
    .B(_02898_));
 sg13g2_a21oi_1 _08539_ (.A1(net183),
    .A2(net185),
    .Y(_02991_),
    .B1(_02531_));
 sg13g2_nor2_1 _08540_ (.A(_02567_),
    .B(net184),
    .Y(_02992_));
 sg13g2_nor2_1 _08541_ (.A(net226),
    .B(net185),
    .Y(_02993_));
 sg13g2_mux2_1 _08542_ (.A0(_02992_),
    .A1(_02993_),
    .S(_02488_),
    .X(_02994_));
 sg13g2_a22oi_1 _08543_ (.Y(_02995_),
    .B1(_02991_),
    .B2(_02994_),
    .A2(_02990_),
    .A1(_02989_));
 sg13g2_nor3_1 _08544_ (.A(net244),
    .B(net226),
    .C(_02606_),
    .Y(_02996_));
 sg13g2_o21ai_1 _08545_ (.B1(_02996_),
    .Y(_02997_),
    .A1(_02411_),
    .A2(_02565_));
 sg13g2_nand3_1 _08546_ (.B(net194),
    .C(_02639_),
    .A(_02446_),
    .Y(_02998_));
 sg13g2_o21ai_1 _08547_ (.B1(_02998_),
    .Y(_02999_),
    .A1(_02610_),
    .A2(_02997_));
 sg13g2_nand2_1 _08548_ (.Y(_03000_),
    .A(net150),
    .B(_02613_));
 sg13g2_o21ai_1 _08549_ (.B1(_03000_),
    .Y(_03001_),
    .A1(net158),
    .A2(_02613_));
 sg13g2_a22oi_1 _08550_ (.Y(_03002_),
    .B1(_03001_),
    .B2(_02657_),
    .A2(net144),
    .A1(_02565_));
 sg13g2_a22oi_1 _08551_ (.Y(_03003_),
    .B1(_02999_),
    .B2(_03002_),
    .A2(_02995_),
    .A1(_02988_));
 sg13g2_a21o_1 _08552_ (.A2(_02598_),
    .A1(_02425_),
    .B1(_02605_),
    .X(_03004_));
 sg13g2_nand3_1 _08553_ (.B(_02639_),
    .C(_03004_),
    .A(net148),
    .Y(_03005_));
 sg13g2_nor3_1 _08554_ (.A(net188),
    .B(net191),
    .C(_02581_),
    .Y(_03006_));
 sg13g2_o21ai_1 _08555_ (.B1(_03006_),
    .Y(_03007_),
    .A1(_02778_),
    .A2(_02880_));
 sg13g2_nand3_1 _08556_ (.B(_03005_),
    .C(_03007_),
    .A(_02928_),
    .Y(_03008_));
 sg13g2_xnor2_1 _08557_ (.Y(_03009_),
    .A(net193),
    .B(_02514_));
 sg13g2_nand3_1 _08558_ (.B(_02889_),
    .C(_03009_),
    .A(net186),
    .Y(_03010_));
 sg13g2_nand2_1 _08559_ (.Y(_03011_),
    .A(_02889_),
    .B(_02875_));
 sg13g2_nand3_1 _08560_ (.B(_03010_),
    .C(_03011_),
    .A(_02626_),
    .Y(_03012_));
 sg13g2_nor3_1 _08561_ (.A(net149),
    .B(_02443_),
    .C(_02776_),
    .Y(_03013_));
 sg13g2_a21oi_1 _08562_ (.A1(_02563_),
    .A2(_02820_),
    .Y(_03014_),
    .B1(net186));
 sg13g2_nor3_1 _08563_ (.A(_02531_),
    .B(_03013_),
    .C(_03014_),
    .Y(_03015_));
 sg13g2_nor4_1 _08564_ (.A(net156),
    .B(_02563_),
    .C(net186),
    .D(_02422_),
    .Y(_03016_));
 sg13g2_a22oi_1 _08565_ (.Y(_03017_),
    .B1(_02419_),
    .B2(net226),
    .A2(net195),
    .A1(_02450_));
 sg13g2_a21oi_1 _08566_ (.A1(net149),
    .A2(_02540_),
    .Y(_03018_),
    .B1(_03017_));
 sg13g2_nor4_1 _08567_ (.A(_02721_),
    .B(_02667_),
    .C(_03016_),
    .D(_03018_),
    .Y(_03019_));
 sg13g2_a221oi_1 _08568_ (.B2(_02785_),
    .C1(_03019_),
    .B1(_03015_),
    .A1(_03008_),
    .Y(_03020_),
    .A2(_03012_));
 sg13g2_nand3_1 _08569_ (.B(_03003_),
    .C(_03020_),
    .A(_02982_),
    .Y(_03021_));
 sg13g2_o21ai_1 _08570_ (.B1(_02309_),
    .Y(_03022_),
    .A1(net190),
    .A2(net229));
 sg13g2_a221oi_1 _08571_ (.B2(net162),
    .C1(net181),
    .B1(_03022_),
    .A1(_02371_),
    .Y(_03023_),
    .A2(net184));
 sg13g2_o21ai_1 _08572_ (.B1(net197),
    .Y(_03024_),
    .A1(_02409_),
    .A2(net228));
 sg13g2_a221oi_1 _08573_ (.B2(_02427_),
    .C1(net226),
    .B1(_03024_),
    .A1(_02450_),
    .Y(_03025_),
    .A2(_02570_));
 sg13g2_mux2_1 _08574_ (.A0(_02757_),
    .A1(_02761_),
    .S(_02427_),
    .X(_03026_));
 sg13g2_o21ai_1 _08575_ (.B1(_03026_),
    .Y(_03027_),
    .A1(_03023_),
    .A2(_03025_));
 sg13g2_nand3_1 _08576_ (.B(net152),
    .C(_02732_),
    .A(net225),
    .Y(_03028_));
 sg13g2_o21ai_1 _08577_ (.B1(_03028_),
    .Y(_03029_),
    .A1(_02645_),
    .A2(_02736_));
 sg13g2_o21ai_1 _08578_ (.B1(net180),
    .Y(_03030_),
    .A1(net159),
    .A2(_02833_));
 sg13g2_o21ai_1 _08579_ (.B1(net144),
    .Y(_03031_),
    .A1(net162),
    .A2(_02894_));
 sg13g2_and2_1 _08580_ (.A(_03030_),
    .B(_03031_),
    .X(_03032_));
 sg13g2_nand3b_1 _08581_ (.B(net227),
    .C(net163),
    .Y(_03033_),
    .A_N(_02442_));
 sg13g2_a21o_1 _08582_ (.A2(_03033_),
    .A1(_02678_),
    .B1(_02708_),
    .X(_03034_));
 sg13g2_nor3_1 _08583_ (.A(net163),
    .B(net227),
    .C(net160),
    .Y(_03035_));
 sg13g2_o21ai_1 _08584_ (.B1(_02639_),
    .Y(_03036_),
    .A1(_02677_),
    .A2(_03035_));
 sg13g2_a22oi_1 _08585_ (.Y(_03037_),
    .B1(_03036_),
    .B2(_02905_),
    .A2(_03034_),
    .A1(_02710_));
 sg13g2_a221oi_1 _08586_ (.B2(_02900_),
    .C1(_03037_),
    .B1(_03032_),
    .A1(_03027_),
    .Y(_03038_),
    .A2(_03029_));
 sg13g2_nor2_1 _08587_ (.A(net240),
    .B(_03038_),
    .Y(_03039_));
 sg13g2_a21oi_1 _08588_ (.A1(_02886_),
    .A2(_02907_),
    .Y(_03040_),
    .B1(_02867_));
 sg13g2_a22oi_1 _08589_ (.Y(_03041_),
    .B1(_03040_),
    .B2(_02966_),
    .A2(_03039_),
    .A1(_03021_));
 sg13g2_buf_1 _08590_ (.A(_03041_),
    .X(_03042_));
 sg13g2_nor2_1 _08591_ (.A(net219),
    .B(_02867_),
    .Y(_03043_));
 sg13g2_nor2_1 _08592_ (.A(_02869_),
    .B(net240),
    .Y(_03044_));
 sg13g2_inv_1 _08593_ (.Y(_03045_),
    .A(_03044_));
 sg13g2_a221oi_1 _08594_ (.B2(_02713_),
    .C1(_03045_),
    .B1(_02693_),
    .A1(_02591_),
    .Y(_03046_),
    .A2(_02642_));
 sg13g2_a221oi_1 _08595_ (.B2(_02845_),
    .C1(_03046_),
    .B1(_03043_),
    .A1(net219),
    .Y(_03047_),
    .A2(_03042_));
 sg13g2_buf_2 _08596_ (.A(_03047_),
    .X(_03048_));
 sg13g2_xnor2_1 _08597_ (.Y(_03049_),
    .A(net166),
    .B(_03048_));
 sg13g2_buf_2 _08598_ (.A(_03049_),
    .X(_03050_));
 sg13g2_mux2_1 _08599_ (.A0(\dtop.vtop.dphases[0][2] ),
    .A1(_03050_),
    .S(_02861_),
    .X(_00177_));
 sg13g2_and2_1 _08600_ (.A(_02263_),
    .B(_02275_),
    .X(_03051_));
 sg13g2_buf_1 _08601_ (.A(_03051_),
    .X(_03052_));
 sg13g2_nand2_1 _08602_ (.Y(_03053_),
    .A(_03052_),
    .B(_02283_));
 sg13g2_buf_1 _08603_ (.A(_03053_),
    .X(_03054_));
 sg13g2_nand3_1 _08604_ (.B(net176),
    .C(net220),
    .A(net248),
    .Y(_03055_));
 sg13g2_nand2_1 _08605_ (.Y(_03056_),
    .A(net219),
    .B(net176));
 sg13g2_nand2_1 _08606_ (.Y(_03057_),
    .A(net219),
    .B(_02286_));
 sg13g2_nand4_1 _08607_ (.B(_02982_),
    .C(_03003_),
    .A(_02856_),
    .Y(_03058_),
    .D(_03020_));
 sg13g2_nand2_1 _08608_ (.Y(_03059_),
    .A(net220),
    .B(_03038_));
 sg13g2_nand2_1 _08609_ (.Y(_03060_),
    .A(net189),
    .B(_02663_));
 sg13g2_nand3_1 _08610_ (.B(net224),
    .C(_03060_),
    .A(net98),
    .Y(_03061_));
 sg13g2_o21ai_1 _08611_ (.B1(net181),
    .Y(_03062_),
    .A1(net156),
    .A2(net157));
 sg13g2_nand4_1 _08612_ (.B(net147),
    .C(_02892_),
    .A(net188),
    .Y(_03063_),
    .D(_03062_));
 sg13g2_nor3_1 _08613_ (.A(net244),
    .B(net192),
    .C(_02633_),
    .Y(_03064_));
 sg13g2_nor3_1 _08614_ (.A(net142),
    .B(_02560_),
    .C(_03064_),
    .Y(_03065_));
 sg13g2_a21oi_1 _08615_ (.A1(_02699_),
    .A2(_02894_),
    .Y(_03066_),
    .B1(net179));
 sg13g2_a22oi_1 _08616_ (.Y(_03067_),
    .B1(_03066_),
    .B2(_02681_),
    .A2(_03065_),
    .A1(_03063_));
 sg13g2_a22oi_1 _08617_ (.Y(_03068_),
    .B1(_02493_),
    .B2(net160),
    .A2(net157),
    .A1(_02573_));
 sg13g2_o21ai_1 _08618_ (.B1(net118),
    .Y(_03069_),
    .A1(_02451_),
    .A2(_02493_));
 sg13g2_nand2b_1 _08619_ (.Y(_03070_),
    .B(net150),
    .A_N(_02573_));
 sg13g2_nand2_1 _08620_ (.Y(_03071_),
    .A(net113),
    .B(_03070_));
 sg13g2_nand3_1 _08621_ (.B(_03069_),
    .C(_03071_),
    .A(_03068_),
    .Y(_03072_));
 sg13g2_nand4_1 _08622_ (.B(net228),
    .C(_02332_),
    .A(net190),
    .Y(_03073_),
    .D(_02350_));
 sg13g2_nand3_1 _08623_ (.B(net124),
    .C(_03073_),
    .A(_02461_),
    .Y(_03074_));
 sg13g2_a221oi_1 _08624_ (.B2(_02833_),
    .C1(net152),
    .B1(net149),
    .A1(net242),
    .Y(_03075_),
    .A2(net241));
 sg13g2_a221oi_1 _08625_ (.B2(_03074_),
    .C1(_03075_),
    .B1(_02645_),
    .A1(net114),
    .Y(_03076_),
    .A2(net180));
 sg13g2_a22oi_1 _08626_ (.Y(_03077_),
    .B1(_03072_),
    .B2(_03076_),
    .A2(_03067_),
    .A1(_03061_));
 sg13g2_buf_1 _08627_ (.A(_03077_),
    .X(_03078_));
 sg13g2_xnor2_1 _08628_ (.Y(_03079_),
    .A(net244),
    .B(net197));
 sg13g2_nor3_1 _08629_ (.A(net225),
    .B(net161),
    .C(net226),
    .Y(_03080_));
 sg13g2_a221oi_1 _08630_ (.B2(_03079_),
    .C1(_03080_),
    .B1(_02699_),
    .A1(net225),
    .Y(_03081_),
    .A2(net144));
 sg13g2_nor2_1 _08631_ (.A(_02473_),
    .B(net198),
    .Y(_03082_));
 sg13g2_nor2_1 _08632_ (.A(net244),
    .B(net184),
    .Y(_03083_));
 sg13g2_or3_1 _08633_ (.A(_02782_),
    .B(_03082_),
    .C(_03083_),
    .X(_03084_));
 sg13g2_nand3_1 _08634_ (.B(_03081_),
    .C(_03084_),
    .A(net179),
    .Y(_03085_));
 sg13g2_o21ai_1 _08635_ (.B1(_03079_),
    .Y(_03086_),
    .A1(net161),
    .A2(_02682_));
 sg13g2_nor2_1 _08636_ (.A(net225),
    .B(_02596_),
    .Y(_03087_));
 sg13g2_a21oi_1 _08637_ (.A1(net225),
    .A2(_02633_),
    .Y(_03088_),
    .B1(_03087_));
 sg13g2_mux2_1 _08638_ (.A0(net149),
    .A1(net185),
    .S(net244),
    .X(_03089_));
 sg13g2_nand2_1 _08639_ (.Y(_03090_),
    .A(net178),
    .B(_03089_));
 sg13g2_nand4_1 _08640_ (.B(_03086_),
    .C(_03088_),
    .A(_02561_),
    .Y(_03091_),
    .D(_03090_));
 sg13g2_a22oi_1 _08641_ (.Y(_03092_),
    .B1(_03091_),
    .B2(_02626_),
    .A2(_03085_),
    .A1(_02928_));
 sg13g2_buf_1 _08642_ (.A(_03092_),
    .X(_03093_));
 sg13g2_nand2_1 _08643_ (.Y(_03094_),
    .A(net144),
    .B(_02894_));
 sg13g2_nand4_1 _08644_ (.B(net180),
    .C(net222),
    .A(net118),
    .Y(_03095_),
    .D(_02833_));
 sg13g2_o21ai_1 _08645_ (.B1(_03095_),
    .Y(_03096_),
    .A1(_02691_),
    .A2(_03094_));
 sg13g2_buf_1 _08646_ (.A(_03096_),
    .X(_03097_));
 sg13g2_o21ai_1 _08647_ (.B1(net120),
    .Y(_03098_),
    .A1(_02461_),
    .A2(_02678_));
 sg13g2_nand4_1 _08648_ (.B(net122),
    .C(net147),
    .A(_02474_),
    .Y(_03099_),
    .D(_02700_));
 sg13g2_nand3_1 _08649_ (.B(net147),
    .C(net178),
    .A(net189),
    .Y(_03100_));
 sg13g2_nand4_1 _08650_ (.B(_03098_),
    .C(_03099_),
    .A(net114),
    .Y(_03101_),
    .D(_03100_));
 sg13g2_buf_1 _08651_ (.A(_03101_),
    .X(_03102_));
 sg13g2_nand2_1 _08652_ (.Y(_03103_),
    .A(net125),
    .B(_02682_));
 sg13g2_nand2_1 _08653_ (.Y(_03104_),
    .A(net181),
    .B(net143));
 sg13g2_a221oi_1 _08654_ (.B2(_03082_),
    .C1(net158),
    .B1(_03104_),
    .A1(net242),
    .Y(_03105_),
    .A2(net241));
 sg13g2_a21oi_1 _08655_ (.A1(net148),
    .A2(net143),
    .Y(_03106_),
    .B1(_02596_));
 sg13g2_a221oi_1 _08656_ (.B2(_02743_),
    .C1(_02742_),
    .B1(_03106_),
    .A1(_03103_),
    .Y(_03107_),
    .A2(_03105_));
 sg13g2_buf_1 _08657_ (.A(_03107_),
    .X(_03108_));
 sg13g2_a221oi_1 _08658_ (.B2(_03108_),
    .C1(net240),
    .B1(_03102_),
    .A1(_02900_),
    .Y(_03109_),
    .A2(_03097_));
 sg13g2_o21ai_1 _08659_ (.B1(_03109_),
    .Y(_03110_),
    .A1(_03078_),
    .A2(_03093_));
 sg13g2_nand3_1 _08660_ (.B(_03059_),
    .C(_03110_),
    .A(_03058_),
    .Y(_03111_));
 sg13g2_mux2_1 _08661_ (.A0(_03056_),
    .A1(_03057_),
    .S(_03111_),
    .X(_03112_));
 sg13g2_o21ai_1 _08662_ (.B1(_03112_),
    .Y(_03113_),
    .A1(_02715_),
    .A2(_03055_));
 sg13g2_nand2_1 _08663_ (.Y(_03114_),
    .A(_02286_),
    .B(net240));
 sg13g2_nor2_1 _08664_ (.A(_02871_),
    .B(_03114_),
    .Y(_03115_));
 sg13g2_nand2_1 _08665_ (.Y(_03116_),
    .A(_02286_),
    .B(_02867_));
 sg13g2_nor2_1 _08666_ (.A(net219),
    .B(_03116_),
    .Y(_03117_));
 sg13g2_nand2_1 _08667_ (.Y(_03118_),
    .A(_03053_),
    .B(_02867_));
 sg13g2_nor2_1 _08668_ (.A(_02870_),
    .B(_03118_),
    .Y(_03119_));
 sg13g2_mux2_1 _08669_ (.A0(_03117_),
    .A1(_03119_),
    .S(_02968_),
    .X(_03120_));
 sg13g2_a21o_1 _08670_ (.A2(_03115_),
    .A1(_02715_),
    .B1(_03120_),
    .X(_03121_));
 sg13g2_or2_1 _08671_ (.X(_03122_),
    .B(_03121_),
    .A(_03113_));
 sg13g2_buf_8 _08672_ (.A(_03122_),
    .X(_03123_));
 sg13g2_nand2_1 _08673_ (.Y(_03124_),
    .A(\dtop.vtop.dphases[0][3] ),
    .B(net239));
 sg13g2_o21ai_1 _08674_ (.B1(_03124_),
    .Y(_00178_),
    .A1(net239),
    .A2(_03123_));
 sg13g2_a221oi_1 _08675_ (.B2(_03108_),
    .C1(_02867_),
    .B1(_03102_),
    .A1(_02900_),
    .Y(_03125_),
    .A2(_03097_));
 sg13g2_o21ai_1 _08676_ (.B1(_03125_),
    .Y(_03126_),
    .A1(_03078_),
    .A2(_03093_));
 sg13g2_nand4_1 _08677_ (.B(_02695_),
    .C(net221),
    .A(net114),
    .Y(_03127_),
    .D(_02639_));
 sg13g2_nand4_1 _08678_ (.B(net120),
    .C(net222),
    .A(net113),
    .Y(_03128_),
    .D(_02889_));
 sg13g2_nand2_1 _08679_ (.Y(_03129_),
    .A(_03127_),
    .B(_03128_));
 sg13g2_nand3_1 _08680_ (.B(_02625_),
    .C(_02898_),
    .A(net153),
    .Y(_03130_));
 sg13g2_nor2_1 _08681_ (.A(net188),
    .B(_02625_),
    .Y(_03131_));
 sg13g2_nand4_1 _08682_ (.B(net223),
    .C(_03073_),
    .A(net152),
    .Y(_03132_),
    .D(_03131_));
 sg13g2_a221oi_1 _08683_ (.B2(_03132_),
    .C1(_03075_),
    .B1(_03130_),
    .A1(_02548_),
    .Y(_03133_),
    .A2(net180));
 sg13g2_buf_1 _08684_ (.A(_03133_),
    .X(_03134_));
 sg13g2_nor3_1 _08685_ (.A(_02549_),
    .B(net117),
    .C(net143),
    .Y(_03135_));
 sg13g2_nor2_1 _08686_ (.A(_02565_),
    .B(_02766_),
    .Y(_03136_));
 sg13g2_a22oi_1 _08687_ (.Y(_03137_),
    .B1(_03136_),
    .B2(_02952_),
    .A2(_02873_),
    .A1(_03135_));
 sg13g2_a21oi_1 _08688_ (.A1(net192),
    .A2(_02782_),
    .Y(_03138_),
    .B1(net193));
 sg13g2_mux2_1 _08689_ (.A0(_03070_),
    .A1(_03138_),
    .S(net179),
    .X(_03139_));
 sg13g2_nor3_1 _08690_ (.A(net155),
    .B(net114),
    .C(net221),
    .Y(_03140_));
 sg13g2_a22oi_1 _08691_ (.Y(_03141_),
    .B1(_02551_),
    .B2(_02558_),
    .A2(net241),
    .A1(net242));
 sg13g2_o21ai_1 _08692_ (.B1(_03141_),
    .Y(_03142_),
    .A1(net147),
    .A2(net178));
 sg13g2_o21ai_1 _08693_ (.B1(net223),
    .Y(_03143_),
    .A1(_02451_),
    .A2(_02493_));
 sg13g2_nand2_1 _08694_ (.Y(_03144_),
    .A(net155),
    .B(net221));
 sg13g2_a221oi_1 _08695_ (.B2(_03143_),
    .C1(_03144_),
    .B1(_03142_),
    .A1(_02647_),
    .Y(_03145_),
    .A2(_02648_));
 sg13g2_a21o_1 _08696_ (.A2(_03140_),
    .A1(_03139_),
    .B1(_03145_),
    .X(_03146_));
 sg13g2_a221oi_1 _08697_ (.B2(_03137_),
    .C1(_03146_),
    .B1(_03134_),
    .A1(_02684_),
    .Y(_03147_),
    .A2(_03129_));
 sg13g2_nor2_1 _08698_ (.A(net121),
    .B(net115),
    .Y(_03148_));
 sg13g2_nor2_1 _08699_ (.A(net223),
    .B(_02625_),
    .Y(_03149_));
 sg13g2_nand3_1 _08700_ (.B(_02677_),
    .C(_03149_),
    .A(net98),
    .Y(_03150_));
 sg13g2_o21ai_1 _08701_ (.B1(_03150_),
    .Y(_03151_),
    .A1(_02742_),
    .A2(_03148_));
 sg13g2_o21ai_1 _08702_ (.B1(net120),
    .Y(_03152_),
    .A1(net147),
    .A2(_02782_));
 sg13g2_o21ai_1 _08703_ (.B1(_02596_),
    .Y(_03153_),
    .A1(_02443_),
    .A2(_02776_));
 sg13g2_a21o_1 _08704_ (.A2(_03152_),
    .A1(net113),
    .B1(_03153_),
    .X(_03154_));
 sg13g2_nor3_1 _08705_ (.A(net121),
    .B(net98),
    .C(_02437_),
    .Y(_03155_));
 sg13g2_a21oi_1 _08706_ (.A1(net121),
    .A2(_03154_),
    .Y(_03156_),
    .B1(_03155_));
 sg13g2_a21oi_1 _08707_ (.A1(_03151_),
    .A2(_03156_),
    .Y(_03157_),
    .B1(_02856_));
 sg13g2_a21oi_1 _08708_ (.A1(_03147_),
    .A2(_03157_),
    .Y(_03158_),
    .B1(net248));
 sg13g2_nand2_1 _08709_ (.Y(_03159_),
    .A(_03126_),
    .B(_03158_));
 sg13g2_o21ai_1 _08710_ (.B1(_03159_),
    .Y(_03160_),
    .A1(net177),
    .A2(_03042_));
 sg13g2_xnor2_1 _08711_ (.Y(_03161_),
    .A(_02287_),
    .B(_03160_));
 sg13g2_buf_2 _08712_ (.A(_03161_),
    .X(_03162_));
 sg13g2_mux2_1 _08713_ (.A0(\dtop.vtop.dphases[0][4] ),
    .A1(_03162_),
    .S(_02861_),
    .X(_00179_));
 sg13g2_a221oi_1 _08714_ (.B2(_03128_),
    .C1(_02683_),
    .B1(_03127_),
    .A1(_02681_),
    .Y(_03163_),
    .A2(_02682_));
 sg13g2_o21ai_1 _08715_ (.B1(net240),
    .Y(_03164_),
    .A1(_03163_),
    .A2(_03146_));
 sg13g2_nand3_1 _08716_ (.B(_03134_),
    .C(_03137_),
    .A(net240),
    .Y(_03165_));
 sg13g2_nand3_1 _08717_ (.B(_03151_),
    .C(_03156_),
    .A(_02855_),
    .Y(_03166_));
 sg13g2_a221oi_1 _08718_ (.B2(_03153_),
    .C1(net221),
    .B1(_02889_),
    .A1(_02647_),
    .Y(_03167_),
    .A2(_02648_));
 sg13g2_nor2_1 _08719_ (.A(_02620_),
    .B(net269),
    .Y(_03168_));
 sg13g2_buf_1 _08720_ (.A(_02465_),
    .X(_03169_));
 sg13g2_nor2_1 _08721_ (.A(_02622_),
    .B(net254),
    .Y(_03170_));
 sg13g2_o21ai_1 _08722_ (.B1(net270),
    .Y(_03171_),
    .A1(_03168_),
    .A2(_03170_));
 sg13g2_nand2_1 _08723_ (.Y(_03172_),
    .A(_02621_),
    .B(net254));
 sg13g2_nand2_1 _08724_ (.Y(_03173_),
    .A(_00055_),
    .B(net269));
 sg13g2_nand3_1 _08725_ (.B(_03172_),
    .C(_03173_),
    .A(net271),
    .Y(_03174_));
 sg13g2_o21ai_1 _08726_ (.B1(net149),
    .Y(_03175_),
    .A1(net226),
    .A2(net160));
 sg13g2_nor3_1 _08727_ (.A(net188),
    .B(net156),
    .C(net223),
    .Y(_03176_));
 sg13g2_a221oi_1 _08728_ (.B2(_03176_),
    .C1(net118),
    .B1(_03175_),
    .A1(_03171_),
    .Y(_03177_),
    .A2(_03174_));
 sg13g2_or2_1 _08729_ (.X(_03178_),
    .B(_03177_),
    .A(_03167_));
 sg13g2_or3_1 _08730_ (.A(net155),
    .B(net118),
    .C(_03138_),
    .X(_03179_));
 sg13g2_o21ai_1 _08731_ (.B1(net161),
    .Y(_03180_),
    .A1(net192),
    .A2(net178));
 sg13g2_nand3_1 _08732_ (.B(net114),
    .C(_03180_),
    .A(net155),
    .Y(_03181_));
 sg13g2_nand2_1 _08733_ (.Y(_03182_),
    .A(net113),
    .B(_02732_));
 sg13g2_nand2_1 _08734_ (.Y(_03183_),
    .A(net114),
    .B(_03149_));
 sg13g2_a22oi_1 _08735_ (.Y(_03184_),
    .B1(_03182_),
    .B2(_03183_),
    .A2(_03181_),
    .A1(_03179_));
 sg13g2_or4_1 _08736_ (.A(_02855_),
    .B(_03134_),
    .C(_03178_),
    .D(_03184_),
    .X(_03185_));
 sg13g2_nand4_1 _08737_ (.B(_03165_),
    .C(_03166_),
    .A(_03164_),
    .Y(_03186_),
    .D(_03185_));
 sg13g2_mux2_1 _08738_ (.A0(_03056_),
    .A1(_03057_),
    .S(_03186_),
    .X(_03187_));
 sg13g2_nor2_1 _08739_ (.A(_02870_),
    .B(net176),
    .Y(_03188_));
 sg13g2_nand4_1 _08740_ (.B(_03059_),
    .C(_03110_),
    .A(_03058_),
    .Y(_03189_),
    .D(_03188_));
 sg13g2_nand2_1 _08741_ (.Y(_03190_),
    .A(net248),
    .B(_03054_));
 sg13g2_or2_1 _08742_ (.X(_03191_),
    .B(_03190_),
    .A(_03110_));
 sg13g2_a21o_1 _08743_ (.A2(_03059_),
    .A1(_03058_),
    .B1(_03190_),
    .X(_03192_));
 sg13g2_and4_1 _08744_ (.A(_03187_),
    .B(_03189_),
    .C(_03191_),
    .D(_03192_),
    .X(_03193_));
 sg13g2_buf_1 _08745_ (.A(_03193_),
    .X(_03194_));
 sg13g2_nand2_1 _08746_ (.Y(_03195_),
    .A(\dtop.vtop.dphases[0][5] ),
    .B(_02864_));
 sg13g2_o21ai_1 _08747_ (.B1(_03195_),
    .Y(_00180_),
    .A1(_02864_),
    .A2(_03194_));
 sg13g2_nand3_1 _08748_ (.B(_03147_),
    .C(_03157_),
    .A(_02286_),
    .Y(_03196_));
 sg13g2_a221oi_1 _08749_ (.B2(_03108_),
    .C1(_03114_),
    .B1(_03102_),
    .A1(_02900_),
    .Y(_03197_),
    .A2(_03097_));
 sg13g2_o21ai_1 _08750_ (.B1(_03197_),
    .Y(_03198_),
    .A1(_03078_),
    .A2(_03093_));
 sg13g2_a21o_1 _08751_ (.A2(_03198_),
    .A1(_03196_),
    .B1(_02871_),
    .X(_03199_));
 sg13g2_a221oi_1 _08752_ (.B2(_03181_),
    .C1(_03116_),
    .B1(_03179_),
    .A1(_02942_),
    .Y(_03200_),
    .A2(_02629_));
 sg13g2_xnor2_1 _08753_ (.Y(_03201_),
    .A(net97),
    .B(net222));
 sg13g2_nor3_1 _08754_ (.A(_02950_),
    .B(_03116_),
    .C(_03201_),
    .Y(_03202_));
 sg13g2_xnor2_1 _08755_ (.Y(_03203_),
    .A(net98),
    .B(net222));
 sg13g2_nor2_1 _08756_ (.A(_03118_),
    .B(_03203_),
    .Y(_03204_));
 sg13g2_nor3_1 _08757_ (.A(net121),
    .B(net97),
    .C(_03138_),
    .Y(_03205_));
 sg13g2_and3_1 _08758_ (.X(_03206_),
    .A(net155),
    .B(net114),
    .C(_03180_));
 sg13g2_buf_1 _08759_ (.A(_03206_),
    .X(_03207_));
 sg13g2_nor4_1 _08760_ (.A(_02962_),
    .B(_03118_),
    .C(_03205_),
    .D(_03207_),
    .Y(_03208_));
 sg13g2_or4_1 _08761_ (.A(_03200_),
    .B(_03202_),
    .C(_03204_),
    .D(_03208_),
    .X(_03209_));
 sg13g2_nor2_1 _08762_ (.A(_03167_),
    .B(_03177_),
    .Y(_03210_));
 sg13g2_mux2_1 _08763_ (.A0(_02732_),
    .A1(_03149_),
    .S(net97),
    .X(_03211_));
 sg13g2_o21ai_1 _08764_ (.B1(_03211_),
    .Y(_03212_),
    .A1(_03205_),
    .A2(_03207_));
 sg13g2_nand2_1 _08765_ (.Y(_03213_),
    .A(_03053_),
    .B(net240));
 sg13g2_a21oi_1 _08766_ (.A1(_03210_),
    .A2(_03212_),
    .Y(_03214_),
    .B1(_03213_));
 sg13g2_nor4_1 _08767_ (.A(_03114_),
    .B(_03134_),
    .C(_03178_),
    .D(_03184_),
    .Y(_03215_));
 sg13g2_nor2b_1 _08768_ (.A(_03213_),
    .B_N(_03134_),
    .Y(_03216_));
 sg13g2_nor4_1 _08769_ (.A(_03209_),
    .B(_03214_),
    .C(_03215_),
    .D(_03216_),
    .Y(_03217_));
 sg13g2_a21oi_1 _08770_ (.A1(_03147_),
    .A2(_03157_),
    .Y(_03218_),
    .B1(_03190_));
 sg13g2_a22oi_1 _08771_ (.Y(_03219_),
    .B1(_03218_),
    .B2(_03126_),
    .A2(_03217_),
    .A1(net219));
 sg13g2_and2_1 _08772_ (.A(_03199_),
    .B(_03219_),
    .X(_03220_));
 sg13g2_buf_2 _08773_ (.A(_03220_),
    .X(_03221_));
 sg13g2_mux2_1 _08774_ (.A0(\dtop.vtop.dphases[0][6] ),
    .A1(_03221_),
    .S(_02861_),
    .X(_00181_));
 sg13g2_xnor2_1 _08775_ (.Y(_03222_),
    .A(_03054_),
    .B(_03186_));
 sg13g2_nor3_1 _08776_ (.A(_02962_),
    .B(_03205_),
    .C(_03207_),
    .Y(_03223_));
 sg13g2_nor2_1 _08777_ (.A(_03201_),
    .B(_03223_),
    .Y(_03224_));
 sg13g2_xnor2_1 _08778_ (.Y(_03225_),
    .A(net166),
    .B(_03224_));
 sg13g2_nand2_1 _08779_ (.Y(_03226_),
    .A(net220),
    .B(_03225_));
 sg13g2_o21ai_1 _08780_ (.B1(_03226_),
    .Y(_03227_),
    .A1(net247),
    .A2(net220));
 sg13g2_nand2_1 _08781_ (.Y(_03228_),
    .A(net177),
    .B(_03227_));
 sg13g2_o21ai_1 _08782_ (.B1(_03228_),
    .Y(_03229_),
    .A1(net177),
    .A2(_03222_));
 sg13g2_buf_1 _08783_ (.A(_03229_),
    .X(_03230_));
 sg13g2_mux2_1 _08784_ (.A0(\dtop.vtop.dphases[0][7] ),
    .A1(net33),
    .S(_02861_),
    .X(_00182_));
 sg13g2_nand2_1 _08785_ (.Y(_03231_),
    .A(net177),
    .B(_03052_));
 sg13g2_o21ai_1 _08786_ (.B1(_03231_),
    .Y(_03232_),
    .A1(net177),
    .A2(_03217_));
 sg13g2_buf_1 _08787_ (.A(_03232_),
    .X(_03233_));
 sg13g2_inv_1 _08788_ (.Y(_03234_),
    .A(_03233_));
 sg13g2_nand2_1 _08789_ (.Y(_03235_),
    .A(\dtop.vtop.dphases[0][8] ),
    .B(net239));
 sg13g2_o21ai_1 _08790_ (.B1(_03235_),
    .Y(_00183_),
    .A1(net239),
    .A2(_03234_));
 sg13g2_nand2_1 _08791_ (.Y(_03236_),
    .A(\dtop.vtop.dphases[0][9] ),
    .B(net239));
 sg13g2_o21ai_1 _08792_ (.B1(_03236_),
    .Y(_00184_),
    .A1(net247),
    .A2(net239));
 sg13g2_nor2_1 _08793_ (.A(_05405_),
    .B(_01315_),
    .Y(_03237_));
 sg13g2_buf_2 _08794_ (.A(_03237_),
    .X(_03238_));
 sg13g2_buf_1 _08795_ (.A(_03238_),
    .X(_03239_));
 sg13g2_mux2_1 _08796_ (.A0(\dtop.vtop.dphases[1][0] ),
    .A1(_02859_),
    .S(_03239_),
    .X(_00185_));
 sg13g2_buf_1 _08797_ (.A(_03052_),
    .X(_03240_));
 sg13g2_mux2_1 _08798_ (.A0(\dtop.vtop.dphases[1][10] ),
    .A1(_03240_),
    .S(net218),
    .X(_00186_));
 sg13g2_inv_1 _08799_ (.Y(_03241_),
    .A(\dtop.vtop.dphases[1][1] ));
 sg13g2_nand2_1 _08800_ (.Y(_03242_),
    .A(_02974_),
    .B(_03238_));
 sg13g2_o21ai_1 _08801_ (.B1(_03242_),
    .Y(_00187_),
    .A1(_03241_),
    .A2(net218));
 sg13g2_inv_1 _08802_ (.Y(_03243_),
    .A(\dtop.vtop.dphases[1][2] ));
 sg13g2_nand2_1 _08803_ (.Y(_03244_),
    .A(_03050_),
    .B(_03238_));
 sg13g2_o21ai_1 _08804_ (.B1(_03244_),
    .Y(_00188_),
    .A1(_03243_),
    .A2(net218));
 sg13g2_inv_1 _08805_ (.Y(_03245_),
    .A(\dtop.vtop.dphases[1][3] ));
 sg13g2_nand2b_1 _08806_ (.Y(_03246_),
    .B(_03238_),
    .A_N(_03123_));
 sg13g2_o21ai_1 _08807_ (.B1(_03246_),
    .Y(_00189_),
    .A1(_03245_),
    .A2(_03239_));
 sg13g2_mux2_1 _08808_ (.A0(\dtop.vtop.dphases[1][4] ),
    .A1(_03162_),
    .S(net218),
    .X(_00190_));
 sg13g2_nand4_1 _08809_ (.B(_03189_),
    .C(_03191_),
    .A(_03187_),
    .Y(_03247_),
    .D(_03192_));
 sg13g2_buf_2 _08810_ (.A(_03247_),
    .X(_03248_));
 sg13g2_mux2_1 _08811_ (.A0(\dtop.vtop.dphases[1][5] ),
    .A1(_03248_),
    .S(net218),
    .X(_00191_));
 sg13g2_mux2_1 _08812_ (.A0(\dtop.vtop.dphases[1][6] ),
    .A1(_03221_),
    .S(net218),
    .X(_00192_));
 sg13g2_mux2_1 _08813_ (.A0(\dtop.vtop.dphases[1][7] ),
    .A1(net33),
    .S(net218),
    .X(_00193_));
 sg13g2_mux2_1 _08814_ (.A0(\dtop.vtop.dphases[1][8] ),
    .A1(_03233_),
    .S(_03238_),
    .X(_00194_));
 sg13g2_nor2_1 _08815_ (.A(_02277_),
    .B(_03043_),
    .Y(_03249_));
 sg13g2_a21oi_1 _08816_ (.A1(_03043_),
    .A2(_03225_),
    .Y(_03250_),
    .B1(_03249_));
 sg13g2_buf_2 _08817_ (.A(_03250_),
    .X(_03251_));
 sg13g2_nor2_1 _08818_ (.A(\dtop.vtop.dphases[1][9] ),
    .B(_03238_),
    .Y(_03252_));
 sg13g2_a21oi_1 _08819_ (.A1(net218),
    .A2(_03251_),
    .Y(_00195_),
    .B1(_03252_));
 sg13g2_nor2_1 _08820_ (.A(_01453_),
    .B(_05405_),
    .Y(_03253_));
 sg13g2_buf_2 _08821_ (.A(_03253_),
    .X(_03254_));
 sg13g2_mux2_1 _08822_ (.A0(\dtop.vtop.dphases[2][0] ),
    .A1(_02859_),
    .S(_03254_),
    .X(_00196_));
 sg13g2_nand3_1 _08823_ (.B(_05163_),
    .C(net277),
    .A(net426),
    .Y(_03255_));
 sg13g2_buf_1 _08824_ (.A(_03255_),
    .X(_03256_));
 sg13g2_nor2_1 _08825_ (.A(net247),
    .B(net253),
    .Y(_03257_));
 sg13g2_a21o_1 _08826_ (.A2(net253),
    .A1(\dtop.vtop.dphases[2][10] ),
    .B1(_03257_),
    .X(_00197_));
 sg13g2_inv_1 _08827_ (.Y(_03258_),
    .A(\dtop.vtop.dphases[2][1] ));
 sg13g2_nand2_1 _08828_ (.Y(_03259_),
    .A(_02974_),
    .B(_03254_));
 sg13g2_o21ai_1 _08829_ (.B1(_03259_),
    .Y(_00198_),
    .A1(_03258_),
    .A2(_03254_));
 sg13g2_inv_1 _08830_ (.Y(_03260_),
    .A(\dtop.vtop.dphases[2][2] ));
 sg13g2_nand2_1 _08831_ (.Y(_03261_),
    .A(_03050_),
    .B(_03254_));
 sg13g2_o21ai_1 _08832_ (.B1(_03261_),
    .Y(_00199_),
    .A1(_03260_),
    .A2(_03254_));
 sg13g2_nand2_1 _08833_ (.Y(_03262_),
    .A(\dtop.vtop.dphases[2][3] ),
    .B(net253));
 sg13g2_o21ai_1 _08834_ (.B1(_03262_),
    .Y(_00200_),
    .A1(_03123_),
    .A2(_03256_));
 sg13g2_mux2_1 _08835_ (.A0(\dtop.vtop.dphases[2][4] ),
    .A1(_03162_),
    .S(_03254_),
    .X(_00201_));
 sg13g2_nand2_1 _08836_ (.Y(_03263_),
    .A(\dtop.vtop.dphases[2][5] ),
    .B(net253));
 sg13g2_o21ai_1 _08837_ (.B1(_03263_),
    .Y(_00202_),
    .A1(_03194_),
    .A2(net253));
 sg13g2_mux2_1 _08838_ (.A0(\dtop.vtop.dphases[2][6] ),
    .A1(_03221_),
    .S(_03254_),
    .X(_00203_));
 sg13g2_mux2_1 _08839_ (.A0(\dtop.vtop.dphases[2][7] ),
    .A1(_03230_),
    .S(_03254_),
    .X(_00204_));
 sg13g2_nand2_1 _08840_ (.Y(_03264_),
    .A(\dtop.vtop.dphases[2][8] ),
    .B(net253));
 sg13g2_o21ai_1 _08841_ (.B1(_03264_),
    .Y(_00205_),
    .A1(_03234_),
    .A2(net253));
 sg13g2_a21o_1 _08842_ (.A2(net253),
    .A1(\dtop.vtop.dphases[2][9] ),
    .B1(_03257_),
    .X(_00206_));
 sg13g2_nand2b_1 _08843_ (.Y(_03265_),
    .B(_05229_),
    .A_N(_01193_));
 sg13g2_nor2_1 _08844_ (.A(_05137_),
    .B(_05264_),
    .Y(_03266_));
 sg13g2_o21ai_1 _08845_ (.B1(net390),
    .Y(_03267_),
    .A1(_01201_),
    .A2(_03266_));
 sg13g2_o21ai_1 _08846_ (.B1(_03267_),
    .Y(_03268_),
    .A1(_05406_),
    .A2(_03265_));
 sg13g2_buf_1 _08847_ (.A(_03268_),
    .X(_03269_));
 sg13g2_xnor2_1 _08848_ (.Y(_03270_),
    .A(_02846_),
    .B(_03269_));
 sg13g2_nor2_1 _08849_ (.A(_02251_),
    .B(_03270_),
    .Y(_03271_));
 sg13g2_nor2_1 _08850_ (.A(_05265_),
    .B(_02848_),
    .Y(_03272_));
 sg13g2_buf_2 _08851_ (.A(_03272_),
    .X(_03273_));
 sg13g2_buf_1 _08852_ (.A(\dtop.vtop.pipeline.zg[5] ),
    .X(_03274_));
 sg13g2_inv_1 _08853_ (.Y(_03275_),
    .A(_03274_));
 sg13g2_buf_1 _08854_ (.A(\dtop.vtop.pipeline.z[11] ),
    .X(_03276_));
 sg13g2_buf_2 _08855_ (.A(\dtop.vtop.pipeline.zg[6] ),
    .X(_03277_));
 sg13g2_nand2b_1 _08856_ (.Y(_03278_),
    .B(_03277_),
    .A_N(_03276_));
 sg13g2_and2_1 _08857_ (.A(_03275_),
    .B(_03278_),
    .X(_03279_));
 sg13g2_buf_1 _08858_ (.A(\dtop.vtop.pipeline.z[10] ),
    .X(_03280_));
 sg13g2_and2_1 _08859_ (.A(net409),
    .B(_03278_),
    .X(_03281_));
 sg13g2_buf_1 _08860_ (.A(\dtop.vtop.pipeline.z[8] ),
    .X(_03282_));
 sg13g2_buf_1 _08861_ (.A(\dtop.vtop.pipeline.zg[3] ),
    .X(_03283_));
 sg13g2_inv_1 _08862_ (.Y(_03284_),
    .A(_03283_));
 sg13g2_buf_1 _08863_ (.A(\dtop.vtop.pipeline.z[7] ),
    .X(_03285_));
 sg13g2_inv_1 _08864_ (.Y(_03286_),
    .A(\dtop.vtop.pipeline.zg[2] ));
 sg13g2_inv_1 _08865_ (.Y(_03287_),
    .A(_03285_));
 sg13g2_buf_1 _08866_ (.A(\dtop.vtop.pipeline.z[6] ),
    .X(_03288_));
 sg13g2_nand2b_1 _08867_ (.Y(_03289_),
    .B(_03288_),
    .A_N(\dtop.vtop.pipeline.zg[1] ));
 sg13g2_nor2b_1 _08868_ (.A(\dtop.vtop.pipeline.z[5] ),
    .B_N(\dtop.vtop.pipeline.zg[0] ),
    .Y(_03290_));
 sg13g2_nor2b_1 _08869_ (.A(_03288_),
    .B_N(\dtop.vtop.pipeline.zg[1] ),
    .Y(_03291_));
 sg13g2_a221oi_1 _08870_ (.B2(_03290_),
    .C1(_03291_),
    .B1(_03289_),
    .A1(_03287_),
    .Y(_03292_),
    .A2(\dtop.vtop.pipeline.zg[2] ));
 sg13g2_a221oi_1 _08871_ (.B2(_03286_),
    .C1(_03292_),
    .B1(_03285_),
    .A1(_03282_),
    .Y(_03293_),
    .A2(_03284_));
 sg13g2_buf_2 _08872_ (.A(\dtop.vtop.pipeline.z[9] ),
    .X(_03294_));
 sg13g2_inv_1 _08873_ (.Y(_03295_),
    .A(_03294_));
 sg13g2_buf_1 _08874_ (.A(\dtop.vtop.pipeline.zg[4] ),
    .X(_03296_));
 sg13g2_nand2_1 _08875_ (.Y(_03297_),
    .A(_03295_),
    .B(net408));
 sg13g2_o21ai_1 _08876_ (.B1(_03297_),
    .Y(_03298_),
    .A1(_03282_),
    .A2(_03284_));
 sg13g2_nand2b_1 _08877_ (.Y(_03299_),
    .B(_03294_),
    .A_N(net408));
 sg13g2_o21ai_1 _08878_ (.B1(_03299_),
    .Y(_03300_),
    .A1(_03293_),
    .A2(_03298_));
 sg13g2_o21ai_1 _08879_ (.B1(_03300_),
    .Y(_03301_),
    .A1(_03279_),
    .A2(_03281_));
 sg13g2_nor2b_1 _08880_ (.A(_03274_),
    .B_N(_03280_),
    .Y(_03302_));
 sg13g2_nor2b_1 _08881_ (.A(_03277_),
    .B_N(_03276_),
    .Y(_03303_));
 sg13g2_a21oi_1 _08882_ (.A1(_03278_),
    .A2(_03302_),
    .Y(_03304_),
    .B1(_03303_));
 sg13g2_buf_1 _08883_ (.A(\dtop.vtop.pipeline.zg[9] ),
    .X(_03305_));
 sg13g2_inv_1 _08884_ (.Y(_03306_),
    .A(_03305_));
 sg13g2_buf_1 _08885_ (.A(\dtop.vtop.pipeline.z[12] ),
    .X(_03307_));
 sg13g2_inv_1 _08886_ (.Y(_03308_),
    .A(_03307_));
 sg13g2_buf_2 _08887_ (.A(\dtop.vtop.pipeline.zg[7] ),
    .X(_03309_));
 sg13g2_buf_1 _08888_ (.A(\dtop.vtop.pipeline.z[13] ),
    .X(_03310_));
 sg13g2_buf_2 _08889_ (.A(\dtop.vtop.pipeline.zg[8] ),
    .X(_03311_));
 sg13g2_nor2b_1 _08890_ (.A(_03310_),
    .B_N(_03311_),
    .Y(_03312_));
 sg13g2_a21oi_1 _08891_ (.A1(_03308_),
    .A2(_03309_),
    .Y(_03313_),
    .B1(_03312_));
 sg13g2_nand2_1 _08892_ (.Y(_03314_),
    .A(_03306_),
    .B(_03313_));
 sg13g2_nand2_1 _08893_ (.Y(_03315_),
    .A(\dtop.vtop.pipeline.z[14] ),
    .B(_03313_));
 sg13g2_a22oi_1 _08894_ (.Y(_03316_),
    .B1(_03314_),
    .B2(_03315_),
    .A2(_03304_),
    .A1(_03301_));
 sg13g2_buf_2 _08895_ (.A(_03316_),
    .X(_03317_));
 sg13g2_inv_1 _08896_ (.Y(_03318_),
    .A(\dtop.vtop.pipeline.z[14] ));
 sg13g2_nand2b_1 _08897_ (.Y(_03319_),
    .B(_03307_),
    .A_N(_03309_));
 sg13g2_nand2b_1 _08898_ (.Y(_03320_),
    .B(_03310_),
    .A_N(_03311_));
 sg13g2_o21ai_1 _08899_ (.B1(_03320_),
    .Y(_03321_),
    .A1(_03312_),
    .A2(_03319_));
 sg13g2_o21ai_1 _08900_ (.B1(_03321_),
    .Y(_03322_),
    .A1(\dtop.vtop.pipeline.z[14] ),
    .A2(_03306_));
 sg13g2_o21ai_1 _08901_ (.B1(_03322_),
    .Y(_03323_),
    .A1(_03318_),
    .A2(_03305_));
 sg13g2_buf_2 _08902_ (.A(_03323_),
    .X(_03324_));
 sg13g2_or2_1 _08903_ (.X(_03325_),
    .B(_03324_),
    .A(_03317_));
 sg13g2_buf_2 _08904_ (.A(_03325_),
    .X(_03326_));
 sg13g2_nand3_1 _08905_ (.B(_03273_),
    .C(_03326_),
    .A(\dtop.vtop.pipeline.zg_valid ),
    .Y(_03327_));
 sg13g2_buf_1 _08906_ (.A(_03327_),
    .X(_03328_));
 sg13g2_nand2_1 _08907_ (.Y(_03329_),
    .A(_03271_),
    .B(_03328_));
 sg13g2_buf_1 _08908_ (.A(_03329_),
    .X(_03330_));
 sg13g2_buf_1 _08909_ (.A(net112),
    .X(_03331_));
 sg13g2_nand2_1 _08910_ (.Y(_03332_),
    .A(net98),
    .B(net120));
 sg13g2_nand2_1 _08911_ (.Y(_03333_),
    .A(net97),
    .B(net115));
 sg13g2_nand2_1 _08912_ (.Y(_03334_),
    .A(_03332_),
    .B(_03333_));
 sg13g2_inv_1 _08913_ (.Y(_03335_),
    .A(\dtop.vtop.pipeline.cosappr_acc[1] ));
 sg13g2_buf_1 _08914_ (.A(\dtop.vtop.pipeline.cosappr_acc[0] ),
    .X(_03336_));
 sg13g2_xnor2_1 _08915_ (.Y(_03337_),
    .A(net97),
    .B(net165));
 sg13g2_buf_2 _08916_ (.A(_03337_),
    .X(_03338_));
 sg13g2_a21oi_1 _08917_ (.A1(_03336_),
    .A2(_03338_),
    .Y(_03339_),
    .B1(_02477_));
 sg13g2_nand3_1 _08918_ (.B(_02477_),
    .C(_03338_),
    .A(_03336_),
    .Y(_03340_));
 sg13g2_o21ai_1 _08919_ (.B1(_03340_),
    .Y(_03341_),
    .A1(_03335_),
    .A2(_03339_));
 sg13g2_buf_1 _08920_ (.A(_03341_),
    .X(_03342_));
 sg13g2_xnor2_1 _08921_ (.Y(_03343_),
    .A(net97),
    .B(net116));
 sg13g2_buf_1 _08922_ (.A(_03343_),
    .X(_03344_));
 sg13g2_nand2_1 _08923_ (.Y(_03345_),
    .A(_03342_),
    .B(_03344_));
 sg13g2_o21ai_1 _08924_ (.B1(\dtop.vtop.pipeline.cosappr_acc[2] ),
    .Y(_03346_),
    .A1(_03342_),
    .A2(_03344_));
 sg13g2_nor2_1 _08925_ (.A(_02249_),
    .B(_02250_),
    .Y(_03347_));
 sg13g2_a21oi_1 _08926_ (.A1(_03345_),
    .A2(_03346_),
    .Y(_03348_),
    .B1(_03347_));
 sg13g2_xnor2_1 _08927_ (.Y(_03349_),
    .A(_03334_),
    .B(_03348_));
 sg13g2_nand2_1 _08928_ (.Y(_03350_),
    .A(_02846_),
    .B(_02251_));
 sg13g2_buf_1 _08929_ (.A(_03350_),
    .X(_03351_));
 sg13g2_nand2_1 _08930_ (.Y(_03352_),
    .A(\dtop.vtop.pipeline.cosappr_acc[3] ),
    .B(net306));
 sg13g2_xnor2_1 _08931_ (.Y(_03353_),
    .A(_03349_),
    .B(_03352_));
 sg13g2_buf_1 _08932_ (.A(\dtop.vtop.color[6] ),
    .X(_03354_));
 sg13g2_nand2_1 _08933_ (.Y(_03355_),
    .A(_03354_),
    .B(net96));
 sg13g2_o21ai_1 _08934_ (.B1(_03355_),
    .Y(_00207_),
    .A1(net96),
    .A2(_03353_));
 sg13g2_buf_1 _08935_ (.A(\dtop.vtop.color[7] ),
    .X(_03356_));
 sg13g2_inv_1 _08936_ (.Y(_03357_),
    .A(_03356_));
 sg13g2_nand2b_1 _08937_ (.Y(_03358_),
    .B(_02250_),
    .A_N(_03270_));
 sg13g2_buf_1 _08938_ (.A(_03358_),
    .X(_03359_));
 sg13g2_buf_1 _08939_ (.A(_03326_),
    .X(_03360_));
 sg13g2_and3_1 _08940_ (.X(_03361_),
    .A(\dtop.vtop.pipeline.zg_valid ),
    .B(_03273_),
    .C(_03360_));
 sg13g2_buf_1 _08941_ (.A(_03361_),
    .X(_03362_));
 sg13g2_nor2_1 _08942_ (.A(_03359_),
    .B(_03362_),
    .Y(_03363_));
 sg13g2_buf_1 _08943_ (.A(_03363_),
    .X(_03364_));
 sg13g2_buf_1 _08944_ (.A(net95),
    .X(_03365_));
 sg13g2_buf_1 _08945_ (.A(_03347_),
    .X(_03366_));
 sg13g2_buf_1 _08946_ (.A(\dtop.vtop.pipeline.cosappr_acc[4] ),
    .X(_03367_));
 sg13g2_a221oi_1 _08947_ (.B2(_03346_),
    .C1(net338),
    .B1(_03345_),
    .A1(_03332_),
    .Y(_03368_),
    .A2(_03333_));
 sg13g2_o21ai_1 _08948_ (.B1(\dtop.vtop.pipeline.cosappr_acc[3] ),
    .Y(_03369_),
    .A1(_03334_),
    .A2(_03348_));
 sg13g2_nand2b_1 _08949_ (.Y(_03370_),
    .B(_03369_),
    .A_N(_03368_));
 sg13g2_xnor2_1 _08950_ (.Y(_03371_),
    .A(_03367_),
    .B(_03370_));
 sg13g2_nor2_1 _08951_ (.A(net338),
    .B(_03371_),
    .Y(_03372_));
 sg13g2_xnor2_1 _08952_ (.Y(_03373_),
    .A(_02796_),
    .B(_03372_));
 sg13g2_nand2_1 _08953_ (.Y(_03374_),
    .A(net84),
    .B(_03373_));
 sg13g2_o21ai_1 _08954_ (.B1(_03374_),
    .Y(_00208_),
    .A1(_03357_),
    .A2(net84));
 sg13g2_nor2_1 _08955_ (.A(_03367_),
    .B(_02817_),
    .Y(_03375_));
 sg13g2_o21ai_1 _08956_ (.B1(_03367_),
    .Y(_03376_),
    .A1(_02817_),
    .A2(_03368_));
 sg13g2_o21ai_1 _08957_ (.B1(_03376_),
    .Y(_03377_),
    .A1(_03369_),
    .A2(_03375_));
 sg13g2_and2_1 _08958_ (.A(_02817_),
    .B(_03368_),
    .X(_03378_));
 sg13g2_a21o_1 _08959_ (.A2(_03377_),
    .A1(_03351_),
    .B1(_03378_),
    .X(_03379_));
 sg13g2_buf_1 _08960_ (.A(_03379_),
    .X(_03380_));
 sg13g2_xnor2_1 _08961_ (.Y(_03381_),
    .A(_02950_),
    .B(_03380_));
 sg13g2_nand2_1 _08962_ (.Y(_03382_),
    .A(\dtop.vtop.pipeline.cosappr_acc[5] ),
    .B(net306));
 sg13g2_xor2_1 _08963_ (.B(_03382_),
    .A(_03381_),
    .X(_03383_));
 sg13g2_buf_1 _08964_ (.A(\dtop.vtop.color[8] ),
    .X(_03384_));
 sg13g2_nand2_1 _08965_ (.Y(_03385_),
    .A(_03384_),
    .B(net96));
 sg13g2_o21ai_1 _08966_ (.B1(_03385_),
    .Y(_00209_),
    .A1(_03331_),
    .A2(_03383_));
 sg13g2_inv_1 _08967_ (.Y(_03386_),
    .A(\dtop.vtop.color[9] ));
 sg13g2_o21ai_1 _08968_ (.B1(\dtop.vtop.pipeline.cosappr_acc[5] ),
    .Y(_03387_),
    .A1(_02962_),
    .A2(_03380_));
 sg13g2_nand2_1 _08969_ (.Y(_03388_),
    .A(_02962_),
    .B(_03380_));
 sg13g2_nand2_1 _08970_ (.Y(_03389_),
    .A(_03387_),
    .B(_03388_));
 sg13g2_xnor2_1 _08971_ (.Y(_03390_),
    .A(\dtop.vtop.pipeline.cosappr_acc[6] ),
    .B(_03389_));
 sg13g2_nor2_1 _08972_ (.A(_03366_),
    .B(_03390_),
    .Y(_03391_));
 sg13g2_xnor2_1 _08973_ (.Y(_03392_),
    .A(_03201_),
    .B(_03391_));
 sg13g2_nand2_1 _08974_ (.Y(_03393_),
    .A(net95),
    .B(_03392_));
 sg13g2_o21ai_1 _08975_ (.B1(_03393_),
    .Y(_00210_),
    .A1(_03386_),
    .A2(_03365_));
 sg13g2_a21oi_1 _08976_ (.A1(net306),
    .A2(_03389_),
    .Y(_03394_),
    .B1(_03203_));
 sg13g2_a21oi_1 _08977_ (.A1(_03203_),
    .A2(_03389_),
    .Y(_03395_),
    .B1(\dtop.vtop.pipeline.cosappr_acc[6] ));
 sg13g2_nor3_1 _08978_ (.A(_03366_),
    .B(_03394_),
    .C(_03395_),
    .Y(_03396_));
 sg13g2_nand2_1 _08979_ (.Y(_03397_),
    .A(\dtop.vtop.pipeline.cosappr_acc[7] ),
    .B(_03396_));
 sg13g2_a21o_1 _08980_ (.A2(net306),
    .A1(\dtop.vtop.pipeline.cosappr_acc[7] ),
    .B1(_03396_),
    .X(_03398_));
 sg13g2_nand2_1 _08981_ (.Y(_03399_),
    .A(_03397_),
    .B(_03398_));
 sg13g2_buf_2 _08982_ (.A(\dtop.vtop.color[10] ),
    .X(_03400_));
 sg13g2_nand2_1 _08983_ (.Y(_03401_),
    .A(_03400_),
    .B(_03331_));
 sg13g2_o21ai_1 _08984_ (.B1(_03401_),
    .Y(_00211_),
    .A1(net96),
    .A2(_03399_));
 sg13g2_xor2_1 _08985_ (.B(_03397_),
    .A(\dtop.vtop.pipeline.cosappr_acc[8] ),
    .X(_03402_));
 sg13g2_nor2_1 _08986_ (.A(net338),
    .B(_03402_),
    .Y(_03403_));
 sg13g2_mux2_1 _08987_ (.A0(\dtop.vtop.color[11] ),
    .A1(_03403_),
    .S(_03365_),
    .X(_00212_));
 sg13g2_buf_1 _08988_ (.A(\dtop.vtop.pipeline.nstep_zg[0] ),
    .X(_03404_));
 sg13g2_buf_1 _08989_ (.A(_03404_),
    .X(_03405_));
 sg13g2_buf_1 _08990_ (.A(\dtop.vtop.pipeline.nstep[0] ),
    .X(_03406_));
 sg13g2_buf_1 _08991_ (.A(net406),
    .X(_03407_));
 sg13g2_buf_1 _08992_ (.A(net268),
    .X(_03408_));
 sg13g2_nor2_1 _08993_ (.A(net252),
    .B(_03330_),
    .Y(_03409_));
 sg13g2_mux2_1 _08994_ (.A0(net368),
    .A1(_03407_),
    .S(_03409_),
    .X(_00248_));
 sg13g2_buf_1 _08995_ (.A(\dtop.vtop.pipeline.nstep_zg[1] ),
    .X(_03410_));
 sg13g2_buf_1 _08996_ (.A(net405),
    .X(_03411_));
 sg13g2_buf_2 _08997_ (.A(\dtop.vtop.pipeline.nstep[1] ),
    .X(_03412_));
 sg13g2_buf_1 _08998_ (.A(_03412_),
    .X(_03413_));
 sg13g2_mux2_1 _08999_ (.A0(_03411_),
    .A1(net365),
    .S(_03409_),
    .X(_00249_));
 sg13g2_nand2_1 _09000_ (.Y(_03414_),
    .A(_05282_),
    .B(_01450_));
 sg13g2_nand2_1 _09001_ (.Y(_03415_),
    .A(net278),
    .B(net338));
 sg13g2_and2_1 _09002_ (.A(_03414_),
    .B(_03415_),
    .X(_03416_));
 sg13g2_buf_1 _09003_ (.A(_03416_),
    .X(_03417_));
 sg13g2_buf_1 _09004_ (.A(net278),
    .X(_03418_));
 sg13g2_inv_1 _09005_ (.Y(_03419_),
    .A(\dtop.vtop.pipeline.phases[2][0] ));
 sg13g2_mux2_1 _09006_ (.A0(_03419_),
    .A1(_00030_),
    .S(net269),
    .X(_03420_));
 sg13g2_nor2_1 _09007_ (.A(_02257_),
    .B(_02340_),
    .Y(_03421_));
 sg13g2_nand2b_1 _09008_ (.Y(_03422_),
    .B(_05185_),
    .A_N(_05194_));
 sg13g2_nor4_1 _09009_ (.A(_05170_),
    .B(_05173_),
    .C(_05175_),
    .D(_03422_),
    .Y(_03423_));
 sg13g2_a21o_1 _09010_ (.A2(_03421_),
    .A1(_05178_),
    .B1(_03423_),
    .X(_03424_));
 sg13g2_buf_1 _09011_ (.A(_03424_),
    .X(_03425_));
 sg13g2_nand2_1 _09012_ (.Y(_03426_),
    .A(\dtop.vtop.pipeline.phases[1][0] ),
    .B(net266));
 sg13g2_o21ai_1 _09013_ (.B1(_03426_),
    .Y(_03427_),
    .A1(net270),
    .A2(_03420_));
 sg13g2_buf_2 _09014_ (.A(_03427_),
    .X(_03428_));
 sg13g2_inv_1 _09015_ (.Y(_03429_),
    .A(\dtop.vtop.pipeline.nstep[0] ));
 sg13g2_buf_1 _09016_ (.A(_03429_),
    .X(_03430_));
 sg13g2_nand2b_1 _09017_ (.Y(_03431_),
    .B(net266),
    .A_N(\dtop.vtop.dphases[1][0] ));
 sg13g2_nand2b_1 _09018_ (.Y(_03432_),
    .B(net275),
    .A_N(\dtop.vtop.dphases[2][0] ));
 sg13g2_a21oi_1 _09019_ (.A1(_05178_),
    .A2(_03421_),
    .Y(_03433_),
    .B1(_03423_));
 sg13g2_nand3_1 _09020_ (.B(_02469_),
    .C(_03433_),
    .A(_00032_),
    .Y(_03434_));
 sg13g2_and3_1 _09021_ (.X(_03435_),
    .A(_03431_),
    .B(_03432_),
    .C(_03434_));
 sg13g2_buf_1 _09022_ (.A(_03435_),
    .X(_03436_));
 sg13g2_nand3_1 _09023_ (.B(_00031_),
    .C(_03436_),
    .A(_03430_),
    .Y(_03437_));
 sg13g2_xnor2_1 _09024_ (.Y(_03438_),
    .A(_03428_),
    .B(_03437_));
 sg13g2_nand2_1 _09025_ (.Y(_03439_),
    .A(net267),
    .B(_03438_));
 sg13g2_nand2_1 _09026_ (.Y(_03440_),
    .A(\dtop.vtop.pipeline.phases[0][0] ),
    .B(_03417_));
 sg13g2_o21ai_1 _09027_ (.B1(_03440_),
    .Y(_00250_),
    .A1(_03417_),
    .A2(_03439_));
 sg13g2_nand2_1 _09028_ (.Y(_03441_),
    .A(_03414_),
    .B(_03415_));
 sg13g2_buf_1 _09029_ (.A(_03441_),
    .X(_03442_));
 sg13g2_nor2_1 _09030_ (.A(net275),
    .B(net266),
    .Y(_03443_));
 sg13g2_buf_2 _09031_ (.A(_03443_),
    .X(_03444_));
 sg13g2_buf_1 _09032_ (.A(_03425_),
    .X(_03445_));
 sg13g2_nand2b_1 _09033_ (.Y(_03446_),
    .B(net251),
    .A_N(\dtop.vtop.dphases[1][5] ));
 sg13g2_o21ai_1 _09034_ (.B1(_03446_),
    .Y(_03447_),
    .A1(\dtop.vtop.dphases[2][5] ),
    .A2(net255));
 sg13g2_a21oi_1 _09035_ (.A1(_00042_),
    .A2(_03444_),
    .Y(_03448_),
    .B1(_03447_));
 sg13g2_nand2b_1 _09036_ (.Y(_03449_),
    .B(net251),
    .A_N(\dtop.vtop.dphases[1][6] ));
 sg13g2_o21ai_1 _09037_ (.B1(_03449_),
    .Y(_03450_),
    .A1(\dtop.vtop.dphases[2][6] ),
    .A2(net255));
 sg13g2_a21oi_1 _09038_ (.A1(_00043_),
    .A2(_03444_),
    .Y(_03451_),
    .B1(_03450_));
 sg13g2_mux2_1 _09039_ (.A0(_03448_),
    .A1(_03451_),
    .S(net364),
    .X(_03452_));
 sg13g2_nand2b_1 _09040_ (.Y(_03453_),
    .B(net251),
    .A_N(\dtop.vtop.dphases[1][8] ));
 sg13g2_o21ai_1 _09041_ (.B1(_03453_),
    .Y(_03454_),
    .A1(\dtop.vtop.dphases[2][8] ),
    .A2(net255));
 sg13g2_a21o_1 _09042_ (.A2(_03444_),
    .A1(_00048_),
    .B1(_03454_),
    .X(_03455_));
 sg13g2_nand2b_1 _09043_ (.Y(_03456_),
    .B(net251),
    .A_N(\dtop.vtop.dphases[1][7] ));
 sg13g2_o21ai_1 _09044_ (.B1(_03456_),
    .Y(_03457_),
    .A1(\dtop.vtop.dphases[2][7] ),
    .A2(net255));
 sg13g2_a21o_1 _09045_ (.A2(_03444_),
    .A1(_00045_),
    .B1(_03457_),
    .X(_03458_));
 sg13g2_or2_1 _09046_ (.X(_03459_),
    .B(_03458_),
    .A(net364));
 sg13g2_o21ai_1 _09047_ (.B1(_03459_),
    .Y(_03460_),
    .A1(net406),
    .A2(_03455_));
 sg13g2_inv_2 _09048_ (.Y(_03461_),
    .A(_03412_));
 sg13g2_mux2_1 _09049_ (.A0(_03452_),
    .A1(_03460_),
    .S(_03461_),
    .X(_03462_));
 sg13g2_nor2_1 _09050_ (.A(net151),
    .B(_03462_),
    .Y(_03463_));
 sg13g2_nor2_1 _09051_ (.A(_00039_),
    .B(net254),
    .Y(_03464_));
 sg13g2_a21oi_1 _09052_ (.A1(\dtop.vtop.pipeline.phases[2][4] ),
    .A2(net254),
    .Y(_03465_),
    .B1(_03464_));
 sg13g2_nand2_1 _09053_ (.Y(_03466_),
    .A(\dtop.vtop.pipeline.phases[1][4] ),
    .B(net251));
 sg13g2_o21ai_1 _09054_ (.B1(_03466_),
    .Y(_03467_),
    .A1(net270),
    .A2(_03465_));
 sg13g2_buf_1 _09055_ (.A(_03467_),
    .X(_03468_));
 sg13g2_a22oi_1 _09056_ (.Y(_03469_),
    .B1(net266),
    .B2(_03241_),
    .A2(net275),
    .A1(_03258_));
 sg13g2_nand3_1 _09057_ (.B(_02469_),
    .C(_03433_),
    .A(_00034_),
    .Y(_03470_));
 sg13g2_nand2_1 _09058_ (.Y(_03471_),
    .A(_03469_),
    .B(_03470_));
 sg13g2_a22oi_1 _09059_ (.Y(_03472_),
    .B1(net266),
    .B2(_03243_),
    .A2(net275),
    .A1(_03260_));
 sg13g2_nand3_1 _09060_ (.B(net255),
    .C(_03433_),
    .A(_00036_),
    .Y(_03473_));
 sg13g2_nand3_1 _09061_ (.B(_03472_),
    .C(_03473_),
    .A(_03429_),
    .Y(_03474_));
 sg13g2_o21ai_1 _09062_ (.B1(_03474_),
    .Y(_03475_),
    .A1(_03429_),
    .A2(_03471_));
 sg13g2_nand3_1 _09063_ (.B(_03432_),
    .C(_03434_),
    .A(_03431_),
    .Y(_03476_));
 sg13g2_o21ai_1 _09064_ (.B1(_03412_),
    .Y(_03477_),
    .A1(_03406_),
    .A2(_03476_));
 sg13g2_o21ai_1 _09065_ (.B1(_03477_),
    .Y(_03478_),
    .A1(_03412_),
    .A2(_03475_));
 sg13g2_nor2_1 _09066_ (.A(_00035_),
    .B(net254),
    .Y(_03479_));
 sg13g2_a21oi_1 _09067_ (.A1(\dtop.vtop.pipeline.phases[2][2] ),
    .A2(net254),
    .Y(_03480_),
    .B1(_03479_));
 sg13g2_nand2_1 _09068_ (.Y(_03481_),
    .A(\dtop.vtop.pipeline.phases[1][2] ),
    .B(net251));
 sg13g2_o21ai_1 _09069_ (.B1(_03481_),
    .Y(_03482_),
    .A1(net270),
    .A2(_03480_));
 sg13g2_inv_1 _09070_ (.Y(_03483_),
    .A(_03482_));
 sg13g2_nor2_1 _09071_ (.A(_03478_),
    .B(_03483_),
    .Y(_03484_));
 sg13g2_inv_1 _09072_ (.Y(_03485_),
    .A(_00033_));
 sg13g2_mux2_1 _09073_ (.A0(\dtop.vtop.pipeline.phases[2][1] ),
    .A1(_03485_),
    .S(net269),
    .X(_03486_));
 sg13g2_a22oi_1 _09074_ (.Y(_03487_),
    .B1(_03486_),
    .B2(_02454_),
    .A2(net266),
    .A1(\dtop.vtop.pipeline.phases[1][1] ));
 sg13g2_nor2_1 _09075_ (.A(_03476_),
    .B(_03487_),
    .Y(_03488_));
 sg13g2_o21ai_1 _09076_ (.B1(_03488_),
    .Y(_03489_),
    .A1(_03406_),
    .A2(_03428_));
 sg13g2_nand2_1 _09077_ (.Y(_03490_),
    .A(_03428_),
    .B(_03436_));
 sg13g2_nand3_1 _09078_ (.B(_03469_),
    .C(_03470_),
    .A(net364),
    .Y(_03491_));
 sg13g2_a21o_1 _09079_ (.A2(_03490_),
    .A1(_03487_),
    .B1(_03491_),
    .X(_03492_));
 sg13g2_inv_1 _09080_ (.Y(_03493_),
    .A(_00031_));
 sg13g2_a221oi_1 _09081_ (.B2(_03492_),
    .C1(_03493_),
    .B1(_03489_),
    .A1(_03478_),
    .Y(_03494_),
    .A2(_03483_));
 sg13g2_nor2_1 _09082_ (.A(_00037_),
    .B(net254),
    .Y(_03495_));
 sg13g2_a21oi_1 _09083_ (.A1(\dtop.vtop.pipeline.phases[2][3] ),
    .A2(net254),
    .Y(_03496_),
    .B1(_03495_));
 sg13g2_nand2_1 _09084_ (.Y(_03497_),
    .A(\dtop.vtop.pipeline.phases[1][3] ),
    .B(_03445_));
 sg13g2_o21ai_1 _09085_ (.B1(_03497_),
    .Y(_03498_),
    .A1(net270),
    .A2(_03496_));
 sg13g2_o21ai_1 _09086_ (.B1(_03498_),
    .Y(_03499_),
    .A1(_03484_),
    .A2(_03494_));
 sg13g2_nand2b_1 _09087_ (.Y(_03500_),
    .B(net266),
    .A_N(\dtop.vtop.dphases[1][3] ));
 sg13g2_o21ai_1 _09088_ (.B1(_03500_),
    .Y(_03501_),
    .A1(\dtop.vtop.dphases[2][3] ),
    .A2(net255));
 sg13g2_a21oi_1 _09089_ (.A1(_00038_),
    .A2(_03444_),
    .Y(_03502_),
    .B1(_03501_));
 sg13g2_and3_1 _09090_ (.X(_03503_),
    .A(net406),
    .B(_03472_),
    .C(_03473_));
 sg13g2_a21o_1 _09091_ (.A2(_03502_),
    .A1(net364),
    .B1(_03503_),
    .X(_03504_));
 sg13g2_nand2_1 _09092_ (.Y(_03505_),
    .A(net406),
    .B(_03436_));
 sg13g2_nand3_1 _09093_ (.B(_03491_),
    .C(_03505_),
    .A(_03412_),
    .Y(_03506_));
 sg13g2_o21ai_1 _09094_ (.B1(_03506_),
    .Y(_03507_),
    .A1(_03412_),
    .A2(_03504_));
 sg13g2_nor3_1 _09095_ (.A(_03484_),
    .B(_03494_),
    .C(_03498_),
    .Y(_03508_));
 sg13g2_a21oi_2 _09096_ (.B1(_03508_),
    .Y(_03509_),
    .A2(_03507_),
    .A1(_03499_));
 sg13g2_nand2b_1 _09097_ (.Y(_03510_),
    .B(net266),
    .A_N(\dtop.vtop.dphases[1][4] ));
 sg13g2_o21ai_1 _09098_ (.B1(_03510_),
    .Y(_03511_),
    .A1(\dtop.vtop.dphases[2][4] ),
    .A2(_02508_));
 sg13g2_a21oi_1 _09099_ (.A1(_00040_),
    .A2(_03444_),
    .Y(_03512_),
    .B1(_03511_));
 sg13g2_and2_1 _09100_ (.A(net406),
    .B(_03502_),
    .X(_03513_));
 sg13g2_a21oi_1 _09101_ (.A1(net364),
    .A2(_03512_),
    .Y(_03514_),
    .B1(_03513_));
 sg13g2_nor2_1 _09102_ (.A(_03461_),
    .B(_03475_),
    .Y(_03515_));
 sg13g2_a21o_1 _09103_ (.A2(_03514_),
    .A1(_03461_),
    .B1(_03515_),
    .X(_03516_));
 sg13g2_inv_1 _09104_ (.Y(_03517_),
    .A(_03516_));
 sg13g2_a21oi_1 _09105_ (.A1(_03468_),
    .A2(_03509_),
    .Y(_03518_),
    .B1(_03517_));
 sg13g2_nor2_1 _09106_ (.A(_03412_),
    .B(_03452_),
    .Y(_03519_));
 sg13g2_a21o_1 _09107_ (.A2(_03514_),
    .A1(_03412_),
    .B1(_03519_),
    .X(_03520_));
 sg13g2_buf_1 _09108_ (.A(_03520_),
    .X(_03521_));
 sg13g2_mux2_1 _09109_ (.A0(_03448_),
    .A1(_03512_),
    .S(net406),
    .X(_03522_));
 sg13g2_mux2_1 _09110_ (.A0(_03504_),
    .A1(_03522_),
    .S(_03461_),
    .X(_03523_));
 sg13g2_buf_1 _09111_ (.A(_03523_),
    .X(_03524_));
 sg13g2_inv_1 _09112_ (.Y(_03525_),
    .A(_03524_));
 sg13g2_nand2_1 _09113_ (.Y(_03526_),
    .A(\dtop.vtop.pipeline.phases[2][5] ),
    .B(_03169_));
 sg13g2_o21ai_1 _09114_ (.B1(_03526_),
    .Y(_03527_),
    .A1(_00041_),
    .A2(_03169_));
 sg13g2_a22oi_1 _09115_ (.Y(_03528_),
    .B1(_03527_),
    .B2(_02454_),
    .A2(_03445_),
    .A1(\dtop.vtop.pipeline.phases[1][5] ));
 sg13g2_buf_1 _09116_ (.A(_03528_),
    .X(_03529_));
 sg13g2_a22oi_1 _09117_ (.Y(_03530_),
    .B1(_03525_),
    .B2(_03529_),
    .A2(_03521_),
    .A1(net119));
 sg13g2_o21ai_1 _09118_ (.B1(_03530_),
    .Y(_03531_),
    .A1(_03468_),
    .A2(_03509_));
 sg13g2_nand2_1 _09119_ (.Y(_03532_),
    .A(net119),
    .B(_03521_));
 sg13g2_nor2_1 _09120_ (.A(_03525_),
    .B(_03529_),
    .Y(_03533_));
 sg13g2_nor2_1 _09121_ (.A(net119),
    .B(_03521_),
    .Y(_03534_));
 sg13g2_a21oi_1 _09122_ (.A1(_03532_),
    .A2(_03533_),
    .Y(_03535_),
    .B1(_03534_));
 sg13g2_o21ai_1 _09123_ (.B1(_03535_),
    .Y(_03536_),
    .A1(_03518_),
    .A2(_03531_));
 sg13g2_nand2_1 _09124_ (.Y(_03537_),
    .A(net406),
    .B(_03451_));
 sg13g2_o21ai_1 _09125_ (.B1(_03537_),
    .Y(_03538_),
    .A1(net406),
    .A2(_03458_));
 sg13g2_or2_1 _09126_ (.X(_03539_),
    .B(_03522_),
    .A(_03461_));
 sg13g2_o21ai_1 _09127_ (.B1(_03539_),
    .Y(_03540_),
    .A1(net365),
    .A2(_03538_));
 sg13g2_nand2_1 _09128_ (.Y(_03541_),
    .A(net145),
    .B(_03540_));
 sg13g2_nor2_1 _09129_ (.A(net145),
    .B(_03540_),
    .Y(_03542_));
 sg13g2_a221oi_1 _09130_ (.B2(_03541_),
    .C1(_03542_),
    .B1(_03536_),
    .A1(net151),
    .Y(_03543_),
    .A2(_03462_));
 sg13g2_nand2b_1 _09131_ (.Y(_03544_),
    .B(net251),
    .A_N(\dtop.vtop.dphases[1][9] ));
 sg13g2_o21ai_1 _09132_ (.B1(_03544_),
    .Y(_03545_),
    .A1(\dtop.vtop.dphases[2][9] ),
    .A2(net255));
 sg13g2_a21o_1 _09133_ (.A2(_03444_),
    .A1(_00050_),
    .B1(_03545_),
    .X(_03546_));
 sg13g2_or2_1 _09134_ (.X(_03547_),
    .B(_03455_),
    .A(net364));
 sg13g2_o21ai_1 _09135_ (.B1(_03547_),
    .Y(_03548_),
    .A1(_03407_),
    .A2(_03546_));
 sg13g2_or2_1 _09136_ (.X(_03549_),
    .B(_03538_),
    .A(_03461_));
 sg13g2_o21ai_1 _09137_ (.B1(_03549_),
    .Y(_03550_),
    .A1(net365),
    .A2(_03548_));
 sg13g2_buf_2 _09138_ (.A(_03550_),
    .X(_03551_));
 sg13g2_nor3_1 _09139_ (.A(_03463_),
    .B(_03543_),
    .C(_03551_),
    .Y(_03552_));
 sg13g2_o21ai_1 _09140_ (.B1(_03551_),
    .Y(_03553_),
    .A1(_03463_),
    .A2(_03543_));
 sg13g2_o21ai_1 _09141_ (.B1(_03553_),
    .Y(_03554_),
    .A1(net116),
    .A2(_03552_));
 sg13g2_nand2b_1 _09142_ (.Y(_03555_),
    .B(net251),
    .A_N(\dtop.vtop.dphases[1][10] ));
 sg13g2_o21ai_1 _09143_ (.B1(_03555_),
    .Y(_03556_),
    .A1(\dtop.vtop.dphases[2][10] ),
    .A2(net255));
 sg13g2_a21o_1 _09144_ (.A2(_03444_),
    .A1(_00052_),
    .B1(_03556_),
    .X(_03557_));
 sg13g2_buf_1 _09145_ (.A(_03557_),
    .X(_03558_));
 sg13g2_mux2_1 _09146_ (.A0(_03546_),
    .A1(_03558_),
    .S(net364),
    .X(_03559_));
 sg13g2_nand2_1 _09147_ (.Y(_03560_),
    .A(net365),
    .B(_03460_));
 sg13g2_o21ai_1 _09148_ (.B1(_03560_),
    .Y(_03561_),
    .A1(net365),
    .A2(_03559_));
 sg13g2_buf_2 _09149_ (.A(_03561_),
    .X(_03562_));
 sg13g2_xnor2_1 _09150_ (.Y(_03563_),
    .A(net120),
    .B(_03562_));
 sg13g2_xnor2_1 _09151_ (.Y(_03564_),
    .A(_03554_),
    .B(_03563_));
 sg13g2_buf_1 _09152_ (.A(_05179_),
    .X(_03565_));
 sg13g2_nand2_1 _09153_ (.Y(_03566_),
    .A(_05353_),
    .B(_05358_));
 sg13g2_xnor2_1 _09154_ (.Y(_03567_),
    .A(_00755_),
    .B(_03566_));
 sg13g2_nor2_1 _09155_ (.A(net262),
    .B(_03567_),
    .Y(_03568_));
 sg13g2_xnor2_1 _09156_ (.Y(_03569_),
    .A(_05374_),
    .B(_03568_));
 sg13g2_nor2_1 _09157_ (.A(_03565_),
    .B(_03569_),
    .Y(_03570_));
 sg13g2_a21oi_1 _09158_ (.A1(net267),
    .A2(_03564_),
    .Y(_03571_),
    .B1(_03570_));
 sg13g2_buf_1 _09159_ (.A(_03441_),
    .X(_03572_));
 sg13g2_nor2_1 _09160_ (.A(\dtop.vtop.pipeline.phases[0][10] ),
    .B(_03572_),
    .Y(_03573_));
 sg13g2_a21oi_1 _09161_ (.A1(net238),
    .A2(_03571_),
    .Y(_00251_),
    .B1(_03573_));
 sg13g2_nand2_1 _09162_ (.Y(_03574_),
    .A(net115),
    .B(_03562_));
 sg13g2_nor2_1 _09163_ (.A(net115),
    .B(_03562_),
    .Y(_03575_));
 sg13g2_a21oi_1 _09164_ (.A1(_03554_),
    .A2(_03574_),
    .Y(_03576_),
    .B1(_03575_));
 sg13g2_nor2_1 _09165_ (.A(net365),
    .B(_03558_),
    .Y(_03577_));
 sg13g2_a21oi_1 _09166_ (.A1(net365),
    .A2(_03548_),
    .Y(_03578_),
    .B1(_03577_));
 sg13g2_xnor2_1 _09167_ (.Y(_03579_),
    .A(net121),
    .B(_03578_));
 sg13g2_xnor2_1 _09168_ (.Y(_03580_),
    .A(_03576_),
    .B(_03579_));
 sg13g2_a21o_1 _09169_ (.A2(_03566_),
    .A1(_05374_),
    .B1(net384),
    .X(_03581_));
 sg13g2_o21ai_1 _09170_ (.B1(_03581_),
    .Y(_03582_),
    .A1(_05374_),
    .A2(_03566_));
 sg13g2_xnor2_1 _09171_ (.Y(_03583_),
    .A(_05360_),
    .B(_03582_));
 sg13g2_nor2_1 _09172_ (.A(net262),
    .B(_03583_),
    .Y(_03584_));
 sg13g2_xnor2_1 _09173_ (.Y(_03585_),
    .A(_05363_),
    .B(_03584_));
 sg13g2_nand2_1 _09174_ (.Y(_03586_),
    .A(net268),
    .B(_03585_));
 sg13g2_o21ai_1 _09175_ (.B1(_03586_),
    .Y(_03587_),
    .A1(net252),
    .A2(_03580_));
 sg13g2_mux2_1 _09176_ (.A0(\dtop.vtop.pipeline.phases[0][11] ),
    .A1(_03587_),
    .S(net238),
    .X(_00252_));
 sg13g2_nor2_1 _09177_ (.A(_03463_),
    .B(_03543_),
    .Y(_03588_));
 sg13g2_buf_2 _09178_ (.A(_03588_),
    .X(_03589_));
 sg13g2_a21o_1 _09179_ (.A2(_03548_),
    .A1(_03413_),
    .B1(_03577_),
    .X(_03590_));
 sg13g2_buf_1 _09180_ (.A(_03590_),
    .X(_03591_));
 sg13g2_a21oi_1 _09181_ (.A1(net117),
    .A2(_03551_),
    .Y(_03592_),
    .B1(_03575_));
 sg13g2_and3_1 _09182_ (.X(_03593_),
    .A(_03589_),
    .B(_03591_),
    .C(_03592_));
 sg13g2_nor2_1 _09183_ (.A(net117),
    .B(_03551_),
    .Y(_03594_));
 sg13g2_o21ai_1 _09184_ (.B1(net115),
    .Y(_03595_),
    .A1(_03562_),
    .A2(_03594_));
 sg13g2_nand2_1 _09185_ (.Y(_03596_),
    .A(_03562_),
    .B(_03594_));
 sg13g2_a21oi_1 _09186_ (.A1(_03595_),
    .A2(_03596_),
    .Y(_03597_),
    .B1(_03578_));
 sg13g2_nor3_1 _09187_ (.A(net121),
    .B(_03593_),
    .C(_03597_),
    .Y(_03598_));
 sg13g2_nand2b_1 _09188_ (.Y(_03599_),
    .B(_03551_),
    .A_N(_03562_));
 sg13g2_nor3_1 _09189_ (.A(_03589_),
    .B(_03591_),
    .C(_03599_),
    .Y(_03600_));
 sg13g2_nor4_1 _09190_ (.A(net116),
    .B(_03589_),
    .C(_03562_),
    .D(_03591_),
    .Y(_03601_));
 sg13g2_nand2_1 _09191_ (.Y(_03602_),
    .A(_03551_),
    .B(_03578_));
 sg13g2_nor3_1 _09192_ (.A(net115),
    .B(_03589_),
    .C(_03602_),
    .Y(_03603_));
 sg13g2_nor3_1 _09193_ (.A(_02766_),
    .B(_03589_),
    .C(_03591_),
    .Y(_03604_));
 sg13g2_or4_1 _09194_ (.A(_03600_),
    .B(_03601_),
    .C(_03603_),
    .D(_03604_),
    .X(_03605_));
 sg13g2_buf_1 _09195_ (.A(_03605_),
    .X(_03606_));
 sg13g2_nor3_1 _09196_ (.A(net116),
    .B(_03591_),
    .C(_03599_),
    .Y(_03607_));
 sg13g2_nor3_1 _09197_ (.A(net115),
    .B(_03562_),
    .C(_03591_),
    .Y(_03608_));
 sg13g2_nor2_1 _09198_ (.A(_03607_),
    .B(_03608_),
    .Y(_03609_));
 sg13g2_o21ai_1 _09199_ (.B1(_03609_),
    .Y(_03610_),
    .A1(_02766_),
    .A2(_03602_));
 sg13g2_nor3_1 _09200_ (.A(_03598_),
    .B(_03606_),
    .C(_03610_),
    .Y(_03611_));
 sg13g2_nand2_1 _09201_ (.Y(_03612_),
    .A(_03413_),
    .B(net367));
 sg13g2_mux2_1 _09202_ (.A0(_03546_),
    .A1(_03558_),
    .S(_03612_),
    .X(_03613_));
 sg13g2_xnor2_1 _09203_ (.Y(_03614_),
    .A(net179),
    .B(_03613_));
 sg13g2_xnor2_1 _09204_ (.Y(_03615_),
    .A(_03611_),
    .B(_03614_));
 sg13g2_mux2_1 _09205_ (.A0(_05382_),
    .A1(_05424_),
    .S(_05384_),
    .X(_03616_));
 sg13g2_nor2_1 _09206_ (.A(net262),
    .B(_03616_),
    .Y(_03617_));
 sg13g2_xnor2_1 _09207_ (.Y(_03618_),
    .A(_05392_),
    .B(_03617_));
 sg13g2_nor2_1 _09208_ (.A(net265),
    .B(_03618_),
    .Y(_03619_));
 sg13g2_a21oi_2 _09209_ (.B1(_03619_),
    .Y(_03620_),
    .A2(_03615_),
    .A1(net267));
 sg13g2_mux2_1 _09210_ (.A0(\dtop.vtop.pipeline.phases[0][12] ),
    .A1(_03620_),
    .S(net238),
    .X(_00253_));
 sg13g2_xor2_1 _09211_ (.B(_05285_),
    .A(_05279_),
    .X(_03621_));
 sg13g2_a21oi_1 _09212_ (.A1(_05382_),
    .A2(_05393_),
    .Y(_03622_),
    .B1(_05394_));
 sg13g2_nor2_1 _09213_ (.A(_05271_),
    .B(_03622_),
    .Y(_03623_));
 sg13g2_xnor2_1 _09214_ (.Y(_03624_),
    .A(_03621_),
    .B(_03623_));
 sg13g2_nor2_1 _09215_ (.A(net224),
    .B(_03613_),
    .Y(_03625_));
 sg13g2_nor4_1 _09216_ (.A(_03598_),
    .B(_03606_),
    .C(_03610_),
    .D(_03613_),
    .Y(_03626_));
 sg13g2_nor4_1 _09217_ (.A(net224),
    .B(_03598_),
    .C(_03606_),
    .D(_03610_),
    .Y(_03627_));
 sg13g2_nor3_2 _09218_ (.A(_03625_),
    .B(_03626_),
    .C(_03627_),
    .Y(_03628_));
 sg13g2_or2_1 _09219_ (.X(_03629_),
    .B(_03558_),
    .A(net221));
 sg13g2_buf_1 _09220_ (.A(_03629_),
    .X(_03630_));
 sg13g2_nand2_1 _09221_ (.Y(_03631_),
    .A(net221),
    .B(_03558_));
 sg13g2_nand2_1 _09222_ (.Y(_03632_),
    .A(_03630_),
    .B(_03631_));
 sg13g2_xnor2_1 _09223_ (.Y(_03633_),
    .A(_03628_),
    .B(_03632_));
 sg13g2_nor2_1 _09224_ (.A(net268),
    .B(_03633_),
    .Y(_03634_));
 sg13g2_a21oi_1 _09225_ (.A1(net252),
    .A2(_03624_),
    .Y(_03635_),
    .B1(_03634_));
 sg13g2_mux2_1 _09226_ (.A0(\dtop.vtop.pipeline.phases[0][13] ),
    .A1(_03635_),
    .S(net238),
    .X(_00254_));
 sg13g2_mux2_1 _09227_ (.A0(_03631_),
    .A1(_03630_),
    .S(_03628_),
    .X(_03636_));
 sg13g2_xor2_1 _09228_ (.B(_03636_),
    .A(_02387_),
    .X(_03637_));
 sg13g2_nor2_1 _09229_ (.A(net265),
    .B(_05415_),
    .Y(_03638_));
 sg13g2_a21oi_1 _09230_ (.A1(net267),
    .A2(_03637_),
    .Y(_03639_),
    .B1(_03638_));
 sg13g2_nor2_1 _09231_ (.A(\dtop.vtop.pipeline.phases[0][14] ),
    .B(net237),
    .Y(_03640_));
 sg13g2_a21oi_1 _09232_ (.A1(net238),
    .A2(_03639_),
    .Y(_00255_),
    .B1(_03640_));
 sg13g2_or2_1 _09233_ (.X(_03641_),
    .B(_03631_),
    .A(_02387_));
 sg13g2_nand2b_1 _09234_ (.Y(_03642_),
    .B(_02387_),
    .A_N(_03630_));
 sg13g2_mux2_1 _09235_ (.A0(_03641_),
    .A1(_03642_),
    .S(_03628_),
    .X(_03643_));
 sg13g2_xnor2_1 _09236_ (.Y(_03644_),
    .A(_03240_),
    .B(_03643_));
 sg13g2_nor2_1 _09237_ (.A(net265),
    .B(_05412_),
    .Y(_03645_));
 sg13g2_a21oi_1 _09238_ (.A1(net267),
    .A2(_03644_),
    .Y(_03646_),
    .B1(_03645_));
 sg13g2_nor2_1 _09239_ (.A(\dtop.vtop.pipeline.phases[0][15] ),
    .B(net237),
    .Y(_03647_));
 sg13g2_a21oi_1 _09240_ (.A1(net238),
    .A2(_03646_),
    .Y(_00256_),
    .B1(_03647_));
 sg13g2_nor2_1 _09241_ (.A(net367),
    .B(_03471_),
    .Y(_03648_));
 sg13g2_a21o_1 _09242_ (.A2(_03471_),
    .A1(_03428_),
    .B1(net367),
    .X(_03649_));
 sg13g2_a22oi_1 _09243_ (.Y(_03650_),
    .B1(_03649_),
    .B2(_03436_),
    .A2(_03490_),
    .A1(_03648_));
 sg13g2_nor2_1 _09244_ (.A(_03493_),
    .B(_03650_),
    .Y(_03651_));
 sg13g2_xor2_1 _09245_ (.B(_03651_),
    .A(_03487_),
    .X(_03652_));
 sg13g2_nor2_1 _09246_ (.A(_05210_),
    .B(net263),
    .Y(_03653_));
 sg13g2_nand3_1 _09247_ (.B(_05240_),
    .C(_03653_),
    .A(net268),
    .Y(_03654_));
 sg13g2_o21ai_1 _09248_ (.B1(_03654_),
    .Y(_03655_),
    .A1(_02862_),
    .A2(_03652_));
 sg13g2_mux2_1 _09249_ (.A0(\dtop.vtop.pipeline.phases[0][1] ),
    .A1(_03655_),
    .S(net237),
    .X(_00257_));
 sg13g2_a21oi_1 _09250_ (.A1(_03489_),
    .A2(_03492_),
    .Y(_03656_),
    .B1(_03493_));
 sg13g2_xnor2_1 _09251_ (.Y(_03657_),
    .A(_03478_),
    .B(_03483_));
 sg13g2_xnor2_1 _09252_ (.Y(_03658_),
    .A(_03656_),
    .B(_03657_));
 sg13g2_nand2_1 _09253_ (.Y(_03659_),
    .A(net265),
    .B(_03658_));
 sg13g2_and2_1 _09254_ (.A(_03654_),
    .B(_03659_),
    .X(_03660_));
 sg13g2_buf_1 _09255_ (.A(_03660_),
    .X(_03661_));
 sg13g2_nor2_1 _09256_ (.A(\dtop.vtop.pipeline.phases[0][2] ),
    .B(net237),
    .Y(_03662_));
 sg13g2_a21oi_1 _09257_ (.A1(net238),
    .A2(_03661_),
    .Y(_00258_),
    .B1(_03662_));
 sg13g2_nor2_1 _09258_ (.A(_03484_),
    .B(_03494_),
    .Y(_03663_));
 sg13g2_xnor2_1 _09259_ (.Y(_03664_),
    .A(_03498_),
    .B(_03507_));
 sg13g2_xnor2_1 _09260_ (.Y(_03665_),
    .A(_03663_),
    .B(_03664_));
 sg13g2_o21ai_1 _09261_ (.B1(_03653_),
    .Y(_03666_),
    .A1(net268),
    .A2(_03665_));
 sg13g2_nand2_1 _09262_ (.Y(_03667_),
    .A(\dtop.vtop.pipeline.phases[0][3] ),
    .B(_03417_));
 sg13g2_o21ai_1 _09263_ (.B1(_03667_),
    .Y(_00259_),
    .A1(_03417_),
    .A2(_03666_));
 sg13g2_xnor2_1 _09264_ (.Y(_03668_),
    .A(_03516_),
    .B(_03468_));
 sg13g2_xnor2_1 _09265_ (.Y(_03669_),
    .A(_03509_),
    .B(_03668_));
 sg13g2_nand2_1 _09266_ (.Y(_03670_),
    .A(net265),
    .B(_03669_));
 sg13g2_nand2_1 _09267_ (.Y(_03671_),
    .A(_05210_),
    .B(_05294_));
 sg13g2_nand3_1 _09268_ (.B(_03670_),
    .C(_03671_),
    .A(net261),
    .Y(_03672_));
 sg13g2_nand2_1 _09269_ (.Y(_03673_),
    .A(\dtop.vtop.pipeline.phases[0][4] ),
    .B(_03417_));
 sg13g2_o21ai_1 _09270_ (.B1(_03673_),
    .Y(_00260_),
    .A1(_03417_),
    .A2(_03672_));
 sg13g2_nor2_1 _09271_ (.A(_03468_),
    .B(_03509_),
    .Y(_03674_));
 sg13g2_nor2_1 _09272_ (.A(_03518_),
    .B(_03674_),
    .Y(_03675_));
 sg13g2_xnor2_1 _09273_ (.Y(_03676_),
    .A(_03524_),
    .B(_03529_));
 sg13g2_xnor2_1 _09274_ (.Y(_03677_),
    .A(_03675_),
    .B(_03676_));
 sg13g2_xnor2_1 _09275_ (.Y(_03678_),
    .A(_05313_),
    .B(_05299_));
 sg13g2_nor2_1 _09276_ (.A(net265),
    .B(_03678_),
    .Y(_03679_));
 sg13g2_a21oi_2 _09277_ (.B1(_03679_),
    .Y(_03680_),
    .A2(_03677_),
    .A1(_03418_));
 sg13g2_mux2_1 _09278_ (.A0(\dtop.vtop.pipeline.phases[0][5] ),
    .A1(_03680_),
    .S(net237),
    .X(_00261_));
 sg13g2_nor2_1 _09279_ (.A(_03524_),
    .B(_03675_),
    .Y(_03681_));
 sg13g2_nor2_1 _09280_ (.A(_03681_),
    .B(_03529_),
    .Y(_03682_));
 sg13g2_a21oi_1 _09281_ (.A1(_03524_),
    .A2(_03675_),
    .Y(_03683_),
    .B1(_03682_));
 sg13g2_xnor2_1 _09282_ (.Y(_03684_),
    .A(net126),
    .B(_03521_));
 sg13g2_xnor2_1 _09283_ (.Y(_03685_),
    .A(_03683_),
    .B(_03684_));
 sg13g2_xnor2_1 _09284_ (.Y(_03686_),
    .A(_05301_),
    .B(_05345_));
 sg13g2_a21oi_1 _09285_ (.A1(net260),
    .A2(_03686_),
    .Y(_03687_),
    .B1(_05311_));
 sg13g2_and3_1 _09286_ (.X(_03688_),
    .A(_05284_),
    .B(_05311_),
    .C(_03686_));
 sg13g2_o21ai_1 _09287_ (.B1(net268),
    .Y(_03689_),
    .A1(_03687_),
    .A2(_03688_));
 sg13g2_o21ai_1 _09288_ (.B1(_03689_),
    .Y(_03690_),
    .A1(_03408_),
    .A2(_03685_));
 sg13g2_nor2_1 _09289_ (.A(\dtop.vtop.pipeline.phases[0][6] ),
    .B(net237),
    .Y(_03691_));
 sg13g2_a21oi_1 _09290_ (.A1(net238),
    .A2(_03690_),
    .Y(_00262_),
    .B1(_03691_));
 sg13g2_xnor2_1 _09291_ (.Y(_03692_),
    .A(net145),
    .B(_03540_));
 sg13g2_xnor2_1 _09292_ (.Y(_03693_),
    .A(_03536_),
    .B(_03692_));
 sg13g2_nor2_1 _09293_ (.A(_05311_),
    .B(_05345_),
    .Y(_03694_));
 sg13g2_nor2_1 _09294_ (.A(_05347_),
    .B(_03694_),
    .Y(_03695_));
 sg13g2_xnor2_1 _09295_ (.Y(_03696_),
    .A(net421),
    .B(_03695_));
 sg13g2_nor2_1 _09296_ (.A(net262),
    .B(_03696_),
    .Y(_03697_));
 sg13g2_xnor2_1 _09297_ (.Y(_03698_),
    .A(_05320_),
    .B(_03697_));
 sg13g2_nor2_1 _09298_ (.A(net265),
    .B(_03698_),
    .Y(_03699_));
 sg13g2_a21oi_1 _09299_ (.A1(_03418_),
    .A2(_03693_),
    .Y(_03700_),
    .B1(_03699_));
 sg13g2_nor2_1 _09300_ (.A(\dtop.vtop.pipeline.phases[0][7] ),
    .B(_03572_),
    .Y(_03701_));
 sg13g2_a21oi_1 _09301_ (.A1(_03442_),
    .A2(_03700_),
    .Y(_00263_),
    .B1(_03701_));
 sg13g2_a21oi_1 _09302_ (.A1(_03536_),
    .A2(_03541_),
    .Y(_03702_),
    .B1(_03542_));
 sg13g2_xnor2_1 _09303_ (.Y(_03703_),
    .A(net151),
    .B(_03462_));
 sg13g2_xnor2_1 _09304_ (.Y(_03704_),
    .A(_03702_),
    .B(_03703_));
 sg13g2_a21oi_1 _09305_ (.A1(_05348_),
    .A2(_03695_),
    .Y(_03705_),
    .B1(net421));
 sg13g2_a21oi_1 _09306_ (.A1(_05312_),
    .A2(_05321_),
    .Y(_03706_),
    .B1(_03705_));
 sg13g2_xor2_1 _09307_ (.B(_03706_),
    .A(net423),
    .X(_03707_));
 sg13g2_nand2_1 _09308_ (.Y(_03708_),
    .A(net260),
    .B(_03707_));
 sg13g2_xnor2_1 _09309_ (.Y(_03709_),
    .A(_05339_),
    .B(_03708_));
 sg13g2_nor2_1 _09310_ (.A(net265),
    .B(_03709_),
    .Y(_03710_));
 sg13g2_a21oi_2 _09311_ (.B1(_03710_),
    .Y(_03711_),
    .A2(_03704_),
    .A1(_03565_));
 sg13g2_mux2_1 _09312_ (.A0(\dtop.vtop.pipeline.phases[0][8] ),
    .A1(_03711_),
    .S(net237),
    .X(_00264_));
 sg13g2_o21ai_1 _09313_ (.B1(_03706_),
    .Y(_03712_),
    .A1(net423),
    .A2(_05339_));
 sg13g2_nand2_1 _09314_ (.Y(_03713_),
    .A(_05356_),
    .B(_03712_));
 sg13g2_xnor2_1 _09315_ (.Y(_03714_),
    .A(_00756_),
    .B(_03713_));
 sg13g2_nand2_1 _09316_ (.Y(_03715_),
    .A(net260),
    .B(_03714_));
 sg13g2_xnor2_1 _09317_ (.Y(_03716_),
    .A(_05329_),
    .B(_03715_));
 sg13g2_xnor2_1 _09318_ (.Y(_03717_),
    .A(net116),
    .B(_03551_));
 sg13g2_xnor2_1 _09319_ (.Y(_03718_),
    .A(_03589_),
    .B(_03717_));
 sg13g2_nor2_1 _09320_ (.A(net268),
    .B(_03718_),
    .Y(_03719_));
 sg13g2_a21oi_2 _09321_ (.B1(_03719_),
    .Y(_03720_),
    .A2(_03716_),
    .A1(_03408_));
 sg13g2_nor2_1 _09322_ (.A(\dtop.vtop.pipeline.phases[0][9] ),
    .B(net237),
    .Y(_03721_));
 sg13g2_a21oi_1 _09323_ (.A1(_03442_),
    .A2(_03720_),
    .Y(_00265_),
    .B1(_03721_));
 sg13g2_inv_1 _09324_ (.Y(_03722_),
    .A(_03439_));
 sg13g2_nand3_1 _09325_ (.B(_02251_),
    .C(net278),
    .A(_02249_),
    .Y(_03723_));
 sg13g2_o21ai_1 _09326_ (.B1(_03723_),
    .Y(_03724_),
    .A1(net278),
    .A2(_01315_));
 sg13g2_buf_1 _09327_ (.A(_03724_),
    .X(_03725_));
 sg13g2_buf_1 _09328_ (.A(_03725_),
    .X(_03726_));
 sg13g2_mux2_1 _09329_ (.A0(\dtop.vtop.pipeline.phases[1][0] ),
    .A1(_03722_),
    .S(net214),
    .X(_00266_));
 sg13g2_buf_1 _09330_ (.A(_03725_),
    .X(_03727_));
 sg13g2_nor2_1 _09331_ (.A(\dtop.vtop.pipeline.phases[1][10] ),
    .B(net213),
    .Y(_03728_));
 sg13g2_a21oi_1 _09332_ (.A1(_03571_),
    .A2(net214),
    .Y(_00267_),
    .B1(_03728_));
 sg13g2_mux2_1 _09333_ (.A0(\dtop.vtop.pipeline.phases[1][11] ),
    .A1(_03587_),
    .S(_03726_),
    .X(_00268_));
 sg13g2_mux2_1 _09334_ (.A0(\dtop.vtop.pipeline.phases[1][12] ),
    .A1(_03620_),
    .S(net214),
    .X(_00269_));
 sg13g2_mux2_1 _09335_ (.A0(\dtop.vtop.pipeline.phases[1][13] ),
    .A1(_03635_),
    .S(net213),
    .X(_00270_));
 sg13g2_nor2_1 _09336_ (.A(\dtop.vtop.pipeline.phases[1][14] ),
    .B(net213),
    .Y(_03729_));
 sg13g2_a21oi_1 _09337_ (.A1(_03639_),
    .A2(net214),
    .Y(_00271_),
    .B1(_03729_));
 sg13g2_nor2_1 _09338_ (.A(\dtop.vtop.pipeline.phases[1][15] ),
    .B(net213),
    .Y(_03730_));
 sg13g2_a21oi_1 _09339_ (.A1(_03646_),
    .A2(net214),
    .Y(_00272_),
    .B1(_03730_));
 sg13g2_mux2_1 _09340_ (.A0(\dtop.vtop.pipeline.phases[1][1] ),
    .A1(_03655_),
    .S(net213),
    .X(_00273_));
 sg13g2_nor2_1 _09341_ (.A(\dtop.vtop.pipeline.phases[1][2] ),
    .B(_03727_),
    .Y(_03731_));
 sg13g2_a21oi_1 _09342_ (.A1(_03661_),
    .A2(_03726_),
    .Y(_00274_),
    .B1(_03731_));
 sg13g2_inv_1 _09343_ (.Y(_03732_),
    .A(_03666_));
 sg13g2_mux2_1 _09344_ (.A0(\dtop.vtop.pipeline.phases[1][3] ),
    .A1(_03732_),
    .S(net213),
    .X(_00275_));
 sg13g2_inv_1 _09345_ (.Y(_03733_),
    .A(_03672_));
 sg13g2_mux2_1 _09346_ (.A0(\dtop.vtop.pipeline.phases[1][4] ),
    .A1(_03733_),
    .S(net213),
    .X(_00276_));
 sg13g2_mux2_1 _09347_ (.A0(\dtop.vtop.pipeline.phases[1][5] ),
    .A1(_03680_),
    .S(_03727_),
    .X(_00277_));
 sg13g2_nor2_1 _09348_ (.A(\dtop.vtop.pipeline.phases[1][6] ),
    .B(_03725_),
    .Y(_03734_));
 sg13g2_a21oi_1 _09349_ (.A1(_03690_),
    .A2(net214),
    .Y(_00278_),
    .B1(_03734_));
 sg13g2_nor2_1 _09350_ (.A(\dtop.vtop.pipeline.phases[1][7] ),
    .B(_03725_),
    .Y(_03735_));
 sg13g2_a21oi_1 _09351_ (.A1(_03700_),
    .A2(net214),
    .Y(_00279_),
    .B1(_03735_));
 sg13g2_mux2_1 _09352_ (.A0(\dtop.vtop.pipeline.phases[1][8] ),
    .A1(_03711_),
    .S(net213),
    .X(_00280_));
 sg13g2_nor2_1 _09353_ (.A(\dtop.vtop.pipeline.phases[1][9] ),
    .B(_03725_),
    .Y(_03736_));
 sg13g2_a21oi_1 _09354_ (.A1(_03720_),
    .A2(net214),
    .Y(_00281_),
    .B1(_03736_));
 sg13g2_a22oi_1 _09355_ (.Y(_03737_),
    .B1(_02252_),
    .B2(_03328_),
    .A2(net268),
    .A1(_05163_));
 sg13g2_buf_1 _09356_ (.A(_03737_),
    .X(_03738_));
 sg13g2_nand2_1 _09357_ (.Y(_03739_),
    .A(\dtop.vtop.pipeline.phases[2][0] ),
    .B(_03738_));
 sg13g2_o21ai_1 _09358_ (.B1(_03739_),
    .Y(_00282_),
    .A1(_03439_),
    .A2(_03738_));
 sg13g2_nand2_1 _09359_ (.Y(_03740_),
    .A(_02252_),
    .B(_03328_));
 sg13g2_o21ai_1 _09360_ (.B1(_03740_),
    .Y(_03741_),
    .A1(_01453_),
    .A2(net278));
 sg13g2_buf_1 _09361_ (.A(_03741_),
    .X(_03742_));
 sg13g2_buf_1 _09362_ (.A(_03742_),
    .X(_03743_));
 sg13g2_buf_1 _09363_ (.A(_03742_),
    .X(_03744_));
 sg13g2_nor2_1 _09364_ (.A(\dtop.vtop.pipeline.phases[2][10] ),
    .B(net82),
    .Y(_03745_));
 sg13g2_a21oi_1 _09365_ (.A1(_03571_),
    .A2(net83),
    .Y(_00283_),
    .B1(_03745_));
 sg13g2_mux2_1 _09366_ (.A0(\dtop.vtop.pipeline.phases[2][11] ),
    .A1(_03587_),
    .S(net83),
    .X(_00284_));
 sg13g2_nand2_1 _09367_ (.Y(_03746_),
    .A(_03620_),
    .B(_03742_));
 sg13g2_o21ai_1 _09368_ (.B1(_03746_),
    .Y(_00285_),
    .A1(_02550_),
    .A2(net83));
 sg13g2_mux2_1 _09369_ (.A0(\dtop.vtop.pipeline.phases[2][13] ),
    .A1(_03635_),
    .S(net82),
    .X(_00286_));
 sg13g2_nor2_1 _09370_ (.A(\dtop.vtop.pipeline.phases[2][14] ),
    .B(net82),
    .Y(_03747_));
 sg13g2_a21oi_1 _09371_ (.A1(_03639_),
    .A2(net83),
    .Y(_00287_),
    .B1(_03747_));
 sg13g2_nor2_1 _09372_ (.A(\dtop.vtop.pipeline.phases[2][15] ),
    .B(net82),
    .Y(_03748_));
 sg13g2_a21oi_1 _09373_ (.A1(_03646_),
    .A2(net83),
    .Y(_00288_),
    .B1(_03748_));
 sg13g2_mux2_1 _09374_ (.A0(\dtop.vtop.pipeline.phases[2][1] ),
    .A1(_03655_),
    .S(net82),
    .X(_00289_));
 sg13g2_nor2_1 _09375_ (.A(\dtop.vtop.pipeline.phases[2][2] ),
    .B(net82),
    .Y(_03749_));
 sg13g2_a21oi_1 _09376_ (.A1(_03661_),
    .A2(net83),
    .Y(_00290_),
    .B1(_03749_));
 sg13g2_nand2_1 _09377_ (.Y(_03750_),
    .A(\dtop.vtop.pipeline.phases[2][3] ),
    .B(_03738_));
 sg13g2_o21ai_1 _09378_ (.B1(_03750_),
    .Y(_00291_),
    .A1(_03666_),
    .A2(_03738_));
 sg13g2_nand2_1 _09379_ (.Y(_03751_),
    .A(\dtop.vtop.pipeline.phases[2][4] ),
    .B(_03738_));
 sg13g2_o21ai_1 _09380_ (.B1(_03751_),
    .Y(_00292_),
    .A1(_03672_),
    .A2(_03738_));
 sg13g2_mux2_1 _09381_ (.A0(\dtop.vtop.pipeline.phases[2][5] ),
    .A1(_03680_),
    .S(net82),
    .X(_00293_));
 sg13g2_nor2_1 _09382_ (.A(\dtop.vtop.pipeline.phases[2][6] ),
    .B(net82),
    .Y(_03752_));
 sg13g2_a21oi_1 _09383_ (.A1(_03690_),
    .A2(net83),
    .Y(_00294_),
    .B1(_03752_));
 sg13g2_nor2_1 _09384_ (.A(\dtop.vtop.pipeline.phases[2][7] ),
    .B(_03744_),
    .Y(_03753_));
 sg13g2_a21oi_1 _09385_ (.A1(_03700_),
    .A2(_03743_),
    .Y(_00295_),
    .B1(_03753_));
 sg13g2_nand2_1 _09386_ (.Y(_03754_),
    .A(_03711_),
    .B(_03742_));
 sg13g2_o21ai_1 _09387_ (.B1(_03754_),
    .Y(_00296_),
    .A1(_02333_),
    .A2(net83));
 sg13g2_nor2_1 _09388_ (.A(\dtop.vtop.pipeline.phases[2][9] ),
    .B(_03744_),
    .Y(_03755_));
 sg13g2_a21oi_1 _09389_ (.A1(_03720_),
    .A2(_03743_),
    .Y(_00297_),
    .B1(_03755_));
 sg13g2_o21ai_1 _09390_ (.B1(_03351_),
    .Y(_03756_),
    .A1(net271),
    .A2(net269));
 sg13g2_buf_1 _09391_ (.A(_03756_),
    .X(_03757_));
 sg13g2_nor2_1 _09392_ (.A(_02357_),
    .B(_03757_),
    .Y(_03758_));
 sg13g2_buf_2 _09393_ (.A(_03758_),
    .X(_03759_));
 sg13g2_xnor2_1 _09394_ (.Y(_03760_),
    .A(_03050_),
    .B(_03759_));
 sg13g2_nand2_1 _09395_ (.Y(_03761_),
    .A(\dtop.vtop.pipeline.zg[0] ),
    .B(net96));
 sg13g2_o21ai_1 _09396_ (.B1(_03761_),
    .Y(_00315_),
    .A1(net96),
    .A2(_03760_));
 sg13g2_buf_1 _09397_ (.A(_03757_),
    .X(_03762_));
 sg13g2_nand2_1 _09398_ (.Y(_03763_),
    .A(_02356_),
    .B(_03050_));
 sg13g2_xnor2_1 _09399_ (.Y(_03764_),
    .A(_02342_),
    .B(_03763_));
 sg13g2_nor2_1 _09400_ (.A(net212),
    .B(_03764_),
    .Y(_03765_));
 sg13g2_xnor2_1 _09401_ (.Y(_03766_),
    .A(_03123_),
    .B(_03765_));
 sg13g2_mux2_1 _09402_ (.A0(\dtop.vtop.pipeline.zg[1] ),
    .A1(_03766_),
    .S(net84),
    .X(_00316_));
 sg13g2_nor2_1 _09403_ (.A(net271),
    .B(net269),
    .Y(_03767_));
 sg13g2_nor2_1 _09404_ (.A(_03347_),
    .B(_03767_),
    .Y(_03768_));
 sg13g2_buf_1 _09405_ (.A(_03768_),
    .X(_03769_));
 sg13g2_a21o_1 _09406_ (.A2(_03763_),
    .A1(_03123_),
    .B1(_02342_),
    .X(_03770_));
 sg13g2_o21ai_1 _09407_ (.B1(_03770_),
    .Y(_03771_),
    .A1(_03123_),
    .A2(_03763_));
 sg13g2_xnor2_1 _09408_ (.Y(_03772_),
    .A(_02299_),
    .B(_03771_));
 sg13g2_nand2_1 _09409_ (.Y(_03773_),
    .A(_03769_),
    .B(_03772_));
 sg13g2_xnor2_1 _09410_ (.Y(_03774_),
    .A(_03162_),
    .B(_03773_));
 sg13g2_nand2_1 _09411_ (.Y(_03775_),
    .A(net95),
    .B(_03774_));
 sg13g2_o21ai_1 _09412_ (.B1(_03775_),
    .Y(_00317_),
    .A1(_03286_),
    .A2(net84));
 sg13g2_nand2_1 _09413_ (.Y(_03776_),
    .A(_02298_),
    .B(_03162_));
 sg13g2_nand2_1 _09414_ (.Y(_03777_),
    .A(net248),
    .B(net220));
 sg13g2_a22oi_1 _09415_ (.Y(_03778_),
    .B1(_03102_),
    .B2(_03108_),
    .A2(_03097_),
    .A1(_02900_));
 sg13g2_o21ai_1 _09416_ (.B1(_03778_),
    .Y(_03779_),
    .A1(_03078_),
    .A2(_03093_));
 sg13g2_nor2_1 _09417_ (.A(_02254_),
    .B(net220),
    .Y(_03780_));
 sg13g2_inv_1 _09418_ (.Y(_03781_),
    .A(_03038_));
 sg13g2_and4_1 _09419_ (.A(net219),
    .B(net220),
    .C(_03021_),
    .D(_03781_),
    .X(_03782_));
 sg13g2_a221oi_1 _09420_ (.B2(_03780_),
    .C1(_03782_),
    .B1(_03779_),
    .A1(_02968_),
    .Y(_03783_),
    .A2(_03044_));
 sg13g2_o21ai_1 _09421_ (.B1(_03783_),
    .Y(_03784_),
    .A1(_02715_),
    .A2(_03777_));
 sg13g2_nand2_2 _09422_ (.Y(_03785_),
    .A(_02356_),
    .B(_03768_));
 sg13g2_nor4_1 _09423_ (.A(net166),
    .B(_03048_),
    .C(_03784_),
    .D(_03785_),
    .Y(_03786_));
 sg13g2_and4_1 _09424_ (.A(net166),
    .B(_03048_),
    .C(_03784_),
    .D(_03759_),
    .X(_03787_));
 sg13g2_nor3_1 _09425_ (.A(_02342_),
    .B(_02286_),
    .C(_03785_),
    .Y(_03788_));
 sg13g2_nor3_1 _09426_ (.A(_02342_),
    .B(net176),
    .C(_03785_),
    .Y(_03789_));
 sg13g2_mux2_1 _09427_ (.A0(_03788_),
    .A1(_03789_),
    .S(_03048_),
    .X(_03790_));
 sg13g2_nor3_1 _09428_ (.A(_02342_),
    .B(_03113_),
    .C(_03121_),
    .Y(_03791_));
 sg13g2_nor4_1 _09429_ (.A(_03786_),
    .B(_03787_),
    .C(_03790_),
    .D(_03791_),
    .Y(_03792_));
 sg13g2_nor2_1 _09430_ (.A(_02298_),
    .B(_03162_),
    .Y(_03793_));
 sg13g2_a21oi_1 _09431_ (.A1(_03776_),
    .A2(_03792_),
    .Y(_03794_),
    .B1(_03793_));
 sg13g2_xnor2_1 _09432_ (.Y(_03795_),
    .A(_02399_),
    .B(_03794_));
 sg13g2_nor2_1 _09433_ (.A(net212),
    .B(_03795_),
    .Y(_03796_));
 sg13g2_xnor2_1 _09434_ (.Y(_03797_),
    .A(_03248_),
    .B(_03796_));
 sg13g2_nand2_1 _09435_ (.Y(_03798_),
    .A(_03283_),
    .B(net112));
 sg13g2_o21ai_1 _09436_ (.B1(_03798_),
    .Y(_00318_),
    .A1(net96),
    .A2(_03797_));
 sg13g2_nor2_1 _09437_ (.A(_03248_),
    .B(_03794_),
    .Y(_03799_));
 sg13g2_nand2_1 _09438_ (.Y(_03800_),
    .A(_03248_),
    .B(_03794_));
 sg13g2_o21ai_1 _09439_ (.B1(_03800_),
    .Y(_03801_),
    .A1(_02400_),
    .A2(_03799_));
 sg13g2_xnor2_1 _09440_ (.Y(_03802_),
    .A(_02455_),
    .B(_03801_));
 sg13g2_nor2_1 _09441_ (.A(net212),
    .B(_03802_),
    .Y(_03803_));
 sg13g2_xor2_1 _09442_ (.B(_03803_),
    .A(_03221_),
    .X(_03804_));
 sg13g2_mux2_1 _09443_ (.A0(net408),
    .A1(_03804_),
    .S(net84),
    .X(_00319_));
 sg13g2_a21o_1 _09444_ (.A2(_03792_),
    .A1(_03776_),
    .B1(_03793_),
    .X(_03805_));
 sg13g2_nand2_1 _09445_ (.Y(_03806_),
    .A(_03248_),
    .B(_03221_));
 sg13g2_a21oi_1 _09446_ (.A1(_02342_),
    .A2(_02299_),
    .Y(_03807_),
    .B1(_03757_));
 sg13g2_nand3_1 _09447_ (.B(_03759_),
    .C(_03807_),
    .A(net176),
    .Y(_03808_));
 sg13g2_or2_1 _09448_ (.X(_03809_),
    .B(_03808_),
    .A(_03048_));
 sg13g2_nand4_1 _09449_ (.B(_03048_),
    .C(_03759_),
    .A(net166),
    .Y(_03810_),
    .D(_03807_));
 sg13g2_nand2_1 _09450_ (.Y(_03811_),
    .A(_02298_),
    .B(_03768_));
 sg13g2_nand4_1 _09451_ (.B(_03809_),
    .C(_03810_),
    .A(_03123_),
    .Y(_03812_),
    .D(_03811_));
 sg13g2_nand3_1 _09452_ (.B(net166),
    .C(_03759_),
    .A(net248),
    .Y(_03813_));
 sg13g2_nand3_1 _09453_ (.B(net176),
    .C(_03759_),
    .A(net248),
    .Y(_03814_));
 sg13g2_mux2_1 _09454_ (.A0(_03813_),
    .A1(_03814_),
    .S(_02857_),
    .X(_03815_));
 sg13g2_nor4_1 _09455_ (.A(net248),
    .B(net176),
    .C(_03042_),
    .D(_03785_),
    .Y(_03816_));
 sg13g2_and4_1 _09456_ (.A(net177),
    .B(net176),
    .C(_03042_),
    .D(_03759_),
    .X(_03817_));
 sg13g2_nor3_1 _09457_ (.A(_03807_),
    .B(_03816_),
    .C(_03817_),
    .Y(_03818_));
 sg13g2_a21o_1 _09458_ (.A2(_03219_),
    .A1(_03199_),
    .B1(_02455_),
    .X(_03819_));
 sg13g2_a22oi_1 _09459_ (.Y(_03820_),
    .B1(_03819_),
    .B2(_02399_),
    .A2(_03248_),
    .A1(_02455_));
 sg13g2_nand2b_1 _09460_ (.Y(_03821_),
    .B(_03162_),
    .A_N(_03820_));
 sg13g2_a21oi_1 _09461_ (.A1(_03815_),
    .A2(_03818_),
    .Y(_03822_),
    .B1(_03821_));
 sg13g2_nor2_1 _09462_ (.A(_03811_),
    .B(_03820_),
    .Y(_03823_));
 sg13g2_or4_1 _09463_ (.A(_03786_),
    .B(_03787_),
    .C(_03790_),
    .D(_03791_),
    .X(_03824_));
 sg13g2_nor2_1 _09464_ (.A(_02400_),
    .B(_03194_),
    .Y(_03825_));
 sg13g2_and2_1 _09465_ (.A(_02455_),
    .B(_03221_),
    .X(_03826_));
 sg13g2_a21o_1 _09466_ (.A2(_03825_),
    .A1(_03819_),
    .B1(_03826_),
    .X(_03827_));
 sg13g2_a221oi_1 _09467_ (.B2(_03824_),
    .C1(_03827_),
    .B1(_03823_),
    .A1(_03812_),
    .Y(_03828_),
    .A2(_03822_));
 sg13g2_o21ai_1 _09468_ (.B1(_03828_),
    .Y(_03829_),
    .A1(_03805_),
    .A2(_03806_));
 sg13g2_buf_1 _09469_ (.A(_03829_),
    .X(_03830_));
 sg13g2_nand2_1 _09470_ (.Y(_03831_),
    .A(net211),
    .B(_03830_));
 sg13g2_xnor2_1 _09471_ (.Y(_03832_),
    .A(net33),
    .B(_03831_));
 sg13g2_nand2_1 _09472_ (.Y(_03833_),
    .A(_02553_),
    .B(net211));
 sg13g2_inv_1 _09473_ (.Y(_03834_),
    .A(_03833_));
 sg13g2_xnor2_1 _09474_ (.Y(_03835_),
    .A(_03832_),
    .B(_03834_));
 sg13g2_nand2_1 _09475_ (.Y(_03836_),
    .A(_03274_),
    .B(net112));
 sg13g2_o21ai_1 _09476_ (.B1(_03836_),
    .Y(_00320_),
    .A1(net96),
    .A2(_03835_));
 sg13g2_o21ai_1 _09477_ (.B1(_03834_),
    .Y(_03837_),
    .A1(net33),
    .A2(_03830_));
 sg13g2_nand3_1 _09478_ (.B(net211),
    .C(_03830_),
    .A(net33),
    .Y(_03838_));
 sg13g2_nand2_1 _09479_ (.Y(_03839_),
    .A(_03837_),
    .B(_03838_));
 sg13g2_nor2_1 _09480_ (.A(_02620_),
    .B(net212),
    .Y(_03840_));
 sg13g2_xnor2_1 _09481_ (.Y(_03841_),
    .A(_03233_),
    .B(_03840_));
 sg13g2_xnor2_1 _09482_ (.Y(_03842_),
    .A(_03839_),
    .B(_03841_));
 sg13g2_mux2_1 _09483_ (.A0(_03277_),
    .A1(_03842_),
    .S(net84),
    .X(_00321_));
 sg13g2_nand2b_1 _09484_ (.Y(_03843_),
    .B(net95),
    .A_N(net410));
 sg13g2_nand3_1 _09485_ (.B(_03363_),
    .C(net211),
    .A(net410),
    .Y(_03844_));
 sg13g2_nand2_1 _09486_ (.Y(_03845_),
    .A(net410),
    .B(net95));
 sg13g2_nor2_1 _09487_ (.A(net410),
    .B(_03757_),
    .Y(_03846_));
 sg13g2_nand2_1 _09488_ (.Y(_03847_),
    .A(net95),
    .B(_03846_));
 sg13g2_nor2_1 _09489_ (.A(net33),
    .B(_03830_),
    .Y(_03848_));
 sg13g2_a21oi_1 _09490_ (.A1(net33),
    .A2(_03830_),
    .Y(_03849_),
    .B1(_02553_));
 sg13g2_nor3_1 _09491_ (.A(_03234_),
    .B(_03848_),
    .C(_03849_),
    .Y(_03850_));
 sg13g2_o21ai_1 _09492_ (.B1(_03234_),
    .Y(_03851_),
    .A1(_03848_),
    .A2(_03849_));
 sg13g2_o21ai_1 _09493_ (.B1(_03851_),
    .Y(_03852_),
    .A1(_02686_),
    .A2(_03850_));
 sg13g2_mux4_1 _09494_ (.S0(_03251_),
    .A0(_03843_),
    .A1(_03844_),
    .A2(_03845_),
    .A3(_03847_),
    .S1(_03852_),
    .X(_03853_));
 sg13g2_nor3_1 _09495_ (.A(_03251_),
    .B(net112),
    .C(net211),
    .Y(_03854_));
 sg13g2_a21oi_1 _09496_ (.A1(_03309_),
    .A2(net112),
    .Y(_03855_),
    .B1(_03854_));
 sg13g2_nand2_1 _09497_ (.Y(_00322_),
    .A(_03853_),
    .B(_03855_));
 sg13g2_nand2_1 _09498_ (.Y(_03856_),
    .A(_03233_),
    .B(_03846_));
 sg13g2_a21oi_1 _09499_ (.A1(net410),
    .A2(_03251_),
    .Y(_03857_),
    .B1(_02620_));
 sg13g2_nand2_1 _09500_ (.Y(_03858_),
    .A(net211),
    .B(_03857_));
 sg13g2_a22oi_1 _09501_ (.Y(_03859_),
    .B1(_03856_),
    .B2(_03858_),
    .A2(_03838_),
    .A1(_03837_));
 sg13g2_or2_1 _09502_ (.X(_03860_),
    .B(_03251_),
    .A(_03234_));
 sg13g2_a21oi_1 _09503_ (.A1(_03837_),
    .A2(_03838_),
    .Y(_03861_),
    .B1(_03860_));
 sg13g2_nor2b_1 _09504_ (.A(_03251_),
    .B_N(_03846_),
    .Y(_03862_));
 sg13g2_nor2_1 _09505_ (.A(_03234_),
    .B(_03858_),
    .Y(_03863_));
 sg13g2_nor4_2 _09506_ (.A(_03859_),
    .B(_03861_),
    .C(_03862_),
    .Y(_03864_),
    .D(_03863_));
 sg13g2_buf_8 _09507_ (.A(_03864_),
    .X(_03865_));
 sg13g2_nor2_1 _09508_ (.A(_00079_),
    .B(_03767_),
    .Y(_03866_));
 sg13g2_nand3_1 _09509_ (.B(_03273_),
    .C(_03767_),
    .A(_02250_),
    .Y(_03867_));
 sg13g2_nand2b_1 _09510_ (.Y(_03868_),
    .B(_03867_),
    .A_N(_03866_));
 sg13g2_a22oi_1 _09511_ (.Y(_03869_),
    .B1(_03868_),
    .B2(_02249_),
    .A2(_03866_),
    .A1(_02250_));
 sg13g2_buf_1 _09512_ (.A(_03869_),
    .X(_03870_));
 sg13g2_xnor2_1 _09513_ (.Y(_03871_),
    .A(net217),
    .B(net141));
 sg13g2_xnor2_1 _09514_ (.Y(_03872_),
    .A(_03865_),
    .B(_03871_));
 sg13g2_mux2_1 _09515_ (.A0(_03311_),
    .A1(_03872_),
    .S(net84),
    .X(_00323_));
 sg13g2_or2_1 _09516_ (.X(_03873_),
    .B(net212),
    .A(\dtop.vtop.pipeline.zg_acc[9] ));
 sg13g2_buf_1 _09517_ (.A(_03873_),
    .X(_03874_));
 sg13g2_nand3_1 _09518_ (.B(net95),
    .C(_03874_),
    .A(net217),
    .Y(_03875_));
 sg13g2_nand3_1 _09519_ (.B(net95),
    .C(_03874_),
    .A(net247),
    .Y(_03876_));
 sg13g2_mux2_1 _09520_ (.A0(_03875_),
    .A1(_03876_),
    .S(_03865_),
    .X(_03877_));
 sg13g2_nor4_1 _09521_ (.A(net217),
    .B(_03329_),
    .C(net141),
    .D(_03874_),
    .Y(_03878_));
 sg13g2_nand2b_1 _09522_ (.Y(_03879_),
    .B(_03878_),
    .A_N(_03865_));
 sg13g2_nor2_1 _09523_ (.A(net247),
    .B(_03874_),
    .Y(_03880_));
 sg13g2_nand4_1 _09524_ (.B(_03865_),
    .C(net141),
    .A(_03364_),
    .Y(_03881_),
    .D(_03880_));
 sg13g2_buf_1 _09525_ (.A(_03305_),
    .X(_03882_));
 sg13g2_nand3b_1 _09526_ (.B(_03874_),
    .C(net217),
    .Y(_03883_),
    .A_N(net141));
 sg13g2_nand3_1 _09527_ (.B(net141),
    .C(_03874_),
    .A(net247),
    .Y(_03884_));
 sg13g2_a21oi_1 _09528_ (.A1(_03883_),
    .A2(_03884_),
    .Y(_03885_),
    .B1(_03330_));
 sg13g2_a21oi_1 _09529_ (.A1(net363),
    .A2(net112),
    .Y(_03886_),
    .B1(_03885_));
 sg13g2_nand4_1 _09530_ (.B(_03879_),
    .C(_03881_),
    .A(_03877_),
    .Y(_00324_),
    .D(_03886_));
 sg13g2_buf_2 _09531_ (.A(\dtop.vtop.rs.scan_y.phase[0] ),
    .X(_03887_));
 sg13g2_buf_1 _09532_ (.A(\dtop.vtop.rs.scan_y.phase[1] ),
    .X(_03888_));
 sg13g2_nor2b_1 _09533_ (.A(_03887_),
    .B_N(_03888_),
    .Y(_03889_));
 sg13g2_buf_1 _09534_ (.A(_00084_),
    .X(_03890_));
 sg13g2_buf_1 _09535_ (.A(\dtop.vtop.rs.x_scan.phase[1] ),
    .X(_03891_));
 sg13g2_nor4_1 _09536_ (.A(net377),
    .B(_03890_),
    .C(_03891_),
    .D(_05261_),
    .Y(_03892_));
 sg13g2_nand3_1 _09537_ (.B(net382),
    .C(_03892_),
    .A(net378),
    .Y(_03893_));
 sg13g2_inv_1 _09538_ (.Y(_03894_),
    .A(_03891_));
 sg13g2_nor4_1 _09539_ (.A(_00516_),
    .B(net382),
    .C(_03894_),
    .D(_05242_),
    .Y(_03895_));
 sg13g2_o21ai_1 _09540_ (.B1(_03895_),
    .Y(_03896_),
    .A1(net377),
    .A2(_03890_));
 sg13g2_buf_2 _09541_ (.A(\dtop.vtop.rs.x_scan.phase[0] ),
    .X(_03897_));
 sg13g2_nand2_1 _09542_ (.Y(_03898_),
    .A(net297),
    .B(_03897_));
 sg13g2_nor2_1 _09543_ (.A(_03890_),
    .B(_03898_),
    .Y(_03899_));
 sg13g2_nor3_1 _09544_ (.A(net297),
    .B(net377),
    .C(_03897_),
    .Y(_03900_));
 sg13g2_xnor2_1 _09545_ (.Y(_03901_),
    .A(_03890_),
    .B(_05188_));
 sg13g2_nor4_1 _09546_ (.A(net345),
    .B(_00411_),
    .C(net308),
    .D(_03901_),
    .Y(_03902_));
 sg13g2_o21ai_1 _09547_ (.B1(_03902_),
    .Y(_03903_),
    .A1(_03899_),
    .A2(_03900_));
 sg13g2_a21oi_2 _09548_ (.B1(_03903_),
    .Y(_03904_),
    .A2(_03896_),
    .A1(_03893_));
 sg13g2_nor2_1 _09549_ (.A(_03894_),
    .B(_03897_),
    .Y(_03905_));
 sg13g2_a21oi_1 _09550_ (.A1(_03904_),
    .A2(_03905_),
    .Y(_03906_),
    .B1(_00085_));
 sg13g2_mux2_1 _09551_ (.A0(_03889_),
    .A1(\dtop.vsync ),
    .S(_03906_),
    .X(_00350_));
 sg13g2_buf_1 _09552_ (.A(net419),
    .X(_03907_));
 sg13g2_buf_1 _09553_ (.A(net362),
    .X(_03908_));
 sg13g2_inv_1 _09554_ (.Y(_03909_),
    .A(net15));
 sg13g2_buf_1 _09555_ (.A(\dtop.ext_control[5] ),
    .X(_03910_));
 sg13g2_nand2_1 _09556_ (.Y(_03911_),
    .A(net419),
    .B(_03910_));
 sg13g2_o21ai_1 _09557_ (.B1(_03911_),
    .Y(_00376_),
    .A1(net337),
    .A2(_03909_));
 sg13g2_nor3_1 _09558_ (.A(net365),
    .B(net367),
    .C(_02850_),
    .Y(_03912_));
 sg13g2_nor2b_1 _09559_ (.A(_03912_),
    .B_N(\dtop.vtop.force_sat0 ),
    .Y(_03913_));
 sg13g2_nor2_1 _09560_ (.A(_01600_),
    .B(_03913_),
    .Y(_03914_));
 sg13g2_nor3_1 _09561_ (.A(net395),
    .B(_00520_),
    .C(_00523_),
    .Y(_03915_));
 sg13g2_nor3_1 _09562_ (.A(_00944_),
    .B(_00515_),
    .C(_03915_),
    .Y(_03916_));
 sg13g2_and2_1 _09563_ (.A(_00443_),
    .B(_00524_),
    .X(_03917_));
 sg13g2_or4_1 _09564_ (.A(_03891_),
    .B(_03897_),
    .C(_03916_),
    .D(_03917_),
    .X(_03918_));
 sg13g2_buf_1 _09565_ (.A(\dtop.vtop.pipeline.dz[7] ),
    .X(_03919_));
 sg13g2_inv_1 _09566_ (.Y(_03920_),
    .A(_03919_));
 sg13g2_xnor2_1 _09567_ (.Y(_03921_),
    .A(\dtop.vtop.pipeline.dz[6] ),
    .B(_00538_));
 sg13g2_xnor2_1 _09568_ (.Y(_03922_),
    .A(_00417_),
    .B(_00422_));
 sg13g2_buf_1 _09569_ (.A(\dtop.vtop.pipeline.dz[4] ),
    .X(_03923_));
 sg13g2_inv_1 _09570_ (.Y(_03924_),
    .A(\dtop.vtop.pipeline.dz[3] ));
 sg13g2_buf_2 _09571_ (.A(_00095_),
    .X(_03925_));
 sg13g2_buf_1 _09572_ (.A(\dtop.vtop.pipeline.dz[2] ),
    .X(_03926_));
 sg13g2_buf_2 _09573_ (.A(\dtop.vtop.pipeline.dz[0] ),
    .X(_03927_));
 sg13g2_buf_1 _09574_ (.A(\dtop.vtop.pipeline.dz[1] ),
    .X(_03928_));
 sg13g2_o21ai_1 _09575_ (.B1(_03928_),
    .Y(_03929_),
    .A1(net299),
    .A2(_03927_));
 sg13g2_nor3_1 _09576_ (.A(net299),
    .B(_03928_),
    .C(_03927_),
    .Y(_03930_));
 sg13g2_a21oi_1 _09577_ (.A1(net354),
    .A2(_03929_),
    .Y(_03931_),
    .B1(_03930_));
 sg13g2_nand2b_1 _09578_ (.Y(_03932_),
    .B(_03931_),
    .A_N(_03926_));
 sg13g2_a21o_1 _09579_ (.A2(_03932_),
    .A1(_03925_),
    .B1(_00445_),
    .X(_03933_));
 sg13g2_nand3_1 _09580_ (.B(_00445_),
    .C(_03931_),
    .A(_03926_),
    .Y(_03934_));
 sg13g2_a22oi_1 _09581_ (.Y(_03935_),
    .B1(_03933_),
    .B2(_03934_),
    .A2(_05228_),
    .A1(_03924_));
 sg13g2_a21oi_1 _09582_ (.A1(\dtop.vtop.pipeline.dz[3] ),
    .A2(_05193_),
    .Y(_03936_),
    .B1(_03935_));
 sg13g2_buf_2 _09583_ (.A(_00094_),
    .X(_03937_));
 sg13g2_o21ai_1 _09584_ (.B1(_03937_),
    .Y(_03938_),
    .A1(_03923_),
    .A2(_03936_));
 sg13g2_inv_1 _09585_ (.Y(_03939_),
    .A(_03923_));
 sg13g2_o21ai_1 _09586_ (.B1(_03922_),
    .Y(_03940_),
    .A1(_03939_),
    .A2(_03936_));
 sg13g2_o21ai_1 _09587_ (.B1(_03940_),
    .Y(_03941_),
    .A1(_03922_),
    .A2(_03938_));
 sg13g2_nand2_1 _09588_ (.Y(_03942_),
    .A(net231),
    .B(_03941_));
 sg13g2_nor2_1 _09589_ (.A(net231),
    .B(_03941_),
    .Y(_03943_));
 sg13g2_a21oi_1 _09590_ (.A1(\dtop.vtop.pipeline.dz[5] ),
    .A2(_03942_),
    .Y(_03944_),
    .B1(_03943_));
 sg13g2_buf_1 _09591_ (.A(_00093_),
    .X(_03945_));
 sg13g2_inv_1 _09592_ (.Y(_03946_),
    .A(_03945_));
 sg13g2_nand2_1 _09593_ (.Y(_03947_),
    .A(_03946_),
    .B(_00538_));
 sg13g2_o21ai_1 _09594_ (.B1(_03947_),
    .Y(_03948_),
    .A1(_03921_),
    .A2(_03944_));
 sg13g2_buf_2 _09595_ (.A(_00092_),
    .X(_03949_));
 sg13g2_inv_1 _09596_ (.Y(_03950_),
    .A(_03949_));
 sg13g2_a21oi_1 _09597_ (.A1(_03920_),
    .A2(_03948_),
    .Y(_03951_),
    .B1(_03950_));
 sg13g2_nand3_1 _09598_ (.B(net137),
    .C(_03948_),
    .A(_03919_),
    .Y(_03952_));
 sg13g2_o21ai_1 _09599_ (.B1(_03952_),
    .Y(_03953_),
    .A1(net110),
    .A2(_03951_));
 sg13g2_buf_1 _09600_ (.A(_00091_),
    .X(_03954_));
 sg13g2_inv_1 _09601_ (.Y(_03955_),
    .A(_03954_));
 sg13g2_o21ai_1 _09602_ (.B1(_03955_),
    .Y(_03956_),
    .A1(_00947_),
    .A2(_03953_));
 sg13g2_nand2_1 _09603_ (.Y(_03957_),
    .A(_00947_),
    .B(_03953_));
 sg13g2_a21oi_1 _09604_ (.A1(_03956_),
    .A2(_03957_),
    .Y(_03958_),
    .B1(_03918_));
 sg13g2_xnor2_1 _09605_ (.Y(_03959_),
    .A(_03919_),
    .B(net93));
 sg13g2_xnor2_1 _09606_ (.Y(_03960_),
    .A(_03923_),
    .B(_00423_));
 sg13g2_xnor2_1 _09607_ (.Y(_03961_),
    .A(_03926_),
    .B(_00445_));
 sg13g2_xor2_1 _09608_ (.B(_03928_),
    .A(net286),
    .X(_03962_));
 sg13g2_xor2_1 _09609_ (.B(_03927_),
    .A(net287),
    .X(_03963_));
 sg13g2_xnor2_1 _09610_ (.Y(_03964_),
    .A(_03924_),
    .B(_05193_));
 sg13g2_nand4_1 _09611_ (.B(_03962_),
    .C(_03963_),
    .A(_03961_),
    .Y(_03965_),
    .D(_03964_));
 sg13g2_xnor2_1 _09612_ (.Y(_03966_),
    .A(\dtop.vtop.pipeline.dz[5] ),
    .B(net201));
 sg13g2_nor4_1 _09613_ (.A(_03921_),
    .B(_03960_),
    .C(_03965_),
    .D(_03966_),
    .Y(_03967_));
 sg13g2_xnor2_1 _09614_ (.Y(_03968_),
    .A(_03954_),
    .B(_00947_));
 sg13g2_nand3_1 _09615_ (.B(_03967_),
    .C(_03968_),
    .A(_03959_),
    .Y(_03969_));
 sg13g2_inv_1 _09616_ (.Y(_03970_),
    .A(_00089_));
 sg13g2_inv_1 _09617_ (.Y(_03971_),
    .A(\dtop.vtop.pipeline.neg_t[4] ));
 sg13g2_xor2_1 _09618_ (.B(_05130_),
    .A(net357),
    .X(_03972_));
 sg13g2_nor4_2 _09619_ (.A(net390),
    .B(net401),
    .C(net393),
    .Y(_03973_),
    .D(_03972_));
 sg13g2_buf_1 _09620_ (.A(_03973_),
    .X(_03974_));
 sg13g2_nand2_1 _09621_ (.Y(_03975_),
    .A(net424),
    .B(_03974_));
 sg13g2_inv_1 _09622_ (.Y(_03976_),
    .A(_00021_));
 sg13g2_inv_1 _09623_ (.Y(_03977_),
    .A(net279));
 sg13g2_buf_1 _09624_ (.A(_00016_),
    .X(_03978_));
 sg13g2_inv_1 _09625_ (.Y(_03979_),
    .A(_03978_));
 sg13g2_buf_1 _09626_ (.A(_00015_),
    .X(_03980_));
 sg13g2_buf_1 _09627_ (.A(_00087_),
    .X(_03981_));
 sg13g2_inv_1 _09628_ (.Y(_03982_),
    .A(_03981_));
 sg13g2_nand3_1 _09629_ (.B(_00467_),
    .C(\dtop.vtop.pipeline.neg_t[0] ),
    .A(_03982_),
    .Y(_03983_));
 sg13g2_and4_1 _09630_ (.A(net425),
    .B(net404),
    .C(_03973_),
    .D(_03983_),
    .X(_03984_));
 sg13g2_nand2b_1 _09631_ (.Y(_03985_),
    .B(_03983_),
    .A_N(net404));
 sg13g2_a21oi_1 _09632_ (.A1(\dtop.vtop.pipeline.neg_t[1] ),
    .A2(_03985_),
    .Y(_03986_),
    .B1(net425));
 sg13g2_a21oi_1 _09633_ (.A1(net404),
    .A2(\dtop.vtop.pipeline.neg_t[1] ),
    .Y(_03987_),
    .B1(_03973_));
 sg13g2_nor3_1 _09634_ (.A(_03984_),
    .B(_03986_),
    .C(_03987_),
    .Y(_03988_));
 sg13g2_buf_1 _09635_ (.A(_00018_),
    .X(_03989_));
 sg13g2_nand2b_1 _09636_ (.Y(_03990_),
    .B(_03989_),
    .A_N(_03988_));
 sg13g2_a22oi_1 _09637_ (.Y(_03991_),
    .B1(_05303_),
    .B2(_03990_),
    .A2(_03979_),
    .A1(_05273_));
 sg13g2_inv_1 _09638_ (.Y(_03992_),
    .A(_03989_));
 sg13g2_nand2_1 _09639_ (.Y(_03993_),
    .A(_05273_),
    .B(_03973_));
 sg13g2_a22oi_1 _09640_ (.Y(_03994_),
    .B1(_03993_),
    .B2(_03978_),
    .A2(_03988_),
    .A1(_03992_));
 sg13g2_o21ai_1 _09641_ (.B1(_03994_),
    .Y(_03995_),
    .A1(_03977_),
    .A2(_03991_));
 sg13g2_a22oi_1 _09642_ (.Y(_03996_),
    .B1(_03995_),
    .B2(_05273_),
    .A2(_03976_),
    .A1(net424));
 sg13g2_nand2b_1 _09643_ (.Y(_03997_),
    .B(_03974_),
    .A_N(_03996_));
 sg13g2_a22oi_1 _09644_ (.Y(_03998_),
    .B1(_03995_),
    .B2(\dtop.vtop.pipeline.neg_t[3] ),
    .A2(_03975_),
    .A1(_00021_));
 sg13g2_a21oi_1 _09645_ (.A1(_05165_),
    .A2(net279),
    .Y(_03999_),
    .B1(\dtop.vtop.pipeline.neg_t[5] ));
 sg13g2_a221oi_1 _09646_ (.B2(_03998_),
    .C1(_03999_),
    .B1(_03997_),
    .A1(_03971_),
    .Y(_04000_),
    .A2(_03975_));
 sg13g2_buf_1 _09647_ (.A(_00025_),
    .X(_04001_));
 sg13g2_buf_2 _09648_ (.A(_00023_),
    .X(_04002_));
 sg13g2_nand3b_1 _09649_ (.B(_05365_),
    .C(_04002_),
    .Y(_04003_),
    .A_N(net427));
 sg13g2_xnor2_1 _09650_ (.Y(_04004_),
    .A(_05365_),
    .B(_04002_));
 sg13g2_nand3_1 _09651_ (.B(net403),
    .C(_04004_),
    .A(net427),
    .Y(_04005_));
 sg13g2_o21ai_1 _09652_ (.B1(_04005_),
    .Y(_04006_),
    .A1(net403),
    .A2(_04003_));
 sg13g2_nor4_1 _09653_ (.A(net427),
    .B(_05365_),
    .C(_04002_),
    .D(net403),
    .Y(_04007_));
 sg13g2_a21oi_1 _09654_ (.A1(net279),
    .A2(_04006_),
    .Y(_04008_),
    .B1(_04007_));
 sg13g2_a21oi_1 _09655_ (.A1(_05165_),
    .A2(\dtop.vtop.pipeline.neg_t[5] ),
    .Y(_04009_),
    .B1(_04008_));
 sg13g2_nor3_1 _09656_ (.A(_04002_),
    .B(net403),
    .C(net279),
    .Y(_04010_));
 sg13g2_nor2_1 _09657_ (.A(_04009_),
    .B(_04010_),
    .Y(_04011_));
 sg13g2_nand2_1 _09658_ (.Y(_04012_),
    .A(_05385_),
    .B(net279));
 sg13g2_nand3_1 _09659_ (.B(net403),
    .C(net279),
    .A(net427),
    .Y(_04013_));
 sg13g2_o21ai_1 _09660_ (.B1(_04013_),
    .Y(_04014_),
    .A1(net427),
    .A2(_04001_));
 sg13g2_nand2_1 _09661_ (.Y(_04015_),
    .A(_05366_),
    .B(_04014_));
 sg13g2_o21ai_1 _09662_ (.B1(_04015_),
    .Y(_04016_),
    .A1(_04001_),
    .A2(net279));
 sg13g2_inv_1 _09663_ (.Y(_04017_),
    .A(\dtop.vtop.pipeline.neg_t[6] ));
 sg13g2_a21oi_1 _09664_ (.A1(net427),
    .A2(net279),
    .Y(_04018_),
    .B1(\dtop.vtop.pipeline.neg_t[7] ));
 sg13g2_a221oi_1 _09665_ (.B2(_04017_),
    .C1(_04018_),
    .B1(_04016_),
    .A1(_00027_),
    .Y(_04019_),
    .A2(_04012_));
 sg13g2_o21ai_1 _09666_ (.B1(_04019_),
    .Y(_04020_),
    .A1(_04000_),
    .A2(_04011_));
 sg13g2_or2_1 _09667_ (.X(_04021_),
    .B(_04012_),
    .A(_00027_));
 sg13g2_buf_1 _09668_ (.A(_00026_),
    .X(_04022_));
 sg13g2_a21oi_1 _09669_ (.A1(_04020_),
    .A2(_04021_),
    .Y(_04023_),
    .B1(_04022_));
 sg13g2_xnor2_1 _09670_ (.Y(_04024_),
    .A(_01509_),
    .B(_04023_));
 sg13g2_nand2_1 _09671_ (.Y(_04025_),
    .A(_03970_),
    .B(_04024_));
 sg13g2_a21oi_1 _09672_ (.A1(_03958_),
    .A2(_03969_),
    .Y(_04026_),
    .B1(_04025_));
 sg13g2_nor4_1 _09673_ (.A(_03891_),
    .B(_03897_),
    .C(_03916_),
    .D(_03917_),
    .Y(_04027_));
 sg13g2_nand2_1 _09674_ (.Y(_04028_),
    .A(_03273_),
    .B(_04027_));
 sg13g2_o21ai_1 _09675_ (.B1(_01487_),
    .Y(_04029_),
    .A1(_04026_),
    .A2(_04028_));
 sg13g2_a21o_1 _09676_ (.A2(_03918_),
    .A1(_03273_),
    .B1(_04029_),
    .X(_04030_));
 sg13g2_nor2_1 _09677_ (.A(\dtop.vtop.force_sat0 ),
    .B(\dtop.ext_control[6] ),
    .Y(_04031_));
 sg13g2_nand2_1 _09678_ (.Y(_04032_),
    .A(\dtop.vtop.logo_d[1] ),
    .B(_04031_));
 sg13g2_nor4_1 _09679_ (.A(_03891_),
    .B(_03897_),
    .C(_03888_),
    .D(_03887_),
    .Y(_04033_));
 sg13g2_o21ai_1 _09680_ (.B1(_04033_),
    .Y(_04034_),
    .A1(_03912_),
    .A2(_04032_));
 sg13g2_a21oi_1 _09681_ (.A1(_03914_),
    .A2(_04030_),
    .Y(_04035_),
    .B1(_04034_));
 sg13g2_buf_2 _09682_ (.A(_04035_),
    .X(_04036_));
 sg13g2_nand2b_1 _09683_ (.Y(_04037_),
    .B(_04036_),
    .A_N(_03911_));
 sg13g2_buf_1 _09684_ (.A(_04037_),
    .X(_04038_));
 sg13g2_nand2b_1 _09685_ (.Y(_04039_),
    .B(\dtop.vtop.force_sat0 ),
    .A_N(_03912_));
 sg13g2_buf_1 _09686_ (.A(\dtop.ext_control[4] ),
    .X(_04040_));
 sg13g2_buf_1 _09687_ (.A(_04040_),
    .X(_04041_));
 sg13g2_nor2_1 _09688_ (.A(net323),
    .B(_04041_),
    .Y(_04042_));
 sg13g2_buf_1 _09689_ (.A(_00013_),
    .X(_04043_));
 sg13g2_xor2_1 _09690_ (.B(_05298_),
    .A(net286),
    .X(_04044_));
 sg13g2_nand2_2 _09691_ (.Y(_04045_),
    .A(_04040_),
    .B(_04044_));
 sg13g2_inv_1 _09692_ (.Y(_04046_),
    .A(_00010_));
 sg13g2_xnor2_1 _09693_ (.Y(_04047_),
    .A(_04046_),
    .B(_04045_));
 sg13g2_and2_1 _09694_ (.A(net287),
    .B(_04040_),
    .X(_04048_));
 sg13g2_buf_1 _09695_ (.A(_04048_),
    .X(_04049_));
 sg13g2_nand3_1 _09696_ (.B(_04047_),
    .C(_04049_),
    .A(_03354_),
    .Y(_04050_));
 sg13g2_o21ai_1 _09697_ (.B1(_04050_),
    .Y(_04051_),
    .A1(_03357_),
    .A2(_04045_));
 sg13g2_a21oi_1 _09698_ (.A1(_04043_),
    .A2(_04051_),
    .Y(_04052_),
    .B1(_03384_));
 sg13g2_inv_1 _09699_ (.Y(_04053_),
    .A(_04043_));
 sg13g2_a21oi_1 _09700_ (.A1(_04053_),
    .A2(_04051_),
    .Y(_04054_),
    .B1(_04042_));
 sg13g2_a21oi_2 _09701_ (.B1(_04054_),
    .Y(_04055_),
    .A2(_04052_),
    .A1(_04042_));
 sg13g2_and2_1 _09702_ (.A(_00012_),
    .B(_04044_),
    .X(_04056_));
 sg13g2_buf_2 _09703_ (.A(_04056_),
    .X(_04057_));
 sg13g2_xnor2_1 _09704_ (.Y(_04058_),
    .A(_00009_),
    .B(_04057_));
 sg13g2_nand2_1 _09705_ (.Y(_04059_),
    .A(_04055_),
    .B(_04058_));
 sg13g2_nand2_1 _09706_ (.Y(_04060_),
    .A(\dtop.vtop.color[9] ),
    .B(_04057_));
 sg13g2_nand2_1 _09707_ (.Y(_04061_),
    .A(_04059_),
    .B(_04060_));
 sg13g2_nand4_1 _09708_ (.B(\dtop.vtop.color[11] ),
    .C(net276),
    .A(_03400_),
    .Y(_04062_),
    .D(_04061_));
 sg13g2_nand2_2 _09709_ (.Y(_04063_),
    .A(_04039_),
    .B(_04062_));
 sg13g2_buf_1 _09710_ (.A(net276),
    .X(_04064_));
 sg13g2_xor2_1 _09711_ (.B(_04061_),
    .A(_00008_),
    .X(_04065_));
 sg13g2_nor2_1 _09712_ (.A(_00514_),
    .B(\dtop.out_sample[6] ),
    .Y(_04066_));
 sg13g2_inv_1 _09713_ (.Y(_04067_),
    .A(\dtop.out_sample[2] ));
 sg13g2_nor2b_1 _09714_ (.A(net287),
    .B_N(\dtop.out_sample[0] ),
    .Y(_04068_));
 sg13g2_nor2_1 _09715_ (.A(\dtop.out_sample[1] ),
    .B(_04068_),
    .Y(_04069_));
 sg13g2_nor2_1 _09716_ (.A(_00465_),
    .B(_04069_),
    .Y(_04070_));
 sg13g2_a221oi_1 _09717_ (.B2(_04068_),
    .C1(_04070_),
    .B1(\dtop.out_sample[1] ),
    .A1(net300),
    .Y(_04071_),
    .A2(\dtop.out_sample[2] ));
 sg13g2_a21oi_1 _09718_ (.A1(_01807_),
    .A2(_04067_),
    .Y(_04072_),
    .B1(_04071_));
 sg13g2_nor2_1 _09719_ (.A(\dtop.out_sample[3] ),
    .B(_04072_),
    .Y(_04073_));
 sg13g2_a21oi_1 _09720_ (.A1(\dtop.out_sample[3] ),
    .A2(_04072_),
    .Y(_04074_),
    .B1(net326));
 sg13g2_nand2b_1 _09721_ (.Y(_04075_),
    .B(\dtop.out_sample[4] ),
    .A_N(net297));
 sg13g2_o21ai_1 _09722_ (.B1(_04075_),
    .Y(_04076_),
    .A1(_04073_),
    .A2(_04074_));
 sg13g2_inv_1 _09723_ (.Y(_04077_),
    .A(\dtop.out_sample[5] ));
 sg13g2_inv_1 _09724_ (.Y(_04078_),
    .A(\dtop.out_sample[4] ));
 sg13g2_a22oi_1 _09725_ (.Y(_04079_),
    .B1(_04078_),
    .B2(_00507_),
    .A2(_04077_),
    .A1(_00539_));
 sg13g2_a22oi_1 _09726_ (.Y(_04080_),
    .B1(_04076_),
    .B2(_04079_),
    .A2(\dtop.out_sample[5] ),
    .A1(_00504_));
 sg13g2_nand2_1 _09727_ (.Y(_04081_),
    .A(_00514_),
    .B(\dtop.out_sample[6] ));
 sg13g2_o21ai_1 _09728_ (.B1(_04081_),
    .Y(_04082_),
    .A1(_04066_),
    .A2(_04080_));
 sg13g2_xnor2_1 _09729_ (.Y(_04083_),
    .A(_05182_),
    .B(_04082_));
 sg13g2_a21oi_1 _09730_ (.A1(_00944_),
    .A2(_04083_),
    .Y(_04084_),
    .B1(net276));
 sg13g2_a21oi_1 _09731_ (.A1(net264),
    .A2(_04065_),
    .Y(_04085_),
    .B1(_04084_));
 sg13g2_nor2_1 _09732_ (.A(_04063_),
    .B(_04085_),
    .Y(_04086_));
 sg13g2_xnor2_1 _09733_ (.Y(_04087_),
    .A(_04043_),
    .B(_04051_));
 sg13g2_a21oi_1 _09734_ (.A1(net264),
    .A2(_04087_),
    .Y(_04088_),
    .B1(_04063_));
 sg13g2_mux2_1 _09735_ (.A0(_04086_),
    .A1(_04088_),
    .S(net361),
    .X(_04089_));
 sg13g2_nand2b_1 _09736_ (.Y(_04090_),
    .B(net16),
    .A_N(net362));
 sg13g2_o21ai_1 _09737_ (.B1(_04090_),
    .Y(_00377_),
    .A1(_04038_),
    .A2(_04089_));
 sg13g2_nand3_1 _09738_ (.B(_04055_),
    .C(_04058_),
    .A(_03400_),
    .Y(_04091_));
 sg13g2_o21ai_1 _09739_ (.B1(_04091_),
    .Y(_04092_),
    .A1(_00008_),
    .A2(_04060_));
 sg13g2_xor2_1 _09740_ (.B(_04092_),
    .A(_00007_),
    .X(_04093_));
 sg13g2_a21oi_1 _09741_ (.A1(_05174_),
    .A2(_04083_),
    .Y(_04094_),
    .B1(_04064_));
 sg13g2_a21oi_1 _09742_ (.A1(net264),
    .A2(_04093_),
    .Y(_04095_),
    .B1(_04094_));
 sg13g2_nor2_1 _09743_ (.A(_04063_),
    .B(_04095_),
    .Y(_04096_));
 sg13g2_xor2_1 _09744_ (.B(_04058_),
    .A(_04055_),
    .X(_04097_));
 sg13g2_a21oi_1 _09745_ (.A1(net264),
    .A2(_04097_),
    .Y(_04098_),
    .B1(_04063_));
 sg13g2_mux2_1 _09746_ (.A0(_04096_),
    .A1(_04098_),
    .S(net361),
    .X(_04099_));
 sg13g2_nand2b_1 _09747_ (.Y(_04100_),
    .B(net17),
    .A_N(net362));
 sg13g2_o21ai_1 _09748_ (.B1(_04100_),
    .Y(_00378_),
    .A1(_04038_),
    .A2(_04099_));
 sg13g2_nand2b_1 _09749_ (.Y(_04101_),
    .B(net18),
    .A_N(net362));
 sg13g2_o21ai_1 _09750_ (.B1(_04101_),
    .Y(_00379_),
    .A1(_04038_),
    .A2(_04086_));
 sg13g2_nand2b_1 _09751_ (.Y(_04102_),
    .B(net19),
    .A_N(net362));
 sg13g2_o21ai_1 _09752_ (.B1(_04102_),
    .Y(_00380_),
    .A1(_04038_),
    .A2(_04096_));
 sg13g2_nand2b_1 _09753_ (.Y(_04103_),
    .B(net20),
    .A_N(net362));
 sg13g2_o21ai_1 _09754_ (.B1(_04103_),
    .Y(_00381_),
    .A1(_03905_),
    .A2(_03911_));
 sg13g2_inv_1 _09755_ (.Y(_04104_),
    .A(net21));
 sg13g2_buf_1 _09756_ (.A(_03910_),
    .X(_04105_));
 sg13g2_nand3_1 _09757_ (.B(net360),
    .C(\uio_out0b[5] ),
    .A(net374),
    .Y(_04106_));
 sg13g2_o21ai_1 _09758_ (.B1(_04106_),
    .Y(_00382_),
    .A1(net337),
    .A2(_04104_));
 sg13g2_nand3_1 _09759_ (.B(_03907_),
    .C(_04083_),
    .A(_00082_),
    .Y(_04107_));
 sg13g2_o21ai_1 _09760_ (.B1(_04107_),
    .Y(_04108_),
    .A1(_01189_),
    .A2(net22));
 sg13g2_inv_1 _09761_ (.Y(_00383_),
    .A(_04108_));
 sg13g2_inv_1 _09762_ (.Y(_04109_),
    .A(net23));
 sg13g2_o21ai_1 _09763_ (.B1(_04107_),
    .Y(_00384_),
    .A1(net337),
    .A2(_04109_));
 sg13g2_inv_1 _09764_ (.Y(_04110_),
    .A(net24));
 sg13g2_nor4_1 _09765_ (.A(_02282_),
    .B(_02280_),
    .C(_02850_),
    .D(_04027_),
    .Y(_04111_));
 sg13g2_o21ai_1 _09766_ (.B1(_03914_),
    .Y(_04112_),
    .A1(_04029_),
    .A2(_04111_));
 sg13g2_nor2b_2 _09767_ (.A(_04034_),
    .B_N(_04112_),
    .Y(_04113_));
 sg13g2_or2_1 _09768_ (.X(_04114_),
    .B(_04083_),
    .A(net276));
 sg13g2_or2_1 _09769_ (.X(_04115_),
    .B(_03305_),
    .A(_03277_));
 sg13g2_buf_1 _09770_ (.A(_04115_),
    .X(_04116_));
 sg13g2_nor2_1 _09771_ (.A(_03882_),
    .B(_03311_),
    .Y(_04117_));
 sg13g2_nor2_2 _09772_ (.A(_03309_),
    .B(net363),
    .Y(_04118_));
 sg13g2_and2_1 _09773_ (.A(_03400_),
    .B(_04118_),
    .X(_04119_));
 sg13g2_nor2_1 _09774_ (.A(_03400_),
    .B(_04118_),
    .Y(_04120_));
 sg13g2_or2_1 _09775_ (.X(_04121_),
    .B(_03384_),
    .A(_03274_));
 sg13g2_nand2b_1 _09776_ (.Y(_04122_),
    .B(_03277_),
    .A_N(\dtop.vtop.color[9] ));
 sg13g2_o21ai_1 _09777_ (.B1(_04122_),
    .Y(_04123_),
    .A1(_03386_),
    .A2(_04116_));
 sg13g2_a22oi_1 _09778_ (.Y(_04124_),
    .B1(_04121_),
    .B2(_04123_),
    .A2(_03386_),
    .A1(net363));
 sg13g2_nor2_1 _09779_ (.A(net408),
    .B(_03305_),
    .Y(_04125_));
 sg13g2_mux2_1 _09780_ (.A0(net408),
    .A1(_04125_),
    .S(_03356_),
    .X(_04126_));
 sg13g2_nand2_1 _09781_ (.Y(_04127_),
    .A(_03284_),
    .B(_00011_));
 sg13g2_and2_1 _09782_ (.A(_00010_),
    .B(_03356_),
    .X(_04128_));
 sg13g2_o21ai_1 _09783_ (.B1(_03384_),
    .Y(_04129_),
    .A1(_03274_),
    .A2(net363));
 sg13g2_o21ai_1 _09784_ (.B1(_04129_),
    .Y(_04130_),
    .A1(_03306_),
    .A2(_04128_));
 sg13g2_a221oi_1 _09785_ (.B2(_04127_),
    .C1(_04130_),
    .B1(_04126_),
    .A1(net408),
    .Y(_04131_),
    .A2(_04046_));
 sg13g2_nand2b_1 _09786_ (.Y(_04132_),
    .B(_04116_),
    .A_N(_00009_));
 sg13g2_o21ai_1 _09787_ (.B1(_04132_),
    .Y(_04133_),
    .A1(_04124_),
    .A2(_04131_));
 sg13g2_o21ai_1 _09788_ (.B1(_04133_),
    .Y(_04134_),
    .A1(_04119_),
    .A2(_04120_));
 sg13g2_or2_1 _09789_ (.X(_04135_),
    .B(_04118_),
    .A(_00008_));
 sg13g2_a221oi_1 _09790_ (.B2(_03309_),
    .C1(_03400_),
    .B1(_04126_),
    .A1(net363),
    .Y(_04136_),
    .A2(_03357_));
 sg13g2_xor2_1 _09791_ (.B(_03356_),
    .A(net408),
    .X(_04137_));
 sg13g2_inv_1 _09792_ (.Y(_04138_),
    .A(_03400_));
 sg13g2_a21oi_1 _09793_ (.A1(_04118_),
    .A2(_04137_),
    .Y(_04139_),
    .B1(_04138_));
 sg13g2_o21ai_1 _09794_ (.B1(net363),
    .Y(_04140_),
    .A1(_03384_),
    .A2(_03354_));
 sg13g2_nor2_1 _09795_ (.A(_03283_),
    .B(net363),
    .Y(_04141_));
 sg13g2_nand2b_1 _09796_ (.Y(_04142_),
    .B(_04141_),
    .A_N(_03354_));
 sg13g2_a22oi_1 _09797_ (.Y(_04143_),
    .B1(_03354_),
    .B2(_03283_),
    .A2(_03384_),
    .A1(_03274_));
 sg13g2_nand3_1 _09798_ (.B(_04142_),
    .C(_04143_),
    .A(_04140_),
    .Y(_04144_));
 sg13g2_nor4_1 _09799_ (.A(_04124_),
    .B(_04136_),
    .C(_04139_),
    .D(_04144_),
    .Y(_04145_));
 sg13g2_a21o_1 _09800_ (.A2(_04135_),
    .A1(_04134_),
    .B1(_04145_),
    .X(_04146_));
 sg13g2_nand2_1 _09801_ (.Y(_04147_),
    .A(_04117_),
    .B(_04146_));
 sg13g2_o21ai_1 _09802_ (.B1(_00007_),
    .Y(_04148_),
    .A1(_04117_),
    .A2(_04146_));
 sg13g2_nand2_1 _09803_ (.Y(_04149_),
    .A(_04147_),
    .B(_04148_));
 sg13g2_buf_2 _09804_ (.A(_04149_),
    .X(_04150_));
 sg13g2_mux2_1 _09805_ (.A0(_04116_),
    .A1(_00009_),
    .S(_04150_),
    .X(_04151_));
 sg13g2_a21oi_1 _09806_ (.A1(_03275_),
    .A2(_03306_),
    .Y(_04152_),
    .B1(_04150_));
 sg13g2_a21oi_2 _09807_ (.B1(_04152_),
    .Y(_04153_),
    .A2(_04150_),
    .A1(_04043_));
 sg13g2_mux2_1 _09808_ (.A0(_04141_),
    .A1(_03354_),
    .S(_04150_),
    .X(_04154_));
 sg13g2_mux2_1 _09809_ (.A0(_04125_),
    .A1(_04046_),
    .S(_04150_),
    .X(_04155_));
 sg13g2_a21oi_1 _09810_ (.A1(_04049_),
    .A2(_04154_),
    .Y(_04156_),
    .B1(_04155_));
 sg13g2_nand3_1 _09811_ (.B(_04154_),
    .C(_04155_),
    .A(_04049_),
    .Y(_04157_));
 sg13g2_o21ai_1 _09812_ (.B1(_04157_),
    .Y(_04158_),
    .A1(_04045_),
    .A2(_04156_));
 sg13g2_nand2_1 _09813_ (.Y(_04159_),
    .A(_04153_),
    .B(_04158_));
 sg13g2_o21ai_1 _09814_ (.B1(_04042_),
    .Y(_04160_),
    .A1(_04153_),
    .A2(_04158_));
 sg13g2_nand3_1 _09815_ (.B(_04159_),
    .C(_04160_),
    .A(_04151_),
    .Y(_04161_));
 sg13g2_a21oi_1 _09816_ (.A1(_04159_),
    .A2(_04160_),
    .Y(_04162_),
    .B1(_04151_));
 sg13g2_a21oi_1 _09817_ (.A1(_04057_),
    .A2(_04161_),
    .Y(_04163_),
    .B1(_04162_));
 sg13g2_mux2_1 _09818_ (.A0(_04118_),
    .A1(_03400_),
    .S(_04150_),
    .X(_04164_));
 sg13g2_nand2b_1 _09819_ (.Y(_04165_),
    .B(_04164_),
    .A_N(_04163_));
 sg13g2_nand2b_1 _09820_ (.Y(_04166_),
    .B(_04117_),
    .A_N(_00007_));
 sg13g2_nand3_1 _09821_ (.B(_04165_),
    .C(_04166_),
    .A(net276),
    .Y(_04167_));
 sg13g2_a21oi_1 _09822_ (.A1(_04114_),
    .A2(_04167_),
    .Y(_04168_),
    .B1(_03913_));
 sg13g2_xor2_1 _09823_ (.B(_04158_),
    .A(_04153_),
    .X(_04169_));
 sg13g2_nand2_1 _09824_ (.Y(_04170_),
    .A(net264),
    .B(_04169_));
 sg13g2_nand2b_1 _09825_ (.Y(_04171_),
    .B(_04163_),
    .A_N(_04164_));
 sg13g2_and3_1 _09826_ (.X(_04172_),
    .A(net264),
    .B(_04165_),
    .C(_04171_));
 sg13g2_nor2_1 _09827_ (.A(net361),
    .B(_04172_),
    .Y(_04173_));
 sg13g2_a21oi_1 _09828_ (.A1(net361),
    .A2(_04170_),
    .Y(_04174_),
    .B1(_04173_));
 sg13g2_o21ai_1 _09829_ (.B1(net276),
    .Y(_04175_),
    .A1(_04165_),
    .A2(_04166_));
 sg13g2_a21o_1 _09830_ (.A2(_04175_),
    .A1(_04114_),
    .B1(_03913_),
    .X(_04176_));
 sg13g2_o21ai_1 _09831_ (.B1(net360),
    .Y(_04177_),
    .A1(_04174_),
    .A2(_04176_));
 sg13g2_o21ai_1 _09832_ (.B1(_04177_),
    .Y(_04178_),
    .A1(net360),
    .A2(_04168_));
 sg13g2_nand3_1 _09833_ (.B(_04113_),
    .C(_04178_),
    .A(net374),
    .Y(_04179_));
 sg13g2_o21ai_1 _09834_ (.B1(_04179_),
    .Y(_00385_),
    .A1(net337),
    .A2(_04110_));
 sg13g2_nand2_1 _09835_ (.Y(_04180_),
    .A(_04159_),
    .B(_04160_));
 sg13g2_xor2_1 _09836_ (.B(_04151_),
    .A(_04057_),
    .X(_04181_));
 sg13g2_xnor2_1 _09837_ (.Y(_04182_),
    .A(_04180_),
    .B(_04181_));
 sg13g2_a21oi_1 _09838_ (.A1(_04064_),
    .A2(_04182_),
    .Y(_04183_),
    .B1(_04176_));
 sg13g2_nor2b_1 _09839_ (.A(net361),
    .B_N(_04168_),
    .Y(_04184_));
 sg13g2_a21oi_1 _09840_ (.A1(_04041_),
    .A2(_04183_),
    .Y(_04185_),
    .B1(_04184_));
 sg13g2_and2_1 _09841_ (.A(_04113_),
    .B(_04185_),
    .X(_04186_));
 sg13g2_nor2_1 _09842_ (.A(net360),
    .B(_04096_),
    .Y(_04187_));
 sg13g2_a22oi_1 _09843_ (.Y(_04188_),
    .B1(_04187_),
    .B2(_04036_),
    .A2(_04186_),
    .A1(net360));
 sg13g2_nor2_1 _09844_ (.A(net374),
    .B(net25),
    .Y(_04189_));
 sg13g2_a21oi_1 _09845_ (.A1(net337),
    .A2(_04188_),
    .Y(_00386_),
    .B1(_04189_));
 sg13g2_o21ai_1 _09846_ (.B1(_04113_),
    .Y(_04190_),
    .A1(_04172_),
    .A2(_04176_));
 sg13g2_o21ai_1 _09847_ (.B1(_04040_),
    .Y(_04191_),
    .A1(net408),
    .A2(_04045_));
 sg13g2_o21ai_1 _09848_ (.B1(_04045_),
    .Y(_04192_),
    .A1(net323),
    .A2(_03296_));
 sg13g2_a22oi_1 _09849_ (.Y(_04193_),
    .B1(_04192_),
    .B2(_03275_),
    .A2(_04191_),
    .A1(net287));
 sg13g2_nor2_1 _09850_ (.A(_03277_),
    .B(_04193_),
    .Y(_04194_));
 sg13g2_nand2_1 _09851_ (.Y(_04195_),
    .A(_04057_),
    .B(_04194_));
 sg13g2_nand2_1 _09852_ (.Y(_04196_),
    .A(_03309_),
    .B(_04195_));
 sg13g2_o21ai_1 _09853_ (.B1(_04196_),
    .Y(_04197_),
    .A1(_04057_),
    .A2(_04194_));
 sg13g2_or2_1 _09854_ (.X(_04198_),
    .B(_04197_),
    .A(_03311_));
 sg13g2_and3_1 _09855_ (.X(_04199_),
    .A(_03882_),
    .B(net264),
    .C(_04198_));
 sg13g2_o21ai_1 _09856_ (.B1(_04039_),
    .Y(_04200_),
    .A1(_04094_),
    .A2(_04199_));
 sg13g2_nand2_1 _09857_ (.Y(_04201_),
    .A(_04036_),
    .B(_04200_));
 sg13g2_inv_1 _09858_ (.Y(_04202_),
    .A(net360));
 sg13g2_mux2_1 _09859_ (.A0(_04190_),
    .A1(_04201_),
    .S(_04202_),
    .X(_04203_));
 sg13g2_nor2_1 _09860_ (.A(net374),
    .B(net26),
    .Y(_04204_));
 sg13g2_a21oi_1 _09861_ (.A1(net337),
    .A2(_04203_),
    .Y(_00387_),
    .B1(_04204_));
 sg13g2_nor2_1 _09862_ (.A(_04202_),
    .B(_04168_),
    .Y(_04205_));
 sg13g2_a22oi_1 _09863_ (.Y(_04206_),
    .B1(_04113_),
    .B2(_04205_),
    .A2(\uio_out0b[5] ),
    .A1(_04202_));
 sg13g2_nor2_1 _09864_ (.A(net374),
    .B(net27),
    .Y(_04207_));
 sg13g2_a21oi_1 _09865_ (.A1(net337),
    .A2(_04206_),
    .Y(_00388_),
    .B1(_04207_));
 sg13g2_nand2_1 _09866_ (.Y(_04208_),
    .A(_03311_),
    .B(_04197_));
 sg13g2_a21oi_1 _09867_ (.A1(_04198_),
    .A2(_04208_),
    .Y(_04209_),
    .B1(_01600_));
 sg13g2_nor4_1 _09868_ (.A(net363),
    .B(_03311_),
    .C(_01600_),
    .D(_04197_),
    .Y(_04210_));
 sg13g2_nor2_1 _09869_ (.A(_03913_),
    .B(_04210_),
    .Y(_04211_));
 sg13g2_o21ai_1 _09870_ (.B1(_04211_),
    .Y(_04212_),
    .A1(_04084_),
    .A2(_04209_));
 sg13g2_xnor2_1 _09871_ (.Y(_04213_),
    .A(_03277_),
    .B(_04193_));
 sg13g2_o21ai_1 _09872_ (.B1(_04211_),
    .Y(_04214_),
    .A1(_01600_),
    .A2(_04213_));
 sg13g2_mux2_1 _09873_ (.A0(_04212_),
    .A1(_04214_),
    .S(net361),
    .X(_04215_));
 sg13g2_nand3_1 _09874_ (.B(_04036_),
    .C(_04215_),
    .A(net360),
    .Y(_04216_));
 sg13g2_o21ai_1 _09875_ (.B1(_04216_),
    .Y(_04217_),
    .A1(_04105_),
    .A2(_04190_));
 sg13g2_mux2_1 _09876_ (.A0(net28),
    .A1(_04217_),
    .S(_01189_),
    .X(_00389_));
 sg13g2_inv_1 _09877_ (.Y(_04218_),
    .A(net29));
 sg13g2_xor2_1 _09878_ (.B(_04057_),
    .A(_03309_),
    .X(_04219_));
 sg13g2_xnor2_1 _09879_ (.Y(_04220_),
    .A(_04194_),
    .B(_04219_));
 sg13g2_nand2_1 _09880_ (.Y(_04221_),
    .A(net264),
    .B(_04220_));
 sg13g2_nand3_1 _09881_ (.B(_04211_),
    .C(_04221_),
    .A(net361),
    .Y(_04222_));
 sg13g2_o21ai_1 _09882_ (.B1(_04222_),
    .Y(_04223_),
    .A1(net361),
    .A2(_04200_));
 sg13g2_nor3_1 _09883_ (.A(_03910_),
    .B(_04063_),
    .C(_04085_),
    .Y(_04224_));
 sg13g2_a21oi_1 _09884_ (.A1(net360),
    .A2(_04223_),
    .Y(_04225_),
    .B1(_04224_));
 sg13g2_nand3_1 _09885_ (.B(_04036_),
    .C(_04225_),
    .A(net362),
    .Y(_04226_));
 sg13g2_o21ai_1 _09886_ (.B1(_04226_),
    .Y(_00390_),
    .A1(net337),
    .A2(_04218_));
 sg13g2_inv_1 _09887_ (.Y(_04227_),
    .A(net30));
 sg13g2_nand3_1 _09888_ (.B(_04036_),
    .C(_04212_),
    .A(net362),
    .Y(_04228_));
 sg13g2_o21ai_1 _09889_ (.B1(_04228_),
    .Y(_00391_),
    .A1(_03908_),
    .A2(_04227_));
 sg13g2_mux2_1 _09890_ (.A0(_03905_),
    .A1(_04201_),
    .S(_04105_),
    .X(_04229_));
 sg13g2_nor2_1 _09891_ (.A(net374),
    .B(net31),
    .Y(_04230_));
 sg13g2_a21oi_1 _09892_ (.A1(_03908_),
    .A2(_04229_),
    .Y(_00392_),
    .B1(_04230_));
 sg13g2_mux2_1 _09893_ (.A0(_01188_),
    .A1(\dtop.vtop.force_sat0 ),
    .S(net374),
    .X(_00097_));
 sg13g2_buf_1 _09894_ (.A(net216),
    .X(_04231_));
 sg13g2_nand3_1 _09895_ (.B(net306),
    .C(_03338_),
    .A(_03336_),
    .Y(_04232_));
 sg13g2_o21ai_1 _09896_ (.B1(_04232_),
    .Y(_04233_),
    .A1(net306),
    .A2(_03338_));
 sg13g2_buf_1 _09897_ (.A(net216),
    .X(_04234_));
 sg13g2_a21oi_1 _09898_ (.A1(net174),
    .A2(_03338_),
    .Y(_04235_),
    .B1(_03336_));
 sg13g2_a21oi_1 _09899_ (.A1(net175),
    .A2(_04233_),
    .Y(_00213_),
    .B1(_04235_));
 sg13g2_nand2_1 _09900_ (.Y(_04236_),
    .A(net306),
    .B(_03339_));
 sg13g2_nand3_1 _09901_ (.B(_03340_),
    .C(_04236_),
    .A(net174),
    .Y(_04237_));
 sg13g2_nand2_1 _09902_ (.Y(_04238_),
    .A(_03336_),
    .B(_03338_));
 sg13g2_nor2_1 _09903_ (.A(_02477_),
    .B(_04232_),
    .Y(_04239_));
 sg13g2_a21oi_1 _09904_ (.A1(_02477_),
    .A2(_04238_),
    .Y(_04240_),
    .B1(_04239_));
 sg13g2_nand2_1 _09905_ (.Y(_04241_),
    .A(_02477_),
    .B(net338));
 sg13g2_o21ai_1 _09906_ (.B1(_04241_),
    .Y(_04242_),
    .A1(\dtop.vtop.pipeline.cosappr_acc[1] ),
    .A2(_04240_));
 sg13g2_a22oi_1 _09907_ (.Y(_04243_),
    .B1(_04242_),
    .B2(net175),
    .A2(_04237_),
    .A1(\dtop.vtop.pipeline.cosappr_acc[1] ));
 sg13g2_inv_1 _09908_ (.Y(_00214_),
    .A(_04243_));
 sg13g2_buf_1 _09909_ (.A(_03271_),
    .X(_04244_));
 sg13g2_nor2_1 _09910_ (.A(net338),
    .B(_03344_),
    .Y(_04245_));
 sg13g2_mux2_1 _09911_ (.A0(_03344_),
    .A1(_04245_),
    .S(_03342_),
    .X(_04246_));
 sg13g2_inv_1 _09912_ (.Y(_04247_),
    .A(\dtop.vtop.pipeline.cosappr_acc[2] ));
 sg13g2_a22oi_1 _09913_ (.Y(_04248_),
    .B1(_04246_),
    .B2(_04247_),
    .A2(_03344_),
    .A1(net338));
 sg13g2_nor3_1 _09914_ (.A(net338),
    .B(_03342_),
    .C(_03344_),
    .Y(_04249_));
 sg13g2_nand2_1 _09915_ (.Y(_04250_),
    .A(net216),
    .B(_03345_));
 sg13g2_o21ai_1 _09916_ (.B1(\dtop.vtop.pipeline.cosappr_acc[2] ),
    .Y(_04251_),
    .A1(_04249_),
    .A2(_04250_));
 sg13g2_o21ai_1 _09917_ (.B1(_04251_),
    .Y(_00215_),
    .A1(net210),
    .A2(_04248_));
 sg13g2_nand2_1 _09918_ (.Y(_04252_),
    .A(net174),
    .B(_03352_));
 sg13g2_a21oi_1 _09919_ (.A1(net306),
    .A2(_03349_),
    .Y(_04253_),
    .B1(net210));
 sg13g2_nand2b_1 _09920_ (.Y(_04254_),
    .B(\dtop.vtop.pipeline.cosappr_acc[3] ),
    .A_N(_04253_));
 sg13g2_o21ai_1 _09921_ (.B1(_04254_),
    .Y(_00216_),
    .A1(_03349_),
    .A2(_04252_));
 sg13g2_mux2_1 _09922_ (.A0(_03367_),
    .A1(_03373_),
    .S(_04231_),
    .X(_00217_));
 sg13g2_and2_1 _09923_ (.A(_03359_),
    .B(_03382_),
    .X(_04255_));
 sg13g2_a22oi_1 _09924_ (.Y(_04256_),
    .B1(_03381_),
    .B2(_04255_),
    .A2(_04244_),
    .A1(\dtop.vtop.pipeline.cosappr_acc[5] ));
 sg13g2_o21ai_1 _09925_ (.B1(_04256_),
    .Y(_00218_),
    .A1(_03381_),
    .A2(_03382_));
 sg13g2_mux2_1 _09926_ (.A0(\dtop.vtop.pipeline.cosappr_acc[6] ),
    .A1(_03392_),
    .S(_04231_),
    .X(_00219_));
 sg13g2_nand2_1 _09927_ (.Y(_04257_),
    .A(\dtop.vtop.pipeline.cosappr_acc[7] ),
    .B(net210));
 sg13g2_o21ai_1 _09928_ (.B1(_04257_),
    .Y(_00220_),
    .A1(net210),
    .A2(_03399_));
 sg13g2_mux2_1 _09929_ (.A0(\dtop.vtop.pipeline.cosappr_acc[8] ),
    .A1(_03403_),
    .S(net175),
    .X(_00221_));
 sg13g2_nor2_1 _09930_ (.A(net210),
    .B(_03759_),
    .Y(_04258_));
 sg13g2_a22oi_1 _09931_ (.Y(_04259_),
    .B1(_04258_),
    .B2(_03050_),
    .A2(net210),
    .A1(_02356_));
 sg13g2_o21ai_1 _09932_ (.B1(_04259_),
    .Y(_00325_),
    .A1(_03050_),
    .A2(_03785_));
 sg13g2_mux2_1 _09933_ (.A0(\dtop.vtop.pipeline.zg_acc[1] ),
    .A1(_03766_),
    .S(net175),
    .X(_00326_));
 sg13g2_nand2_1 _09934_ (.Y(_04260_),
    .A(net174),
    .B(_03774_));
 sg13g2_o21ai_1 _09935_ (.B1(_04260_),
    .Y(_00327_),
    .A1(_02299_),
    .A2(net175));
 sg13g2_nor2_1 _09936_ (.A(_04244_),
    .B(_03799_),
    .Y(_04261_));
 sg13g2_o21ai_1 _09937_ (.B1(_04261_),
    .Y(_04262_),
    .A1(_03762_),
    .A2(_03800_));
 sg13g2_nand3_1 _09938_ (.B(_03769_),
    .C(_03805_),
    .A(_03248_),
    .Y(_04263_));
 sg13g2_o21ai_1 _09939_ (.B1(_04263_),
    .Y(_04264_),
    .A1(_03248_),
    .A2(_03805_));
 sg13g2_a22oi_1 _09940_ (.Y(_04265_),
    .B1(_04264_),
    .B2(_02399_),
    .A2(_03762_),
    .A1(_03194_));
 sg13g2_inv_1 _09941_ (.Y(_04266_),
    .A(_04265_));
 sg13g2_a22oi_1 _09942_ (.Y(_00328_),
    .B1(_04266_),
    .B2(net175),
    .A2(_04262_),
    .A1(_02400_));
 sg13g2_mux2_1 _09943_ (.A0(_02455_),
    .A1(_03804_),
    .S(net174),
    .X(_00329_));
 sg13g2_nand2_1 _09944_ (.Y(_04267_),
    .A(_03832_),
    .B(_03834_));
 sg13g2_o21ai_1 _09945_ (.B1(_04267_),
    .Y(_04268_),
    .A1(net33),
    .A2(net211));
 sg13g2_a21oi_1 _09946_ (.A1(_04234_),
    .A2(_03832_),
    .Y(_04269_),
    .B1(_02553_));
 sg13g2_a21oi_1 _09947_ (.A1(net175),
    .A2(_04268_),
    .Y(_00330_),
    .B1(_04269_));
 sg13g2_mux2_1 _09948_ (.A0(\dtop.vtop.pipeline.zg_acc[6] ),
    .A1(_03842_),
    .S(net174),
    .X(_00331_));
 sg13g2_and3_1 _09949_ (.X(_04270_),
    .A(net410),
    .B(net216),
    .C(net211));
 sg13g2_nor2_1 _09950_ (.A(net410),
    .B(net210),
    .Y(_04271_));
 sg13g2_and2_1 _09951_ (.A(net216),
    .B(_03846_),
    .X(_04272_));
 sg13g2_and2_1 _09952_ (.A(net410),
    .B(net216),
    .X(_04273_));
 sg13g2_mux4_1 _09953_ (.S0(_03251_),
    .A0(_04270_),
    .A1(_04271_),
    .A2(_04272_),
    .A3(_04273_),
    .S1(_03852_),
    .X(_04274_));
 sg13g2_nand3_1 _09954_ (.B(net216),
    .C(net212),
    .A(_03251_),
    .Y(_04275_));
 sg13g2_o21ai_1 _09955_ (.B1(_04275_),
    .Y(_04276_),
    .A1(\dtop.vtop.pipeline.zg_acc[7] ),
    .A2(net174));
 sg13g2_nor2_1 _09956_ (.A(_04274_),
    .B(_04276_),
    .Y(_00332_));
 sg13g2_mux2_1 _09957_ (.A0(\dtop.vtop.pipeline.zg_acc[8] ),
    .A1(_03872_),
    .S(_04234_),
    .X(_00333_));
 sg13g2_nor2_1 _09958_ (.A(net217),
    .B(net141),
    .Y(_04277_));
 sg13g2_and2_1 _09959_ (.A(net217),
    .B(net141),
    .X(_04278_));
 sg13g2_mux2_1 _09960_ (.A0(_04277_),
    .A1(_04278_),
    .S(_03865_),
    .X(_04279_));
 sg13g2_nor2_1 _09961_ (.A(\dtop.vtop.pipeline.zg_acc[9] ),
    .B(net212),
    .Y(_04280_));
 sg13g2_a21oi_1 _09962_ (.A1(\dtop.vtop.pipeline.zg_acc[9] ),
    .A2(net210),
    .Y(_04281_),
    .B1(_04280_));
 sg13g2_or3_1 _09963_ (.A(net217),
    .B(_03271_),
    .C(_03870_),
    .X(_04282_));
 sg13g2_nand3_1 _09964_ (.B(net216),
    .C(net141),
    .A(net217),
    .Y(_04283_));
 sg13g2_mux2_1 _09965_ (.A0(_04282_),
    .A1(_04283_),
    .S(_03865_),
    .X(_04284_));
 sg13g2_a21oi_1 _09966_ (.A1(net174),
    .A2(net212),
    .Y(_04285_),
    .B1(\dtop.vtop.pipeline.zg_acc[9] ));
 sg13g2_a22oi_1 _09967_ (.Y(_00334_),
    .B1(_04284_),
    .B2(_04285_),
    .A2(_04281_),
    .A1(_04279_));
 sg13g2_buf_1 _09968_ (.A(net267),
    .X(_04286_));
 sg13g2_nand4_1 _09969_ (.B(_03970_),
    .C(_03360_),
    .A(\dtop.vtop.pipeline.zg_valid ),
    .Y(_04287_),
    .D(_03958_));
 sg13g2_buf_1 _09970_ (.A(_04287_),
    .X(_04288_));
 sg13g2_buf_1 _09971_ (.A(net40),
    .X(_04289_));
 sg13g2_nand2_1 _09972_ (.Y(_04290_),
    .A(_03927_),
    .B(net37));
 sg13g2_nor2_1 _09973_ (.A(net407),
    .B(_03410_),
    .Y(_04291_));
 sg13g2_xnor2_1 _09974_ (.Y(_04292_),
    .A(_03982_),
    .B(_04291_));
 sg13g2_buf_1 _09975_ (.A(_00088_),
    .X(_04293_));
 sg13g2_o21ai_1 _09976_ (.B1(_04293_),
    .Y(_04294_),
    .A1(_03317_),
    .A2(_03324_));
 sg13g2_o21ai_1 _09977_ (.B1(_04294_),
    .Y(_04295_),
    .A1(net215),
    .A2(_04292_));
 sg13g2_nand2b_1 _09978_ (.Y(_04296_),
    .B(_04295_),
    .A_N(net40));
 sg13g2_nand3_1 _09979_ (.B(_04290_),
    .C(_04296_),
    .A(_04286_),
    .Y(_00222_));
 sg13g2_nand2_1 _09980_ (.Y(_04297_),
    .A(_03981_),
    .B(_04291_));
 sg13g2_o21ai_1 _09981_ (.B1(_04294_),
    .Y(_04298_),
    .A1(_03326_),
    .A2(_04297_));
 sg13g2_buf_1 _09982_ (.A(_04298_),
    .X(_04299_));
 sg13g2_nor2b_1 _09983_ (.A(_03411_),
    .B_N(_03405_),
    .Y(_04300_));
 sg13g2_xnor2_1 _09984_ (.Y(_04301_),
    .A(net404),
    .B(_04300_));
 sg13g2_buf_2 _09985_ (.A(_00067_),
    .X(_04302_));
 sg13g2_nand2_1 _09986_ (.Y(_04303_),
    .A(_04302_),
    .B(net215));
 sg13g2_o21ai_1 _09987_ (.B1(_04303_),
    .Y(_04304_),
    .A1(net215),
    .A2(_04301_));
 sg13g2_xnor2_1 _09988_ (.Y(_04305_),
    .A(_04299_),
    .B(_04304_));
 sg13g2_nand2b_1 _09989_ (.Y(_04306_),
    .B(_04305_),
    .A_N(net37));
 sg13g2_nand2_1 _09990_ (.Y(_04307_),
    .A(_03928_),
    .B(net37));
 sg13g2_nand3_1 _09991_ (.B(_04306_),
    .C(_04307_),
    .A(net250),
    .Y(_00223_));
 sg13g2_nor2_1 _09992_ (.A(_03317_),
    .B(_03324_),
    .Y(_04308_));
 sg13g2_buf_1 _09993_ (.A(_04308_),
    .X(_04309_));
 sg13g2_buf_1 _09994_ (.A(net236),
    .X(_04310_));
 sg13g2_buf_1 _09995_ (.A(net209),
    .X(_04311_));
 sg13g2_nand2_1 _09996_ (.Y(_04312_),
    .A(net404),
    .B(_04299_));
 sg13g2_mux2_1 _09997_ (.A0(_04299_),
    .A1(_04312_),
    .S(net366),
    .X(_04313_));
 sg13g2_nand2b_1 _09998_ (.Y(_04314_),
    .B(net404),
    .A_N(net366));
 sg13g2_nand2b_1 _09999_ (.Y(_04315_),
    .B(net366),
    .A_N(net368));
 sg13g2_nand3_1 _10000_ (.B(_04314_),
    .C(_04315_),
    .A(_04312_),
    .Y(_04316_));
 sg13g2_o21ai_1 _10001_ (.B1(_04316_),
    .Y(_04317_),
    .A1(_03405_),
    .A2(_04313_));
 sg13g2_xnor2_1 _10002_ (.Y(_04318_),
    .A(_03989_),
    .B(_04317_));
 sg13g2_nand2_1 _10003_ (.Y(_04319_),
    .A(_04293_),
    .B(_04302_));
 sg13g2_xor2_1 _10004_ (.B(_04319_),
    .A(_03925_),
    .X(_04320_));
 sg13g2_nor2_1 _10005_ (.A(net173),
    .B(_04320_),
    .Y(_04321_));
 sg13g2_a21oi_1 _10006_ (.A1(net173),
    .A2(_04318_),
    .Y(_04322_),
    .B1(_04321_));
 sg13g2_nand2b_1 _10007_ (.Y(_04323_),
    .B(_04322_),
    .A_N(net40));
 sg13g2_nand2_1 _10008_ (.Y(_04324_),
    .A(_03926_),
    .B(net37));
 sg13g2_nand3_1 _10009_ (.B(_04323_),
    .C(_04324_),
    .A(net250),
    .Y(_00224_));
 sg13g2_nand3_1 _10010_ (.B(_03925_),
    .C(_04302_),
    .A(_04293_),
    .Y(_04325_));
 sg13g2_o21ai_1 _10011_ (.B1(_04300_),
    .Y(_04326_),
    .A1(_03980_),
    .A2(_04299_));
 sg13g2_nand3_1 _10012_ (.B(_04315_),
    .C(_04326_),
    .A(_04312_),
    .Y(_04327_));
 sg13g2_nand3_1 _10013_ (.B(_04309_),
    .C(_04327_),
    .A(_03989_),
    .Y(_04328_));
 sg13g2_o21ai_1 _10014_ (.B1(_04328_),
    .Y(_04329_),
    .A1(_04309_),
    .A2(_04325_));
 sg13g2_buf_1 _10015_ (.A(_04329_),
    .X(_04330_));
 sg13g2_and2_1 _10016_ (.A(net368),
    .B(net366),
    .X(_04331_));
 sg13g2_buf_1 _10017_ (.A(_04331_),
    .X(_04332_));
 sg13g2_xnor2_1 _10018_ (.Y(_04333_),
    .A(_03979_),
    .B(_04332_));
 sg13g2_buf_1 _10019_ (.A(_00068_),
    .X(_04334_));
 sg13g2_and2_1 _10020_ (.A(_04334_),
    .B(_03326_),
    .X(_04335_));
 sg13g2_a21o_1 _10021_ (.A2(_04333_),
    .A1(net173),
    .B1(_04335_),
    .X(_04336_));
 sg13g2_xnor2_1 _10022_ (.Y(_04337_),
    .A(_04330_),
    .B(_04336_));
 sg13g2_nand2b_1 _10023_ (.Y(_04338_),
    .B(_04337_),
    .A_N(net40));
 sg13g2_nand2_1 _10024_ (.Y(_04339_),
    .A(\dtop.vtop.pipeline.dz[3] ),
    .B(net37));
 sg13g2_nand3_1 _10025_ (.B(_04338_),
    .C(_04339_),
    .A(net250),
    .Y(_00225_));
 sg13g2_nand2_1 _10026_ (.Y(_04340_),
    .A(_03923_),
    .B(net37));
 sg13g2_o21ai_1 _10027_ (.B1(_04332_),
    .Y(_04341_),
    .A1(_03978_),
    .A2(_04330_));
 sg13g2_nand2_1 _10028_ (.Y(_04342_),
    .A(_03978_),
    .B(_04330_));
 sg13g2_nand2_1 _10029_ (.Y(_04343_),
    .A(_04341_),
    .B(_04342_));
 sg13g2_a22oi_1 _10030_ (.Y(_04344_),
    .B1(_04343_),
    .B2(net209),
    .A2(_04335_),
    .A1(_04330_));
 sg13g2_buf_1 _10031_ (.A(_04344_),
    .X(_04345_));
 sg13g2_nand2_1 _10032_ (.Y(_04346_),
    .A(_03937_),
    .B(net215));
 sg13g2_o21ai_1 _10033_ (.B1(_04346_),
    .Y(_04347_),
    .A1(_03976_),
    .A2(net215));
 sg13g2_xor2_1 _10034_ (.B(_04347_),
    .A(_04345_),
    .X(_04348_));
 sg13g2_nand2b_1 _10035_ (.Y(_04349_),
    .B(_04348_),
    .A_N(net40));
 sg13g2_nand3_1 _10036_ (.B(_04340_),
    .C(_04349_),
    .A(net250),
    .Y(_00226_));
 sg13g2_nand2_1 _10037_ (.Y(_04350_),
    .A(\dtop.vtop.pipeline.dz[5] ),
    .B(net37));
 sg13g2_buf_1 _10038_ (.A(_00070_),
    .X(_04351_));
 sg13g2_nor2b_1 _10039_ (.A(_04345_),
    .B_N(_03937_),
    .Y(_04352_));
 sg13g2_xnor2_1 _10040_ (.Y(_04353_),
    .A(_04351_),
    .B(_04352_));
 sg13g2_nand2b_1 _10041_ (.Y(_04354_),
    .B(_04353_),
    .A_N(net40));
 sg13g2_nand3_1 _10042_ (.B(_04350_),
    .C(_04354_),
    .A(net250),
    .Y(_00227_));
 sg13g2_nand3_1 _10043_ (.B(_00069_),
    .C(_04310_),
    .A(_00021_),
    .Y(_04355_));
 sg13g2_nand3_1 _10044_ (.B(_04351_),
    .C(_03326_),
    .A(_03937_),
    .Y(_04356_));
 sg13g2_a21oi_2 _10045_ (.B1(_04345_),
    .Y(_04357_),
    .A2(_04356_),
    .A1(_04355_));
 sg13g2_nand2_1 _10046_ (.Y(_04358_),
    .A(_04002_),
    .B(_04310_));
 sg13g2_o21ai_1 _10047_ (.B1(_04358_),
    .Y(_04359_),
    .A1(_03946_),
    .A2(net173));
 sg13g2_xnor2_1 _10048_ (.Y(_04360_),
    .A(_04357_),
    .B(_04359_));
 sg13g2_nand2b_1 _10049_ (.Y(_04361_),
    .B(_04360_),
    .A_N(net40));
 sg13g2_nand2_1 _10050_ (.Y(_04362_),
    .A(\dtop.vtop.pipeline.dz[6] ),
    .B(_04289_));
 sg13g2_nand3_1 _10051_ (.B(_04361_),
    .C(_04362_),
    .A(net250),
    .Y(_00228_));
 sg13g2_nand2_1 _10052_ (.Y(_04363_),
    .A(_03919_),
    .B(_04289_));
 sg13g2_nand2_1 _10053_ (.Y(_04364_),
    .A(_03945_),
    .B(_04357_));
 sg13g2_xnor2_1 _10054_ (.Y(_04365_),
    .A(_03949_),
    .B(_04364_));
 sg13g2_nand2_1 _10055_ (.Y(_04366_),
    .A(_04002_),
    .B(_04357_));
 sg13g2_xor2_1 _10056_ (.B(_04366_),
    .A(net403),
    .X(_04367_));
 sg13g2_nand2_1 _10057_ (.Y(_04368_),
    .A(_04311_),
    .B(_04367_));
 sg13g2_o21ai_1 _10058_ (.B1(_04368_),
    .Y(_04369_),
    .A1(_04311_),
    .A2(_04365_));
 sg13g2_nand2b_1 _10059_ (.Y(_04370_),
    .B(_04369_),
    .A_N(_04288_));
 sg13g2_nand3_1 _10060_ (.B(_04363_),
    .C(_04370_),
    .A(net250),
    .Y(_00229_));
 sg13g2_buf_1 _10061_ (.A(\dtop.vtop.pipeline.dz[8] ),
    .X(_04371_));
 sg13g2_nand2_1 _10062_ (.Y(_04372_),
    .A(_04371_),
    .B(net37));
 sg13g2_nand3_1 _10063_ (.B(net403),
    .C(net209),
    .A(_04002_),
    .Y(_04373_));
 sg13g2_nand3_1 _10064_ (.B(_03945_),
    .C(net215),
    .A(_03949_),
    .Y(_04374_));
 sg13g2_nand2_1 _10065_ (.Y(_04375_),
    .A(_04373_),
    .B(_04374_));
 sg13g2_nand2_1 _10066_ (.Y(_04376_),
    .A(_04357_),
    .B(_04375_));
 sg13g2_mux2_1 _10067_ (.A0(_04371_),
    .A1(\dtop.vtop.pipeline.neg_t[8] ),
    .S(net209),
    .X(_04377_));
 sg13g2_xnor2_1 _10068_ (.Y(_04378_),
    .A(_04376_),
    .B(_04377_));
 sg13g2_nand2b_1 _10069_ (.Y(_04379_),
    .B(_04378_),
    .A_N(net40));
 sg13g2_nand3_1 _10070_ (.B(_04372_),
    .C(_04379_),
    .A(net250),
    .Y(_00230_));
 sg13g2_buf_1 _10071_ (.A(net252),
    .X(_04380_));
 sg13g2_nor2_1 _10072_ (.A(_00089_),
    .B(net215),
    .Y(_04381_));
 sg13g2_buf_1 _10073_ (.A(_04381_),
    .X(_04382_));
 sg13g2_nor2_1 _10074_ (.A(\dtop.vtop.pipeline.neg_t[0] ),
    .B(net140),
    .Y(_04383_));
 sg13g2_nand2_1 _10075_ (.Y(_04384_),
    .A(_03970_),
    .B(net209));
 sg13g2_buf_1 _10076_ (.A(_04384_),
    .X(_04385_));
 sg13g2_nor2_1 _10077_ (.A(_04295_),
    .B(_04385_),
    .Y(_04386_));
 sg13g2_nor3_1 _10078_ (.A(net235),
    .B(_04383_),
    .C(_04386_),
    .Y(_00231_));
 sg13g2_nor2_1 _10079_ (.A(\dtop.vtop.pipeline.neg_t[1] ),
    .B(net140),
    .Y(_04387_));
 sg13g2_nor2_1 _10080_ (.A(_04305_),
    .B(net139),
    .Y(_04388_));
 sg13g2_nor3_1 _10081_ (.A(net235),
    .B(_04387_),
    .C(_04388_),
    .Y(_00232_));
 sg13g2_nor2_1 _10082_ (.A(\dtop.vtop.pipeline.neg_t[2] ),
    .B(net140),
    .Y(_04389_));
 sg13g2_nor2_1 _10083_ (.A(_04322_),
    .B(net139),
    .Y(_04390_));
 sg13g2_nor3_1 _10084_ (.A(net235),
    .B(_04389_),
    .C(_04390_),
    .Y(_00233_));
 sg13g2_nor2_1 _10085_ (.A(\dtop.vtop.pipeline.neg_t[3] ),
    .B(_04382_),
    .Y(_04391_));
 sg13g2_nor2_1 _10086_ (.A(_04337_),
    .B(_04385_),
    .Y(_04392_));
 sg13g2_nor3_1 _10087_ (.A(net235),
    .B(_04391_),
    .C(_04392_),
    .Y(_00234_));
 sg13g2_nand2_1 _10088_ (.Y(_04393_),
    .A(_04348_),
    .B(net140));
 sg13g2_nand2_1 _10089_ (.Y(_04394_),
    .A(\dtop.vtop.pipeline.neg_t[4] ),
    .B(net139));
 sg13g2_buf_1 _10090_ (.A(net252),
    .X(_04395_));
 sg13g2_a21oi_1 _10091_ (.A1(_04393_),
    .A2(_04394_),
    .Y(_00235_),
    .B1(net234));
 sg13g2_nand2_1 _10092_ (.Y(_04396_),
    .A(\dtop.vtop.pipeline.neg_t[5] ),
    .B(net139));
 sg13g2_nor2_1 _10093_ (.A(_03976_),
    .B(_04345_),
    .Y(_04397_));
 sg13g2_xnor2_1 _10094_ (.Y(_04398_),
    .A(_00069_),
    .B(_04397_));
 sg13g2_nand2_1 _10095_ (.Y(_04399_),
    .A(net140),
    .B(_04398_));
 sg13g2_a21oi_1 _10096_ (.A1(_04396_),
    .A2(_04399_),
    .Y(_00236_),
    .B1(_04395_));
 sg13g2_nor2_1 _10097_ (.A(\dtop.vtop.pipeline.neg_t[6] ),
    .B(net140),
    .Y(_04400_));
 sg13g2_nor2_1 _10098_ (.A(_04360_),
    .B(net139),
    .Y(_04401_));
 sg13g2_nor3_1 _10099_ (.A(net235),
    .B(_04400_),
    .C(_04401_),
    .Y(_00237_));
 sg13g2_nand2_1 _10100_ (.Y(_04402_),
    .A(_04369_),
    .B(net140));
 sg13g2_nand2_1 _10101_ (.Y(_04403_),
    .A(\dtop.vtop.pipeline.neg_t[7] ),
    .B(net139));
 sg13g2_a21oi_1 _10102_ (.A1(_04402_),
    .A2(_04403_),
    .Y(_00238_),
    .B1(_04395_));
 sg13g2_buf_1 _10103_ (.A(net252),
    .X(_04404_));
 sg13g2_nor2_1 _10104_ (.A(_04376_),
    .B(net139),
    .Y(_04405_));
 sg13g2_xnor2_1 _10105_ (.Y(_04406_),
    .A(\dtop.vtop.pipeline.neg_t[8] ),
    .B(_04405_));
 sg13g2_nor2_1 _10106_ (.A(net233),
    .B(_04406_),
    .Y(_00239_));
 sg13g2_nand2_1 _10107_ (.Y(_04407_),
    .A(\dtop.vtop.pipeline.neg_t[9] ),
    .B(net139));
 sg13g2_nor2_1 _10108_ (.A(_04376_),
    .B(_04377_),
    .Y(_04408_));
 sg13g2_xnor2_1 _10109_ (.Y(_04409_),
    .A(_04022_),
    .B(_04408_));
 sg13g2_nand2_1 _10110_ (.Y(_04410_),
    .A(net140),
    .B(_04409_));
 sg13g2_a21oi_1 _10111_ (.A1(_04407_),
    .A2(_04410_),
    .Y(_00240_),
    .B1(net235));
 sg13g2_nand2_1 _10112_ (.Y(_04411_),
    .A(\dtop.vtop.pipeline.nstep_counter[0] ),
    .B(net112));
 sg13g2_nand2_1 _10113_ (.Y(_04412_),
    .A(\dtop.vtop.pipeline.next_nstep_counter[0] ),
    .B(_03364_));
 sg13g2_nand3_1 _10114_ (.B(_04411_),
    .C(_04412_),
    .A(net267),
    .Y(_00241_));
 sg13g2_nor3_1 _10115_ (.A(\dtop.vtop.pipeline.nstep_counter[0] ),
    .B(\dtop.vtop.pipeline.nstep_counter[1] ),
    .C(_03329_),
    .Y(_04413_));
 sg13g2_o21ai_1 _10116_ (.B1(\dtop.vtop.pipeline.nstep_counter[1] ),
    .Y(_04414_),
    .A1(\dtop.vtop.pipeline.nstep_counter[0] ),
    .A2(net112));
 sg13g2_nor2b_1 _10117_ (.A(_04413_),
    .B_N(_04414_),
    .Y(_04415_));
 sg13g2_nand2_1 _10118_ (.Y(_00242_),
    .A(_04286_),
    .B(_04415_));
 sg13g2_nor2b_1 _10119_ (.A(\dtop.vtop.pipeline.nstep_counter[2] ),
    .B_N(_04413_),
    .Y(_04416_));
 sg13g2_nor2b_1 _10120_ (.A(_04413_),
    .B_N(\dtop.vtop.pipeline.nstep_counter[2] ),
    .Y(_04417_));
 sg13g2_or3_1 _10121_ (.A(net252),
    .B(_04416_),
    .C(_04417_),
    .X(_00243_));
 sg13g2_nand2b_1 _10122_ (.Y(_04418_),
    .B(_04416_),
    .A_N(\dtop.vtop.pipeline.nstep_counter[3] ));
 sg13g2_nand2b_1 _10123_ (.Y(_04419_),
    .B(\dtop.vtop.pipeline.nstep_counter[3] ),
    .A_N(_04416_));
 sg13g2_nand3_1 _10124_ (.B(_04418_),
    .C(_04419_),
    .A(net267),
    .Y(_00244_));
 sg13g2_a21o_1 _10125_ (.A2(_04418_),
    .A1(\dtop.vtop.pipeline.nstep_counter[4] ),
    .B1(_04380_),
    .X(_00245_));
 sg13g2_xor2_1 _10126_ (.B(net367),
    .A(net351),
    .X(_04420_));
 sg13g2_nor4_1 _10127_ (.A(net399),
    .B(_03493_),
    .C(_03273_),
    .D(_04420_),
    .Y(_04421_));
 sg13g2_nand3_1 _10128_ (.B(net364),
    .C(_02850_),
    .A(net372),
    .Y(_04422_));
 sg13g2_o21ai_1 _10129_ (.B1(_04422_),
    .Y(_04423_),
    .A1(net372),
    .A2(_03430_));
 sg13g2_a22oi_1 _10130_ (.Y(_04424_),
    .B1(_04423_),
    .B2(net399),
    .A2(_03273_),
    .A1(net367));
 sg13g2_nor2_1 _10131_ (.A(_00031_),
    .B(_04424_),
    .Y(_04425_));
 sg13g2_nor4_2 _10132_ (.A(\dtop.vtop.pipeline.nstep_counter[4] ),
    .B(_04418_),
    .C(_04421_),
    .Y(_04426_),
    .D(_04425_));
 sg13g2_xnor2_1 _10133_ (.Y(_04427_),
    .A(net367),
    .B(_04426_));
 sg13g2_nor2_1 _10134_ (.A(_04404_),
    .B(_04427_),
    .Y(_00246_));
 sg13g2_nand2_1 _10135_ (.Y(_04428_),
    .A(net367),
    .B(_04426_));
 sg13g2_xnor2_1 _10136_ (.Y(_04429_),
    .A(_03461_),
    .B(_04428_));
 sg13g2_nor2_1 _10137_ (.A(_04404_),
    .B(_04429_),
    .Y(_00247_));
 sg13g2_nor2_1 _10138_ (.A(_02250_),
    .B(_02264_),
    .Y(_04430_));
 sg13g2_a21oi_1 _10139_ (.A1(_02250_),
    .A2(_03269_),
    .Y(_04431_),
    .B1(_04430_));
 sg13g2_nor3_1 _10140_ (.A(net252),
    .B(net84),
    .C(_04431_),
    .Y(_00298_));
 sg13g2_nand2_1 _10141_ (.Y(_04432_),
    .A(_03269_),
    .B(_03362_));
 sg13g2_o21ai_1 _10142_ (.B1(_02250_),
    .Y(_04433_),
    .A1(_03269_),
    .A2(_03362_));
 sg13g2_a221oi_1 _10143_ (.B2(_02846_),
    .C1(_04380_),
    .B1(_04433_),
    .A1(_02847_),
    .Y(_00299_),
    .A2(_04432_));
 sg13g2_o21ai_1 _10144_ (.B1(\dtop.vtop.pipeline.zg_valid ),
    .Y(_04434_),
    .A1(net209),
    .A2(_03958_));
 sg13g2_buf_1 _10145_ (.A(_04434_),
    .X(_04435_));
 sg13g2_buf_1 _10146_ (.A(_04435_),
    .X(_04436_));
 sg13g2_nand2_1 _10147_ (.Y(_04437_),
    .A(_03927_),
    .B(_04291_));
 sg13g2_nand2_1 _10148_ (.Y(_04438_),
    .A(net173),
    .B(_04437_));
 sg13g2_o21ai_1 _10149_ (.B1(_04438_),
    .Y(_04439_),
    .A1(_03982_),
    .A2(net173));
 sg13g2_nor2_1 _10150_ (.A(_04436_),
    .B(_04439_),
    .Y(_04440_));
 sg13g2_xnor2_1 _10151_ (.Y(_04441_),
    .A(\dtop.vtop.pipeline.z[0] ),
    .B(_04440_));
 sg13g2_nor2_1 _10152_ (.A(net233),
    .B(_04441_),
    .Y(_00300_));
 sg13g2_mux2_1 _10153_ (.A0(_04371_),
    .A1(_03946_),
    .S(net366),
    .X(_04442_));
 sg13g2_nand2_1 _10154_ (.Y(_04443_),
    .A(net368),
    .B(_04442_));
 sg13g2_o21ai_1 _10155_ (.B1(_04443_),
    .Y(_04444_),
    .A1(_03949_),
    .A2(_04315_));
 sg13g2_nor2_1 _10156_ (.A(_03326_),
    .B(_04444_),
    .Y(_04445_));
 sg13g2_a21oi_2 _10157_ (.B1(_04445_),
    .Y(_04446_),
    .A2(_03326_),
    .A1(_04022_));
 sg13g2_inv_1 _10158_ (.Y(_04447_),
    .A(_03282_));
 sg13g2_mux4_1 _10159_ (.S0(net407),
    .A0(_03954_),
    .A1(_03949_),
    .A2(_03945_),
    .A3(_04351_),
    .S1(net405),
    .X(_04448_));
 sg13g2_mux2_1 _10160_ (.A0(_00027_),
    .A1(_04448_),
    .S(net236),
    .X(_04449_));
 sg13g2_buf_1 _10161_ (.A(_04449_),
    .X(_04450_));
 sg13g2_inv_1 _10162_ (.Y(_04451_),
    .A(\dtop.vtop.pipeline.z[4] ));
 sg13g2_mux4_1 _10163_ (.S0(net405),
    .A0(_03937_),
    .A1(_03925_),
    .A2(_04334_),
    .A3(_04302_),
    .S1(net407),
    .X(_04452_));
 sg13g2_mux2_1 _10164_ (.A0(_00021_),
    .A1(_04452_),
    .S(net236),
    .X(_04453_));
 sg13g2_mux4_1 _10165_ (.S0(net405),
    .A0(_04334_),
    .A1(_04302_),
    .A2(_03925_),
    .A3(_04293_),
    .S1(net407),
    .X(_04454_));
 sg13g2_mux2_1 _10166_ (.A0(_03978_),
    .A1(_04454_),
    .S(net236),
    .X(_04455_));
 sg13g2_inv_1 _10167_ (.Y(_04456_),
    .A(_04455_));
 sg13g2_nand2_1 _10168_ (.Y(_04457_),
    .A(\dtop.vtop.pipeline.z[3] ),
    .B(_04456_));
 sg13g2_inv_1 _10169_ (.Y(_04458_),
    .A(\dtop.vtop.pipeline.z[2] ));
 sg13g2_nand2_1 _10170_ (.Y(_04459_),
    .A(net405),
    .B(_03927_));
 sg13g2_o21ai_1 _10171_ (.B1(_04459_),
    .Y(_04460_),
    .A1(net405),
    .A2(_03925_));
 sg13g2_o21ai_1 _10172_ (.B1(net407),
    .Y(_04461_),
    .A1(_03410_),
    .A2(_04302_));
 sg13g2_o21ai_1 _10173_ (.B1(_04461_),
    .Y(_04462_),
    .A1(net407),
    .A2(_04460_));
 sg13g2_mux2_1 _10174_ (.A0(_03989_),
    .A1(_04462_),
    .S(net236),
    .X(_04463_));
 sg13g2_nor2_1 _10175_ (.A(_04458_),
    .B(_04463_),
    .Y(_04464_));
 sg13g2_or4_1 _10176_ (.A(_04302_),
    .B(_03317_),
    .C(_03324_),
    .D(_04437_),
    .X(_04465_));
 sg13g2_nor2_1 _10177_ (.A(_03981_),
    .B(net404),
    .Y(_04466_));
 sg13g2_o21ai_1 _10178_ (.B1(_04466_),
    .Y(_04467_),
    .A1(_03317_),
    .A2(_03324_));
 sg13g2_inv_1 _10179_ (.Y(_04468_),
    .A(\dtop.vtop.pipeline.z[0] ));
 sg13g2_a21o_1 _10180_ (.A2(_04467_),
    .A1(_04465_),
    .B1(_04468_),
    .X(_04469_));
 sg13g2_inv_1 _10181_ (.Y(_04470_),
    .A(\dtop.vtop.pipeline.z[1] ));
 sg13g2_mux2_1 _10182_ (.A0(_04302_),
    .A1(_04293_),
    .S(net407),
    .X(_04471_));
 sg13g2_nor2_1 _10183_ (.A(net405),
    .B(_04471_),
    .Y(_04472_));
 sg13g2_or3_1 _10184_ (.A(_03317_),
    .B(_03324_),
    .C(_04472_),
    .X(_04473_));
 sg13g2_o21ai_1 _10185_ (.B1(net404),
    .Y(_04474_),
    .A1(_03317_),
    .A2(_03324_));
 sg13g2_nor2_1 _10186_ (.A(_03981_),
    .B(_04468_),
    .Y(_04475_));
 sg13g2_nor4_1 _10187_ (.A(_04468_),
    .B(_03317_),
    .C(_03324_),
    .D(_04437_),
    .Y(_04476_));
 sg13g2_a221oi_1 _10188_ (.B2(_03326_),
    .C1(_04476_),
    .B1(_04475_),
    .A1(_04473_),
    .Y(_04477_),
    .A2(_04474_));
 sg13g2_a221oi_1 _10189_ (.B2(_04470_),
    .C1(_04477_),
    .B1(_04469_),
    .A1(_04458_),
    .Y(_04478_),
    .A2(_04463_));
 sg13g2_nand2b_1 _10190_ (.Y(_04479_),
    .B(_04455_),
    .A_N(\dtop.vtop.pipeline.z[3] ));
 sg13g2_o21ai_1 _10191_ (.B1(_04479_),
    .Y(_04480_),
    .A1(_04464_),
    .A2(_04478_));
 sg13g2_a22oi_1 _10192_ (.Y(_04481_),
    .B1(_04457_),
    .B2(_04480_),
    .A2(_04453_),
    .A1(_04451_));
 sg13g2_mux4_1 _10193_ (.S0(net405),
    .A0(_04351_),
    .A1(_04334_),
    .A2(_03937_),
    .A3(_03925_),
    .S1(net407),
    .X(_04482_));
 sg13g2_mux2_1 _10194_ (.A0(_00069_),
    .A1(_04482_),
    .S(net236),
    .X(_04483_));
 sg13g2_inv_1 _10195_ (.Y(_04484_),
    .A(_04453_));
 sg13g2_nand2_1 _10196_ (.Y(_04485_),
    .A(\dtop.vtop.pipeline.z[4] ),
    .B(_04484_));
 sg13g2_nand2_1 _10197_ (.Y(_04486_),
    .A(_04483_),
    .B(_04485_));
 sg13g2_o21ai_1 _10198_ (.B1(\dtop.vtop.pipeline.z[5] ),
    .Y(_04487_),
    .A1(_04481_),
    .A2(_04486_));
 sg13g2_buf_1 _10199_ (.A(_04487_),
    .X(_04488_));
 sg13g2_inv_1 _10200_ (.Y(_04489_),
    .A(_04485_));
 sg13g2_inv_1 _10201_ (.Y(_04490_),
    .A(_04483_));
 sg13g2_o21ai_1 _10202_ (.B1(_04490_),
    .Y(_04491_),
    .A1(_04481_),
    .A2(_04489_));
 sg13g2_buf_1 _10203_ (.A(_04491_),
    .X(_04492_));
 sg13g2_mux4_1 _10204_ (.S0(net368),
    .A0(_03949_),
    .A1(_03945_),
    .A2(_04351_),
    .A3(_03937_),
    .S1(net366),
    .X(_04493_));
 sg13g2_mux2_1 _10205_ (.A0(net403),
    .A1(_04493_),
    .S(net236),
    .X(_04494_));
 sg13g2_mux4_1 _10206_ (.S0(net366),
    .A0(_03945_),
    .A1(_03937_),
    .A2(_04351_),
    .A3(_04334_),
    .S1(net368),
    .X(_04495_));
 sg13g2_mux2_1 _10207_ (.A0(_04002_),
    .A1(_04495_),
    .S(net236),
    .X(_04496_));
 sg13g2_buf_1 _10208_ (.A(_04496_),
    .X(_04497_));
 sg13g2_or2_1 _10209_ (.X(_04498_),
    .B(_04497_),
    .A(_04494_));
 sg13g2_or2_1 _10210_ (.X(_04499_),
    .B(_04497_),
    .A(_03287_));
 sg13g2_and2_1 _10211_ (.A(_04447_),
    .B(_04450_),
    .X(_04500_));
 sg13g2_buf_1 _10212_ (.A(_04500_),
    .X(_04501_));
 sg13g2_a221oi_1 _10213_ (.B2(_04499_),
    .C1(_04501_),
    .B1(_04498_),
    .A1(_04488_),
    .Y(_04502_),
    .A2(_04492_));
 sg13g2_inv_1 _10214_ (.Y(_04503_),
    .A(_04494_));
 sg13g2_nand2_1 _10215_ (.Y(_04504_),
    .A(_03288_),
    .B(_04503_));
 sg13g2_nand2_1 _10216_ (.Y(_04505_),
    .A(_03288_),
    .B(_03285_));
 sg13g2_a221oi_1 _10217_ (.B2(_04505_),
    .C1(_04501_),
    .B1(_04504_),
    .A1(_04488_),
    .Y(_04506_),
    .A2(_04492_));
 sg13g2_inv_1 _10218_ (.Y(_04507_),
    .A(_03288_));
 sg13g2_nor3_1 _10219_ (.A(_04507_),
    .B(_04501_),
    .C(_04498_),
    .Y(_04508_));
 sg13g2_nand2_1 _10220_ (.Y(_04509_),
    .A(_03285_),
    .B(_04503_));
 sg13g2_or2_1 _10221_ (.X(_04510_),
    .B(_04505_),
    .A(_04497_));
 sg13g2_a21oi_1 _10222_ (.A1(_04509_),
    .A2(_04510_),
    .Y(_04511_),
    .B1(_04501_));
 sg13g2_nor4_2 _10223_ (.A(_04502_),
    .B(_04506_),
    .C(_04508_),
    .Y(_04512_),
    .D(_04511_));
 sg13g2_o21ai_1 _10224_ (.B1(_04512_),
    .Y(_04513_),
    .A1(_04447_),
    .A2(_04450_));
 sg13g2_buf_1 _10225_ (.A(_04513_),
    .X(_04514_));
 sg13g2_and2_1 _10226_ (.A(_04446_),
    .B(_04514_),
    .X(_04515_));
 sg13g2_buf_1 _10227_ (.A(_04515_),
    .X(_04516_));
 sg13g2_nor2_2 _10228_ (.A(_04447_),
    .B(_04450_),
    .Y(_04517_));
 sg13g2_nor2_1 _10229_ (.A(_04446_),
    .B(_04517_),
    .Y(_04518_));
 sg13g2_a21oi_1 _10230_ (.A1(_04512_),
    .A2(_04518_),
    .Y(_04519_),
    .B1(_03295_));
 sg13g2_nor2_1 _10231_ (.A(_04516_),
    .B(_04519_),
    .Y(_04520_));
 sg13g2_nor2_1 _10232_ (.A(net368),
    .B(_03954_),
    .Y(_04521_));
 sg13g2_a21oi_1 _10233_ (.A1(net368),
    .A2(_03950_),
    .Y(_04522_),
    .B1(_04521_));
 sg13g2_nor2b_1 _10234_ (.A(_04522_),
    .B_N(net366),
    .Y(_04523_));
 sg13g2_buf_1 _10235_ (.A(_04523_),
    .X(_04524_));
 sg13g2_nor2_1 _10236_ (.A(net215),
    .B(_04524_),
    .Y(_04525_));
 sg13g2_xnor2_1 _10237_ (.Y(_04526_),
    .A(_04520_),
    .B(_04525_));
 sg13g2_nor2_1 _10238_ (.A(net36),
    .B(_04526_),
    .Y(_04527_));
 sg13g2_xnor2_1 _10239_ (.Y(_04528_),
    .A(net409),
    .B(_04527_));
 sg13g2_nor2_1 _10240_ (.A(net233),
    .B(_04528_),
    .Y(_00301_));
 sg13g2_nand2_1 _10241_ (.Y(_04529_),
    .A(_04371_),
    .B(_04332_));
 sg13g2_a21oi_1 _10242_ (.A1(net173),
    .A2(_04529_),
    .Y(_04530_),
    .B1(net409));
 sg13g2_and2_1 _10243_ (.A(_04371_),
    .B(_04332_),
    .X(_04531_));
 sg13g2_buf_1 _10244_ (.A(_04531_),
    .X(_04532_));
 sg13g2_or2_1 _10245_ (.X(_04533_),
    .B(_04524_),
    .A(net409));
 sg13g2_nor3_1 _10246_ (.A(_04446_),
    .B(_04517_),
    .C(_04524_),
    .Y(_04534_));
 sg13g2_nor2_1 _10247_ (.A(_03294_),
    .B(_04524_),
    .Y(_04535_));
 sg13g2_nor2b_1 _10248_ (.A(_04517_),
    .B_N(_04535_),
    .Y(_04536_));
 sg13g2_o21ai_1 _10249_ (.B1(_04512_),
    .Y(_04537_),
    .A1(_04534_),
    .A2(_04536_));
 sg13g2_nor3_1 _10250_ (.A(net409),
    .B(_04446_),
    .C(_04517_),
    .Y(_04538_));
 sg13g2_nor2_1 _10251_ (.A(net409),
    .B(_03294_),
    .Y(_04539_));
 sg13g2_nor2b_1 _10252_ (.A(_04517_),
    .B_N(_04539_),
    .Y(_04540_));
 sg13g2_o21ai_1 _10253_ (.B1(_04512_),
    .Y(_04541_),
    .A1(_04538_),
    .A2(_04540_));
 sg13g2_inv_1 _10254_ (.Y(_04542_),
    .A(_04446_));
 sg13g2_o21ai_1 _10255_ (.B1(_04542_),
    .Y(_04543_),
    .A1(_04535_),
    .A2(_04539_));
 sg13g2_nand4_1 _10256_ (.B(_04537_),
    .C(_04541_),
    .A(_04533_),
    .Y(_04544_),
    .D(_04543_));
 sg13g2_o21ai_1 _10257_ (.B1(net409),
    .Y(_04545_),
    .A1(_04516_),
    .A2(_04519_));
 sg13g2_nand3b_1 _10258_ (.B(_04532_),
    .C(_04545_),
    .Y(_04546_),
    .A_N(_04524_));
 sg13g2_o21ai_1 _10259_ (.B1(_04546_),
    .Y(_04547_),
    .A1(_04532_),
    .A2(_04544_));
 sg13g2_a22oi_1 _10260_ (.Y(_04548_),
    .B1(_04547_),
    .B2(net173),
    .A2(_04530_),
    .A1(_04520_));
 sg13g2_o21ai_1 _10261_ (.B1(_03276_),
    .Y(_04549_),
    .A1(net36),
    .A2(_04548_));
 sg13g2_or3_1 _10262_ (.A(_03276_),
    .B(net36),
    .C(_04548_),
    .X(_04550_));
 sg13g2_a21oi_1 _10263_ (.A1(_04549_),
    .A2(_04550_),
    .Y(_00302_),
    .B1(net235));
 sg13g2_nand2_1 _10264_ (.Y(_04551_),
    .A(_03294_),
    .B(_04514_));
 sg13g2_nor2_1 _10265_ (.A(_03294_),
    .B(_04514_),
    .Y(_04552_));
 sg13g2_a21oi_1 _10266_ (.A1(_04022_),
    .A2(_04551_),
    .Y(_04553_),
    .B1(_04552_));
 sg13g2_or4_1 _10267_ (.A(_03276_),
    .B(net409),
    .C(net209),
    .D(_04553_),
    .X(_04554_));
 sg13g2_buf_1 _10268_ (.A(_04554_),
    .X(_04555_));
 sg13g2_nor2_1 _10269_ (.A(_03276_),
    .B(_04532_),
    .Y(_04556_));
 sg13g2_nand2_1 _10270_ (.Y(_04557_),
    .A(_03276_),
    .B(_04532_));
 sg13g2_o21ai_1 _10271_ (.B1(_04557_),
    .Y(_04558_),
    .A1(_04544_),
    .A2(_04556_));
 sg13g2_nand2_1 _10272_ (.Y(_04559_),
    .A(net209),
    .B(_04558_));
 sg13g2_a21oi_1 _10273_ (.A1(_04555_),
    .A2(_04559_),
    .Y(_04560_),
    .B1(net36));
 sg13g2_xnor2_1 _10274_ (.Y(_04561_),
    .A(_03307_),
    .B(_04560_));
 sg13g2_nor2_1 _10275_ (.A(net233),
    .B(_04561_),
    .Y(_00303_));
 sg13g2_mux2_1 _10276_ (.A0(_04555_),
    .A1(_04559_),
    .S(_03307_),
    .X(_04562_));
 sg13g2_nor2_1 _10277_ (.A(net36),
    .B(_04562_),
    .Y(_04563_));
 sg13g2_xnor2_1 _10278_ (.Y(_04564_),
    .A(_03310_),
    .B(_04563_));
 sg13g2_nor2_1 _10279_ (.A(net233),
    .B(_04564_),
    .Y(_00304_));
 sg13g2_inv_1 _10280_ (.Y(_04565_),
    .A(_03310_));
 sg13g2_nor3_1 _10281_ (.A(_03308_),
    .B(_04565_),
    .C(_04559_),
    .Y(_04566_));
 sg13g2_nor3_1 _10282_ (.A(_03307_),
    .B(_03310_),
    .C(_04555_),
    .Y(_04567_));
 sg13g2_inv_1 _10283_ (.Y(_04568_),
    .A(_04435_));
 sg13g2_o21ai_1 _10284_ (.B1(_04568_),
    .Y(_04569_),
    .A1(_04566_),
    .A2(_04567_));
 sg13g2_xnor2_1 _10285_ (.Y(_04570_),
    .A(_03318_),
    .B(_04569_));
 sg13g2_nor2_1 _10286_ (.A(net233),
    .B(_04570_),
    .Y(_00305_));
 sg13g2_a21oi_1 _10287_ (.A1(_04465_),
    .A2(_04467_),
    .Y(_04571_),
    .B1(_04468_));
 sg13g2_nor3_1 _10288_ (.A(_04435_),
    .B(_04571_),
    .C(_04477_),
    .Y(_04572_));
 sg13g2_xnor2_1 _10289_ (.Y(_04573_),
    .A(\dtop.vtop.pipeline.z[1] ),
    .B(_04572_));
 sg13g2_nor2_1 _10290_ (.A(net233),
    .B(_04573_),
    .Y(_00306_));
 sg13g2_a21oi_1 _10291_ (.A1(_04470_),
    .A2(_04469_),
    .Y(_04574_),
    .B1(_04477_));
 sg13g2_xor2_1 _10292_ (.B(_04574_),
    .A(_04463_),
    .X(_04575_));
 sg13g2_nor2_1 _10293_ (.A(_04436_),
    .B(_04575_),
    .Y(_04576_));
 sg13g2_xnor2_1 _10294_ (.Y(_04577_),
    .A(\dtop.vtop.pipeline.z[2] ),
    .B(_04576_));
 sg13g2_nor2_1 _10295_ (.A(net233),
    .B(_04577_),
    .Y(_00307_));
 sg13g2_nor2_1 _10296_ (.A(_04464_),
    .B(_04478_),
    .Y(_04578_));
 sg13g2_xnor2_1 _10297_ (.Y(_04579_),
    .A(_04456_),
    .B(_04578_));
 sg13g2_nand2_1 _10298_ (.Y(_04580_),
    .A(_04568_),
    .B(_04579_));
 sg13g2_xor2_1 _10299_ (.B(_04580_),
    .A(\dtop.vtop.pipeline.z[3] ),
    .X(_04581_));
 sg13g2_nor2_1 _10300_ (.A(net234),
    .B(_04581_),
    .Y(_00308_));
 sg13g2_nand2_1 _10301_ (.Y(_04582_),
    .A(_04457_),
    .B(_04480_));
 sg13g2_xnor2_1 _10302_ (.Y(_04583_),
    .A(_04484_),
    .B(_04582_));
 sg13g2_nor2_1 _10303_ (.A(net36),
    .B(_04583_),
    .Y(_04584_));
 sg13g2_xnor2_1 _10304_ (.Y(_04585_),
    .A(\dtop.vtop.pipeline.z[4] ),
    .B(_04584_));
 sg13g2_nor2_1 _10305_ (.A(net234),
    .B(_04585_),
    .Y(_00309_));
 sg13g2_or2_1 _10306_ (.X(_04586_),
    .B(_04486_),
    .A(_04481_));
 sg13g2_and3_1 _10307_ (.X(_04587_),
    .A(_04568_),
    .B(_04586_),
    .C(_04492_));
 sg13g2_xnor2_1 _10308_ (.Y(_04588_),
    .A(\dtop.vtop.pipeline.z[5] ),
    .B(_04587_));
 sg13g2_nor2_1 _10309_ (.A(net234),
    .B(_04588_),
    .Y(_00310_));
 sg13g2_and3_1 _10310_ (.X(_04589_),
    .A(_04488_),
    .B(_04492_),
    .C(_04497_));
 sg13g2_a21oi_1 _10311_ (.A1(_04488_),
    .A2(_04492_),
    .Y(_04590_),
    .B1(_04497_));
 sg13g2_nor3_1 _10312_ (.A(_04435_),
    .B(_04589_),
    .C(_04590_),
    .Y(_04591_));
 sg13g2_xnor2_1 _10313_ (.Y(_04592_),
    .A(_03288_),
    .B(_04591_));
 sg13g2_nor2_1 _10314_ (.A(net234),
    .B(_04592_),
    .Y(_00311_));
 sg13g2_nor2_1 _10315_ (.A(_04507_),
    .B(_04589_),
    .Y(_04593_));
 sg13g2_nor2_1 _10316_ (.A(_04593_),
    .B(_04590_),
    .Y(_04594_));
 sg13g2_xnor2_1 _10317_ (.Y(_04595_),
    .A(_04494_),
    .B(_04594_));
 sg13g2_nor2_1 _10318_ (.A(net36),
    .B(_04595_),
    .Y(_04596_));
 sg13g2_xnor2_1 _10319_ (.Y(_04597_),
    .A(_03285_),
    .B(_04596_));
 sg13g2_nor2_1 _10320_ (.A(net234),
    .B(_04597_),
    .Y(_00312_));
 sg13g2_nor2_1 _10321_ (.A(_03285_),
    .B(_04503_),
    .Y(_04598_));
 sg13g2_o21ai_1 _10322_ (.B1(_04509_),
    .Y(_04599_),
    .A1(_04594_),
    .A2(_04598_));
 sg13g2_xor2_1 _10323_ (.B(_04599_),
    .A(_04450_),
    .X(_04600_));
 sg13g2_nor2_1 _10324_ (.A(net36),
    .B(_04600_),
    .Y(_04601_));
 sg13g2_xnor2_1 _10325_ (.Y(_04602_),
    .A(_03282_),
    .B(_04601_));
 sg13g2_nor2_1 _10326_ (.A(net234),
    .B(_04602_),
    .Y(_00313_));
 sg13g2_nor2_1 _10327_ (.A(_04446_),
    .B(_04514_),
    .Y(_04603_));
 sg13g2_nor3_1 _10328_ (.A(_04435_),
    .B(_04516_),
    .C(_04603_),
    .Y(_04604_));
 sg13g2_xnor2_1 _10329_ (.Y(_04605_),
    .A(_03294_),
    .B(_04604_));
 sg13g2_nor2_1 _10330_ (.A(net234),
    .B(_04605_),
    .Y(_00314_));
 sg13g2_a21oi_1 _10331_ (.A1(net175),
    .A2(_03328_),
    .Y(_00335_),
    .B1(net235));
 sg13g2_inv_1 _10332_ (.Y(_04606_),
    .A(_00082_));
 sg13g2_nand2_1 _10333_ (.Y(_04607_),
    .A(_01399_),
    .B(_01400_));
 sg13g2_nor3_2 _10334_ (.A(_00411_),
    .B(_03890_),
    .C(_04607_),
    .Y(_04608_));
 sg13g2_nand3_1 _10335_ (.B(net382),
    .C(_04608_),
    .A(_05168_),
    .Y(_04609_));
 sg13g2_buf_2 _10336_ (.A(_04609_),
    .X(_04610_));
 sg13g2_nor4_1 _10337_ (.A(_05280_),
    .B(_05383_),
    .C(_01769_),
    .D(_05298_),
    .Y(_04611_));
 sg13g2_nand4_1 _10338_ (.B(net421),
    .C(_00645_),
    .A(net423),
    .Y(_04612_),
    .D(_04611_));
 sg13g2_nor4_1 _10339_ (.A(_05322_),
    .B(net422),
    .C(_04610_),
    .D(_04612_),
    .Y(_04613_));
 sg13g2_or2_1 _10340_ (.X(_04614_),
    .B(_04613_),
    .A(_00085_));
 sg13g2_buf_1 _10341_ (.A(_04614_),
    .X(_04615_));
 sg13g2_nor2_2 _10342_ (.A(_00083_),
    .B(_04610_),
    .Y(_04616_));
 sg13g2_and4_1 _10343_ (.A(net423),
    .B(net422),
    .C(net421),
    .D(_04616_),
    .X(_04617_));
 sg13g2_buf_2 _10344_ (.A(_04617_),
    .X(_04618_));
 sg13g2_nand2_1 _10345_ (.Y(_04619_),
    .A(_00928_),
    .B(_04618_));
 sg13g2_nor3_1 _10346_ (.A(net385),
    .B(_05360_),
    .C(_04619_),
    .Y(_04620_));
 sg13g2_nand2_1 _10347_ (.Y(_04621_),
    .A(net389),
    .B(_04620_));
 sg13g2_or4_1 _10348_ (.A(_01753_),
    .B(_04606_),
    .C(_04615_),
    .D(_04621_),
    .X(_04622_));
 sg13g2_nand2_1 _10349_ (.Y(_04623_),
    .A(_00081_),
    .B(_04622_));
 sg13g2_nand2_1 _10350_ (.Y(_04624_),
    .A(_05293_),
    .B(_04623_));
 sg13g2_nor2_1 _10351_ (.A(net425),
    .B(_04624_),
    .Y(_04625_));
 sg13g2_and3_1 _10352_ (.X(_04626_),
    .A(_05272_),
    .B(net352),
    .C(_04625_));
 sg13g2_buf_1 _10353_ (.A(_04626_),
    .X(_04627_));
 sg13g2_and3_1 _10354_ (.X(_04628_),
    .A(net353),
    .B(_00489_),
    .C(_04627_));
 sg13g2_buf_1 _10355_ (.A(_04628_),
    .X(_04629_));
 sg13g2_nor2b_1 _10356_ (.A(net317),
    .B_N(_04629_),
    .Y(_04630_));
 sg13g2_and4_1 _10357_ (.A(_05272_),
    .B(_05293_),
    .C(_05306_),
    .D(_04623_),
    .X(_04631_));
 sg13g2_nand3_1 _10358_ (.B(net352),
    .C(_04631_),
    .A(net353),
    .Y(_04632_));
 sg13g2_or2_1 _10359_ (.X(_04633_),
    .B(_04632_),
    .A(_01126_));
 sg13g2_buf_1 _10360_ (.A(_04633_),
    .X(_04634_));
 sg13g2_nor3_2 _10361_ (.A(net307),
    .B(_02281_),
    .C(_04634_),
    .Y(_04635_));
 sg13g2_o21ai_1 _10362_ (.B1(net357),
    .Y(_04636_),
    .A1(_04630_),
    .A2(_04635_));
 sg13g2_nand3b_1 _10363_ (.B(_04636_),
    .C(net393),
    .Y(_04637_),
    .A_N(_05262_));
 sg13g2_nand2b_1 _10364_ (.Y(_04638_),
    .B(_04629_),
    .A_N(net317));
 sg13g2_nor3_1 _10365_ (.A(net393),
    .B(_05262_),
    .C(_04638_),
    .Y(_04639_));
 sg13g2_and4_1 _10366_ (.A(net393),
    .B(_05262_),
    .C(_04638_),
    .D(_04635_),
    .X(_04640_));
 sg13g2_o21ai_1 _10367_ (.B1(net357),
    .Y(_04641_),
    .A1(_04639_),
    .A2(_04640_));
 sg13g2_nand3_1 _10368_ (.B(_04637_),
    .C(_04641_),
    .A(net411),
    .Y(_04642_));
 sg13g2_o21ai_1 _10369_ (.B1(_00081_),
    .Y(_04643_),
    .A1(_04622_),
    .A2(_04642_));
 sg13g2_nor3_1 _10370_ (.A(_00467_),
    .B(_04623_),
    .C(_04642_),
    .Y(_04644_));
 sg13g2_a21o_1 _10371_ (.A2(_04643_),
    .A1(_00467_),
    .B1(_04644_),
    .X(_00336_));
 sg13g2_and2_1 _10372_ (.A(_00081_),
    .B(_04642_),
    .X(_04645_));
 sg13g2_buf_1 _10373_ (.A(_04645_),
    .X(_04646_));
 sg13g2_buf_1 _10374_ (.A(_04646_),
    .X(_04647_));
 sg13g2_nand3_1 _10375_ (.B(_05154_),
    .C(_04629_),
    .A(net401),
    .Y(_04648_));
 sg13g2_xnor2_1 _10376_ (.Y(_04649_),
    .A(_05268_),
    .B(_04648_));
 sg13g2_nor2_1 _10377_ (.A(net32),
    .B(_04649_),
    .Y(_00337_));
 sg13g2_xnor2_1 _10378_ (.Y(_04650_),
    .A(net357),
    .B(_04635_));
 sg13g2_nor2_1 _10379_ (.A(net32),
    .B(_04650_),
    .Y(_00338_));
 sg13g2_nand2_1 _10380_ (.Y(_04651_),
    .A(net357),
    .B(_04630_));
 sg13g2_xor2_1 _10381_ (.B(_04651_),
    .A(net393),
    .X(_04652_));
 sg13g2_nor2_1 _10382_ (.A(net32),
    .B(_04652_),
    .Y(_00339_));
 sg13g2_nand3_1 _10383_ (.B(net393),
    .C(_04635_),
    .A(net357),
    .Y(_04653_));
 sg13g2_xnor2_1 _10384_ (.Y(_04654_),
    .A(_05262_),
    .B(_04653_));
 sg13g2_nor2_1 _10385_ (.A(net32),
    .B(_04654_),
    .Y(_00340_));
 sg13g2_xor2_1 _10386_ (.B(_04624_),
    .A(_05306_),
    .X(_04655_));
 sg13g2_nor2_1 _10387_ (.A(_04647_),
    .B(_04655_),
    .Y(_00341_));
 sg13g2_xnor2_1 _10388_ (.Y(_04656_),
    .A(_05272_),
    .B(_04625_));
 sg13g2_nor2_1 _10389_ (.A(net32),
    .B(_04656_),
    .Y(_00342_));
 sg13g2_xnor2_1 _10390_ (.Y(_04657_),
    .A(net352),
    .B(_04631_));
 sg13g2_nor2_1 _10391_ (.A(net32),
    .B(_04657_),
    .Y(_00343_));
 sg13g2_xnor2_1 _10392_ (.Y(_04658_),
    .A(_05216_),
    .B(_04627_));
 sg13g2_nor2_1 _10393_ (.A(_04647_),
    .B(_04658_),
    .Y(_00344_));
 sg13g2_xnor2_1 _10394_ (.Y(_04659_),
    .A(_00471_),
    .B(_04632_));
 sg13g2_nor2_1 _10395_ (.A(net32),
    .B(_04659_),
    .Y(_00345_));
 sg13g2_nor2b_1 _10396_ (.A(_01979_),
    .B_N(_04627_),
    .Y(_04660_));
 sg13g2_xnor2_1 _10397_ (.Y(_04661_),
    .A(net391),
    .B(_04660_));
 sg13g2_nor2_1 _10398_ (.A(net32),
    .B(_04661_),
    .Y(_00346_));
 sg13g2_xnor2_1 _10399_ (.Y(_04662_),
    .A(net372),
    .B(_04634_));
 sg13g2_nor2_1 _10400_ (.A(_04646_),
    .B(_04662_),
    .Y(_00347_));
 sg13g2_nand2_1 _10401_ (.Y(_04663_),
    .A(net351),
    .B(_04629_));
 sg13g2_xnor2_1 _10402_ (.Y(_04664_),
    .A(_05229_),
    .B(_04663_));
 sg13g2_nor2_1 _10403_ (.A(_04646_),
    .B(_04664_),
    .Y(_00348_));
 sg13g2_nor2_1 _10404_ (.A(net307),
    .B(_04634_),
    .Y(_04665_));
 sg13g2_xnor2_1 _10405_ (.Y(_04666_),
    .A(net401),
    .B(_04665_));
 sg13g2_nor2_1 _10406_ (.A(_04646_),
    .B(_04666_),
    .Y(_00349_));
 sg13g2_buf_1 _10407_ (.A(_04615_),
    .X(_04667_));
 sg13g2_xnor2_1 _10408_ (.Y(_04668_),
    .A(_05314_),
    .B(_04610_));
 sg13g2_nor2_1 _10409_ (.A(net138),
    .B(_04668_),
    .Y(_00353_));
 sg13g2_xnor2_1 _10410_ (.Y(_04669_),
    .A(net422),
    .B(_04616_));
 sg13g2_nor2_1 _10411_ (.A(net138),
    .B(_04669_),
    .Y(_00354_));
 sg13g2_nand2_1 _10412_ (.Y(_04670_),
    .A(net422),
    .B(_04616_));
 sg13g2_xnor2_1 _10413_ (.Y(_04671_),
    .A(_05351_),
    .B(_04670_));
 sg13g2_nor2_1 _10414_ (.A(net138),
    .B(_04671_),
    .Y(_00355_));
 sg13g2_nand3_1 _10415_ (.B(net421),
    .C(_04616_),
    .A(net422),
    .Y(_04672_));
 sg13g2_xor2_1 _10416_ (.B(_04672_),
    .A(net423),
    .X(_04673_));
 sg13g2_nor2_1 _10417_ (.A(net138),
    .B(_04673_),
    .Y(_00356_));
 sg13g2_xnor2_1 _10418_ (.Y(_04674_),
    .A(net320),
    .B(_04618_));
 sg13g2_nor2_1 _10419_ (.A(net138),
    .B(_04674_),
    .Y(_00357_));
 sg13g2_nand2_1 _10420_ (.Y(_04675_),
    .A(net320),
    .B(_04618_));
 sg13g2_xor2_1 _10421_ (.B(_04675_),
    .A(_00755_),
    .X(_04676_));
 sg13g2_nor2_1 _10422_ (.A(net138),
    .B(_04676_),
    .Y(_00358_));
 sg13g2_xnor2_1 _10423_ (.Y(_04677_),
    .A(_05360_),
    .B(_04619_));
 sg13g2_nor2_1 _10424_ (.A(net138),
    .B(_04677_),
    .Y(_00359_));
 sg13g2_nand3_1 _10425_ (.B(_00928_),
    .C(_04618_),
    .A(net375),
    .Y(_04678_));
 sg13g2_xnor2_1 _10426_ (.Y(_04679_),
    .A(net385),
    .B(_04678_));
 sg13g2_nor2_1 _10427_ (.A(net138),
    .B(_04679_),
    .Y(_00360_));
 sg13g2_xnor2_1 _10428_ (.Y(_04680_),
    .A(net389),
    .B(_04620_));
 sg13g2_nor2_1 _10429_ (.A(_04667_),
    .B(_04680_),
    .Y(_00361_));
 sg13g2_nor2_1 _10430_ (.A(_00411_),
    .B(_04607_),
    .Y(_04681_));
 sg13g2_or2_1 _10431_ (.X(_04682_),
    .B(_04681_),
    .A(_00085_));
 sg13g2_buf_2 _10432_ (.A(_04682_),
    .X(_04683_));
 sg13g2_xnor2_1 _10433_ (.Y(_04684_),
    .A(net287),
    .B(_03907_));
 sg13g2_nor2_1 _10434_ (.A(_04683_),
    .B(_04684_),
    .Y(_00368_));
 sg13g2_nand2_1 _10435_ (.Y(_04685_),
    .A(_00462_),
    .B(net419));
 sg13g2_xnor2_1 _10436_ (.Y(_04686_),
    .A(_05202_),
    .B(_04685_));
 sg13g2_nor2_1 _10437_ (.A(_04683_),
    .B(_04686_),
    .Y(_00369_));
 sg13g2_nor2_1 _10438_ (.A(_05194_),
    .B(_04685_),
    .Y(_04687_));
 sg13g2_xnor2_1 _10439_ (.Y(_04688_),
    .A(_01807_),
    .B(_04687_));
 sg13g2_nor2_1 _10440_ (.A(_04683_),
    .B(_04688_),
    .Y(_00370_));
 sg13g2_nand3_1 _10441_ (.B(_00450_),
    .C(net348),
    .A(net280),
    .Y(_04689_));
 sg13g2_xnor2_1 _10442_ (.Y(_04690_),
    .A(net326),
    .B(_04689_));
 sg13g2_nor2_1 _10443_ (.A(_04683_),
    .B(_04690_),
    .Y(_00371_));
 sg13g2_nor3_1 _10444_ (.A(_05194_),
    .B(net342),
    .C(_04685_),
    .Y(_04691_));
 sg13g2_xnor2_1 _10445_ (.Y(_04692_),
    .A(net297),
    .B(_04691_));
 sg13g2_nor2_1 _10446_ (.A(_04683_),
    .B(_04692_),
    .Y(_00372_));
 sg13g2_nand3_1 _10447_ (.B(_00450_),
    .C(_01249_),
    .A(net297),
    .Y(_04693_));
 sg13g2_xnor2_1 _10448_ (.Y(_04694_),
    .A(net321),
    .B(_04693_));
 sg13g2_nor2_1 _10449_ (.A(_04683_),
    .B(_04694_),
    .Y(_00373_));
 sg13g2_nand3_1 _10450_ (.B(_00507_),
    .C(_04691_),
    .A(_00539_),
    .Y(_04695_));
 sg13g2_xnor2_1 _10451_ (.Y(_04696_),
    .A(net346),
    .B(_04695_));
 sg13g2_nor2_1 _10452_ (.A(_04683_),
    .B(_04696_),
    .Y(_00374_));
 sg13g2_buf_1 _10453_ (.A(net370),
    .X(_04697_));
 sg13g2_nand3_1 _10454_ (.B(_02232_),
    .C(_02246_),
    .A(net411),
    .Y(_04698_));
 sg13g2_buf_1 _10455_ (.A(_04698_),
    .X(_04699_));
 sg13g2_buf_1 _10456_ (.A(_04699_),
    .X(_04700_));
 sg13g2_nand3_1 _10457_ (.B(_01885_),
    .C(net48),
    .A(net336),
    .Y(_04701_));
 sg13g2_buf_1 _10458_ (.A(_04699_),
    .X(_04702_));
 sg13g2_xnor2_1 _10459_ (.Y(_04703_),
    .A(_01930_),
    .B(_01936_));
 sg13g2_nand2b_1 _10460_ (.Y(_04704_),
    .B(_04703_),
    .A_N(net47));
 sg13g2_nand2_1 _10461_ (.Y(_00098_),
    .A(_04701_),
    .B(_04704_));
 sg13g2_o21ai_1 _10462_ (.B1(_01836_),
    .Y(_04705_),
    .A1(_01837_),
    .A2(net272));
 sg13g2_inv_1 _10463_ (.Y(_04706_),
    .A(net272));
 sg13g2_nand2_1 _10464_ (.Y(_04707_),
    .A(_01837_),
    .B(_04706_));
 sg13g2_a22oi_1 _10465_ (.Y(_04708_),
    .B1(net167),
    .B2(net413),
    .A2(net249),
    .A1(net414));
 sg13g2_o21ai_1 _10466_ (.B1(_04708_),
    .Y(_04709_),
    .A1(net371),
    .A2(_04707_));
 sg13g2_a21oi_2 _10467_ (.B1(_04709_),
    .Y(_04710_),
    .A2(_04705_),
    .A1(net371));
 sg13g2_nand2_1 _10468_ (.Y(_04711_),
    .A(net413),
    .B(_01853_));
 sg13g2_xnor2_1 _10469_ (.Y(_04712_),
    .A(net371),
    .B(_01896_));
 sg13g2_nor2_1 _10470_ (.A(_01857_),
    .B(_04712_),
    .Y(_04713_));
 sg13g2_a221oi_1 _10471_ (.B2(_01837_),
    .C1(_04713_),
    .B1(net167),
    .A1(net415),
    .Y(_04714_),
    .A2(net249));
 sg13g2_nand3_1 _10472_ (.B(_01266_),
    .C(_01615_),
    .A(_05387_),
    .Y(_04715_));
 sg13g2_nor2_1 _10473_ (.A(_01482_),
    .B(_04715_),
    .Y(_04716_));
 sg13g2_o21ai_1 _10474_ (.B1(net411),
    .Y(_04717_),
    .A1(_01387_),
    .A2(_01787_));
 sg13g2_nor2b_1 _10475_ (.A(_04716_),
    .B_N(_04717_),
    .Y(_04718_));
 sg13g2_buf_2 _10476_ (.A(_04718_),
    .X(_04719_));
 sg13g2_buf_1 _10477_ (.A(_04719_),
    .X(_04720_));
 sg13g2_inv_1 _10478_ (.Y(_04721_),
    .A(_00071_));
 sg13g2_mux4_1 _10479_ (.S0(net104),
    .A0(_05150_),
    .A1(_05250_),
    .A2(\dtop.player_inst.synth.alu.registers[4][5] ),
    .A3(_04721_),
    .S1(_02153_),
    .X(_04722_));
 sg13g2_mux2_1 _10480_ (.A0(_00059_),
    .A1(_00073_),
    .S(net85),
    .X(_04723_));
 sg13g2_nand2_1 _10481_ (.Y(_04724_),
    .A(_00072_),
    .B(net85));
 sg13g2_o21ai_1 _10482_ (.B1(_04724_),
    .Y(_04725_),
    .A1(_00403_),
    .A2(net85));
 sg13g2_mux2_1 _10483_ (.A0(_04723_),
    .A1(_04725_),
    .S(net102),
    .X(_04726_));
 sg13g2_nand2_1 _10484_ (.Y(_04727_),
    .A(net103),
    .B(_04726_));
 sg13g2_o21ai_1 _10485_ (.B1(_04727_),
    .Y(_04728_),
    .A1(net103),
    .A2(_04722_));
 sg13g2_nand2_1 _10486_ (.Y(_04729_),
    .A(net99),
    .B(_02105_));
 sg13g2_o21ai_1 _10487_ (.B1(_04729_),
    .Y(_04730_),
    .A1(net99),
    .A2(_04728_));
 sg13g2_nand2_1 _10488_ (.Y(_04731_),
    .A(\dtop.player_inst.synth.alu.registers[0][8] ),
    .B(net127));
 sg13g2_a22oi_1 _10489_ (.Y(_04732_),
    .B1(_01770_),
    .B2(_05306_),
    .A2(net281),
    .A1(\dtop.player_inst.synth.alu.registers[1][8] ));
 sg13g2_a21oi_1 _10490_ (.A1(_02033_),
    .A2(_02037_),
    .Y(_04733_),
    .B1(_02091_));
 sg13g2_buf_2 _10491_ (.A(_04733_),
    .X(_04734_));
 sg13g2_nand2_1 _10492_ (.Y(_04735_),
    .A(net296),
    .B(_02001_));
 sg13g2_nor3_2 _10493_ (.A(_02148_),
    .B(_04734_),
    .C(_04735_),
    .Y(_04736_));
 sg13g2_nor4_1 _10494_ (.A(net296),
    .B(_04734_),
    .C(_02137_),
    .D(_02139_),
    .Y(_04737_));
 sg13g2_nor4_1 _10495_ (.A(_02027_),
    .B(_02093_),
    .C(_02004_),
    .D(_04737_),
    .Y(_04738_));
 sg13g2_inv_1 _10496_ (.Y(_04739_),
    .A(_02101_));
 sg13g2_o21ai_1 _10497_ (.B1(_04739_),
    .Y(_04740_),
    .A1(_04736_),
    .A2(_04738_));
 sg13g2_nand4_1 _10498_ (.B(_04731_),
    .C(_04732_),
    .A(_01750_),
    .Y(_04741_),
    .D(_04740_));
 sg13g2_o21ai_1 _10499_ (.B1(_04741_),
    .Y(_04742_),
    .A1(net86),
    .A2(_04730_));
 sg13g2_xnor2_1 _10500_ (.Y(_04743_),
    .A(net81),
    .B(_04742_));
 sg13g2_nand3_1 _10501_ (.B(_04714_),
    .C(_04743_),
    .A(_04711_),
    .Y(_04744_));
 sg13g2_buf_1 _10502_ (.A(_04744_),
    .X(_04745_));
 sg13g2_nor2b_1 _10503_ (.A(_04710_),
    .B_N(_04745_),
    .Y(_04746_));
 sg13g2_mux2_1 _10504_ (.A0(_00074_),
    .A1(_00075_),
    .S(net85),
    .X(_04747_));
 sg13g2_mux2_1 _10505_ (.A0(_04723_),
    .A1(_04747_),
    .S(net104),
    .X(_04748_));
 sg13g2_nor2_1 _10506_ (.A(_05250_),
    .B(net85),
    .Y(_04749_));
 sg13g2_a21oi_1 _10507_ (.A1(_00071_),
    .A2(net85),
    .Y(_04750_),
    .B1(_04749_));
 sg13g2_nor2_1 _10508_ (.A(net102),
    .B(_04725_),
    .Y(_04751_));
 sg13g2_a21oi_1 _10509_ (.A1(net102),
    .A2(_04750_),
    .Y(_04752_),
    .B1(_04751_));
 sg13g2_mux2_1 _10510_ (.A0(_04748_),
    .A1(_04752_),
    .S(net105),
    .X(_04753_));
 sg13g2_inv_1 _10511_ (.Y(_04754_),
    .A(\dtop.player_inst.synth.alu.registers[4][3] ));
 sg13g2_inv_1 _10512_ (.Y(_04755_),
    .A(\dtop.player_inst.synth.alu.registers[4][2] ));
 sg13g2_mux4_1 _10513_ (.S0(_01597_),
    .A0(_05221_),
    .A1(_00471_),
    .A2(_04754_),
    .A3(_04755_),
    .S1(net101),
    .X(_04756_));
 sg13g2_inv_1 _10514_ (.Y(_04757_),
    .A(\dtop.player_inst.synth.alu.registers[4][5] ));
 sg13g2_inv_1 _10515_ (.Y(_04758_),
    .A(\dtop.player_inst.synth.alu.registers[4][4] ));
 sg13g2_mux4_1 _10516_ (.S0(_01597_),
    .A0(_05229_),
    .A1(net372),
    .A2(_04757_),
    .A3(_04758_),
    .S1(_01736_),
    .X(_04759_));
 sg13g2_mux2_1 _10517_ (.A0(_04756_),
    .A1(_04759_),
    .S(net129),
    .X(_04760_));
 sg13g2_and2_1 _10518_ (.A(net99),
    .B(_04760_),
    .X(_04761_));
 sg13g2_a21oi_1 _10519_ (.A1(_01622_),
    .A2(_04753_),
    .Y(_04762_),
    .B1(_04761_));
 sg13g2_nor2_1 _10520_ (.A(_04734_),
    .B(_02140_),
    .Y(_04763_));
 sg13g2_nor2_1 _10521_ (.A(_02027_),
    .B(_04763_),
    .Y(_04764_));
 sg13g2_o21ai_1 _10522_ (.B1(_04739_),
    .Y(_04765_),
    .A1(_04736_),
    .A2(_04764_));
 sg13g2_nand2_1 _10523_ (.Y(_04766_),
    .A(\dtop.player_inst.synth.alu.registers[0][9] ),
    .B(net127));
 sg13g2_a22oi_1 _10524_ (.Y(_04767_),
    .B1(_01770_),
    .B2(_05272_),
    .A2(net281),
    .A1(\dtop.player_inst.synth.alu.registers[1][9] ));
 sg13g2_nand4_1 _10525_ (.B(_04765_),
    .C(_04766_),
    .A(_01750_),
    .Y(_04768_),
    .D(_04767_));
 sg13g2_o21ai_1 _10526_ (.B1(_04768_),
    .Y(_04769_),
    .A1(net86),
    .A2(_04762_));
 sg13g2_xnor2_1 _10527_ (.Y(_04770_),
    .A(net81),
    .B(_04769_));
 sg13g2_nor2b_1 _10528_ (.A(_04770_),
    .B_N(_04745_),
    .Y(_04771_));
 sg13g2_a21oi_1 _10529_ (.A1(_02111_),
    .A2(_01842_),
    .Y(_04772_),
    .B1(_01387_));
 sg13g2_xnor2_1 _10530_ (.Y(_04773_),
    .A(net371),
    .B(_02113_));
 sg13g2_a22oi_1 _10531_ (.Y(_04774_),
    .B1(_04772_),
    .B2(_04773_),
    .A2(_01821_),
    .A1(net272));
 sg13g2_inv_1 _10532_ (.Y(_04775_),
    .A(_04774_));
 sg13g2_o21ai_1 _10533_ (.B1(_01821_),
    .Y(_04776_),
    .A1(net412),
    .A2(_01855_));
 sg13g2_a22oi_1 _10534_ (.Y(_04777_),
    .B1(_04776_),
    .B2(_04772_),
    .A2(_04775_),
    .A1(_01855_));
 sg13g2_and2_1 _10535_ (.A(_02135_),
    .B(_02140_),
    .X(_04778_));
 sg13g2_nand2b_1 _10536_ (.Y(_04779_),
    .B(_02148_),
    .A_N(_02004_));
 sg13g2_a221oi_1 _10537_ (.B2(_04734_),
    .C1(_04779_),
    .B1(_02002_),
    .A1(_02064_),
    .Y(_04780_),
    .A2(_02073_));
 sg13g2_nor3_1 _10538_ (.A(_04736_),
    .B(_04778_),
    .C(_04780_),
    .Y(_04781_));
 sg13g2_o21ai_1 _10539_ (.B1(_04717_),
    .Y(_04782_),
    .A1(_01482_),
    .A2(_04715_));
 sg13g2_buf_1 _10540_ (.A(_04782_),
    .X(_04783_));
 sg13g2_and2_1 _10541_ (.A(_05383_),
    .B(_01772_),
    .X(_04784_));
 sg13g2_a221oi_1 _10542_ (.B2(\dtop.player_inst.synth.alu.registers[2][5] ),
    .C1(_04784_),
    .B1(_01728_),
    .A1(\dtop.player_inst.synth.alu.registers[1][5] ),
    .Y(_04785_),
    .A2(net281));
 sg13g2_a22oi_1 _10543_ (.Y(_04786_),
    .B1(net259),
    .B2(\dtop.player_inst.synth.alu.registers[5][5] ),
    .A2(net273),
    .A1(_05350_));
 sg13g2_a22oi_1 _10544_ (.Y(_04787_),
    .B1(_01768_),
    .B2(\dtop.player_inst.synth.alu.registers[3][5] ),
    .A2(_01760_),
    .A1(\dtop.player_inst.synth.alu.registers[0][5] ));
 sg13g2_and4_1 _10545_ (.A(_01748_),
    .B(_04785_),
    .C(_04786_),
    .D(_04787_),
    .X(_04788_));
 sg13g2_buf_1 _10546_ (.A(_04788_),
    .X(_04789_));
 sg13g2_inv_1 _10547_ (.Y(_04790_),
    .A(_04789_));
 sg13g2_nor2_1 _10548_ (.A(net111),
    .B(_04790_),
    .Y(_04791_));
 sg13g2_or4_1 _10549_ (.A(_04736_),
    .B(_04790_),
    .C(_04778_),
    .D(_04780_),
    .X(_04792_));
 sg13g2_mux4_1 _10550_ (.S0(_01597_),
    .A0(net353),
    .A1(_05333_),
    .A2(\dtop.player_inst.synth.alu.registers[4][1] ),
    .A3(\dtop.player_inst.synth.alu.registers[4][0] ),
    .S1(net101),
    .X(_04793_));
 sg13g2_a221oi_1 _10551_ (.B2(net129),
    .C1(net128),
    .B1(_04793_),
    .A1(_01864_),
    .Y(_04794_),
    .A2(_01865_));
 sg13g2_a21o_1 _10552_ (.A2(_04760_),
    .A1(_01622_),
    .B1(_04794_),
    .X(_04795_));
 sg13g2_a221oi_1 _10553_ (.B2(_02101_),
    .C1(_04719_),
    .B1(_04789_),
    .A1(_01863_),
    .Y(_04796_),
    .A2(_04795_));
 sg13g2_nor2_1 _10554_ (.A(net100),
    .B(net111),
    .Y(_04797_));
 sg13g2_and3_1 _10555_ (.X(_04798_),
    .A(_02101_),
    .B(_04719_),
    .C(_04789_));
 sg13g2_a21o_1 _10556_ (.A2(_04797_),
    .A1(_04795_),
    .B1(_04798_),
    .X(_04799_));
 sg13g2_a221oi_1 _10557_ (.B2(_04796_),
    .C1(_04799_),
    .B1(_04792_),
    .A1(_04781_),
    .Y(_04800_),
    .A2(_04791_));
 sg13g2_buf_1 _10558_ (.A(_04800_),
    .X(_04801_));
 sg13g2_nor2_1 _10559_ (.A(_04777_),
    .B(_04801_),
    .Y(_04802_));
 sg13g2_xnor2_1 _10560_ (.Y(_04803_),
    .A(_02110_),
    .B(net81));
 sg13g2_nor2_1 _10561_ (.A(_02128_),
    .B(net81),
    .Y(_04804_));
 sg13g2_nor2_1 _10562_ (.A(_02128_),
    .B(net111),
    .Y(_04805_));
 sg13g2_mux2_1 _10563_ (.A0(_04804_),
    .A1(_04805_),
    .S(_02159_),
    .X(_04806_));
 sg13g2_nor3_1 _10564_ (.A(_04802_),
    .B(_04803_),
    .C(_04806_),
    .Y(_04807_));
 sg13g2_inv_1 _10565_ (.Y(_04808_),
    .A(_02120_));
 sg13g2_nor3_1 _10566_ (.A(_04808_),
    .B(_04802_),
    .C(_04806_),
    .Y(_04809_));
 sg13g2_a21o_1 _10567_ (.A2(_01892_),
    .A1(_01881_),
    .B1(_04719_),
    .X(_04810_));
 sg13g2_and2_1 _10568_ (.A(_01914_),
    .B(_04719_),
    .X(_04811_));
 sg13g2_nand4_1 _10569_ (.B(_01892_),
    .C(_01929_),
    .A(_01881_),
    .Y(_04812_),
    .D(_04811_));
 sg13g2_nand3_1 _10570_ (.B(_01899_),
    .C(_01900_),
    .A(_01894_),
    .Y(_04813_));
 sg13g2_nand3_1 _10571_ (.B(_01914_),
    .C(_01929_),
    .A(_04813_),
    .Y(_04814_));
 sg13g2_nand3_1 _10572_ (.B(_01892_),
    .C(_04813_),
    .A(_01881_),
    .Y(_04815_));
 sg13g2_nand4_1 _10573_ (.B(_04812_),
    .C(_04814_),
    .A(_04810_),
    .Y(_04816_),
    .D(_04815_));
 sg13g2_buf_1 _10574_ (.A(_04816_),
    .X(_04817_));
 sg13g2_nor2b_1 _10575_ (.A(_01936_),
    .B_N(_01914_),
    .Y(_04818_));
 sg13g2_nor2_1 _10576_ (.A(net100),
    .B(_01902_),
    .Y(_04819_));
 sg13g2_nand4_1 _10577_ (.B(_01872_),
    .C(_01879_),
    .A(_01866_),
    .Y(_04820_),
    .D(_04819_));
 sg13g2_a21o_1 _10578_ (.A2(net111),
    .A1(_01892_),
    .B1(_01902_),
    .X(_04821_));
 sg13g2_and4_1 _10579_ (.A(_01929_),
    .B(_04818_),
    .C(_04820_),
    .D(_04821_),
    .X(_04822_));
 sg13g2_buf_1 _10580_ (.A(_04822_),
    .X(_04823_));
 sg13g2_nand2b_1 _10581_ (.Y(_04824_),
    .B(_04719_),
    .A_N(_01936_));
 sg13g2_a21oi_1 _10582_ (.A1(_01881_),
    .A2(_01892_),
    .Y(_04825_),
    .B1(_04824_));
 sg13g2_nor3_1 _10583_ (.A(_01860_),
    .B(_04823_),
    .C(_04825_),
    .Y(_04826_));
 sg13g2_or2_1 _10584_ (.X(_04827_),
    .B(net111),
    .A(_01870_));
 sg13g2_a21oi_1 _10585_ (.A1(_01762_),
    .A2(_01778_),
    .Y(_04828_),
    .B1(_04827_));
 sg13g2_mux2_1 _10586_ (.A0(_04716_),
    .A1(_04828_),
    .S(_01744_),
    .X(_04829_));
 sg13g2_nor4_1 _10587_ (.A(_01755_),
    .B(_01756_),
    .C(_01780_),
    .D(net111),
    .Y(_04830_));
 sg13g2_nand2_1 _10588_ (.Y(_04831_),
    .A(net100),
    .B(_04719_));
 sg13g2_nand3_1 _10589_ (.B(_01778_),
    .C(net111),
    .A(_01762_),
    .Y(_04832_));
 sg13g2_o21ai_1 _10590_ (.B1(_04832_),
    .Y(_04833_),
    .A1(_01780_),
    .A2(_04831_));
 sg13g2_nor3_2 _10591_ (.A(_04829_),
    .B(_04830_),
    .C(_04833_),
    .Y(_04834_));
 sg13g2_nor2_1 _10592_ (.A(_01860_),
    .B(_04834_),
    .Y(_04835_));
 sg13g2_a21oi_2 _10593_ (.B1(_04835_),
    .Y(_04836_),
    .A2(_04826_),
    .A1(_04817_));
 sg13g2_and2_1 _10594_ (.A(_02151_),
    .B(_02158_),
    .X(_04837_));
 sg13g2_and2_1 _10595_ (.A(_02128_),
    .B(_04719_),
    .X(_04838_));
 sg13g2_nor3_1 _10596_ (.A(_04834_),
    .B(_04823_),
    .C(_04825_),
    .Y(_04839_));
 sg13g2_nand2_1 _10597_ (.Y(_04840_),
    .A(_02128_),
    .B(_04783_));
 sg13g2_a21oi_1 _10598_ (.A1(_02151_),
    .A2(_02158_),
    .Y(_04841_),
    .B1(_04840_));
 sg13g2_a221oi_1 _10599_ (.B2(_04839_),
    .C1(_04841_),
    .B1(_04817_),
    .A1(_04837_),
    .Y(_04842_),
    .A2(_04838_));
 sg13g2_nand2_1 _10600_ (.Y(_04843_),
    .A(_04836_),
    .B(_04842_));
 sg13g2_o21ai_1 _10601_ (.B1(_04843_),
    .Y(_04844_),
    .A1(_04807_),
    .A2(_04809_));
 sg13g2_nor2_1 _10602_ (.A(_04802_),
    .B(_04803_),
    .Y(_04845_));
 sg13g2_a22oi_1 _10603_ (.Y(_04846_),
    .B1(_04845_),
    .B2(_02120_),
    .A2(_04801_),
    .A1(_04777_));
 sg13g2_inv_2 _10604_ (.Y(_04847_),
    .A(_01896_));
 sg13g2_xnor2_1 _10605_ (.Y(_04848_),
    .A(net371),
    .B(_02111_));
 sg13g2_o21ai_1 _10606_ (.B1(_02172_),
    .Y(_04849_),
    .A1(net272),
    .A2(_04848_));
 sg13g2_a221oi_1 _10607_ (.B2(net412),
    .C1(_04849_),
    .B1(net167),
    .A1(_02113_),
    .Y(_04850_),
    .A2(_01838_));
 sg13g2_o21ai_1 _10608_ (.B1(_04850_),
    .Y(_04851_),
    .A1(_04847_),
    .A2(_01836_));
 sg13g2_inv_1 _10609_ (.Y(_04852_),
    .A(_04851_));
 sg13g2_a21o_1 _10610_ (.A2(_04846_),
    .A1(_04844_),
    .B1(_04852_),
    .X(_04853_));
 sg13g2_nor2_1 _10611_ (.A(_02137_),
    .B(_02139_),
    .Y(_04854_));
 sg13g2_nor3_1 _10612_ (.A(_02148_),
    .B(_04734_),
    .C(_04854_),
    .Y(_04855_));
 sg13g2_o21ai_1 _10613_ (.B1(_02148_),
    .Y(_04856_),
    .A1(_04734_),
    .A2(_04854_));
 sg13g2_a221oi_1 _10614_ (.B2(_02005_),
    .C1(_02101_),
    .B1(_04856_),
    .A1(net296),
    .Y(_04857_),
    .A2(_04855_));
 sg13g2_a21oi_1 _10615_ (.A1(_02093_),
    .A2(_02004_),
    .Y(_04858_),
    .B1(_02140_));
 sg13g2_nand2b_1 _10616_ (.Y(_04859_),
    .B(_02148_),
    .A_N(_04858_));
 sg13g2_nand2_1 _10617_ (.Y(_04860_),
    .A(_05281_),
    .B(_01772_));
 sg13g2_a22oi_1 _10618_ (.Y(_04861_),
    .B1(net282),
    .B2(\dtop.player_inst.synth.alu.registers[2][6] ),
    .A2(_01774_),
    .A1(\dtop.player_inst.synth.alu.registers[1][6] ));
 sg13g2_a22oi_1 _10619_ (.Y(_04862_),
    .B1(_01668_),
    .B2(\dtop.player_inst.synth.alu.registers[5][6] ),
    .A2(net273),
    .A1(_05342_));
 sg13g2_nand4_1 _10620_ (.B(_04860_),
    .C(_04861_),
    .A(net86),
    .Y(_04863_),
    .D(_04862_));
 sg13g2_a21o_1 _10621_ (.A2(_01768_),
    .A1(\dtop.player_inst.synth.alu.registers[3][6] ),
    .B1(_04863_),
    .X(_04864_));
 sg13g2_a221oi_1 _10622_ (.B2(_04859_),
    .C1(_04864_),
    .B1(_04857_),
    .A1(\dtop.player_inst.synth.alu.registers[0][6] ),
    .Y(_04865_),
    .A2(net127));
 sg13g2_mux4_1 _10623_ (.S0(net102),
    .A0(_01508_),
    .A1(_05221_),
    .A2(_04758_),
    .A3(_04754_),
    .S1(_02153_),
    .X(_04866_));
 sg13g2_nor2_1 _10624_ (.A(net105),
    .B(_04722_),
    .Y(_04867_));
 sg13g2_a21oi_1 _10625_ (.A1(net105),
    .A2(_04866_),
    .Y(_04868_),
    .B1(_04867_));
 sg13g2_mux2_1 _10626_ (.A0(_01744_),
    .A1(_04868_),
    .S(net128),
    .X(_04869_));
 sg13g2_nor2_1 _10627_ (.A(net86),
    .B(_04869_),
    .Y(_04870_));
 sg13g2_nor2_1 _10628_ (.A(_04865_),
    .B(_04870_),
    .Y(_04871_));
 sg13g2_xnor2_1 _10629_ (.Y(_04872_),
    .A(net81),
    .B(_04871_));
 sg13g2_nand2_1 _10630_ (.Y(_04873_),
    .A(_04851_),
    .B(_04872_));
 sg13g2_inv_1 _10631_ (.Y(_04874_),
    .A(_04872_));
 sg13g2_a21o_1 _10632_ (.A2(_04846_),
    .A1(_04844_),
    .B1(_04874_),
    .X(_04875_));
 sg13g2_and3_1 _10633_ (.X(_04876_),
    .A(_04853_),
    .B(_04873_),
    .C(_04875_));
 sg13g2_inv_1 _10634_ (.Y(_04877_),
    .A(_01837_));
 sg13g2_xnor2_1 _10635_ (.Y(_04878_),
    .A(net371),
    .B(_01933_));
 sg13g2_nor2_1 _10636_ (.A(net272),
    .B(_04878_),
    .Y(_04879_));
 sg13g2_a221oi_1 _10637_ (.B2(_01896_),
    .C1(_04879_),
    .B1(net167),
    .A1(_01782_),
    .Y(_04880_),
    .A2(net249));
 sg13g2_o21ai_1 _10638_ (.B1(_04880_),
    .Y(_04881_),
    .A1(_04877_),
    .A2(_01836_));
 sg13g2_mux2_1 _10639_ (.A0(_04759_),
    .A1(_04752_),
    .S(_01525_),
    .X(_04882_));
 sg13g2_nor2_1 _10640_ (.A(net128),
    .B(_02152_),
    .Y(_04883_));
 sg13g2_a21oi_1 _10641_ (.A1(net128),
    .A2(_04882_),
    .Y(_04884_),
    .B1(_04883_));
 sg13g2_nand2_1 _10642_ (.Y(_04885_),
    .A(_02148_),
    .B(_04734_));
 sg13g2_a21oi_1 _10643_ (.A1(_04854_),
    .A2(_02004_),
    .Y(_04886_),
    .B1(_02002_));
 sg13g2_nand2b_1 _10644_ (.Y(_04887_),
    .B(_02004_),
    .A_N(_04734_));
 sg13g2_o21ai_1 _10645_ (.B1(_04887_),
    .Y(_04888_),
    .A1(_04885_),
    .A2(_04886_));
 sg13g2_or3_1 _10646_ (.A(_01197_),
    .B(_02027_),
    .C(_02001_),
    .X(_04889_));
 sg13g2_nand4_1 _10647_ (.B(_04854_),
    .C(_04735_),
    .A(_04885_),
    .Y(_04890_),
    .D(_04889_));
 sg13g2_nor2b_1 _10648_ (.A(_04888_),
    .B_N(_04890_),
    .Y(_04891_));
 sg13g2_nand2_1 _10649_ (.Y(_04892_),
    .A(\dtop.player_inst.synth.alu.registers[1][7] ),
    .B(_01774_));
 sg13g2_a22oi_1 _10650_ (.Y(_04893_),
    .B1(_01770_),
    .B2(_05293_),
    .A2(_01728_),
    .A1(\dtop.player_inst.synth.alu.registers[2][7] ));
 sg13g2_nand3_1 _10651_ (.B(_04892_),
    .C(_04893_),
    .A(net86),
    .Y(_04894_));
 sg13g2_a221oi_1 _10652_ (.B2(\dtop.player_inst.synth.alu.registers[3][7] ),
    .C1(_04894_),
    .B1(_01768_),
    .A1(\dtop.player_inst.synth.alu.registers[0][7] ),
    .Y(_04895_),
    .A2(_01761_));
 sg13g2_o21ai_1 _10653_ (.B1(_04895_),
    .Y(_04896_),
    .A1(_02101_),
    .A2(_04891_));
 sg13g2_o21ai_1 _10654_ (.B1(_04896_),
    .Y(_04897_),
    .A1(net86),
    .A2(_04884_));
 sg13g2_xnor2_1 _10655_ (.Y(_04898_),
    .A(_04720_),
    .B(_04897_));
 sg13g2_nor2b_1 _10656_ (.A(_04881_),
    .B_N(_04898_),
    .Y(_04899_));
 sg13g2_nand2b_1 _10657_ (.Y(_04900_),
    .B(_04881_),
    .A_N(_04898_));
 sg13g2_o21ai_1 _10658_ (.B1(_04900_),
    .Y(_04901_),
    .A1(_04876_),
    .A2(_04899_));
 sg13g2_o21ai_1 _10659_ (.B1(_04901_),
    .Y(_04902_),
    .A1(_04746_),
    .A2(_04771_));
 sg13g2_a21o_1 _10660_ (.A2(_04714_),
    .A1(_04711_),
    .B1(_04743_),
    .X(_04903_));
 sg13g2_a21o_1 _10661_ (.A2(_04770_),
    .A1(_04710_),
    .B1(_04903_),
    .X(_04904_));
 sg13g2_or2_1 _10662_ (.X(_04905_),
    .B(_04770_),
    .A(_04710_));
 sg13g2_nand3_1 _10663_ (.B(_04904_),
    .C(_04905_),
    .A(_04902_),
    .Y(_04906_));
 sg13g2_mux2_1 _10664_ (.A0(_05262_),
    .A1(_00076_),
    .S(net85),
    .X(_04907_));
 sg13g2_mux4_1 _10665_ (.S0(net102),
    .A0(_04723_),
    .A1(_04725_),
    .A2(_04907_),
    .A3(_04747_),
    .S1(net103),
    .X(_04908_));
 sg13g2_nor2_1 _10666_ (.A(net99),
    .B(_04908_),
    .Y(_04909_));
 sg13g2_a21oi_1 _10667_ (.A1(net99),
    .A2(_04868_),
    .Y(_04910_),
    .B1(_04909_));
 sg13g2_nor2_1 _10668_ (.A(_00060_),
    .B(_01726_),
    .Y(_04911_));
 sg13g2_and2_1 _10669_ (.A(\dtop.player_inst.synth.alu.registers[1][10] ),
    .B(net281),
    .X(_04912_));
 sg13g2_a221oi_1 _10670_ (.B2(_01747_),
    .C1(_04912_),
    .B1(_04911_),
    .A1(\dtop.player_inst.synth.alu.registers[0][10] ),
    .Y(_04913_),
    .A2(net127));
 sg13g2_o21ai_1 _10671_ (.B1(_04913_),
    .Y(_04914_),
    .A1(net86),
    .A2(_04910_));
 sg13g2_xnor2_1 _10672_ (.Y(_04915_),
    .A(_04720_),
    .B(_04914_));
 sg13g2_inv_1 _10673_ (.Y(_04916_),
    .A(net371));
 sg13g2_and4_1 _10674_ (.A(net413),
    .B(_04706_),
    .C(_01821_),
    .D(_01854_),
    .X(_04917_));
 sg13g2_nor4_1 _10675_ (.A(_04916_),
    .B(_01853_),
    .C(net167),
    .D(_04917_),
    .Y(_04918_));
 sg13g2_o21ai_1 _10676_ (.B1(_04916_),
    .Y(_04919_),
    .A1(net413),
    .A2(_01857_));
 sg13g2_nor2b_1 _10677_ (.A(_04918_),
    .B_N(_04919_),
    .Y(_04920_));
 sg13g2_xor2_1 _10678_ (.B(_04920_),
    .A(_04915_),
    .X(_04921_));
 sg13g2_xnor2_1 _10679_ (.Y(_04922_),
    .A(_04906_),
    .B(_04921_));
 sg13g2_nand3_1 _10680_ (.B(_02114_),
    .C(_04702_),
    .A(_04697_),
    .Y(_04923_));
 sg13g2_o21ai_1 _10681_ (.B1(_04923_),
    .Y(_00099_),
    .A1(_04700_),
    .A2(_04922_));
 sg13g2_nand2_1 _10682_ (.Y(_04924_),
    .A(_01926_),
    .B(_01927_));
 sg13g2_nand2_1 _10683_ (.Y(_04925_),
    .A(_01915_),
    .B(_01923_));
 sg13g2_nand3_1 _10684_ (.B(_01936_),
    .C(net81),
    .A(_04925_),
    .Y(_04926_));
 sg13g2_o21ai_1 _10685_ (.B1(_04926_),
    .Y(_04927_),
    .A1(_01936_),
    .A2(net81));
 sg13g2_nand3_1 _10686_ (.B(_04924_),
    .C(_04927_),
    .A(_01914_),
    .Y(_04928_));
 sg13g2_xnor2_1 _10687_ (.Y(_04929_),
    .A(_01893_),
    .B(_04813_));
 sg13g2_xnor2_1 _10688_ (.Y(_04930_),
    .A(_04928_),
    .B(_04929_));
 sg13g2_nand3_1 _10689_ (.B(net414),
    .C(net47),
    .A(net336),
    .Y(_04931_));
 sg13g2_o21ai_1 _10690_ (.B1(_04931_),
    .Y(_00100_),
    .A1(net48),
    .A2(_04930_));
 sg13g2_nor2_1 _10691_ (.A(_04823_),
    .B(_04825_),
    .Y(_04932_));
 sg13g2_nand2_1 _10692_ (.Y(_04933_),
    .A(_04817_),
    .B(_04932_));
 sg13g2_xnor2_1 _10693_ (.Y(_04934_),
    .A(_01860_),
    .B(_04834_));
 sg13g2_xnor2_1 _10694_ (.Y(_04935_),
    .A(_04933_),
    .B(_04934_));
 sg13g2_nand3_1 _10695_ (.B(net415),
    .C(net47),
    .A(net336),
    .Y(_04936_));
 sg13g2_o21ai_1 _10696_ (.B1(_04936_),
    .Y(_00101_),
    .A1(net48),
    .A2(_04935_));
 sg13g2_o21ai_1 _10697_ (.B1(_04836_),
    .Y(_04937_),
    .A1(_04834_),
    .A2(_04933_));
 sg13g2_xnor2_1 _10698_ (.Y(_04938_),
    .A(_02159_),
    .B(net81));
 sg13g2_xnor2_1 _10699_ (.Y(_04939_),
    .A(_02128_),
    .B(_04938_));
 sg13g2_xnor2_1 _10700_ (.Y(_04940_),
    .A(_04937_),
    .B(_04939_));
 sg13g2_nand3_1 _10701_ (.B(_01782_),
    .C(net47),
    .A(net336),
    .Y(_04941_));
 sg13g2_o21ai_1 _10702_ (.B1(_04941_),
    .Y(_00102_),
    .A1(net48),
    .A2(_04940_));
 sg13g2_a21oi_2 _10703_ (.B1(_04806_),
    .Y(_04942_),
    .A2(_04842_),
    .A1(_04836_));
 sg13g2_xnor2_1 _10704_ (.Y(_04943_),
    .A(_02110_),
    .B(net111));
 sg13g2_xnor2_1 _10705_ (.Y(_04944_),
    .A(_04808_),
    .B(_04943_));
 sg13g2_xnor2_1 _10706_ (.Y(_04945_),
    .A(_04942_),
    .B(_04944_));
 sg13g2_nand3_1 _10707_ (.B(_02113_),
    .C(net47),
    .A(net336),
    .Y(_04946_));
 sg13g2_o21ai_1 _10708_ (.B1(_04946_),
    .Y(_00103_),
    .A1(net48),
    .A2(_04945_));
 sg13g2_nand3_1 _10709_ (.B(_02111_),
    .C(net47),
    .A(net336),
    .Y(_04947_));
 sg13g2_a21oi_1 _10710_ (.A1(_04943_),
    .A2(_04942_),
    .Y(_04948_),
    .B1(_02120_));
 sg13g2_nor2_1 _10711_ (.A(_04943_),
    .B(_04942_),
    .Y(_04949_));
 sg13g2_nor2_1 _10712_ (.A(_04948_),
    .B(_04949_),
    .Y(_04950_));
 sg13g2_xnor2_1 _10713_ (.Y(_04951_),
    .A(_04777_),
    .B(_04801_));
 sg13g2_xnor2_1 _10714_ (.Y(_04952_),
    .A(_04950_),
    .B(_04951_));
 sg13g2_nand2b_1 _10715_ (.Y(_04953_),
    .B(_04952_),
    .A_N(net47));
 sg13g2_nand2_1 _10716_ (.Y(_00104_),
    .A(_04947_),
    .B(_04953_));
 sg13g2_and2_1 _10717_ (.A(_04844_),
    .B(_04846_),
    .X(_04954_));
 sg13g2_xnor2_1 _10718_ (.Y(_04955_),
    .A(_04851_),
    .B(_04872_));
 sg13g2_xnor2_1 _10719_ (.Y(_04956_),
    .A(_04954_),
    .B(_04955_));
 sg13g2_nand3_1 _10720_ (.B(net412),
    .C(net47),
    .A(net336),
    .Y(_04957_));
 sg13g2_o21ai_1 _10721_ (.B1(_04957_),
    .Y(_00105_),
    .A1(net48),
    .A2(_04956_));
 sg13g2_nor2b_1 _10722_ (.A(_04899_),
    .B_N(_04900_),
    .Y(_04958_));
 sg13g2_xor2_1 _10723_ (.B(_04958_),
    .A(_04876_),
    .X(_04959_));
 sg13g2_buf_1 _10724_ (.A(net370),
    .X(_04960_));
 sg13g2_nand3_1 _10725_ (.B(_01896_),
    .C(_04702_),
    .A(net335),
    .Y(_04961_));
 sg13g2_o21ai_1 _10726_ (.B1(_04961_),
    .Y(_00106_),
    .A1(net48),
    .A2(_04959_));
 sg13g2_nand2_1 _10727_ (.Y(_04962_),
    .A(_04903_),
    .B(_04745_));
 sg13g2_xor2_1 _10728_ (.B(_04962_),
    .A(_04901_),
    .X(_04963_));
 sg13g2_nand3_1 _10729_ (.B(_01837_),
    .C(_04699_),
    .A(net335),
    .Y(_04964_));
 sg13g2_o21ai_1 _10730_ (.B1(_04964_),
    .Y(_00107_),
    .A1(_04700_),
    .A2(_04963_));
 sg13g2_inv_1 _10731_ (.Y(_04965_),
    .A(_04903_));
 sg13g2_a21oi_1 _10732_ (.A1(_04901_),
    .A2(_04745_),
    .Y(_04966_),
    .B1(_04965_));
 sg13g2_xnor2_1 _10733_ (.Y(_04967_),
    .A(_04710_),
    .B(_04770_));
 sg13g2_xnor2_1 _10734_ (.Y(_04968_),
    .A(_04966_),
    .B(_04967_));
 sg13g2_nand3_1 _10735_ (.B(net413),
    .C(_04699_),
    .A(net335),
    .Y(_04969_));
 sg13g2_o21ai_1 _10736_ (.B1(_04969_),
    .Y(_00108_),
    .A1(net48),
    .A2(_04968_));
 sg13g2_inv_1 _10737_ (.Y(_04970_),
    .A(\dtop.player_inst.synth.alu.carry ));
 sg13g2_nand2b_1 _10738_ (.Y(_04971_),
    .B(_02232_),
    .A_N(_00085_));
 sg13g2_buf_1 _10739_ (.A(_04971_),
    .X(_04972_));
 sg13g2_or2_1 _10740_ (.X(_04973_),
    .B(_04972_),
    .A(_02247_));
 sg13g2_a21oi_1 _10741_ (.A1(_04915_),
    .A2(_04920_),
    .Y(_04974_),
    .B1(_04973_));
 sg13g2_o21ai_1 _10742_ (.B1(_04906_),
    .Y(_04975_),
    .A1(_04915_),
    .A2(_04920_));
 sg13g2_inv_1 _10743_ (.Y(_04976_),
    .A(net411));
 sg13g2_buf_1 _10744_ (.A(_04976_),
    .X(_04977_));
 sg13g2_a221oi_1 _10745_ (.B2(_04975_),
    .C1(net334),
    .B1(_04974_),
    .A1(_04970_),
    .Y(_00109_),
    .A2(_04973_));
 sg13g2_nand2_1 _10746_ (.Y(_04978_),
    .A(_01397_),
    .B(_01405_));
 sg13g2_nand2_1 _10747_ (.Y(_04979_),
    .A(_01686_),
    .B(_01687_));
 sg13g2_nand4_1 _10748_ (.B(net292),
    .C(net310),
    .A(net311),
    .Y(_04980_),
    .D(_01360_));
 sg13g2_nand3_1 _10749_ (.B(_02174_),
    .C(_04980_),
    .A(_01788_),
    .Y(_04981_));
 sg13g2_nor3_1 _10750_ (.A(_01680_),
    .B(_04979_),
    .C(_04981_),
    .Y(_04982_));
 sg13g2_a21oi_1 _10751_ (.A1(_01249_),
    .A2(net295),
    .Y(_04983_),
    .B1(_01316_));
 sg13g2_nand4_1 _10752_ (.B(_01636_),
    .C(_01646_),
    .A(_01644_),
    .Y(_04984_),
    .D(_04983_));
 sg13g2_nand3_1 _10753_ (.B(_01439_),
    .C(_01360_),
    .A(_01322_),
    .Y(_04985_));
 sg13g2_nand3_1 _10754_ (.B(_01240_),
    .C(_01409_),
    .A(_01456_),
    .Y(_04986_));
 sg13g2_a21oi_1 _10755_ (.A1(_04985_),
    .A2(_04986_),
    .Y(_04987_),
    .B1(_00442_));
 sg13g2_nor3_1 _10756_ (.A(_01329_),
    .B(_04984_),
    .C(_04987_),
    .Y(_04988_));
 sg13g2_a21oi_1 _10757_ (.A1(_00465_),
    .A2(net312),
    .Y(_04989_),
    .B1(_01300_));
 sg13g2_o21ai_1 _10758_ (.B1(_01830_),
    .Y(_04990_),
    .A1(_00462_),
    .A2(_04989_));
 sg13g2_a21oi_1 _10759_ (.A1(net283),
    .A2(_04990_),
    .Y(_04991_),
    .B1(_02237_));
 sg13g2_a221oi_1 _10760_ (.B2(net283),
    .C1(_01363_),
    .B1(_01637_),
    .A1(_01218_),
    .Y(_04992_),
    .A2(_01210_));
 sg13g2_nand4_1 _10761_ (.B(_04988_),
    .C(_04991_),
    .A(_04982_),
    .Y(_04993_),
    .D(_04992_));
 sg13g2_nor3_1 _10762_ (.A(_02197_),
    .B(_04978_),
    .C(_04993_),
    .Y(_04994_));
 sg13g2_nand3_1 _10763_ (.B(_02232_),
    .C(_04994_),
    .A(net411),
    .Y(_04995_));
 sg13g2_buf_1 _10764_ (.A(_04995_),
    .X(_04996_));
 sg13g2_buf_1 _10765_ (.A(_04996_),
    .X(_04997_));
 sg13g2_buf_1 _10766_ (.A(_04996_),
    .X(_04998_));
 sg13g2_nand3_1 _10767_ (.B(\dtop.player_inst.synth.alu.registers[0][0] ),
    .C(net45),
    .A(net335),
    .Y(_04999_));
 sg13g2_o21ai_1 _10768_ (.B1(_04999_),
    .Y(_00111_),
    .A1(_01886_),
    .A2(net46));
 sg13g2_nand3_1 _10769_ (.B(\dtop.player_inst.synth.alu.registers[0][10] ),
    .C(net45),
    .A(net335),
    .Y(_05000_));
 sg13g2_o21ai_1 _10770_ (.B1(_05000_),
    .Y(_00112_),
    .A1(_04916_),
    .A2(net46));
 sg13g2_inv_1 _10771_ (.Y(_05001_),
    .A(net414));
 sg13g2_nand3_1 _10772_ (.B(\dtop.player_inst.synth.alu.registers[0][1] ),
    .C(net45),
    .A(net335),
    .Y(_05002_));
 sg13g2_o21ai_1 _10773_ (.B1(_05002_),
    .Y(_00113_),
    .A1(_05001_),
    .A2(net46));
 sg13g2_inv_1 _10774_ (.Y(_05003_),
    .A(net415));
 sg13g2_nand3_1 _10775_ (.B(\dtop.player_inst.synth.alu.registers[0][2] ),
    .C(net45),
    .A(net335),
    .Y(_05004_));
 sg13g2_o21ai_1 _10776_ (.B1(_05004_),
    .Y(_00114_),
    .A1(_05003_),
    .A2(net46));
 sg13g2_nand3_1 _10777_ (.B(\dtop.player_inst.synth.alu.registers[0][3] ),
    .C(_04998_),
    .A(net335),
    .Y(_05005_));
 sg13g2_o21ai_1 _10778_ (.B1(_05005_),
    .Y(_00115_),
    .A1(_01783_),
    .A2(net46));
 sg13g2_nand3_1 _10779_ (.B(\dtop.player_inst.synth.alu.registers[0][4] ),
    .C(net45),
    .A(_04960_),
    .Y(_05006_));
 sg13g2_o21ai_1 _10780_ (.B1(_05006_),
    .Y(_00116_),
    .A1(_02122_),
    .A2(net46));
 sg13g2_nand3_1 _10781_ (.B(\dtop.player_inst.synth.alu.registers[0][5] ),
    .C(net45),
    .A(_04960_),
    .Y(_05007_));
 sg13g2_o21ai_1 _10782_ (.B1(_05007_),
    .Y(_00117_),
    .A1(_02112_),
    .A2(net46));
 sg13g2_inv_1 _10783_ (.Y(_05008_),
    .A(net412));
 sg13g2_buf_1 _10784_ (.A(net370),
    .X(_05009_));
 sg13g2_nand3_1 _10785_ (.B(\dtop.player_inst.synth.alu.registers[0][6] ),
    .C(net45),
    .A(_05009_),
    .Y(_05010_));
 sg13g2_o21ai_1 _10786_ (.B1(_05010_),
    .Y(_00118_),
    .A1(_05008_),
    .A2(_04997_));
 sg13g2_nand3_1 _10787_ (.B(\dtop.player_inst.synth.alu.registers[0][7] ),
    .C(_04998_),
    .A(_05009_),
    .Y(_05011_));
 sg13g2_o21ai_1 _10788_ (.B1(_05011_),
    .Y(_00119_),
    .A1(_04847_),
    .A2(_04997_));
 sg13g2_nand3_1 _10789_ (.B(\dtop.player_inst.synth.alu.registers[0][8] ),
    .C(_04996_),
    .A(net333),
    .Y(_05012_));
 sg13g2_o21ai_1 _10790_ (.B1(_05012_),
    .Y(_00120_),
    .A1(_04877_),
    .A2(net46));
 sg13g2_inv_1 _10791_ (.Y(_05013_),
    .A(_01895_));
 sg13g2_nand3_1 _10792_ (.B(\dtop.player_inst.synth.alu.registers[0][9] ),
    .C(_04996_),
    .A(net333),
    .Y(_05014_));
 sg13g2_o21ai_1 _10793_ (.B1(_05014_),
    .Y(_00121_),
    .A1(_05013_),
    .A2(net45));
 sg13g2_nand4_1 _10794_ (.B(_01333_),
    .C(_01417_),
    .A(net411),
    .Y(_05015_),
    .D(_02232_));
 sg13g2_buf_1 _10795_ (.A(_05015_),
    .X(_05016_));
 sg13g2_buf_1 _10796_ (.A(_05016_),
    .X(_05017_));
 sg13g2_buf_1 _10797_ (.A(_05016_),
    .X(_05018_));
 sg13g2_nand3_1 _10798_ (.B(\dtop.player_inst.synth.alu.registers[1][0] ),
    .C(net43),
    .A(net333),
    .Y(_05019_));
 sg13g2_o21ai_1 _10799_ (.B1(_05019_),
    .Y(_00122_),
    .A1(_01886_),
    .A2(net44));
 sg13g2_nand3_1 _10800_ (.B(\dtop.player_inst.synth.alu.registers[1][10] ),
    .C(net43),
    .A(net333),
    .Y(_05020_));
 sg13g2_o21ai_1 _10801_ (.B1(_05020_),
    .Y(_00123_),
    .A1(_04916_),
    .A2(net44));
 sg13g2_nand3_1 _10802_ (.B(\dtop.player_inst.synth.alu.registers[1][1] ),
    .C(net43),
    .A(net333),
    .Y(_05021_));
 sg13g2_o21ai_1 _10803_ (.B1(_05021_),
    .Y(_00124_),
    .A1(_05001_),
    .A2(net44));
 sg13g2_nand3_1 _10804_ (.B(\dtop.player_inst.synth.alu.registers[1][2] ),
    .C(net43),
    .A(net333),
    .Y(_05022_));
 sg13g2_o21ai_1 _10805_ (.B1(_05022_),
    .Y(_00125_),
    .A1(_05003_),
    .A2(net44));
 sg13g2_nand3_1 _10806_ (.B(\dtop.player_inst.synth.alu.registers[1][3] ),
    .C(net43),
    .A(net333),
    .Y(_05023_));
 sg13g2_o21ai_1 _10807_ (.B1(_05023_),
    .Y(_00126_),
    .A1(_01783_),
    .A2(net44));
 sg13g2_nand3_1 _10808_ (.B(\dtop.player_inst.synth.alu.registers[1][4] ),
    .C(net43),
    .A(net333),
    .Y(_05024_));
 sg13g2_o21ai_1 _10809_ (.B1(_05024_),
    .Y(_00127_),
    .A1(_02122_),
    .A2(net44));
 sg13g2_buf_1 _10810_ (.A(net411),
    .X(_05025_));
 sg13g2_nand3_1 _10811_ (.B(\dtop.player_inst.synth.alu.registers[1][5] ),
    .C(net43),
    .A(net359),
    .Y(_05026_));
 sg13g2_o21ai_1 _10812_ (.B1(_05026_),
    .Y(_00128_),
    .A1(_02112_),
    .A2(net44));
 sg13g2_nand3_1 _10813_ (.B(\dtop.player_inst.synth.alu.registers[1][6] ),
    .C(_05018_),
    .A(net359),
    .Y(_05027_));
 sg13g2_o21ai_1 _10814_ (.B1(_05027_),
    .Y(_00129_),
    .A1(_05008_),
    .A2(_05017_));
 sg13g2_nand3_1 _10815_ (.B(\dtop.player_inst.synth.alu.registers[1][7] ),
    .C(_05018_),
    .A(net359),
    .Y(_05028_));
 sg13g2_o21ai_1 _10816_ (.B1(_05028_),
    .Y(_00130_),
    .A1(_04847_),
    .A2(_05017_));
 sg13g2_nand3_1 _10817_ (.B(\dtop.player_inst.synth.alu.registers[1][8] ),
    .C(_05016_),
    .A(net359),
    .Y(_05029_));
 sg13g2_o21ai_1 _10818_ (.B1(_05029_),
    .Y(_00131_),
    .A1(_04877_),
    .A2(net44));
 sg13g2_nand3_1 _10819_ (.B(\dtop.player_inst.synth.alu.registers[1][9] ),
    .C(_05016_),
    .A(net359),
    .Y(_05030_));
 sg13g2_o21ai_1 _10820_ (.B1(_05030_),
    .Y(_00132_),
    .A1(_05013_),
    .A2(net43));
 sg13g2_buf_1 _10821_ (.A(net370),
    .X(_05031_));
 sg13g2_or2_1 _10822_ (.X(_05032_),
    .B(_04972_),
    .A(_01682_));
 sg13g2_buf_2 _10823_ (.A(_05032_),
    .X(_05033_));
 sg13g2_buf_1 _10824_ (.A(_05033_),
    .X(_05034_));
 sg13g2_nand2_1 _10825_ (.Y(_05035_),
    .A(\dtop.player_inst.synth.alu.registers[2][0] ),
    .B(net35));
 sg13g2_o21ai_1 _10826_ (.B1(_05035_),
    .Y(_05036_),
    .A1(_01886_),
    .A2(net35));
 sg13g2_and2_1 _10827_ (.A(net332),
    .B(_05036_),
    .X(_00133_));
 sg13g2_nand2_1 _10828_ (.Y(_05037_),
    .A(\dtop.player_inst.synth.alu.registers[2][1] ),
    .B(net35));
 sg13g2_o21ai_1 _10829_ (.B1(_05037_),
    .Y(_05038_),
    .A1(_05001_),
    .A2(net35));
 sg13g2_and2_1 _10830_ (.A(net332),
    .B(_05038_),
    .X(_00134_));
 sg13g2_nand2_1 _10831_ (.Y(_05039_),
    .A(\dtop.player_inst.synth.alu.registers[2][2] ),
    .B(_05033_));
 sg13g2_o21ai_1 _10832_ (.B1(_05039_),
    .Y(_05040_),
    .A1(_05003_),
    .A2(net35));
 sg13g2_and2_1 _10833_ (.A(net332),
    .B(_05040_),
    .X(_00135_));
 sg13g2_nand2_1 _10834_ (.Y(_05041_),
    .A(\dtop.player_inst.synth.alu.registers[2][3] ),
    .B(_05033_));
 sg13g2_o21ai_1 _10835_ (.B1(_05041_),
    .Y(_05042_),
    .A1(_01783_),
    .A2(net35));
 sg13g2_and2_1 _10836_ (.A(net332),
    .B(_05042_),
    .X(_00136_));
 sg13g2_nand2_1 _10837_ (.Y(_05043_),
    .A(\dtop.player_inst.synth.alu.registers[2][4] ),
    .B(_05033_));
 sg13g2_o21ai_1 _10838_ (.B1(_05043_),
    .Y(_05044_),
    .A1(_02122_),
    .A2(net35));
 sg13g2_and2_1 _10839_ (.A(net332),
    .B(_05044_),
    .X(_00137_));
 sg13g2_nand2_1 _10840_ (.Y(_05045_),
    .A(\dtop.player_inst.synth.alu.registers[2][5] ),
    .B(_05033_));
 sg13g2_o21ai_1 _10841_ (.B1(_05045_),
    .Y(_05046_),
    .A1(_02112_),
    .A2(_05034_));
 sg13g2_and2_1 _10842_ (.A(net332),
    .B(_05046_),
    .X(_00138_));
 sg13g2_nand2_1 _10843_ (.Y(_05047_),
    .A(\dtop.player_inst.synth.alu.registers[2][6] ),
    .B(_05033_));
 sg13g2_o21ai_1 _10844_ (.B1(_05047_),
    .Y(_05048_),
    .A1(_05008_),
    .A2(net35));
 sg13g2_and2_1 _10845_ (.A(_05031_),
    .B(_05048_),
    .X(_00139_));
 sg13g2_nand2_1 _10846_ (.Y(_05049_),
    .A(\dtop.player_inst.synth.alu.registers[2][7] ),
    .B(_05033_));
 sg13g2_o21ai_1 _10847_ (.B1(_05049_),
    .Y(_05050_),
    .A1(_04847_),
    .A2(_05034_));
 sg13g2_and2_1 _10848_ (.A(_05031_),
    .B(_05050_),
    .X(_00140_));
 sg13g2_nand4_1 _10849_ (.B(net283),
    .C(_01213_),
    .A(_02170_),
    .Y(_05051_),
    .D(_02232_));
 sg13g2_buf_2 _10850_ (.A(_05051_),
    .X(_05052_));
 sg13g2_buf_1 _10851_ (.A(_05052_),
    .X(_05053_));
 sg13g2_nand3_1 _10852_ (.B(\dtop.player_inst.synth.alu.registers[3][0] ),
    .C(net42),
    .A(_05025_),
    .Y(_05054_));
 sg13g2_o21ai_1 _10853_ (.B1(_05054_),
    .Y(_00141_),
    .A1(_01886_),
    .A2(net42));
 sg13g2_nand3_1 _10854_ (.B(\dtop.player_inst.synth.alu.registers[3][1] ),
    .C(_05053_),
    .A(_05025_),
    .Y(_05055_));
 sg13g2_o21ai_1 _10855_ (.B1(_05055_),
    .Y(_00142_),
    .A1(_05001_),
    .A2(_05053_));
 sg13g2_nand3_1 _10856_ (.B(\dtop.player_inst.synth.alu.registers[3][2] ),
    .C(_05052_),
    .A(net359),
    .Y(_05056_));
 sg13g2_o21ai_1 _10857_ (.B1(_05056_),
    .Y(_00143_),
    .A1(_05003_),
    .A2(net42));
 sg13g2_nand3_1 _10858_ (.B(\dtop.player_inst.synth.alu.registers[3][3] ),
    .C(_05052_),
    .A(net359),
    .Y(_05057_));
 sg13g2_o21ai_1 _10859_ (.B1(_05057_),
    .Y(_00144_),
    .A1(_01783_),
    .A2(net42));
 sg13g2_nand3_1 _10860_ (.B(\dtop.player_inst.synth.alu.registers[3][4] ),
    .C(_05052_),
    .A(net359),
    .Y(_05058_));
 sg13g2_o21ai_1 _10861_ (.B1(_05058_),
    .Y(_00145_),
    .A1(_02122_),
    .A2(net42));
 sg13g2_nand3_1 _10862_ (.B(\dtop.player_inst.synth.alu.registers[3][5] ),
    .C(_05052_),
    .A(net370),
    .Y(_05059_));
 sg13g2_o21ai_1 _10863_ (.B1(_05059_),
    .Y(_00146_),
    .A1(_02112_),
    .A2(net42));
 sg13g2_nand3_1 _10864_ (.B(\dtop.player_inst.synth.alu.registers[3][6] ),
    .C(_05052_),
    .A(_02171_),
    .Y(_05060_));
 sg13g2_o21ai_1 _10865_ (.B1(_05060_),
    .Y(_00147_),
    .A1(_05008_),
    .A2(net42));
 sg13g2_nand3_1 _10866_ (.B(\dtop.player_inst.synth.alu.registers[3][7] ),
    .C(_05052_),
    .A(_02171_),
    .Y(_05061_));
 sg13g2_o21ai_1 _10867_ (.B1(_05061_),
    .Y(_00148_),
    .A1(_04847_),
    .A2(net42));
 sg13g2_or2_1 _10868_ (.X(_05062_),
    .B(_04992_),
    .A(_04972_));
 sg13g2_buf_2 _10869_ (.A(_05062_),
    .X(_05063_));
 sg13g2_buf_1 _10870_ (.A(_05063_),
    .X(_05064_));
 sg13g2_mux2_1 _10871_ (.A0(_01885_),
    .A1(\dtop.player_inst.synth.alu.registers[4][0] ),
    .S(net34),
    .X(_05065_));
 sg13g2_and2_1 _10872_ (.A(net332),
    .B(_05065_),
    .X(_00149_));
 sg13g2_buf_1 _10873_ (.A(net370),
    .X(_05066_));
 sg13g2_mux2_1 _10874_ (.A0(_02114_),
    .A1(\dtop.player_inst.synth.alu.registers[4][10] ),
    .S(net34),
    .X(_05067_));
 sg13g2_and2_1 _10875_ (.A(net331),
    .B(_05067_),
    .X(_00150_));
 sg13g2_mux2_1 _10876_ (.A0(net414),
    .A1(\dtop.player_inst.synth.alu.registers[4][1] ),
    .S(net34),
    .X(_05068_));
 sg13g2_and2_1 _10877_ (.A(net331),
    .B(_05068_),
    .X(_00151_));
 sg13g2_mux2_1 _10878_ (.A0(net415),
    .A1(\dtop.player_inst.synth.alu.registers[4][2] ),
    .S(net34),
    .X(_05069_));
 sg13g2_and2_1 _10879_ (.A(net331),
    .B(_05069_),
    .X(_00152_));
 sg13g2_nor2_1 _10880_ (.A(_01783_),
    .B(_05064_),
    .Y(_05070_));
 sg13g2_a21oi_1 _10881_ (.A1(\dtop.player_inst.synth.alu.registers[4][3] ),
    .A2(net34),
    .Y(_05071_),
    .B1(_05070_));
 sg13g2_nor2_1 _10882_ (.A(net334),
    .B(_05071_),
    .Y(_00153_));
 sg13g2_nor2_1 _10883_ (.A(_02122_),
    .B(_05064_),
    .Y(_05072_));
 sg13g2_a21oi_1 _10884_ (.A1(\dtop.player_inst.synth.alu.registers[4][4] ),
    .A2(net34),
    .Y(_05073_),
    .B1(_05072_));
 sg13g2_nor2_1 _10885_ (.A(net334),
    .B(_05073_),
    .Y(_00154_));
 sg13g2_mux2_1 _10886_ (.A0(_02111_),
    .A1(\dtop.player_inst.synth.alu.registers[4][5] ),
    .S(_05063_),
    .X(_05074_));
 sg13g2_and2_1 _10887_ (.A(net331),
    .B(_05074_),
    .X(_00155_));
 sg13g2_mux2_1 _10888_ (.A0(net412),
    .A1(\dtop.player_inst.synth.alu.registers[4][6] ),
    .S(_05063_),
    .X(_05075_));
 sg13g2_and2_1 _10889_ (.A(net331),
    .B(_05075_),
    .X(_00156_));
 sg13g2_nand2_1 _10890_ (.Y(_05076_),
    .A(\dtop.player_inst.synth.alu.registers[4][7] ),
    .B(_05063_));
 sg13g2_o21ai_1 _10891_ (.B1(_05076_),
    .Y(_05077_),
    .A1(_04847_),
    .A2(net34));
 sg13g2_and2_1 _10892_ (.A(net331),
    .B(_05077_),
    .X(_00157_));
 sg13g2_nand2_1 _10893_ (.Y(_05078_),
    .A(\dtop.player_inst.synth.alu.registers[4][8] ),
    .B(_05063_));
 sg13g2_o21ai_1 _10894_ (.B1(_05078_),
    .Y(_05079_),
    .A1(_04877_),
    .A2(net34));
 sg13g2_and2_1 _10895_ (.A(net331),
    .B(_05079_),
    .X(_00158_));
 sg13g2_mux2_1 _10896_ (.A0(net413),
    .A1(\dtop.player_inst.synth.alu.registers[4][9] ),
    .S(_05063_),
    .X(_05080_));
 sg13g2_and2_1 _10897_ (.A(net331),
    .B(_05080_),
    .X(_00159_));
 sg13g2_or2_1 _10898_ (.X(_05081_),
    .B(_04982_),
    .A(_04972_));
 sg13g2_buf_1 _10899_ (.A(_05081_),
    .X(_05082_));
 sg13g2_mux2_1 _10900_ (.A0(_01885_),
    .A1(\dtop.player_inst.synth.alu.registers[5][0] ),
    .S(net39),
    .X(_05083_));
 sg13g2_and2_1 _10901_ (.A(_05066_),
    .B(_05083_),
    .X(_00160_));
 sg13g2_mux2_1 _10902_ (.A0(_01850_),
    .A1(\dtop.player_inst.synth.alu.registers[5][1] ),
    .S(net39),
    .X(_05084_));
 sg13g2_and2_1 _10903_ (.A(_05066_),
    .B(_05084_),
    .X(_00161_));
 sg13g2_buf_1 _10904_ (.A(net370),
    .X(_05085_));
 sg13g2_mux2_1 _10905_ (.A0(net415),
    .A1(\dtop.player_inst.synth.alu.registers[5][2] ),
    .S(net39),
    .X(_05086_));
 sg13g2_and2_1 _10906_ (.A(net330),
    .B(_05086_),
    .X(_00162_));
 sg13g2_nand2_1 _10907_ (.Y(_05087_),
    .A(\dtop.player_inst.synth.alu.registers[5][3] ),
    .B(net39));
 sg13g2_o21ai_1 _10908_ (.B1(_05087_),
    .Y(_05088_),
    .A1(_01783_),
    .A2(net39));
 sg13g2_and2_1 _10909_ (.A(net330),
    .B(_05088_),
    .X(_00163_));
 sg13g2_nand2_1 _10910_ (.Y(_05089_),
    .A(\dtop.player_inst.synth.alu.registers[5][4] ),
    .B(_05082_));
 sg13g2_o21ai_1 _10911_ (.B1(_05089_),
    .Y(_05090_),
    .A1(_02122_),
    .A2(net39));
 sg13g2_and2_1 _10912_ (.A(net330),
    .B(_05090_),
    .X(_00164_));
 sg13g2_mux2_1 _10913_ (.A0(_02111_),
    .A1(\dtop.player_inst.synth.alu.registers[5][5] ),
    .S(net39),
    .X(_05091_));
 sg13g2_and2_1 _10914_ (.A(net330),
    .B(_05091_),
    .X(_00165_));
 sg13g2_mux2_1 _10915_ (.A0(net412),
    .A1(\dtop.player_inst.synth.alu.registers[5][6] ),
    .S(net39),
    .X(_05092_));
 sg13g2_and2_1 _10916_ (.A(net330),
    .B(_05092_),
    .X(_00166_));
 sg13g2_or2_1 _10917_ (.X(_05093_),
    .B(_04972_),
    .A(_04607_));
 sg13g2_buf_1 _10918_ (.A(_05093_),
    .X(_05094_));
 sg13g2_mux2_1 _10919_ (.A0(_01885_),
    .A1(\dtop.out_sample[0] ),
    .S(net38),
    .X(_05095_));
 sg13g2_and2_1 _10920_ (.A(net330),
    .B(_05095_),
    .X(_00167_));
 sg13g2_mux2_1 _10921_ (.A0(net414),
    .A1(\dtop.out_sample[1] ),
    .S(net38),
    .X(_05096_));
 sg13g2_and2_1 _10922_ (.A(net330),
    .B(_05096_),
    .X(_00168_));
 sg13g2_mux2_1 _10923_ (.A0(_01846_),
    .A1(\dtop.out_sample[2] ),
    .S(net38),
    .X(_05097_));
 sg13g2_and2_1 _10924_ (.A(_05085_),
    .B(_05097_),
    .X(_00169_));
 sg13g2_nand2_1 _10925_ (.Y(_05098_),
    .A(\dtop.out_sample[3] ),
    .B(net38));
 sg13g2_o21ai_1 _10926_ (.B1(_05098_),
    .Y(_05099_),
    .A1(_01783_),
    .A2(_05094_));
 sg13g2_and2_1 _10927_ (.A(_05085_),
    .B(_05099_),
    .X(_00170_));
 sg13g2_nor2_1 _10928_ (.A(_02122_),
    .B(net38),
    .Y(_05100_));
 sg13g2_a21oi_1 _10929_ (.A1(\dtop.out_sample[4] ),
    .A2(net38),
    .Y(_05101_),
    .B1(_05100_));
 sg13g2_nor2_1 _10930_ (.A(net334),
    .B(_05101_),
    .Y(_00171_));
 sg13g2_mux2_1 _10931_ (.A0(_02111_),
    .A1(\dtop.out_sample[5] ),
    .S(net38),
    .X(_05102_));
 sg13g2_and2_1 _10932_ (.A(net330),
    .B(_05102_),
    .X(_00172_));
 sg13g2_mux2_1 _10933_ (.A0(net412),
    .A1(\dtop.out_sample[6] ),
    .S(net38),
    .X(_05103_));
 sg13g2_and2_1 _10934_ (.A(_04697_),
    .B(_05103_),
    .X(_00173_));
 sg13g2_nand3b_1 _10935_ (.B(_01769_),
    .C(_00792_),
    .Y(_05104_),
    .A_N(_00083_));
 sg13g2_nor4_1 _10936_ (.A(_00063_),
    .B(_00062_),
    .C(_00061_),
    .D(_05104_),
    .Y(_05105_));
 sg13g2_mux2_1 _10937_ (.A0(_03887_),
    .A1(_03889_),
    .S(net422),
    .X(_05106_));
 sg13g2_nand2_1 _10938_ (.Y(_05107_),
    .A(_00066_),
    .B(_05106_));
 sg13g2_or4_1 _10939_ (.A(_00730_),
    .B(_05301_),
    .C(_03888_),
    .D(_03887_),
    .X(_05108_));
 sg13g2_o21ai_1 _10940_ (.B1(_05108_),
    .Y(_05109_),
    .A1(_00688_),
    .A2(_05107_));
 sg13g2_nand2_1 _10941_ (.Y(_05110_),
    .A(_03888_),
    .B(_03887_));
 sg13g2_nor3_1 _10942_ (.A(net320),
    .B(_05346_),
    .C(_05110_),
    .Y(_05111_));
 sg13g2_a21oi_1 _10943_ (.A1(_05105_),
    .A2(_05109_),
    .Y(_05112_),
    .B1(_05111_));
 sg13g2_and4_1 _10944_ (.A(_01753_),
    .B(_00063_),
    .C(_00062_),
    .D(_00061_),
    .X(_05113_));
 sg13g2_a21oi_1 _10945_ (.A1(_00083_),
    .A2(_05113_),
    .Y(_05114_),
    .B1(_05110_));
 sg13g2_nor3_1 _10946_ (.A(net343),
    .B(_00066_),
    .C(_05114_),
    .Y(_05115_));
 sg13g2_a21oi_1 _10947_ (.A1(net319),
    .A2(_05110_),
    .Y(_05116_),
    .B1(_05115_));
 sg13g2_nor4_2 _10948_ (.A(_00449_),
    .B(_04610_),
    .C(_05112_),
    .Y(_05117_),
    .D(_05116_));
 sg13g2_xnor2_1 _10949_ (.Y(_05118_),
    .A(_03887_),
    .B(_05117_));
 sg13g2_nor2_1 _10950_ (.A(net334),
    .B(_05118_),
    .Y(_00351_));
 sg13g2_nand2_1 _10951_ (.Y(_05119_),
    .A(_03887_),
    .B(_05117_));
 sg13g2_xor2_1 _10952_ (.B(_05119_),
    .A(_03888_),
    .X(_05120_));
 sg13g2_nor2_1 _10953_ (.A(net334),
    .B(_05120_),
    .Y(_00352_));
 sg13g2_xnor2_1 _10954_ (.Y(_05121_),
    .A(_01769_),
    .B(_04621_));
 sg13g2_nor3_1 _10955_ (.A(_04976_),
    .B(_04667_),
    .C(_05121_),
    .Y(_00362_));
 sg13g2_xnor2_1 _10956_ (.Y(_05122_),
    .A(_03897_),
    .B(_03904_));
 sg13g2_nor2_1 _10957_ (.A(net334),
    .B(_05122_),
    .Y(_00363_));
 sg13g2_nand2_1 _10958_ (.Y(_05123_),
    .A(_03897_),
    .B(_03904_));
 sg13g2_xnor2_1 _10959_ (.Y(_05124_),
    .A(_03894_),
    .B(_05123_));
 sg13g2_nand2_1 _10960_ (.Y(_00364_),
    .A(net332),
    .B(_05124_));
 sg13g2_xnor2_1 _10961_ (.Y(_05125_),
    .A(net395),
    .B(_04681_));
 sg13g2_nor2_1 _10962_ (.A(_04977_),
    .B(_05125_),
    .Y(_00365_));
 sg13g2_xnor2_1 _10963_ (.Y(_05126_),
    .A(net378),
    .B(_04608_));
 sg13g2_nor2_1 _10964_ (.A(net334),
    .B(_05126_),
    .Y(_00366_));
 sg13g2_nand2_1 _10965_ (.Y(_05127_),
    .A(net378),
    .B(_04608_));
 sg13g2_xnor2_1 _10966_ (.Y(_05128_),
    .A(_00515_),
    .B(_05127_));
 sg13g2_nor2_1 _10967_ (.A(_04977_),
    .B(_05128_),
    .Y(_00367_));
 sg13g2_and2_1 _10968_ (.A(_00411_),
    .B(net336),
    .X(_00375_));
 sg13g2_dfrbp_1 _10969_ (.CLK(clknet_leaf_17_clk),
    .RESET_B(net430),
    .D(_00096_),
    .Q_N(_05630_),
    .Q(\dtop.vtop.logo_d[1] ));
 sg13g2_dfrbp_1 _10970_ (.CLK(clknet_leaf_16_clk),
    .RESET_B(net431),
    .D(_00097_),
    .Q_N(_05629_),
    .Q(\dtop.vtop.force_sat0 ));
 sg13g2_buf_4 clkbuf_leaf_0_clk (.X(clknet_leaf_0_clk),
    .A(clknet_4_0_0_clk));
 sg13g2_buf_1 _10972_ (.A(net15),
    .X(net10));
 sg13g2_buf_1 _10973_ (.A(net15),
    .X(net11));
 sg13g2_buf_1 _10974_ (.A(net15),
    .X(net12));
 sg13g2_buf_1 _10975_ (.A(net15),
    .X(net13));
 sg13g2_buf_1 _10976_ (.A(net15),
    .X(net14));
 sg13g2_buf_1 _10977_ (.A(net432),
    .X(uio_oe[6]));
 sg13g2_buf_1 _10978_ (.A(net433),
    .X(uio_oe[7]));
 sg13g2_dfrbp_1 \dtop.player_inst.synth.alu.acc[0]$_SDFFE_PN0P_  (.CLK(clknet_leaf_24_clk),
    .RESET_B(net434),
    .D(_00098_),
    .Q_N(_05628_),
    .Q(\dtop.player_inst.synth.alu.acc[0] ));
 sg13g2_dfrbp_1 \dtop.player_inst.synth.alu.acc[10]$_SDFFE_PN0P_  (.CLK(clknet_leaf_27_clk),
    .RESET_B(net435),
    .D(_00099_),
    .Q_N(_00060_),
    .Q(\dtop.player_inst.synth.alu.acc[10] ));
 sg13g2_dfrbp_1 \dtop.player_inst.synth.alu.acc[1]$_SDFFE_PN0P_  (.CLK(clknet_leaf_24_clk),
    .RESET_B(net436),
    .D(_00100_),
    .Q_N(_05627_),
    .Q(\dtop.player_inst.synth.alu.acc[1] ));
 sg13g2_dfrbp_1 \dtop.player_inst.synth.alu.acc[2]$_SDFFE_PN0P_  (.CLK(clknet_leaf_24_clk),
    .RESET_B(net437),
    .D(_00101_),
    .Q_N(_05626_),
    .Q(\dtop.player_inst.synth.alu.acc[2] ));
 sg13g2_dfrbp_1 \dtop.player_inst.synth.alu.acc[3]$_SDFFE_PN0P_  (.CLK(clknet_leaf_24_clk),
    .RESET_B(net438),
    .D(_00102_),
    .Q_N(_05625_),
    .Q(\dtop.player_inst.synth.alu.acc[3] ));
 sg13g2_dfrbp_1 \dtop.player_inst.synth.alu.acc[4]$_SDFFE_PN0P_  (.CLK(clknet_leaf_24_clk),
    .RESET_B(net439),
    .D(_00103_),
    .Q_N(_05624_),
    .Q(\dtop.player_inst.synth.alu.acc[4] ));
 sg13g2_dfrbp_1 \dtop.player_inst.synth.alu.acc[5]$_SDFFE_PN0P_  (.CLK(clknet_leaf_24_clk),
    .RESET_B(net440),
    .D(_00104_),
    .Q_N(_05623_),
    .Q(\dtop.player_inst.synth.alu.acc[5] ));
 sg13g2_dfrbp_1 \dtop.player_inst.synth.alu.acc[6]$_SDFFE_PN0P_  (.CLK(clknet_leaf_18_clk),
    .RESET_B(net441),
    .D(_00105_),
    .Q_N(_05622_),
    .Q(\dtop.player_inst.synth.alu.acc[6] ));
 sg13g2_dfrbp_1 \dtop.player_inst.synth.alu.acc[7]$_SDFFE_PN0P_  (.CLK(clknet_4_13_0_clk),
    .RESET_B(net442),
    .D(_00106_),
    .Q_N(_05621_),
    .Q(\dtop.player_inst.synth.alu.acc[7] ));
 sg13g2_dfrbp_1 \dtop.player_inst.synth.alu.acc[8]$_SDFFE_PN0P_  (.CLK(clknet_leaf_27_clk),
    .RESET_B(net443),
    .D(_00107_),
    .Q_N(_05620_),
    .Q(\dtop.player_inst.synth.alu.acc[8] ));
 sg13g2_dfrbp_1 \dtop.player_inst.synth.alu.acc[9]$_SDFFE_PN0P_  (.CLK(clknet_leaf_27_clk),
    .RESET_B(net444),
    .D(_00108_),
    .Q_N(_05619_),
    .Q(\dtop.player_inst.synth.alu.acc[9] ));
 sg13g2_dfrbp_1 \dtop.player_inst.synth.alu.carry$_SDFFE_PN0P_  (.CLK(clknet_leaf_26_clk),
    .RESET_B(net445),
    .D(_00109_),
    .Q_N(_05618_),
    .Q(\dtop.player_inst.synth.alu.carry ));
 sg13g2_dfrbp_1 \dtop.player_inst.synth.alu.oct_en$_DFFE_PP_  (.CLK(clknet_leaf_26_clk),
    .RESET_B(net446),
    .D(_00110_),
    .Q_N(_05617_),
    .Q(\dtop.player_inst.synth.alu.oct_en ));
 sg13g2_dfrbp_1 \dtop.player_inst.synth.alu.registers[0][0]$_SDFFE_PN0P_  (.CLK(clknet_leaf_27_clk),
    .RESET_B(net447),
    .D(_00111_),
    .Q_N(_05616_),
    .Q(\dtop.player_inst.synth.alu.registers[0][0] ));
 sg13g2_dfrbp_1 \dtop.player_inst.synth.alu.registers[0][10]$_SDFFE_PN0P_  (.CLK(clknet_leaf_27_clk),
    .RESET_B(net448),
    .D(_00112_),
    .Q_N(_05615_),
    .Q(\dtop.player_inst.synth.alu.registers[0][10] ));
 sg13g2_dfrbp_1 \dtop.player_inst.synth.alu.registers[0][1]$_SDFFE_PN0P_  (.CLK(clknet_leaf_28_clk),
    .RESET_B(net449),
    .D(_00113_),
    .Q_N(_05614_),
    .Q(\dtop.player_inst.synth.alu.registers[0][1] ));
 sg13g2_dfrbp_1 \dtop.player_inst.synth.alu.registers[0][2]$_SDFFE_PN0P_  (.CLK(clknet_leaf_28_clk),
    .RESET_B(net450),
    .D(_00114_),
    .Q_N(_05613_),
    .Q(\dtop.player_inst.synth.alu.registers[0][2] ));
 sg13g2_dfrbp_1 \dtop.player_inst.synth.alu.registers[0][3]$_SDFFE_PN0P_  (.CLK(clknet_leaf_28_clk),
    .RESET_B(net451),
    .D(_00115_),
    .Q_N(_05612_),
    .Q(\dtop.player_inst.synth.alu.registers[0][3] ));
 sg13g2_dfrbp_1 \dtop.player_inst.synth.alu.registers[0][4]$_SDFFE_PN0P_  (.CLK(clknet_leaf_28_clk),
    .RESET_B(net452),
    .D(_00116_),
    .Q_N(_05611_),
    .Q(\dtop.player_inst.synth.alu.registers[0][4] ));
 sg13g2_dfrbp_1 \dtop.player_inst.synth.alu.registers[0][5]$_SDFFE_PN0P_  (.CLK(clknet_leaf_27_clk),
    .RESET_B(net453),
    .D(_00117_),
    .Q_N(_05610_),
    .Q(\dtop.player_inst.synth.alu.registers[0][5] ));
 sg13g2_dfrbp_1 \dtop.player_inst.synth.alu.registers[0][6]$_SDFFE_PN0P_  (.CLK(clknet_leaf_29_clk),
    .RESET_B(net454),
    .D(_00118_),
    .Q_N(_05609_),
    .Q(\dtop.player_inst.synth.alu.registers[0][6] ));
 sg13g2_dfrbp_1 \dtop.player_inst.synth.alu.registers[0][7]$_SDFFE_PN0P_  (.CLK(clknet_leaf_29_clk),
    .RESET_B(net455),
    .D(_00119_),
    .Q_N(_05608_),
    .Q(\dtop.player_inst.synth.alu.registers[0][7] ));
 sg13g2_dfrbp_1 \dtop.player_inst.synth.alu.registers[0][8]$_SDFFE_PN0P_  (.CLK(clknet_leaf_27_clk),
    .RESET_B(net456),
    .D(_00120_),
    .Q_N(_05607_),
    .Q(\dtop.player_inst.synth.alu.registers[0][8] ));
 sg13g2_dfrbp_1 \dtop.player_inst.synth.alu.registers[0][9]$_SDFFE_PN0P_  (.CLK(clknet_leaf_26_clk),
    .RESET_B(net457),
    .D(_00121_),
    .Q_N(_05606_),
    .Q(\dtop.player_inst.synth.alu.registers[0][9] ));
 sg13g2_dfrbp_1 \dtop.player_inst.synth.alu.registers[1][0]$_SDFFE_PN0P_  (.CLK(clknet_leaf_31_clk),
    .RESET_B(net458),
    .D(_00122_),
    .Q_N(_05605_),
    .Q(\dtop.player_inst.synth.alu.registers[1][0] ));
 sg13g2_dfrbp_1 \dtop.player_inst.synth.alu.registers[1][10]$_SDFFE_PN0P_  (.CLK(clknet_leaf_26_clk),
    .RESET_B(net459),
    .D(_00123_),
    .Q_N(_05604_),
    .Q(\dtop.player_inst.synth.alu.registers[1][10] ));
 sg13g2_dfrbp_1 \dtop.player_inst.synth.alu.registers[1][1]$_SDFFE_PN0P_  (.CLK(clknet_leaf_31_clk),
    .RESET_B(net460),
    .D(_00124_),
    .Q_N(_05603_),
    .Q(\dtop.player_inst.synth.alu.registers[1][1] ));
 sg13g2_dfrbp_1 \dtop.player_inst.synth.alu.registers[1][2]$_SDFFE_PN0P_  (.CLK(clknet_leaf_30_clk),
    .RESET_B(net461),
    .D(_00125_),
    .Q_N(_05602_),
    .Q(\dtop.player_inst.synth.alu.registers[1][2] ));
 sg13g2_dfrbp_1 \dtop.player_inst.synth.alu.registers[1][3]$_SDFFE_PN0P_  (.CLK(clknet_leaf_31_clk),
    .RESET_B(net462),
    .D(_00126_),
    .Q_N(_05601_),
    .Q(\dtop.player_inst.synth.alu.registers[1][3] ));
 sg13g2_dfrbp_1 \dtop.player_inst.synth.alu.registers[1][4]$_SDFFE_PN0P_  (.CLK(clknet_leaf_31_clk),
    .RESET_B(net463),
    .D(_00127_),
    .Q_N(_05600_),
    .Q(\dtop.player_inst.synth.alu.registers[1][4] ));
 sg13g2_dfrbp_1 \dtop.player_inst.synth.alu.registers[1][5]$_SDFFE_PN0P_  (.CLK(clknet_leaf_31_clk),
    .RESET_B(net464),
    .D(_00128_),
    .Q_N(_05599_),
    .Q(\dtop.player_inst.synth.alu.registers[1][5] ));
 sg13g2_dfrbp_1 \dtop.player_inst.synth.alu.registers[1][6]$_SDFFE_PN0P_  (.CLK(clknet_leaf_29_clk),
    .RESET_B(net465),
    .D(_00129_),
    .Q_N(_05598_),
    .Q(\dtop.player_inst.synth.alu.registers[1][6] ));
 sg13g2_dfrbp_1 \dtop.player_inst.synth.alu.registers[1][7]$_SDFFE_PN0P_  (.CLK(clknet_leaf_29_clk),
    .RESET_B(net466),
    .D(_00130_),
    .Q_N(_05597_),
    .Q(\dtop.player_inst.synth.alu.registers[1][7] ));
 sg13g2_dfrbp_1 \dtop.player_inst.synth.alu.registers[1][8]$_SDFFE_PN0P_  (.CLK(clknet_leaf_26_clk),
    .RESET_B(net467),
    .D(_00131_),
    .Q_N(_05596_),
    .Q(\dtop.player_inst.synth.alu.registers[1][8] ));
 sg13g2_dfrbp_1 \dtop.player_inst.synth.alu.registers[1][9]$_SDFFE_PN0P_  (.CLK(clknet_leaf_26_clk),
    .RESET_B(net468),
    .D(_00132_),
    .Q_N(_05595_),
    .Q(\dtop.player_inst.synth.alu.registers[1][9] ));
 sg13g2_dfrbp_1 \dtop.player_inst.synth.alu.registers[2][0]$_SDFFE_PN0P_  (.CLK(clknet_leaf_30_clk),
    .RESET_B(net469),
    .D(_00133_),
    .Q_N(_05594_),
    .Q(\dtop.player_inst.synth.alu.registers[2][0] ));
 sg13g2_dfrbp_1 \dtop.player_inst.synth.alu.registers[2][1]$_SDFFE_PN0P_  (.CLK(clknet_leaf_30_clk),
    .RESET_B(net470),
    .D(_00134_),
    .Q_N(_05593_),
    .Q(\dtop.player_inst.synth.alu.registers[2][1] ));
 sg13g2_dfrbp_1 \dtop.player_inst.synth.alu.registers[2][2]$_SDFFE_PN0P_  (.CLK(clknet_leaf_30_clk),
    .RESET_B(net471),
    .D(_00135_),
    .Q_N(_05592_),
    .Q(\dtop.player_inst.synth.alu.registers[2][2] ));
 sg13g2_dfrbp_1 \dtop.player_inst.synth.alu.registers[2][3]$_SDFFE_PN0P_  (.CLK(clknet_leaf_30_clk),
    .RESET_B(net472),
    .D(_00136_),
    .Q_N(_05591_),
    .Q(\dtop.player_inst.synth.alu.registers[2][3] ));
 sg13g2_dfrbp_1 \dtop.player_inst.synth.alu.registers[2][4]$_SDFFE_PN0P_  (.CLK(clknet_leaf_30_clk),
    .RESET_B(net473),
    .D(_00137_),
    .Q_N(_05590_),
    .Q(\dtop.player_inst.synth.alu.registers[2][4] ));
 sg13g2_dfrbp_1 \dtop.player_inst.synth.alu.registers[2][5]$_SDFFE_PN0P_  (.CLK(clknet_leaf_30_clk),
    .RESET_B(net474),
    .D(_00138_),
    .Q_N(_05589_),
    .Q(\dtop.player_inst.synth.alu.registers[2][5] ));
 sg13g2_dfrbp_1 \dtop.player_inst.synth.alu.registers[2][6]$_SDFFE_PN0P_  (.CLK(clknet_leaf_29_clk),
    .RESET_B(net475),
    .D(_00139_),
    .Q_N(_05588_),
    .Q(\dtop.player_inst.synth.alu.registers[2][6] ));
 sg13g2_dfrbp_1 \dtop.player_inst.synth.alu.registers[2][7]$_SDFFE_PN0P_  (.CLK(clknet_leaf_30_clk),
    .RESET_B(net476),
    .D(_00140_),
    .Q_N(_05587_),
    .Q(\dtop.player_inst.synth.alu.registers[2][7] ));
 sg13g2_dfrbp_1 \dtop.player_inst.synth.alu.registers[3][0]$_SDFFE_PN0P_  (.CLK(clknet_leaf_29_clk),
    .RESET_B(net477),
    .D(_00141_),
    .Q_N(_05586_),
    .Q(\dtop.player_inst.synth.alu.registers[3][0] ));
 sg13g2_dfrbp_1 \dtop.player_inst.synth.alu.registers[3][1]$_SDFFE_PN0P_  (.CLK(clknet_leaf_29_clk),
    .RESET_B(net478),
    .D(_00142_),
    .Q_N(_05585_),
    .Q(\dtop.player_inst.synth.alu.registers[3][1] ));
 sg13g2_dfrbp_1 \dtop.player_inst.synth.alu.registers[3][2]$_SDFFE_PN0P_  (.CLK(clknet_leaf_29_clk),
    .RESET_B(net479),
    .D(_00143_),
    .Q_N(_05584_),
    .Q(\dtop.player_inst.synth.alu.registers[3][2] ));
 sg13g2_dfrbp_1 \dtop.player_inst.synth.alu.registers[3][3]$_SDFFE_PN0P_  (.CLK(clknet_leaf_28_clk),
    .RESET_B(net480),
    .D(_00144_),
    .Q_N(_05583_),
    .Q(\dtop.player_inst.synth.alu.registers[3][3] ));
 sg13g2_dfrbp_1 \dtop.player_inst.synth.alu.registers[3][4]$_SDFFE_PN0P_  (.CLK(clknet_leaf_28_clk),
    .RESET_B(net481),
    .D(_00145_),
    .Q_N(_05582_),
    .Q(\dtop.player_inst.synth.alu.registers[3][4] ));
 sg13g2_dfrbp_1 \dtop.player_inst.synth.alu.registers[3][5]$_SDFFE_PN0P_  (.CLK(clknet_leaf_28_clk),
    .RESET_B(net482),
    .D(_00146_),
    .Q_N(_05581_),
    .Q(\dtop.player_inst.synth.alu.registers[3][5] ));
 sg13g2_dfrbp_1 \dtop.player_inst.synth.alu.registers[3][6]$_SDFFE_PN0P_  (.CLK(clknet_leaf_27_clk),
    .RESET_B(net483),
    .D(_00147_),
    .Q_N(_05580_),
    .Q(\dtop.player_inst.synth.alu.registers[3][6] ));
 sg13g2_dfrbp_1 \dtop.player_inst.synth.alu.registers[3][7]$_SDFFE_PN0P_  (.CLK(clknet_leaf_28_clk),
    .RESET_B(net484),
    .D(_00148_),
    .Q_N(_05579_),
    .Q(\dtop.player_inst.synth.alu.registers[3][7] ));
 sg13g2_dfrbp_1 \dtop.player_inst.synth.alu.registers[4][0]$_SDFFE_PN0P_  (.CLK(clknet_leaf_24_clk),
    .RESET_B(net485),
    .D(_00149_),
    .Q_N(_05578_),
    .Q(\dtop.player_inst.synth.alu.registers[4][0] ));
 sg13g2_dfrbp_1 \dtop.player_inst.synth.alu.registers[4][10]$_SDFFE_PN0P_  (.CLK(clknet_leaf_17_clk),
    .RESET_B(net486),
    .D(_00150_),
    .Q_N(_00076_),
    .Q(\dtop.player_inst.synth.alu.registers[4][10] ));
 sg13g2_dfrbp_1 \dtop.player_inst.synth.alu.registers[4][1]$_SDFFE_PN0P_  (.CLK(clknet_leaf_19_clk),
    .RESET_B(net487),
    .D(_00151_),
    .Q_N(_05577_),
    .Q(\dtop.player_inst.synth.alu.registers[4][1] ));
 sg13g2_dfrbp_1 \dtop.player_inst.synth.alu.registers[4][2]$_SDFFE_PN0P_  (.CLK(clknet_leaf_19_clk),
    .RESET_B(net488),
    .D(_00152_),
    .Q_N(_05576_),
    .Q(\dtop.player_inst.synth.alu.registers[4][2] ));
 sg13g2_dfrbp_1 \dtop.player_inst.synth.alu.registers[4][3]$_SDFFE_PN0P_  (.CLK(clknet_leaf_19_clk),
    .RESET_B(net489),
    .D(_00153_),
    .Q_N(_05575_),
    .Q(\dtop.player_inst.synth.alu.registers[4][3] ));
 sg13g2_dfrbp_1 \dtop.player_inst.synth.alu.registers[4][4]$_SDFFE_PN0P_  (.CLK(clknet_leaf_19_clk),
    .RESET_B(net490),
    .D(_00154_),
    .Q_N(_05574_),
    .Q(\dtop.player_inst.synth.alu.registers[4][4] ));
 sg13g2_dfrbp_1 \dtop.player_inst.synth.alu.registers[4][5]$_SDFFE_PN0P_  (.CLK(clknet_leaf_18_clk),
    .RESET_B(net491),
    .D(_00155_),
    .Q_N(_05573_),
    .Q(\dtop.player_inst.synth.alu.registers[4][5] ));
 sg13g2_dfrbp_1 \dtop.player_inst.synth.alu.registers[4][6]$_SDFFE_PN0P_  (.CLK(clknet_leaf_18_clk),
    .RESET_B(net492),
    .D(_00156_),
    .Q_N(_00071_),
    .Q(\dtop.player_inst.synth.alu.registers[4][6] ));
 sg13g2_dfrbp_1 \dtop.player_inst.synth.alu.registers[4][7]$_SDFFE_PN0P_  (.CLK(clknet_leaf_17_clk),
    .RESET_B(net493),
    .D(_00157_),
    .Q_N(_00072_),
    .Q(\dtop.player_inst.synth.alu.registers[4][7] ));
 sg13g2_dfrbp_1 \dtop.player_inst.synth.alu.registers[4][8]$_SDFFE_PN0P_  (.CLK(clknet_leaf_17_clk),
    .RESET_B(net494),
    .D(_00158_),
    .Q_N(_00073_),
    .Q(\dtop.player_inst.synth.alu.registers[4][8] ));
 sg13g2_dfrbp_1 \dtop.player_inst.synth.alu.registers[4][9]$_SDFFE_PN0P_  (.CLK(clknet_leaf_17_clk),
    .RESET_B(net495),
    .D(_00159_),
    .Q_N(_00075_),
    .Q(\dtop.player_inst.synth.alu.registers[4][9] ));
 sg13g2_dfrbp_1 \dtop.player_inst.synth.alu.registers[5][0]$_SDFFE_PN0P_  (.CLK(clknet_leaf_31_clk),
    .RESET_B(net496),
    .D(_00160_),
    .Q_N(_05572_),
    .Q(\dtop.player_inst.synth.alu.registers[5][0] ));
 sg13g2_dfrbp_1 \dtop.player_inst.synth.alu.registers[5][1]$_SDFFE_PN0P_  (.CLK(clknet_4_11_0_clk),
    .RESET_B(net497),
    .D(_00161_),
    .Q_N(_05571_),
    .Q(\dtop.player_inst.synth.alu.registers[5][1] ));
 sg13g2_dfrbp_1 \dtop.player_inst.synth.alu.registers[5][2]$_SDFFE_PN0P_  (.CLK(clknet_leaf_33_clk),
    .RESET_B(net498),
    .D(_00162_),
    .Q_N(_05570_),
    .Q(\dtop.player_inst.synth.alu.registers[5][2] ));
 sg13g2_dfrbp_1 \dtop.player_inst.synth.alu.registers[5][3]$_SDFFE_PN0P_  (.CLK(clknet_leaf_33_clk),
    .RESET_B(net499),
    .D(_00163_),
    .Q_N(_05569_),
    .Q(\dtop.player_inst.synth.alu.registers[5][3] ));
 sg13g2_dfrbp_1 \dtop.player_inst.synth.alu.registers[5][4]$_SDFFE_PN0P_  (.CLK(clknet_leaf_33_clk),
    .RESET_B(net500),
    .D(_00164_),
    .Q_N(_05568_),
    .Q(\dtop.player_inst.synth.alu.registers[5][4] ));
 sg13g2_dfrbp_1 \dtop.player_inst.synth.alu.registers[5][5]$_SDFFE_PN0P_  (.CLK(clknet_leaf_33_clk),
    .RESET_B(net501),
    .D(_00165_),
    .Q_N(_05567_),
    .Q(\dtop.player_inst.synth.alu.registers[5][5] ));
 sg13g2_dfrbp_1 \dtop.player_inst.synth.alu.registers[5][6]$_SDFFE_PN0P_  (.CLK(clknet_leaf_31_clk),
    .RESET_B(net502),
    .D(_00166_),
    .Q_N(_05566_),
    .Q(\dtop.player_inst.synth.alu.registers[5][6] ));
 sg13g2_dfrbp_1 \dtop.player_inst.synth.alu.registers[6][0]$_SDFFE_PN0P_  (.CLK(clknet_leaf_34_clk),
    .RESET_B(net503),
    .D(_00167_),
    .Q_N(_05565_),
    .Q(\dtop.out_sample[0] ));
 sg13g2_dfrbp_1 \dtop.player_inst.synth.alu.registers[6][1]$_SDFFE_PN0P_  (.CLK(clknet_leaf_34_clk),
    .RESET_B(net504),
    .D(_00168_),
    .Q_N(_05564_),
    .Q(\dtop.out_sample[1] ));
 sg13g2_dfrbp_1 \dtop.player_inst.synth.alu.registers[6][2]$_SDFFE_PN0P_  (.CLK(clknet_leaf_34_clk),
    .RESET_B(net505),
    .D(_00169_),
    .Q_N(_05563_),
    .Q(\dtop.out_sample[2] ));
 sg13g2_dfrbp_1 \dtop.player_inst.synth.alu.registers[6][3]$_SDFFE_PN0P_  (.CLK(clknet_leaf_33_clk),
    .RESET_B(net506),
    .D(_00170_),
    .Q_N(_05562_),
    .Q(\dtop.out_sample[3] ));
 sg13g2_dfrbp_1 \dtop.player_inst.synth.alu.registers[6][4]$_SDFFE_PN0P_  (.CLK(clknet_leaf_33_clk),
    .RESET_B(net507),
    .D(_00171_),
    .Q_N(_05561_),
    .Q(\dtop.out_sample[4] ));
 sg13g2_dfrbp_1 \dtop.player_inst.synth.alu.registers[6][5]$_SDFFE_PN0P_  (.CLK(clknet_leaf_33_clk),
    .RESET_B(net508),
    .D(_00172_),
    .Q_N(_05560_),
    .Q(\dtop.out_sample[5] ));
 sg13g2_dfrbp_1 \dtop.player_inst.synth.alu.registers[6][6]$_SDFFE_PN0P_  (.CLK(clknet_leaf_33_clk),
    .RESET_B(net509),
    .D(_00173_),
    .Q_N(_05559_),
    .Q(\dtop.out_sample[6] ));
 sg13g2_dfrbp_1 \dtop.vtop.dphases[0][0]$_DFFE_PP_  (.CLK(clknet_leaf_47_clk),
    .RESET_B(net510),
    .D(_00174_),
    .Q_N(_00032_),
    .Q(\dtop.vtop.dphases[0][0] ));
 sg13g2_dfrbp_1 \dtop.vtop.dphases[0][10]$_DFFE_PP_  (.CLK(clknet_leaf_49_clk),
    .RESET_B(net511),
    .D(_00175_),
    .Q_N(_00052_),
    .Q(\dtop.vtop.dphases[0][10] ));
 sg13g2_dfrbp_1 \dtop.vtop.dphases[0][1]$_DFFE_PP_  (.CLK(clknet_leaf_46_clk),
    .RESET_B(net512),
    .D(_00176_),
    .Q_N(_00034_),
    .Q(\dtop.vtop.dphases[0][1] ));
 sg13g2_dfrbp_1 \dtop.vtop.dphases[0][2]$_DFFE_PP_  (.CLK(clknet_leaf_46_clk),
    .RESET_B(net513),
    .D(_00177_),
    .Q_N(_00036_),
    .Q(\dtop.vtop.dphases[0][2] ));
 sg13g2_dfrbp_1 \dtop.vtop.dphases[0][3]$_DFFE_PP_  (.CLK(clknet_leaf_49_clk),
    .RESET_B(net514),
    .D(_00178_),
    .Q_N(_00038_),
    .Q(\dtop.vtop.dphases[0][3] ));
 sg13g2_dfrbp_1 \dtop.vtop.dphases[0][4]$_DFFE_PP_  (.CLK(clknet_leaf_50_clk),
    .RESET_B(net515),
    .D(_00179_),
    .Q_N(_00040_),
    .Q(\dtop.vtop.dphases[0][4] ));
 sg13g2_dfrbp_1 \dtop.vtop.dphases[0][5]$_DFFE_PP_  (.CLK(clknet_leaf_49_clk),
    .RESET_B(net516),
    .D(_00180_),
    .Q_N(_00042_),
    .Q(\dtop.vtop.dphases[0][5] ));
 sg13g2_dfrbp_1 \dtop.vtop.dphases[0][6]$_DFFE_PP_  (.CLK(clknet_leaf_50_clk),
    .RESET_B(net517),
    .D(_00181_),
    .Q_N(_00043_),
    .Q(\dtop.vtop.dphases[0][6] ));
 sg13g2_dfrbp_1 \dtop.vtop.dphases[0][7]$_DFFE_PP_  (.CLK(clknet_leaf_49_clk),
    .RESET_B(net518),
    .D(_00182_),
    .Q_N(_00045_),
    .Q(\dtop.vtop.dphases[0][7] ));
 sg13g2_dfrbp_1 \dtop.vtop.dphases[0][8]$_DFFE_PP_  (.CLK(clknet_leaf_48_clk),
    .RESET_B(net519),
    .D(_00183_),
    .Q_N(_00048_),
    .Q(\dtop.vtop.dphases[0][8] ));
 sg13g2_dfrbp_1 \dtop.vtop.dphases[0][9]$_DFFE_PP_  (.CLK(clknet_leaf_49_clk),
    .RESET_B(net520),
    .D(_00184_),
    .Q_N(_00050_),
    .Q(\dtop.vtop.dphases[0][9] ));
 sg13g2_dfrbp_1 \dtop.vtop.dphases[1][0]$_DFFE_PP_  (.CLK(clknet_leaf_47_clk),
    .RESET_B(net521),
    .D(_00185_),
    .Q_N(_05558_),
    .Q(\dtop.vtop.dphases[1][0] ));
 sg13g2_dfrbp_1 \dtop.vtop.dphases[1][10]$_DFFE_PP_  (.CLK(clknet_leaf_48_clk),
    .RESET_B(net522),
    .D(_00186_),
    .Q_N(_05557_),
    .Q(\dtop.vtop.dphases[1][10] ));
 sg13g2_dfrbp_1 \dtop.vtop.dphases[1][1]$_DFFE_PP_  (.CLK(clknet_leaf_46_clk),
    .RESET_B(net523),
    .D(_00187_),
    .Q_N(_05556_),
    .Q(\dtop.vtop.dphases[1][1] ));
 sg13g2_dfrbp_1 \dtop.vtop.dphases[1][2]$_DFFE_PP_  (.CLK(clknet_leaf_47_clk),
    .RESET_B(net524),
    .D(_00188_),
    .Q_N(_05555_),
    .Q(\dtop.vtop.dphases[1][2] ));
 sg13g2_dfrbp_1 \dtop.vtop.dphases[1][3]$_DFFE_PP_  (.CLK(clknet_leaf_53_clk),
    .RESET_B(net525),
    .D(_00189_),
    .Q_N(_05554_),
    .Q(\dtop.vtop.dphases[1][3] ));
 sg13g2_dfrbp_1 \dtop.vtop.dphases[1][4]$_DFFE_PP_  (.CLK(clknet_4_2_0_clk),
    .RESET_B(net526),
    .D(_00190_),
    .Q_N(_05553_),
    .Q(\dtop.vtop.dphases[1][4] ));
 sg13g2_dfrbp_1 \dtop.vtop.dphases[1][5]$_DFFE_PP_  (.CLK(clknet_leaf_52_clk),
    .RESET_B(net527),
    .D(_00191_),
    .Q_N(_05552_),
    .Q(\dtop.vtop.dphases[1][5] ));
 sg13g2_dfrbp_1 \dtop.vtop.dphases[1][6]$_DFFE_PP_  (.CLK(clknet_leaf_53_clk),
    .RESET_B(net528),
    .D(_00192_),
    .Q_N(_05551_),
    .Q(\dtop.vtop.dphases[1][6] ));
 sg13g2_dfrbp_1 \dtop.vtop.dphases[1][7]$_DFFE_PP_  (.CLK(clknet_leaf_53_clk),
    .RESET_B(net529),
    .D(_00193_),
    .Q_N(_05550_),
    .Q(\dtop.vtop.dphases[1][7] ));
 sg13g2_dfrbp_1 \dtop.vtop.dphases[1][8]$_DFFE_PP_  (.CLK(clknet_leaf_53_clk),
    .RESET_B(net530),
    .D(_00194_),
    .Q_N(_05549_),
    .Q(\dtop.vtop.dphases[1][8] ));
 sg13g2_dfrbp_1 \dtop.vtop.dphases[1][9]$_DFFE_PP_  (.CLK(clknet_leaf_48_clk),
    .RESET_B(net531),
    .D(_00195_),
    .Q_N(_05548_),
    .Q(\dtop.vtop.dphases[1][9] ));
 sg13g2_dfrbp_1 \dtop.vtop.dphases[2][0]$_DFFE_PP_  (.CLK(clknet_leaf_8_clk),
    .RESET_B(net532),
    .D(_00196_),
    .Q_N(_05547_),
    .Q(\dtop.vtop.dphases[2][0] ));
 sg13g2_dfrbp_1 \dtop.vtop.dphases[2][10]$_DFFE_PP_  (.CLK(clknet_leaf_47_clk),
    .RESET_B(net533),
    .D(_00197_),
    .Q_N(_05546_),
    .Q(\dtop.vtop.dphases[2][10] ));
 sg13g2_dfrbp_1 \dtop.vtop.dphases[2][1]$_DFFE_PP_  (.CLK(clknet_leaf_46_clk),
    .RESET_B(net534),
    .D(_00198_),
    .Q_N(_05545_),
    .Q(\dtop.vtop.dphases[2][1] ));
 sg13g2_dfrbp_1 \dtop.vtop.dphases[2][2]$_DFFE_PP_  (.CLK(clknet_leaf_46_clk),
    .RESET_B(net535),
    .D(_00199_),
    .Q_N(_05544_),
    .Q(\dtop.vtop.dphases[2][2] ));
 sg13g2_dfrbp_1 \dtop.vtop.dphases[2][3]$_DFFE_PP_  (.CLK(clknet_leaf_49_clk),
    .RESET_B(net536),
    .D(_00200_),
    .Q_N(_05543_),
    .Q(\dtop.vtop.dphases[2][3] ));
 sg13g2_dfrbp_1 \dtop.vtop.dphases[2][4]$_DFFE_PP_  (.CLK(clknet_leaf_50_clk),
    .RESET_B(net537),
    .D(_00201_),
    .Q_N(_05542_),
    .Q(\dtop.vtop.dphases[2][4] ));
 sg13g2_dfrbp_1 \dtop.vtop.dphases[2][5]$_DFFE_PP_  (.CLK(clknet_leaf_49_clk),
    .RESET_B(net538),
    .D(_00202_),
    .Q_N(_05541_),
    .Q(\dtop.vtop.dphases[2][5] ));
 sg13g2_dfrbp_1 \dtop.vtop.dphases[2][6]$_DFFE_PP_  (.CLK(clknet_leaf_53_clk),
    .RESET_B(net539),
    .D(_00203_),
    .Q_N(_05540_),
    .Q(\dtop.vtop.dphases[2][6] ));
 sg13g2_dfrbp_1 \dtop.vtop.dphases[2][7]$_DFFE_PP_  (.CLK(clknet_leaf_53_clk),
    .RESET_B(net540),
    .D(_00204_),
    .Q_N(_05539_),
    .Q(\dtop.vtop.dphases[2][7] ));
 sg13g2_dfrbp_1 \dtop.vtop.dphases[2][8]$_DFFE_PP_  (.CLK(clknet_leaf_48_clk),
    .RESET_B(net541),
    .D(_00205_),
    .Q_N(_05538_),
    .Q(\dtop.vtop.dphases[2][8] ));
 sg13g2_dfrbp_1 \dtop.vtop.dphases[2][9]$_DFFE_PP_  (.CLK(clknet_leaf_48_clk),
    .RESET_B(net542),
    .D(_00206_),
    .Q_N(_05537_),
    .Q(\dtop.vtop.dphases[2][9] ));
 sg13g2_dfrbp_1 \dtop.vtop.pipeline.cosappr[3]$_DFFE_PP_  (.CLK(clknet_leaf_7_clk),
    .RESET_B(net543),
    .D(_00207_),
    .Q_N(_00011_),
    .Q(\dtop.vtop.color[6] ));
 sg13g2_dfrbp_1 \dtop.vtop.pipeline.cosappr[4]$_DFFE_PP_  (.CLK(clknet_leaf_7_clk),
    .RESET_B(net544),
    .D(_00208_),
    .Q_N(_00010_),
    .Q(\dtop.vtop.color[7] ));
 sg13g2_dfrbp_1 \dtop.vtop.pipeline.cosappr[5]$_DFFE_PP_  (.CLK(clknet_leaf_7_clk),
    .RESET_B(net545),
    .D(_00209_),
    .Q_N(_00013_),
    .Q(\dtop.vtop.color[8] ));
 sg13g2_dfrbp_1 \dtop.vtop.pipeline.cosappr[6]$_DFFE_PP_  (.CLK(clknet_leaf_6_clk),
    .RESET_B(net546),
    .D(_00210_),
    .Q_N(_00009_),
    .Q(\dtop.vtop.color[9] ));
 sg13g2_dfrbp_1 \dtop.vtop.pipeline.cosappr[7]$_DFFE_PP_  (.CLK(clknet_leaf_7_clk),
    .RESET_B(net547),
    .D(_00211_),
    .Q_N(_00008_),
    .Q(\dtop.vtop.color[10] ));
 sg13g2_dfrbp_1 \dtop.vtop.pipeline.cosappr[8]$_DFFE_PP_  (.CLK(clknet_leaf_6_clk),
    .RESET_B(net548),
    .D(_00212_),
    .Q_N(_00007_),
    .Q(\dtop.vtop.color[11] ));
 sg13g2_dfrbp_1 \dtop.vtop.pipeline.cosappr_acc[0]$_DFFE_PN_  (.CLK(clknet_leaf_56_clk),
    .RESET_B(net549),
    .D(_00213_),
    .Q_N(_05536_),
    .Q(\dtop.vtop.pipeline.cosappr_acc[0] ));
 sg13g2_dfrbp_1 \dtop.vtop.pipeline.cosappr_acc[1]$_DFFE_PN_  (.CLK(clknet_leaf_56_clk),
    .RESET_B(net550),
    .D(_00214_),
    .Q_N(_05535_),
    .Q(\dtop.vtop.pipeline.cosappr_acc[1] ));
 sg13g2_dfrbp_1 \dtop.vtop.pipeline.cosappr_acc[2]$_DFFE_PN_  (.CLK(clknet_leaf_56_clk),
    .RESET_B(net551),
    .D(_00215_),
    .Q_N(_05534_),
    .Q(\dtop.vtop.pipeline.cosappr_acc[2] ));
 sg13g2_dfrbp_1 \dtop.vtop.pipeline.cosappr_acc[3]$_DFFE_PN_  (.CLK(clknet_leaf_52_clk),
    .RESET_B(net552),
    .D(_00216_),
    .Q_N(_05533_),
    .Q(\dtop.vtop.pipeline.cosappr_acc[3] ));
 sg13g2_dfrbp_1 \dtop.vtop.pipeline.cosappr_acc[4]$_DFFE_PN_  (.CLK(clknet_leaf_52_clk),
    .RESET_B(net553),
    .D(_00217_),
    .Q_N(_05532_),
    .Q(\dtop.vtop.pipeline.cosappr_acc[4] ));
 sg13g2_dfrbp_1 \dtop.vtop.pipeline.cosappr_acc[5]$_DFFE_PN_  (.CLK(clknet_leaf_51_clk),
    .RESET_B(net554),
    .D(_00218_),
    .Q_N(_05531_),
    .Q(\dtop.vtop.pipeline.cosappr_acc[5] ));
 sg13g2_dfrbp_1 \dtop.vtop.pipeline.cosappr_acc[6]$_DFFE_PN_  (.CLK(clknet_leaf_51_clk),
    .RESET_B(net555),
    .D(_00219_),
    .Q_N(_05530_),
    .Q(\dtop.vtop.pipeline.cosappr_acc[6] ));
 sg13g2_dfrbp_1 \dtop.vtop.pipeline.cosappr_acc[7]$_DFFE_PN_  (.CLK(clknet_leaf_56_clk),
    .RESET_B(net556),
    .D(_00220_),
    .Q_N(_05529_),
    .Q(\dtop.vtop.pipeline.cosappr_acc[7] ));
 sg13g2_dfrbp_1 \dtop.vtop.pipeline.cosappr_acc[8]$_DFFE_PN_  (.CLK(clknet_leaf_56_clk),
    .RESET_B(net557),
    .D(_00221_),
    .Q_N(_05528_),
    .Q(\dtop.vtop.pipeline.cosappr_acc[8] ));
 sg13g2_dfrbp_1 \dtop.vtop.pipeline.dz[0]$_SDFFE_PP1P_  (.CLK(clknet_leaf_3_clk),
    .RESET_B(net558),
    .D(_00222_),
    .Q_N(_00088_),
    .Q(\dtop.vtop.pipeline.dz[0] ));
 sg13g2_dfrbp_1 \dtop.vtop.pipeline.dz[1]$_SDFFE_PP1P_  (.CLK(clknet_leaf_6_clk),
    .RESET_B(net559),
    .D(_00223_),
    .Q_N(_00067_),
    .Q(\dtop.vtop.pipeline.dz[1] ));
 sg13g2_dfrbp_1 \dtop.vtop.pipeline.dz[2]$_SDFFE_PP1P_  (.CLK(clknet_leaf_6_clk),
    .RESET_B(net560),
    .D(_00224_),
    .Q_N(_00095_),
    .Q(\dtop.vtop.pipeline.dz[2] ));
 sg13g2_dfrbp_1 \dtop.vtop.pipeline.dz[3]$_SDFFE_PP1P_  (.CLK(clknet_leaf_12_clk),
    .RESET_B(net561),
    .D(_00225_),
    .Q_N(_00068_),
    .Q(\dtop.vtop.pipeline.dz[3] ));
 sg13g2_dfrbp_1 \dtop.vtop.pipeline.dz[4]$_SDFFE_PP1P_  (.CLK(clknet_leaf_12_clk),
    .RESET_B(net562),
    .D(_00226_),
    .Q_N(_00094_),
    .Q(\dtop.vtop.pipeline.dz[4] ));
 sg13g2_dfrbp_1 \dtop.vtop.pipeline.dz[5]$_SDFFE_PP1P_  (.CLK(clknet_leaf_12_clk),
    .RESET_B(net563),
    .D(_00227_),
    .Q_N(_00070_),
    .Q(\dtop.vtop.pipeline.dz[5] ));
 sg13g2_dfrbp_1 \dtop.vtop.pipeline.dz[6]$_SDFFE_PP1P_  (.CLK(clknet_leaf_5_clk),
    .RESET_B(net564),
    .D(_00228_),
    .Q_N(_00093_),
    .Q(\dtop.vtop.pipeline.dz[6] ));
 sg13g2_dfrbp_1 \dtop.vtop.pipeline.dz[7]$_SDFFE_PP1P_  (.CLK(clknet_leaf_12_clk),
    .RESET_B(net565),
    .D(_00229_),
    .Q_N(_00092_),
    .Q(\dtop.vtop.pipeline.dz[7] ));
 sg13g2_dfrbp_1 \dtop.vtop.pipeline.dz[8]$_SDFFE_PP1P_  (.CLK(clknet_leaf_4_clk),
    .RESET_B(net566),
    .D(_00230_),
    .Q_N(_00091_),
    .Q(\dtop.vtop.pipeline.dz[8] ));
 sg13g2_dfrbp_1 \dtop.vtop.pipeline.neg_t[0]$_SDFFE_PP0P_  (.CLK(clknet_leaf_6_clk),
    .RESET_B(net567),
    .D(_00231_),
    .Q_N(_00087_),
    .Q(\dtop.vtop.pipeline.neg_t[0] ));
 sg13g2_dfrbp_1 \dtop.vtop.pipeline.neg_t[1]$_SDFFE_PP0P_  (.CLK(clknet_leaf_6_clk),
    .RESET_B(net568),
    .D(_00232_),
    .Q_N(_00015_),
    .Q(\dtop.vtop.pipeline.neg_t[1] ));
 sg13g2_dfrbp_1 \dtop.vtop.pipeline.neg_t[2]$_SDFFE_PP0P_  (.CLK(clknet_leaf_5_clk),
    .RESET_B(net569),
    .D(_00233_),
    .Q_N(_00018_),
    .Q(\dtop.vtop.pipeline.neg_t[2] ));
 sg13g2_dfrbp_1 \dtop.vtop.pipeline.neg_t[3]$_SDFFE_PP0P_  (.CLK(clknet_leaf_5_clk),
    .RESET_B(net570),
    .D(_00234_),
    .Q_N(_00016_),
    .Q(\dtop.vtop.pipeline.neg_t[3] ));
 sg13g2_dfrbp_1 \dtop.vtop.pipeline.neg_t[4]$_SDFFE_PP0P_  (.CLK(clknet_leaf_12_clk),
    .RESET_B(net571),
    .D(_00235_),
    .Q_N(_00021_),
    .Q(\dtop.vtop.pipeline.neg_t[4] ));
 sg13g2_dfrbp_1 \dtop.vtop.pipeline.neg_t[5]$_SDFFE_PP0P_  (.CLK(clknet_leaf_5_clk),
    .RESET_B(net572),
    .D(_00236_),
    .Q_N(_00069_),
    .Q(\dtop.vtop.pipeline.neg_t[5] ));
 sg13g2_dfrbp_1 \dtop.vtop.pipeline.neg_t[6]$_SDFFE_PP0P_  (.CLK(clknet_leaf_5_clk),
    .RESET_B(net573),
    .D(_00237_),
    .Q_N(_00023_),
    .Q(\dtop.vtop.pipeline.neg_t[6] ));
 sg13g2_dfrbp_1 \dtop.vtop.pipeline.neg_t[7]$_SDFFE_PP0P_  (.CLK(clknet_leaf_12_clk),
    .RESET_B(net574),
    .D(_00238_),
    .Q_N(_00025_),
    .Q(\dtop.vtop.pipeline.neg_t[7] ));
 sg13g2_dfrbp_1 \dtop.vtop.pipeline.neg_t[8]$_SDFFE_PP0P_  (.CLK(clknet_leaf_4_clk),
    .RESET_B(net575),
    .D(_00239_),
    .Q_N(_00027_),
    .Q(\dtop.vtop.pipeline.neg_t[8] ));
 sg13g2_dfrbp_1 \dtop.vtop.pipeline.neg_t[9]$_SDFFE_PP0P_  (.CLK(clknet_leaf_4_clk),
    .RESET_B(net576),
    .D(_00240_),
    .Q_N(_00026_),
    .Q(\dtop.vtop.pipeline.neg_t[9] ));
 sg13g2_dfrbp_1 \dtop.vtop.pipeline.nstep_counter[0]$_SDFFE_PP1P_  (.CLK(clknet_leaf_3_clk),
    .RESET_B(net577),
    .D(_00241_),
    .Q_N(\dtop.vtop.pipeline.next_nstep_counter[0] ),
    .Q(\dtop.vtop.pipeline.nstep_counter[0] ));
 sg13g2_dfrbp_1 \dtop.vtop.pipeline.nstep_counter[1]$_SDFFE_PP1P_  (.CLK(clknet_leaf_7_clk),
    .RESET_B(net578),
    .D(_00242_),
    .Q_N(_05527_),
    .Q(\dtop.vtop.pipeline.nstep_counter[1] ));
 sg13g2_dfrbp_1 \dtop.vtop.pipeline.nstep_counter[2]$_SDFFE_PP1P_  (.CLK(clknet_leaf_8_clk),
    .RESET_B(net579),
    .D(_00243_),
    .Q_N(_05526_),
    .Q(\dtop.vtop.pipeline.nstep_counter[2] ));
 sg13g2_dfrbp_1 \dtop.vtop.pipeline.nstep_counter[3]$_SDFFE_PP1P_  (.CLK(clknet_leaf_8_clk),
    .RESET_B(net580),
    .D(_00244_),
    .Q_N(_05525_),
    .Q(\dtop.vtop.pipeline.nstep_counter[3] ));
 sg13g2_dfrbp_1 \dtop.vtop.pipeline.nstep_counter[4]$_SDFFE_PP1P_  (.CLK(clknet_leaf_8_clk),
    .RESET_B(net581),
    .D(_00245_),
    .Q_N(_05524_),
    .Q(\dtop.vtop.pipeline.nstep_counter[4] ));
 sg13g2_dfrbp_1 \dtop.vtop.pipeline.nstep_reg[0]$_SDFF_PP0_  (.CLK(clknet_leaf_47_clk),
    .RESET_B(net582),
    .D(_00246_),
    .Q_N(_05523_),
    .Q(\dtop.vtop.pipeline.nstep[0] ));
 sg13g2_dfrbp_1 \dtop.vtop.pipeline.nstep_reg[1]$_SDFF_PP0_  (.CLK(clknet_leaf_8_clk),
    .RESET_B(net583),
    .D(_00247_),
    .Q_N(_00031_),
    .Q(\dtop.vtop.pipeline.nstep[1] ));
 sg13g2_dfrbp_1 \dtop.vtop.pipeline.nstep_zg[0]$_DFFE_PP_  (.CLK(clknet_leaf_7_clk),
    .RESET_B(net584),
    .D(_00248_),
    .Q_N(_05522_),
    .Q(\dtop.vtop.pipeline.nstep_zg[0] ));
 sg13g2_dfrbp_1 \dtop.vtop.pipeline.nstep_zg[1]$_DFFE_PP_  (.CLK(clknet_leaf_3_clk),
    .RESET_B(net585),
    .D(_00249_),
    .Q_N(_05521_),
    .Q(\dtop.vtop.pipeline.nstep_zg[1] ));
 sg13g2_dfrbp_1 \dtop.vtop.pipeline.phases[0][0]$_DFFE_PP_  (.CLK(clknet_leaf_45_clk),
    .RESET_B(net586),
    .D(_00250_),
    .Q_N(_00030_),
    .Q(\dtop.vtop.pipeline.phases[0][0] ));
 sg13g2_dfrbp_1 \dtop.vtop.pipeline.phases[0][10]$_DFFE_PP_  (.CLK(clknet_leaf_42_clk),
    .RESET_B(net587),
    .D(_00251_),
    .Q_N(_00051_),
    .Q(\dtop.vtop.pipeline.phases[0][10] ));
 sg13g2_dfrbp_1 \dtop.vtop.pipeline.phases[0][11]$_DFFE_PP_  (.CLK(clknet_leaf_42_clk),
    .RESET_B(net588),
    .D(_00252_),
    .Q_N(_00053_),
    .Q(\dtop.vtop.pipeline.phases[0][11] ));
 sg13g2_dfrbp_1 \dtop.vtop.pipeline.phases[0][12]$_DFFE_PP_  (.CLK(clknet_leaf_42_clk),
    .RESET_B(net589),
    .D(_00253_),
    .Q_N(_00054_),
    .Q(\dtop.vtop.pipeline.phases[0][12] ));
 sg13g2_dfrbp_1 \dtop.vtop.pipeline.phases[0][13]$_DFFE_PP_  (.CLK(clknet_leaf_44_clk),
    .RESET_B(net590),
    .D(_00254_),
    .Q_N(_00055_),
    .Q(\dtop.vtop.pipeline.phases[0][13] ));
 sg13g2_dfrbp_1 \dtop.vtop.pipeline.phases[0][14]$_DFFE_PP_  (.CLK(clknet_leaf_39_clk),
    .RESET_B(net591),
    .D(_00255_),
    .Q_N(_00057_),
    .Q(\dtop.vtop.pipeline.phases[0][14] ));
 sg13g2_dfrbp_1 \dtop.vtop.pipeline.phases[0][15]$_DFFE_PP_  (.CLK(clknet_leaf_44_clk),
    .RESET_B(net592),
    .D(_00256_),
    .Q_N(_00003_),
    .Q(\dtop.vtop.pipeline.phases[0][15] ));
 sg13g2_dfrbp_1 \dtop.vtop.pipeline.phases[0][1]$_DFFE_PP_  (.CLK(clknet_leaf_37_clk),
    .RESET_B(net593),
    .D(_00257_),
    .Q_N(_00033_),
    .Q(\dtop.vtop.pipeline.phases[0][1] ));
 sg13g2_dfrbp_1 \dtop.vtop.pipeline.phases[0][2]$_DFFE_PP_  (.CLK(clknet_leaf_39_clk),
    .RESET_B(net594),
    .D(_00258_),
    .Q_N(_00035_),
    .Q(\dtop.vtop.pipeline.phases[0][2] ));
 sg13g2_dfrbp_1 \dtop.vtop.pipeline.phases[0][3]$_DFFE_PP_  (.CLK(clknet_leaf_45_clk),
    .RESET_B(net595),
    .D(_00259_),
    .Q_N(_00037_),
    .Q(\dtop.vtop.pipeline.phases[0][3] ));
 sg13g2_dfrbp_1 \dtop.vtop.pipeline.phases[0][4]$_DFFE_PP_  (.CLK(clknet_leaf_36_clk),
    .RESET_B(net596),
    .D(_00260_),
    .Q_N(_00039_),
    .Q(\dtop.vtop.pipeline.phases[0][4] ));
 sg13g2_dfrbp_1 \dtop.vtop.pipeline.phases[0][5]$_DFFE_PP_  (.CLK(clknet_leaf_39_clk),
    .RESET_B(net597),
    .D(_00261_),
    .Q_N(_00041_),
    .Q(\dtop.vtop.pipeline.phases[0][5] ));
 sg13g2_dfrbp_1 \dtop.vtop.pipeline.phases[0][6]$_DFFE_PP_  (.CLK(clknet_leaf_38_clk),
    .RESET_B(net598),
    .D(_00262_),
    .Q_N(_05520_),
    .Q(\dtop.vtop.pipeline.phases[0][6] ));
 sg13g2_dfrbp_1 \dtop.vtop.pipeline.phases[0][7]$_DFFE_PP_  (.CLK(clknet_leaf_39_clk),
    .RESET_B(net599),
    .D(_00263_),
    .Q_N(_00044_),
    .Q(\dtop.vtop.pipeline.phases[0][7] ));
 sg13g2_dfrbp_1 \dtop.vtop.pipeline.phases[0][8]$_DFFE_PP_  (.CLK(clknet_leaf_37_clk),
    .RESET_B(net600),
    .D(_00264_),
    .Q_N(_00046_),
    .Q(\dtop.vtop.pipeline.phases[0][8] ));
 sg13g2_dfrbp_1 \dtop.vtop.pipeline.phases[0][9]$_DFFE_PP_  (.CLK(clknet_leaf_42_clk),
    .RESET_B(net601),
    .D(_00265_),
    .Q_N(_00049_),
    .Q(\dtop.vtop.pipeline.phases[0][9] ));
 sg13g2_dfrbp_1 \dtop.vtop.pipeline.phases[1][0]$_DFFE_PP_  (.CLK(clknet_leaf_45_clk),
    .RESET_B(net602),
    .D(_00266_),
    .Q_N(_05519_),
    .Q(\dtop.vtop.pipeline.phases[1][0] ));
 sg13g2_dfrbp_1 \dtop.vtop.pipeline.phases[1][10]$_DFFE_PP_  (.CLK(clknet_leaf_39_clk),
    .RESET_B(net603),
    .D(_00267_),
    .Q_N(_05518_),
    .Q(\dtop.vtop.pipeline.phases[1][10] ));
 sg13g2_dfrbp_1 \dtop.vtop.pipeline.phases[1][11]$_DFFE_PP_  (.CLK(clknet_leaf_39_clk),
    .RESET_B(net604),
    .D(_00268_),
    .Q_N(_05517_),
    .Q(\dtop.vtop.pipeline.phases[1][11] ));
 sg13g2_dfrbp_1 \dtop.vtop.pipeline.phases[1][12]$_DFFE_PP_  (.CLK(clknet_leaf_44_clk),
    .RESET_B(net605),
    .D(_00269_),
    .Q_N(_05516_),
    .Q(\dtop.vtop.pipeline.phases[1][12] ));
 sg13g2_dfrbp_1 \dtop.vtop.pipeline.phases[1][13]$_DFFE_PP_  (.CLK(clknet_leaf_44_clk),
    .RESET_B(net606),
    .D(_00270_),
    .Q_N(_05515_),
    .Q(\dtop.vtop.pipeline.phases[1][13] ));
 sg13g2_dfrbp_1 \dtop.vtop.pipeline.phases[1][14]$_DFFE_PP_  (.CLK(clknet_leaf_40_clk),
    .RESET_B(net607),
    .D(_00271_),
    .Q_N(_05514_),
    .Q(\dtop.vtop.pipeline.phases[1][14] ));
 sg13g2_dfrbp_1 \dtop.vtop.pipeline.phases[1][15]$_DFFE_PP_  (.CLK(clknet_leaf_44_clk),
    .RESET_B(net608),
    .D(_00272_),
    .Q_N(_05513_),
    .Q(\dtop.vtop.pipeline.phases[1][15] ));
 sg13g2_dfrbp_1 \dtop.vtop.pipeline.phases[1][1]$_DFFE_PP_  (.CLK(clknet_leaf_37_clk),
    .RESET_B(net609),
    .D(_00273_),
    .Q_N(_05512_),
    .Q(\dtop.vtop.pipeline.phases[1][1] ));
 sg13g2_dfrbp_1 \dtop.vtop.pipeline.phases[1][2]$_DFFE_PP_  (.CLK(clknet_leaf_39_clk),
    .RESET_B(net610),
    .D(_00274_),
    .Q_N(_05511_),
    .Q(\dtop.vtop.pipeline.phases[1][2] ));
 sg13g2_dfrbp_1 \dtop.vtop.pipeline.phases[1][3]$_DFFE_PP_  (.CLK(clknet_leaf_36_clk),
    .RESET_B(net611),
    .D(_00275_),
    .Q_N(_05510_),
    .Q(\dtop.vtop.pipeline.phases[1][3] ));
 sg13g2_dfrbp_1 \dtop.vtop.pipeline.phases[1][4]$_DFFE_PP_  (.CLK(clknet_leaf_37_clk),
    .RESET_B(net612),
    .D(_00276_),
    .Q_N(_05509_),
    .Q(\dtop.vtop.pipeline.phases[1][4] ));
 sg13g2_dfrbp_1 \dtop.vtop.pipeline.phases[1][5]$_DFFE_PP_  (.CLK(clknet_leaf_40_clk),
    .RESET_B(net613),
    .D(_00277_),
    .Q_N(_05508_),
    .Q(\dtop.vtop.pipeline.phases[1][5] ));
 sg13g2_dfrbp_1 \dtop.vtop.pipeline.phases[1][6]$_DFFE_PP_  (.CLK(clknet_leaf_38_clk),
    .RESET_B(net614),
    .D(_00278_),
    .Q_N(_05507_),
    .Q(\dtop.vtop.pipeline.phases[1][6] ));
 sg13g2_dfrbp_1 \dtop.vtop.pipeline.phases[1][7]$_DFFE_PP_  (.CLK(clknet_leaf_38_clk),
    .RESET_B(net615),
    .D(_00279_),
    .Q_N(_05506_),
    .Q(\dtop.vtop.pipeline.phases[1][7] ));
 sg13g2_dfrbp_1 \dtop.vtop.pipeline.phases[1][8]$_DFFE_PP_  (.CLK(clknet_leaf_37_clk),
    .RESET_B(net616),
    .D(_00280_),
    .Q_N(_05505_),
    .Q(\dtop.vtop.pipeline.phases[1][8] ));
 sg13g2_dfrbp_1 \dtop.vtop.pipeline.phases[1][9]$_DFFE_PP_  (.CLK(clknet_leaf_44_clk),
    .RESET_B(net617),
    .D(_00281_),
    .Q_N(_05504_),
    .Q(\dtop.vtop.pipeline.phases[1][9] ));
 sg13g2_dfrbp_1 \dtop.vtop.pipeline.phases[2][0]$_DFFE_PP_  (.CLK(clknet_leaf_45_clk),
    .RESET_B(net618),
    .D(_00282_),
    .Q_N(_05503_),
    .Q(\dtop.vtop.pipeline.phases[2][0] ));
 sg13g2_dfrbp_1 \dtop.vtop.pipeline.phases[2][10]$_DFFE_PP_  (.CLK(clknet_leaf_41_clk),
    .RESET_B(net619),
    .D(_00283_),
    .Q_N(_05502_),
    .Q(\dtop.vtop.pipeline.phases[2][10] ));
 sg13g2_dfrbp_1 \dtop.vtop.pipeline.phases[2][11]$_DFFE_PP_  (.CLK(clknet_leaf_42_clk),
    .RESET_B(net620),
    .D(_00284_),
    .Q_N(_05501_),
    .Q(\dtop.vtop.pipeline.phases[2][11] ));
 sg13g2_dfrbp_1 \dtop.vtop.pipeline.phases[2][12]$_DFFE_PP_  (.CLK(clknet_leaf_41_clk),
    .RESET_B(net621),
    .D(_00285_),
    .Q_N(_05500_),
    .Q(\dtop.vtop.pipeline.phases[2][12] ));
 sg13g2_dfrbp_1 \dtop.vtop.pipeline.phases[2][13]$_DFFE_PP_  (.CLK(clknet_leaf_44_clk),
    .RESET_B(net622),
    .D(_00286_),
    .Q_N(_05499_),
    .Q(\dtop.vtop.pipeline.phases[2][13] ));
 sg13g2_dfrbp_1 \dtop.vtop.pipeline.phases[2][14]$_DFFE_PP_  (.CLK(clknet_leaf_39_clk),
    .RESET_B(net623),
    .D(_00287_),
    .Q_N(_05498_),
    .Q(\dtop.vtop.pipeline.phases[2][14] ));
 sg13g2_dfrbp_1 \dtop.vtop.pipeline.phases[2][15]$_DFFE_PP_  (.CLK(clknet_leaf_44_clk),
    .RESET_B(net624),
    .D(_00288_),
    .Q_N(_05497_),
    .Q(\dtop.vtop.pipeline.phases[2][15] ));
 sg13g2_dfrbp_1 \dtop.vtop.pipeline.phases[2][1]$_DFFE_PP_  (.CLK(clknet_leaf_37_clk),
    .RESET_B(net625),
    .D(_00289_),
    .Q_N(_05496_),
    .Q(\dtop.vtop.pipeline.phases[2][1] ));
 sg13g2_dfrbp_1 \dtop.vtop.pipeline.phases[2][2]$_DFFE_PP_  (.CLK(clknet_leaf_40_clk),
    .RESET_B(net626),
    .D(_00290_),
    .Q_N(_05495_),
    .Q(\dtop.vtop.pipeline.phases[2][2] ));
 sg13g2_dfrbp_1 \dtop.vtop.pipeline.phases[2][3]$_DFFE_PP_  (.CLK(clknet_leaf_45_clk),
    .RESET_B(net627),
    .D(_00291_),
    .Q_N(_05494_),
    .Q(\dtop.vtop.pipeline.phases[2][3] ));
 sg13g2_dfrbp_1 \dtop.vtop.pipeline.phases[2][4]$_DFFE_PP_  (.CLK(clknet_leaf_36_clk),
    .RESET_B(net628),
    .D(_00292_),
    .Q_N(_05493_),
    .Q(\dtop.vtop.pipeline.phases[2][4] ));
 sg13g2_dfrbp_1 \dtop.vtop.pipeline.phases[2][5]$_DFFE_PP_  (.CLK(clknet_leaf_40_clk),
    .RESET_B(net629),
    .D(_00293_),
    .Q_N(_05492_),
    .Q(\dtop.vtop.pipeline.phases[2][5] ));
 sg13g2_dfrbp_1 \dtop.vtop.pipeline.phases[2][6]$_DFFE_PP_  (.CLK(clknet_leaf_38_clk),
    .RESET_B(net630),
    .D(_00294_),
    .Q_N(_05491_),
    .Q(\dtop.vtop.pipeline.phases[2][6] ));
 sg13g2_dfrbp_1 \dtop.vtop.pipeline.phases[2][7]$_DFFE_PP_  (.CLK(clknet_leaf_42_clk),
    .RESET_B(net631),
    .D(_00295_),
    .Q_N(_05490_),
    .Q(\dtop.vtop.pipeline.phases[2][7] ));
 sg13g2_dfrbp_1 \dtop.vtop.pipeline.phases[2][8]$_DFFE_PP_  (.CLK(clknet_leaf_38_clk),
    .RESET_B(net632),
    .D(_00296_),
    .Q_N(_05489_),
    .Q(\dtop.vtop.pipeline.phases[2][8] ));
 sg13g2_dfrbp_1 \dtop.vtop.pipeline.phases[2][9]$_DFFE_PP_  (.CLK(clknet_leaf_42_clk),
    .RESET_B(net633),
    .D(_00297_),
    .Q_N(_05488_),
    .Q(\dtop.vtop.pipeline.phases[2][9] ));
 sg13g2_dfrbp_1 \dtop.vtop.pipeline.wave_index[0]$_SDFF_PP0_  (.CLK(clknet_leaf_7_clk),
    .RESET_B(net634),
    .D(_00298_),
    .Q_N(_00004_),
    .Q(\dtop.vtop.pipeline.wave_index[0] ));
 sg13g2_dfrbp_1 \dtop.vtop.pipeline.wave_index[1]$_SDFF_PP0_  (.CLK(clknet_leaf_47_clk),
    .RESET_B(net635),
    .D(_00299_),
    .Q_N(_00006_),
    .Q(\dtop.vtop.pipeline.wave_index[1] ));
 sg13g2_dfrbp_1 \dtop.vtop.pipeline.z[0]$_SDFFE_PP0P_  (.CLK(clknet_leaf_3_clk),
    .RESET_B(net636),
    .D(_00300_),
    .Q_N(_05487_),
    .Q(\dtop.vtop.pipeline.z[0] ));
 sg13g2_dfrbp_1 \dtop.vtop.pipeline.z[10]$_SDFFE_PP0P_  (.CLK(clknet_leaf_1_clk),
    .RESET_B(net637),
    .D(_00301_),
    .Q_N(_05486_),
    .Q(\dtop.vtop.pipeline.z[10] ));
 sg13g2_dfrbp_1 \dtop.vtop.pipeline.z[11]$_SDFFE_PP0P_  (.CLK(clknet_leaf_1_clk),
    .RESET_B(net638),
    .D(_00302_),
    .Q_N(_05485_),
    .Q(\dtop.vtop.pipeline.z[11] ));
 sg13g2_dfrbp_1 \dtop.vtop.pipeline.z[12]$_SDFFE_PP0P_  (.CLK(clknet_leaf_2_clk),
    .RESET_B(net639),
    .D(_00303_),
    .Q_N(_05484_),
    .Q(\dtop.vtop.pipeline.z[12] ));
 sg13g2_dfrbp_1 \dtop.vtop.pipeline.z[13]$_SDFFE_PP0P_  (.CLK(clknet_leaf_2_clk),
    .RESET_B(net640),
    .D(_00304_),
    .Q_N(_05483_),
    .Q(\dtop.vtop.pipeline.z[13] ));
 sg13g2_dfrbp_1 \dtop.vtop.pipeline.z[14]$_SDFFE_PP0P_  (.CLK(clknet_leaf_3_clk),
    .RESET_B(net641),
    .D(_00305_),
    .Q_N(_05482_),
    .Q(\dtop.vtop.pipeline.z[14] ));
 sg13g2_dfrbp_1 \dtop.vtop.pipeline.z[1]$_SDFFE_PP0P_  (.CLK(clknet_leaf_4_clk),
    .RESET_B(net642),
    .D(_00306_),
    .Q_N(_05481_),
    .Q(\dtop.vtop.pipeline.z[1] ));
 sg13g2_dfrbp_1 \dtop.vtop.pipeline.z[2]$_SDFFE_PP0P_  (.CLK(clknet_leaf_4_clk),
    .RESET_B(net643),
    .D(_00307_),
    .Q_N(_05480_),
    .Q(\dtop.vtop.pipeline.z[2] ));
 sg13g2_dfrbp_1 \dtop.vtop.pipeline.z[3]$_SDFFE_PP0P_  (.CLK(clknet_leaf_1_clk),
    .RESET_B(net644),
    .D(_00308_),
    .Q_N(_05479_),
    .Q(\dtop.vtop.pipeline.z[3] ));
 sg13g2_dfrbp_1 \dtop.vtop.pipeline.z[4]$_SDFFE_PP0P_  (.CLK(clknet_leaf_0_clk),
    .RESET_B(net645),
    .D(_00309_),
    .Q_N(_05478_),
    .Q(\dtop.vtop.pipeline.z[4] ));
 sg13g2_dfrbp_1 \dtop.vtop.pipeline.z[5]$_SDFFE_PP0P_  (.CLK(clknet_leaf_0_clk),
    .RESET_B(net646),
    .D(_00310_),
    .Q_N(_05477_),
    .Q(\dtop.vtop.pipeline.z[5] ));
 sg13g2_dfrbp_1 \dtop.vtop.pipeline.z[6]$_SDFFE_PP0P_  (.CLK(clknet_leaf_57_clk),
    .RESET_B(net647),
    .D(_00311_),
    .Q_N(_05476_),
    .Q(\dtop.vtop.pipeline.z[6] ));
 sg13g2_dfrbp_1 \dtop.vtop.pipeline.z[7]$_SDFFE_PP0P_  (.CLK(clknet_leaf_57_clk),
    .RESET_B(net648),
    .D(_00312_),
    .Q_N(_05475_),
    .Q(\dtop.vtop.pipeline.z[7] ));
 sg13g2_dfrbp_1 \dtop.vtop.pipeline.z[8]$_SDFFE_PP0P_  (.CLK(clknet_leaf_57_clk),
    .RESET_B(net649),
    .D(_00313_),
    .Q_N(_05474_),
    .Q(\dtop.vtop.pipeline.z[8] ));
 sg13g2_dfrbp_1 \dtop.vtop.pipeline.z[9]$_SDFFE_PP0P_  (.CLK(clknet_leaf_0_clk),
    .RESET_B(net650),
    .D(_00314_),
    .Q_N(_05473_),
    .Q(\dtop.vtop.pipeline.z[9] ));
 sg13g2_dfrbp_1 \dtop.vtop.pipeline.zg[0]$_DFFE_PP_  (.CLK(clknet_leaf_55_clk),
    .RESET_B(net651),
    .D(_00315_),
    .Q_N(_05472_),
    .Q(\dtop.vtop.pipeline.zg[0] ));
 sg13g2_dfrbp_1 \dtop.vtop.pipeline.zg[1]$_DFFE_PP_  (.CLK(clknet_leaf_57_clk),
    .RESET_B(net652),
    .D(_00316_),
    .Q_N(_05471_),
    .Q(\dtop.vtop.pipeline.zg[1] ));
 sg13g2_dfrbp_1 \dtop.vtop.pipeline.zg[2]$_DFFE_PP_  (.CLK(clknet_leaf_57_clk),
    .RESET_B(net653),
    .D(_00317_),
    .Q_N(_05470_),
    .Q(\dtop.vtop.pipeline.zg[2] ));
 sg13g2_dfrbp_1 \dtop.vtop.pipeline.zg[3]$_DFFE_PP_  (.CLK(clknet_leaf_53_clk),
    .RESET_B(net654),
    .D(_00318_),
    .Q_N(_05469_),
    .Q(\dtop.vtop.pipeline.zg[3] ));
 sg13g2_dfrbp_1 \dtop.vtop.pipeline.zg[4]$_DFFE_PP_  (.CLK(clknet_leaf_56_clk),
    .RESET_B(net655),
    .D(_00319_),
    .Q_N(_05468_),
    .Q(\dtop.vtop.pipeline.zg[4] ));
 sg13g2_dfrbp_1 \dtop.vtop.pipeline.zg[5]$_DFFE_PP_  (.CLK(clknet_leaf_2_clk),
    .RESET_B(net656),
    .D(_00320_),
    .Q_N(_05467_),
    .Q(\dtop.vtop.pipeline.zg[5] ));
 sg13g2_dfrbp_1 \dtop.vtop.pipeline.zg[6]$_DFFE_PP_  (.CLK(clknet_leaf_0_clk),
    .RESET_B(net657),
    .D(_00321_),
    .Q_N(_05466_),
    .Q(\dtop.vtop.pipeline.zg[6] ));
 sg13g2_dfrbp_1 \dtop.vtop.pipeline.zg[7]$_DFFE_PP_  (.CLK(clknet_leaf_2_clk),
    .RESET_B(net658),
    .D(_00322_),
    .Q_N(_05465_),
    .Q(\dtop.vtop.pipeline.zg[7] ));
 sg13g2_dfrbp_1 \dtop.vtop.pipeline.zg[8]$_DFFE_PP_  (.CLK(clknet_leaf_2_clk),
    .RESET_B(net659),
    .D(_00323_),
    .Q_N(_05464_),
    .Q(\dtop.vtop.pipeline.zg[8] ));
 sg13g2_dfrbp_1 \dtop.vtop.pipeline.zg[9]$_DFFE_PP_  (.CLK(clknet_leaf_7_clk),
    .RESET_B(net660),
    .D(_00324_),
    .Q_N(_05463_),
    .Q(\dtop.vtop.pipeline.zg[9] ));
 sg13g2_dfrbp_1 \dtop.vtop.pipeline.zg_acc[0]$_DFFE_PN_  (.CLK(clknet_leaf_52_clk),
    .RESET_B(net661),
    .D(_00325_),
    .Q_N(_05462_),
    .Q(\dtop.vtop.pipeline.zg_acc[0] ));
 sg13g2_dfrbp_1 \dtop.vtop.pipeline.zg_acc[1]$_DFFE_PN_  (.CLK(clknet_leaf_55_clk),
    .RESET_B(net662),
    .D(_00326_),
    .Q_N(_00047_),
    .Q(\dtop.vtop.pipeline.zg_acc[1] ));
 sg13g2_dfrbp_1 \dtop.vtop.pipeline.zg_acc[2]$_DFFE_PN_  (.CLK(clknet_leaf_55_clk),
    .RESET_B(net663),
    .D(_00327_),
    .Q_N(_05461_),
    .Q(\dtop.vtop.pipeline.zg_acc[2] ));
 sg13g2_dfrbp_1 \dtop.vtop.pipeline.zg_acc[3]$_DFFE_PN_  (.CLK(clknet_leaf_52_clk),
    .RESET_B(net664),
    .D(_00328_),
    .Q_N(_05460_),
    .Q(\dtop.vtop.pipeline.zg_acc[3] ));
 sg13g2_dfrbp_1 \dtop.vtop.pipeline.zg_acc[4]$_DFFE_PN_  (.CLK(clknet_leaf_55_clk),
    .RESET_B(net665),
    .D(_00329_),
    .Q_N(_05459_),
    .Q(\dtop.vtop.pipeline.zg_acc[4] ));
 sg13g2_dfrbp_1 \dtop.vtop.pipeline.zg_acc[5]$_DFFE_PN_  (.CLK(clknet_leaf_2_clk),
    .RESET_B(net666),
    .D(_00330_),
    .Q_N(_05458_),
    .Q(\dtop.vtop.pipeline.zg_acc[5] ));
 sg13g2_dfrbp_1 \dtop.vtop.pipeline.zg_acc[6]$_DFFE_PN_  (.CLK(clknet_leaf_55_clk),
    .RESET_B(net667),
    .D(_00331_),
    .Q_N(_00056_),
    .Q(\dtop.vtop.pipeline.zg_acc[6] ));
 sg13g2_dfrbp_1 \dtop.vtop.pipeline.zg_acc[7]$_DFFE_PN_  (.CLK(clknet_leaf_55_clk),
    .RESET_B(net668),
    .D(_00332_),
    .Q_N(_00058_),
    .Q(\dtop.vtop.pipeline.zg_acc[7] ));
 sg13g2_dfrbp_1 \dtop.vtop.pipeline.zg_acc[8]$_DFFE_PN_  (.CLK(clknet_leaf_48_clk),
    .RESET_B(net669),
    .D(_00333_),
    .Q_N(_00079_),
    .Q(\dtop.vtop.pipeline.zg_acc[8] ));
 sg13g2_dfrbp_1 \dtop.vtop.pipeline.zg_acc[9]$_DFFE_PN_  (.CLK(clknet_4_6_0_clk),
    .RESET_B(net670),
    .D(_00334_),
    .Q_N(_05457_),
    .Q(\dtop.vtop.pipeline.zg_acc[9] ));
 sg13g2_dfrbp_1 \dtop.vtop.pipeline.zg_valid$_SDFFE_PP0P_  (.CLK(clknet_leaf_3_clk),
    .RESET_B(net671),
    .D(_00335_),
    .Q_N(_00089_),
    .Q(\dtop.vtop.pipeline.zg_valid ));
 sg13g2_dfrbp_1 \dtop.vtop.r_frame_counter[0]$_SDFF_PP0_  (.CLK(clknet_leaf_20_clk),
    .RESET_B(net672),
    .D(_00336_),
    .Q_N(_00014_),
    .Q(\dtop.detune_counter[4] ));
 sg13g2_dfrbp_1 \dtop.vtop.r_frame_counter[10]$_SDFF_PP0_  (.CLK(clknet_leaf_22_clk),
    .RESET_B(net673),
    .D(_00337_),
    .Q_N(_00029_),
    .Q(\dtop.detune_counter[14] ));
 sg13g2_dfrbp_1 \dtop.vtop.r_frame_counter[11]$_SDFF_PP0_  (.CLK(clknet_leaf_10_clk),
    .RESET_B(net674),
    .D(_00338_),
    .Q_N(_00059_),
    .Q(\dtop.detune_counter[15] ));
 sg13g2_dfrbp_1 \dtop.vtop.r_frame_counter[12]$_SDFF_PP0_  (.CLK(clknet_leaf_20_clk),
    .RESET_B(net675),
    .D(_00339_),
    .Q_N(_00074_),
    .Q(\dtop.detune_counter[16] ));
 sg13g2_dfrbp_1 \dtop.vtop.r_frame_counter[13]$_SDFF_PP0_  (.CLK(clknet_leaf_10_clk),
    .RESET_B(net676),
    .D(_00340_),
    .Q_N(_00086_),
    .Q(\dtop.detune_counter[17] ));
 sg13g2_dfrbp_1 \dtop.vtop.r_frame_counter[1]$_SDFF_PP0_  (.CLK(clknet_leaf_20_clk),
    .RESET_B(net677),
    .D(_00341_),
    .Q_N(_00080_),
    .Q(\dtop.detune_counter[5] ));
 sg13g2_dfrbp_1 \dtop.vtop.r_frame_counter[2]$_SDFF_PP0_  (.CLK(clknet_leaf_20_clk),
    .RESET_B(net678),
    .D(_00342_),
    .Q_N(_00019_),
    .Q(\dtop.detune_counter[6] ));
 sg13g2_dfrbp_1 \dtop.vtop.r_frame_counter[3]$_SDFF_PP0_  (.CLK(clknet_leaf_20_clk),
    .RESET_B(net679),
    .D(_00343_),
    .Q_N(_00017_),
    .Q(\dtop.detune_counter[7] ));
 sg13g2_dfrbp_1 \dtop.vtop.r_frame_counter[4]$_SDFF_PP0_  (.CLK(clknet_leaf_22_clk),
    .RESET_B(net680),
    .D(_00344_),
    .Q_N(_00022_),
    .Q(\dtop.detune_counter[8] ));
 sg13g2_dfrbp_1 \dtop.vtop.r_frame_counter[5]$_SDFF_PP0_  (.CLK(clknet_leaf_21_clk),
    .RESET_B(net681),
    .D(_00345_),
    .Q_N(_00020_),
    .Q(\dtop.detune_counter[9] ));
 sg13g2_dfrbp_1 \dtop.vtop.r_frame_counter[6]$_SDFF_PP0_  (.CLK(clknet_leaf_21_clk),
    .RESET_B(net682),
    .D(_00346_),
    .Q_N(_00024_),
    .Q(\dtop.detune_counter[10] ));
 sg13g2_dfrbp_1 \dtop.vtop.r_frame_counter[7]$_SDFF_PP0_  (.CLK(clknet_leaf_10_clk),
    .RESET_B(net683),
    .D(_00347_),
    .Q_N(_00001_),
    .Q(\dtop.detune_counter[11] ));
 sg13g2_dfrbp_1 \dtop.vtop.r_frame_counter[8]$_SDFF_PP0_  (.CLK(clknet_leaf_10_clk),
    .RESET_B(net684),
    .D(_00348_),
    .Q_N(_00028_),
    .Q(\dtop.detune_counter[12] ));
 sg13g2_dfrbp_1 \dtop.vtop.r_frame_counter[9]$_SDFF_PP0_  (.CLK(clknet_leaf_10_clk),
    .RESET_B(net685),
    .D(_00349_),
    .Q_N(_00000_),
    .Q(\dtop.detune_counter[13] ));
 sg13g2_dfrbp_1 \dtop.vtop.rs.r_vsync$_DFFE_PP_  (.CLK(clknet_leaf_16_clk),
    .RESET_B(net686),
    .D(_00350_),
    .Q_N(\uio_out0b[5] ),
    .Q(\dtop.vsync ));
 sg13g2_dfrbp_1 \dtop.vtop.rs.scan_y.phase[0]$_SDFF_PN0_  (.CLK(clknet_leaf_11_clk),
    .RESET_B(net687),
    .D(_00351_),
    .Q_N(_05456_),
    .Q(\dtop.vtop.rs.scan_y.phase[0] ));
 sg13g2_dfrbp_1 \dtop.vtop.rs.scan_y.phase[1]$_SDFF_PN0_  (.CLK(clknet_leaf_11_clk),
    .RESET_B(net688),
    .D(_00352_),
    .Q_N(_05455_),
    .Q(\dtop.vtop.rs.scan_y.phase[1] ));
 sg13g2_dfrbp_1 \dtop.vtop.rs.scan_y.y[0]$_SDFF_PP0_  (.CLK(clknet_leaf_10_clk),
    .RESET_B(net689),
    .D(_00353_),
    .Q_N(_00083_),
    .Q(\dtop.player_inst.oct_counter[3] ));
 sg13g2_dfrbp_1 \dtop.vtop.rs.scan_y.y[1]$_SDFF_PP0_  (.CLK(clknet_leaf_10_clk),
    .RESET_B(net690),
    .D(_00354_),
    .Q_N(_05454_),
    .Q(\dtop.player_inst.oct_counter[4] ));
 sg13g2_dfrbp_1 \dtop.vtop.rs.scan_y.y[2]$_SDFF_PP0_  (.CLK(clknet_leaf_11_clk),
    .RESET_B(net691),
    .D(_00355_),
    .Q_N(_00066_),
    .Q(\dtop.player_inst.oct_counter[5] ));
 sg13g2_dfrbp_1 \dtop.vtop.rs.scan_y.y[3]$_SDFF_PP0_  (.CLK(clknet_leaf_11_clk),
    .RESET_B(net692),
    .D(_00356_),
    .Q_N(_00065_),
    .Q(\dtop.player_inst.oct_counter[6] ));
 sg13g2_dfrbp_1 \dtop.vtop.rs.scan_y.y[4]$_SDFF_PP0_  (.CLK(clknet_leaf_21_clk),
    .RESET_B(net693),
    .D(_00357_),
    .Q_N(_00064_),
    .Q(\dtop.vtop.logo.addr[7] ));
 sg13g2_dfrbp_1 \dtop.vtop.rs.scan_y.y[5]$_SDFF_PP0_  (.CLK(clknet_leaf_16_clk),
    .RESET_B(net694),
    .D(_00358_),
    .Q_N(_05453_),
    .Q(\dtop.vtop.logo.addr[8] ));
 sg13g2_dfrbp_1 \dtop.vtop.rs.scan_y.y[6]$_SDFF_PP0_  (.CLK(clknet_leaf_15_clk),
    .RESET_B(net695),
    .D(_00359_),
    .Q_N(_00063_),
    .Q(\dtop.vtop.logo.addr[9] ));
 sg13g2_dfrbp_1 \dtop.vtop.rs.scan_y.y[7]$_SDFF_PP0_  (.CLK(clknet_leaf_15_clk),
    .RESET_B(net696),
    .D(_00360_),
    .Q_N(_00062_),
    .Q(\dtop.vtop.logo.addr[10] ));
 sg13g2_dfrbp_1 \dtop.vtop.rs.scan_y.y[8]$_SDFF_PP0_  (.CLK(clknet_leaf_15_clk),
    .RESET_B(net697),
    .D(_00361_),
    .Q_N(_00061_),
    .Q(\dtop.vtop.logo.addr[11] ));
 sg13g2_dfrbp_1 \dtop.vtop.rs.scan_y.y[9]$_SDFF_PN0_  (.CLK(clknet_leaf_15_clk),
    .RESET_B(net698),
    .D(_00362_),
    .Q_N(_05452_),
    .Q(\dtop.vtop.rs.saturated ));
 sg13g2_dfrbp_1 \dtop.vtop.rs.x_scan.phase[0]$_SDFF_PN0_  (.CLK(clknet_leaf_10_clk),
    .RESET_B(net699),
    .D(_00363_),
    .Q_N(_05451_),
    .Q(\dtop.vtop.rs.x_scan.phase[0] ));
 sg13g2_dfrbp_1 \dtop.vtop.rs.x_scan.phase[1]$_SDFF_PN1_  (.CLK(clknet_leaf_23_clk),
    .RESET_B(net700),
    .D(_00364_),
    .Q_N(_05450_),
    .Q(\dtop.vtop.rs.x_scan.phase[1] ));
 sg13g2_dfrbp_1 \dtop.vtop.rs.x_scan.r_coarse[0]$_SDFF_PN0_  (.CLK(clknet_leaf_36_clk),
    .RESET_B(net701),
    .D(_00365_),
    .Q_N(_00084_),
    .Q(\dtop.player_inst.oct_counter[0] ));
 sg13g2_dfrbp_1 \dtop.vtop.rs.x_scan.r_coarse[1]$_SDFF_PN0_  (.CLK(clknet_leaf_36_clk),
    .RESET_B(net702),
    .D(_00366_),
    .Q_N(_05449_),
    .Q(\dtop.player_inst.oct_counter[1] ));
 sg13g2_dfrbp_1 \dtop.vtop.rs.x_scan.r_coarse[2]$_SDFF_PN0_  (.CLK(clknet_leaf_36_clk),
    .RESET_B(net703),
    .D(_00367_),
    .Q_N(_00077_),
    .Q(\dtop.player_inst.oct_counter[2] ));
 sg13g2_dfrbp_1 \dtop.vtop.rs.x_scan.r_fine[0]$_SDFF_PP0_  (.CLK(clknet_4_11_0_clk),
    .RESET_B(net704),
    .D(_00368_),
    .Q_N(_05448_),
    .Q(\dtop.player_inst.program_addr[0] ));
 sg13g2_dfrbp_1 \dtop.vtop.rs.x_scan.r_fine[1]$_SDFF_PP0_  (.CLK(clknet_leaf_40_clk),
    .RESET_B(net705),
    .D(_00369_),
    .Q_N(_00005_),
    .Q(\dtop.player_inst.program_addr[1] ));
 sg13g2_dfrbp_1 \dtop.vtop.rs.x_scan.r_fine[2]$_SDFF_PP0_  (.CLK(clknet_leaf_40_clk),
    .RESET_B(net706),
    .D(_00370_),
    .Q_N(_00090_),
    .Q(\dtop.player_inst.program_addr[2] ));
 sg13g2_dfrbp_1 \dtop.vtop.rs.x_scan.r_fine[3]$_SDFF_PP0_  (.CLK(clknet_leaf_37_clk),
    .RESET_B(net707),
    .D(_00371_),
    .Q_N(_00002_),
    .Q(\dtop.player_inst.program_addr[3] ));
 sg13g2_dfrbp_1 \dtop.vtop.rs.x_scan.r_fine[4]$_SDFF_PP0_  (.CLK(clknet_leaf_41_clk),
    .RESET_B(net708),
    .D(_00372_),
    .Q_N(_05447_),
    .Q(\dtop.player_inst.program_addr[4] ));
 sg13g2_dfrbp_1 \dtop.vtop.rs.x_scan.r_fine[5]$_SDFF_PP0_  (.CLK(clknet_leaf_37_clk),
    .RESET_B(net709),
    .D(_00373_),
    .Q_N(_05446_),
    .Q(\dtop.player_inst.program_addr[5] ));
 sg13g2_dfrbp_1 \dtop.vtop.rs.x_scan.r_fine[6]$_SDFF_PP0_  (.CLK(clknet_leaf_41_clk),
    .RESET_B(net710),
    .D(_00374_),
    .Q_N(_00078_),
    .Q(\dtop.player_inst.program_addr[6] ));
 sg13g2_dfrbp_1 \dtop.vtop.xfrac_counter$_SDFF_PN0_  (.CLK(clknet_leaf_23_clk),
    .RESET_B(net711),
    .D(_00375_),
    .Q_N(_05428_),
    .Q(\dtop.enable ));
 sg13g2_dfrbp_1 \rst_n_reg$_DFF_P_  (.CLK(clknet_leaf_15_clk),
    .RESET_B(net712),
    .D(net1),
    .Q_N(_00085_),
    .Q(rst_n_reg));
 sg13g2_dfrbp_1 \ui_in_reg[0]$_DFF_P_  (.CLK(clknet_leaf_18_clk),
    .RESET_B(net713),
    .D(net2),
    .Q_N(_05631_),
    .Q(\dtop.ext_control[0] ));
 sg13g2_dfrbp_1 \ui_in_reg[1]$_DFF_P_  (.CLK(clknet_leaf_18_clk),
    .RESET_B(net714),
    .D(net3),
    .Q_N(_05632_),
    .Q(\dtop.ext_control[1] ));
 sg13g2_dfrbp_1 \ui_in_reg[2]$_DFF_P_  (.CLK(clknet_leaf_18_clk),
    .RESET_B(net715),
    .D(net4),
    .Q_N(_05633_),
    .Q(\dtop.ext_control[2] ));
 sg13g2_dfrbp_1 \ui_in_reg[3]$_DFF_P_  (.CLK(clknet_leaf_18_clk),
    .RESET_B(net716),
    .D(net5),
    .Q_N(_00082_),
    .Q(\dtop.ext_control[3] ));
 sg13g2_dfrbp_1 \ui_in_reg[4]$_DFF_P_  (.CLK(clknet_4_6_0_clk),
    .RESET_B(net717),
    .D(net6),
    .Q_N(_00012_),
    .Q(\dtop.ext_control[4] ));
 sg13g2_dfrbp_1 \ui_in_reg[5]$_DFF_P_  (.CLK(clknet_leaf_17_clk),
    .RESET_B(net718),
    .D(net7),
    .Q_N(_05634_),
    .Q(\dtop.ext_control[5] ));
 sg13g2_dfrbp_1 \ui_in_reg[6]$_DFF_P_  (.CLK(clknet_leaf_17_clk),
    .RESET_B(net719),
    .D(net8),
    .Q_N(_05635_),
    .Q(\dtop.ext_control[6] ));
 sg13g2_dfrbp_1 \ui_in_reg[7]$_DFF_P_  (.CLK(clknet_leaf_18_clk),
    .RESET_B(net720),
    .D(net9),
    .Q_N(_00081_),
    .Q(advance_frame));
 sg13g2_dfrbp_1 \uio_oe1[4]$_DFFE_PP_  (.CLK(clknet_leaf_13_clk),
    .RESET_B(net721),
    .D(_00376_),
    .Q_N(_05445_),
    .Q(net15));
 sg13g2_dfrbp_1 \uio_out1[0]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_14_clk),
    .RESET_B(net722),
    .D(_00377_),
    .Q_N(_05444_),
    .Q(net16));
 sg13g2_dfrbp_1 \uio_out1[1]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_14_clk),
    .RESET_B(net723),
    .D(_00378_),
    .Q_N(_05443_),
    .Q(net17));
 sg13g2_dfrbp_1 \uio_out1[2]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_14_clk),
    .RESET_B(net724),
    .D(_00379_),
    .Q_N(_05442_),
    .Q(net18));
 sg13g2_dfrbp_1 \uio_out1[3]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_13_clk),
    .RESET_B(net725),
    .D(_00380_),
    .Q_N(_05441_),
    .Q(net19));
 sg13g2_dfrbp_1 \uio_out1[4]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_13_clk),
    .RESET_B(net726),
    .D(_00381_),
    .Q_N(_05440_),
    .Q(net20));
 sg13g2_dfrbp_1 \uio_out1[5]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_13_clk),
    .RESET_B(net727),
    .D(_00382_),
    .Q_N(_05439_),
    .Q(net21));
 sg13g2_dfrbp_1 \uio_out1[6]$_DFFE_PP_  (.CLK(clknet_leaf_13_clk),
    .RESET_B(net728),
    .D(_00383_),
    .Q_N(_05438_),
    .Q(net22));
 sg13g2_dfrbp_1 \uio_out1[7]$_DFFE_PP_  (.CLK(clknet_leaf_13_clk),
    .RESET_B(net729),
    .D(_00384_),
    .Q_N(_05437_),
    .Q(net23));
 sg13g2_dfrbp_1 \uo_out1[0]$_DFFE_PP_  (.CLK(clknet_leaf_16_clk),
    .RESET_B(net730),
    .D(_00385_),
    .Q_N(_05436_),
    .Q(net24));
 sg13g2_dfrbp_1 \uo_out1[1]$_DFFE_PP_  (.CLK(clknet_leaf_16_clk),
    .RESET_B(net731),
    .D(_00386_),
    .Q_N(_05435_),
    .Q(net25));
 sg13g2_dfrbp_1 \uo_out1[2]$_DFFE_PP_  (.CLK(clknet_leaf_17_clk),
    .RESET_B(net732),
    .D(_00387_),
    .Q_N(_05434_),
    .Q(net26));
 sg13g2_dfrbp_1 \uo_out1[3]$_DFFE_PP_  (.CLK(clknet_leaf_16_clk),
    .RESET_B(net733),
    .D(_00388_),
    .Q_N(_05433_),
    .Q(net27));
 sg13g2_dfrbp_1 \uo_out1[4]$_DFFE_PP_  (.CLK(clknet_leaf_16_clk),
    .RESET_B(net734),
    .D(_00389_),
    .Q_N(_05432_),
    .Q(net28));
 sg13g2_dfrbp_1 \uo_out1[5]$_DFFE_PP_  (.CLK(clknet_leaf_14_clk),
    .RESET_B(net735),
    .D(_00390_),
    .Q_N(_05431_),
    .Q(net29));
 sg13g2_dfrbp_1 \uo_out1[6]$_DFFE_PP_  (.CLK(clknet_leaf_14_clk),
    .RESET_B(net736),
    .D(_00391_),
    .Q_N(_05430_),
    .Q(net30));
 sg13g2_dfrbp_1 \uo_out1[7]$_DFFE_PP_  (.CLK(clknet_leaf_16_clk),
    .RESET_B(net737),
    .D(_00392_),
    .Q_N(_05429_),
    .Q(net31));
 sg13g2_buf_1 input1 (.A(rst_n),
    .X(net1));
 sg13g2_buf_1 input2 (.A(ui_in[0]),
    .X(net2));
 sg13g2_buf_1 input3 (.A(ui_in[1]),
    .X(net3));
 sg13g2_buf_1 input4 (.A(ui_in[2]),
    .X(net4));
 sg13g2_buf_1 input5 (.A(ui_in[3]),
    .X(net5));
 sg13g2_buf_1 input6 (.A(ui_in[4]),
    .X(net6));
 sg13g2_buf_1 input7 (.A(ui_in[5]),
    .X(net7));
 sg13g2_buf_1 input8 (.A(ui_in[6]),
    .X(net8));
 sg13g2_buf_1 input9 (.A(ui_in[7]),
    .X(net9));
 sg13g2_buf_1 output10 (.A(net10),
    .X(uio_oe[0]));
 sg13g2_buf_1 output11 (.A(net11),
    .X(uio_oe[1]));
 sg13g2_buf_1 output12 (.A(net12),
    .X(uio_oe[2]));
 sg13g2_buf_1 output13 (.A(net13),
    .X(uio_oe[3]));
 sg13g2_buf_1 output14 (.A(net14),
    .X(uio_oe[4]));
 sg13g2_buf_1 output15 (.A(net15),
    .X(uio_oe[5]));
 sg13g2_buf_1 output16 (.A(net16),
    .X(uio_out[0]));
 sg13g2_buf_1 output17 (.A(net17),
    .X(uio_out[1]));
 sg13g2_buf_1 output18 (.A(net18),
    .X(uio_out[2]));
 sg13g2_buf_1 output19 (.A(net19),
    .X(uio_out[3]));
 sg13g2_buf_1 output20 (.A(net20),
    .X(uio_out[4]));
 sg13g2_buf_1 output21 (.A(net21),
    .X(uio_out[5]));
 sg13g2_buf_1 output22 (.A(net22),
    .X(uio_out[6]));
 sg13g2_buf_1 output23 (.A(net23),
    .X(uio_out[7]));
 sg13g2_buf_1 output24 (.A(net24),
    .X(uo_out[0]));
 sg13g2_buf_1 output25 (.A(net25),
    .X(uo_out[1]));
 sg13g2_buf_1 output26 (.A(net26),
    .X(uo_out[2]));
 sg13g2_buf_1 output27 (.A(net27),
    .X(uo_out[3]));
 sg13g2_buf_1 output28 (.A(net28),
    .X(uo_out[4]));
 sg13g2_buf_1 output29 (.A(net29),
    .X(uo_out[5]));
 sg13g2_buf_1 output30 (.A(net30),
    .X(uo_out[6]));
 sg13g2_buf_1 output31 (.A(net31),
    .X(uo_out[7]));
 sg13g2_buf_2 fanout32 (.A(_04647_),
    .X(net32));
 sg13g2_buf_2 fanout33 (.A(_03230_),
    .X(net33));
 sg13g2_buf_2 fanout34 (.A(_05064_),
    .X(net34));
 sg13g2_buf_2 fanout35 (.A(_05034_),
    .X(net35));
 sg13g2_buf_2 fanout36 (.A(_04436_),
    .X(net36));
 sg13g2_buf_2 fanout37 (.A(_04289_),
    .X(net37));
 sg13g2_buf_2 fanout38 (.A(_05094_),
    .X(net38));
 sg13g2_buf_2 fanout39 (.A(_05082_),
    .X(net39));
 sg13g2_buf_2 fanout40 (.A(_04288_),
    .X(net40));
 sg13g2_buf_2 fanout41 (.A(_00699_),
    .X(net41));
 sg13g2_buf_2 fanout42 (.A(_05053_),
    .X(net42));
 sg13g2_buf_2 fanout43 (.A(_05018_),
    .X(net43));
 sg13g2_buf_2 fanout44 (.A(_05017_),
    .X(net44));
 sg13g2_buf_2 fanout45 (.A(_04998_),
    .X(net45));
 sg13g2_buf_2 fanout46 (.A(_04997_),
    .X(net46));
 sg13g2_buf_2 fanout47 (.A(_04702_),
    .X(net47));
 sg13g2_buf_2 fanout48 (.A(_04700_),
    .X(net48));
 sg13g2_buf_2 fanout49 (.A(_00665_),
    .X(net49));
 sg13g2_buf_2 fanout50 (.A(_00652_),
    .X(net50));
 sg13g2_buf_2 fanout51 (.A(_00500_),
    .X(net51));
 sg13g2_buf_2 fanout52 (.A(_00687_),
    .X(net52));
 sg13g2_buf_2 fanout53 (.A(_00673_),
    .X(net53));
 sg13g2_buf_2 fanout54 (.A(_00671_),
    .X(net54));
 sg13g2_buf_2 fanout55 (.A(_00654_),
    .X(net55));
 sg13g2_buf_2 fanout56 (.A(_00651_),
    .X(net56));
 sg13g2_buf_2 fanout57 (.A(_00640_),
    .X(net57));
 sg13g2_buf_2 fanout58 (.A(_00607_),
    .X(net58));
 sg13g2_buf_2 fanout59 (.A(_00581_),
    .X(net59));
 sg13g2_buf_2 fanout60 (.A(_00499_),
    .X(net60));
 sg13g2_buf_2 fanout61 (.A(_00719_),
    .X(net61));
 sg13g2_buf_2 fanout62 (.A(_00670_),
    .X(net62));
 sg13g2_buf_2 fanout63 (.A(_00668_),
    .X(net63));
 sg13g2_buf_2 fanout64 (.A(_00666_),
    .X(net64));
 sg13g2_buf_2 fanout65 (.A(_00606_),
    .X(net65));
 sg13g2_buf_2 fanout66 (.A(_00597_),
    .X(net66));
 sg13g2_buf_2 fanout67 (.A(_00567_),
    .X(net67));
 sg13g2_buf_2 fanout68 (.A(_00734_),
    .X(net68));
 sg13g2_buf_2 fanout69 (.A(_00716_),
    .X(net69));
 sg13g2_buf_2 fanout70 (.A(_00596_),
    .X(net70));
 sg13g2_buf_2 fanout71 (.A(_00591_),
    .X(net71));
 sg13g2_buf_2 fanout72 (.A(_00566_),
    .X(net72));
 sg13g2_buf_2 fanout73 (.A(_00536_),
    .X(net73));
 sg13g2_buf_2 fanout74 (.A(_00800_),
    .X(net74));
 sg13g2_buf_2 fanout75 (.A(_00762_),
    .X(net75));
 sg13g2_buf_2 fanout76 (.A(_00638_),
    .X(net76));
 sg13g2_buf_2 fanout77 (.A(_00602_),
    .X(net77));
 sg13g2_buf_2 fanout78 (.A(_00595_),
    .X(net78));
 sg13g2_buf_2 fanout79 (.A(_00584_),
    .X(net79));
 sg13g2_buf_2 fanout80 (.A(_00532_),
    .X(net80));
 sg13g2_buf_2 fanout81 (.A(_04720_),
    .X(net81));
 sg13g2_buf_2 fanout82 (.A(_03744_),
    .X(net82));
 sg13g2_buf_2 fanout83 (.A(_03743_),
    .X(net83));
 sg13g2_buf_2 fanout84 (.A(_03365_),
    .X(net84));
 sg13g2_buf_2 fanout85 (.A(_02153_),
    .X(net85));
 sg13g2_buf_2 fanout86 (.A(_01750_),
    .X(net86));
 sg13g2_buf_2 fanout87 (.A(_00799_),
    .X(net87));
 sg13g2_buf_2 fanout88 (.A(_00659_),
    .X(net88));
 sg13g2_buf_2 fanout89 (.A(_00583_),
    .X(net89));
 sg13g2_buf_2 fanout90 (.A(_00580_),
    .X(net90));
 sg13g2_buf_2 fanout91 (.A(_00574_),
    .X(net91));
 sg13g2_buf_2 fanout92 (.A(_00563_),
    .X(net92));
 sg13g2_buf_2 fanout93 (.A(_00531_),
    .X(net93));
 sg13g2_buf_2 fanout94 (.A(_00494_),
    .X(net94));
 sg13g2_buf_2 fanout95 (.A(_03364_),
    .X(net95));
 sg13g2_buf_2 fanout96 (.A(_03331_),
    .X(net96));
 sg13g2_buf_2 fanout97 (.A(_02549_),
    .X(net97));
 sg13g2_buf_2 fanout98 (.A(_02546_),
    .X(net98));
 sg13g2_buf_2 fanout99 (.A(_01870_),
    .X(net99));
 sg13g2_buf_2 fanout100 (.A(_01749_),
    .X(net100));
 sg13g2_buf_2 fanout101 (.A(_01739_),
    .X(net101));
 sg13g2_buf_4 fanout102 (.X(net102),
    .A(_01598_));
 sg13g2_buf_2 fanout103 (.A(_01525_),
    .X(net103));
 sg13g2_buf_4 fanout104 (.X(net104),
    .A(_01517_));
 sg13g2_buf_2 fanout105 (.A(_01485_),
    .X(net105));
 sg13g2_buf_2 fanout106 (.A(_00744_),
    .X(net106));
 sg13g2_buf_2 fanout107 (.A(_00710_),
    .X(net107));
 sg13g2_buf_2 fanout108 (.A(_00613_),
    .X(net108));
 sg13g2_buf_2 fanout109 (.A(_00579_),
    .X(net109));
 sg13g2_buf_2 fanout110 (.A(_00530_),
    .X(net110));
 sg13g2_buf_2 fanout111 (.A(_04783_),
    .X(net111));
 sg13g2_buf_2 fanout112 (.A(_03330_),
    .X(net112));
 sg13g2_buf_2 fanout113 (.A(_02721_),
    .X(net113));
 sg13g2_buf_2 fanout114 (.A(_02717_),
    .X(net114));
 sg13g2_buf_2 fanout115 (.A(_02695_),
    .X(net115));
 sg13g2_buf_2 fanout116 (.A(_02657_),
    .X(net116));
 sg13g2_buf_2 fanout117 (.A(_02564_),
    .X(net117));
 sg13g2_buf_2 fanout118 (.A(_02548_),
    .X(net118));
 sg13g2_buf_2 fanout119 (.A(_02533_),
    .X(net119));
 sg13g2_buf_2 fanout120 (.A(_02484_),
    .X(net120));
 sg13g2_buf_2 fanout121 (.A(_02475_),
    .X(net121));
 sg13g2_buf_2 fanout122 (.A(_02451_),
    .X(net122));
 sg13g2_buf_2 fanout123 (.A(_02446_),
    .X(net123));
 sg13g2_buf_2 fanout124 (.A(_02393_),
    .X(net124));
 sg13g2_buf_2 fanout125 (.A(_02378_),
    .X(net125));
 sg13g2_buf_2 fanout126 (.A(_02374_),
    .X(net126));
 sg13g2_buf_2 fanout127 (.A(_01761_),
    .X(net127));
 sg13g2_buf_2 fanout128 (.A(_01622_),
    .X(net128));
 sg13g2_buf_2 fanout129 (.A(_01524_),
    .X(net129));
 sg13g2_buf_2 fanout130 (.A(_00866_),
    .X(net130));
 sg13g2_buf_2 fanout131 (.A(_00737_),
    .X(net131));
 sg13g2_buf_2 fanout132 (.A(_00612_),
    .X(net132));
 sg13g2_buf_2 fanout133 (.A(_00587_),
    .X(net133));
 sg13g2_buf_2 fanout134 (.A(_00578_),
    .X(net134));
 sg13g2_buf_2 fanout135 (.A(_00561_),
    .X(net135));
 sg13g2_buf_2 fanout136 (.A(_00547_),
    .X(net136));
 sg13g2_buf_2 fanout137 (.A(_00529_),
    .X(net137));
 sg13g2_buf_2 fanout138 (.A(_04667_),
    .X(net138));
 sg13g2_buf_2 fanout139 (.A(_04385_),
    .X(net139));
 sg13g2_buf_2 fanout140 (.A(_04382_),
    .X(net140));
 sg13g2_buf_2 fanout141 (.A(_03870_),
    .X(net141));
 sg13g2_buf_2 fanout142 (.A(_02658_),
    .X(net142));
 sg13g2_buf_2 fanout143 (.A(_02613_),
    .X(net143));
 sg13g2_buf_2 fanout144 (.A(_02606_),
    .X(net144));
 sg13g2_buf_2 fanout145 (.A(_02602_),
    .X(net145));
 sg13g2_buf_2 fanout146 (.A(_02568_),
    .X(net146));
 sg13g2_buf_2 fanout147 (.A(_02563_),
    .X(net147));
 sg13g2_buf_2 fanout148 (.A(_02540_),
    .X(net148));
 sg13g2_buf_2 fanout149 (.A(_02538_),
    .X(net149));
 sg13g2_buf_2 fanout150 (.A(_02536_),
    .X(net150));
 sg13g2_buf_2 fanout151 (.A(_02517_),
    .X(net151));
 sg13g2_buf_2 fanout152 (.A(_02488_),
    .X(net152));
 sg13g2_buf_2 fanout153 (.A(_02485_),
    .X(net153));
 sg13g2_buf_2 fanout154 (.A(_02479_),
    .X(net154));
 sg13g2_buf_2 fanout155 (.A(_02474_),
    .X(net155));
 sg13g2_buf_2 fanout156 (.A(_02450_),
    .X(net156));
 sg13g2_buf_2 fanout157 (.A(_02443_),
    .X(net157));
 sg13g2_buf_2 fanout158 (.A(_02440_),
    .X(net158));
 sg13g2_buf_2 fanout159 (.A(_02427_),
    .X(net159));
 sg13g2_buf_2 fanout160 (.A(_02422_),
    .X(net160));
 sg13g2_buf_2 fanout161 (.A(_02411_),
    .X(net161));
 sg13g2_buf_2 fanout162 (.A(_02392_),
    .X(net162));
 sg13g2_buf_2 fanout163 (.A(_02377_),
    .X(net163));
 sg13g2_buf_2 fanout164 (.A(_02373_),
    .X(net164));
 sg13g2_buf_2 fanout165 (.A(_02372_),
    .X(net165));
 sg13g2_buf_2 fanout166 (.A(_02287_),
    .X(net166));
 sg13g2_buf_2 fanout167 (.A(_01845_),
    .X(net167));
 sg13g2_buf_2 fanout168 (.A(_00674_),
    .X(net168));
 sg13g2_buf_2 fanout169 (.A(_00611_),
    .X(net169));
 sg13g2_buf_2 fanout170 (.A(_00585_),
    .X(net170));
 sg13g2_buf_2 fanout171 (.A(_00577_),
    .X(net171));
 sg13g2_buf_2 fanout172 (.A(_00571_),
    .X(net172));
 sg13g2_buf_2 fanout173 (.A(_04311_),
    .X(net173));
 sg13g2_buf_2 fanout174 (.A(_04234_),
    .X(net174));
 sg13g2_buf_2 fanout175 (.A(_04231_),
    .X(net175));
 sg13g2_buf_2 fanout176 (.A(_03054_),
    .X(net176));
 sg13g2_buf_2 fanout177 (.A(_02871_),
    .X(net177));
 sg13g2_buf_2 fanout178 (.A(_02697_),
    .X(net178));
 sg13g2_buf_2 fanout179 (.A(_02618_),
    .X(net179));
 sg13g2_buf_2 fanout180 (.A(_02599_),
    .X(net180));
 sg13g2_buf_2 fanout181 (.A(_02567_),
    .X(net181));
 sg13g2_buf_2 fanout182 (.A(_02539_),
    .X(net182));
 sg13g2_buf_2 fanout183 (.A(_02537_),
    .X(net183));
 sg13g2_buf_2 fanout184 (.A(_02529_),
    .X(net184));
 sg13g2_buf_2 fanout185 (.A(_02526_),
    .X(net185));
 sg13g2_buf_2 fanout186 (.A(_02516_),
    .X(net186));
 sg13g2_buf_2 fanout187 (.A(_02478_),
    .X(net187));
 sg13g2_buf_2 fanout188 (.A(_02473_),
    .X(net188));
 sg13g2_buf_2 fanout189 (.A(_02462_),
    .X(net189));
 sg13g2_buf_2 fanout190 (.A(_02449_),
    .X(net190));
 sg13g2_buf_2 fanout191 (.A(_02425_),
    .X(net191));
 sg13g2_buf_2 fanout192 (.A(_02419_),
    .X(net192));
 sg13g2_buf_2 fanout193 (.A(_02410_),
    .X(net193));
 sg13g2_buf_2 fanout194 (.A(_02376_),
    .X(net194));
 sg13g2_buf_2 fanout195 (.A(_02371_),
    .X(net195));
 sg13g2_buf_2 fanout196 (.A(_02367_),
    .X(net196));
 sg13g2_buf_2 fanout197 (.A(_02329_),
    .X(net197));
 sg13g2_buf_2 fanout198 (.A(_02309_),
    .X(net198));
 sg13g2_buf_2 fanout199 (.A(_01965_),
    .X(net199));
 sg13g2_buf_2 fanout200 (.A(_01746_),
    .X(net200));
 sg13g2_buf_2 fanout201 (.A(_00913_),
    .X(net201));
 sg13g2_buf_2 fanout202 (.A(_00610_),
    .X(net202));
 sg13g2_buf_2 fanout203 (.A(_00576_),
    .X(net203));
 sg13g2_buf_2 fanout204 (.A(_00570_),
    .X(net204));
 sg13g2_buf_2 fanout205 (.A(_00559_),
    .X(net205));
 sg13g2_buf_2 fanout206 (.A(_05240_),
    .X(net206));
 sg13g2_buf_2 fanout207 (.A(_05224_),
    .X(net207));
 sg13g2_buf_2 fanout208 (.A(_05213_),
    .X(net208));
 sg13g2_buf_2 fanout209 (.A(_04310_),
    .X(net209));
 sg13g2_buf_2 fanout210 (.A(_04244_),
    .X(net210));
 sg13g2_buf_2 fanout211 (.A(_03769_),
    .X(net211));
 sg13g2_buf_2 fanout212 (.A(_03762_),
    .X(net212));
 sg13g2_buf_2 fanout213 (.A(_03727_),
    .X(net213));
 sg13g2_buf_2 fanout214 (.A(_03726_),
    .X(net214));
 sg13g2_buf_2 fanout215 (.A(_03360_),
    .X(net215));
 sg13g2_buf_2 fanout216 (.A(_03359_),
    .X(net216));
 sg13g2_buf_2 fanout217 (.A(_03240_),
    .X(net217));
 sg13g2_buf_2 fanout218 (.A(_03239_),
    .X(net218));
 sg13g2_buf_2 fanout219 (.A(_02870_),
    .X(net219));
 sg13g2_buf_2 fanout220 (.A(_02856_),
    .X(net220));
 sg13g2_buf_2 fanout221 (.A(_02690_),
    .X(net221));
 sg13g2_buf_2 fanout222 (.A(_02628_),
    .X(net222));
 sg13g2_buf_2 fanout223 (.A(_02581_),
    .X(net223));
 sg13g2_buf_2 fanout224 (.A(_02561_),
    .X(net224));
 sg13g2_buf_2 fanout225 (.A(_02461_),
    .X(net225));
 sg13g2_buf_2 fanout226 (.A(_02423_),
    .X(net226));
 sg13g2_buf_2 fanout227 (.A(_02375_),
    .X(net227));
 sg13g2_buf_2 fanout228 (.A(_02370_),
    .X(net228));
 sg13g2_buf_2 fanout229 (.A(_02366_),
    .X(net229));
 sg13g2_buf_2 fanout230 (.A(_02325_),
    .X(net230));
 sg13g2_buf_2 fanout231 (.A(_00906_),
    .X(net231));
 sg13g2_buf_2 fanout232 (.A(_05239_),
    .X(net232));
 sg13g2_buf_2 fanout233 (.A(_04404_),
    .X(net233));
 sg13g2_buf_2 fanout234 (.A(_04395_),
    .X(net234));
 sg13g2_buf_2 fanout235 (.A(_04380_),
    .X(net235));
 sg13g2_buf_2 fanout236 (.A(_04309_),
    .X(net236));
 sg13g2_buf_2 fanout237 (.A(_03572_),
    .X(net237));
 sg13g2_buf_2 fanout238 (.A(_03442_),
    .X(net238));
 sg13g2_buf_2 fanout239 (.A(_02864_),
    .X(net239));
 sg13g2_buf_2 fanout240 (.A(_02855_),
    .X(net240));
 sg13g2_buf_2 fanout241 (.A(_02594_),
    .X(net241));
 sg13g2_buf_2 fanout242 (.A(_02593_),
    .X(net242));
 sg13g2_buf_2 fanout243 (.A(_02491_),
    .X(net243));
 sg13g2_buf_2 fanout244 (.A(_02460_),
    .X(net244));
 sg13g2_buf_2 fanout245 (.A(_02330_),
    .X(net245));
 sg13g2_buf_2 fanout246 (.A(_02327_),
    .X(net246));
 sg13g2_buf_2 fanout247 (.A(_02277_),
    .X(net247));
 sg13g2_buf_2 fanout248 (.A(_02254_),
    .X(net248));
 sg13g2_buf_2 fanout249 (.A(_01838_),
    .X(net249));
 sg13g2_buf_2 fanout250 (.A(_04286_),
    .X(net250));
 sg13g2_buf_2 fanout251 (.A(_03445_),
    .X(net251));
 sg13g2_buf_2 fanout252 (.A(_03408_),
    .X(net252));
 sg13g2_buf_2 fanout253 (.A(_03256_),
    .X(net253));
 sg13g2_buf_2 fanout254 (.A(_03169_),
    .X(net254));
 sg13g2_buf_2 fanout255 (.A(_02508_),
    .X(net255));
 sg13g2_buf_2 fanout256 (.A(_02364_),
    .X(net256));
 sg13g2_buf_2 fanout257 (.A(_02354_),
    .X(net257));
 sg13g2_buf_2 fanout258 (.A(_02323_),
    .X(net258));
 sg13g2_buf_2 fanout259 (.A(_01668_),
    .X(net259));
 sg13g2_buf_2 fanout260 (.A(_05284_),
    .X(net260));
 sg13g2_buf_2 fanout261 (.A(_05277_),
    .X(net261));
 sg13g2_buf_2 fanout262 (.A(_05271_),
    .X(net262));
 sg13g2_buf_2 fanout263 (.A(_05248_),
    .X(net263));
 sg13g2_buf_2 fanout264 (.A(_04064_),
    .X(net264));
 sg13g2_buf_2 fanout265 (.A(_03565_),
    .X(net265));
 sg13g2_buf_2 fanout266 (.A(_03425_),
    .X(net266));
 sg13g2_buf_2 fanout267 (.A(_03418_),
    .X(net267));
 sg13g2_buf_2 fanout268 (.A(_02862_),
    .X(net268));
 sg13g2_buf_2 fanout269 (.A(_02623_),
    .X(net269));
 sg13g2_buf_2 fanout270 (.A(_02500_),
    .X(net270));
 sg13g2_buf_4 fanout271 (.X(net271),
    .A(_02454_));
 sg13g2_buf_2 fanout272 (.A(_01857_),
    .X(net272));
 sg13g2_buf_2 fanout273 (.A(_01657_),
    .X(net273));
 sg13g2_buf_2 fanout274 (.A(_01225_),
    .X(net274));
 sg13g2_buf_2 fanout275 (.A(_02292_),
    .X(net275));
 sg13g2_buf_2 fanout276 (.A(_01589_),
    .X(net276));
 sg13g2_buf_2 fanout277 (.A(_05282_),
    .X(net277));
 sg13g2_buf_2 fanout278 (.A(_05179_),
    .X(net278));
 sg13g2_buf_2 fanout279 (.A(_03974_),
    .X(net279));
 sg13g2_buf_2 fanout280 (.A(_01807_),
    .X(net280));
 sg13g2_buf_2 fanout281 (.A(_01774_),
    .X(net281));
 sg13g2_buf_2 fanout282 (.A(_01728_),
    .X(net282));
 sg13g2_buf_2 fanout283 (.A(_01462_),
    .X(net283));
 sg13g2_buf_2 fanout284 (.A(_01333_),
    .X(net284));
 sg13g2_buf_2 fanout285 (.A(_01218_),
    .X(net285));
 sg13g2_buf_2 fanout286 (.A(_00465_),
    .X(net286));
 sg13g2_buf_2 fanout287 (.A(_00462_),
    .X(net287));
 sg13g2_buf_2 fanout288 (.A(_05244_),
    .X(net288));
 sg13g2_buf_2 fanout289 (.A(_05236_),
    .X(net289));
 sg13g2_buf_2 fanout290 (.A(_05178_),
    .X(net290));
 sg13g2_buf_2 fanout291 (.A(_05143_),
    .X(net291));
 sg13g2_buf_2 fanout292 (.A(_01456_),
    .X(net292));
 sg13g2_buf_2 fanout293 (.A(_01349_),
    .X(net293));
 sg13g2_buf_2 fanout294 (.A(_01287_),
    .X(net294));
 sg13g2_buf_2 fanout295 (.A(_01273_),
    .X(net295));
 sg13g2_buf_2 fanout296 (.A(_01197_),
    .X(net296));
 sg13g2_buf_2 fanout297 (.A(_00507_),
    .X(net297));
 sg13g2_buf_2 fanout298 (.A(_00464_),
    .X(net298));
 sg13g2_buf_2 fanout299 (.A(_00461_),
    .X(net299));
 sg13g2_buf_2 fanout300 (.A(_00442_),
    .X(net300));
 sg13g2_buf_2 fanout301 (.A(_05235_),
    .X(net301));
 sg13g2_buf_2 fanout302 (.A(_05204_),
    .X(net302));
 sg13g2_buf_2 fanout303 (.A(_05177_),
    .X(net303));
 sg13g2_buf_2 fanout304 (.A(_05142_),
    .X(net304));
 sg13g2_buf_2 fanout305 (.A(_05135_),
    .X(net305));
 sg13g2_buf_2 fanout306 (.A(_03351_),
    .X(net306));
 sg13g2_buf_2 fanout307 (.A(_01580_),
    .X(net307));
 sg13g2_buf_2 fanout308 (.A(_01398_),
    .X(net308));
 sg13g2_buf_2 fanout309 (.A(_01368_),
    .X(net309));
 sg13g2_buf_2 fanout310 (.A(_01358_),
    .X(net310));
 sg13g2_buf_2 fanout311 (.A(_01340_),
    .X(net311));
 sg13g2_buf_2 fanout312 (.A(_01303_),
    .X(net312));
 sg13g2_buf_2 fanout313 (.A(_01290_),
    .X(net313));
 sg13g2_buf_2 fanout314 (.A(_01278_),
    .X(net314));
 sg13g2_buf_2 fanout315 (.A(_01272_),
    .X(net315));
 sg13g2_buf_2 fanout316 (.A(_01235_),
    .X(net316));
 sg13g2_buf_2 fanout317 (.A(_01229_),
    .X(net317));
 sg13g2_buf_2 fanout318 (.A(_01203_),
    .X(net318));
 sg13g2_buf_2 fanout319 (.A(_00756_),
    .X(net319));
 sg13g2_buf_2 fanout320 (.A(_00688_),
    .X(net320));
 sg13g2_buf_2 fanout321 (.A(_00504_),
    .X(net321));
 sg13g2_buf_2 fanout322 (.A(_00460_),
    .X(net322));
 sg13g2_buf_2 fanout323 (.A(_00435_),
    .X(net323));
 sg13g2_buf_2 fanout324 (.A(_00420_),
    .X(net324));
 sg13g2_buf_2 fanout325 (.A(_05205_),
    .X(net325));
 sg13g2_buf_2 fanout326 (.A(_05181_),
    .X(net326));
 sg13g2_buf_2 fanout327 (.A(_05161_),
    .X(net327));
 sg13g2_buf_2 fanout328 (.A(_05147_),
    .X(net328));
 sg13g2_buf_2 fanout329 (.A(_05141_),
    .X(net329));
 sg13g2_buf_2 fanout330 (.A(_05085_),
    .X(net330));
 sg13g2_buf_2 fanout331 (.A(_05066_),
    .X(net331));
 sg13g2_buf_2 fanout332 (.A(_05031_),
    .X(net332));
 sg13g2_buf_2 fanout333 (.A(_05009_),
    .X(net333));
 sg13g2_buf_2 fanout334 (.A(_04977_),
    .X(net334));
 sg13g2_buf_2 fanout335 (.A(_04960_),
    .X(net335));
 sg13g2_buf_2 fanout336 (.A(_04697_),
    .X(net336));
 sg13g2_buf_2 fanout337 (.A(_03908_),
    .X(net337));
 sg13g2_buf_2 fanout338 (.A(_03366_),
    .X(net338));
 sg13g2_buf_2 fanout339 (.A(_01565_),
    .X(net339));
 sg13g2_buf_2 fanout340 (.A(_01322_),
    .X(net340));
 sg13g2_buf_2 fanout341 (.A(_01293_),
    .X(net341));
 sg13g2_buf_2 fanout342 (.A(_01207_),
    .X(net342));
 sg13g2_buf_2 fanout343 (.A(_00755_),
    .X(net343));
 sg13g2_buf_2 fanout344 (.A(_00642_),
    .X(net344));
 sg13g2_buf_2 fanout345 (.A(_00539_),
    .X(net345));
 sg13g2_buf_2 fanout346 (.A(_00514_),
    .X(net346));
 sg13g2_buf_2 fanout347 (.A(_00459_),
    .X(net347));
 sg13g2_buf_2 fanout348 (.A(_00438_),
    .X(net348));
 sg13g2_buf_2 fanout349 (.A(_00419_),
    .X(net349));
 sg13g2_buf_2 fanout350 (.A(_00407_),
    .X(net350));
 sg13g2_buf_2 fanout351 (.A(_05387_),
    .X(net351));
 sg13g2_buf_2 fanout352 (.A(_05333_),
    .X(net352));
 sg13g2_buf_2 fanout353 (.A(_05216_),
    .X(net353));
 sg13g2_buf_2 fanout354 (.A(_05202_),
    .X(net354));
 sg13g2_buf_2 fanout355 (.A(_05160_),
    .X(net355));
 sg13g2_buf_2 fanout356 (.A(_05157_),
    .X(net356));
 sg13g2_buf_2 fanout357 (.A(_05144_),
    .X(net357));
 sg13g2_buf_2 fanout358 (.A(_05140_),
    .X(net358));
 sg13g2_buf_2 fanout359 (.A(_05025_),
    .X(net359));
 sg13g2_buf_2 fanout360 (.A(_04105_),
    .X(net360));
 sg13g2_buf_2 fanout361 (.A(_04041_),
    .X(net361));
 sg13g2_buf_1 fanout362 (.A(_03907_),
    .X(net362));
 sg13g2_buf_2 fanout363 (.A(_03882_),
    .X(net363));
 sg13g2_buf_2 fanout364 (.A(_03430_),
    .X(net364));
 sg13g2_buf_2 fanout365 (.A(_03413_),
    .X(net365));
 sg13g2_buf_2 fanout366 (.A(_03411_),
    .X(net366));
 sg13g2_buf_2 fanout367 (.A(_03407_),
    .X(net367));
 sg13g2_buf_2 fanout368 (.A(_03405_),
    .X(net368));
 sg13g2_buf_2 fanout369 (.A(_02296_),
    .X(net369));
 sg13g2_buf_2 fanout370 (.A(_02171_),
    .X(net370));
 sg13g2_buf_4 fanout371 (.X(net371),
    .A(_02114_));
 sg13g2_buf_2 fanout372 (.A(_01508_),
    .X(net372));
 sg13g2_buf_2 fanout373 (.A(_01214_),
    .X(net373));
 sg13g2_buf_2 fanout374 (.A(_01189_),
    .X(net374));
 sg13g2_buf_2 fanout375 (.A(_00779_),
    .X(net375));
 sg13g2_buf_2 fanout376 (.A(_00629_),
    .X(net376));
 sg13g2_buf_2 fanout377 (.A(_00522_),
    .X(net377));
 sg13g2_buf_2 fanout378 (.A(_00516_),
    .X(net378));
 sg13g2_buf_2 fanout379 (.A(_00513_),
    .X(net379));
 sg13g2_buf_2 fanout380 (.A(_00502_),
    .X(net380));
 sg13g2_buf_2 fanout381 (.A(_00433_),
    .X(net381));
 sg13g2_buf_2 fanout382 (.A(_00421_),
    .X(net382));
 sg13g2_buf_2 fanout383 (.A(_00418_),
    .X(net383));
 sg13g2_buf_2 fanout384 (.A(_05421_),
    .X(net384));
 sg13g2_buf_2 fanout385 (.A(_05384_),
    .X(net385));
 sg13g2_buf_2 fanout386 (.A(_05368_),
    .X(net386));
 sg13g2_buf_2 fanout387 (.A(_05354_),
    .X(net387));
 sg13g2_buf_2 fanout388 (.A(_05332_),
    .X(net388));
 sg13g2_buf_2 fanout389 (.A(_05281_),
    .X(net389));
 sg13g2_buf_2 fanout390 (.A(_05254_),
    .X(net390));
 sg13g2_buf_2 fanout391 (.A(_05220_),
    .X(net391));
 sg13g2_buf_2 fanout392 (.A(_05215_),
    .X(net392));
 sg13g2_buf_2 fanout393 (.A(_05197_),
    .X(net393));
 sg13g2_buf_2 fanout394 (.A(_05188_),
    .X(net394));
 sg13g2_buf_2 fanout395 (.A(_05182_),
    .X(net395));
 sg13g2_buf_2 fanout396 (.A(_05159_),
    .X(net396));
 sg13g2_buf_2 fanout397 (.A(_05156_),
    .X(net397));
 sg13g2_buf_2 fanout398 (.A(_05152_),
    .X(net398));
 sg13g2_buf_2 fanout399 (.A(_05150_),
    .X(net399));
 sg13g2_buf_2 fanout400 (.A(_05139_),
    .X(net400));
 sg13g2_buf_2 fanout401 (.A(_05137_),
    .X(net401));
 sg13g2_buf_2 fanout402 (.A(_05132_),
    .X(net402));
 sg13g2_buf_2 fanout403 (.A(_04001_),
    .X(net403));
 sg13g2_buf_2 fanout404 (.A(_03980_),
    .X(net404));
 sg13g2_buf_4 fanout405 (.X(net405),
    .A(_03410_));
 sg13g2_buf_2 fanout406 (.A(_03406_),
    .X(net406));
 sg13g2_buf_2 fanout407 (.A(_03404_),
    .X(net407));
 sg13g2_buf_2 fanout408 (.A(_03296_),
    .X(net408));
 sg13g2_buf_2 fanout409 (.A(_03280_),
    .X(net409));
 sg13g2_buf_2 fanout410 (.A(_02381_),
    .X(net410));
 sg13g2_buf_2 fanout411 (.A(_02170_),
    .X(net411));
 sg13g2_buf_2 fanout412 (.A(_01933_),
    .X(net412));
 sg13g2_buf_2 fanout413 (.A(_01895_),
    .X(net413));
 sg13g2_buf_2 fanout414 (.A(_01850_),
    .X(net414));
 sg13g2_buf_2 fanout415 (.A(_01846_),
    .X(net415));
 sg13g2_buf_2 fanout416 (.A(_00521_),
    .X(net416));
 sg13g2_buf_2 fanout417 (.A(_00512_),
    .X(net417));
 sg13g2_buf_2 fanout418 (.A(_00501_),
    .X(net418));
 sg13g2_buf_2 fanout419 (.A(_00450_),
    .X(net419));
 sg13g2_buf_2 fanout420 (.A(_05367_),
    .X(net420));
 sg13g2_buf_2 fanout421 (.A(_05350_),
    .X(net421));
 sg13g2_buf_2 fanout422 (.A(_05346_),
    .X(net422));
 sg13g2_buf_2 fanout423 (.A(_05342_),
    .X(net423));
 sg13g2_buf_2 fanout424 (.A(_05334_),
    .X(net424));
 sg13g2_buf_2 fanout425 (.A(_05290_),
    .X(net425));
 sg13g2_buf_2 fanout426 (.A(_05242_),
    .X(net426));
 sg13g2_buf_2 fanout427 (.A(_05225_),
    .X(net427));
 sg13g2_buf_2 fanout428 (.A(_05185_),
    .X(net428));
 sg13g2_buf_2 fanout429 (.A(_05155_),
    .X(net429));
 sg13g2_tiehi _10969__430 (.L_HI(net430));
 sg13g2_tiehi _10970__431 (.L_HI(net431));
 sg13g2_tiehi _10977__432 (.L_HI(net432));
 sg13g2_tiehi _10978__433 (.L_HI(net433));
 sg13g2_tiehi \dtop.player_inst.synth.alu.acc[0]$_SDFFE_PN0P__434  (.L_HI(net434));
 sg13g2_tiehi \dtop.player_inst.synth.alu.acc[10]$_SDFFE_PN0P__435  (.L_HI(net435));
 sg13g2_tiehi \dtop.player_inst.synth.alu.acc[1]$_SDFFE_PN0P__436  (.L_HI(net436));
 sg13g2_tiehi \dtop.player_inst.synth.alu.acc[2]$_SDFFE_PN0P__437  (.L_HI(net437));
 sg13g2_tiehi \dtop.player_inst.synth.alu.acc[3]$_SDFFE_PN0P__438  (.L_HI(net438));
 sg13g2_tiehi \dtop.player_inst.synth.alu.acc[4]$_SDFFE_PN0P__439  (.L_HI(net439));
 sg13g2_tiehi \dtop.player_inst.synth.alu.acc[5]$_SDFFE_PN0P__440  (.L_HI(net440));
 sg13g2_tiehi \dtop.player_inst.synth.alu.acc[6]$_SDFFE_PN0P__441  (.L_HI(net441));
 sg13g2_tiehi \dtop.player_inst.synth.alu.acc[7]$_SDFFE_PN0P__442  (.L_HI(net442));
 sg13g2_tiehi \dtop.player_inst.synth.alu.acc[8]$_SDFFE_PN0P__443  (.L_HI(net443));
 sg13g2_tiehi \dtop.player_inst.synth.alu.acc[9]$_SDFFE_PN0P__444  (.L_HI(net444));
 sg13g2_tiehi \dtop.player_inst.synth.alu.carry$_SDFFE_PN0P__445  (.L_HI(net445));
 sg13g2_tiehi \dtop.player_inst.synth.alu.oct_en$_DFFE_PP__446  (.L_HI(net446));
 sg13g2_tiehi \dtop.player_inst.synth.alu.registers[0][0]$_SDFFE_PN0P__447  (.L_HI(net447));
 sg13g2_tiehi \dtop.player_inst.synth.alu.registers[0][10]$_SDFFE_PN0P__448  (.L_HI(net448));
 sg13g2_tiehi \dtop.player_inst.synth.alu.registers[0][1]$_SDFFE_PN0P__449  (.L_HI(net449));
 sg13g2_tiehi \dtop.player_inst.synth.alu.registers[0][2]$_SDFFE_PN0P__450  (.L_HI(net450));
 sg13g2_tiehi \dtop.player_inst.synth.alu.registers[0][3]$_SDFFE_PN0P__451  (.L_HI(net451));
 sg13g2_tiehi \dtop.player_inst.synth.alu.registers[0][4]$_SDFFE_PN0P__452  (.L_HI(net452));
 sg13g2_tiehi \dtop.player_inst.synth.alu.registers[0][5]$_SDFFE_PN0P__453  (.L_HI(net453));
 sg13g2_tiehi \dtop.player_inst.synth.alu.registers[0][6]$_SDFFE_PN0P__454  (.L_HI(net454));
 sg13g2_tiehi \dtop.player_inst.synth.alu.registers[0][7]$_SDFFE_PN0P__455  (.L_HI(net455));
 sg13g2_tiehi \dtop.player_inst.synth.alu.registers[0][8]$_SDFFE_PN0P__456  (.L_HI(net456));
 sg13g2_tiehi \dtop.player_inst.synth.alu.registers[0][9]$_SDFFE_PN0P__457  (.L_HI(net457));
 sg13g2_tiehi \dtop.player_inst.synth.alu.registers[1][0]$_SDFFE_PN0P__458  (.L_HI(net458));
 sg13g2_tiehi \dtop.player_inst.synth.alu.registers[1][10]$_SDFFE_PN0P__459  (.L_HI(net459));
 sg13g2_tiehi \dtop.player_inst.synth.alu.registers[1][1]$_SDFFE_PN0P__460  (.L_HI(net460));
 sg13g2_tiehi \dtop.player_inst.synth.alu.registers[1][2]$_SDFFE_PN0P__461  (.L_HI(net461));
 sg13g2_tiehi \dtop.player_inst.synth.alu.registers[1][3]$_SDFFE_PN0P__462  (.L_HI(net462));
 sg13g2_tiehi \dtop.player_inst.synth.alu.registers[1][4]$_SDFFE_PN0P__463  (.L_HI(net463));
 sg13g2_tiehi \dtop.player_inst.synth.alu.registers[1][5]$_SDFFE_PN0P__464  (.L_HI(net464));
 sg13g2_tiehi \dtop.player_inst.synth.alu.registers[1][6]$_SDFFE_PN0P__465  (.L_HI(net465));
 sg13g2_tiehi \dtop.player_inst.synth.alu.registers[1][7]$_SDFFE_PN0P__466  (.L_HI(net466));
 sg13g2_tiehi \dtop.player_inst.synth.alu.registers[1][8]$_SDFFE_PN0P__467  (.L_HI(net467));
 sg13g2_tiehi \dtop.player_inst.synth.alu.registers[1][9]$_SDFFE_PN0P__468  (.L_HI(net468));
 sg13g2_tiehi \dtop.player_inst.synth.alu.registers[2][0]$_SDFFE_PN0P__469  (.L_HI(net469));
 sg13g2_tiehi \dtop.player_inst.synth.alu.registers[2][1]$_SDFFE_PN0P__470  (.L_HI(net470));
 sg13g2_tiehi \dtop.player_inst.synth.alu.registers[2][2]$_SDFFE_PN0P__471  (.L_HI(net471));
 sg13g2_tiehi \dtop.player_inst.synth.alu.registers[2][3]$_SDFFE_PN0P__472  (.L_HI(net472));
 sg13g2_tiehi \dtop.player_inst.synth.alu.registers[2][4]$_SDFFE_PN0P__473  (.L_HI(net473));
 sg13g2_tiehi \dtop.player_inst.synth.alu.registers[2][5]$_SDFFE_PN0P__474  (.L_HI(net474));
 sg13g2_tiehi \dtop.player_inst.synth.alu.registers[2][6]$_SDFFE_PN0P__475  (.L_HI(net475));
 sg13g2_tiehi \dtop.player_inst.synth.alu.registers[2][7]$_SDFFE_PN0P__476  (.L_HI(net476));
 sg13g2_tiehi \dtop.player_inst.synth.alu.registers[3][0]$_SDFFE_PN0P__477  (.L_HI(net477));
 sg13g2_tiehi \dtop.player_inst.synth.alu.registers[3][1]$_SDFFE_PN0P__478  (.L_HI(net478));
 sg13g2_tiehi \dtop.player_inst.synth.alu.registers[3][2]$_SDFFE_PN0P__479  (.L_HI(net479));
 sg13g2_tiehi \dtop.player_inst.synth.alu.registers[3][3]$_SDFFE_PN0P__480  (.L_HI(net480));
 sg13g2_tiehi \dtop.player_inst.synth.alu.registers[3][4]$_SDFFE_PN0P__481  (.L_HI(net481));
 sg13g2_tiehi \dtop.player_inst.synth.alu.registers[3][5]$_SDFFE_PN0P__482  (.L_HI(net482));
 sg13g2_tiehi \dtop.player_inst.synth.alu.registers[3][6]$_SDFFE_PN0P__483  (.L_HI(net483));
 sg13g2_tiehi \dtop.player_inst.synth.alu.registers[3][7]$_SDFFE_PN0P__484  (.L_HI(net484));
 sg13g2_tiehi \dtop.player_inst.synth.alu.registers[4][0]$_SDFFE_PN0P__485  (.L_HI(net485));
 sg13g2_tiehi \dtop.player_inst.synth.alu.registers[4][10]$_SDFFE_PN0P__486  (.L_HI(net486));
 sg13g2_tiehi \dtop.player_inst.synth.alu.registers[4][1]$_SDFFE_PN0P__487  (.L_HI(net487));
 sg13g2_tiehi \dtop.player_inst.synth.alu.registers[4][2]$_SDFFE_PN0P__488  (.L_HI(net488));
 sg13g2_tiehi \dtop.player_inst.synth.alu.registers[4][3]$_SDFFE_PN0P__489  (.L_HI(net489));
 sg13g2_tiehi \dtop.player_inst.synth.alu.registers[4][4]$_SDFFE_PN0P__490  (.L_HI(net490));
 sg13g2_tiehi \dtop.player_inst.synth.alu.registers[4][5]$_SDFFE_PN0P__491  (.L_HI(net491));
 sg13g2_tiehi \dtop.player_inst.synth.alu.registers[4][6]$_SDFFE_PN0P__492  (.L_HI(net492));
 sg13g2_tiehi \dtop.player_inst.synth.alu.registers[4][7]$_SDFFE_PN0P__493  (.L_HI(net493));
 sg13g2_tiehi \dtop.player_inst.synth.alu.registers[4][8]$_SDFFE_PN0P__494  (.L_HI(net494));
 sg13g2_tiehi \dtop.player_inst.synth.alu.registers[4][9]$_SDFFE_PN0P__495  (.L_HI(net495));
 sg13g2_tiehi \dtop.player_inst.synth.alu.registers[5][0]$_SDFFE_PN0P__496  (.L_HI(net496));
 sg13g2_tiehi \dtop.player_inst.synth.alu.registers[5][1]$_SDFFE_PN0P__497  (.L_HI(net497));
 sg13g2_tiehi \dtop.player_inst.synth.alu.registers[5][2]$_SDFFE_PN0P__498  (.L_HI(net498));
 sg13g2_tiehi \dtop.player_inst.synth.alu.registers[5][3]$_SDFFE_PN0P__499  (.L_HI(net499));
 sg13g2_tiehi \dtop.player_inst.synth.alu.registers[5][4]$_SDFFE_PN0P__500  (.L_HI(net500));
 sg13g2_tiehi \dtop.player_inst.synth.alu.registers[5][5]$_SDFFE_PN0P__501  (.L_HI(net501));
 sg13g2_tiehi \dtop.player_inst.synth.alu.registers[5][6]$_SDFFE_PN0P__502  (.L_HI(net502));
 sg13g2_tiehi \dtop.player_inst.synth.alu.registers[6][0]$_SDFFE_PN0P__503  (.L_HI(net503));
 sg13g2_tiehi \dtop.player_inst.synth.alu.registers[6][1]$_SDFFE_PN0P__504  (.L_HI(net504));
 sg13g2_tiehi \dtop.player_inst.synth.alu.registers[6][2]$_SDFFE_PN0P__505  (.L_HI(net505));
 sg13g2_tiehi \dtop.player_inst.synth.alu.registers[6][3]$_SDFFE_PN0P__506  (.L_HI(net506));
 sg13g2_tiehi \dtop.player_inst.synth.alu.registers[6][4]$_SDFFE_PN0P__507  (.L_HI(net507));
 sg13g2_tiehi \dtop.player_inst.synth.alu.registers[6][5]$_SDFFE_PN0P__508  (.L_HI(net508));
 sg13g2_tiehi \dtop.player_inst.synth.alu.registers[6][6]$_SDFFE_PN0P__509  (.L_HI(net509));
 sg13g2_tiehi \dtop.vtop.dphases[0][0]$_DFFE_PP__510  (.L_HI(net510));
 sg13g2_tiehi \dtop.vtop.dphases[0][10]$_DFFE_PP__511  (.L_HI(net511));
 sg13g2_tiehi \dtop.vtop.dphases[0][1]$_DFFE_PP__512  (.L_HI(net512));
 sg13g2_tiehi \dtop.vtop.dphases[0][2]$_DFFE_PP__513  (.L_HI(net513));
 sg13g2_tiehi \dtop.vtop.dphases[0][3]$_DFFE_PP__514  (.L_HI(net514));
 sg13g2_tiehi \dtop.vtop.dphases[0][4]$_DFFE_PP__515  (.L_HI(net515));
 sg13g2_tiehi \dtop.vtop.dphases[0][5]$_DFFE_PP__516  (.L_HI(net516));
 sg13g2_tiehi \dtop.vtop.dphases[0][6]$_DFFE_PP__517  (.L_HI(net517));
 sg13g2_tiehi \dtop.vtop.dphases[0][7]$_DFFE_PP__518  (.L_HI(net518));
 sg13g2_tiehi \dtop.vtop.dphases[0][8]$_DFFE_PP__519  (.L_HI(net519));
 sg13g2_tiehi \dtop.vtop.dphases[0][9]$_DFFE_PP__520  (.L_HI(net520));
 sg13g2_tiehi \dtop.vtop.dphases[1][0]$_DFFE_PP__521  (.L_HI(net521));
 sg13g2_tiehi \dtop.vtop.dphases[1][10]$_DFFE_PP__522  (.L_HI(net522));
 sg13g2_tiehi \dtop.vtop.dphases[1][1]$_DFFE_PP__523  (.L_HI(net523));
 sg13g2_tiehi \dtop.vtop.dphases[1][2]$_DFFE_PP__524  (.L_HI(net524));
 sg13g2_tiehi \dtop.vtop.dphases[1][3]$_DFFE_PP__525  (.L_HI(net525));
 sg13g2_tiehi \dtop.vtop.dphases[1][4]$_DFFE_PP__526  (.L_HI(net526));
 sg13g2_tiehi \dtop.vtop.dphases[1][5]$_DFFE_PP__527  (.L_HI(net527));
 sg13g2_tiehi \dtop.vtop.dphases[1][6]$_DFFE_PP__528  (.L_HI(net528));
 sg13g2_tiehi \dtop.vtop.dphases[1][7]$_DFFE_PP__529  (.L_HI(net529));
 sg13g2_tiehi \dtop.vtop.dphases[1][8]$_DFFE_PP__530  (.L_HI(net530));
 sg13g2_tiehi \dtop.vtop.dphases[1][9]$_DFFE_PP__531  (.L_HI(net531));
 sg13g2_tiehi \dtop.vtop.dphases[2][0]$_DFFE_PP__532  (.L_HI(net532));
 sg13g2_tiehi \dtop.vtop.dphases[2][10]$_DFFE_PP__533  (.L_HI(net533));
 sg13g2_tiehi \dtop.vtop.dphases[2][1]$_DFFE_PP__534  (.L_HI(net534));
 sg13g2_tiehi \dtop.vtop.dphases[2][2]$_DFFE_PP__535  (.L_HI(net535));
 sg13g2_tiehi \dtop.vtop.dphases[2][3]$_DFFE_PP__536  (.L_HI(net536));
 sg13g2_tiehi \dtop.vtop.dphases[2][4]$_DFFE_PP__537  (.L_HI(net537));
 sg13g2_tiehi \dtop.vtop.dphases[2][5]$_DFFE_PP__538  (.L_HI(net538));
 sg13g2_tiehi \dtop.vtop.dphases[2][6]$_DFFE_PP__539  (.L_HI(net539));
 sg13g2_tiehi \dtop.vtop.dphases[2][7]$_DFFE_PP__540  (.L_HI(net540));
 sg13g2_tiehi \dtop.vtop.dphases[2][8]$_DFFE_PP__541  (.L_HI(net541));
 sg13g2_tiehi \dtop.vtop.dphases[2][9]$_DFFE_PP__542  (.L_HI(net542));
 sg13g2_tiehi \dtop.vtop.pipeline.cosappr[3]$_DFFE_PP__543  (.L_HI(net543));
 sg13g2_tiehi \dtop.vtop.pipeline.cosappr[4]$_DFFE_PP__544  (.L_HI(net544));
 sg13g2_tiehi \dtop.vtop.pipeline.cosappr[5]$_DFFE_PP__545  (.L_HI(net545));
 sg13g2_tiehi \dtop.vtop.pipeline.cosappr[6]$_DFFE_PP__546  (.L_HI(net546));
 sg13g2_tiehi \dtop.vtop.pipeline.cosappr[7]$_DFFE_PP__547  (.L_HI(net547));
 sg13g2_tiehi \dtop.vtop.pipeline.cosappr[8]$_DFFE_PP__548  (.L_HI(net548));
 sg13g2_tiehi \dtop.vtop.pipeline.cosappr_acc[0]$_DFFE_PN__549  (.L_HI(net549));
 sg13g2_tiehi \dtop.vtop.pipeline.cosappr_acc[1]$_DFFE_PN__550  (.L_HI(net550));
 sg13g2_tiehi \dtop.vtop.pipeline.cosappr_acc[2]$_DFFE_PN__551  (.L_HI(net551));
 sg13g2_tiehi \dtop.vtop.pipeline.cosappr_acc[3]$_DFFE_PN__552  (.L_HI(net552));
 sg13g2_tiehi \dtop.vtop.pipeline.cosappr_acc[4]$_DFFE_PN__553  (.L_HI(net553));
 sg13g2_tiehi \dtop.vtop.pipeline.cosappr_acc[5]$_DFFE_PN__554  (.L_HI(net554));
 sg13g2_tiehi \dtop.vtop.pipeline.cosappr_acc[6]$_DFFE_PN__555  (.L_HI(net555));
 sg13g2_tiehi \dtop.vtop.pipeline.cosappr_acc[7]$_DFFE_PN__556  (.L_HI(net556));
 sg13g2_tiehi \dtop.vtop.pipeline.cosappr_acc[8]$_DFFE_PN__557  (.L_HI(net557));
 sg13g2_tiehi \dtop.vtop.pipeline.dz[0]$_SDFFE_PP1P__558  (.L_HI(net558));
 sg13g2_tiehi \dtop.vtop.pipeline.dz[1]$_SDFFE_PP1P__559  (.L_HI(net559));
 sg13g2_tiehi \dtop.vtop.pipeline.dz[2]$_SDFFE_PP1P__560  (.L_HI(net560));
 sg13g2_tiehi \dtop.vtop.pipeline.dz[3]$_SDFFE_PP1P__561  (.L_HI(net561));
 sg13g2_tiehi \dtop.vtop.pipeline.dz[4]$_SDFFE_PP1P__562  (.L_HI(net562));
 sg13g2_tiehi \dtop.vtop.pipeline.dz[5]$_SDFFE_PP1P__563  (.L_HI(net563));
 sg13g2_tiehi \dtop.vtop.pipeline.dz[6]$_SDFFE_PP1P__564  (.L_HI(net564));
 sg13g2_tiehi \dtop.vtop.pipeline.dz[7]$_SDFFE_PP1P__565  (.L_HI(net565));
 sg13g2_tiehi \dtop.vtop.pipeline.dz[8]$_SDFFE_PP1P__566  (.L_HI(net566));
 sg13g2_tiehi \dtop.vtop.pipeline.neg_t[0]$_SDFFE_PP0P__567  (.L_HI(net567));
 sg13g2_tiehi \dtop.vtop.pipeline.neg_t[1]$_SDFFE_PP0P__568  (.L_HI(net568));
 sg13g2_tiehi \dtop.vtop.pipeline.neg_t[2]$_SDFFE_PP0P__569  (.L_HI(net569));
 sg13g2_tiehi \dtop.vtop.pipeline.neg_t[3]$_SDFFE_PP0P__570  (.L_HI(net570));
 sg13g2_tiehi \dtop.vtop.pipeline.neg_t[4]$_SDFFE_PP0P__571  (.L_HI(net571));
 sg13g2_tiehi \dtop.vtop.pipeline.neg_t[5]$_SDFFE_PP0P__572  (.L_HI(net572));
 sg13g2_tiehi \dtop.vtop.pipeline.neg_t[6]$_SDFFE_PP0P__573  (.L_HI(net573));
 sg13g2_tiehi \dtop.vtop.pipeline.neg_t[7]$_SDFFE_PP0P__574  (.L_HI(net574));
 sg13g2_tiehi \dtop.vtop.pipeline.neg_t[8]$_SDFFE_PP0P__575  (.L_HI(net575));
 sg13g2_tiehi \dtop.vtop.pipeline.neg_t[9]$_SDFFE_PP0P__576  (.L_HI(net576));
 sg13g2_tiehi \dtop.vtop.pipeline.nstep_counter[0]$_SDFFE_PP1P__577  (.L_HI(net577));
 sg13g2_tiehi \dtop.vtop.pipeline.nstep_counter[1]$_SDFFE_PP1P__578  (.L_HI(net578));
 sg13g2_tiehi \dtop.vtop.pipeline.nstep_counter[2]$_SDFFE_PP1P__579  (.L_HI(net579));
 sg13g2_tiehi \dtop.vtop.pipeline.nstep_counter[3]$_SDFFE_PP1P__580  (.L_HI(net580));
 sg13g2_tiehi \dtop.vtop.pipeline.nstep_counter[4]$_SDFFE_PP1P__581  (.L_HI(net581));
 sg13g2_tiehi \dtop.vtop.pipeline.nstep_reg[0]$_SDFF_PP0__582  (.L_HI(net582));
 sg13g2_tiehi \dtop.vtop.pipeline.nstep_reg[1]$_SDFF_PP0__583  (.L_HI(net583));
 sg13g2_tiehi \dtop.vtop.pipeline.nstep_zg[0]$_DFFE_PP__584  (.L_HI(net584));
 sg13g2_tiehi \dtop.vtop.pipeline.nstep_zg[1]$_DFFE_PP__585  (.L_HI(net585));
 sg13g2_tiehi \dtop.vtop.pipeline.phases[0][0]$_DFFE_PP__586  (.L_HI(net586));
 sg13g2_tiehi \dtop.vtop.pipeline.phases[0][10]$_DFFE_PP__587  (.L_HI(net587));
 sg13g2_tiehi \dtop.vtop.pipeline.phases[0][11]$_DFFE_PP__588  (.L_HI(net588));
 sg13g2_tiehi \dtop.vtop.pipeline.phases[0][12]$_DFFE_PP__589  (.L_HI(net589));
 sg13g2_tiehi \dtop.vtop.pipeline.phases[0][13]$_DFFE_PP__590  (.L_HI(net590));
 sg13g2_tiehi \dtop.vtop.pipeline.phases[0][14]$_DFFE_PP__591  (.L_HI(net591));
 sg13g2_tiehi \dtop.vtop.pipeline.phases[0][15]$_DFFE_PP__592  (.L_HI(net592));
 sg13g2_tiehi \dtop.vtop.pipeline.phases[0][1]$_DFFE_PP__593  (.L_HI(net593));
 sg13g2_tiehi \dtop.vtop.pipeline.phases[0][2]$_DFFE_PP__594  (.L_HI(net594));
 sg13g2_tiehi \dtop.vtop.pipeline.phases[0][3]$_DFFE_PP__595  (.L_HI(net595));
 sg13g2_tiehi \dtop.vtop.pipeline.phases[0][4]$_DFFE_PP__596  (.L_HI(net596));
 sg13g2_tiehi \dtop.vtop.pipeline.phases[0][5]$_DFFE_PP__597  (.L_HI(net597));
 sg13g2_tiehi \dtop.vtop.pipeline.phases[0][6]$_DFFE_PP__598  (.L_HI(net598));
 sg13g2_tiehi \dtop.vtop.pipeline.phases[0][7]$_DFFE_PP__599  (.L_HI(net599));
 sg13g2_tiehi \dtop.vtop.pipeline.phases[0][8]$_DFFE_PP__600  (.L_HI(net600));
 sg13g2_tiehi \dtop.vtop.pipeline.phases[0][9]$_DFFE_PP__601  (.L_HI(net601));
 sg13g2_tiehi \dtop.vtop.pipeline.phases[1][0]$_DFFE_PP__602  (.L_HI(net602));
 sg13g2_tiehi \dtop.vtop.pipeline.phases[1][10]$_DFFE_PP__603  (.L_HI(net603));
 sg13g2_tiehi \dtop.vtop.pipeline.phases[1][11]$_DFFE_PP__604  (.L_HI(net604));
 sg13g2_tiehi \dtop.vtop.pipeline.phases[1][12]$_DFFE_PP__605  (.L_HI(net605));
 sg13g2_tiehi \dtop.vtop.pipeline.phases[1][13]$_DFFE_PP__606  (.L_HI(net606));
 sg13g2_tiehi \dtop.vtop.pipeline.phases[1][14]$_DFFE_PP__607  (.L_HI(net607));
 sg13g2_tiehi \dtop.vtop.pipeline.phases[1][15]$_DFFE_PP__608  (.L_HI(net608));
 sg13g2_tiehi \dtop.vtop.pipeline.phases[1][1]$_DFFE_PP__609  (.L_HI(net609));
 sg13g2_tiehi \dtop.vtop.pipeline.phases[1][2]$_DFFE_PP__610  (.L_HI(net610));
 sg13g2_tiehi \dtop.vtop.pipeline.phases[1][3]$_DFFE_PP__611  (.L_HI(net611));
 sg13g2_tiehi \dtop.vtop.pipeline.phases[1][4]$_DFFE_PP__612  (.L_HI(net612));
 sg13g2_tiehi \dtop.vtop.pipeline.phases[1][5]$_DFFE_PP__613  (.L_HI(net613));
 sg13g2_tiehi \dtop.vtop.pipeline.phases[1][6]$_DFFE_PP__614  (.L_HI(net614));
 sg13g2_tiehi \dtop.vtop.pipeline.phases[1][7]$_DFFE_PP__615  (.L_HI(net615));
 sg13g2_tiehi \dtop.vtop.pipeline.phases[1][8]$_DFFE_PP__616  (.L_HI(net616));
 sg13g2_tiehi \dtop.vtop.pipeline.phases[1][9]$_DFFE_PP__617  (.L_HI(net617));
 sg13g2_tiehi \dtop.vtop.pipeline.phases[2][0]$_DFFE_PP__618  (.L_HI(net618));
 sg13g2_tiehi \dtop.vtop.pipeline.phases[2][10]$_DFFE_PP__619  (.L_HI(net619));
 sg13g2_tiehi \dtop.vtop.pipeline.phases[2][11]$_DFFE_PP__620  (.L_HI(net620));
 sg13g2_tiehi \dtop.vtop.pipeline.phases[2][12]$_DFFE_PP__621  (.L_HI(net621));
 sg13g2_tiehi \dtop.vtop.pipeline.phases[2][13]$_DFFE_PP__622  (.L_HI(net622));
 sg13g2_tiehi \dtop.vtop.pipeline.phases[2][14]$_DFFE_PP__623  (.L_HI(net623));
 sg13g2_tiehi \dtop.vtop.pipeline.phases[2][15]$_DFFE_PP__624  (.L_HI(net624));
 sg13g2_tiehi \dtop.vtop.pipeline.phases[2][1]$_DFFE_PP__625  (.L_HI(net625));
 sg13g2_tiehi \dtop.vtop.pipeline.phases[2][2]$_DFFE_PP__626  (.L_HI(net626));
 sg13g2_tiehi \dtop.vtop.pipeline.phases[2][3]$_DFFE_PP__627  (.L_HI(net627));
 sg13g2_tiehi \dtop.vtop.pipeline.phases[2][4]$_DFFE_PP__628  (.L_HI(net628));
 sg13g2_tiehi \dtop.vtop.pipeline.phases[2][5]$_DFFE_PP__629  (.L_HI(net629));
 sg13g2_tiehi \dtop.vtop.pipeline.phases[2][6]$_DFFE_PP__630  (.L_HI(net630));
 sg13g2_tiehi \dtop.vtop.pipeline.phases[2][7]$_DFFE_PP__631  (.L_HI(net631));
 sg13g2_tiehi \dtop.vtop.pipeline.phases[2][8]$_DFFE_PP__632  (.L_HI(net632));
 sg13g2_tiehi \dtop.vtop.pipeline.phases[2][9]$_DFFE_PP__633  (.L_HI(net633));
 sg13g2_tiehi \dtop.vtop.pipeline.wave_index[0]$_SDFF_PP0__634  (.L_HI(net634));
 sg13g2_tiehi \dtop.vtop.pipeline.wave_index[1]$_SDFF_PP0__635  (.L_HI(net635));
 sg13g2_tiehi \dtop.vtop.pipeline.z[0]$_SDFFE_PP0P__636  (.L_HI(net636));
 sg13g2_tiehi \dtop.vtop.pipeline.z[10]$_SDFFE_PP0P__637  (.L_HI(net637));
 sg13g2_tiehi \dtop.vtop.pipeline.z[11]$_SDFFE_PP0P__638  (.L_HI(net638));
 sg13g2_tiehi \dtop.vtop.pipeline.z[12]$_SDFFE_PP0P__639  (.L_HI(net639));
 sg13g2_tiehi \dtop.vtop.pipeline.z[13]$_SDFFE_PP0P__640  (.L_HI(net640));
 sg13g2_tiehi \dtop.vtop.pipeline.z[14]$_SDFFE_PP0P__641  (.L_HI(net641));
 sg13g2_tiehi \dtop.vtop.pipeline.z[1]$_SDFFE_PP0P__642  (.L_HI(net642));
 sg13g2_tiehi \dtop.vtop.pipeline.z[2]$_SDFFE_PP0P__643  (.L_HI(net643));
 sg13g2_tiehi \dtop.vtop.pipeline.z[3]$_SDFFE_PP0P__644  (.L_HI(net644));
 sg13g2_tiehi \dtop.vtop.pipeline.z[4]$_SDFFE_PP0P__645  (.L_HI(net645));
 sg13g2_tiehi \dtop.vtop.pipeline.z[5]$_SDFFE_PP0P__646  (.L_HI(net646));
 sg13g2_tiehi \dtop.vtop.pipeline.z[6]$_SDFFE_PP0P__647  (.L_HI(net647));
 sg13g2_tiehi \dtop.vtop.pipeline.z[7]$_SDFFE_PP0P__648  (.L_HI(net648));
 sg13g2_tiehi \dtop.vtop.pipeline.z[8]$_SDFFE_PP0P__649  (.L_HI(net649));
 sg13g2_tiehi \dtop.vtop.pipeline.z[9]$_SDFFE_PP0P__650  (.L_HI(net650));
 sg13g2_tiehi \dtop.vtop.pipeline.zg[0]$_DFFE_PP__651  (.L_HI(net651));
 sg13g2_tiehi \dtop.vtop.pipeline.zg[1]$_DFFE_PP__652  (.L_HI(net652));
 sg13g2_tiehi \dtop.vtop.pipeline.zg[2]$_DFFE_PP__653  (.L_HI(net653));
 sg13g2_tiehi \dtop.vtop.pipeline.zg[3]$_DFFE_PP__654  (.L_HI(net654));
 sg13g2_tiehi \dtop.vtop.pipeline.zg[4]$_DFFE_PP__655  (.L_HI(net655));
 sg13g2_tiehi \dtop.vtop.pipeline.zg[5]$_DFFE_PP__656  (.L_HI(net656));
 sg13g2_tiehi \dtop.vtop.pipeline.zg[6]$_DFFE_PP__657  (.L_HI(net657));
 sg13g2_tiehi \dtop.vtop.pipeline.zg[7]$_DFFE_PP__658  (.L_HI(net658));
 sg13g2_tiehi \dtop.vtop.pipeline.zg[8]$_DFFE_PP__659  (.L_HI(net659));
 sg13g2_tiehi \dtop.vtop.pipeline.zg[9]$_DFFE_PP__660  (.L_HI(net660));
 sg13g2_tiehi \dtop.vtop.pipeline.zg_acc[0]$_DFFE_PN__661  (.L_HI(net661));
 sg13g2_tiehi \dtop.vtop.pipeline.zg_acc[1]$_DFFE_PN__662  (.L_HI(net662));
 sg13g2_tiehi \dtop.vtop.pipeline.zg_acc[2]$_DFFE_PN__663  (.L_HI(net663));
 sg13g2_tiehi \dtop.vtop.pipeline.zg_acc[3]$_DFFE_PN__664  (.L_HI(net664));
 sg13g2_tiehi \dtop.vtop.pipeline.zg_acc[4]$_DFFE_PN__665  (.L_HI(net665));
 sg13g2_tiehi \dtop.vtop.pipeline.zg_acc[5]$_DFFE_PN__666  (.L_HI(net666));
 sg13g2_tiehi \dtop.vtop.pipeline.zg_acc[6]$_DFFE_PN__667  (.L_HI(net667));
 sg13g2_tiehi \dtop.vtop.pipeline.zg_acc[7]$_DFFE_PN__668  (.L_HI(net668));
 sg13g2_tiehi \dtop.vtop.pipeline.zg_acc[8]$_DFFE_PN__669  (.L_HI(net669));
 sg13g2_tiehi \dtop.vtop.pipeline.zg_acc[9]$_DFFE_PN__670  (.L_HI(net670));
 sg13g2_tiehi \dtop.vtop.pipeline.zg_valid$_SDFFE_PP0P__671  (.L_HI(net671));
 sg13g2_tiehi \dtop.vtop.r_frame_counter[0]$_SDFF_PP0__672  (.L_HI(net672));
 sg13g2_tiehi \dtop.vtop.r_frame_counter[10]$_SDFF_PP0__673  (.L_HI(net673));
 sg13g2_tiehi \dtop.vtop.r_frame_counter[11]$_SDFF_PP0__674  (.L_HI(net674));
 sg13g2_tiehi \dtop.vtop.r_frame_counter[12]$_SDFF_PP0__675  (.L_HI(net675));
 sg13g2_tiehi \dtop.vtop.r_frame_counter[13]$_SDFF_PP0__676  (.L_HI(net676));
 sg13g2_tiehi \dtop.vtop.r_frame_counter[1]$_SDFF_PP0__677  (.L_HI(net677));
 sg13g2_tiehi \dtop.vtop.r_frame_counter[2]$_SDFF_PP0__678  (.L_HI(net678));
 sg13g2_tiehi \dtop.vtop.r_frame_counter[3]$_SDFF_PP0__679  (.L_HI(net679));
 sg13g2_tiehi \dtop.vtop.r_frame_counter[4]$_SDFF_PP0__680  (.L_HI(net680));
 sg13g2_tiehi \dtop.vtop.r_frame_counter[5]$_SDFF_PP0__681  (.L_HI(net681));
 sg13g2_tiehi \dtop.vtop.r_frame_counter[6]$_SDFF_PP0__682  (.L_HI(net682));
 sg13g2_tiehi \dtop.vtop.r_frame_counter[7]$_SDFF_PP0__683  (.L_HI(net683));
 sg13g2_tiehi \dtop.vtop.r_frame_counter[8]$_SDFF_PP0__684  (.L_HI(net684));
 sg13g2_tiehi \dtop.vtop.r_frame_counter[9]$_SDFF_PP0__685  (.L_HI(net685));
 sg13g2_tiehi \dtop.vtop.rs.r_vsync$_DFFE_PP__686  (.L_HI(net686));
 sg13g2_tiehi \dtop.vtop.rs.scan_y.phase[0]$_SDFF_PN0__687  (.L_HI(net687));
 sg13g2_tiehi \dtop.vtop.rs.scan_y.phase[1]$_SDFF_PN0__688  (.L_HI(net688));
 sg13g2_tiehi \dtop.vtop.rs.scan_y.y[0]$_SDFF_PP0__689  (.L_HI(net689));
 sg13g2_tiehi \dtop.vtop.rs.scan_y.y[1]$_SDFF_PP0__690  (.L_HI(net690));
 sg13g2_tiehi \dtop.vtop.rs.scan_y.y[2]$_SDFF_PP0__691  (.L_HI(net691));
 sg13g2_tiehi \dtop.vtop.rs.scan_y.y[3]$_SDFF_PP0__692  (.L_HI(net692));
 sg13g2_tiehi \dtop.vtop.rs.scan_y.y[4]$_SDFF_PP0__693  (.L_HI(net693));
 sg13g2_tiehi \dtop.vtop.rs.scan_y.y[5]$_SDFF_PP0__694  (.L_HI(net694));
 sg13g2_tiehi \dtop.vtop.rs.scan_y.y[6]$_SDFF_PP0__695  (.L_HI(net695));
 sg13g2_tiehi \dtop.vtop.rs.scan_y.y[7]$_SDFF_PP0__696  (.L_HI(net696));
 sg13g2_tiehi \dtop.vtop.rs.scan_y.y[8]$_SDFF_PP0__697  (.L_HI(net697));
 sg13g2_tiehi \dtop.vtop.rs.scan_y.y[9]$_SDFF_PN0__698  (.L_HI(net698));
 sg13g2_tiehi \dtop.vtop.rs.x_scan.phase[0]$_SDFF_PN0__699  (.L_HI(net699));
 sg13g2_tiehi \dtop.vtop.rs.x_scan.phase[1]$_SDFF_PN1__700  (.L_HI(net700));
 sg13g2_tiehi \dtop.vtop.rs.x_scan.r_coarse[0]$_SDFF_PN0__701  (.L_HI(net701));
 sg13g2_tiehi \dtop.vtop.rs.x_scan.r_coarse[1]$_SDFF_PN0__702  (.L_HI(net702));
 sg13g2_tiehi \dtop.vtop.rs.x_scan.r_coarse[2]$_SDFF_PN0__703  (.L_HI(net703));
 sg13g2_tiehi \dtop.vtop.rs.x_scan.r_fine[0]$_SDFF_PP0__704  (.L_HI(net704));
 sg13g2_tiehi \dtop.vtop.rs.x_scan.r_fine[1]$_SDFF_PP0__705  (.L_HI(net705));
 sg13g2_tiehi \dtop.vtop.rs.x_scan.r_fine[2]$_SDFF_PP0__706  (.L_HI(net706));
 sg13g2_tiehi \dtop.vtop.rs.x_scan.r_fine[3]$_SDFF_PP0__707  (.L_HI(net707));
 sg13g2_tiehi \dtop.vtop.rs.x_scan.r_fine[4]$_SDFF_PP0__708  (.L_HI(net708));
 sg13g2_tiehi \dtop.vtop.rs.x_scan.r_fine[5]$_SDFF_PP0__709  (.L_HI(net709));
 sg13g2_tiehi \dtop.vtop.rs.x_scan.r_fine[6]$_SDFF_PP0__710  (.L_HI(net710));
 sg13g2_tiehi \dtop.vtop.xfrac_counter$_SDFF_PN0__711  (.L_HI(net711));
 sg13g2_tiehi \rst_n_reg$_DFF_P__712  (.L_HI(net712));
 sg13g2_tiehi \ui_in_reg[0]$_DFF_P__713  (.L_HI(net713));
 sg13g2_tiehi \ui_in_reg[1]$_DFF_P__714  (.L_HI(net714));
 sg13g2_tiehi \ui_in_reg[2]$_DFF_P__715  (.L_HI(net715));
 sg13g2_tiehi \ui_in_reg[3]$_DFF_P__716  (.L_HI(net716));
 sg13g2_tiehi \ui_in_reg[4]$_DFF_P__717  (.L_HI(net717));
 sg13g2_tiehi \ui_in_reg[5]$_DFF_P__718  (.L_HI(net718));
 sg13g2_tiehi \ui_in_reg[6]$_DFF_P__719  (.L_HI(net719));
 sg13g2_tiehi \ui_in_reg[7]$_DFF_P__720  (.L_HI(net720));
 sg13g2_tiehi \uio_oe1[4]$_DFFE_PP__721  (.L_HI(net721));
 sg13g2_tiehi \uio_out1[0]$_SDFFCE_PN0P__722  (.L_HI(net722));
 sg13g2_tiehi \uio_out1[1]$_SDFFCE_PN0P__723  (.L_HI(net723));
 sg13g2_tiehi \uio_out1[2]$_SDFFCE_PN0P__724  (.L_HI(net724));
 sg13g2_tiehi \uio_out1[3]$_SDFFCE_PN0P__725  (.L_HI(net725));
 sg13g2_tiehi \uio_out1[4]$_SDFFCE_PN0P__726  (.L_HI(net726));
 sg13g2_tiehi \uio_out1[5]$_SDFFCE_PN0P__727  (.L_HI(net727));
 sg13g2_tiehi \uio_out1[6]$_DFFE_PP__728  (.L_HI(net728));
 sg13g2_tiehi \uio_out1[7]$_DFFE_PP__729  (.L_HI(net729));
 sg13g2_tiehi \uo_out1[0]$_DFFE_PP__730  (.L_HI(net730));
 sg13g2_tiehi \uo_out1[1]$_DFFE_PP__731  (.L_HI(net731));
 sg13g2_tiehi \uo_out1[2]$_DFFE_PP__732  (.L_HI(net732));
 sg13g2_tiehi \uo_out1[3]$_DFFE_PP__733  (.L_HI(net733));
 sg13g2_tiehi \uo_out1[4]$_DFFE_PP__734  (.L_HI(net734));
 sg13g2_tiehi \uo_out1[5]$_DFFE_PP__735  (.L_HI(net735));
 sg13g2_tiehi \uo_out1[6]$_DFFE_PP__736  (.L_HI(net736));
 sg13g2_tiehi \uo_out1[7]$_DFFE_PP__737  (.L_HI(net737));
 sg13g2_buf_4 clkbuf_leaf_1_clk (.X(clknet_leaf_1_clk),
    .A(clknet_4_1_0_clk));
 sg13g2_buf_4 clkbuf_leaf_2_clk (.X(clknet_leaf_2_clk),
    .A(clknet_4_1_0_clk));
 sg13g2_buf_4 clkbuf_leaf_3_clk (.X(clknet_leaf_3_clk),
    .A(clknet_4_4_0_clk));
 sg13g2_buf_4 clkbuf_leaf_4_clk (.X(clknet_leaf_4_clk),
    .A(clknet_4_4_0_clk));
 sg13g2_buf_4 clkbuf_leaf_5_clk (.X(clknet_leaf_5_clk),
    .A(clknet_4_4_0_clk));
 sg13g2_buf_4 clkbuf_leaf_6_clk (.X(clknet_leaf_6_clk),
    .A(clknet_4_4_0_clk));
 sg13g2_buf_4 clkbuf_leaf_7_clk (.X(clknet_leaf_7_clk),
    .A(clknet_4_6_0_clk));
 sg13g2_buf_4 clkbuf_leaf_8_clk (.X(clknet_leaf_8_clk),
    .A(clknet_4_6_0_clk));
 sg13g2_buf_4 clkbuf_leaf_10_clk (.X(clknet_leaf_10_clk),
    .A(clknet_4_9_0_clk));
 sg13g2_buf_4 clkbuf_leaf_11_clk (.X(clknet_leaf_11_clk),
    .A(clknet_4_7_0_clk));
 sg13g2_buf_4 clkbuf_leaf_12_clk (.X(clknet_leaf_12_clk),
    .A(clknet_4_5_0_clk));
 sg13g2_buf_4 clkbuf_leaf_13_clk (.X(clknet_leaf_13_clk),
    .A(clknet_4_5_0_clk));
 sg13g2_buf_4 clkbuf_leaf_14_clk (.X(clknet_leaf_14_clk),
    .A(clknet_4_5_0_clk));
 sg13g2_buf_4 clkbuf_leaf_15_clk (.X(clknet_leaf_15_clk),
    .A(clknet_4_7_0_clk));
 sg13g2_buf_4 clkbuf_leaf_16_clk (.X(clknet_leaf_16_clk),
    .A(clknet_4_7_0_clk));
 sg13g2_buf_4 clkbuf_leaf_17_clk (.X(clknet_leaf_17_clk),
    .A(clknet_4_13_0_clk));
 sg13g2_buf_4 clkbuf_leaf_18_clk (.X(clknet_leaf_18_clk),
    .A(clknet_4_13_0_clk));
 sg13g2_buf_4 clkbuf_leaf_19_clk (.X(clknet_leaf_19_clk),
    .A(clknet_4_12_0_clk));
 sg13g2_buf_4 clkbuf_leaf_20_clk (.X(clknet_leaf_20_clk),
    .A(clknet_4_12_0_clk));
 sg13g2_buf_4 clkbuf_leaf_21_clk (.X(clknet_leaf_21_clk),
    .A(clknet_4_12_0_clk));
 sg13g2_buf_4 clkbuf_leaf_22_clk (.X(clknet_leaf_22_clk),
    .A(clknet_4_9_0_clk));
 sg13g2_buf_4 clkbuf_leaf_23_clk (.X(clknet_leaf_23_clk),
    .A(clknet_4_9_0_clk));
 sg13g2_buf_4 clkbuf_leaf_24_clk (.X(clknet_leaf_24_clk),
    .A(clknet_4_12_0_clk));
 sg13g2_buf_4 clkbuf_leaf_26_clk (.X(clknet_leaf_26_clk),
    .A(clknet_4_14_0_clk));
 sg13g2_buf_4 clkbuf_leaf_27_clk (.X(clknet_leaf_27_clk),
    .A(clknet_4_15_0_clk));
 sg13g2_buf_4 clkbuf_leaf_28_clk (.X(clknet_leaf_28_clk),
    .A(clknet_4_15_0_clk));
 sg13g2_buf_4 clkbuf_leaf_29_clk (.X(clknet_leaf_29_clk),
    .A(clknet_4_15_0_clk));
 sg13g2_buf_4 clkbuf_leaf_30_clk (.X(clknet_leaf_30_clk),
    .A(clknet_4_14_0_clk));
 sg13g2_buf_4 clkbuf_leaf_31_clk (.X(clknet_leaf_31_clk),
    .A(clknet_4_14_0_clk));
 sg13g2_buf_4 clkbuf_leaf_33_clk (.X(clknet_leaf_33_clk),
    .A(clknet_4_14_0_clk));
 sg13g2_buf_4 clkbuf_leaf_34_clk (.X(clknet_leaf_34_clk),
    .A(clknet_4_11_0_clk));
 sg13g2_buf_4 clkbuf_leaf_36_clk (.X(clknet_leaf_36_clk),
    .A(clknet_4_9_0_clk));
 sg13g2_buf_4 clkbuf_leaf_37_clk (.X(clknet_leaf_37_clk),
    .A(clknet_4_8_0_clk));
 sg13g2_buf_4 clkbuf_leaf_38_clk (.X(clknet_leaf_38_clk),
    .A(clknet_4_8_0_clk));
 sg13g2_buf_4 clkbuf_leaf_39_clk (.X(clknet_leaf_39_clk),
    .A(clknet_4_10_0_clk));
 sg13g2_buf_4 clkbuf_leaf_40_clk (.X(clknet_leaf_40_clk),
    .A(clknet_4_10_0_clk));
 sg13g2_buf_4 clkbuf_leaf_41_clk (.X(clknet_leaf_41_clk),
    .A(clknet_4_10_0_clk));
 sg13g2_buf_4 clkbuf_leaf_42_clk (.X(clknet_leaf_42_clk),
    .A(clknet_4_10_0_clk));
 sg13g2_buf_4 clkbuf_leaf_44_clk (.X(clknet_leaf_44_clk),
    .A(clknet_4_8_0_clk));
 sg13g2_buf_4 clkbuf_leaf_45_clk (.X(clknet_leaf_45_clk),
    .A(clknet_4_8_0_clk));
 sg13g2_buf_4 clkbuf_leaf_46_clk (.X(clknet_leaf_46_clk),
    .A(clknet_4_3_0_clk));
 sg13g2_buf_4 clkbuf_leaf_47_clk (.X(clknet_leaf_47_clk),
    .A(clknet_4_3_0_clk));
 sg13g2_buf_4 clkbuf_leaf_48_clk (.X(clknet_leaf_48_clk),
    .A(clknet_4_1_0_clk));
 sg13g2_buf_4 clkbuf_leaf_49_clk (.X(clknet_leaf_49_clk),
    .A(clknet_4_3_0_clk));
 sg13g2_buf_4 clkbuf_leaf_50_clk (.X(clknet_leaf_50_clk),
    .A(clknet_4_2_0_clk));
 sg13g2_buf_4 clkbuf_leaf_51_clk (.X(clknet_leaf_51_clk),
    .A(clknet_4_2_0_clk));
 sg13g2_buf_4 clkbuf_leaf_52_clk (.X(clknet_leaf_52_clk),
    .A(clknet_4_2_0_clk));
 sg13g2_buf_4 clkbuf_leaf_53_clk (.X(clknet_leaf_53_clk),
    .A(clknet_4_1_0_clk));
 sg13g2_buf_4 clkbuf_leaf_55_clk (.X(clknet_leaf_55_clk),
    .A(clknet_4_0_0_clk));
 sg13g2_buf_4 clkbuf_leaf_56_clk (.X(clknet_leaf_56_clk),
    .A(clknet_4_0_0_clk));
 sg13g2_buf_4 clkbuf_leaf_57_clk (.X(clknet_leaf_57_clk),
    .A(clknet_4_0_0_clk));
 sg13g2_buf_2 clkbuf_0_clk (.A(clk),
    .X(clknet_0_clk));
 sg13g2_buf_4 clkbuf_4_0_0_clk (.X(clknet_4_0_0_clk),
    .A(clknet_0_clk));
 sg13g2_buf_4 clkbuf_4_1_0_clk (.X(clknet_4_1_0_clk),
    .A(clknet_0_clk));
 sg13g2_buf_4 clkbuf_4_2_0_clk (.X(clknet_4_2_0_clk),
    .A(clknet_0_clk));
 sg13g2_buf_4 clkbuf_4_3_0_clk (.X(clknet_4_3_0_clk),
    .A(clknet_0_clk));
 sg13g2_buf_4 clkbuf_4_4_0_clk (.X(clknet_4_4_0_clk),
    .A(clknet_0_clk));
 sg13g2_buf_4 clkbuf_4_5_0_clk (.X(clknet_4_5_0_clk),
    .A(clknet_0_clk));
 sg13g2_buf_4 clkbuf_4_6_0_clk (.X(clknet_4_6_0_clk),
    .A(clknet_0_clk));
 sg13g2_buf_4 clkbuf_4_7_0_clk (.X(clknet_4_7_0_clk),
    .A(clknet_0_clk));
 sg13g2_buf_4 clkbuf_4_8_0_clk (.X(clknet_4_8_0_clk),
    .A(clknet_0_clk));
 sg13g2_buf_4 clkbuf_4_9_0_clk (.X(clknet_4_9_0_clk),
    .A(clknet_0_clk));
 sg13g2_buf_4 clkbuf_4_10_0_clk (.X(clknet_4_10_0_clk),
    .A(clknet_0_clk));
 sg13g2_buf_4 clkbuf_4_11_0_clk (.X(clknet_4_11_0_clk),
    .A(clknet_0_clk));
 sg13g2_buf_4 clkbuf_4_12_0_clk (.X(clknet_4_12_0_clk),
    .A(clknet_0_clk));
 sg13g2_buf_4 clkbuf_4_13_0_clk (.X(clknet_4_13_0_clk),
    .A(clknet_0_clk));
 sg13g2_buf_4 clkbuf_4_14_0_clk (.X(clknet_4_14_0_clk),
    .A(clknet_0_clk));
 sg13g2_buf_4 clkbuf_4_15_0_clk (.X(clknet_4_15_0_clk),
    .A(clknet_0_clk));
 sg13g2_buf_1 clkload0 (.A(clknet_4_2_0_clk));
 sg13g2_buf_4 clkload1 (.A(clknet_4_3_0_clk));
 sg13g2_buf_4 clkload2 (.A(clknet_4_5_0_clk));
 sg13g2_buf_1 clkload3 (.A(clknet_4_6_0_clk));
 sg13g2_buf_4 clkload4 (.A(clknet_4_7_0_clk));
 sg13g2_inv_2 clkload5 (.A(clknet_4_11_0_clk));
 sg13g2_inv_2 clkload6 (.A(clknet_4_13_0_clk));
 sg13g2_buf_4 clkload7 (.A(clknet_4_15_0_clk));
 sg13g2_inv_2 clkload8 (.A(clknet_leaf_0_clk));
 sg13g2_inv_1 clkload9 (.A(clknet_leaf_57_clk));
 sg13g2_inv_4 clkload10 (.A(clknet_leaf_1_clk));
 sg13g2_inv_1 clkload11 (.A(clknet_leaf_2_clk));
 sg13g2_inv_1 clkload12 (.A(clknet_leaf_48_clk));
 sg13g2_inv_2 clkload13 (.A(clknet_leaf_50_clk));
 sg13g2_buf_8 clkload14 (.A(clknet_leaf_51_clk));
 sg13g2_inv_2 clkload15 (.A(clknet_leaf_46_clk));
 sg13g2_inv_1 clkload16 (.A(clknet_leaf_47_clk));
 sg13g2_inv_1 clkload17 (.A(clknet_leaf_4_clk));
 sg13g2_inv_1 clkload18 (.A(clknet_leaf_5_clk));
 sg13g2_inv_1 clkload19 (.A(clknet_leaf_14_clk));
 sg13g2_buf_8 clkload20 (.A(clknet_leaf_8_clk));
 sg13g2_inv_4 clkload21 (.A(clknet_leaf_11_clk));
 sg13g2_buf_8 clkload22 (.A(clknet_leaf_15_clk));
 sg13g2_buf_8 clkload23 (.A(clknet_leaf_38_clk));
 sg13g2_buf_8 clkload24 (.A(clknet_leaf_45_clk));
 sg13g2_buf_16 clkload25 (.A(clknet_leaf_22_clk));
 sg13g2_buf_16 clkload26 (.A(clknet_leaf_23_clk));
 sg13g2_inv_2 clkload27 (.A(clknet_leaf_36_clk));
 sg13g2_inv_2 clkload28 (.A(clknet_leaf_40_clk));
 sg13g2_inv_4 clkload29 (.A(clknet_leaf_41_clk));
 sg13g2_inv_1 clkload30 (.A(clknet_leaf_42_clk));
 sg13g2_buf_8 clkload31 (.A(clknet_leaf_19_clk));
 sg13g2_inv_2 clkload32 (.A(clknet_leaf_20_clk));
 sg13g2_inv_4 clkload33 (.A(clknet_leaf_21_clk));
 sg13g2_inv_2 clkload34 (.A(clknet_leaf_26_clk));
 sg13g2_inv_1 clkload35 (.A(clknet_leaf_31_clk));
 sg13g2_antennanp ANTENNA_1 (.A(_02381_));
 sg13g2_antennanp ANTENNA_2 (.A(_02381_));
 sg13g2_antennanp ANTENNA_3 (.A(_02381_));
 sg13g2_antennanp ANTENNA_4 (.A(_05346_));
 sg13g2_antennanp ANTENNA_5 (.A(_05346_));
 sg13g2_antennanp ANTENNA_6 (.A(_05346_));
 sg13g2_antennanp ANTENNA_7 (.A(_05376_));
 sg13g2_antennanp ANTENNA_8 (.A(_05376_));
 sg13g2_antennanp ANTENNA_9 (.A(_05376_));
 sg13g2_antennanp ANTENNA_10 (.A(_05376_));
 sg13g2_antennanp ANTENNA_11 (.A(_05376_));
 sg13g2_antennanp ANTENNA_12 (.A(_05376_));
 sg13g2_antennanp ANTENNA_13 (.A(_05376_));
 sg13g2_antennanp ANTENNA_14 (.A(net6));
 sg13g2_antennanp ANTENNA_15 (.A(net332));
 sg13g2_antennanp ANTENNA_16 (.A(net332));
 sg13g2_antennanp ANTENNA_17 (.A(net332));
 sg13g2_antennanp ANTENNA_18 (.A(net332));
 sg13g2_antennanp ANTENNA_19 (.A(net332));
 sg13g2_antennanp ANTENNA_20 (.A(net332));
 sg13g2_antennanp ANTENNA_21 (.A(net332));
 sg13g2_antennanp ANTENNA_22 (.A(net332));
 sg13g2_antennanp ANTENNA_23 (.A(_05346_));
 sg13g2_antennanp ANTENNA_24 (.A(_05346_));
 sg13g2_antennanp ANTENNA_25 (.A(_05346_));
 sg13g2_antennanp ANTENNA_26 (.A(net6));
 sg13g2_antennanp ANTENNA_27 (.A(net332));
 sg13g2_antennanp ANTENNA_28 (.A(net332));
 sg13g2_antennanp ANTENNA_29 (.A(net332));
 sg13g2_antennanp ANTENNA_30 (.A(net332));
 sg13g2_antennanp ANTENNA_31 (.A(net332));
 sg13g2_antennanp ANTENNA_32 (.A(net332));
 sg13g2_antennanp ANTENNA_33 (.A(net332));
 sg13g2_antennanp ANTENNA_34 (.A(net332));
 sg13g2_antennanp ANTENNA_35 (.A(net6));
 sg13g2_antennanp ANTENNA_36 (.A(net332));
 sg13g2_antennanp ANTENNA_37 (.A(net332));
 sg13g2_antennanp ANTENNA_38 (.A(net332));
 sg13g2_antennanp ANTENNA_39 (.A(net332));
 sg13g2_antennanp ANTENNA_40 (.A(net332));
 sg13g2_antennanp ANTENNA_41 (.A(net332));
 sg13g2_antennanp ANTENNA_42 (.A(net332));
 sg13g2_antennanp ANTENNA_43 (.A(net332));
 sg13g2_antennanp ANTENNA_44 (.A(net332));
 sg13g2_antennanp ANTENNA_45 (.A(net6));
 sg13g2_antennanp ANTENNA_46 (.A(net332));
 sg13g2_antennanp ANTENNA_47 (.A(net332));
 sg13g2_antennanp ANTENNA_48 (.A(net332));
 sg13g2_antennanp ANTENNA_49 (.A(net332));
 sg13g2_antennanp ANTENNA_50 (.A(net332));
 sg13g2_antennanp ANTENNA_51 (.A(net332));
 sg13g2_antennanp ANTENNA_52 (.A(net332));
 sg13g2_antennanp ANTENNA_53 (.A(net332));
 sg13g2_antennanp ANTENNA_54 (.A(net332));
 sg13g2_antennanp ANTENNA_55 (.A(net6));
 sg13g2_antennanp ANTENNA_56 (.A(net332));
 sg13g2_antennanp ANTENNA_57 (.A(net332));
 sg13g2_antennanp ANTENNA_58 (.A(net332));
 sg13g2_antennanp ANTENNA_59 (.A(net332));
 sg13g2_antennanp ANTENNA_60 (.A(net332));
 sg13g2_antennanp ANTENNA_61 (.A(net332));
 sg13g2_antennanp ANTENNA_62 (.A(net332));
 sg13g2_antennanp ANTENNA_63 (.A(net332));
 sg13g2_antennanp ANTENNA_64 (.A(net332));
 sg13g2_decap_8 FILLER_0_0 ();
 sg13g2_decap_8 FILLER_0_7 ();
 sg13g2_decap_8 FILLER_0_14 ();
 sg13g2_decap_8 FILLER_0_21 ();
 sg13g2_decap_8 FILLER_0_28 ();
 sg13g2_decap_8 FILLER_0_35 ();
 sg13g2_decap_8 FILLER_0_42 ();
 sg13g2_decap_8 FILLER_0_49 ();
 sg13g2_decap_8 FILLER_0_56 ();
 sg13g2_decap_8 FILLER_0_63 ();
 sg13g2_decap_8 FILLER_0_70 ();
 sg13g2_decap_8 FILLER_0_77 ();
 sg13g2_decap_8 FILLER_0_84 ();
 sg13g2_decap_8 FILLER_0_91 ();
 sg13g2_decap_8 FILLER_0_98 ();
 sg13g2_decap_8 FILLER_0_105 ();
 sg13g2_decap_4 FILLER_0_112 ();
 sg13g2_fill_1 FILLER_0_116 ();
 sg13g2_fill_2 FILLER_0_146 ();
 sg13g2_fill_1 FILLER_0_148 ();
 sg13g2_fill_2 FILLER_0_158 ();
 sg13g2_fill_1 FILLER_0_160 ();
 sg13g2_decap_8 FILLER_0_175 ();
 sg13g2_decap_8 FILLER_0_182 ();
 sg13g2_decap_8 FILLER_0_189 ();
 sg13g2_decap_8 FILLER_0_196 ();
 sg13g2_decap_8 FILLER_0_233 ();
 sg13g2_fill_2 FILLER_0_240 ();
 sg13g2_fill_2 FILLER_0_272 ();
 sg13g2_fill_1 FILLER_0_274 ();
 sg13g2_decap_8 FILLER_0_280 ();
 sg13g2_fill_1 FILLER_0_287 ();
 sg13g2_fill_1 FILLER_0_293 ();
 sg13g2_decap_8 FILLER_0_302 ();
 sg13g2_decap_4 FILLER_0_309 ();
 sg13g2_fill_2 FILLER_0_313 ();
 sg13g2_decap_8 FILLER_0_319 ();
 sg13g2_decap_4 FILLER_0_326 ();
 sg13g2_fill_2 FILLER_0_330 ();
 sg13g2_decap_8 FILLER_0_341 ();
 sg13g2_decap_4 FILLER_0_348 ();
 sg13g2_fill_1 FILLER_0_352 ();
 sg13g2_fill_1 FILLER_0_396 ();
 sg13g2_decap_8 FILLER_0_423 ();
 sg13g2_decap_8 FILLER_0_430 ();
 sg13g2_fill_2 FILLER_0_437 ();
 sg13g2_decap_8 FILLER_0_443 ();
 sg13g2_decap_8 FILLER_0_450 ();
 sg13g2_decap_8 FILLER_0_457 ();
 sg13g2_decap_8 FILLER_0_464 ();
 sg13g2_decap_8 FILLER_0_471 ();
 sg13g2_decap_8 FILLER_0_478 ();
 sg13g2_decap_8 FILLER_0_485 ();
 sg13g2_decap_8 FILLER_0_492 ();
 sg13g2_decap_8 FILLER_0_499 ();
 sg13g2_decap_8 FILLER_0_506 ();
 sg13g2_decap_8 FILLER_0_513 ();
 sg13g2_decap_8 FILLER_0_520 ();
 sg13g2_decap_8 FILLER_0_527 ();
 sg13g2_decap_4 FILLER_0_534 ();
 sg13g2_decap_8 FILLER_0_551 ();
 sg13g2_decap_8 FILLER_0_558 ();
 sg13g2_decap_8 FILLER_0_565 ();
 sg13g2_decap_8 FILLER_0_572 ();
 sg13g2_decap_8 FILLER_0_579 ();
 sg13g2_decap_4 FILLER_0_586 ();
 sg13g2_fill_2 FILLER_0_590 ();
 sg13g2_decap_8 FILLER_0_604 ();
 sg13g2_decap_8 FILLER_0_611 ();
 sg13g2_decap_8 FILLER_0_618 ();
 sg13g2_decap_8 FILLER_0_625 ();
 sg13g2_fill_2 FILLER_0_632 ();
 sg13g2_decap_8 FILLER_0_643 ();
 sg13g2_decap_8 FILLER_0_650 ();
 sg13g2_decap_8 FILLER_0_657 ();
 sg13g2_decap_8 FILLER_0_664 ();
 sg13g2_decap_8 FILLER_0_671 ();
 sg13g2_decap_4 FILLER_0_678 ();
 sg13g2_fill_2 FILLER_0_682 ();
 sg13g2_decap_8 FILLER_0_689 ();
 sg13g2_decap_8 FILLER_0_696 ();
 sg13g2_decap_8 FILLER_0_703 ();
 sg13g2_decap_8 FILLER_0_710 ();
 sg13g2_decap_8 FILLER_0_722 ();
 sg13g2_decap_8 FILLER_0_768 ();
 sg13g2_decap_8 FILLER_0_775 ();
 sg13g2_decap_8 FILLER_0_782 ();
 sg13g2_decap_8 FILLER_0_789 ();
 sg13g2_decap_8 FILLER_0_796 ();
 sg13g2_decap_8 FILLER_0_803 ();
 sg13g2_decap_8 FILLER_0_810 ();
 sg13g2_decap_8 FILLER_0_817 ();
 sg13g2_decap_8 FILLER_0_824 ();
 sg13g2_decap_8 FILLER_0_831 ();
 sg13g2_decap_8 FILLER_0_838 ();
 sg13g2_decap_8 FILLER_0_845 ();
 sg13g2_decap_8 FILLER_0_852 ();
 sg13g2_decap_8 FILLER_0_859 ();
 sg13g2_decap_8 FILLER_0_866 ();
 sg13g2_decap_4 FILLER_0_873 ();
 sg13g2_fill_1 FILLER_0_877 ();
 sg13g2_decap_8 FILLER_1_0 ();
 sg13g2_decap_8 FILLER_1_7 ();
 sg13g2_decap_8 FILLER_1_14 ();
 sg13g2_decap_8 FILLER_1_21 ();
 sg13g2_decap_8 FILLER_1_28 ();
 sg13g2_decap_8 FILLER_1_35 ();
 sg13g2_decap_8 FILLER_1_42 ();
 sg13g2_decap_8 FILLER_1_49 ();
 sg13g2_decap_8 FILLER_1_56 ();
 sg13g2_decap_8 FILLER_1_63 ();
 sg13g2_decap_8 FILLER_1_70 ();
 sg13g2_decap_8 FILLER_1_77 ();
 sg13g2_decap_8 FILLER_1_84 ();
 sg13g2_decap_8 FILLER_1_91 ();
 sg13g2_decap_8 FILLER_1_98 ();
 sg13g2_decap_8 FILLER_1_105 ();
 sg13g2_decap_8 FILLER_1_112 ();
 sg13g2_decap_8 FILLER_1_119 ();
 sg13g2_fill_1 FILLER_1_126 ();
 sg13g2_decap_8 FILLER_1_131 ();
 sg13g2_decap_8 FILLER_1_138 ();
 sg13g2_decap_4 FILLER_1_145 ();
 sg13g2_fill_1 FILLER_1_149 ();
 sg13g2_fill_1 FILLER_1_161 ();
 sg13g2_fill_2 FILLER_1_170 ();
 sg13g2_decap_8 FILLER_1_180 ();
 sg13g2_fill_1 FILLER_1_187 ();
 sg13g2_fill_1 FILLER_1_197 ();
 sg13g2_decap_4 FILLER_1_202 ();
 sg13g2_fill_1 FILLER_1_206 ();
 sg13g2_fill_2 FILLER_1_212 ();
 sg13g2_fill_1 FILLER_1_214 ();
 sg13g2_fill_1 FILLER_1_220 ();
 sg13g2_fill_2 FILLER_1_225 ();
 sg13g2_decap_8 FILLER_1_232 ();
 sg13g2_fill_2 FILLER_1_239 ();
 sg13g2_fill_1 FILLER_1_241 ();
 sg13g2_fill_1 FILLER_1_246 ();
 sg13g2_fill_1 FILLER_1_252 ();
 sg13g2_fill_2 FILLER_1_258 ();
 sg13g2_fill_1 FILLER_1_260 ();
 sg13g2_decap_4 FILLER_1_266 ();
 sg13g2_fill_1 FILLER_1_286 ();
 sg13g2_fill_1 FILLER_1_291 ();
 sg13g2_fill_2 FILLER_1_296 ();
 sg13g2_fill_2 FILLER_1_306 ();
 sg13g2_fill_2 FILLER_1_343 ();
 sg13g2_decap_4 FILLER_1_352 ();
 sg13g2_decap_8 FILLER_1_361 ();
 sg13g2_decap_4 FILLER_1_368 ();
 sg13g2_fill_2 FILLER_1_372 ();
 sg13g2_fill_2 FILLER_1_378 ();
 sg13g2_decap_4 FILLER_1_428 ();
 sg13g2_fill_1 FILLER_1_432 ();
 sg13g2_decap_8 FILLER_1_459 ();
 sg13g2_decap_4 FILLER_1_466 ();
 sg13g2_fill_2 FILLER_1_470 ();
 sg13g2_decap_8 FILLER_1_476 ();
 sg13g2_decap_8 FILLER_1_483 ();
 sg13g2_decap_8 FILLER_1_490 ();
 sg13g2_decap_4 FILLER_1_497 ();
 sg13g2_decap_8 FILLER_1_509 ();
 sg13g2_decap_8 FILLER_1_521 ();
 sg13g2_decap_4 FILLER_1_528 ();
 sg13g2_decap_8 FILLER_1_540 ();
 sg13g2_decap_8 FILLER_1_547 ();
 sg13g2_decap_8 FILLER_1_554 ();
 sg13g2_decap_8 FILLER_1_561 ();
 sg13g2_fill_1 FILLER_1_572 ();
 sg13g2_fill_2 FILLER_1_586 ();
 sg13g2_fill_1 FILLER_1_588 ();
 sg13g2_fill_2 FILLER_1_610 ();
 sg13g2_fill_1 FILLER_1_612 ();
 sg13g2_decap_8 FILLER_1_623 ();
 sg13g2_fill_2 FILLER_1_630 ();
 sg13g2_decap_8 FILLER_1_647 ();
 sg13g2_fill_1 FILLER_1_654 ();
 sg13g2_decap_8 FILLER_1_659 ();
 sg13g2_fill_1 FILLER_1_666 ();
 sg13g2_decap_8 FILLER_1_694 ();
 sg13g2_fill_2 FILLER_1_701 ();
 sg13g2_fill_1 FILLER_1_703 ();
 sg13g2_fill_2 FILLER_1_716 ();
 sg13g2_fill_1 FILLER_1_718 ();
 sg13g2_decap_8 FILLER_1_724 ();
 sg13g2_fill_2 FILLER_1_731 ();
 sg13g2_fill_1 FILLER_1_733 ();
 sg13g2_decap_8 FILLER_1_747 ();
 sg13g2_decap_8 FILLER_1_763 ();
 sg13g2_decap_8 FILLER_1_770 ();
 sg13g2_decap_8 FILLER_1_777 ();
 sg13g2_decap_8 FILLER_1_784 ();
 sg13g2_decap_8 FILLER_1_791 ();
 sg13g2_decap_8 FILLER_1_798 ();
 sg13g2_decap_8 FILLER_1_805 ();
 sg13g2_decap_8 FILLER_1_812 ();
 sg13g2_decap_8 FILLER_1_819 ();
 sg13g2_decap_8 FILLER_1_826 ();
 sg13g2_decap_8 FILLER_1_833 ();
 sg13g2_decap_8 FILLER_1_840 ();
 sg13g2_decap_8 FILLER_1_847 ();
 sg13g2_decap_8 FILLER_1_854 ();
 sg13g2_decap_8 FILLER_1_861 ();
 sg13g2_decap_8 FILLER_1_868 ();
 sg13g2_fill_2 FILLER_1_875 ();
 sg13g2_fill_1 FILLER_1_877 ();
 sg13g2_decap_8 FILLER_2_0 ();
 sg13g2_decap_8 FILLER_2_7 ();
 sg13g2_decap_8 FILLER_2_14 ();
 sg13g2_decap_8 FILLER_2_21 ();
 sg13g2_decap_8 FILLER_2_28 ();
 sg13g2_decap_8 FILLER_2_35 ();
 sg13g2_decap_8 FILLER_2_42 ();
 sg13g2_decap_8 FILLER_2_49 ();
 sg13g2_decap_8 FILLER_2_56 ();
 sg13g2_decap_8 FILLER_2_63 ();
 sg13g2_decap_8 FILLER_2_70 ();
 sg13g2_decap_8 FILLER_2_77 ();
 sg13g2_decap_8 FILLER_2_84 ();
 sg13g2_decap_8 FILLER_2_91 ();
 sg13g2_decap_8 FILLER_2_98 ();
 sg13g2_decap_4 FILLER_2_105 ();
 sg13g2_fill_2 FILLER_2_135 ();
 sg13g2_fill_1 FILLER_2_137 ();
 sg13g2_decap_4 FILLER_2_142 ();
 sg13g2_decap_8 FILLER_2_171 ();
 sg13g2_decap_8 FILLER_2_178 ();
 sg13g2_decap_8 FILLER_2_185 ();
 sg13g2_decap_4 FILLER_2_192 ();
 sg13g2_decap_4 FILLER_2_229 ();
 sg13g2_decap_8 FILLER_2_250 ();
 sg13g2_decap_8 FILLER_2_257 ();
 sg13g2_decap_8 FILLER_2_264 ();
 sg13g2_fill_1 FILLER_2_271 ();
 sg13g2_decap_8 FILLER_2_277 ();
 sg13g2_decap_8 FILLER_2_288 ();
 sg13g2_decap_4 FILLER_2_295 ();
 sg13g2_fill_1 FILLER_2_299 ();
 sg13g2_decap_8 FILLER_2_310 ();
 sg13g2_decap_8 FILLER_2_322 ();
 sg13g2_decap_4 FILLER_2_329 ();
 sg13g2_fill_2 FILLER_2_333 ();
 sg13g2_decap_8 FILLER_2_340 ();
 sg13g2_decap_4 FILLER_2_347 ();
 sg13g2_fill_2 FILLER_2_351 ();
 sg13g2_fill_1 FILLER_2_359 ();
 sg13g2_decap_8 FILLER_2_364 ();
 sg13g2_decap_8 FILLER_2_371 ();
 sg13g2_fill_1 FILLER_2_378 ();
 sg13g2_fill_1 FILLER_2_396 ();
 sg13g2_decap_8 FILLER_2_406 ();
 sg13g2_decap_8 FILLER_2_413 ();
 sg13g2_decap_8 FILLER_2_420 ();
 sg13g2_decap_8 FILLER_2_427 ();
 sg13g2_decap_8 FILLER_2_438 ();
 sg13g2_decap_8 FILLER_2_445 ();
 sg13g2_decap_4 FILLER_2_452 ();
 sg13g2_fill_1 FILLER_2_456 ();
 sg13g2_decap_8 FILLER_2_473 ();
 sg13g2_decap_8 FILLER_2_480 ();
 sg13g2_decap_8 FILLER_2_487 ();
 sg13g2_decap_8 FILLER_2_494 ();
 sg13g2_decap_8 FILLER_2_501 ();
 sg13g2_decap_4 FILLER_2_508 ();
 sg13g2_decap_8 FILLER_2_535 ();
 sg13g2_decap_8 FILLER_2_542 ();
 sg13g2_decap_4 FILLER_2_549 ();
 sg13g2_fill_1 FILLER_2_558 ();
 sg13g2_decap_8 FILLER_2_569 ();
 sg13g2_fill_1 FILLER_2_576 ();
 sg13g2_decap_4 FILLER_2_621 ();
 sg13g2_fill_2 FILLER_2_638 ();
 sg13g2_fill_1 FILLER_2_640 ();
 sg13g2_decap_4 FILLER_2_645 ();
 sg13g2_decap_8 FILLER_2_659 ();
 sg13g2_fill_1 FILLER_2_666 ();
 sg13g2_decap_8 FILLER_2_671 ();
 sg13g2_decap_8 FILLER_2_678 ();
 sg13g2_fill_2 FILLER_2_685 ();
 sg13g2_fill_1 FILLER_2_702 ();
 sg13g2_decap_8 FILLER_2_708 ();
 sg13g2_fill_1 FILLER_2_715 ();
 sg13g2_fill_2 FILLER_2_721 ();
 sg13g2_decap_8 FILLER_2_743 ();
 sg13g2_decap_4 FILLER_2_750 ();
 sg13g2_decap_8 FILLER_2_767 ();
 sg13g2_decap_8 FILLER_2_774 ();
 sg13g2_decap_8 FILLER_2_781 ();
 sg13g2_decap_8 FILLER_2_788 ();
 sg13g2_decap_8 FILLER_2_795 ();
 sg13g2_decap_8 FILLER_2_802 ();
 sg13g2_decap_8 FILLER_2_809 ();
 sg13g2_decap_8 FILLER_2_816 ();
 sg13g2_decap_8 FILLER_2_823 ();
 sg13g2_decap_8 FILLER_2_830 ();
 sg13g2_decap_8 FILLER_2_837 ();
 sg13g2_decap_8 FILLER_2_844 ();
 sg13g2_decap_8 FILLER_2_851 ();
 sg13g2_decap_8 FILLER_2_858 ();
 sg13g2_decap_8 FILLER_2_865 ();
 sg13g2_decap_4 FILLER_2_872 ();
 sg13g2_fill_2 FILLER_2_876 ();
 sg13g2_decap_8 FILLER_3_0 ();
 sg13g2_decap_8 FILLER_3_7 ();
 sg13g2_decap_8 FILLER_3_14 ();
 sg13g2_decap_8 FILLER_3_21 ();
 sg13g2_decap_8 FILLER_3_28 ();
 sg13g2_decap_8 FILLER_3_35 ();
 sg13g2_decap_8 FILLER_3_42 ();
 sg13g2_decap_8 FILLER_3_49 ();
 sg13g2_decap_8 FILLER_3_56 ();
 sg13g2_decap_8 FILLER_3_63 ();
 sg13g2_decap_8 FILLER_3_70 ();
 sg13g2_decap_8 FILLER_3_77 ();
 sg13g2_decap_8 FILLER_3_84 ();
 sg13g2_decap_8 FILLER_3_91 ();
 sg13g2_decap_8 FILLER_3_98 ();
 sg13g2_decap_8 FILLER_3_105 ();
 sg13g2_fill_2 FILLER_3_112 ();
 sg13g2_fill_1 FILLER_3_114 ();
 sg13g2_decap_8 FILLER_3_119 ();
 sg13g2_decap_8 FILLER_3_126 ();
 sg13g2_decap_8 FILLER_3_133 ();
 sg13g2_decap_8 FILLER_3_140 ();
 sg13g2_fill_2 FILLER_3_147 ();
 sg13g2_fill_1 FILLER_3_149 ();
 sg13g2_fill_2 FILLER_3_158 ();
 sg13g2_decap_8 FILLER_3_197 ();
 sg13g2_decap_8 FILLER_3_204 ();
 sg13g2_decap_8 FILLER_3_211 ();
 sg13g2_decap_4 FILLER_3_218 ();
 sg13g2_decap_8 FILLER_3_226 ();
 sg13g2_fill_1 FILLER_3_233 ();
 sg13g2_decap_8 FILLER_3_238 ();
 sg13g2_decap_8 FILLER_3_245 ();
 sg13g2_decap_4 FILLER_3_252 ();
 sg13g2_decap_8 FILLER_3_264 ();
 sg13g2_decap_8 FILLER_3_271 ();
 sg13g2_decap_8 FILLER_3_278 ();
 sg13g2_fill_1 FILLER_3_285 ();
 sg13g2_decap_8 FILLER_3_294 ();
 sg13g2_decap_8 FILLER_3_301 ();
 sg13g2_decap_4 FILLER_3_308 ();
 sg13g2_fill_1 FILLER_3_312 ();
 sg13g2_decap_8 FILLER_3_339 ();
 sg13g2_decap_4 FILLER_3_346 ();
 sg13g2_fill_1 FILLER_3_350 ();
 sg13g2_decap_8 FILLER_3_364 ();
 sg13g2_decap_8 FILLER_3_371 ();
 sg13g2_decap_8 FILLER_3_378 ();
 sg13g2_decap_8 FILLER_3_385 ();
 sg13g2_fill_1 FILLER_3_392 ();
 sg13g2_decap_4 FILLER_3_397 ();
 sg13g2_fill_1 FILLER_3_401 ();
 sg13g2_decap_8 FILLER_3_407 ();
 sg13g2_decap_8 FILLER_3_414 ();
 sg13g2_decap_4 FILLER_3_431 ();
 sg13g2_fill_1 FILLER_3_435 ();
 sg13g2_decap_8 FILLER_3_444 ();
 sg13g2_decap_8 FILLER_3_451 ();
 sg13g2_decap_4 FILLER_3_458 ();
 sg13g2_fill_2 FILLER_3_471 ();
 sg13g2_decap_4 FILLER_3_477 ();
 sg13g2_decap_4 FILLER_3_492 ();
 sg13g2_fill_1 FILLER_3_496 ();
 sg13g2_decap_4 FILLER_3_507 ();
 sg13g2_fill_1 FILLER_3_511 ();
 sg13g2_fill_2 FILLER_3_557 ();
 sg13g2_decap_4 FILLER_3_563 ();
 sg13g2_fill_1 FILLER_3_567 ();
 sg13g2_fill_2 FILLER_3_591 ();
 sg13g2_fill_1 FILLER_3_593 ();
 sg13g2_fill_2 FILLER_3_598 ();
 sg13g2_fill_1 FILLER_3_600 ();
 sg13g2_decap_8 FILLER_3_605 ();
 sg13g2_decap_8 FILLER_3_612 ();
 sg13g2_decap_8 FILLER_3_634 ();
 sg13g2_fill_2 FILLER_3_641 ();
 sg13g2_decap_4 FILLER_3_647 ();
 sg13g2_fill_1 FILLER_3_651 ();
 sg13g2_decap_8 FILLER_3_656 ();
 sg13g2_fill_2 FILLER_3_663 ();
 sg13g2_fill_2 FILLER_3_674 ();
 sg13g2_fill_2 FILLER_3_708 ();
 sg13g2_decap_4 FILLER_3_725 ();
 sg13g2_fill_2 FILLER_3_729 ();
 sg13g2_fill_1 FILLER_3_753 ();
 sg13g2_decap_4 FILLER_3_772 ();
 sg13g2_fill_2 FILLER_3_780 ();
 sg13g2_fill_1 FILLER_3_787 ();
 sg13g2_decap_8 FILLER_3_792 ();
 sg13g2_decap_8 FILLER_3_803 ();
 sg13g2_decap_4 FILLER_3_810 ();
 sg13g2_decap_8 FILLER_3_818 ();
 sg13g2_fill_1 FILLER_3_825 ();
 sg13g2_decap_8 FILLER_3_830 ();
 sg13g2_decap_8 FILLER_3_837 ();
 sg13g2_decap_8 FILLER_3_844 ();
 sg13g2_decap_8 FILLER_3_851 ();
 sg13g2_decap_8 FILLER_3_858 ();
 sg13g2_decap_8 FILLER_3_865 ();
 sg13g2_decap_4 FILLER_3_872 ();
 sg13g2_fill_2 FILLER_3_876 ();
 sg13g2_decap_8 FILLER_4_0 ();
 sg13g2_decap_8 FILLER_4_7 ();
 sg13g2_decap_8 FILLER_4_14 ();
 sg13g2_decap_8 FILLER_4_21 ();
 sg13g2_decap_8 FILLER_4_28 ();
 sg13g2_fill_2 FILLER_4_35 ();
 sg13g2_fill_1 FILLER_4_37 ();
 sg13g2_decap_8 FILLER_4_42 ();
 sg13g2_decap_8 FILLER_4_49 ();
 sg13g2_decap_8 FILLER_4_56 ();
 sg13g2_decap_4 FILLER_4_63 ();
 sg13g2_decap_4 FILLER_4_97 ();
 sg13g2_fill_2 FILLER_4_101 ();
 sg13g2_decap_8 FILLER_4_107 ();
 sg13g2_fill_2 FILLER_4_114 ();
 sg13g2_fill_1 FILLER_4_116 ();
 sg13g2_decap_4 FILLER_4_173 ();
 sg13g2_fill_2 FILLER_4_177 ();
 sg13g2_fill_1 FILLER_4_192 ();
 sg13g2_decap_8 FILLER_4_229 ();
 sg13g2_fill_1 FILLER_4_236 ();
 sg13g2_fill_2 FILLER_4_247 ();
 sg13g2_decap_4 FILLER_4_280 ();
 sg13g2_fill_1 FILLER_4_284 ();
 sg13g2_decap_8 FILLER_4_325 ();
 sg13g2_fill_1 FILLER_4_350 ();
 sg13g2_decap_4 FILLER_4_384 ();
 sg13g2_fill_2 FILLER_4_428 ();
 sg13g2_decap_8 FILLER_4_445 ();
 sg13g2_decap_8 FILLER_4_452 ();
 sg13g2_decap_4 FILLER_4_459 ();
 sg13g2_fill_2 FILLER_4_475 ();
 sg13g2_decap_8 FILLER_4_485 ();
 sg13g2_decap_8 FILLER_4_492 ();
 sg13g2_fill_2 FILLER_4_499 ();
 sg13g2_decap_8 FILLER_4_517 ();
 sg13g2_decap_8 FILLER_4_524 ();
 sg13g2_decap_8 FILLER_4_531 ();
 sg13g2_decap_8 FILLER_4_538 ();
 sg13g2_decap_4 FILLER_4_545 ();
 sg13g2_decap_8 FILLER_4_554 ();
 sg13g2_fill_2 FILLER_4_561 ();
 sg13g2_fill_1 FILLER_4_563 ();
 sg13g2_fill_1 FILLER_4_579 ();
 sg13g2_decap_4 FILLER_4_584 ();
 sg13g2_fill_2 FILLER_4_588 ();
 sg13g2_fill_1 FILLER_4_604 ();
 sg13g2_fill_1 FILLER_4_615 ();
 sg13g2_fill_2 FILLER_4_625 ();
 sg13g2_decap_4 FILLER_4_631 ();
 sg13g2_fill_1 FILLER_4_635 ();
 sg13g2_fill_2 FILLER_4_640 ();
 sg13g2_fill_1 FILLER_4_642 ();
 sg13g2_decap_4 FILLER_4_661 ();
 sg13g2_fill_1 FILLER_4_665 ();
 sg13g2_fill_1 FILLER_4_671 ();
 sg13g2_fill_1 FILLER_4_682 ();
 sg13g2_fill_2 FILLER_4_710 ();
 sg13g2_fill_1 FILLER_4_712 ();
 sg13g2_decap_8 FILLER_4_719 ();
 sg13g2_decap_4 FILLER_4_730 ();
 sg13g2_fill_1 FILLER_4_739 ();
 sg13g2_fill_2 FILLER_4_781 ();
 sg13g2_fill_1 FILLER_4_783 ();
 sg13g2_fill_2 FILLER_4_788 ();
 sg13g2_fill_1 FILLER_4_790 ();
 sg13g2_fill_2 FILLER_4_795 ();
 sg13g2_fill_2 FILLER_4_801 ();
 sg13g2_fill_1 FILLER_4_803 ();
 sg13g2_fill_2 FILLER_4_809 ();
 sg13g2_fill_1 FILLER_4_811 ();
 sg13g2_fill_2 FILLER_4_817 ();
 sg13g2_fill_1 FILLER_4_819 ();
 sg13g2_decap_8 FILLER_4_824 ();
 sg13g2_decap_8 FILLER_4_831 ();
 sg13g2_decap_8 FILLER_4_838 ();
 sg13g2_decap_8 FILLER_4_845 ();
 sg13g2_decap_8 FILLER_4_852 ();
 sg13g2_decap_8 FILLER_4_859 ();
 sg13g2_decap_8 FILLER_4_866 ();
 sg13g2_decap_4 FILLER_4_873 ();
 sg13g2_fill_1 FILLER_4_877 ();
 sg13g2_decap_8 FILLER_5_0 ();
 sg13g2_decap_8 FILLER_5_7 ();
 sg13g2_decap_8 FILLER_5_14 ();
 sg13g2_decap_8 FILLER_5_21 ();
 sg13g2_fill_2 FILLER_5_28 ();
 sg13g2_fill_1 FILLER_5_30 ();
 sg13g2_decap_8 FILLER_5_61 ();
 sg13g2_fill_1 FILLER_5_68 ();
 sg13g2_fill_1 FILLER_5_73 ();
 sg13g2_decap_8 FILLER_5_82 ();
 sg13g2_fill_2 FILLER_5_89 ();
 sg13g2_fill_1 FILLER_5_91 ();
 sg13g2_decap_8 FILLER_5_132 ();
 sg13g2_decap_8 FILLER_5_139 ();
 sg13g2_decap_8 FILLER_5_146 ();
 sg13g2_decap_8 FILLER_5_153 ();
 sg13g2_decap_8 FILLER_5_160 ();
 sg13g2_decap_8 FILLER_5_167 ();
 sg13g2_decap_8 FILLER_5_174 ();
 sg13g2_fill_1 FILLER_5_181 ();
 sg13g2_decap_4 FILLER_5_208 ();
 sg13g2_decap_8 FILLER_5_216 ();
 sg13g2_decap_8 FILLER_5_223 ();
 sg13g2_decap_4 FILLER_5_230 ();
 sg13g2_fill_1 FILLER_5_234 ();
 sg13g2_decap_8 FILLER_5_265 ();
 sg13g2_decap_4 FILLER_5_272 ();
 sg13g2_fill_1 FILLER_5_276 ();
 sg13g2_decap_8 FILLER_5_281 ();
 sg13g2_decap_4 FILLER_5_288 ();
 sg13g2_fill_2 FILLER_5_292 ();
 sg13g2_decap_4 FILLER_5_301 ();
 sg13g2_fill_1 FILLER_5_305 ();
 sg13g2_decap_8 FILLER_5_310 ();
 sg13g2_decap_8 FILLER_5_317 ();
 sg13g2_decap_8 FILLER_5_324 ();
 sg13g2_decap_8 FILLER_5_331 ();
 sg13g2_decap_8 FILLER_5_338 ();
 sg13g2_decap_8 FILLER_5_345 ();
 sg13g2_decap_8 FILLER_5_352 ();
 sg13g2_fill_1 FILLER_5_359 ();
 sg13g2_decap_8 FILLER_5_374 ();
 sg13g2_decap_4 FILLER_5_391 ();
 sg13g2_fill_2 FILLER_5_395 ();
 sg13g2_fill_1 FILLER_5_402 ();
 sg13g2_decap_4 FILLER_5_418 ();
 sg13g2_fill_1 FILLER_5_422 ();
 sg13g2_decap_8 FILLER_5_439 ();
 sg13g2_decap_4 FILLER_5_446 ();
 sg13g2_decap_8 FILLER_5_467 ();
 sg13g2_fill_2 FILLER_5_474 ();
 sg13g2_fill_1 FILLER_5_476 ();
 sg13g2_decap_8 FILLER_5_481 ();
 sg13g2_decap_8 FILLER_5_488 ();
 sg13g2_decap_8 FILLER_5_495 ();
 sg13g2_fill_1 FILLER_5_502 ();
 sg13g2_decap_4 FILLER_5_518 ();
 sg13g2_decap_8 FILLER_5_526 ();
 sg13g2_decap_4 FILLER_5_533 ();
 sg13g2_fill_2 FILLER_5_537 ();
 sg13g2_fill_2 FILLER_5_549 ();
 sg13g2_fill_1 FILLER_5_595 ();
 sg13g2_fill_2 FILLER_5_602 ();
 sg13g2_fill_2 FILLER_5_614 ();
 sg13g2_fill_2 FILLER_5_624 ();
 sg13g2_fill_1 FILLER_5_640 ();
 sg13g2_decap_8 FILLER_5_685 ();
 sg13g2_fill_1 FILLER_5_700 ();
 sg13g2_fill_2 FILLER_5_714 ();
 sg13g2_fill_1 FILLER_5_716 ();
 sg13g2_decap_4 FILLER_5_722 ();
 sg13g2_fill_2 FILLER_5_726 ();
 sg13g2_fill_1 FILLER_5_761 ();
 sg13g2_decap_8 FILLER_5_768 ();
 sg13g2_decap_4 FILLER_5_775 ();
 sg13g2_fill_1 FILLER_5_779 ();
 sg13g2_fill_1 FILLER_5_793 ();
 sg13g2_fill_1 FILLER_5_804 ();
 sg13g2_fill_1 FILLER_5_814 ();
 sg13g2_decap_8 FILLER_5_824 ();
 sg13g2_decap_8 FILLER_5_831 ();
 sg13g2_decap_8 FILLER_5_838 ();
 sg13g2_decap_8 FILLER_5_845 ();
 sg13g2_decap_8 FILLER_5_852 ();
 sg13g2_decap_8 FILLER_5_859 ();
 sg13g2_decap_8 FILLER_5_866 ();
 sg13g2_decap_4 FILLER_5_873 ();
 sg13g2_fill_1 FILLER_5_877 ();
 sg13g2_decap_8 FILLER_6_0 ();
 sg13g2_decap_8 FILLER_6_7 ();
 sg13g2_decap_4 FILLER_6_14 ();
 sg13g2_fill_2 FILLER_6_18 ();
 sg13g2_decap_8 FILLER_6_24 ();
 sg13g2_fill_2 FILLER_6_31 ();
 sg13g2_fill_2 FILLER_6_49 ();
 sg13g2_fill_1 FILLER_6_59 ();
 sg13g2_fill_2 FILLER_6_88 ();
 sg13g2_fill_1 FILLER_6_90 ();
 sg13g2_decap_8 FILLER_6_101 ();
 sg13g2_decap_8 FILLER_6_108 ();
 sg13g2_fill_2 FILLER_6_115 ();
 sg13g2_fill_1 FILLER_6_117 ();
 sg13g2_decap_8 FILLER_6_127 ();
 sg13g2_decap_8 FILLER_6_134 ();
 sg13g2_fill_2 FILLER_6_141 ();
 sg13g2_decap_8 FILLER_6_169 ();
 sg13g2_fill_2 FILLER_6_176 ();
 sg13g2_fill_1 FILLER_6_178 ();
 sg13g2_decap_8 FILLER_6_189 ();
 sg13g2_fill_1 FILLER_6_196 ();
 sg13g2_decap_8 FILLER_6_206 ();
 sg13g2_fill_1 FILLER_6_213 ();
 sg13g2_decap_8 FILLER_6_218 ();
 sg13g2_decap_8 FILLER_6_225 ();
 sg13g2_decap_8 FILLER_6_232 ();
 sg13g2_decap_8 FILLER_6_239 ();
 sg13g2_fill_2 FILLER_6_246 ();
 sg13g2_decap_4 FILLER_6_264 ();
 sg13g2_fill_2 FILLER_6_268 ();
 sg13g2_decap_4 FILLER_6_290 ();
 sg13g2_fill_1 FILLER_6_294 ();
 sg13g2_decap_8 FILLER_6_320 ();
 sg13g2_decap_4 FILLER_6_327 ();
 sg13g2_fill_1 FILLER_6_331 ();
 sg13g2_fill_2 FILLER_6_344 ();
 sg13g2_decap_4 FILLER_6_356 ();
 sg13g2_fill_2 FILLER_6_360 ();
 sg13g2_decap_8 FILLER_6_376 ();
 sg13g2_decap_8 FILLER_6_383 ();
 sg13g2_decap_8 FILLER_6_390 ();
 sg13g2_decap_4 FILLER_6_397 ();
 sg13g2_decap_8 FILLER_6_406 ();
 sg13g2_decap_4 FILLER_6_413 ();
 sg13g2_fill_2 FILLER_6_417 ();
 sg13g2_fill_1 FILLER_6_432 ();
 sg13g2_decap_8 FILLER_6_438 ();
 sg13g2_decap_8 FILLER_6_445 ();
 sg13g2_decap_4 FILLER_6_452 ();
 sg13g2_decap_4 FILLER_6_471 ();
 sg13g2_fill_2 FILLER_6_479 ();
 sg13g2_fill_2 FILLER_6_492 ();
 sg13g2_fill_1 FILLER_6_494 ();
 sg13g2_decap_8 FILLER_6_500 ();
 sg13g2_decap_8 FILLER_6_517 ();
 sg13g2_decap_8 FILLER_6_524 ();
 sg13g2_decap_8 FILLER_6_531 ();
 sg13g2_fill_1 FILLER_6_538 ();
 sg13g2_fill_2 FILLER_6_543 ();
 sg13g2_fill_2 FILLER_6_564 ();
 sg13g2_fill_1 FILLER_6_581 ();
 sg13g2_fill_2 FILLER_6_603 ();
 sg13g2_fill_2 FILLER_6_613 ();
 sg13g2_decap_8 FILLER_6_620 ();
 sg13g2_decap_8 FILLER_6_627 ();
 sg13g2_decap_4 FILLER_6_634 ();
 sg13g2_fill_1 FILLER_6_638 ();
 sg13g2_decap_8 FILLER_6_655 ();
 sg13g2_decap_8 FILLER_6_662 ();
 sg13g2_decap_4 FILLER_6_669 ();
 sg13g2_fill_2 FILLER_6_677 ();
 sg13g2_fill_1 FILLER_6_690 ();
 sg13g2_fill_1 FILLER_6_701 ();
 sg13g2_fill_1 FILLER_6_708 ();
 sg13g2_decap_8 FILLER_6_713 ();
 sg13g2_decap_8 FILLER_6_720 ();
 sg13g2_decap_8 FILLER_6_727 ();
 sg13g2_decap_8 FILLER_6_734 ();
 sg13g2_fill_1 FILLER_6_746 ();
 sg13g2_fill_1 FILLER_6_758 ();
 sg13g2_decap_4 FILLER_6_774 ();
 sg13g2_fill_2 FILLER_6_778 ();
 sg13g2_fill_2 FILLER_6_789 ();
 sg13g2_fill_2 FILLER_6_802 ();
 sg13g2_fill_1 FILLER_6_804 ();
 sg13g2_fill_2 FILLER_6_813 ();
 sg13g2_fill_1 FILLER_6_815 ();
 sg13g2_fill_1 FILLER_6_825 ();
 sg13g2_decap_8 FILLER_6_834 ();
 sg13g2_decap_8 FILLER_6_841 ();
 sg13g2_decap_8 FILLER_6_848 ();
 sg13g2_decap_8 FILLER_6_855 ();
 sg13g2_decap_8 FILLER_6_862 ();
 sg13g2_decap_8 FILLER_6_869 ();
 sg13g2_fill_2 FILLER_6_876 ();
 sg13g2_fill_1 FILLER_7_26 ();
 sg13g2_decap_8 FILLER_7_31 ();
 sg13g2_fill_2 FILLER_7_38 ();
 sg13g2_fill_1 FILLER_7_40 ();
 sg13g2_fill_2 FILLER_7_49 ();
 sg13g2_fill_2 FILLER_7_65 ();
 sg13g2_fill_1 FILLER_7_67 ();
 sg13g2_fill_2 FILLER_7_81 ();
 sg13g2_fill_1 FILLER_7_87 ();
 sg13g2_decap_4 FILLER_7_91 ();
 sg13g2_fill_2 FILLER_7_95 ();
 sg13g2_fill_2 FILLER_7_105 ();
 sg13g2_fill_1 FILLER_7_110 ();
 sg13g2_fill_2 FILLER_7_137 ();
 sg13g2_decap_8 FILLER_7_153 ();
 sg13g2_decap_8 FILLER_7_160 ();
 sg13g2_decap_8 FILLER_7_167 ();
 sg13g2_decap_4 FILLER_7_188 ();
 sg13g2_fill_1 FILLER_7_192 ();
 sg13g2_fill_2 FILLER_7_197 ();
 sg13g2_fill_1 FILLER_7_234 ();
 sg13g2_decap_8 FILLER_7_259 ();
 sg13g2_decap_8 FILLER_7_315 ();
 sg13g2_fill_1 FILLER_7_322 ();
 sg13g2_decap_4 FILLER_7_338 ();
 sg13g2_fill_1 FILLER_7_342 ();
 sg13g2_fill_1 FILLER_7_365 ();
 sg13g2_decap_8 FILLER_7_372 ();
 sg13g2_decap_8 FILLER_7_379 ();
 sg13g2_decap_8 FILLER_7_386 ();
 sg13g2_decap_8 FILLER_7_393 ();
 sg13g2_fill_2 FILLER_7_400 ();
 sg13g2_decap_8 FILLER_7_412 ();
 sg13g2_decap_4 FILLER_7_419 ();
 sg13g2_decap_8 FILLER_7_431 ();
 sg13g2_fill_2 FILLER_7_438 ();
 sg13g2_fill_1 FILLER_7_440 ();
 sg13g2_fill_1 FILLER_7_446 ();
 sg13g2_fill_2 FILLER_7_451 ();
 sg13g2_fill_1 FILLER_7_461 ();
 sg13g2_fill_2 FILLER_7_470 ();
 sg13g2_fill_1 FILLER_7_472 ();
 sg13g2_fill_1 FILLER_7_483 ();
 sg13g2_fill_1 FILLER_7_489 ();
 sg13g2_decap_4 FILLER_7_508 ();
 sg13g2_fill_2 FILLER_7_512 ();
 sg13g2_decap_8 FILLER_7_525 ();
 sg13g2_decap_8 FILLER_7_532 ();
 sg13g2_fill_1 FILLER_7_539 ();
 sg13g2_fill_1 FILLER_7_552 ();
 sg13g2_fill_2 FILLER_7_557 ();
 sg13g2_fill_1 FILLER_7_564 ();
 sg13g2_fill_2 FILLER_7_570 ();
 sg13g2_decap_4 FILLER_7_593 ();
 sg13g2_fill_1 FILLER_7_597 ();
 sg13g2_decap_4 FILLER_7_602 ();
 sg13g2_fill_2 FILLER_7_612 ();
 sg13g2_decap_8 FILLER_7_620 ();
 sg13g2_decap_4 FILLER_7_627 ();
 sg13g2_fill_2 FILLER_7_636 ();
 sg13g2_fill_2 FILLER_7_655 ();
 sg13g2_fill_1 FILLER_7_676 ();
 sg13g2_fill_1 FILLER_7_682 ();
 sg13g2_fill_1 FILLER_7_688 ();
 sg13g2_fill_1 FILLER_7_699 ();
 sg13g2_decap_8 FILLER_7_704 ();
 sg13g2_decap_8 FILLER_7_711 ();
 sg13g2_fill_1 FILLER_7_718 ();
 sg13g2_fill_2 FILLER_7_729 ();
 sg13g2_fill_1 FILLER_7_741 ();
 sg13g2_fill_1 FILLER_7_747 ();
 sg13g2_fill_1 FILLER_7_759 ();
 sg13g2_decap_4 FILLER_7_775 ();
 sg13g2_decap_4 FILLER_7_792 ();
 sg13g2_fill_2 FILLER_7_796 ();
 sg13g2_fill_2 FILLER_7_817 ();
 sg13g2_decap_4 FILLER_7_826 ();
 sg13g2_decap_8 FILLER_7_835 ();
 sg13g2_decap_8 FILLER_7_842 ();
 sg13g2_decap_8 FILLER_7_849 ();
 sg13g2_decap_8 FILLER_7_856 ();
 sg13g2_decap_8 FILLER_7_863 ();
 sg13g2_decap_8 FILLER_7_870 ();
 sg13g2_fill_1 FILLER_7_877 ();
 sg13g2_decap_4 FILLER_8_0 ();
 sg13g2_decap_8 FILLER_8_8 ();
 sg13g2_decap_8 FILLER_8_15 ();
 sg13g2_decap_8 FILLER_8_22 ();
 sg13g2_decap_8 FILLER_8_29 ();
 sg13g2_decap_8 FILLER_8_36 ();
 sg13g2_decap_4 FILLER_8_43 ();
 sg13g2_fill_1 FILLER_8_47 ();
 sg13g2_decap_4 FILLER_8_62 ();
 sg13g2_decap_8 FILLER_8_84 ();
 sg13g2_decap_8 FILLER_8_91 ();
 sg13g2_fill_2 FILLER_8_98 ();
 sg13g2_fill_1 FILLER_8_100 ();
 sg13g2_decap_8 FILLER_8_109 ();
 sg13g2_decap_8 FILLER_8_116 ();
 sg13g2_decap_4 FILLER_8_123 ();
 sg13g2_fill_1 FILLER_8_127 ();
 sg13g2_fill_1 FILLER_8_132 ();
 sg13g2_decap_8 FILLER_8_141 ();
 sg13g2_decap_8 FILLER_8_148 ();
 sg13g2_decap_4 FILLER_8_155 ();
 sg13g2_fill_2 FILLER_8_159 ();
 sg13g2_decap_8 FILLER_8_199 ();
 sg13g2_decap_8 FILLER_8_206 ();
 sg13g2_decap_8 FILLER_8_213 ();
 sg13g2_decap_8 FILLER_8_220 ();
 sg13g2_fill_2 FILLER_8_227 ();
 sg13g2_decap_8 FILLER_8_239 ();
 sg13g2_fill_2 FILLER_8_246 ();
 sg13g2_fill_1 FILLER_8_248 ();
 sg13g2_decap_8 FILLER_8_261 ();
 sg13g2_decap_4 FILLER_8_268 ();
 sg13g2_fill_2 FILLER_8_284 ();
 sg13g2_fill_1 FILLER_8_286 ();
 sg13g2_fill_2 FILLER_8_292 ();
 sg13g2_decap_8 FILLER_8_302 ();
 sg13g2_decap_8 FILLER_8_309 ();
 sg13g2_decap_4 FILLER_8_316 ();
 sg13g2_fill_2 FILLER_8_320 ();
 sg13g2_fill_1 FILLER_8_342 ();
 sg13g2_fill_2 FILLER_8_353 ();
 sg13g2_decap_4 FILLER_8_365 ();
 sg13g2_fill_2 FILLER_8_377 ();
 sg13g2_decap_8 FILLER_8_393 ();
 sg13g2_fill_2 FILLER_8_400 ();
 sg13g2_decap_4 FILLER_8_423 ();
 sg13g2_decap_4 FILLER_8_431 ();
 sg13g2_decap_4 FILLER_8_445 ();
 sg13g2_fill_2 FILLER_8_449 ();
 sg13g2_fill_2 FILLER_8_459 ();
 sg13g2_decap_8 FILLER_8_469 ();
 sg13g2_fill_1 FILLER_8_476 ();
 sg13g2_fill_2 FILLER_8_480 ();
 sg13g2_fill_1 FILLER_8_482 ();
 sg13g2_decap_4 FILLER_8_488 ();
 sg13g2_fill_1 FILLER_8_492 ();
 sg13g2_fill_1 FILLER_8_498 ();
 sg13g2_fill_1 FILLER_8_515 ();
 sg13g2_decap_8 FILLER_8_540 ();
 sg13g2_decap_8 FILLER_8_547 ();
 sg13g2_decap_8 FILLER_8_554 ();
 sg13g2_decap_8 FILLER_8_561 ();
 sg13g2_decap_8 FILLER_8_568 ();
 sg13g2_decap_4 FILLER_8_579 ();
 sg13g2_fill_1 FILLER_8_583 ();
 sg13g2_decap_8 FILLER_8_595 ();
 sg13g2_decap_8 FILLER_8_602 ();
 sg13g2_decap_8 FILLER_8_609 ();
 sg13g2_decap_8 FILLER_8_616 ();
 sg13g2_decap_4 FILLER_8_623 ();
 sg13g2_fill_1 FILLER_8_627 ();
 sg13g2_decap_8 FILLER_8_642 ();
 sg13g2_decap_4 FILLER_8_649 ();
 sg13g2_decap_4 FILLER_8_659 ();
 sg13g2_fill_1 FILLER_8_663 ();
 sg13g2_fill_2 FILLER_8_679 ();
 sg13g2_fill_1 FILLER_8_681 ();
 sg13g2_fill_2 FILLER_8_712 ();
 sg13g2_fill_1 FILLER_8_719 ();
 sg13g2_decap_8 FILLER_8_728 ();
 sg13g2_decap_4 FILLER_8_735 ();
 sg13g2_fill_1 FILLER_8_739 ();
 sg13g2_decap_8 FILLER_8_749 ();
 sg13g2_fill_2 FILLER_8_756 ();
 sg13g2_fill_2 FILLER_8_791 ();
 sg13g2_fill_1 FILLER_8_793 ();
 sg13g2_fill_1 FILLER_8_825 ();
 sg13g2_decap_8 FILLER_8_831 ();
 sg13g2_decap_8 FILLER_8_838 ();
 sg13g2_decap_8 FILLER_8_845 ();
 sg13g2_decap_8 FILLER_8_852 ();
 sg13g2_decap_8 FILLER_8_859 ();
 sg13g2_decap_8 FILLER_8_866 ();
 sg13g2_decap_4 FILLER_8_873 ();
 sg13g2_fill_1 FILLER_8_877 ();
 sg13g2_fill_1 FILLER_9_0 ();
 sg13g2_fill_2 FILLER_9_27 ();
 sg13g2_decap_8 FILLER_9_33 ();
 sg13g2_decap_8 FILLER_9_40 ();
 sg13g2_fill_1 FILLER_9_58 ();
 sg13g2_fill_1 FILLER_9_64 ();
 sg13g2_decap_8 FILLER_9_83 ();
 sg13g2_decap_8 FILLER_9_90 ();
 sg13g2_fill_1 FILLER_9_97 ();
 sg13g2_decap_8 FILLER_9_103 ();
 sg13g2_fill_2 FILLER_9_110 ();
 sg13g2_decap_8 FILLER_9_116 ();
 sg13g2_fill_1 FILLER_9_123 ();
 sg13g2_fill_1 FILLER_9_154 ();
 sg13g2_decap_8 FILLER_9_160 ();
 sg13g2_fill_2 FILLER_9_167 ();
 sg13g2_fill_1 FILLER_9_169 ();
 sg13g2_decap_4 FILLER_9_180 ();
 sg13g2_decap_8 FILLER_9_192 ();
 sg13g2_decap_8 FILLER_9_199 ();
 sg13g2_fill_1 FILLER_9_206 ();
 sg13g2_fill_2 FILLER_9_211 ();
 sg13g2_fill_2 FILLER_9_239 ();
 sg13g2_fill_1 FILLER_9_241 ();
 sg13g2_decap_8 FILLER_9_247 ();
 sg13g2_decap_8 FILLER_9_254 ();
 sg13g2_fill_2 FILLER_9_261 ();
 sg13g2_decap_4 FILLER_9_268 ();
 sg13g2_fill_2 FILLER_9_276 ();
 sg13g2_decap_4 FILLER_9_286 ();
 sg13g2_decap_8 FILLER_9_302 ();
 sg13g2_decap_8 FILLER_9_309 ();
 sg13g2_fill_2 FILLER_9_316 ();
 sg13g2_fill_2 FILLER_9_323 ();
 sg13g2_fill_1 FILLER_9_337 ();
 sg13g2_fill_2 FILLER_9_350 ();
 sg13g2_decap_8 FILLER_9_360 ();
 sg13g2_decap_8 FILLER_9_367 ();
 sg13g2_fill_2 FILLER_9_374 ();
 sg13g2_fill_1 FILLER_9_376 ();
 sg13g2_fill_2 FILLER_9_395 ();
 sg13g2_fill_2 FILLER_9_409 ();
 sg13g2_fill_2 FILLER_9_424 ();
 sg13g2_decap_8 FILLER_9_453 ();
 sg13g2_decap_8 FILLER_9_460 ();
 sg13g2_fill_2 FILLER_9_467 ();
 sg13g2_fill_1 FILLER_9_469 ();
 sg13g2_fill_2 FILLER_9_474 ();
 sg13g2_fill_1 FILLER_9_476 ();
 sg13g2_decap_8 FILLER_9_486 ();
 sg13g2_decap_8 FILLER_9_493 ();
 sg13g2_fill_2 FILLER_9_500 ();
 sg13g2_decap_8 FILLER_9_507 ();
 sg13g2_decap_8 FILLER_9_518 ();
 sg13g2_decap_8 FILLER_9_525 ();
 sg13g2_fill_1 FILLER_9_532 ();
 sg13g2_decap_4 FILLER_9_543 ();
 sg13g2_fill_2 FILLER_9_547 ();
 sg13g2_decap_8 FILLER_9_554 ();
 sg13g2_decap_8 FILLER_9_561 ();
 sg13g2_decap_4 FILLER_9_568 ();
 sg13g2_decap_8 FILLER_9_582 ();
 sg13g2_fill_2 FILLER_9_589 ();
 sg13g2_fill_1 FILLER_9_591 ();
 sg13g2_fill_1 FILLER_9_597 ();
 sg13g2_fill_1 FILLER_9_602 ();
 sg13g2_fill_1 FILLER_9_612 ();
 sg13g2_fill_2 FILLER_9_618 ();
 sg13g2_fill_1 FILLER_9_620 ();
 sg13g2_decap_8 FILLER_9_626 ();
 sg13g2_decap_8 FILLER_9_638 ();
 sg13g2_decap_4 FILLER_9_645 ();
 sg13g2_fill_2 FILLER_9_654 ();
 sg13g2_fill_1 FILLER_9_656 ();
 sg13g2_fill_2 FILLER_9_670 ();
 sg13g2_decap_4 FILLER_9_685 ();
 sg13g2_fill_2 FILLER_9_689 ();
 sg13g2_fill_2 FILLER_9_695 ();
 sg13g2_decap_8 FILLER_9_706 ();
 sg13g2_decap_8 FILLER_9_713 ();
 sg13g2_decap_8 FILLER_9_720 ();
 sg13g2_fill_1 FILLER_9_727 ();
 sg13g2_fill_1 FILLER_9_748 ();
 sg13g2_fill_2 FILLER_9_754 ();
 sg13g2_fill_1 FILLER_9_756 ();
 sg13g2_fill_1 FILLER_9_767 ();
 sg13g2_decap_4 FILLER_9_778 ();
 sg13g2_fill_1 FILLER_9_786 ();
 sg13g2_fill_1 FILLER_9_795 ();
 sg13g2_decap_4 FILLER_9_809 ();
 sg13g2_fill_2 FILLER_9_813 ();
 sg13g2_decap_8 FILLER_9_840 ();
 sg13g2_decap_8 FILLER_9_847 ();
 sg13g2_decap_8 FILLER_9_854 ();
 sg13g2_decap_8 FILLER_9_861 ();
 sg13g2_decap_8 FILLER_9_868 ();
 sg13g2_fill_2 FILLER_9_875 ();
 sg13g2_fill_1 FILLER_9_877 ();
 sg13g2_decap_8 FILLER_10_0 ();
 sg13g2_decap_8 FILLER_10_11 ();
 sg13g2_decap_8 FILLER_10_18 ();
 sg13g2_decap_4 FILLER_10_25 ();
 sg13g2_fill_2 FILLER_10_62 ();
 sg13g2_fill_1 FILLER_10_64 ();
 sg13g2_decap_4 FILLER_10_81 ();
 sg13g2_decap_8 FILLER_10_89 ();
 sg13g2_fill_1 FILLER_10_96 ();
 sg13g2_decap_4 FILLER_10_100 ();
 sg13g2_fill_2 FILLER_10_104 ();
 sg13g2_fill_2 FILLER_10_132 ();
 sg13g2_decap_8 FILLER_10_139 ();
 sg13g2_decap_8 FILLER_10_156 ();
 sg13g2_decap_8 FILLER_10_163 ();
 sg13g2_decap_8 FILLER_10_178 ();
 sg13g2_decap_4 FILLER_10_185 ();
 sg13g2_fill_1 FILLER_10_189 ();
 sg13g2_decap_4 FILLER_10_198 ();
 sg13g2_fill_2 FILLER_10_202 ();
 sg13g2_fill_2 FILLER_10_208 ();
 sg13g2_fill_1 FILLER_10_210 ();
 sg13g2_fill_2 FILLER_10_220 ();
 sg13g2_fill_1 FILLER_10_222 ();
 sg13g2_decap_8 FILLER_10_238 ();
 sg13g2_decap_8 FILLER_10_245 ();
 sg13g2_decap_8 FILLER_10_252 ();
 sg13g2_fill_1 FILLER_10_259 ();
 sg13g2_decap_8 FILLER_10_274 ();
 sg13g2_decap_4 FILLER_10_281 ();
 sg13g2_fill_1 FILLER_10_285 ();
 sg13g2_decap_8 FILLER_10_300 ();
 sg13g2_decap_4 FILLER_10_307 ();
 sg13g2_decap_4 FILLER_10_325 ();
 sg13g2_fill_2 FILLER_10_329 ();
 sg13g2_decap_8 FILLER_10_341 ();
 sg13g2_decap_4 FILLER_10_348 ();
 sg13g2_fill_1 FILLER_10_352 ();
 sg13g2_decap_8 FILLER_10_357 ();
 sg13g2_decap_8 FILLER_10_364 ();
 sg13g2_decap_8 FILLER_10_371 ();
 sg13g2_decap_8 FILLER_10_382 ();
 sg13g2_decap_8 FILLER_10_389 ();
 sg13g2_decap_4 FILLER_10_396 ();
 sg13g2_fill_1 FILLER_10_400 ();
 sg13g2_fill_1 FILLER_10_414 ();
 sg13g2_decap_4 FILLER_10_420 ();
 sg13g2_decap_8 FILLER_10_429 ();
 sg13g2_fill_2 FILLER_10_436 ();
 sg13g2_decap_8 FILLER_10_447 ();
 sg13g2_decap_8 FILLER_10_454 ();
 sg13g2_decap_4 FILLER_10_461 ();
 sg13g2_fill_1 FILLER_10_465 ();
 sg13g2_fill_2 FILLER_10_471 ();
 sg13g2_decap_8 FILLER_10_494 ();
 sg13g2_fill_1 FILLER_10_501 ();
 sg13g2_decap_4 FILLER_10_510 ();
 sg13g2_fill_2 FILLER_10_518 ();
 sg13g2_fill_1 FILLER_10_530 ();
 sg13g2_fill_2 FILLER_10_549 ();
 sg13g2_fill_1 FILLER_10_551 ();
 sg13g2_fill_1 FILLER_10_563 ();
 sg13g2_fill_2 FILLER_10_589 ();
 sg13g2_fill_2 FILLER_10_617 ();
 sg13g2_fill_2 FILLER_10_631 ();
 sg13g2_decap_8 FILLER_10_650 ();
 sg13g2_fill_2 FILLER_10_657 ();
 sg13g2_decap_8 FILLER_10_663 ();
 sg13g2_decap_4 FILLER_10_670 ();
 sg13g2_fill_2 FILLER_10_674 ();
 sg13g2_fill_1 FILLER_10_681 ();
 sg13g2_decap_8 FILLER_10_687 ();
 sg13g2_decap_4 FILLER_10_694 ();
 sg13g2_decap_8 FILLER_10_708 ();
 sg13g2_fill_2 FILLER_10_715 ();
 sg13g2_decap_8 FILLER_10_722 ();
 sg13g2_decap_4 FILLER_10_729 ();
 sg13g2_fill_1 FILLER_10_733 ();
 sg13g2_fill_2 FILLER_10_752 ();
 sg13g2_fill_2 FILLER_10_774 ();
 sg13g2_fill_1 FILLER_10_776 ();
 sg13g2_fill_1 FILLER_10_788 ();
 sg13g2_decap_4 FILLER_10_798 ();
 sg13g2_fill_1 FILLER_10_802 ();
 sg13g2_decap_4 FILLER_10_823 ();
 sg13g2_fill_1 FILLER_10_827 ();
 sg13g2_decap_8 FILLER_10_833 ();
 sg13g2_decap_8 FILLER_10_840 ();
 sg13g2_decap_8 FILLER_10_847 ();
 sg13g2_decap_8 FILLER_10_854 ();
 sg13g2_decap_8 FILLER_10_861 ();
 sg13g2_decap_8 FILLER_10_868 ();
 sg13g2_fill_2 FILLER_10_875 ();
 sg13g2_fill_1 FILLER_10_877 ();
 sg13g2_decap_8 FILLER_11_0 ();
 sg13g2_decap_8 FILLER_11_7 ();
 sg13g2_decap_8 FILLER_11_14 ();
 sg13g2_decap_8 FILLER_11_21 ();
 sg13g2_fill_2 FILLER_11_28 ();
 sg13g2_fill_1 FILLER_11_42 ();
 sg13g2_decap_4 FILLER_11_67 ();
 sg13g2_decap_4 FILLER_11_75 ();
 sg13g2_decap_8 FILLER_11_105 ();
 sg13g2_fill_2 FILLER_11_112 ();
 sg13g2_fill_1 FILLER_11_114 ();
 sg13g2_decap_4 FILLER_11_169 ();
 sg13g2_fill_1 FILLER_11_173 ();
 sg13g2_decap_8 FILLER_11_183 ();
 sg13g2_decap_8 FILLER_11_190 ();
 sg13g2_decap_4 FILLER_11_197 ();
 sg13g2_fill_1 FILLER_11_201 ();
 sg13g2_fill_1 FILLER_11_223 ();
 sg13g2_fill_2 FILLER_11_232 ();
 sg13g2_fill_2 FILLER_11_238 ();
 sg13g2_fill_2 FILLER_11_245 ();
 sg13g2_fill_2 FILLER_11_273 ();
 sg13g2_fill_1 FILLER_11_275 ();
 sg13g2_fill_2 FILLER_11_302 ();
 sg13g2_fill_1 FILLER_11_304 ();
 sg13g2_decap_8 FILLER_11_331 ();
 sg13g2_decap_4 FILLER_11_364 ();
 sg13g2_decap_8 FILLER_11_411 ();
 sg13g2_decap_8 FILLER_11_418 ();
 sg13g2_decap_8 FILLER_11_425 ();
 sg13g2_decap_8 FILLER_11_432 ();
 sg13g2_decap_8 FILLER_11_439 ();
 sg13g2_decap_8 FILLER_11_446 ();
 sg13g2_decap_8 FILLER_11_453 ();
 sg13g2_decap_4 FILLER_11_460 ();
 sg13g2_fill_1 FILLER_11_464 ();
 sg13g2_fill_2 FILLER_11_475 ();
 sg13g2_fill_1 FILLER_11_477 ();
 sg13g2_fill_2 FILLER_11_491 ();
 sg13g2_fill_1 FILLER_11_493 ();
 sg13g2_fill_1 FILLER_11_500 ();
 sg13g2_fill_2 FILLER_11_506 ();
 sg13g2_decap_4 FILLER_11_528 ();
 sg13g2_fill_1 FILLER_11_536 ();
 sg13g2_decap_4 FILLER_11_544 ();
 sg13g2_fill_2 FILLER_11_548 ();
 sg13g2_decap_8 FILLER_11_559 ();
 sg13g2_fill_2 FILLER_11_584 ();
 sg13g2_fill_1 FILLER_11_586 ();
 sg13g2_fill_2 FILLER_11_593 ();
 sg13g2_fill_2 FILLER_11_605 ();
 sg13g2_fill_1 FILLER_11_615 ();
 sg13g2_fill_2 FILLER_11_621 ();
 sg13g2_fill_2 FILLER_11_631 ();
 sg13g2_decap_4 FILLER_11_641 ();
 sg13g2_fill_2 FILLER_11_653 ();
 sg13g2_fill_1 FILLER_11_665 ();
 sg13g2_decap_4 FILLER_11_675 ();
 sg13g2_fill_2 FILLER_11_702 ();
 sg13g2_fill_1 FILLER_11_709 ();
 sg13g2_decap_8 FILLER_11_715 ();
 sg13g2_decap_8 FILLER_11_722 ();
 sg13g2_decap_4 FILLER_11_729 ();
 sg13g2_fill_1 FILLER_11_733 ();
 sg13g2_fill_1 FILLER_11_758 ();
 sg13g2_fill_1 FILLER_11_767 ();
 sg13g2_fill_2 FILLER_11_801 ();
 sg13g2_fill_1 FILLER_11_803 ();
 sg13g2_fill_2 FILLER_11_808 ();
 sg13g2_fill_1 FILLER_11_810 ();
 sg13g2_fill_2 FILLER_11_815 ();
 sg13g2_decap_8 FILLER_11_829 ();
 sg13g2_decap_8 FILLER_11_836 ();
 sg13g2_decap_8 FILLER_11_843 ();
 sg13g2_decap_8 FILLER_11_850 ();
 sg13g2_decap_8 FILLER_11_857 ();
 sg13g2_decap_8 FILLER_11_864 ();
 sg13g2_decap_8 FILLER_11_871 ();
 sg13g2_fill_1 FILLER_12_26 ();
 sg13g2_decap_4 FILLER_12_31 ();
 sg13g2_fill_1 FILLER_12_46 ();
 sg13g2_decap_8 FILLER_12_54 ();
 sg13g2_decap_4 FILLER_12_61 ();
 sg13g2_fill_2 FILLER_12_65 ();
 sg13g2_fill_2 FILLER_12_83 ();
 sg13g2_fill_1 FILLER_12_85 ();
 sg13g2_decap_8 FILLER_12_90 ();
 sg13g2_decap_8 FILLER_12_117 ();
 sg13g2_decap_8 FILLER_12_128 ();
 sg13g2_decap_8 FILLER_12_135 ();
 sg13g2_fill_2 FILLER_12_165 ();
 sg13g2_fill_1 FILLER_12_167 ();
 sg13g2_fill_1 FILLER_12_173 ();
 sg13g2_fill_2 FILLER_12_180 ();
 sg13g2_fill_1 FILLER_12_182 ();
 sg13g2_fill_1 FILLER_12_187 ();
 sg13g2_fill_1 FILLER_12_197 ();
 sg13g2_fill_1 FILLER_12_210 ();
 sg13g2_decap_4 FILLER_12_216 ();
 sg13g2_decap_8 FILLER_12_224 ();
 sg13g2_fill_2 FILLER_12_231 ();
 sg13g2_fill_1 FILLER_12_233 ();
 sg13g2_decap_8 FILLER_12_244 ();
 sg13g2_decap_8 FILLER_12_268 ();
 sg13g2_decap_8 FILLER_12_275 ();
 sg13g2_fill_2 FILLER_12_282 ();
 sg13g2_decap_8 FILLER_12_288 ();
 sg13g2_decap_8 FILLER_12_295 ();
 sg13g2_fill_2 FILLER_12_302 ();
 sg13g2_fill_2 FILLER_12_309 ();
 sg13g2_fill_1 FILLER_12_311 ();
 sg13g2_fill_2 FILLER_12_317 ();
 sg13g2_fill_1 FILLER_12_319 ();
 sg13g2_decap_8 FILLER_12_325 ();
 sg13g2_decap_8 FILLER_12_332 ();
 sg13g2_fill_1 FILLER_12_344 ();
 sg13g2_decap_8 FILLER_12_349 ();
 sg13g2_fill_2 FILLER_12_361 ();
 sg13g2_decap_8 FILLER_12_393 ();
 sg13g2_decap_8 FILLER_12_400 ();
 sg13g2_decap_4 FILLER_12_407 ();
 sg13g2_decap_8 FILLER_12_447 ();
 sg13g2_decap_8 FILLER_12_454 ();
 sg13g2_decap_8 FILLER_12_461 ();
 sg13g2_decap_8 FILLER_12_468 ();
 sg13g2_decap_8 FILLER_12_483 ();
 sg13g2_decap_4 FILLER_12_490 ();
 sg13g2_decap_8 FILLER_12_498 ();
 sg13g2_decap_8 FILLER_12_505 ();
 sg13g2_decap_4 FILLER_12_512 ();
 sg13g2_decap_4 FILLER_12_520 ();
 sg13g2_fill_1 FILLER_12_524 ();
 sg13g2_decap_8 FILLER_12_535 ();
 sg13g2_fill_2 FILLER_12_542 ();
 sg13g2_decap_4 FILLER_12_559 ();
 sg13g2_fill_2 FILLER_12_579 ();
 sg13g2_fill_1 FILLER_12_581 ();
 sg13g2_decap_4 FILLER_12_597 ();
 sg13g2_decap_8 FILLER_12_633 ();
 sg13g2_fill_1 FILLER_12_640 ();
 sg13g2_decap_8 FILLER_12_647 ();
 sg13g2_decap_4 FILLER_12_654 ();
 sg13g2_fill_1 FILLER_12_658 ();
 sg13g2_decap_8 FILLER_12_664 ();
 sg13g2_decap_4 FILLER_12_671 ();
 sg13g2_fill_2 FILLER_12_683 ();
 sg13g2_fill_1 FILLER_12_685 ();
 sg13g2_decap_8 FILLER_12_694 ();
 sg13g2_decap_8 FILLER_12_701 ();
 sg13g2_fill_1 FILLER_12_712 ();
 sg13g2_decap_8 FILLER_12_717 ();
 sg13g2_fill_2 FILLER_12_740 ();
 sg13g2_fill_1 FILLER_12_760 ();
 sg13g2_fill_2 FILLER_12_765 ();
 sg13g2_fill_1 FILLER_12_773 ();
 sg13g2_decap_4 FILLER_12_783 ();
 sg13g2_fill_1 FILLER_12_787 ();
 sg13g2_fill_1 FILLER_12_792 ();
 sg13g2_fill_2 FILLER_12_798 ();
 sg13g2_fill_2 FILLER_12_804 ();
 sg13g2_fill_1 FILLER_12_806 ();
 sg13g2_fill_1 FILLER_12_816 ();
 sg13g2_fill_2 FILLER_12_821 ();
 sg13g2_decap_8 FILLER_12_828 ();
 sg13g2_decap_8 FILLER_12_835 ();
 sg13g2_decap_8 FILLER_12_842 ();
 sg13g2_decap_8 FILLER_12_849 ();
 sg13g2_decap_8 FILLER_12_856 ();
 sg13g2_decap_8 FILLER_12_863 ();
 sg13g2_decap_8 FILLER_12_870 ();
 sg13g2_fill_1 FILLER_12_877 ();
 sg13g2_decap_8 FILLER_13_0 ();
 sg13g2_decap_8 FILLER_13_11 ();
 sg13g2_decap_8 FILLER_13_18 ();
 sg13g2_decap_8 FILLER_13_25 ();
 sg13g2_decap_4 FILLER_13_32 ();
 sg13g2_decap_8 FILLER_13_49 ();
 sg13g2_decap_8 FILLER_13_56 ();
 sg13g2_decap_8 FILLER_13_83 ();
 sg13g2_decap_8 FILLER_13_90 ();
 sg13g2_decap_4 FILLER_13_97 ();
 sg13g2_fill_2 FILLER_13_101 ();
 sg13g2_fill_1 FILLER_13_106 ();
 sg13g2_decap_8 FILLER_13_111 ();
 sg13g2_fill_1 FILLER_13_118 ();
 sg13g2_decap_4 FILLER_13_145 ();
 sg13g2_fill_1 FILLER_13_149 ();
 sg13g2_fill_1 FILLER_13_155 ();
 sg13g2_decap_8 FILLER_13_160 ();
 sg13g2_decap_4 FILLER_13_167 ();
 sg13g2_fill_2 FILLER_13_171 ();
 sg13g2_fill_1 FILLER_13_178 ();
 sg13g2_fill_2 FILLER_13_183 ();
 sg13g2_fill_1 FILLER_13_185 ();
 sg13g2_decap_4 FILLER_13_191 ();
 sg13g2_fill_1 FILLER_13_200 ();
 sg13g2_fill_2 FILLER_13_205 ();
 sg13g2_decap_4 FILLER_13_211 ();
 sg13g2_fill_2 FILLER_13_215 ();
 sg13g2_decap_8 FILLER_13_226 ();
 sg13g2_decap_4 FILLER_13_233 ();
 sg13g2_fill_1 FILLER_13_237 ();
 sg13g2_decap_8 FILLER_13_243 ();
 sg13g2_fill_2 FILLER_13_317 ();
 sg13g2_fill_2 FILLER_13_324 ();
 sg13g2_decap_8 FILLER_13_330 ();
 sg13g2_decap_4 FILLER_13_337 ();
 sg13g2_fill_2 FILLER_13_341 ();
 sg13g2_decap_4 FILLER_13_348 ();
 sg13g2_decap_4 FILLER_13_383 ();
 sg13g2_fill_1 FILLER_13_387 ();
 sg13g2_decap_4 FILLER_13_393 ();
 sg13g2_fill_2 FILLER_13_397 ();
 sg13g2_fill_1 FILLER_13_403 ();
 sg13g2_fill_1 FILLER_13_409 ();
 sg13g2_fill_2 FILLER_13_414 ();
 sg13g2_fill_2 FILLER_13_421 ();
 sg13g2_fill_1 FILLER_13_423 ();
 sg13g2_fill_1 FILLER_13_429 ();
 sg13g2_decap_8 FILLER_13_434 ();
 sg13g2_fill_2 FILLER_13_441 ();
 sg13g2_fill_1 FILLER_13_443 ();
 sg13g2_decap_4 FILLER_13_449 ();
 sg13g2_fill_1 FILLER_13_453 ();
 sg13g2_fill_1 FILLER_13_458 ();
 sg13g2_decap_8 FILLER_13_467 ();
 sg13g2_decap_8 FILLER_13_474 ();
 sg13g2_decap_8 FILLER_13_481 ();
 sg13g2_decap_8 FILLER_13_488 ();
 sg13g2_decap_8 FILLER_13_495 ();
 sg13g2_decap_8 FILLER_13_502 ();
 sg13g2_decap_8 FILLER_13_509 ();
 sg13g2_decap_4 FILLER_13_520 ();
 sg13g2_fill_2 FILLER_13_536 ();
 sg13g2_fill_2 FILLER_13_542 ();
 sg13g2_fill_1 FILLER_13_555 ();
 sg13g2_fill_1 FILLER_13_572 ();
 sg13g2_fill_1 FILLER_13_583 ();
 sg13g2_fill_1 FILLER_13_595 ();
 sg13g2_decap_4 FILLER_13_604 ();
 sg13g2_fill_1 FILLER_13_608 ();
 sg13g2_fill_2 FILLER_13_614 ();
 sg13g2_fill_1 FILLER_13_616 ();
 sg13g2_fill_2 FILLER_13_621 ();
 sg13g2_fill_1 FILLER_13_623 ();
 sg13g2_fill_2 FILLER_13_635 ();
 sg13g2_fill_1 FILLER_13_637 ();
 sg13g2_fill_1 FILLER_13_642 ();
 sg13g2_decap_4 FILLER_13_653 ();
 sg13g2_fill_1 FILLER_13_657 ();
 sg13g2_decap_8 FILLER_13_670 ();
 sg13g2_decap_4 FILLER_13_677 ();
 sg13g2_fill_2 FILLER_13_689 ();
 sg13g2_fill_1 FILLER_13_691 ();
 sg13g2_decap_8 FILLER_13_697 ();
 sg13g2_fill_1 FILLER_13_709 ();
 sg13g2_decap_8 FILLER_13_715 ();
 sg13g2_decap_8 FILLER_13_722 ();
 sg13g2_decap_4 FILLER_13_729 ();
 sg13g2_fill_2 FILLER_13_762 ();
 sg13g2_decap_4 FILLER_13_770 ();
 sg13g2_fill_2 FILLER_13_774 ();
 sg13g2_fill_2 FILLER_13_786 ();
 sg13g2_decap_4 FILLER_13_794 ();
 sg13g2_decap_4 FILLER_13_808 ();
 sg13g2_fill_2 FILLER_13_812 ();
 sg13g2_decap_8 FILLER_13_829 ();
 sg13g2_decap_8 FILLER_13_836 ();
 sg13g2_decap_8 FILLER_13_843 ();
 sg13g2_decap_8 FILLER_13_850 ();
 sg13g2_decap_8 FILLER_13_857 ();
 sg13g2_decap_8 FILLER_13_864 ();
 sg13g2_decap_8 FILLER_13_871 ();
 sg13g2_decap_4 FILLER_14_0 ();
 sg13g2_decap_8 FILLER_14_51 ();
 sg13g2_fill_1 FILLER_14_58 ();
 sg13g2_fill_1 FILLER_14_81 ();
 sg13g2_decap_8 FILLER_14_86 ();
 sg13g2_decap_8 FILLER_14_119 ();
 sg13g2_fill_2 FILLER_14_126 ();
 sg13g2_fill_1 FILLER_14_128 ();
 sg13g2_decap_8 FILLER_14_133 ();
 sg13g2_decap_4 FILLER_14_140 ();
 sg13g2_fill_2 FILLER_14_148 ();
 sg13g2_fill_1 FILLER_14_150 ();
 sg13g2_decap_8 FILLER_14_155 ();
 sg13g2_decap_8 FILLER_14_162 ();
 sg13g2_decap_4 FILLER_14_169 ();
 sg13g2_fill_1 FILLER_14_173 ();
 sg13g2_decap_4 FILLER_14_191 ();
 sg13g2_fill_1 FILLER_14_195 ();
 sg13g2_decap_8 FILLER_14_243 ();
 sg13g2_decap_4 FILLER_14_250 ();
 sg13g2_fill_2 FILLER_14_254 ();
 sg13g2_decap_4 FILLER_14_260 ();
 sg13g2_fill_2 FILLER_14_264 ();
 sg13g2_decap_8 FILLER_14_274 ();
 sg13g2_fill_2 FILLER_14_281 ();
 sg13g2_decap_8 FILLER_14_287 ();
 sg13g2_decap_8 FILLER_14_294 ();
 sg13g2_decap_4 FILLER_14_301 ();
 sg13g2_fill_1 FILLER_14_305 ();
 sg13g2_decap_4 FILLER_14_311 ();
 sg13g2_fill_1 FILLER_14_315 ();
 sg13g2_decap_8 FILLER_14_346 ();
 sg13g2_decap_4 FILLER_14_353 ();
 sg13g2_fill_1 FILLER_14_357 ();
 sg13g2_decap_4 FILLER_14_362 ();
 sg13g2_decap_8 FILLER_14_373 ();
 sg13g2_decap_4 FILLER_14_380 ();
 sg13g2_fill_2 FILLER_14_384 ();
 sg13g2_fill_2 FILLER_14_391 ();
 sg13g2_fill_1 FILLER_14_393 ();
 sg13g2_decap_8 FILLER_14_420 ();
 sg13g2_decap_4 FILLER_14_427 ();
 sg13g2_fill_2 FILLER_14_436 ();
 sg13g2_fill_1 FILLER_14_442 ();
 sg13g2_decap_8 FILLER_14_453 ();
 sg13g2_fill_2 FILLER_14_460 ();
 sg13g2_decap_8 FILLER_14_487 ();
 sg13g2_decap_8 FILLER_14_494 ();
 sg13g2_decap_8 FILLER_14_510 ();
 sg13g2_decap_8 FILLER_14_517 ();
 sg13g2_decap_4 FILLER_14_524 ();
 sg13g2_decap_8 FILLER_14_548 ();
 sg13g2_fill_1 FILLER_14_555 ();
 sg13g2_fill_2 FILLER_14_564 ();
 sg13g2_fill_1 FILLER_14_566 ();
 sg13g2_decap_8 FILLER_14_573 ();
 sg13g2_fill_1 FILLER_14_580 ();
 sg13g2_decap_4 FILLER_14_592 ();
 sg13g2_fill_1 FILLER_14_596 ();
 sg13g2_fill_2 FILLER_14_605 ();
 sg13g2_fill_1 FILLER_14_607 ();
 sg13g2_fill_1 FILLER_14_619 ();
 sg13g2_fill_2 FILLER_14_625 ();
 sg13g2_fill_1 FILLER_14_627 ();
 sg13g2_decap_4 FILLER_14_633 ();
 sg13g2_decap_8 FILLER_14_645 ();
 sg13g2_decap_8 FILLER_14_652 ();
 sg13g2_fill_1 FILLER_14_659 ();
 sg13g2_fill_1 FILLER_14_672 ();
 sg13g2_fill_2 FILLER_14_678 ();
 sg13g2_fill_2 FILLER_14_694 ();
 sg13g2_fill_1 FILLER_14_749 ();
 sg13g2_decap_4 FILLER_14_754 ();
 sg13g2_decap_4 FILLER_14_767 ();
 sg13g2_decap_4 FILLER_14_781 ();
 sg13g2_fill_1 FILLER_14_785 ();
 sg13g2_fill_2 FILLER_14_793 ();
 sg13g2_fill_2 FILLER_14_799 ();
 sg13g2_fill_1 FILLER_14_801 ();
 sg13g2_fill_2 FILLER_14_815 ();
 sg13g2_fill_1 FILLER_14_817 ();
 sg13g2_fill_2 FILLER_14_822 ();
 sg13g2_fill_1 FILLER_14_824 ();
 sg13g2_decap_8 FILLER_14_829 ();
 sg13g2_decap_8 FILLER_14_836 ();
 sg13g2_decap_8 FILLER_14_843 ();
 sg13g2_decap_8 FILLER_14_850 ();
 sg13g2_decap_8 FILLER_14_857 ();
 sg13g2_decap_8 FILLER_14_864 ();
 sg13g2_decap_8 FILLER_14_871 ();
 sg13g2_decap_8 FILLER_15_0 ();
 sg13g2_decap_4 FILLER_15_7 ();
 sg13g2_decap_8 FILLER_15_15 ();
 sg13g2_decap_8 FILLER_15_22 ();
 sg13g2_decap_4 FILLER_15_29 ();
 sg13g2_fill_2 FILLER_15_33 ();
 sg13g2_decap_8 FILLER_15_55 ();
 sg13g2_fill_2 FILLER_15_62 ();
 sg13g2_fill_1 FILLER_15_76 ();
 sg13g2_decap_8 FILLER_15_82 ();
 sg13g2_decap_4 FILLER_15_89 ();
 sg13g2_fill_1 FILLER_15_93 ();
 sg13g2_decap_4 FILLER_15_98 ();
 sg13g2_decap_4 FILLER_15_106 ();
 sg13g2_decap_4 FILLER_15_114 ();
 sg13g2_decap_4 FILLER_15_163 ();
 sg13g2_fill_1 FILLER_15_167 ();
 sg13g2_fill_1 FILLER_15_172 ();
 sg13g2_decap_8 FILLER_15_191 ();
 sg13g2_decap_4 FILLER_15_203 ();
 sg13g2_fill_2 FILLER_15_207 ();
 sg13g2_decap_4 FILLER_15_218 ();
 sg13g2_fill_2 FILLER_15_222 ();
 sg13g2_decap_8 FILLER_15_228 ();
 sg13g2_decap_4 FILLER_15_235 ();
 sg13g2_decap_4 FILLER_15_243 ();
 sg13g2_fill_2 FILLER_15_252 ();
 sg13g2_fill_2 FILLER_15_259 ();
 sg13g2_fill_1 FILLER_15_261 ();
 sg13g2_decap_8 FILLER_15_266 ();
 sg13g2_decap_8 FILLER_15_273 ();
 sg13g2_decap_8 FILLER_15_280 ();
 sg13g2_fill_2 FILLER_15_287 ();
 sg13g2_fill_1 FILLER_15_289 ();
 sg13g2_decap_8 FILLER_15_294 ();
 sg13g2_fill_2 FILLER_15_301 ();
 sg13g2_fill_1 FILLER_15_303 ();
 sg13g2_fill_1 FILLER_15_313 ();
 sg13g2_fill_2 FILLER_15_319 ();
 sg13g2_fill_2 FILLER_15_326 ();
 sg13g2_decap_4 FILLER_15_332 ();
 sg13g2_decap_8 FILLER_15_340 ();
 sg13g2_fill_1 FILLER_15_365 ();
 sg13g2_fill_1 FILLER_15_371 ();
 sg13g2_fill_2 FILLER_15_376 ();
 sg13g2_decap_4 FILLER_15_383 ();
 sg13g2_fill_2 FILLER_15_392 ();
 sg13g2_fill_1 FILLER_15_394 ();
 sg13g2_fill_2 FILLER_15_399 ();
 sg13g2_decap_8 FILLER_15_405 ();
 sg13g2_decap_8 FILLER_15_412 ();
 sg13g2_decap_4 FILLER_15_419 ();
 sg13g2_fill_2 FILLER_15_423 ();
 sg13g2_decap_4 FILLER_15_444 ();
 sg13g2_decap_4 FILLER_15_455 ();
 sg13g2_fill_1 FILLER_15_459 ();
 sg13g2_fill_2 FILLER_15_465 ();
 sg13g2_decap_4 FILLER_15_477 ();
 sg13g2_fill_1 FILLER_15_481 ();
 sg13g2_decap_8 FILLER_15_488 ();
 sg13g2_decap_8 FILLER_15_495 ();
 sg13g2_decap_4 FILLER_15_507 ();
 sg13g2_decap_8 FILLER_15_519 ();
 sg13g2_decap_8 FILLER_15_526 ();
 sg13g2_fill_2 FILLER_15_533 ();
 sg13g2_fill_1 FILLER_15_535 ();
 sg13g2_fill_1 FILLER_15_540 ();
 sg13g2_fill_2 FILLER_15_546 ();
 sg13g2_fill_2 FILLER_15_553 ();
 sg13g2_decap_8 FILLER_15_559 ();
 sg13g2_decap_8 FILLER_15_566 ();
 sg13g2_fill_1 FILLER_15_573 ();
 sg13g2_decap_4 FILLER_15_609 ();
 sg13g2_fill_2 FILLER_15_613 ();
 sg13g2_decap_4 FILLER_15_620 ();
 sg13g2_fill_2 FILLER_15_629 ();
 sg13g2_fill_1 FILLER_15_631 ();
 sg13g2_fill_2 FILLER_15_636 ();
 sg13g2_fill_1 FILLER_15_638 ();
 sg13g2_fill_2 FILLER_15_645 ();
 sg13g2_fill_1 FILLER_15_652 ();
 sg13g2_decap_8 FILLER_15_658 ();
 sg13g2_fill_2 FILLER_15_671 ();
 sg13g2_fill_1 FILLER_15_673 ();
 sg13g2_fill_1 FILLER_15_682 ();
 sg13g2_fill_1 FILLER_15_692 ();
 sg13g2_fill_1 FILLER_15_697 ();
 sg13g2_fill_2 FILLER_15_703 ();
 sg13g2_decap_8 FILLER_15_712 ();
 sg13g2_decap_4 FILLER_15_719 ();
 sg13g2_fill_2 FILLER_15_723 ();
 sg13g2_fill_1 FILLER_15_730 ();
 sg13g2_decap_4 FILLER_15_745 ();
 sg13g2_fill_1 FILLER_15_749 ();
 sg13g2_fill_2 FILLER_15_760 ();
 sg13g2_fill_1 FILLER_15_762 ();
 sg13g2_decap_4 FILLER_15_768 ();
 sg13g2_fill_1 FILLER_15_772 ();
 sg13g2_fill_1 FILLER_15_785 ();
 sg13g2_decap_8 FILLER_15_794 ();
 sg13g2_fill_2 FILLER_15_808 ();
 sg13g2_decap_8 FILLER_15_815 ();
 sg13g2_decap_8 FILLER_15_822 ();
 sg13g2_decap_8 FILLER_15_829 ();
 sg13g2_decap_8 FILLER_15_836 ();
 sg13g2_decap_8 FILLER_15_843 ();
 sg13g2_decap_8 FILLER_15_850 ();
 sg13g2_decap_8 FILLER_15_857 ();
 sg13g2_decap_8 FILLER_15_864 ();
 sg13g2_decap_8 FILLER_15_871 ();
 sg13g2_decap_8 FILLER_16_0 ();
 sg13g2_fill_1 FILLER_16_7 ();
 sg13g2_decap_8 FILLER_16_20 ();
 sg13g2_decap_8 FILLER_16_27 ();
 sg13g2_fill_2 FILLER_16_34 ();
 sg13g2_fill_1 FILLER_16_36 ();
 sg13g2_decap_8 FILLER_16_49 ();
 sg13g2_fill_2 FILLER_16_56 ();
 sg13g2_fill_2 FILLER_16_77 ();
 sg13g2_decap_8 FILLER_16_84 ();
 sg13g2_fill_2 FILLER_16_91 ();
 sg13g2_fill_1 FILLER_16_93 ();
 sg13g2_fill_1 FILLER_16_102 ();
 sg13g2_decap_8 FILLER_16_149 ();
 sg13g2_fill_1 FILLER_16_156 ();
 sg13g2_decap_4 FILLER_16_162 ();
 sg13g2_fill_2 FILLER_16_166 ();
 sg13g2_decap_8 FILLER_16_173 ();
 sg13g2_decap_8 FILLER_16_180 ();
 sg13g2_decap_8 FILLER_16_187 ();
 sg13g2_decap_4 FILLER_16_194 ();
 sg13g2_decap_4 FILLER_16_202 ();
 sg13g2_decap_4 FILLER_16_220 ();
 sg13g2_decap_8 FILLER_16_228 ();
 sg13g2_decap_8 FILLER_16_235 ();
 sg13g2_decap_4 FILLER_16_242 ();
 sg13g2_fill_2 FILLER_16_281 ();
 sg13g2_decap_8 FILLER_16_309 ();
 sg13g2_decap_4 FILLER_16_316 ();
 sg13g2_fill_2 FILLER_16_353 ();
 sg13g2_fill_1 FILLER_16_355 ();
 sg13g2_fill_1 FILLER_16_382 ();
 sg13g2_decap_8 FILLER_16_414 ();
 sg13g2_fill_1 FILLER_16_421 ();
 sg13g2_fill_2 FILLER_16_427 ();
 sg13g2_decap_8 FILLER_16_448 ();
 sg13g2_fill_2 FILLER_16_455 ();
 sg13g2_fill_1 FILLER_16_465 ();
 sg13g2_decap_4 FILLER_16_470 ();
 sg13g2_fill_2 FILLER_16_484 ();
 sg13g2_decap_8 FILLER_16_499 ();
 sg13g2_decap_8 FILLER_16_506 ();
 sg13g2_decap_8 FILLER_16_513 ();
 sg13g2_decap_8 FILLER_16_520 ();
 sg13g2_fill_1 FILLER_16_527 ();
 sg13g2_decap_8 FILLER_16_558 ();
 sg13g2_decap_8 FILLER_16_565 ();
 sg13g2_decap_4 FILLER_16_572 ();
 sg13g2_fill_1 FILLER_16_576 ();
 sg13g2_decap_8 FILLER_16_582 ();
 sg13g2_fill_2 FILLER_16_589 ();
 sg13g2_decap_8 FILLER_16_596 ();
 sg13g2_fill_2 FILLER_16_603 ();
 sg13g2_fill_1 FILLER_16_605 ();
 sg13g2_decap_8 FILLER_16_618 ();
 sg13g2_fill_1 FILLER_16_625 ();
 sg13g2_fill_2 FILLER_16_637 ();
 sg13g2_fill_1 FILLER_16_639 ();
 sg13g2_fill_1 FILLER_16_653 ();
 sg13g2_decap_4 FILLER_16_659 ();
 sg13g2_fill_2 FILLER_16_663 ();
 sg13g2_fill_2 FILLER_16_679 ();
 sg13g2_fill_1 FILLER_16_681 ();
 sg13g2_fill_1 FILLER_16_694 ();
 sg13g2_fill_2 FILLER_16_707 ();
 sg13g2_decap_8 FILLER_16_728 ();
 sg13g2_decap_4 FILLER_16_735 ();
 sg13g2_decap_4 FILLER_16_743 ();
 sg13g2_fill_2 FILLER_16_747 ();
 sg13g2_decap_4 FILLER_16_754 ();
 sg13g2_fill_2 FILLER_16_758 ();
 sg13g2_decap_8 FILLER_16_768 ();
 sg13g2_fill_2 FILLER_16_775 ();
 sg13g2_fill_1 FILLER_16_777 ();
 sg13g2_decap_8 FILLER_16_796 ();
 sg13g2_decap_4 FILLER_16_803 ();
 sg13g2_fill_2 FILLER_16_807 ();
 sg13g2_fill_1 FILLER_16_813 ();
 sg13g2_decap_8 FILLER_16_822 ();
 sg13g2_decap_8 FILLER_16_829 ();
 sg13g2_decap_8 FILLER_16_836 ();
 sg13g2_decap_8 FILLER_16_843 ();
 sg13g2_decap_8 FILLER_16_850 ();
 sg13g2_decap_8 FILLER_16_857 ();
 sg13g2_decap_8 FILLER_16_864 ();
 sg13g2_decap_8 FILLER_16_871 ();
 sg13g2_decap_4 FILLER_17_0 ();
 sg13g2_fill_1 FILLER_17_34 ();
 sg13g2_decap_4 FILLER_17_39 ();
 sg13g2_decap_8 FILLER_17_47 ();
 sg13g2_decap_8 FILLER_17_54 ();
 sg13g2_decap_4 FILLER_17_61 ();
 sg13g2_decap_8 FILLER_17_81 ();
 sg13g2_decap_4 FILLER_17_88 ();
 sg13g2_fill_1 FILLER_17_92 ();
 sg13g2_decap_8 FILLER_17_108 ();
 sg13g2_decap_8 FILLER_17_115 ();
 sg13g2_decap_4 FILLER_17_122 ();
 sg13g2_fill_2 FILLER_17_126 ();
 sg13g2_decap_8 FILLER_17_138 ();
 sg13g2_decap_8 FILLER_17_145 ();
 sg13g2_decap_8 FILLER_17_152 ();
 sg13g2_decap_8 FILLER_17_159 ();
 sg13g2_decap_8 FILLER_17_166 ();
 sg13g2_decap_8 FILLER_17_173 ();
 sg13g2_decap_8 FILLER_17_180 ();
 sg13g2_fill_1 FILLER_17_187 ();
 sg13g2_fill_1 FILLER_17_198 ();
 sg13g2_fill_1 FILLER_17_209 ();
 sg13g2_decap_8 FILLER_17_242 ();
 sg13g2_decap_8 FILLER_17_249 ();
 sg13g2_decap_4 FILLER_17_256 ();
 sg13g2_decap_4 FILLER_17_269 ();
 sg13g2_fill_1 FILLER_17_277 ();
 sg13g2_decap_8 FILLER_17_289 ();
 sg13g2_decap_8 FILLER_17_296 ();
 sg13g2_decap_8 FILLER_17_303 ();
 sg13g2_decap_8 FILLER_17_310 ();
 sg13g2_decap_8 FILLER_17_317 ();
 sg13g2_decap_4 FILLER_17_324 ();
 sg13g2_fill_1 FILLER_17_328 ();
 sg13g2_fill_1 FILLER_17_334 ();
 sg13g2_decap_8 FILLER_17_339 ();
 sg13g2_decap_8 FILLER_17_346 ();
 sg13g2_decap_8 FILLER_17_353 ();
 sg13g2_fill_2 FILLER_17_360 ();
 sg13g2_fill_1 FILLER_17_362 ();
 sg13g2_decap_8 FILLER_17_367 ();
 sg13g2_decap_8 FILLER_17_374 ();
 sg13g2_decap_4 FILLER_17_381 ();
 sg13g2_fill_1 FILLER_17_385 ();
 sg13g2_decap_8 FILLER_17_391 ();
 sg13g2_fill_2 FILLER_17_398 ();
 sg13g2_fill_1 FILLER_17_400 ();
 sg13g2_decap_8 FILLER_17_406 ();
 sg13g2_decap_8 FILLER_17_413 ();
 sg13g2_decap_8 FILLER_17_424 ();
 sg13g2_decap_8 FILLER_17_431 ();
 sg13g2_decap_4 FILLER_17_438 ();
 sg13g2_decap_8 FILLER_17_450 ();
 sg13g2_fill_1 FILLER_17_457 ();
 sg13g2_fill_2 FILLER_17_463 ();
 sg13g2_decap_4 FILLER_17_482 ();
 sg13g2_decap_8 FILLER_17_494 ();
 sg13g2_decap_4 FILLER_17_501 ();
 sg13g2_fill_2 FILLER_17_505 ();
 sg13g2_decap_8 FILLER_17_512 ();
 sg13g2_fill_2 FILLER_17_519 ();
 sg13g2_decap_8 FILLER_17_526 ();
 sg13g2_decap_8 FILLER_17_533 ();
 sg13g2_fill_2 FILLER_17_540 ();
 sg13g2_fill_2 FILLER_17_555 ();
 sg13g2_decap_8 FILLER_17_562 ();
 sg13g2_decap_8 FILLER_17_569 ();
 sg13g2_decap_8 FILLER_17_576 ();
 sg13g2_decap_8 FILLER_17_583 ();
 sg13g2_decap_4 FILLER_17_607 ();
 sg13g2_fill_1 FILLER_17_620 ();
 sg13g2_fill_2 FILLER_17_625 ();
 sg13g2_decap_8 FILLER_17_631 ();
 sg13g2_fill_1 FILLER_17_638 ();
 sg13g2_fill_1 FILLER_17_645 ();
 sg13g2_decap_4 FILLER_17_650 ();
 sg13g2_decap_8 FILLER_17_664 ();
 sg13g2_fill_1 FILLER_17_671 ();
 sg13g2_decap_8 FILLER_17_681 ();
 sg13g2_decap_8 FILLER_17_688 ();
 sg13g2_decap_4 FILLER_17_695 ();
 sg13g2_fill_1 FILLER_17_699 ();
 sg13g2_decap_8 FILLER_17_719 ();
 sg13g2_decap_8 FILLER_17_726 ();
 sg13g2_decap_8 FILLER_17_733 ();
 sg13g2_fill_2 FILLER_17_740 ();
 sg13g2_decap_4 FILLER_17_755 ();
 sg13g2_fill_2 FILLER_17_759 ();
 sg13g2_decap_8 FILLER_17_765 ();
 sg13g2_fill_2 FILLER_17_772 ();
 sg13g2_decap_8 FILLER_17_779 ();
 sg13g2_decap_8 FILLER_17_786 ();
 sg13g2_decap_4 FILLER_17_793 ();
 sg13g2_fill_2 FILLER_17_797 ();
 sg13g2_decap_8 FILLER_17_803 ();
 sg13g2_fill_2 FILLER_17_810 ();
 sg13g2_fill_1 FILLER_17_812 ();
 sg13g2_fill_1 FILLER_17_817 ();
 sg13g2_decap_8 FILLER_17_823 ();
 sg13g2_decap_8 FILLER_17_830 ();
 sg13g2_decap_8 FILLER_17_837 ();
 sg13g2_decap_8 FILLER_17_844 ();
 sg13g2_decap_8 FILLER_17_851 ();
 sg13g2_decap_8 FILLER_17_858 ();
 sg13g2_decap_8 FILLER_17_865 ();
 sg13g2_decap_4 FILLER_17_872 ();
 sg13g2_fill_2 FILLER_17_876 ();
 sg13g2_decap_8 FILLER_18_0 ();
 sg13g2_fill_1 FILLER_18_7 ();
 sg13g2_decap_8 FILLER_18_18 ();
 sg13g2_decap_4 FILLER_18_25 ();
 sg13g2_fill_2 FILLER_18_29 ();
 sg13g2_fill_2 FILLER_18_40 ();
 sg13g2_decap_8 FILLER_18_59 ();
 sg13g2_decap_8 FILLER_18_66 ();
 sg13g2_fill_1 FILLER_18_73 ();
 sg13g2_decap_8 FILLER_18_82 ();
 sg13g2_fill_2 FILLER_18_89 ();
 sg13g2_fill_1 FILLER_18_91 ();
 sg13g2_fill_1 FILLER_18_96 ();
 sg13g2_fill_1 FILLER_18_102 ();
 sg13g2_fill_1 FILLER_18_108 ();
 sg13g2_decap_4 FILLER_18_112 ();
 sg13g2_decap_4 FILLER_18_119 ();
 sg13g2_fill_1 FILLER_18_123 ();
 sg13g2_decap_4 FILLER_18_134 ();
 sg13g2_decap_4 FILLER_18_174 ();
 sg13g2_fill_2 FILLER_18_178 ();
 sg13g2_decap_8 FILLER_18_221 ();
 sg13g2_decap_8 FILLER_18_228 ();
 sg13g2_fill_2 FILLER_18_235 ();
 sg13g2_decap_4 FILLER_18_241 ();
 sg13g2_fill_1 FILLER_18_245 ();
 sg13g2_decap_8 FILLER_18_250 ();
 sg13g2_fill_2 FILLER_18_257 ();
 sg13g2_fill_1 FILLER_18_285 ();
 sg13g2_fill_2 FILLER_18_312 ();
 sg13g2_fill_1 FILLER_18_319 ();
 sg13g2_fill_2 FILLER_18_325 ();
 sg13g2_fill_2 FILLER_18_364 ();
 sg13g2_decap_8 FILLER_18_396 ();
 sg13g2_decap_8 FILLER_18_424 ();
 sg13g2_decap_8 FILLER_18_431 ();
 sg13g2_fill_2 FILLER_18_438 ();
 sg13g2_fill_1 FILLER_18_466 ();
 sg13g2_fill_2 FILLER_18_484 ();
 sg13g2_decap_8 FILLER_18_489 ();
 sg13g2_fill_1 FILLER_18_496 ();
 sg13g2_decap_8 FILLER_18_525 ();
 sg13g2_decap_4 FILLER_18_532 ();
 sg13g2_fill_1 FILLER_18_536 ();
 sg13g2_decap_8 FILLER_18_547 ();
 sg13g2_fill_2 FILLER_18_554 ();
 sg13g2_decap_8 FILLER_18_581 ();
 sg13g2_fill_1 FILLER_18_588 ();
 sg13g2_decap_8 FILLER_18_604 ();
 sg13g2_decap_8 FILLER_18_611 ();
 sg13g2_decap_8 FILLER_18_618 ();
 sg13g2_decap_8 FILLER_18_625 ();
 sg13g2_fill_2 FILLER_18_632 ();
 sg13g2_fill_1 FILLER_18_634 ();
 sg13g2_decap_4 FILLER_18_644 ();
 sg13g2_fill_1 FILLER_18_648 ();
 sg13g2_decap_8 FILLER_18_658 ();
 sg13g2_decap_8 FILLER_18_665 ();
 sg13g2_decap_8 FILLER_18_672 ();
 sg13g2_decap_4 FILLER_18_679 ();
 sg13g2_decap_8 FILLER_18_687 ();
 sg13g2_fill_1 FILLER_18_694 ();
 sg13g2_fill_1 FILLER_18_705 ();
 sg13g2_decap_4 FILLER_18_739 ();
 sg13g2_fill_1 FILLER_18_743 ();
 sg13g2_fill_2 FILLER_18_754 ();
 sg13g2_decap_8 FILLER_18_767 ();
 sg13g2_decap_4 FILLER_18_774 ();
 sg13g2_fill_1 FILLER_18_778 ();
 sg13g2_fill_1 FILLER_18_788 ();
 sg13g2_fill_1 FILLER_18_795 ();
 sg13g2_fill_1 FILLER_18_802 ();
 sg13g2_decap_8 FILLER_18_814 ();
 sg13g2_decap_8 FILLER_18_821 ();
 sg13g2_decap_8 FILLER_18_828 ();
 sg13g2_decap_8 FILLER_18_835 ();
 sg13g2_decap_8 FILLER_18_842 ();
 sg13g2_decap_8 FILLER_18_849 ();
 sg13g2_decap_8 FILLER_18_856 ();
 sg13g2_decap_8 FILLER_18_863 ();
 sg13g2_decap_8 FILLER_18_870 ();
 sg13g2_fill_1 FILLER_18_877 ();
 sg13g2_decap_4 FILLER_19_26 ();
 sg13g2_fill_2 FILLER_19_30 ();
 sg13g2_fill_2 FILLER_19_44 ();
 sg13g2_fill_2 FILLER_19_52 ();
 sg13g2_fill_1 FILLER_19_54 ();
 sg13g2_fill_1 FILLER_19_81 ();
 sg13g2_decap_4 FILLER_19_90 ();
 sg13g2_decap_8 FILLER_19_98 ();
 sg13g2_fill_2 FILLER_19_105 ();
 sg13g2_decap_8 FILLER_19_112 ();
 sg13g2_decap_8 FILLER_19_119 ();
 sg13g2_decap_4 FILLER_19_126 ();
 sg13g2_fill_2 FILLER_19_135 ();
 sg13g2_fill_1 FILLER_19_137 ();
 sg13g2_fill_1 FILLER_19_143 ();
 sg13g2_decap_4 FILLER_19_149 ();
 sg13g2_fill_2 FILLER_19_153 ();
 sg13g2_decap_8 FILLER_19_159 ();
 sg13g2_fill_1 FILLER_19_166 ();
 sg13g2_decap_8 FILLER_19_172 ();
 sg13g2_decap_4 FILLER_19_179 ();
 sg13g2_fill_1 FILLER_19_183 ();
 sg13g2_decap_8 FILLER_19_194 ();
 sg13g2_decap_8 FILLER_19_201 ();
 sg13g2_decap_4 FILLER_19_213 ();
 sg13g2_fill_2 FILLER_19_217 ();
 sg13g2_decap_8 FILLER_19_255 ();
 sg13g2_decap_8 FILLER_19_262 ();
 sg13g2_fill_2 FILLER_19_269 ();
 sg13g2_fill_1 FILLER_19_271 ();
 sg13g2_decap_4 FILLER_19_276 ();
 sg13g2_fill_1 FILLER_19_280 ();
 sg13g2_decap_8 FILLER_19_284 ();
 sg13g2_fill_1 FILLER_19_291 ();
 sg13g2_decap_4 FILLER_19_296 ();
 sg13g2_fill_2 FILLER_19_300 ();
 sg13g2_fill_1 FILLER_19_309 ();
 sg13g2_decap_8 FILLER_19_314 ();
 sg13g2_decap_8 FILLER_19_321 ();
 sg13g2_decap_4 FILLER_19_349 ();
 sg13g2_fill_2 FILLER_19_353 ();
 sg13g2_decap_4 FILLER_19_360 ();
 sg13g2_decap_8 FILLER_19_374 ();
 sg13g2_decap_8 FILLER_19_381 ();
 sg13g2_decap_8 FILLER_19_388 ();
 sg13g2_decap_8 FILLER_19_395 ();
 sg13g2_fill_1 FILLER_19_402 ();
 sg13g2_decap_8 FILLER_19_407 ();
 sg13g2_fill_1 FILLER_19_414 ();
 sg13g2_decap_4 FILLER_19_420 ();
 sg13g2_decap_8 FILLER_19_429 ();
 sg13g2_decap_4 FILLER_19_436 ();
 sg13g2_fill_2 FILLER_19_440 ();
 sg13g2_decap_4 FILLER_19_456 ();
 sg13g2_fill_2 FILLER_19_460 ();
 sg13g2_decap_4 FILLER_19_475 ();
 sg13g2_decap_8 FILLER_19_484 ();
 sg13g2_decap_8 FILLER_19_491 ();
 sg13g2_decap_4 FILLER_19_498 ();
 sg13g2_decap_4 FILLER_19_523 ();
 sg13g2_fill_1 FILLER_19_527 ();
 sg13g2_decap_4 FILLER_19_532 ();
 sg13g2_fill_2 FILLER_19_536 ();
 sg13g2_decap_8 FILLER_19_547 ();
 sg13g2_decap_8 FILLER_19_554 ();
 sg13g2_decap_8 FILLER_19_561 ();
 sg13g2_decap_8 FILLER_19_568 ();
 sg13g2_decap_8 FILLER_19_575 ();
 sg13g2_decap_8 FILLER_19_582 ();
 sg13g2_fill_1 FILLER_19_589 ();
 sg13g2_fill_2 FILLER_19_594 ();
 sg13g2_decap_8 FILLER_19_601 ();
 sg13g2_decap_8 FILLER_19_608 ();
 sg13g2_decap_8 FILLER_19_615 ();
 sg13g2_decap_8 FILLER_19_622 ();
 sg13g2_decap_4 FILLER_19_629 ();
 sg13g2_fill_2 FILLER_19_633 ();
 sg13g2_fill_1 FILLER_19_639 ();
 sg13g2_fill_2 FILLER_19_648 ();
 sg13g2_fill_1 FILLER_19_663 ();
 sg13g2_decap_8 FILLER_19_669 ();
 sg13g2_fill_2 FILLER_19_676 ();
 sg13g2_fill_1 FILLER_19_678 ();
 sg13g2_fill_1 FILLER_19_683 ();
 sg13g2_fill_1 FILLER_19_688 ();
 sg13g2_decap_8 FILLER_19_694 ();
 sg13g2_decap_8 FILLER_19_701 ();
 sg13g2_fill_1 FILLER_19_708 ();
 sg13g2_decap_4 FILLER_19_715 ();
 sg13g2_fill_1 FILLER_19_719 ();
 sg13g2_fill_1 FILLER_19_733 ();
 sg13g2_fill_2 FILLER_19_739 ();
 sg13g2_fill_1 FILLER_19_741 ();
 sg13g2_decap_8 FILLER_19_753 ();
 sg13g2_fill_1 FILLER_19_760 ();
 sg13g2_decap_4 FILLER_19_767 ();
 sg13g2_fill_1 FILLER_19_777 ();
 sg13g2_decap_8 FILLER_19_815 ();
 sg13g2_decap_8 FILLER_19_822 ();
 sg13g2_decap_8 FILLER_19_829 ();
 sg13g2_decap_8 FILLER_19_836 ();
 sg13g2_decap_8 FILLER_19_843 ();
 sg13g2_decap_8 FILLER_19_850 ();
 sg13g2_decap_8 FILLER_19_857 ();
 sg13g2_decap_8 FILLER_19_864 ();
 sg13g2_decap_8 FILLER_19_871 ();
 sg13g2_decap_8 FILLER_20_0 ();
 sg13g2_decap_4 FILLER_20_7 ();
 sg13g2_fill_1 FILLER_20_11 ();
 sg13g2_decap_8 FILLER_20_16 ();
 sg13g2_fill_1 FILLER_20_23 ();
 sg13g2_decap_4 FILLER_20_28 ();
 sg13g2_decap_8 FILLER_20_37 ();
 sg13g2_decap_4 FILLER_20_44 ();
 sg13g2_fill_1 FILLER_20_48 ();
 sg13g2_fill_2 FILLER_20_54 ();
 sg13g2_fill_1 FILLER_20_56 ();
 sg13g2_decap_8 FILLER_20_61 ();
 sg13g2_fill_2 FILLER_20_68 ();
 sg13g2_fill_1 FILLER_20_70 ();
 sg13g2_decap_8 FILLER_20_75 ();
 sg13g2_decap_8 FILLER_20_82 ();
 sg13g2_decap_8 FILLER_20_89 ();
 sg13g2_fill_1 FILLER_20_96 ();
 sg13g2_fill_1 FILLER_20_109 ();
 sg13g2_decap_8 FILLER_20_114 ();
 sg13g2_fill_2 FILLER_20_121 ();
 sg13g2_decap_8 FILLER_20_126 ();
 sg13g2_decap_4 FILLER_20_133 ();
 sg13g2_fill_2 FILLER_20_157 ();
 sg13g2_decap_8 FILLER_20_167 ();
 sg13g2_decap_4 FILLER_20_174 ();
 sg13g2_fill_1 FILLER_20_178 ();
 sg13g2_decap_8 FILLER_20_215 ();
 sg13g2_decap_8 FILLER_20_222 ();
 sg13g2_fill_1 FILLER_20_229 ();
 sg13g2_decap_8 FILLER_20_235 ();
 sg13g2_decap_4 FILLER_20_242 ();
 sg13g2_fill_1 FILLER_20_250 ();
 sg13g2_fill_1 FILLER_20_255 ();
 sg13g2_fill_2 FILLER_20_260 ();
 sg13g2_fill_1 FILLER_20_262 ();
 sg13g2_fill_2 FILLER_20_311 ();
 sg13g2_fill_1 FILLER_20_313 ();
 sg13g2_fill_2 FILLER_20_324 ();
 sg13g2_fill_1 FILLER_20_326 ();
 sg13g2_decap_4 FILLER_20_360 ();
 sg13g2_fill_2 FILLER_20_368 ();
 sg13g2_fill_2 FILLER_20_379 ();
 sg13g2_decap_4 FILLER_20_395 ();
 sg13g2_fill_2 FILLER_20_409 ();
 sg13g2_fill_1 FILLER_20_411 ();
 sg13g2_decap_4 FILLER_20_417 ();
 sg13g2_decap_4 FILLER_20_425 ();
 sg13g2_fill_2 FILLER_20_429 ();
 sg13g2_decap_8 FILLER_20_448 ();
 sg13g2_decap_8 FILLER_20_455 ();
 sg13g2_decap_4 FILLER_20_462 ();
 sg13g2_fill_1 FILLER_20_466 ();
 sg13g2_decap_4 FILLER_20_471 ();
 sg13g2_decap_8 FILLER_20_490 ();
 sg13g2_decap_8 FILLER_20_497 ();
 sg13g2_fill_2 FILLER_20_504 ();
 sg13g2_fill_1 FILLER_20_506 ();
 sg13g2_decap_4 FILLER_20_510 ();
 sg13g2_decap_8 FILLER_20_517 ();
 sg13g2_decap_8 FILLER_20_524 ();
 sg13g2_decap_8 FILLER_20_531 ();
 sg13g2_fill_2 FILLER_20_543 ();
 sg13g2_decap_8 FILLER_20_549 ();
 sg13g2_fill_2 FILLER_20_556 ();
 sg13g2_fill_1 FILLER_20_558 ();
 sg13g2_fill_1 FILLER_20_569 ();
 sg13g2_decap_4 FILLER_20_574 ();
 sg13g2_decap_8 FILLER_20_586 ();
 sg13g2_decap_8 FILLER_20_593 ();
 sg13g2_decap_8 FILLER_20_600 ();
 sg13g2_decap_4 FILLER_20_607 ();
 sg13g2_decap_8 FILLER_20_615 ();
 sg13g2_decap_4 FILLER_20_622 ();
 sg13g2_fill_1 FILLER_20_626 ();
 sg13g2_decap_4 FILLER_20_631 ();
 sg13g2_fill_1 FILLER_20_635 ();
 sg13g2_fill_2 FILLER_20_640 ();
 sg13g2_fill_2 FILLER_20_647 ();
 sg13g2_fill_2 FILLER_20_658 ();
 sg13g2_decap_4 FILLER_20_664 ();
 sg13g2_decap_8 FILLER_20_680 ();
 sg13g2_decap_8 FILLER_20_687 ();
 sg13g2_fill_2 FILLER_20_694 ();
 sg13g2_fill_1 FILLER_20_696 ();
 sg13g2_decap_8 FILLER_20_705 ();
 sg13g2_fill_1 FILLER_20_712 ();
 sg13g2_fill_1 FILLER_20_718 ();
 sg13g2_decap_8 FILLER_20_729 ();
 sg13g2_fill_2 FILLER_20_736 ();
 sg13g2_decap_4 FILLER_20_743 ();
 sg13g2_fill_1 FILLER_20_755 ();
 sg13g2_fill_2 FILLER_20_760 ();
 sg13g2_fill_1 FILLER_20_762 ();
 sg13g2_fill_2 FILLER_20_771 ();
 sg13g2_fill_1 FILLER_20_773 ();
 sg13g2_decap_4 FILLER_20_778 ();
 sg13g2_fill_1 FILLER_20_786 ();
 sg13g2_decap_4 FILLER_20_805 ();
 sg13g2_fill_2 FILLER_20_809 ();
 sg13g2_decap_8 FILLER_20_816 ();
 sg13g2_decap_8 FILLER_20_823 ();
 sg13g2_decap_8 FILLER_20_830 ();
 sg13g2_decap_8 FILLER_20_837 ();
 sg13g2_decap_8 FILLER_20_844 ();
 sg13g2_decap_8 FILLER_20_851 ();
 sg13g2_decap_8 FILLER_20_858 ();
 sg13g2_decap_8 FILLER_20_865 ();
 sg13g2_decap_4 FILLER_20_872 ();
 sg13g2_fill_2 FILLER_20_876 ();
 sg13g2_fill_1 FILLER_21_0 ();
 sg13g2_fill_2 FILLER_21_35 ();
 sg13g2_decap_4 FILLER_21_44 ();
 sg13g2_fill_1 FILLER_21_48 ();
 sg13g2_fill_1 FILLER_21_58 ();
 sg13g2_decap_8 FILLER_21_89 ();
 sg13g2_fill_2 FILLER_21_96 ();
 sg13g2_fill_1 FILLER_21_98 ();
 sg13g2_decap_8 FILLER_21_149 ();
 sg13g2_decap_8 FILLER_21_156 ();
 sg13g2_decap_8 FILLER_21_163 ();
 sg13g2_decap_8 FILLER_21_170 ();
 sg13g2_decap_4 FILLER_21_177 ();
 sg13g2_fill_2 FILLER_21_181 ();
 sg13g2_fill_2 FILLER_21_198 ();
 sg13g2_fill_1 FILLER_21_200 ();
 sg13g2_fill_2 FILLER_21_207 ();
 sg13g2_fill_1 FILLER_21_209 ();
 sg13g2_decap_8 FILLER_21_220 ();
 sg13g2_decap_8 FILLER_21_227 ();
 sg13g2_decap_8 FILLER_21_234 ();
 sg13g2_fill_2 FILLER_21_241 ();
 sg13g2_fill_1 FILLER_21_243 ();
 sg13g2_decap_8 FILLER_21_265 ();
 sg13g2_fill_1 FILLER_21_276 ();
 sg13g2_decap_8 FILLER_21_281 ();
 sg13g2_fill_2 FILLER_21_288 ();
 sg13g2_decap_8 FILLER_21_320 ();
 sg13g2_decap_4 FILLER_21_327 ();
 sg13g2_fill_2 FILLER_21_331 ();
 sg13g2_decap_8 FILLER_21_345 ();
 sg13g2_decap_4 FILLER_21_352 ();
 sg13g2_fill_2 FILLER_21_356 ();
 sg13g2_decap_8 FILLER_21_363 ();
 sg13g2_decap_8 FILLER_21_370 ();
 sg13g2_decap_4 FILLER_21_377 ();
 sg13g2_fill_2 FILLER_21_381 ();
 sg13g2_decap_8 FILLER_21_393 ();
 sg13g2_fill_1 FILLER_21_400 ();
 sg13g2_decap_8 FILLER_21_415 ();
 sg13g2_decap_8 FILLER_21_422 ();
 sg13g2_decap_4 FILLER_21_437 ();
 sg13g2_decap_8 FILLER_21_449 ();
 sg13g2_decap_8 FILLER_21_456 ();
 sg13g2_fill_2 FILLER_21_463 ();
 sg13g2_decap_8 FILLER_21_477 ();
 sg13g2_decap_8 FILLER_21_484 ();
 sg13g2_decap_8 FILLER_21_491 ();
 sg13g2_decap_4 FILLER_21_498 ();
 sg13g2_fill_1 FILLER_21_502 ();
 sg13g2_decap_8 FILLER_21_524 ();
 sg13g2_decap_8 FILLER_21_531 ();
 sg13g2_decap_8 FILLER_21_538 ();
 sg13g2_decap_8 FILLER_21_545 ();
 sg13g2_fill_2 FILLER_21_552 ();
 sg13g2_fill_1 FILLER_21_554 ();
 sg13g2_decap_4 FILLER_21_576 ();
 sg13g2_fill_1 FILLER_21_580 ();
 sg13g2_decap_8 FILLER_21_601 ();
 sg13g2_decap_4 FILLER_21_608 ();
 sg13g2_fill_2 FILLER_21_612 ();
 sg13g2_decap_8 FILLER_21_618 ();
 sg13g2_decap_4 FILLER_21_625 ();
 sg13g2_fill_2 FILLER_21_645 ();
 sg13g2_decap_4 FILLER_21_661 ();
 sg13g2_decap_8 FILLER_21_675 ();
 sg13g2_decap_8 FILLER_21_682 ();
 sg13g2_decap_4 FILLER_21_689 ();
 sg13g2_fill_2 FILLER_21_693 ();
 sg13g2_fill_2 FILLER_21_700 ();
 sg13g2_decap_8 FILLER_21_706 ();
 sg13g2_decap_8 FILLER_21_713 ();
 sg13g2_fill_2 FILLER_21_720 ();
 sg13g2_decap_8 FILLER_21_730 ();
 sg13g2_fill_2 FILLER_21_737 ();
 sg13g2_decap_4 FILLER_21_743 ();
 sg13g2_fill_2 FILLER_21_747 ();
 sg13g2_decap_4 FILLER_21_753 ();
 sg13g2_fill_1 FILLER_21_757 ();
 sg13g2_decap_8 FILLER_21_766 ();
 sg13g2_decap_8 FILLER_21_773 ();
 sg13g2_decap_8 FILLER_21_780 ();
 sg13g2_decap_4 FILLER_21_795 ();
 sg13g2_decap_8 FILLER_21_816 ();
 sg13g2_decap_8 FILLER_21_823 ();
 sg13g2_decap_8 FILLER_21_830 ();
 sg13g2_decap_8 FILLER_21_837 ();
 sg13g2_decap_8 FILLER_21_844 ();
 sg13g2_decap_8 FILLER_21_851 ();
 sg13g2_decap_8 FILLER_21_858 ();
 sg13g2_decap_8 FILLER_21_865 ();
 sg13g2_decap_4 FILLER_21_872 ();
 sg13g2_fill_2 FILLER_21_876 ();
 sg13g2_decap_8 FILLER_22_0 ();
 sg13g2_decap_8 FILLER_22_11 ();
 sg13g2_decap_8 FILLER_22_18 ();
 sg13g2_fill_2 FILLER_22_25 ();
 sg13g2_decap_4 FILLER_22_32 ();
 sg13g2_fill_1 FILLER_22_36 ();
 sg13g2_decap_8 FILLER_22_53 ();
 sg13g2_decap_8 FILLER_22_60 ();
 sg13g2_fill_1 FILLER_22_67 ();
 sg13g2_decap_4 FILLER_22_72 ();
 sg13g2_fill_1 FILLER_22_76 ();
 sg13g2_fill_2 FILLER_22_88 ();
 sg13g2_decap_8 FILLER_22_94 ();
 sg13g2_fill_2 FILLER_22_101 ();
 sg13g2_decap_8 FILLER_22_108 ();
 sg13g2_decap_4 FILLER_22_115 ();
 sg13g2_fill_2 FILLER_22_124 ();
 sg13g2_decap_4 FILLER_22_131 ();
 sg13g2_decap_8 FILLER_22_140 ();
 sg13g2_decap_8 FILLER_22_147 ();
 sg13g2_decap_8 FILLER_22_154 ();
 sg13g2_decap_4 FILLER_22_161 ();
 sg13g2_fill_1 FILLER_22_165 ();
 sg13g2_decap_4 FILLER_22_173 ();
 sg13g2_decap_4 FILLER_22_181 ();
 sg13g2_fill_1 FILLER_22_185 ();
 sg13g2_fill_2 FILLER_22_198 ();
 sg13g2_fill_2 FILLER_22_234 ();
 sg13g2_fill_2 FILLER_22_239 ();
 sg13g2_fill_1 FILLER_22_241 ();
 sg13g2_fill_1 FILLER_22_246 ();
 sg13g2_fill_1 FILLER_22_252 ();
 sg13g2_decap_8 FILLER_22_260 ();
 sg13g2_decap_4 FILLER_22_267 ();
 sg13g2_fill_1 FILLER_22_271 ();
 sg13g2_decap_4 FILLER_22_276 ();
 sg13g2_fill_1 FILLER_22_280 ();
 sg13g2_decap_8 FILLER_22_286 ();
 sg13g2_fill_2 FILLER_22_293 ();
 sg13g2_decap_8 FILLER_22_299 ();
 sg13g2_fill_1 FILLER_22_306 ();
 sg13g2_decap_8 FILLER_22_311 ();
 sg13g2_decap_8 FILLER_22_318 ();
 sg13g2_fill_1 FILLER_22_325 ();
 sg13g2_fill_2 FILLER_22_356 ();
 sg13g2_decap_4 FILLER_22_362 ();
 sg13g2_fill_1 FILLER_22_366 ();
 sg13g2_decap_8 FILLER_22_371 ();
 sg13g2_fill_2 FILLER_22_378 ();
 sg13g2_fill_1 FILLER_22_380 ();
 sg13g2_fill_2 FILLER_22_391 ();
 sg13g2_fill_1 FILLER_22_393 ();
 sg13g2_fill_1 FILLER_22_398 ();
 sg13g2_decap_8 FILLER_22_403 ();
 sg13g2_fill_1 FILLER_22_410 ();
 sg13g2_decap_8 FILLER_22_415 ();
 sg13g2_decap_8 FILLER_22_422 ();
 sg13g2_decap_4 FILLER_22_437 ();
 sg13g2_fill_1 FILLER_22_441 ();
 sg13g2_decap_4 FILLER_22_450 ();
 sg13g2_decap_8 FILLER_22_466 ();
 sg13g2_fill_1 FILLER_22_473 ();
 sg13g2_fill_2 FILLER_22_484 ();
 sg13g2_fill_1 FILLER_22_486 ();
 sg13g2_decap_8 FILLER_22_516 ();
 sg13g2_decap_8 FILLER_22_523 ();
 sg13g2_fill_2 FILLER_22_530 ();
 sg13g2_fill_1 FILLER_22_532 ();
 sg13g2_fill_1 FILLER_22_548 ();
 sg13g2_decap_4 FILLER_22_562 ();
 sg13g2_decap_4 FILLER_22_571 ();
 sg13g2_fill_2 FILLER_22_575 ();
 sg13g2_decap_4 FILLER_22_582 ();
 sg13g2_fill_2 FILLER_22_586 ();
 sg13g2_fill_2 FILLER_22_606 ();
 sg13g2_decap_4 FILLER_22_618 ();
 sg13g2_decap_4 FILLER_22_637 ();
 sg13g2_fill_1 FILLER_22_641 ();
 sg13g2_fill_2 FILLER_22_665 ();
 sg13g2_fill_1 FILLER_22_667 ();
 sg13g2_decap_8 FILLER_22_675 ();
 sg13g2_decap_8 FILLER_22_682 ();
 sg13g2_decap_8 FILLER_22_704 ();
 sg13g2_decap_8 FILLER_22_711 ();
 sg13g2_decap_8 FILLER_22_718 ();
 sg13g2_decap_8 FILLER_22_725 ();
 sg13g2_fill_2 FILLER_22_732 ();
 sg13g2_fill_1 FILLER_22_734 ();
 sg13g2_decap_8 FILLER_22_745 ();
 sg13g2_decap_4 FILLER_22_752 ();
 sg13g2_fill_1 FILLER_22_756 ();
 sg13g2_decap_8 FILLER_22_771 ();
 sg13g2_decap_8 FILLER_22_782 ();
 sg13g2_decap_8 FILLER_22_789 ();
 sg13g2_decap_8 FILLER_22_796 ();
 sg13g2_decap_8 FILLER_22_803 ();
 sg13g2_decap_8 FILLER_22_810 ();
 sg13g2_decap_8 FILLER_22_817 ();
 sg13g2_decap_8 FILLER_22_824 ();
 sg13g2_decap_8 FILLER_22_831 ();
 sg13g2_decap_8 FILLER_22_838 ();
 sg13g2_decap_8 FILLER_22_845 ();
 sg13g2_decap_8 FILLER_22_852 ();
 sg13g2_decap_8 FILLER_22_859 ();
 sg13g2_decap_8 FILLER_22_866 ();
 sg13g2_decap_4 FILLER_22_873 ();
 sg13g2_fill_1 FILLER_22_877 ();
 sg13g2_decap_8 FILLER_23_0 ();
 sg13g2_fill_1 FILLER_23_7 ();
 sg13g2_decap_4 FILLER_23_12 ();
 sg13g2_fill_2 FILLER_23_20 ();
 sg13g2_decap_4 FILLER_23_30 ();
 sg13g2_fill_2 FILLER_23_34 ();
 sg13g2_decap_4 FILLER_23_52 ();
 sg13g2_fill_1 FILLER_23_56 ();
 sg13g2_fill_2 FILLER_23_74 ();
 sg13g2_decap_4 FILLER_23_88 ();
 sg13g2_fill_1 FILLER_23_92 ();
 sg13g2_decap_4 FILLER_23_98 ();
 sg13g2_decap_4 FILLER_23_111 ();
 sg13g2_fill_2 FILLER_23_115 ();
 sg13g2_decap_8 FILLER_23_134 ();
 sg13g2_decap_4 FILLER_23_141 ();
 sg13g2_decap_8 FILLER_23_154 ();
 sg13g2_fill_1 FILLER_23_161 ();
 sg13g2_fill_2 FILLER_23_197 ();
 sg13g2_fill_2 FILLER_23_204 ();
 sg13g2_fill_1 FILLER_23_206 ();
 sg13g2_fill_2 FILLER_23_211 ();
 sg13g2_decap_8 FILLER_23_218 ();
 sg13g2_decap_8 FILLER_23_225 ();
 sg13g2_decap_4 FILLER_23_236 ();
 sg13g2_fill_1 FILLER_23_264 ();
 sg13g2_decap_4 FILLER_23_291 ();
 sg13g2_fill_2 FILLER_23_333 ();
 sg13g2_fill_1 FILLER_23_335 ();
 sg13g2_decap_8 FILLER_23_341 ();
 sg13g2_fill_2 FILLER_23_348 ();
 sg13g2_fill_1 FILLER_23_350 ();
 sg13g2_fill_1 FILLER_23_360 ();
 sg13g2_fill_2 FILLER_23_390 ();
 sg13g2_fill_1 FILLER_23_392 ();
 sg13g2_fill_1 FILLER_23_398 ();
 sg13g2_decap_8 FILLER_23_433 ();
 sg13g2_fill_2 FILLER_23_440 ();
 sg13g2_decap_8 FILLER_23_459 ();
 sg13g2_decap_4 FILLER_23_466 ();
 sg13g2_fill_1 FILLER_23_470 ();
 sg13g2_decap_8 FILLER_23_479 ();
 sg13g2_decap_8 FILLER_23_486 ();
 sg13g2_fill_1 FILLER_23_493 ();
 sg13g2_fill_1 FILLER_23_498 ();
 sg13g2_fill_1 FILLER_23_503 ();
 sg13g2_fill_2 FILLER_23_514 ();
 sg13g2_fill_2 FILLER_23_526 ();
 sg13g2_fill_1 FILLER_23_528 ();
 sg13g2_decap_4 FILLER_23_543 ();
 sg13g2_decap_8 FILLER_23_551 ();
 sg13g2_decap_8 FILLER_23_558 ();
 sg13g2_decap_8 FILLER_23_565 ();
 sg13g2_decap_8 FILLER_23_572 ();
 sg13g2_fill_1 FILLER_23_584 ();
 sg13g2_fill_1 FILLER_23_590 ();
 sg13g2_fill_1 FILLER_23_596 ();
 sg13g2_fill_1 FILLER_23_602 ();
 sg13g2_decap_8 FILLER_23_613 ();
 sg13g2_fill_1 FILLER_23_620 ();
 sg13g2_decap_8 FILLER_23_633 ();
 sg13g2_decap_4 FILLER_23_640 ();
 sg13g2_fill_2 FILLER_23_644 ();
 sg13g2_fill_1 FILLER_23_656 ();
 sg13g2_fill_1 FILLER_23_661 ();
 sg13g2_decap_8 FILLER_23_666 ();
 sg13g2_decap_8 FILLER_23_673 ();
 sg13g2_fill_2 FILLER_23_680 ();
 sg13g2_decap_8 FILLER_23_687 ();
 sg13g2_fill_1 FILLER_23_698 ();
 sg13g2_decap_8 FILLER_23_713 ();
 sg13g2_fill_1 FILLER_23_720 ();
 sg13g2_decap_8 FILLER_23_726 ();
 sg13g2_fill_2 FILLER_23_733 ();
 sg13g2_decap_8 FILLER_23_744 ();
 sg13g2_decap_8 FILLER_23_751 ();
 sg13g2_decap_4 FILLER_23_758 ();
 sg13g2_fill_2 FILLER_23_762 ();
 sg13g2_decap_8 FILLER_23_775 ();
 sg13g2_fill_1 FILLER_23_782 ();
 sg13g2_decap_8 FILLER_23_819 ();
 sg13g2_decap_8 FILLER_23_826 ();
 sg13g2_decap_8 FILLER_23_833 ();
 sg13g2_decap_8 FILLER_23_840 ();
 sg13g2_decap_8 FILLER_23_847 ();
 sg13g2_decap_8 FILLER_23_854 ();
 sg13g2_decap_8 FILLER_23_861 ();
 sg13g2_decap_8 FILLER_23_868 ();
 sg13g2_fill_2 FILLER_23_875 ();
 sg13g2_fill_1 FILLER_23_877 ();
 sg13g2_fill_1 FILLER_24_0 ();
 sg13g2_decap_8 FILLER_24_27 ();
 sg13g2_decap_8 FILLER_24_34 ();
 sg13g2_decap_8 FILLER_24_41 ();
 sg13g2_decap_8 FILLER_24_48 ();
 sg13g2_decap_8 FILLER_24_55 ();
 sg13g2_fill_2 FILLER_24_62 ();
 sg13g2_fill_1 FILLER_24_64 ();
 sg13g2_decap_4 FILLER_24_74 ();
 sg13g2_fill_2 FILLER_24_82 ();
 sg13g2_fill_1 FILLER_24_100 ();
 sg13g2_fill_1 FILLER_24_106 ();
 sg13g2_decap_4 FILLER_24_138 ();
 sg13g2_fill_1 FILLER_24_142 ();
 sg13g2_fill_1 FILLER_24_160 ();
 sg13g2_decap_8 FILLER_24_165 ();
 sg13g2_fill_2 FILLER_24_172 ();
 sg13g2_fill_1 FILLER_24_174 ();
 sg13g2_fill_2 FILLER_24_180 ();
 sg13g2_fill_1 FILLER_24_182 ();
 sg13g2_fill_1 FILLER_24_187 ();
 sg13g2_fill_2 FILLER_24_203 ();
 sg13g2_fill_2 FILLER_24_209 ();
 sg13g2_fill_1 FILLER_24_211 ();
 sg13g2_decap_8 FILLER_24_246 ();
 sg13g2_decap_8 FILLER_24_253 ();
 sg13g2_decap_4 FILLER_24_260 ();
 sg13g2_fill_1 FILLER_24_264 ();
 sg13g2_decap_8 FILLER_24_269 ();
 sg13g2_fill_2 FILLER_24_276 ();
 sg13g2_decap_8 FILLER_24_281 ();
 sg13g2_fill_1 FILLER_24_288 ();
 sg13g2_decap_8 FILLER_24_298 ();
 sg13g2_fill_1 FILLER_24_305 ();
 sg13g2_decap_8 FILLER_24_317 ();
 sg13g2_decap_8 FILLER_24_324 ();
 sg13g2_fill_1 FILLER_24_341 ();
 sg13g2_decap_8 FILLER_24_346 ();
 sg13g2_fill_2 FILLER_24_353 ();
 sg13g2_fill_1 FILLER_24_355 ();
 sg13g2_decap_8 FILLER_24_377 ();
 sg13g2_fill_2 FILLER_24_390 ();
 sg13g2_decap_8 FILLER_24_402 ();
 sg13g2_decap_8 FILLER_24_409 ();
 sg13g2_decap_8 FILLER_24_416 ();
 sg13g2_decap_8 FILLER_24_423 ();
 sg13g2_fill_1 FILLER_24_430 ();
 sg13g2_decap_8 FILLER_24_457 ();
 sg13g2_decap_8 FILLER_24_464 ();
 sg13g2_decap_8 FILLER_24_471 ();
 sg13g2_fill_2 FILLER_24_478 ();
 sg13g2_decap_8 FILLER_24_514 ();
 sg13g2_fill_2 FILLER_24_521 ();
 sg13g2_fill_1 FILLER_24_523 ();
 sg13g2_fill_1 FILLER_24_538 ();
 sg13g2_decap_8 FILLER_24_549 ();
 sg13g2_decap_8 FILLER_24_556 ();
 sg13g2_decap_8 FILLER_24_563 ();
 sg13g2_decap_8 FILLER_24_583 ();
 sg13g2_fill_1 FILLER_24_590 ();
 sg13g2_fill_2 FILLER_24_610 ();
 sg13g2_decap_4 FILLER_24_617 ();
 sg13g2_fill_2 FILLER_24_621 ();
 sg13g2_fill_2 FILLER_24_636 ();
 sg13g2_fill_1 FILLER_24_638 ();
 sg13g2_fill_2 FILLER_24_644 ();
 sg13g2_fill_1 FILLER_24_661 ();
 sg13g2_decap_8 FILLER_24_674 ();
 sg13g2_decap_4 FILLER_24_681 ();
 sg13g2_fill_2 FILLER_24_685 ();
 sg13g2_decap_8 FILLER_24_691 ();
 sg13g2_fill_2 FILLER_24_698 ();
 sg13g2_fill_1 FILLER_24_700 ();
 sg13g2_decap_4 FILLER_24_705 ();
 sg13g2_decap_4 FILLER_24_712 ();
 sg13g2_decap_8 FILLER_24_730 ();
 sg13g2_fill_1 FILLER_24_737 ();
 sg13g2_decap_8 FILLER_24_742 ();
 sg13g2_fill_1 FILLER_24_749 ();
 sg13g2_fill_2 FILLER_24_754 ();
 sg13g2_decap_4 FILLER_24_778 ();
 sg13g2_fill_1 FILLER_24_782 ();
 sg13g2_decap_8 FILLER_24_793 ();
 sg13g2_decap_8 FILLER_24_804 ();
 sg13g2_fill_2 FILLER_24_811 ();
 sg13g2_decap_8 FILLER_24_817 ();
 sg13g2_decap_8 FILLER_24_824 ();
 sg13g2_decap_8 FILLER_24_831 ();
 sg13g2_decap_8 FILLER_24_838 ();
 sg13g2_decap_8 FILLER_24_845 ();
 sg13g2_decap_8 FILLER_24_852 ();
 sg13g2_decap_8 FILLER_24_859 ();
 sg13g2_decap_8 FILLER_24_866 ();
 sg13g2_decap_4 FILLER_24_873 ();
 sg13g2_fill_1 FILLER_24_877 ();
 sg13g2_decap_8 FILLER_25_0 ();
 sg13g2_fill_2 FILLER_25_7 ();
 sg13g2_fill_1 FILLER_25_9 ();
 sg13g2_fill_2 FILLER_25_21 ();
 sg13g2_fill_1 FILLER_25_23 ();
 sg13g2_fill_1 FILLER_25_54 ();
 sg13g2_decap_8 FILLER_25_60 ();
 sg13g2_decap_8 FILLER_25_67 ();
 sg13g2_decap_8 FILLER_25_74 ();
 sg13g2_fill_2 FILLER_25_81 ();
 sg13g2_fill_1 FILLER_25_83 ();
 sg13g2_decap_4 FILLER_25_106 ();
 sg13g2_fill_2 FILLER_25_116 ();
 sg13g2_decap_8 FILLER_25_125 ();
 sg13g2_decap_4 FILLER_25_132 ();
 sg13g2_fill_2 FILLER_25_172 ();
 sg13g2_fill_1 FILLER_25_174 ();
 sg13g2_decap_4 FILLER_25_201 ();
 sg13g2_fill_2 FILLER_25_205 ();
 sg13g2_decap_8 FILLER_25_212 ();
 sg13g2_decap_4 FILLER_25_219 ();
 sg13g2_decap_8 FILLER_25_227 ();
 sg13g2_decap_8 FILLER_25_234 ();
 sg13g2_decap_8 FILLER_25_241 ();
 sg13g2_decap_8 FILLER_25_248 ();
 sg13g2_decap_4 FILLER_25_260 ();
 sg13g2_fill_2 FILLER_25_264 ();
 sg13g2_decap_4 FILLER_25_270 ();
 sg13g2_fill_1 FILLER_25_274 ();
 sg13g2_decap_4 FILLER_25_279 ();
 sg13g2_fill_1 FILLER_25_283 ();
 sg13g2_fill_1 FILLER_25_288 ();
 sg13g2_fill_2 FILLER_25_292 ();
 sg13g2_fill_2 FILLER_25_304 ();
 sg13g2_fill_2 FILLER_25_332 ();
 sg13g2_fill_1 FILLER_25_334 ();
 sg13g2_decap_4 FILLER_25_361 ();
 sg13g2_decap_4 FILLER_25_398 ();
 sg13g2_decap_8 FILLER_25_407 ();
 sg13g2_decap_8 FILLER_25_414 ();
 sg13g2_decap_8 FILLER_25_421 ();
 sg13g2_fill_2 FILLER_25_433 ();
 sg13g2_fill_1 FILLER_25_443 ();
 sg13g2_fill_1 FILLER_25_449 ();
 sg13g2_decap_4 FILLER_25_454 ();
 sg13g2_fill_2 FILLER_25_458 ();
 sg13g2_decap_4 FILLER_25_465 ();
 sg13g2_fill_2 FILLER_25_469 ();
 sg13g2_decap_8 FILLER_25_475 ();
 sg13g2_decap_8 FILLER_25_482 ();
 sg13g2_decap_8 FILLER_25_489 ();
 sg13g2_decap_8 FILLER_25_496 ();
 sg13g2_decap_8 FILLER_25_513 ();
 sg13g2_decap_8 FILLER_25_520 ();
 sg13g2_fill_2 FILLER_25_552 ();
 sg13g2_decap_8 FILLER_25_580 ();
 sg13g2_decap_8 FILLER_25_587 ();
 sg13g2_decap_8 FILLER_25_594 ();
 sg13g2_decap_4 FILLER_25_601 ();
 sg13g2_fill_1 FILLER_25_605 ();
 sg13g2_decap_8 FILLER_25_611 ();
 sg13g2_fill_1 FILLER_25_618 ();
 sg13g2_fill_1 FILLER_25_623 ();
 sg13g2_fill_1 FILLER_25_634 ();
 sg13g2_fill_2 FILLER_25_644 ();
 sg13g2_fill_1 FILLER_25_646 ();
 sg13g2_fill_1 FILLER_25_652 ();
 sg13g2_decap_8 FILLER_25_662 ();
 sg13g2_decap_8 FILLER_25_669 ();
 sg13g2_decap_8 FILLER_25_676 ();
 sg13g2_decap_8 FILLER_25_683 ();
 sg13g2_decap_8 FILLER_25_690 ();
 sg13g2_decap_8 FILLER_25_697 ();
 sg13g2_fill_2 FILLER_25_704 ();
 sg13g2_fill_1 FILLER_25_706 ();
 sg13g2_decap_8 FILLER_25_711 ();
 sg13g2_decap_4 FILLER_25_718 ();
 sg13g2_fill_1 FILLER_25_722 ();
 sg13g2_decap_4 FILLER_25_727 ();
 sg13g2_fill_2 FILLER_25_731 ();
 sg13g2_fill_1 FILLER_25_751 ();
 sg13g2_fill_1 FILLER_25_762 ();
 sg13g2_fill_2 FILLER_25_767 ();
 sg13g2_decap_8 FILLER_25_799 ();
 sg13g2_decap_8 FILLER_25_832 ();
 sg13g2_decap_8 FILLER_25_839 ();
 sg13g2_decap_8 FILLER_25_846 ();
 sg13g2_decap_8 FILLER_25_853 ();
 sg13g2_decap_8 FILLER_25_860 ();
 sg13g2_decap_8 FILLER_25_867 ();
 sg13g2_decap_4 FILLER_25_874 ();
 sg13g2_fill_1 FILLER_26_0 ();
 sg13g2_decap_4 FILLER_26_27 ();
 sg13g2_fill_1 FILLER_26_31 ();
 sg13g2_decap_8 FILLER_26_36 ();
 sg13g2_fill_1 FILLER_26_43 ();
 sg13g2_fill_1 FILLER_26_52 ();
 sg13g2_decap_8 FILLER_26_58 ();
 sg13g2_decap_4 FILLER_26_65 ();
 sg13g2_fill_1 FILLER_26_78 ();
 sg13g2_fill_2 FILLER_26_95 ();
 sg13g2_fill_1 FILLER_26_101 ();
 sg13g2_decap_8 FILLER_26_107 ();
 sg13g2_fill_1 FILLER_26_114 ();
 sg13g2_fill_2 FILLER_26_119 ();
 sg13g2_decap_8 FILLER_26_125 ();
 sg13g2_decap_8 FILLER_26_132 ();
 sg13g2_fill_2 FILLER_26_139 ();
 sg13g2_fill_1 FILLER_26_141 ();
 sg13g2_fill_1 FILLER_26_152 ();
 sg13g2_decap_8 FILLER_26_157 ();
 sg13g2_decap_8 FILLER_26_164 ();
 sg13g2_decap_8 FILLER_26_171 ();
 sg13g2_fill_2 FILLER_26_178 ();
 sg13g2_fill_1 FILLER_26_180 ();
 sg13g2_decap_4 FILLER_26_185 ();
 sg13g2_fill_1 FILLER_26_189 ();
 sg13g2_decap_8 FILLER_26_195 ();
 sg13g2_fill_2 FILLER_26_202 ();
 sg13g2_fill_1 FILLER_26_208 ();
 sg13g2_decap_8 FILLER_26_221 ();
 sg13g2_decap_8 FILLER_26_228 ();
 sg13g2_decap_8 FILLER_26_235 ();
 sg13g2_decap_4 FILLER_26_242 ();
 sg13g2_fill_1 FILLER_26_246 ();
 sg13g2_fill_2 FILLER_26_256 ();
 sg13g2_fill_1 FILLER_26_258 ();
 sg13g2_decap_8 FILLER_26_293 ();
 sg13g2_fill_2 FILLER_26_300 ();
 sg13g2_decap_8 FILLER_26_316 ();
 sg13g2_decap_4 FILLER_26_323 ();
 sg13g2_decap_8 FILLER_26_341 ();
 sg13g2_fill_2 FILLER_26_348 ();
 sg13g2_decap_8 FILLER_26_355 ();
 sg13g2_fill_2 FILLER_26_362 ();
 sg13g2_fill_1 FILLER_26_364 ();
 sg13g2_fill_2 FILLER_26_370 ();
 sg13g2_fill_1 FILLER_26_379 ();
 sg13g2_fill_2 FILLER_26_384 ();
 sg13g2_decap_4 FILLER_26_391 ();
 sg13g2_fill_1 FILLER_26_395 ();
 sg13g2_decap_8 FILLER_26_401 ();
 sg13g2_decap_8 FILLER_26_408 ();
 sg13g2_fill_1 FILLER_26_415 ();
 sg13g2_decap_8 FILLER_26_421 ();
 sg13g2_fill_2 FILLER_26_428 ();
 sg13g2_decap_8 FILLER_26_434 ();
 sg13g2_fill_1 FILLER_26_441 ();
 sg13g2_fill_2 FILLER_26_458 ();
 sg13g2_fill_1 FILLER_26_460 ();
 sg13g2_fill_1 FILLER_26_466 ();
 sg13g2_fill_1 FILLER_26_472 ();
 sg13g2_fill_1 FILLER_26_478 ();
 sg13g2_decap_4 FILLER_26_519 ();
 sg13g2_decap_4 FILLER_26_567 ();
 sg13g2_decap_8 FILLER_26_622 ();
 sg13g2_fill_1 FILLER_26_629 ();
 sg13g2_fill_2 FILLER_26_635 ();
 sg13g2_fill_2 FILLER_26_670 ();
 sg13g2_fill_2 FILLER_26_713 ();
 sg13g2_decap_8 FILLER_26_745 ();
 sg13g2_decap_4 FILLER_26_752 ();
 sg13g2_decap_8 FILLER_26_807 ();
 sg13g2_decap_8 FILLER_26_814 ();
 sg13g2_decap_8 FILLER_26_821 ();
 sg13g2_decap_8 FILLER_26_828 ();
 sg13g2_decap_8 FILLER_26_835 ();
 sg13g2_decap_8 FILLER_26_842 ();
 sg13g2_decap_8 FILLER_26_849 ();
 sg13g2_decap_8 FILLER_26_856 ();
 sg13g2_decap_8 FILLER_26_863 ();
 sg13g2_decap_8 FILLER_26_870 ();
 sg13g2_fill_1 FILLER_26_877 ();
 sg13g2_decap_8 FILLER_27_0 ();
 sg13g2_fill_1 FILLER_27_7 ();
 sg13g2_decap_8 FILLER_27_24 ();
 sg13g2_decap_8 FILLER_27_31 ();
 sg13g2_fill_1 FILLER_27_38 ();
 sg13g2_decap_8 FILLER_27_48 ();
 sg13g2_decap_4 FILLER_27_55 ();
 sg13g2_decap_8 FILLER_27_69 ();
 sg13g2_decap_4 FILLER_27_76 ();
 sg13g2_fill_1 FILLER_27_80 ();
 sg13g2_fill_1 FILLER_27_91 ();
 sg13g2_fill_1 FILLER_27_100 ();
 sg13g2_fill_2 FILLER_27_105 ();
 sg13g2_fill_1 FILLER_27_111 ();
 sg13g2_fill_2 FILLER_27_122 ();
 sg13g2_decap_4 FILLER_27_128 ();
 sg13g2_decap_4 FILLER_27_140 ();
 sg13g2_decap_4 FILLER_27_148 ();
 sg13g2_decap_4 FILLER_27_178 ();
 sg13g2_fill_1 FILLER_27_182 ();
 sg13g2_decap_8 FILLER_27_196 ();
 sg13g2_decap_8 FILLER_27_233 ();
 sg13g2_fill_2 FILLER_27_240 ();
 sg13g2_fill_1 FILLER_27_242 ();
 sg13g2_fill_2 FILLER_27_248 ();
 sg13g2_fill_1 FILLER_27_250 ();
 sg13g2_decap_8 FILLER_27_255 ();
 sg13g2_decap_8 FILLER_27_262 ();
 sg13g2_decap_8 FILLER_27_269 ();
 sg13g2_decap_4 FILLER_27_276 ();
 sg13g2_fill_1 FILLER_27_284 ();
 sg13g2_decap_4 FILLER_27_315 ();
 sg13g2_decap_8 FILLER_27_345 ();
 sg13g2_fill_1 FILLER_27_352 ();
 sg13g2_fill_2 FILLER_27_363 ();
 sg13g2_fill_1 FILLER_27_365 ();
 sg13g2_fill_1 FILLER_27_373 ();
 sg13g2_fill_1 FILLER_27_388 ();
 sg13g2_fill_1 FILLER_27_396 ();
 sg13g2_decap_4 FILLER_27_401 ();
 sg13g2_decap_8 FILLER_27_409 ();
 sg13g2_decap_8 FILLER_27_416 ();
 sg13g2_decap_8 FILLER_27_423 ();
 sg13g2_fill_1 FILLER_27_430 ();
 sg13g2_fill_2 FILLER_27_436 ();
 sg13g2_fill_1 FILLER_27_443 ();
 sg13g2_decap_8 FILLER_27_467 ();
 sg13g2_decap_4 FILLER_27_474 ();
 sg13g2_decap_4 FILLER_27_482 ();
 sg13g2_decap_8 FILLER_27_494 ();
 sg13g2_decap_8 FILLER_27_501 ();
 sg13g2_decap_4 FILLER_27_508 ();
 sg13g2_fill_2 FILLER_27_512 ();
 sg13g2_decap_8 FILLER_27_523 ();
 sg13g2_decap_8 FILLER_27_535 ();
 sg13g2_decap_8 FILLER_27_542 ();
 sg13g2_decap_4 FILLER_27_549 ();
 sg13g2_fill_1 FILLER_27_553 ();
 sg13g2_decap_4 FILLER_27_571 ();
 sg13g2_decap_8 FILLER_27_579 ();
 sg13g2_decap_4 FILLER_27_586 ();
 sg13g2_decap_8 FILLER_27_594 ();
 sg13g2_decap_8 FILLER_27_601 ();
 sg13g2_decap_8 FILLER_27_608 ();
 sg13g2_decap_4 FILLER_27_615 ();
 sg13g2_fill_1 FILLER_27_619 ();
 sg13g2_decap_4 FILLER_27_630 ();
 sg13g2_fill_1 FILLER_27_634 ();
 sg13g2_fill_1 FILLER_27_646 ();
 sg13g2_decap_8 FILLER_27_651 ();
 sg13g2_fill_1 FILLER_27_658 ();
 sg13g2_decap_8 FILLER_27_662 ();
 sg13g2_fill_2 FILLER_27_669 ();
 sg13g2_decap_8 FILLER_27_677 ();
 sg13g2_decap_8 FILLER_27_684 ();
 sg13g2_fill_1 FILLER_27_691 ();
 sg13g2_decap_8 FILLER_27_696 ();
 sg13g2_decap_8 FILLER_27_703 ();
 sg13g2_decap_8 FILLER_27_710 ();
 sg13g2_decap_8 FILLER_27_726 ();
 sg13g2_decap_4 FILLER_27_733 ();
 sg13g2_fill_1 FILLER_27_737 ();
 sg13g2_fill_1 FILLER_27_747 ();
 sg13g2_decap_4 FILLER_27_774 ();
 sg13g2_decap_8 FILLER_27_789 ();
 sg13g2_decap_8 FILLER_27_796 ();
 sg13g2_decap_8 FILLER_27_803 ();
 sg13g2_decap_8 FILLER_27_810 ();
 sg13g2_decap_8 FILLER_27_817 ();
 sg13g2_decap_8 FILLER_27_824 ();
 sg13g2_decap_8 FILLER_27_831 ();
 sg13g2_decap_8 FILLER_27_838 ();
 sg13g2_decap_8 FILLER_27_845 ();
 sg13g2_decap_8 FILLER_27_852 ();
 sg13g2_decap_8 FILLER_27_859 ();
 sg13g2_decap_8 FILLER_27_866 ();
 sg13g2_decap_4 FILLER_27_873 ();
 sg13g2_fill_1 FILLER_27_877 ();
 sg13g2_decap_8 FILLER_28_0 ();
 sg13g2_fill_2 FILLER_28_7 ();
 sg13g2_fill_1 FILLER_28_9 ();
 sg13g2_decap_8 FILLER_28_37 ();
 sg13g2_decap_8 FILLER_28_44 ();
 sg13g2_fill_1 FILLER_28_51 ();
 sg13g2_decap_8 FILLER_28_66 ();
 sg13g2_decap_4 FILLER_28_73 ();
 sg13g2_decap_4 FILLER_28_81 ();
 sg13g2_fill_1 FILLER_28_85 ();
 sg13g2_fill_1 FILLER_28_111 ();
 sg13g2_decap_8 FILLER_28_162 ();
 sg13g2_decap_8 FILLER_28_169 ();
 sg13g2_decap_8 FILLER_28_206 ();
 sg13g2_fill_2 FILLER_28_213 ();
 sg13g2_fill_1 FILLER_28_215 ();
 sg13g2_decap_8 FILLER_28_231 ();
 sg13g2_decap_4 FILLER_28_238 ();
 sg13g2_fill_1 FILLER_28_242 ();
 sg13g2_decap_8 FILLER_28_269 ();
 sg13g2_decap_8 FILLER_28_276 ();
 sg13g2_decap_8 FILLER_28_283 ();
 sg13g2_decap_4 FILLER_28_290 ();
 sg13g2_fill_1 FILLER_28_294 ();
 sg13g2_decap_8 FILLER_28_299 ();
 sg13g2_decap_8 FILLER_28_306 ();
 sg13g2_decap_8 FILLER_28_313 ();
 sg13g2_decap_8 FILLER_28_320 ();
 sg13g2_fill_2 FILLER_28_327 ();
 sg13g2_decap_8 FILLER_28_333 ();
 sg13g2_decap_4 FILLER_28_340 ();
 sg13g2_fill_1 FILLER_28_344 ();
 sg13g2_fill_2 FILLER_28_349 ();
 sg13g2_fill_1 FILLER_28_351 ();
 sg13g2_decap_8 FILLER_28_373 ();
 sg13g2_fill_2 FILLER_28_384 ();
 sg13g2_fill_2 FILLER_28_393 ();
 sg13g2_decap_8 FILLER_28_405 ();
 sg13g2_decap_8 FILLER_28_412 ();
 sg13g2_fill_1 FILLER_28_419 ();
 sg13g2_fill_1 FILLER_28_430 ();
 sg13g2_fill_2 FILLER_28_453 ();
 sg13g2_fill_1 FILLER_28_455 ();
 sg13g2_fill_2 FILLER_28_461 ();
 sg13g2_decap_4 FILLER_28_473 ();
 sg13g2_decap_8 FILLER_28_481 ();
 sg13g2_fill_2 FILLER_28_488 ();
 sg13g2_fill_1 FILLER_28_490 ();
 sg13g2_decap_4 FILLER_28_517 ();
 sg13g2_decap_4 FILLER_28_525 ();
 sg13g2_fill_2 FILLER_28_560 ();
 sg13g2_fill_1 FILLER_28_562 ();
 sg13g2_fill_2 FILLER_28_589 ();
 sg13g2_decap_8 FILLER_28_595 ();
 sg13g2_fill_2 FILLER_28_602 ();
 sg13g2_fill_1 FILLER_28_604 ();
 sg13g2_fill_1 FILLER_28_609 ();
 sg13g2_decap_8 FILLER_28_615 ();
 sg13g2_decap_4 FILLER_28_622 ();
 sg13g2_decap_4 FILLER_28_633 ();
 sg13g2_fill_2 FILLER_28_637 ();
 sg13g2_decap_8 FILLER_28_644 ();
 sg13g2_fill_2 FILLER_28_651 ();
 sg13g2_decap_4 FILLER_28_683 ();
 sg13g2_decap_8 FILLER_28_691 ();
 sg13g2_decap_8 FILLER_28_698 ();
 sg13g2_decap_8 FILLER_28_705 ();
 sg13g2_fill_1 FILLER_28_717 ();
 sg13g2_decap_8 FILLER_28_726 ();
 sg13g2_fill_2 FILLER_28_733 ();
 sg13g2_decap_4 FILLER_28_744 ();
 sg13g2_fill_1 FILLER_28_748 ();
 sg13g2_fill_1 FILLER_28_754 ();
 sg13g2_decap_8 FILLER_28_763 ();
 sg13g2_decap_8 FILLER_28_770 ();
 sg13g2_fill_2 FILLER_28_777 ();
 sg13g2_fill_1 FILLER_28_779 ();
 sg13g2_decap_8 FILLER_28_788 ();
 sg13g2_fill_2 FILLER_28_795 ();
 sg13g2_fill_1 FILLER_28_797 ();
 sg13g2_decap_8 FILLER_28_802 ();
 sg13g2_decap_8 FILLER_28_809 ();
 sg13g2_decap_8 FILLER_28_816 ();
 sg13g2_decap_8 FILLER_28_823 ();
 sg13g2_decap_8 FILLER_28_830 ();
 sg13g2_decap_8 FILLER_28_837 ();
 sg13g2_decap_8 FILLER_28_844 ();
 sg13g2_decap_8 FILLER_28_851 ();
 sg13g2_decap_8 FILLER_28_858 ();
 sg13g2_decap_8 FILLER_28_865 ();
 sg13g2_decap_4 FILLER_28_872 ();
 sg13g2_fill_2 FILLER_28_876 ();
 sg13g2_decap_8 FILLER_29_0 ();
 sg13g2_fill_2 FILLER_29_7 ();
 sg13g2_fill_2 FILLER_29_13 ();
 sg13g2_fill_1 FILLER_29_15 ();
 sg13g2_fill_2 FILLER_29_20 ();
 sg13g2_fill_1 FILLER_29_27 ();
 sg13g2_decap_8 FILLER_29_33 ();
 sg13g2_fill_2 FILLER_29_40 ();
 sg13g2_decap_8 FILLER_29_68 ();
 sg13g2_decap_4 FILLER_29_75 ();
 sg13g2_fill_1 FILLER_29_79 ();
 sg13g2_decap_8 FILLER_29_89 ();
 sg13g2_decap_4 FILLER_29_96 ();
 sg13g2_fill_2 FILLER_29_105 ();
 sg13g2_fill_2 FILLER_29_111 ();
 sg13g2_fill_1 FILLER_29_113 ();
 sg13g2_decap_4 FILLER_29_123 ();
 sg13g2_decap_8 FILLER_29_130 ();
 sg13g2_decap_8 FILLER_29_137 ();
 sg13g2_decap_4 FILLER_29_144 ();
 sg13g2_fill_2 FILLER_29_148 ();
 sg13g2_decap_8 FILLER_29_154 ();
 sg13g2_decap_8 FILLER_29_161 ();
 sg13g2_decap_8 FILLER_29_168 ();
 sg13g2_fill_2 FILLER_29_175 ();
 sg13g2_fill_1 FILLER_29_177 ();
 sg13g2_decap_4 FILLER_29_183 ();
 sg13g2_fill_2 FILLER_29_196 ();
 sg13g2_fill_1 FILLER_29_198 ();
 sg13g2_decap_8 FILLER_29_209 ();
 sg13g2_fill_1 FILLER_29_216 ();
 sg13g2_fill_2 FILLER_29_237 ();
 sg13g2_fill_1 FILLER_29_247 ();
 sg13g2_decap_8 FILLER_29_251 ();
 sg13g2_fill_2 FILLER_29_258 ();
 sg13g2_fill_1 FILLER_29_260 ();
 sg13g2_fill_1 FILLER_29_270 ();
 sg13g2_decap_4 FILLER_29_276 ();
 sg13g2_decap_8 FILLER_29_284 ();
 sg13g2_decap_8 FILLER_29_291 ();
 sg13g2_fill_2 FILLER_29_307 ();
 sg13g2_fill_2 FILLER_29_317 ();
 sg13g2_fill_1 FILLER_29_319 ();
 sg13g2_decap_8 FILLER_29_346 ();
 sg13g2_fill_2 FILLER_29_353 ();
 sg13g2_fill_1 FILLER_29_355 ();
 sg13g2_fill_2 FILLER_29_364 ();
 sg13g2_fill_2 FILLER_29_389 ();
 sg13g2_fill_1 FILLER_29_391 ();
 sg13g2_decap_4 FILLER_29_397 ();
 sg13g2_fill_2 FILLER_29_401 ();
 sg13g2_fill_2 FILLER_29_407 ();
 sg13g2_fill_2 FILLER_29_417 ();
 sg13g2_fill_1 FILLER_29_419 ();
 sg13g2_decap_8 FILLER_29_463 ();
 sg13g2_decap_8 FILLER_29_470 ();
 sg13g2_decap_4 FILLER_29_477 ();
 sg13g2_fill_2 FILLER_29_481 ();
 sg13g2_decap_8 FILLER_29_488 ();
 sg13g2_fill_1 FILLER_29_495 ();
 sg13g2_fill_1 FILLER_29_500 ();
 sg13g2_decap_8 FILLER_29_505 ();
 sg13g2_decap_8 FILLER_29_512 ();
 sg13g2_decap_8 FILLER_29_519 ();
 sg13g2_decap_8 FILLER_29_526 ();
 sg13g2_fill_2 FILLER_29_533 ();
 sg13g2_decap_8 FILLER_29_539 ();
 sg13g2_fill_2 FILLER_29_546 ();
 sg13g2_fill_2 FILLER_29_561 ();
 sg13g2_fill_1 FILLER_29_563 ();
 sg13g2_fill_2 FILLER_29_573 ();
 sg13g2_fill_1 FILLER_29_575 ();
 sg13g2_fill_1 FILLER_29_585 ();
 sg13g2_fill_2 FILLER_29_596 ();
 sg13g2_fill_2 FILLER_29_624 ();
 sg13g2_fill_1 FILLER_29_626 ();
 sg13g2_decap_8 FILLER_29_632 ();
 sg13g2_decap_8 FILLER_29_639 ();
 sg13g2_decap_4 FILLER_29_646 ();
 sg13g2_decap_4 FILLER_29_653 ();
 sg13g2_fill_2 FILLER_29_657 ();
 sg13g2_fill_2 FILLER_29_672 ();
 sg13g2_fill_2 FILLER_29_679 ();
 sg13g2_fill_2 FILLER_29_707 ();
 sg13g2_fill_1 FILLER_29_709 ();
 sg13g2_fill_1 FILLER_29_736 ();
 sg13g2_fill_1 FILLER_29_763 ();
 sg13g2_fill_1 FILLER_29_773 ();
 sg13g2_decap_8 FILLER_29_778 ();
 sg13g2_decap_4 FILLER_29_785 ();
 sg13g2_fill_2 FILLER_29_789 ();
 sg13g2_decap_8 FILLER_29_817 ();
 sg13g2_decap_8 FILLER_29_824 ();
 sg13g2_decap_8 FILLER_29_831 ();
 sg13g2_decap_8 FILLER_29_838 ();
 sg13g2_decap_8 FILLER_29_845 ();
 sg13g2_decap_8 FILLER_29_852 ();
 sg13g2_decap_8 FILLER_29_859 ();
 sg13g2_decap_8 FILLER_29_866 ();
 sg13g2_decap_4 FILLER_29_873 ();
 sg13g2_fill_1 FILLER_29_877 ();
 sg13g2_decap_8 FILLER_30_0 ();
 sg13g2_decap_8 FILLER_30_28 ();
 sg13g2_decap_8 FILLER_30_35 ();
 sg13g2_fill_2 FILLER_30_42 ();
 sg13g2_decap_8 FILLER_30_54 ();
 sg13g2_decap_8 FILLER_30_61 ();
 sg13g2_decap_8 FILLER_30_68 ();
 sg13g2_decap_4 FILLER_30_75 ();
 sg13g2_decap_4 FILLER_30_84 ();
 sg13g2_fill_2 FILLER_30_88 ();
 sg13g2_fill_1 FILLER_30_110 ();
 sg13g2_fill_1 FILLER_30_120 ();
 sg13g2_fill_1 FILLER_30_130 ();
 sg13g2_decap_8 FILLER_30_157 ();
 sg13g2_decap_4 FILLER_30_164 ();
 sg13g2_fill_2 FILLER_30_168 ();
 sg13g2_decap_8 FILLER_30_174 ();
 sg13g2_fill_2 FILLER_30_181 ();
 sg13g2_fill_1 FILLER_30_183 ();
 sg13g2_fill_2 FILLER_30_197 ();
 sg13g2_decap_8 FILLER_30_210 ();
 sg13g2_decap_4 FILLER_30_217 ();
 sg13g2_decap_8 FILLER_30_224 ();
 sg13g2_fill_1 FILLER_30_231 ();
 sg13g2_decap_8 FILLER_30_244 ();
 sg13g2_decap_8 FILLER_30_251 ();
 sg13g2_decap_8 FILLER_30_258 ();
 sg13g2_fill_1 FILLER_30_265 ();
 sg13g2_fill_1 FILLER_30_307 ();
 sg13g2_fill_1 FILLER_30_317 ();
 sg13g2_fill_1 FILLER_30_322 ();
 sg13g2_decap_8 FILLER_30_327 ();
 sg13g2_decap_8 FILLER_30_334 ();
 sg13g2_decap_8 FILLER_30_341 ();
 sg13g2_decap_8 FILLER_30_348 ();
 sg13g2_decap_4 FILLER_30_355 ();
 sg13g2_decap_4 FILLER_30_370 ();
 sg13g2_fill_1 FILLER_30_374 ();
 sg13g2_decap_8 FILLER_30_385 ();
 sg13g2_decap_8 FILLER_30_392 ();
 sg13g2_decap_8 FILLER_30_399 ();
 sg13g2_decap_8 FILLER_30_406 ();
 sg13g2_fill_2 FILLER_30_413 ();
 sg13g2_fill_1 FILLER_30_415 ();
 sg13g2_decap_8 FILLER_30_424 ();
 sg13g2_fill_1 FILLER_30_431 ();
 sg13g2_decap_8 FILLER_30_454 ();
 sg13g2_fill_2 FILLER_30_478 ();
 sg13g2_fill_1 FILLER_30_480 ();
 sg13g2_decap_8 FILLER_30_516 ();
 sg13g2_decap_8 FILLER_30_523 ();
 sg13g2_decap_4 FILLER_30_530 ();
 sg13g2_fill_2 FILLER_30_534 ();
 sg13g2_decap_4 FILLER_30_540 ();
 sg13g2_fill_1 FILLER_30_544 ();
 sg13g2_decap_8 FILLER_30_613 ();
 sg13g2_decap_4 FILLER_30_620 ();
 sg13g2_fill_2 FILLER_30_628 ();
 sg13g2_fill_2 FILLER_30_656 ();
 sg13g2_fill_1 FILLER_30_658 ();
 sg13g2_decap_8 FILLER_30_672 ();
 sg13g2_decap_8 FILLER_30_679 ();
 sg13g2_decap_8 FILLER_30_686 ();
 sg13g2_decap_4 FILLER_30_693 ();
 sg13g2_decap_8 FILLER_30_705 ();
 sg13g2_decap_8 FILLER_30_712 ();
 sg13g2_fill_2 FILLER_30_719 ();
 sg13g2_fill_1 FILLER_30_721 ();
 sg13g2_decap_8 FILLER_30_727 ();
 sg13g2_fill_1 FILLER_30_734 ();
 sg13g2_fill_1 FILLER_30_752 ();
 sg13g2_decap_8 FILLER_30_757 ();
 sg13g2_fill_2 FILLER_30_764 ();
 sg13g2_fill_1 FILLER_30_766 ();
 sg13g2_decap_8 FILLER_30_793 ();
 sg13g2_decap_8 FILLER_30_800 ();
 sg13g2_decap_8 FILLER_30_807 ();
 sg13g2_decap_8 FILLER_30_814 ();
 sg13g2_decap_8 FILLER_30_821 ();
 sg13g2_decap_8 FILLER_30_828 ();
 sg13g2_decap_8 FILLER_30_835 ();
 sg13g2_decap_8 FILLER_30_842 ();
 sg13g2_decap_8 FILLER_30_849 ();
 sg13g2_decap_8 FILLER_30_856 ();
 sg13g2_decap_8 FILLER_30_863 ();
 sg13g2_decap_8 FILLER_30_870 ();
 sg13g2_fill_1 FILLER_30_877 ();
 sg13g2_fill_1 FILLER_31_0 ();
 sg13g2_fill_2 FILLER_31_27 ();
 sg13g2_fill_2 FILLER_31_50 ();
 sg13g2_fill_2 FILLER_31_62 ();
 sg13g2_fill_1 FILLER_31_85 ();
 sg13g2_decap_8 FILLER_31_101 ();
 sg13g2_decap_4 FILLER_31_108 ();
 sg13g2_fill_1 FILLER_31_117 ();
 sg13g2_fill_1 FILLER_31_123 ();
 sg13g2_fill_1 FILLER_31_128 ();
 sg13g2_decap_4 FILLER_31_134 ();
 sg13g2_decap_8 FILLER_31_142 ();
 sg13g2_decap_8 FILLER_31_149 ();
 sg13g2_decap_4 FILLER_31_156 ();
 sg13g2_fill_1 FILLER_31_160 ();
 sg13g2_decap_8 FILLER_31_187 ();
 sg13g2_fill_2 FILLER_31_199 ();
 sg13g2_decap_4 FILLER_31_211 ();
 sg13g2_decap_8 FILLER_31_252 ();
 sg13g2_decap_8 FILLER_31_259 ();
 sg13g2_decap_4 FILLER_31_266 ();
 sg13g2_fill_1 FILLER_31_270 ();
 sg13g2_fill_2 FILLER_31_309 ();
 sg13g2_fill_1 FILLER_31_311 ();
 sg13g2_decap_4 FILLER_31_338 ();
 sg13g2_fill_1 FILLER_31_342 ();
 sg13g2_decap_8 FILLER_31_348 ();
 sg13g2_fill_2 FILLER_31_355 ();
 sg13g2_fill_1 FILLER_31_357 ();
 sg13g2_fill_2 FILLER_31_363 ();
 sg13g2_fill_1 FILLER_31_365 ();
 sg13g2_fill_1 FILLER_31_372 ();
 sg13g2_decap_4 FILLER_31_384 ();
 sg13g2_fill_1 FILLER_31_388 ();
 sg13g2_decap_4 FILLER_31_397 ();
 sg13g2_decap_4 FILLER_31_409 ();
 sg13g2_fill_2 FILLER_31_413 ();
 sg13g2_decap_8 FILLER_31_420 ();
 sg13g2_decap_8 FILLER_31_427 ();
 sg13g2_decap_4 FILLER_31_434 ();
 sg13g2_fill_1 FILLER_31_438 ();
 sg13g2_fill_2 FILLER_31_443 ();
 sg13g2_fill_1 FILLER_31_445 ();
 sg13g2_decap_4 FILLER_31_454 ();
 sg13g2_fill_1 FILLER_31_458 ();
 sg13g2_decap_8 FILLER_31_463 ();
 sg13g2_decap_8 FILLER_31_470 ();
 sg13g2_fill_2 FILLER_31_477 ();
 sg13g2_fill_2 FILLER_31_488 ();
 sg13g2_fill_1 FILLER_31_490 ();
 sg13g2_fill_1 FILLER_31_495 ();
 sg13g2_decap_4 FILLER_31_502 ();
 sg13g2_fill_1 FILLER_31_506 ();
 sg13g2_fill_2 FILLER_31_512 ();
 sg13g2_fill_1 FILLER_31_514 ();
 sg13g2_decap_8 FILLER_31_555 ();
 sg13g2_decap_8 FILLER_31_562 ();
 sg13g2_fill_2 FILLER_31_574 ();
 sg13g2_fill_1 FILLER_31_576 ();
 sg13g2_decap_8 FILLER_31_607 ();
 sg13g2_decap_8 FILLER_31_614 ();
 sg13g2_decap_8 FILLER_31_621 ();
 sg13g2_decap_8 FILLER_31_628 ();
 sg13g2_decap_4 FILLER_31_635 ();
 sg13g2_decap_8 FILLER_31_643 ();
 sg13g2_decap_8 FILLER_31_650 ();
 sg13g2_fill_1 FILLER_31_721 ();
 sg13g2_decap_8 FILLER_31_748 ();
 sg13g2_fill_2 FILLER_31_755 ();
 sg13g2_decap_4 FILLER_31_762 ();
 sg13g2_fill_1 FILLER_31_766 ();
 sg13g2_decap_8 FILLER_31_771 ();
 sg13g2_decap_8 FILLER_31_778 ();
 sg13g2_decap_8 FILLER_31_785 ();
 sg13g2_decap_8 FILLER_31_792 ();
 sg13g2_decap_8 FILLER_31_799 ();
 sg13g2_decap_8 FILLER_31_806 ();
 sg13g2_decap_8 FILLER_31_813 ();
 sg13g2_decap_8 FILLER_31_820 ();
 sg13g2_decap_8 FILLER_31_827 ();
 sg13g2_decap_8 FILLER_31_834 ();
 sg13g2_decap_8 FILLER_31_841 ();
 sg13g2_decap_8 FILLER_31_848 ();
 sg13g2_decap_8 FILLER_31_855 ();
 sg13g2_decap_8 FILLER_31_862 ();
 sg13g2_decap_8 FILLER_31_869 ();
 sg13g2_fill_2 FILLER_31_876 ();
 sg13g2_decap_8 FILLER_32_0 ();
 sg13g2_decap_8 FILLER_32_11 ();
 sg13g2_fill_1 FILLER_32_18 ();
 sg13g2_decap_8 FILLER_32_23 ();
 sg13g2_fill_2 FILLER_32_30 ();
 sg13g2_fill_1 FILLER_32_32 ();
 sg13g2_decap_4 FILLER_32_75 ();
 sg13g2_fill_1 FILLER_32_79 ();
 sg13g2_decap_8 FILLER_32_101 ();
 sg13g2_fill_1 FILLER_32_108 ();
 sg13g2_fill_2 FILLER_32_129 ();
 sg13g2_decap_8 FILLER_32_148 ();
 sg13g2_fill_1 FILLER_32_155 ();
 sg13g2_decap_8 FILLER_32_161 ();
 sg13g2_decap_8 FILLER_32_168 ();
 sg13g2_decap_8 FILLER_32_175 ();
 sg13g2_decap_8 FILLER_32_182 ();
 sg13g2_decap_8 FILLER_32_189 ();
 sg13g2_fill_2 FILLER_32_196 ();
 sg13g2_decap_8 FILLER_32_214 ();
 sg13g2_decap_8 FILLER_32_225 ();
 sg13g2_decap_8 FILLER_32_232 ();
 sg13g2_decap_8 FILLER_32_249 ();
 sg13g2_fill_2 FILLER_32_256 ();
 sg13g2_fill_1 FILLER_32_258 ();
 sg13g2_fill_2 FILLER_32_328 ();
 sg13g2_fill_2 FILLER_32_346 ();
 sg13g2_decap_4 FILLER_32_351 ();
 sg13g2_fill_2 FILLER_32_355 ();
 sg13g2_fill_1 FILLER_32_367 ();
 sg13g2_fill_1 FILLER_32_385 ();
 sg13g2_fill_2 FILLER_32_398 ();
 sg13g2_fill_1 FILLER_32_400 ();
 sg13g2_fill_2 FILLER_32_415 ();
 sg13g2_decap_8 FILLER_32_425 ();
 sg13g2_decap_8 FILLER_32_432 ();
 sg13g2_decap_8 FILLER_32_439 ();
 sg13g2_decap_4 FILLER_32_446 ();
 sg13g2_fill_2 FILLER_32_458 ();
 sg13g2_fill_1 FILLER_32_460 ();
 sg13g2_fill_2 FILLER_32_495 ();
 sg13g2_fill_1 FILLER_32_497 ();
 sg13g2_decap_8 FILLER_32_508 ();
 sg13g2_decap_8 FILLER_32_515 ();
 sg13g2_fill_2 FILLER_32_522 ();
 sg13g2_fill_1 FILLER_32_524 ();
 sg13g2_decap_8 FILLER_32_530 ();
 sg13g2_decap_8 FILLER_32_537 ();
 sg13g2_decap_8 FILLER_32_544 ();
 sg13g2_decap_8 FILLER_32_551 ();
 sg13g2_decap_8 FILLER_32_558 ();
 sg13g2_decap_4 FILLER_32_565 ();
 sg13g2_decap_8 FILLER_32_575 ();
 sg13g2_fill_2 FILLER_32_582 ();
 sg13g2_fill_2 FILLER_32_594 ();
 sg13g2_decap_4 FILLER_32_600 ();
 sg13g2_decap_4 FILLER_32_640 ();
 sg13g2_fill_2 FILLER_32_644 ();
 sg13g2_decap_8 FILLER_32_652 ();
 sg13g2_fill_1 FILLER_32_659 ();
 sg13g2_fill_1 FILLER_32_663 ();
 sg13g2_decap_8 FILLER_32_682 ();
 sg13g2_fill_1 FILLER_32_689 ();
 sg13g2_decap_8 FILLER_32_694 ();
 sg13g2_decap_8 FILLER_32_705 ();
 sg13g2_decap_8 FILLER_32_712 ();
 sg13g2_decap_8 FILLER_32_719 ();
 sg13g2_fill_2 FILLER_32_726 ();
 sg13g2_fill_2 FILLER_32_732 ();
 sg13g2_fill_1 FILLER_32_734 ();
 sg13g2_decap_8 FILLER_32_744 ();
 sg13g2_decap_4 FILLER_32_751 ();
 sg13g2_fill_1 FILLER_32_755 ();
 sg13g2_decap_8 FILLER_32_786 ();
 sg13g2_decap_8 FILLER_32_793 ();
 sg13g2_decap_8 FILLER_32_800 ();
 sg13g2_decap_8 FILLER_32_807 ();
 sg13g2_decap_8 FILLER_32_814 ();
 sg13g2_decap_8 FILLER_32_821 ();
 sg13g2_decap_8 FILLER_32_828 ();
 sg13g2_decap_8 FILLER_32_835 ();
 sg13g2_decap_8 FILLER_32_842 ();
 sg13g2_decap_8 FILLER_32_849 ();
 sg13g2_decap_8 FILLER_32_856 ();
 sg13g2_decap_8 FILLER_32_863 ();
 sg13g2_decap_8 FILLER_32_870 ();
 sg13g2_fill_1 FILLER_32_877 ();
 sg13g2_decap_8 FILLER_33_0 ();
 sg13g2_fill_1 FILLER_33_7 ();
 sg13g2_decap_4 FILLER_33_21 ();
 sg13g2_fill_1 FILLER_33_25 ();
 sg13g2_decap_8 FILLER_33_30 ();
 sg13g2_decap_4 FILLER_33_37 ();
 sg13g2_fill_2 FILLER_33_46 ();
 sg13g2_fill_2 FILLER_33_58 ();
 sg13g2_fill_1 FILLER_33_60 ();
 sg13g2_decap_8 FILLER_33_71 ();
 sg13g2_decap_4 FILLER_33_78 ();
 sg13g2_fill_2 FILLER_33_82 ();
 sg13g2_decap_8 FILLER_33_99 ();
 sg13g2_decap_8 FILLER_33_106 ();
 sg13g2_decap_8 FILLER_33_113 ();
 sg13g2_decap_8 FILLER_33_120 ();
 sg13g2_decap_4 FILLER_33_127 ();
 sg13g2_fill_2 FILLER_33_131 ();
 sg13g2_fill_2 FILLER_33_141 ();
 sg13g2_decap_8 FILLER_33_148 ();
 sg13g2_decap_8 FILLER_33_155 ();
 sg13g2_decap_8 FILLER_33_162 ();
 sg13g2_fill_2 FILLER_33_169 ();
 sg13g2_fill_1 FILLER_33_171 ();
 sg13g2_decap_4 FILLER_33_186 ();
 sg13g2_fill_2 FILLER_33_190 ();
 sg13g2_fill_2 FILLER_33_202 ();
 sg13g2_decap_4 FILLER_33_210 ();
 sg13g2_fill_1 FILLER_33_214 ();
 sg13g2_fill_2 FILLER_33_225 ();
 sg13g2_fill_2 FILLER_33_232 ();
 sg13g2_fill_2 FILLER_33_244 ();
 sg13g2_fill_1 FILLER_33_246 ();
 sg13g2_decap_8 FILLER_33_255 ();
 sg13g2_fill_2 FILLER_33_262 ();
 sg13g2_decap_8 FILLER_33_268 ();
 sg13g2_decap_8 FILLER_33_275 ();
 sg13g2_decap_8 FILLER_33_282 ();
 sg13g2_decap_8 FILLER_33_289 ();
 sg13g2_fill_1 FILLER_33_296 ();
 sg13g2_decap_8 FILLER_33_301 ();
 sg13g2_decap_8 FILLER_33_308 ();
 sg13g2_decap_8 FILLER_33_315 ();
 sg13g2_decap_8 FILLER_33_322 ();
 sg13g2_fill_2 FILLER_33_329 ();
 sg13g2_decap_8 FILLER_33_339 ();
 sg13g2_decap_8 FILLER_33_346 ();
 sg13g2_decap_8 FILLER_33_353 ();
 sg13g2_decap_8 FILLER_33_360 ();
 sg13g2_decap_8 FILLER_33_367 ();
 sg13g2_decap_8 FILLER_33_374 ();
 sg13g2_decap_8 FILLER_33_381 ();
 sg13g2_decap_4 FILLER_33_388 ();
 sg13g2_decap_8 FILLER_33_416 ();
 sg13g2_decap_4 FILLER_33_466 ();
 sg13g2_fill_2 FILLER_33_470 ();
 sg13g2_fill_2 FILLER_33_476 ();
 sg13g2_fill_1 FILLER_33_478 ();
 sg13g2_fill_2 FILLER_33_483 ();
 sg13g2_fill_2 FILLER_33_506 ();
 sg13g2_fill_2 FILLER_33_513 ();
 sg13g2_fill_2 FILLER_33_520 ();
 sg13g2_fill_1 FILLER_33_522 ();
 sg13g2_decap_8 FILLER_33_531 ();
 sg13g2_fill_1 FILLER_33_538 ();
 sg13g2_fill_1 FILLER_33_575 ();
 sg13g2_decap_4 FILLER_33_617 ();
 sg13g2_decap_4 FILLER_33_661 ();
 sg13g2_fill_1 FILLER_33_665 ();
 sg13g2_fill_2 FILLER_33_680 ();
 sg13g2_fill_1 FILLER_33_682 ();
 sg13g2_fill_1 FILLER_33_709 ();
 sg13g2_fill_2 FILLER_33_733 ();
 sg13g2_fill_1 FILLER_33_735 ();
 sg13g2_decap_8 FILLER_33_746 ();
 sg13g2_decap_8 FILLER_33_757 ();
 sg13g2_decap_8 FILLER_33_764 ();
 sg13g2_decap_4 FILLER_33_771 ();
 sg13g2_fill_2 FILLER_33_775 ();
 sg13g2_decap_8 FILLER_33_791 ();
 sg13g2_decap_8 FILLER_33_798 ();
 sg13g2_decap_8 FILLER_33_805 ();
 sg13g2_decap_8 FILLER_33_812 ();
 sg13g2_decap_8 FILLER_33_819 ();
 sg13g2_decap_8 FILLER_33_826 ();
 sg13g2_decap_8 FILLER_33_833 ();
 sg13g2_decap_8 FILLER_33_840 ();
 sg13g2_decap_8 FILLER_33_847 ();
 sg13g2_decap_8 FILLER_33_854 ();
 sg13g2_decap_8 FILLER_33_861 ();
 sg13g2_decap_8 FILLER_33_868 ();
 sg13g2_fill_2 FILLER_33_875 ();
 sg13g2_fill_1 FILLER_33_877 ();
 sg13g2_decap_8 FILLER_34_0 ();
 sg13g2_fill_2 FILLER_34_7 ();
 sg13g2_fill_1 FILLER_34_9 ();
 sg13g2_fill_2 FILLER_34_18 ();
 sg13g2_decap_8 FILLER_34_24 ();
 sg13g2_decap_8 FILLER_34_31 ();
 sg13g2_decap_4 FILLER_34_38 ();
 sg13g2_fill_2 FILLER_34_42 ();
 sg13g2_fill_1 FILLER_34_48 ();
 sg13g2_decap_8 FILLER_34_59 ();
 sg13g2_decap_8 FILLER_34_66 ();
 sg13g2_decap_4 FILLER_34_73 ();
 sg13g2_decap_8 FILLER_34_94 ();
 sg13g2_decap_4 FILLER_34_101 ();
 sg13g2_fill_1 FILLER_34_105 ();
 sg13g2_fill_1 FILLER_34_110 ();
 sg13g2_fill_1 FILLER_34_119 ();
 sg13g2_decap_8 FILLER_34_128 ();
 sg13g2_decap_8 FILLER_34_135 ();
 sg13g2_fill_1 FILLER_34_142 ();
 sg13g2_decap_8 FILLER_34_156 ();
 sg13g2_fill_2 FILLER_34_163 ();
 sg13g2_fill_1 FILLER_34_204 ();
 sg13g2_decap_4 FILLER_34_210 ();
 sg13g2_fill_2 FILLER_34_214 ();
 sg13g2_decap_8 FILLER_34_229 ();
 sg13g2_fill_1 FILLER_34_236 ();
 sg13g2_decap_8 FILLER_34_257 ();
 sg13g2_decap_8 FILLER_34_264 ();
 sg13g2_decap_8 FILLER_34_271 ();
 sg13g2_decap_4 FILLER_34_278 ();
 sg13g2_fill_2 FILLER_34_282 ();
 sg13g2_decap_8 FILLER_34_292 ();
 sg13g2_fill_1 FILLER_34_299 ();
 sg13g2_decap_4 FILLER_34_316 ();
 sg13g2_fill_1 FILLER_34_320 ();
 sg13g2_decap_8 FILLER_34_333 ();
 sg13g2_decap_8 FILLER_34_340 ();
 sg13g2_decap_8 FILLER_34_347 ();
 sg13g2_decap_8 FILLER_34_354 ();
 sg13g2_decap_8 FILLER_34_361 ();
 sg13g2_decap_8 FILLER_34_368 ();
 sg13g2_decap_8 FILLER_34_375 ();
 sg13g2_decap_8 FILLER_34_382 ();
 sg13g2_decap_4 FILLER_34_389 ();
 sg13g2_decap_8 FILLER_34_397 ();
 sg13g2_fill_2 FILLER_34_404 ();
 sg13g2_decap_8 FILLER_34_416 ();
 sg13g2_decap_8 FILLER_34_423 ();
 sg13g2_fill_1 FILLER_34_430 ();
 sg13g2_decap_4 FILLER_34_440 ();
 sg13g2_decap_4 FILLER_34_452 ();
 sg13g2_fill_1 FILLER_34_456 ();
 sg13g2_decap_8 FILLER_34_461 ();
 sg13g2_decap_8 FILLER_34_468 ();
 sg13g2_fill_1 FILLER_34_475 ();
 sg13g2_fill_1 FILLER_34_507 ();
 sg13g2_fill_2 FILLER_34_511 ();
 sg13g2_fill_1 FILLER_34_513 ();
 sg13g2_fill_1 FILLER_34_524 ();
 sg13g2_decap_4 FILLER_34_551 ();
 sg13g2_fill_2 FILLER_34_555 ();
 sg13g2_decap_4 FILLER_34_561 ();
 sg13g2_fill_2 FILLER_34_565 ();
 sg13g2_fill_2 FILLER_34_577 ();
 sg13g2_fill_1 FILLER_34_579 ();
 sg13g2_fill_1 FILLER_34_584 ();
 sg13g2_fill_2 FILLER_34_593 ();
 sg13g2_decap_8 FILLER_34_602 ();
 sg13g2_decap_8 FILLER_34_609 ();
 sg13g2_decap_8 FILLER_34_616 ();
 sg13g2_decap_4 FILLER_34_623 ();
 sg13g2_fill_1 FILLER_34_627 ();
 sg13g2_decap_8 FILLER_34_633 ();
 sg13g2_fill_2 FILLER_34_640 ();
 sg13g2_decap_8 FILLER_34_659 ();
 sg13g2_decap_8 FILLER_34_666 ();
 sg13g2_decap_8 FILLER_34_699 ();
 sg13g2_fill_2 FILLER_34_706 ();
 sg13g2_fill_2 FILLER_34_734 ();
 sg13g2_decap_4 FILLER_34_740 ();
 sg13g2_fill_2 FILLER_34_744 ();
 sg13g2_decap_8 FILLER_34_772 ();
 sg13g2_decap_8 FILLER_34_779 ();
 sg13g2_decap_8 FILLER_34_786 ();
 sg13g2_decap_8 FILLER_34_793 ();
 sg13g2_decap_8 FILLER_34_800 ();
 sg13g2_decap_8 FILLER_34_807 ();
 sg13g2_decap_8 FILLER_34_814 ();
 sg13g2_decap_8 FILLER_34_821 ();
 sg13g2_decap_8 FILLER_34_828 ();
 sg13g2_decap_8 FILLER_34_835 ();
 sg13g2_decap_8 FILLER_34_842 ();
 sg13g2_decap_8 FILLER_34_849 ();
 sg13g2_decap_8 FILLER_34_856 ();
 sg13g2_decap_8 FILLER_34_863 ();
 sg13g2_decap_8 FILLER_34_870 ();
 sg13g2_fill_1 FILLER_34_877 ();
 sg13g2_decap_8 FILLER_35_0 ();
 sg13g2_decap_4 FILLER_35_7 ();
 sg13g2_fill_2 FILLER_35_11 ();
 sg13g2_decap_8 FILLER_35_30 ();
 sg13g2_decap_4 FILLER_35_37 ();
 sg13g2_fill_2 FILLER_35_41 ();
 sg13g2_decap_8 FILLER_35_59 ();
 sg13g2_decap_8 FILLER_35_66 ();
 sg13g2_decap_8 FILLER_35_95 ();
 sg13g2_fill_2 FILLER_35_102 ();
 sg13g2_fill_1 FILLER_35_104 ();
 sg13g2_fill_1 FILLER_35_121 ();
 sg13g2_fill_1 FILLER_35_127 ();
 sg13g2_fill_1 FILLER_35_133 ();
 sg13g2_fill_1 FILLER_35_139 ();
 sg13g2_decap_8 FILLER_35_166 ();
 sg13g2_fill_2 FILLER_35_173 ();
 sg13g2_fill_1 FILLER_35_175 ();
 sg13g2_decap_4 FILLER_35_184 ();
 sg13g2_decap_8 FILLER_35_200 ();
 sg13g2_decap_8 FILLER_35_207 ();
 sg13g2_decap_4 FILLER_35_214 ();
 sg13g2_fill_1 FILLER_35_218 ();
 sg13g2_fill_2 FILLER_35_232 ();
 sg13g2_fill_1 FILLER_35_239 ();
 sg13g2_decap_8 FILLER_35_261 ();
 sg13g2_decap_8 FILLER_35_268 ();
 sg13g2_fill_2 FILLER_35_275 ();
 sg13g2_fill_2 FILLER_35_305 ();
 sg13g2_decap_4 FILLER_35_317 ();
 sg13g2_decap_8 FILLER_35_325 ();
 sg13g2_decap_8 FILLER_35_332 ();
 sg13g2_fill_1 FILLER_35_339 ();
 sg13g2_fill_1 FILLER_35_365 ();
 sg13g2_decap_8 FILLER_35_378 ();
 sg13g2_decap_4 FILLER_35_385 ();
 sg13g2_fill_1 FILLER_35_389 ();
 sg13g2_fill_2 FILLER_35_394 ();
 sg13g2_fill_2 FILLER_35_421 ();
 sg13g2_fill_1 FILLER_35_423 ();
 sg13g2_decap_4 FILLER_35_428 ();
 sg13g2_fill_2 FILLER_35_440 ();
 sg13g2_fill_2 FILLER_35_451 ();
 sg13g2_decap_8 FILLER_35_461 ();
 sg13g2_decap_8 FILLER_35_468 ();
 sg13g2_decap_4 FILLER_35_475 ();
 sg13g2_fill_1 FILLER_35_479 ();
 sg13g2_fill_1 FILLER_35_484 ();
 sg13g2_fill_2 FILLER_35_490 ();
 sg13g2_decap_4 FILLER_35_496 ();
 sg13g2_fill_2 FILLER_35_500 ();
 sg13g2_decap_8 FILLER_35_511 ();
 sg13g2_decap_4 FILLER_35_518 ();
 sg13g2_decap_4 FILLER_35_539 ();
 sg13g2_fill_1 FILLER_35_543 ();
 sg13g2_fill_2 FILLER_35_570 ();
 sg13g2_fill_2 FILLER_35_598 ();
 sg13g2_fill_1 FILLER_35_600 ();
 sg13g2_fill_2 FILLER_35_614 ();
 sg13g2_fill_1 FILLER_35_616 ();
 sg13g2_fill_2 FILLER_35_622 ();
 sg13g2_fill_1 FILLER_35_624 ();
 sg13g2_fill_2 FILLER_35_630 ();
 sg13g2_fill_1 FILLER_35_632 ();
 sg13g2_fill_2 FILLER_35_646 ();
 sg13g2_decap_8 FILLER_35_652 ();
 sg13g2_decap_8 FILLER_35_659 ();
 sg13g2_decap_8 FILLER_35_666 ();
 sg13g2_decap_4 FILLER_35_673 ();
 sg13g2_fill_2 FILLER_35_677 ();
 sg13g2_decap_8 FILLER_35_683 ();
 sg13g2_decap_8 FILLER_35_690 ();
 sg13g2_fill_2 FILLER_35_697 ();
 sg13g2_fill_1 FILLER_35_699 ();
 sg13g2_decap_8 FILLER_35_704 ();
 sg13g2_fill_2 FILLER_35_711 ();
 sg13g2_fill_1 FILLER_35_713 ();
 sg13g2_fill_1 FILLER_35_722 ();
 sg13g2_fill_2 FILLER_35_736 ();
 sg13g2_fill_1 FILLER_35_738 ();
 sg13g2_decap_8 FILLER_35_744 ();
 sg13g2_decap_8 FILLER_35_751 ();
 sg13g2_decap_4 FILLER_35_758 ();
 sg13g2_fill_2 FILLER_35_762 ();
 sg13g2_decap_8 FILLER_35_790 ();
 sg13g2_decap_8 FILLER_35_797 ();
 sg13g2_decap_8 FILLER_35_804 ();
 sg13g2_decap_8 FILLER_35_811 ();
 sg13g2_decap_8 FILLER_35_818 ();
 sg13g2_decap_8 FILLER_35_825 ();
 sg13g2_decap_8 FILLER_35_832 ();
 sg13g2_decap_8 FILLER_35_839 ();
 sg13g2_decap_8 FILLER_35_846 ();
 sg13g2_decap_8 FILLER_35_853 ();
 sg13g2_decap_8 FILLER_35_860 ();
 sg13g2_decap_8 FILLER_35_867 ();
 sg13g2_decap_4 FILLER_35_874 ();
 sg13g2_decap_8 FILLER_36_0 ();
 sg13g2_decap_8 FILLER_36_7 ();
 sg13g2_fill_2 FILLER_36_18 ();
 sg13g2_fill_2 FILLER_36_24 ();
 sg13g2_decap_8 FILLER_36_35 ();
 sg13g2_decap_8 FILLER_36_50 ();
 sg13g2_fill_2 FILLER_36_57 ();
 sg13g2_fill_1 FILLER_36_59 ();
 sg13g2_decap_4 FILLER_36_72 ();
 sg13g2_fill_1 FILLER_36_76 ();
 sg13g2_decap_8 FILLER_36_96 ();
 sg13g2_decap_8 FILLER_36_103 ();
 sg13g2_decap_8 FILLER_36_110 ();
 sg13g2_fill_2 FILLER_36_121 ();
 sg13g2_decap_4 FILLER_36_127 ();
 sg13g2_fill_2 FILLER_36_135 ();
 sg13g2_fill_1 FILLER_36_146 ();
 sg13g2_decap_8 FILLER_36_151 ();
 sg13g2_decap_4 FILLER_36_158 ();
 sg13g2_fill_1 FILLER_36_162 ();
 sg13g2_decap_8 FILLER_36_167 ();
 sg13g2_decap_4 FILLER_36_174 ();
 sg13g2_fill_2 FILLER_36_178 ();
 sg13g2_fill_2 FILLER_36_185 ();
 sg13g2_fill_1 FILLER_36_187 ();
 sg13g2_decap_8 FILLER_36_202 ();
 sg13g2_decap_4 FILLER_36_209 ();
 sg13g2_fill_1 FILLER_36_213 ();
 sg13g2_decap_4 FILLER_36_222 ();
 sg13g2_fill_1 FILLER_36_226 ();
 sg13g2_fill_1 FILLER_36_236 ();
 sg13g2_fill_2 FILLER_36_245 ();
 sg13g2_decap_8 FILLER_36_258 ();
 sg13g2_decap_8 FILLER_36_265 ();
 sg13g2_fill_2 FILLER_36_272 ();
 sg13g2_fill_2 FILLER_36_281 ();
 sg13g2_fill_1 FILLER_36_283 ();
 sg13g2_fill_2 FILLER_36_289 ();
 sg13g2_fill_1 FILLER_36_295 ();
 sg13g2_decap_8 FILLER_36_302 ();
 sg13g2_fill_2 FILLER_36_309 ();
 sg13g2_fill_1 FILLER_36_311 ();
 sg13g2_decap_8 FILLER_36_321 ();
 sg13g2_decap_8 FILLER_36_328 ();
 sg13g2_fill_1 FILLER_36_335 ();
 sg13g2_fill_2 FILLER_36_340 ();
 sg13g2_fill_1 FILLER_36_342 ();
 sg13g2_decap_4 FILLER_36_347 ();
 sg13g2_decap_4 FILLER_36_379 ();
 sg13g2_fill_2 FILLER_36_393 ();
 sg13g2_fill_1 FILLER_36_400 ();
 sg13g2_decap_8 FILLER_36_414 ();
 sg13g2_decap_4 FILLER_36_426 ();
 sg13g2_fill_1 FILLER_36_430 ();
 sg13g2_decap_4 FILLER_36_439 ();
 sg13g2_decap_4 FILLER_36_447 ();
 sg13g2_fill_2 FILLER_36_459 ();
 sg13g2_fill_1 FILLER_36_461 ();
 sg13g2_decap_8 FILLER_36_467 ();
 sg13g2_fill_1 FILLER_36_474 ();
 sg13g2_decap_8 FILLER_36_501 ();
 sg13g2_fill_2 FILLER_36_508 ();
 sg13g2_decap_8 FILLER_36_519 ();
 sg13g2_decap_8 FILLER_36_526 ();
 sg13g2_decap_8 FILLER_36_533 ();
 sg13g2_decap_8 FILLER_36_540 ();
 sg13g2_decap_4 FILLER_36_547 ();
 sg13g2_decap_8 FILLER_36_555 ();
 sg13g2_decap_8 FILLER_36_562 ();
 sg13g2_decap_8 FILLER_36_569 ();
 sg13g2_fill_2 FILLER_36_576 ();
 sg13g2_fill_1 FILLER_36_578 ();
 sg13g2_decap_8 FILLER_36_583 ();
 sg13g2_decap_8 FILLER_36_590 ();
 sg13g2_decap_8 FILLER_36_597 ();
 sg13g2_decap_8 FILLER_36_604 ();
 sg13g2_decap_8 FILLER_36_611 ();
 sg13g2_decap_4 FILLER_36_618 ();
 sg13g2_fill_2 FILLER_36_639 ();
 sg13g2_decap_8 FILLER_36_658 ();
 sg13g2_decap_8 FILLER_36_665 ();
 sg13g2_decap_8 FILLER_36_672 ();
 sg13g2_decap_8 FILLER_36_679 ();
 sg13g2_fill_2 FILLER_36_686 ();
 sg13g2_fill_1 FILLER_36_688 ();
 sg13g2_decap_4 FILLER_36_719 ();
 sg13g2_decap_4 FILLER_36_753 ();
 sg13g2_decap_8 FILLER_36_761 ();
 sg13g2_decap_4 FILLER_36_768 ();
 sg13g2_fill_1 FILLER_36_772 ();
 sg13g2_decap_8 FILLER_36_777 ();
 sg13g2_decap_4 FILLER_36_784 ();
 sg13g2_fill_2 FILLER_36_788 ();
 sg13g2_decap_8 FILLER_36_803 ();
 sg13g2_decap_8 FILLER_36_810 ();
 sg13g2_decap_8 FILLER_36_817 ();
 sg13g2_decap_8 FILLER_36_824 ();
 sg13g2_decap_8 FILLER_36_831 ();
 sg13g2_decap_8 FILLER_36_838 ();
 sg13g2_decap_8 FILLER_36_845 ();
 sg13g2_decap_8 FILLER_36_852 ();
 sg13g2_decap_8 FILLER_36_859 ();
 sg13g2_decap_8 FILLER_36_866 ();
 sg13g2_decap_4 FILLER_36_873 ();
 sg13g2_fill_1 FILLER_36_877 ();
 sg13g2_fill_2 FILLER_37_26 ();
 sg13g2_fill_2 FILLER_37_33 ();
 sg13g2_fill_1 FILLER_37_35 ();
 sg13g2_decap_8 FILLER_37_67 ();
 sg13g2_decap_8 FILLER_37_74 ();
 sg13g2_decap_4 FILLER_37_81 ();
 sg13g2_fill_1 FILLER_37_85 ();
 sg13g2_decap_4 FILLER_37_90 ();
 sg13g2_decap_8 FILLER_37_134 ();
 sg13g2_decap_8 FILLER_37_141 ();
 sg13g2_fill_1 FILLER_37_148 ();
 sg13g2_decap_8 FILLER_37_153 ();
 sg13g2_decap_8 FILLER_37_160 ();
 sg13g2_decap_8 FILLER_37_167 ();
 sg13g2_fill_2 FILLER_37_174 ();
 sg13g2_fill_1 FILLER_37_176 ();
 sg13g2_fill_2 FILLER_37_201 ();
 sg13g2_decap_8 FILLER_37_209 ();
 sg13g2_fill_2 FILLER_37_216 ();
 sg13g2_fill_1 FILLER_37_218 ();
 sg13g2_fill_1 FILLER_37_240 ();
 sg13g2_fill_1 FILLER_37_246 ();
 sg13g2_decap_8 FILLER_37_265 ();
 sg13g2_decap_4 FILLER_37_272 ();
 sg13g2_fill_2 FILLER_37_276 ();
 sg13g2_fill_1 FILLER_37_291 ();
 sg13g2_decap_8 FILLER_37_304 ();
 sg13g2_decap_4 FILLER_37_315 ();
 sg13g2_decap_4 FILLER_37_327 ();
 sg13g2_fill_1 FILLER_37_331 ();
 sg13g2_fill_1 FILLER_37_340 ();
 sg13g2_fill_2 FILLER_37_349 ();
 sg13g2_fill_2 FILLER_37_355 ();
 sg13g2_fill_2 FILLER_37_365 ();
 sg13g2_fill_1 FILLER_37_367 ();
 sg13g2_decap_4 FILLER_37_372 ();
 sg13g2_fill_2 FILLER_37_376 ();
 sg13g2_fill_2 FILLER_37_382 ();
 sg13g2_fill_1 FILLER_37_403 ();
 sg13g2_fill_2 FILLER_37_430 ();
 sg13g2_fill_1 FILLER_37_432 ();
 sg13g2_decap_8 FILLER_37_461 ();
 sg13g2_decap_8 FILLER_37_468 ();
 sg13g2_decap_8 FILLER_37_475 ();
 sg13g2_decap_4 FILLER_37_482 ();
 sg13g2_decap_8 FILLER_37_499 ();
 sg13g2_fill_2 FILLER_37_506 ();
 sg13g2_fill_1 FILLER_37_508 ();
 sg13g2_decap_8 FILLER_37_544 ();
 sg13g2_decap_4 FILLER_37_551 ();
 sg13g2_fill_1 FILLER_37_555 ();
 sg13g2_decap_8 FILLER_37_560 ();
 sg13g2_decap_8 FILLER_37_567 ();
 sg13g2_decap_8 FILLER_37_574 ();
 sg13g2_decap_8 FILLER_37_581 ();
 sg13g2_fill_1 FILLER_37_588 ();
 sg13g2_decap_8 FILLER_37_615 ();
 sg13g2_decap_8 FILLER_37_622 ();
 sg13g2_decap_4 FILLER_37_629 ();
 sg13g2_decap_8 FILLER_37_638 ();
 sg13g2_decap_8 FILLER_37_645 ();
 sg13g2_decap_8 FILLER_37_652 ();
 sg13g2_decap_8 FILLER_37_659 ();
 sg13g2_decap_8 FILLER_37_666 ();
 sg13g2_decap_8 FILLER_37_673 ();
 sg13g2_decap_8 FILLER_37_692 ();
 sg13g2_decap_8 FILLER_37_699 ();
 sg13g2_decap_8 FILLER_37_706 ();
 sg13g2_decap_4 FILLER_37_713 ();
 sg13g2_decap_8 FILLER_37_725 ();
 sg13g2_fill_2 FILLER_37_732 ();
 sg13g2_decap_8 FILLER_37_738 ();
 sg13g2_decap_8 FILLER_37_750 ();
 sg13g2_decap_8 FILLER_37_757 ();
 sg13g2_decap_8 FILLER_37_764 ();
 sg13g2_decap_8 FILLER_37_771 ();
 sg13g2_fill_2 FILLER_37_778 ();
 sg13g2_decap_4 FILLER_37_785 ();
 sg13g2_fill_2 FILLER_37_789 ();
 sg13g2_decap_8 FILLER_37_804 ();
 sg13g2_decap_8 FILLER_37_811 ();
 sg13g2_decap_8 FILLER_37_818 ();
 sg13g2_decap_8 FILLER_37_825 ();
 sg13g2_decap_8 FILLER_37_832 ();
 sg13g2_decap_8 FILLER_37_839 ();
 sg13g2_decap_8 FILLER_37_846 ();
 sg13g2_decap_8 FILLER_37_853 ();
 sg13g2_decap_8 FILLER_37_860 ();
 sg13g2_decap_8 FILLER_37_867 ();
 sg13g2_decap_4 FILLER_37_874 ();
 sg13g2_decap_8 FILLER_38_0 ();
 sg13g2_decap_8 FILLER_38_11 ();
 sg13g2_decap_4 FILLER_38_18 ();
 sg13g2_fill_2 FILLER_38_22 ();
 sg13g2_decap_8 FILLER_38_33 ();
 sg13g2_fill_2 FILLER_38_40 ();
 sg13g2_fill_1 FILLER_38_42 ();
 sg13g2_fill_1 FILLER_38_47 ();
 sg13g2_fill_2 FILLER_38_59 ();
 sg13g2_fill_2 FILLER_38_78 ();
 sg13g2_fill_1 FILLER_38_80 ();
 sg13g2_decap_4 FILLER_38_86 ();
 sg13g2_decap_4 FILLER_38_94 ();
 sg13g2_fill_2 FILLER_38_102 ();
 sg13g2_fill_1 FILLER_38_104 ();
 sg13g2_fill_2 FILLER_38_117 ();
 sg13g2_fill_1 FILLER_38_119 ();
 sg13g2_decap_8 FILLER_38_125 ();
 sg13g2_fill_1 FILLER_38_132 ();
 sg13g2_decap_8 FILLER_38_168 ();
 sg13g2_decap_8 FILLER_38_175 ();
 sg13g2_decap_8 FILLER_38_182 ();
 sg13g2_decap_8 FILLER_38_201 ();
 sg13g2_fill_2 FILLER_38_208 ();
 sg13g2_fill_1 FILLER_38_218 ();
 sg13g2_fill_2 FILLER_38_239 ();
 sg13g2_fill_2 FILLER_38_245 ();
 sg13g2_decap_8 FILLER_38_264 ();
 sg13g2_decap_8 FILLER_38_271 ();
 sg13g2_fill_1 FILLER_38_278 ();
 sg13g2_fill_1 FILLER_38_287 ();
 sg13g2_fill_1 FILLER_38_293 ();
 sg13g2_decap_8 FILLER_38_302 ();
 sg13g2_fill_1 FILLER_38_309 ();
 sg13g2_fill_2 FILLER_38_318 ();
 sg13g2_fill_1 FILLER_38_320 ();
 sg13g2_decap_8 FILLER_38_334 ();
 sg13g2_fill_2 FILLER_38_351 ();
 sg13g2_decap_8 FILLER_38_362 ();
 sg13g2_fill_2 FILLER_38_369 ();
 sg13g2_decap_8 FILLER_38_375 ();
 sg13g2_decap_8 FILLER_38_382 ();
 sg13g2_fill_2 FILLER_38_389 ();
 sg13g2_fill_1 FILLER_38_391 ();
 sg13g2_fill_1 FILLER_38_399 ();
 sg13g2_decap_8 FILLER_38_417 ();
 sg13g2_fill_2 FILLER_38_424 ();
 sg13g2_decap_4 FILLER_38_431 ();
 sg13g2_fill_1 FILLER_38_435 ();
 sg13g2_decap_4 FILLER_38_440 ();
 sg13g2_fill_1 FILLER_38_444 ();
 sg13g2_decap_8 FILLER_38_461 ();
 sg13g2_decap_8 FILLER_38_468 ();
 sg13g2_decap_8 FILLER_38_475 ();
 sg13g2_fill_2 FILLER_38_482 ();
 sg13g2_decap_8 FILLER_38_510 ();
 sg13g2_decap_4 FILLER_38_517 ();
 sg13g2_fill_1 FILLER_38_521 ();
 sg13g2_decap_8 FILLER_38_529 ();
 sg13g2_fill_2 FILLER_38_536 ();
 sg13g2_fill_1 FILLER_38_538 ();
 sg13g2_decap_4 FILLER_38_543 ();
 sg13g2_fill_2 FILLER_38_547 ();
 sg13g2_decap_8 FILLER_38_575 ();
 sg13g2_decap_4 FILLER_38_582 ();
 sg13g2_fill_2 FILLER_38_586 ();
 sg13g2_fill_1 FILLER_38_592 ();
 sg13g2_decap_8 FILLER_38_610 ();
 sg13g2_decap_8 FILLER_38_622 ();
 sg13g2_decap_8 FILLER_38_629 ();
 sg13g2_decap_4 FILLER_38_636 ();
 sg13g2_fill_1 FILLER_38_640 ();
 sg13g2_decap_8 FILLER_38_654 ();
 sg13g2_decap_8 FILLER_38_661 ();
 sg13g2_decap_8 FILLER_38_668 ();
 sg13g2_decap_8 FILLER_38_675 ();
 sg13g2_decap_8 FILLER_38_686 ();
 sg13g2_decap_4 FILLER_38_693 ();
 sg13g2_decap_8 FILLER_38_702 ();
 sg13g2_decap_8 FILLER_38_709 ();
 sg13g2_fill_2 FILLER_38_716 ();
 sg13g2_decap_8 FILLER_38_742 ();
 sg13g2_decap_4 FILLER_38_749 ();
 sg13g2_fill_2 FILLER_38_765 ();
 sg13g2_fill_1 FILLER_38_767 ();
 sg13g2_decap_4 FILLER_38_811 ();
 sg13g2_fill_2 FILLER_38_815 ();
 sg13g2_decap_8 FILLER_38_830 ();
 sg13g2_fill_2 FILLER_38_837 ();
 sg13g2_fill_1 FILLER_38_839 ();
 sg13g2_decap_8 FILLER_38_844 ();
 sg13g2_decap_8 FILLER_38_851 ();
 sg13g2_decap_8 FILLER_38_858 ();
 sg13g2_decap_8 FILLER_38_865 ();
 sg13g2_decap_4 FILLER_38_872 ();
 sg13g2_fill_2 FILLER_38_876 ();
 sg13g2_decap_8 FILLER_39_30 ();
 sg13g2_decap_8 FILLER_39_37 ();
 sg13g2_fill_2 FILLER_39_52 ();
 sg13g2_decap_8 FILLER_39_59 ();
 sg13g2_fill_2 FILLER_39_66 ();
 sg13g2_fill_1 FILLER_39_68 ();
 sg13g2_decap_4 FILLER_39_77 ();
 sg13g2_fill_2 FILLER_39_81 ();
 sg13g2_decap_8 FILLER_39_109 ();
 sg13g2_decap_4 FILLER_39_116 ();
 sg13g2_fill_2 FILLER_39_120 ();
 sg13g2_fill_1 FILLER_39_127 ();
 sg13g2_fill_2 FILLER_39_132 ();
 sg13g2_decap_8 FILLER_39_138 ();
 sg13g2_decap_4 FILLER_39_145 ();
 sg13g2_decap_8 FILLER_39_168 ();
 sg13g2_fill_2 FILLER_39_175 ();
 sg13g2_decap_8 FILLER_39_185 ();
 sg13g2_fill_2 FILLER_39_192 ();
 sg13g2_decap_8 FILLER_39_202 ();
 sg13g2_decap_8 FILLER_39_209 ();
 sg13g2_fill_2 FILLER_39_216 ();
 sg13g2_decap_8 FILLER_39_262 ();
 sg13g2_decap_8 FILLER_39_269 ();
 sg13g2_fill_1 FILLER_39_284 ();
 sg13g2_fill_1 FILLER_39_295 ();
 sg13g2_fill_1 FILLER_39_301 ();
 sg13g2_fill_1 FILLER_39_316 ();
 sg13g2_fill_1 FILLER_39_321 ();
 sg13g2_fill_2 FILLER_39_340 ();
 sg13g2_decap_4 FILLER_39_347 ();
 sg13g2_fill_1 FILLER_39_351 ();
 sg13g2_decap_4 FILLER_39_360 ();
 sg13g2_decap_8 FILLER_39_397 ();
 sg13g2_decap_8 FILLER_39_404 ();
 sg13g2_fill_1 FILLER_39_411 ();
 sg13g2_fill_2 FILLER_39_421 ();
 sg13g2_fill_1 FILLER_39_423 ();
 sg13g2_fill_2 FILLER_39_428 ();
 sg13g2_decap_8 FILLER_39_441 ();
 sg13g2_decap_8 FILLER_39_448 ();
 sg13g2_decap_8 FILLER_39_465 ();
 sg13g2_decap_8 FILLER_39_472 ();
 sg13g2_fill_1 FILLER_39_505 ();
 sg13g2_fill_2 FILLER_39_549 ();
 sg13g2_fill_1 FILLER_39_551 ();
 sg13g2_decap_8 FILLER_39_556 ();
 sg13g2_decap_8 FILLER_39_563 ();
 sg13g2_decap_8 FILLER_39_570 ();
 sg13g2_decap_8 FILLER_39_577 ();
 sg13g2_fill_1 FILLER_39_584 ();
 sg13g2_decap_4 FILLER_39_589 ();
 sg13g2_fill_2 FILLER_39_593 ();
 sg13g2_decap_8 FILLER_39_599 ();
 sg13g2_fill_1 FILLER_39_606 ();
 sg13g2_decap_8 FILLER_39_612 ();
 sg13g2_fill_2 FILLER_39_619 ();
 sg13g2_fill_1 FILLER_39_621 ();
 sg13g2_decap_8 FILLER_39_627 ();
 sg13g2_decap_4 FILLER_39_634 ();
 sg13g2_fill_1 FILLER_39_638 ();
 sg13g2_decap_8 FILLER_39_648 ();
 sg13g2_fill_2 FILLER_39_655 ();
 sg13g2_decap_4 FILLER_39_675 ();
 sg13g2_fill_2 FILLER_39_679 ();
 sg13g2_decap_8 FILLER_39_691 ();
 sg13g2_decap_8 FILLER_39_707 ();
 sg13g2_decap_8 FILLER_39_714 ();
 sg13g2_fill_2 FILLER_39_721 ();
 sg13g2_fill_1 FILLER_39_723 ();
 sg13g2_fill_1 FILLER_39_729 ();
 sg13g2_fill_2 FILLER_39_773 ();
 sg13g2_fill_1 FILLER_39_775 ();
 sg13g2_fill_1 FILLER_39_780 ();
 sg13g2_fill_1 FILLER_39_794 ();
 sg13g2_decap_8 FILLER_39_808 ();
 sg13g2_fill_2 FILLER_39_815 ();
 sg13g2_decap_8 FILLER_39_827 ();
 sg13g2_decap_8 FILLER_39_834 ();
 sg13g2_fill_1 FILLER_39_841 ();
 sg13g2_decap_8 FILLER_39_846 ();
 sg13g2_decap_8 FILLER_39_853 ();
 sg13g2_decap_8 FILLER_39_860 ();
 sg13g2_decap_8 FILLER_39_867 ();
 sg13g2_decap_4 FILLER_39_874 ();
 sg13g2_decap_8 FILLER_40_0 ();
 sg13g2_fill_2 FILLER_40_7 ();
 sg13g2_fill_1 FILLER_40_9 ();
 sg13g2_fill_2 FILLER_40_14 ();
 sg13g2_fill_1 FILLER_40_16 ();
 sg13g2_decap_4 FILLER_40_31 ();
 sg13g2_fill_2 FILLER_40_35 ();
 sg13g2_fill_1 FILLER_40_42 ();
 sg13g2_fill_2 FILLER_40_52 ();
 sg13g2_fill_2 FILLER_40_59 ();
 sg13g2_fill_1 FILLER_40_65 ();
 sg13g2_decap_8 FILLER_40_70 ();
 sg13g2_decap_8 FILLER_40_77 ();
 sg13g2_fill_2 FILLER_40_84 ();
 sg13g2_decap_8 FILLER_40_103 ();
 sg13g2_decap_8 FILLER_40_110 ();
 sg13g2_decap_4 FILLER_40_117 ();
 sg13g2_fill_1 FILLER_40_121 ();
 sg13g2_fill_1 FILLER_40_152 ();
 sg13g2_decap_8 FILLER_40_166 ();
 sg13g2_decap_8 FILLER_40_173 ();
 sg13g2_fill_2 FILLER_40_180 ();
 sg13g2_fill_2 FILLER_40_190 ();
 sg13g2_fill_1 FILLER_40_192 ();
 sg13g2_decap_8 FILLER_40_210 ();
 sg13g2_fill_2 FILLER_40_217 ();
 sg13g2_fill_1 FILLER_40_219 ();
 sg13g2_fill_2 FILLER_40_230 ();
 sg13g2_fill_1 FILLER_40_232 ();
 sg13g2_fill_1 FILLER_40_238 ();
 sg13g2_decap_8 FILLER_40_247 ();
 sg13g2_decap_8 FILLER_40_258 ();
 sg13g2_decap_8 FILLER_40_265 ();
 sg13g2_fill_2 FILLER_40_272 ();
 sg13g2_fill_2 FILLER_40_296 ();
 sg13g2_fill_1 FILLER_40_306 ();
 sg13g2_decap_8 FILLER_40_312 ();
 sg13g2_decap_4 FILLER_40_319 ();
 sg13g2_fill_2 FILLER_40_323 ();
 sg13g2_fill_2 FILLER_40_329 ();
 sg13g2_fill_1 FILLER_40_331 ();
 sg13g2_decap_8 FILLER_40_342 ();
 sg13g2_decap_4 FILLER_40_349 ();
 sg13g2_decap_8 FILLER_40_357 ();
 sg13g2_decap_4 FILLER_40_364 ();
 sg13g2_fill_1 FILLER_40_368 ();
 sg13g2_decap_4 FILLER_40_402 ();
 sg13g2_fill_2 FILLER_40_406 ();
 sg13g2_fill_2 FILLER_40_418 ();
 sg13g2_fill_1 FILLER_40_420 ();
 sg13g2_decap_4 FILLER_40_426 ();
 sg13g2_fill_1 FILLER_40_430 ();
 sg13g2_decap_4 FILLER_40_440 ();
 sg13g2_fill_1 FILLER_40_444 ();
 sg13g2_decap_8 FILLER_40_458 ();
 sg13g2_decap_8 FILLER_40_465 ();
 sg13g2_decap_4 FILLER_40_472 ();
 sg13g2_fill_2 FILLER_40_476 ();
 sg13g2_fill_1 FILLER_40_482 ();
 sg13g2_decap_8 FILLER_40_495 ();
 sg13g2_fill_1 FILLER_40_502 ();
 sg13g2_fill_2 FILLER_40_516 ();
 sg13g2_fill_1 FILLER_40_518 ();
 sg13g2_decap_4 FILLER_40_523 ();
 sg13g2_decap_8 FILLER_40_531 ();
 sg13g2_fill_2 FILLER_40_538 ();
 sg13g2_fill_1 FILLER_40_540 ();
 sg13g2_decap_8 FILLER_40_545 ();
 sg13g2_decap_8 FILLER_40_552 ();
 sg13g2_decap_8 FILLER_40_559 ();
 sg13g2_decap_8 FILLER_40_566 ();
 sg13g2_decap_8 FILLER_40_573 ();
 sg13g2_fill_2 FILLER_40_580 ();
 sg13g2_decap_8 FILLER_40_590 ();
 sg13g2_decap_4 FILLER_40_597 ();
 sg13g2_fill_1 FILLER_40_601 ();
 sg13g2_decap_8 FILLER_40_606 ();
 sg13g2_fill_1 FILLER_40_631 ();
 sg13g2_fill_1 FILLER_40_647 ();
 sg13g2_fill_2 FILLER_40_653 ();
 sg13g2_fill_2 FILLER_40_675 ();
 sg13g2_fill_1 FILLER_40_686 ();
 sg13g2_decap_4 FILLER_40_696 ();
 sg13g2_decap_4 FILLER_40_705 ();
 sg13g2_fill_1 FILLER_40_709 ();
 sg13g2_decap_8 FILLER_40_717 ();
 sg13g2_decap_8 FILLER_40_724 ();
 sg13g2_fill_1 FILLER_40_731 ();
 sg13g2_decap_8 FILLER_40_738 ();
 sg13g2_fill_1 FILLER_40_745 ();
 sg13g2_decap_4 FILLER_40_751 ();
 sg13g2_fill_1 FILLER_40_755 ();
 sg13g2_decap_4 FILLER_40_765 ();
 sg13g2_fill_1 FILLER_40_779 ();
 sg13g2_fill_2 FILLER_40_784 ();
 sg13g2_decap_4 FILLER_40_790 ();
 sg13g2_fill_2 FILLER_40_794 ();
 sg13g2_decap_4 FILLER_40_801 ();
 sg13g2_fill_2 FILLER_40_819 ();
 sg13g2_fill_1 FILLER_40_821 ();
 sg13g2_fill_2 FILLER_40_837 ();
 sg13g2_fill_1 FILLER_40_839 ();
 sg13g2_decap_8 FILLER_40_844 ();
 sg13g2_decap_8 FILLER_40_851 ();
 sg13g2_decap_8 FILLER_40_858 ();
 sg13g2_decap_8 FILLER_40_865 ();
 sg13g2_decap_4 FILLER_40_872 ();
 sg13g2_fill_2 FILLER_40_876 ();
 sg13g2_decap_8 FILLER_41_0 ();
 sg13g2_decap_8 FILLER_41_7 ();
 sg13g2_decap_4 FILLER_41_14 ();
 sg13g2_fill_1 FILLER_41_18 ();
 sg13g2_decap_8 FILLER_41_28 ();
 sg13g2_decap_4 FILLER_41_35 ();
 sg13g2_fill_1 FILLER_41_39 ();
 sg13g2_fill_2 FILLER_41_66 ();
 sg13g2_fill_1 FILLER_41_68 ();
 sg13g2_decap_8 FILLER_41_72 ();
 sg13g2_decap_8 FILLER_41_79 ();
 sg13g2_fill_1 FILLER_41_86 ();
 sg13g2_fill_2 FILLER_41_97 ();
 sg13g2_fill_1 FILLER_41_99 ();
 sg13g2_fill_2 FILLER_41_110 ();
 sg13g2_fill_1 FILLER_41_112 ();
 sg13g2_decap_8 FILLER_41_117 ();
 sg13g2_fill_2 FILLER_41_124 ();
 sg13g2_fill_1 FILLER_41_126 ();
 sg13g2_decap_4 FILLER_41_131 ();
 sg13g2_fill_2 FILLER_41_135 ();
 sg13g2_decap_8 FILLER_41_142 ();
 sg13g2_fill_2 FILLER_41_159 ();
 sg13g2_fill_1 FILLER_41_161 ();
 sg13g2_fill_1 FILLER_41_167 ();
 sg13g2_decap_8 FILLER_41_173 ();
 sg13g2_decap_8 FILLER_41_180 ();
 sg13g2_decap_4 FILLER_41_187 ();
 sg13g2_fill_2 FILLER_41_191 ();
 sg13g2_decap_8 FILLER_41_208 ();
 sg13g2_decap_8 FILLER_41_215 ();
 sg13g2_fill_2 FILLER_41_222 ();
 sg13g2_decap_8 FILLER_41_239 ();
 sg13g2_decap_8 FILLER_41_246 ();
 sg13g2_decap_8 FILLER_41_253 ();
 sg13g2_decap_4 FILLER_41_260 ();
 sg13g2_fill_2 FILLER_41_264 ();
 sg13g2_decap_8 FILLER_41_270 ();
 sg13g2_fill_2 FILLER_41_277 ();
 sg13g2_fill_1 FILLER_41_279 ();
 sg13g2_fill_1 FILLER_41_283 ();
 sg13g2_decap_4 FILLER_41_287 ();
 sg13g2_fill_2 FILLER_41_291 ();
 sg13g2_decap_8 FILLER_41_298 ();
 sg13g2_decap_8 FILLER_41_305 ();
 sg13g2_fill_1 FILLER_41_312 ();
 sg13g2_decap_8 FILLER_41_322 ();
 sg13g2_fill_2 FILLER_41_329 ();
 sg13g2_fill_1 FILLER_41_331 ();
 sg13g2_decap_8 FILLER_41_342 ();
 sg13g2_fill_2 FILLER_41_349 ();
 sg13g2_fill_1 FILLER_41_351 ();
 sg13g2_fill_2 FILLER_41_382 ();
 sg13g2_decap_4 FILLER_41_388 ();
 sg13g2_decap_8 FILLER_41_397 ();
 sg13g2_decap_4 FILLER_41_404 ();
 sg13g2_fill_2 FILLER_41_408 ();
 sg13g2_decap_4 FILLER_41_414 ();
 sg13g2_fill_2 FILLER_41_418 ();
 sg13g2_fill_2 FILLER_41_424 ();
 sg13g2_fill_1 FILLER_41_426 ();
 sg13g2_fill_1 FILLER_41_431 ();
 sg13g2_fill_1 FILLER_41_437 ();
 sg13g2_fill_1 FILLER_41_445 ();
 sg13g2_fill_1 FILLER_41_451 ();
 sg13g2_decap_4 FILLER_41_462 ();
 sg13g2_decap_4 FILLER_41_482 ();
 sg13g2_fill_2 FILLER_41_486 ();
 sg13g2_fill_2 FILLER_41_492 ();
 sg13g2_decap_8 FILLER_41_523 ();
 sg13g2_decap_4 FILLER_41_530 ();
 sg13g2_fill_1 FILLER_41_534 ();
 sg13g2_decap_8 FILLER_41_540 ();
 sg13g2_decap_8 FILLER_41_547 ();
 sg13g2_decap_4 FILLER_41_554 ();
 sg13g2_fill_1 FILLER_41_558 ();
 sg13g2_fill_1 FILLER_41_571 ();
 sg13g2_decap_8 FILLER_41_598 ();
 sg13g2_decap_4 FILLER_41_638 ();
 sg13g2_fill_2 FILLER_41_642 ();
 sg13g2_fill_1 FILLER_41_649 ();
 sg13g2_decap_8 FILLER_41_655 ();
 sg13g2_fill_1 FILLER_41_662 ();
 sg13g2_decap_8 FILLER_41_668 ();
 sg13g2_decap_4 FILLER_41_675 ();
 sg13g2_fill_1 FILLER_41_679 ();
 sg13g2_decap_8 FILLER_41_689 ();
 sg13g2_fill_2 FILLER_41_696 ();
 sg13g2_fill_1 FILLER_41_698 ();
 sg13g2_decap_8 FILLER_41_703 ();
 sg13g2_decap_4 FILLER_41_710 ();
 sg13g2_fill_2 FILLER_41_718 ();
 sg13g2_decap_4 FILLER_41_743 ();
 sg13g2_fill_2 FILLER_41_747 ();
 sg13g2_fill_2 FILLER_41_776 ();
 sg13g2_decap_4 FILLER_41_782 ();
 sg13g2_fill_1 FILLER_41_797 ();
 sg13g2_decap_8 FILLER_41_814 ();
 sg13g2_decap_4 FILLER_41_821 ();
 sg13g2_fill_2 FILLER_41_825 ();
 sg13g2_decap_8 FILLER_41_840 ();
 sg13g2_decap_4 FILLER_41_847 ();
 sg13g2_fill_2 FILLER_41_851 ();
 sg13g2_decap_8 FILLER_41_857 ();
 sg13g2_decap_8 FILLER_41_864 ();
 sg13g2_decap_8 FILLER_41_871 ();
 sg13g2_fill_1 FILLER_42_0 ();
 sg13g2_decap_4 FILLER_42_32 ();
 sg13g2_fill_2 FILLER_42_41 ();
 sg13g2_fill_1 FILLER_42_43 ();
 sg13g2_fill_2 FILLER_42_48 ();
 sg13g2_fill_1 FILLER_42_50 ();
 sg13g2_decap_8 FILLER_42_55 ();
 sg13g2_fill_1 FILLER_42_67 ();
 sg13g2_decap_4 FILLER_42_77 ();
 sg13g2_fill_2 FILLER_42_81 ();
 sg13g2_fill_2 FILLER_42_91 ();
 sg13g2_fill_1 FILLER_42_93 ();
 sg13g2_decap_4 FILLER_42_100 ();
 sg13g2_fill_2 FILLER_42_104 ();
 sg13g2_fill_2 FILLER_42_132 ();
 sg13g2_fill_1 FILLER_42_134 ();
 sg13g2_fill_2 FILLER_42_140 ();
 sg13g2_fill_1 FILLER_42_158 ();
 sg13g2_fill_1 FILLER_42_167 ();
 sg13g2_decap_8 FILLER_42_178 ();
 sg13g2_fill_2 FILLER_42_193 ();
 sg13g2_decap_8 FILLER_42_208 ();
 sg13g2_decap_8 FILLER_42_215 ();
 sg13g2_fill_2 FILLER_42_222 ();
 sg13g2_fill_1 FILLER_42_224 ();
 sg13g2_decap_8 FILLER_42_245 ();
 sg13g2_decap_8 FILLER_42_252 ();
 sg13g2_fill_1 FILLER_42_259 ();
 sg13g2_decap_8 FILLER_42_290 ();
 sg13g2_decap_8 FILLER_42_297 ();
 sg13g2_fill_2 FILLER_42_304 ();
 sg13g2_fill_1 FILLER_42_306 ();
 sg13g2_decap_8 FILLER_42_310 ();
 sg13g2_fill_1 FILLER_42_317 ();
 sg13g2_decap_4 FILLER_42_323 ();
 sg13g2_decap_4 FILLER_42_334 ();
 sg13g2_fill_1 FILLER_42_338 ();
 sg13g2_fill_2 FILLER_42_359 ();
 sg13g2_fill_1 FILLER_42_361 ();
 sg13g2_fill_2 FILLER_42_376 ();
 sg13g2_fill_1 FILLER_42_378 ();
 sg13g2_decap_4 FILLER_42_384 ();
 sg13g2_fill_2 FILLER_42_392 ();
 sg13g2_fill_1 FILLER_42_394 ();
 sg13g2_decap_8 FILLER_42_414 ();
 sg13g2_decap_4 FILLER_42_431 ();
 sg13g2_decap_8 FILLER_42_439 ();
 sg13g2_decap_8 FILLER_42_446 ();
 sg13g2_decap_8 FILLER_42_453 ();
 sg13g2_decap_8 FILLER_42_460 ();
 sg13g2_decap_8 FILLER_42_467 ();
 sg13g2_fill_1 FILLER_42_474 ();
 sg13g2_fill_2 FILLER_42_488 ();
 sg13g2_decap_4 FILLER_42_517 ();
 sg13g2_decap_4 FILLER_42_527 ();
 sg13g2_fill_2 FILLER_42_535 ();
 sg13g2_decap_4 FILLER_42_554 ();
 sg13g2_fill_1 FILLER_42_558 ();
 sg13g2_decap_8 FILLER_42_564 ();
 sg13g2_decap_8 FILLER_42_571 ();
 sg13g2_fill_1 FILLER_42_578 ();
 sg13g2_fill_1 FILLER_42_606 ();
 sg13g2_fill_1 FILLER_42_611 ();
 sg13g2_decap_8 FILLER_42_621 ();
 sg13g2_fill_1 FILLER_42_628 ();
 sg13g2_fill_2 FILLER_42_634 ();
 sg13g2_fill_1 FILLER_42_636 ();
 sg13g2_decap_4 FILLER_42_658 ();
 sg13g2_fill_1 FILLER_42_662 ();
 sg13g2_fill_2 FILLER_42_667 ();
 sg13g2_fill_1 FILLER_42_669 ();
 sg13g2_fill_2 FILLER_42_691 ();
 sg13g2_fill_2 FILLER_42_698 ();
 sg13g2_fill_1 FILLER_42_700 ();
 sg13g2_fill_2 FILLER_42_719 ();
 sg13g2_decap_8 FILLER_42_730 ();
 sg13g2_decap_8 FILLER_42_740 ();
 sg13g2_fill_1 FILLER_42_762 ();
 sg13g2_fill_1 FILLER_42_768 ();
 sg13g2_fill_2 FILLER_42_789 ();
 sg13g2_fill_1 FILLER_42_791 ();
 sg13g2_fill_2 FILLER_42_801 ();
 sg13g2_decap_8 FILLER_42_808 ();
 sg13g2_decap_8 FILLER_42_815 ();
 sg13g2_decap_8 FILLER_42_822 ();
 sg13g2_decap_8 FILLER_42_829 ();
 sg13g2_fill_1 FILLER_42_836 ();
 sg13g2_decap_4 FILLER_42_842 ();
 sg13g2_fill_1 FILLER_42_846 ();
 sg13g2_decap_4 FILLER_42_873 ();
 sg13g2_fill_1 FILLER_42_877 ();
 sg13g2_decap_8 FILLER_43_0 ();
 sg13g2_decap_4 FILLER_43_7 ();
 sg13g2_decap_4 FILLER_43_15 ();
 sg13g2_fill_2 FILLER_43_19 ();
 sg13g2_fill_2 FILLER_43_25 ();
 sg13g2_fill_1 FILLER_43_27 ();
 sg13g2_fill_2 FILLER_43_66 ();
 sg13g2_fill_2 FILLER_43_76 ();
 sg13g2_decap_4 FILLER_43_84 ();
 sg13g2_fill_2 FILLER_43_88 ();
 sg13g2_decap_8 FILLER_43_95 ();
 sg13g2_decap_4 FILLER_43_102 ();
 sg13g2_fill_1 FILLER_43_106 ();
 sg13g2_decap_8 FILLER_43_116 ();
 sg13g2_decap_4 FILLER_43_123 ();
 sg13g2_decap_8 FILLER_43_132 ();
 sg13g2_fill_2 FILLER_43_139 ();
 sg13g2_decap_4 FILLER_43_163 ();
 sg13g2_fill_1 FILLER_43_167 ();
 sg13g2_decap_8 FILLER_43_176 ();
 sg13g2_decap_8 FILLER_43_183 ();
 sg13g2_decap_4 FILLER_43_195 ();
 sg13g2_decap_8 FILLER_43_215 ();
 sg13g2_decap_4 FILLER_43_222 ();
 sg13g2_decap_8 FILLER_43_253 ();
 sg13g2_decap_4 FILLER_43_260 ();
 sg13g2_fill_1 FILLER_43_264 ();
 sg13g2_decap_8 FILLER_43_270 ();
 sg13g2_decap_8 FILLER_43_277 ();
 sg13g2_fill_2 FILLER_43_284 ();
 sg13g2_decap_4 FILLER_43_290 ();
 sg13g2_decap_8 FILLER_43_307 ();
 sg13g2_decap_4 FILLER_43_314 ();
 sg13g2_fill_2 FILLER_43_318 ();
 sg13g2_decap_8 FILLER_43_335 ();
 sg13g2_fill_2 FILLER_43_342 ();
 sg13g2_fill_2 FILLER_43_354 ();
 sg13g2_fill_1 FILLER_43_356 ();
 sg13g2_decap_4 FILLER_43_377 ();
 sg13g2_fill_1 FILLER_43_416 ();
 sg13g2_decap_8 FILLER_43_420 ();
 sg13g2_decap_8 FILLER_43_427 ();
 sg13g2_decap_8 FILLER_43_434 ();
 sg13g2_decap_8 FILLER_43_441 ();
 sg13g2_decap_8 FILLER_43_448 ();
 sg13g2_decap_8 FILLER_43_455 ();
 sg13g2_decap_8 FILLER_43_462 ();
 sg13g2_decap_8 FILLER_43_469 ();
 sg13g2_fill_1 FILLER_43_476 ();
 sg13g2_fill_1 FILLER_43_490 ();
 sg13g2_fill_1 FILLER_43_494 ();
 sg13g2_fill_1 FILLER_43_505 ();
 sg13g2_fill_1 FILLER_43_511 ();
 sg13g2_fill_2 FILLER_43_519 ();
 sg13g2_decap_4 FILLER_43_526 ();
 sg13g2_decap_8 FILLER_43_540 ();
 sg13g2_decap_8 FILLER_43_547 ();
 sg13g2_decap_8 FILLER_43_554 ();
 sg13g2_decap_8 FILLER_43_561 ();
 sg13g2_fill_2 FILLER_43_568 ();
 sg13g2_fill_2 FILLER_43_575 ();
 sg13g2_fill_1 FILLER_43_581 ();
 sg13g2_decap_4 FILLER_43_617 ();
 sg13g2_decap_4 FILLER_43_625 ();
 sg13g2_fill_1 FILLER_43_629 ();
 sg13g2_fill_2 FILLER_43_643 ();
 sg13g2_fill_1 FILLER_43_645 ();
 sg13g2_decap_8 FILLER_43_650 ();
 sg13g2_decap_4 FILLER_43_657 ();
 sg13g2_fill_2 FILLER_43_661 ();
 sg13g2_fill_2 FILLER_43_685 ();
 sg13g2_fill_1 FILLER_43_699 ();
 sg13g2_fill_2 FILLER_43_713 ();
 sg13g2_fill_1 FILLER_43_720 ();
 sg13g2_decap_8 FILLER_43_742 ();
 sg13g2_decap_4 FILLER_43_749 ();
 sg13g2_decap_8 FILLER_43_774 ();
 sg13g2_fill_1 FILLER_43_781 ();
 sg13g2_decap_4 FILLER_43_801 ();
 sg13g2_fill_1 FILLER_43_810 ();
 sg13g2_decap_4 FILLER_43_835 ();
 sg13g2_decap_8 FILLER_43_852 ();
 sg13g2_fill_1 FILLER_43_859 ();
 sg13g2_decap_8 FILLER_43_865 ();
 sg13g2_decap_4 FILLER_43_872 ();
 sg13g2_fill_2 FILLER_43_876 ();
 sg13g2_decap_8 FILLER_44_0 ();
 sg13g2_decap_8 FILLER_44_11 ();
 sg13g2_decap_4 FILLER_44_23 ();
 sg13g2_decap_4 FILLER_44_32 ();
 sg13g2_fill_1 FILLER_44_36 ();
 sg13g2_decap_4 FILLER_44_44 ();
 sg13g2_fill_2 FILLER_44_48 ();
 sg13g2_decap_8 FILLER_44_53 ();
 sg13g2_decap_8 FILLER_44_60 ();
 sg13g2_decap_8 FILLER_44_67 ();
 sg13g2_fill_2 FILLER_44_74 ();
 sg13g2_fill_2 FILLER_44_85 ();
 sg13g2_decap_4 FILLER_44_121 ();
 sg13g2_fill_2 FILLER_44_125 ();
 sg13g2_decap_8 FILLER_44_135 ();
 sg13g2_decap_8 FILLER_44_142 ();
 sg13g2_decap_8 FILLER_44_157 ();
 sg13g2_decap_8 FILLER_44_164 ();
 sg13g2_decap_8 FILLER_44_171 ();
 sg13g2_decap_4 FILLER_44_178 ();
 sg13g2_fill_2 FILLER_44_191 ();
 sg13g2_fill_1 FILLER_44_193 ();
 sg13g2_decap_8 FILLER_44_214 ();
 sg13g2_decap_8 FILLER_44_221 ();
 sg13g2_fill_2 FILLER_44_228 ();
 sg13g2_decap_4 FILLER_44_240 ();
 sg13g2_fill_1 FILLER_44_244 ();
 sg13g2_fill_1 FILLER_44_253 ();
 sg13g2_decap_4 FILLER_44_275 ();
 sg13g2_fill_1 FILLER_44_279 ();
 sg13g2_decap_8 FILLER_44_285 ();
 sg13g2_decap_8 FILLER_44_311 ();
 sg13g2_decap_8 FILLER_44_318 ();
 sg13g2_decap_8 FILLER_44_325 ();
 sg13g2_decap_8 FILLER_44_332 ();
 sg13g2_decap_8 FILLER_44_339 ();
 sg13g2_decap_8 FILLER_44_346 ();
 sg13g2_decap_4 FILLER_44_353 ();
 sg13g2_fill_2 FILLER_44_367 ();
 sg13g2_decap_4 FILLER_44_377 ();
 sg13g2_fill_2 FILLER_44_381 ();
 sg13g2_fill_1 FILLER_44_403 ();
 sg13g2_decap_8 FILLER_44_413 ();
 sg13g2_decap_8 FILLER_44_420 ();
 sg13g2_decap_8 FILLER_44_427 ();
 sg13g2_decap_8 FILLER_44_434 ();
 sg13g2_fill_1 FILLER_44_441 ();
 sg13g2_decap_8 FILLER_44_457 ();
 sg13g2_decap_4 FILLER_44_464 ();
 sg13g2_fill_2 FILLER_44_468 ();
 sg13g2_fill_1 FILLER_44_475 ();
 sg13g2_fill_2 FILLER_44_510 ();
 sg13g2_fill_2 FILLER_44_517 ();
 sg13g2_decap_8 FILLER_44_527 ();
 sg13g2_decap_8 FILLER_44_538 ();
 sg13g2_decap_4 FILLER_44_545 ();
 sg13g2_fill_1 FILLER_44_549 ();
 sg13g2_decap_8 FILLER_44_555 ();
 sg13g2_decap_8 FILLER_44_562 ();
 sg13g2_decap_8 FILLER_44_569 ();
 sg13g2_fill_2 FILLER_44_576 ();
 sg13g2_fill_1 FILLER_44_585 ();
 sg13g2_decap_4 FILLER_44_596 ();
 sg13g2_fill_2 FILLER_44_625 ();
 sg13g2_decap_8 FILLER_44_645 ();
 sg13g2_fill_1 FILLER_44_656 ();
 sg13g2_decap_4 FILLER_44_666 ();
 sg13g2_fill_1 FILLER_44_670 ();
 sg13g2_fill_2 FILLER_44_705 ();
 sg13g2_decap_4 FILLER_44_714 ();
 sg13g2_fill_2 FILLER_44_723 ();
 sg13g2_fill_1 FILLER_44_725 ();
 sg13g2_decap_8 FILLER_44_749 ();
 sg13g2_decap_8 FILLER_44_761 ();
 sg13g2_decap_4 FILLER_44_768 ();
 sg13g2_fill_1 FILLER_44_780 ();
 sg13g2_fill_2 FILLER_44_790 ();
 sg13g2_fill_2 FILLER_44_796 ();
 sg13g2_fill_1 FILLER_44_798 ();
 sg13g2_decap_8 FILLER_44_803 ();
 sg13g2_decap_8 FILLER_44_810 ();
 sg13g2_fill_2 FILLER_44_817 ();
 sg13g2_fill_1 FILLER_44_824 ();
 sg13g2_fill_1 FILLER_44_830 ();
 sg13g2_decap_4 FILLER_44_836 ();
 sg13g2_fill_2 FILLER_44_845 ();
 sg13g2_fill_1 FILLER_44_847 ();
 sg13g2_decap_8 FILLER_44_853 ();
 sg13g2_decap_8 FILLER_44_860 ();
 sg13g2_decap_8 FILLER_44_867 ();
 sg13g2_decap_4 FILLER_44_874 ();
 sg13g2_fill_2 FILLER_45_26 ();
 sg13g2_fill_2 FILLER_45_32 ();
 sg13g2_fill_2 FILLER_45_52 ();
 sg13g2_fill_1 FILLER_45_82 ();
 sg13g2_decap_8 FILLER_45_87 ();
 sg13g2_decap_8 FILLER_45_94 ();
 sg13g2_decap_8 FILLER_45_101 ();
 sg13g2_decap_8 FILLER_45_108 ();
 sg13g2_decap_8 FILLER_45_115 ();
 sg13g2_decap_8 FILLER_45_122 ();
 sg13g2_decap_8 FILLER_45_134 ();
 sg13g2_decap_4 FILLER_45_141 ();
 sg13g2_decap_8 FILLER_45_157 ();
 sg13g2_fill_1 FILLER_45_164 ();
 sg13g2_decap_4 FILLER_45_173 ();
 sg13g2_fill_1 FILLER_45_177 ();
 sg13g2_decap_8 FILLER_45_188 ();
 sg13g2_decap_8 FILLER_45_195 ();
 sg13g2_fill_2 FILLER_45_202 ();
 sg13g2_decap_8 FILLER_45_214 ();
 sg13g2_decap_8 FILLER_45_221 ();
 sg13g2_fill_1 FILLER_45_228 ();
 sg13g2_fill_2 FILLER_45_233 ();
 sg13g2_fill_1 FILLER_45_235 ();
 sg13g2_decap_8 FILLER_45_241 ();
 sg13g2_decap_8 FILLER_45_248 ();
 sg13g2_fill_1 FILLER_45_259 ();
 sg13g2_fill_2 FILLER_45_269 ();
 sg13g2_decap_4 FILLER_45_275 ();
 sg13g2_decap_8 FILLER_45_283 ();
 sg13g2_decap_8 FILLER_45_290 ();
 sg13g2_decap_8 FILLER_45_297 ();
 sg13g2_decap_8 FILLER_45_304 ();
 sg13g2_fill_2 FILLER_45_311 ();
 sg13g2_decap_8 FILLER_45_317 ();
 sg13g2_fill_2 FILLER_45_324 ();
 sg13g2_fill_1 FILLER_45_326 ();
 sg13g2_decap_8 FILLER_45_332 ();
 sg13g2_fill_1 FILLER_45_339 ();
 sg13g2_decap_4 FILLER_45_345 ();
 sg13g2_fill_1 FILLER_45_349 ();
 sg13g2_decap_4 FILLER_45_354 ();
 sg13g2_decap_4 FILLER_45_364 ();
 sg13g2_fill_1 FILLER_45_368 ();
 sg13g2_decap_4 FILLER_45_374 ();
 sg13g2_fill_1 FILLER_45_378 ();
 sg13g2_fill_1 FILLER_45_383 ();
 sg13g2_fill_2 FILLER_45_393 ();
 sg13g2_decap_8 FILLER_45_400 ();
 sg13g2_decap_8 FILLER_45_407 ();
 sg13g2_fill_2 FILLER_45_414 ();
 sg13g2_decap_8 FILLER_45_422 ();
 sg13g2_decap_4 FILLER_45_429 ();
 sg13g2_decap_8 FILLER_45_453 ();
 sg13g2_decap_8 FILLER_45_460 ();
 sg13g2_decap_4 FILLER_45_480 ();
 sg13g2_fill_2 FILLER_45_488 ();
 sg13g2_fill_1 FILLER_45_490 ();
 sg13g2_fill_1 FILLER_45_495 ();
 sg13g2_fill_2 FILLER_45_502 ();
 sg13g2_decap_8 FILLER_45_513 ();
 sg13g2_decap_8 FILLER_45_520 ();
 sg13g2_decap_4 FILLER_45_527 ();
 sg13g2_fill_1 FILLER_45_531 ();
 sg13g2_fill_1 FILLER_45_536 ();
 sg13g2_decap_8 FILLER_45_540 ();
 sg13g2_fill_1 FILLER_45_547 ();
 sg13g2_decap_4 FILLER_45_552 ();
 sg13g2_fill_2 FILLER_45_556 ();
 sg13g2_decap_8 FILLER_45_574 ();
 sg13g2_fill_2 FILLER_45_581 ();
 sg13g2_fill_2 FILLER_45_595 ();
 sg13g2_fill_1 FILLER_45_597 ();
 sg13g2_fill_1 FILLER_45_608 ();
 sg13g2_fill_2 FILLER_45_614 ();
 sg13g2_fill_1 FILLER_45_625 ();
 sg13g2_fill_2 FILLER_45_633 ();
 sg13g2_fill_1 FILLER_45_635 ();
 sg13g2_decap_8 FILLER_45_640 ();
 sg13g2_fill_1 FILLER_45_647 ();
 sg13g2_fill_1 FILLER_45_653 ();
 sg13g2_decap_8 FILLER_45_658 ();
 sg13g2_decap_8 FILLER_45_665 ();
 sg13g2_decap_8 FILLER_45_691 ();
 sg13g2_decap_4 FILLER_45_698 ();
 sg13g2_fill_1 FILLER_45_706 ();
 sg13g2_fill_2 FILLER_45_720 ();
 sg13g2_decap_4 FILLER_45_734 ();
 sg13g2_fill_1 FILLER_45_738 ();
 sg13g2_decap_4 FILLER_45_743 ();
 sg13g2_fill_2 FILLER_45_752 ();
 sg13g2_fill_2 FILLER_45_772 ();
 sg13g2_fill_1 FILLER_45_774 ();
 sg13g2_decap_4 FILLER_45_785 ();
 sg13g2_decap_4 FILLER_45_793 ();
 sg13g2_fill_1 FILLER_45_797 ();
 sg13g2_decap_4 FILLER_45_802 ();
 sg13g2_fill_2 FILLER_45_815 ();
 sg13g2_fill_1 FILLER_45_833 ();
 sg13g2_fill_1 FILLER_45_847 ();
 sg13g2_decap_8 FILLER_45_853 ();
 sg13g2_decap_8 FILLER_45_860 ();
 sg13g2_decap_8 FILLER_45_867 ();
 sg13g2_decap_4 FILLER_45_874 ();
 sg13g2_decap_8 FILLER_46_0 ();
 sg13g2_decap_8 FILLER_46_7 ();
 sg13g2_decap_8 FILLER_46_47 ();
 sg13g2_decap_8 FILLER_46_54 ();
 sg13g2_decap_8 FILLER_46_61 ();
 sg13g2_decap_4 FILLER_46_68 ();
 sg13g2_fill_1 FILLER_46_72 ();
 sg13g2_decap_8 FILLER_46_78 ();
 sg13g2_fill_1 FILLER_46_85 ();
 sg13g2_decap_8 FILLER_46_97 ();
 sg13g2_fill_2 FILLER_46_104 ();
 sg13g2_decap_8 FILLER_46_118 ();
 sg13g2_decap_8 FILLER_46_125 ();
 sg13g2_fill_1 FILLER_46_132 ();
 sg13g2_fill_2 FILLER_46_141 ();
 sg13g2_fill_1 FILLER_46_143 ();
 sg13g2_decap_8 FILLER_46_156 ();
 sg13g2_decap_4 FILLER_46_163 ();
 sg13g2_fill_1 FILLER_46_167 ();
 sg13g2_decap_8 FILLER_46_176 ();
 sg13g2_decap_4 FILLER_46_183 ();
 sg13g2_fill_2 FILLER_46_206 ();
 sg13g2_decap_8 FILLER_46_213 ();
 sg13g2_decap_8 FILLER_46_224 ();
 sg13g2_decap_4 FILLER_46_231 ();
 sg13g2_fill_2 FILLER_46_235 ();
 sg13g2_decap_8 FILLER_46_242 ();
 sg13g2_fill_2 FILLER_46_249 ();
 sg13g2_fill_2 FILLER_46_270 ();
 sg13g2_fill_1 FILLER_46_272 ();
 sg13g2_fill_2 FILLER_46_304 ();
 sg13g2_fill_1 FILLER_46_306 ();
 sg13g2_fill_2 FILLER_46_341 ();
 sg13g2_fill_2 FILLER_46_347 ();
 sg13g2_decap_8 FILLER_46_354 ();
 sg13g2_decap_4 FILLER_46_361 ();
 sg13g2_fill_2 FILLER_46_381 ();
 sg13g2_fill_1 FILLER_46_383 ();
 sg13g2_fill_2 FILLER_46_389 ();
 sg13g2_fill_2 FILLER_46_395 ();
 sg13g2_decap_8 FILLER_46_400 ();
 sg13g2_fill_1 FILLER_46_407 ();
 sg13g2_decap_8 FILLER_46_450 ();
 sg13g2_decap_8 FILLER_46_471 ();
 sg13g2_decap_4 FILLER_46_478 ();
 sg13g2_decap_8 FILLER_46_514 ();
 sg13g2_decap_4 FILLER_46_521 ();
 sg13g2_decap_8 FILLER_46_551 ();
 sg13g2_decap_4 FILLER_46_558 ();
 sg13g2_fill_1 FILLER_46_562 ();
 sg13g2_decap_8 FILLER_46_567 ();
 sg13g2_decap_4 FILLER_46_574 ();
 sg13g2_decap_8 FILLER_46_583 ();
 sg13g2_fill_1 FILLER_46_590 ();
 sg13g2_decap_4 FILLER_46_599 ();
 sg13g2_fill_2 FILLER_46_603 ();
 sg13g2_fill_2 FILLER_46_620 ();
 sg13g2_fill_1 FILLER_46_622 ();
 sg13g2_fill_2 FILLER_46_641 ();
 sg13g2_fill_1 FILLER_46_643 ();
 sg13g2_fill_2 FILLER_46_653 ();
 sg13g2_fill_1 FILLER_46_655 ();
 sg13g2_decap_4 FILLER_46_666 ();
 sg13g2_fill_2 FILLER_46_670 ();
 sg13g2_decap_8 FILLER_46_688 ();
 sg13g2_decap_4 FILLER_46_695 ();
 sg13g2_fill_2 FILLER_46_699 ();
 sg13g2_fill_2 FILLER_46_706 ();
 sg13g2_fill_1 FILLER_46_708 ();
 sg13g2_fill_2 FILLER_46_714 ();
 sg13g2_fill_1 FILLER_46_716 ();
 sg13g2_decap_8 FILLER_46_740 ();
 sg13g2_fill_1 FILLER_46_747 ();
 sg13g2_fill_2 FILLER_46_763 ();
 sg13g2_fill_1 FILLER_46_769 ();
 sg13g2_fill_1 FILLER_46_780 ();
 sg13g2_fill_1 FILLER_46_786 ();
 sg13g2_decap_8 FILLER_46_792 ();
 sg13g2_decap_8 FILLER_46_819 ();
 sg13g2_decap_4 FILLER_46_826 ();
 sg13g2_fill_1 FILLER_46_830 ();
 sg13g2_fill_2 FILLER_46_836 ();
 sg13g2_decap_8 FILLER_46_852 ();
 sg13g2_decap_8 FILLER_46_859 ();
 sg13g2_decap_8 FILLER_46_866 ();
 sg13g2_decap_4 FILLER_46_873 ();
 sg13g2_fill_1 FILLER_46_877 ();
 sg13g2_decap_8 FILLER_47_0 ();
 sg13g2_decap_8 FILLER_47_7 ();
 sg13g2_fill_2 FILLER_47_14 ();
 sg13g2_fill_1 FILLER_47_16 ();
 sg13g2_fill_1 FILLER_47_27 ();
 sg13g2_fill_1 FILLER_47_40 ();
 sg13g2_fill_1 FILLER_47_49 ();
 sg13g2_decap_8 FILLER_47_59 ();
 sg13g2_fill_2 FILLER_47_66 ();
 sg13g2_fill_2 FILLER_47_77 ();
 sg13g2_fill_1 FILLER_47_79 ();
 sg13g2_fill_1 FILLER_47_84 ();
 sg13g2_fill_2 FILLER_47_96 ();
 sg13g2_fill_2 FILLER_47_107 ();
 sg13g2_fill_1 FILLER_47_109 ();
 sg13g2_decap_4 FILLER_47_120 ();
 sg13g2_decap_4 FILLER_47_137 ();
 sg13g2_decap_8 FILLER_47_157 ();
 sg13g2_fill_2 FILLER_47_164 ();
 sg13g2_fill_1 FILLER_47_166 ();
 sg13g2_decap_4 FILLER_47_193 ();
 sg13g2_fill_1 FILLER_47_197 ();
 sg13g2_decap_4 FILLER_47_202 ();
 sg13g2_fill_2 FILLER_47_206 ();
 sg13g2_decap_4 FILLER_47_212 ();
 sg13g2_decap_8 FILLER_47_251 ();
 sg13g2_decap_8 FILLER_47_269 ();
 sg13g2_fill_2 FILLER_47_276 ();
 sg13g2_fill_1 FILLER_47_281 ();
 sg13g2_decap_8 FILLER_47_287 ();
 sg13g2_fill_2 FILLER_47_294 ();
 sg13g2_fill_1 FILLER_47_296 ();
 sg13g2_decap_4 FILLER_47_306 ();
 sg13g2_fill_2 FILLER_47_310 ();
 sg13g2_decap_8 FILLER_47_316 ();
 sg13g2_decap_4 FILLER_47_323 ();
 sg13g2_fill_2 FILLER_47_335 ();
 sg13g2_fill_1 FILLER_47_337 ();
 sg13g2_fill_2 FILLER_47_354 ();
 sg13g2_fill_2 FILLER_47_364 ();
 sg13g2_fill_1 FILLER_47_366 ();
 sg13g2_fill_2 FILLER_47_371 ();
 sg13g2_fill_2 FILLER_47_377 ();
 sg13g2_fill_1 FILLER_47_379 ();
 sg13g2_decap_4 FILLER_47_390 ();
 sg13g2_decap_8 FILLER_47_397 ();
 sg13g2_decap_8 FILLER_47_404 ();
 sg13g2_fill_1 FILLER_47_411 ();
 sg13g2_decap_8 FILLER_47_426 ();
 sg13g2_decap_8 FILLER_47_451 ();
 sg13g2_decap_8 FILLER_47_458 ();
 sg13g2_decap_8 FILLER_47_465 ();
 sg13g2_decap_8 FILLER_47_472 ();
 sg13g2_fill_2 FILLER_47_479 ();
 sg13g2_fill_2 FILLER_47_506 ();
 sg13g2_fill_2 FILLER_47_516 ();
 sg13g2_decap_8 FILLER_47_542 ();
 sg13g2_decap_8 FILLER_47_549 ();
 sg13g2_fill_2 FILLER_47_556 ();
 sg13g2_fill_1 FILLER_47_558 ();
 sg13g2_decap_4 FILLER_47_568 ();
 sg13g2_fill_1 FILLER_47_572 ();
 sg13g2_decap_4 FILLER_47_588 ();
 sg13g2_fill_2 FILLER_47_592 ();
 sg13g2_fill_2 FILLER_47_597 ();
 sg13g2_fill_1 FILLER_47_599 ();
 sg13g2_fill_2 FILLER_47_605 ();
 sg13g2_fill_2 FILLER_47_613 ();
 sg13g2_fill_2 FILLER_47_620 ();
 sg13g2_decap_4 FILLER_47_627 ();
 sg13g2_fill_1 FILLER_47_636 ();
 sg13g2_fill_2 FILLER_47_642 ();
 sg13g2_fill_1 FILLER_47_644 ();
 sg13g2_fill_2 FILLER_47_655 ();
 sg13g2_fill_1 FILLER_47_657 ();
 sg13g2_decap_8 FILLER_47_663 ();
 sg13g2_fill_1 FILLER_47_670 ();
 sg13g2_decap_4 FILLER_47_677 ();
 sg13g2_fill_2 FILLER_47_681 ();
 sg13g2_fill_1 FILLER_47_695 ();
 sg13g2_decap_8 FILLER_47_725 ();
 sg13g2_fill_1 FILLER_47_737 ();
 sg13g2_decap_8 FILLER_47_743 ();
 sg13g2_decap_4 FILLER_47_750 ();
 sg13g2_fill_1 FILLER_47_754 ();
 sg13g2_decap_8 FILLER_47_760 ();
 sg13g2_fill_2 FILLER_47_767 ();
 sg13g2_decap_4 FILLER_47_786 ();
 sg13g2_decap_4 FILLER_47_815 ();
 sg13g2_fill_1 FILLER_47_829 ();
 sg13g2_fill_2 FILLER_47_838 ();
 sg13g2_fill_1 FILLER_47_840 ();
 sg13g2_decap_8 FILLER_47_849 ();
 sg13g2_decap_8 FILLER_47_856 ();
 sg13g2_decap_8 FILLER_47_863 ();
 sg13g2_decap_8 FILLER_47_870 ();
 sg13g2_fill_1 FILLER_47_877 ();
 sg13g2_decap_8 FILLER_48_0 ();
 sg13g2_decap_8 FILLER_48_7 ();
 sg13g2_decap_8 FILLER_48_14 ();
 sg13g2_decap_8 FILLER_48_21 ();
 sg13g2_decap_8 FILLER_48_28 ();
 sg13g2_decap_8 FILLER_48_35 ();
 sg13g2_decap_4 FILLER_48_42 ();
 sg13g2_fill_2 FILLER_48_49 ();
 sg13g2_decap_8 FILLER_48_66 ();
 sg13g2_fill_1 FILLER_48_73 ();
 sg13g2_decap_8 FILLER_48_90 ();
 sg13g2_decap_4 FILLER_48_97 ();
 sg13g2_decap_8 FILLER_48_105 ();
 sg13g2_decap_8 FILLER_48_112 ();
 sg13g2_decap_8 FILLER_48_119 ();
 sg13g2_decap_8 FILLER_48_126 ();
 sg13g2_decap_8 FILLER_48_133 ();
 sg13g2_fill_2 FILLER_48_140 ();
 sg13g2_decap_8 FILLER_48_156 ();
 sg13g2_decap_8 FILLER_48_163 ();
 sg13g2_fill_1 FILLER_48_170 ();
 sg13g2_fill_2 FILLER_48_230 ();
 sg13g2_decap_8 FILLER_48_244 ();
 sg13g2_fill_2 FILLER_48_251 ();
 sg13g2_fill_1 FILLER_48_253 ();
 sg13g2_fill_1 FILLER_48_292 ();
 sg13g2_decap_4 FILLER_48_319 ();
 sg13g2_fill_2 FILLER_48_323 ();
 sg13g2_decap_8 FILLER_48_329 ();
 sg13g2_fill_1 FILLER_48_336 ();
 sg13g2_fill_1 FILLER_48_350 ();
 sg13g2_fill_2 FILLER_48_381 ();
 sg13g2_fill_1 FILLER_48_383 ();
 sg13g2_fill_1 FILLER_48_388 ();
 sg13g2_fill_2 FILLER_48_402 ();
 sg13g2_fill_1 FILLER_48_409 ();
 sg13g2_decap_8 FILLER_48_414 ();
 sg13g2_decap_4 FILLER_48_450 ();
 sg13g2_fill_2 FILLER_48_454 ();
 sg13g2_fill_2 FILLER_48_465 ();
 sg13g2_decap_4 FILLER_48_477 ();
 sg13g2_decap_8 FILLER_48_498 ();
 sg13g2_fill_2 FILLER_48_505 ();
 sg13g2_fill_1 FILLER_48_507 ();
 sg13g2_fill_1 FILLER_48_518 ();
 sg13g2_fill_1 FILLER_48_525 ();
 sg13g2_decap_8 FILLER_48_535 ();
 sg13g2_decap_4 FILLER_48_542 ();
 sg13g2_fill_1 FILLER_48_546 ();
 sg13g2_decap_8 FILLER_48_552 ();
 sg13g2_decap_4 FILLER_48_559 ();
 sg13g2_fill_1 FILLER_48_563 ();
 sg13g2_fill_1 FILLER_48_580 ();
 sg13g2_decap_8 FILLER_48_595 ();
 sg13g2_fill_1 FILLER_48_602 ();
 sg13g2_decap_4 FILLER_48_613 ();
 sg13g2_fill_1 FILLER_48_617 ();
 sg13g2_fill_1 FILLER_48_622 ();
 sg13g2_decap_4 FILLER_48_628 ();
 sg13g2_decap_8 FILLER_48_642 ();
 sg13g2_decap_8 FILLER_48_649 ();
 sg13g2_decap_8 FILLER_48_672 ();
 sg13g2_fill_2 FILLER_48_679 ();
 sg13g2_fill_1 FILLER_48_681 ();
 sg13g2_fill_2 FILLER_48_688 ();
 sg13g2_decap_4 FILLER_48_705 ();
 sg13g2_fill_2 FILLER_48_723 ();
 sg13g2_fill_1 FILLER_48_747 ();
 sg13g2_decap_8 FILLER_48_756 ();
 sg13g2_decap_8 FILLER_48_763 ();
 sg13g2_fill_2 FILLER_48_770 ();
 sg13g2_fill_1 FILLER_48_772 ();
 sg13g2_fill_1 FILLER_48_784 ();
 sg13g2_fill_2 FILLER_48_789 ();
 sg13g2_fill_2 FILLER_48_797 ();
 sg13g2_fill_1 FILLER_48_799 ();
 sg13g2_fill_2 FILLER_48_806 ();
 sg13g2_fill_1 FILLER_48_808 ();
 sg13g2_decap_8 FILLER_48_813 ();
 sg13g2_decap_8 FILLER_48_835 ();
 sg13g2_fill_2 FILLER_48_842 ();
 sg13g2_fill_1 FILLER_48_844 ();
 sg13g2_decap_8 FILLER_48_849 ();
 sg13g2_decap_8 FILLER_48_856 ();
 sg13g2_decap_8 FILLER_48_863 ();
 sg13g2_decap_8 FILLER_48_870 ();
 sg13g2_fill_1 FILLER_48_877 ();
 sg13g2_decap_8 FILLER_49_0 ();
 sg13g2_decap_8 FILLER_49_7 ();
 sg13g2_decap_4 FILLER_49_14 ();
 sg13g2_decap_8 FILLER_49_23 ();
 sg13g2_decap_8 FILLER_49_30 ();
 sg13g2_decap_4 FILLER_49_42 ();
 sg13g2_fill_2 FILLER_49_46 ();
 sg13g2_fill_2 FILLER_49_52 ();
 sg13g2_decap_8 FILLER_49_58 ();
 sg13g2_fill_2 FILLER_49_65 ();
 sg13g2_fill_1 FILLER_49_67 ();
 sg13g2_decap_8 FILLER_49_76 ();
 sg13g2_fill_2 FILLER_49_106 ();
 sg13g2_fill_1 FILLER_49_108 ();
 sg13g2_fill_1 FILLER_49_121 ();
 sg13g2_fill_1 FILLER_49_130 ();
 sg13g2_decap_4 FILLER_49_135 ();
 sg13g2_fill_2 FILLER_49_139 ();
 sg13g2_decap_8 FILLER_49_153 ();
 sg13g2_decap_8 FILLER_49_160 ();
 sg13g2_fill_2 FILLER_49_167 ();
 sg13g2_decap_4 FILLER_49_177 ();
 sg13g2_decap_8 FILLER_49_185 ();
 sg13g2_decap_8 FILLER_49_192 ();
 sg13g2_decap_8 FILLER_49_199 ();
 sg13g2_decap_8 FILLER_49_206 ();
 sg13g2_decap_4 FILLER_49_213 ();
 sg13g2_decap_8 FILLER_49_221 ();
 sg13g2_fill_2 FILLER_49_228 ();
 sg13g2_decap_8 FILLER_49_243 ();
 sg13g2_decap_8 FILLER_49_250 ();
 sg13g2_decap_4 FILLER_49_257 ();
 sg13g2_decap_8 FILLER_49_277 ();
 sg13g2_decap_4 FILLER_49_292 ();
 sg13g2_fill_2 FILLER_49_300 ();
 sg13g2_fill_1 FILLER_49_302 ();
 sg13g2_decap_8 FILLER_49_311 ();
 sg13g2_fill_1 FILLER_49_318 ();
 sg13g2_decap_8 FILLER_49_323 ();
 sg13g2_decap_8 FILLER_49_330 ();
 sg13g2_decap_4 FILLER_49_337 ();
 sg13g2_fill_1 FILLER_49_341 ();
 sg13g2_decap_8 FILLER_49_347 ();
 sg13g2_decap_8 FILLER_49_361 ();
 sg13g2_fill_1 FILLER_49_368 ();
 sg13g2_decap_8 FILLER_49_379 ();
 sg13g2_decap_4 FILLER_49_386 ();
 sg13g2_fill_2 FILLER_49_394 ();
 sg13g2_decap_4 FILLER_49_404 ();
 sg13g2_decap_8 FILLER_49_412 ();
 sg13g2_decap_4 FILLER_49_419 ();
 sg13g2_fill_1 FILLER_49_423 ();
 sg13g2_decap_8 FILLER_49_428 ();
 sg13g2_decap_8 FILLER_49_435 ();
 sg13g2_fill_2 FILLER_49_442 ();
 sg13g2_decap_8 FILLER_49_486 ();
 sg13g2_decap_8 FILLER_49_493 ();
 sg13g2_decap_4 FILLER_49_500 ();
 sg13g2_decap_8 FILLER_49_509 ();
 sg13g2_decap_8 FILLER_49_516 ();
 sg13g2_decap_8 FILLER_49_523 ();
 sg13g2_fill_2 FILLER_49_530 ();
 sg13g2_fill_1 FILLER_49_532 ();
 sg13g2_decap_8 FILLER_49_542 ();
 sg13g2_decap_8 FILLER_49_549 ();
 sg13g2_decap_8 FILLER_49_556 ();
 sg13g2_decap_4 FILLER_49_563 ();
 sg13g2_fill_1 FILLER_49_567 ();
 sg13g2_decap_8 FILLER_49_591 ();
 sg13g2_fill_2 FILLER_49_598 ();
 sg13g2_decap_8 FILLER_49_605 ();
 sg13g2_fill_2 FILLER_49_627 ();
 sg13g2_fill_1 FILLER_49_629 ();
 sg13g2_fill_1 FILLER_49_635 ();
 sg13g2_fill_2 FILLER_49_641 ();
 sg13g2_fill_1 FILLER_49_643 ();
 sg13g2_decap_4 FILLER_49_655 ();
 sg13g2_fill_1 FILLER_49_659 ();
 sg13g2_fill_2 FILLER_49_676 ();
 sg13g2_fill_1 FILLER_49_678 ();
 sg13g2_decap_8 FILLER_49_685 ();
 sg13g2_decap_8 FILLER_49_696 ();
 sg13g2_decap_4 FILLER_49_703 ();
 sg13g2_fill_2 FILLER_49_714 ();
 sg13g2_decap_4 FILLER_49_721 ();
 sg13g2_decap_4 FILLER_49_756 ();
 sg13g2_fill_1 FILLER_49_760 ();
 sg13g2_fill_2 FILLER_49_766 ();
 sg13g2_fill_2 FILLER_49_773 ();
 sg13g2_fill_1 FILLER_49_775 ();
 sg13g2_fill_1 FILLER_49_786 ();
 sg13g2_fill_2 FILLER_49_819 ();
 sg13g2_fill_1 FILLER_49_821 ();
 sg13g2_decap_4 FILLER_49_833 ();
 sg13g2_fill_1 FILLER_49_837 ();
 sg13g2_fill_2 FILLER_49_875 ();
 sg13g2_fill_1 FILLER_49_877 ();
 sg13g2_decap_8 FILLER_50_0 ();
 sg13g2_decap_8 FILLER_50_7 ();
 sg13g2_fill_2 FILLER_50_14 ();
 sg13g2_decap_4 FILLER_50_36 ();
 sg13g2_fill_1 FILLER_50_47 ();
 sg13g2_fill_2 FILLER_50_71 ();
 sg13g2_fill_2 FILLER_50_78 ();
 sg13g2_fill_1 FILLER_50_87 ();
 sg13g2_fill_1 FILLER_50_93 ();
 sg13g2_fill_1 FILLER_50_99 ();
 sg13g2_fill_2 FILLER_50_110 ();
 sg13g2_fill_2 FILLER_50_117 ();
 sg13g2_fill_1 FILLER_50_119 ();
 sg13g2_fill_1 FILLER_50_125 ();
 sg13g2_decap_4 FILLER_50_131 ();
 sg13g2_fill_1 FILLER_50_135 ();
 sg13g2_fill_2 FILLER_50_141 ();
 sg13g2_fill_1 FILLER_50_143 ();
 sg13g2_decap_8 FILLER_50_152 ();
 sg13g2_decap_8 FILLER_50_159 ();
 sg13g2_decap_8 FILLER_50_166 ();
 sg13g2_fill_2 FILLER_50_189 ();
 sg13g2_fill_2 FILLER_50_195 ();
 sg13g2_fill_1 FILLER_50_197 ();
 sg13g2_decap_4 FILLER_50_212 ();
 sg13g2_fill_1 FILLER_50_216 ();
 sg13g2_decap_8 FILLER_50_227 ();
 sg13g2_decap_4 FILLER_50_234 ();
 sg13g2_decap_8 FILLER_50_246 ();
 sg13g2_decap_8 FILLER_50_253 ();
 sg13g2_decap_4 FILLER_50_260 ();
 sg13g2_fill_1 FILLER_50_264 ();
 sg13g2_decap_8 FILLER_50_270 ();
 sg13g2_decap_8 FILLER_50_277 ();
 sg13g2_fill_1 FILLER_50_284 ();
 sg13g2_decap_4 FILLER_50_290 ();
 sg13g2_fill_2 FILLER_50_302 ();
 sg13g2_fill_1 FILLER_50_304 ();
 sg13g2_decap_8 FILLER_50_339 ();
 sg13g2_fill_1 FILLER_50_346 ();
 sg13g2_decap_8 FILLER_50_360 ();
 sg13g2_decap_4 FILLER_50_367 ();
 sg13g2_fill_2 FILLER_50_371 ();
 sg13g2_decap_8 FILLER_50_381 ();
 sg13g2_decap_8 FILLER_50_388 ();
 sg13g2_fill_2 FILLER_50_395 ();
 sg13g2_fill_1 FILLER_50_410 ();
 sg13g2_fill_2 FILLER_50_415 ();
 sg13g2_fill_2 FILLER_50_421 ();
 sg13g2_fill_1 FILLER_50_432 ();
 sg13g2_fill_1 FILLER_50_437 ();
 sg13g2_fill_1 FILLER_50_443 ();
 sg13g2_decap_4 FILLER_50_450 ();
 sg13g2_fill_1 FILLER_50_454 ();
 sg13g2_fill_2 FILLER_50_471 ();
 sg13g2_fill_1 FILLER_50_473 ();
 sg13g2_fill_1 FILLER_50_487 ();
 sg13g2_decap_4 FILLER_50_514 ();
 sg13g2_fill_1 FILLER_50_518 ();
 sg13g2_decap_8 FILLER_50_524 ();
 sg13g2_decap_8 FILLER_50_531 ();
 sg13g2_fill_2 FILLER_50_538 ();
 sg13g2_decap_8 FILLER_50_544 ();
 sg13g2_decap_8 FILLER_50_551 ();
 sg13g2_decap_8 FILLER_50_558 ();
 sg13g2_decap_8 FILLER_50_565 ();
 sg13g2_decap_4 FILLER_50_595 ();
 sg13g2_fill_1 FILLER_50_599 ();
 sg13g2_decap_8 FILLER_50_604 ();
 sg13g2_decap_4 FILLER_50_611 ();
 sg13g2_decap_8 FILLER_50_620 ();
 sg13g2_fill_1 FILLER_50_631 ();
 sg13g2_decap_8 FILLER_50_645 ();
 sg13g2_decap_8 FILLER_50_652 ();
 sg13g2_fill_1 FILLER_50_659 ();
 sg13g2_decap_4 FILLER_50_665 ();
 sg13g2_fill_1 FILLER_50_669 ();
 sg13g2_decap_4 FILLER_50_674 ();
 sg13g2_fill_2 FILLER_50_688 ();
 sg13g2_decap_8 FILLER_50_699 ();
 sg13g2_fill_1 FILLER_50_706 ();
 sg13g2_decap_4 FILLER_50_713 ();
 sg13g2_decap_4 FILLER_50_740 ();
 sg13g2_fill_1 FILLER_50_744 ();
 sg13g2_decap_8 FILLER_50_757 ();
 sg13g2_decap_4 FILLER_50_764 ();
 sg13g2_fill_1 FILLER_50_768 ();
 sg13g2_fill_1 FILLER_50_779 ();
 sg13g2_decap_4 FILLER_50_785 ();
 sg13g2_fill_1 FILLER_50_789 ();
 sg13g2_fill_1 FILLER_50_808 ();
 sg13g2_fill_2 FILLER_50_814 ();
 sg13g2_fill_1 FILLER_50_816 ();
 sg13g2_decap_4 FILLER_50_822 ();
 sg13g2_fill_2 FILLER_50_826 ();
 sg13g2_decap_8 FILLER_50_840 ();
 sg13g2_decap_8 FILLER_50_847 ();
 sg13g2_decap_8 FILLER_50_854 ();
 sg13g2_decap_8 FILLER_50_861 ();
 sg13g2_decap_8 FILLER_50_868 ();
 sg13g2_fill_2 FILLER_50_875 ();
 sg13g2_fill_1 FILLER_50_877 ();
 sg13g2_decap_8 FILLER_51_0 ();
 sg13g2_decap_8 FILLER_51_7 ();
 sg13g2_decap_8 FILLER_51_14 ();
 sg13g2_fill_1 FILLER_51_34 ();
 sg13g2_fill_2 FILLER_51_57 ();
 sg13g2_fill_2 FILLER_51_64 ();
 sg13g2_fill_2 FILLER_51_71 ();
 sg13g2_fill_1 FILLER_51_73 ();
 sg13g2_fill_2 FILLER_51_79 ();
 sg13g2_fill_1 FILLER_51_81 ();
 sg13g2_fill_2 FILLER_51_92 ();
 sg13g2_fill_1 FILLER_51_94 ();
 sg13g2_fill_1 FILLER_51_118 ();
 sg13g2_fill_1 FILLER_51_123 ();
 sg13g2_fill_1 FILLER_51_128 ();
 sg13g2_decap_4 FILLER_51_133 ();
 sg13g2_decap_8 FILLER_51_141 ();
 sg13g2_decap_8 FILLER_51_154 ();
 sg13g2_decap_8 FILLER_51_161 ();
 sg13g2_decap_8 FILLER_51_168 ();
 sg13g2_decap_8 FILLER_51_175 ();
 sg13g2_fill_2 FILLER_51_182 ();
 sg13g2_fill_1 FILLER_51_184 ();
 sg13g2_fill_2 FILLER_51_189 ();
 sg13g2_decap_4 FILLER_51_211 ();
 sg13g2_fill_2 FILLER_51_222 ();
 sg13g2_fill_2 FILLER_51_238 ();
 sg13g2_fill_1 FILLER_51_240 ();
 sg13g2_decap_8 FILLER_51_261 ();
 sg13g2_decap_8 FILLER_51_268 ();
 sg13g2_fill_2 FILLER_51_275 ();
 sg13g2_decap_8 FILLER_51_282 ();
 sg13g2_fill_2 FILLER_51_289 ();
 sg13g2_fill_1 FILLER_51_291 ();
 sg13g2_decap_4 FILLER_51_300 ();
 sg13g2_decap_8 FILLER_51_321 ();
 sg13g2_decap_8 FILLER_51_328 ();
 sg13g2_decap_8 FILLER_51_335 ();
 sg13g2_fill_1 FILLER_51_342 ();
 sg13g2_fill_1 FILLER_51_361 ();
 sg13g2_fill_2 FILLER_51_371 ();
 sg13g2_fill_1 FILLER_51_377 ();
 sg13g2_decap_4 FILLER_51_383 ();
 sg13g2_fill_2 FILLER_51_387 ();
 sg13g2_fill_1 FILLER_51_402 ();
 sg13g2_fill_1 FILLER_51_408 ();
 sg13g2_fill_1 FILLER_51_414 ();
 sg13g2_fill_1 FILLER_51_420 ();
 sg13g2_fill_2 FILLER_51_426 ();
 sg13g2_fill_2 FILLER_51_433 ();
 sg13g2_fill_1 FILLER_51_435 ();
 sg13g2_decap_8 FILLER_51_450 ();
 sg13g2_fill_1 FILLER_51_457 ();
 sg13g2_decap_8 FILLER_51_463 ();
 sg13g2_decap_8 FILLER_51_470 ();
 sg13g2_fill_2 FILLER_51_477 ();
 sg13g2_decap_8 FILLER_51_508 ();
 sg13g2_fill_1 FILLER_51_515 ();
 sg13g2_decap_8 FILLER_51_539 ();
 sg13g2_decap_8 FILLER_51_546 ();
 sg13g2_decap_8 FILLER_51_553 ();
 sg13g2_fill_1 FILLER_51_560 ();
 sg13g2_fill_2 FILLER_51_569 ();
 sg13g2_fill_1 FILLER_51_571 ();
 sg13g2_fill_1 FILLER_51_577 ();
 sg13g2_fill_2 FILLER_51_584 ();
 sg13g2_fill_1 FILLER_51_586 ();
 sg13g2_fill_2 FILLER_51_592 ();
 sg13g2_fill_1 FILLER_51_594 ();
 sg13g2_decap_4 FILLER_51_601 ();
 sg13g2_fill_1 FILLER_51_605 ();
 sg13g2_fill_1 FILLER_51_611 ();
 sg13g2_decap_4 FILLER_51_637 ();
 sg13g2_fill_2 FILLER_51_641 ();
 sg13g2_fill_2 FILLER_51_657 ();
 sg13g2_fill_1 FILLER_51_659 ();
 sg13g2_decap_4 FILLER_51_665 ();
 sg13g2_fill_1 FILLER_51_674 ();
 sg13g2_fill_2 FILLER_51_680 ();
 sg13g2_fill_1 FILLER_51_682 ();
 sg13g2_decap_4 FILLER_51_688 ();
 sg13g2_fill_2 FILLER_51_692 ();
 sg13g2_decap_8 FILLER_51_704 ();
 sg13g2_decap_8 FILLER_51_711 ();
 sg13g2_fill_2 FILLER_51_726 ();
 sg13g2_decap_8 FILLER_51_744 ();
 sg13g2_fill_1 FILLER_51_751 ();
 sg13g2_fill_1 FILLER_51_767 ();
 sg13g2_fill_2 FILLER_51_795 ();
 sg13g2_decap_4 FILLER_51_801 ();
 sg13g2_fill_1 FILLER_51_805 ();
 sg13g2_fill_2 FILLER_51_810 ();
 sg13g2_fill_1 FILLER_51_812 ();
 sg13g2_decap_8 FILLER_51_818 ();
 sg13g2_fill_1 FILLER_51_825 ();
 sg13g2_decap_8 FILLER_51_834 ();
 sg13g2_decap_8 FILLER_51_841 ();
 sg13g2_decap_8 FILLER_51_848 ();
 sg13g2_fill_1 FILLER_51_855 ();
 sg13g2_decap_8 FILLER_51_860 ();
 sg13g2_decap_8 FILLER_51_867 ();
 sg13g2_decap_4 FILLER_51_874 ();
 sg13g2_decap_8 FILLER_52_0 ();
 sg13g2_decap_8 FILLER_52_7 ();
 sg13g2_decap_8 FILLER_52_14 ();
 sg13g2_fill_2 FILLER_52_21 ();
 sg13g2_fill_1 FILLER_52_23 ();
 sg13g2_fill_2 FILLER_52_29 ();
 sg13g2_fill_1 FILLER_52_31 ();
 sg13g2_fill_2 FILLER_52_49 ();
 sg13g2_fill_2 FILLER_52_75 ();
 sg13g2_fill_2 FILLER_52_83 ();
 sg13g2_fill_1 FILLER_52_85 ();
 sg13g2_fill_1 FILLER_52_91 ();
 sg13g2_fill_2 FILLER_52_97 ();
 sg13g2_fill_1 FILLER_52_99 ();
 sg13g2_fill_1 FILLER_52_113 ();
 sg13g2_fill_2 FILLER_52_135 ();
 sg13g2_decap_8 FILLER_52_149 ();
 sg13g2_decap_8 FILLER_52_161 ();
 sg13g2_decap_8 FILLER_52_168 ();
 sg13g2_decap_4 FILLER_52_175 ();
 sg13g2_fill_2 FILLER_52_179 ();
 sg13g2_decap_4 FILLER_52_198 ();
 sg13g2_fill_1 FILLER_52_202 ();
 sg13g2_fill_1 FILLER_52_233 ();
 sg13g2_decap_4 FILLER_52_239 ();
 sg13g2_fill_1 FILLER_52_243 ();
 sg13g2_decap_8 FILLER_52_270 ();
 sg13g2_decap_8 FILLER_52_277 ();
 sg13g2_decap_4 FILLER_52_284 ();
 sg13g2_fill_2 FILLER_52_288 ();
 sg13g2_fill_2 FILLER_52_311 ();
 sg13g2_fill_1 FILLER_52_313 ();
 sg13g2_decap_8 FILLER_52_322 ();
 sg13g2_decap_4 FILLER_52_397 ();
 sg13g2_decap_8 FILLER_52_406 ();
 sg13g2_decap_8 FILLER_52_413 ();
 sg13g2_fill_2 FILLER_52_425 ();
 sg13g2_fill_2 FILLER_52_431 ();
 sg13g2_fill_1 FILLER_52_446 ();
 sg13g2_fill_1 FILLER_52_451 ();
 sg13g2_fill_1 FILLER_52_457 ();
 sg13g2_fill_1 FILLER_52_463 ();
 sg13g2_fill_2 FILLER_52_469 ();
 sg13g2_fill_2 FILLER_52_475 ();
 sg13g2_fill_1 FILLER_52_482 ();
 sg13g2_decap_8 FILLER_52_488 ();
 sg13g2_decap_8 FILLER_52_495 ();
 sg13g2_decap_8 FILLER_52_502 ();
 sg13g2_decap_8 FILLER_52_509 ();
 sg13g2_decap_4 FILLER_52_516 ();
 sg13g2_decap_4 FILLER_52_525 ();
 sg13g2_fill_2 FILLER_52_529 ();
 sg13g2_decap_4 FILLER_52_546 ();
 sg13g2_fill_1 FILLER_52_550 ();
 sg13g2_decap_8 FILLER_52_556 ();
 sg13g2_decap_8 FILLER_52_563 ();
 sg13g2_decap_4 FILLER_52_570 ();
 sg13g2_fill_1 FILLER_52_574 ();
 sg13g2_fill_1 FILLER_52_584 ();
 sg13g2_fill_2 FILLER_52_591 ();
 sg13g2_fill_2 FILLER_52_598 ();
 sg13g2_fill_2 FILLER_52_604 ();
 sg13g2_fill_2 FILLER_52_611 ();
 sg13g2_fill_1 FILLER_52_613 ();
 sg13g2_fill_1 FILLER_52_619 ();
 sg13g2_fill_2 FILLER_52_626 ();
 sg13g2_fill_1 FILLER_52_628 ();
 sg13g2_decap_4 FILLER_52_656 ();
 sg13g2_fill_1 FILLER_52_660 ();
 sg13g2_decap_4 FILLER_52_685 ();
 sg13g2_decap_8 FILLER_52_702 ();
 sg13g2_fill_2 FILLER_52_709 ();
 sg13g2_decap_4 FILLER_52_719 ();
 sg13g2_fill_1 FILLER_52_729 ();
 sg13g2_decap_4 FILLER_52_746 ();
 sg13g2_fill_1 FILLER_52_750 ();
 sg13g2_fill_1 FILLER_52_764 ();
 sg13g2_fill_2 FILLER_52_769 ();
 sg13g2_fill_1 FILLER_52_771 ();
 sg13g2_decap_4 FILLER_52_777 ();
 sg13g2_fill_1 FILLER_52_781 ();
 sg13g2_decap_4 FILLER_52_787 ();
 sg13g2_fill_1 FILLER_52_791 ();
 sg13g2_decap_4 FILLER_52_797 ();
 sg13g2_decap_8 FILLER_52_805 ();
 sg13g2_decap_8 FILLER_52_812 ();
 sg13g2_decap_4 FILLER_52_819 ();
 sg13g2_fill_2 FILLER_52_836 ();
 sg13g2_decap_4 FILLER_52_843 ();
 sg13g2_fill_2 FILLER_52_847 ();
 sg13g2_fill_2 FILLER_52_875 ();
 sg13g2_fill_1 FILLER_52_877 ();
 sg13g2_decap_8 FILLER_53_0 ();
 sg13g2_fill_2 FILLER_53_7 ();
 sg13g2_fill_1 FILLER_53_9 ();
 sg13g2_decap_8 FILLER_53_19 ();
 sg13g2_decap_8 FILLER_53_26 ();
 sg13g2_fill_1 FILLER_53_38 ();
 sg13g2_fill_1 FILLER_53_47 ();
 sg13g2_fill_2 FILLER_53_75 ();
 sg13g2_fill_1 FILLER_53_77 ();
 sg13g2_decap_4 FILLER_53_89 ();
 sg13g2_decap_4 FILLER_53_119 ();
 sg13g2_fill_1 FILLER_53_123 ();
 sg13g2_fill_1 FILLER_53_154 ();
 sg13g2_fill_2 FILLER_53_178 ();
 sg13g2_fill_1 FILLER_53_180 ();
 sg13g2_decap_8 FILLER_53_185 ();
 sg13g2_fill_1 FILLER_53_192 ();
 sg13g2_fill_2 FILLER_53_202 ();
 sg13g2_fill_1 FILLER_53_204 ();
 sg13g2_decap_8 FILLER_53_209 ();
 sg13g2_fill_2 FILLER_53_216 ();
 sg13g2_fill_1 FILLER_53_218 ();
 sg13g2_decap_8 FILLER_53_223 ();
 sg13g2_decap_4 FILLER_53_230 ();
 sg13g2_fill_2 FILLER_53_238 ();
 sg13g2_fill_2 FILLER_53_262 ();
 sg13g2_fill_2 FILLER_53_304 ();
 sg13g2_fill_1 FILLER_53_306 ();
 sg13g2_decap_8 FILLER_53_324 ();
 sg13g2_decap_4 FILLER_53_331 ();
 sg13g2_fill_2 FILLER_53_335 ();
 sg13g2_decap_4 FILLER_53_347 ();
 sg13g2_fill_1 FILLER_53_360 ();
 sg13g2_fill_2 FILLER_53_378 ();
 sg13g2_fill_1 FILLER_53_380 ();
 sg13g2_fill_2 FILLER_53_385 ();
 sg13g2_fill_1 FILLER_53_398 ();
 sg13g2_fill_2 FILLER_53_410 ();
 sg13g2_decap_8 FILLER_53_427 ();
 sg13g2_fill_1 FILLER_53_434 ();
 sg13g2_fill_2 FILLER_53_449 ();
 sg13g2_fill_1 FILLER_53_464 ();
 sg13g2_fill_2 FILLER_53_470 ();
 sg13g2_fill_1 FILLER_53_472 ();
 sg13g2_decap_8 FILLER_53_508 ();
 sg13g2_decap_8 FILLER_53_515 ();
 sg13g2_decap_8 FILLER_53_522 ();
 sg13g2_fill_2 FILLER_53_529 ();
 sg13g2_fill_2 FILLER_53_537 ();
 sg13g2_decap_8 FILLER_53_544 ();
 sg13g2_decap_8 FILLER_53_551 ();
 sg13g2_decap_4 FILLER_53_558 ();
 sg13g2_fill_2 FILLER_53_562 ();
 sg13g2_decap_8 FILLER_53_569 ();
 sg13g2_decap_4 FILLER_53_576 ();
 sg13g2_fill_2 FILLER_53_580 ();
 sg13g2_fill_2 FILLER_53_587 ();
 sg13g2_fill_2 FILLER_53_601 ();
 sg13g2_fill_1 FILLER_53_603 ();
 sg13g2_fill_2 FILLER_53_610 ();
 sg13g2_fill_1 FILLER_53_612 ();
 sg13g2_fill_2 FILLER_53_619 ();
 sg13g2_decap_8 FILLER_53_629 ();
 sg13g2_fill_2 FILLER_53_636 ();
 sg13g2_decap_8 FILLER_53_645 ();
 sg13g2_fill_2 FILLER_53_652 ();
 sg13g2_fill_2 FILLER_53_663 ();
 sg13g2_fill_1 FILLER_53_684 ();
 sg13g2_fill_2 FILLER_53_715 ();
 sg13g2_fill_2 FILLER_53_722 ();
 sg13g2_fill_1 FILLER_53_724 ();
 sg13g2_fill_2 FILLER_53_751 ();
 sg13g2_fill_1 FILLER_53_753 ();
 sg13g2_decap_8 FILLER_53_772 ();
 sg13g2_fill_2 FILLER_53_779 ();
 sg13g2_decap_4 FILLER_53_786 ();
 sg13g2_fill_2 FILLER_53_790 ();
 sg13g2_decap_8 FILLER_53_798 ();
 sg13g2_decap_8 FILLER_53_805 ();
 sg13g2_decap_8 FILLER_53_812 ();
 sg13g2_decap_8 FILLER_53_819 ();
 sg13g2_decap_8 FILLER_53_826 ();
 sg13g2_decap_8 FILLER_53_841 ();
 sg13g2_fill_2 FILLER_53_848 ();
 sg13g2_decap_8 FILLER_53_862 ();
 sg13g2_decap_8 FILLER_53_869 ();
 sg13g2_fill_2 FILLER_53_876 ();
 sg13g2_decap_8 FILLER_54_0 ();
 sg13g2_decap_8 FILLER_54_7 ();
 sg13g2_fill_2 FILLER_54_14 ();
 sg13g2_decap_8 FILLER_54_20 ();
 sg13g2_fill_2 FILLER_54_42 ();
 sg13g2_fill_2 FILLER_54_48 ();
 sg13g2_fill_2 FILLER_54_55 ();
 sg13g2_decap_4 FILLER_54_67 ();
 sg13g2_fill_1 FILLER_54_71 ();
 sg13g2_fill_2 FILLER_54_82 ();
 sg13g2_fill_1 FILLER_54_84 ();
 sg13g2_fill_1 FILLER_54_90 ();
 sg13g2_fill_1 FILLER_54_101 ();
 sg13g2_decap_8 FILLER_54_110 ();
 sg13g2_decap_8 FILLER_54_117 ();
 sg13g2_fill_2 FILLER_54_124 ();
 sg13g2_decap_8 FILLER_54_149 ();
 sg13g2_decap_8 FILLER_54_156 ();
 sg13g2_decap_4 FILLER_54_163 ();
 sg13g2_fill_1 FILLER_54_167 ();
 sg13g2_fill_2 FILLER_54_173 ();
 sg13g2_fill_1 FILLER_54_175 ();
 sg13g2_fill_1 FILLER_54_184 ();
 sg13g2_decap_8 FILLER_54_205 ();
 sg13g2_decap_8 FILLER_54_212 ();
 sg13g2_fill_2 FILLER_54_219 ();
 sg13g2_decap_8 FILLER_54_225 ();
 sg13g2_fill_2 FILLER_54_238 ();
 sg13g2_decap_8 FILLER_54_256 ();
 sg13g2_decap_8 FILLER_54_263 ();
 sg13g2_fill_1 FILLER_54_270 ();
 sg13g2_fill_2 FILLER_54_275 ();
 sg13g2_fill_1 FILLER_54_277 ();
 sg13g2_decap_8 FILLER_54_283 ();
 sg13g2_decap_4 FILLER_54_290 ();
 sg13g2_fill_1 FILLER_54_294 ();
 sg13g2_fill_2 FILLER_54_318 ();
 sg13g2_fill_1 FILLER_54_324 ();
 sg13g2_decap_8 FILLER_54_335 ();
 sg13g2_fill_1 FILLER_54_350 ();
 sg13g2_fill_2 FILLER_54_356 ();
 sg13g2_fill_2 FILLER_54_370 ();
 sg13g2_decap_8 FILLER_54_381 ();
 sg13g2_fill_2 FILLER_54_388 ();
 sg13g2_fill_1 FILLER_54_390 ();
 sg13g2_fill_2 FILLER_54_412 ();
 sg13g2_fill_1 FILLER_54_414 ();
 sg13g2_fill_1 FILLER_54_419 ();
 sg13g2_decap_8 FILLER_54_446 ();
 sg13g2_decap_8 FILLER_54_453 ();
 sg13g2_decap_8 FILLER_54_460 ();
 sg13g2_decap_8 FILLER_54_467 ();
 sg13g2_decap_4 FILLER_54_474 ();
 sg13g2_fill_1 FILLER_54_496 ();
 sg13g2_fill_1 FILLER_54_502 ();
 sg13g2_decap_8 FILLER_54_507 ();
 sg13g2_decap_8 FILLER_54_518 ();
 sg13g2_decap_4 FILLER_54_525 ();
 sg13g2_decap_8 FILLER_54_557 ();
 sg13g2_decap_8 FILLER_54_564 ();
 sg13g2_decap_4 FILLER_54_571 ();
 sg13g2_fill_1 FILLER_54_575 ();
 sg13g2_fill_1 FILLER_54_580 ();
 sg13g2_decap_4 FILLER_54_588 ();
 sg13g2_fill_2 FILLER_54_592 ();
 sg13g2_fill_2 FILLER_54_598 ();
 sg13g2_fill_2 FILLER_54_618 ();
 sg13g2_fill_1 FILLER_54_620 ();
 sg13g2_fill_2 FILLER_54_637 ();
 sg13g2_fill_1 FILLER_54_639 ();
 sg13g2_decap_8 FILLER_54_644 ();
 sg13g2_decap_8 FILLER_54_651 ();
 sg13g2_decap_4 FILLER_54_674 ();
 sg13g2_fill_1 FILLER_54_678 ();
 sg13g2_decap_8 FILLER_54_683 ();
 sg13g2_fill_1 FILLER_54_690 ();
 sg13g2_decap_4 FILLER_54_696 ();
 sg13g2_fill_1 FILLER_54_700 ();
 sg13g2_fill_1 FILLER_54_716 ();
 sg13g2_decap_8 FILLER_54_726 ();
 sg13g2_fill_2 FILLER_54_733 ();
 sg13g2_fill_1 FILLER_54_735 ();
 sg13g2_decap_8 FILLER_54_740 ();
 sg13g2_decap_4 FILLER_54_747 ();
 sg13g2_fill_1 FILLER_54_751 ();
 sg13g2_decap_8 FILLER_54_761 ();
 sg13g2_fill_2 FILLER_54_768 ();
 sg13g2_fill_1 FILLER_54_770 ();
 sg13g2_decap_4 FILLER_54_775 ();
 sg13g2_decap_4 FILLER_54_788 ();
 sg13g2_fill_1 FILLER_54_801 ();
 sg13g2_decap_8 FILLER_54_805 ();
 sg13g2_fill_1 FILLER_54_812 ();
 sg13g2_fill_2 FILLER_54_832 ();
 sg13g2_decap_8 FILLER_54_844 ();
 sg13g2_fill_1 FILLER_54_851 ();
 sg13g2_decap_8 FILLER_55_0 ();
 sg13g2_decap_8 FILLER_55_7 ();
 sg13g2_decap_8 FILLER_55_14 ();
 sg13g2_fill_1 FILLER_55_21 ();
 sg13g2_decap_4 FILLER_55_27 ();
 sg13g2_fill_1 FILLER_55_57 ();
 sg13g2_fill_2 FILLER_55_83 ();
 sg13g2_decap_4 FILLER_55_90 ();
 sg13g2_fill_2 FILLER_55_102 ();
 sg13g2_decap_8 FILLER_55_135 ();
 sg13g2_decap_8 FILLER_55_142 ();
 sg13g2_decap_8 FILLER_55_149 ();
 sg13g2_decap_8 FILLER_55_156 ();
 sg13g2_decap_8 FILLER_55_163 ();
 sg13g2_decap_8 FILLER_55_170 ();
 sg13g2_fill_1 FILLER_55_177 ();
 sg13g2_decap_4 FILLER_55_184 ();
 sg13g2_fill_2 FILLER_55_188 ();
 sg13g2_decap_8 FILLER_55_200 ();
 sg13g2_decap_8 FILLER_55_207 ();
 sg13g2_decap_8 FILLER_55_253 ();
 sg13g2_fill_2 FILLER_55_260 ();
 sg13g2_fill_1 FILLER_55_262 ();
 sg13g2_fill_1 FILLER_55_271 ();
 sg13g2_decap_8 FILLER_55_277 ();
 sg13g2_decap_8 FILLER_55_284 ();
 sg13g2_decap_8 FILLER_55_291 ();
 sg13g2_decap_8 FILLER_55_298 ();
 sg13g2_fill_2 FILLER_55_305 ();
 sg13g2_decap_4 FILLER_55_314 ();
 sg13g2_decap_4 FILLER_55_326 ();
 sg13g2_fill_2 FILLER_55_330 ();
 sg13g2_decap_8 FILLER_55_336 ();
 sg13g2_decap_4 FILLER_55_343 ();
 sg13g2_fill_2 FILLER_55_347 ();
 sg13g2_decap_8 FILLER_55_353 ();
 sg13g2_decap_8 FILLER_55_360 ();
 sg13g2_decap_8 FILLER_55_367 ();
 sg13g2_fill_1 FILLER_55_374 ();
 sg13g2_decap_8 FILLER_55_383 ();
 sg13g2_fill_2 FILLER_55_390 ();
 sg13g2_fill_1 FILLER_55_392 ();
 sg13g2_decap_4 FILLER_55_397 ();
 sg13g2_decap_8 FILLER_55_405 ();
 sg13g2_decap_8 FILLER_55_412 ();
 sg13g2_decap_4 FILLER_55_419 ();
 sg13g2_fill_2 FILLER_55_428 ();
 sg13g2_decap_4 FILLER_55_443 ();
 sg13g2_decap_4 FILLER_55_456 ();
 sg13g2_fill_1 FILLER_55_464 ();
 sg13g2_decap_8 FILLER_55_503 ();
 sg13g2_decap_8 FILLER_55_510 ();
 sg13g2_decap_4 FILLER_55_517 ();
 sg13g2_fill_2 FILLER_55_521 ();
 sg13g2_fill_2 FILLER_55_552 ();
 sg13g2_fill_1 FILLER_55_554 ();
 sg13g2_decap_8 FILLER_55_560 ();
 sg13g2_decap_8 FILLER_55_574 ();
 sg13g2_decap_8 FILLER_55_581 ();
 sg13g2_decap_8 FILLER_55_588 ();
 sg13g2_fill_1 FILLER_55_595 ();
 sg13g2_decap_8 FILLER_55_604 ();
 sg13g2_decap_8 FILLER_55_611 ();
 sg13g2_fill_2 FILLER_55_618 ();
 sg13g2_fill_2 FILLER_55_644 ();
 sg13g2_decap_8 FILLER_55_668 ();
 sg13g2_decap_4 FILLER_55_675 ();
 sg13g2_fill_2 FILLER_55_679 ();
 sg13g2_decap_4 FILLER_55_697 ();
 sg13g2_fill_2 FILLER_55_701 ();
 sg13g2_fill_2 FILLER_55_709 ();
 sg13g2_fill_1 FILLER_55_711 ();
 sg13g2_decap_8 FILLER_55_717 ();
 sg13g2_decap_4 FILLER_55_724 ();
 sg13g2_fill_2 FILLER_55_728 ();
 sg13g2_decap_8 FILLER_55_735 ();
 sg13g2_decap_8 FILLER_55_742 ();
 sg13g2_decap_8 FILLER_55_749 ();
 sg13g2_decap_8 FILLER_55_756 ();
 sg13g2_decap_8 FILLER_55_763 ();
 sg13g2_decap_8 FILLER_55_770 ();
 sg13g2_fill_1 FILLER_55_777 ();
 sg13g2_decap_8 FILLER_55_783 ();
 sg13g2_decap_8 FILLER_55_790 ();
 sg13g2_decap_8 FILLER_55_797 ();
 sg13g2_fill_1 FILLER_55_804 ();
 sg13g2_decap_8 FILLER_55_809 ();
 sg13g2_decap_4 FILLER_55_816 ();
 sg13g2_decap_8 FILLER_55_840 ();
 sg13g2_decap_8 FILLER_55_847 ();
 sg13g2_fill_1 FILLER_55_854 ();
 sg13g2_decap_8 FILLER_55_859 ();
 sg13g2_decap_8 FILLER_55_866 ();
 sg13g2_decap_4 FILLER_55_873 ();
 sg13g2_fill_1 FILLER_55_877 ();
 sg13g2_decap_8 FILLER_56_0 ();
 sg13g2_decap_8 FILLER_56_7 ();
 sg13g2_decap_4 FILLER_56_14 ();
 sg13g2_fill_1 FILLER_56_18 ();
 sg13g2_decap_4 FILLER_56_23 ();
 sg13g2_fill_2 FILLER_56_51 ();
 sg13g2_fill_1 FILLER_56_53 ();
 sg13g2_decap_4 FILLER_56_73 ();
 sg13g2_fill_2 FILLER_56_82 ();
 sg13g2_fill_1 FILLER_56_84 ();
 sg13g2_fill_2 FILLER_56_97 ();
 sg13g2_fill_1 FILLER_56_99 ();
 sg13g2_decap_4 FILLER_56_104 ();
 sg13g2_fill_1 FILLER_56_108 ();
 sg13g2_fill_2 FILLER_56_114 ();
 sg13g2_fill_1 FILLER_56_116 ();
 sg13g2_fill_2 FILLER_56_126 ();
 sg13g2_fill_1 FILLER_56_128 ();
 sg13g2_decap_8 FILLER_56_133 ();
 sg13g2_decap_8 FILLER_56_140 ();
 sg13g2_decap_8 FILLER_56_147 ();
 sg13g2_decap_8 FILLER_56_154 ();
 sg13g2_decap_8 FILLER_56_161 ();
 sg13g2_decap_8 FILLER_56_168 ();
 sg13g2_fill_2 FILLER_56_175 ();
 sg13g2_fill_1 FILLER_56_177 ();
 sg13g2_fill_2 FILLER_56_193 ();
 sg13g2_fill_1 FILLER_56_198 ();
 sg13g2_decap_8 FILLER_56_203 ();
 sg13g2_decap_8 FILLER_56_210 ();
 sg13g2_decap_8 FILLER_56_217 ();
 sg13g2_decap_4 FILLER_56_224 ();
 sg13g2_fill_2 FILLER_56_228 ();
 sg13g2_decap_8 FILLER_56_234 ();
 sg13g2_fill_1 FILLER_56_241 ();
 sg13g2_fill_1 FILLER_56_254 ();
 sg13g2_fill_2 FILLER_56_259 ();
 sg13g2_fill_1 FILLER_56_291 ();
 sg13g2_fill_1 FILLER_56_296 ();
 sg13g2_fill_1 FILLER_56_305 ();
 sg13g2_fill_1 FILLER_56_311 ();
 sg13g2_decap_4 FILLER_56_322 ();
 sg13g2_fill_1 FILLER_56_326 ();
 sg13g2_fill_1 FILLER_56_334 ();
 sg13g2_fill_1 FILLER_56_361 ();
 sg13g2_fill_1 FILLER_56_366 ();
 sg13g2_fill_1 FILLER_56_373 ();
 sg13g2_fill_1 FILLER_56_379 ();
 sg13g2_fill_2 FILLER_56_386 ();
 sg13g2_decap_8 FILLER_56_394 ();
 sg13g2_fill_1 FILLER_56_401 ();
 sg13g2_decap_4 FILLER_56_406 ();
 sg13g2_fill_1 FILLER_56_410 ();
 sg13g2_decap_8 FILLER_56_421 ();
 sg13g2_decap_8 FILLER_56_428 ();
 sg13g2_decap_8 FILLER_56_435 ();
 sg13g2_decap_8 FILLER_56_442 ();
 sg13g2_fill_1 FILLER_56_449 ();
 sg13g2_decap_8 FILLER_56_455 ();
 sg13g2_decap_4 FILLER_56_462 ();
 sg13g2_fill_2 FILLER_56_466 ();
 sg13g2_decap_8 FILLER_56_480 ();
 sg13g2_decap_4 FILLER_56_487 ();
 sg13g2_fill_1 FILLER_56_491 ();
 sg13g2_decap_8 FILLER_56_496 ();
 sg13g2_decap_8 FILLER_56_503 ();
 sg13g2_decap_4 FILLER_56_510 ();
 sg13g2_fill_2 FILLER_56_514 ();
 sg13g2_decap_8 FILLER_56_521 ();
 sg13g2_fill_1 FILLER_56_528 ();
 sg13g2_decap_4 FILLER_56_533 ();
 sg13g2_fill_1 FILLER_56_537 ();
 sg13g2_decap_8 FILLER_56_550 ();
 sg13g2_fill_2 FILLER_56_570 ();
 sg13g2_fill_1 FILLER_56_572 ();
 sg13g2_decap_8 FILLER_56_580 ();
 sg13g2_decap_8 FILLER_56_602 ();
 sg13g2_decap_4 FILLER_56_609 ();
 sg13g2_decap_8 FILLER_56_618 ();
 sg13g2_decap_8 FILLER_56_625 ();
 sg13g2_decap_4 FILLER_56_632 ();
 sg13g2_fill_2 FILLER_56_636 ();
 sg13g2_fill_2 FILLER_56_649 ();
 sg13g2_fill_1 FILLER_56_651 ();
 sg13g2_decap_8 FILLER_56_661 ();
 sg13g2_decap_8 FILLER_56_668 ();
 sg13g2_fill_1 FILLER_56_675 ();
 sg13g2_decap_8 FILLER_56_694 ();
 sg13g2_decap_8 FILLER_56_701 ();
 sg13g2_decap_8 FILLER_56_708 ();
 sg13g2_fill_2 FILLER_56_715 ();
 sg13g2_fill_2 FILLER_56_721 ();
 sg13g2_decap_8 FILLER_56_732 ();
 sg13g2_fill_2 FILLER_56_739 ();
 sg13g2_decap_8 FILLER_56_745 ();
 sg13g2_decap_8 FILLER_56_752 ();
 sg13g2_decap_8 FILLER_56_759 ();
 sg13g2_decap_8 FILLER_56_766 ();
 sg13g2_fill_1 FILLER_56_773 ();
 sg13g2_decap_8 FILLER_56_778 ();
 sg13g2_decap_8 FILLER_56_785 ();
 sg13g2_fill_2 FILLER_56_792 ();
 sg13g2_decap_8 FILLER_56_824 ();
 sg13g2_fill_1 FILLER_56_831 ();
 sg13g2_decap_4 FILLER_56_873 ();
 sg13g2_fill_1 FILLER_56_877 ();
 sg13g2_decap_8 FILLER_57_0 ();
 sg13g2_decap_4 FILLER_57_7 ();
 sg13g2_fill_1 FILLER_57_11 ();
 sg13g2_decap_4 FILLER_57_17 ();
 sg13g2_fill_2 FILLER_57_25 ();
 sg13g2_fill_1 FILLER_57_34 ();
 sg13g2_fill_1 FILLER_57_48 ();
 sg13g2_fill_1 FILLER_57_55 ();
 sg13g2_fill_2 FILLER_57_62 ();
 sg13g2_fill_1 FILLER_57_69 ();
 sg13g2_fill_2 FILLER_57_77 ();
 sg13g2_fill_2 FILLER_57_85 ();
 sg13g2_fill_2 FILLER_57_93 ();
 sg13g2_fill_1 FILLER_57_95 ();
 sg13g2_fill_2 FILLER_57_115 ();
 sg13g2_fill_1 FILLER_57_117 ();
 sg13g2_fill_2 FILLER_57_126 ();
 sg13g2_decap_4 FILLER_57_144 ();
 sg13g2_decap_8 FILLER_57_153 ();
 sg13g2_decap_8 FILLER_57_160 ();
 sg13g2_decap_4 FILLER_57_167 ();
 sg13g2_decap_4 FILLER_57_181 ();
 sg13g2_fill_1 FILLER_57_189 ();
 sg13g2_fill_1 FILLER_57_194 ();
 sg13g2_decap_8 FILLER_57_209 ();
 sg13g2_decap_4 FILLER_57_216 ();
 sg13g2_fill_1 FILLER_57_220 ();
 sg13g2_decap_8 FILLER_57_237 ();
 sg13g2_fill_1 FILLER_57_244 ();
 sg13g2_decap_8 FILLER_57_271 ();
 sg13g2_fill_2 FILLER_57_278 ();
 sg13g2_decap_8 FILLER_57_285 ();
 sg13g2_decap_8 FILLER_57_292 ();
 sg13g2_decap_8 FILLER_57_299 ();
 sg13g2_fill_2 FILLER_57_306 ();
 sg13g2_fill_1 FILLER_57_312 ();
 sg13g2_fill_1 FILLER_57_318 ();
 sg13g2_fill_2 FILLER_57_327 ();
 sg13g2_decap_4 FILLER_57_338 ();
 sg13g2_fill_1 FILLER_57_342 ();
 sg13g2_fill_1 FILLER_57_351 ();
 sg13g2_decap_4 FILLER_57_356 ();
 sg13g2_fill_2 FILLER_57_360 ();
 sg13g2_fill_2 FILLER_57_370 ();
 sg13g2_fill_1 FILLER_57_377 ();
 sg13g2_decap_8 FILLER_57_387 ();
 sg13g2_fill_1 FILLER_57_394 ();
 sg13g2_fill_1 FILLER_57_405 ();
 sg13g2_fill_2 FILLER_57_410 ();
 sg13g2_fill_2 FILLER_57_417 ();
 sg13g2_decap_4 FILLER_57_424 ();
 sg13g2_decap_4 FILLER_57_433 ();
 sg13g2_fill_2 FILLER_57_441 ();
 sg13g2_decap_8 FILLER_57_453 ();
 sg13g2_decap_8 FILLER_57_460 ();
 sg13g2_decap_4 FILLER_57_467 ();
 sg13g2_fill_2 FILLER_57_471 ();
 sg13g2_fill_2 FILLER_57_482 ();
 sg13g2_decap_4 FILLER_57_494 ();
 sg13g2_decap_8 FILLER_57_502 ();
 sg13g2_fill_2 FILLER_57_509 ();
 sg13g2_decap_4 FILLER_57_521 ();
 sg13g2_fill_1 FILLER_57_525 ();
 sg13g2_fill_1 FILLER_57_530 ();
 sg13g2_fill_1 FILLER_57_536 ();
 sg13g2_fill_2 FILLER_57_542 ();
 sg13g2_decap_8 FILLER_57_554 ();
 sg13g2_fill_1 FILLER_57_561 ();
 sg13g2_fill_2 FILLER_57_567 ();
 sg13g2_fill_1 FILLER_57_569 ();
 sg13g2_decap_8 FILLER_57_578 ();
 sg13g2_decap_8 FILLER_57_585 ();
 sg13g2_decap_8 FILLER_57_592 ();
 sg13g2_decap_8 FILLER_57_599 ();
 sg13g2_decap_8 FILLER_57_606 ();
 sg13g2_decap_8 FILLER_57_613 ();
 sg13g2_decap_8 FILLER_57_620 ();
 sg13g2_decap_4 FILLER_57_627 ();
 sg13g2_fill_2 FILLER_57_631 ();
 sg13g2_decap_8 FILLER_57_645 ();
 sg13g2_decap_8 FILLER_57_652 ();
 sg13g2_decap_8 FILLER_57_659 ();
 sg13g2_decap_4 FILLER_57_666 ();
 sg13g2_fill_2 FILLER_57_674 ();
 sg13g2_fill_1 FILLER_57_676 ();
 sg13g2_decap_4 FILLER_57_682 ();
 sg13g2_fill_2 FILLER_57_686 ();
 sg13g2_decap_4 FILLER_57_693 ();
 sg13g2_fill_1 FILLER_57_697 ();
 sg13g2_fill_1 FILLER_57_708 ();
 sg13g2_fill_1 FILLER_57_713 ();
 sg13g2_fill_1 FILLER_57_719 ();
 sg13g2_fill_1 FILLER_57_730 ();
 sg13g2_decap_4 FILLER_57_738 ();
 sg13g2_fill_1 FILLER_57_742 ();
 sg13g2_decap_8 FILLER_57_747 ();
 sg13g2_decap_4 FILLER_57_754 ();
 sg13g2_fill_1 FILLER_57_758 ();
 sg13g2_decap_8 FILLER_57_809 ();
 sg13g2_decap_8 FILLER_57_829 ();
 sg13g2_fill_2 FILLER_57_836 ();
 sg13g2_decap_8 FILLER_57_869 ();
 sg13g2_fill_2 FILLER_57_876 ();
 sg13g2_decap_8 FILLER_58_0 ();
 sg13g2_fill_2 FILLER_58_7 ();
 sg13g2_fill_1 FILLER_58_15 ();
 sg13g2_fill_1 FILLER_58_21 ();
 sg13g2_fill_2 FILLER_58_27 ();
 sg13g2_fill_2 FILLER_58_33 ();
 sg13g2_decap_8 FILLER_58_48 ();
 sg13g2_fill_2 FILLER_58_55 ();
 sg13g2_fill_1 FILLER_58_61 ();
 sg13g2_decap_4 FILLER_58_67 ();
 sg13g2_decap_8 FILLER_58_75 ();
 sg13g2_fill_1 FILLER_58_82 ();
 sg13g2_decap_4 FILLER_58_97 ();
 sg13g2_fill_1 FILLER_58_101 ();
 sg13g2_decap_4 FILLER_58_107 ();
 sg13g2_fill_1 FILLER_58_111 ();
 sg13g2_decap_4 FILLER_58_117 ();
 sg13g2_fill_2 FILLER_58_121 ();
 sg13g2_fill_2 FILLER_58_128 ();
 sg13g2_fill_1 FILLER_58_130 ();
 sg13g2_fill_1 FILLER_58_141 ();
 sg13g2_decap_8 FILLER_58_146 ();
 sg13g2_decap_4 FILLER_58_153 ();
 sg13g2_fill_1 FILLER_58_157 ();
 sg13g2_decap_8 FILLER_58_162 ();
 sg13g2_decap_4 FILLER_58_169 ();
 sg13g2_fill_1 FILLER_58_173 ();
 sg13g2_decap_4 FILLER_58_193 ();
 sg13g2_fill_1 FILLER_58_197 ();
 sg13g2_decap_4 FILLER_58_207 ();
 sg13g2_decap_8 FILLER_58_215 ();
 sg13g2_decap_8 FILLER_58_222 ();
 sg13g2_decap_4 FILLER_58_229 ();
 sg13g2_fill_1 FILLER_58_242 ();
 sg13g2_fill_2 FILLER_58_253 ();
 sg13g2_fill_2 FILLER_58_260 ();
 sg13g2_decap_8 FILLER_58_288 ();
 sg13g2_decap_8 FILLER_58_295 ();
 sg13g2_fill_1 FILLER_58_302 ();
 sg13g2_fill_2 FILLER_58_307 ();
 sg13g2_fill_1 FILLER_58_309 ();
 sg13g2_decap_4 FILLER_58_318 ();
 sg13g2_decap_4 FILLER_58_343 ();
 sg13g2_fill_1 FILLER_58_347 ();
 sg13g2_decap_4 FILLER_58_364 ();
 sg13g2_fill_2 FILLER_58_376 ();
 sg13g2_fill_1 FILLER_58_378 ();
 sg13g2_fill_1 FILLER_58_384 ();
 sg13g2_fill_1 FILLER_58_393 ();
 sg13g2_decap_8 FILLER_58_399 ();
 sg13g2_fill_1 FILLER_58_406 ();
 sg13g2_decap_4 FILLER_58_438 ();
 sg13g2_fill_2 FILLER_58_442 ();
 sg13g2_fill_1 FILLER_58_449 ();
 sg13g2_fill_2 FILLER_58_459 ();
 sg13g2_fill_1 FILLER_58_461 ();
 sg13g2_decap_4 FILLER_58_467 ();
 sg13g2_fill_1 FILLER_58_475 ();
 sg13g2_fill_2 FILLER_58_484 ();
 sg13g2_fill_1 FILLER_58_492 ();
 sg13g2_decap_4 FILLER_58_510 ();
 sg13g2_fill_2 FILLER_58_529 ();
 sg13g2_fill_1 FILLER_58_531 ();
 sg13g2_decap_8 FILLER_58_537 ();
 sg13g2_decap_8 FILLER_58_544 ();
 sg13g2_fill_1 FILLER_58_551 ();
 sg13g2_decap_8 FILLER_58_579 ();
 sg13g2_fill_2 FILLER_58_586 ();
 sg13g2_fill_1 FILLER_58_588 ();
 sg13g2_fill_2 FILLER_58_603 ();
 sg13g2_fill_1 FILLER_58_605 ();
 sg13g2_decap_8 FILLER_58_617 ();
 sg13g2_decap_8 FILLER_58_624 ();
 sg13g2_decap_4 FILLER_58_631 ();
 sg13g2_fill_2 FILLER_58_635 ();
 sg13g2_fill_2 FILLER_58_654 ();
 sg13g2_fill_1 FILLER_58_656 ();
 sg13g2_decap_8 FILLER_58_663 ();
 sg13g2_decap_4 FILLER_58_670 ();
 sg13g2_fill_1 FILLER_58_674 ();
 sg13g2_decap_8 FILLER_58_687 ();
 sg13g2_decap_4 FILLER_58_694 ();
 sg13g2_fill_2 FILLER_58_698 ();
 sg13g2_decap_8 FILLER_58_729 ();
 sg13g2_decap_8 FILLER_58_736 ();
 sg13g2_decap_8 FILLER_58_752 ();
 sg13g2_decap_4 FILLER_58_759 ();
 sg13g2_fill_1 FILLER_58_763 ();
 sg13g2_fill_1 FILLER_58_774 ();
 sg13g2_decap_8 FILLER_58_779 ();
 sg13g2_decap_8 FILLER_58_786 ();
 sg13g2_fill_2 FILLER_58_793 ();
 sg13g2_fill_1 FILLER_58_795 ();
 sg13g2_fill_2 FILLER_58_806 ();
 sg13g2_fill_1 FILLER_58_808 ();
 sg13g2_decap_8 FILLER_58_835 ();
 sg13g2_decap_8 FILLER_58_842 ();
 sg13g2_fill_2 FILLER_58_849 ();
 sg13g2_fill_1 FILLER_58_851 ();
 sg13g2_decap_4 FILLER_58_856 ();
 sg13g2_decap_8 FILLER_58_864 ();
 sg13g2_decap_8 FILLER_58_871 ();
 sg13g2_decap_8 FILLER_59_0 ();
 sg13g2_decap_4 FILLER_59_7 ();
 sg13g2_fill_2 FILLER_59_11 ();
 sg13g2_fill_2 FILLER_59_26 ();
 sg13g2_fill_2 FILLER_59_45 ();
 sg13g2_fill_1 FILLER_59_47 ();
 sg13g2_fill_1 FILLER_59_52 ();
 sg13g2_fill_1 FILLER_59_66 ();
 sg13g2_decap_4 FILLER_59_73 ();
 sg13g2_fill_2 FILLER_59_77 ();
 sg13g2_fill_2 FILLER_59_83 ();
 sg13g2_decap_8 FILLER_59_91 ();
 sg13g2_fill_1 FILLER_59_98 ();
 sg13g2_fill_1 FILLER_59_113 ();
 sg13g2_fill_2 FILLER_59_119 ();
 sg13g2_decap_4 FILLER_59_126 ();
 sg13g2_fill_1 FILLER_59_139 ();
 sg13g2_decap_8 FILLER_59_153 ();
 sg13g2_decap_8 FILLER_59_160 ();
 sg13g2_fill_1 FILLER_59_167 ();
 sg13g2_decap_4 FILLER_59_190 ();
 sg13g2_fill_1 FILLER_59_194 ();
 sg13g2_fill_1 FILLER_59_208 ();
 sg13g2_fill_1 FILLER_59_218 ();
 sg13g2_decap_8 FILLER_59_223 ();
 sg13g2_decap_8 FILLER_59_230 ();
 sg13g2_decap_4 FILLER_59_237 ();
 sg13g2_fill_2 FILLER_59_251 ();
 sg13g2_fill_1 FILLER_59_253 ();
 sg13g2_decap_8 FILLER_59_278 ();
 sg13g2_decap_8 FILLER_59_285 ();
 sg13g2_decap_8 FILLER_59_292 ();
 sg13g2_decap_4 FILLER_59_299 ();
 sg13g2_fill_2 FILLER_59_303 ();
 sg13g2_fill_2 FILLER_59_318 ();
 sg13g2_fill_1 FILLER_59_320 ();
 sg13g2_fill_2 FILLER_59_340 ();
 sg13g2_fill_2 FILLER_59_351 ();
 sg13g2_fill_1 FILLER_59_353 ();
 sg13g2_fill_1 FILLER_59_373 ();
 sg13g2_fill_1 FILLER_59_378 ();
 sg13g2_fill_2 FILLER_59_387 ();
 sg13g2_decap_4 FILLER_59_407 ();
 sg13g2_fill_2 FILLER_59_411 ();
 sg13g2_fill_1 FILLER_59_417 ();
 sg13g2_fill_1 FILLER_59_423 ();
 sg13g2_fill_2 FILLER_59_429 ();
 sg13g2_fill_1 FILLER_59_435 ();
 sg13g2_fill_2 FILLER_59_446 ();
 sg13g2_fill_1 FILLER_59_448 ();
 sg13g2_decap_8 FILLER_59_464 ();
 sg13g2_fill_2 FILLER_59_471 ();
 sg13g2_decap_8 FILLER_59_478 ();
 sg13g2_decap_8 FILLER_59_485 ();
 sg13g2_fill_2 FILLER_59_492 ();
 sg13g2_fill_1 FILLER_59_494 ();
 sg13g2_fill_1 FILLER_59_507 ();
 sg13g2_fill_1 FILLER_59_513 ();
 sg13g2_decap_4 FILLER_59_522 ();
 sg13g2_fill_2 FILLER_59_526 ();
 sg13g2_decap_8 FILLER_59_532 ();
 sg13g2_fill_2 FILLER_59_539 ();
 sg13g2_decap_8 FILLER_59_546 ();
 sg13g2_decap_8 FILLER_59_553 ();
 sg13g2_decap_8 FILLER_59_560 ();
 sg13g2_decap_8 FILLER_59_567 ();
 sg13g2_decap_8 FILLER_59_574 ();
 sg13g2_decap_4 FILLER_59_581 ();
 sg13g2_fill_1 FILLER_59_585 ();
 sg13g2_fill_2 FILLER_59_623 ();
 sg13g2_fill_1 FILLER_59_625 ();
 sg13g2_decap_4 FILLER_59_630 ();
 sg13g2_fill_1 FILLER_59_634 ();
 sg13g2_fill_2 FILLER_59_639 ();
 sg13g2_decap_8 FILLER_59_666 ();
 sg13g2_decap_4 FILLER_59_673 ();
 sg13g2_decap_4 FILLER_59_691 ();
 sg13g2_fill_1 FILLER_59_695 ();
 sg13g2_fill_2 FILLER_59_700 ();
 sg13g2_decap_4 FILLER_59_714 ();
 sg13g2_decap_8 FILLER_59_728 ();
 sg13g2_fill_1 FILLER_59_741 ();
 sg13g2_decap_8 FILLER_59_790 ();
 sg13g2_fill_2 FILLER_59_797 ();
 sg13g2_fill_2 FILLER_59_803 ();
 sg13g2_fill_2 FILLER_59_810 ();
 sg13g2_fill_1 FILLER_59_812 ();
 sg13g2_fill_2 FILLER_59_826 ();
 sg13g2_decap_8 FILLER_59_843 ();
 sg13g2_fill_1 FILLER_59_850 ();
 sg13g2_fill_1 FILLER_59_877 ();
 sg13g2_decap_8 FILLER_60_0 ();
 sg13g2_decap_4 FILLER_60_7 ();
 sg13g2_decap_4 FILLER_60_19 ();
 sg13g2_fill_2 FILLER_60_27 ();
 sg13g2_fill_2 FILLER_60_39 ();
 sg13g2_fill_1 FILLER_60_41 ();
 sg13g2_fill_2 FILLER_60_46 ();
 sg13g2_fill_1 FILLER_60_48 ();
 sg13g2_fill_1 FILLER_60_58 ();
 sg13g2_fill_1 FILLER_60_68 ();
 sg13g2_decap_4 FILLER_60_80 ();
 sg13g2_fill_1 FILLER_60_84 ();
 sg13g2_decap_4 FILLER_60_109 ();
 sg13g2_fill_2 FILLER_60_113 ();
 sg13g2_decap_8 FILLER_60_134 ();
 sg13g2_decap_8 FILLER_60_141 ();
 sg13g2_decap_8 FILLER_60_148 ();
 sg13g2_decap_8 FILLER_60_155 ();
 sg13g2_decap_8 FILLER_60_162 ();
 sg13g2_fill_1 FILLER_60_169 ();
 sg13g2_fill_1 FILLER_60_179 ();
 sg13g2_decap_4 FILLER_60_189 ();
 sg13g2_fill_1 FILLER_60_193 ();
 sg13g2_decap_8 FILLER_60_203 ();
 sg13g2_fill_1 FILLER_60_210 ();
 sg13g2_decap_8 FILLER_60_225 ();
 sg13g2_decap_8 FILLER_60_232 ();
 sg13g2_fill_1 FILLER_60_243 ();
 sg13g2_fill_1 FILLER_60_252 ();
 sg13g2_decap_4 FILLER_60_257 ();
 sg13g2_fill_2 FILLER_60_261 ();
 sg13g2_decap_8 FILLER_60_267 ();
 sg13g2_decap_4 FILLER_60_274 ();
 sg13g2_decap_8 FILLER_60_289 ();
 sg13g2_decap_8 FILLER_60_296 ();
 sg13g2_decap_8 FILLER_60_303 ();
 sg13g2_fill_2 FILLER_60_310 ();
 sg13g2_fill_1 FILLER_60_312 ();
 sg13g2_fill_1 FILLER_60_317 ();
 sg13g2_decap_4 FILLER_60_333 ();
 sg13g2_fill_1 FILLER_60_356 ();
 sg13g2_fill_2 FILLER_60_367 ();
 sg13g2_fill_1 FILLER_60_369 ();
 sg13g2_fill_1 FILLER_60_379 ();
 sg13g2_fill_2 FILLER_60_385 ();
 sg13g2_fill_1 FILLER_60_397 ();
 sg13g2_decap_4 FILLER_60_403 ();
 sg13g2_fill_2 FILLER_60_407 ();
 sg13g2_fill_1 FILLER_60_413 ();
 sg13g2_fill_2 FILLER_60_419 ();
 sg13g2_fill_2 FILLER_60_430 ();
 sg13g2_decap_8 FILLER_60_460 ();
 sg13g2_decap_8 FILLER_60_467 ();
 sg13g2_decap_8 FILLER_60_474 ();
 sg13g2_decap_8 FILLER_60_481 ();
 sg13g2_decap_8 FILLER_60_488 ();
 sg13g2_decap_8 FILLER_60_495 ();
 sg13g2_decap_4 FILLER_60_502 ();
 sg13g2_fill_2 FILLER_60_506 ();
 sg13g2_decap_8 FILLER_60_520 ();
 sg13g2_fill_2 FILLER_60_527 ();
 sg13g2_fill_2 FILLER_60_543 ();
 sg13g2_fill_1 FILLER_60_545 ();
 sg13g2_fill_1 FILLER_60_568 ();
 sg13g2_decap_8 FILLER_60_573 ();
 sg13g2_fill_1 FILLER_60_580 ();
 sg13g2_fill_1 FILLER_60_590 ();
 sg13g2_fill_2 FILLER_60_603 ();
 sg13g2_decap_4 FILLER_60_613 ();
 sg13g2_decap_4 FILLER_60_622 ();
 sg13g2_fill_2 FILLER_60_635 ();
 sg13g2_fill_1 FILLER_60_637 ();
 sg13g2_fill_1 FILLER_60_646 ();
 sg13g2_fill_2 FILLER_60_653 ();
 sg13g2_decap_4 FILLER_60_669 ();
 sg13g2_decap_8 FILLER_60_692 ();
 sg13g2_decap_4 FILLER_60_699 ();
 sg13g2_fill_2 FILLER_60_703 ();
 sg13g2_decap_8 FILLER_60_710 ();
 sg13g2_decap_8 FILLER_60_717 ();
 sg13g2_decap_8 FILLER_60_724 ();
 sg13g2_decap_8 FILLER_60_731 ();
 sg13g2_decap_8 FILLER_60_738 ();
 sg13g2_decap_8 FILLER_60_774 ();
 sg13g2_fill_2 FILLER_60_786 ();
 sg13g2_fill_1 FILLER_60_793 ();
 sg13g2_decap_8 FILLER_60_820 ();
 sg13g2_fill_1 FILLER_60_827 ();
 sg13g2_fill_2 FILLER_60_833 ();
 sg13g2_fill_1 FILLER_60_840 ();
 sg13g2_decap_8 FILLER_60_867 ();
 sg13g2_decap_4 FILLER_60_874 ();
 sg13g2_decap_8 FILLER_61_0 ();
 sg13g2_decap_8 FILLER_61_7 ();
 sg13g2_fill_1 FILLER_61_22 ();
 sg13g2_fill_2 FILLER_61_43 ();
 sg13g2_fill_1 FILLER_61_45 ();
 sg13g2_fill_1 FILLER_61_59 ();
 sg13g2_fill_2 FILLER_61_74 ();
 sg13g2_decap_4 FILLER_61_81 ();
 sg13g2_fill_1 FILLER_61_85 ();
 sg13g2_fill_2 FILLER_61_97 ();
 sg13g2_fill_1 FILLER_61_104 ();
 sg13g2_fill_1 FILLER_61_111 ();
 sg13g2_fill_1 FILLER_61_121 ();
 sg13g2_fill_1 FILLER_61_128 ();
 sg13g2_decap_4 FILLER_61_139 ();
 sg13g2_fill_1 FILLER_61_143 ();
 sg13g2_decap_8 FILLER_61_149 ();
 sg13g2_decap_8 FILLER_61_156 ();
 sg13g2_fill_1 FILLER_61_167 ();
 sg13g2_decap_4 FILLER_61_174 ();
 sg13g2_decap_8 FILLER_61_183 ();
 sg13g2_fill_2 FILLER_61_190 ();
 sg13g2_decap_4 FILLER_61_197 ();
 sg13g2_decap_8 FILLER_61_206 ();
 sg13g2_decap_8 FILLER_61_213 ();
 sg13g2_fill_2 FILLER_61_220 ();
 sg13g2_decap_8 FILLER_61_226 ();
 sg13g2_fill_1 FILLER_61_233 ();
 sg13g2_decap_8 FILLER_61_271 ();
 sg13g2_decap_8 FILLER_61_278 ();
 sg13g2_fill_1 FILLER_61_285 ();
 sg13g2_decap_8 FILLER_61_290 ();
 sg13g2_decap_4 FILLER_61_297 ();
 sg13g2_fill_1 FILLER_61_305 ();
 sg13g2_decap_4 FILLER_61_315 ();
 sg13g2_decap_8 FILLER_61_332 ();
 sg13g2_decap_4 FILLER_61_339 ();
 sg13g2_fill_1 FILLER_61_343 ();
 sg13g2_fill_2 FILLER_61_349 ();
 sg13g2_fill_2 FILLER_61_382 ();
 sg13g2_decap_4 FILLER_61_402 ();
 sg13g2_fill_2 FILLER_61_416 ();
 sg13g2_decap_8 FILLER_61_432 ();
 sg13g2_decap_8 FILLER_61_452 ();
 sg13g2_decap_8 FILLER_61_459 ();
 sg13g2_fill_1 FILLER_61_466 ();
 sg13g2_decap_8 FILLER_61_476 ();
 sg13g2_decap_8 FILLER_61_483 ();
 sg13g2_decap_8 FILLER_61_490 ();
 sg13g2_decap_8 FILLER_61_497 ();
 sg13g2_decap_8 FILLER_61_504 ();
 sg13g2_decap_4 FILLER_61_511 ();
 sg13g2_fill_1 FILLER_61_515 ();
 sg13g2_fill_2 FILLER_61_535 ();
 sg13g2_decap_8 FILLER_61_541 ();
 sg13g2_decap_8 FILLER_61_548 ();
 sg13g2_fill_2 FILLER_61_555 ();
 sg13g2_fill_1 FILLER_61_557 ();
 sg13g2_fill_2 FILLER_61_570 ();
 sg13g2_fill_2 FILLER_61_578 ();
 sg13g2_fill_1 FILLER_61_580 ();
 sg13g2_fill_1 FILLER_61_586 ();
 sg13g2_fill_2 FILLER_61_594 ();
 sg13g2_fill_1 FILLER_61_604 ();
 sg13g2_fill_1 FILLER_61_610 ();
 sg13g2_decap_8 FILLER_61_616 ();
 sg13g2_decap_8 FILLER_61_623 ();
 sg13g2_decap_4 FILLER_61_630 ();
 sg13g2_fill_1 FILLER_61_634 ();
 sg13g2_decap_4 FILLER_61_643 ();
 sg13g2_decap_8 FILLER_61_652 ();
 sg13g2_decap_8 FILLER_61_659 ();
 sg13g2_fill_1 FILLER_61_666 ();
 sg13g2_decap_8 FILLER_61_680 ();
 sg13g2_decap_8 FILLER_61_687 ();
 sg13g2_decap_8 FILLER_61_694 ();
 sg13g2_fill_2 FILLER_61_747 ();
 sg13g2_fill_2 FILLER_61_755 ();
 sg13g2_fill_1 FILLER_61_757 ();
 sg13g2_fill_2 FILLER_61_768 ();
 sg13g2_fill_1 FILLER_61_770 ();
 sg13g2_decap_4 FILLER_61_801 ();
 sg13g2_fill_2 FILLER_61_805 ();
 sg13g2_fill_2 FILLER_61_826 ();
 sg13g2_decap_8 FILLER_61_832 ();
 sg13g2_fill_2 FILLER_61_843 ();
 sg13g2_fill_2 FILLER_61_848 ();
 sg13g2_fill_2 FILLER_61_857 ();
 sg13g2_decap_4 FILLER_61_872 ();
 sg13g2_fill_2 FILLER_61_876 ();
 sg13g2_decap_8 FILLER_62_0 ();
 sg13g2_decap_8 FILLER_62_7 ();
 sg13g2_fill_1 FILLER_62_14 ();
 sg13g2_decap_8 FILLER_62_20 ();
 sg13g2_fill_2 FILLER_62_27 ();
 sg13g2_fill_1 FILLER_62_35 ();
 sg13g2_fill_1 FILLER_62_40 ();
 sg13g2_fill_2 FILLER_62_46 ();
 sg13g2_fill_1 FILLER_62_48 ();
 sg13g2_fill_2 FILLER_62_60 ();
 sg13g2_fill_2 FILLER_62_67 ();
 sg13g2_fill_1 FILLER_62_77 ();
 sg13g2_fill_2 FILLER_62_86 ();
 sg13g2_fill_2 FILLER_62_97 ();
 sg13g2_fill_2 FILLER_62_104 ();
 sg13g2_fill_1 FILLER_62_119 ();
 sg13g2_fill_1 FILLER_62_129 ();
 sg13g2_decap_8 FILLER_62_134 ();
 sg13g2_fill_2 FILLER_62_141 ();
 sg13g2_fill_1 FILLER_62_153 ();
 sg13g2_fill_1 FILLER_62_165 ();
 sg13g2_decap_8 FILLER_62_170 ();
 sg13g2_decap_8 FILLER_62_177 ();
 sg13g2_decap_8 FILLER_62_184 ();
 sg13g2_fill_2 FILLER_62_191 ();
 sg13g2_decap_8 FILLER_62_213 ();
 sg13g2_decap_8 FILLER_62_220 ();
 sg13g2_decap_8 FILLER_62_227 ();
 sg13g2_decap_8 FILLER_62_234 ();
 sg13g2_fill_2 FILLER_62_241 ();
 sg13g2_fill_1 FILLER_62_243 ();
 sg13g2_decap_8 FILLER_62_249 ();
 sg13g2_fill_2 FILLER_62_261 ();
 sg13g2_fill_1 FILLER_62_263 ();
 sg13g2_fill_1 FILLER_62_276 ();
 sg13g2_decap_4 FILLER_62_283 ();
 sg13g2_fill_1 FILLER_62_287 ();
 sg13g2_fill_2 FILLER_62_292 ();
 sg13g2_fill_1 FILLER_62_324 ();
 sg13g2_decap_8 FILLER_62_333 ();
 sg13g2_decap_8 FILLER_62_340 ();
 sg13g2_fill_2 FILLER_62_347 ();
 sg13g2_fill_1 FILLER_62_349 ();
 sg13g2_decap_8 FILLER_62_354 ();
 sg13g2_decap_8 FILLER_62_375 ();
 sg13g2_decap_4 FILLER_62_382 ();
 sg13g2_fill_2 FILLER_62_386 ();
 sg13g2_decap_8 FILLER_62_393 ();
 sg13g2_decap_8 FILLER_62_400 ();
 sg13g2_decap_8 FILLER_62_407 ();
 sg13g2_decap_4 FILLER_62_414 ();
 sg13g2_decap_8 FILLER_62_423 ();
 sg13g2_decap_8 FILLER_62_430 ();
 sg13g2_decap_8 FILLER_62_437 ();
 sg13g2_decap_8 FILLER_62_444 ();
 sg13g2_decap_8 FILLER_62_451 ();
 sg13g2_decap_4 FILLER_62_458 ();
 sg13g2_fill_1 FILLER_62_466 ();
 sg13g2_decap_8 FILLER_62_471 ();
 sg13g2_decap_8 FILLER_62_478 ();
 sg13g2_decap_8 FILLER_62_485 ();
 sg13g2_decap_4 FILLER_62_492 ();
 sg13g2_fill_2 FILLER_62_496 ();
 sg13g2_fill_1 FILLER_62_507 ();
 sg13g2_decap_4 FILLER_62_515 ();
 sg13g2_fill_1 FILLER_62_519 ();
 sg13g2_decap_4 FILLER_62_530 ();
 sg13g2_fill_2 FILLER_62_534 ();
 sg13g2_fill_1 FILLER_62_541 ();
 sg13g2_decap_8 FILLER_62_547 ();
 sg13g2_decap_8 FILLER_62_554 ();
 sg13g2_fill_2 FILLER_62_561 ();
 sg13g2_fill_1 FILLER_62_563 ();
 sg13g2_decap_4 FILLER_62_573 ();
 sg13g2_fill_2 FILLER_62_581 ();
 sg13g2_fill_1 FILLER_62_583 ();
 sg13g2_fill_2 FILLER_62_588 ();
 sg13g2_fill_1 FILLER_62_590 ();
 sg13g2_decap_8 FILLER_62_609 ();
 sg13g2_fill_2 FILLER_62_616 ();
 sg13g2_fill_1 FILLER_62_618 ();
 sg13g2_decap_8 FILLER_62_628 ();
 sg13g2_decap_8 FILLER_62_635 ();
 sg13g2_decap_8 FILLER_62_642 ();
 sg13g2_decap_8 FILLER_62_649 ();
 sg13g2_decap_8 FILLER_62_656 ();
 sg13g2_decap_4 FILLER_62_663 ();
 sg13g2_decap_4 FILLER_62_698 ();
 sg13g2_fill_2 FILLER_62_712 ();
 sg13g2_decap_8 FILLER_62_726 ();
 sg13g2_fill_2 FILLER_62_733 ();
 sg13g2_decap_8 FILLER_62_739 ();
 sg13g2_fill_2 FILLER_62_746 ();
 sg13g2_fill_2 FILLER_62_754 ();
 sg13g2_decap_8 FILLER_62_760 ();
 sg13g2_decap_4 FILLER_62_772 ();
 sg13g2_fill_1 FILLER_62_776 ();
 sg13g2_decap_8 FILLER_62_781 ();
 sg13g2_decap_8 FILLER_62_788 ();
 sg13g2_decap_8 FILLER_62_795 ();
 sg13g2_fill_2 FILLER_62_838 ();
 sg13g2_fill_2 FILLER_62_850 ();
 sg13g2_decap_8 FILLER_63_0 ();
 sg13g2_decap_8 FILLER_63_7 ();
 sg13g2_fill_1 FILLER_63_14 ();
 sg13g2_fill_2 FILLER_63_32 ();
 sg13g2_fill_2 FILLER_63_39 ();
 sg13g2_fill_2 FILLER_63_51 ();
 sg13g2_fill_2 FILLER_63_57 ();
 sg13g2_fill_1 FILLER_63_59 ();
 sg13g2_fill_2 FILLER_63_68 ();
 sg13g2_decap_4 FILLER_63_74 ();
 sg13g2_fill_1 FILLER_63_88 ();
 sg13g2_fill_2 FILLER_63_98 ();
 sg13g2_fill_1 FILLER_63_100 ();
 sg13g2_fill_1 FILLER_63_113 ();
 sg13g2_fill_1 FILLER_63_123 ();
 sg13g2_fill_1 FILLER_63_140 ();
 sg13g2_decap_4 FILLER_63_145 ();
 sg13g2_decap_4 FILLER_63_154 ();
 sg13g2_fill_2 FILLER_63_158 ();
 sg13g2_fill_1 FILLER_63_169 ();
 sg13g2_decap_4 FILLER_63_174 ();
 sg13g2_decap_8 FILLER_63_184 ();
 sg13g2_decap_8 FILLER_63_191 ();
 sg13g2_decap_8 FILLER_63_198 ();
 sg13g2_decap_8 FILLER_63_205 ();
 sg13g2_decap_8 FILLER_63_212 ();
 sg13g2_decap_4 FILLER_63_219 ();
 sg13g2_decap_8 FILLER_63_227 ();
 sg13g2_decap_4 FILLER_63_234 ();
 sg13g2_fill_2 FILLER_63_238 ();
 sg13g2_fill_1 FILLER_63_266 ();
 sg13g2_fill_1 FILLER_63_277 ();
 sg13g2_decap_8 FILLER_63_284 ();
 sg13g2_decap_8 FILLER_63_291 ();
 sg13g2_fill_2 FILLER_63_298 ();
 sg13g2_fill_1 FILLER_63_300 ();
 sg13g2_fill_1 FILLER_63_306 ();
 sg13g2_decap_8 FILLER_63_311 ();
 sg13g2_decap_4 FILLER_63_318 ();
 sg13g2_fill_1 FILLER_63_322 ();
 sg13g2_decap_4 FILLER_63_334 ();
 sg13g2_decap_8 FILLER_63_343 ();
 sg13g2_decap_8 FILLER_63_350 ();
 sg13g2_decap_8 FILLER_63_357 ();
 sg13g2_decap_8 FILLER_63_364 ();
 sg13g2_decap_4 FILLER_63_371 ();
 sg13g2_decap_8 FILLER_63_400 ();
 sg13g2_fill_2 FILLER_63_407 ();
 sg13g2_fill_1 FILLER_63_423 ();
 sg13g2_decap_4 FILLER_63_429 ();
 sg13g2_decap_4 FILLER_63_453 ();
 sg13g2_fill_1 FILLER_63_457 ();
 sg13g2_decap_8 FILLER_63_472 ();
 sg13g2_decap_8 FILLER_63_479 ();
 sg13g2_fill_2 FILLER_63_486 ();
 sg13g2_fill_1 FILLER_63_488 ();
 sg13g2_fill_1 FILLER_63_493 ();
 sg13g2_fill_2 FILLER_63_502 ();
 sg13g2_fill_1 FILLER_63_504 ();
 sg13g2_fill_1 FILLER_63_523 ();
 sg13g2_decap_8 FILLER_63_548 ();
 sg13g2_decap_8 FILLER_63_555 ();
 sg13g2_decap_4 FILLER_63_562 ();
 sg13g2_fill_2 FILLER_63_566 ();
 sg13g2_decap_4 FILLER_63_572 ();
 sg13g2_fill_2 FILLER_63_601 ();
 sg13g2_fill_1 FILLER_63_614 ();
 sg13g2_fill_2 FILLER_63_621 ();
 sg13g2_fill_1 FILLER_63_633 ();
 sg13g2_decap_8 FILLER_63_639 ();
 sg13g2_fill_2 FILLER_63_655 ();
 sg13g2_fill_1 FILLER_63_657 ();
 sg13g2_fill_2 FILLER_63_664 ();
 sg13g2_decap_4 FILLER_63_671 ();
 sg13g2_fill_2 FILLER_63_679 ();
 sg13g2_decap_8 FILLER_63_686 ();
 sg13g2_decap_8 FILLER_63_693 ();
 sg13g2_fill_2 FILLER_63_700 ();
 sg13g2_fill_1 FILLER_63_702 ();
 sg13g2_fill_1 FILLER_63_707 ();
 sg13g2_fill_2 FILLER_63_712 ();
 sg13g2_decap_8 FILLER_63_718 ();
 sg13g2_decap_8 FILLER_63_725 ();
 sg13g2_fill_2 FILLER_63_732 ();
 sg13g2_fill_1 FILLER_63_740 ();
 sg13g2_decap_8 FILLER_63_749 ();
 sg13g2_decap_8 FILLER_63_756 ();
 sg13g2_decap_8 FILLER_63_763 ();
 sg13g2_decap_4 FILLER_63_806 ();
 sg13g2_decap_8 FILLER_63_819 ();
 sg13g2_decap_8 FILLER_63_826 ();
 sg13g2_decap_8 FILLER_63_833 ();
 sg13g2_decap_4 FILLER_63_840 ();
 sg13g2_decap_8 FILLER_63_867 ();
 sg13g2_decap_4 FILLER_63_874 ();
 sg13g2_decap_8 FILLER_64_0 ();
 sg13g2_decap_8 FILLER_64_7 ();
 sg13g2_decap_4 FILLER_64_14 ();
 sg13g2_fill_2 FILLER_64_18 ();
 sg13g2_decap_4 FILLER_64_25 ();
 sg13g2_fill_1 FILLER_64_29 ();
 sg13g2_decap_4 FILLER_64_45 ();
 sg13g2_fill_1 FILLER_64_49 ();
 sg13g2_decap_4 FILLER_64_55 ();
 sg13g2_decap_8 FILLER_64_64 ();
 sg13g2_decap_8 FILLER_64_71 ();
 sg13g2_fill_2 FILLER_64_78 ();
 sg13g2_fill_1 FILLER_64_80 ();
 sg13g2_decap_8 FILLER_64_91 ();
 sg13g2_fill_2 FILLER_64_108 ();
 sg13g2_decap_8 FILLER_64_114 ();
 sg13g2_decap_4 FILLER_64_121 ();
 sg13g2_fill_2 FILLER_64_125 ();
 sg13g2_fill_1 FILLER_64_136 ();
 sg13g2_fill_2 FILLER_64_143 ();
 sg13g2_fill_2 FILLER_64_150 ();
 sg13g2_decap_8 FILLER_64_184 ();
 sg13g2_decap_4 FILLER_64_191 ();
 sg13g2_fill_2 FILLER_64_195 ();
 sg13g2_decap_4 FILLER_64_207 ();
 sg13g2_fill_2 FILLER_64_214 ();
 sg13g2_fill_1 FILLER_64_216 ();
 sg13g2_decap_8 FILLER_64_223 ();
 sg13g2_decap_8 FILLER_64_230 ();
 sg13g2_fill_1 FILLER_64_249 ();
 sg13g2_decap_8 FILLER_64_254 ();
 sg13g2_decap_8 FILLER_64_269 ();
 sg13g2_decap_8 FILLER_64_276 ();
 sg13g2_decap_8 FILLER_64_283 ();
 sg13g2_decap_4 FILLER_64_290 ();
 sg13g2_decap_8 FILLER_64_313 ();
 sg13g2_fill_2 FILLER_64_320 ();
 sg13g2_fill_1 FILLER_64_322 ();
 sg13g2_decap_8 FILLER_64_339 ();
 sg13g2_decap_8 FILLER_64_346 ();
 sg13g2_decap_4 FILLER_64_353 ();
 sg13g2_fill_2 FILLER_64_390 ();
 sg13g2_fill_1 FILLER_64_392 ();
 sg13g2_decap_4 FILLER_64_402 ();
 sg13g2_fill_2 FILLER_64_411 ();
 sg13g2_decap_8 FILLER_64_423 ();
 sg13g2_decap_8 FILLER_64_430 ();
 sg13g2_decap_8 FILLER_64_437 ();
 sg13g2_decap_4 FILLER_64_454 ();
 sg13g2_fill_1 FILLER_64_474 ();
 sg13g2_decap_8 FILLER_64_485 ();
 sg13g2_decap_4 FILLER_64_492 ();
 sg13g2_fill_1 FILLER_64_496 ();
 sg13g2_decap_8 FILLER_64_533 ();
 sg13g2_decap_8 FILLER_64_540 ();
 sg13g2_decap_8 FILLER_64_547 ();
 sg13g2_decap_8 FILLER_64_554 ();
 sg13g2_decap_8 FILLER_64_561 ();
 sg13g2_decap_4 FILLER_64_568 ();
 sg13g2_decap_8 FILLER_64_581 ();
 sg13g2_decap_4 FILLER_64_588 ();
 sg13g2_fill_2 FILLER_64_598 ();
 sg13g2_decap_4 FILLER_64_604 ();
 sg13g2_fill_1 FILLER_64_608 ();
 sg13g2_fill_1 FILLER_64_623 ();
 sg13g2_decap_8 FILLER_64_629 ();
 sg13g2_decap_8 FILLER_64_636 ();
 sg13g2_decap_8 FILLER_64_643 ();
 sg13g2_decap_8 FILLER_64_650 ();
 sg13g2_decap_4 FILLER_64_657 ();
 sg13g2_decap_4 FILLER_64_697 ();
 sg13g2_fill_1 FILLER_64_701 ();
 sg13g2_decap_4 FILLER_64_707 ();
 sg13g2_fill_1 FILLER_64_711 ();
 sg13g2_fill_1 FILLER_64_727 ();
 sg13g2_decap_4 FILLER_64_733 ();
 sg13g2_fill_2 FILLER_64_773 ();
 sg13g2_fill_1 FILLER_64_775 ();
 sg13g2_fill_1 FILLER_64_781 ();
 sg13g2_fill_1 FILLER_64_787 ();
 sg13g2_fill_2 FILLER_64_797 ();
 sg13g2_decap_8 FILLER_64_805 ();
 sg13g2_decap_8 FILLER_64_812 ();
 sg13g2_decap_8 FILLER_64_823 ();
 sg13g2_fill_2 FILLER_64_834 ();
 sg13g2_fill_1 FILLER_64_849 ();
 sg13g2_fill_2 FILLER_64_876 ();
 sg13g2_decap_8 FILLER_65_0 ();
 sg13g2_decap_8 FILLER_65_7 ();
 sg13g2_fill_2 FILLER_65_14 ();
 sg13g2_fill_2 FILLER_65_20 ();
 sg13g2_decap_4 FILLER_65_32 ();
 sg13g2_decap_8 FILLER_65_50 ();
 sg13g2_fill_2 FILLER_65_62 ();
 sg13g2_decap_4 FILLER_65_82 ();
 sg13g2_decap_4 FILLER_65_96 ();
 sg13g2_decap_4 FILLER_65_113 ();
 sg13g2_fill_2 FILLER_65_117 ();
 sg13g2_decap_8 FILLER_65_124 ();
 sg13g2_fill_1 FILLER_65_136 ();
 sg13g2_fill_1 FILLER_65_145 ();
 sg13g2_fill_1 FILLER_65_156 ();
 sg13g2_fill_1 FILLER_65_180 ();
 sg13g2_fill_2 FILLER_65_186 ();
 sg13g2_fill_1 FILLER_65_192 ();
 sg13g2_fill_2 FILLER_65_202 ();
 sg13g2_fill_2 FILLER_65_209 ();
 sg13g2_fill_1 FILLER_65_211 ();
 sg13g2_decap_8 FILLER_65_223 ();
 sg13g2_fill_2 FILLER_65_230 ();
 sg13g2_fill_1 FILLER_65_232 ();
 sg13g2_fill_2 FILLER_65_267 ();
 sg13g2_fill_1 FILLER_65_269 ();
 sg13g2_fill_1 FILLER_65_274 ();
 sg13g2_decap_4 FILLER_65_283 ();
 sg13g2_fill_2 FILLER_65_287 ();
 sg13g2_decap_4 FILLER_65_297 ();
 sg13g2_decap_4 FILLER_65_308 ();
 sg13g2_fill_1 FILLER_65_312 ();
 sg13g2_decap_4 FILLER_65_317 ();
 sg13g2_decap_8 FILLER_65_333 ();
 sg13g2_fill_2 FILLER_65_340 ();
 sg13g2_fill_1 FILLER_65_342 ();
 sg13g2_decap_8 FILLER_65_374 ();
 sg13g2_fill_2 FILLER_65_381 ();
 sg13g2_fill_1 FILLER_65_383 ();
 sg13g2_decap_8 FILLER_65_388 ();
 sg13g2_fill_1 FILLER_65_395 ();
 sg13g2_decap_8 FILLER_65_400 ();
 sg13g2_decap_4 FILLER_65_407 ();
 sg13g2_fill_2 FILLER_65_411 ();
 sg13g2_fill_2 FILLER_65_432 ();
 sg13g2_fill_1 FILLER_65_434 ();
 sg13g2_fill_2 FILLER_65_448 ();
 sg13g2_fill_1 FILLER_65_450 ();
 sg13g2_decap_8 FILLER_65_455 ();
 sg13g2_decap_4 FILLER_65_473 ();
 sg13g2_fill_2 FILLER_65_481 ();
 sg13g2_fill_2 FILLER_65_493 ();
 sg13g2_fill_1 FILLER_65_495 ();
 sg13g2_decap_8 FILLER_65_506 ();
 sg13g2_fill_2 FILLER_65_513 ();
 sg13g2_fill_1 FILLER_65_515 ();
 sg13g2_decap_8 FILLER_65_524 ();
 sg13g2_decap_4 FILLER_65_531 ();
 sg13g2_decap_8 FILLER_65_545 ();
 sg13g2_decap_8 FILLER_65_552 ();
 sg13g2_decap_8 FILLER_65_559 ();
 sg13g2_decap_4 FILLER_65_566 ();
 sg13g2_fill_2 FILLER_65_579 ();
 sg13g2_fill_1 FILLER_65_581 ();
 sg13g2_fill_1 FILLER_65_587 ();
 sg13g2_fill_1 FILLER_65_593 ();
 sg13g2_fill_1 FILLER_65_600 ();
 sg13g2_fill_1 FILLER_65_606 ();
 sg13g2_fill_1 FILLER_65_611 ();
 sg13g2_decap_8 FILLER_65_629 ();
 sg13g2_decap_4 FILLER_65_636 ();
 sg13g2_fill_2 FILLER_65_640 ();
 sg13g2_decap_8 FILLER_65_646 ();
 sg13g2_decap_8 FILLER_65_653 ();
 sg13g2_decap_8 FILLER_65_660 ();
 sg13g2_decap_8 FILLER_65_667 ();
 sg13g2_fill_2 FILLER_65_674 ();
 sg13g2_fill_1 FILLER_65_676 ();
 sg13g2_decap_4 FILLER_65_686 ();
 sg13g2_decap_4 FILLER_65_694 ();
 sg13g2_fill_1 FILLER_65_702 ();
 sg13g2_decap_8 FILLER_65_715 ();
 sg13g2_decap_8 FILLER_65_722 ();
 sg13g2_decap_8 FILLER_65_729 ();
 sg13g2_decap_8 FILLER_65_736 ();
 sg13g2_fill_1 FILLER_65_743 ();
 sg13g2_fill_2 FILLER_65_752 ();
 sg13g2_decap_4 FILLER_65_758 ();
 sg13g2_fill_2 FILLER_65_783 ();
 sg13g2_decap_8 FILLER_65_791 ();
 sg13g2_fill_2 FILLER_65_798 ();
 sg13g2_fill_1 FILLER_65_836 ();
 sg13g2_fill_2 FILLER_65_875 ();
 sg13g2_fill_1 FILLER_65_877 ();
 sg13g2_decap_4 FILLER_66_0 ();
 sg13g2_fill_2 FILLER_66_4 ();
 sg13g2_decap_8 FILLER_66_15 ();
 sg13g2_fill_1 FILLER_66_32 ();
 sg13g2_fill_2 FILLER_66_47 ();
 sg13g2_fill_1 FILLER_66_49 ();
 sg13g2_decap_8 FILLER_66_69 ();
 sg13g2_fill_1 FILLER_66_76 ();
 sg13g2_decap_8 FILLER_66_100 ();
 sg13g2_fill_2 FILLER_66_107 ();
 sg13g2_fill_2 FILLER_66_115 ();
 sg13g2_fill_1 FILLER_66_117 ();
 sg13g2_fill_2 FILLER_66_143 ();
 sg13g2_fill_1 FILLER_66_145 ();
 sg13g2_fill_1 FILLER_66_158 ();
 sg13g2_decap_8 FILLER_66_164 ();
 sg13g2_decap_8 FILLER_66_171 ();
 sg13g2_decap_8 FILLER_66_178 ();
 sg13g2_decap_4 FILLER_66_185 ();
 sg13g2_fill_1 FILLER_66_202 ();
 sg13g2_decap_8 FILLER_66_208 ();
 sg13g2_decap_8 FILLER_66_224 ();
 sg13g2_decap_4 FILLER_66_231 ();
 sg13g2_fill_1 FILLER_66_235 ();
 sg13g2_fill_2 FILLER_66_244 ();
 sg13g2_fill_2 FILLER_66_250 ();
 sg13g2_fill_1 FILLER_66_252 ();
 sg13g2_decap_4 FILLER_66_260 ();
 sg13g2_fill_2 FILLER_66_276 ();
 sg13g2_fill_1 FILLER_66_278 ();
 sg13g2_decap_8 FILLER_66_292 ();
 sg13g2_decap_8 FILLER_66_299 ();
 sg13g2_fill_1 FILLER_66_310 ();
 sg13g2_fill_1 FILLER_66_320 ();
 sg13g2_decap_8 FILLER_66_333 ();
 sg13g2_fill_2 FILLER_66_340 ();
 sg13g2_fill_2 FILLER_66_347 ();
 sg13g2_decap_8 FILLER_66_353 ();
 sg13g2_decap_8 FILLER_66_360 ();
 sg13g2_decap_8 FILLER_66_367 ();
 sg13g2_decap_4 FILLER_66_374 ();
 sg13g2_fill_2 FILLER_66_378 ();
 sg13g2_decap_8 FILLER_66_409 ();
 sg13g2_decap_8 FILLER_66_416 ();
 sg13g2_decap_4 FILLER_66_423 ();
 sg13g2_decap_8 FILLER_66_462 ();
 sg13g2_fill_2 FILLER_66_469 ();
 sg13g2_decap_4 FILLER_66_493 ();
 sg13g2_fill_1 FILLER_66_501 ();
 sg13g2_decap_8 FILLER_66_511 ();
 sg13g2_decap_4 FILLER_66_518 ();
 sg13g2_fill_1 FILLER_66_522 ();
 sg13g2_decap_4 FILLER_66_533 ();
 sg13g2_fill_1 FILLER_66_548 ();
 sg13g2_fill_2 FILLER_66_553 ();
 sg13g2_decap_8 FILLER_66_560 ();
 sg13g2_fill_1 FILLER_66_567 ();
 sg13g2_decap_8 FILLER_66_579 ();
 sg13g2_decap_4 FILLER_66_586 ();
 sg13g2_decap_8 FILLER_66_595 ();
 sg13g2_decap_8 FILLER_66_602 ();
 sg13g2_decap_4 FILLER_66_609 ();
 sg13g2_decap_8 FILLER_66_618 ();
 sg13g2_fill_2 FILLER_66_625 ();
 sg13g2_fill_1 FILLER_66_627 ();
 sg13g2_decap_8 FILLER_66_642 ();
 sg13g2_decap_8 FILLER_66_649 ();
 sg13g2_decap_4 FILLER_66_656 ();
 sg13g2_fill_2 FILLER_66_660 ();
 sg13g2_fill_2 FILLER_66_691 ();
 sg13g2_fill_1 FILLER_66_697 ();
 sg13g2_fill_2 FILLER_66_711 ();
 sg13g2_fill_2 FILLER_66_718 ();
 sg13g2_fill_1 FILLER_66_720 ();
 sg13g2_fill_2 FILLER_66_725 ();
 sg13g2_fill_1 FILLER_66_731 ();
 sg13g2_decap_4 FILLER_66_737 ();
 sg13g2_decap_8 FILLER_66_758 ();
 sg13g2_decap_8 FILLER_66_791 ();
 sg13g2_fill_2 FILLER_66_798 ();
 sg13g2_decap_8 FILLER_66_806 ();
 sg13g2_fill_2 FILLER_66_813 ();
 sg13g2_fill_1 FILLER_66_815 ();
 sg13g2_decap_8 FILLER_66_820 ();
 sg13g2_decap_4 FILLER_66_827 ();
 sg13g2_fill_2 FILLER_66_831 ();
 sg13g2_fill_2 FILLER_66_840 ();
 sg13g2_decap_8 FILLER_66_855 ();
 sg13g2_decap_8 FILLER_66_862 ();
 sg13g2_decap_8 FILLER_66_869 ();
 sg13g2_fill_2 FILLER_66_876 ();
 sg13g2_decap_8 FILLER_67_0 ();
 sg13g2_decap_4 FILLER_67_7 ();
 sg13g2_fill_1 FILLER_67_11 ();
 sg13g2_fill_2 FILLER_67_51 ();
 sg13g2_fill_1 FILLER_67_57 ();
 sg13g2_fill_2 FILLER_67_63 ();
 sg13g2_decap_8 FILLER_67_76 ();
 sg13g2_fill_1 FILLER_67_83 ();
 sg13g2_decap_4 FILLER_67_112 ();
 sg13g2_fill_2 FILLER_67_116 ();
 sg13g2_decap_4 FILLER_67_134 ();
 sg13g2_decap_4 FILLER_67_142 ();
 sg13g2_fill_1 FILLER_67_151 ();
 sg13g2_fill_1 FILLER_67_159 ();
 sg13g2_decap_4 FILLER_67_177 ();
 sg13g2_fill_1 FILLER_67_181 ();
 sg13g2_fill_1 FILLER_67_186 ();
 sg13g2_fill_2 FILLER_67_192 ();
 sg13g2_fill_2 FILLER_67_199 ();
 sg13g2_fill_1 FILLER_67_201 ();
 sg13g2_decap_4 FILLER_67_219 ();
 sg13g2_fill_1 FILLER_67_223 ();
 sg13g2_decap_8 FILLER_67_230 ();
 sg13g2_decap_4 FILLER_67_241 ();
 sg13g2_fill_1 FILLER_67_245 ();
 sg13g2_fill_2 FILLER_67_262 ();
 sg13g2_fill_1 FILLER_67_264 ();
 sg13g2_fill_2 FILLER_67_285 ();
 sg13g2_fill_2 FILLER_67_325 ();
 sg13g2_fill_1 FILLER_67_353 ();
 sg13g2_decap_8 FILLER_67_359 ();
 sg13g2_decap_8 FILLER_67_395 ();
 sg13g2_decap_8 FILLER_67_426 ();
 sg13g2_decap_4 FILLER_67_448 ();
 sg13g2_fill_2 FILLER_67_452 ();
 sg13g2_decap_4 FILLER_67_458 ();
 sg13g2_fill_2 FILLER_67_462 ();
 sg13g2_fill_2 FILLER_67_475 ();
 sg13g2_fill_1 FILLER_67_477 ();
 sg13g2_decap_8 FILLER_67_491 ();
 sg13g2_decap_8 FILLER_67_498 ();
 sg13g2_decap_8 FILLER_67_515 ();
 sg13g2_decap_4 FILLER_67_533 ();
 sg13g2_decap_8 FILLER_67_543 ();
 sg13g2_decap_8 FILLER_67_550 ();
 sg13g2_fill_1 FILLER_67_566 ();
 sg13g2_decap_8 FILLER_67_571 ();
 sg13g2_fill_2 FILLER_67_586 ();
 sg13g2_fill_1 FILLER_67_588 ();
 sg13g2_fill_1 FILLER_67_600 ();
 sg13g2_fill_2 FILLER_67_606 ();
 sg13g2_fill_1 FILLER_67_611 ();
 sg13g2_fill_2 FILLER_67_617 ();
 sg13g2_fill_1 FILLER_67_623 ();
 sg13g2_decap_8 FILLER_67_644 ();
 sg13g2_decap_8 FILLER_67_651 ();
 sg13g2_fill_2 FILLER_67_658 ();
 sg13g2_fill_1 FILLER_67_660 ();
 sg13g2_fill_2 FILLER_67_673 ();
 sg13g2_decap_4 FILLER_67_680 ();
 sg13g2_fill_1 FILLER_67_684 ();
 sg13g2_fill_2 FILLER_67_721 ();
 sg13g2_fill_1 FILLER_67_723 ();
 sg13g2_decap_4 FILLER_67_736 ();
 sg13g2_decap_4 FILLER_67_752 ();
 sg13g2_fill_1 FILLER_67_756 ();
 sg13g2_decap_4 FILLER_67_765 ();
 sg13g2_fill_1 FILLER_67_769 ();
 sg13g2_decap_8 FILLER_67_774 ();
 sg13g2_decap_8 FILLER_67_781 ();
 sg13g2_decap_8 FILLER_67_788 ();
 sg13g2_decap_4 FILLER_67_795 ();
 sg13g2_fill_1 FILLER_67_840 ();
 sg13g2_fill_2 FILLER_67_875 ();
 sg13g2_fill_1 FILLER_67_877 ();
 sg13g2_decap_8 FILLER_68_0 ();
 sg13g2_decap_8 FILLER_68_7 ();
 sg13g2_fill_2 FILLER_68_14 ();
 sg13g2_fill_2 FILLER_68_35 ();
 sg13g2_fill_2 FILLER_68_51 ();
 sg13g2_fill_1 FILLER_68_53 ();
 sg13g2_decap_8 FILLER_68_58 ();
 sg13g2_fill_1 FILLER_68_65 ();
 sg13g2_decap_4 FILLER_68_71 ();
 sg13g2_decap_8 FILLER_68_88 ();
 sg13g2_decap_8 FILLER_68_95 ();
 sg13g2_fill_2 FILLER_68_102 ();
 sg13g2_fill_1 FILLER_68_104 ();
 sg13g2_fill_2 FILLER_68_116 ();
 sg13g2_fill_1 FILLER_68_118 ();
 sg13g2_decap_8 FILLER_68_145 ();
 sg13g2_fill_2 FILLER_68_152 ();
 sg13g2_fill_1 FILLER_68_168 ();
 sg13g2_decap_8 FILLER_68_179 ();
 sg13g2_fill_2 FILLER_68_192 ();
 sg13g2_fill_2 FILLER_68_199 ();
 sg13g2_decap_4 FILLER_68_206 ();
 sg13g2_fill_1 FILLER_68_210 ();
 sg13g2_decap_8 FILLER_68_215 ();
 sg13g2_decap_8 FILLER_68_222 ();
 sg13g2_decap_8 FILLER_68_229 ();
 sg13g2_fill_2 FILLER_68_236 ();
 sg13g2_fill_2 FILLER_68_282 ();
 sg13g2_fill_1 FILLER_68_284 ();
 sg13g2_fill_2 FILLER_68_331 ();
 sg13g2_decap_4 FILLER_68_337 ();
 sg13g2_fill_1 FILLER_68_341 ();
 sg13g2_decap_8 FILLER_68_346 ();
 sg13g2_decap_8 FILLER_68_353 ();
 sg13g2_decap_8 FILLER_68_360 ();
 sg13g2_decap_8 FILLER_68_367 ();
 sg13g2_fill_1 FILLER_68_374 ();
 sg13g2_decap_8 FILLER_68_399 ();
 sg13g2_fill_2 FILLER_68_406 ();
 sg13g2_decap_4 FILLER_68_411 ();
 sg13g2_fill_2 FILLER_68_415 ();
 sg13g2_decap_4 FILLER_68_440 ();
 sg13g2_fill_2 FILLER_68_444 ();
 sg13g2_decap_4 FILLER_68_467 ();
 sg13g2_fill_2 FILLER_68_471 ();
 sg13g2_decap_4 FILLER_68_477 ();
 sg13g2_fill_2 FILLER_68_488 ();
 sg13g2_decap_4 FILLER_68_494 ();
 sg13g2_fill_1 FILLER_68_498 ();
 sg13g2_fill_2 FILLER_68_504 ();
 sg13g2_fill_2 FILLER_68_518 ();
 sg13g2_fill_2 FILLER_68_524 ();
 sg13g2_fill_1 FILLER_68_526 ();
 sg13g2_fill_2 FILLER_68_532 ();
 sg13g2_fill_1 FILLER_68_534 ();
 sg13g2_fill_2 FILLER_68_540 ();
 sg13g2_fill_1 FILLER_68_542 ();
 sg13g2_decap_4 FILLER_68_553 ();
 sg13g2_fill_1 FILLER_68_557 ();
 sg13g2_fill_2 FILLER_68_563 ();
 sg13g2_fill_1 FILLER_68_584 ();
 sg13g2_decap_8 FILLER_68_597 ();
 sg13g2_decap_8 FILLER_68_604 ();
 sg13g2_decap_8 FILLER_68_611 ();
 sg13g2_decap_8 FILLER_68_618 ();
 sg13g2_fill_2 FILLER_68_625 ();
 sg13g2_fill_2 FILLER_68_632 ();
 sg13g2_decap_8 FILLER_68_652 ();
 sg13g2_decap_4 FILLER_68_659 ();
 sg13g2_fill_2 FILLER_68_663 ();
 sg13g2_decap_8 FILLER_68_670 ();
 sg13g2_decap_8 FILLER_68_677 ();
 sg13g2_fill_2 FILLER_68_684 ();
 sg13g2_fill_2 FILLER_68_692 ();
 sg13g2_fill_1 FILLER_68_694 ();
 sg13g2_decap_4 FILLER_68_705 ();
 sg13g2_fill_2 FILLER_68_709 ();
 sg13g2_decap_8 FILLER_68_715 ();
 sg13g2_decap_8 FILLER_68_722 ();
 sg13g2_decap_8 FILLER_68_734 ();
 sg13g2_fill_2 FILLER_68_741 ();
 sg13g2_fill_1 FILLER_68_743 ();
 sg13g2_decap_4 FILLER_68_770 ();
 sg13g2_decap_8 FILLER_68_805 ();
 sg13g2_decap_8 FILLER_68_812 ();
 sg13g2_decap_8 FILLER_68_819 ();
 sg13g2_decap_8 FILLER_68_826 ();
 sg13g2_fill_2 FILLER_68_833 ();
 sg13g2_fill_1 FILLER_68_835 ();
 sg13g2_fill_1 FILLER_68_840 ();
 sg13g2_fill_2 FILLER_68_844 ();
 sg13g2_decap_8 FILLER_68_869 ();
 sg13g2_fill_2 FILLER_68_876 ();
 sg13g2_decap_8 FILLER_69_0 ();
 sg13g2_decap_4 FILLER_69_7 ();
 sg13g2_fill_1 FILLER_69_11 ();
 sg13g2_fill_2 FILLER_69_21 ();
 sg13g2_fill_1 FILLER_69_23 ();
 sg13g2_fill_2 FILLER_69_40 ();
 sg13g2_fill_2 FILLER_69_47 ();
 sg13g2_fill_1 FILLER_69_49 ();
 sg13g2_fill_2 FILLER_69_55 ();
 sg13g2_decap_4 FILLER_69_76 ();
 sg13g2_fill_2 FILLER_69_89 ();
 sg13g2_fill_2 FILLER_69_99 ();
 sg13g2_fill_1 FILLER_69_101 ();
 sg13g2_fill_1 FILLER_69_106 ();
 sg13g2_fill_2 FILLER_69_117 ();
 sg13g2_fill_1 FILLER_69_119 ();
 sg13g2_fill_2 FILLER_69_124 ();
 sg13g2_decap_4 FILLER_69_130 ();
 sg13g2_decap_4 FILLER_69_139 ();
 sg13g2_fill_1 FILLER_69_143 ();
 sg13g2_fill_1 FILLER_69_162 ();
 sg13g2_fill_2 FILLER_69_167 ();
 sg13g2_fill_1 FILLER_69_169 ();
 sg13g2_fill_1 FILLER_69_180 ();
 sg13g2_fill_1 FILLER_69_186 ();
 sg13g2_fill_2 FILLER_69_193 ();
 sg13g2_fill_2 FILLER_69_200 ();
 sg13g2_decap_8 FILLER_69_215 ();
 sg13g2_decap_8 FILLER_69_222 ();
 sg13g2_decap_8 FILLER_69_229 ();
 sg13g2_decap_8 FILLER_69_236 ();
 sg13g2_fill_1 FILLER_69_243 ();
 sg13g2_fill_2 FILLER_69_257 ();
 sg13g2_decap_8 FILLER_69_267 ();
 sg13g2_decap_8 FILLER_69_274 ();
 sg13g2_decap_4 FILLER_69_281 ();
 sg13g2_fill_2 FILLER_69_285 ();
 sg13g2_decap_4 FILLER_69_292 ();
 sg13g2_fill_2 FILLER_69_296 ();
 sg13g2_decap_8 FILLER_69_302 ();
 sg13g2_decap_8 FILLER_69_309 ();
 sg13g2_fill_1 FILLER_69_316 ();
 sg13g2_decap_8 FILLER_69_343 ();
 sg13g2_decap_8 FILLER_69_350 ();
 sg13g2_decap_8 FILLER_69_357 ();
 sg13g2_decap_8 FILLER_69_364 ();
 sg13g2_decap_8 FILLER_69_371 ();
 sg13g2_decap_8 FILLER_69_378 ();
 sg13g2_fill_2 FILLER_69_385 ();
 sg13g2_fill_1 FILLER_69_392 ();
 sg13g2_decap_8 FILLER_69_397 ();
 sg13g2_fill_2 FILLER_69_404 ();
 sg13g2_decap_8 FILLER_69_421 ();
 sg13g2_decap_4 FILLER_69_428 ();
 sg13g2_fill_2 FILLER_69_432 ();
 sg13g2_fill_2 FILLER_69_455 ();
 sg13g2_fill_1 FILLER_69_457 ();
 sg13g2_decap_8 FILLER_69_463 ();
 sg13g2_decap_8 FILLER_69_470 ();
 sg13g2_fill_1 FILLER_69_477 ();
 sg13g2_decap_8 FILLER_69_488 ();
 sg13g2_decap_8 FILLER_69_495 ();
 sg13g2_decap_8 FILLER_69_502 ();
 sg13g2_fill_2 FILLER_69_509 ();
 sg13g2_decap_8 FILLER_69_516 ();
 sg13g2_fill_2 FILLER_69_523 ();
 sg13g2_decap_4 FILLER_69_535 ();
 sg13g2_fill_2 FILLER_69_553 ();
 sg13g2_fill_1 FILLER_69_555 ();
 sg13g2_fill_2 FILLER_69_561 ();
 sg13g2_fill_2 FILLER_69_568 ();
 sg13g2_decap_4 FILLER_69_576 ();
 sg13g2_decap_8 FILLER_69_584 ();
 sg13g2_decap_4 FILLER_69_591 ();
 sg13g2_decap_8 FILLER_69_599 ();
 sg13g2_fill_1 FILLER_69_606 ();
 sg13g2_fill_2 FILLER_69_619 ();
 sg13g2_fill_1 FILLER_69_621 ();
 sg13g2_fill_1 FILLER_69_632 ();
 sg13g2_fill_2 FILLER_69_642 ();
 sg13g2_fill_1 FILLER_69_644 ();
 sg13g2_decap_4 FILLER_69_653 ();
 sg13g2_decap_4 FILLER_69_661 ();
 sg13g2_decap_8 FILLER_69_675 ();
 sg13g2_decap_8 FILLER_69_682 ();
 sg13g2_fill_2 FILLER_69_689 ();
 sg13g2_fill_1 FILLER_69_729 ();
 sg13g2_decap_8 FILLER_69_738 ();
 sg13g2_fill_1 FILLER_69_755 ();
 sg13g2_decap_8 FILLER_69_766 ();
 sg13g2_decap_4 FILLER_69_773 ();
 sg13g2_fill_1 FILLER_69_777 ();
 sg13g2_decap_4 FILLER_69_783 ();
 sg13g2_decap_8 FILLER_69_791 ();
 sg13g2_fill_1 FILLER_69_798 ();
 sg13g2_fill_1 FILLER_69_840 ();
 sg13g2_fill_2 FILLER_69_846 ();
 sg13g2_decap_4 FILLER_69_874 ();
 sg13g2_decap_8 FILLER_70_0 ();
 sg13g2_decap_4 FILLER_70_7 ();
 sg13g2_decap_8 FILLER_70_16 ();
 sg13g2_fill_2 FILLER_70_23 ();
 sg13g2_fill_1 FILLER_70_48 ();
 sg13g2_decap_8 FILLER_70_79 ();
 sg13g2_decap_8 FILLER_70_86 ();
 sg13g2_fill_2 FILLER_70_93 ();
 sg13g2_decap_8 FILLER_70_100 ();
 sg13g2_fill_1 FILLER_70_107 ();
 sg13g2_decap_8 FILLER_70_118 ();
 sg13g2_fill_2 FILLER_70_129 ();
 sg13g2_fill_1 FILLER_70_135 ();
 sg13g2_decap_8 FILLER_70_140 ();
 sg13g2_decap_8 FILLER_70_147 ();
 sg13g2_fill_1 FILLER_70_154 ();
 sg13g2_fill_2 FILLER_70_163 ();
 sg13g2_decap_4 FILLER_70_171 ();
 sg13g2_decap_4 FILLER_70_180 ();
 sg13g2_fill_2 FILLER_70_184 ();
 sg13g2_decap_8 FILLER_70_213 ();
 sg13g2_decap_8 FILLER_70_220 ();
 sg13g2_decap_4 FILLER_70_227 ();
 sg13g2_fill_2 FILLER_70_231 ();
 sg13g2_fill_1 FILLER_70_238 ();
 sg13g2_fill_2 FILLER_70_243 ();
 sg13g2_decap_8 FILLER_70_255 ();
 sg13g2_decap_4 FILLER_70_262 ();
 sg13g2_fill_1 FILLER_70_266 ();
 sg13g2_decap_4 FILLER_70_271 ();
 sg13g2_fill_1 FILLER_70_275 ();
 sg13g2_decap_8 FILLER_70_280 ();
 sg13g2_decap_4 FILLER_70_287 ();
 sg13g2_fill_2 FILLER_70_321 ();
 sg13g2_decap_4 FILLER_70_327 ();
 sg13g2_fill_2 FILLER_70_331 ();
 sg13g2_decap_8 FILLER_70_343 ();
 sg13g2_decap_8 FILLER_70_350 ();
 sg13g2_decap_4 FILLER_70_367 ();
 sg13g2_fill_1 FILLER_70_371 ();
 sg13g2_fill_2 FILLER_70_393 ();
 sg13g2_fill_2 FILLER_70_399 ();
 sg13g2_fill_1 FILLER_70_401 ();
 sg13g2_fill_2 FILLER_70_407 ();
 sg13g2_fill_1 FILLER_70_409 ();
 sg13g2_fill_2 FILLER_70_420 ();
 sg13g2_fill_1 FILLER_70_422 ();
 sg13g2_decap_8 FILLER_70_433 ();
 sg13g2_fill_2 FILLER_70_461 ();
 sg13g2_decap_4 FILLER_70_476 ();
 sg13g2_fill_1 FILLER_70_480 ();
 sg13g2_decap_4 FILLER_70_486 ();
 sg13g2_fill_1 FILLER_70_490 ();
 sg13g2_fill_2 FILLER_70_501 ();
 sg13g2_fill_1 FILLER_70_515 ();
 sg13g2_decap_8 FILLER_70_521 ();
 sg13g2_fill_1 FILLER_70_528 ();
 sg13g2_fill_1 FILLER_70_533 ();
 sg13g2_fill_1 FILLER_70_539 ();
 sg13g2_decap_4 FILLER_70_544 ();
 sg13g2_fill_2 FILLER_70_548 ();
 sg13g2_fill_2 FILLER_70_554 ();
 sg13g2_fill_2 FILLER_70_561 ();
 sg13g2_decap_8 FILLER_70_567 ();
 sg13g2_decap_8 FILLER_70_574 ();
 sg13g2_decap_8 FILLER_70_585 ();
 sg13g2_fill_2 FILLER_70_592 ();
 sg13g2_decap_8 FILLER_70_599 ();
 sg13g2_decap_8 FILLER_70_606 ();
 sg13g2_decap_8 FILLER_70_613 ();
 sg13g2_decap_8 FILLER_70_620 ();
 sg13g2_decap_4 FILLER_70_627 ();
 sg13g2_fill_2 FILLER_70_631 ();
 sg13g2_fill_2 FILLER_70_642 ();
 sg13g2_decap_8 FILLER_70_652 ();
 sg13g2_decap_8 FILLER_70_659 ();
 sg13g2_decap_4 FILLER_70_666 ();
 sg13g2_fill_2 FILLER_70_670 ();
 sg13g2_decap_4 FILLER_70_677 ();
 sg13g2_fill_1 FILLER_70_681 ();
 sg13g2_decap_4 FILLER_70_694 ();
 sg13g2_fill_2 FILLER_70_711 ();
 sg13g2_fill_1 FILLER_70_713 ();
 sg13g2_fill_1 FILLER_70_728 ();
 sg13g2_decap_8 FILLER_70_738 ();
 sg13g2_decap_4 FILLER_70_745 ();
 sg13g2_fill_2 FILLER_70_749 ();
 sg13g2_decap_8 FILLER_70_762 ();
 sg13g2_fill_2 FILLER_70_769 ();
 sg13g2_fill_2 FILLER_70_796 ();
 sg13g2_decap_8 FILLER_70_803 ();
 sg13g2_decap_4 FILLER_70_810 ();
 sg13g2_fill_2 FILLER_70_814 ();
 sg13g2_decap_8 FILLER_70_820 ();
 sg13g2_fill_1 FILLER_70_840 ();
 sg13g2_fill_2 FILLER_70_849 ();
 sg13g2_fill_1 FILLER_70_877 ();
 sg13g2_decap_8 FILLER_71_0 ();
 sg13g2_decap_4 FILLER_71_7 ();
 sg13g2_fill_2 FILLER_71_25 ();
 sg13g2_fill_1 FILLER_71_27 ();
 sg13g2_fill_2 FILLER_71_53 ();
 sg13g2_fill_1 FILLER_71_55 ();
 sg13g2_decap_8 FILLER_71_61 ();
 sg13g2_fill_1 FILLER_71_83 ();
 sg13g2_decap_8 FILLER_71_89 ();
 sg13g2_decap_8 FILLER_71_107 ();
 sg13g2_fill_1 FILLER_71_122 ();
 sg13g2_fill_1 FILLER_71_127 ();
 sg13g2_decap_4 FILLER_71_136 ();
 sg13g2_decap_4 FILLER_71_154 ();
 sg13g2_decap_8 FILLER_71_167 ();
 sg13g2_fill_2 FILLER_71_174 ();
 sg13g2_fill_2 FILLER_71_185 ();
 sg13g2_fill_1 FILLER_71_187 ();
 sg13g2_fill_1 FILLER_71_193 ();
 sg13g2_fill_1 FILLER_71_200 ();
 sg13g2_decap_4 FILLER_71_209 ();
 sg13g2_decap_8 FILLER_71_217 ();
 sg13g2_fill_2 FILLER_71_224 ();
 sg13g2_fill_1 FILLER_71_226 ();
 sg13g2_decap_8 FILLER_71_258 ();
 sg13g2_fill_2 FILLER_71_265 ();
 sg13g2_fill_1 FILLER_71_267 ();
 sg13g2_decap_4 FILLER_71_294 ();
 sg13g2_decap_8 FILLER_71_302 ();
 sg13g2_decap_8 FILLER_71_309 ();
 sg13g2_decap_8 FILLER_71_316 ();
 sg13g2_decap_8 FILLER_71_323 ();
 sg13g2_decap_4 FILLER_71_330 ();
 sg13g2_decap_4 FILLER_71_344 ();
 sg13g2_fill_1 FILLER_71_369 ();
 sg13g2_fill_1 FILLER_71_374 ();
 sg13g2_fill_2 FILLER_71_386 ();
 sg13g2_fill_1 FILLER_71_397 ();
 sg13g2_decap_8 FILLER_71_403 ();
 sg13g2_decap_8 FILLER_71_410 ();
 sg13g2_decap_8 FILLER_71_417 ();
 sg13g2_decap_8 FILLER_71_424 ();
 sg13g2_decap_8 FILLER_71_431 ();
 sg13g2_decap_8 FILLER_71_438 ();
 sg13g2_fill_2 FILLER_71_445 ();
 sg13g2_fill_1 FILLER_71_447 ();
 sg13g2_fill_1 FILLER_71_471 ();
 sg13g2_decap_4 FILLER_71_477 ();
 sg13g2_fill_2 FILLER_71_481 ();
 sg13g2_fill_1 FILLER_71_487 ();
 sg13g2_decap_4 FILLER_71_493 ();
 sg13g2_fill_2 FILLER_71_516 ();
 sg13g2_decap_4 FILLER_71_531 ();
 sg13g2_fill_1 FILLER_71_535 ();
 sg13g2_decap_8 FILLER_71_547 ();
 sg13g2_decap_8 FILLER_71_554 ();
 sg13g2_fill_2 FILLER_71_561 ();
 sg13g2_fill_1 FILLER_71_563 ();
 sg13g2_fill_2 FILLER_71_568 ();
 sg13g2_fill_1 FILLER_71_570 ();
 sg13g2_decap_4 FILLER_71_580 ();
 sg13g2_fill_2 FILLER_71_592 ();
 sg13g2_fill_1 FILLER_71_594 ();
 sg13g2_fill_2 FILLER_71_603 ();
 sg13g2_fill_1 FILLER_71_605 ();
 sg13g2_fill_2 FILLER_71_614 ();
 sg13g2_fill_2 FILLER_71_620 ();
 sg13g2_fill_1 FILLER_71_622 ();
 sg13g2_fill_1 FILLER_71_631 ();
 sg13g2_fill_1 FILLER_71_638 ();
 sg13g2_decap_8 FILLER_71_643 ();
 sg13g2_decap_4 FILLER_71_650 ();
 sg13g2_fill_1 FILLER_71_659 ();
 sg13g2_fill_1 FILLER_71_668 ();
 sg13g2_fill_1 FILLER_71_677 ();
 sg13g2_fill_2 FILLER_71_683 ();
 sg13g2_fill_2 FILLER_71_689 ();
 sg13g2_decap_4 FILLER_71_695 ();
 sg13g2_decap_8 FILLER_71_743 ();
 sg13g2_fill_2 FILLER_71_750 ();
 sg13g2_decap_8 FILLER_71_763 ();
 sg13g2_decap_4 FILLER_71_770 ();
 sg13g2_fill_1 FILLER_71_774 ();
 sg13g2_fill_1 FILLER_71_840 ();
 sg13g2_decap_4 FILLER_71_853 ();
 sg13g2_fill_2 FILLER_71_857 ();
 sg13g2_decap_8 FILLER_71_863 ();
 sg13g2_decap_8 FILLER_71_870 ();
 sg13g2_fill_1 FILLER_71_877 ();
 sg13g2_decap_8 FILLER_72_0 ();
 sg13g2_decap_4 FILLER_72_7 ();
 sg13g2_fill_1 FILLER_72_11 ();
 sg13g2_decap_4 FILLER_72_16 ();
 sg13g2_fill_2 FILLER_72_20 ();
 sg13g2_fill_1 FILLER_72_38 ();
 sg13g2_fill_2 FILLER_72_43 ();
 sg13g2_fill_1 FILLER_72_45 ();
 sg13g2_fill_2 FILLER_72_57 ();
 sg13g2_decap_8 FILLER_72_68 ();
 sg13g2_decap_4 FILLER_72_83 ();
 sg13g2_fill_2 FILLER_72_96 ();
 sg13g2_fill_1 FILLER_72_98 ();
 sg13g2_decap_8 FILLER_72_116 ();
 sg13g2_decap_8 FILLER_72_123 ();
 sg13g2_decap_4 FILLER_72_136 ();
 sg13g2_fill_2 FILLER_72_140 ();
 sg13g2_fill_2 FILLER_72_147 ();
 sg13g2_fill_1 FILLER_72_149 ();
 sg13g2_fill_1 FILLER_72_160 ();
 sg13g2_fill_2 FILLER_72_165 ();
 sg13g2_fill_2 FILLER_72_188 ();
 sg13g2_decap_4 FILLER_72_194 ();
 sg13g2_decap_8 FILLER_72_203 ();
 sg13g2_decap_8 FILLER_72_210 ();
 sg13g2_decap_8 FILLER_72_217 ();
 sg13g2_decap_8 FILLER_72_224 ();
 sg13g2_decap_4 FILLER_72_231 ();
 sg13g2_fill_1 FILLER_72_235 ();
 sg13g2_decap_8 FILLER_72_250 ();
 sg13g2_decap_8 FILLER_72_257 ();
 sg13g2_decap_8 FILLER_72_264 ();
 sg13g2_decap_8 FILLER_72_271 ();
 sg13g2_decap_8 FILLER_72_278 ();
 sg13g2_fill_1 FILLER_72_289 ();
 sg13g2_fill_2 FILLER_72_294 ();
 sg13g2_fill_1 FILLER_72_296 ();
 sg13g2_decap_8 FILLER_72_301 ();
 sg13g2_decap_8 FILLER_72_308 ();
 sg13g2_decap_8 FILLER_72_315 ();
 sg13g2_decap_8 FILLER_72_322 ();
 sg13g2_decap_4 FILLER_72_329 ();
 sg13g2_decap_8 FILLER_72_342 ();
 sg13g2_fill_1 FILLER_72_349 ();
 sg13g2_decap_8 FILLER_72_370 ();
 sg13g2_decap_8 FILLER_72_377 ();
 sg13g2_decap_8 FILLER_72_393 ();
 sg13g2_fill_2 FILLER_72_400 ();
 sg13g2_decap_8 FILLER_72_407 ();
 sg13g2_decap_8 FILLER_72_414 ();
 sg13g2_fill_2 FILLER_72_421 ();
 sg13g2_fill_1 FILLER_72_423 ();
 sg13g2_fill_1 FILLER_72_433 ();
 sg13g2_decap_4 FILLER_72_438 ();
 sg13g2_fill_1 FILLER_72_442 ();
 sg13g2_decap_8 FILLER_72_467 ();
 sg13g2_decap_8 FILLER_72_474 ();
 sg13g2_decap_8 FILLER_72_481 ();
 sg13g2_decap_8 FILLER_72_488 ();
 sg13g2_decap_4 FILLER_72_495 ();
 sg13g2_fill_2 FILLER_72_499 ();
 sg13g2_fill_2 FILLER_72_515 ();
 sg13g2_fill_1 FILLER_72_521 ();
 sg13g2_decap_8 FILLER_72_551 ();
 sg13g2_decap_4 FILLER_72_558 ();
 sg13g2_decap_8 FILLER_72_572 ();
 sg13g2_decap_4 FILLER_72_579 ();
 sg13g2_fill_1 FILLER_72_583 ();
 sg13g2_decap_8 FILLER_72_592 ();
 sg13g2_decap_8 FILLER_72_599 ();
 sg13g2_fill_1 FILLER_72_606 ();
 sg13g2_fill_2 FILLER_72_612 ();
 sg13g2_fill_1 FILLER_72_614 ();
 sg13g2_decap_4 FILLER_72_628 ();
 sg13g2_fill_1 FILLER_72_632 ();
 sg13g2_fill_2 FILLER_72_672 ();
 sg13g2_fill_2 FILLER_72_682 ();
 sg13g2_fill_1 FILLER_72_684 ();
 sg13g2_decap_8 FILLER_72_689 ();
 sg13g2_fill_2 FILLER_72_696 ();
 sg13g2_fill_2 FILLER_72_708 ();
 sg13g2_fill_1 FILLER_72_710 ();
 sg13g2_fill_2 FILLER_72_720 ();
 sg13g2_fill_1 FILLER_72_722 ();
 sg13g2_fill_2 FILLER_72_731 ();
 sg13g2_decap_8 FILLER_72_737 ();
 sg13g2_fill_1 FILLER_72_744 ();
 sg13g2_decap_8 FILLER_72_750 ();
 sg13g2_fill_2 FILLER_72_757 ();
 sg13g2_decap_4 FILLER_72_763 ();
 sg13g2_decap_8 FILLER_72_770 ();
 sg13g2_decap_4 FILLER_72_777 ();
 sg13g2_decap_8 FILLER_72_785 ();
 sg13g2_decap_8 FILLER_72_792 ();
 sg13g2_decap_8 FILLER_72_799 ();
 sg13g2_fill_1 FILLER_72_806 ();
 sg13g2_decap_4 FILLER_72_838 ();
 sg13g2_fill_1 FILLER_72_842 ();
 sg13g2_fill_2 FILLER_72_848 ();
 sg13g2_fill_1 FILLER_72_850 ();
 sg13g2_fill_1 FILLER_72_877 ();
 sg13g2_decap_8 FILLER_73_0 ();
 sg13g2_decap_8 FILLER_73_7 ();
 sg13g2_fill_2 FILLER_73_14 ();
 sg13g2_fill_2 FILLER_73_20 ();
 sg13g2_fill_1 FILLER_73_30 ();
 sg13g2_fill_1 FILLER_73_35 ();
 sg13g2_fill_2 FILLER_73_42 ();
 sg13g2_fill_1 FILLER_73_54 ();
 sg13g2_fill_2 FILLER_73_68 ();
 sg13g2_fill_1 FILLER_73_70 ();
 sg13g2_decap_8 FILLER_73_76 ();
 sg13g2_decap_4 FILLER_73_83 ();
 sg13g2_decap_4 FILLER_73_102 ();
 sg13g2_fill_2 FILLER_73_110 ();
 sg13g2_fill_1 FILLER_73_117 ();
 sg13g2_decap_8 FILLER_73_122 ();
 sg13g2_decap_8 FILLER_73_129 ();
 sg13g2_decap_8 FILLER_73_136 ();
 sg13g2_fill_1 FILLER_73_143 ();
 sg13g2_fill_1 FILLER_73_153 ();
 sg13g2_fill_1 FILLER_73_159 ();
 sg13g2_decap_8 FILLER_73_171 ();
 sg13g2_decap_8 FILLER_73_178 ();
 sg13g2_decap_4 FILLER_73_185 ();
 sg13g2_fill_2 FILLER_73_189 ();
 sg13g2_fill_2 FILLER_73_195 ();
 sg13g2_decap_8 FILLER_73_201 ();
 sg13g2_fill_2 FILLER_73_208 ();
 sg13g2_fill_1 FILLER_73_210 ();
 sg13g2_fill_1 FILLER_73_234 ();
 sg13g2_fill_1 FILLER_73_244 ();
 sg13g2_fill_2 FILLER_73_256 ();
 sg13g2_fill_1 FILLER_73_258 ();
 sg13g2_fill_1 FILLER_73_268 ();
 sg13g2_decap_4 FILLER_73_305 ();
 sg13g2_fill_1 FILLER_73_309 ();
 sg13g2_fill_2 FILLER_73_341 ();
 sg13g2_decap_8 FILLER_73_352 ();
 sg13g2_decap_8 FILLER_73_359 ();
 sg13g2_decap_8 FILLER_73_371 ();
 sg13g2_fill_1 FILLER_73_413 ();
 sg13g2_decap_8 FILLER_73_444 ();
 sg13g2_fill_2 FILLER_73_451 ();
 sg13g2_decap_8 FILLER_73_479 ();
 sg13g2_decap_8 FILLER_73_486 ();
 sg13g2_fill_1 FILLER_73_493 ();
 sg13g2_decap_4 FILLER_73_502 ();
 sg13g2_fill_1 FILLER_73_506 ();
 sg13g2_decap_8 FILLER_73_524 ();
 sg13g2_fill_2 FILLER_73_531 ();
 sg13g2_fill_2 FILLER_73_565 ();
 sg13g2_decap_8 FILLER_73_571 ();
 sg13g2_decap_8 FILLER_73_578 ();
 sg13g2_decap_8 FILLER_73_585 ();
 sg13g2_decap_8 FILLER_73_592 ();
 sg13g2_fill_2 FILLER_73_609 ();
 sg13g2_fill_1 FILLER_73_611 ();
 sg13g2_fill_1 FILLER_73_616 ();
 sg13g2_fill_2 FILLER_73_632 ();
 sg13g2_decap_8 FILLER_73_654 ();
 sg13g2_decap_4 FILLER_73_661 ();
 sg13g2_fill_2 FILLER_73_665 ();
 sg13g2_decap_8 FILLER_73_679 ();
 sg13g2_decap_8 FILLER_73_686 ();
 sg13g2_decap_4 FILLER_73_693 ();
 sg13g2_fill_2 FILLER_73_697 ();
 sg13g2_fill_2 FILLER_73_746 ();
 sg13g2_fill_2 FILLER_73_762 ();
 sg13g2_fill_2 FILLER_73_800 ();
 sg13g2_decap_8 FILLER_73_812 ();
 sg13g2_fill_1 FILLER_73_827 ();
 sg13g2_decap_8 FILLER_73_832 ();
 sg13g2_decap_8 FILLER_73_839 ();
 sg13g2_decap_8 FILLER_73_846 ();
 sg13g2_decap_4 FILLER_73_853 ();
 sg13g2_fill_1 FILLER_73_857 ();
 sg13g2_decap_8 FILLER_73_862 ();
 sg13g2_decap_8 FILLER_73_869 ();
 sg13g2_fill_2 FILLER_73_876 ();
 sg13g2_decap_8 FILLER_74_0 ();
 sg13g2_decap_8 FILLER_74_7 ();
 sg13g2_fill_1 FILLER_74_14 ();
 sg13g2_decap_4 FILLER_74_29 ();
 sg13g2_fill_2 FILLER_74_41 ();
 sg13g2_decap_4 FILLER_74_48 ();
 sg13g2_fill_1 FILLER_74_66 ();
 sg13g2_decap_8 FILLER_74_83 ();
 sg13g2_decap_4 FILLER_74_90 ();
 sg13g2_fill_1 FILLER_74_94 ();
 sg13g2_fill_1 FILLER_74_103 ();
 sg13g2_fill_1 FILLER_74_124 ();
 sg13g2_fill_2 FILLER_74_146 ();
 sg13g2_decap_8 FILLER_74_169 ();
 sg13g2_decap_8 FILLER_74_176 ();
 sg13g2_decap_8 FILLER_74_183 ();
 sg13g2_decap_4 FILLER_74_190 ();
 sg13g2_fill_2 FILLER_74_194 ();
 sg13g2_decap_4 FILLER_74_201 ();
 sg13g2_fill_1 FILLER_74_205 ();
 sg13g2_decap_8 FILLER_74_226 ();
 sg13g2_decap_8 FILLER_74_233 ();
 sg13g2_fill_1 FILLER_74_240 ();
 sg13g2_decap_8 FILLER_74_251 ();
 sg13g2_decap_8 FILLER_74_258 ();
 sg13g2_decap_8 FILLER_74_265 ();
 sg13g2_fill_2 FILLER_74_272 ();
 sg13g2_fill_1 FILLER_74_274 ();
 sg13g2_decap_4 FILLER_74_285 ();
 sg13g2_decap_8 FILLER_74_293 ();
 sg13g2_decap_8 FILLER_74_300 ();
 sg13g2_decap_8 FILLER_74_307 ();
 sg13g2_decap_8 FILLER_74_374 ();
 sg13g2_decap_8 FILLER_74_381 ();
 sg13g2_fill_1 FILLER_74_388 ();
 sg13g2_decap_8 FILLER_74_393 ();
 sg13g2_decap_8 FILLER_74_400 ();
 sg13g2_fill_1 FILLER_74_407 ();
 sg13g2_fill_2 FILLER_74_412 ();
 sg13g2_fill_1 FILLER_74_414 ();
 sg13g2_decap_8 FILLER_74_432 ();
 sg13g2_decap_8 FILLER_74_439 ();
 sg13g2_decap_8 FILLER_74_446 ();
 sg13g2_decap_4 FILLER_74_453 ();
 sg13g2_decap_8 FILLER_74_461 ();
 sg13g2_decap_8 FILLER_74_468 ();
 sg13g2_decap_8 FILLER_74_475 ();
 sg13g2_decap_8 FILLER_74_487 ();
 sg13g2_fill_1 FILLER_74_494 ();
 sg13g2_decap_4 FILLER_74_500 ();
 sg13g2_fill_2 FILLER_74_504 ();
 sg13g2_fill_2 FILLER_74_514 ();
 sg13g2_fill_1 FILLER_74_542 ();
 sg13g2_decap_8 FILLER_74_551 ();
 sg13g2_fill_1 FILLER_74_558 ();
 sg13g2_fill_1 FILLER_74_567 ();
 sg13g2_decap_8 FILLER_74_580 ();
 sg13g2_decap_4 FILLER_74_587 ();
 sg13g2_fill_1 FILLER_74_591 ();
 sg13g2_fill_2 FILLER_74_613 ();
 sg13g2_fill_1 FILLER_74_615 ();
 sg13g2_decap_8 FILLER_74_624 ();
 sg13g2_decap_4 FILLER_74_631 ();
 sg13g2_fill_2 FILLER_74_635 ();
 sg13g2_fill_1 FILLER_74_646 ();
 sg13g2_decap_4 FILLER_74_655 ();
 sg13g2_decap_8 FILLER_74_662 ();
 sg13g2_decap_8 FILLER_74_677 ();
 sg13g2_fill_2 FILLER_74_684 ();
 sg13g2_decap_8 FILLER_74_691 ();
 sg13g2_decap_4 FILLER_74_698 ();
 sg13g2_decap_4 FILLER_74_747 ();
 sg13g2_decap_4 FILLER_74_755 ();
 sg13g2_fill_2 FILLER_74_767 ();
 sg13g2_fill_2 FILLER_74_779 ();
 sg13g2_decap_8 FILLER_74_785 ();
 sg13g2_decap_4 FILLER_74_792 ();
 sg13g2_fill_1 FILLER_74_796 ();
 sg13g2_fill_1 FILLER_74_807 ();
 sg13g2_decap_4 FILLER_74_834 ();
 sg13g2_fill_2 FILLER_74_838 ();
 sg13g2_fill_2 FILLER_74_850 ();
 sg13g2_decap_8 FILLER_75_0 ();
 sg13g2_decap_4 FILLER_75_7 ();
 sg13g2_fill_1 FILLER_75_21 ();
 sg13g2_fill_1 FILLER_75_26 ();
 sg13g2_fill_2 FILLER_75_37 ();
 sg13g2_fill_1 FILLER_75_39 ();
 sg13g2_fill_1 FILLER_75_53 ();
 sg13g2_decap_8 FILLER_75_60 ();
 sg13g2_fill_1 FILLER_75_67 ();
 sg13g2_decap_4 FILLER_75_72 ();
 sg13g2_fill_2 FILLER_75_76 ();
 sg13g2_decap_8 FILLER_75_94 ();
 sg13g2_fill_1 FILLER_75_101 ();
 sg13g2_decap_4 FILLER_75_108 ();
 sg13g2_fill_2 FILLER_75_129 ();
 sg13g2_fill_1 FILLER_75_139 ();
 sg13g2_decap_4 FILLER_75_157 ();
 sg13g2_decap_8 FILLER_75_170 ();
 sg13g2_decap_8 FILLER_75_177 ();
 sg13g2_fill_2 FILLER_75_193 ();
 sg13g2_fill_1 FILLER_75_195 ();
 sg13g2_decap_8 FILLER_75_201 ();
 sg13g2_decap_8 FILLER_75_208 ();
 sg13g2_fill_2 FILLER_75_215 ();
 sg13g2_fill_2 FILLER_75_226 ();
 sg13g2_fill_2 FILLER_75_232 ();
 sg13g2_decap_8 FILLER_75_270 ();
 sg13g2_decap_4 FILLER_75_277 ();
 sg13g2_fill_1 FILLER_75_281 ();
 sg13g2_decap_8 FILLER_75_308 ();
 sg13g2_decap_8 FILLER_75_315 ();
 sg13g2_decap_4 FILLER_75_322 ();
 sg13g2_fill_1 FILLER_75_326 ();
 sg13g2_decap_4 FILLER_75_331 ();
 sg13g2_fill_1 FILLER_75_335 ();
 sg13g2_fill_2 FILLER_75_356 ();
 sg13g2_fill_1 FILLER_75_362 ();
 sg13g2_fill_2 FILLER_75_368 ();
 sg13g2_fill_2 FILLER_75_374 ();
 sg13g2_fill_1 FILLER_75_376 ();
 sg13g2_fill_2 FILLER_75_403 ();
 sg13g2_fill_1 FILLER_75_405 ();
 sg13g2_decap_4 FILLER_75_440 ();
 sg13g2_decap_4 FILLER_75_470 ();
 sg13g2_fill_1 FILLER_75_492 ();
 sg13g2_fill_1 FILLER_75_497 ();
 sg13g2_decap_8 FILLER_75_503 ();
 sg13g2_decap_8 FILLER_75_510 ();
 sg13g2_fill_1 FILLER_75_517 ();
 sg13g2_decap_4 FILLER_75_523 ();
 sg13g2_fill_2 FILLER_75_527 ();
 sg13g2_fill_1 FILLER_75_545 ();
 sg13g2_decap_8 FILLER_75_554 ();
 sg13g2_fill_2 FILLER_75_561 ();
 sg13g2_fill_1 FILLER_75_563 ();
 sg13g2_decap_8 FILLER_75_574 ();
 sg13g2_decap_8 FILLER_75_581 ();
 sg13g2_fill_2 FILLER_75_596 ();
 sg13g2_fill_1 FILLER_75_598 ();
 sg13g2_fill_1 FILLER_75_604 ();
 sg13g2_decap_8 FILLER_75_622 ();
 sg13g2_decap_4 FILLER_75_629 ();
 sg13g2_fill_1 FILLER_75_633 ();
 sg13g2_fill_2 FILLER_75_638 ();
 sg13g2_fill_1 FILLER_75_640 ();
 sg13g2_fill_1 FILLER_75_646 ();
 sg13g2_fill_2 FILLER_75_653 ();
 sg13g2_fill_1 FILLER_75_655 ();
 sg13g2_decap_4 FILLER_75_674 ();
 sg13g2_decap_8 FILLER_75_704 ();
 sg13g2_decap_8 FILLER_75_711 ();
 sg13g2_decap_8 FILLER_75_722 ();
 sg13g2_decap_8 FILLER_75_729 ();
 sg13g2_decap_8 FILLER_75_736 ();
 sg13g2_decap_4 FILLER_75_743 ();
 sg13g2_fill_2 FILLER_75_758 ();
 sg13g2_decap_8 FILLER_75_768 ();
 sg13g2_fill_1 FILLER_75_775 ();
 sg13g2_decap_8 FILLER_75_806 ();
 sg13g2_fill_1 FILLER_75_813 ();
 sg13g2_decap_8 FILLER_75_821 ();
 sg13g2_decap_8 FILLER_75_828 ();
 sg13g2_decap_8 FILLER_75_835 ();
 sg13g2_fill_1 FILLER_75_842 ();
 sg13g2_decap_8 FILLER_75_847 ();
 sg13g2_decap_4 FILLER_75_854 ();
 sg13g2_decap_8 FILLER_75_862 ();
 sg13g2_decap_8 FILLER_75_869 ();
 sg13g2_fill_2 FILLER_75_876 ();
 sg13g2_decap_8 FILLER_76_0 ();
 sg13g2_decap_8 FILLER_76_7 ();
 sg13g2_decap_4 FILLER_76_14 ();
 sg13g2_fill_1 FILLER_76_18 ();
 sg13g2_fill_2 FILLER_76_33 ();
 sg13g2_fill_2 FILLER_76_60 ();
 sg13g2_fill_1 FILLER_76_62 ();
 sg13g2_fill_2 FILLER_76_68 ();
 sg13g2_fill_2 FILLER_76_78 ();
 sg13g2_fill_1 FILLER_76_80 ();
 sg13g2_decap_4 FILLER_76_86 ();
 sg13g2_decap_4 FILLER_76_101 ();
 sg13g2_fill_1 FILLER_76_111 ();
 sg13g2_decap_8 FILLER_76_128 ();
 sg13g2_decap_8 FILLER_76_135 ();
 sg13g2_decap_8 FILLER_76_142 ();
 sg13g2_decap_8 FILLER_76_149 ();
 sg13g2_decap_8 FILLER_76_156 ();
 sg13g2_decap_8 FILLER_76_163 ();
 sg13g2_decap_8 FILLER_76_170 ();
 sg13g2_fill_2 FILLER_76_177 ();
 sg13g2_decap_8 FILLER_76_210 ();
 sg13g2_fill_2 FILLER_76_243 ();
 sg13g2_fill_1 FILLER_76_249 ();
 sg13g2_fill_2 FILLER_76_262 ();
 sg13g2_fill_1 FILLER_76_264 ();
 sg13g2_fill_2 FILLER_76_270 ();
 sg13g2_decap_8 FILLER_76_298 ();
 sg13g2_decap_8 FILLER_76_305 ();
 sg13g2_fill_2 FILLER_76_312 ();
 sg13g2_decap_4 FILLER_76_322 ();
 sg13g2_fill_1 FILLER_76_326 ();
 sg13g2_decap_8 FILLER_76_331 ();
 sg13g2_decap_8 FILLER_76_338 ();
 sg13g2_fill_1 FILLER_76_355 ();
 sg13g2_fill_1 FILLER_76_366 ();
 sg13g2_decap_4 FILLER_76_377 ();
 sg13g2_fill_2 FILLER_76_386 ();
 sg13g2_fill_2 FILLER_76_392 ();
 sg13g2_fill_1 FILLER_76_394 ();
 sg13g2_decap_8 FILLER_76_405 ();
 sg13g2_fill_2 FILLER_76_412 ();
 sg13g2_fill_1 FILLER_76_414 ();
 sg13g2_fill_2 FILLER_76_430 ();
 sg13g2_fill_2 FILLER_76_442 ();
 sg13g2_fill_2 FILLER_76_449 ();
 sg13g2_fill_1 FILLER_76_451 ();
 sg13g2_fill_2 FILLER_76_456 ();
 sg13g2_fill_1 FILLER_76_458 ();
 sg13g2_fill_2 FILLER_76_485 ();
 sg13g2_decap_8 FILLER_76_492 ();
 sg13g2_fill_1 FILLER_76_499 ();
 sg13g2_fill_2 FILLER_76_504 ();
 sg13g2_fill_1 FILLER_76_506 ();
 sg13g2_decap_8 FILLER_76_516 ();
 sg13g2_decap_4 FILLER_76_523 ();
 sg13g2_fill_1 FILLER_76_527 ();
 sg13g2_decap_8 FILLER_76_536 ();
 sg13g2_decap_8 FILLER_76_543 ();
 sg13g2_decap_4 FILLER_76_550 ();
 sg13g2_fill_2 FILLER_76_570 ();
 sg13g2_decap_8 FILLER_76_576 ();
 sg13g2_decap_8 FILLER_76_583 ();
 sg13g2_fill_1 FILLER_76_590 ();
 sg13g2_fill_1 FILLER_76_599 ();
 sg13g2_fill_2 FILLER_76_604 ();
 sg13g2_fill_1 FILLER_76_610 ();
 sg13g2_fill_2 FILLER_76_619 ();
 sg13g2_decap_8 FILLER_76_634 ();
 sg13g2_decap_8 FILLER_76_664 ();
 sg13g2_decap_8 FILLER_76_671 ();
 sg13g2_fill_2 FILLER_76_678 ();
 sg13g2_decap_8 FILLER_76_687 ();
 sg13g2_decap_8 FILLER_76_694 ();
 sg13g2_fill_2 FILLER_76_701 ();
 sg13g2_fill_1 FILLER_76_703 ();
 sg13g2_fill_2 FILLER_76_740 ();
 sg13g2_fill_1 FILLER_76_742 ();
 sg13g2_fill_1 FILLER_76_757 ();
 sg13g2_decap_4 FILLER_76_768 ();
 sg13g2_fill_2 FILLER_76_772 ();
 sg13g2_fill_1 FILLER_76_779 ();
 sg13g2_decap_8 FILLER_76_787 ();
 sg13g2_decap_8 FILLER_76_794 ();
 sg13g2_decap_8 FILLER_76_801 ();
 sg13g2_fill_1 FILLER_76_808 ();
 sg13g2_fill_1 FILLER_76_819 ();
 sg13g2_decap_8 FILLER_76_824 ();
 sg13g2_decap_4 FILLER_76_831 ();
 sg13g2_decap_8 FILLER_76_850 ();
 sg13g2_fill_2 FILLER_76_857 ();
 sg13g2_decap_8 FILLER_76_863 ();
 sg13g2_decap_8 FILLER_76_870 ();
 sg13g2_fill_1 FILLER_76_877 ();
 sg13g2_decap_8 FILLER_77_0 ();
 sg13g2_decap_8 FILLER_77_7 ();
 sg13g2_decap_8 FILLER_77_14 ();
 sg13g2_decap_8 FILLER_77_21 ();
 sg13g2_decap_8 FILLER_77_36 ();
 sg13g2_fill_1 FILLER_77_43 ();
 sg13g2_decap_8 FILLER_77_48 ();
 sg13g2_decap_8 FILLER_77_59 ();
 sg13g2_decap_8 FILLER_77_66 ();
 sg13g2_fill_1 FILLER_77_73 ();
 sg13g2_decap_8 FILLER_77_86 ();
 sg13g2_decap_4 FILLER_77_103 ();
 sg13g2_decap_8 FILLER_77_118 ();
 sg13g2_decap_8 FILLER_77_125 ();
 sg13g2_decap_8 FILLER_77_132 ();
 sg13g2_fill_2 FILLER_77_139 ();
 sg13g2_fill_1 FILLER_77_141 ();
 sg13g2_decap_4 FILLER_77_146 ();
 sg13g2_decap_4 FILLER_77_185 ();
 sg13g2_decap_8 FILLER_77_193 ();
 sg13g2_decap_8 FILLER_77_200 ();
 sg13g2_decap_8 FILLER_77_228 ();
 sg13g2_decap_8 FILLER_77_235 ();
 sg13g2_decap_8 FILLER_77_242 ();
 sg13g2_decap_8 FILLER_77_249 ();
 sg13g2_fill_2 FILLER_77_256 ();
 sg13g2_fill_1 FILLER_77_258 ();
 sg13g2_decap_8 FILLER_77_267 ();
 sg13g2_decap_4 FILLER_77_274 ();
 sg13g2_fill_2 FILLER_77_278 ();
 sg13g2_fill_2 FILLER_77_289 ();
 sg13g2_fill_1 FILLER_77_291 ();
 sg13g2_decap_4 FILLER_77_295 ();
 sg13g2_fill_1 FILLER_77_299 ();
 sg13g2_decap_8 FILLER_77_304 ();
 sg13g2_decap_4 FILLER_77_311 ();
 sg13g2_fill_1 FILLER_77_315 ();
 sg13g2_decap_8 FILLER_77_347 ();
 sg13g2_fill_1 FILLER_77_354 ();
 sg13g2_decap_8 FILLER_77_381 ();
 sg13g2_decap_8 FILLER_77_388 ();
 sg13g2_decap_8 FILLER_77_395 ();
 sg13g2_decap_8 FILLER_77_402 ();
 sg13g2_decap_8 FILLER_77_440 ();
 sg13g2_decap_4 FILLER_77_447 ();
 sg13g2_fill_2 FILLER_77_451 ();
 sg13g2_decap_8 FILLER_77_457 ();
 sg13g2_fill_2 FILLER_77_464 ();
 sg13g2_decap_4 FILLER_77_470 ();
 sg13g2_fill_1 FILLER_77_487 ();
 sg13g2_decap_4 FILLER_77_493 ();
 sg13g2_fill_2 FILLER_77_505 ();
 sg13g2_fill_1 FILLER_77_507 ();
 sg13g2_fill_1 FILLER_77_512 ();
 sg13g2_fill_2 FILLER_77_521 ();
 sg13g2_fill_1 FILLER_77_523 ();
 sg13g2_decap_8 FILLER_77_549 ();
 sg13g2_decap_8 FILLER_77_585 ();
 sg13g2_decap_8 FILLER_77_592 ();
 sg13g2_fill_1 FILLER_77_599 ();
 sg13g2_fill_2 FILLER_77_613 ();
 sg13g2_decap_8 FILLER_77_632 ();
 sg13g2_decap_4 FILLER_77_639 ();
 sg13g2_fill_1 FILLER_77_643 ();
 sg13g2_decap_4 FILLER_77_669 ();
 sg13g2_fill_2 FILLER_77_673 ();
 sg13g2_decap_8 FILLER_77_687 ();
 sg13g2_fill_2 FILLER_77_694 ();
 sg13g2_fill_1 FILLER_77_696 ();
 sg13g2_decap_8 FILLER_77_702 ();
 sg13g2_decap_8 FILLER_77_709 ();
 sg13g2_fill_1 FILLER_77_716 ();
 sg13g2_fill_1 FILLER_77_725 ();
 sg13g2_decap_8 FILLER_77_734 ();
 sg13g2_decap_4 FILLER_77_741 ();
 sg13g2_fill_2 FILLER_77_745 ();
 sg13g2_fill_2 FILLER_77_773 ();
 sg13g2_fill_2 FILLER_77_806 ();
 sg13g2_fill_1 FILLER_77_808 ();
 sg13g2_fill_2 FILLER_77_812 ();
 sg13g2_fill_2 FILLER_77_850 ();
 sg13g2_decap_8 FILLER_78_0 ();
 sg13g2_decap_8 FILLER_78_7 ();
 sg13g2_decap_8 FILLER_78_14 ();
 sg13g2_decap_8 FILLER_78_21 ();
 sg13g2_decap_8 FILLER_78_28 ();
 sg13g2_decap_4 FILLER_78_35 ();
 sg13g2_decap_8 FILLER_78_42 ();
 sg13g2_decap_8 FILLER_78_49 ();
 sg13g2_decap_8 FILLER_78_56 ();
 sg13g2_decap_8 FILLER_78_63 ();
 sg13g2_decap_8 FILLER_78_70 ();
 sg13g2_decap_4 FILLER_78_77 ();
 sg13g2_decap_8 FILLER_78_89 ();
 sg13g2_decap_8 FILLER_78_96 ();
 sg13g2_decap_8 FILLER_78_103 ();
 sg13g2_decap_8 FILLER_78_110 ();
 sg13g2_decap_8 FILLER_78_117 ();
 sg13g2_decap_8 FILLER_78_124 ();
 sg13g2_decap_4 FILLER_78_131 ();
 sg13g2_decap_4 FILLER_78_202 ();
 sg13g2_decap_4 FILLER_78_237 ();
 sg13g2_fill_2 FILLER_78_241 ();
 sg13g2_decap_8 FILLER_78_278 ();
 sg13g2_decap_4 FILLER_78_285 ();
 sg13g2_decap_4 FILLER_78_319 ();
 sg13g2_decap_8 FILLER_78_349 ();
 sg13g2_decap_8 FILLER_78_356 ();
 sg13g2_decap_8 FILLER_78_367 ();
 sg13g2_decap_4 FILLER_78_374 ();
 sg13g2_fill_2 FILLER_78_382 ();
 sg13g2_fill_1 FILLER_78_384 ();
 sg13g2_decap_4 FILLER_78_411 ();
 sg13g2_fill_1 FILLER_78_415 ();
 sg13g2_decap_8 FILLER_78_420 ();
 sg13g2_decap_8 FILLER_78_427 ();
 sg13g2_decap_4 FILLER_78_434 ();
 sg13g2_fill_2 FILLER_78_438 ();
 sg13g2_fill_2 FILLER_78_444 ();
 sg13g2_fill_1 FILLER_78_446 ();
 sg13g2_fill_2 FILLER_78_473 ();
 sg13g2_fill_1 FILLER_78_475 ();
 sg13g2_fill_1 FILLER_78_484 ();
 sg13g2_decap_8 FILLER_78_490 ();
 sg13g2_decap_8 FILLER_78_497 ();
 sg13g2_decap_4 FILLER_78_504 ();
 sg13g2_decap_8 FILLER_78_516 ();
 sg13g2_decap_8 FILLER_78_523 ();
 sg13g2_fill_2 FILLER_78_530 ();
 sg13g2_fill_1 FILLER_78_532 ();
 sg13g2_decap_8 FILLER_78_546 ();
 sg13g2_fill_2 FILLER_78_553 ();
 sg13g2_decap_8 FILLER_78_563 ();
 sg13g2_decap_8 FILLER_78_570 ();
 sg13g2_fill_1 FILLER_78_577 ();
 sg13g2_decap_8 FILLER_78_591 ();
 sg13g2_fill_1 FILLER_78_598 ();
 sg13g2_decap_8 FILLER_78_614 ();
 sg13g2_decap_8 FILLER_78_621 ();
 sg13g2_decap_8 FILLER_78_628 ();
 sg13g2_decap_8 FILLER_78_635 ();
 sg13g2_decap_8 FILLER_78_642 ();
 sg13g2_decap_4 FILLER_78_649 ();
 sg13g2_fill_2 FILLER_78_657 ();
 sg13g2_fill_1 FILLER_78_667 ();
 sg13g2_fill_2 FILLER_78_673 ();
 sg13g2_decap_4 FILLER_78_736 ();
 sg13g2_fill_1 FILLER_78_740 ();
 sg13g2_fill_1 FILLER_78_746 ();
 sg13g2_fill_1 FILLER_78_756 ();
 sg13g2_decap_4 FILLER_78_762 ();
 sg13g2_fill_2 FILLER_78_771 ();
 sg13g2_decap_8 FILLER_78_778 ();
 sg13g2_fill_2 FILLER_78_789 ();
 sg13g2_fill_2 FILLER_78_796 ();
 sg13g2_fill_1 FILLER_78_798 ();
 sg13g2_fill_2 FILLER_78_804 ();
 sg13g2_fill_1 FILLER_78_806 ();
 sg13g2_fill_2 FILLER_78_812 ();
 sg13g2_decap_8 FILLER_78_827 ();
 sg13g2_decap_8 FILLER_78_834 ();
 sg13g2_fill_1 FILLER_78_841 ();
 sg13g2_decap_4 FILLER_78_872 ();
 sg13g2_fill_2 FILLER_78_876 ();
 sg13g2_decap_8 FILLER_79_0 ();
 sg13g2_decap_4 FILLER_79_7 ();
 sg13g2_fill_1 FILLER_79_11 ();
 sg13g2_fill_1 FILLER_79_16 ();
 sg13g2_fill_2 FILLER_79_72 ();
 sg13g2_fill_1 FILLER_79_74 ();
 sg13g2_fill_2 FILLER_79_84 ();
 sg13g2_fill_1 FILLER_79_91 ();
 sg13g2_decap_8 FILLER_79_126 ();
 sg13g2_decap_8 FILLER_79_133 ();
 sg13g2_fill_1 FILLER_79_140 ();
 sg13g2_decap_4 FILLER_79_145 ();
 sg13g2_decap_8 FILLER_79_153 ();
 sg13g2_decap_4 FILLER_79_160 ();
 sg13g2_fill_2 FILLER_79_168 ();
 sg13g2_decap_8 FILLER_79_196 ();
 sg13g2_fill_2 FILLER_79_203 ();
 sg13g2_fill_2 FILLER_79_209 ();
 sg13g2_fill_1 FILLER_79_214 ();
 sg13g2_fill_1 FILLER_79_219 ();
 sg13g2_decap_8 FILLER_79_224 ();
 sg13g2_fill_2 FILLER_79_240 ();
 sg13g2_fill_1 FILLER_79_242 ();
 sg13g2_fill_1 FILLER_79_247 ();
 sg13g2_fill_2 FILLER_79_252 ();
 sg13g2_decap_4 FILLER_79_262 ();
 sg13g2_decap_4 FILLER_79_271 ();
 sg13g2_fill_2 FILLER_79_275 ();
 sg13g2_decap_8 FILLER_79_281 ();
 sg13g2_decap_8 FILLER_79_288 ();
 sg13g2_decap_8 FILLER_79_295 ();
 sg13g2_decap_4 FILLER_79_302 ();
 sg13g2_decap_8 FILLER_79_310 ();
 sg13g2_decap_8 FILLER_79_317 ();
 sg13g2_decap_8 FILLER_79_324 ();
 sg13g2_decap_8 FILLER_79_335 ();
 sg13g2_decap_4 FILLER_79_342 ();
 sg13g2_decap_4 FILLER_79_396 ();
 sg13g2_fill_2 FILLER_79_400 ();
 sg13g2_decap_8 FILLER_79_406 ();
 sg13g2_decap_8 FILLER_79_413 ();
 sg13g2_decap_8 FILLER_79_420 ();
 sg13g2_decap_4 FILLER_79_427 ();
 sg13g2_fill_1 FILLER_79_431 ();
 sg13g2_fill_1 FILLER_79_458 ();
 sg13g2_fill_2 FILLER_79_463 ();
 sg13g2_fill_2 FILLER_79_469 ();
 sg13g2_fill_2 FILLER_79_476 ();
 sg13g2_fill_1 FILLER_79_478 ();
 sg13g2_decap_8 FILLER_79_498 ();
 sg13g2_fill_1 FILLER_79_515 ();
 sg13g2_fill_2 FILLER_79_525 ();
 sg13g2_decap_4 FILLER_79_558 ();
 sg13g2_decap_4 FILLER_79_606 ();
 sg13g2_decap_4 FILLER_79_618 ();
 sg13g2_fill_2 FILLER_79_632 ();
 sg13g2_decap_4 FILLER_79_638 ();
 sg13g2_decap_8 FILLER_79_647 ();
 sg13g2_fill_2 FILLER_79_654 ();
 sg13g2_fill_2 FILLER_79_661 ();
 sg13g2_fill_1 FILLER_79_663 ();
 sg13g2_decap_8 FILLER_79_679 ();
 sg13g2_fill_1 FILLER_79_686 ();
 sg13g2_decap_4 FILLER_79_692 ();
 sg13g2_fill_2 FILLER_79_696 ();
 sg13g2_fill_1 FILLER_79_703 ();
 sg13g2_decap_8 FILLER_79_709 ();
 sg13g2_fill_2 FILLER_79_716 ();
 sg13g2_decap_4 FILLER_79_722 ();
 sg13g2_fill_2 FILLER_79_726 ();
 sg13g2_decap_8 FILLER_79_754 ();
 sg13g2_decap_4 FILLER_79_761 ();
 sg13g2_decap_8 FILLER_79_817 ();
 sg13g2_decap_8 FILLER_79_824 ();
 sg13g2_decap_8 FILLER_79_831 ();
 sg13g2_decap_8 FILLER_79_838 ();
 sg13g2_decap_8 FILLER_79_845 ();
 sg13g2_decap_8 FILLER_79_852 ();
 sg13g2_decap_8 FILLER_79_859 ();
 sg13g2_decap_8 FILLER_79_866 ();
 sg13g2_decap_4 FILLER_79_873 ();
 sg13g2_fill_1 FILLER_79_877 ();
 sg13g2_decap_8 FILLER_80_0 ();
 sg13g2_decap_8 FILLER_80_7 ();
 sg13g2_decap_4 FILLER_80_14 ();
 sg13g2_fill_1 FILLER_80_18 ();
 sg13g2_fill_2 FILLER_80_23 ();
 sg13g2_decap_8 FILLER_80_55 ();
 sg13g2_fill_2 FILLER_80_62 ();
 sg13g2_fill_1 FILLER_80_64 ();
 sg13g2_fill_2 FILLER_80_89 ();
 sg13g2_fill_1 FILLER_80_91 ();
 sg13g2_fill_1 FILLER_80_170 ();
 sg13g2_fill_2 FILLER_80_175 ();
 sg13g2_fill_2 FILLER_80_181 ();
 sg13g2_decap_4 FILLER_80_187 ();
 sg13g2_fill_2 FILLER_80_191 ();
 sg13g2_fill_2 FILLER_80_268 ();
 sg13g2_fill_2 FILLER_80_296 ();
 sg13g2_fill_1 FILLER_80_298 ();
 sg13g2_decap_4 FILLER_80_325 ();
 sg13g2_decap_4 FILLER_80_341 ();
 sg13g2_fill_2 FILLER_80_345 ();
 sg13g2_fill_1 FILLER_80_359 ();
 sg13g2_decap_8 FILLER_80_416 ();
 sg13g2_decap_8 FILLER_80_423 ();
 sg13g2_decap_8 FILLER_80_430 ();
 sg13g2_decap_8 FILLER_80_437 ();
 sg13g2_decap_8 FILLER_80_444 ();
 sg13g2_decap_8 FILLER_80_477 ();
 sg13g2_decap_8 FILLER_80_484 ();
 sg13g2_fill_2 FILLER_80_491 ();
 sg13g2_decap_8 FILLER_80_523 ();
 sg13g2_decap_8 FILLER_80_530 ();
 sg13g2_decap_4 FILLER_80_537 ();
 sg13g2_decap_8 FILLER_80_545 ();
 sg13g2_decap_4 FILLER_80_552 ();
 sg13g2_fill_2 FILLER_80_556 ();
 sg13g2_decap_8 FILLER_80_563 ();
 sg13g2_decap_8 FILLER_80_570 ();
 sg13g2_decap_8 FILLER_80_577 ();
 sg13g2_decap_8 FILLER_80_584 ();
 sg13g2_decap_8 FILLER_80_591 ();
 sg13g2_decap_8 FILLER_80_598 ();
 sg13g2_decap_8 FILLER_80_605 ();
 sg13g2_decap_8 FILLER_80_612 ();
 sg13g2_decap_4 FILLER_80_619 ();
 sg13g2_fill_1 FILLER_80_623 ();
 sg13g2_decap_8 FILLER_80_650 ();
 sg13g2_decap_8 FILLER_80_657 ();
 sg13g2_decap_4 FILLER_80_664 ();
 sg13g2_fill_1 FILLER_80_681 ();
 sg13g2_decap_4 FILLER_80_690 ();
 sg13g2_fill_1 FILLER_80_694 ();
 sg13g2_decap_8 FILLER_80_700 ();
 sg13g2_decap_4 FILLER_80_737 ();
 sg13g2_decap_8 FILLER_80_745 ();
 sg13g2_decap_8 FILLER_80_752 ();
 sg13g2_decap_8 FILLER_80_759 ();
 sg13g2_decap_8 FILLER_80_766 ();
 sg13g2_decap_8 FILLER_80_777 ();
 sg13g2_decap_8 FILLER_80_784 ();
 sg13g2_decap_8 FILLER_80_791 ();
 sg13g2_fill_2 FILLER_80_798 ();
 sg13g2_decap_8 FILLER_80_804 ();
 sg13g2_decap_4 FILLER_80_811 ();
 sg13g2_fill_2 FILLER_80_815 ();
 sg13g2_decap_8 FILLER_80_847 ();
 sg13g2_decap_8 FILLER_80_854 ();
 sg13g2_decap_8 FILLER_80_861 ();
 sg13g2_decap_8 FILLER_80_868 ();
 sg13g2_fill_2 FILLER_80_875 ();
 sg13g2_fill_1 FILLER_80_877 ();
endmodule
