module tt_um_rebeccargb_colorbars (clk,
    ena,
    rst_n,
    ui_in,
    uio_in,
    uio_oe,
    uio_out,
    uo_out);
 input clk;
 input ena;
 input rst_n;
 input [7:0] ui_in;
 input [7:0] uio_in;
 output [7:0] uio_oe;
 output [7:0] uio_out;
 output [7:0] uo_out;

 wire _0000_;
 wire _0001_;
 wire _0002_;
 wire _0003_;
 wire _0004_;
 wire _0005_;
 wire _0006_;
 wire _0007_;
 wire _0008_;
 wire _0009_;
 wire _0010_;
 wire _0011_;
 wire _0012_;
 wire _0013_;
 wire _0014_;
 wire _0015_;
 wire _0016_;
 wire _0017_;
 wire _0018_;
 wire _0019_;
 wire _0020_;
 wire _0021_;
 wire _0022_;
 wire _0023_;
 wire _0024_;
 wire _0025_;
 wire _0026_;
 wire _0027_;
 wire _0028_;
 wire _0029_;
 wire _0030_;
 wire _0031_;
 wire _0032_;
 wire _0033_;
 wire _0034_;
 wire _0035_;
 wire _0036_;
 wire _0037_;
 wire _0038_;
 wire _0039_;
 wire _0040_;
 wire _0041_;
 wire _0042_;
 wire _0043_;
 wire _0044_;
 wire _0045_;
 wire _0046_;
 wire _0047_;
 wire _0048_;
 wire _0049_;
 wire _0050_;
 wire _0051_;
 wire _0052_;
 wire _0053_;
 wire _0054_;
 wire _0055_;
 wire _0056_;
 wire _0057_;
 wire _0058_;
 wire _0059_;
 wire _0060_;
 wire _0061_;
 wire _0062_;
 wire _0063_;
 wire _0064_;
 wire _0065_;
 wire _0066_;
 wire _0067_;
 wire _0068_;
 wire _0069_;
 wire _0070_;
 wire _0071_;
 wire _0072_;
 wire _0073_;
 wire _0074_;
 wire _0075_;
 wire _0076_;
 wire _0077_;
 wire _0078_;
 wire _0079_;
 wire _0080_;
 wire _0081_;
 wire _0082_;
 wire _0083_;
 wire _0084_;
 wire _0085_;
 wire _0086_;
 wire _0087_;
 wire _0088_;
 wire _0089_;
 wire _0090_;
 wire _0091_;
 wire _0092_;
 wire _0093_;
 wire _0094_;
 wire _0095_;
 wire _0096_;
 wire _0097_;
 wire _0098_;
 wire _0099_;
 wire _0100_;
 wire _0101_;
 wire _0102_;
 wire _0103_;
 wire _0104_;
 wire _0105_;
 wire _0106_;
 wire _0107_;
 wire _0108_;
 wire _0109_;
 wire _0110_;
 wire _0111_;
 wire _0112_;
 wire _0113_;
 wire _0114_;
 wire _0115_;
 wire _0116_;
 wire _0117_;
 wire _0118_;
 wire _0119_;
 wire _0120_;
 wire _0121_;
 wire _0122_;
 wire _0123_;
 wire _0124_;
 wire _0125_;
 wire _0126_;
 wire _0127_;
 wire _0128_;
 wire _0129_;
 wire _0130_;
 wire _0131_;
 wire _0132_;
 wire _0133_;
 wire _0134_;
 wire _0135_;
 wire _0136_;
 wire _0137_;
 wire _0138_;
 wire _0139_;
 wire _0140_;
 wire _0141_;
 wire _0142_;
 wire _0143_;
 wire _0144_;
 wire _0145_;
 wire _0146_;
 wire _0147_;
 wire _0148_;
 wire _0149_;
 wire _0150_;
 wire _0151_;
 wire _0152_;
 wire _0153_;
 wire _0154_;
 wire _0155_;
 wire _0156_;
 wire _0157_;
 wire _0158_;
 wire _0159_;
 wire _0160_;
 wire _0161_;
 wire _0162_;
 wire _0163_;
 wire _0164_;
 wire _0165_;
 wire _0166_;
 wire _0167_;
 wire _0168_;
 wire _0169_;
 wire _0170_;
 wire _0171_;
 wire _0172_;
 wire _0173_;
 wire _0174_;
 wire _0175_;
 wire _0176_;
 wire _0177_;
 wire _0178_;
 wire _0179_;
 wire _0180_;
 wire _0181_;
 wire _0182_;
 wire _0183_;
 wire _0184_;
 wire _0185_;
 wire _0186_;
 wire _0187_;
 wire _0188_;
 wire _0189_;
 wire _0190_;
 wire _0191_;
 wire _0192_;
 wire _0193_;
 wire _0194_;
 wire _0195_;
 wire _0196_;
 wire _0197_;
 wire _0198_;
 wire _0199_;
 wire _0200_;
 wire _0201_;
 wire _0202_;
 wire _0203_;
 wire _0204_;
 wire _0205_;
 wire _0206_;
 wire _0207_;
 wire _0208_;
 wire _0209_;
 wire _0210_;
 wire _0211_;
 wire _0212_;
 wire _0213_;
 wire _0214_;
 wire _0215_;
 wire _0216_;
 wire _0217_;
 wire _0218_;
 wire _0219_;
 wire _0220_;
 wire _0221_;
 wire _0222_;
 wire _0223_;
 wire _0224_;
 wire _0225_;
 wire _0226_;
 wire _0227_;
 wire _0228_;
 wire _0229_;
 wire _0230_;
 wire _0231_;
 wire _0232_;
 wire _0233_;
 wire _0234_;
 wire _0235_;
 wire _0236_;
 wire _0237_;
 wire _0238_;
 wire _0239_;
 wire _0240_;
 wire _0241_;
 wire _0242_;
 wire _0243_;
 wire _0244_;
 wire _0245_;
 wire _0246_;
 wire _0247_;
 wire _0248_;
 wire _0249_;
 wire _0250_;
 wire _0251_;
 wire _0252_;
 wire _0253_;
 wire _0254_;
 wire _0255_;
 wire _0256_;
 wire _0257_;
 wire _0258_;
 wire _0259_;
 wire _0260_;
 wire _0261_;
 wire _0262_;
 wire _0263_;
 wire _0264_;
 wire _0265_;
 wire _0266_;
 wire _0267_;
 wire _0268_;
 wire _0269_;
 wire _0270_;
 wire _0271_;
 wire _0272_;
 wire _0273_;
 wire _0274_;
 wire _0275_;
 wire _0276_;
 wire _0277_;
 wire _0278_;
 wire _0279_;
 wire _0280_;
 wire _0281_;
 wire _0282_;
 wire _0283_;
 wire _0284_;
 wire _0285_;
 wire _0286_;
 wire _0287_;
 wire _0288_;
 wire _0289_;
 wire _0290_;
 wire _0291_;
 wire _0292_;
 wire _0293_;
 wire _0294_;
 wire _0295_;
 wire _0296_;
 wire _0297_;
 wire _0298_;
 wire _0299_;
 wire _0300_;
 wire _0301_;
 wire _0302_;
 wire _0303_;
 wire _0304_;
 wire _0305_;
 wire _0306_;
 wire _0307_;
 wire _0308_;
 wire _0309_;
 wire _0310_;
 wire _0311_;
 wire _0312_;
 wire _0313_;
 wire _0314_;
 wire _0315_;
 wire _0316_;
 wire _0317_;
 wire _0318_;
 wire _0319_;
 wire _0320_;
 wire _0321_;
 wire _0322_;
 wire _0323_;
 wire _0324_;
 wire _0325_;
 wire _0326_;
 wire _0327_;
 wire _0328_;
 wire _0329_;
 wire _0330_;
 wire _0331_;
 wire _0332_;
 wire _0333_;
 wire _0334_;
 wire _0335_;
 wire _0336_;
 wire _0337_;
 wire _0338_;
 wire _0339_;
 wire _0340_;
 wire _0341_;
 wire _0342_;
 wire _0343_;
 wire _0344_;
 wire _0345_;
 wire _0346_;
 wire _0347_;
 wire _0348_;
 wire _0349_;
 wire _0350_;
 wire _0351_;
 wire _0352_;
 wire _0353_;
 wire _0354_;
 wire _0355_;
 wire _0356_;
 wire _0357_;
 wire _0358_;
 wire _0359_;
 wire _0360_;
 wire _0361_;
 wire _0362_;
 wire _0363_;
 wire _0364_;
 wire _0365_;
 wire _0366_;
 wire _0367_;
 wire _0368_;
 wire _0369_;
 wire _0370_;
 wire _0371_;
 wire _0372_;
 wire _0373_;
 wire _0374_;
 wire _0375_;
 wire _0376_;
 wire _0377_;
 wire _0378_;
 wire _0379_;
 wire _0380_;
 wire _0381_;
 wire _0382_;
 wire _0383_;
 wire _0384_;
 wire _0385_;
 wire _0386_;
 wire _0387_;
 wire _0388_;
 wire _0389_;
 wire _0390_;
 wire _0391_;
 wire _0392_;
 wire _0393_;
 wire _0394_;
 wire _0395_;
 wire _0396_;
 wire _0397_;
 wire _0398_;
 wire _0399_;
 wire _0400_;
 wire _0401_;
 wire _0402_;
 wire _0403_;
 wire _0404_;
 wire _0405_;
 wire _0406_;
 wire _0407_;
 wire _0408_;
 wire _0409_;
 wire _0410_;
 wire _0411_;
 wire _0412_;
 wire _0413_;
 wire _0414_;
 wire _0415_;
 wire _0416_;
 wire _0417_;
 wire _0418_;
 wire _0419_;
 wire _0420_;
 wire _0421_;
 wire _0422_;
 wire _0423_;
 wire _0424_;
 wire _0425_;
 wire _0426_;
 wire _0427_;
 wire _0428_;
 wire _0429_;
 wire _0430_;
 wire _0431_;
 wire _0432_;
 wire _0433_;
 wire _0434_;
 wire _0435_;
 wire _0436_;
 wire _0437_;
 wire _0438_;
 wire _0439_;
 wire _0440_;
 wire _0441_;
 wire _0442_;
 wire _0443_;
 wire _0444_;
 wire _0445_;
 wire _0446_;
 wire _0447_;
 wire _0448_;
 wire _0449_;
 wire _0450_;
 wire _0451_;
 wire _0452_;
 wire _0453_;
 wire _0454_;
 wire _0455_;
 wire _0456_;
 wire _0457_;
 wire _0458_;
 wire _0459_;
 wire _0460_;
 wire _0461_;
 wire _0462_;
 wire _0463_;
 wire _0464_;
 wire _0465_;
 wire _0466_;
 wire _0467_;
 wire _0468_;
 wire _0469_;
 wire _0470_;
 wire _0471_;
 wire _0472_;
 wire _0473_;
 wire _0474_;
 wire _0475_;
 wire _0476_;
 wire _0477_;
 wire _0478_;
 wire _0479_;
 wire _0480_;
 wire _0481_;
 wire _0482_;
 wire _0483_;
 wire _0484_;
 wire _0485_;
 wire _0486_;
 wire _0487_;
 wire _0488_;
 wire _0489_;
 wire _0490_;
 wire _0491_;
 wire _0492_;
 wire _0493_;
 wire _0494_;
 wire _0495_;
 wire _0496_;
 wire _0497_;
 wire _0498_;
 wire _0499_;
 wire _0500_;
 wire _0501_;
 wire _0502_;
 wire _0503_;
 wire _0504_;
 wire _0505_;
 wire _0506_;
 wire _0507_;
 wire _0508_;
 wire _0509_;
 wire _0510_;
 wire _0511_;
 wire _0512_;
 wire _0513_;
 wire _0514_;
 wire _0515_;
 wire _0516_;
 wire _0517_;
 wire _0518_;
 wire _0519_;
 wire _0520_;
 wire _0521_;
 wire _0522_;
 wire _0523_;
 wire _0524_;
 wire _0525_;
 wire _0526_;
 wire _0527_;
 wire _0528_;
 wire _0529_;
 wire _0530_;
 wire _0531_;
 wire _0532_;
 wire _0533_;
 wire _0534_;
 wire _0535_;
 wire _0536_;
 wire _0537_;
 wire _0538_;
 wire _0539_;
 wire _0540_;
 wire _0541_;
 wire _0542_;
 wire _0543_;
 wire _0544_;
 wire _0545_;
 wire _0546_;
 wire _0547_;
 wire _0548_;
 wire _0549_;
 wire _0550_;
 wire _0551_;
 wire _0552_;
 wire _0553_;
 wire _0554_;
 wire _0555_;
 wire _0556_;
 wire _0557_;
 wire _0558_;
 wire _0559_;
 wire _0560_;
 wire _0561_;
 wire _0562_;
 wire _0563_;
 wire _0564_;
 wire _0565_;
 wire _0566_;
 wire _0567_;
 wire _0568_;
 wire _0569_;
 wire _0570_;
 wire _0571_;
 wire _0572_;
 wire _0573_;
 wire _0574_;
 wire _0575_;
 wire _0576_;
 wire _0577_;
 wire _0578_;
 wire _0579_;
 wire _0580_;
 wire _0581_;
 wire _0582_;
 wire _0583_;
 wire _0584_;
 wire _0585_;
 wire _0586_;
 wire _0587_;
 wire _0588_;
 wire _0589_;
 wire _0590_;
 wire _0591_;
 wire _0592_;
 wire _0593_;
 wire _0594_;
 wire _0595_;
 wire _0596_;
 wire _0597_;
 wire _0598_;
 wire _0599_;
 wire _0600_;
 wire _0601_;
 wire _0602_;
 wire _0603_;
 wire _0604_;
 wire _0605_;
 wire _0606_;
 wire _0607_;
 wire _0608_;
 wire _0609_;
 wire _0610_;
 wire _0611_;
 wire _0612_;
 wire _0613_;
 wire _0614_;
 wire _0615_;
 wire _0616_;
 wire _0617_;
 wire _0618_;
 wire _0619_;
 wire _0620_;
 wire _0621_;
 wire _0622_;
 wire _0623_;
 wire _0624_;
 wire _0625_;
 wire _0626_;
 wire _0627_;
 wire _0628_;
 wire _0629_;
 wire _0630_;
 wire _0631_;
 wire _0632_;
 wire _0633_;
 wire _0634_;
 wire _0635_;
 wire _0636_;
 wire _0637_;
 wire _0638_;
 wire _0639_;
 wire _0640_;
 wire _0641_;
 wire _0642_;
 wire _0643_;
 wire _0644_;
 wire _0645_;
 wire _0646_;
 wire _0647_;
 wire _0648_;
 wire _0649_;
 wire _0650_;
 wire _0651_;
 wire _0652_;
 wire _0653_;
 wire _0654_;
 wire _0655_;
 wire _0656_;
 wire _0657_;
 wire _0658_;
 wire _0659_;
 wire _0660_;
 wire _0661_;
 wire _0662_;
 wire _0663_;
 wire _0664_;
 wire _0665_;
 wire _0666_;
 wire _0667_;
 wire _0668_;
 wire _0669_;
 wire _0670_;
 wire _0671_;
 wire _0672_;
 wire _0673_;
 wire _0674_;
 wire _0675_;
 wire _0676_;
 wire _0677_;
 wire _0678_;
 wire _0679_;
 wire _0680_;
 wire _0681_;
 wire _0682_;
 wire _0683_;
 wire _0684_;
 wire _0685_;
 wire _0686_;
 wire _0687_;
 wire _0688_;
 wire _0689_;
 wire _0690_;
 wire _0691_;
 wire _0692_;
 wire _0693_;
 wire _0694_;
 wire _0695_;
 wire _0696_;
 wire _0697_;
 wire _0698_;
 wire _0699_;
 wire _0700_;
 wire _0701_;
 wire _0702_;
 wire _0703_;
 wire _0704_;
 wire _0705_;
 wire _0706_;
 wire _0707_;
 wire _0708_;
 wire _0709_;
 wire _0710_;
 wire _0711_;
 wire _0712_;
 wire _0713_;
 wire _0714_;
 wire _0715_;
 wire _0716_;
 wire _0717_;
 wire _0718_;
 wire _0719_;
 wire _0720_;
 wire _0721_;
 wire _0722_;
 wire _0723_;
 wire _0724_;
 wire _0725_;
 wire _0726_;
 wire _0727_;
 wire _0728_;
 wire _0729_;
 wire _0730_;
 wire _0731_;
 wire _0732_;
 wire _0733_;
 wire _0734_;
 wire _0735_;
 wire _0736_;
 wire _0737_;
 wire _0738_;
 wire _0739_;
 wire _0740_;
 wire _0741_;
 wire _0742_;
 wire _0743_;
 wire _0744_;
 wire _0745_;
 wire _0746_;
 wire _0747_;
 wire _0748_;
 wire _0749_;
 wire _0750_;
 wire _0751_;
 wire _0752_;
 wire _0753_;
 wire _0754_;
 wire _0755_;
 wire _0756_;
 wire _0757_;
 wire _0758_;
 wire _0759_;
 wire _0760_;
 wire _0761_;
 wire _0762_;
 wire _0763_;
 wire _0764_;
 wire _0765_;
 wire _0766_;
 wire _0767_;
 wire _0768_;
 wire _0769_;
 wire _0770_;
 wire _0771_;
 wire _0772_;
 wire _0773_;
 wire _0774_;
 wire _0775_;
 wire _0776_;
 wire _0777_;
 wire _0778_;
 wire _0779_;
 wire _0780_;
 wire _0781_;
 wire _0782_;
 wire _0783_;
 wire _0784_;
 wire _0785_;
 wire _0786_;
 wire _0787_;
 wire _0788_;
 wire _0789_;
 wire _0790_;
 wire _0791_;
 wire _0792_;
 wire _0793_;
 wire _0794_;
 wire _0795_;
 wire _0796_;
 wire _0797_;
 wire _0798_;
 wire _0799_;
 wire _0800_;
 wire _0801_;
 wire _0802_;
 wire _0803_;
 wire _0804_;
 wire _0805_;
 wire _0806_;
 wire _0807_;
 wire _0808_;
 wire _0809_;
 wire _0810_;
 wire _0811_;
 wire _0812_;
 wire _0813_;
 wire _0814_;
 wire _0815_;
 wire _0816_;
 wire _0817_;
 wire _0818_;
 wire _0819_;
 wire _0820_;
 wire _0821_;
 wire _0822_;
 wire _0823_;
 wire _0824_;
 wire _0825_;
 wire _0826_;
 wire _0827_;
 wire _0828_;
 wire _0829_;
 wire _0830_;
 wire _0831_;
 wire _0832_;
 wire _0833_;
 wire _0834_;
 wire _0835_;
 wire _0836_;
 wire _0837_;
 wire _0838_;
 wire _0839_;
 wire _0840_;
 wire _0841_;
 wire _0842_;
 wire _0843_;
 wire _0844_;
 wire _0845_;
 wire _0846_;
 wire _0847_;
 wire _0848_;
 wire _0849_;
 wire _0850_;
 wire _0851_;
 wire _0852_;
 wire _0853_;
 wire _0854_;
 wire _0855_;
 wire _0856_;
 wire _0857_;
 wire _0858_;
 wire _0859_;
 wire _0860_;
 wire _0861_;
 wire _0862_;
 wire _0863_;
 wire _0864_;
 wire _0865_;
 wire _0866_;
 wire _0867_;
 wire _0868_;
 wire _0869_;
 wire _0870_;
 wire _0871_;
 wire _0872_;
 wire _0873_;
 wire _0874_;
 wire _0875_;
 wire _0876_;
 wire _0877_;
 wire _0878_;
 wire _0879_;
 wire _0880_;
 wire _0881_;
 wire _0882_;
 wire _0883_;
 wire _0884_;
 wire _0885_;
 wire _0886_;
 wire _0887_;
 wire _0888_;
 wire _0889_;
 wire _0890_;
 wire _0891_;
 wire _0892_;
 wire _0893_;
 wire _0894_;
 wire _0895_;
 wire _0896_;
 wire _0897_;
 wire _0898_;
 wire _0899_;
 wire _0900_;
 wire _0901_;
 wire _0902_;
 wire _0903_;
 wire _0904_;
 wire _0905_;
 wire _0906_;
 wire _0907_;
 wire _0908_;
 wire _0909_;
 wire _0910_;
 wire _0911_;
 wire _0912_;
 wire _0913_;
 wire _0914_;
 wire _0915_;
 wire _0916_;
 wire _0917_;
 wire _0918_;
 wire _0919_;
 wire _0920_;
 wire _0921_;
 wire _0922_;
 wire _0923_;
 wire _0924_;
 wire _0925_;
 wire _0926_;
 wire _0927_;
 wire _0928_;
 wire _0929_;
 wire _0930_;
 wire _0931_;
 wire _0932_;
 wire _0933_;
 wire _0934_;
 wire _0935_;
 wire _0936_;
 wire _0937_;
 wire _0938_;
 wire _0939_;
 wire _0940_;
 wire _0941_;
 wire _0942_;
 wire _0943_;
 wire _0944_;
 wire _0945_;
 wire _0946_;
 wire _0947_;
 wire _0948_;
 wire _0949_;
 wire _0950_;
 wire _0951_;
 wire _0952_;
 wire _0953_;
 wire _0954_;
 wire _0955_;
 wire _0956_;
 wire _0957_;
 wire _0958_;
 wire _0959_;
 wire _0960_;
 wire _0961_;
 wire _0962_;
 wire _0963_;
 wire _0964_;
 wire _0965_;
 wire _0966_;
 wire _0967_;
 wire _0968_;
 wire _0969_;
 wire _0970_;
 wire _0971_;
 wire _0972_;
 wire _0973_;
 wire _0974_;
 wire _0975_;
 wire _0976_;
 wire _0977_;
 wire _0978_;
 wire _0979_;
 wire _0980_;
 wire _0981_;
 wire _0982_;
 wire _0983_;
 wire _0984_;
 wire _0985_;
 wire _0986_;
 wire _0987_;
 wire _0988_;
 wire _0989_;
 wire _0990_;
 wire _0991_;
 wire _0992_;
 wire _0993_;
 wire _0994_;
 wire _0995_;
 wire _0996_;
 wire _0997_;
 wire _0998_;
 wire _0999_;
 wire _1000_;
 wire _1001_;
 wire _1002_;
 wire _1003_;
 wire _1004_;
 wire _1005_;
 wire _1006_;
 wire _1007_;
 wire _1008_;
 wire _1009_;
 wire _1010_;
 wire _1011_;
 wire _1012_;
 wire _1013_;
 wire _1014_;
 wire _1015_;
 wire _1016_;
 wire _1017_;
 wire _1018_;
 wire _1019_;
 wire _1020_;
 wire _1021_;
 wire _1022_;
 wire _1023_;
 wire _1024_;
 wire _1025_;
 wire _1026_;
 wire _1027_;
 wire _1028_;
 wire _1029_;
 wire _1030_;
 wire _1031_;
 wire _1032_;
 wire _1033_;
 wire _1034_;
 wire _1035_;
 wire _1036_;
 wire _1037_;
 wire _1038_;
 wire _1039_;
 wire _1040_;
 wire _1041_;
 wire _1042_;
 wire _1043_;
 wire _1044_;
 wire _1045_;
 wire _1046_;
 wire _1047_;
 wire _1048_;
 wire _1049_;
 wire _1050_;
 wire _1051_;
 wire _1052_;
 wire _1053_;
 wire _1054_;
 wire _1055_;
 wire _1056_;
 wire _1057_;
 wire _1058_;
 wire _1059_;
 wire _1060_;
 wire _1061_;
 wire _1062_;
 wire _1063_;
 wire _1064_;
 wire _1065_;
 wire _1066_;
 wire _1067_;
 wire _1068_;
 wire _1069_;
 wire _1070_;
 wire _1071_;
 wire _1072_;
 wire _1073_;
 wire _1074_;
 wire _1075_;
 wire _1076_;
 wire _1077_;
 wire _1078_;
 wire _1079_;
 wire _1080_;
 wire _1081_;
 wire _1082_;
 wire _1083_;
 wire _1084_;
 wire _1085_;
 wire _1086_;
 wire _1087_;
 wire _1088_;
 wire _1089_;
 wire _1090_;
 wire _1091_;
 wire _1092_;
 wire _1093_;
 wire _1094_;
 wire _1095_;
 wire _1096_;
 wire _1097_;
 wire _1098_;
 wire _1099_;
 wire _1100_;
 wire _1101_;
 wire _1102_;
 wire _1103_;
 wire _1104_;
 wire _1105_;
 wire _1106_;
 wire _1107_;
 wire _1108_;
 wire _1109_;
 wire _1110_;
 wire _1111_;
 wire _1112_;
 wire _1113_;
 wire _1114_;
 wire _1115_;
 wire _1116_;
 wire _1117_;
 wire _1118_;
 wire _1119_;
 wire _1120_;
 wire _1121_;
 wire _1122_;
 wire _1123_;
 wire _1124_;
 wire _1125_;
 wire _1126_;
 wire _1127_;
 wire _1128_;
 wire _1129_;
 wire _1130_;
 wire _1131_;
 wire _1132_;
 wire _1133_;
 wire _1134_;
 wire _1135_;
 wire _1136_;
 wire _1137_;
 wire _1138_;
 wire _1139_;
 wire _1140_;
 wire _1141_;
 wire _1142_;
 wire _1143_;
 wire _1144_;
 wire _1145_;
 wire _1146_;
 wire _1147_;
 wire _1148_;
 wire _1149_;
 wire _1150_;
 wire _1151_;
 wire _1152_;
 wire _1153_;
 wire _1154_;
 wire _1155_;
 wire _1156_;
 wire _1157_;
 wire _1158_;
 wire _1159_;
 wire _1160_;
 wire _1161_;
 wire _1162_;
 wire _1163_;
 wire _1164_;
 wire _1165_;
 wire _1166_;
 wire _1167_;
 wire _1168_;
 wire _1169_;
 wire _1170_;
 wire _1171_;
 wire _1172_;
 wire _1173_;
 wire _1174_;
 wire _1175_;
 wire _1176_;
 wire _1177_;
 wire _1178_;
 wire _1179_;
 wire _1180_;
 wire _1181_;
 wire _1182_;
 wire _1183_;
 wire _1184_;
 wire _1185_;
 wire _1186_;
 wire _1187_;
 wire _1188_;
 wire _1189_;
 wire _1190_;
 wire _1191_;
 wire _1192_;
 wire _1193_;
 wire _1194_;
 wire _1195_;
 wire _1196_;
 wire _1197_;
 wire _1198_;
 wire _1199_;
 wire _1200_;
 wire _1201_;
 wire _1202_;
 wire _1203_;
 wire _1204_;
 wire _1205_;
 wire _1206_;
 wire _1207_;
 wire _1208_;
 wire _1209_;
 wire _1210_;
 wire _1211_;
 wire _1212_;
 wire _1213_;
 wire _1214_;
 wire _1215_;
 wire _1216_;
 wire _1217_;
 wire _1218_;
 wire _1219_;
 wire _1220_;
 wire _1221_;
 wire _1222_;
 wire _1223_;
 wire _1224_;
 wire _1225_;
 wire _1226_;
 wire _1227_;
 wire _1228_;
 wire _1229_;
 wire _1230_;
 wire _1231_;
 wire _1232_;
 wire _1233_;
 wire _1234_;
 wire _1235_;
 wire _1236_;
 wire _1237_;
 wire _1238_;
 wire _1239_;
 wire _1240_;
 wire _1241_;
 wire _1242_;
 wire _1243_;
 wire _1244_;
 wire _1245_;
 wire _1246_;
 wire _1247_;
 wire _1248_;
 wire _1249_;
 wire _1250_;
 wire _1251_;
 wire _1252_;
 wire _1253_;
 wire _1254_;
 wire _1255_;
 wire _1256_;
 wire _1257_;
 wire _1258_;
 wire _1259_;
 wire _1260_;
 wire _1261_;
 wire _1262_;
 wire _1263_;
 wire _1264_;
 wire _1265_;
 wire _1266_;
 wire _1267_;
 wire _1268_;
 wire _1269_;
 wire _1270_;
 wire _1271_;
 wire _1272_;
 wire _1273_;
 wire clknet_0_clk;
 wire \counter[0] ;
 wire \counter[1] ;
 wire \counter[2] ;
 wire \counter[3] ;
 wire \counter[4] ;
 wire \counter[5] ;
 wire \counter[6] ;
 wire \counter[7] ;
 wire \counter[8] ;
 wire \counter[9] ;
 wire hsync;
 wire \hvsync_gen.hpos[0] ;
 wire \hvsync_gen.hpos[1] ;
 wire \hvsync_gen.hpos[2] ;
 wire \hvsync_gen.hpos[3] ;
 wire \hvsync_gen.hpos[4] ;
 wire \hvsync_gen.hpos[5] ;
 wire \hvsync_gen.hpos[6] ;
 wire \hvsync_gen.hpos[7] ;
 wire \hvsync_gen.hpos[8] ;
 wire \hvsync_gen.hpos[9] ;
 wire \hvsync_gen.vpos[0] ;
 wire \hvsync_gen.vpos[1] ;
 wire \hvsync_gen.vpos[2] ;
 wire \hvsync_gen.vpos[3] ;
 wire \hvsync_gen.vpos[4] ;
 wire \hvsync_gen.vpos[5] ;
 wire \hvsync_gen.vpos[6] ;
 wire \hvsync_gen.vpos[7] ;
 wire \hvsync_gen.vpos[8] ;
 wire \hvsync_gen.vpos[9] ;
 wire \hvsync_gen.vsync ;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net130;
 wire net131;
 wire net132;
 wire clknet_2_0__leaf_clk;
 wire clknet_2_1__leaf_clk;
 wire clknet_2_2__leaf_clk;
 wire clknet_2_3__leaf_clk;

 sg13g2_buf_1 _1275_ (.A(\hvsync_gen.vpos[9] ),
    .X(_0079_));
 sg13g2_buf_1 _1276_ (.A(\hvsync_gen.vpos[8] ),
    .X(_0090_));
 sg13g2_buf_1 _1277_ (.A(_0090_),
    .X(_0101_));
 sg13g2_buf_1 _1278_ (.A(\hvsync_gen.vpos[7] ),
    .X(_0112_));
 sg13g2_buf_8 _1279_ (.A(\hvsync_gen.vpos[6] ),
    .X(_0123_));
 sg13g2_buf_1 _1280_ (.A(_0123_),
    .X(_0134_));
 sg13g2_buf_1 _1281_ (.A(\hvsync_gen.vpos[5] ),
    .X(_0145_));
 sg13g2_nand4_1 _1282_ (.B(net89),
    .C(net79),
    .A(net80),
    .Y(_0156_),
    .D(net88));
 sg13g2_buf_1 _1283_ (.A(\hvsync_gen.vpos[3] ),
    .X(_0167_));
 sg13g2_buf_1 _1284_ (.A(_0167_),
    .X(_0178_));
 sg13g2_buf_1 _1285_ (.A(\hvsync_gen.vpos[1] ),
    .X(_0189_));
 sg13g2_nand2_1 _1286_ (.Y(_0200_),
    .A(net78),
    .B(net87));
 sg13g2_buf_8 _1287_ (.A(\hvsync_gen.vpos[4] ),
    .X(_0211_));
 sg13g2_buf_1 _1288_ (.A(_0211_),
    .X(_0222_));
 sg13g2_inv_1 _1289_ (.Y(_0233_),
    .A(net77));
 sg13g2_buf_2 _1290_ (.A(\hvsync_gen.vpos[2] ),
    .X(_0244_));
 sg13g2_inv_1 _1291_ (.Y(_0255_),
    .A(_0244_));
 sg13g2_buf_1 _1292_ (.A(_0255_),
    .X(_0266_));
 sg13g2_nand2_1 _1293_ (.Y(_0277_),
    .A(_0233_),
    .B(net59));
 sg13g2_nor4_1 _1294_ (.A(net90),
    .B(_0156_),
    .C(_0200_),
    .D(_0277_),
    .Y(_0001_));
 sg13g2_buf_2 _1295_ (.A(\hvsync_gen.hpos[9] ),
    .X(_0298_));
 sg13g2_inv_2 _1296_ (.Y(_0309_),
    .A(_0298_));
 sg13g2_buf_1 _1297_ (.A(\hvsync_gen.hpos[7] ),
    .X(_0320_));
 sg13g2_buf_1 _1298_ (.A(_0320_),
    .X(_0331_));
 sg13g2_buf_1 _1299_ (.A(\hvsync_gen.hpos[6] ),
    .X(_0342_));
 sg13g2_buf_1 _1300_ (.A(_0342_),
    .X(_0353_));
 sg13g2_inv_2 _1301_ (.Y(_0364_),
    .A(_0353_));
 sg13g2_buf_2 _1302_ (.A(\hvsync_gen.hpos[5] ),
    .X(_0375_));
 sg13g2_inv_2 _1303_ (.Y(_0386_),
    .A(_0375_));
 sg13g2_buf_1 _1304_ (.A(\hvsync_gen.hpos[4] ),
    .X(_0397_));
 sg13g2_inv_2 _1305_ (.Y(_0408_),
    .A(net86));
 sg13g2_nand3_1 _1306_ (.B(_0386_),
    .C(_0408_),
    .A(_0364_),
    .Y(_0419_));
 sg13g2_buf_2 _1307_ (.A(\hvsync_gen.hpos[8] ),
    .X(_0428_));
 sg13g2_buf_1 _1308_ (.A(_0428_),
    .X(_0434_));
 sg13g2_buf_1 _1309_ (.A(_0434_),
    .X(_0435_));
 sg13g2_a21oi_1 _1310_ (.A1(net76),
    .A2(_0419_),
    .Y(_0436_),
    .B1(net58));
 sg13g2_buf_1 _1311_ (.A(_0375_),
    .X(_0437_));
 sg13g2_and3_1 _1312_ (.X(_0438_),
    .A(net76),
    .B(net75),
    .C(_0437_));
 sg13g2_buf_1 _1313_ (.A(_0438_),
    .X(_0439_));
 sg13g2_a21oi_1 _1314_ (.A1(net86),
    .A2(_0439_),
    .Y(_0440_),
    .B1(net58));
 sg13g2_nor2_1 _1315_ (.A(_0006_),
    .B(_0440_),
    .Y(_0441_));
 sg13g2_nor3_1 _1316_ (.A(_0309_),
    .B(_0436_),
    .C(_0441_),
    .Y(_0000_));
 sg13g2_buf_1 _1317_ (.A(ui_in[2]),
    .X(_0442_));
 sg13g2_inv_1 _1318_ (.Y(_0443_),
    .A(_0442_));
 sg13g2_inv_2 _1319_ (.Y(_0444_),
    .A(_0015_));
 sg13g2_nand3_1 _1320_ (.B(_0298_),
    .C(_0444_),
    .A(net85),
    .Y(_0445_));
 sg13g2_buf_1 _1321_ (.A(_0442_),
    .X(_0446_));
 sg13g2_inv_2 _1322_ (.Y(_0447_),
    .A(_0428_));
 sg13g2_nor2_1 _1323_ (.A(net84),
    .B(_0447_),
    .Y(_0448_));
 sg13g2_buf_1 _1324_ (.A(\counter[4] ),
    .X(_0449_));
 sg13g2_nand2_1 _1325_ (.Y(_0450_),
    .A(net72),
    .B(net86));
 sg13g2_nor2_1 _1326_ (.A(net72),
    .B(\hvsync_gen.hpos[4] ),
    .Y(_0451_));
 sg13g2_nor2_1 _1327_ (.A(\counter[3] ),
    .B(\hvsync_gen.hpos[3] ),
    .Y(_0452_));
 sg13g2_or2_1 _1328_ (.X(_0453_),
    .B(_0452_),
    .A(_0451_));
 sg13g2_nand2_1 _1329_ (.Y(_0454_),
    .A(_0450_),
    .B(_0453_));
 sg13g2_buf_2 _1330_ (.A(\counter[2] ),
    .X(_0455_));
 sg13g2_buf_1 _1331_ (.A(\hvsync_gen.hpos[2] ),
    .X(_0456_));
 sg13g2_buf_2 _1332_ (.A(\hvsync_gen.hpos[0] ),
    .X(_0457_));
 sg13g2_buf_2 _1333_ (.A(\hvsync_gen.hpos[1] ),
    .X(_0458_));
 sg13g2_a21o_1 _1334_ (.A2(_0457_),
    .A1(\counter[0] ),
    .B1(_0458_),
    .X(_0459_));
 sg13g2_buf_1 _1335_ (.A(\counter[1] ),
    .X(_0460_));
 sg13g2_buf_1 _1336_ (.A(\counter[0] ),
    .X(_0461_));
 sg13g2_and3_1 _1337_ (.X(_0462_),
    .A(net69),
    .B(_0458_),
    .C(_0457_));
 sg13g2_a221oi_1 _1338_ (.B2(net70),
    .C1(_0462_),
    .B1(_0459_),
    .A1(net71),
    .Y(_0463_),
    .A2(_0456_));
 sg13g2_buf_2 _1339_ (.A(_0463_),
    .X(_0464_));
 sg13g2_nor2_2 _1340_ (.A(_0455_),
    .B(_0456_),
    .Y(_0465_));
 sg13g2_buf_1 _1341_ (.A(\hvsync_gen.hpos[3] ),
    .X(_0466_));
 sg13g2_a22oi_1 _1342_ (.Y(_0467_),
    .B1(_0449_),
    .B2(\hvsync_gen.hpos[4] ),
    .A2(net83),
    .A1(\counter[3] ));
 sg13g2_o21ai_1 _1343_ (.B1(_0467_),
    .Y(_0468_),
    .A1(_0464_),
    .A2(_0465_));
 sg13g2_buf_1 _1344_ (.A(\counter[5] ),
    .X(_0469_));
 sg13g2_nand2_1 _1345_ (.Y(_0470_),
    .A(net68),
    .B(_0375_));
 sg13g2_nor2_1 _1346_ (.A(\counter[6] ),
    .B(_0342_),
    .Y(_0471_));
 sg13g2_nand2_1 _1347_ (.Y(_0472_),
    .A(\counter[6] ),
    .B(_0342_));
 sg13g2_o21ai_1 _1348_ (.B1(_0472_),
    .Y(_0473_),
    .A1(_0470_),
    .A2(net67));
 sg13g2_xor2_1 _1349_ (.B(_0320_),
    .A(\counter[7] ),
    .X(_0474_));
 sg13g2_xnor2_1 _1350_ (.Y(_0475_),
    .A(_0473_),
    .B(_0474_));
 sg13g2_a21oi_1 _1351_ (.A1(_0454_),
    .A2(_0468_),
    .Y(_0476_),
    .B1(_0475_));
 sg13g2_nor2_2 _1352_ (.A(net68),
    .B(_0375_),
    .Y(_0477_));
 sg13g2_a21oi_1 _1353_ (.A1(_0477_),
    .A2(_0472_),
    .Y(_0478_),
    .B1(net67));
 sg13g2_xor2_1 _1354_ (.B(_0474_),
    .A(_0478_),
    .X(_0479_));
 sg13g2_and3_1 _1355_ (.X(_0480_),
    .A(_0454_),
    .B(_0468_),
    .C(_0479_));
 sg13g2_buf_2 _1356_ (.A(\counter[9] ),
    .X(_0481_));
 sg13g2_xnor2_1 _1357_ (.Y(_0482_),
    .A(_0481_),
    .B(_0298_));
 sg13g2_inv_1 _1358_ (.Y(_0483_),
    .A(_0482_));
 sg13g2_buf_1 _1359_ (.A(\counter[8] ),
    .X(_0484_));
 sg13g2_buf_1 _1360_ (.A(\counter[7] ),
    .X(_0485_));
 sg13g2_nor2_1 _1361_ (.A(net66),
    .B(_0320_),
    .Y(_0486_));
 sg13g2_nor2_1 _1362_ (.A(_0484_),
    .B(_0428_),
    .Y(_0487_));
 sg13g2_nor2_1 _1363_ (.A(_0486_),
    .B(_0487_),
    .Y(_0488_));
 sg13g2_a21o_1 _1364_ (.A2(_0428_),
    .A1(_0484_),
    .B1(_0488_),
    .X(_0489_));
 sg13g2_xnor2_1 _1365_ (.Y(_0490_),
    .A(_0483_),
    .B(_0489_));
 sg13g2_or3_1 _1366_ (.A(_0476_),
    .B(_0480_),
    .C(_0490_),
    .X(_0491_));
 sg13g2_buf_1 _1367_ (.A(_0491_),
    .X(_0492_));
 sg13g2_nand2_1 _1368_ (.Y(_0493_),
    .A(\counter[3] ),
    .B(net83));
 sg13g2_nor3_1 _1369_ (.A(_0477_),
    .B(_0451_),
    .C(_0493_),
    .Y(_0494_));
 sg13g2_o21ai_1 _1370_ (.B1(_0470_),
    .Y(_0495_),
    .A1(_0477_),
    .A2(_0450_));
 sg13g2_a22oi_1 _1371_ (.Y(_0496_),
    .B1(_0484_),
    .B2(_0428_),
    .A2(_0320_),
    .A1(\counter[7] ));
 sg13g2_nand2_1 _1372_ (.Y(_0497_),
    .A(_0481_),
    .B(_0298_));
 sg13g2_o21ai_1 _1373_ (.B1(_0497_),
    .Y(_0498_),
    .A1(_0487_),
    .A2(_0496_));
 sg13g2_nor4_1 _1374_ (.A(_0342_),
    .B(_0494_),
    .C(_0495_),
    .D(_0498_),
    .Y(_0499_));
 sg13g2_buf_1 _1375_ (.A(\counter[6] ),
    .X(_0500_));
 sg13g2_nor4_1 _1376_ (.A(net65),
    .B(_0494_),
    .C(_0495_),
    .D(_0498_),
    .Y(_0501_));
 sg13g2_or4_1 _1377_ (.A(_0477_),
    .B(_0464_),
    .C(_0453_),
    .D(_0465_),
    .X(_0502_));
 sg13g2_o21ai_1 _1378_ (.B1(_0502_),
    .Y(_0503_),
    .A1(_0499_),
    .A2(_0501_));
 sg13g2_or2_1 _1379_ (.X(_0504_),
    .B(_0342_),
    .A(net65));
 sg13g2_a21o_1 _1380_ (.A2(_0488_),
    .A1(_0504_),
    .B1(_0498_),
    .X(_0505_));
 sg13g2_or2_1 _1381_ (.X(_0506_),
    .B(_0298_),
    .A(_0481_));
 sg13g2_nand3_1 _1382_ (.B(_0505_),
    .C(_0506_),
    .A(_0503_),
    .Y(_0507_));
 sg13g2_and3_1 _1383_ (.X(_0508_),
    .A(net84),
    .B(_0492_),
    .C(_0507_));
 sg13g2_and3_1 _1384_ (.X(_0509_),
    .A(_0503_),
    .B(_0505_),
    .C(_0506_));
 sg13g2_buf_2 _1385_ (.A(_0509_),
    .X(_0510_));
 sg13g2_nor2_1 _1386_ (.A(_0487_),
    .B(_0496_),
    .Y(_0511_));
 sg13g2_xnor2_1 _1387_ (.Y(_0512_),
    .A(_0483_),
    .B(_0511_));
 sg13g2_o21ai_1 _1388_ (.B1(_0512_),
    .Y(_0513_),
    .A1(_0476_),
    .A2(_0480_));
 sg13g2_buf_1 _1389_ (.A(_0513_),
    .X(_0514_));
 sg13g2_and3_1 _1390_ (.X(_0515_),
    .A(net84),
    .B(_0510_),
    .C(_0514_));
 sg13g2_xnor2_1 _1391_ (.Y(_0516_),
    .A(_0484_),
    .B(_0434_));
 sg13g2_or2_1 _1392_ (.X(_0517_),
    .B(_0375_),
    .A(net68));
 sg13g2_buf_1 _1393_ (.A(_0517_),
    .X(_0518_));
 sg13g2_o21ai_1 _1394_ (.B1(_0470_),
    .Y(_0519_),
    .A1(_0451_),
    .A2(_0467_));
 sg13g2_buf_1 _1395_ (.A(_0519_),
    .X(_0520_));
 sg13g2_or2_1 _1396_ (.X(_0521_),
    .B(_0342_),
    .A(_0320_));
 sg13g2_buf_1 _1397_ (.A(_0521_),
    .X(_0522_));
 sg13g2_or2_1 _1398_ (.X(_0523_),
    .B(_0342_),
    .A(net66));
 sg13g2_nor4_2 _1399_ (.A(_0477_),
    .B(_0464_),
    .C(_0453_),
    .Y(_0524_),
    .D(_0465_));
 sg13g2_a221oi_1 _1400_ (.B2(_0523_),
    .C1(_0524_),
    .B1(_0522_),
    .A1(_0518_),
    .Y(_0525_),
    .A2(_0520_));
 sg13g2_or2_1 _1401_ (.X(_0526_),
    .B(net65),
    .A(_0331_));
 sg13g2_or2_1 _1402_ (.X(_0527_),
    .B(\counter[6] ),
    .A(net66));
 sg13g2_a221oi_1 _1403_ (.B2(_0527_),
    .C1(_0524_),
    .B1(_0526_),
    .A1(_0518_),
    .Y(_0528_),
    .A2(_0520_));
 sg13g2_a21oi_1 _1404_ (.A1(_0526_),
    .A2(_0527_),
    .Y(_0529_),
    .B1(net75));
 sg13g2_or4_1 _1405_ (.A(_0486_),
    .B(_0525_),
    .C(_0528_),
    .D(_0529_),
    .X(_0530_));
 sg13g2_xnor2_1 _1406_ (.Y(_0531_),
    .A(_0516_),
    .B(_0530_));
 sg13g2_mux2_1 _1407_ (.A0(_0508_),
    .A1(_0515_),
    .S(_0531_),
    .X(_0532_));
 sg13g2_a21o_1 _1408_ (.A2(_0520_),
    .A1(_0518_),
    .B1(_0524_),
    .X(_0533_));
 sg13g2_xor2_1 _1409_ (.B(_0533_),
    .A(net65),
    .X(_0534_));
 sg13g2_nand2_1 _1410_ (.Y(_0535_),
    .A(_0442_),
    .B(_0534_));
 sg13g2_xnor2_1 _1411_ (.Y(_0536_),
    .A(_0364_),
    .B(_0535_));
 sg13g2_o21ai_1 _1412_ (.B1(_0536_),
    .Y(_0537_),
    .A1(_0448_),
    .A2(_0532_));
 sg13g2_nand2_1 _1413_ (.Y(_0538_),
    .A(_0445_),
    .B(_0537_));
 sg13g2_nand2_1 _1414_ (.Y(_0539_),
    .A(_0503_),
    .B(_0505_));
 sg13g2_or2_1 _1415_ (.X(_0540_),
    .B(_0539_),
    .A(_0492_));
 sg13g2_or2_1 _1416_ (.X(_0541_),
    .B(_0514_),
    .A(_0539_));
 sg13g2_mux2_1 _1417_ (.A0(_0540_),
    .A1(_0541_),
    .S(_0531_),
    .X(_0542_));
 sg13g2_nor2_1 _1418_ (.A(_0492_),
    .B(_0510_),
    .Y(_0543_));
 sg13g2_a21oi_1 _1419_ (.A1(_0531_),
    .A2(_0543_),
    .Y(_0544_),
    .B1(net85));
 sg13g2_a21oi_1 _1420_ (.A1(_0531_),
    .A2(_0543_),
    .Y(_0545_),
    .B1(_0506_));
 sg13g2_a221oi_1 _1421_ (.B2(_0544_),
    .C1(_0545_),
    .B1(_0542_),
    .A1(net85),
    .Y(_0546_),
    .A2(_0309_));
 sg13g2_buf_1 _1422_ (.A(_0546_),
    .X(_0547_));
 sg13g2_buf_2 _1423_ (.A(_0547_),
    .X(_0548_));
 sg13g2_buf_1 _1424_ (.A(_0484_),
    .X(_0549_));
 sg13g2_a221oi_1 _1425_ (.B2(_0520_),
    .C1(_0524_),
    .B1(_0518_),
    .A1(_0500_),
    .Y(_0550_),
    .A2(net75));
 sg13g2_buf_1 _1426_ (.A(_0550_),
    .X(_0551_));
 sg13g2_nor3_2 _1427_ (.A(_0485_),
    .B(_0331_),
    .C(_0428_),
    .Y(_0552_));
 sg13g2_nand2_1 _1428_ (.Y(_0553_),
    .A(_0485_),
    .B(net76));
 sg13g2_nor3_1 _1429_ (.A(_0447_),
    .B(net67),
    .C(_0553_),
    .Y(_0554_));
 sg13g2_nor2_1 _1430_ (.A(_0447_),
    .B(_0553_),
    .Y(_0555_));
 sg13g2_nand2b_1 _1431_ (.Y(_0556_),
    .B(_0555_),
    .A_N(_0472_));
 sg13g2_nand2_1 _1432_ (.Y(_0557_),
    .A(net67),
    .B(_0552_));
 sg13g2_nand3_1 _1433_ (.B(_0556_),
    .C(_0557_),
    .A(_0482_),
    .Y(_0558_));
 sg13g2_a221oi_1 _1434_ (.B2(_0533_),
    .C1(_0558_),
    .B1(_0554_),
    .A1(_0551_),
    .Y(_0559_),
    .A2(_0552_));
 sg13g2_nor3_1 _1435_ (.A(_0549_),
    .B(_0507_),
    .C(_0559_),
    .Y(_0560_));
 sg13g2_or2_1 _1436_ (.X(_0561_),
    .B(_0482_),
    .A(_0474_));
 sg13g2_nor4_1 _1437_ (.A(net67),
    .B(_0551_),
    .C(_0552_),
    .D(_0561_),
    .Y(_0562_));
 sg13g2_or2_1 _1438_ (.X(_0563_),
    .B(_0552_),
    .A(_0482_));
 sg13g2_nor4_1 _1439_ (.A(net74),
    .B(net67),
    .C(_0551_),
    .D(_0563_),
    .Y(_0564_));
 sg13g2_a21oi_1 _1440_ (.A1(_0518_),
    .A2(_0520_),
    .Y(_0565_),
    .B1(_0500_));
 sg13g2_a21oi_1 _1441_ (.A1(_0518_),
    .A2(_0520_),
    .Y(_0566_),
    .B1(net75));
 sg13g2_o21ai_1 _1442_ (.B1(_0502_),
    .Y(_0567_),
    .A1(_0565_),
    .A2(_0566_));
 sg13g2_nand3_1 _1443_ (.B(_0483_),
    .C(_0553_),
    .A(net74),
    .Y(_0568_));
 sg13g2_or2_1 _1444_ (.X(_0569_),
    .B(_0561_),
    .A(_0555_));
 sg13g2_a22oi_1 _1445_ (.Y(_0570_),
    .B1(_0568_),
    .B2(_0569_),
    .A2(_0567_),
    .A1(_0504_));
 sg13g2_nor3_1 _1446_ (.A(_0562_),
    .B(_0564_),
    .C(_0570_),
    .Y(_0571_));
 sg13g2_o21ai_1 _1447_ (.B1(_0514_),
    .Y(_0572_),
    .A1(_0492_),
    .A2(_0510_));
 sg13g2_xor2_1 _1448_ (.B(_0530_),
    .A(_0516_),
    .X(_0573_));
 sg13g2_a221oi_1 _1449_ (.B2(_0573_),
    .C1(net85),
    .B1(_0572_),
    .A1(_0560_),
    .Y(_0574_),
    .A2(_0571_));
 sg13g2_nor2_1 _1450_ (.A(net74),
    .B(_0553_),
    .Y(_0575_));
 sg13g2_a21oi_1 _1451_ (.A1(net74),
    .A2(_0486_),
    .Y(_0576_),
    .B1(_0575_));
 sg13g2_nor2_1 _1452_ (.A(_0482_),
    .B(_0576_),
    .Y(_0577_));
 sg13g2_o21ai_1 _1453_ (.B1(_0577_),
    .Y(_0578_),
    .A1(net67),
    .A2(_0551_));
 sg13g2_or4_1 _1454_ (.A(net67),
    .B(_0551_),
    .C(_0483_),
    .D(_0576_),
    .X(_0579_));
 sg13g2_and3_1 _1455_ (.X(_0580_),
    .A(_0447_),
    .B(_0474_),
    .C(_0483_));
 sg13g2_nand3_1 _1456_ (.B(_0567_),
    .C(_0580_),
    .A(_0504_),
    .Y(_0581_));
 sg13g2_and3_1 _1457_ (.X(_0582_),
    .A(net74),
    .B(_0474_),
    .C(_0482_));
 sg13g2_o21ai_1 _1458_ (.B1(_0582_),
    .Y(_0583_),
    .A1(_0471_),
    .A2(_0551_));
 sg13g2_nand4_1 _1459_ (.B(_0579_),
    .C(_0581_),
    .A(_0578_),
    .Y(_0584_),
    .D(_0583_));
 sg13g2_and2_1 _1460_ (.A(_0549_),
    .B(_0510_),
    .X(_0585_));
 sg13g2_nor2_1 _1461_ (.A(_0510_),
    .B(_0514_),
    .Y(_0586_));
 sg13g2_a21oi_1 _1462_ (.A1(_0584_),
    .A2(_0585_),
    .Y(_0587_),
    .B1(_0586_));
 sg13g2_nor2_1 _1463_ (.A(_0446_),
    .B(_0444_),
    .Y(_0588_));
 sg13g2_a21oi_2 _1464_ (.B1(_0588_),
    .Y(_0589_),
    .A2(_0587_),
    .A1(_0574_));
 sg13g2_nor2_1 _1465_ (.A(net41),
    .B(_0589_),
    .Y(_0590_));
 sg13g2_a21o_1 _1466_ (.A2(_0587_),
    .A1(_0574_),
    .B1(_0588_),
    .X(_0591_));
 sg13g2_buf_1 _1467_ (.A(_0591_),
    .X(_0592_));
 sg13g2_nand2_2 _1468_ (.Y(_0593_),
    .A(net85),
    .B(net74));
 sg13g2_nand3_1 _1469_ (.B(_0492_),
    .C(_0507_),
    .A(_0446_),
    .Y(_0594_));
 sg13g2_nand3_1 _1470_ (.B(_0510_),
    .C(_0514_),
    .A(_0442_),
    .Y(_0595_));
 sg13g2_mux2_1 _1471_ (.A0(_0594_),
    .A1(_0595_),
    .S(_0531_),
    .X(_0596_));
 sg13g2_xnor2_1 _1472_ (.Y(_0597_),
    .A(net75),
    .B(_0535_));
 sg13g2_a21oi_2 _1473_ (.B1(_0597_),
    .Y(_0598_),
    .A2(_0596_),
    .A1(_0593_));
 sg13g2_o21ai_1 _1474_ (.B1(_0598_),
    .Y(_0599_),
    .A1(net41),
    .A2(_0592_));
 sg13g2_o21ai_1 _1475_ (.B1(_0599_),
    .Y(_0600_),
    .A1(_0538_),
    .A2(_0590_));
 sg13g2_nand2_1 _1476_ (.Y(_0601_),
    .A(_0492_),
    .B(_0507_));
 sg13g2_nand2_1 _1477_ (.Y(_0602_),
    .A(_0510_),
    .B(_0514_));
 sg13g2_mux2_1 _1478_ (.A0(_0601_),
    .A1(_0602_),
    .S(_0531_),
    .X(_0603_));
 sg13g2_xnor2_1 _1479_ (.Y(_0604_),
    .A(_0353_),
    .B(_0534_));
 sg13g2_nor2_1 _1480_ (.A(net85),
    .B(_0604_),
    .Y(_0605_));
 sg13g2_nor3_1 _1481_ (.A(net84),
    .B(_0364_),
    .C(net74),
    .Y(_0606_));
 sg13g2_a21o_1 _1482_ (.A2(_0605_),
    .A1(_0603_),
    .B1(_0606_),
    .X(_0607_));
 sg13g2_buf_1 _1483_ (.A(_0607_),
    .X(_0608_));
 sg13g2_nand2_1 _1484_ (.Y(_0609_),
    .A(_0454_),
    .B(_0468_));
 sg13g2_xnor2_1 _1485_ (.Y(_0610_),
    .A(_0469_),
    .B(_0609_));
 sg13g2_nand2_1 _1486_ (.Y(_0611_),
    .A(net84),
    .B(_0610_));
 sg13g2_xnor2_1 _1487_ (.Y(_0612_),
    .A(_0375_),
    .B(_0611_));
 sg13g2_buf_1 _1488_ (.A(_0612_),
    .X(_0613_));
 sg13g2_nor4_1 _1489_ (.A(net42),
    .B(_0592_),
    .C(_0608_),
    .D(net44),
    .Y(_0614_));
 sg13g2_nand2_2 _1490_ (.Y(_0615_),
    .A(_0443_),
    .B(_0444_));
 sg13g2_xnor2_1 _1491_ (.Y(_0616_),
    .A(_0386_),
    .B(_0611_));
 sg13g2_buf_1 _1492_ (.A(_0616_),
    .X(_0617_));
 sg13g2_nand4_1 _1493_ (.B(_0598_),
    .C(net41),
    .A(_0615_),
    .Y(_0618_),
    .D(net43));
 sg13g2_nor2b_1 _1494_ (.A(_0614_),
    .B_N(_0618_),
    .Y(_0619_));
 sg13g2_nand2_2 _1495_ (.Y(_0620_),
    .A(_0600_),
    .B(_0619_));
 sg13g2_inv_1 _1496_ (.Y(_0621_),
    .A(_0620_));
 sg13g2_buf_1 _1497_ (.A(_0621_),
    .X(net9));
 sg13g2_nand2_1 _1498_ (.Y(_0622_),
    .A(_0593_),
    .B(_0596_));
 sg13g2_nand2_1 _1499_ (.Y(_0623_),
    .A(_0615_),
    .B(net41));
 sg13g2_nor2_1 _1500_ (.A(net41),
    .B(_0592_),
    .Y(_0624_));
 sg13g2_a21oi_1 _1501_ (.A1(_0597_),
    .A2(_0623_),
    .Y(_0625_),
    .B1(_0624_));
 sg13g2_a21oi_1 _1502_ (.A1(_0615_),
    .A2(net41),
    .Y(_0626_),
    .B1(_0622_));
 sg13g2_a21o_1 _1503_ (.A2(_0625_),
    .A1(_0622_),
    .B1(_0626_),
    .X(_0627_));
 sg13g2_buf_1 _1504_ (.A(_0627_),
    .X(_0628_));
 sg13g2_inv_1 _1505_ (.Y(_0629_),
    .A(_0628_));
 sg13g2_buf_1 _1506_ (.A(_0629_),
    .X(net10));
 sg13g2_a21oi_1 _1507_ (.A1(_0603_),
    .A2(_0605_),
    .Y(_0630_),
    .B1(_0606_));
 sg13g2_buf_1 _1508_ (.A(\counter[3] ),
    .X(_0631_));
 sg13g2_nor3_1 _1509_ (.A(_0464_),
    .B(_0452_),
    .C(_0465_),
    .Y(_0632_));
 sg13g2_a21oi_1 _1510_ (.A1(_0631_),
    .A2(net83),
    .Y(_0633_),
    .B1(_0632_));
 sg13g2_xnor2_1 _1511_ (.Y(_0634_),
    .A(_0449_),
    .B(_0633_));
 sg13g2_nand2_1 _1512_ (.Y(_0635_),
    .A(net84),
    .B(_0634_));
 sg13g2_xnor2_1 _1513_ (.Y(_0636_),
    .A(_0397_),
    .B(_0635_));
 sg13g2_nand3_1 _1514_ (.B(net42),
    .C(_0636_),
    .A(_0537_),
    .Y(_0637_));
 sg13g2_nand2_1 _1515_ (.Y(_0638_),
    .A(_0630_),
    .B(_0637_));
 sg13g2_nor2_1 _1516_ (.A(_0608_),
    .B(net44),
    .Y(_0639_));
 sg13g2_xnor2_1 _1517_ (.Y(_0640_),
    .A(_0408_),
    .B(_0635_));
 sg13g2_nand2_1 _1518_ (.Y(_0641_),
    .A(_0616_),
    .B(_0640_));
 sg13g2_nor2_1 _1519_ (.A(net42),
    .B(_0641_),
    .Y(_0642_));
 sg13g2_nor3_1 _1520_ (.A(_0589_),
    .B(_0639_),
    .C(_0642_),
    .Y(_0643_));
 sg13g2_a21o_1 _1521_ (.A2(net42),
    .A1(_0615_),
    .B1(_0597_),
    .X(_0644_));
 sg13g2_nand2_1 _1522_ (.Y(_0645_),
    .A(_0536_),
    .B(_0616_));
 sg13g2_nand3b_1 _1523_ (.B(_0589_),
    .C(_0645_),
    .Y(_0646_),
    .A_N(net42));
 sg13g2_o21ai_1 _1524_ (.B1(_0536_),
    .Y(_0647_),
    .A1(net42),
    .A2(_0592_));
 sg13g2_a22oi_1 _1525_ (.Y(_0648_),
    .B1(_0646_),
    .B2(_0647_),
    .A2(_0644_),
    .A1(net44));
 sg13g2_nor2_1 _1526_ (.A(net43),
    .B(_0640_),
    .Y(_0649_));
 sg13g2_a21oi_1 _1527_ (.A1(net42),
    .A2(_0641_),
    .Y(_0650_),
    .B1(_0649_));
 sg13g2_a21oi_1 _1528_ (.A1(_0593_),
    .A2(_0596_),
    .Y(_0651_),
    .B1(_0636_));
 sg13g2_or4_1 _1529_ (.A(net42),
    .B(_0592_),
    .C(_0645_),
    .D(_0651_),
    .X(_0652_));
 sg13g2_o21ai_1 _1530_ (.B1(_0652_),
    .Y(_0653_),
    .A1(_0630_),
    .A2(_0650_));
 sg13g2_a221oi_1 _1531_ (.B2(_0622_),
    .C1(_0653_),
    .B1(_0648_),
    .A1(_0638_),
    .Y(_0654_),
    .A2(_0643_));
 sg13g2_buf_2 _1532_ (.A(_0654_),
    .X(_0655_));
 sg13g2_inv_1 _1533_ (.Y(_0656_),
    .A(_0655_));
 sg13g2_buf_1 _1534_ (.A(_0656_),
    .X(net8));
 sg13g2_o21ai_1 _1535_ (.B1(_0445_),
    .Y(_0657_),
    .A1(_0547_),
    .A2(_0589_));
 sg13g2_or3_1 _1536_ (.A(_0598_),
    .B(_0614_),
    .C(_0657_),
    .X(_0658_));
 sg13g2_nand3_1 _1537_ (.B(net41),
    .C(net43),
    .A(_0615_),
    .Y(_0659_));
 sg13g2_nand3b_1 _1538_ (.B(_0659_),
    .C(_0598_),
    .Y(_0660_),
    .A_N(_0624_));
 sg13g2_a21oi_1 _1539_ (.A1(_0443_),
    .A2(_0309_),
    .Y(_0661_),
    .B1(_0545_));
 sg13g2_nand2_1 _1540_ (.Y(_0662_),
    .A(_0542_),
    .B(_0544_));
 sg13g2_a221oi_1 _1541_ (.B2(_0598_),
    .C1(_0608_),
    .B1(_0589_),
    .A1(_0661_),
    .Y(_0663_),
    .A2(_0662_));
 sg13g2_nand3_1 _1542_ (.B(_0593_),
    .C(_0596_),
    .A(_0536_),
    .Y(_0664_));
 sg13g2_o21ai_1 _1543_ (.B1(_0597_),
    .Y(_0665_),
    .A1(_0448_),
    .A2(_0532_));
 sg13g2_and4_1 _1544_ (.A(_0615_),
    .B(_0546_),
    .C(_0664_),
    .D(_0665_),
    .X(_0666_));
 sg13g2_nor2_1 _1545_ (.A(_0445_),
    .B(_0608_),
    .Y(_0667_));
 sg13g2_nor3_1 _1546_ (.A(_0663_),
    .B(_0666_),
    .C(_0667_),
    .Y(_0668_));
 sg13g2_buf_1 _1547_ (.A(_0668_),
    .X(_0669_));
 sg13g2_a21oi_1 _1548_ (.A1(_0658_),
    .A2(_0660_),
    .Y(_0670_),
    .B1(net39));
 sg13g2_inv_2 _1549_ (.Y(_0671_),
    .A(_0466_));
 sg13g2_nor2_1 _1550_ (.A(_0464_),
    .B(_0465_),
    .Y(_0672_));
 sg13g2_xnor2_1 _1551_ (.Y(_0673_),
    .A(_0631_),
    .B(_0672_));
 sg13g2_nor2_1 _1552_ (.A(net85),
    .B(_0673_),
    .Y(_0674_));
 sg13g2_xnor2_1 _1553_ (.Y(_0675_),
    .A(_0671_),
    .B(_0674_));
 sg13g2_a21oi_1 _1554_ (.A1(_0636_),
    .A2(_0675_),
    .Y(_0676_),
    .B1(net44));
 sg13g2_or3_1 _1555_ (.A(_0663_),
    .B(_0666_),
    .C(_0667_),
    .X(_0677_));
 sg13g2_buf_1 _1556_ (.A(_0677_),
    .X(_0678_));
 sg13g2_nor2_1 _1557_ (.A(_0640_),
    .B(_0678_),
    .Y(_0679_));
 sg13g2_nand3b_1 _1558_ (.B(_0589_),
    .C(_0608_),
    .Y(_0680_),
    .A_N(_0548_));
 sg13g2_nand3_1 _1559_ (.B(_0537_),
    .C(_0548_),
    .A(_0615_),
    .Y(_0681_));
 sg13g2_a21oi_1 _1560_ (.A1(_0680_),
    .A2(_0681_),
    .Y(_0682_),
    .B1(_0613_));
 sg13g2_xnor2_1 _1561_ (.Y(_0683_),
    .A(_0598_),
    .B(_0617_));
 sg13g2_nor4_1 _1562_ (.A(_0537_),
    .B(net41),
    .C(_0592_),
    .D(_0617_),
    .Y(_0684_));
 sg13g2_a21o_1 _1563_ (.A2(_0683_),
    .A1(_0657_),
    .B1(_0684_),
    .X(_0685_));
 sg13g2_nor2_2 _1564_ (.A(_0682_),
    .B(_0685_),
    .Y(_0686_));
 sg13g2_a21oi_1 _1565_ (.A1(_0636_),
    .A2(_0675_),
    .Y(_0687_),
    .B1(net43));
 sg13g2_and4_1 _1566_ (.A(_0658_),
    .B(_0660_),
    .C(net39),
    .D(_0687_),
    .X(_0688_));
 sg13g2_a221oi_1 _1567_ (.B2(_0686_),
    .C1(_0688_),
    .B1(_0679_),
    .A1(_0670_),
    .Y(_0689_),
    .A2(_0676_));
 sg13g2_buf_2 _1568_ (.A(_0689_),
    .X(_0690_));
 sg13g2_or3_1 _1569_ (.A(_0668_),
    .B(_0682_),
    .C(_0685_),
    .X(_0691_));
 sg13g2_nor2_2 _1570_ (.A(_0636_),
    .B(_0675_),
    .Y(_0692_));
 sg13g2_nand4_1 _1571_ (.B(_0600_),
    .C(_0619_),
    .A(net43),
    .Y(_0693_),
    .D(_0692_));
 sg13g2_nand3_1 _1572_ (.B(_0692_),
    .C(_0678_),
    .A(net44),
    .Y(_0694_));
 sg13g2_and4_1 _1573_ (.A(_0655_),
    .B(_0691_),
    .C(_0693_),
    .D(_0694_),
    .X(_0695_));
 sg13g2_buf_2 _1574_ (.A(_0695_),
    .X(_0696_));
 sg13g2_a21oi_2 _1575_ (.B1(_0696_),
    .Y(_0697_),
    .A2(_0690_),
    .A1(_0656_));
 sg13g2_inv_4 _1576_ (.A(_0697_),
    .Y(_0698_));
 sg13g2_buf_1 _1577_ (.A(_0698_),
    .X(net7));
 sg13g2_buf_2 _1578_ (.A(\hvsync_gen.vpos[0] ),
    .X(_0699_));
 sg13g2_buf_2 _1579_ (.A(rst_n),
    .X(_0700_));
 sg13g2_buf_1 _1580_ (.A(_0456_),
    .X(_0701_));
 sg13g2_and2_1 _1581_ (.A(_0458_),
    .B(_0457_),
    .X(_0702_));
 sg13g2_nand3_1 _1582_ (.B(net83),
    .C(_0702_),
    .A(net63),
    .Y(_0703_));
 sg13g2_nor2_2 _1583_ (.A(_0408_),
    .B(_0703_),
    .Y(_0704_));
 sg13g2_nor2_1 _1584_ (.A(_0309_),
    .B(_0522_),
    .Y(_0705_));
 sg13g2_nand4_1 _1585_ (.B(net58),
    .C(_0704_),
    .A(_0386_),
    .Y(_0706_),
    .D(_0705_));
 sg13g2_buf_1 _1586_ (.A(_0706_),
    .X(_0707_));
 sg13g2_and2_1 _1587_ (.A(_0700_),
    .B(_0707_),
    .X(_0708_));
 sg13g2_buf_2 _1588_ (.A(_0708_),
    .X(_0709_));
 sg13g2_inv_1 _1589_ (.Y(_0710_),
    .A(_0699_));
 sg13g2_or2_1 _1590_ (.X(_0711_),
    .B(_0123_),
    .A(_0112_));
 sg13g2_buf_1 _1591_ (.A(_0711_),
    .X(_0712_));
 sg13g2_nor2_1 _1592_ (.A(_0145_),
    .B(_0712_),
    .Y(_0713_));
 sg13g2_inv_1 _1593_ (.Y(_0714_),
    .A(net90));
 sg13g2_nor4_1 _1594_ (.A(_0101_),
    .B(_0714_),
    .C(_0222_),
    .D(net87),
    .Y(_0715_));
 sg13g2_inv_1 _1595_ (.Y(_0716_),
    .A(net78));
 sg13g2_buf_1 _1596_ (.A(_0716_),
    .X(_0717_));
 sg13g2_nor2_1 _1597_ (.A(net54),
    .B(_0255_),
    .Y(_0718_));
 sg13g2_nand4_1 _1598_ (.B(_0713_),
    .C(_0715_),
    .A(_0710_),
    .Y(_0719_),
    .D(_0718_));
 sg13g2_nand2_1 _1599_ (.Y(_0720_),
    .A(_0700_),
    .B(_0719_));
 sg13g2_nor2_1 _1600_ (.A(_0707_),
    .B(net50),
    .Y(_0721_));
 sg13g2_buf_1 _1601_ (.A(_0721_),
    .X(_0722_));
 sg13g2_a22oi_1 _1602_ (.Y(_0723_),
    .B1(net48),
    .B2(_0018_),
    .A2(_0709_),
    .A1(_0699_));
 sg13g2_inv_1 _1603_ (.Y(_0039_),
    .A(_0723_));
 sg13g2_inv_1 _1604_ (.Y(_0724_),
    .A(_0189_));
 sg13g2_a21oi_1 _1605_ (.A1(_0710_),
    .A2(net48),
    .Y(_0725_),
    .B1(_0709_));
 sg13g2_nand3_1 _1606_ (.B(_0699_),
    .C(_0722_),
    .A(net62),
    .Y(_0726_));
 sg13g2_o21ai_1 _1607_ (.B1(_0726_),
    .Y(_0040_),
    .A1(net62),
    .A2(_0725_));
 sg13g2_nand4_1 _1608_ (.B(net59),
    .C(_0699_),
    .A(net87),
    .Y(_0727_),
    .D(_0700_));
 sg13g2_a21oi_1 _1609_ (.A1(net87),
    .A2(_0699_),
    .Y(_0728_),
    .B1(net50));
 sg13g2_buf_1 _1610_ (.A(_0244_),
    .X(_0729_));
 sg13g2_o21ai_1 _1611_ (.B1(net61),
    .Y(_0730_),
    .A1(_0709_),
    .A2(_0728_));
 sg13g2_o21ai_1 _1612_ (.B1(_0730_),
    .Y(_0041_),
    .A1(_0707_),
    .A2(_0727_));
 sg13g2_buf_1 _1613_ (.A(_0178_),
    .X(_0731_));
 sg13g2_nor3_1 _1614_ (.A(net62),
    .B(net59),
    .C(_0018_),
    .Y(_0732_));
 sg13g2_nand2_1 _1615_ (.Y(_0733_),
    .A(_0722_),
    .B(_0732_));
 sg13g2_nor2_1 _1616_ (.A(net50),
    .B(_0732_),
    .Y(_0734_));
 sg13g2_o21ai_1 _1617_ (.B1(net56),
    .Y(_0735_),
    .A1(_0709_),
    .A2(_0734_));
 sg13g2_o21ai_1 _1618_ (.B1(_0735_),
    .Y(_0042_),
    .A1(net56),
    .A2(_0733_));
 sg13g2_nor3_1 _1619_ (.A(net59),
    .B(_0710_),
    .C(_0200_),
    .Y(_0736_));
 sg13g2_nand2_2 _1620_ (.Y(_0737_),
    .A(_0700_),
    .B(_0707_));
 sg13g2_o21ai_1 _1621_ (.B1(_0737_),
    .Y(_0738_),
    .A1(net50),
    .A2(_0736_));
 sg13g2_and2_1 _1622_ (.A(_0233_),
    .B(_0736_),
    .X(_0739_));
 sg13g2_a22oi_1 _1623_ (.Y(_0740_),
    .B1(_0739_),
    .B2(net48),
    .A2(_0738_),
    .A1(_0222_));
 sg13g2_inv_1 _1624_ (.Y(_0043_),
    .A(_0740_));
 sg13g2_and2_1 _1625_ (.A(_0211_),
    .B(_0167_),
    .X(_0741_));
 sg13g2_and4_1 _1626_ (.A(net87),
    .B(net61),
    .C(_0699_),
    .D(_0741_),
    .X(_0742_));
 sg13g2_buf_1 _1627_ (.A(_0742_),
    .X(_0743_));
 sg13g2_nand2_1 _1628_ (.Y(_0744_),
    .A(net48),
    .B(_0743_));
 sg13g2_nor2_1 _1629_ (.A(net50),
    .B(_0743_),
    .Y(_0745_));
 sg13g2_o21ai_1 _1630_ (.B1(net88),
    .Y(_0746_),
    .A1(_0709_),
    .A2(_0745_));
 sg13g2_o21ai_1 _1631_ (.B1(_0746_),
    .Y(_0044_),
    .A1(net88),
    .A2(_0744_));
 sg13g2_nand3_1 _1632_ (.B(net48),
    .C(_0743_),
    .A(net88),
    .Y(_0747_));
 sg13g2_a21oi_1 _1633_ (.A1(net88),
    .A2(_0743_),
    .Y(_0748_),
    .B1(net50));
 sg13g2_o21ai_1 _1634_ (.B1(net79),
    .Y(_0749_),
    .A1(_0709_),
    .A2(_0748_));
 sg13g2_o21ai_1 _1635_ (.B1(_0749_),
    .Y(_0045_),
    .A1(net79),
    .A2(_0747_));
 sg13g2_and4_1 _1636_ (.A(_0134_),
    .B(net88),
    .C(_0732_),
    .D(_0741_),
    .X(_0750_));
 sg13g2_o21ai_1 _1637_ (.B1(_0737_),
    .Y(_0751_),
    .A1(net50),
    .A2(_0750_));
 sg13g2_inv_1 _1638_ (.Y(_0752_),
    .A(net89));
 sg13g2_and2_1 _1639_ (.A(_0752_),
    .B(_0750_),
    .X(_0753_));
 sg13g2_a22oi_1 _1640_ (.Y(_0754_),
    .B1(_0753_),
    .B2(net48),
    .A2(_0751_),
    .A1(_0112_));
 sg13g2_inv_1 _1641_ (.Y(_0046_),
    .A(_0754_));
 sg13g2_and2_1 _1642_ (.A(net89),
    .B(_0123_),
    .X(_0755_));
 sg13g2_and3_1 _1643_ (.X(_0756_),
    .A(net88),
    .B(_0743_),
    .C(_0755_));
 sg13g2_nand2_1 _1644_ (.Y(_0757_),
    .A(net48),
    .B(_0756_));
 sg13g2_o21ai_1 _1645_ (.B1(_0737_),
    .Y(_0758_),
    .A1(net50),
    .A2(_0756_));
 sg13g2_nand2_1 _1646_ (.Y(_0759_),
    .A(_0101_),
    .B(_0758_));
 sg13g2_o21ai_1 _1647_ (.B1(_0759_),
    .Y(_0047_),
    .A1(net80),
    .A2(_0757_));
 sg13g2_nor2b_1 _1648_ (.A(_0156_),
    .B_N(_0743_),
    .Y(_0760_));
 sg13g2_nand2_1 _1649_ (.Y(_0761_),
    .A(net48),
    .B(_0760_));
 sg13g2_nor3_1 _1650_ (.A(_0707_),
    .B(_0720_),
    .C(_0760_),
    .Y(_0762_));
 sg13g2_o21ai_1 _1651_ (.B1(_0079_),
    .Y(_0763_),
    .A1(_0709_),
    .A2(_0762_));
 sg13g2_o21ai_1 _1652_ (.B1(_0763_),
    .Y(_0048_),
    .A1(net90),
    .A2(_0761_));
 sg13g2_and2_1 _1653_ (.A(_0017_),
    .B(_0709_),
    .X(_0029_));
 sg13g2_xnor2_1 _1654_ (.Y(_0764_),
    .A(_0458_),
    .B(_0457_));
 sg13g2_nor2_1 _1655_ (.A(_0737_),
    .B(_0764_),
    .Y(_0030_));
 sg13g2_inv_1 _1656_ (.Y(_0765_),
    .A(_0700_));
 sg13g2_buf_1 _1657_ (.A(_0765_),
    .X(_0766_));
 sg13g2_xnor2_1 _1658_ (.Y(_0767_),
    .A(net63),
    .B(_0702_));
 sg13g2_nor2_1 _1659_ (.A(net60),
    .B(_0767_),
    .Y(_0031_));
 sg13g2_nand2_1 _1660_ (.Y(_0768_),
    .A(net63),
    .B(_0702_));
 sg13g2_xnor2_1 _1661_ (.Y(_0769_),
    .A(_0671_),
    .B(_0768_));
 sg13g2_nor2_1 _1662_ (.A(net60),
    .B(_0769_),
    .Y(_0032_));
 sg13g2_xnor2_1 _1663_ (.Y(_0770_),
    .A(_0408_),
    .B(_0703_));
 sg13g2_nor2_1 _1664_ (.A(net60),
    .B(_0770_),
    .Y(_0033_));
 sg13g2_xnor2_1 _1665_ (.Y(_0771_),
    .A(net73),
    .B(_0704_));
 sg13g2_nor2_1 _1666_ (.A(_0737_),
    .B(_0771_),
    .Y(_0034_));
 sg13g2_nand2_1 _1667_ (.Y(_0772_),
    .A(net73),
    .B(_0704_));
 sg13g2_xnor2_1 _1668_ (.Y(_0773_),
    .A(_0364_),
    .B(_0772_));
 sg13g2_nor2_1 _1669_ (.A(_0766_),
    .B(_0773_),
    .Y(_0035_));
 sg13g2_nand3_1 _1670_ (.B(net73),
    .C(_0704_),
    .A(net75),
    .Y(_0774_));
 sg13g2_xor2_1 _1671_ (.B(_0774_),
    .A(net76),
    .X(_0775_));
 sg13g2_nor2_1 _1672_ (.A(_0766_),
    .B(_0775_),
    .Y(_0036_));
 sg13g2_nand2_1 _1673_ (.Y(_0776_),
    .A(_0439_),
    .B(_0704_));
 sg13g2_xnor2_1 _1674_ (.Y(_0777_),
    .A(_0447_),
    .B(_0776_));
 sg13g2_nor2_1 _1675_ (.A(_0737_),
    .B(_0777_),
    .Y(_0037_));
 sg13g2_nand3_1 _1676_ (.B(net75),
    .C(net58),
    .A(net76),
    .Y(_0778_));
 sg13g2_nor2_1 _1677_ (.A(_0772_),
    .B(_0778_),
    .Y(_0779_));
 sg13g2_xnor2_1 _1678_ (.Y(_0780_),
    .A(_0298_),
    .B(_0779_));
 sg13g2_nor2_1 _1679_ (.A(_0737_),
    .B(_0780_),
    .Y(_0038_));
 sg13g2_buf_2 _1680_ (.A(_0009_),
    .X(_0781_));
 sg13g2_and4_1 _1681_ (.A(net64),
    .B(net65),
    .C(net68),
    .D(net72),
    .X(_0782_));
 sg13g2_nand2_1 _1682_ (.Y(_0783_),
    .A(net70),
    .B(net69));
 sg13g2_o21ai_1 _1683_ (.B1(_0007_),
    .Y(_0784_),
    .A1(net71),
    .A2(_0783_));
 sg13g2_nand4_1 _1684_ (.B(net57),
    .C(_0782_),
    .A(net66),
    .Y(_0785_),
    .D(_0784_));
 sg13g2_buf_1 _1685_ (.A(_0785_),
    .X(_0786_));
 sg13g2_nor2_1 _1686_ (.A(_0781_),
    .B(net53),
    .Y(_0787_));
 sg13g2_nand2b_1 _1687_ (.Y(_0788_),
    .B(_0783_),
    .A_N(net71));
 sg13g2_nand3_1 _1688_ (.B(_0782_),
    .C(_0788_),
    .A(net66),
    .Y(_0789_));
 sg13g2_buf_1 _1689_ (.A(_0789_),
    .X(_0790_));
 sg13g2_buf_1 _1690_ (.A(_0481_),
    .X(_0791_));
 sg13g2_nand2_1 _1691_ (.Y(_0792_),
    .A(net55),
    .B(net57));
 sg13g2_nor3_1 _1692_ (.A(_0787_),
    .B(net52),
    .C(_0792_),
    .Y(_0793_));
 sg13g2_nand2_1 _1693_ (.Y(_0794_),
    .A(_0010_),
    .B(_0793_));
 sg13g2_o21ai_1 _1694_ (.B1(_0794_),
    .Y(_0795_),
    .A1(net69),
    .A2(_0793_));
 sg13g2_and2_1 _1695_ (.A(_0700_),
    .B(_0795_),
    .X(_0019_));
 sg13g2_xnor2_1 _1696_ (.Y(_0796_),
    .A(net70),
    .B(net69));
 sg13g2_nor2_1 _1697_ (.A(net60),
    .B(_0796_),
    .Y(_0020_));
 sg13g2_nand3_1 _1698_ (.B(net69),
    .C(net71),
    .A(net70),
    .Y(_0797_));
 sg13g2_a21oi_1 _1699_ (.A1(_0788_),
    .A2(_0797_),
    .Y(_0021_),
    .B1(net60));
 sg13g2_xnor2_1 _1700_ (.Y(_0798_),
    .A(net64),
    .B(_0784_));
 sg13g2_nor2_1 _1701_ (.A(net60),
    .B(_0798_),
    .Y(_0022_));
 sg13g2_nand2_1 _1702_ (.Y(_0799_),
    .A(net64),
    .B(_0788_));
 sg13g2_xor2_1 _1703_ (.B(_0799_),
    .A(net72),
    .X(_0800_));
 sg13g2_nor2_1 _1704_ (.A(net60),
    .B(_0800_),
    .Y(_0023_));
 sg13g2_nand3_1 _1705_ (.B(net72),
    .C(_0784_),
    .A(net64),
    .Y(_0801_));
 sg13g2_xor2_1 _1706_ (.B(_0801_),
    .A(net68),
    .X(_0802_));
 sg13g2_nor2_1 _1707_ (.A(net60),
    .B(_0802_),
    .Y(_0024_));
 sg13g2_nand4_1 _1708_ (.B(net68),
    .C(net72),
    .A(net64),
    .Y(_0803_),
    .D(_0788_));
 sg13g2_xnor2_1 _1709_ (.Y(_0804_),
    .A(net65),
    .B(_0803_));
 sg13g2_and2_1 _1710_ (.A(_0700_),
    .B(_0804_),
    .X(_0025_));
 sg13g2_xnor2_1 _1711_ (.Y(_0805_),
    .A(net53),
    .B(net52));
 sg13g2_inv_1 _1712_ (.Y(_0806_),
    .A(net52));
 sg13g2_nor3_1 _1713_ (.A(net55),
    .B(net53),
    .C(_0806_),
    .Y(_0807_));
 sg13g2_a21oi_1 _1714_ (.A1(net55),
    .A2(_0805_),
    .Y(_0808_),
    .B1(_0807_));
 sg13g2_inv_2 _1715_ (.Y(_0809_),
    .A(_0781_));
 sg13g2_nand2_1 _1716_ (.Y(_0810_),
    .A(_0782_),
    .B(_0784_));
 sg13g2_xnor2_1 _1717_ (.Y(_0811_),
    .A(_0008_),
    .B(_0810_));
 sg13g2_o21ai_1 _1718_ (.B1(_0811_),
    .Y(_0812_),
    .A1(_0809_),
    .A2(net52));
 sg13g2_nand2b_1 _1719_ (.Y(_0813_),
    .B(net53),
    .A_N(net55));
 sg13g2_nand3_1 _1720_ (.B(_0812_),
    .C(_0813_),
    .A(_0792_),
    .Y(_0814_));
 sg13g2_o21ai_1 _1721_ (.B1(_0814_),
    .Y(_0815_),
    .A1(_0781_),
    .A2(_0808_));
 sg13g2_nand3_1 _1722_ (.B(_0781_),
    .C(net53),
    .A(_0791_),
    .Y(_0816_));
 sg13g2_nand2b_1 _1723_ (.Y(_0817_),
    .B(_0816_),
    .A_N(_0811_));
 sg13g2_nand2_1 _1724_ (.Y(_0818_),
    .A(_0811_),
    .B(_0815_));
 sg13g2_o21ai_1 _1725_ (.B1(_0818_),
    .Y(_0819_),
    .A1(_0815_),
    .A2(_0817_));
 sg13g2_and2_1 _1726_ (.A(_0700_),
    .B(_0819_),
    .X(_0026_));
 sg13g2_nor3_1 _1727_ (.A(net57),
    .B(_0781_),
    .C(net52),
    .Y(_0820_));
 sg13g2_nor2_1 _1728_ (.A(_0809_),
    .B(_0806_),
    .Y(_0821_));
 sg13g2_a21o_1 _1729_ (.A2(net52),
    .A1(_0786_),
    .B1(_0781_),
    .X(_0822_));
 sg13g2_nor3_1 _1730_ (.A(_0786_),
    .B(net52),
    .C(_0811_),
    .Y(_0823_));
 sg13g2_or2_1 _1731_ (.X(_0824_),
    .B(_0823_),
    .A(_0781_));
 sg13g2_a22oi_1 _1732_ (.Y(_0825_),
    .B1(_0824_),
    .B2(net57),
    .A2(_0822_),
    .A1(_0811_));
 sg13g2_nor2_1 _1733_ (.A(_0781_),
    .B(_0790_),
    .Y(_0826_));
 sg13g2_nor2b_1 _1734_ (.A(net53),
    .B_N(_0811_),
    .Y(_0827_));
 sg13g2_nor3_1 _1735_ (.A(net55),
    .B(_0826_),
    .C(_0827_),
    .Y(_0828_));
 sg13g2_a21oi_1 _1736_ (.A1(net55),
    .A2(_0825_),
    .Y(_0829_),
    .B1(_0828_));
 sg13g2_nor4_1 _1737_ (.A(_0765_),
    .B(_0820_),
    .C(_0821_),
    .D(_0829_),
    .Y(_0027_));
 sg13g2_nor2_1 _1738_ (.A(net57),
    .B(net52),
    .Y(_0830_));
 sg13g2_xnor2_1 _1739_ (.Y(_0831_),
    .A(_0809_),
    .B(_0830_));
 sg13g2_and3_1 _1740_ (.X(_0832_),
    .A(net55),
    .B(net53),
    .C(_0831_));
 sg13g2_nor2_1 _1741_ (.A(_0826_),
    .B(_0821_),
    .Y(_0833_));
 sg13g2_nor3_1 _1742_ (.A(net55),
    .B(net53),
    .C(_0833_),
    .Y(_0834_));
 sg13g2_o21ai_1 _1743_ (.B1(_0811_),
    .Y(_0835_),
    .A1(_0832_),
    .A2(_0834_));
 sg13g2_nand4_1 _1744_ (.B(net57),
    .C(_0809_),
    .A(_0791_),
    .Y(_0836_),
    .D(_0823_));
 sg13g2_a21oi_1 _1745_ (.A1(_0835_),
    .A2(_0836_),
    .Y(_0028_),
    .B1(_0765_));
 sg13g2_inv_2 _1746_ (.Y(_0837_),
    .A(_0123_));
 sg13g2_nor2_2 _1747_ (.A(_0244_),
    .B(_0004_),
    .Y(_0838_));
 sg13g2_buf_2 _1748_ (.A(_0003_),
    .X(_0839_));
 sg13g2_and2_1 _1749_ (.A(_0167_),
    .B(_0839_),
    .X(_0840_));
 sg13g2_buf_2 _1750_ (.A(_0840_),
    .X(_0841_));
 sg13g2_and2_1 _1751_ (.A(_0838_),
    .B(_0841_),
    .X(_0842_));
 sg13g2_nor3_1 _1752_ (.A(net80),
    .B(net90),
    .C(net77),
    .Y(_0843_));
 sg13g2_nand4_1 _1753_ (.B(_0837_),
    .C(_0842_),
    .A(_0752_),
    .Y(_0844_),
    .D(_0843_));
 sg13g2_nand2_1 _1754_ (.Y(_0845_),
    .A(_0838_),
    .B(_0841_));
 sg13g2_buf_1 _1755_ (.A(_0002_),
    .X(_0846_));
 sg13g2_nor2_1 _1756_ (.A(net82),
    .B(_0712_),
    .Y(_0847_));
 sg13g2_a21oi_1 _1757_ (.A1(net82),
    .A2(_0755_),
    .Y(_0848_),
    .B1(_0847_));
 sg13g2_nand2_2 _1758_ (.Y(_0849_),
    .A(\hvsync_gen.vpos[7] ),
    .B(_0123_));
 sg13g2_nor2_2 _1759_ (.A(_0090_),
    .B(\hvsync_gen.vpos[9] ),
    .Y(_0850_));
 sg13g2_a21oi_1 _1760_ (.A1(_0849_),
    .A2(_0850_),
    .Y(_0851_),
    .B1(_0716_));
 sg13g2_xnor2_1 _1761_ (.Y(_0852_),
    .A(net77),
    .B(_0851_));
 sg13g2_nor4_1 _1762_ (.A(\hvsync_gen.vpos[7] ),
    .B(_0211_),
    .C(_0244_),
    .D(_0004_),
    .Y(_0853_));
 sg13g2_nand3_1 _1763_ (.B(_0841_),
    .C(_0853_),
    .A(_0850_),
    .Y(_0854_));
 sg13g2_nor3_2 _1764_ (.A(\hvsync_gen.vpos[5] ),
    .B(_0211_),
    .C(_0167_),
    .Y(_0855_));
 sg13g2_nor2_1 _1765_ (.A(_0837_),
    .B(_0855_),
    .Y(_0856_));
 sg13g2_or2_1 _1766_ (.X(_0857_),
    .B(\hvsync_gen.vpos[9] ),
    .A(_0090_));
 sg13g2_buf_1 _1767_ (.A(_0857_),
    .X(_0858_));
 sg13g2_nor3_1 _1768_ (.A(_0123_),
    .B(_0211_),
    .C(_0858_),
    .Y(_0859_));
 sg13g2_or3_1 _1769_ (.A(\hvsync_gen.vpos[5] ),
    .B(_0211_),
    .C(_0167_),
    .X(_0860_));
 sg13g2_buf_2 _1770_ (.A(_0860_),
    .X(_0861_));
 sg13g2_nor2_1 _1771_ (.A(_0123_),
    .B(_0861_),
    .Y(_0862_));
 sg13g2_a221oi_1 _1772_ (.B2(_0842_),
    .C1(_0862_),
    .B1(_0859_),
    .A1(_0854_),
    .Y(_0863_),
    .A2(_0856_));
 sg13g2_or4_1 _1773_ (.A(_0845_),
    .B(_0848_),
    .C(_0852_),
    .D(_0863_),
    .X(_0864_));
 sg13g2_nor2_2 _1774_ (.A(_0849_),
    .B(_0855_),
    .Y(_0865_));
 sg13g2_nand4_1 _1775_ (.B(net90),
    .C(_0846_),
    .A(net80),
    .Y(_0866_),
    .D(_0865_));
 sg13g2_a21oi_1 _1776_ (.A1(_0755_),
    .A2(_0861_),
    .Y(_0867_),
    .B1(_0846_));
 sg13g2_inv_1 _1777_ (.Y(_0868_),
    .A(_0002_));
 sg13g2_nor4_1 _1778_ (.A(net80),
    .B(_0868_),
    .C(_0849_),
    .D(_0855_),
    .Y(_0869_));
 sg13g2_o21ai_1 _1779_ (.B1(_0714_),
    .Y(_0870_),
    .A1(_0867_),
    .A2(_0869_));
 sg13g2_o21ai_1 _1780_ (.B1(_0850_),
    .Y(_0871_),
    .A1(_0849_),
    .A2(_0855_));
 sg13g2_buf_2 _1781_ (.A(_0871_),
    .X(_0872_));
 sg13g2_nand3_1 _1782_ (.B(_0741_),
    .C(_0838_),
    .A(_0839_),
    .Y(_0873_));
 sg13g2_or2_1 _1783_ (.X(_0874_),
    .B(_0873_),
    .A(_0872_));
 sg13g2_xnor2_1 _1784_ (.Y(_0875_),
    .A(_0211_),
    .B(net78));
 sg13g2_a21oi_1 _1785_ (.A1(_0712_),
    .A2(_0849_),
    .Y(_0876_),
    .B1(_0875_));
 sg13g2_nand2_1 _1786_ (.Y(_0877_),
    .A(_0842_),
    .B(_0876_));
 sg13g2_a221oi_1 _1787_ (.B2(_0874_),
    .C1(_0877_),
    .B1(_0863_),
    .A1(_0866_),
    .Y(_0878_),
    .A2(_0870_));
 sg13g2_nand2_1 _1788_ (.Y(_0879_),
    .A(_0090_),
    .B(_0002_));
 sg13g2_mux2_1 _1789_ (.A0(_0002_),
    .A1(_0879_),
    .S(_0714_),
    .X(_0880_));
 sg13g2_inv_1 _1790_ (.Y(_0881_),
    .A(_0090_));
 sg13g2_nand4_1 _1791_ (.B(net90),
    .C(_0755_),
    .A(_0881_),
    .Y(_0882_),
    .D(_0861_));
 sg13g2_nor2_1 _1792_ (.A(net80),
    .B(_0002_),
    .Y(_0883_));
 sg13g2_o21ai_1 _1793_ (.B1(_0883_),
    .Y(_0884_),
    .A1(_0849_),
    .A2(_0855_));
 sg13g2_and3_1 _1794_ (.X(_0885_),
    .A(_0880_),
    .B(_0882_),
    .C(_0884_));
 sg13g2_buf_1 _1795_ (.A(_0885_),
    .X(_0886_));
 sg13g2_a21oi_1 _1796_ (.A1(_0864_),
    .A2(_0878_),
    .Y(_0887_),
    .B1(_0886_));
 sg13g2_nand2_1 _1797_ (.Y(_0888_),
    .A(net82),
    .B(_0858_));
 sg13g2_mux2_1 _1798_ (.A0(_0888_),
    .A1(net82),
    .S(_0865_),
    .X(_0889_));
 sg13g2_buf_2 _1799_ (.A(_0889_),
    .X(_0890_));
 sg13g2_nand4_1 _1800_ (.B(_0839_),
    .C(_0244_),
    .A(net78),
    .Y(_0891_),
    .D(_0004_));
 sg13g2_nor2_2 _1801_ (.A(net77),
    .B(_0891_),
    .Y(_0892_));
 sg13g2_a21oi_1 _1802_ (.A1(_0850_),
    .A2(_0892_),
    .Y(_0893_),
    .B1(_0856_));
 sg13g2_nor3_1 _1803_ (.A(net77),
    .B(_0850_),
    .C(_0891_),
    .Y(_0894_));
 sg13g2_nor4_1 _1804_ (.A(net89),
    .B(_0837_),
    .C(_0855_),
    .D(_0894_),
    .Y(_0895_));
 sg13g2_a21oi_2 _1805_ (.B1(_0895_),
    .Y(_0896_),
    .A2(_0893_),
    .A1(net89));
 sg13g2_and4_1 _1806_ (.A(_0844_),
    .B(net49),
    .C(_0890_),
    .D(_0896_),
    .X(_0897_));
 sg13g2_buf_1 _1807_ (.A(_0897_),
    .X(_0898_));
 sg13g2_nand2_1 _1808_ (.Y(_0899_),
    .A(_0850_),
    .B(_0841_));
 sg13g2_and2_1 _1809_ (.A(_0244_),
    .B(_0004_),
    .X(_0900_));
 sg13g2_a21oi_1 _1810_ (.A1(net77),
    .A2(_0838_),
    .Y(_0901_),
    .B1(_0900_));
 sg13g2_nor3_1 _1811_ (.A(net89),
    .B(_0899_),
    .C(_0901_),
    .Y(_0902_));
 sg13g2_nor3_1 _1812_ (.A(_0837_),
    .B(_0855_),
    .C(_0902_),
    .Y(_0903_));
 sg13g2_or2_1 _1813_ (.X(_0904_),
    .B(_0901_),
    .A(_0899_));
 sg13g2_a21oi_1 _1814_ (.A1(_0861_),
    .A2(_0904_),
    .Y(_0905_),
    .B1(net79));
 sg13g2_or2_1 _1815_ (.X(_0906_),
    .B(_0905_),
    .A(_0903_));
 sg13g2_nand4_1 _1816_ (.B(_0838_),
    .C(_0841_),
    .A(_0837_),
    .Y(_0907_),
    .D(_0843_));
 sg13g2_a221oi_1 _1817_ (.B2(net82),
    .C1(net89),
    .B1(_0858_),
    .A1(_0123_),
    .Y(_0908_),
    .A2(_0861_));
 sg13g2_a22oi_1 _1818_ (.Y(_0909_),
    .B1(_0907_),
    .B2(_0908_),
    .A2(_0865_),
    .A1(net82));
 sg13g2_nand4_1 _1819_ (.B(_0850_),
    .C(_0841_),
    .A(_0837_),
    .Y(_0910_),
    .D(_0853_));
 sg13g2_nand4_1 _1820_ (.B(_0882_),
    .C(_0884_),
    .A(_0880_),
    .Y(_0911_),
    .D(_0910_));
 sg13g2_nand3_1 _1821_ (.B(_0911_),
    .C(_0892_),
    .A(_0909_),
    .Y(_0912_));
 sg13g2_nand2_1 _1822_ (.Y(_0913_),
    .A(_0909_),
    .B(_0911_));
 sg13g2_inv_1 _1823_ (.Y(_0914_),
    .A(_0892_));
 sg13g2_nor4_1 _1824_ (.A(net51),
    .B(_0914_),
    .C(_0903_),
    .D(_0905_),
    .Y(_0915_));
 sg13g2_a21o_1 _1825_ (.A2(_0912_),
    .A1(_0906_),
    .B1(_0915_),
    .X(_0916_));
 sg13g2_buf_1 _1826_ (.A(_0916_),
    .X(_0917_));
 sg13g2_and2_1 _1827_ (.A(_0898_),
    .B(_0917_),
    .X(_0918_));
 sg13g2_nor2_1 _1828_ (.A(_0886_),
    .B(_0890_),
    .Y(_0919_));
 sg13g2_o21ai_1 _1829_ (.B1(_0911_),
    .Y(_0920_),
    .A1(_0886_),
    .A2(_0896_));
 sg13g2_a22oi_1 _1830_ (.Y(_0921_),
    .B1(_0920_),
    .B2(_0890_),
    .A2(_0896_),
    .A1(_0919_));
 sg13g2_xnor2_1 _1831_ (.Y(_0922_),
    .A(_0752_),
    .B(_0856_));
 sg13g2_nor2_1 _1832_ (.A(net79),
    .B(_0854_),
    .Y(_0923_));
 sg13g2_nor3_1 _1833_ (.A(_0922_),
    .B(_0923_),
    .C(_0919_),
    .Y(_0924_));
 sg13g2_a21o_1 _1834_ (.A2(_0922_),
    .A1(net49),
    .B1(_0924_),
    .X(_0925_));
 sg13g2_buf_1 _1835_ (.A(_0925_),
    .X(_0926_));
 sg13g2_a21oi_1 _1836_ (.A1(_0917_),
    .A2(_0921_),
    .Y(_0927_),
    .B1(_0926_));
 sg13g2_nor2_1 _1837_ (.A(_0918_),
    .B(_0927_),
    .Y(_0928_));
 sg13g2_nor2_2 _1838_ (.A(net77),
    .B(_0178_),
    .Y(_0929_));
 sg13g2_xor2_1 _1839_ (.B(_0929_),
    .A(_0839_),
    .X(_0930_));
 sg13g2_nand2_1 _1840_ (.Y(_0931_),
    .A(_0928_),
    .B(_0930_));
 sg13g2_a21oi_1 _1841_ (.A1(net49),
    .A2(_0922_),
    .Y(_0932_),
    .B1(_0924_));
 sg13g2_o21ai_1 _1842_ (.B1(_0917_),
    .Y(_0933_),
    .A1(_0932_),
    .A2(_0898_));
 sg13g2_a21oi_1 _1843_ (.A1(net82),
    .A2(_0858_),
    .Y(_0934_),
    .B1(net89));
 sg13g2_and4_1 _1844_ (.A(_0868_),
    .B(_0838_),
    .C(_0841_),
    .D(_0843_),
    .X(_0935_));
 sg13g2_o21ai_1 _1845_ (.B1(_0861_),
    .Y(_0936_),
    .A1(net79),
    .A2(_0935_));
 sg13g2_a22oi_1 _1846_ (.Y(_0937_),
    .B1(_0934_),
    .B2(_0936_),
    .A2(_0865_),
    .A1(net82));
 sg13g2_and2_1 _1847_ (.A(net77),
    .B(_0937_),
    .X(_0938_));
 sg13g2_a22oi_1 _1848_ (.Y(_0939_),
    .B1(_0938_),
    .B2(_0887_),
    .A2(_0913_),
    .A1(_0233_));
 sg13g2_o21ai_1 _1849_ (.B1(_0921_),
    .Y(_0940_),
    .A1(_0891_),
    .A2(_0939_));
 sg13g2_mux2_1 _1850_ (.A0(_0933_),
    .A1(_0917_),
    .S(_0940_),
    .X(_0941_));
 sg13g2_xnor2_1 _1851_ (.Y(_0942_),
    .A(_0839_),
    .B(_0929_));
 sg13g2_nand2_1 _1852_ (.Y(_0943_),
    .A(_0837_),
    .B(_0892_));
 sg13g2_nand2_1 _1853_ (.Y(_0944_),
    .A(net79),
    .B(_0892_));
 sg13g2_nand4_1 _1854_ (.B(_0861_),
    .C(_0850_),
    .A(_0849_),
    .Y(_0945_),
    .D(_0873_));
 sg13g2_mux2_1 _1855_ (.A0(_0943_),
    .A1(_0944_),
    .S(_0945_),
    .X(_0946_));
 sg13g2_o21ai_1 _1856_ (.B1(_0922_),
    .Y(_0947_),
    .A1(_0946_),
    .A2(_0890_));
 sg13g2_and2_1 _1857_ (.A(net49),
    .B(_0947_),
    .X(_0948_));
 sg13g2_inv_1 _1858_ (.Y(_0949_),
    .A(_0946_));
 sg13g2_and2_1 _1859_ (.A(_0844_),
    .B(_0890_),
    .X(_0950_));
 sg13g2_inv_1 _1860_ (.Y(_0951_),
    .A(_0950_));
 sg13g2_a21oi_1 _1861_ (.A1(net49),
    .A2(_0949_),
    .Y(_0952_),
    .B1(_0951_));
 sg13g2_o21ai_1 _1862_ (.B1(net79),
    .Y(_0953_),
    .A1(_0855_),
    .A2(_0902_));
 sg13g2_nand3_1 _1863_ (.B(_0861_),
    .C(_0904_),
    .A(_0837_),
    .Y(_0954_));
 sg13g2_nor2_1 _1864_ (.A(_0886_),
    .B(_0891_),
    .Y(_0955_));
 sg13g2_a221oi_1 _1865_ (.B2(_0937_),
    .C1(_0892_),
    .B1(_0955_),
    .A1(_0953_),
    .Y(_0956_),
    .A2(_0954_));
 sg13g2_nor2_1 _1866_ (.A(net51),
    .B(_0946_),
    .Y(_0957_));
 sg13g2_or2_1 _1867_ (.X(_0958_),
    .B(_0957_),
    .A(_0956_));
 sg13g2_nor4_2 _1868_ (.A(_0948_),
    .B(_0952_),
    .C(_0932_),
    .Y(_0959_),
    .D(_0958_));
 sg13g2_nor2_1 _1869_ (.A(_0956_),
    .B(_0957_),
    .Y(_0960_));
 sg13g2_nand4_1 _1870_ (.B(net49),
    .C(_0890_),
    .A(_0844_),
    .Y(_0961_),
    .D(_0896_));
 sg13g2_a21oi_2 _1871_ (.B1(_0961_),
    .Y(_0962_),
    .A2(_0960_),
    .A1(_0926_));
 sg13g2_nor2_2 _1872_ (.A(_0959_),
    .B(_0962_),
    .Y(_0963_));
 sg13g2_nand3b_1 _1873_ (.B(_0942_),
    .C(_0963_),
    .Y(_0964_),
    .A_N(_0941_));
 sg13g2_nand2_1 _1874_ (.Y(_0965_),
    .A(net78),
    .B(_0900_));
 sg13g2_or2_1 _1875_ (.X(_0966_),
    .B(_0004_),
    .A(_0244_));
 sg13g2_o21ai_1 _1876_ (.B1(net78),
    .Y(_0967_),
    .A1(_0966_),
    .A2(_0872_));
 sg13g2_xnor2_1 _1877_ (.Y(_0968_),
    .A(_0233_),
    .B(_0967_));
 sg13g2_or2_1 _1878_ (.X(_0969_),
    .B(_0968_),
    .A(_0965_));
 sg13g2_or3_1 _1879_ (.A(_0969_),
    .B(net51),
    .C(_0898_),
    .X(_0970_));
 sg13g2_nand3_1 _1880_ (.B(net51),
    .C(_0961_),
    .A(_0968_),
    .Y(_0971_));
 sg13g2_a221oi_1 _1881_ (.B2(_0960_),
    .C1(_0952_),
    .B1(_0926_),
    .A1(net49),
    .Y(_0972_),
    .A2(_0947_));
 sg13g2_a21o_1 _1882_ (.A2(_0971_),
    .A1(_0970_),
    .B1(_0972_),
    .X(_0973_));
 sg13g2_nor2b_2 _1883_ (.A(_0969_),
    .B_N(net51),
    .Y(_0974_));
 sg13g2_nor2b_1 _1884_ (.A(net51),
    .B_N(_0968_),
    .Y(_0975_));
 sg13g2_o21ai_1 _1885_ (.B1(_0972_),
    .Y(_0976_),
    .A1(_0974_),
    .A2(_0975_));
 sg13g2_a22oi_1 _1886_ (.Y(_0977_),
    .B1(_0898_),
    .B2(_0974_),
    .A2(_0968_),
    .A1(_0965_));
 sg13g2_nand3_1 _1887_ (.B(_0976_),
    .C(_0977_),
    .A(_0973_),
    .Y(_0978_));
 sg13g2_buf_2 _1888_ (.A(_0978_),
    .X(_0979_));
 sg13g2_a21o_1 _1889_ (.A2(_0964_),
    .A1(_0931_),
    .B1(_0979_),
    .X(_0980_));
 sg13g2_buf_2 _1890_ (.A(_0980_),
    .X(_0981_));
 sg13g2_or2_1 _1891_ (.X(_0982_),
    .B(_0927_),
    .A(_0918_));
 sg13g2_nor2_1 _1892_ (.A(_0926_),
    .B(_0917_),
    .Y(_0983_));
 sg13g2_mux2_1 _1893_ (.A0(_0918_),
    .A1(_0983_),
    .S(_0940_),
    .X(_0984_));
 sg13g2_or3_1 _1894_ (.A(_0959_),
    .B(_0962_),
    .C(_0942_),
    .X(_0985_));
 sg13g2_o21ai_1 _1895_ (.B1(_0942_),
    .Y(_0986_),
    .A1(_0959_),
    .A2(_0962_));
 sg13g2_o21ai_1 _1896_ (.B1(_0986_),
    .Y(_0987_),
    .A1(_0984_),
    .A2(_0985_));
 sg13g2_a22oi_1 _1897_ (.Y(_0988_),
    .B1(_0987_),
    .B2(_0979_),
    .A2(_0942_),
    .A1(_0982_));
 sg13g2_buf_2 _1898_ (.A(_0988_),
    .X(_0989_));
 sg13g2_a21oi_2 _1899_ (.B1(net56),
    .Y(_0990_),
    .A2(_0989_),
    .A1(_0981_));
 sg13g2_nand2_1 _1900_ (.Y(_0991_),
    .A(net87),
    .B(_0990_));
 sg13g2_and2_1 _1901_ (.A(_0981_),
    .B(_0989_),
    .X(_0992_));
 sg13g2_buf_2 _1902_ (.A(_0992_),
    .X(_0993_));
 sg13g2_nand3_1 _1903_ (.B(_0928_),
    .C(_0941_),
    .A(_0963_),
    .Y(_0994_));
 sg13g2_nor2_1 _1904_ (.A(_0716_),
    .B(_0966_),
    .Y(_0995_));
 sg13g2_a21oi_1 _1905_ (.A1(_0984_),
    .A2(_0930_),
    .Y(_0996_),
    .B1(_0995_));
 sg13g2_nand3_1 _1906_ (.B(_0942_),
    .C(_0941_),
    .A(_0982_),
    .Y(_0997_));
 sg13g2_nand4_1 _1907_ (.B(_0994_),
    .C(_0996_),
    .A(_0979_),
    .Y(_0998_),
    .D(_0997_));
 sg13g2_buf_1 _1908_ (.A(_0998_),
    .X(_0999_));
 sg13g2_nand2_1 _1909_ (.Y(_1000_),
    .A(net78),
    .B(_0838_));
 sg13g2_and4_1 _1910_ (.A(_0982_),
    .B(_0930_),
    .C(_0941_),
    .D(_1000_),
    .X(_1001_));
 sg13g2_nor2_1 _1911_ (.A(_0963_),
    .B(_0995_),
    .Y(_1002_));
 sg13g2_nand2_1 _1912_ (.Y(_1003_),
    .A(_0932_),
    .B(_0917_));
 sg13g2_nand2b_1 _1913_ (.Y(_1004_),
    .B(_0926_),
    .A_N(_0917_));
 sg13g2_mux2_1 _1914_ (.A0(_1003_),
    .A1(_1004_),
    .S(_0940_),
    .X(_1005_));
 sg13g2_nor3_1 _1915_ (.A(_0930_),
    .B(_0995_),
    .C(_1005_),
    .Y(_1006_));
 sg13g2_or4_1 _1916_ (.A(_0979_),
    .B(_1001_),
    .C(_1002_),
    .D(_1006_),
    .X(_1007_));
 sg13g2_buf_2 _1917_ (.A(_1007_),
    .X(_1008_));
 sg13g2_a21oi_2 _1918_ (.B1(net54),
    .Y(_1009_),
    .A2(_1008_),
    .A1(_0999_));
 sg13g2_nand3_1 _1919_ (.B(net51),
    .C(_0961_),
    .A(_0875_),
    .Y(_1010_));
 sg13g2_a21o_1 _1920_ (.A2(_1010_),
    .A1(_0970_),
    .B1(_0972_),
    .X(_1011_));
 sg13g2_nor2b_1 _1921_ (.A(net51),
    .B_N(_0875_),
    .Y(_1012_));
 sg13g2_o21ai_1 _1922_ (.B1(_0972_),
    .Y(_1013_),
    .A1(_0974_),
    .A2(_1012_));
 sg13g2_a22oi_1 _1923_ (.Y(_1014_),
    .B1(_0898_),
    .B2(_0974_),
    .A2(_0875_),
    .A1(_0965_));
 sg13g2_nand3_1 _1924_ (.B(_1013_),
    .C(_1014_),
    .A(_1011_),
    .Y(_1015_));
 sg13g2_nor3_1 _1925_ (.A(_0959_),
    .B(_0962_),
    .C(_0995_),
    .Y(_1016_));
 sg13g2_a221oi_1 _1926_ (.B2(_1016_),
    .C1(_1005_),
    .B1(_1015_),
    .A1(_0963_),
    .Y(_1017_),
    .A2(_0942_));
 sg13g2_and4_1 _1927_ (.A(net49),
    .B(_0922_),
    .C(_0949_),
    .D(_0890_),
    .X(_1018_));
 sg13g2_a21o_1 _1928_ (.A2(_1015_),
    .A1(_1001_),
    .B1(_1018_),
    .X(_1019_));
 sg13g2_nand2_1 _1929_ (.Y(_1020_),
    .A(_0984_),
    .B(_0942_));
 sg13g2_a21oi_1 _1930_ (.A1(_1000_),
    .A2(_1015_),
    .Y(_1021_),
    .B1(_1020_));
 sg13g2_nor2_1 _1931_ (.A(_0963_),
    .B(_0930_),
    .Y(_1022_));
 sg13g2_and3_1 _1932_ (.X(_1023_),
    .A(_1022_),
    .B(_1000_),
    .C(_1015_));
 sg13g2_or4_1 _1933_ (.A(_1017_),
    .B(_1019_),
    .C(_1021_),
    .D(_1023_),
    .X(_1024_));
 sg13g2_a21oi_1 _1934_ (.A1(_0993_),
    .A2(_1009_),
    .Y(_1025_),
    .B1(_1024_));
 sg13g2_inv_1 _1935_ (.Y(_1026_),
    .A(_0200_));
 sg13g2_nor4_1 _1936_ (.A(_1017_),
    .B(_1019_),
    .C(_1021_),
    .D(_1023_),
    .Y(_1027_));
 sg13g2_buf_1 _1937_ (.A(_1027_),
    .X(_1028_));
 sg13g2_o21ai_1 _1938_ (.B1(net61),
    .Y(_1029_),
    .A1(_1026_),
    .A2(_1028_));
 sg13g2_a21o_1 _1939_ (.A2(_1025_),
    .A1(_0991_),
    .B1(_1029_),
    .X(_1030_));
 sg13g2_nand2_2 _1940_ (.Y(_1031_),
    .A(_0981_),
    .B(_0989_));
 sg13g2_nand2_1 _1941_ (.Y(_1032_),
    .A(_1031_),
    .B(net38));
 sg13g2_nand2_1 _1942_ (.Y(_1033_),
    .A(net54),
    .B(_0255_));
 sg13g2_nand3_1 _1943_ (.B(_0999_),
    .C(_1008_),
    .A(_0718_),
    .Y(_1034_));
 sg13g2_o21ai_1 _1944_ (.B1(_1034_),
    .Y(_1035_),
    .A1(net38),
    .A2(_1033_));
 sg13g2_nor2_2 _1945_ (.A(net54),
    .B(net61),
    .Y(_1036_));
 sg13g2_nor2_1 _1946_ (.A(net78),
    .B(_0255_),
    .Y(_1037_));
 sg13g2_mux2_1 _1947_ (.A0(_1036_),
    .A1(_1037_),
    .S(_1031_),
    .X(_1038_));
 sg13g2_nand2_1 _1948_ (.Y(_1039_),
    .A(_0999_),
    .B(_1008_));
 sg13g2_a221oi_1 _1949_ (.B2(net36),
    .C1(_1018_),
    .B1(_1038_),
    .A1(_1032_),
    .Y(_1040_),
    .A2(_1035_));
 sg13g2_and4_1 _1950_ (.A(_0979_),
    .B(_0994_),
    .C(_0996_),
    .D(_0997_),
    .X(_1041_));
 sg13g2_buf_2 _1951_ (.A(_1041_),
    .X(_1042_));
 sg13g2_nor4_2 _1952_ (.A(_0979_),
    .B(_1001_),
    .C(_1002_),
    .Y(_1043_),
    .D(_1006_));
 sg13g2_nor2_1 _1953_ (.A(_1042_),
    .B(_1043_),
    .Y(_1044_));
 sg13g2_nor2_1 _1954_ (.A(_0993_),
    .B(_1044_),
    .Y(_1045_));
 sg13g2_nor3_1 _1955_ (.A(net56),
    .B(net62),
    .C(net61),
    .Y(_1046_));
 sg13g2_nor3_2 _1956_ (.A(_0729_),
    .B(_1042_),
    .C(_1043_),
    .Y(_1047_));
 sg13g2_nor2_1 _1957_ (.A(_0717_),
    .B(net87),
    .Y(_1048_));
 sg13g2_a21oi_1 _1958_ (.A1(_0993_),
    .A2(_1048_),
    .Y(_1049_),
    .B1(_0990_));
 sg13g2_a22oi_1 _1959_ (.Y(_1050_),
    .B1(_1047_),
    .B2(_1049_),
    .A2(_1046_),
    .A1(_1045_));
 sg13g2_and3_1 _1960_ (.X(_1051_),
    .A(_1030_),
    .B(_1040_),
    .C(_1050_));
 sg13g2_buf_8 _1961_ (.A(_1051_),
    .X(_1052_));
 sg13g2_a21oi_1 _1962_ (.A1(_0999_),
    .A2(_1008_),
    .Y(_1053_),
    .B1(_0255_));
 sg13g2_xnor2_1 _1963_ (.Y(_1054_),
    .A(net56),
    .B(_1028_));
 sg13g2_nand3_1 _1964_ (.B(_1053_),
    .C(_1054_),
    .A(net87),
    .Y(_1055_));
 sg13g2_nand2_1 _1965_ (.Y(_1056_),
    .A(_0990_),
    .B(_1047_));
 sg13g2_buf_1 _1966_ (.A(_1024_),
    .X(_1057_));
 sg13g2_nand2_1 _1967_ (.Y(_1058_),
    .A(net37),
    .B(_1036_));
 sg13g2_buf_1 _1968_ (.A(_0993_),
    .X(_1059_));
 sg13g2_nor3_1 _1969_ (.A(net54),
    .B(net31),
    .C(net37),
    .Y(_1060_));
 sg13g2_nor2_1 _1970_ (.A(net56),
    .B(_1031_),
    .Y(_1061_));
 sg13g2_o21ai_1 _1971_ (.B1(_0729_),
    .Y(_1062_),
    .A1(_1042_),
    .A2(_1043_));
 sg13g2_nand2_1 _1972_ (.Y(_1063_),
    .A(net62),
    .B(_1062_));
 sg13g2_o21ai_1 _1973_ (.B1(_1063_),
    .Y(_1064_),
    .A1(_1060_),
    .A2(_1061_));
 sg13g2_and4_1 _1974_ (.A(_1055_),
    .B(_1056_),
    .C(_1058_),
    .D(_1064_),
    .X(_1065_));
 sg13g2_buf_1 _1975_ (.A(_1065_),
    .X(_1066_));
 sg13g2_nor2_1 _1976_ (.A(_1052_),
    .B(_1066_),
    .Y(_1067_));
 sg13g2_buf_2 _1977_ (.A(_0005_),
    .X(_1068_));
 sg13g2_inv_4 _1978_ (.A(_1052_),
    .Y(_1069_));
 sg13g2_nor3_1 _1979_ (.A(net56),
    .B(_1042_),
    .C(_1043_),
    .Y(_1070_));
 sg13g2_o21ai_1 _1980_ (.B1(net59),
    .Y(_1071_),
    .A1(net37),
    .A2(_1070_));
 sg13g2_a21oi_1 _1981_ (.A1(net38),
    .A2(_1053_),
    .Y(_1072_),
    .B1(_0993_));
 sg13g2_o21ai_1 _1982_ (.B1(_1036_),
    .Y(_1073_),
    .A1(_1042_),
    .A2(_1043_));
 sg13g2_o21ai_1 _1983_ (.B1(_1037_),
    .Y(_1074_),
    .A1(_1042_),
    .A2(_1043_));
 sg13g2_and3_1 _1984_ (.X(_1075_),
    .A(_1034_),
    .B(_1073_),
    .C(_1074_));
 sg13g2_a22oi_1 _1985_ (.Y(_1076_),
    .B1(_1075_),
    .B2(_1059_),
    .A2(_1072_),
    .A1(_1071_));
 sg13g2_nand2_1 _1986_ (.Y(_1077_),
    .A(_0699_),
    .B(_1076_));
 sg13g2_a21oi_1 _1987_ (.A1(_1068_),
    .A2(_1069_),
    .Y(_1078_),
    .B1(_1077_));
 sg13g2_nor3_1 _1988_ (.A(net54),
    .B(_1031_),
    .C(net36),
    .Y(_1079_));
 sg13g2_mux2_1 _1989_ (.A0(_0990_),
    .A1(_1009_),
    .S(_1057_),
    .X(_1080_));
 sg13g2_o21ai_1 _1990_ (.B1(net62),
    .Y(_1081_),
    .A1(_1079_),
    .A2(_1080_));
 sg13g2_nand3_1 _1991_ (.B(net37),
    .C(_1044_),
    .A(_1026_),
    .Y(_1082_));
 sg13g2_nor2_1 _1992_ (.A(_1068_),
    .B(_1018_),
    .Y(_1083_));
 sg13g2_o21ai_1 _1993_ (.B1(net37),
    .Y(_1084_),
    .A1(net56),
    .A2(_1053_));
 sg13g2_a221oi_1 _1994_ (.B2(net38),
    .C1(_1047_),
    .B1(_0990_),
    .A1(_0718_),
    .Y(_1085_),
    .A2(net31));
 sg13g2_a22oi_1 _1995_ (.Y(_1086_),
    .B1(_1084_),
    .B2(_1085_),
    .A2(_1083_),
    .A1(_1082_));
 sg13g2_nand3b_1 _1996_ (.B(_1081_),
    .C(_1086_),
    .Y(_1087_),
    .A_N(_1076_));
 sg13g2_buf_2 _1997_ (.A(_1087_),
    .X(_1088_));
 sg13g2_nand3_1 _1998_ (.B(net61),
    .C(net37),
    .A(_0731_),
    .Y(_1089_));
 sg13g2_nand3_1 _1999_ (.B(_0999_),
    .C(_1008_),
    .A(net59),
    .Y(_1090_));
 sg13g2_nand4_1 _2000_ (.B(net38),
    .C(_1062_),
    .A(_0990_),
    .Y(_1091_),
    .D(_1090_));
 sg13g2_nand3_1 _2001_ (.B(_1044_),
    .C(_1036_),
    .A(net31),
    .Y(_1092_));
 sg13g2_nand3_1 _2002_ (.B(_1091_),
    .C(_1092_),
    .A(_1089_),
    .Y(_1093_));
 sg13g2_nor3_1 _2003_ (.A(net54),
    .B(net59),
    .C(_1068_),
    .Y(_1094_));
 sg13g2_nand4_1 _2004_ (.B(net38),
    .C(net36),
    .A(_1031_),
    .Y(_1095_),
    .D(_1094_));
 sg13g2_inv_1 _2005_ (.Y(_1096_),
    .A(_1068_));
 sg13g2_nand4_1 _2006_ (.B(net37),
    .C(net36),
    .A(_1096_),
    .Y(_1097_),
    .D(_1036_));
 sg13g2_or4_1 _2007_ (.A(_1068_),
    .B(net31),
    .C(net36),
    .D(_1033_),
    .X(_1098_));
 sg13g2_nand4_1 _2008_ (.B(net31),
    .C(net36),
    .A(_1096_),
    .Y(_1099_),
    .D(_1037_));
 sg13g2_nand4_1 _2009_ (.B(_1097_),
    .C(_1098_),
    .A(_1095_),
    .Y(_1100_),
    .D(_1099_));
 sg13g2_a21oi_1 _2010_ (.A1(net62),
    .A2(_1093_),
    .Y(_1101_),
    .B1(_1100_));
 sg13g2_nand2_2 _2011_ (.Y(_1102_),
    .A(_1088_),
    .B(_1101_));
 sg13g2_nor3_2 _2012_ (.A(_1067_),
    .B(net24),
    .C(_1102_),
    .Y(_1103_));
 sg13g2_inv_1 _2013_ (.Y(net11),
    .A(_1103_));
 sg13g2_buf_1 _2014_ (.A(_1069_),
    .X(net12));
 sg13g2_nand3_1 _2015_ (.B(_0981_),
    .C(_0989_),
    .A(_0255_),
    .Y(_1104_));
 sg13g2_a21oi_1 _2016_ (.A1(_0981_),
    .A2(_0989_),
    .Y(_1105_),
    .B1(net59));
 sg13g2_a21oi_1 _2017_ (.A1(net54),
    .A2(_1104_),
    .Y(_1106_),
    .B1(_1105_));
 sg13g2_nor2_1 _2018_ (.A(_1039_),
    .B(_1106_),
    .Y(_1107_));
 sg13g2_nor2b_1 _2019_ (.A(_1107_),
    .B_N(_1025_),
    .Y(_1108_));
 sg13g2_buf_2 _2020_ (.A(_1108_),
    .X(_1109_));
 sg13g2_inv_1 _2021_ (.Y(_1110_),
    .A(_1109_));
 sg13g2_buf_1 _2022_ (.A(_1110_),
    .X(net13));
 sg13g2_nor2_1 _2023_ (.A(_1031_),
    .B(_1009_),
    .Y(_1111_));
 sg13g2_nor2_2 _2024_ (.A(_1057_),
    .B(_1111_),
    .Y(_1112_));
 sg13g2_inv_1 _2025_ (.Y(net14),
    .A(_1112_));
 sg13g2_buf_1 _2026_ (.A(ui_in[3]),
    .X(_1113_));
 sg13g2_buf_1 _2027_ (.A(_1113_),
    .X(_1114_));
 sg13g2_nor3_1 _2028_ (.A(net71),
    .B(net64),
    .C(net72),
    .Y(_1115_));
 sg13g2_nor2b_1 _2029_ (.A(net68),
    .B_N(_1115_),
    .Y(_1116_));
 sg13g2_nor2_1 _2030_ (.A(net70),
    .B(net69),
    .Y(_1117_));
 sg13g2_nand2_1 _2031_ (.Y(_1118_),
    .A(_1116_),
    .B(_1117_));
 sg13g2_xor2_1 _2032_ (.B(_1118_),
    .A(net65),
    .X(_1119_));
 sg13g2_xnor2_1 _2033_ (.Y(_1120_),
    .A(_0364_),
    .B(_1119_));
 sg13g2_inv_1 _2034_ (.Y(_1121_),
    .A(_1120_));
 sg13g2_nor2b_1 _2035_ (.A(net70),
    .B_N(_0010_),
    .Y(_1122_));
 sg13g2_nand2_1 _2036_ (.Y(_1123_),
    .A(_1115_),
    .B(_1122_));
 sg13g2_xor2_1 _2037_ (.B(_1123_),
    .A(net68),
    .X(_1124_));
 sg13g2_inv_1 _2038_ (.Y(_1125_),
    .A(_0016_));
 sg13g2_nor2b_1 _2039_ (.A(_0458_),
    .B_N(_0457_),
    .Y(_1126_));
 sg13g2_o21ai_1 _2040_ (.B1(net69),
    .Y(_1127_),
    .A1(_1125_),
    .A2(_1126_));
 sg13g2_inv_1 _2041_ (.Y(_1128_),
    .A(_0461_));
 sg13g2_a21oi_1 _2042_ (.A1(_1128_),
    .A2(_1125_),
    .Y(_1129_),
    .B1(_0462_));
 sg13g2_mux2_1 _2043_ (.A0(_1127_),
    .A1(_1129_),
    .S(net70),
    .X(_1130_));
 sg13g2_xnor2_1 _2044_ (.Y(_1131_),
    .A(_0455_),
    .B(_1117_));
 sg13g2_xnor2_1 _2045_ (.Y(_1132_),
    .A(_0456_),
    .B(_1131_));
 sg13g2_nand2b_1 _2046_ (.Y(_1133_),
    .B(_1131_),
    .A_N(_0014_));
 sg13g2_o21ai_1 _2047_ (.B1(_1133_),
    .Y(_1134_),
    .A1(_1130_),
    .A2(_1132_));
 sg13g2_nor2b_1 _2048_ (.A(net71),
    .B_N(_1122_),
    .Y(_1135_));
 sg13g2_xnor2_1 _2049_ (.Y(_1136_),
    .A(net64),
    .B(_1135_));
 sg13g2_xnor2_1 _2050_ (.Y(_1137_),
    .A(_0671_),
    .B(_1136_));
 sg13g2_inv_1 _2051_ (.Y(_1138_),
    .A(_0013_));
 sg13g2_and2_1 _2052_ (.A(_1138_),
    .B(_1136_),
    .X(_1139_));
 sg13g2_a21o_1 _2053_ (.A2(_1137_),
    .A1(_1134_),
    .B1(_1139_),
    .X(_1140_));
 sg13g2_nor4_1 _2054_ (.A(net70),
    .B(net69),
    .C(net71),
    .D(net64),
    .Y(_1141_));
 sg13g2_xnor2_1 _2055_ (.Y(_1142_),
    .A(net72),
    .B(_1141_));
 sg13g2_xnor2_1 _2056_ (.Y(_1143_),
    .A(net86),
    .B(_1142_));
 sg13g2_inv_1 _2057_ (.Y(_1144_),
    .A(_1143_));
 sg13g2_nor2b_1 _2058_ (.A(_0012_),
    .B_N(_1142_),
    .Y(_1145_));
 sg13g2_a21o_1 _2059_ (.A2(_1144_),
    .A1(_1140_),
    .B1(_1145_),
    .X(_1146_));
 sg13g2_nor2_1 _2060_ (.A(_1124_),
    .B(_1146_),
    .Y(_1147_));
 sg13g2_a21oi_1 _2061_ (.A1(_1124_),
    .A2(_1146_),
    .Y(_1148_),
    .B1(_0375_));
 sg13g2_or3_1 _2062_ (.A(_1121_),
    .B(_1147_),
    .C(_1148_),
    .X(_1149_));
 sg13g2_nand2b_1 _2063_ (.Y(_1150_),
    .B(_1119_),
    .A_N(_0011_));
 sg13g2_nor2b_1 _2064_ (.A(net65),
    .B_N(_1116_),
    .Y(_1151_));
 sg13g2_nand2_1 _2065_ (.Y(_1152_),
    .A(_1151_),
    .B(_1122_));
 sg13g2_xor2_1 _2066_ (.B(_1152_),
    .A(_0008_),
    .X(_1153_));
 sg13g2_xnor2_1 _2067_ (.Y(_1154_),
    .A(net76),
    .B(_1153_));
 sg13g2_a21oi_1 _2068_ (.A1(_1149_),
    .A2(_1150_),
    .Y(_1155_),
    .B1(_1154_));
 sg13g2_and2_1 _2069_ (.A(_0444_),
    .B(_1153_),
    .X(_1156_));
 sg13g2_nand2_1 _2070_ (.Y(_1157_),
    .A(_1151_),
    .B(_1117_));
 sg13g2_nand2_1 _2071_ (.Y(_1158_),
    .A(net66),
    .B(_1157_));
 sg13g2_xnor2_1 _2072_ (.Y(_1159_),
    .A(_0809_),
    .B(_1158_));
 sg13g2_xnor2_1 _2073_ (.Y(_1160_),
    .A(net74),
    .B(_1159_));
 sg13g2_o21ai_1 _2074_ (.B1(_1160_),
    .Y(_1161_),
    .A1(_1155_),
    .A2(_1156_));
 sg13g2_or3_1 _2075_ (.A(_1155_),
    .B(_1156_),
    .C(_1160_),
    .X(_1162_));
 sg13g2_buf_1 _2076_ (.A(_1162_),
    .X(_1163_));
 sg13g2_and2_1 _2077_ (.A(_1161_),
    .B(_1163_),
    .X(_1164_));
 sg13g2_a21o_1 _2078_ (.A2(_1150_),
    .A1(_1149_),
    .B1(_1154_),
    .X(_1165_));
 sg13g2_buf_1 _2079_ (.A(_1165_),
    .X(_1166_));
 sg13g2_nand2_1 _2080_ (.Y(_1167_),
    .A(_0444_),
    .B(_1153_));
 sg13g2_nor2_1 _2081_ (.A(net58),
    .B(_1159_),
    .Y(_1168_));
 sg13g2_a21oi_2 _2082_ (.B1(_1168_),
    .Y(_1169_),
    .A2(_1167_),
    .A1(_1166_));
 sg13g2_and2_1 _2083_ (.A(net58),
    .B(_1159_),
    .X(_1170_));
 sg13g2_nor2_2 _2084_ (.A(_1169_),
    .B(_1170_),
    .Y(_1171_));
 sg13g2_a21oi_1 _2085_ (.A1(net66),
    .A2(_1152_),
    .Y(_1172_),
    .B1(net57));
 sg13g2_xnor2_1 _2086_ (.Y(_1173_),
    .A(_0481_),
    .B(_1172_));
 sg13g2_xnor2_1 _2087_ (.Y(_1174_),
    .A(_0309_),
    .B(_1173_));
 sg13g2_buf_1 _2088_ (.A(_1174_),
    .X(_1175_));
 sg13g2_nand3_1 _2089_ (.B(_1150_),
    .C(_1154_),
    .A(_1149_),
    .Y(_1176_));
 sg13g2_nor2_2 _2090_ (.A(_0006_),
    .B(_1173_),
    .Y(_1177_));
 sg13g2_a21oi_2 _2091_ (.B1(_1177_),
    .Y(_1178_),
    .A2(_1176_),
    .A1(_1166_));
 sg13g2_and3_1 _2092_ (.X(_1179_),
    .A(_1166_),
    .B(_1176_),
    .C(_1177_));
 sg13g2_a21oi_1 _2093_ (.A1(net66),
    .A2(_1157_),
    .Y(_1180_),
    .B1(net57));
 sg13g2_nand2b_1 _2094_ (.Y(_1181_),
    .B(_0481_),
    .A_N(_1180_));
 sg13g2_buf_1 _2095_ (.A(_1181_),
    .X(_1182_));
 sg13g2_mux2_1 _2096_ (.A0(_1178_),
    .A1(_1179_),
    .S(_1182_),
    .X(_1183_));
 sg13g2_nand3_1 _2097_ (.B(net46),
    .C(_1183_),
    .A(_1171_),
    .Y(_1184_));
 sg13g2_a21o_1 _2098_ (.A2(_1167_),
    .A1(_1166_),
    .B1(_1168_),
    .X(_1185_));
 sg13g2_buf_1 _2099_ (.A(_1185_),
    .X(_1186_));
 sg13g2_nand2_2 _2100_ (.Y(_1187_),
    .A(net58),
    .B(_1159_));
 sg13g2_nand2_2 _2101_ (.Y(_1188_),
    .A(_1186_),
    .B(_1187_));
 sg13g2_inv_1 _2102_ (.Y(_1189_),
    .A(net46));
 sg13g2_and2_1 _2103_ (.A(_1166_),
    .B(_1176_),
    .X(_1190_));
 sg13g2_buf_1 _2104_ (.A(_1190_),
    .X(_1191_));
 sg13g2_nand4_1 _2105_ (.B(_1189_),
    .C(net47),
    .A(_1188_),
    .Y(_1192_),
    .D(net40));
 sg13g2_nand2_1 _2106_ (.Y(_1193_),
    .A(_1184_),
    .B(_1192_));
 sg13g2_nand2_2 _2107_ (.Y(_1194_),
    .A(_1161_),
    .B(_1163_));
 sg13g2_inv_1 _2108_ (.Y(_1195_),
    .A(net40));
 sg13g2_nand3_1 _2109_ (.B(_1195_),
    .C(_1177_),
    .A(_1182_),
    .Y(_1196_));
 sg13g2_nor3_1 _2110_ (.A(net47),
    .B(_1178_),
    .C(_1179_),
    .Y(_1197_));
 sg13g2_nor2_1 _2111_ (.A(_1194_),
    .B(_1197_),
    .Y(_1198_));
 sg13g2_nand2_1 _2112_ (.Y(_1199_),
    .A(net47),
    .B(_1178_));
 sg13g2_a22oi_1 _2113_ (.Y(_1200_),
    .B1(_1198_),
    .B2(_1199_),
    .A2(_1196_),
    .A1(_1194_));
 sg13g2_xnor2_1 _2114_ (.Y(_1201_),
    .A(_1171_),
    .B(_1189_));
 sg13g2_a22oi_1 _2115_ (.Y(_1202_),
    .B1(_1200_),
    .B2(_1201_),
    .A2(_1193_),
    .A1(_1164_));
 sg13g2_nor2b_1 _2116_ (.A(net81),
    .B_N(_0006_),
    .Y(_1203_));
 sg13g2_a21o_1 _2117_ (.A2(_1202_),
    .A1(net81),
    .B1(_1203_),
    .X(_1204_));
 sg13g2_buf_1 _2118_ (.A(_1204_),
    .X(_1205_));
 sg13g2_nor3_1 _2119_ (.A(_1169_),
    .B(_1170_),
    .C(_1177_),
    .Y(_1206_));
 sg13g2_or2_1 _2120_ (.X(_1207_),
    .B(_1173_),
    .A(_0006_));
 sg13g2_buf_1 _2121_ (.A(_1207_),
    .X(_1208_));
 sg13g2_a21oi_1 _2122_ (.A1(_1186_),
    .A2(_1187_),
    .Y(_1209_),
    .B1(_1208_));
 sg13g2_nor2b_2 _2123_ (.A(_1180_),
    .B_N(_0481_),
    .Y(_1210_));
 sg13g2_o21ai_1 _2124_ (.B1(_1210_),
    .Y(_1211_),
    .A1(_1206_),
    .A2(_1209_));
 sg13g2_nand2_1 _2125_ (.Y(_1212_),
    .A(net46),
    .B(_1208_));
 sg13g2_nor2_1 _2126_ (.A(_1210_),
    .B(_1212_),
    .Y(_1213_));
 sg13g2_a21oi_1 _2127_ (.A1(_1188_),
    .A2(_1213_),
    .Y(_1214_),
    .B1(_1164_));
 sg13g2_nor3_1 _2128_ (.A(_1169_),
    .B(_1170_),
    .C(_1208_),
    .Y(_1215_));
 sg13g2_a21oi_1 _2129_ (.A1(_1186_),
    .A2(_1187_),
    .Y(_1216_),
    .B1(net47));
 sg13g2_a221oi_1 _2130_ (.B2(_1208_),
    .C1(_1194_),
    .B1(_1216_),
    .A1(net47),
    .Y(_1217_),
    .A2(_1215_));
 sg13g2_a21o_1 _2131_ (.A2(_1214_),
    .A1(_1211_),
    .B1(_1217_),
    .X(_1218_));
 sg13g2_inv_2 _2132_ (.Y(_1219_),
    .A(_1113_));
 sg13g2_nor3_1 _2133_ (.A(_1219_),
    .B(_1189_),
    .C(net40),
    .Y(_1220_));
 sg13g2_nand2_1 _2134_ (.Y(_1221_),
    .A(_1218_),
    .B(_1220_));
 sg13g2_and2_1 _2135_ (.A(_1164_),
    .B(_1178_),
    .X(_1222_));
 sg13g2_nor2_1 _2136_ (.A(_1188_),
    .B(net47),
    .Y(_1223_));
 sg13g2_nand2_1 _2137_ (.Y(_1224_),
    .A(_1114_),
    .B(_1189_));
 sg13g2_a221oi_1 _2138_ (.B2(_1223_),
    .C1(_1224_),
    .B1(_1222_),
    .A1(net40),
    .Y(_1225_),
    .A2(_1216_));
 sg13g2_xnor2_1 _2139_ (.Y(_1226_),
    .A(_1210_),
    .B(_1177_));
 sg13g2_nand3_1 _2140_ (.B(_1187_),
    .C(_1226_),
    .A(_1186_),
    .Y(_1227_));
 sg13g2_nand2_1 _2141_ (.Y(_1228_),
    .A(_1210_),
    .B(_1208_));
 sg13g2_and4_1 _2142_ (.A(_1186_),
    .B(_1187_),
    .C(net40),
    .D(_1228_),
    .X(_1229_));
 sg13g2_a21oi_1 _2143_ (.A1(_1195_),
    .A2(_1227_),
    .Y(_1230_),
    .B1(_1229_));
 sg13g2_nor2b_1 _2144_ (.A(net40),
    .B_N(_1212_),
    .Y(_1231_));
 sg13g2_mux2_1 _2145_ (.A0(_1179_),
    .A1(_1231_),
    .S(_1188_),
    .X(_1232_));
 sg13g2_nor2_1 _2146_ (.A(_1194_),
    .B(_1210_),
    .Y(_1233_));
 sg13g2_a22oi_1 _2147_ (.Y(_1234_),
    .B1(_1232_),
    .B2(_1233_),
    .A2(_1230_),
    .A1(_1194_));
 sg13g2_and3_1 _2148_ (.X(_1235_),
    .A(_1186_),
    .B(_1187_),
    .C(_1228_));
 sg13g2_nand3_1 _2149_ (.B(net46),
    .C(net40),
    .A(_1114_),
    .Y(_1236_));
 sg13g2_a221oi_1 _2150_ (.B2(_1194_),
    .C1(_1236_),
    .B1(_1235_),
    .A1(_1171_),
    .Y(_1237_),
    .A2(_1226_));
 sg13g2_a21oi_1 _2151_ (.A1(_1161_),
    .A2(_1163_),
    .Y(_1238_),
    .B1(_1228_));
 sg13g2_and4_1 _2152_ (.A(_1161_),
    .B(_1163_),
    .C(net47),
    .D(_1212_),
    .X(_1239_));
 sg13g2_o21ai_1 _2153_ (.B1(_1188_),
    .Y(_1240_),
    .A1(_1238_),
    .A2(_1239_));
 sg13g2_nor2_1 _2154_ (.A(_0444_),
    .B(net81),
    .Y(_1241_));
 sg13g2_a21o_1 _2155_ (.A2(_1240_),
    .A1(_1237_),
    .B1(_1241_),
    .X(_1242_));
 sg13g2_a21oi_1 _2156_ (.A1(_1225_),
    .A2(_1234_),
    .Y(_1243_),
    .B1(_1242_));
 sg13g2_nand2_1 _2157_ (.Y(_1244_),
    .A(_1221_),
    .B(_1243_));
 sg13g2_nor2_1 _2158_ (.A(_1147_),
    .B(_1148_),
    .Y(_1245_));
 sg13g2_xnor2_1 _2159_ (.Y(_1246_),
    .A(_1121_),
    .B(_1245_));
 sg13g2_nand2_1 _2160_ (.Y(_1247_),
    .A(_0011_),
    .B(_1219_));
 sg13g2_o21ai_1 _2161_ (.B1(_1247_),
    .Y(_1248_),
    .A1(_1219_),
    .A2(_1246_));
 sg13g2_buf_1 _2162_ (.A(_1248_),
    .X(_1249_));
 sg13g2_nand2_1 _2163_ (.Y(_1250_),
    .A(_1124_),
    .B(_1146_));
 sg13g2_nand3b_1 _2164_ (.B(net81),
    .C(_1250_),
    .Y(_1251_),
    .A_N(_1147_));
 sg13g2_xnor2_1 _2165_ (.Y(_1252_),
    .A(_0386_),
    .B(_1251_));
 sg13g2_xnor2_1 _2166_ (.Y(_1253_),
    .A(_1134_),
    .B(_1137_));
 sg13g2_nor2_1 _2167_ (.A(_1138_),
    .B(net81),
    .Y(_1254_));
 sg13g2_a21oi_1 _2168_ (.A1(net81),
    .A2(_1253_),
    .Y(_1255_),
    .B1(_1254_));
 sg13g2_xnor2_1 _2169_ (.Y(_1256_),
    .A(_0460_),
    .B(_0458_));
 sg13g2_nor2_1 _2170_ (.A(_1128_),
    .B(_0457_),
    .Y(_1257_));
 sg13g2_xnor2_1 _2171_ (.Y(_1258_),
    .A(_1256_),
    .B(_1257_));
 sg13g2_nor2_1 _2172_ (.A(_0016_),
    .B(_1113_),
    .Y(_0049_));
 sg13g2_a21oi_1 _2173_ (.A1(_1113_),
    .A2(_1258_),
    .Y(_0050_),
    .B1(_0049_));
 sg13g2_xnor2_1 _2174_ (.Y(_0051_),
    .A(_1130_),
    .B(_1132_));
 sg13g2_mux2_1 _2175_ (.A0(_0014_),
    .A1(_0051_),
    .S(_1113_),
    .X(_0052_));
 sg13g2_nand2_1 _2176_ (.Y(_0053_),
    .A(_0050_),
    .B(_0052_));
 sg13g2_xnor2_1 _2177_ (.Y(_0054_),
    .A(_1140_),
    .B(_1143_));
 sg13g2_nor2_1 _2178_ (.A(_1219_),
    .B(_0054_),
    .Y(_0055_));
 sg13g2_a21oi_2 _2179_ (.B1(_0055_),
    .Y(_0056_),
    .A2(_1219_),
    .A1(_0012_));
 sg13g2_o21ai_1 _2180_ (.B1(_0056_),
    .Y(_0057_),
    .A1(_1255_),
    .A2(_0053_));
 sg13g2_nand4_1 _2181_ (.B(_1249_),
    .C(_1252_),
    .A(_1244_),
    .Y(_0058_),
    .D(_0057_));
 sg13g2_o21ai_1 _2182_ (.B1(net40),
    .Y(_0059_),
    .A1(_1188_),
    .A2(net46));
 sg13g2_nor2_1 _2183_ (.A(net46),
    .B(_1191_),
    .Y(_0060_));
 sg13g2_a21o_1 _2184_ (.A2(_1177_),
    .A1(net46),
    .B1(_0060_),
    .X(_0061_));
 sg13g2_a22oi_1 _2185_ (.Y(_0062_),
    .B1(_0061_),
    .B2(_1188_),
    .A2(_0059_),
    .A1(_1177_));
 sg13g2_nand2_1 _2186_ (.Y(_0063_),
    .A(_1175_),
    .B(_1191_));
 sg13g2_o21ai_1 _2187_ (.B1(_0063_),
    .Y(_0064_),
    .A1(_1188_),
    .A2(_0060_));
 sg13g2_nor2_1 _2188_ (.A(_1164_),
    .B(_1177_),
    .Y(_0065_));
 sg13g2_a21oi_1 _2189_ (.A1(_0064_),
    .A2(_0065_),
    .Y(_0066_),
    .B1(_1210_));
 sg13g2_o21ai_1 _2190_ (.B1(_0066_),
    .Y(_0067_),
    .A1(_1194_),
    .A2(_0062_));
 sg13g2_nor2_1 _2191_ (.A(_1171_),
    .B(net46),
    .Y(_0068_));
 sg13g2_nor2_1 _2192_ (.A(_1189_),
    .B(_1178_),
    .Y(_0069_));
 sg13g2_a21o_1 _2193_ (.A2(_0069_),
    .A1(_1171_),
    .B1(_1179_),
    .X(_0070_));
 sg13g2_o21ai_1 _2194_ (.B1(_1194_),
    .Y(_0071_),
    .A1(_0068_),
    .A2(_0070_));
 sg13g2_a21oi_1 _2195_ (.A1(_1201_),
    .A2(_1222_),
    .Y(_0072_),
    .B1(net47));
 sg13g2_a21oi_1 _2196_ (.A1(_0071_),
    .A2(_0072_),
    .Y(_0073_),
    .B1(_1219_));
 sg13g2_a22oi_1 _2197_ (.Y(_0074_),
    .B1(_0067_),
    .B2(_0073_),
    .A2(_1219_),
    .A1(net58));
 sg13g2_inv_1 _2198_ (.Y(_0075_),
    .A(_0074_));
 sg13g2_nand2_1 _2199_ (.Y(_0076_),
    .A(_0058_),
    .B(_0075_));
 sg13g2_a21oi_1 _2200_ (.A1(_1205_),
    .A2(_0076_),
    .Y(_0077_),
    .B1(_0872_));
 sg13g2_nor3_1 _2201_ (.A(_0145_),
    .B(_0712_),
    .C(_0741_),
    .Y(_0078_));
 sg13g2_nor2b_1 _2202_ (.A(net90),
    .B_N(net1),
    .Y(_0080_));
 sg13g2_o21ai_1 _2203_ (.B1(_0080_),
    .Y(_0081_),
    .A1(_0881_),
    .A2(_0078_));
 sg13g2_buf_1 _2204_ (.A(_0675_),
    .X(_0082_));
 sg13g2_a21oi_1 _2205_ (.A1(_0460_),
    .A2(_0459_),
    .Y(_0083_),
    .B1(_0462_));
 sg13g2_xor2_1 _2206_ (.B(_0083_),
    .A(net71),
    .X(_0084_));
 sg13g2_nor2_1 _2207_ (.A(net85),
    .B(_0084_),
    .Y(_0085_));
 sg13g2_xnor2_1 _2208_ (.Y(_0086_),
    .A(net63),
    .B(_0085_));
 sg13g2_nand2_1 _2209_ (.Y(_0087_),
    .A(_0461_),
    .B(_0457_));
 sg13g2_xnor2_1 _2210_ (.Y(_0088_),
    .A(_0087_),
    .B(_1256_));
 sg13g2_nand2_1 _2211_ (.Y(_0089_),
    .A(net84),
    .B(_0088_));
 sg13g2_o21ai_1 _2212_ (.B1(_0089_),
    .Y(_0091_),
    .A1(net84),
    .A2(_1125_));
 sg13g2_nor2_1 _2213_ (.A(_0086_),
    .B(_0091_),
    .Y(_0092_));
 sg13g2_nand2_1 _2214_ (.Y(_0093_),
    .A(net45),
    .B(_0092_));
 sg13g2_xnor2_1 _2215_ (.Y(_0094_),
    .A(_0640_),
    .B(_0655_));
 sg13g2_nand3_1 _2216_ (.B(_0686_),
    .C(_0094_),
    .A(net45),
    .Y(_0095_));
 sg13g2_o21ai_1 _2217_ (.B1(_0095_),
    .Y(_0096_),
    .A1(_0698_),
    .A2(_0093_));
 sg13g2_inv_1 _2218_ (.Y(_0097_),
    .A(_0086_));
 sg13g2_nor2_1 _2219_ (.A(_0097_),
    .B(_0094_),
    .Y(_0098_));
 sg13g2_nor2_1 _2220_ (.A(net45),
    .B(_0094_),
    .Y(_0099_));
 sg13g2_o21ai_1 _2221_ (.B1(_0698_),
    .Y(_0100_),
    .A1(_0098_),
    .A2(_0099_));
 sg13g2_nor2_1 _2222_ (.A(net45),
    .B(_0686_),
    .Y(_0102_));
 sg13g2_nor2b_1 _2223_ (.A(_0082_),
    .B_N(_0092_),
    .Y(_0103_));
 sg13g2_nor3_1 _2224_ (.A(_0082_),
    .B(_0097_),
    .C(_0094_),
    .Y(_0104_));
 sg13g2_a221oi_1 _2225_ (.B2(_0698_),
    .C1(_0104_),
    .B1(_0103_),
    .A1(_0094_),
    .Y(_0105_),
    .A2(_0102_));
 sg13g2_nand3b_1 _2226_ (.B(_0100_),
    .C(_0105_),
    .Y(_0106_),
    .A_N(_0096_));
 sg13g2_buf_2 _2227_ (.A(_0106_),
    .X(_0107_));
 sg13g2_mux2_1 _2228_ (.A0(net5),
    .A1(net6),
    .S(_0107_),
    .X(_0108_));
 sg13g2_inv_1 _2229_ (.Y(_0109_),
    .A(net45));
 sg13g2_nor2_1 _2230_ (.A(_0109_),
    .B(_0086_),
    .Y(_0110_));
 sg13g2_buf_1 _2231_ (.A(_0655_),
    .X(_0111_));
 sg13g2_a22oi_1 _2232_ (.Y(_0113_),
    .B1(_0110_),
    .B2(net35),
    .A2(_0686_),
    .A1(_0678_));
 sg13g2_or2_1 _2233_ (.X(_0114_),
    .B(_0113_),
    .A(_0640_));
 sg13g2_nor2_1 _2234_ (.A(_0636_),
    .B(net35),
    .Y(_0115_));
 sg13g2_nand2_1 _2235_ (.Y(_0116_),
    .A(_0110_),
    .B(_0115_));
 sg13g2_a21oi_1 _2236_ (.A1(_0655_),
    .A2(net45),
    .Y(_0117_),
    .B1(_0636_));
 sg13g2_nor2_1 _2237_ (.A(net35),
    .B(net45),
    .Y(_0118_));
 sg13g2_inv_1 _2238_ (.Y(_0119_),
    .A(_0686_));
 sg13g2_o21ai_1 _2239_ (.B1(_0119_),
    .Y(_0120_),
    .A1(_0117_),
    .A2(_0118_));
 sg13g2_nand3_1 _2240_ (.B(net39),
    .C(_0686_),
    .A(net35),
    .Y(_0121_));
 sg13g2_nand4_1 _2241_ (.B(_0116_),
    .C(_0120_),
    .A(_0114_),
    .Y(_0122_),
    .D(_0121_));
 sg13g2_nand2_1 _2242_ (.Y(_0124_),
    .A(_0086_),
    .B(_0091_));
 sg13g2_xnor2_1 _2243_ (.Y(_0125_),
    .A(_0109_),
    .B(_0697_));
 sg13g2_or3_1 _2244_ (.A(_0122_),
    .B(_0124_),
    .C(_0125_),
    .X(_0126_));
 sg13g2_and2_1 _2245_ (.A(_0107_),
    .B(_0126_),
    .X(_0127_));
 sg13g2_mux2_1 _2246_ (.A0(net3),
    .A1(net4),
    .S(_0127_),
    .X(_0128_));
 sg13g2_nand2_1 _2247_ (.Y(_0129_),
    .A(_0697_),
    .B(_0104_));
 sg13g2_nand2_2 _2248_ (.Y(_0130_),
    .A(_0122_),
    .B(_0129_));
 sg13g2_mux2_1 _2249_ (.A0(_0108_),
    .A1(_0128_),
    .S(_0130_),
    .X(_0131_));
 sg13g2_nor2b_1 _2250_ (.A(_0131_),
    .B_N(net2),
    .Y(_0132_));
 sg13g2_nor2_1 _2251_ (.A(_0081_),
    .B(_0132_),
    .Y(_0133_));
 sg13g2_a221oi_1 _2252_ (.B2(_1059_),
    .C1(_0710_),
    .B1(_1075_),
    .A1(_1071_),
    .Y(_0135_),
    .A2(_1072_));
 sg13g2_o21ai_1 _2253_ (.B1(_0135_),
    .Y(_0136_),
    .A1(_1096_),
    .A2(_1052_));
 sg13g2_nand2_1 _2254_ (.Y(_0137_),
    .A(net62),
    .B(_1093_));
 sg13g2_and3_1 _2255_ (.X(_0138_),
    .A(_1066_),
    .B(_1088_),
    .C(_0137_));
 sg13g2_buf_1 _2256_ (.A(_1052_),
    .X(_0139_));
 sg13g2_a21oi_1 _2257_ (.A1(_0136_),
    .A2(_0138_),
    .Y(_0140_),
    .B1(net25));
 sg13g2_nor2_1 _2258_ (.A(_0621_),
    .B(_0628_),
    .Y(_0141_));
 sg13g2_nand3_1 _2259_ (.B(_0140_),
    .C(_0141_),
    .A(net27),
    .Y(_0142_));
 sg13g2_buf_1 _2260_ (.A(_0620_),
    .X(_0143_));
 sg13g2_buf_1 _2261_ (.A(_0628_),
    .X(_0144_));
 sg13g2_nand3_1 _2262_ (.B(_1088_),
    .C(_0137_),
    .A(_1066_),
    .Y(_0146_));
 sg13g2_nor4_1 _2263_ (.A(net34),
    .B(net30),
    .C(net24),
    .D(_0146_),
    .Y(_0147_));
 sg13g2_nand2_1 _2264_ (.Y(_0148_),
    .A(_0699_),
    .B(_1068_));
 sg13g2_a221oi_1 _2265_ (.B2(net31),
    .C1(_0148_),
    .B1(_1075_),
    .A1(_1071_),
    .Y(_0149_),
    .A2(_1072_));
 sg13g2_xnor2_1 _2266_ (.Y(_0150_),
    .A(_0731_),
    .B(_1031_));
 sg13g2_mux2_1 _2267_ (.A0(net38),
    .A1(net36),
    .S(_0266_),
    .X(_0151_));
 sg13g2_a22oi_1 _2268_ (.Y(_0152_),
    .B1(_0150_),
    .B2(_0151_),
    .A2(_1047_),
    .A1(_0990_));
 sg13g2_or3_1 _2269_ (.A(_1100_),
    .B(_0149_),
    .C(_0152_),
    .X(_0153_));
 sg13g2_buf_1 _2270_ (.A(_0153_),
    .X(_0154_));
 sg13g2_nand2_1 _2271_ (.Y(_0155_),
    .A(net34),
    .B(net28));
 sg13g2_a21oi_1 _2272_ (.A1(_0154_),
    .A2(_0155_),
    .Y(_0157_),
    .B1(_0697_));
 sg13g2_buf_1 _2273_ (.A(net35),
    .X(_0158_));
 sg13g2_o21ai_1 _2274_ (.B1(net29),
    .Y(_0159_),
    .A1(_0147_),
    .A2(_0157_));
 sg13g2_nor2_1 _2275_ (.A(_0629_),
    .B(_0690_),
    .Y(_0160_));
 sg13g2_inv_1 _2276_ (.Y(_0161_),
    .A(_0160_));
 sg13g2_nor2_1 _2277_ (.A(net33),
    .B(_0161_),
    .Y(_0162_));
 sg13g2_nor2_1 _2278_ (.A(net26),
    .B(_0162_),
    .Y(_0163_));
 sg13g2_nand2_1 _2279_ (.Y(_0164_),
    .A(_0144_),
    .B(_0697_));
 sg13g2_nand2_1 _2280_ (.Y(_0165_),
    .A(net33),
    .B(net29));
 sg13g2_a21oi_1 _2281_ (.A1(net28),
    .A2(net23),
    .Y(_0166_),
    .B1(_0165_));
 sg13g2_o21ai_1 _2282_ (.B1(_0166_),
    .Y(_0168_),
    .A1(_0140_),
    .A2(_0164_));
 sg13g2_nand4_1 _2283_ (.B(_0159_),
    .C(_0163_),
    .A(_0142_),
    .Y(_0169_),
    .D(_0168_));
 sg13g2_nor3_1 _2284_ (.A(_0139_),
    .B(net24),
    .C(_0146_),
    .Y(_0170_));
 sg13g2_nand4_1 _2285_ (.B(_0691_),
    .C(_0693_),
    .A(net35),
    .Y(_0171_),
    .D(_0694_));
 sg13g2_buf_2 _2286_ (.A(_0171_),
    .X(_0172_));
 sg13g2_nor3_2 _2287_ (.A(_0621_),
    .B(_0629_),
    .C(_0172_),
    .Y(_0173_));
 sg13g2_a21oi_1 _2288_ (.A1(_0170_),
    .A2(_0173_),
    .Y(_0174_),
    .B1(_1109_));
 sg13g2_nor2_1 _2289_ (.A(_1112_),
    .B(_0174_),
    .Y(_0175_));
 sg13g2_a221oi_1 _2290_ (.B2(_0724_),
    .C1(_1100_),
    .B1(_1093_),
    .A1(_1068_),
    .Y(_0176_),
    .A2(_0135_));
 sg13g2_a21oi_1 _2291_ (.A1(_1088_),
    .A2(_0176_),
    .Y(_0177_),
    .B1(net23));
 sg13g2_nor2_1 _2292_ (.A(_0620_),
    .B(_0628_),
    .Y(_0179_));
 sg13g2_nor2_1 _2293_ (.A(net27),
    .B(_0179_),
    .Y(_0180_));
 sg13g2_xnor2_1 _2294_ (.Y(_0181_),
    .A(net32),
    .B(_0180_));
 sg13g2_mux2_1 _2295_ (.A0(_0676_),
    .A1(net44),
    .S(_0111_),
    .X(_0182_));
 sg13g2_nor2_1 _2296_ (.A(net39),
    .B(_0182_),
    .Y(_0183_));
 sg13g2_a21oi_1 _2297_ (.A1(net39),
    .A2(_0115_),
    .Y(_0184_),
    .B1(_0183_));
 sg13g2_nor2_1 _2298_ (.A(_0143_),
    .B(_0184_),
    .Y(_0185_));
 sg13g2_a221oi_1 _2299_ (.B2(_0678_),
    .C1(net32),
    .B1(net28),
    .A1(_0600_),
    .Y(_0186_),
    .A2(_0619_));
 sg13g2_nand3_1 _2300_ (.B(_0158_),
    .C(_0692_),
    .A(_0621_),
    .Y(_0187_));
 sg13g2_or2_1 _2301_ (.X(_0188_),
    .B(net35),
    .A(_0640_));
 sg13g2_a21oi_1 _2302_ (.A1(_0187_),
    .A2(_0188_),
    .Y(_0190_),
    .B1(net44));
 sg13g2_o21ai_1 _2303_ (.B1(_0669_),
    .Y(_0191_),
    .A1(_0688_),
    .A2(_0190_));
 sg13g2_and2_1 _2304_ (.A(_0111_),
    .B(_0678_),
    .X(_0192_));
 sg13g2_nand2_1 _2305_ (.Y(_0193_),
    .A(_0620_),
    .B(_0692_));
 sg13g2_nand3_1 _2306_ (.B(_0192_),
    .C(_0193_),
    .A(_0613_),
    .Y(_0194_));
 sg13g2_a21oi_1 _2307_ (.A1(_0191_),
    .A2(_0194_),
    .Y(_0195_),
    .B1(net30));
 sg13g2_nor4_1 _2308_ (.A(_0154_),
    .B(_0185_),
    .C(_0186_),
    .D(_0195_),
    .Y(_0196_));
 sg13g2_a21oi_1 _2309_ (.A1(_0177_),
    .A2(_0181_),
    .Y(_0197_),
    .B1(_0196_));
 sg13g2_nor2_1 _2310_ (.A(net34),
    .B(net32),
    .Y(_0198_));
 sg13g2_a21oi_1 _2311_ (.A1(net32),
    .A2(_0679_),
    .Y(_0199_),
    .B1(_0192_));
 sg13g2_inv_1 _2312_ (.Y(_0201_),
    .A(_0199_));
 sg13g2_nor2_1 _2313_ (.A(net43),
    .B(net39),
    .Y(_0202_));
 sg13g2_a21oi_1 _2314_ (.A1(net43),
    .A2(_0621_),
    .Y(_0203_),
    .B1(_0202_));
 sg13g2_nand2_1 _2315_ (.Y(_0204_),
    .A(net35),
    .B(_0692_));
 sg13g2_a21oi_1 _2316_ (.A1(_0670_),
    .A2(_0676_),
    .Y(_0205_),
    .B1(_0688_));
 sg13g2_o21ai_1 _2317_ (.B1(_0205_),
    .Y(_0206_),
    .A1(_0203_),
    .A2(_0204_));
 sg13g2_o21ai_1 _2318_ (.B1(_0144_),
    .Y(_0207_),
    .A1(_0201_),
    .A2(_0206_));
 sg13g2_nor2_1 _2319_ (.A(_0621_),
    .B(_0656_),
    .Y(_0208_));
 sg13g2_nand2_1 _2320_ (.Y(_0209_),
    .A(_0109_),
    .B(_0669_));
 sg13g2_a22oi_1 _2321_ (.Y(_0210_),
    .B1(_0209_),
    .B2(net29),
    .A2(net39),
    .A1(_0641_));
 sg13g2_nand2_1 _2322_ (.Y(_0212_),
    .A(_0636_),
    .B(net45));
 sg13g2_a21oi_1 _2323_ (.A1(_0620_),
    .A2(_0212_),
    .Y(_0213_),
    .B1(net43));
 sg13g2_nor3_1 _2324_ (.A(_0208_),
    .B(_0210_),
    .C(_0213_),
    .Y(_0214_));
 sg13g2_o21ai_1 _2325_ (.B1(_0629_),
    .Y(_0215_),
    .A1(net44),
    .A2(net39));
 sg13g2_nor3_1 _2326_ (.A(net32),
    .B(_0206_),
    .C(_0215_),
    .Y(_0216_));
 sg13g2_or2_1 _2327_ (.X(_0217_),
    .B(_0216_),
    .A(_0214_));
 sg13g2_a21o_1 _2328_ (.A2(_0207_),
    .A1(_0198_),
    .B1(_0217_),
    .X(_0218_));
 sg13g2_a22oi_1 _2329_ (.Y(_0219_),
    .B1(_0218_),
    .B2(net23),
    .A2(_0170_),
    .A1(_0160_));
 sg13g2_nand3_1 _2330_ (.B(_0197_),
    .C(_0219_),
    .A(net26),
    .Y(_0220_));
 sg13g2_a21oi_1 _2331_ (.A1(_0173_),
    .A2(_0177_),
    .Y(_0221_),
    .B1(net26));
 sg13g2_nor2_1 _2332_ (.A(net14),
    .B(_0221_),
    .Y(_0223_));
 sg13g2_a221oi_1 _2333_ (.B2(_0223_),
    .C1(_0130_),
    .B1(_0220_),
    .A1(_0169_),
    .Y(_0224_),
    .A2(_0175_));
 sg13g2_o21ai_1 _2334_ (.B1(_0198_),
    .Y(_0225_),
    .A1(_1078_),
    .A2(_1102_));
 sg13g2_nand2_1 _2335_ (.Y(_0226_),
    .A(_0165_),
    .B(_0697_));
 sg13g2_or4_1 _2336_ (.A(_1067_),
    .B(net24),
    .C(_1102_),
    .D(_0226_),
    .X(_0227_));
 sg13g2_and4_1 _2337_ (.A(_1030_),
    .B(_1040_),
    .C(_1050_),
    .D(_1110_),
    .X(_0228_));
 sg13g2_and2_1 _2338_ (.A(net28),
    .B(_0228_),
    .X(_0229_));
 sg13g2_inv_1 _2339_ (.Y(_0230_),
    .A(_0229_));
 sg13g2_a21oi_1 _2340_ (.A1(_0225_),
    .A2(_0227_),
    .Y(_0231_),
    .B1(_0230_));
 sg13g2_nor4_1 _2341_ (.A(net33),
    .B(_1069_),
    .C(_1110_),
    .D(_0161_),
    .Y(_0232_));
 sg13g2_o21ai_1 _2342_ (.B1(_0232_),
    .Y(_0234_),
    .A1(net24),
    .A2(_1102_));
 sg13g2_a21oi_1 _2343_ (.A1(net33),
    .A2(_0172_),
    .Y(_0235_),
    .B1(_0208_));
 sg13g2_nor2_1 _2344_ (.A(_1052_),
    .B(_1110_),
    .Y(_0236_));
 sg13g2_a22oi_1 _2345_ (.Y(_0237_),
    .B1(_0236_),
    .B2(_0173_),
    .A2(_0229_),
    .A1(_0235_));
 sg13g2_and4_1 _2346_ (.A(_1112_),
    .B(_0130_),
    .C(_0234_),
    .D(_0237_),
    .X(_0238_));
 sg13g2_inv_1 _2347_ (.Y(_0239_),
    .A(_0185_));
 sg13g2_a21oi_1 _2348_ (.A1(net29),
    .A2(_0172_),
    .Y(_0240_),
    .B1(_0628_));
 sg13g2_nor2_1 _2349_ (.A(net33),
    .B(_0240_),
    .Y(_0241_));
 sg13g2_nand2_1 _2350_ (.Y(_0242_),
    .A(net32),
    .B(_0179_));
 sg13g2_nand2_1 _2351_ (.Y(_0243_),
    .A(net30),
    .B(net29));
 sg13g2_nand3_1 _2352_ (.B(_0242_),
    .C(_0243_),
    .A(net26),
    .Y(_0245_));
 sg13g2_nor3_1 _2353_ (.A(net25),
    .B(_0241_),
    .C(_0245_),
    .Y(_0246_));
 sg13g2_o21ai_1 _2354_ (.B1(_0246_),
    .Y(_0247_),
    .A1(_1103_),
    .A2(_0239_));
 sg13g2_nand3b_1 _2355_ (.B(_0238_),
    .C(_0247_),
    .Y(_0248_),
    .A_N(_0231_));
 sg13g2_nand3_1 _2356_ (.B(net30),
    .C(net32),
    .A(net33),
    .Y(_0249_));
 sg13g2_nand2_1 _2357_ (.Y(_0250_),
    .A(net27),
    .B(_0208_));
 sg13g2_a21o_1 _2358_ (.A2(_0250_),
    .A1(_0249_),
    .B1(_1103_),
    .X(_0251_));
 sg13g2_nor3_1 _2359_ (.A(_0143_),
    .B(net10),
    .C(net8),
    .Y(_0252_));
 sg13g2_nor2_1 _2360_ (.A(_0697_),
    .B(_0249_),
    .Y(_0253_));
 sg13g2_a21oi_1 _2361_ (.A1(_1103_),
    .A2(_0252_),
    .Y(_0254_),
    .B1(_0253_));
 sg13g2_nand2_1 _2362_ (.Y(_0256_),
    .A(_0139_),
    .B(net26));
 sg13g2_a21oi_1 _2363_ (.A1(_0251_),
    .A2(_0254_),
    .Y(_0257_),
    .B1(_0256_));
 sg13g2_nand3_1 _2364_ (.B(_0136_),
    .C(_0138_),
    .A(net23),
    .Y(_0258_));
 sg13g2_nor2_1 _2365_ (.A(net34),
    .B(net28),
    .Y(_0259_));
 sg13g2_nand2_1 _2366_ (.Y(_0260_),
    .A(_0172_),
    .B(_0690_));
 sg13g2_a22oi_1 _2367_ (.Y(_0261_),
    .B1(_0240_),
    .B2(net34),
    .A2(_0260_),
    .A1(_0259_));
 sg13g2_nand4_1 _2368_ (.B(_1088_),
    .C(_0176_),
    .A(net34),
    .Y(_0262_),
    .D(_0240_));
 sg13g2_o21ai_1 _2369_ (.B1(_0262_),
    .Y(_0263_),
    .A1(net25),
    .A2(_0261_));
 sg13g2_nand2_1 _2370_ (.Y(_0264_),
    .A(net29),
    .B(_0179_));
 sg13g2_a21oi_1 _2371_ (.A1(_0161_),
    .A2(_0264_),
    .Y(_0265_),
    .B1(_0154_));
 sg13g2_a21oi_1 _2372_ (.A1(_0258_),
    .A2(_0263_),
    .Y(_0267_),
    .B1(_0265_));
 sg13g2_nand2_1 _2373_ (.Y(_0268_),
    .A(_1109_),
    .B(_0127_));
 sg13g2_a21oi_1 _2374_ (.A1(net28),
    .A2(net29),
    .Y(_0269_),
    .B1(net34));
 sg13g2_o21ai_1 _2375_ (.B1(_0269_),
    .Y(_0270_),
    .A1(net28),
    .A2(_0690_));
 sg13g2_nand3b_1 _2376_ (.B(_0270_),
    .C(_1109_),
    .Y(_0271_),
    .A_N(_0241_));
 sg13g2_nor4_1 _2377_ (.A(net25),
    .B(net24),
    .C(_0146_),
    .D(_0271_),
    .Y(_0272_));
 sg13g2_a21o_1 _2378_ (.A2(_0176_),
    .A1(_1088_),
    .B1(net23),
    .X(_0273_));
 sg13g2_a221oi_1 _2379_ (.B2(_0228_),
    .C1(_1112_),
    .B1(_0173_),
    .A1(_0122_),
    .Y(_0274_),
    .A2(_0129_));
 sg13g2_o21ai_1 _2380_ (.B1(_0274_),
    .Y(_0275_),
    .A1(_0273_),
    .A2(_0271_));
 sg13g2_o21ai_1 _2381_ (.B1(_0127_),
    .Y(_0276_),
    .A1(_0272_),
    .A2(_0275_));
 sg13g2_o21ai_1 _2382_ (.B1(_0276_),
    .Y(_0278_),
    .A1(_0267_),
    .A2(_0268_));
 sg13g2_o21ai_1 _2383_ (.B1(_0278_),
    .Y(_0279_),
    .A1(_0248_),
    .A2(_0257_));
 sg13g2_a221oi_1 _2384_ (.B2(_0173_),
    .C1(_1109_),
    .B1(_0170_),
    .A1(net25),
    .Y(_0280_),
    .A2(_0162_));
 sg13g2_nor4_1 _2385_ (.A(_1112_),
    .B(_0130_),
    .C(_0107_),
    .D(_0280_),
    .Y(_0281_));
 sg13g2_o21ai_1 _2386_ (.B1(_1068_),
    .Y(_0282_),
    .A1(_1069_),
    .A2(_1077_));
 sg13g2_nand4_1 _2387_ (.B(net61),
    .C(net31),
    .A(_0717_),
    .Y(_0283_),
    .D(net36));
 sg13g2_nor2_1 _2388_ (.A(net61),
    .B(net38),
    .Y(_0284_));
 sg13g2_nor3_1 _2389_ (.A(_0266_),
    .B(net31),
    .C(net37),
    .Y(_0285_));
 sg13g2_o21ai_1 _2390_ (.B1(_1009_),
    .Y(_0286_),
    .A1(_0284_),
    .A2(_0285_));
 sg13g2_nand4_1 _2391_ (.B(_1056_),
    .C(_0283_),
    .A(_1096_),
    .Y(_0287_),
    .D(_0286_));
 sg13g2_a21o_1 _2392_ (.A2(_0135_),
    .A1(_1069_),
    .B1(_0287_),
    .X(_0288_));
 sg13g2_nand4_1 _2393_ (.B(_1066_),
    .C(_1088_),
    .A(net27),
    .Y(_0289_),
    .D(_0137_));
 sg13g2_a21o_1 _2394_ (.A2(_0288_),
    .A1(_0282_),
    .B1(_0289_),
    .X(_0290_));
 sg13g2_a21oi_1 _2395_ (.A1(net27),
    .A2(net25),
    .Y(_0291_),
    .B1(net30));
 sg13g2_nand4_1 _2396_ (.B(_1066_),
    .C(_1088_),
    .A(_0696_),
    .Y(_0292_),
    .D(_0137_));
 sg13g2_a21oi_1 _2397_ (.A1(_0282_),
    .A2(_0288_),
    .Y(_0293_),
    .B1(_0292_));
 sg13g2_a221oi_1 _2398_ (.B2(_0291_),
    .C1(_0293_),
    .B1(_0290_),
    .A1(_0696_),
    .Y(_0294_),
    .A2(net25));
 sg13g2_o21ai_1 _2399_ (.B1(_0690_),
    .Y(_0295_),
    .A1(net30),
    .A2(_0172_));
 sg13g2_a21o_1 _2400_ (.A2(_0295_),
    .A1(_0154_),
    .B1(net33),
    .X(_0296_));
 sg13g2_nand2_1 _2401_ (.Y(_0297_),
    .A(_0136_),
    .B(_0138_));
 sg13g2_nor2_1 _2402_ (.A(net25),
    .B(_0264_),
    .Y(_0299_));
 sg13g2_o21ai_1 _2403_ (.B1(_1109_),
    .Y(_0300_),
    .A1(net27),
    .A2(_0242_));
 sg13g2_a21oi_1 _2404_ (.A1(_0297_),
    .A2(_0299_),
    .Y(_0301_),
    .B1(_0300_));
 sg13g2_o21ai_1 _2405_ (.B1(_0301_),
    .Y(_0302_),
    .A1(_0294_),
    .A2(_0296_));
 sg13g2_nor4_1 _2406_ (.A(_0690_),
    .B(net23),
    .C(net24),
    .D(_1102_),
    .Y(_0303_));
 sg13g2_and2_1 _2407_ (.A(net26),
    .B(_0259_),
    .X(_0304_));
 sg13g2_o21ai_1 _2408_ (.B1(_0304_),
    .Y(_0305_),
    .A1(net29),
    .A2(_0303_));
 sg13g2_and2_1 _2409_ (.A(_1112_),
    .B(_0234_),
    .X(_0306_));
 sg13g2_nand4_1 _2410_ (.B(_0696_),
    .C(net26),
    .A(net30),
    .Y(_0307_),
    .D(_0258_));
 sg13g2_nand4_1 _2411_ (.B(net23),
    .C(net11),
    .A(net27),
    .Y(_0308_),
    .D(_0304_));
 sg13g2_nand4_1 _2412_ (.B(_0306_),
    .C(_0307_),
    .A(_0305_),
    .Y(_0310_),
    .D(_0308_));
 sg13g2_nand2_1 _2413_ (.Y(_0311_),
    .A(_0107_),
    .B(_0126_));
 sg13g2_nand2_1 _2414_ (.Y(_0312_),
    .A(net26),
    .B(_0162_));
 sg13g2_nor2_1 _2415_ (.A(net34),
    .B(_0690_),
    .Y(_0313_));
 sg13g2_nor2_1 _2416_ (.A(net9),
    .B(_0260_),
    .Y(_0314_));
 sg13g2_nor3_1 _2417_ (.A(net28),
    .B(_0313_),
    .C(_0314_),
    .Y(_0315_));
 sg13g2_a21oi_1 _2418_ (.A1(_1109_),
    .A2(_0315_),
    .Y(_0316_),
    .B1(_1112_));
 sg13g2_o21ai_1 _2419_ (.B1(_0316_),
    .Y(_0317_),
    .A1(_0140_),
    .A2(_0312_));
 sg13g2_and3_1 _2420_ (.X(_0318_),
    .A(_0130_),
    .B(_0311_),
    .C(_0317_));
 sg13g2_a221oi_1 _2421_ (.B2(_0177_),
    .C1(net13),
    .B1(_0173_),
    .A1(net23),
    .Y(_0319_),
    .A2(_0162_));
 sg13g2_nor4_1 _2422_ (.A(net14),
    .B(_0130_),
    .C(_0107_),
    .D(_0319_),
    .Y(_0321_));
 sg13g2_nor2_1 _2423_ (.A(net24),
    .B(_0146_),
    .Y(_0322_));
 sg13g2_nand4_1 _2424_ (.B(net7),
    .C(net12),
    .A(net8),
    .Y(_0323_),
    .D(_0141_));
 sg13g2_nand2_1 _2425_ (.Y(_0324_),
    .A(_0158_),
    .B(_0141_));
 sg13g2_a21oi_1 _2426_ (.A1(_0242_),
    .A2(_0324_),
    .Y(_0325_),
    .B1(net7));
 sg13g2_a21oi_1 _2427_ (.A1(net9),
    .A2(_0698_),
    .Y(_0326_),
    .B1(net30));
 sg13g2_mux2_1 _2428_ (.A0(_0326_),
    .A1(_0173_),
    .S(_0154_),
    .X(_0327_));
 sg13g2_nor3_1 _2429_ (.A(_1109_),
    .B(_0325_),
    .C(_0327_),
    .Y(_0328_));
 sg13g2_o21ai_1 _2430_ (.B1(_0328_),
    .Y(_0329_),
    .A1(_0322_),
    .A2(_0323_));
 sg13g2_a21o_1 _2431_ (.A2(_0329_),
    .A1(_0321_),
    .B1(net2),
    .X(_0330_));
 sg13g2_a221oi_1 _2432_ (.B2(_0318_),
    .C1(_0330_),
    .B1(_0310_),
    .A1(_0281_),
    .Y(_0332_),
    .A2(_0302_));
 sg13g2_o21ai_1 _2433_ (.B1(_0332_),
    .Y(_0333_),
    .A1(_0224_),
    .A2(_0279_));
 sg13g2_a21o_1 _2434_ (.A2(_1253_),
    .A1(net81),
    .B1(_1254_),
    .X(_0334_));
 sg13g2_or2_1 _2435_ (.X(_0335_),
    .B(_0052_),
    .A(_0050_));
 sg13g2_nand2_1 _2436_ (.Y(_0336_),
    .A(_0334_),
    .B(_0335_));
 sg13g2_xnor2_1 _2437_ (.Y(_0337_),
    .A(net73),
    .B(_1251_));
 sg13g2_o21ai_1 _2438_ (.B1(_0337_),
    .Y(_0338_),
    .A1(_0056_),
    .A2(_0336_));
 sg13g2_and4_1 _2439_ (.A(_1244_),
    .B(_1249_),
    .C(_0074_),
    .D(_0338_),
    .X(_0339_));
 sg13g2_nand2_1 _2440_ (.Y(_0340_),
    .A(_0134_),
    .B(net88));
 sg13g2_o21ai_1 _2441_ (.B1(_0752_),
    .Y(_0341_),
    .A1(_0340_),
    .A2(_0929_));
 sg13g2_a21o_1 _2442_ (.A2(_0341_),
    .A1(net80),
    .B1(_0079_),
    .X(_0343_));
 sg13g2_a21oi_1 _2443_ (.A1(net81),
    .A2(_1202_),
    .Y(_0344_),
    .B1(_1203_));
 sg13g2_nor2_1 _2444_ (.A(_0334_),
    .B(_0335_),
    .Y(_0345_));
 sg13g2_o21ai_1 _2445_ (.B1(_0337_),
    .Y(_0346_),
    .A1(_0056_),
    .A2(_0345_));
 sg13g2_or2_1 _2446_ (.X(_0347_),
    .B(_0346_),
    .A(_1249_));
 sg13g2_a21oi_1 _2447_ (.A1(_1255_),
    .A2(_0053_),
    .Y(_0348_),
    .B1(_0056_));
 sg13g2_a21oi_1 _2448_ (.A1(_1252_),
    .A2(_0348_),
    .Y(_0349_),
    .B1(_1249_));
 sg13g2_a221oi_1 _2449_ (.B2(_1234_),
    .C1(_1242_),
    .B1(_1225_),
    .A1(_1218_),
    .Y(_0350_),
    .A2(_1220_));
 sg13g2_mux2_1 _2450_ (.A0(_0347_),
    .A1(_0349_),
    .S(_0350_),
    .X(_0351_));
 sg13g2_nor3_1 _2451_ (.A(_0344_),
    .B(_0074_),
    .C(_0351_),
    .Y(_0352_));
 sg13g2_nor2_1 _2452_ (.A(_0343_),
    .B(_0352_),
    .Y(_0354_));
 sg13g2_o21ai_1 _2453_ (.B1(_0354_),
    .Y(_0355_),
    .A1(_1205_),
    .A2(_0339_));
 sg13g2_o21ai_1 _2454_ (.B1(_0013_),
    .Y(_0356_),
    .A1(net83),
    .A2(_0768_));
 sg13g2_a21o_1 _2455_ (.A2(_0356_),
    .A1(net86),
    .B1(net73),
    .X(_0357_));
 sg13g2_a21oi_1 _2456_ (.A1(net75),
    .A2(_0357_),
    .Y(_0358_),
    .B1(net76));
 sg13g2_o21ai_1 _2457_ (.B1(_0309_),
    .Y(_0359_),
    .A1(_0447_),
    .A2(_0358_));
 sg13g2_a21oi_2 _2458_ (.B1(net90),
    .Y(_0360_),
    .A2(_0712_),
    .A1(net80));
 sg13g2_a21oi_1 _2459_ (.A1(_0343_),
    .A2(_0359_),
    .Y(_0361_),
    .B1(_0360_));
 sg13g2_nand2_1 _2460_ (.Y(_0362_),
    .A(_0081_),
    .B(_0360_));
 sg13g2_nor2_1 _2461_ (.A(_0344_),
    .B(_0362_),
    .Y(_0363_));
 sg13g2_a22oi_1 _2462_ (.Y(_0365_),
    .B1(_0363_),
    .B2(_0076_),
    .A2(_0361_),
    .A1(_0355_));
 sg13g2_nand2_1 _2463_ (.Y(_0366_),
    .A(_0872_),
    .B(_0365_));
 sg13g2_a21oi_1 _2464_ (.A1(_0133_),
    .A2(_0333_),
    .Y(_0367_),
    .B1(_0366_));
 sg13g2_nand4_1 _2465_ (.B(_0058_),
    .C(_0075_),
    .A(_1205_),
    .Y(_0368_),
    .D(_0351_));
 sg13g2_nand3_1 _2466_ (.B(_0056_),
    .C(_0336_),
    .A(_0337_),
    .Y(_0369_));
 sg13g2_a21o_1 _2467_ (.A2(_0369_),
    .A1(_1249_),
    .B1(_1244_),
    .X(_0370_));
 sg13g2_nand3_1 _2468_ (.B(_0074_),
    .C(_0370_),
    .A(_1205_),
    .Y(_0371_));
 sg13g2_nand2_1 _2469_ (.Y(_0372_),
    .A(_0344_),
    .B(_0339_));
 sg13g2_nand3_1 _2470_ (.B(_0371_),
    .C(_0372_),
    .A(_0368_),
    .Y(_0373_));
 sg13g2_nand3_1 _2471_ (.B(_1255_),
    .C(_0053_),
    .A(_0056_),
    .Y(_0374_));
 sg13g2_a21o_1 _2472_ (.A2(_0374_),
    .A1(_1252_),
    .B1(_1249_),
    .X(_0376_));
 sg13g2_nand4_1 _2473_ (.B(_1244_),
    .C(_0074_),
    .A(_1205_),
    .Y(_0377_),
    .D(_0376_));
 sg13g2_inv_1 _2474_ (.Y(_0378_),
    .A(_0377_));
 sg13g2_a21oi_1 _2475_ (.A1(_0872_),
    .A2(_0362_),
    .Y(_0379_),
    .B1(_0378_));
 sg13g2_nand3_1 _2476_ (.B(net86),
    .C(_0522_),
    .A(_0437_),
    .Y(_0380_));
 sg13g2_nor4_1 _2477_ (.A(_1125_),
    .B(net63),
    .C(_0466_),
    .D(_1126_),
    .Y(_0381_));
 sg13g2_nand2_1 _2478_ (.Y(_0382_),
    .A(_0309_),
    .B(_0447_));
 sg13g2_nor2_1 _2479_ (.A(net76),
    .B(_0382_),
    .Y(_0383_));
 sg13g2_o21ai_1 _2480_ (.B1(_0383_),
    .Y(_0384_),
    .A1(_0380_),
    .A2(_0381_));
 sg13g2_and2_1 _2481_ (.A(_0343_),
    .B(_0384_),
    .X(_0385_));
 sg13g2_nor2_1 _2482_ (.A(net83),
    .B(net86),
    .Y(_0387_));
 sg13g2_nand2b_1 _2483_ (.Y(_0388_),
    .B(_0387_),
    .A_N(_0701_));
 sg13g2_a21oi_1 _2484_ (.A1(_0439_),
    .A2(_0388_),
    .Y(_0389_),
    .B1(_0382_));
 sg13g2_nor2_1 _2485_ (.A(_1125_),
    .B(net63),
    .Y(_0390_));
 sg13g2_a21oi_1 _2486_ (.A1(net83),
    .A2(_0390_),
    .Y(_0391_),
    .B1(_0013_));
 sg13g2_o21ai_1 _2487_ (.B1(net73),
    .Y(_0392_),
    .A1(net86),
    .A2(_0391_));
 sg13g2_nor4_1 _2488_ (.A(_0701_),
    .B(_0671_),
    .C(_0397_),
    .D(_0447_),
    .Y(_0393_));
 sg13g2_nand3_1 _2489_ (.B(_1126_),
    .C(_0393_),
    .A(_0439_),
    .Y(_0394_));
 sg13g2_o21ai_1 _2490_ (.B1(net83),
    .Y(_0395_),
    .A1(_0458_),
    .A2(net63));
 sg13g2_nand3_1 _2491_ (.B(_0408_),
    .C(_0395_),
    .A(_0386_),
    .Y(_0396_));
 sg13g2_nor2_1 _2492_ (.A(_0298_),
    .B(_0778_),
    .Y(_0398_));
 sg13g2_nand4_1 _2493_ (.B(_0394_),
    .C(_0396_),
    .A(_0392_),
    .Y(_0399_),
    .D(_0398_));
 sg13g2_a21oi_1 _2494_ (.A1(_0768_),
    .A2(_0387_),
    .Y(_0400_),
    .B1(net73));
 sg13g2_nand2_1 _2495_ (.Y(_0401_),
    .A(net73),
    .B(_0387_));
 sg13g2_a21oi_1 _2496_ (.A1(_0458_),
    .A2(net63),
    .Y(_0402_),
    .B1(_0401_));
 sg13g2_nor3_1 _2497_ (.A(_0309_),
    .B(_0435_),
    .C(_0522_),
    .Y(_0403_));
 sg13g2_o21ai_1 _2498_ (.B1(_0403_),
    .Y(_0404_),
    .A1(_0400_),
    .A2(_0402_));
 sg13g2_nand3b_1 _2499_ (.B(_0399_),
    .C(_0404_),
    .Y(_0405_),
    .A_N(_0389_));
 sg13g2_a22oi_1 _2500_ (.Y(_0406_),
    .B1(_0385_),
    .B2(_0405_),
    .A2(_0379_),
    .A1(_0373_));
 sg13g2_nand2_1 _2501_ (.Y(_0407_),
    .A(_0350_),
    .B(_0349_));
 sg13g2_nand4_1 _2502_ (.B(_0058_),
    .C(_0075_),
    .A(_1205_),
    .Y(_0409_),
    .D(_0407_));
 sg13g2_a221oi_1 _2503_ (.B2(_0399_),
    .C1(_0360_),
    .B1(_0385_),
    .A1(_0354_),
    .Y(_0410_),
    .A2(_0377_));
 sg13g2_a21oi_1 _2504_ (.A1(_0379_),
    .A2(_0409_),
    .Y(_0411_),
    .B1(_0410_));
 sg13g2_nand2b_1 _2505_ (.Y(_0412_),
    .B(_0411_),
    .A_N(_0406_));
 sg13g2_inv_1 _2506_ (.Y(_0413_),
    .A(_0412_));
 sg13g2_o21ai_1 _2507_ (.B1(_0413_),
    .Y(_0414_),
    .A1(_0077_),
    .A2(_0367_));
 sg13g2_o21ai_1 _2508_ (.B1(_0298_),
    .Y(_0415_),
    .A1(_0435_),
    .A2(_0444_));
 sg13g2_nand3_1 _2509_ (.B(_0156_),
    .C(_0415_),
    .A(_0714_),
    .Y(_0416_));
 sg13g2_a21oi_1 _2510_ (.A1(_0373_),
    .A2(_0377_),
    .Y(_0417_),
    .B1(_0343_));
 sg13g2_a21oi_1 _2511_ (.A1(_0385_),
    .A2(_0389_),
    .Y(_0418_),
    .B1(_0360_));
 sg13g2_nand2b_1 _2512_ (.Y(_0420_),
    .B(_0418_),
    .A_N(_0417_));
 sg13g2_inv_1 _2513_ (.Y(_0421_),
    .A(_0872_));
 sg13g2_a221oi_1 _2514_ (.B2(_0081_),
    .C1(_0421_),
    .B1(_0420_),
    .A1(_0133_),
    .Y(_0422_),
    .A2(_0333_));
 sg13g2_buf_2 _2515_ (.A(_0422_),
    .X(_0423_));
 sg13g2_nor2_1 _2516_ (.A(_0416_),
    .B(_0423_),
    .Y(_0424_));
 sg13g2_inv_1 _2517_ (.Y(_0425_),
    .A(_0411_));
 sg13g2_nand2_1 _2518_ (.Y(_0426_),
    .A(_0406_),
    .B(_0425_));
 sg13g2_and3_1 _2519_ (.X(net15),
    .A(_0414_),
    .B(_0424_),
    .C(_0426_));
 sg13g2_o21ai_1 _2520_ (.B1(_0412_),
    .Y(_0427_),
    .A1(_0077_),
    .A2(_0367_));
 sg13g2_and2_1 _2521_ (.A(_0424_),
    .B(_0427_),
    .X(net16));
 sg13g2_nand2b_1 _2522_ (.Y(_0429_),
    .B(_0406_),
    .A_N(_0423_));
 sg13g2_nand2b_1 _2523_ (.Y(_0430_),
    .B(_0411_),
    .A_N(_0365_));
 sg13g2_a21oi_1 _2524_ (.A1(_0429_),
    .A2(_0430_),
    .Y(net17),
    .B1(_0416_));
 sg13g2_or3_1 _2525_ (.A(_0077_),
    .B(_0367_),
    .C(_0416_),
    .X(_0431_));
 sg13g2_xor2_1 _2526_ (.B(_0423_),
    .A(_0406_),
    .X(_0432_));
 sg13g2_nor3_1 _2527_ (.A(_0425_),
    .B(_0431_),
    .C(_0432_),
    .Y(net19));
 sg13g2_nor2_1 _2528_ (.A(_0412_),
    .B(_0431_),
    .Y(net20));
 sg13g2_mux2_1 _2529_ (.A0(_0412_),
    .A1(_0426_),
    .S(_0423_),
    .X(_0433_));
 sg13g2_nor2_1 _2530_ (.A(_0431_),
    .B(_0433_),
    .Y(net21));
 sg13g2_buf_1 clkbuf_0_clk (.A(clk),
    .X(clknet_0_clk));
 sg13g2_buf_1 _2532_ (.A(net93),
    .X(uio_oe[0]));
 sg13g2_buf_1 _2533_ (.A(net94),
    .X(uio_oe[1]));
 sg13g2_buf_1 _2534_ (.A(net95),
    .X(uio_oe[2]));
 sg13g2_buf_1 _2535_ (.A(net96),
    .X(uio_oe[3]));
 sg13g2_buf_1 _2536_ (.A(net97),
    .X(uio_oe[4]));
 sg13g2_buf_1 _2537_ (.A(net98),
    .X(uio_oe[5]));
 sg13g2_buf_1 _2538_ (.A(net99),
    .X(uio_oe[6]));
 sg13g2_buf_1 _2539_ (.A(net100),
    .X(uio_oe[7]));
 sg13g2_buf_1 _2540_ (.A(net92),
    .X(net18));
 sg13g2_buf_1 _2541_ (.A(hsync),
    .X(net22));
 sg13g2_dfrbp_1 \counter[0]$_SDFF_PN0_  (.CLK(net91),
    .RESET_B(net101),
    .D(_0019_),
    .Q_N(_0010_),
    .Q(\counter[0] ));
 sg13g2_dfrbp_1 \counter[1]$_SDFF_PN0_  (.CLK(net91),
    .RESET_B(net102),
    .D(_0020_),
    .Q_N(_1272_),
    .Q(\counter[1] ));
 sg13g2_dfrbp_1 \counter[2]$_SDFF_PN0_  (.CLK(net91),
    .RESET_B(net103),
    .D(_0021_),
    .Q_N(_0007_),
    .Q(\counter[2] ));
 sg13g2_dfrbp_1 \counter[3]$_SDFF_PN0_  (.CLK(net92),
    .RESET_B(net104),
    .D(_0022_),
    .Q_N(_1271_),
    .Q(\counter[3] ));
 sg13g2_dfrbp_1 \counter[4]$_SDFF_PN0_  (.CLK(net91),
    .RESET_B(net105),
    .D(_0023_),
    .Q_N(_1270_),
    .Q(\counter[4] ));
 sg13g2_dfrbp_1 \counter[5]$_SDFF_PN0_  (.CLK(net91),
    .RESET_B(net106),
    .D(_0024_),
    .Q_N(_1269_),
    .Q(\counter[5] ));
 sg13g2_dfrbp_1 \counter[6]$_SDFF_PN0_  (.CLK(net91),
    .RESET_B(net107),
    .D(_0025_),
    .Q_N(_1268_),
    .Q(\counter[6] ));
 sg13g2_dfrbp_1 \counter[7]$_SDFF_PN0_  (.CLK(net91),
    .RESET_B(net108),
    .D(_0026_),
    .Q_N(_0008_),
    .Q(\counter[7] ));
 sg13g2_dfrbp_1 \counter[8]$_SDFF_PN0_  (.CLK(net91),
    .RESET_B(net109),
    .D(_0027_),
    .Q_N(_0009_),
    .Q(\counter[8] ));
 sg13g2_dfrbp_1 \counter[9]$_SDFF_PN0_  (.CLK(net92),
    .RESET_B(net110),
    .D(_0028_),
    .Q_N(_1267_),
    .Q(\counter[9] ));
 sg13g2_dfrbp_1 \hvsync_gen.hpos[0]$_SDFF_PP0_  (.CLK(clknet_2_0__leaf_clk),
    .RESET_B(net111),
    .D(_0029_),
    .Q_N(_0017_),
    .Q(\hvsync_gen.hpos[0] ));
 sg13g2_dfrbp_1 \hvsync_gen.hpos[1]$_SDFF_PP0_  (.CLK(clknet_2_1__leaf_clk),
    .RESET_B(net112),
    .D(_0030_),
    .Q_N(_0016_),
    .Q(\hvsync_gen.hpos[1] ));
 sg13g2_dfrbp_1 \hvsync_gen.hpos[2]$_SDFF_PP0_  (.CLK(clknet_2_0__leaf_clk),
    .RESET_B(net113),
    .D(_0031_),
    .Q_N(_0014_),
    .Q(\hvsync_gen.hpos[2] ));
 sg13g2_dfrbp_1 \hvsync_gen.hpos[3]$_SDFF_PP0_  (.CLK(clknet_2_2__leaf_clk),
    .RESET_B(net114),
    .D(_0032_),
    .Q_N(_0013_),
    .Q(\hvsync_gen.hpos[3] ));
 sg13g2_dfrbp_1 \hvsync_gen.hpos[4]$_SDFF_PP0_  (.CLK(clknet_2_2__leaf_clk),
    .RESET_B(net115),
    .D(_0033_),
    .Q_N(_0012_),
    .Q(\hvsync_gen.hpos[4] ));
 sg13g2_dfrbp_1 \hvsync_gen.hpos[5]$_SDFF_PP0_  (.CLK(clknet_2_2__leaf_clk),
    .RESET_B(net116),
    .D(_0034_),
    .Q_N(_1266_),
    .Q(\hvsync_gen.hpos[5] ));
 sg13g2_dfrbp_1 \hvsync_gen.hpos[6]$_SDFF_PP0_  (.CLK(clknet_2_2__leaf_clk),
    .RESET_B(net117),
    .D(_0035_),
    .Q_N(_0011_),
    .Q(\hvsync_gen.hpos[6] ));
 sg13g2_dfrbp_1 \hvsync_gen.hpos[7]$_SDFF_PP0_  (.CLK(clknet_2_2__leaf_clk),
    .RESET_B(net118),
    .D(_0036_),
    .Q_N(_0015_),
    .Q(\hvsync_gen.hpos[7] ));
 sg13g2_dfrbp_1 \hvsync_gen.hpos[8]$_SDFF_PP0_  (.CLK(clknet_2_3__leaf_clk),
    .RESET_B(net119),
    .D(_0037_),
    .Q_N(_1265_),
    .Q(\hvsync_gen.hpos[8] ));
 sg13g2_dfrbp_1 \hvsync_gen.hpos[9]$_SDFF_PP0_  (.CLK(clknet_2_2__leaf_clk),
    .RESET_B(net120),
    .D(_0038_),
    .Q_N(_0006_),
    .Q(\hvsync_gen.hpos[9] ));
 sg13g2_dfrbp_1 \hvsync_gen.hsync$_DFF_P_  (.CLK(clknet_2_3__leaf_clk),
    .RESET_B(net121),
    .D(_0000_),
    .Q_N(_1264_),
    .Q(hsync));
 sg13g2_dfrbp_1 \hvsync_gen.vpos[0]$_SDFFCE_PP0P_  (.CLK(clknet_2_3__leaf_clk),
    .RESET_B(net122),
    .D(_0039_),
    .Q_N(_0018_),
    .Q(\hvsync_gen.vpos[0] ));
 sg13g2_dfrbp_1 \hvsync_gen.vpos[1]$_SDFFCE_PP0P_  (.CLK(clknet_2_3__leaf_clk),
    .RESET_B(net123),
    .D(_0040_),
    .Q_N(_0005_),
    .Q(\hvsync_gen.vpos[1] ));
 sg13g2_dfrbp_1 \hvsync_gen.vpos[2]$_SDFFCE_PP0P_  (.CLK(clknet_2_1__leaf_clk),
    .RESET_B(net124),
    .D(_0041_),
    .Q_N(_0004_),
    .Q(\hvsync_gen.vpos[2] ));
 sg13g2_dfrbp_1 \hvsync_gen.vpos[3]$_SDFFCE_PP0P_  (.CLK(clknet_2_1__leaf_clk),
    .RESET_B(net125),
    .D(_0042_),
    .Q_N(_1263_),
    .Q(\hvsync_gen.vpos[3] ));
 sg13g2_dfrbp_1 \hvsync_gen.vpos[4]$_SDFFCE_PP0P_  (.CLK(clknet_2_0__leaf_clk),
    .RESET_B(net126),
    .D(_0043_),
    .Q_N(_1262_),
    .Q(\hvsync_gen.vpos[4] ));
 sg13g2_dfrbp_1 \hvsync_gen.vpos[5]$_SDFFCE_PP0P_  (.CLK(clknet_2_0__leaf_clk),
    .RESET_B(net127),
    .D(_0044_),
    .Q_N(_0003_),
    .Q(\hvsync_gen.vpos[5] ));
 sg13g2_dfrbp_1 \hvsync_gen.vpos[6]$_SDFFCE_PP0P_  (.CLK(clknet_2_0__leaf_clk),
    .RESET_B(net128),
    .D(_0045_),
    .Q_N(_1261_),
    .Q(\hvsync_gen.vpos[6] ));
 sg13g2_dfrbp_1 \hvsync_gen.vpos[7]$_SDFFCE_PP0P_  (.CLK(clknet_2_1__leaf_clk),
    .RESET_B(net129),
    .D(_0046_),
    .Q_N(_1260_),
    .Q(\hvsync_gen.vpos[7] ));
 sg13g2_dfrbp_1 \hvsync_gen.vpos[8]$_SDFFCE_PP0P_  (.CLK(clknet_2_0__leaf_clk),
    .RESET_B(net130),
    .D(_0047_),
    .Q_N(_0002_),
    .Q(\hvsync_gen.vpos[8] ));
 sg13g2_dfrbp_1 \hvsync_gen.vpos[9]$_SDFFCE_PP0P_  (.CLK(clknet_2_1__leaf_clk),
    .RESET_B(net131),
    .D(_0048_),
    .Q_N(_1273_),
    .Q(\hvsync_gen.vpos[9] ));
 sg13g2_dfrbp_1 \hvsync_gen.vsync$_DFF_P_  (.CLK(clknet_2_3__leaf_clk),
    .RESET_B(net132),
    .D(_0001_),
    .Q_N(_1259_),
    .Q(\hvsync_gen.vsync ));
 sg13g2_buf_1 input1 (.A(ui_in[0]),
    .X(net1));
 sg13g2_buf_1 input2 (.A(ui_in[1]),
    .X(net2));
 sg13g2_buf_1 input3 (.A(ui_in[4]),
    .X(net3));
 sg13g2_buf_1 input4 (.A(ui_in[5]),
    .X(net4));
 sg13g2_buf_1 input5 (.A(ui_in[6]),
    .X(net5));
 sg13g2_buf_1 input6 (.A(ui_in[7]),
    .X(net6));
 sg13g2_buf_1 output7 (.A(net27),
    .X(uio_out[0]));
 sg13g2_buf_1 output8 (.A(net32),
    .X(uio_out[1]));
 sg13g2_buf_1 output9 (.A(net33),
    .X(uio_out[2]));
 sg13g2_buf_1 output10 (.A(net10),
    .X(uio_out[3]));
 sg13g2_buf_1 output11 (.A(net11),
    .X(uio_out[4]));
 sg13g2_buf_1 output12 (.A(net12),
    .X(uio_out[5]));
 sg13g2_buf_1 output13 (.A(net13),
    .X(uio_out[6]));
 sg13g2_buf_1 output14 (.A(net14),
    .X(uio_out[7]));
 sg13g2_buf_1 output15 (.A(net15),
    .X(uo_out[0]));
 sg13g2_buf_1 output16 (.A(net16),
    .X(uo_out[1]));
 sg13g2_buf_1 output17 (.A(net17),
    .X(uo_out[2]));
 sg13g2_buf_1 output18 (.A(net18),
    .X(uo_out[3]));
 sg13g2_buf_1 output19 (.A(net19),
    .X(uo_out[4]));
 sg13g2_buf_1 output20 (.A(net20),
    .X(uo_out[5]));
 sg13g2_buf_1 output21 (.A(net21),
    .X(uo_out[6]));
 sg13g2_buf_1 output22 (.A(net22),
    .X(uo_out[7]));
 sg13g2_buf_2 fanout23 (.A(net12),
    .X(net23));
 sg13g2_buf_2 fanout24 (.A(_1078_),
    .X(net24));
 sg13g2_buf_2 fanout25 (.A(_0139_),
    .X(net25));
 sg13g2_buf_2 fanout26 (.A(net13),
    .X(net26));
 sg13g2_buf_2 fanout27 (.A(net7),
    .X(net27));
 sg13g2_buf_2 fanout28 (.A(net10),
    .X(net28));
 sg13g2_buf_2 fanout29 (.A(_0158_),
    .X(net29));
 sg13g2_buf_2 fanout30 (.A(_0144_),
    .X(net30));
 sg13g2_buf_2 fanout31 (.A(_1059_),
    .X(net31));
 sg13g2_buf_2 fanout32 (.A(net8),
    .X(net32));
 sg13g2_buf_2 fanout33 (.A(net9),
    .X(net33));
 sg13g2_buf_2 fanout34 (.A(_0143_),
    .X(net34));
 sg13g2_buf_2 fanout35 (.A(_0111_),
    .X(net35));
 sg13g2_buf_2 fanout36 (.A(_1039_),
    .X(net36));
 sg13g2_buf_2 fanout37 (.A(_1057_),
    .X(net37));
 sg13g2_buf_2 fanout38 (.A(_1028_),
    .X(net38));
 sg13g2_buf_2 fanout39 (.A(_0669_),
    .X(net39));
 sg13g2_buf_2 fanout40 (.A(_1191_),
    .X(net40));
 sg13g2_buf_2 fanout41 (.A(_0548_),
    .X(net41));
 sg13g2_buf_2 fanout42 (.A(_0547_),
    .X(net42));
 sg13g2_buf_2 fanout43 (.A(_0617_),
    .X(net43));
 sg13g2_buf_2 fanout44 (.A(_0613_),
    .X(net44));
 sg13g2_buf_2 fanout45 (.A(_0082_),
    .X(net45));
 sg13g2_buf_2 fanout46 (.A(_1175_),
    .X(net46));
 sg13g2_buf_2 fanout47 (.A(_1182_),
    .X(net47));
 sg13g2_buf_2 fanout48 (.A(_0722_),
    .X(net48));
 sg13g2_buf_2 fanout49 (.A(_0887_),
    .X(net49));
 sg13g2_buf_2 fanout50 (.A(_0720_),
    .X(net50));
 sg13g2_buf_2 fanout51 (.A(_0913_),
    .X(net51));
 sg13g2_buf_2 fanout52 (.A(_0790_),
    .X(net52));
 sg13g2_buf_2 fanout53 (.A(_0786_),
    .X(net53));
 sg13g2_buf_2 fanout54 (.A(_0717_),
    .X(net54));
 sg13g2_buf_2 fanout55 (.A(_0791_),
    .X(net55));
 sg13g2_buf_2 fanout56 (.A(_0731_),
    .X(net56));
 sg13g2_buf_2 fanout57 (.A(_0549_),
    .X(net57));
 sg13g2_buf_2 fanout58 (.A(_0435_),
    .X(net58));
 sg13g2_buf_2 fanout59 (.A(_0266_),
    .X(net59));
 sg13g2_buf_2 fanout60 (.A(_0766_),
    .X(net60));
 sg13g2_buf_2 fanout61 (.A(_0729_),
    .X(net61));
 sg13g2_buf_2 fanout62 (.A(_0724_),
    .X(net62));
 sg13g2_buf_2 fanout63 (.A(_0701_),
    .X(net63));
 sg13g2_buf_2 fanout64 (.A(_0631_),
    .X(net64));
 sg13g2_buf_2 fanout65 (.A(_0500_),
    .X(net65));
 sg13g2_buf_2 fanout66 (.A(_0485_),
    .X(net66));
 sg13g2_buf_2 fanout67 (.A(_0471_),
    .X(net67));
 sg13g2_buf_2 fanout68 (.A(_0469_),
    .X(net68));
 sg13g2_buf_2 fanout69 (.A(_0461_),
    .X(net69));
 sg13g2_buf_2 fanout70 (.A(_0460_),
    .X(net70));
 sg13g2_buf_2 fanout71 (.A(_0455_),
    .X(net71));
 sg13g2_buf_2 fanout72 (.A(_0449_),
    .X(net72));
 sg13g2_buf_2 fanout73 (.A(_0437_),
    .X(net73));
 sg13g2_buf_2 fanout74 (.A(_0434_),
    .X(net74));
 sg13g2_buf_2 fanout75 (.A(_0353_),
    .X(net75));
 sg13g2_buf_2 fanout76 (.A(_0331_),
    .X(net76));
 sg13g2_buf_2 fanout77 (.A(_0222_),
    .X(net77));
 sg13g2_buf_2 fanout78 (.A(_0178_),
    .X(net78));
 sg13g2_buf_2 fanout79 (.A(_0134_),
    .X(net79));
 sg13g2_buf_2 fanout80 (.A(_0101_),
    .X(net80));
 sg13g2_buf_2 fanout81 (.A(_1114_),
    .X(net81));
 sg13g2_buf_2 fanout82 (.A(_0846_),
    .X(net82));
 sg13g2_buf_2 fanout83 (.A(_0466_),
    .X(net83));
 sg13g2_buf_2 fanout84 (.A(_0446_),
    .X(net84));
 sg13g2_buf_2 fanout85 (.A(_0443_),
    .X(net85));
 sg13g2_buf_2 fanout86 (.A(_0397_),
    .X(net86));
 sg13g2_buf_2 fanout87 (.A(_0189_),
    .X(net87));
 sg13g2_buf_2 fanout88 (.A(_0145_),
    .X(net88));
 sg13g2_buf_2 fanout89 (.A(_0112_),
    .X(net89));
 sg13g2_buf_2 fanout90 (.A(_0079_),
    .X(net90));
 sg13g2_buf_2 fanout91 (.A(net92),
    .X(net91));
 sg13g2_buf_1 fanout92 (.A(\hvsync_gen.vsync ),
    .X(net92));
 sg13g2_tiehi _2532__93 (.L_HI(net93));
 sg13g2_tiehi _2533__94 (.L_HI(net94));
 sg13g2_tiehi _2534__95 (.L_HI(net95));
 sg13g2_tiehi _2535__96 (.L_HI(net96));
 sg13g2_tiehi _2536__97 (.L_HI(net97));
 sg13g2_tiehi _2537__98 (.L_HI(net98));
 sg13g2_tiehi _2538__99 (.L_HI(net99));
 sg13g2_tiehi _2539__100 (.L_HI(net100));
 sg13g2_tiehi \counter[0]$_SDFF_PN0__101  (.L_HI(net101));
 sg13g2_tiehi \counter[1]$_SDFF_PN0__102  (.L_HI(net102));
 sg13g2_tiehi \counter[2]$_SDFF_PN0__103  (.L_HI(net103));
 sg13g2_tiehi \counter[3]$_SDFF_PN0__104  (.L_HI(net104));
 sg13g2_tiehi \counter[4]$_SDFF_PN0__105  (.L_HI(net105));
 sg13g2_tiehi \counter[5]$_SDFF_PN0__106  (.L_HI(net106));
 sg13g2_tiehi \counter[6]$_SDFF_PN0__107  (.L_HI(net107));
 sg13g2_tiehi \counter[7]$_SDFF_PN0__108  (.L_HI(net108));
 sg13g2_tiehi \counter[8]$_SDFF_PN0__109  (.L_HI(net109));
 sg13g2_tiehi \counter[9]$_SDFF_PN0__110  (.L_HI(net110));
 sg13g2_tiehi \hvsync_gen.hpos[0]$_SDFF_PP0__111  (.L_HI(net111));
 sg13g2_tiehi \hvsync_gen.hpos[1]$_SDFF_PP0__112  (.L_HI(net112));
 sg13g2_tiehi \hvsync_gen.hpos[2]$_SDFF_PP0__113  (.L_HI(net113));
 sg13g2_tiehi \hvsync_gen.hpos[3]$_SDFF_PP0__114  (.L_HI(net114));
 sg13g2_tiehi \hvsync_gen.hpos[4]$_SDFF_PP0__115  (.L_HI(net115));
 sg13g2_tiehi \hvsync_gen.hpos[5]$_SDFF_PP0__116  (.L_HI(net116));
 sg13g2_tiehi \hvsync_gen.hpos[6]$_SDFF_PP0__117  (.L_HI(net117));
 sg13g2_tiehi \hvsync_gen.hpos[7]$_SDFF_PP0__118  (.L_HI(net118));
 sg13g2_tiehi \hvsync_gen.hpos[8]$_SDFF_PP0__119  (.L_HI(net119));
 sg13g2_tiehi \hvsync_gen.hpos[9]$_SDFF_PP0__120  (.L_HI(net120));
 sg13g2_tiehi \hvsync_gen.hsync$_DFF_P__121  (.L_HI(net121));
 sg13g2_tiehi \hvsync_gen.vpos[0]$_SDFFCE_PP0P__122  (.L_HI(net122));
 sg13g2_tiehi \hvsync_gen.vpos[1]$_SDFFCE_PP0P__123  (.L_HI(net123));
 sg13g2_tiehi \hvsync_gen.vpos[2]$_SDFFCE_PP0P__124  (.L_HI(net124));
 sg13g2_tiehi \hvsync_gen.vpos[3]$_SDFFCE_PP0P__125  (.L_HI(net125));
 sg13g2_tiehi \hvsync_gen.vpos[4]$_SDFFCE_PP0P__126  (.L_HI(net126));
 sg13g2_tiehi \hvsync_gen.vpos[5]$_SDFFCE_PP0P__127  (.L_HI(net127));
 sg13g2_tiehi \hvsync_gen.vpos[6]$_SDFFCE_PP0P__128  (.L_HI(net128));
 sg13g2_tiehi \hvsync_gen.vpos[7]$_SDFFCE_PP0P__129  (.L_HI(net129));
 sg13g2_tiehi \hvsync_gen.vpos[8]$_SDFFCE_PP0P__130  (.L_HI(net130));
 sg13g2_tiehi \hvsync_gen.vpos[9]$_SDFFCE_PP0P__131  (.L_HI(net131));
 sg13g2_tiehi \hvsync_gen.vsync$_DFF_P__132  (.L_HI(net132));
 sg13g2_buf_1 clkbuf_2_0__f_clk (.A(clknet_0_clk),
    .X(clknet_2_0__leaf_clk));
 sg13g2_buf_1 clkbuf_2_1__f_clk (.A(clknet_0_clk),
    .X(clknet_2_1__leaf_clk));
 sg13g2_buf_1 clkbuf_2_2__f_clk (.A(clknet_0_clk),
    .X(clknet_2_2__leaf_clk));
 sg13g2_buf_1 clkbuf_2_3__f_clk (.A(clknet_0_clk),
    .X(clknet_2_3__leaf_clk));
 sg13g2_inv_1 clkload0 (.A(clknet_2_1__leaf_clk));
 sg13g2_inv_1 clkload1 (.A(clknet_2_3__leaf_clk));
 sg13g2_decap_8 FILLER_0_0 ();
 sg13g2_decap_8 FILLER_0_7 ();
 sg13g2_decap_8 FILLER_0_14 ();
 sg13g2_decap_8 FILLER_0_21 ();
 sg13g2_decap_8 FILLER_0_28 ();
 sg13g2_decap_8 FILLER_0_35 ();
 sg13g2_decap_8 FILLER_0_42 ();
 sg13g2_decap_8 FILLER_0_49 ();
 sg13g2_decap_8 FILLER_0_56 ();
 sg13g2_decap_8 FILLER_0_63 ();
 sg13g2_decap_8 FILLER_0_70 ();
 sg13g2_decap_8 FILLER_0_77 ();
 sg13g2_decap_8 FILLER_0_84 ();
 sg13g2_decap_8 FILLER_0_91 ();
 sg13g2_decap_8 FILLER_0_98 ();
 sg13g2_decap_8 FILLER_0_105 ();
 sg13g2_decap_8 FILLER_0_112 ();
 sg13g2_decap_8 FILLER_0_119 ();
 sg13g2_decap_8 FILLER_0_126 ();
 sg13g2_decap_8 FILLER_0_133 ();
 sg13g2_decap_8 FILLER_0_140 ();
 sg13g2_decap_8 FILLER_0_147 ();
 sg13g2_decap_8 FILLER_0_154 ();
 sg13g2_decap_8 FILLER_0_161 ();
 sg13g2_decap_8 FILLER_0_168 ();
 sg13g2_decap_8 FILLER_0_175 ();
 sg13g2_decap_8 FILLER_0_182 ();
 sg13g2_decap_8 FILLER_0_189 ();
 sg13g2_decap_8 FILLER_0_196 ();
 sg13g2_decap_8 FILLER_0_203 ();
 sg13g2_decap_8 FILLER_0_210 ();
 sg13g2_decap_8 FILLER_0_217 ();
 sg13g2_decap_8 FILLER_0_224 ();
 sg13g2_decap_8 FILLER_0_231 ();
 sg13g2_decap_8 FILLER_0_238 ();
 sg13g2_decap_8 FILLER_0_245 ();
 sg13g2_decap_8 FILLER_0_252 ();
 sg13g2_decap_8 FILLER_0_259 ();
 sg13g2_decap_8 FILLER_0_266 ();
 sg13g2_decap_8 FILLER_0_273 ();
 sg13g2_decap_8 FILLER_0_280 ();
 sg13g2_decap_8 FILLER_0_287 ();
 sg13g2_decap_8 FILLER_0_294 ();
 sg13g2_decap_8 FILLER_0_301 ();
 sg13g2_decap_8 FILLER_0_308 ();
 sg13g2_decap_8 FILLER_0_315 ();
 sg13g2_decap_8 FILLER_0_322 ();
 sg13g2_decap_8 FILLER_0_329 ();
 sg13g2_decap_8 FILLER_0_336 ();
 sg13g2_decap_8 FILLER_0_343 ();
 sg13g2_decap_8 FILLER_0_350 ();
 sg13g2_decap_8 FILLER_0_357 ();
 sg13g2_decap_8 FILLER_0_364 ();
 sg13g2_decap_8 FILLER_0_371 ();
 sg13g2_decap_8 FILLER_0_378 ();
 sg13g2_decap_8 FILLER_0_385 ();
 sg13g2_decap_8 FILLER_0_392 ();
 sg13g2_decap_8 FILLER_0_399 ();
 sg13g2_decap_8 FILLER_0_406 ();
 sg13g2_decap_8 FILLER_0_413 ();
 sg13g2_decap_8 FILLER_0_420 ();
 sg13g2_fill_2 FILLER_0_427 ();
 sg13g2_fill_1 FILLER_0_429 ();
 sg13g2_decap_8 FILLER_1_0 ();
 sg13g2_decap_8 FILLER_1_7 ();
 sg13g2_decap_8 FILLER_1_14 ();
 sg13g2_decap_8 FILLER_1_21 ();
 sg13g2_decap_8 FILLER_1_28 ();
 sg13g2_decap_8 FILLER_1_35 ();
 sg13g2_decap_8 FILLER_1_42 ();
 sg13g2_decap_8 FILLER_1_49 ();
 sg13g2_decap_8 FILLER_1_56 ();
 sg13g2_decap_8 FILLER_1_63 ();
 sg13g2_decap_8 FILLER_1_70 ();
 sg13g2_decap_8 FILLER_1_77 ();
 sg13g2_decap_8 FILLER_1_84 ();
 sg13g2_decap_8 FILLER_1_91 ();
 sg13g2_decap_8 FILLER_1_98 ();
 sg13g2_decap_8 FILLER_1_105 ();
 sg13g2_decap_8 FILLER_1_112 ();
 sg13g2_decap_8 FILLER_1_119 ();
 sg13g2_decap_8 FILLER_1_126 ();
 sg13g2_decap_8 FILLER_1_133 ();
 sg13g2_decap_8 FILLER_1_140 ();
 sg13g2_decap_8 FILLER_1_147 ();
 sg13g2_decap_8 FILLER_1_154 ();
 sg13g2_decap_8 FILLER_1_161 ();
 sg13g2_decap_8 FILLER_1_168 ();
 sg13g2_decap_8 FILLER_1_175 ();
 sg13g2_decap_8 FILLER_1_182 ();
 sg13g2_decap_8 FILLER_1_189 ();
 sg13g2_decap_8 FILLER_1_196 ();
 sg13g2_decap_8 FILLER_1_203 ();
 sg13g2_decap_8 FILLER_1_210 ();
 sg13g2_decap_8 FILLER_1_217 ();
 sg13g2_decap_8 FILLER_1_224 ();
 sg13g2_decap_8 FILLER_1_231 ();
 sg13g2_decap_8 FILLER_1_238 ();
 sg13g2_decap_8 FILLER_1_245 ();
 sg13g2_decap_8 FILLER_1_252 ();
 sg13g2_decap_8 FILLER_1_259 ();
 sg13g2_decap_8 FILLER_1_266 ();
 sg13g2_decap_8 FILLER_1_273 ();
 sg13g2_decap_8 FILLER_1_280 ();
 sg13g2_decap_8 FILLER_1_287 ();
 sg13g2_decap_8 FILLER_1_294 ();
 sg13g2_decap_8 FILLER_1_301 ();
 sg13g2_decap_8 FILLER_1_308 ();
 sg13g2_decap_8 FILLER_1_315 ();
 sg13g2_decap_8 FILLER_1_322 ();
 sg13g2_decap_8 FILLER_1_329 ();
 sg13g2_decap_8 FILLER_1_336 ();
 sg13g2_decap_8 FILLER_1_343 ();
 sg13g2_decap_8 FILLER_1_350 ();
 sg13g2_decap_8 FILLER_1_357 ();
 sg13g2_decap_8 FILLER_1_364 ();
 sg13g2_decap_8 FILLER_1_371 ();
 sg13g2_decap_8 FILLER_1_378 ();
 sg13g2_decap_8 FILLER_1_385 ();
 sg13g2_decap_8 FILLER_1_392 ();
 sg13g2_decap_8 FILLER_1_399 ();
 sg13g2_decap_8 FILLER_1_406 ();
 sg13g2_decap_8 FILLER_1_413 ();
 sg13g2_decap_8 FILLER_1_420 ();
 sg13g2_fill_2 FILLER_1_427 ();
 sg13g2_fill_1 FILLER_1_429 ();
 sg13g2_decap_8 FILLER_2_0 ();
 sg13g2_decap_8 FILLER_2_7 ();
 sg13g2_decap_8 FILLER_2_14 ();
 sg13g2_decap_8 FILLER_2_21 ();
 sg13g2_decap_8 FILLER_2_28 ();
 sg13g2_decap_8 FILLER_2_35 ();
 sg13g2_decap_8 FILLER_2_42 ();
 sg13g2_decap_8 FILLER_2_49 ();
 sg13g2_decap_8 FILLER_2_56 ();
 sg13g2_decap_8 FILLER_2_63 ();
 sg13g2_decap_8 FILLER_2_70 ();
 sg13g2_decap_8 FILLER_2_77 ();
 sg13g2_decap_8 FILLER_2_84 ();
 sg13g2_decap_8 FILLER_2_91 ();
 sg13g2_decap_8 FILLER_2_98 ();
 sg13g2_decap_8 FILLER_2_105 ();
 sg13g2_decap_8 FILLER_2_112 ();
 sg13g2_decap_8 FILLER_2_119 ();
 sg13g2_decap_8 FILLER_2_126 ();
 sg13g2_decap_8 FILLER_2_133 ();
 sg13g2_decap_8 FILLER_2_140 ();
 sg13g2_decap_8 FILLER_2_147 ();
 sg13g2_decap_8 FILLER_2_154 ();
 sg13g2_decap_8 FILLER_2_161 ();
 sg13g2_decap_8 FILLER_2_168 ();
 sg13g2_decap_8 FILLER_2_175 ();
 sg13g2_decap_8 FILLER_2_182 ();
 sg13g2_decap_8 FILLER_2_189 ();
 sg13g2_decap_8 FILLER_2_196 ();
 sg13g2_decap_8 FILLER_2_203 ();
 sg13g2_decap_8 FILLER_2_210 ();
 sg13g2_decap_8 FILLER_2_217 ();
 sg13g2_decap_8 FILLER_2_224 ();
 sg13g2_decap_8 FILLER_2_231 ();
 sg13g2_decap_8 FILLER_2_238 ();
 sg13g2_decap_8 FILLER_2_245 ();
 sg13g2_decap_8 FILLER_2_252 ();
 sg13g2_decap_8 FILLER_2_259 ();
 sg13g2_decap_8 FILLER_2_266 ();
 sg13g2_decap_8 FILLER_2_273 ();
 sg13g2_decap_8 FILLER_2_280 ();
 sg13g2_decap_8 FILLER_2_287 ();
 sg13g2_decap_8 FILLER_2_294 ();
 sg13g2_decap_8 FILLER_2_301 ();
 sg13g2_decap_8 FILLER_2_308 ();
 sg13g2_decap_8 FILLER_2_315 ();
 sg13g2_decap_8 FILLER_2_322 ();
 sg13g2_decap_8 FILLER_2_329 ();
 sg13g2_decap_8 FILLER_2_336 ();
 sg13g2_decap_8 FILLER_2_343 ();
 sg13g2_decap_8 FILLER_2_350 ();
 sg13g2_decap_8 FILLER_2_357 ();
 sg13g2_decap_8 FILLER_2_364 ();
 sg13g2_decap_8 FILLER_2_371 ();
 sg13g2_decap_8 FILLER_2_378 ();
 sg13g2_decap_8 FILLER_2_385 ();
 sg13g2_decap_8 FILLER_2_392 ();
 sg13g2_decap_8 FILLER_2_399 ();
 sg13g2_decap_8 FILLER_2_406 ();
 sg13g2_decap_8 FILLER_2_413 ();
 sg13g2_decap_8 FILLER_2_420 ();
 sg13g2_fill_2 FILLER_2_427 ();
 sg13g2_fill_1 FILLER_2_429 ();
 sg13g2_decap_8 FILLER_3_0 ();
 sg13g2_decap_8 FILLER_3_7 ();
 sg13g2_decap_8 FILLER_3_14 ();
 sg13g2_decap_8 FILLER_3_21 ();
 sg13g2_decap_8 FILLER_3_28 ();
 sg13g2_decap_8 FILLER_3_35 ();
 sg13g2_decap_8 FILLER_3_42 ();
 sg13g2_decap_8 FILLER_3_49 ();
 sg13g2_decap_8 FILLER_3_56 ();
 sg13g2_decap_8 FILLER_3_63 ();
 sg13g2_decap_8 FILLER_3_70 ();
 sg13g2_decap_8 FILLER_3_77 ();
 sg13g2_decap_8 FILLER_3_84 ();
 sg13g2_decap_8 FILLER_3_91 ();
 sg13g2_decap_8 FILLER_3_98 ();
 sg13g2_decap_8 FILLER_3_105 ();
 sg13g2_decap_8 FILLER_3_112 ();
 sg13g2_decap_8 FILLER_3_119 ();
 sg13g2_decap_8 FILLER_3_126 ();
 sg13g2_decap_8 FILLER_3_133 ();
 sg13g2_decap_8 FILLER_3_140 ();
 sg13g2_decap_8 FILLER_3_147 ();
 sg13g2_decap_8 FILLER_3_154 ();
 sg13g2_decap_8 FILLER_3_161 ();
 sg13g2_decap_8 FILLER_3_168 ();
 sg13g2_decap_8 FILLER_3_175 ();
 sg13g2_decap_8 FILLER_3_182 ();
 sg13g2_decap_8 FILLER_3_189 ();
 sg13g2_decap_8 FILLER_3_196 ();
 sg13g2_decap_8 FILLER_3_203 ();
 sg13g2_decap_8 FILLER_3_210 ();
 sg13g2_decap_8 FILLER_3_217 ();
 sg13g2_decap_8 FILLER_3_224 ();
 sg13g2_decap_8 FILLER_3_231 ();
 sg13g2_decap_8 FILLER_3_238 ();
 sg13g2_decap_8 FILLER_3_245 ();
 sg13g2_decap_8 FILLER_3_252 ();
 sg13g2_decap_8 FILLER_3_259 ();
 sg13g2_decap_8 FILLER_3_266 ();
 sg13g2_decap_8 FILLER_3_273 ();
 sg13g2_decap_8 FILLER_3_280 ();
 sg13g2_decap_8 FILLER_3_287 ();
 sg13g2_decap_8 FILLER_3_294 ();
 sg13g2_decap_8 FILLER_3_301 ();
 sg13g2_decap_8 FILLER_3_308 ();
 sg13g2_decap_8 FILLER_3_315 ();
 sg13g2_decap_8 FILLER_3_330 ();
 sg13g2_decap_4 FILLER_3_344 ();
 sg13g2_fill_1 FILLER_3_348 ();
 sg13g2_decap_4 FILLER_3_354 ();
 sg13g2_fill_1 FILLER_3_358 ();
 sg13g2_decap_8 FILLER_3_363 ();
 sg13g2_decap_8 FILLER_3_370 ();
 sg13g2_decap_8 FILLER_3_377 ();
 sg13g2_decap_8 FILLER_3_384 ();
 sg13g2_decap_8 FILLER_3_391 ();
 sg13g2_decap_8 FILLER_3_398 ();
 sg13g2_decap_8 FILLER_3_405 ();
 sg13g2_decap_8 FILLER_3_412 ();
 sg13g2_decap_8 FILLER_3_419 ();
 sg13g2_decap_4 FILLER_3_426 ();
 sg13g2_decap_8 FILLER_4_0 ();
 sg13g2_decap_8 FILLER_4_7 ();
 sg13g2_decap_8 FILLER_4_14 ();
 sg13g2_decap_8 FILLER_4_21 ();
 sg13g2_decap_8 FILLER_4_28 ();
 sg13g2_decap_8 FILLER_4_35 ();
 sg13g2_decap_8 FILLER_4_42 ();
 sg13g2_decap_8 FILLER_4_49 ();
 sg13g2_decap_8 FILLER_4_56 ();
 sg13g2_decap_8 FILLER_4_63 ();
 sg13g2_decap_8 FILLER_4_70 ();
 sg13g2_decap_8 FILLER_4_77 ();
 sg13g2_decap_8 FILLER_4_84 ();
 sg13g2_decap_8 FILLER_4_91 ();
 sg13g2_decap_8 FILLER_4_98 ();
 sg13g2_decap_8 FILLER_4_105 ();
 sg13g2_decap_8 FILLER_4_112 ();
 sg13g2_decap_8 FILLER_4_119 ();
 sg13g2_decap_8 FILLER_4_126 ();
 sg13g2_decap_8 FILLER_4_133 ();
 sg13g2_decap_8 FILLER_4_140 ();
 sg13g2_decap_8 FILLER_4_147 ();
 sg13g2_decap_8 FILLER_4_154 ();
 sg13g2_decap_8 FILLER_4_161 ();
 sg13g2_decap_8 FILLER_4_168 ();
 sg13g2_decap_8 FILLER_4_175 ();
 sg13g2_decap_8 FILLER_4_182 ();
 sg13g2_decap_8 FILLER_4_189 ();
 sg13g2_decap_8 FILLER_4_196 ();
 sg13g2_decap_8 FILLER_4_203 ();
 sg13g2_decap_8 FILLER_4_210 ();
 sg13g2_decap_8 FILLER_4_217 ();
 sg13g2_decap_8 FILLER_4_224 ();
 sg13g2_decap_8 FILLER_4_231 ();
 sg13g2_decap_8 FILLER_4_238 ();
 sg13g2_decap_8 FILLER_4_245 ();
 sg13g2_decap_8 FILLER_4_252 ();
 sg13g2_decap_8 FILLER_4_259 ();
 sg13g2_decap_8 FILLER_4_266 ();
 sg13g2_decap_8 FILLER_4_273 ();
 sg13g2_decap_8 FILLER_4_280 ();
 sg13g2_decap_8 FILLER_4_287 ();
 sg13g2_fill_1 FILLER_4_294 ();
 sg13g2_fill_2 FILLER_4_323 ();
 sg13g2_decap_4 FILLER_4_370 ();
 sg13g2_fill_1 FILLER_4_374 ();
 sg13g2_decap_8 FILLER_4_380 ();
 sg13g2_decap_8 FILLER_4_413 ();
 sg13g2_decap_8 FILLER_4_420 ();
 sg13g2_fill_2 FILLER_4_427 ();
 sg13g2_fill_1 FILLER_4_429 ();
 sg13g2_decap_8 FILLER_5_0 ();
 sg13g2_decap_8 FILLER_5_7 ();
 sg13g2_decap_8 FILLER_5_14 ();
 sg13g2_decap_8 FILLER_5_21 ();
 sg13g2_decap_8 FILLER_5_28 ();
 sg13g2_decap_8 FILLER_5_35 ();
 sg13g2_decap_8 FILLER_5_42 ();
 sg13g2_decap_8 FILLER_5_49 ();
 sg13g2_decap_8 FILLER_5_56 ();
 sg13g2_decap_8 FILLER_5_63 ();
 sg13g2_decap_8 FILLER_5_70 ();
 sg13g2_decap_8 FILLER_5_77 ();
 sg13g2_decap_8 FILLER_5_84 ();
 sg13g2_decap_8 FILLER_5_91 ();
 sg13g2_decap_8 FILLER_5_98 ();
 sg13g2_decap_8 FILLER_5_105 ();
 sg13g2_decap_8 FILLER_5_112 ();
 sg13g2_decap_8 FILLER_5_119 ();
 sg13g2_decap_8 FILLER_5_126 ();
 sg13g2_decap_8 FILLER_5_133 ();
 sg13g2_decap_8 FILLER_5_140 ();
 sg13g2_decap_8 FILLER_5_147 ();
 sg13g2_decap_8 FILLER_5_154 ();
 sg13g2_decap_8 FILLER_5_161 ();
 sg13g2_decap_8 FILLER_5_168 ();
 sg13g2_decap_4 FILLER_5_175 ();
 sg13g2_fill_1 FILLER_5_179 ();
 sg13g2_fill_1 FILLER_5_214 ();
 sg13g2_decap_4 FILLER_5_241 ();
 sg13g2_fill_2 FILLER_5_245 ();
 sg13g2_decap_8 FILLER_5_251 ();
 sg13g2_decap_8 FILLER_5_258 ();
 sg13g2_decap_8 FILLER_5_265 ();
 sg13g2_decap_8 FILLER_5_272 ();
 sg13g2_decap_8 FILLER_5_279 ();
 sg13g2_decap_8 FILLER_5_286 ();
 sg13g2_decap_8 FILLER_5_293 ();
 sg13g2_fill_2 FILLER_5_300 ();
 sg13g2_decap_4 FILLER_5_314 ();
 sg13g2_decap_4 FILLER_5_343 ();
 sg13g2_decap_8 FILLER_5_352 ();
 sg13g2_decap_8 FILLER_5_359 ();
 sg13g2_fill_2 FILLER_5_366 ();
 sg13g2_fill_2 FILLER_5_373 ();
 sg13g2_fill_1 FILLER_5_385 ();
 sg13g2_fill_2 FILLER_5_390 ();
 sg13g2_fill_1 FILLER_5_396 ();
 sg13g2_fill_2 FILLER_5_402 ();
 sg13g2_fill_1 FILLER_5_410 ();
 sg13g2_decap_8 FILLER_5_418 ();
 sg13g2_decap_4 FILLER_5_425 ();
 sg13g2_fill_1 FILLER_5_429 ();
 sg13g2_decap_8 FILLER_6_0 ();
 sg13g2_decap_8 FILLER_6_7 ();
 sg13g2_decap_8 FILLER_6_14 ();
 sg13g2_decap_8 FILLER_6_21 ();
 sg13g2_decap_8 FILLER_6_28 ();
 sg13g2_decap_8 FILLER_6_35 ();
 sg13g2_decap_8 FILLER_6_42 ();
 sg13g2_decap_8 FILLER_6_49 ();
 sg13g2_decap_8 FILLER_6_56 ();
 sg13g2_decap_8 FILLER_6_63 ();
 sg13g2_decap_8 FILLER_6_70 ();
 sg13g2_decap_8 FILLER_6_77 ();
 sg13g2_decap_8 FILLER_6_84 ();
 sg13g2_decap_8 FILLER_6_91 ();
 sg13g2_decap_8 FILLER_6_98 ();
 sg13g2_decap_8 FILLER_6_105 ();
 sg13g2_decap_8 FILLER_6_112 ();
 sg13g2_decap_8 FILLER_6_119 ();
 sg13g2_decap_8 FILLER_6_126 ();
 sg13g2_decap_8 FILLER_6_133 ();
 sg13g2_decap_8 FILLER_6_140 ();
 sg13g2_decap_8 FILLER_6_147 ();
 sg13g2_decap_8 FILLER_6_154 ();
 sg13g2_decap_8 FILLER_6_161 ();
 sg13g2_decap_8 FILLER_6_168 ();
 sg13g2_decap_8 FILLER_6_175 ();
 sg13g2_decap_4 FILLER_6_182 ();
 sg13g2_fill_1 FILLER_6_186 ();
 sg13g2_decap_4 FILLER_6_190 ();
 sg13g2_fill_1 FILLER_6_194 ();
 sg13g2_fill_1 FILLER_6_199 ();
 sg13g2_fill_2 FILLER_6_226 ();
 sg13g2_fill_1 FILLER_6_228 ();
 sg13g2_decap_8 FILLER_6_234 ();
 sg13g2_fill_1 FILLER_6_241 ();
 sg13g2_decap_8 FILLER_6_277 ();
 sg13g2_decap_8 FILLER_6_284 ();
 sg13g2_fill_2 FILLER_6_291 ();
 sg13g2_fill_1 FILLER_6_293 ();
 sg13g2_decap_4 FILLER_6_299 ();
 sg13g2_fill_2 FILLER_6_308 ();
 sg13g2_fill_2 FILLER_6_314 ();
 sg13g2_fill_2 FILLER_6_322 ();
 sg13g2_fill_1 FILLER_6_333 ();
 sg13g2_fill_1 FILLER_6_342 ();
 sg13g2_fill_1 FILLER_6_347 ();
 sg13g2_fill_2 FILLER_6_366 ();
 sg13g2_fill_1 FILLER_6_391 ();
 sg13g2_decap_4 FILLER_6_400 ();
 sg13g2_decap_8 FILLER_6_409 ();
 sg13g2_decap_8 FILLER_6_416 ();
 sg13g2_decap_8 FILLER_6_423 ();
 sg13g2_decap_8 FILLER_7_0 ();
 sg13g2_decap_8 FILLER_7_7 ();
 sg13g2_decap_8 FILLER_7_14 ();
 sg13g2_decap_8 FILLER_7_21 ();
 sg13g2_decap_8 FILLER_7_28 ();
 sg13g2_decap_8 FILLER_7_35 ();
 sg13g2_decap_8 FILLER_7_42 ();
 sg13g2_decap_8 FILLER_7_49 ();
 sg13g2_decap_8 FILLER_7_56 ();
 sg13g2_decap_8 FILLER_7_63 ();
 sg13g2_decap_8 FILLER_7_70 ();
 sg13g2_decap_8 FILLER_7_77 ();
 sg13g2_decap_8 FILLER_7_84 ();
 sg13g2_decap_8 FILLER_7_91 ();
 sg13g2_decap_8 FILLER_7_98 ();
 sg13g2_decap_8 FILLER_7_105 ();
 sg13g2_decap_8 FILLER_7_112 ();
 sg13g2_decap_8 FILLER_7_119 ();
 sg13g2_decap_8 FILLER_7_126 ();
 sg13g2_decap_8 FILLER_7_133 ();
 sg13g2_decap_8 FILLER_7_140 ();
 sg13g2_decap_4 FILLER_7_147 ();
 sg13g2_fill_2 FILLER_7_151 ();
 sg13g2_decap_8 FILLER_7_157 ();
 sg13g2_decap_8 FILLER_7_164 ();
 sg13g2_decap_8 FILLER_7_171 ();
 sg13g2_fill_1 FILLER_7_178 ();
 sg13g2_fill_2 FILLER_7_192 ();
 sg13g2_decap_4 FILLER_7_208 ();
 sg13g2_fill_1 FILLER_7_212 ();
 sg13g2_fill_1 FILLER_7_218 ();
 sg13g2_fill_2 FILLER_7_230 ();
 sg13g2_decap_8 FILLER_7_241 ();
 sg13g2_decap_8 FILLER_7_248 ();
 sg13g2_fill_1 FILLER_7_255 ();
 sg13g2_fill_1 FILLER_7_273 ();
 sg13g2_decap_4 FILLER_7_282 ();
 sg13g2_fill_2 FILLER_7_286 ();
 sg13g2_fill_2 FILLER_7_334 ();
 sg13g2_fill_1 FILLER_7_336 ();
 sg13g2_decap_4 FILLER_7_357 ();
 sg13g2_decap_4 FILLER_7_383 ();
 sg13g2_fill_1 FILLER_7_387 ();
 sg13g2_fill_2 FILLER_7_406 ();
 sg13g2_decap_8 FILLER_7_416 ();
 sg13g2_decap_8 FILLER_7_423 ();
 sg13g2_decap_8 FILLER_8_0 ();
 sg13g2_decap_8 FILLER_8_7 ();
 sg13g2_decap_8 FILLER_8_14 ();
 sg13g2_decap_8 FILLER_8_21 ();
 sg13g2_decap_8 FILLER_8_28 ();
 sg13g2_decap_8 FILLER_8_35 ();
 sg13g2_decap_8 FILLER_8_42 ();
 sg13g2_decap_8 FILLER_8_49 ();
 sg13g2_decap_8 FILLER_8_56 ();
 sg13g2_decap_8 FILLER_8_63 ();
 sg13g2_decap_8 FILLER_8_70 ();
 sg13g2_decap_8 FILLER_8_77 ();
 sg13g2_decap_8 FILLER_8_84 ();
 sg13g2_decap_8 FILLER_8_91 ();
 sg13g2_decap_8 FILLER_8_98 ();
 sg13g2_decap_8 FILLER_8_105 ();
 sg13g2_decap_8 FILLER_8_112 ();
 sg13g2_decap_8 FILLER_8_119 ();
 sg13g2_decap_8 FILLER_8_126 ();
 sg13g2_decap_8 FILLER_8_133 ();
 sg13g2_decap_4 FILLER_8_140 ();
 sg13g2_fill_2 FILLER_8_144 ();
 sg13g2_fill_1 FILLER_8_176 ();
 sg13g2_fill_2 FILLER_8_200 ();
 sg13g2_fill_1 FILLER_8_202 ();
 sg13g2_decap_4 FILLER_8_208 ();
 sg13g2_fill_2 FILLER_8_212 ();
 sg13g2_fill_1 FILLER_8_223 ();
 sg13g2_fill_1 FILLER_8_229 ();
 sg13g2_decap_8 FILLER_8_256 ();
 sg13g2_decap_4 FILLER_8_263 ();
 sg13g2_fill_2 FILLER_8_267 ();
 sg13g2_decap_8 FILLER_8_274 ();
 sg13g2_decap_8 FILLER_8_281 ();
 sg13g2_decap_4 FILLER_8_288 ();
 sg13g2_fill_2 FILLER_8_292 ();
 sg13g2_decap_8 FILLER_8_299 ();
 sg13g2_decap_8 FILLER_8_306 ();
 sg13g2_fill_2 FILLER_8_325 ();
 sg13g2_fill_1 FILLER_8_327 ();
 sg13g2_fill_1 FILLER_8_356 ();
 sg13g2_fill_1 FILLER_8_369 ();
 sg13g2_decap_8 FILLER_8_377 ();
 sg13g2_decap_8 FILLER_8_384 ();
 sg13g2_decap_8 FILLER_8_398 ();
 sg13g2_decap_8 FILLER_8_405 ();
 sg13g2_decap_8 FILLER_8_412 ();
 sg13g2_decap_8 FILLER_8_419 ();
 sg13g2_decap_4 FILLER_8_426 ();
 sg13g2_decap_8 FILLER_9_0 ();
 sg13g2_decap_8 FILLER_9_7 ();
 sg13g2_decap_8 FILLER_9_14 ();
 sg13g2_decap_8 FILLER_9_21 ();
 sg13g2_decap_8 FILLER_9_28 ();
 sg13g2_decap_8 FILLER_9_35 ();
 sg13g2_decap_8 FILLER_9_42 ();
 sg13g2_decap_8 FILLER_9_49 ();
 sg13g2_decap_8 FILLER_9_56 ();
 sg13g2_decap_8 FILLER_9_63 ();
 sg13g2_decap_8 FILLER_9_70 ();
 sg13g2_decap_8 FILLER_9_77 ();
 sg13g2_decap_8 FILLER_9_84 ();
 sg13g2_decap_8 FILLER_9_91 ();
 sg13g2_decap_8 FILLER_9_98 ();
 sg13g2_decap_8 FILLER_9_105 ();
 sg13g2_decap_8 FILLER_9_112 ();
 sg13g2_decap_8 FILLER_9_119 ();
 sg13g2_decap_4 FILLER_9_126 ();
 sg13g2_decap_4 FILLER_9_160 ();
 sg13g2_fill_2 FILLER_9_164 ();
 sg13g2_fill_1 FILLER_9_170 ();
 sg13g2_fill_1 FILLER_9_179 ();
 sg13g2_fill_2 FILLER_9_185 ();
 sg13g2_fill_2 FILLER_9_192 ();
 sg13g2_fill_2 FILLER_9_198 ();
 sg13g2_fill_1 FILLER_9_200 ();
 sg13g2_decap_4 FILLER_9_205 ();
 sg13g2_fill_2 FILLER_9_209 ();
 sg13g2_decap_8 FILLER_9_216 ();
 sg13g2_fill_2 FILLER_9_223 ();
 sg13g2_decap_4 FILLER_9_228 ();
 sg13g2_fill_2 FILLER_9_232 ();
 sg13g2_decap_8 FILLER_9_239 ();
 sg13g2_fill_1 FILLER_9_246 ();
 sg13g2_decap_8 FILLER_9_251 ();
 sg13g2_decap_4 FILLER_9_258 ();
 sg13g2_fill_1 FILLER_9_262 ();
 sg13g2_decap_4 FILLER_9_275 ();
 sg13g2_fill_2 FILLER_9_279 ();
 sg13g2_fill_2 FILLER_9_305 ();
 sg13g2_fill_1 FILLER_9_307 ();
 sg13g2_fill_1 FILLER_9_317 ();
 sg13g2_decap_8 FILLER_9_333 ();
 sg13g2_decap_4 FILLER_9_340 ();
 sg13g2_fill_1 FILLER_9_344 ();
 sg13g2_decap_8 FILLER_9_350 ();
 sg13g2_fill_2 FILLER_9_369 ();
 sg13g2_fill_1 FILLER_9_371 ();
 sg13g2_decap_8 FILLER_9_376 ();
 sg13g2_decap_8 FILLER_9_383 ();
 sg13g2_decap_8 FILLER_9_390 ();
 sg13g2_decap_8 FILLER_9_397 ();
 sg13g2_decap_8 FILLER_9_404 ();
 sg13g2_fill_2 FILLER_9_411 ();
 sg13g2_decap_8 FILLER_9_419 ();
 sg13g2_decap_4 FILLER_9_426 ();
 sg13g2_decap_8 FILLER_10_0 ();
 sg13g2_decap_8 FILLER_10_7 ();
 sg13g2_decap_8 FILLER_10_14 ();
 sg13g2_decap_8 FILLER_10_21 ();
 sg13g2_decap_8 FILLER_10_28 ();
 sg13g2_decap_8 FILLER_10_35 ();
 sg13g2_decap_8 FILLER_10_42 ();
 sg13g2_decap_8 FILLER_10_49 ();
 sg13g2_decap_8 FILLER_10_56 ();
 sg13g2_decap_8 FILLER_10_63 ();
 sg13g2_decap_8 FILLER_10_70 ();
 sg13g2_decap_8 FILLER_10_77 ();
 sg13g2_decap_8 FILLER_10_84 ();
 sg13g2_decap_8 FILLER_10_91 ();
 sg13g2_decap_8 FILLER_10_98 ();
 sg13g2_decap_8 FILLER_10_105 ();
 sg13g2_decap_8 FILLER_10_112 ();
 sg13g2_decap_8 FILLER_10_119 ();
 sg13g2_decap_8 FILLER_10_126 ();
 sg13g2_fill_2 FILLER_10_133 ();
 sg13g2_decap_8 FILLER_10_139 ();
 sg13g2_decap_8 FILLER_10_146 ();
 sg13g2_fill_1 FILLER_10_157 ();
 sg13g2_fill_2 FILLER_10_206 ();
 sg13g2_fill_1 FILLER_10_208 ();
 sg13g2_decap_4 FILLER_10_225 ();
 sg13g2_fill_1 FILLER_10_229 ();
 sg13g2_fill_2 FILLER_10_238 ();
 sg13g2_decap_8 FILLER_10_266 ();
 sg13g2_decap_4 FILLER_10_273 ();
 sg13g2_decap_4 FILLER_10_282 ();
 sg13g2_fill_2 FILLER_10_286 ();
 sg13g2_fill_2 FILLER_10_292 ();
 sg13g2_fill_1 FILLER_10_298 ();
 sg13g2_fill_1 FILLER_10_308 ();
 sg13g2_fill_1 FILLER_10_314 ();
 sg13g2_fill_2 FILLER_10_334 ();
 sg13g2_fill_1 FILLER_10_336 ();
 sg13g2_fill_1 FILLER_10_341 ();
 sg13g2_fill_2 FILLER_10_358 ();
 sg13g2_fill_1 FILLER_10_360 ();
 sg13g2_decap_8 FILLER_10_365 ();
 sg13g2_decap_8 FILLER_10_372 ();
 sg13g2_decap_8 FILLER_10_379 ();
 sg13g2_fill_2 FILLER_10_394 ();
 sg13g2_fill_1 FILLER_10_396 ();
 sg13g2_fill_1 FILLER_10_406 ();
 sg13g2_fill_1 FILLER_10_416 ();
 sg13g2_decap_8 FILLER_10_422 ();
 sg13g2_fill_1 FILLER_10_429 ();
 sg13g2_decap_8 FILLER_11_0 ();
 sg13g2_decap_8 FILLER_11_7 ();
 sg13g2_decap_8 FILLER_11_14 ();
 sg13g2_decap_8 FILLER_11_21 ();
 sg13g2_decap_8 FILLER_11_28 ();
 sg13g2_decap_8 FILLER_11_35 ();
 sg13g2_decap_8 FILLER_11_42 ();
 sg13g2_decap_8 FILLER_11_49 ();
 sg13g2_decap_8 FILLER_11_56 ();
 sg13g2_decap_8 FILLER_11_63 ();
 sg13g2_decap_8 FILLER_11_70 ();
 sg13g2_decap_8 FILLER_11_77 ();
 sg13g2_decap_8 FILLER_11_84 ();
 sg13g2_decap_8 FILLER_11_91 ();
 sg13g2_decap_8 FILLER_11_98 ();
 sg13g2_decap_8 FILLER_11_105 ();
 sg13g2_decap_8 FILLER_11_112 ();
 sg13g2_decap_8 FILLER_11_119 ();
 sg13g2_decap_8 FILLER_11_126 ();
 sg13g2_decap_8 FILLER_11_133 ();
 sg13g2_decap_8 FILLER_11_140 ();
 sg13g2_decap_8 FILLER_11_147 ();
 sg13g2_fill_2 FILLER_11_154 ();
 sg13g2_decap_8 FILLER_11_186 ();
 sg13g2_fill_2 FILLER_11_193 ();
 sg13g2_fill_1 FILLER_11_195 ();
 sg13g2_decap_8 FILLER_11_209 ();
 sg13g2_fill_2 FILLER_11_216 ();
 sg13g2_decap_8 FILLER_11_223 ();
 sg13g2_decap_8 FILLER_11_256 ();
 sg13g2_decap_8 FILLER_11_263 ();
 sg13g2_fill_2 FILLER_11_270 ();
 sg13g2_fill_1 FILLER_11_302 ();
 sg13g2_fill_2 FILLER_11_311 ();
 sg13g2_fill_2 FILLER_11_321 ();
 sg13g2_fill_1 FILLER_11_323 ();
 sg13g2_fill_2 FILLER_11_355 ();
 sg13g2_fill_1 FILLER_11_361 ();
 sg13g2_fill_2 FILLER_11_380 ();
 sg13g2_fill_1 FILLER_11_382 ();
 sg13g2_fill_1 FILLER_11_392 ();
 sg13g2_fill_2 FILLER_11_396 ();
 sg13g2_fill_1 FILLER_11_398 ();
 sg13g2_decap_4 FILLER_11_424 ();
 sg13g2_fill_2 FILLER_11_428 ();
 sg13g2_decap_8 FILLER_12_0 ();
 sg13g2_decap_8 FILLER_12_7 ();
 sg13g2_decap_8 FILLER_12_14 ();
 sg13g2_decap_8 FILLER_12_21 ();
 sg13g2_decap_8 FILLER_12_28 ();
 sg13g2_decap_8 FILLER_12_35 ();
 sg13g2_decap_8 FILLER_12_42 ();
 sg13g2_decap_8 FILLER_12_49 ();
 sg13g2_decap_8 FILLER_12_56 ();
 sg13g2_decap_8 FILLER_12_63 ();
 sg13g2_decap_8 FILLER_12_70 ();
 sg13g2_decap_8 FILLER_12_77 ();
 sg13g2_decap_8 FILLER_12_84 ();
 sg13g2_decap_8 FILLER_12_91 ();
 sg13g2_decap_8 FILLER_12_98 ();
 sg13g2_decap_8 FILLER_12_105 ();
 sg13g2_decap_8 FILLER_12_112 ();
 sg13g2_fill_2 FILLER_12_119 ();
 sg13g2_fill_1 FILLER_12_147 ();
 sg13g2_decap_4 FILLER_12_152 ();
 sg13g2_fill_1 FILLER_12_156 ();
 sg13g2_fill_2 FILLER_12_162 ();
 sg13g2_fill_1 FILLER_12_164 ();
 sg13g2_fill_1 FILLER_12_170 ();
 sg13g2_fill_2 FILLER_12_176 ();
 sg13g2_fill_1 FILLER_12_178 ();
 sg13g2_decap_4 FILLER_12_192 ();
 sg13g2_decap_4 FILLER_12_209 ();
 sg13g2_decap_4 FILLER_12_226 ();
 sg13g2_decap_8 FILLER_12_238 ();
 sg13g2_fill_1 FILLER_12_245 ();
 sg13g2_decap_4 FILLER_12_253 ();
 sg13g2_fill_1 FILLER_12_273 ();
 sg13g2_fill_1 FILLER_12_278 ();
 sg13g2_fill_1 FILLER_12_283 ();
 sg13g2_decap_8 FILLER_12_289 ();
 sg13g2_decap_8 FILLER_12_296 ();
 sg13g2_decap_8 FILLER_12_303 ();
 sg13g2_decap_8 FILLER_12_310 ();
 sg13g2_decap_8 FILLER_12_317 ();
 sg13g2_decap_8 FILLER_12_324 ();
 sg13g2_fill_1 FILLER_12_331 ();
 sg13g2_fill_2 FILLER_12_350 ();
 sg13g2_fill_1 FILLER_12_352 ();
 sg13g2_decap_4 FILLER_12_358 ();
 sg13g2_fill_2 FILLER_12_362 ();
 sg13g2_fill_1 FILLER_12_372 ();
 sg13g2_decap_4 FILLER_12_377 ();
 sg13g2_fill_2 FILLER_12_395 ();
 sg13g2_fill_1 FILLER_12_397 ();
 sg13g2_decap_4 FILLER_12_402 ();
 sg13g2_decap_8 FILLER_12_423 ();
 sg13g2_decap_8 FILLER_13_0 ();
 sg13g2_decap_8 FILLER_13_7 ();
 sg13g2_decap_8 FILLER_13_14 ();
 sg13g2_decap_8 FILLER_13_21 ();
 sg13g2_decap_8 FILLER_13_28 ();
 sg13g2_decap_8 FILLER_13_35 ();
 sg13g2_decap_8 FILLER_13_42 ();
 sg13g2_decap_8 FILLER_13_49 ();
 sg13g2_decap_8 FILLER_13_56 ();
 sg13g2_decap_8 FILLER_13_63 ();
 sg13g2_decap_8 FILLER_13_70 ();
 sg13g2_decap_8 FILLER_13_77 ();
 sg13g2_decap_8 FILLER_13_84 ();
 sg13g2_decap_8 FILLER_13_91 ();
 sg13g2_decap_8 FILLER_13_98 ();
 sg13g2_decap_8 FILLER_13_105 ();
 sg13g2_decap_8 FILLER_13_112 ();
 sg13g2_decap_8 FILLER_13_119 ();
 sg13g2_fill_1 FILLER_13_126 ();
 sg13g2_decap_8 FILLER_13_131 ();
 sg13g2_decap_8 FILLER_13_138 ();
 sg13g2_fill_2 FILLER_13_149 ();
 sg13g2_decap_4 FILLER_13_159 ();
 sg13g2_decap_8 FILLER_13_172 ();
 sg13g2_decap_4 FILLER_13_179 ();
 sg13g2_fill_2 FILLER_13_187 ();
 sg13g2_decap_8 FILLER_13_198 ();
 sg13g2_decap_8 FILLER_13_205 ();
 sg13g2_decap_4 FILLER_13_212 ();
 sg13g2_fill_1 FILLER_13_216 ();
 sg13g2_fill_1 FILLER_13_230 ();
 sg13g2_fill_1 FILLER_13_235 ();
 sg13g2_fill_2 FILLER_13_240 ();
 sg13g2_fill_1 FILLER_13_242 ();
 sg13g2_decap_8 FILLER_13_260 ();
 sg13g2_fill_1 FILLER_13_267 ();
 sg13g2_fill_2 FILLER_13_298 ();
 sg13g2_fill_1 FILLER_13_304 ();
 sg13g2_decap_4 FILLER_13_310 ();
 sg13g2_decap_4 FILLER_13_322 ();
 sg13g2_fill_1 FILLER_13_326 ();
 sg13g2_fill_2 FILLER_13_351 ();
 sg13g2_fill_2 FILLER_13_366 ();
 sg13g2_decap_4 FILLER_13_375 ();
 sg13g2_fill_2 FILLER_13_387 ();
 sg13g2_decap_4 FILLER_13_397 ();
 sg13g2_decap_8 FILLER_13_422 ();
 sg13g2_fill_1 FILLER_13_429 ();
 sg13g2_decap_8 FILLER_14_0 ();
 sg13g2_decap_8 FILLER_14_7 ();
 sg13g2_decap_8 FILLER_14_14 ();
 sg13g2_decap_8 FILLER_14_21 ();
 sg13g2_decap_8 FILLER_14_28 ();
 sg13g2_decap_8 FILLER_14_35 ();
 sg13g2_decap_8 FILLER_14_42 ();
 sg13g2_decap_8 FILLER_14_49 ();
 sg13g2_decap_8 FILLER_14_56 ();
 sg13g2_decap_8 FILLER_14_63 ();
 sg13g2_decap_8 FILLER_14_70 ();
 sg13g2_decap_8 FILLER_14_77 ();
 sg13g2_decap_8 FILLER_14_84 ();
 sg13g2_decap_8 FILLER_14_91 ();
 sg13g2_decap_8 FILLER_14_98 ();
 sg13g2_decap_8 FILLER_14_105 ();
 sg13g2_decap_8 FILLER_14_112 ();
 sg13g2_decap_8 FILLER_14_119 ();
 sg13g2_decap_8 FILLER_14_126 ();
 sg13g2_decap_8 FILLER_14_133 ();
 sg13g2_decap_8 FILLER_14_140 ();
 sg13g2_decap_4 FILLER_14_147 ();
 sg13g2_fill_2 FILLER_14_151 ();
 sg13g2_decap_8 FILLER_14_158 ();
 sg13g2_fill_1 FILLER_14_179 ();
 sg13g2_fill_1 FILLER_14_184 ();
 sg13g2_decap_8 FILLER_14_211 ();
 sg13g2_decap_4 FILLER_14_229 ();
 sg13g2_fill_2 FILLER_14_233 ();
 sg13g2_fill_2 FILLER_14_242 ();
 sg13g2_decap_8 FILLER_14_249 ();
 sg13g2_fill_1 FILLER_14_256 ();
 sg13g2_decap_8 FILLER_14_261 ();
 sg13g2_decap_4 FILLER_14_268 ();
 sg13g2_decap_8 FILLER_14_276 ();
 sg13g2_decap_8 FILLER_14_283 ();
 sg13g2_fill_1 FILLER_14_320 ();
 sg13g2_fill_1 FILLER_14_326 ();
 sg13g2_decap_4 FILLER_14_332 ();
 sg13g2_fill_1 FILLER_14_336 ();
 sg13g2_decap_8 FILLER_14_342 ();
 sg13g2_fill_1 FILLER_14_349 ();
 sg13g2_fill_1 FILLER_14_355 ();
 sg13g2_fill_1 FILLER_14_361 ();
 sg13g2_decap_4 FILLER_14_382 ();
 sg13g2_decap_8 FILLER_14_391 ();
 sg13g2_decap_8 FILLER_14_405 ();
 sg13g2_decap_8 FILLER_14_412 ();
 sg13g2_decap_8 FILLER_14_419 ();
 sg13g2_decap_4 FILLER_14_426 ();
 sg13g2_decap_8 FILLER_15_0 ();
 sg13g2_decap_8 FILLER_15_7 ();
 sg13g2_decap_8 FILLER_15_14 ();
 sg13g2_decap_8 FILLER_15_21 ();
 sg13g2_decap_8 FILLER_15_28 ();
 sg13g2_decap_8 FILLER_15_35 ();
 sg13g2_decap_8 FILLER_15_42 ();
 sg13g2_decap_8 FILLER_15_49 ();
 sg13g2_decap_8 FILLER_15_56 ();
 sg13g2_decap_8 FILLER_15_63 ();
 sg13g2_decap_8 FILLER_15_70 ();
 sg13g2_decap_8 FILLER_15_77 ();
 sg13g2_decap_8 FILLER_15_84 ();
 sg13g2_decap_8 FILLER_15_91 ();
 sg13g2_decap_8 FILLER_15_98 ();
 sg13g2_decap_8 FILLER_15_105 ();
 sg13g2_decap_8 FILLER_15_112 ();
 sg13g2_decap_8 FILLER_15_119 ();
 sg13g2_decap_8 FILLER_15_126 ();
 sg13g2_fill_2 FILLER_15_133 ();
 sg13g2_fill_2 FILLER_15_161 ();
 sg13g2_fill_1 FILLER_15_163 ();
 sg13g2_fill_2 FILLER_15_169 ();
 sg13g2_fill_1 FILLER_15_171 ();
 sg13g2_fill_2 FILLER_15_178 ();
 sg13g2_fill_2 FILLER_15_188 ();
 sg13g2_fill_1 FILLER_15_190 ();
 sg13g2_fill_2 FILLER_15_199 ();
 sg13g2_fill_1 FILLER_15_201 ();
 sg13g2_fill_2 FILLER_15_207 ();
 sg13g2_fill_1 FILLER_15_217 ();
 sg13g2_fill_2 FILLER_15_223 ();
 sg13g2_decap_4 FILLER_15_237 ();
 sg13g2_fill_1 FILLER_15_241 ();
 sg13g2_decap_4 FILLER_15_284 ();
 sg13g2_fill_1 FILLER_15_288 ();
 sg13g2_fill_1 FILLER_15_294 ();
 sg13g2_fill_1 FILLER_15_303 ();
 sg13g2_fill_1 FILLER_15_329 ();
 sg13g2_decap_8 FILLER_15_334 ();
 sg13g2_decap_8 FILLER_15_341 ();
 sg13g2_fill_1 FILLER_15_348 ();
 sg13g2_decap_8 FILLER_15_365 ();
 sg13g2_decap_8 FILLER_15_372 ();
 sg13g2_decap_4 FILLER_15_379 ();
 sg13g2_decap_8 FILLER_15_398 ();
 sg13g2_fill_2 FILLER_15_405 ();
 sg13g2_fill_1 FILLER_15_407 ();
 sg13g2_decap_8 FILLER_15_419 ();
 sg13g2_decap_4 FILLER_15_426 ();
 sg13g2_decap_8 FILLER_16_0 ();
 sg13g2_decap_8 FILLER_16_7 ();
 sg13g2_decap_8 FILLER_16_14 ();
 sg13g2_decap_8 FILLER_16_21 ();
 sg13g2_decap_8 FILLER_16_28 ();
 sg13g2_decap_8 FILLER_16_35 ();
 sg13g2_decap_8 FILLER_16_42 ();
 sg13g2_decap_8 FILLER_16_49 ();
 sg13g2_decap_8 FILLER_16_56 ();
 sg13g2_decap_8 FILLER_16_63 ();
 sg13g2_decap_8 FILLER_16_70 ();
 sg13g2_decap_8 FILLER_16_77 ();
 sg13g2_decap_8 FILLER_16_84 ();
 sg13g2_decap_8 FILLER_16_91 ();
 sg13g2_decap_8 FILLER_16_98 ();
 sg13g2_decap_8 FILLER_16_105 ();
 sg13g2_decap_8 FILLER_16_112 ();
 sg13g2_decap_8 FILLER_16_119 ();
 sg13g2_decap_8 FILLER_16_126 ();
 sg13g2_decap_8 FILLER_16_133 ();
 sg13g2_fill_1 FILLER_16_140 ();
 sg13g2_decap_8 FILLER_16_145 ();
 sg13g2_decap_4 FILLER_16_152 ();
 sg13g2_fill_1 FILLER_16_156 ();
 sg13g2_fill_1 FILLER_16_166 ();
 sg13g2_decap_8 FILLER_16_180 ();
 sg13g2_decap_4 FILLER_16_187 ();
 sg13g2_fill_2 FILLER_16_191 ();
 sg13g2_decap_4 FILLER_16_212 ();
 sg13g2_fill_1 FILLER_16_227 ();
 sg13g2_decap_8 FILLER_16_259 ();
 sg13g2_fill_2 FILLER_16_266 ();
 sg13g2_fill_2 FILLER_16_277 ();
 sg13g2_fill_1 FILLER_16_279 ();
 sg13g2_decap_4 FILLER_16_288 ();
 sg13g2_decap_8 FILLER_16_302 ();
 sg13g2_fill_2 FILLER_16_309 ();
 sg13g2_fill_1 FILLER_16_311 ();
 sg13g2_fill_2 FILLER_16_316 ();
 sg13g2_fill_2 FILLER_16_326 ();
 sg13g2_fill_2 FILLER_16_340 ();
 sg13g2_fill_1 FILLER_16_342 ();
 sg13g2_fill_2 FILLER_16_347 ();
 sg13g2_decap_8 FILLER_16_361 ();
 sg13g2_decap_8 FILLER_16_368 ();
 sg13g2_decap_4 FILLER_16_375 ();
 sg13g2_decap_8 FILLER_16_390 ();
 sg13g2_fill_2 FILLER_16_397 ();
 sg13g2_fill_2 FILLER_16_413 ();
 sg13g2_decap_8 FILLER_16_420 ();
 sg13g2_fill_2 FILLER_16_427 ();
 sg13g2_fill_1 FILLER_16_429 ();
 sg13g2_decap_8 FILLER_17_0 ();
 sg13g2_decap_8 FILLER_17_7 ();
 sg13g2_decap_8 FILLER_17_14 ();
 sg13g2_decap_8 FILLER_17_21 ();
 sg13g2_decap_8 FILLER_17_28 ();
 sg13g2_decap_8 FILLER_17_35 ();
 sg13g2_decap_8 FILLER_17_42 ();
 sg13g2_decap_8 FILLER_17_49 ();
 sg13g2_decap_8 FILLER_17_56 ();
 sg13g2_decap_8 FILLER_17_63 ();
 sg13g2_decap_8 FILLER_17_70 ();
 sg13g2_decap_8 FILLER_17_77 ();
 sg13g2_decap_8 FILLER_17_84 ();
 sg13g2_decap_8 FILLER_17_91 ();
 sg13g2_decap_8 FILLER_17_98 ();
 sg13g2_decap_8 FILLER_17_105 ();
 sg13g2_fill_2 FILLER_17_112 ();
 sg13g2_fill_1 FILLER_17_148 ();
 sg13g2_fill_1 FILLER_17_164 ();
 sg13g2_decap_8 FILLER_17_172 ();
 sg13g2_fill_1 FILLER_17_179 ();
 sg13g2_decap_8 FILLER_17_205 ();
 sg13g2_fill_2 FILLER_17_212 ();
 sg13g2_decap_8 FILLER_17_222 ();
 sg13g2_fill_2 FILLER_17_241 ();
 sg13g2_fill_1 FILLER_17_243 ();
 sg13g2_fill_2 FILLER_17_253 ();
 sg13g2_fill_1 FILLER_17_255 ();
 sg13g2_fill_1 FILLER_17_264 ();
 sg13g2_fill_2 FILLER_17_271 ();
 sg13g2_fill_1 FILLER_17_273 ();
 sg13g2_fill_1 FILLER_17_287 ();
 sg13g2_decap_8 FILLER_17_300 ();
 sg13g2_decap_8 FILLER_17_307 ();
 sg13g2_fill_1 FILLER_17_314 ();
 sg13g2_decap_8 FILLER_17_319 ();
 sg13g2_decap_4 FILLER_17_326 ();
 sg13g2_decap_8 FILLER_17_334 ();
 sg13g2_decap_8 FILLER_17_341 ();
 sg13g2_fill_2 FILLER_17_352 ();
 sg13g2_fill_1 FILLER_17_354 ();
 sg13g2_fill_2 FILLER_17_363 ();
 sg13g2_fill_1 FILLER_17_389 ();
 sg13g2_fill_2 FILLER_17_394 ();
 sg13g2_fill_2 FILLER_17_409 ();
 sg13g2_decap_8 FILLER_17_421 ();
 sg13g2_fill_2 FILLER_17_428 ();
 sg13g2_decap_8 FILLER_18_0 ();
 sg13g2_decap_8 FILLER_18_7 ();
 sg13g2_decap_8 FILLER_18_14 ();
 sg13g2_decap_8 FILLER_18_21 ();
 sg13g2_decap_8 FILLER_18_28 ();
 sg13g2_decap_8 FILLER_18_35 ();
 sg13g2_decap_8 FILLER_18_42 ();
 sg13g2_decap_8 FILLER_18_49 ();
 sg13g2_decap_8 FILLER_18_56 ();
 sg13g2_decap_8 FILLER_18_63 ();
 sg13g2_decap_8 FILLER_18_70 ();
 sg13g2_decap_8 FILLER_18_77 ();
 sg13g2_fill_2 FILLER_18_84 ();
 sg13g2_fill_1 FILLER_18_86 ();
 sg13g2_decap_8 FILLER_18_91 ();
 sg13g2_decap_4 FILLER_18_98 ();
 sg13g2_decap_4 FILLER_18_115 ();
 sg13g2_fill_1 FILLER_18_119 ();
 sg13g2_decap_8 FILLER_18_124 ();
 sg13g2_decap_8 FILLER_18_131 ();
 sg13g2_decap_4 FILLER_18_138 ();
 sg13g2_fill_1 FILLER_18_142 ();
 sg13g2_fill_1 FILLER_18_164 ();
 sg13g2_decap_4 FILLER_18_168 ();
 sg13g2_fill_2 FILLER_18_172 ();
 sg13g2_fill_1 FILLER_18_179 ();
 sg13g2_fill_2 FILLER_18_190 ();
 sg13g2_fill_1 FILLER_18_192 ();
 sg13g2_decap_4 FILLER_18_206 ();
 sg13g2_fill_1 FILLER_18_222 ();
 sg13g2_decap_4 FILLER_18_227 ();
 sg13g2_fill_2 FILLER_18_231 ();
 sg13g2_fill_2 FILLER_18_245 ();
 sg13g2_fill_2 FILLER_18_256 ();
 sg13g2_fill_1 FILLER_18_258 ();
 sg13g2_fill_2 FILLER_18_264 ();
 sg13g2_fill_1 FILLER_18_266 ();
 sg13g2_fill_1 FILLER_18_273 ();
 sg13g2_fill_2 FILLER_18_278 ();
 sg13g2_decap_8 FILLER_18_291 ();
 sg13g2_fill_2 FILLER_18_298 ();
 sg13g2_fill_1 FILLER_18_300 ();
 sg13g2_decap_4 FILLER_18_306 ();
 sg13g2_fill_1 FILLER_18_310 ();
 sg13g2_decap_8 FILLER_18_315 ();
 sg13g2_decap_4 FILLER_18_322 ();
 sg13g2_fill_2 FILLER_18_326 ();
 sg13g2_decap_8 FILLER_18_340 ();
 sg13g2_fill_1 FILLER_18_347 ();
 sg13g2_decap_8 FILLER_18_352 ();
 sg13g2_decap_4 FILLER_18_368 ();
 sg13g2_fill_2 FILLER_18_390 ();
 sg13g2_fill_1 FILLER_18_392 ();
 sg13g2_fill_1 FILLER_18_429 ();
 sg13g2_decap_8 FILLER_19_0 ();
 sg13g2_decap_8 FILLER_19_7 ();
 sg13g2_decap_8 FILLER_19_14 ();
 sg13g2_decap_8 FILLER_19_21 ();
 sg13g2_decap_8 FILLER_19_28 ();
 sg13g2_decap_8 FILLER_19_35 ();
 sg13g2_decap_8 FILLER_19_42 ();
 sg13g2_decap_8 FILLER_19_49 ();
 sg13g2_decap_8 FILLER_19_56 ();
 sg13g2_fill_1 FILLER_19_63 ();
 sg13g2_decap_8 FILLER_19_68 ();
 sg13g2_decap_4 FILLER_19_75 ();
 sg13g2_fill_1 FILLER_19_79 ();
 sg13g2_fill_2 FILLER_19_106 ();
 sg13g2_fill_2 FILLER_19_111 ();
 sg13g2_fill_1 FILLER_19_113 ();
 sg13g2_decap_4 FILLER_19_145 ();
 sg13g2_fill_1 FILLER_19_149 ();
 sg13g2_decap_8 FILLER_19_166 ();
 sg13g2_decap_4 FILLER_19_173 ();
 sg13g2_decap_4 FILLER_19_192 ();
 sg13g2_decap_4 FILLER_19_206 ();
 sg13g2_fill_1 FILLER_19_210 ();
 sg13g2_decap_4 FILLER_19_224 ();
 sg13g2_fill_1 FILLER_19_244 ();
 sg13g2_fill_1 FILLER_19_249 ();
 sg13g2_fill_1 FILLER_19_255 ();
 sg13g2_fill_1 FILLER_19_267 ();
 sg13g2_fill_1 FILLER_19_273 ();
 sg13g2_fill_1 FILLER_19_285 ();
 sg13g2_fill_2 FILLER_19_295 ();
 sg13g2_decap_4 FILLER_19_305 ();
 sg13g2_fill_1 FILLER_19_309 ();
 sg13g2_decap_4 FILLER_19_320 ();
 sg13g2_decap_4 FILLER_19_328 ();
 sg13g2_decap_8 FILLER_19_340 ();
 sg13g2_decap_8 FILLER_19_347 ();
 sg13g2_fill_1 FILLER_19_363 ();
 sg13g2_fill_1 FILLER_19_380 ();
 sg13g2_decap_4 FILLER_19_408 ();
 sg13g2_decap_8 FILLER_19_421 ();
 sg13g2_fill_2 FILLER_19_428 ();
 sg13g2_decap_8 FILLER_20_0 ();
 sg13g2_decap_8 FILLER_20_7 ();
 sg13g2_decap_8 FILLER_20_14 ();
 sg13g2_decap_8 FILLER_20_21 ();
 sg13g2_decap_8 FILLER_20_28 ();
 sg13g2_decap_8 FILLER_20_35 ();
 sg13g2_decap_8 FILLER_20_42 ();
 sg13g2_decap_8 FILLER_20_49 ();
 sg13g2_fill_1 FILLER_20_56 ();
 sg13g2_decap_8 FILLER_20_83 ();
 sg13g2_decap_8 FILLER_20_90 ();
 sg13g2_fill_1 FILLER_20_97 ();
 sg13g2_fill_2 FILLER_20_102 ();
 sg13g2_decap_8 FILLER_20_109 ();
 sg13g2_decap_4 FILLER_20_116 ();
 sg13g2_fill_1 FILLER_20_120 ();
 sg13g2_fill_2 FILLER_20_129 ();
 sg13g2_decap_8 FILLER_20_136 ();
 sg13g2_decap_8 FILLER_20_143 ();
 sg13g2_decap_4 FILLER_20_150 ();
 sg13g2_decap_8 FILLER_20_205 ();
 sg13g2_decap_4 FILLER_20_212 ();
 sg13g2_fill_1 FILLER_20_216 ();
 sg13g2_decap_8 FILLER_20_224 ();
 sg13g2_decap_8 FILLER_20_231 ();
 sg13g2_decap_4 FILLER_20_238 ();
 sg13g2_decap_8 FILLER_20_261 ();
 sg13g2_decap_4 FILLER_20_268 ();
 sg13g2_fill_1 FILLER_20_286 ();
 sg13g2_fill_1 FILLER_20_292 ();
 sg13g2_fill_1 FILLER_20_297 ();
 sg13g2_fill_2 FILLER_20_306 ();
 sg13g2_decap_8 FILLER_20_313 ();
 sg13g2_fill_1 FILLER_20_320 ();
 sg13g2_fill_1 FILLER_20_325 ();
 sg13g2_fill_2 FILLER_20_335 ();
 sg13g2_decap_8 FILLER_20_341 ();
 sg13g2_decap_8 FILLER_20_364 ();
 sg13g2_fill_2 FILLER_20_387 ();
 sg13g2_fill_1 FILLER_20_389 ();
 sg13g2_fill_2 FILLER_20_395 ();
 sg13g2_fill_1 FILLER_20_397 ();
 sg13g2_fill_2 FILLER_20_402 ();
 sg13g2_decap_8 FILLER_20_421 ();
 sg13g2_fill_2 FILLER_20_428 ();
 sg13g2_decap_8 FILLER_21_0 ();
 sg13g2_decap_8 FILLER_21_7 ();
 sg13g2_decap_8 FILLER_21_14 ();
 sg13g2_decap_8 FILLER_21_21 ();
 sg13g2_decap_8 FILLER_21_28 ();
 sg13g2_decap_8 FILLER_21_35 ();
 sg13g2_decap_8 FILLER_21_42 ();
 sg13g2_decap_8 FILLER_21_49 ();
 sg13g2_fill_1 FILLER_21_56 ();
 sg13g2_decap_8 FILLER_21_61 ();
 sg13g2_decap_8 FILLER_21_68 ();
 sg13g2_fill_2 FILLER_21_75 ();
 sg13g2_fill_1 FILLER_21_77 ();
 sg13g2_decap_8 FILLER_21_117 ();
 sg13g2_decap_8 FILLER_21_144 ();
 sg13g2_decap_8 FILLER_21_151 ();
 sg13g2_fill_2 FILLER_21_158 ();
 sg13g2_decap_4 FILLER_21_164 ();
 sg13g2_fill_2 FILLER_21_168 ();
 sg13g2_decap_8 FILLER_21_174 ();
 sg13g2_decap_8 FILLER_21_181 ();
 sg13g2_fill_2 FILLER_21_188 ();
 sg13g2_decap_8 FILLER_21_194 ();
 sg13g2_fill_2 FILLER_21_201 ();
 sg13g2_decap_8 FILLER_21_212 ();
 sg13g2_fill_1 FILLER_21_219 ();
 sg13g2_decap_8 FILLER_21_228 ();
 sg13g2_fill_1 FILLER_21_235 ();
 sg13g2_decap_8 FILLER_21_244 ();
 sg13g2_fill_1 FILLER_21_256 ();
 sg13g2_fill_1 FILLER_21_261 ();
 sg13g2_fill_2 FILLER_21_267 ();
 sg13g2_fill_1 FILLER_21_269 ();
 sg13g2_fill_1 FILLER_21_278 ();
 sg13g2_decap_4 FILLER_21_284 ();
 sg13g2_fill_2 FILLER_21_297 ();
 sg13g2_decap_8 FILLER_21_304 ();
 sg13g2_decap_4 FILLER_21_311 ();
 sg13g2_fill_1 FILLER_21_315 ();
 sg13g2_decap_8 FILLER_21_332 ();
 sg13g2_decap_8 FILLER_21_339 ();
 sg13g2_fill_2 FILLER_21_354 ();
 sg13g2_decap_8 FILLER_21_361 ();
 sg13g2_fill_1 FILLER_21_368 ();
 sg13g2_fill_1 FILLER_21_382 ();
 sg13g2_fill_1 FILLER_21_393 ();
 sg13g2_fill_1 FILLER_21_399 ();
 sg13g2_decap_8 FILLER_21_419 ();
 sg13g2_decap_4 FILLER_21_426 ();
 sg13g2_decap_8 FILLER_22_0 ();
 sg13g2_decap_8 FILLER_22_7 ();
 sg13g2_decap_8 FILLER_22_14 ();
 sg13g2_decap_8 FILLER_22_21 ();
 sg13g2_decap_8 FILLER_22_28 ();
 sg13g2_fill_1 FILLER_22_35 ();
 sg13g2_fill_2 FILLER_22_40 ();
 sg13g2_fill_1 FILLER_22_47 ();
 sg13g2_fill_2 FILLER_22_78 ();
 sg13g2_decap_4 FILLER_22_84 ();
 sg13g2_fill_2 FILLER_22_88 ();
 sg13g2_fill_2 FILLER_22_116 ();
 sg13g2_fill_1 FILLER_22_122 ();
 sg13g2_fill_1 FILLER_22_137 ();
 sg13g2_fill_2 FILLER_22_143 ();
 sg13g2_decap_4 FILLER_22_149 ();
 sg13g2_fill_2 FILLER_22_153 ();
 sg13g2_decap_8 FILLER_22_181 ();
 sg13g2_decap_8 FILLER_22_188 ();
 sg13g2_decap_8 FILLER_22_195 ();
 sg13g2_decap_8 FILLER_22_202 ();
 sg13g2_decap_8 FILLER_22_209 ();
 sg13g2_fill_2 FILLER_22_216 ();
 sg13g2_fill_1 FILLER_22_218 ();
 sg13g2_fill_1 FILLER_22_234 ();
 sg13g2_fill_1 FILLER_22_240 ();
 sg13g2_decap_4 FILLER_22_249 ();
 sg13g2_decap_8 FILLER_22_260 ();
 sg13g2_decap_4 FILLER_22_267 ();
 sg13g2_fill_2 FILLER_22_271 ();
 sg13g2_fill_1 FILLER_22_288 ();
 sg13g2_fill_1 FILLER_22_297 ();
 sg13g2_decap_4 FILLER_22_302 ();
 sg13g2_fill_1 FILLER_22_306 ();
 sg13g2_decap_8 FILLER_22_311 ();
 sg13g2_fill_1 FILLER_22_318 ();
 sg13g2_decap_8 FILLER_22_324 ();
 sg13g2_fill_1 FILLER_22_331 ();
 sg13g2_decap_8 FILLER_22_340 ();
 sg13g2_fill_2 FILLER_22_347 ();
 sg13g2_fill_1 FILLER_22_349 ();
 sg13g2_fill_2 FILLER_22_365 ();
 sg13g2_fill_1 FILLER_22_372 ();
 sg13g2_fill_2 FILLER_22_377 ();
 sg13g2_decap_8 FILLER_22_387 ();
 sg13g2_decap_8 FILLER_22_394 ();
 sg13g2_fill_1 FILLER_22_401 ();
 sg13g2_decap_8 FILLER_22_422 ();
 sg13g2_fill_1 FILLER_22_429 ();
 sg13g2_decap_8 FILLER_23_0 ();
 sg13g2_decap_8 FILLER_23_7 ();
 sg13g2_decap_8 FILLER_23_14 ();
 sg13g2_fill_2 FILLER_23_21 ();
 sg13g2_fill_2 FILLER_23_36 ();
 sg13g2_fill_1 FILLER_23_38 ();
 sg13g2_fill_1 FILLER_23_53 ();
 sg13g2_decap_8 FILLER_23_64 ();
 sg13g2_decap_8 FILLER_23_71 ();
 sg13g2_fill_1 FILLER_23_78 ();
 sg13g2_fill_2 FILLER_23_82 ();
 sg13g2_decap_4 FILLER_23_93 ();
 sg13g2_fill_1 FILLER_23_97 ();
 sg13g2_fill_2 FILLER_23_102 ();
 sg13g2_fill_1 FILLER_23_104 ();
 sg13g2_fill_2 FILLER_23_112 ();
 sg13g2_fill_1 FILLER_23_114 ();
 sg13g2_decap_8 FILLER_23_140 ();
 sg13g2_decap_4 FILLER_23_147 ();
 sg13g2_fill_2 FILLER_23_151 ();
 sg13g2_decap_8 FILLER_23_166 ();
 sg13g2_fill_2 FILLER_23_173 ();
 sg13g2_fill_1 FILLER_23_175 ();
 sg13g2_decap_8 FILLER_23_180 ();
 sg13g2_fill_1 FILLER_23_192 ();
 sg13g2_decap_8 FILLER_23_198 ();
 sg13g2_decap_4 FILLER_23_205 ();
 sg13g2_fill_1 FILLER_23_209 ();
 sg13g2_fill_1 FILLER_23_214 ();
 sg13g2_fill_2 FILLER_23_225 ();
 sg13g2_decap_4 FILLER_23_232 ();
 sg13g2_fill_2 FILLER_23_246 ();
 sg13g2_fill_1 FILLER_23_248 ();
 sg13g2_fill_1 FILLER_23_256 ();
 sg13g2_decap_8 FILLER_23_265 ();
 sg13g2_decap_8 FILLER_23_272 ();
 sg13g2_decap_4 FILLER_23_279 ();
 sg13g2_fill_1 FILLER_23_283 ();
 sg13g2_fill_2 FILLER_23_297 ();
 sg13g2_fill_1 FILLER_23_299 ();
 sg13g2_decap_4 FILLER_23_326 ();
 sg13g2_decap_8 FILLER_23_342 ();
 sg13g2_decap_8 FILLER_23_349 ();
 sg13g2_fill_2 FILLER_23_362 ();
 sg13g2_fill_1 FILLER_23_364 ();
 sg13g2_fill_2 FILLER_23_372 ();
 sg13g2_decap_8 FILLER_23_388 ();
 sg13g2_fill_2 FILLER_23_395 ();
 sg13g2_decap_8 FILLER_23_423 ();
 sg13g2_decap_8 FILLER_24_0 ();
 sg13g2_fill_2 FILLER_24_7 ();
 sg13g2_fill_1 FILLER_24_9 ();
 sg13g2_fill_2 FILLER_24_33 ();
 sg13g2_decap_4 FILLER_24_40 ();
 sg13g2_fill_1 FILLER_24_73 ();
 sg13g2_fill_1 FILLER_24_79 ();
 sg13g2_fill_2 FILLER_24_91 ();
 sg13g2_fill_1 FILLER_24_93 ();
 sg13g2_fill_1 FILLER_24_120 ();
 sg13g2_fill_1 FILLER_24_127 ();
 sg13g2_fill_2 FILLER_24_134 ();
 sg13g2_decap_8 FILLER_24_141 ();
 sg13g2_fill_2 FILLER_24_148 ();
 sg13g2_fill_1 FILLER_24_150 ();
 sg13g2_decap_8 FILLER_24_166 ();
 sg13g2_decap_8 FILLER_24_208 ();
 sg13g2_fill_2 FILLER_24_215 ();
 sg13g2_fill_1 FILLER_24_217 ();
 sg13g2_fill_2 FILLER_24_239 ();
 sg13g2_decap_8 FILLER_24_261 ();
 sg13g2_fill_2 FILLER_24_268 ();
 sg13g2_fill_1 FILLER_24_270 ();
 sg13g2_decap_4 FILLER_24_275 ();
 sg13g2_fill_2 FILLER_24_295 ();
 sg13g2_fill_1 FILLER_24_297 ();
 sg13g2_decap_8 FILLER_24_329 ();
 sg13g2_decap_4 FILLER_24_336 ();
 sg13g2_fill_1 FILLER_24_340 ();
 sg13g2_fill_1 FILLER_24_345 ();
 sg13g2_fill_2 FILLER_24_350 ();
 sg13g2_fill_1 FILLER_24_362 ();
 sg13g2_fill_1 FILLER_24_367 ();
 sg13g2_fill_1 FILLER_24_372 ();
 sg13g2_fill_2 FILLER_24_387 ();
 sg13g2_fill_1 FILLER_24_389 ();
 sg13g2_fill_2 FILLER_24_401 ();
 sg13g2_decap_8 FILLER_24_415 ();
 sg13g2_decap_8 FILLER_24_422 ();
 sg13g2_fill_1 FILLER_24_429 ();
 sg13g2_decap_8 FILLER_25_0 ();
 sg13g2_decap_4 FILLER_25_7 ();
 sg13g2_fill_1 FILLER_25_11 ();
 sg13g2_decap_4 FILLER_25_18 ();
 sg13g2_fill_2 FILLER_25_33 ();
 sg13g2_decap_4 FILLER_25_53 ();
 sg13g2_fill_1 FILLER_25_57 ();
 sg13g2_decap_4 FILLER_25_64 ();
 sg13g2_fill_2 FILLER_25_68 ();
 sg13g2_decap_4 FILLER_25_75 ();
 sg13g2_decap_4 FILLER_25_85 ();
 sg13g2_fill_2 FILLER_25_98 ();
 sg13g2_decap_8 FILLER_25_105 ();
 sg13g2_decap_8 FILLER_25_112 ();
 sg13g2_fill_1 FILLER_25_119 ();
 sg13g2_fill_2 FILLER_25_124 ();
 sg13g2_fill_2 FILLER_25_139 ();
 sg13g2_fill_1 FILLER_25_149 ();
 sg13g2_decap_4 FILLER_25_162 ();
 sg13g2_decap_8 FILLER_25_192 ();
 sg13g2_decap_8 FILLER_25_203 ();
 sg13g2_decap_8 FILLER_25_210 ();
 sg13g2_decap_8 FILLER_25_217 ();
 sg13g2_fill_2 FILLER_25_224 ();
 sg13g2_fill_2 FILLER_25_231 ();
 sg13g2_fill_1 FILLER_25_237 ();
 sg13g2_fill_2 FILLER_25_248 ();
 sg13g2_fill_1 FILLER_25_256 ();
 sg13g2_decap_8 FILLER_25_280 ();
 sg13g2_decap_8 FILLER_25_287 ();
 sg13g2_fill_1 FILLER_25_294 ();
 sg13g2_decap_4 FILLER_25_299 ();
 sg13g2_fill_1 FILLER_25_303 ();
 sg13g2_decap_4 FILLER_25_308 ();
 sg13g2_fill_1 FILLER_25_312 ();
 sg13g2_decap_8 FILLER_25_317 ();
 sg13g2_decap_8 FILLER_25_324 ();
 sg13g2_decap_8 FILLER_25_331 ();
 sg13g2_decap_4 FILLER_25_338 ();
 sg13g2_fill_1 FILLER_25_342 ();
 sg13g2_fill_1 FILLER_25_356 ();
 sg13g2_decap_8 FILLER_25_365 ();
 sg13g2_decap_8 FILLER_25_390 ();
 sg13g2_fill_2 FILLER_25_397 ();
 sg13g2_decap_8 FILLER_25_423 ();
 sg13g2_decap_8 FILLER_26_0 ();
 sg13g2_decap_8 FILLER_26_7 ();
 sg13g2_fill_2 FILLER_26_14 ();
 sg13g2_fill_1 FILLER_26_29 ();
 sg13g2_fill_2 FILLER_26_34 ();
 sg13g2_fill_1 FILLER_26_36 ();
 sg13g2_decap_4 FILLER_26_57 ();
 sg13g2_decap_4 FILLER_26_66 ();
 sg13g2_fill_1 FILLER_26_70 ();
 sg13g2_fill_2 FILLER_26_80 ();
 sg13g2_fill_1 FILLER_26_87 ();
 sg13g2_fill_2 FILLER_26_93 ();
 sg13g2_decap_8 FILLER_26_100 ();
 sg13g2_decap_4 FILLER_26_107 ();
 sg13g2_fill_1 FILLER_26_111 ();
 sg13g2_decap_4 FILLER_26_115 ();
 sg13g2_fill_2 FILLER_26_124 ();
 sg13g2_fill_2 FILLER_26_133 ();
 sg13g2_fill_2 FILLER_26_143 ();
 sg13g2_decap_4 FILLER_26_149 ();
 sg13g2_fill_1 FILLER_26_153 ();
 sg13g2_fill_2 FILLER_26_159 ();
 sg13g2_decap_8 FILLER_26_165 ();
 sg13g2_decap_8 FILLER_26_172 ();
 sg13g2_decap_8 FILLER_26_179 ();
 sg13g2_decap_4 FILLER_26_215 ();
 sg13g2_fill_1 FILLER_26_219 ();
 sg13g2_decap_8 FILLER_26_224 ();
 sg13g2_decap_8 FILLER_26_231 ();
 sg13g2_decap_8 FILLER_26_238 ();
 sg13g2_fill_1 FILLER_26_266 ();
 sg13g2_decap_8 FILLER_26_287 ();
 sg13g2_decap_8 FILLER_26_294 ();
 sg13g2_fill_1 FILLER_26_301 ();
 sg13g2_decap_8 FILLER_26_328 ();
 sg13g2_decap_8 FILLER_26_335 ();
 sg13g2_fill_1 FILLER_26_342 ();
 sg13g2_decap_8 FILLER_26_353 ();
 sg13g2_fill_1 FILLER_26_367 ();
 sg13g2_decap_4 FILLER_26_373 ();
 sg13g2_fill_1 FILLER_26_377 ();
 sg13g2_fill_2 FILLER_26_391 ();
 sg13g2_decap_4 FILLER_26_400 ();
 sg13g2_fill_2 FILLER_26_404 ();
 sg13g2_decap_8 FILLER_26_417 ();
 sg13g2_decap_4 FILLER_26_424 ();
 sg13g2_fill_2 FILLER_26_428 ();
 sg13g2_decap_8 FILLER_27_0 ();
 sg13g2_decap_4 FILLER_27_7 ();
 sg13g2_fill_2 FILLER_27_11 ();
 sg13g2_fill_1 FILLER_27_25 ();
 sg13g2_fill_1 FILLER_27_34 ();
 sg13g2_fill_2 FILLER_27_47 ();
 sg13g2_fill_1 FILLER_27_49 ();
 sg13g2_fill_2 FILLER_27_66 ();
 sg13g2_fill_2 FILLER_27_80 ();
 sg13g2_fill_1 FILLER_27_87 ();
 sg13g2_fill_2 FILLER_27_94 ();
 sg13g2_fill_1 FILLER_27_96 ();
 sg13g2_decap_4 FILLER_27_102 ();
 sg13g2_fill_2 FILLER_27_106 ();
 sg13g2_fill_1 FILLER_27_117 ();
 sg13g2_fill_1 FILLER_27_142 ();
 sg13g2_fill_2 FILLER_27_153 ();
 sg13g2_fill_1 FILLER_27_161 ();
 sg13g2_decap_8 FILLER_27_170 ();
 sg13g2_fill_2 FILLER_27_177 ();
 sg13g2_fill_2 FILLER_27_190 ();
 sg13g2_decap_8 FILLER_27_201 ();
 sg13g2_fill_1 FILLER_27_208 ();
 sg13g2_fill_2 FILLER_27_240 ();
 sg13g2_fill_1 FILLER_27_242 ();
 sg13g2_fill_1 FILLER_27_267 ();
 sg13g2_decap_8 FILLER_27_273 ();
 sg13g2_decap_8 FILLER_27_280 ();
 sg13g2_fill_2 FILLER_27_287 ();
 sg13g2_fill_1 FILLER_27_289 ();
 sg13g2_decap_8 FILLER_27_316 ();
 sg13g2_decap_4 FILLER_27_323 ();
 sg13g2_fill_2 FILLER_27_327 ();
 sg13g2_decap_8 FILLER_27_339 ();
 sg13g2_fill_2 FILLER_27_355 ();
 sg13g2_decap_4 FILLER_27_362 ();
 sg13g2_fill_1 FILLER_27_366 ();
 sg13g2_decap_4 FILLER_27_390 ();
 sg13g2_fill_1 FILLER_27_394 ();
 sg13g2_decap_4 FILLER_27_400 ();
 sg13g2_fill_2 FILLER_27_404 ();
 sg13g2_decap_8 FILLER_27_419 ();
 sg13g2_decap_4 FILLER_27_426 ();
 sg13g2_decap_8 FILLER_28_0 ();
 sg13g2_decap_4 FILLER_28_7 ();
 sg13g2_fill_1 FILLER_28_11 ();
 sg13g2_decap_4 FILLER_28_16 ();
 sg13g2_decap_4 FILLER_28_25 ();
 sg13g2_fill_2 FILLER_28_42 ();
 sg13g2_fill_1 FILLER_28_44 ();
 sg13g2_fill_2 FILLER_28_50 ();
 sg13g2_fill_1 FILLER_28_52 ();
 sg13g2_decap_4 FILLER_28_58 ();
 sg13g2_fill_1 FILLER_28_62 ();
 sg13g2_fill_2 FILLER_28_71 ();
 sg13g2_fill_1 FILLER_28_73 ();
 sg13g2_decap_8 FILLER_28_80 ();
 sg13g2_decap_8 FILLER_28_87 ();
 sg13g2_decap_8 FILLER_28_94 ();
 sg13g2_decap_8 FILLER_28_101 ();
 sg13g2_fill_1 FILLER_28_108 ();
 sg13g2_fill_2 FILLER_28_112 ();
 sg13g2_fill_1 FILLER_28_114 ();
 sg13g2_decap_4 FILLER_28_141 ();
 sg13g2_fill_2 FILLER_28_145 ();
 sg13g2_fill_2 FILLER_28_163 ();
 sg13g2_fill_1 FILLER_28_170 ();
 sg13g2_fill_2 FILLER_28_189 ();
 sg13g2_decap_4 FILLER_28_196 ();
 sg13g2_fill_2 FILLER_28_200 ();
 sg13g2_decap_4 FILLER_28_232 ();
 sg13g2_fill_1 FILLER_28_236 ();
 sg13g2_decap_8 FILLER_28_241 ();
 sg13g2_decap_8 FILLER_28_248 ();
 sg13g2_fill_2 FILLER_28_255 ();
 sg13g2_fill_1 FILLER_28_257 ();
 sg13g2_decap_8 FILLER_28_263 ();
 sg13g2_decap_4 FILLER_28_270 ();
 sg13g2_decap_8 FILLER_28_278 ();
 sg13g2_decap_8 FILLER_28_285 ();
 sg13g2_decap_8 FILLER_28_292 ();
 sg13g2_decap_8 FILLER_28_303 ();
 sg13g2_decap_8 FILLER_28_310 ();
 sg13g2_decap_8 FILLER_28_317 ();
 sg13g2_decap_8 FILLER_28_324 ();
 sg13g2_decap_4 FILLER_28_331 ();
 sg13g2_fill_1 FILLER_28_339 ();
 sg13g2_fill_1 FILLER_28_345 ();
 sg13g2_fill_1 FILLER_28_358 ();
 sg13g2_fill_1 FILLER_28_364 ();
 sg13g2_decap_8 FILLER_28_383 ();
 sg13g2_decap_8 FILLER_28_412 ();
 sg13g2_decap_8 FILLER_28_419 ();
 sg13g2_decap_4 FILLER_28_426 ();
 sg13g2_decap_4 FILLER_29_0 ();
 sg13g2_fill_1 FILLER_29_4 ();
 sg13g2_fill_2 FILLER_29_19 ();
 sg13g2_fill_2 FILLER_29_41 ();
 sg13g2_fill_1 FILLER_29_43 ();
 sg13g2_fill_1 FILLER_29_63 ();
 sg13g2_fill_2 FILLER_29_69 ();
 sg13g2_fill_2 FILLER_29_79 ();
 sg13g2_fill_2 FILLER_29_86 ();
 sg13g2_fill_1 FILLER_29_88 ();
 sg13g2_decap_8 FILLER_29_100 ();
 sg13g2_fill_2 FILLER_29_107 ();
 sg13g2_decap_8 FILLER_29_115 ();
 sg13g2_decap_8 FILLER_29_122 ();
 sg13g2_decap_4 FILLER_29_129 ();
 sg13g2_fill_1 FILLER_29_133 ();
 sg13g2_fill_2 FILLER_29_143 ();
 sg13g2_fill_2 FILLER_29_154 ();
 sg13g2_fill_1 FILLER_29_156 ();
 sg13g2_decap_4 FILLER_29_160 ();
 sg13g2_fill_2 FILLER_29_178 ();
 sg13g2_decap_4 FILLER_29_185 ();
 sg13g2_fill_1 FILLER_29_189 ();
 sg13g2_decap_8 FILLER_29_194 ();
 sg13g2_decap_8 FILLER_29_201 ();
 sg13g2_fill_2 FILLER_29_208 ();
 sg13g2_fill_2 FILLER_29_214 ();
 sg13g2_decap_8 FILLER_29_224 ();
 sg13g2_decap_8 FILLER_29_231 ();
 sg13g2_fill_1 FILLER_29_238 ();
 sg13g2_fill_1 FILLER_29_243 ();
 sg13g2_decap_8 FILLER_29_249 ();
 sg13g2_decap_8 FILLER_29_256 ();
 sg13g2_fill_2 FILLER_29_263 ();
 sg13g2_decap_4 FILLER_29_270 ();
 sg13g2_fill_2 FILLER_29_278 ();
 sg13g2_decap_8 FILLER_29_293 ();
 sg13g2_decap_8 FILLER_29_300 ();
 sg13g2_decap_8 FILLER_29_307 ();
 sg13g2_fill_2 FILLER_29_314 ();
 sg13g2_decap_4 FILLER_29_332 ();
 sg13g2_fill_1 FILLER_29_336 ();
 sg13g2_decap_8 FILLER_29_355 ();
 sg13g2_fill_2 FILLER_29_367 ();
 sg13g2_fill_1 FILLER_29_377 ();
 sg13g2_fill_1 FILLER_29_386 ();
 sg13g2_fill_2 FILLER_29_414 ();
 sg13g2_fill_1 FILLER_29_416 ();
 sg13g2_decap_8 FILLER_29_421 ();
 sg13g2_fill_2 FILLER_29_428 ();
 sg13g2_decap_8 FILLER_30_0 ();
 sg13g2_decap_4 FILLER_30_7 ();
 sg13g2_fill_1 FILLER_30_11 ();
 sg13g2_fill_1 FILLER_30_20 ();
 sg13g2_decap_4 FILLER_30_25 ();
 sg13g2_decap_8 FILLER_30_57 ();
 sg13g2_decap_8 FILLER_30_68 ();
 sg13g2_fill_2 FILLER_30_75 ();
 sg13g2_fill_1 FILLER_30_77 ();
 sg13g2_fill_2 FILLER_30_83 ();
 sg13g2_decap_8 FILLER_30_101 ();
 sg13g2_decap_4 FILLER_30_108 ();
 sg13g2_decap_4 FILLER_30_117 ();
 sg13g2_decap_4 FILLER_30_126 ();
 sg13g2_fill_2 FILLER_30_141 ();
 sg13g2_fill_2 FILLER_30_147 ();
 sg13g2_fill_1 FILLER_30_164 ();
 sg13g2_decap_4 FILLER_30_180 ();
 sg13g2_fill_1 FILLER_30_184 ();
 sg13g2_decap_8 FILLER_30_201 ();
 sg13g2_decap_8 FILLER_30_212 ();
 sg13g2_decap_8 FILLER_30_219 ();
 sg13g2_decap_4 FILLER_30_226 ();
 sg13g2_fill_2 FILLER_30_230 ();
 sg13g2_decap_4 FILLER_30_237 ();
 sg13g2_decap_4 FILLER_30_256 ();
 sg13g2_fill_2 FILLER_30_269 ();
 sg13g2_fill_2 FILLER_30_278 ();
 sg13g2_fill_2 FILLER_30_286 ();
 sg13g2_fill_1 FILLER_30_293 ();
 sg13g2_decap_8 FILLER_30_303 ();
 sg13g2_fill_2 FILLER_30_323 ();
 sg13g2_fill_1 FILLER_30_366 ();
 sg13g2_fill_2 FILLER_30_372 ();
 sg13g2_fill_1 FILLER_30_374 ();
 sg13g2_fill_1 FILLER_30_399 ();
 sg13g2_fill_1 FILLER_30_410 ();
 sg13g2_decap_8 FILLER_30_420 ();
 sg13g2_fill_2 FILLER_30_427 ();
 sg13g2_fill_1 FILLER_30_429 ();
 sg13g2_decap_8 FILLER_31_0 ();
 sg13g2_fill_1 FILLER_31_7 ();
 sg13g2_decap_4 FILLER_31_41 ();
 sg13g2_decap_8 FILLER_31_56 ();
 sg13g2_decap_8 FILLER_31_63 ();
 sg13g2_decap_4 FILLER_31_70 ();
 sg13g2_fill_1 FILLER_31_74 ();
 sg13g2_decap_4 FILLER_31_88 ();
 sg13g2_fill_2 FILLER_31_92 ();
 sg13g2_decap_8 FILLER_31_98 ();
 sg13g2_decap_8 FILLER_31_105 ();
 sg13g2_decap_4 FILLER_31_112 ();
 sg13g2_fill_2 FILLER_31_116 ();
 sg13g2_fill_1 FILLER_31_128 ();
 sg13g2_fill_1 FILLER_31_134 ();
 sg13g2_fill_1 FILLER_31_140 ();
 sg13g2_fill_2 FILLER_31_145 ();
 sg13g2_decap_4 FILLER_31_198 ();
 sg13g2_fill_1 FILLER_31_202 ();
 sg13g2_fill_1 FILLER_31_210 ();
 sg13g2_fill_1 FILLER_31_216 ();
 sg13g2_fill_2 FILLER_31_222 ();
 sg13g2_fill_2 FILLER_31_231 ();
 sg13g2_fill_2 FILLER_31_238 ();
 sg13g2_fill_1 FILLER_31_240 ();
 sg13g2_decap_8 FILLER_31_253 ();
 sg13g2_fill_2 FILLER_31_260 ();
 sg13g2_fill_1 FILLER_31_262 ();
 sg13g2_fill_1 FILLER_31_313 ();
 sg13g2_fill_1 FILLER_31_319 ();
 sg13g2_fill_1 FILLER_31_325 ();
 sg13g2_fill_1 FILLER_31_347 ();
 sg13g2_fill_1 FILLER_31_357 ();
 sg13g2_fill_2 FILLER_31_362 ();
 sg13g2_fill_2 FILLER_31_368 ();
 sg13g2_decap_4 FILLER_31_392 ();
 sg13g2_fill_1 FILLER_31_415 ();
 sg13g2_decap_8 FILLER_31_421 ();
 sg13g2_fill_2 FILLER_31_428 ();
 sg13g2_decap_8 FILLER_32_0 ();
 sg13g2_decap_8 FILLER_32_7 ();
 sg13g2_fill_1 FILLER_32_14 ();
 sg13g2_fill_2 FILLER_32_25 ();
 sg13g2_fill_1 FILLER_32_27 ();
 sg13g2_fill_2 FILLER_32_36 ();
 sg13g2_fill_2 FILLER_32_44 ();
 sg13g2_decap_4 FILLER_32_51 ();
 sg13g2_fill_1 FILLER_32_55 ();
 sg13g2_decap_8 FILLER_32_73 ();
 sg13g2_decap_8 FILLER_32_84 ();
 sg13g2_fill_2 FILLER_32_91 ();
 sg13g2_fill_1 FILLER_32_93 ();
 sg13g2_fill_2 FILLER_32_102 ();
 sg13g2_decap_8 FILLER_32_112 ();
 sg13g2_fill_1 FILLER_32_119 ();
 sg13g2_decap_4 FILLER_32_125 ();
 sg13g2_fill_2 FILLER_32_133 ();
 sg13g2_fill_1 FILLER_32_149 ();
 sg13g2_fill_1 FILLER_32_161 ();
 sg13g2_decap_8 FILLER_32_196 ();
 sg13g2_decap_8 FILLER_32_203 ();
 sg13g2_decap_8 FILLER_32_210 ();
 sg13g2_fill_2 FILLER_32_217 ();
 sg13g2_decap_4 FILLER_32_231 ();
 sg13g2_fill_2 FILLER_32_235 ();
 sg13g2_decap_4 FILLER_32_241 ();
 sg13g2_decap_4 FILLER_32_257 ();
 sg13g2_fill_2 FILLER_32_261 ();
 sg13g2_fill_1 FILLER_32_272 ();
 sg13g2_decap_8 FILLER_32_294 ();
 sg13g2_fill_1 FILLER_32_301 ();
 sg13g2_decap_8 FILLER_32_307 ();
 sg13g2_fill_1 FILLER_32_314 ();
 sg13g2_fill_1 FILLER_32_320 ();
 sg13g2_fill_1 FILLER_32_355 ();
 sg13g2_fill_1 FILLER_32_366 ();
 sg13g2_fill_1 FILLER_32_375 ();
 sg13g2_decap_8 FILLER_32_380 ();
 sg13g2_decap_4 FILLER_32_387 ();
 sg13g2_fill_2 FILLER_32_391 ();
 sg13g2_decap_8 FILLER_32_420 ();
 sg13g2_fill_2 FILLER_32_427 ();
 sg13g2_fill_1 FILLER_32_429 ();
 sg13g2_decap_8 FILLER_33_0 ();
 sg13g2_decap_4 FILLER_33_7 ();
 sg13g2_decap_4 FILLER_33_22 ();
 sg13g2_fill_1 FILLER_33_26 ();
 sg13g2_fill_2 FILLER_33_41 ();
 sg13g2_fill_2 FILLER_33_57 ();
 sg13g2_fill_1 FILLER_33_70 ();
 sg13g2_decap_8 FILLER_33_76 ();
 sg13g2_decap_8 FILLER_33_83 ();
 sg13g2_decap_8 FILLER_33_90 ();
 sg13g2_decap_8 FILLER_33_97 ();
 sg13g2_decap_8 FILLER_33_104 ();
 sg13g2_decap_4 FILLER_33_111 ();
 sg13g2_fill_2 FILLER_33_130 ();
 sg13g2_fill_1 FILLER_33_132 ();
 sg13g2_fill_2 FILLER_33_141 ();
 sg13g2_decap_4 FILLER_33_149 ();
 sg13g2_fill_2 FILLER_33_159 ();
 sg13g2_decap_4 FILLER_33_166 ();
 sg13g2_fill_2 FILLER_33_174 ();
 sg13g2_fill_1 FILLER_33_176 ();
 sg13g2_fill_2 FILLER_33_192 ();
 sg13g2_fill_2 FILLER_33_200 ();
 sg13g2_decap_4 FILLER_33_209 ();
 sg13g2_fill_1 FILLER_33_225 ();
 sg13g2_fill_2 FILLER_33_231 ();
 sg13g2_fill_1 FILLER_33_233 ();
 sg13g2_decap_4 FILLER_33_240 ();
 sg13g2_fill_2 FILLER_33_244 ();
 sg13g2_decap_4 FILLER_33_252 ();
 sg13g2_decap_4 FILLER_33_260 ();
 sg13g2_fill_2 FILLER_33_264 ();
 sg13g2_decap_4 FILLER_33_276 ();
 sg13g2_fill_1 FILLER_33_286 ();
 sg13g2_fill_2 FILLER_33_294 ();
 sg13g2_fill_1 FILLER_33_296 ();
 sg13g2_decap_4 FILLER_33_312 ();
 sg13g2_fill_2 FILLER_33_316 ();
 sg13g2_decap_8 FILLER_33_328 ();
 sg13g2_fill_2 FILLER_33_335 ();
 sg13g2_fill_1 FILLER_33_337 ();
 sg13g2_decap_8 FILLER_33_382 ();
 sg13g2_decap_8 FILLER_33_389 ();
 sg13g2_decap_4 FILLER_33_396 ();
 sg13g2_fill_2 FILLER_33_400 ();
 sg13g2_fill_1 FILLER_33_416 ();
 sg13g2_decap_8 FILLER_33_421 ();
 sg13g2_fill_2 FILLER_33_428 ();
 sg13g2_decap_8 FILLER_34_0 ();
 sg13g2_decap_8 FILLER_34_7 ();
 sg13g2_fill_1 FILLER_34_22 ();
 sg13g2_decap_4 FILLER_34_27 ();
 sg13g2_decap_4 FILLER_34_39 ();
 sg13g2_fill_1 FILLER_34_43 ();
 sg13g2_fill_1 FILLER_34_72 ();
 sg13g2_decap_4 FILLER_34_78 ();
 sg13g2_fill_1 FILLER_34_82 ();
 sg13g2_fill_1 FILLER_34_92 ();
 sg13g2_decap_8 FILLER_34_118 ();
 sg13g2_decap_4 FILLER_34_125 ();
 sg13g2_fill_1 FILLER_34_150 ();
 sg13g2_fill_1 FILLER_34_157 ();
 sg13g2_decap_4 FILLER_34_163 ();
 sg13g2_decap_4 FILLER_34_171 ();
 sg13g2_fill_1 FILLER_34_180 ();
 sg13g2_fill_1 FILLER_34_190 ();
 sg13g2_fill_2 FILLER_34_196 ();
 sg13g2_decap_8 FILLER_34_203 ();
 sg13g2_decap_8 FILLER_34_213 ();
 sg13g2_decap_8 FILLER_34_220 ();
 sg13g2_decap_8 FILLER_34_227 ();
 sg13g2_decap_4 FILLER_34_238 ();
 sg13g2_fill_2 FILLER_34_242 ();
 sg13g2_fill_1 FILLER_34_250 ();
 sg13g2_fill_2 FILLER_34_256 ();
 sg13g2_fill_2 FILLER_34_263 ();
 sg13g2_fill_2 FILLER_34_274 ();
 sg13g2_fill_2 FILLER_34_287 ();
 sg13g2_fill_1 FILLER_34_289 ();
 sg13g2_fill_1 FILLER_34_296 ();
 sg13g2_decap_8 FILLER_34_329 ();
 sg13g2_decap_8 FILLER_34_336 ();
 sg13g2_fill_1 FILLER_34_356 ();
 sg13g2_fill_1 FILLER_34_361 ();
 sg13g2_fill_2 FILLER_34_367 ();
 sg13g2_fill_1 FILLER_34_369 ();
 sg13g2_decap_8 FILLER_34_380 ();
 sg13g2_decap_8 FILLER_34_387 ();
 sg13g2_fill_1 FILLER_34_394 ();
 sg13g2_fill_2 FILLER_34_406 ();
 sg13g2_fill_1 FILLER_34_408 ();
 sg13g2_decap_8 FILLER_34_413 ();
 sg13g2_decap_8 FILLER_34_420 ();
 sg13g2_fill_2 FILLER_34_427 ();
 sg13g2_fill_1 FILLER_34_429 ();
 sg13g2_decap_8 FILLER_35_0 ();
 sg13g2_fill_2 FILLER_35_7 ();
 sg13g2_fill_2 FILLER_35_30 ();
 sg13g2_fill_1 FILLER_35_36 ();
 sg13g2_decap_8 FILLER_35_45 ();
 sg13g2_decap_8 FILLER_35_52 ();
 sg13g2_fill_1 FILLER_35_59 ();
 sg13g2_decap_8 FILLER_35_65 ();
 sg13g2_fill_2 FILLER_35_72 ();
 sg13g2_fill_1 FILLER_35_74 ();
 sg13g2_fill_2 FILLER_35_89 ();
 sg13g2_fill_1 FILLER_35_91 ();
 sg13g2_fill_1 FILLER_35_96 ();
 sg13g2_decap_8 FILLER_35_111 ();
 sg13g2_fill_1 FILLER_35_118 ();
 sg13g2_decap_4 FILLER_35_123 ();
 sg13g2_fill_1 FILLER_35_135 ();
 sg13g2_fill_2 FILLER_35_140 ();
 sg13g2_fill_1 FILLER_35_142 ();
 sg13g2_fill_1 FILLER_35_148 ();
 sg13g2_fill_1 FILLER_35_155 ();
 sg13g2_fill_1 FILLER_35_177 ();
 sg13g2_fill_2 FILLER_35_183 ();
 sg13g2_fill_2 FILLER_35_190 ();
 sg13g2_fill_2 FILLER_35_199 ();
 sg13g2_fill_1 FILLER_35_201 ();
 sg13g2_fill_2 FILLER_35_210 ();
 sg13g2_fill_1 FILLER_35_212 ();
 sg13g2_decap_4 FILLER_35_226 ();
 sg13g2_decap_8 FILLER_35_234 ();
 sg13g2_decap_4 FILLER_35_241 ();
 sg13g2_fill_1 FILLER_35_245 ();
 sg13g2_decap_4 FILLER_35_250 ();
 sg13g2_fill_2 FILLER_35_254 ();
 sg13g2_fill_2 FILLER_35_260 ();
 sg13g2_fill_1 FILLER_35_262 ();
 sg13g2_fill_2 FILLER_35_271 ();
 sg13g2_fill_1 FILLER_35_273 ();
 sg13g2_fill_2 FILLER_35_285 ();
 sg13g2_fill_1 FILLER_35_287 ();
 sg13g2_fill_1 FILLER_35_293 ();
 sg13g2_fill_1 FILLER_35_302 ();
 sg13g2_fill_1 FILLER_35_309 ();
 sg13g2_fill_2 FILLER_35_315 ();
 sg13g2_decap_4 FILLER_35_334 ();
 sg13g2_fill_2 FILLER_35_354 ();
 sg13g2_fill_1 FILLER_35_356 ();
 sg13g2_fill_1 FILLER_35_362 ();
 sg13g2_decap_8 FILLER_35_388 ();
 sg13g2_fill_2 FILLER_35_395 ();
 sg13g2_fill_1 FILLER_35_410 ();
 sg13g2_decap_4 FILLER_35_424 ();
 sg13g2_fill_2 FILLER_35_428 ();
 sg13g2_decap_8 FILLER_36_0 ();
 sg13g2_fill_2 FILLER_36_7 ();
 sg13g2_fill_1 FILLER_36_9 ();
 sg13g2_fill_2 FILLER_36_15 ();
 sg13g2_fill_1 FILLER_36_44 ();
 sg13g2_fill_2 FILLER_36_50 ();
 sg13g2_fill_1 FILLER_36_52 ();
 sg13g2_fill_1 FILLER_36_59 ();
 sg13g2_fill_2 FILLER_36_65 ();
 sg13g2_decap_4 FILLER_36_116 ();
 sg13g2_fill_1 FILLER_36_120 ();
 sg13g2_decap_4 FILLER_36_125 ();
 sg13g2_fill_2 FILLER_36_129 ();
 sg13g2_fill_2 FILLER_36_136 ();
 sg13g2_fill_1 FILLER_36_138 ();
 sg13g2_decap_4 FILLER_36_160 ();
 sg13g2_fill_2 FILLER_36_169 ();
 sg13g2_decap_8 FILLER_36_200 ();
 sg13g2_decap_8 FILLER_36_207 ();
 sg13g2_decap_8 FILLER_36_214 ();
 sg13g2_decap_4 FILLER_36_221 ();
 sg13g2_fill_2 FILLER_36_225 ();
 sg13g2_decap_4 FILLER_36_237 ();
 sg13g2_fill_1 FILLER_36_241 ();
 sg13g2_decap_8 FILLER_36_250 ();
 sg13g2_fill_1 FILLER_36_257 ();
 sg13g2_fill_2 FILLER_36_263 ();
 sg13g2_fill_1 FILLER_36_265 ();
 sg13g2_fill_1 FILLER_36_269 ();
 sg13g2_decap_8 FILLER_36_278 ();
 sg13g2_decap_8 FILLER_36_285 ();
 sg13g2_fill_2 FILLER_36_292 ();
 sg13g2_decap_4 FILLER_36_309 ();
 sg13g2_fill_1 FILLER_36_317 ();
 sg13g2_fill_1 FILLER_36_323 ();
 sg13g2_decap_4 FILLER_36_337 ();
 sg13g2_fill_1 FILLER_36_341 ();
 sg13g2_decap_8 FILLER_36_348 ();
 sg13g2_decap_8 FILLER_36_360 ();
 sg13g2_decap_8 FILLER_36_367 ();
 sg13g2_fill_2 FILLER_36_374 ();
 sg13g2_decap_8 FILLER_36_380 ();
 sg13g2_decap_8 FILLER_36_387 ();
 sg13g2_decap_8 FILLER_36_394 ();
 sg13g2_fill_1 FILLER_36_413 ();
 sg13g2_decap_8 FILLER_36_423 ();
 sg13g2_fill_2 FILLER_37_0 ();
 sg13g2_fill_1 FILLER_37_2 ();
 sg13g2_decap_4 FILLER_37_26 ();
 sg13g2_fill_1 FILLER_37_30 ();
 sg13g2_fill_1 FILLER_37_54 ();
 sg13g2_fill_2 FILLER_37_67 ();
 sg13g2_decap_4 FILLER_37_75 ();
 sg13g2_fill_1 FILLER_37_79 ();
 sg13g2_decap_4 FILLER_37_85 ();
 sg13g2_decap_8 FILLER_37_107 ();
 sg13g2_decap_4 FILLER_37_114 ();
 sg13g2_fill_2 FILLER_37_127 ();
 sg13g2_fill_1 FILLER_37_129 ();
 sg13g2_fill_1 FILLER_37_141 ();
 sg13g2_decap_8 FILLER_37_147 ();
 sg13g2_fill_2 FILLER_37_154 ();
 sg13g2_fill_1 FILLER_37_156 ();
 sg13g2_fill_2 FILLER_37_162 ();
 sg13g2_fill_2 FILLER_37_177 ();
 sg13g2_fill_1 FILLER_37_184 ();
 sg13g2_fill_2 FILLER_37_189 ();
 sg13g2_fill_1 FILLER_37_191 ();
 sg13g2_fill_1 FILLER_37_202 ();
 sg13g2_fill_2 FILLER_37_207 ();
 sg13g2_fill_1 FILLER_37_209 ();
 sg13g2_fill_2 FILLER_37_214 ();
 sg13g2_fill_2 FILLER_37_235 ();
 sg13g2_fill_1 FILLER_37_289 ();
 sg13g2_fill_1 FILLER_37_295 ();
 sg13g2_decap_4 FILLER_37_300 ();
 sg13g2_fill_2 FILLER_37_304 ();
 sg13g2_fill_2 FILLER_37_311 ();
 sg13g2_fill_1 FILLER_37_364 ();
 sg13g2_decap_4 FILLER_37_370 ();
 sg13g2_decap_8 FILLER_37_378 ();
 sg13g2_decap_8 FILLER_37_385 ();
 sg13g2_decap_8 FILLER_37_392 ();
 sg13g2_decap_4 FILLER_37_399 ();
 sg13g2_fill_2 FILLER_37_403 ();
 sg13g2_fill_1 FILLER_37_409 ();
 sg13g2_decap_8 FILLER_37_423 ();
 sg13g2_decap_8 FILLER_38_0 ();
 sg13g2_decap_8 FILLER_38_7 ();
 sg13g2_decap_8 FILLER_38_14 ();
 sg13g2_fill_1 FILLER_38_21 ();
 sg13g2_decap_8 FILLER_38_32 ();
 sg13g2_decap_8 FILLER_38_39 ();
 sg13g2_decap_8 FILLER_38_46 ();
 sg13g2_decap_8 FILLER_38_53 ();
 sg13g2_decap_8 FILLER_38_60 ();
 sg13g2_fill_2 FILLER_38_67 ();
 sg13g2_decap_4 FILLER_38_93 ();
 sg13g2_fill_1 FILLER_38_133 ();
 sg13g2_decap_8 FILLER_38_139 ();
 sg13g2_fill_2 FILLER_38_155 ();
 sg13g2_decap_8 FILLER_38_166 ();
 sg13g2_decap_8 FILLER_38_173 ();
 sg13g2_fill_2 FILLER_38_184 ();
 sg13g2_fill_2 FILLER_38_192 ();
 sg13g2_fill_1 FILLER_38_194 ();
 sg13g2_decap_4 FILLER_38_203 ();
 sg13g2_fill_2 FILLER_38_214 ();
 sg13g2_fill_1 FILLER_38_216 ();
 sg13g2_fill_1 FILLER_38_221 ();
 sg13g2_fill_1 FILLER_38_239 ();
 sg13g2_fill_2 FILLER_38_244 ();
 sg13g2_decap_8 FILLER_38_275 ();
 sg13g2_decap_8 FILLER_38_282 ();
 sg13g2_decap_8 FILLER_38_289 ();
 sg13g2_decap_8 FILLER_38_296 ();
 sg13g2_decap_4 FILLER_38_303 ();
 sg13g2_fill_1 FILLER_38_307 ();
 sg13g2_decap_8 FILLER_38_312 ();
 sg13g2_decap_4 FILLER_38_319 ();
 sg13g2_fill_1 FILLER_38_329 ();
 sg13g2_fill_1 FILLER_38_378 ();
 sg13g2_fill_1 FILLER_38_387 ();
 sg13g2_decap_8 FILLER_38_393 ();
 sg13g2_fill_2 FILLER_38_400 ();
 sg13g2_fill_1 FILLER_38_402 ();
 sg13g2_fill_2 FILLER_38_413 ();
 sg13g2_fill_1 FILLER_38_415 ();
 sg13g2_decap_8 FILLER_38_423 ();
endmodule
