module tt_um_htfab_rotfpga2_ff (clk,
    ena,
    rst_n,
    ui_in,
    uio_in,
    uio_oe,
    uio_out,
    uo_out);
 input clk;
 input ena;
 input rst_n;
 input [7:0] ui_in;
 input [7:0] uio_in;
 output [7:0] uio_oe;
 output [7:0] uio_out;
 output [7:0] uo_out;

 wire _0000_;
 wire _0001_;
 wire _0002_;
 wire _0003_;
 wire _0004_;
 wire _0005_;
 wire _0006_;
 wire _0007_;
 wire _0008_;
 wire _0009_;
 wire _0010_;
 wire _0011_;
 wire _0012_;
 wire _0013_;
 wire _0014_;
 wire _0015_;
 wire _0016_;
 wire _0017_;
 wire _0018_;
 wire _0019_;
 wire _0020_;
 wire _0021_;
 wire _0022_;
 wire _0023_;
 wire _0024_;
 wire _0025_;
 wire _0026_;
 wire _0027_;
 wire _0028_;
 wire _0029_;
 wire _0030_;
 wire _0031_;
 wire _0032_;
 wire _0033_;
 wire _0034_;
 wire _0035_;
 wire _0036_;
 wire _0037_;
 wire _0038_;
 wire _0039_;
 wire _0040_;
 wire _0041_;
 wire _0042_;
 wire _0043_;
 wire _0044_;
 wire _0045_;
 wire _0046_;
 wire _0047_;
 wire _0048_;
 wire _0049_;
 wire _0050_;
 wire _0051_;
 wire _0052_;
 wire _0053_;
 wire _0054_;
 wire _0055_;
 wire _0056_;
 wire _0057_;
 wire _0058_;
 wire _0059_;
 wire _0060_;
 wire _0061_;
 wire _0062_;
 wire _0063_;
 wire _0064_;
 wire _0065_;
 wire _0066_;
 wire _0067_;
 wire _0068_;
 wire _0069_;
 wire _0070_;
 wire _0071_;
 wire _0072_;
 wire _0073_;
 wire _0074_;
 wire _0075_;
 wire _0076_;
 wire _0077_;
 wire _0078_;
 wire _0079_;
 wire _0080_;
 wire _0081_;
 wire _0082_;
 wire _0083_;
 wire _0084_;
 wire _0085_;
 wire _0086_;
 wire _0087_;
 wire _0088_;
 wire _0089_;
 wire _0090_;
 wire _0091_;
 wire _0092_;
 wire _0093_;
 wire _0094_;
 wire _0095_;
 wire _0096_;
 wire _0097_;
 wire _0098_;
 wire _0099_;
 wire _0100_;
 wire _0101_;
 wire _0102_;
 wire _0103_;
 wire _0104_;
 wire _0105_;
 wire _0106_;
 wire _0107_;
 wire _0108_;
 wire _0109_;
 wire _0110_;
 wire _0111_;
 wire _0112_;
 wire _0113_;
 wire _0114_;
 wire _0115_;
 wire _0116_;
 wire _0117_;
 wire _0118_;
 wire _0119_;
 wire _0120_;
 wire _0121_;
 wire _0122_;
 wire _0123_;
 wire _0124_;
 wire _0125_;
 wire _0126_;
 wire _0127_;
 wire _0128_;
 wire _0129_;
 wire _0130_;
 wire _0131_;
 wire _0132_;
 wire _0133_;
 wire _0134_;
 wire _0135_;
 wire _0136_;
 wire _0137_;
 wire _0138_;
 wire _0139_;
 wire _0140_;
 wire _0141_;
 wire _0142_;
 wire _0143_;
 wire _0144_;
 wire _0145_;
 wire _0146_;
 wire _0147_;
 wire _0148_;
 wire _0149_;
 wire _0150_;
 wire _0151_;
 wire _0152_;
 wire _0153_;
 wire _0154_;
 wire _0155_;
 wire _0156_;
 wire _0157_;
 wire _0158_;
 wire _0159_;
 wire _0160_;
 wire _0161_;
 wire _0162_;
 wire _0163_;
 wire _0164_;
 wire _0165_;
 wire _0166_;
 wire _0167_;
 wire _0168_;
 wire _0169_;
 wire _0170_;
 wire _0171_;
 wire _0172_;
 wire _0173_;
 wire _0174_;
 wire _0175_;
 wire _0176_;
 wire _0177_;
 wire _0178_;
 wire _0179_;
 wire _0180_;
 wire _0181_;
 wire _0182_;
 wire _0183_;
 wire _0184_;
 wire _0185_;
 wire _0186_;
 wire _0187_;
 wire _0188_;
 wire _0189_;
 wire _0190_;
 wire _0191_;
 wire _0192_;
 wire _0193_;
 wire _0194_;
 wire _0195_;
 wire _0196_;
 wire _0197_;
 wire _0198_;
 wire _0199_;
 wire _0200_;
 wire _0201_;
 wire _0202_;
 wire _0203_;
 wire _0204_;
 wire _0205_;
 wire _0206_;
 wire _0207_;
 wire _0208_;
 wire _0209_;
 wire _0210_;
 wire _0211_;
 wire _0212_;
 wire _0213_;
 wire _0214_;
 wire _0215_;
 wire _0216_;
 wire _0217_;
 wire _0218_;
 wire _0219_;
 wire _0220_;
 wire _0221_;
 wire _0222_;
 wire _0223_;
 wire _0224_;
 wire _0225_;
 wire _0226_;
 wire _0227_;
 wire _0228_;
 wire _0229_;
 wire _0230_;
 wire _0231_;
 wire _0232_;
 wire _0233_;
 wire _0234_;
 wire _0235_;
 wire _0236_;
 wire _0237_;
 wire _0238_;
 wire _0239_;
 wire _0240_;
 wire _0241_;
 wire _0242_;
 wire _0243_;
 wire _0244_;
 wire _0245_;
 wire _0246_;
 wire _0247_;
 wire _0248_;
 wire _0249_;
 wire _0250_;
 wire _0251_;
 wire _0252_;
 wire _0253_;
 wire _0254_;
 wire _0255_;
 wire _0256_;
 wire _0257_;
 wire _0258_;
 wire _0259_;
 wire _0260_;
 wire _0261_;
 wire _0262_;
 wire _0263_;
 wire _0264_;
 wire _0265_;
 wire _0266_;
 wire _0267_;
 wire _0268_;
 wire _0269_;
 wire _0270_;
 wire _0271_;
 wire _0272_;
 wire _0273_;
 wire _0274_;
 wire _0275_;
 wire _0276_;
 wire _0277_;
 wire _0278_;
 wire _0279_;
 wire _0280_;
 wire _0281_;
 wire _0282_;
 wire _0283_;
 wire _0284_;
 wire _0285_;
 wire _0286_;
 wire _0287_;
 wire _0288_;
 wire _0289_;
 wire _0290_;
 wire _0291_;
 wire _0292_;
 wire _0293_;
 wire _0294_;
 wire _0295_;
 wire _0296_;
 wire _0297_;
 wire _0298_;
 wire _0299_;
 wire _0300_;
 wire _0301_;
 wire _0302_;
 wire _0303_;
 wire _0304_;
 wire _0305_;
 wire _0306_;
 wire _0307_;
 wire _0308_;
 wire _0309_;
 wire _0310_;
 wire _0311_;
 wire _0312_;
 wire _0313_;
 wire _0314_;
 wire _0315_;
 wire _0316_;
 wire _0317_;
 wire _0318_;
 wire _0319_;
 wire _0320_;
 wire _0321_;
 wire _0322_;
 wire _0323_;
 wire _0324_;
 wire _0325_;
 wire _0326_;
 wire _0327_;
 wire _0328_;
 wire _0329_;
 wire _0330_;
 wire _0331_;
 wire _0332_;
 wire _0333_;
 wire _0334_;
 wire _0335_;
 wire _0336_;
 wire _0337_;
 wire _0338_;
 wire _0339_;
 wire _0340_;
 wire _0341_;
 wire _0342_;
 wire _0343_;
 wire _0344_;
 wire _0345_;
 wire _0346_;
 wire _0347_;
 wire _0348_;
 wire _0349_;
 wire _0350_;
 wire _0351_;
 wire _0352_;
 wire _0353_;
 wire _0354_;
 wire _0355_;
 wire _0356_;
 wire _0357_;
 wire _0358_;
 wire _0359_;
 wire _0360_;
 wire _0361_;
 wire _0362_;
 wire _0363_;
 wire _0364_;
 wire _0365_;
 wire _0366_;
 wire _0367_;
 wire _0368_;
 wire _0369_;
 wire _0370_;
 wire _0371_;
 wire _0372_;
 wire _0373_;
 wire _0374_;
 wire _0375_;
 wire _0376_;
 wire _0377_;
 wire _0378_;
 wire _0379_;
 wire _0380_;
 wire _0381_;
 wire _0382_;
 wire _0383_;
 wire _0384_;
 wire _0385_;
 wire _0386_;
 wire _0387_;
 wire _0388_;
 wire _0389_;
 wire _0390_;
 wire _0391_;
 wire _0392_;
 wire _0393_;
 wire _0394_;
 wire _0395_;
 wire _0396_;
 wire _0397_;
 wire _0398_;
 wire _0399_;
 wire _0400_;
 wire _0401_;
 wire _0402_;
 wire _0403_;
 wire _0404_;
 wire _0405_;
 wire _0406_;
 wire _0407_;
 wire _0408_;
 wire _0409_;
 wire _0410_;
 wire _0411_;
 wire _0412_;
 wire _0413_;
 wire _0414_;
 wire _0415_;
 wire _0416_;
 wire _0417_;
 wire _0418_;
 wire _0419_;
 wire _0420_;
 wire _0421_;
 wire _0422_;
 wire _0423_;
 wire _0424_;
 wire _0425_;
 wire _0426_;
 wire _0427_;
 wire _0428_;
 wire _0429_;
 wire _0430_;
 wire _0431_;
 wire _0432_;
 wire _0433_;
 wire _0434_;
 wire _0435_;
 wire _0436_;
 wire _0437_;
 wire _0438_;
 wire _0439_;
 wire _0440_;
 wire _0441_;
 wire _0442_;
 wire _0443_;
 wire _0444_;
 wire _0445_;
 wire _0446_;
 wire _0447_;
 wire _0448_;
 wire _0449_;
 wire _0450_;
 wire _0451_;
 wire _0452_;
 wire _0453_;
 wire _0454_;
 wire _0455_;
 wire _0456_;
 wire _0457_;
 wire _0458_;
 wire _0459_;
 wire _0460_;
 wire _0461_;
 wire _0462_;
 wire _0463_;
 wire _0464_;
 wire _0465_;
 wire _0466_;
 wire _0467_;
 wire _0468_;
 wire _0469_;
 wire _0470_;
 wire _0471_;
 wire _0472_;
 wire _0473_;
 wire _0474_;
 wire _0475_;
 wire _0476_;
 wire _0477_;
 wire _0478_;
 wire _0479_;
 wire _0480_;
 wire _0481_;
 wire _0482_;
 wire _0483_;
 wire _0484_;
 wire _0485_;
 wire _0486_;
 wire _0487_;
 wire _0488_;
 wire _0489_;
 wire _0490_;
 wire _0491_;
 wire _0492_;
 wire _0493_;
 wire _0494_;
 wire _0495_;
 wire _0496_;
 wire _0497_;
 wire _0498_;
 wire _0499_;
 wire _0500_;
 wire _0501_;
 wire _0502_;
 wire _0503_;
 wire _0504_;
 wire _0505_;
 wire _0506_;
 wire _0507_;
 wire _0508_;
 wire _0509_;
 wire _0510_;
 wire _0511_;
 wire _0512_;
 wire _0513_;
 wire _0514_;
 wire _0515_;
 wire _0516_;
 wire _0517_;
 wire _0518_;
 wire _0519_;
 wire _0520_;
 wire _0521_;
 wire _0522_;
 wire _0523_;
 wire _0524_;
 wire _0525_;
 wire _0526_;
 wire _0527_;
 wire _0528_;
 wire _0529_;
 wire _0530_;
 wire _0531_;
 wire _0532_;
 wire _0533_;
 wire _0534_;
 wire _0535_;
 wire _0536_;
 wire _0537_;
 wire _0538_;
 wire _0539_;
 wire _0540_;
 wire _0541_;
 wire _0542_;
 wire _0543_;
 wire _0544_;
 wire _0545_;
 wire _0546_;
 wire _0547_;
 wire _0548_;
 wire _0549_;
 wire _0550_;
 wire _0551_;
 wire _0552_;
 wire _0553_;
 wire _0554_;
 wire _0555_;
 wire _0556_;
 wire _0557_;
 wire _0558_;
 wire _0559_;
 wire _0560_;
 wire _0561_;
 wire _0562_;
 wire _0563_;
 wire _0564_;
 wire _0565_;
 wire _0566_;
 wire _0567_;
 wire _0568_;
 wire _0569_;
 wire _0570_;
 wire _0571_;
 wire _0572_;
 wire _0573_;
 wire _0574_;
 wire _0575_;
 wire _0576_;
 wire _0577_;
 wire _0578_;
 wire _0579_;
 wire _0580_;
 wire _0581_;
 wire _0582_;
 wire _0583_;
 wire _0584_;
 wire _0585_;
 wire _0586_;
 wire _0587_;
 wire _0588_;
 wire _0589_;
 wire _0590_;
 wire _0591_;
 wire _0592_;
 wire _0593_;
 wire _0594_;
 wire _0595_;
 wire _0596_;
 wire _0597_;
 wire _0598_;
 wire _0599_;
 wire _0600_;
 wire _0601_;
 wire _0602_;
 wire _0603_;
 wire _0604_;
 wire _0605_;
 wire _0606_;
 wire _0607_;
 wire _0608_;
 wire _0609_;
 wire _0610_;
 wire _0611_;
 wire _0612_;
 wire _0613_;
 wire _0614_;
 wire _0615_;
 wire _0616_;
 wire _0617_;
 wire _0618_;
 wire _0619_;
 wire _0620_;
 wire _0621_;
 wire _0622_;
 wire _0623_;
 wire _0624_;
 wire _0625_;
 wire _0626_;
 wire _0627_;
 wire _0628_;
 wire _0629_;
 wire _0630_;
 wire _0631_;
 wire _0632_;
 wire _0633_;
 wire _0634_;
 wire _0635_;
 wire _0636_;
 wire _0637_;
 wire _0638_;
 wire _0639_;
 wire _0640_;
 wire _0641_;
 wire _0642_;
 wire _0643_;
 wire _0644_;
 wire _0645_;
 wire _0646_;
 wire _0647_;
 wire _0648_;
 wire _0649_;
 wire _0650_;
 wire _0651_;
 wire _0652_;
 wire _0653_;
 wire _0654_;
 wire _0655_;
 wire _0656_;
 wire _0657_;
 wire _0658_;
 wire _0659_;
 wire _0660_;
 wire _0661_;
 wire _0662_;
 wire _0663_;
 wire _0664_;
 wire _0665_;
 wire _0666_;
 wire _0667_;
 wire _0668_;
 wire _0669_;
 wire _0670_;
 wire _0671_;
 wire _0672_;
 wire _0673_;
 wire _0674_;
 wire _0675_;
 wire _0676_;
 wire _0677_;
 wire _0678_;
 wire _0679_;
 wire _0680_;
 wire _0681_;
 wire _0682_;
 wire _0683_;
 wire _0684_;
 wire _0685_;
 wire _0686_;
 wire _0687_;
 wire _0688_;
 wire _0689_;
 wire _0690_;
 wire _0691_;
 wire _0692_;
 wire _0693_;
 wire _0694_;
 wire _0695_;
 wire _0696_;
 wire _0697_;
 wire _0698_;
 wire _0699_;
 wire _0700_;
 wire _0701_;
 wire _0702_;
 wire _0703_;
 wire _0704_;
 wire _0705_;
 wire _0706_;
 wire _0707_;
 wire _0708_;
 wire _0709_;
 wire _0710_;
 wire _0711_;
 wire _0712_;
 wire _0713_;
 wire _0714_;
 wire _0715_;
 wire _0716_;
 wire _0717_;
 wire _0718_;
 wire _0719_;
 wire _0720_;
 wire _0721_;
 wire _0722_;
 wire _0723_;
 wire _0724_;
 wire _0725_;
 wire _0726_;
 wire _0727_;
 wire _0728_;
 wire _0729_;
 wire _0730_;
 wire _0731_;
 wire _0732_;
 wire _0733_;
 wire _0734_;
 wire _0735_;
 wire _0736_;
 wire _0737_;
 wire _0738_;
 wire _0739_;
 wire _0740_;
 wire _0741_;
 wire _0742_;
 wire _0743_;
 wire _0744_;
 wire _0745_;
 wire _0746_;
 wire _0747_;
 wire _0748_;
 wire _0749_;
 wire _0750_;
 wire _0751_;
 wire _0752_;
 wire _0753_;
 wire _0754_;
 wire _0755_;
 wire _0756_;
 wire _0757_;
 wire _0758_;
 wire _0759_;
 wire _0760_;
 wire _0761_;
 wire _0762_;
 wire _0763_;
 wire _0764_;
 wire _0765_;
 wire _0766_;
 wire _0767_;
 wire _0768_;
 wire _0769_;
 wire _0770_;
 wire _0771_;
 wire _0772_;
 wire _0773_;
 wire _0774_;
 wire _0775_;
 wire _0776_;
 wire _0777_;
 wire _0778_;
 wire _0779_;
 wire _0780_;
 wire _0781_;
 wire _0782_;
 wire _0783_;
 wire _0784_;
 wire _0785_;
 wire _0786_;
 wire _0787_;
 wire _0788_;
 wire _0789_;
 wire _0790_;
 wire _0791_;
 wire _0792_;
 wire _0793_;
 wire _0794_;
 wire _0795_;
 wire _0796_;
 wire _0797_;
 wire _0798_;
 wire _0799_;
 wire _0800_;
 wire _0801_;
 wire _0802_;
 wire _0803_;
 wire _0804_;
 wire _0805_;
 wire _0806_;
 wire _0807_;
 wire _0808_;
 wire _0809_;
 wire _0810_;
 wire _0811_;
 wire _0812_;
 wire _0813_;
 wire _0814_;
 wire _0815_;
 wire _0816_;
 wire _0817_;
 wire _0818_;
 wire _0819_;
 wire _0820_;
 wire _0821_;
 wire _0822_;
 wire _0823_;
 wire _0824_;
 wire _0825_;
 wire _0826_;
 wire _0827_;
 wire _0828_;
 wire _0829_;
 wire _0830_;
 wire _0831_;
 wire _0832_;
 wire _0833_;
 wire _0834_;
 wire _0835_;
 wire _0836_;
 wire _0837_;
 wire _0838_;
 wire _0839_;
 wire _0840_;
 wire _0841_;
 wire _0842_;
 wire _0843_;
 wire _0844_;
 wire _0845_;
 wire _0846_;
 wire _0847_;
 wire _0848_;
 wire _0849_;
 wire _0850_;
 wire _0851_;
 wire _0852_;
 wire _0853_;
 wire _0854_;
 wire _0855_;
 wire _0856_;
 wire _0857_;
 wire _0858_;
 wire _0859_;
 wire _0860_;
 wire _0861_;
 wire _0862_;
 wire _0863_;
 wire _0864_;
 wire _0865_;
 wire _0866_;
 wire _0867_;
 wire _0868_;
 wire _0869_;
 wire _0870_;
 wire _0871_;
 wire _0872_;
 wire _0873_;
 wire _0874_;
 wire _0875_;
 wire _0876_;
 wire _0877_;
 wire _0878_;
 wire _0879_;
 wire _0880_;
 wire _0881_;
 wire _0882_;
 wire _0883_;
 wire _0884_;
 wire _0885_;
 wire _0886_;
 wire _0887_;
 wire _0888_;
 wire _0889_;
 wire _0890_;
 wire _0891_;
 wire _0892_;
 wire _0893_;
 wire _0894_;
 wire _0895_;
 wire _0896_;
 wire _0897_;
 wire _0898_;
 wire _0899_;
 wire _0900_;
 wire _0901_;
 wire _0902_;
 wire _0903_;
 wire _0904_;
 wire _0905_;
 wire _0906_;
 wire _0907_;
 wire _0908_;
 wire _0909_;
 wire _0910_;
 wire _0911_;
 wire _0912_;
 wire _0913_;
 wire _0914_;
 wire _0915_;
 wire _0916_;
 wire _0917_;
 wire _0918_;
 wire _0919_;
 wire _0920_;
 wire _0921_;
 wire _0922_;
 wire _0923_;
 wire _0924_;
 wire _0925_;
 wire _0926_;
 wire _0927_;
 wire _0928_;
 wire _0929_;
 wire _0930_;
 wire _0931_;
 wire _0932_;
 wire _0933_;
 wire _0934_;
 wire _0935_;
 wire _0936_;
 wire _0937_;
 wire _0938_;
 wire _0939_;
 wire _0940_;
 wire _0941_;
 wire _0942_;
 wire _0943_;
 wire _0944_;
 wire _0945_;
 wire _0946_;
 wire _0947_;
 wire _0948_;
 wire _0949_;
 wire _0950_;
 wire _0951_;
 wire _0952_;
 wire _0953_;
 wire _0954_;
 wire _0955_;
 wire _0956_;
 wire _0957_;
 wire _0958_;
 wire _0959_;
 wire _0960_;
 wire _0961_;
 wire _0962_;
 wire _0963_;
 wire _0964_;
 wire _0965_;
 wire _0966_;
 wire _0967_;
 wire _0968_;
 wire _0969_;
 wire _0970_;
 wire _0971_;
 wire _0972_;
 wire _0973_;
 wire _0974_;
 wire _0975_;
 wire _0976_;
 wire _0977_;
 wire _0978_;
 wire _0979_;
 wire _0980_;
 wire _0981_;
 wire _0982_;
 wire _0983_;
 wire _0984_;
 wire _0985_;
 wire _0986_;
 wire _0987_;
 wire _0988_;
 wire _0989_;
 wire _0990_;
 wire _0991_;
 wire _0992_;
 wire _0993_;
 wire _0994_;
 wire _0995_;
 wire _0996_;
 wire _0997_;
 wire _0998_;
 wire _0999_;
 wire _1000_;
 wire _1001_;
 wire _1002_;
 wire _1003_;
 wire _1004_;
 wire _1005_;
 wire _1006_;
 wire _1007_;
 wire _1008_;
 wire _1009_;
 wire _1010_;
 wire _1011_;
 wire _1012_;
 wire _1013_;
 wire _1014_;
 wire _1015_;
 wire _1016_;
 wire _1017_;
 wire _1018_;
 wire _1019_;
 wire _1020_;
 wire _1021_;
 wire _1022_;
 wire _1023_;
 wire _1024_;
 wire _1025_;
 wire _1026_;
 wire _1027_;
 wire _1028_;
 wire _1029_;
 wire _1030_;
 wire _1031_;
 wire _1032_;
 wire _1033_;
 wire _1034_;
 wire _1035_;
 wire _1036_;
 wire _1037_;
 wire _1038_;
 wire _1039_;
 wire _1040_;
 wire _1041_;
 wire _1042_;
 wire _1043_;
 wire _1044_;
 wire _1045_;
 wire _1046_;
 wire _1047_;
 wire _1048_;
 wire _1049_;
 wire _1050_;
 wire _1051_;
 wire _1052_;
 wire _1053_;
 wire _1054_;
 wire _1055_;
 wire _1056_;
 wire _1057_;
 wire _1058_;
 wire _1059_;
 wire _1060_;
 wire _1061_;
 wire _1062_;
 wire _1063_;
 wire _1064_;
 wire _1065_;
 wire _1066_;
 wire _1067_;
 wire _1068_;
 wire _1069_;
 wire _1070_;
 wire _1071_;
 wire _1072_;
 wire _1073_;
 wire _1074_;
 wire _1075_;
 wire _1076_;
 wire _1077_;
 wire _1078_;
 wire _1079_;
 wire _1080_;
 wire _1081_;
 wire _1082_;
 wire _1083_;
 wire _1084_;
 wire _1085_;
 wire _1086_;
 wire _1087_;
 wire _1088_;
 wire _1089_;
 wire _1090_;
 wire _1091_;
 wire _1092_;
 wire _1093_;
 wire _1094_;
 wire _1095_;
 wire _1096_;
 wire _1097_;
 wire _1098_;
 wire _1099_;
 wire _1100_;
 wire _1101_;
 wire _1102_;
 wire _1103_;
 wire _1104_;
 wire _1105_;
 wire _1106_;
 wire _1107_;
 wire _1108_;
 wire _1109_;
 wire _1110_;
 wire _1111_;
 wire _1112_;
 wire _1113_;
 wire _1114_;
 wire _1115_;
 wire _1116_;
 wire _1117_;
 wire _1118_;
 wire _1119_;
 wire _1120_;
 wire _1121_;
 wire _1122_;
 wire _1123_;
 wire _1124_;
 wire _1125_;
 wire _1126_;
 wire _1127_;
 wire _1128_;
 wire _1129_;
 wire _1130_;
 wire _1131_;
 wire _1132_;
 wire _1133_;
 wire _1134_;
 wire _1135_;
 wire _1136_;
 wire _1137_;
 wire _1138_;
 wire _1139_;
 wire _1140_;
 wire _1141_;
 wire _1142_;
 wire _1143_;
 wire _1144_;
 wire _1145_;
 wire _1146_;
 wire _1147_;
 wire _1148_;
 wire _1149_;
 wire _1150_;
 wire _1151_;
 wire _1152_;
 wire _1153_;
 wire _1154_;
 wire _1155_;
 wire _1156_;
 wire _1157_;
 wire _1158_;
 wire _1159_;
 wire _1160_;
 wire _1161_;
 wire _1162_;
 wire _1163_;
 wire _1164_;
 wire _1165_;
 wire _1166_;
 wire _1167_;
 wire _1168_;
 wire _1169_;
 wire _1170_;
 wire _1171_;
 wire _1172_;
 wire _1173_;
 wire _1174_;
 wire _1175_;
 wire _1176_;
 wire _1177_;
 wire _1178_;
 wire _1179_;
 wire _1180_;
 wire _1181_;
 wire _1182_;
 wire _1183_;
 wire _1184_;
 wire _1185_;
 wire _1186_;
 wire _1187_;
 wire _1188_;
 wire _1189_;
 wire _1190_;
 wire _1191_;
 wire _1192_;
 wire _1193_;
 wire _1194_;
 wire _1195_;
 wire _1196_;
 wire _1197_;
 wire _1198_;
 wire _1199_;
 wire _1200_;
 wire _1201_;
 wire _1202_;
 wire _1203_;
 wire _1204_;
 wire _1205_;
 wire _1206_;
 wire _1207_;
 wire _1208_;
 wire _1209_;
 wire _1210_;
 wire _1211_;
 wire _1212_;
 wire _1213_;
 wire _1214_;
 wire _1215_;
 wire _1216_;
 wire _1217_;
 wire _1218_;
 wire _1219_;
 wire _1220_;
 wire _1221_;
 wire _1222_;
 wire _1223_;
 wire _1224_;
 wire _1225_;
 wire _1226_;
 wire _1227_;
 wire _1228_;
 wire _1229_;
 wire _1230_;
 wire _1231_;
 wire _1232_;
 wire _1233_;
 wire _1234_;
 wire _1235_;
 wire _1236_;
 wire _1237_;
 wire _1238_;
 wire _1239_;
 wire _1240_;
 wire _1241_;
 wire _1242_;
 wire _1243_;
 wire _1244_;
 wire _1245_;
 wire _1246_;
 wire _1247_;
 wire _1248_;
 wire _1249_;
 wire _1250_;
 wire _1251_;
 wire _1252_;
 wire _1253_;
 wire _1254_;
 wire _1255_;
 wire _1256_;
 wire _1257_;
 wire _1258_;
 wire _1259_;
 wire _1260_;
 wire _1261_;
 wire _1262_;
 wire _1263_;
 wire _1264_;
 wire _1265_;
 wire _1266_;
 wire _1267_;
 wire _1268_;
 wire _1269_;
 wire _1270_;
 wire _1271_;
 wire _1272_;
 wire _1273_;
 wire _1274_;
 wire _1275_;
 wire _1276_;
 wire _1277_;
 wire _1278_;
 wire _1279_;
 wire _1280_;
 wire _1281_;
 wire _1282_;
 wire _1283_;
 wire _1284_;
 wire _1285_;
 wire _1286_;
 wire _1287_;
 wire _1288_;
 wire _1289_;
 wire _1290_;
 wire _1291_;
 wire _1292_;
 wire _1293_;
 wire _1294_;
 wire _1295_;
 wire _1296_;
 wire _1297_;
 wire _1298_;
 wire _1299_;
 wire _1300_;
 wire _1301_;
 wire _1302_;
 wire _1303_;
 wire _1304_;
 wire _1305_;
 wire _1306_;
 wire _1307_;
 wire _1308_;
 wire _1309_;
 wire _1310_;
 wire _1311_;
 wire _1312_;
 wire _1313_;
 wire _1314_;
 wire _1315_;
 wire _1316_;
 wire _1317_;
 wire _1318_;
 wire _1319_;
 wire _1320_;
 wire _1321_;
 wire _1322_;
 wire _1323_;
 wire _1324_;
 wire _1325_;
 wire _1326_;
 wire _1327_;
 wire _1328_;
 wire _1329_;
 wire _1330_;
 wire _1331_;
 wire _1332_;
 wire _1333_;
 wire _1334_;
 wire _1335_;
 wire _1336_;
 wire _1337_;
 wire _1338_;
 wire _1339_;
 wire _1340_;
 wire _1341_;
 wire _1342_;
 wire _1343_;
 wire _1344_;
 wire _1345_;
 wire _1346_;
 wire _1347_;
 wire _1348_;
 wire _1349_;
 wire _1350_;
 wire _1351_;
 wire _1352_;
 wire _1353_;
 wire _1354_;
 wire _1355_;
 wire _1356_;
 wire _1357_;
 wire _1358_;
 wire _1359_;
 wire _1360_;
 wire _1361_;
 wire _1362_;
 wire _1363_;
 wire _1364_;
 wire _1365_;
 wire _1366_;
 wire _1367_;
 wire _1368_;
 wire _1369_;
 wire _1370_;
 wire _1371_;
 wire _1372_;
 wire _1373_;
 wire _1374_;
 wire _1375_;
 wire _1376_;
 wire _1377_;
 wire _1378_;
 wire _1379_;
 wire _1380_;
 wire _1381_;
 wire _1382_;
 wire _1383_;
 wire _1384_;
 wire _1385_;
 wire _1386_;
 wire _1387_;
 wire _1388_;
 wire _1389_;
 wire _1390_;
 wire _1391_;
 wire _1392_;
 wire _1393_;
 wire _1394_;
 wire _1395_;
 wire _1396_;
 wire _1397_;
 wire _1398_;
 wire _1399_;
 wire _1400_;
 wire _1401_;
 wire _1402_;
 wire _1403_;
 wire _1404_;
 wire _1405_;
 wire _1406_;
 wire _1407_;
 wire _1408_;
 wire _1409_;
 wire _1410_;
 wire _1411_;
 wire _1412_;
 wire _1413_;
 wire _1414_;
 wire _1415_;
 wire _1416_;
 wire _1417_;
 wire _1418_;
 wire _1419_;
 wire _1420_;
 wire _1421_;
 wire _1422_;
 wire _1423_;
 wire _1424_;
 wire _1425_;
 wire _1426_;
 wire _1427_;
 wire _1428_;
 wire _1429_;
 wire _1430_;
 wire _1431_;
 wire _1432_;
 wire _1433_;
 wire _1434_;
 wire _1435_;
 wire _1436_;
 wire _1437_;
 wire _1438_;
 wire _1439_;
 wire _1440_;
 wire _1441_;
 wire _1442_;
 wire _1443_;
 wire _1444_;
 wire _1445_;
 wire _1446_;
 wire _1447_;
 wire _1448_;
 wire _1449_;
 wire _1450_;
 wire _1451_;
 wire _1452_;
 wire _1453_;
 wire _1454_;
 wire _1455_;
 wire _1456_;
 wire _1457_;
 wire _1458_;
 wire _1459_;
 wire _1460_;
 wire _1461_;
 wire _1462_;
 wire _1463_;
 wire _1464_;
 wire _1465_;
 wire _1466_;
 wire _1467_;
 wire _1468_;
 wire _1469_;
 wire _1470_;
 wire _1471_;
 wire _1472_;
 wire _1473_;
 wire _1474_;
 wire _1475_;
 wire _1476_;
 wire _1477_;
 wire _1478_;
 wire _1479_;
 wire _1480_;
 wire _1481_;
 wire _1482_;
 wire _1483_;
 wire _1484_;
 wire _1485_;
 wire _1486_;
 wire _1487_;
 wire _1488_;
 wire _1489_;
 wire _1490_;
 wire _1491_;
 wire _1492_;
 wire _1493_;
 wire _1494_;
 wire _1495_;
 wire _1496_;
 wire _1497_;
 wire _1498_;
 wire _1499_;
 wire _1500_;
 wire _1501_;
 wire _1502_;
 wire _1503_;
 wire _1504_;
 wire _1505_;
 wire _1506_;
 wire _1507_;
 wire _1508_;
 wire _1509_;
 wire _1510_;
 wire _1511_;
 wire _1512_;
 wire _1513_;
 wire _1514_;
 wire _1515_;
 wire _1516_;
 wire _1517_;
 wire _1518_;
 wire _1519_;
 wire _1520_;
 wire _1521_;
 wire _1522_;
 wire _1523_;
 wire _1524_;
 wire _1525_;
 wire _1526_;
 wire _1527_;
 wire _1528_;
 wire _1529_;
 wire _1530_;
 wire _1531_;
 wire _1532_;
 wire _1533_;
 wire _1534_;
 wire _1535_;
 wire _1536_;
 wire _1537_;
 wire _1538_;
 wire _1539_;
 wire _1540_;
 wire _1541_;
 wire _1542_;
 wire _1543_;
 wire _1544_;
 wire _1545_;
 wire _1546_;
 wire _1547_;
 wire _1548_;
 wire _1549_;
 wire _1550_;
 wire _1551_;
 wire _1552_;
 wire _1553_;
 wire _1554_;
 wire _1555_;
 wire _1556_;
 wire _1557_;
 wire _1558_;
 wire _1559_;
 wire _1560_;
 wire _1561_;
 wire _1562_;
 wire _1563_;
 wire _1564_;
 wire _1565_;
 wire _1566_;
 wire _1567_;
 wire _1568_;
 wire _1569_;
 wire _1570_;
 wire _1571_;
 wire _1572_;
 wire _1573_;
 wire _1574_;
 wire _1575_;
 wire _1576_;
 wire _1577_;
 wire _1578_;
 wire _1579_;
 wire _1580_;
 wire _1581_;
 wire _1582_;
 wire _1583_;
 wire _1584_;
 wire _1585_;
 wire _1586_;
 wire _1587_;
 wire _1588_;
 wire _1589_;
 wire _1590_;
 wire _1591_;
 wire _1592_;
 wire _1593_;
 wire _1594_;
 wire _1595_;
 wire _1596_;
 wire _1597_;
 wire _1598_;
 wire _1599_;
 wire _1600_;
 wire _1601_;
 wire _1602_;
 wire _1603_;
 wire _1604_;
 wire _1605_;
 wire _1606_;
 wire _1607_;
 wire _1608_;
 wire _1609_;
 wire _1610_;
 wire _1611_;
 wire _1612_;
 wire _1613_;
 wire _1614_;
 wire _1615_;
 wire _1616_;
 wire _1617_;
 wire _1618_;
 wire _1619_;
 wire _1620_;
 wire _1621_;
 wire _1622_;
 wire _1623_;
 wire _1624_;
 wire _1625_;
 wire _1626_;
 wire _1627_;
 wire _1628_;
 wire _1629_;
 wire _1630_;
 wire _1631_;
 wire _1632_;
 wire _1633_;
 wire _1634_;
 wire _1635_;
 wire _1636_;
 wire _1637_;
 wire _1638_;
 wire _1639_;
 wire _1640_;
 wire _1641_;
 wire _1642_;
 wire _1643_;
 wire _1644_;
 wire _1645_;
 wire _1646_;
 wire _1647_;
 wire _1648_;
 wire _1649_;
 wire _1650_;
 wire _1651_;
 wire _1652_;
 wire _1653_;
 wire _1654_;
 wire _1655_;
 wire _1656_;
 wire _1657_;
 wire _1658_;
 wire _1659_;
 wire _1660_;
 wire _1661_;
 wire _1662_;
 wire _1663_;
 wire _1664_;
 wire _1665_;
 wire _1666_;
 wire _1667_;
 wire _1668_;
 wire _1669_;
 wire _1670_;
 wire _1671_;
 wire _1672_;
 wire _1673_;
 wire _1674_;
 wire _1675_;
 wire _1676_;
 wire _1677_;
 wire _1678_;
 wire _1679_;
 wire _1680_;
 wire _1681_;
 wire _1682_;
 wire _1683_;
 wire _1684_;
 wire _1685_;
 wire _1686_;
 wire _1687_;
 wire _1688_;
 wire _1689_;
 wire _1690_;
 wire _1691_;
 wire _1692_;
 wire _1693_;
 wire _1694_;
 wire _1695_;
 wire _1696_;
 wire _1697_;
 wire _1698_;
 wire _1699_;
 wire _1700_;
 wire _1701_;
 wire _1702_;
 wire _1703_;
 wire _1704_;
 wire _1705_;
 wire _1706_;
 wire _1707_;
 wire _1708_;
 wire _1709_;
 wire _1710_;
 wire _1711_;
 wire _1712_;
 wire _1713_;
 wire _1714_;
 wire _1715_;
 wire _1716_;
 wire _1717_;
 wire _1718_;
 wire _1719_;
 wire _1720_;
 wire _1721_;
 wire _1722_;
 wire _1723_;
 wire _1724_;
 wire _1725_;
 wire _1726_;
 wire _1727_;
 wire _1728_;
 wire _1729_;
 wire _1730_;
 wire _1731_;
 wire _1732_;
 wire _1733_;
 wire _1734_;
 wire _1735_;
 wire _1736_;
 wire _1737_;
 wire _1738_;
 wire _1739_;
 wire _1740_;
 wire _1741_;
 wire _1742_;
 wire _1743_;
 wire _1744_;
 wire _1745_;
 wire _1746_;
 wire _1747_;
 wire _1748_;
 wire _1749_;
 wire _1750_;
 wire _1751_;
 wire _1752_;
 wire _1753_;
 wire _1754_;
 wire _1755_;
 wire _1756_;
 wire _1757_;
 wire _1758_;
 wire _1759_;
 wire _1760_;
 wire _1761_;
 wire _1762_;
 wire _1763_;
 wire _1764_;
 wire _1765_;
 wire _1766_;
 wire _1767_;
 wire _1768_;
 wire _1769_;
 wire _1770_;
 wire _1771_;
 wire _1772_;
 wire _1773_;
 wire _1774_;
 wire _1775_;
 wire _1776_;
 wire _1777_;
 wire _1778_;
 wire _1779_;
 wire _1780_;
 wire _1781_;
 wire _1782_;
 wire _1783_;
 wire _1784_;
 wire _1785_;
 wire _1786_;
 wire _1787_;
 wire _1788_;
 wire _1789_;
 wire _1790_;
 wire _1791_;
 wire _1792_;
 wire _1793_;
 wire _1794_;
 wire _1795_;
 wire _1796_;
 wire _1797_;
 wire _1798_;
 wire _1799_;
 wire _1800_;
 wire _1801_;
 wire _1802_;
 wire _1803_;
 wire _1804_;
 wire _1805_;
 wire _1806_;
 wire _1807_;
 wire _1808_;
 wire _1809_;
 wire _1810_;
 wire _1811_;
 wire _1812_;
 wire _1813_;
 wire _1814_;
 wire _1815_;
 wire _1816_;
 wire _1817_;
 wire _1818_;
 wire _1819_;
 wire _1820_;
 wire _1821_;
 wire _1822_;
 wire _1823_;
 wire _1824_;
 wire _1825_;
 wire _1826_;
 wire _1827_;
 wire _1828_;
 wire _1829_;
 wire _1830_;
 wire _1831_;
 wire _1832_;
 wire _1833_;
 wire _1834_;
 wire _1835_;
 wire _1836_;
 wire _1837_;
 wire _1838_;
 wire _1839_;
 wire _1840_;
 wire _1841_;
 wire _1842_;
 wire _1843_;
 wire _1844_;
 wire _1845_;
 wire _1846_;
 wire _1847_;
 wire _1848_;
 wire _1849_;
 wire _1850_;
 wire _1851_;
 wire _1852_;
 wire _1853_;
 wire _1854_;
 wire _1855_;
 wire _1856_;
 wire _1857_;
 wire _1858_;
 wire _1859_;
 wire _1860_;
 wire _1861_;
 wire _1862_;
 wire _1863_;
 wire _1864_;
 wire _1865_;
 wire _1866_;
 wire _1867_;
 wire _1868_;
 wire _1869_;
 wire _1870_;
 wire _1871_;
 wire _1872_;
 wire _1873_;
 wire _1874_;
 wire _1875_;
 wire _1876_;
 wire _1877_;
 wire _1878_;
 wire _1879_;
 wire _1880_;
 wire _1881_;
 wire _1882_;
 wire _1883_;
 wire _1884_;
 wire _1885_;
 wire _1886_;
 wire _1887_;
 wire _1888_;
 wire _1889_;
 wire _1890_;
 wire _1891_;
 wire _1892_;
 wire _1893_;
 wire _1894_;
 wire _1895_;
 wire _1896_;
 wire _1897_;
 wire _1898_;
 wire _1899_;
 wire _1900_;
 wire _1901_;
 wire _1902_;
 wire _1903_;
 wire _1904_;
 wire _1905_;
 wire _1906_;
 wire _1907_;
 wire _1908_;
 wire _1909_;
 wire _1910_;
 wire _1911_;
 wire _1912_;
 wire _1913_;
 wire _1914_;
 wire _1915_;
 wire _1916_;
 wire _1917_;
 wire _1918_;
 wire _1919_;
 wire _1920_;
 wire _1921_;
 wire _1922_;
 wire _1923_;
 wire _1924_;
 wire _1925_;
 wire _1926_;
 wire _1927_;
 wire _1928_;
 wire _1929_;
 wire _1930_;
 wire _1931_;
 wire _1932_;
 wire _1933_;
 wire _1934_;
 wire _1935_;
 wire _1936_;
 wire _1937_;
 wire _1938_;
 wire _1939_;
 wire _1940_;
 wire _1941_;
 wire _1942_;
 wire _1943_;
 wire _1944_;
 wire _1945_;
 wire _1946_;
 wire _1947_;
 wire _1948_;
 wire _1949_;
 wire _1950_;
 wire _1951_;
 wire _1952_;
 wire _1953_;
 wire _1954_;
 wire _1955_;
 wire _1956_;
 wire _1957_;
 wire _1958_;
 wire _1959_;
 wire _1960_;
 wire _1961_;
 wire _1962_;
 wire _1963_;
 wire _1964_;
 wire _1965_;
 wire _1966_;
 wire _1967_;
 wire _1968_;
 wire _1969_;
 wire _1970_;
 wire _1971_;
 wire _1972_;
 wire _1973_;
 wire _1974_;
 wire _1975_;
 wire _1976_;
 wire _1977_;
 wire _1978_;
 wire _1979_;
 wire _1980_;
 wire _1981_;
 wire _1982_;
 wire _1983_;
 wire _1984_;
 wire _1985_;
 wire _1986_;
 wire _1987_;
 wire _1988_;
 wire _1989_;
 wire _1990_;
 wire _1991_;
 wire _1992_;
 wire _1993_;
 wire _1994_;
 wire _1995_;
 wire _1996_;
 wire _1997_;
 wire _1998_;
 wire _1999_;
 wire _2000_;
 wire _2001_;
 wire _2002_;
 wire _2003_;
 wire _2004_;
 wire _2005_;
 wire _2006_;
 wire _2007_;
 wire _2008_;
 wire _2009_;
 wire _2010_;
 wire _2011_;
 wire _2012_;
 wire _2013_;
 wire _2014_;
 wire _2015_;
 wire _2016_;
 wire _2017_;
 wire _2018_;
 wire _2019_;
 wire _2020_;
 wire _2021_;
 wire _2022_;
 wire _2023_;
 wire _2024_;
 wire _2025_;
 wire _2026_;
 wire _2027_;
 wire _2028_;
 wire _2029_;
 wire _2030_;
 wire _2031_;
 wire _2032_;
 wire _2033_;
 wire _2034_;
 wire _2035_;
 wire _2036_;
 wire _2037_;
 wire _2038_;
 wire _2039_;
 wire _2040_;
 wire _2041_;
 wire _2042_;
 wire _2043_;
 wire _2044_;
 wire _2045_;
 wire _2046_;
 wire _2047_;
 wire _2048_;
 wire _2049_;
 wire _2050_;
 wire _2051_;
 wire _2052_;
 wire _2053_;
 wire _2054_;
 wire _2055_;
 wire _2056_;
 wire _2057_;
 wire _2058_;
 wire _2059_;
 wire _2060_;
 wire _2061_;
 wire _2062_;
 wire _2063_;
 wire _2064_;
 wire _2065_;
 wire _2066_;
 wire _2067_;
 wire _2068_;
 wire _2069_;
 wire _2070_;
 wire _2071_;
 wire _2072_;
 wire _2073_;
 wire _2074_;
 wire _2075_;
 wire _2076_;
 wire _2077_;
 wire _2078_;
 wire _2079_;
 wire _2080_;
 wire _2081_;
 wire _2082_;
 wire _2083_;
 wire _2084_;
 wire _2085_;
 wire _2086_;
 wire _2087_;
 wire _2088_;
 wire _2089_;
 wire _2090_;
 wire _2091_;
 wire _2092_;
 wire _2093_;
 wire _2094_;
 wire _2095_;
 wire _2096_;
 wire _2097_;
 wire _2098_;
 wire _2099_;
 wire _2100_;
 wire _2101_;
 wire _2102_;
 wire _2103_;
 wire _2104_;
 wire _2105_;
 wire _2106_;
 wire _2107_;
 wire _2108_;
 wire _2109_;
 wire _2110_;
 wire _2111_;
 wire _2112_;
 wire _2113_;
 wire _2114_;
 wire _2115_;
 wire _2116_;
 wire _2117_;
 wire _2118_;
 wire _2119_;
 wire _2120_;
 wire _2121_;
 wire _2122_;
 wire _2123_;
 wire _2124_;
 wire _2125_;
 wire _2126_;
 wire _2127_;
 wire _2128_;
 wire _2129_;
 wire _2130_;
 wire _2131_;
 wire _2132_;
 wire _2133_;
 wire _2134_;
 wire _2135_;
 wire _2136_;
 wire _2137_;
 wire _2138_;
 wire _2139_;
 wire _2140_;
 wire _2141_;
 wire _2142_;
 wire _2143_;
 wire _2144_;
 wire _2145_;
 wire _2146_;
 wire _2147_;
 wire _2148_;
 wire _2149_;
 wire _2150_;
 wire _2151_;
 wire _2152_;
 wire _2153_;
 wire _2154_;
 wire _2155_;
 wire _2156_;
 wire _2157_;
 wire _2158_;
 wire _2159_;
 wire _2160_;
 wire _2161_;
 wire _2162_;
 wire _2163_;
 wire _2164_;
 wire _2165_;
 wire _2166_;
 wire _2167_;
 wire _2168_;
 wire _2169_;
 wire _2170_;
 wire _2171_;
 wire _2172_;
 wire _2173_;
 wire _2174_;
 wire _2175_;
 wire _2176_;
 wire _2177_;
 wire _2178_;
 wire _2179_;
 wire _2180_;
 wire _2181_;
 wire _2182_;
 wire _2183_;
 wire _2184_;
 wire _2185_;
 wire _2186_;
 wire _2187_;
 wire _2188_;
 wire _2189_;
 wire _2190_;
 wire _2191_;
 wire _2192_;
 wire _2193_;
 wire _2194_;
 wire _2195_;
 wire _2196_;
 wire _2197_;
 wire _2198_;
 wire _2199_;
 wire _2200_;
 wire _2201_;
 wire _2202_;
 wire _2203_;
 wire _2204_;
 wire _2205_;
 wire _2206_;
 wire _2207_;
 wire _2208_;
 wire _2209_;
 wire _2210_;
 wire _2211_;
 wire _2212_;
 wire _2213_;
 wire _2214_;
 wire _2215_;
 wire _2216_;
 wire _2217_;
 wire _2218_;
 wire _2219_;
 wire _2220_;
 wire _2221_;
 wire _2222_;
 wire _2223_;
 wire _2224_;
 wire _2225_;
 wire _2226_;
 wire _2227_;
 wire _2228_;
 wire _2229_;
 wire _2230_;
 wire _2231_;
 wire _2232_;
 wire _2233_;
 wire _2234_;
 wire _2235_;
 wire _2236_;
 wire _2237_;
 wire _2238_;
 wire _2239_;
 wire _2240_;
 wire _2241_;
 wire _2242_;
 wire _2243_;
 wire _2244_;
 wire _2245_;
 wire _2246_;
 wire _2247_;
 wire _2248_;
 wire _2249_;
 wire _2250_;
 wire _2251_;
 wire _2252_;
 wire _2253_;
 wire _2254_;
 wire _2255_;
 wire _2256_;
 wire _2257_;
 wire _2258_;
 wire _2259_;
 wire _2260_;
 wire _2261_;
 wire _2262_;
 wire _2263_;
 wire _2264_;
 wire _2265_;
 wire _2266_;
 wire _2267_;
 wire _2268_;
 wire _2269_;
 wire _2270_;
 wire _2271_;
 wire _2272_;
 wire _2273_;
 wire _2274_;
 wire _2275_;
 wire _2276_;
 wire _2277_;
 wire _2278_;
 wire _2279_;
 wire _2280_;
 wire _2281_;
 wire _2282_;
 wire _2283_;
 wire _2284_;
 wire _2285_;
 wire _2286_;
 wire _2287_;
 wire _2288_;
 wire _2289_;
 wire _2290_;
 wire _2291_;
 wire _2292_;
 wire _2293_;
 wire _2294_;
 wire _2295_;
 wire _2296_;
 wire _2297_;
 wire _2298_;
 wire _2299_;
 wire _2300_;
 wire _2301_;
 wire _2302_;
 wire _2303_;
 wire _2304_;
 wire _2305_;
 wire _2306_;
 wire _2307_;
 wire _2308_;
 wire _2309_;
 wire _2310_;
 wire _2311_;
 wire _2312_;
 wire _2313_;
 wire _2314_;
 wire _2315_;
 wire _2316_;
 wire _2317_;
 wire _2318_;
 wire _2319_;
 wire _2320_;
 wire _2321_;
 wire _2322_;
 wire _2323_;
 wire _2324_;
 wire _2325_;
 wire _2326_;
 wire _2327_;
 wire _2328_;
 wire _2329_;
 wire _2330_;
 wire _2331_;
 wire _2332_;
 wire _2333_;
 wire _2334_;
 wire _2335_;
 wire _2336_;
 wire _2337_;
 wire _2338_;
 wire _2339_;
 wire _2340_;
 wire _2341_;
 wire _2342_;
 wire _2343_;
 wire _2344_;
 wire _2345_;
 wire _2346_;
 wire _2347_;
 wire _2348_;
 wire _2349_;
 wire _2350_;
 wire _2351_;
 wire _2352_;
 wire _2353_;
 wire _2354_;
 wire _2355_;
 wire _2356_;
 wire _2357_;
 wire _2358_;
 wire _2359_;
 wire _2360_;
 wire _2361_;
 wire _2362_;
 wire _2363_;
 wire _2364_;
 wire _2365_;
 wire _2366_;
 wire _2367_;
 wire _2368_;
 wire _2369_;
 wire _2370_;
 wire _2371_;
 wire _2372_;
 wire _2373_;
 wire _2374_;
 wire _2375_;
 wire _2376_;
 wire _2377_;
 wire _2378_;
 wire _2379_;
 wire _2380_;
 wire _2381_;
 wire _2382_;
 wire _2383_;
 wire _2384_;
 wire _2385_;
 wire _2386_;
 wire _2387_;
 wire _2388_;
 wire _2389_;
 wire _2390_;
 wire _2391_;
 wire _2392_;
 wire _2393_;
 wire _2394_;
 wire _2395_;
 wire _2396_;
 wire _2397_;
 wire _2398_;
 wire _2399_;
 wire _2400_;
 wire _2401_;
 wire _2402_;
 wire _2403_;
 wire _2404_;
 wire _2405_;
 wire _2406_;
 wire _2407_;
 wire _2408_;
 wire _2409_;
 wire _2410_;
 wire _2411_;
 wire _2412_;
 wire _2413_;
 wire _2414_;
 wire _2415_;
 wire _2416_;
 wire _2417_;
 wire _2418_;
 wire _2419_;
 wire _2420_;
 wire _2421_;
 wire _2422_;
 wire _2423_;
 wire _2424_;
 wire _2425_;
 wire _2426_;
 wire _2427_;
 wire _2428_;
 wire _2429_;
 wire _2430_;
 wire _2431_;
 wire _2432_;
 wire _2433_;
 wire _2434_;
 wire _2435_;
 wire _2436_;
 wire _2437_;
 wire _2438_;
 wire _2439_;
 wire _2440_;
 wire _2441_;
 wire _2442_;
 wire _2443_;
 wire _2444_;
 wire _2445_;
 wire _2446_;
 wire _2447_;
 wire _2448_;
 wire _2449_;
 wire _2450_;
 wire _2451_;
 wire _2452_;
 wire _2453_;
 wire _2454_;
 wire _2455_;
 wire _2456_;
 wire _2457_;
 wire _2458_;
 wire _2459_;
 wire _2460_;
 wire _2461_;
 wire _2462_;
 wire _2463_;
 wire _2464_;
 wire _2465_;
 wire _2466_;
 wire _2467_;
 wire _2468_;
 wire _2469_;
 wire _2470_;
 wire _2471_;
 wire _2472_;
 wire _2473_;
 wire _2474_;
 wire _2475_;
 wire _2476_;
 wire _2477_;
 wire _2478_;
 wire _2479_;
 wire _2480_;
 wire _2481_;
 wire _2482_;
 wire _2483_;
 wire _2484_;
 wire _2485_;
 wire _2486_;
 wire _2487_;
 wire _2488_;
 wire _2489_;
 wire _2490_;
 wire _2491_;
 wire _2492_;
 wire _2493_;
 wire _2494_;
 wire _2495_;
 wire _2496_;
 wire _2497_;
 wire _2498_;
 wire _2499_;
 wire _2500_;
 wire _2501_;
 wire _2502_;
 wire _2503_;
 wire _2504_;
 wire _2505_;
 wire _2506_;
 wire _2507_;
 wire _2508_;
 wire _2509_;
 wire _2510_;
 wire _2511_;
 wire _2512_;
 wire _2513_;
 wire _2514_;
 wire _2515_;
 wire _2516_;
 wire _2517_;
 wire _2518_;
 wire _2519_;
 wire _2520_;
 wire _2521_;
 wire _2522_;
 wire _2523_;
 wire _2524_;
 wire _2525_;
 wire _2526_;
 wire _2527_;
 wire _2528_;
 wire _2529_;
 wire _2530_;
 wire _2531_;
 wire _2532_;
 wire _2533_;
 wire _2534_;
 wire _2535_;
 wire _2536_;
 wire _2537_;
 wire _2538_;
 wire _2539_;
 wire _2540_;
 wire _2541_;
 wire _2542_;
 wire _2543_;
 wire _2544_;
 wire _2545_;
 wire _2546_;
 wire _2547_;
 wire _2548_;
 wire _2549_;
 wire _2550_;
 wire _2551_;
 wire _2552_;
 wire _2553_;
 wire _2554_;
 wire _2555_;
 wire _2556_;
 wire _2557_;
 wire _2558_;
 wire _2559_;
 wire _2560_;
 wire _2561_;
 wire _2562_;
 wire _2563_;
 wire _2564_;
 wire _2565_;
 wire _2566_;
 wire _2567_;
 wire _2568_;
 wire _2569_;
 wire _2570_;
 wire _2571_;
 wire _2572_;
 wire _2573_;
 wire _2574_;
 wire _2575_;
 wire _2576_;
 wire _2577_;
 wire _2578_;
 wire _2579_;
 wire _2580_;
 wire _2581_;
 wire _2582_;
 wire _2583_;
 wire _2584_;
 wire _2585_;
 wire _2586_;
 wire _2587_;
 wire _2588_;
 wire _2589_;
 wire _2590_;
 wire _2591_;
 wire _2592_;
 wire _2593_;
 wire _2594_;
 wire _2595_;
 wire _2596_;
 wire _2597_;
 wire _2598_;
 wire _2599_;
 wire _2600_;
 wire _2601_;
 wire _2602_;
 wire _2603_;
 wire _2604_;
 wire _2605_;
 wire _2606_;
 wire _2607_;
 wire _2608_;
 wire _2609_;
 wire _2610_;
 wire _2611_;
 wire _2612_;
 wire _2613_;
 wire _2614_;
 wire _2615_;
 wire _2616_;
 wire _2617_;
 wire _2618_;
 wire _2619_;
 wire _2620_;
 wire _2621_;
 wire _2622_;
 wire _2623_;
 wire _2624_;
 wire _2625_;
 wire _2626_;
 wire _2627_;
 wire _2628_;
 wire _2629_;
 wire _2630_;
 wire _2631_;
 wire _2632_;
 wire _2633_;
 wire _2634_;
 wire _2635_;
 wire _2636_;
 wire _2637_;
 wire _2638_;
 wire _2639_;
 wire _2640_;
 wire _2641_;
 wire _2642_;
 wire _2643_;
 wire _2644_;
 wire _2645_;
 wire _2646_;
 wire _2647_;
 wire _2648_;
 wire _2649_;
 wire _2650_;
 wire _2651_;
 wire _2652_;
 wire _2653_;
 wire _2654_;
 wire _2655_;
 wire _2656_;
 wire _2657_;
 wire _2658_;
 wire _2659_;
 wire _2660_;
 wire _2661_;
 wire _2662_;
 wire _2663_;
 wire _2664_;
 wire _2665_;
 wire _2666_;
 wire _2667_;
 wire _2668_;
 wire _2669_;
 wire _2670_;
 wire _2671_;
 wire _2672_;
 wire _2673_;
 wire _2674_;
 wire _2675_;
 wire _2676_;
 wire _2677_;
 wire _2678_;
 wire _2679_;
 wire _2680_;
 wire _2681_;
 wire _2682_;
 wire _2683_;
 wire _2684_;
 wire _2685_;
 wire _2686_;
 wire _2687_;
 wire _2688_;
 wire _2689_;
 wire _2690_;
 wire _2691_;
 wire _2692_;
 wire _2693_;
 wire _2694_;
 wire _2695_;
 wire _2696_;
 wire _2697_;
 wire _2698_;
 wire _2699_;
 wire _2700_;
 wire _2701_;
 wire _2702_;
 wire _2703_;
 wire _2704_;
 wire _2705_;
 wire _2706_;
 wire _2707_;
 wire _2708_;
 wire _2709_;
 wire _2710_;
 wire _2711_;
 wire _2712_;
 wire _2713_;
 wire _2714_;
 wire _2715_;
 wire _2716_;
 wire _2717_;
 wire _2718_;
 wire _2719_;
 wire _2720_;
 wire _2721_;
 wire _2722_;
 wire _2723_;
 wire _2724_;
 wire _2725_;
 wire _2726_;
 wire _2727_;
 wire _2728_;
 wire _2729_;
 wire _2730_;
 wire _2731_;
 wire _2732_;
 wire _2733_;
 wire _2734_;
 wire _2735_;
 wire _2736_;
 wire _2737_;
 wire _2738_;
 wire _2739_;
 wire _2740_;
 wire _2741_;
 wire _2742_;
 wire _2743_;
 wire _2744_;
 wire _2745_;
 wire _2746_;
 wire _2747_;
 wire _2748_;
 wire _2749_;
 wire _2750_;
 wire _2751_;
 wire _2752_;
 wire _2753_;
 wire _2754_;
 wire _2755_;
 wire _2756_;
 wire _2757_;
 wire _2758_;
 wire _2759_;
 wire _2760_;
 wire _2761_;
 wire _2762_;
 wire _2763_;
 wire _2764_;
 wire _2765_;
 wire _2766_;
 wire _2767_;
 wire _2768_;
 wire _2769_;
 wire _2770_;
 wire _2771_;
 wire _2772_;
 wire _2773_;
 wire _2774_;
 wire _2775_;
 wire _2776_;
 wire _2777_;
 wire _2778_;
 wire _2779_;
 wire _2780_;
 wire _2781_;
 wire _2782_;
 wire _2783_;
 wire _2784_;
 wire _2785_;
 wire _2786_;
 wire _2787_;
 wire _2788_;
 wire _2789_;
 wire _2790_;
 wire _2791_;
 wire _2792_;
 wire _2793_;
 wire _2794_;
 wire _2795_;
 wire _2796_;
 wire _2797_;
 wire _2798_;
 wire _2799_;
 wire _2800_;
 wire _2801_;
 wire _2802_;
 wire _2803_;
 wire _2804_;
 wire _2805_;
 wire _2806_;
 wire _2807_;
 wire _2808_;
 wire _2809_;
 wire _2810_;
 wire _2811_;
 wire _2812_;
 wire _2813_;
 wire _2814_;
 wire _2815_;
 wire _2816_;
 wire _2817_;
 wire _2818_;
 wire _2819_;
 wire _2820_;
 wire _2821_;
 wire _2822_;
 wire _2823_;
 wire _2824_;
 wire _2825_;
 wire _2826_;
 wire _2827_;
 wire _2828_;
 wire _2829_;
 wire _2830_;
 wire _2831_;
 wire _2832_;
 wire _2833_;
 wire _2834_;
 wire _2835_;
 wire _2836_;
 wire _2837_;
 wire _2838_;
 wire _2839_;
 wire _2840_;
 wire _2841_;
 wire _2842_;
 wire _2843_;
 wire _2844_;
 wire _2845_;
 wire _2846_;
 wire _2847_;
 wire _2848_;
 wire _2849_;
 wire _2850_;
 wire _2851_;
 wire _2852_;
 wire _2853_;
 wire _2854_;
 wire _2855_;
 wire _2856_;
 wire _2857_;
 wire _2858_;
 wire _2859_;
 wire _2860_;
 wire _2861_;
 wire _2862_;
 wire _2863_;
 wire _2864_;
 wire _2865_;
 wire _2866_;
 wire _2867_;
 wire _2868_;
 wire _2869_;
 wire _2870_;
 wire _2871_;
 wire _2872_;
 wire _2873_;
 wire _2874_;
 wire _2875_;
 wire _2876_;
 wire _2877_;
 wire _2878_;
 wire _2879_;
 wire _2880_;
 wire _2881_;
 wire _2882_;
 wire _2883_;
 wire _2884_;
 wire _2885_;
 wire _2886_;
 wire _2887_;
 wire _2888_;
 wire _2889_;
 wire _2890_;
 wire _2891_;
 wire _2892_;
 wire _2893_;
 wire _2894_;
 wire _2895_;
 wire _2896_;
 wire _2897_;
 wire _2898_;
 wire _2899_;
 wire _2900_;
 wire _2901_;
 wire _2902_;
 wire _2903_;
 wire _2904_;
 wire _2905_;
 wire _2906_;
 wire _2907_;
 wire _2908_;
 wire _2909_;
 wire _2910_;
 wire _2911_;
 wire _2912_;
 wire _2913_;
 wire _2914_;
 wire _2915_;
 wire _2916_;
 wire _2917_;
 wire _2918_;
 wire _2919_;
 wire _2920_;
 wire _2921_;
 wire _2922_;
 wire _2923_;
 wire _2924_;
 wire _2925_;
 wire _2926_;
 wire _2927_;
 wire _2928_;
 wire _2929_;
 wire _2930_;
 wire _2931_;
 wire _2932_;
 wire _2933_;
 wire _2934_;
 wire _2935_;
 wire _2936_;
 wire _2937_;
 wire _2938_;
 wire _2939_;
 wire _2940_;
 wire _2941_;
 wire _2942_;
 wire _2943_;
 wire _2944_;
 wire _2945_;
 wire _2946_;
 wire _2947_;
 wire _2948_;
 wire _2949_;
 wire _2950_;
 wire _2951_;
 wire _2952_;
 wire _2953_;
 wire _2954_;
 wire _2955_;
 wire _2956_;
 wire _2957_;
 wire _2958_;
 wire _2959_;
 wire _2960_;
 wire _2961_;
 wire _2962_;
 wire _2963_;
 wire _2964_;
 wire _2965_;
 wire _2966_;
 wire _2967_;
 wire _2968_;
 wire _2969_;
 wire _2970_;
 wire _2971_;
 wire _2972_;
 wire _2973_;
 wire _2974_;
 wire _2975_;
 wire _2976_;
 wire _2977_;
 wire _2978_;
 wire _2979_;
 wire _2980_;
 wire _2981_;
 wire _2982_;
 wire _2983_;
 wire _2984_;
 wire _2985_;
 wire _2986_;
 wire _2987_;
 wire _2988_;
 wire _2989_;
 wire _2990_;
 wire _2991_;
 wire _2992_;
 wire _2993_;
 wire _2994_;
 wire _2995_;
 wire _2996_;
 wire _2997_;
 wire _2998_;
 wire _2999_;
 wire _3000_;
 wire _3001_;
 wire _3002_;
 wire _3003_;
 wire _3004_;
 wire _3005_;
 wire _3006_;
 wire _3007_;
 wire _3008_;
 wire _3009_;
 wire _3010_;
 wire _3011_;
 wire _3012_;
 wire _3013_;
 wire _3014_;
 wire _3015_;
 wire _3016_;
 wire _3017_;
 wire _3018_;
 wire _3019_;
 wire _3020_;
 wire _3021_;
 wire _3022_;
 wire _3023_;
 wire _3024_;
 wire _3025_;
 wire _3026_;
 wire _3027_;
 wire _3028_;
 wire _3029_;
 wire _3030_;
 wire _3031_;
 wire _3032_;
 wire _3033_;
 wire _3034_;
 wire _3035_;
 wire _3036_;
 wire _3037_;
 wire _3038_;
 wire _3039_;
 wire _3040_;
 wire _3041_;
 wire _3042_;
 wire _3043_;
 wire _3044_;
 wire _3045_;
 wire _3046_;
 wire _3047_;
 wire _3048_;
 wire _3049_;
 wire _3050_;
 wire _3051_;
 wire _3052_;
 wire _3053_;
 wire _3054_;
 wire _3055_;
 wire _3056_;
 wire _3057_;
 wire _3058_;
 wire _3059_;
 wire _3060_;
 wire _3061_;
 wire _3062_;
 wire _3063_;
 wire _3064_;
 wire _3065_;
 wire _3066_;
 wire _3067_;
 wire _3068_;
 wire _3069_;
 wire _3070_;
 wire _3071_;
 wire _3072_;
 wire _3073_;
 wire _3074_;
 wire _3075_;
 wire _3076_;
 wire _3077_;
 wire _3078_;
 wire _3079_;
 wire _3080_;
 wire _3081_;
 wire _3082_;
 wire _3083_;
 wire _3084_;
 wire _3085_;
 wire _3086_;
 wire _3087_;
 wire _3088_;
 wire _3089_;
 wire _3090_;
 wire _3091_;
 wire _3092_;
 wire _3093_;
 wire _3094_;
 wire _3095_;
 wire _3096_;
 wire _3097_;
 wire _3098_;
 wire _3099_;
 wire _3100_;
 wire _3101_;
 wire _3102_;
 wire _3103_;
 wire _3104_;
 wire _3105_;
 wire _3106_;
 wire _3107_;
 wire _3108_;
 wire _3109_;
 wire _3110_;
 wire _3111_;
 wire _3112_;
 wire _3113_;
 wire _3114_;
 wire _3115_;
 wire _3116_;
 wire _3117_;
 wire _3118_;
 wire _3119_;
 wire _3120_;
 wire _3121_;
 wire _3122_;
 wire _3123_;
 wire _3124_;
 wire _3125_;
 wire _3126_;
 wire _3127_;
 wire _3128_;
 wire _3129_;
 wire _3130_;
 wire _3131_;
 wire _3132_;
 wire _3133_;
 wire _3134_;
 wire _3135_;
 wire _3136_;
 wire _3137_;
 wire _3138_;
 wire _3139_;
 wire _3140_;
 wire _3141_;
 wire _3142_;
 wire _3143_;
 wire _3144_;
 wire _3145_;
 wire _3146_;
 wire _3147_;
 wire _3148_;
 wire _3149_;
 wire _3150_;
 wire _3151_;
 wire _3152_;
 wire _3153_;
 wire _3154_;
 wire _3155_;
 wire _3156_;
 wire _3157_;
 wire _3158_;
 wire _3159_;
 wire _3160_;
 wire _3161_;
 wire _3162_;
 wire _3163_;
 wire _3164_;
 wire _3165_;
 wire _3166_;
 wire _3167_;
 wire _3168_;
 wire _3169_;
 wire _3170_;
 wire _3171_;
 wire _3172_;
 wire _3173_;
 wire _3174_;
 wire _3175_;
 wire _3176_;
 wire _3177_;
 wire _3178_;
 wire _3179_;
 wire _3180_;
 wire _3181_;
 wire _3182_;
 wire _3183_;
 wire _3184_;
 wire _3185_;
 wire _3186_;
 wire _3187_;
 wire _3188_;
 wire _3189_;
 wire _3190_;
 wire _3191_;
 wire _3192_;
 wire _3193_;
 wire _3194_;
 wire _3195_;
 wire _3196_;
 wire _3197_;
 wire _3198_;
 wire _3199_;
 wire _3200_;
 wire _3201_;
 wire _3202_;
 wire _3203_;
 wire _3204_;
 wire _3205_;
 wire _3206_;
 wire _3207_;
 wire _3208_;
 wire _3209_;
 wire _3210_;
 wire _3211_;
 wire _3212_;
 wire _3213_;
 wire _3214_;
 wire _3215_;
 wire _3216_;
 wire _3217_;
 wire clknet_leaf_0_clk;
 wire net199;
 wire \g.g_y[0].g_x[0].t.out_sc ;
 wire \g.g_y[0].g_x[0].t.r_d ;
 wire \g.g_y[0].g_x[0].t.r_ghl ;
 wire \g.g_y[0].g_x[0].t.r_gnl ;
 wire \g.g_y[0].g_x[0].t.r_h ;
 wire \g.g_y[0].g_x[0].t.r_v ;
 wire \g.g_y[0].g_x[1].t.out_sc ;
 wire \g.g_y[0].g_x[1].t.r_d ;
 wire \g.g_y[0].g_x[1].t.r_h ;
 wire \g.g_y[0].g_x[1].t.r_v ;
 wire \g.g_y[0].g_x[2].t.out_sc ;
 wire \g.g_y[0].g_x[2].t.r_d ;
 wire \g.g_y[0].g_x[2].t.r_ghl ;
 wire \g.g_y[0].g_x[2].t.r_gnl ;
 wire \g.g_y[0].g_x[2].t.r_h ;
 wire \g.g_y[0].g_x[2].t.r_v ;
 wire \g.g_y[0].g_x[3].t.out_sc ;
 wire \g.g_y[0].g_x[3].t.r_d ;
 wire \g.g_y[0].g_x[3].t.r_h ;
 wire \g.g_y[0].g_x[3].t.r_v ;
 wire \g.g_y[0].g_x[4].t.out_sc ;
 wire \g.g_y[0].g_x[4].t.r_d ;
 wire \g.g_y[0].g_x[4].t.r_ghl ;
 wire \g.g_y[0].g_x[4].t.r_gnl ;
 wire \g.g_y[0].g_x[4].t.r_h ;
 wire \g.g_y[0].g_x[4].t.r_v ;
 wire \g.g_y[0].g_x[5].t.out_sc ;
 wire \g.g_y[0].g_x[5].t.r_d ;
 wire \g.g_y[0].g_x[5].t.r_h ;
 wire \g.g_y[0].g_x[5].t.r_v ;
 wire \g.g_y[0].g_x[6].t.out_sc ;
 wire \g.g_y[0].g_x[6].t.r_d ;
 wire \g.g_y[0].g_x[6].t.r_ghl ;
 wire \g.g_y[0].g_x[6].t.r_gnl ;
 wire \g.g_y[0].g_x[6].t.r_h ;
 wire \g.g_y[0].g_x[6].t.r_v ;
 wire \g.g_y[0].g_x[7].t.out_r ;
 wire \g.g_y[0].g_x[7].t.out_sc ;
 wire \g.g_y[0].g_x[7].t.r_d ;
 wire \g.g_y[0].g_x[7].t.r_h ;
 wire \g.g_y[0].g_x[7].t.r_v ;
 wire \g.g_y[1].g_x[0].t.out_sc ;
 wire \g.g_y[1].g_x[0].t.r_d ;
 wire \g.g_y[1].g_x[0].t.r_h ;
 wire \g.g_y[1].g_x[0].t.r_v ;
 wire \g.g_y[1].g_x[1].t.out_sc ;
 wire \g.g_y[1].g_x[1].t.r_d ;
 wire \g.g_y[1].g_x[1].t.r_ghl ;
 wire \g.g_y[1].g_x[1].t.r_gnl ;
 wire \g.g_y[1].g_x[1].t.r_h ;
 wire \g.g_y[1].g_x[1].t.r_v ;
 wire \g.g_y[1].g_x[2].t.out_sc ;
 wire \g.g_y[1].g_x[2].t.r_d ;
 wire \g.g_y[1].g_x[2].t.r_h ;
 wire \g.g_y[1].g_x[2].t.r_v ;
 wire \g.g_y[1].g_x[3].t.out_sc ;
 wire \g.g_y[1].g_x[3].t.r_d ;
 wire \g.g_y[1].g_x[3].t.r_ghl ;
 wire \g.g_y[1].g_x[3].t.r_gnl ;
 wire \g.g_y[1].g_x[3].t.r_h ;
 wire \g.g_y[1].g_x[3].t.r_v ;
 wire \g.g_y[1].g_x[4].t.out_sc ;
 wire \g.g_y[1].g_x[4].t.r_d ;
 wire \g.g_y[1].g_x[4].t.r_h ;
 wire \g.g_y[1].g_x[4].t.r_v ;
 wire \g.g_y[1].g_x[5].t.out_sc ;
 wire \g.g_y[1].g_x[5].t.r_d ;
 wire \g.g_y[1].g_x[5].t.r_ghl ;
 wire \g.g_y[1].g_x[5].t.r_gnl ;
 wire \g.g_y[1].g_x[5].t.r_h ;
 wire \g.g_y[1].g_x[5].t.r_v ;
 wire \g.g_y[1].g_x[6].t.out_sc ;
 wire \g.g_y[1].g_x[6].t.r_d ;
 wire \g.g_y[1].g_x[6].t.r_h ;
 wire \g.g_y[1].g_x[6].t.r_v ;
 wire \g.g_y[1].g_x[7].t.out_r ;
 wire \g.g_y[1].g_x[7].t.out_sc ;
 wire \g.g_y[1].g_x[7].t.r_d ;
 wire \g.g_y[1].g_x[7].t.r_ghl ;
 wire \g.g_y[1].g_x[7].t.r_gnl ;
 wire \g.g_y[1].g_x[7].t.r_h ;
 wire \g.g_y[1].g_x[7].t.r_v ;
 wire \g.g_y[2].g_x[0].t.out_sc ;
 wire \g.g_y[2].g_x[0].t.r_d ;
 wire \g.g_y[2].g_x[0].t.r_ghl ;
 wire \g.g_y[2].g_x[0].t.r_gnl ;
 wire \g.g_y[2].g_x[0].t.r_h ;
 wire \g.g_y[2].g_x[0].t.r_v ;
 wire \g.g_y[2].g_x[1].t.out_sc ;
 wire \g.g_y[2].g_x[1].t.r_d ;
 wire \g.g_y[2].g_x[1].t.r_h ;
 wire \g.g_y[2].g_x[1].t.r_v ;
 wire \g.g_y[2].g_x[2].t.out_sc ;
 wire \g.g_y[2].g_x[2].t.r_d ;
 wire \g.g_y[2].g_x[2].t.r_ghl ;
 wire \g.g_y[2].g_x[2].t.r_gnl ;
 wire \g.g_y[2].g_x[2].t.r_h ;
 wire \g.g_y[2].g_x[2].t.r_v ;
 wire \g.g_y[2].g_x[3].t.out_sc ;
 wire \g.g_y[2].g_x[3].t.r_d ;
 wire \g.g_y[2].g_x[3].t.r_h ;
 wire \g.g_y[2].g_x[3].t.r_v ;
 wire \g.g_y[2].g_x[4].t.out_sc ;
 wire \g.g_y[2].g_x[4].t.r_d ;
 wire \g.g_y[2].g_x[4].t.r_ghl ;
 wire \g.g_y[2].g_x[4].t.r_gnl ;
 wire \g.g_y[2].g_x[4].t.r_h ;
 wire \g.g_y[2].g_x[4].t.r_v ;
 wire \g.g_y[2].g_x[5].t.out_sc ;
 wire \g.g_y[2].g_x[5].t.r_d ;
 wire \g.g_y[2].g_x[5].t.r_h ;
 wire \g.g_y[2].g_x[5].t.r_v ;
 wire \g.g_y[2].g_x[6].t.out_sc ;
 wire \g.g_y[2].g_x[6].t.r_d ;
 wire \g.g_y[2].g_x[6].t.r_ghl ;
 wire \g.g_y[2].g_x[6].t.r_gnl ;
 wire \g.g_y[2].g_x[6].t.r_h ;
 wire \g.g_y[2].g_x[6].t.r_v ;
 wire \g.g_y[2].g_x[7].t.out_r ;
 wire \g.g_y[2].g_x[7].t.out_sc ;
 wire \g.g_y[2].g_x[7].t.r_d ;
 wire \g.g_y[2].g_x[7].t.r_h ;
 wire \g.g_y[2].g_x[7].t.r_v ;
 wire \g.g_y[3].g_x[0].t.out_sc ;
 wire \g.g_y[3].g_x[0].t.r_d ;
 wire \g.g_y[3].g_x[0].t.r_h ;
 wire \g.g_y[3].g_x[0].t.r_v ;
 wire \g.g_y[3].g_x[1].t.out_sc ;
 wire \g.g_y[3].g_x[1].t.r_d ;
 wire \g.g_y[3].g_x[1].t.r_ghl ;
 wire \g.g_y[3].g_x[1].t.r_gnl ;
 wire \g.g_y[3].g_x[1].t.r_h ;
 wire \g.g_y[3].g_x[1].t.r_v ;
 wire \g.g_y[3].g_x[2].t.out_sc ;
 wire \g.g_y[3].g_x[2].t.r_d ;
 wire \g.g_y[3].g_x[2].t.r_h ;
 wire \g.g_y[3].g_x[2].t.r_v ;
 wire \g.g_y[3].g_x[3].t.out_sc ;
 wire \g.g_y[3].g_x[3].t.r_d ;
 wire \g.g_y[3].g_x[3].t.r_ghl ;
 wire \g.g_y[3].g_x[3].t.r_gnl ;
 wire \g.g_y[3].g_x[3].t.r_h ;
 wire \g.g_y[3].g_x[3].t.r_v ;
 wire \g.g_y[3].g_x[4].t.out_sc ;
 wire \g.g_y[3].g_x[4].t.r_d ;
 wire \g.g_y[3].g_x[4].t.r_h ;
 wire \g.g_y[3].g_x[4].t.r_v ;
 wire \g.g_y[3].g_x[5].t.out_sc ;
 wire \g.g_y[3].g_x[5].t.r_d ;
 wire \g.g_y[3].g_x[5].t.r_ghl ;
 wire \g.g_y[3].g_x[5].t.r_gnl ;
 wire \g.g_y[3].g_x[5].t.r_h ;
 wire \g.g_y[3].g_x[5].t.r_v ;
 wire \g.g_y[3].g_x[6].t.out_sc ;
 wire \g.g_y[3].g_x[6].t.r_d ;
 wire \g.g_y[3].g_x[6].t.r_h ;
 wire \g.g_y[3].g_x[6].t.r_v ;
 wire \g.g_y[3].g_x[7].t.out_r ;
 wire \g.g_y[3].g_x[7].t.out_sc ;
 wire \g.g_y[3].g_x[7].t.r_d ;
 wire \g.g_y[3].g_x[7].t.r_ghl ;
 wire \g.g_y[3].g_x[7].t.r_gnl ;
 wire \g.g_y[3].g_x[7].t.r_h ;
 wire \g.g_y[3].g_x[7].t.r_v ;
 wire \g.g_y[4].g_x[0].t.out_sc ;
 wire \g.g_y[4].g_x[0].t.r_d ;
 wire \g.g_y[4].g_x[0].t.r_ghl ;
 wire \g.g_y[4].g_x[0].t.r_gnl ;
 wire \g.g_y[4].g_x[0].t.r_h ;
 wire \g.g_y[4].g_x[0].t.r_v ;
 wire \g.g_y[4].g_x[1].t.out_sc ;
 wire \g.g_y[4].g_x[1].t.r_d ;
 wire \g.g_y[4].g_x[1].t.r_h ;
 wire \g.g_y[4].g_x[1].t.r_v ;
 wire \g.g_y[4].g_x[2].t.out_sc ;
 wire \g.g_y[4].g_x[2].t.r_d ;
 wire \g.g_y[4].g_x[2].t.r_ghl ;
 wire \g.g_y[4].g_x[2].t.r_gnl ;
 wire \g.g_y[4].g_x[2].t.r_h ;
 wire \g.g_y[4].g_x[2].t.r_v ;
 wire \g.g_y[4].g_x[3].t.out_sc ;
 wire \g.g_y[4].g_x[3].t.r_d ;
 wire \g.g_y[4].g_x[3].t.r_h ;
 wire \g.g_y[4].g_x[3].t.r_v ;
 wire \g.g_y[4].g_x[4].t.out_sc ;
 wire \g.g_y[4].g_x[4].t.r_d ;
 wire \g.g_y[4].g_x[4].t.r_ghl ;
 wire \g.g_y[4].g_x[4].t.r_gnl ;
 wire \g.g_y[4].g_x[4].t.r_h ;
 wire \g.g_y[4].g_x[4].t.r_v ;
 wire \g.g_y[4].g_x[5].t.out_sc ;
 wire \g.g_y[4].g_x[5].t.r_d ;
 wire \g.g_y[4].g_x[5].t.r_h ;
 wire \g.g_y[4].g_x[5].t.r_v ;
 wire \g.g_y[4].g_x[6].t.out_sc ;
 wire \g.g_y[4].g_x[6].t.r_d ;
 wire \g.g_y[4].g_x[6].t.r_ghl ;
 wire \g.g_y[4].g_x[6].t.r_gnl ;
 wire \g.g_y[4].g_x[6].t.r_h ;
 wire \g.g_y[4].g_x[6].t.r_v ;
 wire \g.g_y[4].g_x[7].t.out_r ;
 wire \g.g_y[4].g_x[7].t.out_sc ;
 wire \g.g_y[4].g_x[7].t.r_d ;
 wire \g.g_y[4].g_x[7].t.r_h ;
 wire \g.g_y[4].g_x[7].t.r_v ;
 wire \g.g_y[5].g_x[0].t.out_sc ;
 wire \g.g_y[5].g_x[0].t.r_d ;
 wire \g.g_y[5].g_x[0].t.r_h ;
 wire \g.g_y[5].g_x[0].t.r_v ;
 wire \g.g_y[5].g_x[1].t.out_sc ;
 wire \g.g_y[5].g_x[1].t.r_d ;
 wire \g.g_y[5].g_x[1].t.r_ghl ;
 wire \g.g_y[5].g_x[1].t.r_gnl ;
 wire \g.g_y[5].g_x[1].t.r_h ;
 wire \g.g_y[5].g_x[1].t.r_v ;
 wire \g.g_y[5].g_x[2].t.out_sc ;
 wire \g.g_y[5].g_x[2].t.r_d ;
 wire \g.g_y[5].g_x[2].t.r_h ;
 wire \g.g_y[5].g_x[2].t.r_v ;
 wire \g.g_y[5].g_x[3].t.out_sc ;
 wire \g.g_y[5].g_x[3].t.r_d ;
 wire \g.g_y[5].g_x[3].t.r_ghl ;
 wire \g.g_y[5].g_x[3].t.r_gnl ;
 wire \g.g_y[5].g_x[3].t.r_h ;
 wire \g.g_y[5].g_x[3].t.r_v ;
 wire \g.g_y[5].g_x[4].t.out_sc ;
 wire \g.g_y[5].g_x[4].t.r_d ;
 wire \g.g_y[5].g_x[4].t.r_h ;
 wire \g.g_y[5].g_x[4].t.r_v ;
 wire \g.g_y[5].g_x[5].t.out_sc ;
 wire \g.g_y[5].g_x[5].t.r_d ;
 wire \g.g_y[5].g_x[5].t.r_ghl ;
 wire \g.g_y[5].g_x[5].t.r_gnl ;
 wire \g.g_y[5].g_x[5].t.r_h ;
 wire \g.g_y[5].g_x[5].t.r_v ;
 wire \g.g_y[5].g_x[6].t.out_sc ;
 wire \g.g_y[5].g_x[6].t.r_d ;
 wire \g.g_y[5].g_x[6].t.r_h ;
 wire \g.g_y[5].g_x[6].t.r_v ;
 wire \g.g_y[5].g_x[7].t.out_r ;
 wire \g.g_y[5].g_x[7].t.out_sc ;
 wire \g.g_y[5].g_x[7].t.r_d ;
 wire \g.g_y[5].g_x[7].t.r_ghl ;
 wire \g.g_y[5].g_x[7].t.r_gnl ;
 wire \g.g_y[5].g_x[7].t.r_h ;
 wire \g.g_y[5].g_x[7].t.r_v ;
 wire \g.g_y[6].g_x[0].t.out_sc ;
 wire \g.g_y[6].g_x[0].t.r_d ;
 wire \g.g_y[6].g_x[0].t.r_ghl ;
 wire \g.g_y[6].g_x[0].t.r_gnl ;
 wire \g.g_y[6].g_x[0].t.r_h ;
 wire \g.g_y[6].g_x[0].t.r_v ;
 wire \g.g_y[6].g_x[1].t.out_sc ;
 wire \g.g_y[6].g_x[1].t.r_d ;
 wire \g.g_y[6].g_x[1].t.r_h ;
 wire \g.g_y[6].g_x[1].t.r_v ;
 wire \g.g_y[6].g_x[2].t.out_sc ;
 wire \g.g_y[6].g_x[2].t.r_d ;
 wire \g.g_y[6].g_x[2].t.r_ghl ;
 wire \g.g_y[6].g_x[2].t.r_gnl ;
 wire \g.g_y[6].g_x[2].t.r_h ;
 wire \g.g_y[6].g_x[2].t.r_v ;
 wire \g.g_y[6].g_x[3].t.out_sc ;
 wire \g.g_y[6].g_x[3].t.r_d ;
 wire \g.g_y[6].g_x[3].t.r_h ;
 wire \g.g_y[6].g_x[3].t.r_v ;
 wire \g.g_y[6].g_x[4].t.out_sc ;
 wire \g.g_y[6].g_x[4].t.r_d ;
 wire \g.g_y[6].g_x[4].t.r_ghl ;
 wire \g.g_y[6].g_x[4].t.r_gnl ;
 wire \g.g_y[6].g_x[4].t.r_h ;
 wire \g.g_y[6].g_x[4].t.r_v ;
 wire \g.g_y[6].g_x[5].t.out_sc ;
 wire \g.g_y[6].g_x[5].t.r_d ;
 wire \g.g_y[6].g_x[5].t.r_h ;
 wire \g.g_y[6].g_x[5].t.r_v ;
 wire \g.g_y[6].g_x[6].t.out_sc ;
 wire \g.g_y[6].g_x[6].t.r_d ;
 wire \g.g_y[6].g_x[6].t.r_ghl ;
 wire \g.g_y[6].g_x[6].t.r_gnl ;
 wire \g.g_y[6].g_x[6].t.r_h ;
 wire \g.g_y[6].g_x[6].t.r_v ;
 wire \g.g_y[6].g_x[7].t.out_r ;
 wire \g.g_y[6].g_x[7].t.out_sc ;
 wire \g.g_y[6].g_x[7].t.r_d ;
 wire \g.g_y[6].g_x[7].t.r_h ;
 wire \g.g_y[6].g_x[7].t.r_v ;
 wire \g.g_y[7].g_x[0].t.out_sc ;
 wire \g.g_y[7].g_x[0].t.r_d ;
 wire \g.g_y[7].g_x[0].t.r_h ;
 wire \g.g_y[7].g_x[0].t.r_v ;
 wire \g.g_y[7].g_x[1].t.out_sc ;
 wire \g.g_y[7].g_x[1].t.r_d ;
 wire \g.g_y[7].g_x[1].t.r_ghl ;
 wire \g.g_y[7].g_x[1].t.r_gnl ;
 wire \g.g_y[7].g_x[1].t.r_h ;
 wire \g.g_y[7].g_x[1].t.r_v ;
 wire \g.g_y[7].g_x[2].t.out_sc ;
 wire \g.g_y[7].g_x[2].t.r_d ;
 wire \g.g_y[7].g_x[2].t.r_h ;
 wire \g.g_y[7].g_x[2].t.r_v ;
 wire \g.g_y[7].g_x[3].t.out_sc ;
 wire \g.g_y[7].g_x[3].t.r_d ;
 wire \g.g_y[7].g_x[3].t.r_ghl ;
 wire \g.g_y[7].g_x[3].t.r_gnl ;
 wire \g.g_y[7].g_x[3].t.r_h ;
 wire \g.g_y[7].g_x[3].t.r_v ;
 wire \g.g_y[7].g_x[4].t.out_sc ;
 wire \g.g_y[7].g_x[4].t.r_d ;
 wire \g.g_y[7].g_x[4].t.r_h ;
 wire \g.g_y[7].g_x[4].t.r_v ;
 wire \g.g_y[7].g_x[5].t.out_sc ;
 wire \g.g_y[7].g_x[5].t.r_d ;
 wire \g.g_y[7].g_x[5].t.r_ghl ;
 wire \g.g_y[7].g_x[5].t.r_gnl ;
 wire \g.g_y[7].g_x[5].t.r_h ;
 wire \g.g_y[7].g_x[5].t.r_v ;
 wire \g.g_y[7].g_x[6].t.out_sc ;
 wire \g.g_y[7].g_x[6].t.r_d ;
 wire \g.g_y[7].g_x[6].t.r_h ;
 wire \g.g_y[7].g_x[6].t.r_v ;
 wire \g.g_y[7].g_x[7].t.out_r ;
 wire \g.g_y[7].g_x[7].t.out_sc ;
 wire \g.g_y[7].g_x[7].t.r_d ;
 wire \g.g_y[7].g_x[7].t.r_ghl ;
 wire \g.g_y[7].g_x[7].t.r_gnl ;
 wire \g.g_y[7].g_x[7].t.r_h ;
 wire \g.g_y[7].g_x[7].t.r_v ;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net180;
 wire net181;
 wire net182;
 wire net183;
 wire net184;
 wire net185;
 wire net186;
 wire net187;
 wire net188;
 wire net189;
 wire net190;
 wire net191;
 wire net192;
 wire net193;
 wire net194;
 wire net195;
 wire net196;
 wire net197;
 wire net198;
 wire net200;
 wire net201;
 wire net202;
 wire net203;
 wire net204;
 wire net205;
 wire net206;
 wire net207;
 wire net208;
 wire net209;
 wire net210;
 wire net211;
 wire net212;
 wire net213;
 wire net214;
 wire net215;
 wire net216;
 wire net217;
 wire net218;
 wire net219;
 wire net220;
 wire net221;
 wire net222;
 wire net223;
 wire net224;
 wire net225;
 wire net226;
 wire net227;
 wire net228;
 wire net229;
 wire net230;
 wire net231;
 wire net232;
 wire net233;
 wire net234;
 wire net235;
 wire net236;
 wire net237;
 wire net238;
 wire net239;
 wire net240;
 wire net241;
 wire net242;
 wire net243;
 wire net244;
 wire net245;
 wire net246;
 wire net247;
 wire net248;
 wire net249;
 wire net250;
 wire net251;
 wire net252;
 wire net253;
 wire net254;
 wire net255;
 wire net256;
 wire net257;
 wire net258;
 wire net259;
 wire net260;
 wire net261;
 wire net262;
 wire net263;
 wire net264;
 wire net265;
 wire net266;
 wire net267;
 wire net268;
 wire net269;
 wire net270;
 wire net271;
 wire net272;
 wire net273;
 wire net274;
 wire net275;
 wire net276;
 wire net277;
 wire net278;
 wire net279;
 wire net280;
 wire net281;
 wire net282;
 wire net283;
 wire net284;
 wire net285;
 wire net286;
 wire net287;
 wire net288;
 wire net289;
 wire net290;
 wire net291;
 wire net292;
 wire net293;
 wire net294;
 wire net295;
 wire net296;
 wire net297;
 wire net298;
 wire net299;
 wire net300;
 wire net301;
 wire net302;
 wire net303;
 wire net304;
 wire net305;
 wire net306;
 wire net307;
 wire net308;
 wire net309;
 wire net310;
 wire net311;
 wire net312;
 wire net313;
 wire net314;
 wire net315;
 wire net316;
 wire net317;
 wire net318;
 wire net319;
 wire net320;
 wire net321;
 wire net322;
 wire net323;
 wire net324;
 wire net325;
 wire net326;
 wire net327;
 wire net328;
 wire net329;
 wire net330;
 wire net331;
 wire net332;
 wire net333;
 wire net334;
 wire net335;
 wire net336;
 wire net337;
 wire net338;
 wire net339;
 wire net340;
 wire net341;
 wire net342;
 wire net343;
 wire net344;
 wire net345;
 wire net346;
 wire net347;
 wire net348;
 wire net349;
 wire net350;
 wire net351;
 wire net352;
 wire net353;
 wire net354;
 wire net355;
 wire net356;
 wire net357;
 wire net358;
 wire net359;
 wire net360;
 wire net361;
 wire net362;
 wire net363;
 wire net364;
 wire net365;
 wire net366;
 wire net367;
 wire net368;
 wire net369;
 wire net370;
 wire net371;
 wire net372;
 wire net373;
 wire net374;
 wire net375;
 wire net376;
 wire net377;
 wire net378;
 wire net379;
 wire net380;
 wire net381;
 wire net382;
 wire net383;
 wire net384;
 wire net385;
 wire net386;
 wire net387;
 wire net388;
 wire net389;
 wire net390;
 wire net391;
 wire net392;
 wire net393;
 wire net394;
 wire net395;
 wire net396;
 wire net397;
 wire net398;
 wire net399;
 wire net400;
 wire net401;
 wire net402;
 wire net403;
 wire net404;
 wire net405;
 wire net406;
 wire net407;
 wire net408;
 wire net409;
 wire net410;
 wire net411;
 wire net412;
 wire net413;
 wire net414;
 wire net415;
 wire net416;
 wire net417;
 wire net418;
 wire net419;
 wire net420;
 wire net421;
 wire net422;
 wire net423;
 wire net424;
 wire net425;
 wire net426;
 wire net427;
 wire net428;
 wire net429;
 wire net430;
 wire net431;
 wire net432;
 wire net433;
 wire net434;
 wire net435;
 wire net436;
 wire net437;
 wire net438;
 wire net439;
 wire net440;
 wire net441;
 wire net442;
 wire net443;
 wire net444;
 wire net445;
 wire net446;
 wire net447;
 wire net448;
 wire net449;
 wire net450;
 wire net451;
 wire net452;
 wire net453;
 wire net454;
 wire net455;
 wire net456;
 wire net457;
 wire net458;
 wire net459;
 wire net460;
 wire net461;
 wire net462;
 wire net463;
 wire net464;
 wire net465;
 wire net466;
 wire net467;
 wire net468;
 wire net469;
 wire net470;
 wire net471;
 wire net472;
 wire net473;
 wire net474;
 wire net475;
 wire net476;
 wire net477;
 wire net478;
 wire net479;
 wire net480;
 wire net481;
 wire net482;
 wire net483;
 wire net484;
 wire net485;
 wire net486;
 wire net487;
 wire net488;
 wire net489;
 wire net490;
 wire net491;
 wire net492;
 wire net493;
 wire net494;
 wire net495;
 wire net496;
 wire net497;
 wire net498;
 wire net499;
 wire net500;
 wire net501;
 wire net502;
 wire net503;
 wire net504;
 wire net505;
 wire net506;
 wire net507;
 wire net508;
 wire net509;
 wire net510;
 wire net511;
 wire net512;
 wire net513;
 wire net514;
 wire net515;
 wire net516;
 wire net517;
 wire net518;
 wire net519;
 wire clknet_leaf_1_clk;
 wire clknet_leaf_2_clk;
 wire clknet_leaf_3_clk;
 wire clknet_leaf_4_clk;
 wire clknet_leaf_5_clk;
 wire clknet_leaf_6_clk;
 wire clknet_leaf_7_clk;
 wire clknet_leaf_8_clk;
 wire clknet_leaf_9_clk;
 wire clknet_leaf_10_clk;
 wire clknet_leaf_11_clk;
 wire clknet_leaf_12_clk;
 wire clknet_leaf_13_clk;
 wire clknet_leaf_14_clk;
 wire clknet_leaf_15_clk;
 wire clknet_leaf_16_clk;
 wire clknet_leaf_17_clk;
 wire clknet_leaf_18_clk;
 wire clknet_leaf_19_clk;
 wire clknet_leaf_20_clk;
 wire clknet_leaf_21_clk;
 wire clknet_leaf_22_clk;
 wire clknet_leaf_23_clk;
 wire clknet_leaf_24_clk;
 wire clknet_leaf_25_clk;
 wire clknet_leaf_26_clk;
 wire clknet_leaf_27_clk;
 wire clknet_leaf_28_clk;
 wire clknet_leaf_29_clk;
 wire clknet_leaf_30_clk;
 wire clknet_leaf_31_clk;
 wire clknet_leaf_32_clk;
 wire clknet_leaf_33_clk;
 wire clknet_leaf_34_clk;
 wire clknet_leaf_35_clk;
 wire clknet_leaf_36_clk;
 wire clknet_leaf_37_clk;
 wire clknet_leaf_38_clk;
 wire clknet_leaf_39_clk;
 wire clknet_0_clk;
 wire clknet_3_0__leaf_clk;
 wire clknet_3_1__leaf_clk;
 wire clknet_3_2__leaf_clk;
 wire clknet_3_3__leaf_clk;
 wire clknet_3_4__leaf_clk;
 wire clknet_3_5__leaf_clk;
 wire clknet_3_6__leaf_clk;
 wire clknet_3_7__leaf_clk;

 sg13g2_buf_1 _3220_ (.A(rst_n),
    .X(_2581_));
 sg13g2_buf_1 _3221_ (.A(net184),
    .X(_2582_));
 sg13g2_buf_1 _3222_ (.A(net181),
    .X(_2583_));
 sg13g2_buf_2 _3223_ (.A(\g.g_y[0].g_x[0].t.out_sc ),
    .X(_2584_));
 sg13g2_buf_2 _3224_ (.A(\g.g_y[0].g_x[0].t.r_d ),
    .X(_2585_));
 sg13g2_buf_1 _3225_ (.A(uio_in[0]),
    .X(_2586_));
 sg13g2_buf_1 _3226_ (.A(uio_in[6]),
    .X(_2587_));
 sg13g2_nand2_1 _3227_ (.Y(_2588_),
    .A(net183),
    .B(net182));
 sg13g2_buf_2 _3228_ (.A(_2588_),
    .X(_2589_));
 sg13g2_nand2_1 _3229_ (.Y(_2590_),
    .A(net10),
    .B(net11));
 sg13g2_or2_1 _3230_ (.X(_2591_),
    .B(_2590_),
    .A(_2589_));
 sg13g2_buf_1 _3231_ (.A(_2591_),
    .X(_2592_));
 sg13g2_buf_1 _3232_ (.A(_2592_),
    .X(_2593_));
 sg13g2_mux2_1 _3233_ (.A0(_2584_),
    .A1(_2585_),
    .S(net47),
    .X(_2594_));
 sg13g2_and2_1 _3234_ (.A(net131),
    .B(_2594_),
    .X(_0000_));
 sg13g2_inv_1 _3235_ (.Y(_2595_),
    .A(net183));
 sg13g2_o21ai_1 _3236_ (.B1(_2595_),
    .Y(_2596_),
    .A1(net10),
    .A2(net11));
 sg13g2_and2_1 _3237_ (.A(net182),
    .B(_2596_),
    .X(_2597_));
 sg13g2_buf_2 _3238_ (.A(_2597_),
    .X(_2598_));
 sg13g2_buf_1 _3239_ (.A(_2598_),
    .X(_2599_));
 sg13g2_buf_1 _3240_ (.A(\g.g_y[0].g_x[0].t.r_h ),
    .X(_2600_));
 sg13g2_buf_1 _3241_ (.A(\g.g_y[0].g_x[1].t.r_d ),
    .X(_2601_));
 sg13g2_buf_1 _3242_ (.A(\g.g_y[7].g_x[1].t.r_ghl ),
    .X(_2602_));
 sg13g2_buf_2 _3243_ (.A(\g.g_y[7].g_x[1].t.out_sc ),
    .X(_2603_));
 sg13g2_buf_2 _3244_ (.A(\g.g_y[7].g_x[1].t.r_d ),
    .X(_2604_));
 sg13g2_mux2_1 _3245_ (.A0(\g.g_y[7].g_x[1].t.r_gnl ),
    .A1(_2603_),
    .S(_2604_),
    .X(_2605_));
 sg13g2_buf_2 _3246_ (.A(\g.g_y[7].g_x[1].t.r_v ),
    .X(_2606_));
 sg13g2_mux2_1 _3247_ (.A0(_2602_),
    .A1(_2605_),
    .S(_2606_),
    .X(_2607_));
 sg13g2_buf_2 _3248_ (.A(\g.g_y[1].g_x[1].t.out_sc ),
    .X(_2608_));
 sg13g2_buf_2 _3249_ (.A(\g.g_y[1].g_x[1].t.r_d ),
    .X(_2609_));
 sg13g2_mux2_1 _3250_ (.A0(\g.g_y[1].g_x[1].t.r_gnl ),
    .A1(_2608_),
    .S(_2609_),
    .X(_2610_));
 sg13g2_buf_1 _3251_ (.A(\g.g_y[1].g_x[1].t.r_ghl ),
    .X(_2611_));
 sg13g2_buf_2 _3252_ (.A(\g.g_y[1].g_x[1].t.r_v ),
    .X(_2612_));
 sg13g2_mux2_1 _3253_ (.A0(_2610_),
    .A1(_2611_),
    .S(_2612_),
    .X(_2613_));
 sg13g2_buf_1 _3254_ (.A(\g.g_y[0].g_x[1].t.r_v ),
    .X(_2614_));
 sg13g2_inv_1 _3255_ (.Y(_2615_),
    .A(_2614_));
 sg13g2_mux2_1 _3256_ (.A0(_2607_),
    .A1(_2613_),
    .S(_2615_),
    .X(_2616_));
 sg13g2_buf_1 _3257_ (.A(\g.g_y[0].g_x[0].t.r_ghl ),
    .X(_2617_));
 sg13g2_mux2_1 _3258_ (.A0(_2584_),
    .A1(\g.g_y[0].g_x[0].t.r_gnl ),
    .S(_2585_),
    .X(_2618_));
 sg13g2_mux2_1 _3259_ (.A0(_2617_),
    .A1(_2618_),
    .S(net180),
    .X(_2619_));
 sg13g2_buf_2 _3260_ (.A(\g.g_y[0].g_x[2].t.out_sc ),
    .X(_2620_));
 sg13g2_buf_2 _3261_ (.A(\g.g_y[0].g_x[2].t.r_d ),
    .X(_2621_));
 sg13g2_mux2_1 _3262_ (.A0(_2620_),
    .A1(\g.g_y[0].g_x[2].t.r_gnl ),
    .S(_2621_),
    .X(_2622_));
 sg13g2_buf_1 _3263_ (.A(\g.g_y[0].g_x[2].t.r_ghl ),
    .X(_2623_));
 sg13g2_buf_2 _3264_ (.A(\g.g_y[0].g_x[2].t.r_h ),
    .X(_2624_));
 sg13g2_mux2_1 _3265_ (.A0(_2622_),
    .A1(_2623_),
    .S(_2624_),
    .X(_2625_));
 sg13g2_buf_1 _3266_ (.A(\g.g_y[0].g_x[1].t.r_h ),
    .X(_2626_));
 sg13g2_inv_1 _3267_ (.Y(_2627_),
    .A(_2626_));
 sg13g2_mux2_1 _3268_ (.A0(_2619_),
    .A1(_2625_),
    .S(_2627_),
    .X(_2628_));
 sg13g2_nand3_1 _3269_ (.B(_2616_),
    .C(_2628_),
    .A(_2601_),
    .Y(_2629_));
 sg13g2_buf_2 _3270_ (.A(\g.g_y[0].g_x[1].t.out_sc ),
    .X(_2630_));
 sg13g2_nor2_1 _3271_ (.A(_2630_),
    .B(net179),
    .Y(_2631_));
 sg13g2_nor2_1 _3272_ (.A(_2626_),
    .B(_2631_),
    .Y(_2632_));
 sg13g2_mux2_1 _3273_ (.A0(_2607_),
    .A1(_2613_),
    .S(_2614_),
    .X(_2633_));
 sg13g2_mux2_1 _3274_ (.A0(_2625_),
    .A1(_2633_),
    .S(net179),
    .X(_2634_));
 sg13g2_a22oi_1 _3275_ (.Y(_2635_),
    .B1(_2634_),
    .B2(_2626_),
    .A2(_2632_),
    .A1(_2629_));
 sg13g2_nor2_1 _3276_ (.A(net180),
    .B(net1),
    .Y(_2636_));
 sg13g2_a21o_1 _3277_ (.A2(_2635_),
    .A1(net180),
    .B1(_2636_),
    .X(_2637_));
 sg13g2_buf_1 _3278_ (.A(\g.g_y[7].g_x[0].t.r_d ),
    .X(_2638_));
 sg13g2_buf_1 _3279_ (.A(_2638_),
    .X(_2639_));
 sg13g2_mux2_1 _3280_ (.A0(_2603_),
    .A1(\g.g_y[7].g_x[1].t.r_gnl ),
    .S(_2604_),
    .X(_2640_));
 sg13g2_buf_2 _3281_ (.A(\g.g_y[7].g_x[1].t.r_h ),
    .X(_2641_));
 sg13g2_mux2_1 _3282_ (.A0(_2640_),
    .A1(_2602_),
    .S(_2641_),
    .X(_2642_));
 sg13g2_buf_1 _3283_ (.A(_2642_),
    .X(_2643_));
 sg13g2_buf_2 _3284_ (.A(\g.g_y[7].g_x[0].t.r_h ),
    .X(_2644_));
 sg13g2_mux2_1 _3285_ (.A0(net8),
    .A1(_2643_),
    .S(_2644_),
    .X(_2645_));
 sg13g2_or2_1 _3286_ (.X(_2646_),
    .B(_2645_),
    .A(net130));
 sg13g2_buf_1 _3287_ (.A(\g.g_y[6].g_x[0].t.r_v ),
    .X(_2647_));
 sg13g2_buf_2 _3288_ (.A(\g.g_y[6].g_x[0].t.out_sc ),
    .X(_2648_));
 sg13g2_buf_2 _3289_ (.A(\g.g_y[6].g_x[0].t.r_d ),
    .X(_2649_));
 sg13g2_mux2_1 _3290_ (.A0(\g.g_y[6].g_x[0].t.r_gnl ),
    .A1(_2648_),
    .S(_2649_),
    .X(_2650_));
 sg13g2_buf_1 _3291_ (.A(_2650_),
    .X(_2651_));
 sg13g2_buf_1 _3292_ (.A(\g.g_y[6].g_x[0].t.r_ghl ),
    .X(_2652_));
 sg13g2_nor2b_1 _3293_ (.A(net178),
    .B_N(_2652_),
    .Y(_2653_));
 sg13g2_a21oi_1 _3294_ (.A1(net178),
    .A2(_2651_),
    .Y(_2654_),
    .B1(_2653_));
 sg13g2_buf_2 _3295_ (.A(\g.g_y[7].g_x[0].t.r_v ),
    .X(_2655_));
 sg13g2_a21oi_1 _3296_ (.A1(net130),
    .A2(_2654_),
    .Y(_2656_),
    .B1(_2655_));
 sg13g2_mux2_1 _3297_ (.A0(_2643_),
    .A1(net8),
    .S(_2644_),
    .X(_2657_));
 sg13g2_nor2_1 _3298_ (.A(_2638_),
    .B(_2654_),
    .Y(_2658_));
 sg13g2_buf_2 _3299_ (.A(\g.g_y[7].g_x[0].t.out_sc ),
    .X(_2659_));
 sg13g2_nor2b_1 _3300_ (.A(_2659_),
    .B_N(_2638_),
    .Y(_2660_));
 sg13g2_a21oi_1 _3301_ (.A1(_2657_),
    .A2(_2658_),
    .Y(_2661_),
    .B1(_2660_));
 sg13g2_a22oi_1 _3302_ (.Y(_2662_),
    .B1(_2661_),
    .B2(_2655_),
    .A2(_2656_),
    .A1(_2646_));
 sg13g2_buf_2 _3303_ (.A(\g.g_y[1].g_x[0].t.r_v ),
    .X(_2663_));
 sg13g2_mux2_1 _3304_ (.A0(_2608_),
    .A1(\g.g_y[1].g_x[1].t.r_gnl ),
    .S(_2609_),
    .X(_2664_));
 sg13g2_buf_2 _3305_ (.A(\g.g_y[1].g_x[1].t.r_h ),
    .X(_2665_));
 sg13g2_mux2_1 _3306_ (.A0(_2664_),
    .A1(_2611_),
    .S(_2665_),
    .X(_2666_));
 sg13g2_buf_1 _3307_ (.A(_2666_),
    .X(_2667_));
 sg13g2_buf_2 _3308_ (.A(\g.g_y[1].g_x[0].t.r_h ),
    .X(_2668_));
 sg13g2_mux2_1 _3309_ (.A0(net2),
    .A1(_2667_),
    .S(_2668_),
    .X(_2669_));
 sg13g2_buf_2 _3310_ (.A(\g.g_y[2].g_x[0].t.out_sc ),
    .X(_2670_));
 sg13g2_buf_2 _3311_ (.A(\g.g_y[2].g_x[0].t.r_d ),
    .X(_2671_));
 sg13g2_mux2_1 _3312_ (.A0(\g.g_y[2].g_x[0].t.r_gnl ),
    .A1(_2670_),
    .S(_2671_),
    .X(_2672_));
 sg13g2_buf_1 _3313_ (.A(\g.g_y[2].g_x[0].t.r_ghl ),
    .X(_2673_));
 sg13g2_buf_2 _3314_ (.A(\g.g_y[2].g_x[0].t.r_v ),
    .X(_2674_));
 sg13g2_mux2_1 _3315_ (.A0(_2672_),
    .A1(_2673_),
    .S(_2674_),
    .X(_2675_));
 sg13g2_buf_1 _3316_ (.A(_2675_),
    .X(_2676_));
 sg13g2_buf_2 _3317_ (.A(\g.g_y[1].g_x[0].t.r_d ),
    .X(_2677_));
 sg13g2_mux2_1 _3318_ (.A0(_2669_),
    .A1(_2676_),
    .S(_2677_),
    .X(_2678_));
 sg13g2_inv_2 _3319_ (.Y(_2679_),
    .A(_2677_));
 sg13g2_mux2_1 _3320_ (.A0(_2667_),
    .A1(net2),
    .S(_2668_),
    .X(_2680_));
 sg13g2_nand3_1 _3321_ (.B(_2676_),
    .C(_2680_),
    .A(_2679_),
    .Y(_2681_));
 sg13g2_buf_2 _3322_ (.A(\g.g_y[1].g_x[0].t.out_sc ),
    .X(_2682_));
 sg13g2_nor2_1 _3323_ (.A(_2679_),
    .B(_2682_),
    .Y(_2683_));
 sg13g2_nor2_1 _3324_ (.A(_2663_),
    .B(_2683_),
    .Y(_2684_));
 sg13g2_a22oi_1 _3325_ (.Y(_2685_),
    .B1(_2681_),
    .B2(_2684_),
    .A2(_2678_),
    .A1(_2663_));
 sg13g2_buf_2 _3326_ (.A(\g.g_y[0].g_x[0].t.r_v ),
    .X(_2686_));
 sg13g2_mux2_1 _3327_ (.A0(_2662_),
    .A1(_2685_),
    .S(_2686_),
    .X(_2687_));
 sg13g2_mux2_1 _3328_ (.A0(_2637_),
    .A1(_2687_),
    .S(_2585_),
    .X(_2688_));
 sg13g2_buf_1 _3329_ (.A(_2598_),
    .X(_2689_));
 sg13g2_buf_1 _3330_ (.A(net184),
    .X(_2690_));
 sg13g2_o21ai_1 _3331_ (.B1(net177),
    .Y(_2691_),
    .A1(_2617_),
    .A2(net45));
 sg13g2_a21oi_1 _3332_ (.A1(net46),
    .A2(_2688_),
    .Y(_0001_),
    .B1(_2691_));
 sg13g2_nor2b_1 _3333_ (.A(net1),
    .B_N(net180),
    .Y(_2692_));
 sg13g2_nor2b_1 _3334_ (.A(_2600_),
    .B_N(_2635_),
    .Y(_2693_));
 sg13g2_mux2_1 _3335_ (.A0(_2685_),
    .A1(_2662_),
    .S(_2686_),
    .X(_2694_));
 sg13g2_nor3_1 _3336_ (.A(_2692_),
    .B(_2693_),
    .C(_2694_),
    .Y(_2695_));
 sg13g2_buf_1 _3337_ (.A(_2581_),
    .X(_2696_));
 sg13g2_o21ai_1 _3338_ (.B1(net176),
    .Y(_2697_),
    .A1(\g.g_y[0].g_x[0].t.r_gnl ),
    .A2(_2689_));
 sg13g2_a21oi_1 _3339_ (.A1(net46),
    .A2(_2695_),
    .Y(_0002_),
    .B1(_2697_));
 sg13g2_nand2b_1 _3340_ (.Y(_2698_),
    .B(net11),
    .A_N(net10));
 sg13g2_buf_1 _3341_ (.A(_2698_),
    .X(_2699_));
 sg13g2_nor2_1 _3342_ (.A(_2589_),
    .B(_2699_),
    .Y(_2700_));
 sg13g2_buf_2 _3343_ (.A(_2700_),
    .X(_2701_));
 sg13g2_buf_1 _3344_ (.A(net66),
    .X(_2702_));
 sg13g2_nand2_1 _3345_ (.Y(_2703_),
    .A(_2584_),
    .B(net44));
 sg13g2_buf_1 _3346_ (.A(_2589_),
    .X(_2704_));
 sg13g2_buf_1 _3347_ (.A(net99),
    .X(_2705_));
 sg13g2_buf_1 _3348_ (.A(_2699_),
    .X(_2706_));
 sg13g2_buf_1 _3349_ (.A(_2706_),
    .X(_2707_));
 sg13g2_o21ai_1 _3350_ (.B1(net180),
    .Y(_2708_),
    .A1(net65),
    .A2(net98));
 sg13g2_inv_2 _3351_ (.Y(_2709_),
    .A(net184));
 sg13g2_buf_1 _3352_ (.A(_2709_),
    .X(_2710_));
 sg13g2_buf_1 _3353_ (.A(net128),
    .X(_2711_));
 sg13g2_a21oi_1 _3354_ (.A1(_2703_),
    .A2(_2708_),
    .Y(_0003_),
    .B1(net97));
 sg13g2_buf_1 _3355_ (.A(uio_in[5]),
    .X(_2712_));
 sg13g2_nand2_2 _3356_ (.Y(_2713_),
    .A(_2712_),
    .B(net184));
 sg13g2_nand2b_1 _3357_ (.Y(_2714_),
    .B(_2595_),
    .A_N(_2713_));
 sg13g2_buf_2 _3358_ (.A(_2714_),
    .X(_2715_));
 sg13g2_buf_1 _3359_ (.A(_2715_),
    .X(_2716_));
 sg13g2_mux2_1 _3360_ (.A0(_2687_),
    .A1(_2637_),
    .S(_2585_),
    .X(_2717_));
 sg13g2_nor2_1 _3361_ (.A(_2712_),
    .B(_2709_),
    .Y(_2718_));
 sg13g2_buf_8 _3362_ (.A(_2718_),
    .X(_2719_));
 sg13g2_buf_8 _3363_ (.A(_2719_),
    .X(_2720_));
 sg13g2_nor2_1 _3364_ (.A(_2595_),
    .B(_2713_),
    .Y(_2721_));
 sg13g2_buf_1 _3365_ (.A(_2721_),
    .X(_2722_));
 sg13g2_buf_1 _3366_ (.A(net96),
    .X(_2723_));
 sg13g2_a22oi_1 _3367_ (.Y(_2724_),
    .B1(net62),
    .B2(net9),
    .A2(net63),
    .A1(_2584_));
 sg13g2_o21ai_1 _3368_ (.B1(_2724_),
    .Y(_0004_),
    .A1(net64),
    .A2(_2717_));
 sg13g2_nand2b_1 _3369_ (.Y(_2725_),
    .B(net10),
    .A_N(net11));
 sg13g2_buf_1 _3370_ (.A(_2725_),
    .X(_2726_));
 sg13g2_nor2_1 _3371_ (.A(_2589_),
    .B(_2726_),
    .Y(_2727_));
 sg13g2_buf_2 _3372_ (.A(_2727_),
    .X(_2728_));
 sg13g2_buf_1 _3373_ (.A(_2728_),
    .X(_2729_));
 sg13g2_nand2_1 _3374_ (.Y(_2730_),
    .A(_2584_),
    .B(net43));
 sg13g2_buf_1 _3375_ (.A(_2726_),
    .X(_2731_));
 sg13g2_buf_1 _3376_ (.A(net127),
    .X(_2732_));
 sg13g2_o21ai_1 _3377_ (.B1(_2686_),
    .Y(_2733_),
    .A1(net65),
    .A2(net95));
 sg13g2_a21oi_1 _3378_ (.A1(_2730_),
    .A2(_2733_),
    .Y(_0005_),
    .B1(net97));
 sg13g2_mux2_1 _3379_ (.A0(_2630_),
    .A1(net179),
    .S(net47),
    .X(_2734_));
 sg13g2_and2_1 _3380_ (.A(net131),
    .B(_2734_),
    .X(_0006_));
 sg13g2_nand2_1 _3381_ (.Y(_2735_),
    .A(_2630_),
    .B(net44));
 sg13g2_o21ai_1 _3382_ (.B1(_2626_),
    .Y(_2736_),
    .A1(net65),
    .A2(net98));
 sg13g2_a21oi_1 _3383_ (.A1(_2735_),
    .A2(_2736_),
    .Y(_0007_),
    .B1(net97));
 sg13g2_buf_1 _3384_ (.A(_2709_),
    .X(_2737_));
 sg13g2_buf_1 _3385_ (.A(net126),
    .X(_2738_));
 sg13g2_buf_1 _3386_ (.A(_2712_),
    .X(_2739_));
 sg13g2_buf_1 _3387_ (.A(net175),
    .X(_2740_));
 sg13g2_mux2_1 _3388_ (.A0(_2619_),
    .A1(_2625_),
    .S(_2626_),
    .X(_2741_));
 sg13g2_mux2_1 _3389_ (.A0(_2633_),
    .A1(_2741_),
    .S(net179),
    .X(_2742_));
 sg13g2_buf_1 _3390_ (.A(_2595_),
    .X(_2743_));
 sg13g2_mux2_1 _3391_ (.A0(_2584_),
    .A1(_2742_),
    .S(net124),
    .X(_2744_));
 sg13g2_buf_1 _3392_ (.A(net175),
    .X(_2745_));
 sg13g2_nor2b_1 _3393_ (.A(net123),
    .B_N(_2630_),
    .Y(_2746_));
 sg13g2_a21oi_1 _3394_ (.A1(net125),
    .A2(_2744_),
    .Y(_2747_),
    .B1(_2746_));
 sg13g2_nor2_1 _3395_ (.A(net94),
    .B(_2747_),
    .Y(_0008_));
 sg13g2_nand2_1 _3396_ (.Y(_2748_),
    .A(_2630_),
    .B(_2729_));
 sg13g2_o21ai_1 _3397_ (.B1(_2614_),
    .Y(_2749_),
    .A1(_2705_),
    .A2(_2732_));
 sg13g2_a21oi_1 _3398_ (.A1(_2748_),
    .A2(_2749_),
    .Y(_0009_),
    .B1(net97));
 sg13g2_mux2_1 _3399_ (.A0(_2620_),
    .A1(_2621_),
    .S(_2593_),
    .X(_2750_));
 sg13g2_and2_1 _3400_ (.A(_2583_),
    .B(_2750_),
    .X(_0010_));
 sg13g2_o21ai_1 _3401_ (.B1(net12),
    .Y(_2751_),
    .A1(_2586_),
    .A2(_2590_));
 sg13g2_and2_1 _3402_ (.A(net182),
    .B(_2751_),
    .X(_2752_));
 sg13g2_buf_2 _3403_ (.A(_2752_),
    .X(_2753_));
 sg13g2_buf_1 _3404_ (.A(_2753_),
    .X(_2754_));
 sg13g2_nor2_1 _3405_ (.A(_2627_),
    .B(_2631_),
    .Y(_2755_));
 sg13g2_mux2_1 _3406_ (.A0(_2619_),
    .A1(_2633_),
    .S(net179),
    .X(_2756_));
 sg13g2_a22oi_1 _3407_ (.Y(_2757_),
    .B1(_2756_),
    .B2(_2627_),
    .A2(_2755_),
    .A1(_2629_));
 sg13g2_buf_2 _3408_ (.A(\g.g_y[0].g_x[3].t.r_d ),
    .X(_2758_));
 sg13g2_buf_2 _3409_ (.A(\g.g_y[7].g_x[3].t.r_v ),
    .X(_2759_));
 sg13g2_buf_2 _3410_ (.A(\g.g_y[7].g_x[3].t.out_sc ),
    .X(_2760_));
 sg13g2_buf_2 _3411_ (.A(\g.g_y[7].g_x[3].t.r_d ),
    .X(_2761_));
 sg13g2_mux2_1 _3412_ (.A0(\g.g_y[7].g_x[3].t.r_gnl ),
    .A1(_2760_),
    .S(_2761_),
    .X(_2762_));
 sg13g2_buf_1 _3413_ (.A(\g.g_y[7].g_x[3].t.r_ghl ),
    .X(_2763_));
 sg13g2_nor2b_1 _3414_ (.A(_2759_),
    .B_N(_2763_),
    .Y(_2764_));
 sg13g2_a21o_1 _3415_ (.A2(_2762_),
    .A1(_2759_),
    .B1(_2764_),
    .X(_2765_));
 sg13g2_buf_2 _3416_ (.A(\g.g_y[1].g_x[3].t.out_sc ),
    .X(_2766_));
 sg13g2_buf_2 _3417_ (.A(\g.g_y[1].g_x[3].t.r_d ),
    .X(_2767_));
 sg13g2_mux2_1 _3418_ (.A0(\g.g_y[1].g_x[3].t.r_gnl ),
    .A1(_2766_),
    .S(_2767_),
    .X(_2768_));
 sg13g2_buf_1 _3419_ (.A(_2768_),
    .X(_2769_));
 sg13g2_buf_1 _3420_ (.A(\g.g_y[1].g_x[3].t.r_ghl ),
    .X(_2770_));
 sg13g2_buf_1 _3421_ (.A(\g.g_y[1].g_x[3].t.r_v ),
    .X(_2771_));
 sg13g2_mux2_1 _3422_ (.A0(_2769_),
    .A1(_2770_),
    .S(_2771_),
    .X(_2772_));
 sg13g2_buf_1 _3423_ (.A(\g.g_y[0].g_x[3].t.r_v ),
    .X(_2773_));
 sg13g2_inv_1 _3424_ (.Y(_2774_),
    .A(_2773_));
 sg13g2_mux2_1 _3425_ (.A0(_2765_),
    .A1(_2772_),
    .S(_2774_),
    .X(_2775_));
 sg13g2_buf_2 _3426_ (.A(\g.g_y[0].g_x[4].t.out_sc ),
    .X(_2776_));
 sg13g2_buf_2 _3427_ (.A(\g.g_y[0].g_x[4].t.r_d ),
    .X(_2777_));
 sg13g2_mux2_1 _3428_ (.A0(_2776_),
    .A1(\g.g_y[0].g_x[4].t.r_gnl ),
    .S(_2777_),
    .X(_2778_));
 sg13g2_buf_1 _3429_ (.A(_2778_),
    .X(_2779_));
 sg13g2_buf_1 _3430_ (.A(\g.g_y[0].g_x[4].t.r_ghl ),
    .X(_2780_));
 sg13g2_buf_1 _3431_ (.A(\g.g_y[0].g_x[4].t.r_h ),
    .X(_2781_));
 sg13g2_mux2_1 _3432_ (.A0(_2779_),
    .A1(_2780_),
    .S(net174),
    .X(_2782_));
 sg13g2_nor2b_1 _3433_ (.A(_2624_),
    .B_N(_2623_),
    .Y(_2783_));
 sg13g2_a21o_1 _3434_ (.A2(_2622_),
    .A1(_2624_),
    .B1(_2783_),
    .X(_2784_));
 sg13g2_buf_2 _3435_ (.A(\g.g_y[0].g_x[3].t.r_h ),
    .X(_2785_));
 sg13g2_mux2_1 _3436_ (.A0(_2782_),
    .A1(_2784_),
    .S(_2785_),
    .X(_2786_));
 sg13g2_nand3_1 _3437_ (.B(_2775_),
    .C(_2786_),
    .A(_2758_),
    .Y(_2787_));
 sg13g2_buf_2 _3438_ (.A(\g.g_y[0].g_x[3].t.out_sc ),
    .X(_2788_));
 sg13g2_nor2_1 _3439_ (.A(_2788_),
    .B(_2758_),
    .Y(_2789_));
 sg13g2_nor2_1 _3440_ (.A(_2785_),
    .B(_2789_),
    .Y(_2790_));
 sg13g2_a21oi_1 _3441_ (.A1(_2759_),
    .A2(_2762_),
    .Y(_2791_),
    .B1(_2764_));
 sg13g2_nand2b_1 _3442_ (.Y(_2792_),
    .B(_2771_),
    .A_N(_2770_));
 sg13g2_o21ai_1 _3443_ (.B1(_2792_),
    .Y(_2793_),
    .A1(_2771_),
    .A2(_2769_));
 sg13g2_mux2_1 _3444_ (.A0(_2791_),
    .A1(_2793_),
    .S(_2773_),
    .X(_2794_));
 sg13g2_nand2_1 _3445_ (.Y(_2795_),
    .A(_2758_),
    .B(_2794_));
 sg13g2_o21ai_1 _3446_ (.B1(_2785_),
    .Y(_2796_),
    .A1(_2758_),
    .A2(_2782_));
 sg13g2_inv_1 _3447_ (.Y(_2797_),
    .A(_2796_));
 sg13g2_a22oi_1 _3448_ (.Y(_2798_),
    .B1(_2795_),
    .B2(_2797_),
    .A2(_2790_),
    .A1(_2787_));
 sg13g2_mux2_1 _3449_ (.A0(_2757_),
    .A1(_2798_),
    .S(_2624_),
    .X(_2799_));
 sg13g2_buf_2 _3450_ (.A(\g.g_y[6].g_x[2].t.r_v ),
    .X(_2800_));
 sg13g2_buf_2 _3451_ (.A(\g.g_y[6].g_x[2].t.out_sc ),
    .X(_2801_));
 sg13g2_buf_2 _3452_ (.A(\g.g_y[6].g_x[2].t.r_d ),
    .X(_2802_));
 sg13g2_mux2_1 _3453_ (.A0(\g.g_y[6].g_x[2].t.r_gnl ),
    .A1(_2801_),
    .S(_2802_),
    .X(_2803_));
 sg13g2_buf_1 _3454_ (.A(\g.g_y[6].g_x[2].t.r_ghl ),
    .X(_2804_));
 sg13g2_nor2b_1 _3455_ (.A(_2800_),
    .B_N(_2804_),
    .Y(_2805_));
 sg13g2_a21oi_1 _3456_ (.A1(_2800_),
    .A2(_2803_),
    .Y(_2806_),
    .B1(_2805_));
 sg13g2_buf_1 _3457_ (.A(\g.g_y[0].g_x[2].t.r_v ),
    .X(_2807_));
 sg13g2_mux2_1 _3458_ (.A0(\g.g_y[0].g_x[2].t.r_gnl ),
    .A1(_2620_),
    .S(_2621_),
    .X(_2808_));
 sg13g2_buf_1 _3459_ (.A(_2808_),
    .X(_2809_));
 sg13g2_nand2b_1 _3460_ (.Y(_2810_),
    .B(net173),
    .A_N(_2623_));
 sg13g2_o21ai_1 _3461_ (.B1(_2810_),
    .Y(_2811_),
    .A1(net173),
    .A2(_2809_));
 sg13g2_buf_2 _3462_ (.A(\g.g_y[7].g_x[2].t.r_v ),
    .X(_2812_));
 sg13g2_mux2_1 _3463_ (.A0(_2806_),
    .A1(_2811_),
    .S(_2812_),
    .X(_2813_));
 sg13g2_nor2b_1 _3464_ (.A(_2641_),
    .B_N(_2602_),
    .Y(_2814_));
 sg13g2_a21oi_1 _3465_ (.A1(_2641_),
    .A2(_2640_),
    .Y(_2815_),
    .B1(_2814_));
 sg13g2_buf_2 _3466_ (.A(\g.g_y[7].g_x[3].t.r_h ),
    .X(_2816_));
 sg13g2_mux2_1 _3467_ (.A0(_2760_),
    .A1(\g.g_y[7].g_x[3].t.r_gnl ),
    .S(_2761_),
    .X(_2817_));
 sg13g2_nand2b_1 _3468_ (.Y(_2818_),
    .B(_2816_),
    .A_N(_2763_));
 sg13g2_o21ai_1 _3469_ (.B1(_2818_),
    .Y(_2819_),
    .A1(_2816_),
    .A2(_2817_));
 sg13g2_buf_2 _3470_ (.A(\g.g_y[7].g_x[2].t.r_h ),
    .X(_2820_));
 sg13g2_mux2_1 _3471_ (.A0(_2815_),
    .A1(_2819_),
    .S(_2820_),
    .X(_2821_));
 sg13g2_buf_1 _3472_ (.A(\g.g_y[7].g_x[2].t.r_d ),
    .X(_2822_));
 sg13g2_inv_1 _3473_ (.Y(_2823_),
    .A(net172));
 sg13g2_mux2_1 _3474_ (.A0(_2813_),
    .A1(_2821_),
    .S(_2823_),
    .X(_2824_));
 sg13g2_mux2_1 _3475_ (.A0(_2811_),
    .A1(_2806_),
    .S(_2812_),
    .X(_2825_));
 sg13g2_mux2_1 _3476_ (.A0(_2817_),
    .A1(_2763_),
    .S(_2816_),
    .X(_2826_));
 sg13g2_nor2_1 _3477_ (.A(_2820_),
    .B(_2822_),
    .Y(_2827_));
 sg13g2_nor2b_1 _3478_ (.A(net172),
    .B_N(_2820_),
    .Y(_2828_));
 sg13g2_a21o_1 _3479_ (.A2(_2640_),
    .A1(_2641_),
    .B1(_2814_),
    .X(_2829_));
 sg13g2_a22oi_1 _3480_ (.Y(_2830_),
    .B1(_2828_),
    .B2(_2829_),
    .A2(_2827_),
    .A1(_2826_));
 sg13g2_buf_2 _3481_ (.A(\g.g_y[7].g_x[2].t.out_sc ),
    .X(_2831_));
 sg13g2_nand2b_1 _3482_ (.Y(_2832_),
    .B(net172),
    .A_N(_2831_));
 sg13g2_o21ai_1 _3483_ (.B1(_2832_),
    .Y(_2833_),
    .A1(_2825_),
    .A2(_2830_));
 sg13g2_mux2_1 _3484_ (.A0(_2824_),
    .A1(_2833_),
    .S(_2812_),
    .X(_2834_));
 sg13g2_buf_1 _3485_ (.A(\g.g_y[1].g_x[2].t.r_d ),
    .X(_2835_));
 sg13g2_nor2b_1 _3486_ (.A(net173),
    .B_N(_2623_),
    .Y(_2836_));
 sg13g2_a21o_1 _3487_ (.A2(_2809_),
    .A1(net173),
    .B1(_2836_),
    .X(_2837_));
 sg13g2_buf_2 _3488_ (.A(\g.g_y[2].g_x[2].t.out_sc ),
    .X(_2838_));
 sg13g2_buf_2 _3489_ (.A(\g.g_y[2].g_x[2].t.r_d ),
    .X(_2839_));
 sg13g2_mux2_1 _3490_ (.A0(\g.g_y[2].g_x[2].t.r_gnl ),
    .A1(_2838_),
    .S(_2839_),
    .X(_2840_));
 sg13g2_buf_1 _3491_ (.A(\g.g_y[2].g_x[2].t.r_ghl ),
    .X(_2841_));
 sg13g2_buf_2 _3492_ (.A(\g.g_y[2].g_x[2].t.r_v ),
    .X(_2842_));
 sg13g2_mux2_1 _3493_ (.A0(_2840_),
    .A1(_2841_),
    .S(_2842_),
    .X(_2843_));
 sg13g2_buf_1 _3494_ (.A(\g.g_y[1].g_x[2].t.r_v ),
    .X(_2844_));
 sg13g2_inv_1 _3495_ (.Y(_2845_),
    .A(_2844_));
 sg13g2_mux2_1 _3496_ (.A0(_2837_),
    .A1(_2843_),
    .S(_2845_),
    .X(_2846_));
 sg13g2_nor2b_1 _3497_ (.A(_2665_),
    .B_N(_2611_),
    .Y(_2847_));
 sg13g2_a21o_1 _3498_ (.A2(_2664_),
    .A1(_2665_),
    .B1(_2847_),
    .X(_2848_));
 sg13g2_mux2_1 _3499_ (.A0(_2766_),
    .A1(\g.g_y[1].g_x[3].t.r_gnl ),
    .S(_2767_),
    .X(_2849_));
 sg13g2_buf_2 _3500_ (.A(_2849_),
    .X(_2850_));
 sg13g2_inv_1 _3501_ (.Y(_2851_),
    .A(\g.g_y[1].g_x[3].t.r_h ));
 sg13g2_mux2_1 _3502_ (.A0(_2770_),
    .A1(_2850_),
    .S(_2851_),
    .X(_2852_));
 sg13g2_buf_2 _3503_ (.A(\g.g_y[1].g_x[2].t.r_h ),
    .X(_2853_));
 sg13g2_inv_1 _3504_ (.Y(_2854_),
    .A(_2853_));
 sg13g2_mux2_1 _3505_ (.A0(_2848_),
    .A1(_2852_),
    .S(_2854_),
    .X(_2855_));
 sg13g2_nand3b_1 _3506_ (.B(_2846_),
    .C(_2855_),
    .Y(_2856_),
    .A_N(_2835_));
 sg13g2_buf_1 _3507_ (.A(_2835_),
    .X(_2857_));
 sg13g2_buf_1 _3508_ (.A(\g.g_y[1].g_x[2].t.out_sc ),
    .X(_2858_));
 sg13g2_inv_1 _3509_ (.Y(_2859_),
    .A(_2858_));
 sg13g2_a21oi_1 _3510_ (.A1(_2857_),
    .A2(_2859_),
    .Y(_2860_),
    .B1(_2844_));
 sg13g2_a21oi_1 _3511_ (.A1(_2665_),
    .A2(_2664_),
    .Y(_2861_),
    .B1(_2847_));
 sg13g2_buf_1 _3512_ (.A(\g.g_y[1].g_x[3].t.r_h ),
    .X(_2862_));
 sg13g2_nand2b_1 _3513_ (.Y(_2863_),
    .B(net171),
    .A_N(_2770_));
 sg13g2_o21ai_1 _3514_ (.B1(_2863_),
    .Y(_2864_),
    .A1(_2862_),
    .A2(_2850_));
 sg13g2_mux2_1 _3515_ (.A0(_2861_),
    .A1(_2864_),
    .S(_2853_),
    .X(_2865_));
 sg13g2_nand2b_1 _3516_ (.Y(_2866_),
    .B(_2865_),
    .A_N(net122));
 sg13g2_nand2b_1 _3517_ (.Y(_2867_),
    .B(_2842_),
    .A_N(_2841_));
 sg13g2_o21ai_1 _3518_ (.B1(_2867_),
    .Y(_2868_),
    .A1(_2842_),
    .A2(_2840_));
 sg13g2_a21oi_1 _3519_ (.A1(net122),
    .A2(_2868_),
    .Y(_2869_),
    .B1(_2845_));
 sg13g2_a22oi_1 _3520_ (.Y(_2870_),
    .B1(_2866_),
    .B2(_2869_),
    .A2(_2860_),
    .A1(_2856_));
 sg13g2_mux2_1 _3521_ (.A0(_2834_),
    .A1(_2870_),
    .S(net173),
    .X(_2871_));
 sg13g2_mux2_1 _3522_ (.A0(_2799_),
    .A1(_2871_),
    .S(_2621_),
    .X(_2872_));
 sg13g2_buf_1 _3523_ (.A(_2753_),
    .X(_2873_));
 sg13g2_o21ai_1 _3524_ (.B1(net176),
    .Y(_2874_),
    .A1(_2623_),
    .A2(net59));
 sg13g2_a21oi_1 _3525_ (.A1(net60),
    .A2(_2872_),
    .Y(_0011_),
    .B1(_2874_));
 sg13g2_nand2b_1 _3526_ (.Y(_2875_),
    .B(_2807_),
    .A_N(_2834_));
 sg13g2_or2_1 _3527_ (.X(_2876_),
    .B(_2870_),
    .A(net173));
 sg13g2_nor2b_1 _3528_ (.A(_2624_),
    .B_N(_2798_),
    .Y(_2877_));
 sg13g2_a221oi_1 _3529_ (.B2(_2876_),
    .C1(_2877_),
    .B1(_2875_),
    .A1(_2624_),
    .Y(_2878_),
    .A2(_2757_));
 sg13g2_o21ai_1 _3530_ (.B1(_2696_),
    .Y(_2879_),
    .A1(\g.g_y[0].g_x[2].t.r_gnl ),
    .A2(net59));
 sg13g2_a21oi_1 _3531_ (.A1(net60),
    .A2(_2878_),
    .Y(_0012_),
    .B1(_2879_));
 sg13g2_nand2_1 _3532_ (.Y(_2880_),
    .A(_2620_),
    .B(_2702_));
 sg13g2_o21ai_1 _3533_ (.B1(_2624_),
    .Y(_2881_),
    .A1(net65),
    .A2(_2707_));
 sg13g2_a21oi_1 _3534_ (.A1(_2880_),
    .A2(_2881_),
    .Y(_0013_),
    .B1(_2711_));
 sg13g2_mux2_1 _3535_ (.A0(_2871_),
    .A1(_2799_),
    .S(_2621_),
    .X(_2882_));
 sg13g2_a22oi_1 _3536_ (.Y(_2883_),
    .B1(net62),
    .B2(_2630_),
    .A2(net63),
    .A1(_2620_));
 sg13g2_o21ai_1 _3537_ (.B1(_2883_),
    .Y(_0014_),
    .A1(_2716_),
    .A2(_2882_));
 sg13g2_nand2_1 _3538_ (.Y(_2884_),
    .A(_2620_),
    .B(_2729_));
 sg13g2_o21ai_1 _3539_ (.B1(_2807_),
    .Y(_2885_),
    .A1(_2705_),
    .A2(_2732_));
 sg13g2_a21oi_1 _3540_ (.A1(_2884_),
    .A2(_2885_),
    .Y(_0015_),
    .B1(_2711_));
 sg13g2_mux2_1 _3541_ (.A0(_2788_),
    .A1(_2758_),
    .S(_2593_),
    .X(_2886_));
 sg13g2_and2_1 _3542_ (.A(_2583_),
    .B(_2886_),
    .X(_0016_));
 sg13g2_nand2_1 _3543_ (.Y(_2887_),
    .A(_2788_),
    .B(net44));
 sg13g2_o21ai_1 _3544_ (.B1(_2785_),
    .Y(_2888_),
    .A1(net65),
    .A2(_2707_));
 sg13g2_buf_1 _3545_ (.A(_2737_),
    .X(_2889_));
 sg13g2_a21oi_1 _3546_ (.A1(_2887_),
    .A2(_2888_),
    .Y(_0017_),
    .B1(net93));
 sg13g2_buf_1 _3547_ (.A(net128),
    .X(_2890_));
 sg13g2_buf_1 _3548_ (.A(net175),
    .X(_2891_));
 sg13g2_nor2_1 _3549_ (.A(_2788_),
    .B(net121),
    .Y(_2892_));
 sg13g2_inv_1 _3550_ (.Y(_2893_),
    .A(net175));
 sg13g2_buf_1 _3551_ (.A(_2893_),
    .X(_2894_));
 sg13g2_buf_1 _3552_ (.A(net183),
    .X(_2895_));
 sg13g2_buf_1 _3553_ (.A(_2895_),
    .X(_2896_));
 sg13g2_a21oi_1 _3554_ (.A1(_2624_),
    .A2(_2622_),
    .Y(_2897_),
    .B1(_2783_));
 sg13g2_nand2b_1 _3555_ (.Y(_0320_),
    .B(net174),
    .A_N(_2780_));
 sg13g2_o21ai_1 _3556_ (.B1(_0320_),
    .Y(_0321_),
    .A1(net174),
    .A2(_2779_));
 sg13g2_mux2_1 _3557_ (.A0(_2897_),
    .A1(_0321_),
    .S(_2785_),
    .X(_0322_));
 sg13g2_mux2_1 _3558_ (.A0(_2794_),
    .A1(_0322_),
    .S(_2758_),
    .X(_0323_));
 sg13g2_buf_1 _3559_ (.A(net183),
    .X(_0324_));
 sg13g2_nand2_1 _3560_ (.Y(_0325_),
    .A(net169),
    .B(_2620_));
 sg13g2_o21ai_1 _3561_ (.B1(_0325_),
    .Y(_0326_),
    .A1(_2896_),
    .A2(_0323_));
 sg13g2_nor2_1 _3562_ (.A(net91),
    .B(_0326_),
    .Y(_0327_));
 sg13g2_nor3_1 _3563_ (.A(net92),
    .B(_2892_),
    .C(_0327_),
    .Y(_0018_));
 sg13g2_nand2_1 _3564_ (.Y(_0328_),
    .A(_2788_),
    .B(net43));
 sg13g2_o21ai_1 _3565_ (.B1(_2773_),
    .Y(_0329_),
    .A1(net65),
    .A2(net95));
 sg13g2_a21oi_1 _3566_ (.A1(_0328_),
    .A2(_0329_),
    .Y(_0019_),
    .B1(net93));
 sg13g2_mux2_1 _3567_ (.A0(_2776_),
    .A1(_2777_),
    .S(net47),
    .X(_0330_));
 sg13g2_and2_1 _3568_ (.A(net131),
    .B(_0330_),
    .X(_0020_));
 sg13g2_nor2b_1 _3569_ (.A(_2789_),
    .B_N(_2785_),
    .Y(_0331_));
 sg13g2_inv_1 _3570_ (.Y(_0332_),
    .A(_2758_));
 sg13g2_a21oi_1 _3571_ (.A1(_0332_),
    .A2(_2897_),
    .Y(_0333_),
    .B1(_2785_));
 sg13g2_a22oi_1 _3572_ (.Y(_0334_),
    .B1(_0333_),
    .B2(_2795_),
    .A2(_0331_),
    .A1(_2787_));
 sg13g2_buf_2 _3573_ (.A(\g.g_y[1].g_x[5].t.r_v ),
    .X(_0335_));
 sg13g2_buf_2 _3574_ (.A(\g.g_y[1].g_x[5].t.out_sc ),
    .X(_0336_));
 sg13g2_buf_8 _3575_ (.A(\g.g_y[1].g_x[5].t.r_d ),
    .X(_0337_));
 sg13g2_mux2_1 _3576_ (.A0(\g.g_y[1].g_x[5].t.r_gnl ),
    .A1(_0336_),
    .S(_0337_),
    .X(_0338_));
 sg13g2_buf_1 _3577_ (.A(_0338_),
    .X(_0339_));
 sg13g2_buf_1 _3578_ (.A(\g.g_y[1].g_x[5].t.r_ghl ),
    .X(_0340_));
 sg13g2_nand2b_1 _3579_ (.Y(_0341_),
    .B(_0335_),
    .A_N(_0340_));
 sg13g2_o21ai_1 _3580_ (.B1(_0341_),
    .Y(_0342_),
    .A1(_0335_),
    .A2(_0339_));
 sg13g2_buf_2 _3581_ (.A(\g.g_y[7].g_x[5].t.r_v ),
    .X(_0343_));
 sg13g2_inv_1 _3582_ (.Y(_0344_),
    .A(_0343_));
 sg13g2_buf_2 _3583_ (.A(\g.g_y[7].g_x[5].t.out_sc ),
    .X(_0345_));
 sg13g2_buf_2 _3584_ (.A(\g.g_y[7].g_x[5].t.r_d ),
    .X(_0346_));
 sg13g2_mux2_1 _3585_ (.A0(\g.g_y[7].g_x[5].t.r_gnl ),
    .A1(_0345_),
    .S(_0346_),
    .X(_0347_));
 sg13g2_buf_1 _3586_ (.A(_0347_),
    .X(_0348_));
 sg13g2_buf_1 _3587_ (.A(\g.g_y[7].g_x[5].t.r_ghl ),
    .X(_0349_));
 sg13g2_or2_1 _3588_ (.X(_0350_),
    .B(_0343_),
    .A(_0349_));
 sg13g2_o21ai_1 _3589_ (.B1(_0350_),
    .Y(_0351_),
    .A1(_0344_),
    .A2(_0348_));
 sg13g2_buf_2 _3590_ (.A(\g.g_y[0].g_x[5].t.r_v ),
    .X(_0352_));
 sg13g2_mux2_1 _3591_ (.A0(_0342_),
    .A1(_0351_),
    .S(_0352_),
    .X(_0353_));
 sg13g2_buf_2 _3592_ (.A(\g.g_y[0].g_x[6].t.out_sc ),
    .X(_0354_));
 sg13g2_buf_2 _3593_ (.A(\g.g_y[0].g_x[6].t.r_d ),
    .X(_0355_));
 sg13g2_mux2_1 _3594_ (.A0(_0354_),
    .A1(\g.g_y[0].g_x[6].t.r_gnl ),
    .S(_0355_),
    .X(_0356_));
 sg13g2_buf_1 _3595_ (.A(_0356_),
    .X(_0357_));
 sg13g2_buf_1 _3596_ (.A(\g.g_y[0].g_x[6].t.r_ghl ),
    .X(_0358_));
 sg13g2_buf_1 _3597_ (.A(\g.g_y[0].g_x[6].t.r_h ),
    .X(_0359_));
 sg13g2_mux2_1 _3598_ (.A0(_0357_),
    .A1(_0358_),
    .S(net168),
    .X(_0360_));
 sg13g2_buf_1 _3599_ (.A(\g.g_y[0].g_x[5].t.r_d ),
    .X(_0361_));
 sg13g2_nand3b_1 _3600_ (.B(_0360_),
    .C(net167),
    .Y(_0362_),
    .A_N(_0353_));
 sg13g2_buf_2 _3601_ (.A(\g.g_y[0].g_x[5].t.r_h ),
    .X(_0363_));
 sg13g2_buf_2 _3602_ (.A(\g.g_y[0].g_x[5].t.out_sc ),
    .X(_0364_));
 sg13g2_nor2_1 _3603_ (.A(_0364_),
    .B(net167),
    .Y(_0365_));
 sg13g2_nor2_1 _3604_ (.A(_0363_),
    .B(_0365_),
    .Y(_0366_));
 sg13g2_inv_1 _3605_ (.Y(_0367_),
    .A(\g.g_y[0].g_x[5].t.r_d ));
 sg13g2_nand2b_1 _3606_ (.Y(_0368_),
    .B(net168),
    .A_N(_0358_));
 sg13g2_o21ai_1 _3607_ (.B1(_0368_),
    .Y(_0369_),
    .A1(net168),
    .A2(_0357_));
 sg13g2_inv_1 _3608_ (.Y(_0370_),
    .A(_0335_));
 sg13g2_mux2_1 _3609_ (.A0(_0340_),
    .A1(_0339_),
    .S(_0370_),
    .X(_0371_));
 sg13g2_or2_1 _3610_ (.X(_0372_),
    .B(_0348_),
    .A(_0344_));
 sg13g2_nor2b_1 _3611_ (.A(_0352_),
    .B_N(_0350_),
    .Y(_0373_));
 sg13g2_a221oi_1 _3612_ (.B2(_0373_),
    .C1(_0367_),
    .B1(_0372_),
    .A1(_0352_),
    .Y(_0374_),
    .A2(_0371_));
 sg13g2_a21oi_1 _3613_ (.A1(_0367_),
    .A2(_0369_),
    .Y(_0375_),
    .B1(_0374_));
 sg13g2_a22oi_1 _3614_ (.Y(_0376_),
    .B1(_0375_),
    .B2(_0363_),
    .A2(_0366_),
    .A1(_0362_));
 sg13g2_mux2_1 _3615_ (.A0(_0334_),
    .A1(_0376_),
    .S(net174),
    .X(_0377_));
 sg13g2_buf_1 _3616_ (.A(\g.g_y[1].g_x[4].t.r_v ),
    .X(_0378_));
 sg13g2_buf_1 _3617_ (.A(\g.g_y[1].g_x[4].t.r_d ),
    .X(_0379_));
 sg13g2_buf_1 _3618_ (.A(\g.g_y[1].g_x[4].t.out_sc ),
    .X(_0380_));
 sg13g2_inv_1 _3619_ (.Y(_0381_),
    .A(_0380_));
 sg13g2_nand2_1 _3620_ (.Y(_0382_),
    .A(_0379_),
    .B(_0381_));
 sg13g2_buf_2 _3621_ (.A(\g.g_y[0].g_x[4].t.r_v ),
    .X(_0383_));
 sg13g2_o21ai_1 _3622_ (.B1(_0383_),
    .Y(_0384_),
    .A1(_0378_),
    .A2(_0382_));
 sg13g2_buf_1 _3623_ (.A(\g.g_y[7].g_x[4].t.r_v ),
    .X(_0385_));
 sg13g2_buf_1 _3624_ (.A(\g.g_y[7].g_x[4].t.r_d ),
    .X(_0386_));
 sg13g2_buf_1 _3625_ (.A(_0386_),
    .X(_0387_));
 sg13g2_mux2_1 _3626_ (.A0(_0345_),
    .A1(\g.g_y[7].g_x[5].t.r_gnl ),
    .S(_0346_),
    .X(_0388_));
 sg13g2_buf_2 _3627_ (.A(\g.g_y[7].g_x[5].t.r_h ),
    .X(_0389_));
 sg13g2_mux2_1 _3628_ (.A0(_0388_),
    .A1(_0349_),
    .S(_0389_),
    .X(_0390_));
 sg13g2_buf_2 _3629_ (.A(_0390_),
    .X(_0391_));
 sg13g2_mux2_1 _3630_ (.A0(_2763_),
    .A1(_2817_),
    .S(_2816_),
    .X(_0392_));
 sg13g2_buf_1 _3631_ (.A(\g.g_y[7].g_x[4].t.r_h ),
    .X(_0393_));
 sg13g2_inv_1 _3632_ (.Y(_0394_),
    .A(_0393_));
 sg13g2_mux2_1 _3633_ (.A0(_0391_),
    .A1(_0392_),
    .S(_0394_),
    .X(_0395_));
 sg13g2_buf_1 _3634_ (.A(_0395_),
    .X(_0396_));
 sg13g2_or3_1 _3635_ (.A(net166),
    .B(net119),
    .C(_0396_),
    .X(_0397_));
 sg13g2_buf_2 _3636_ (.A(\g.g_y[7].g_x[4].t.out_sc ),
    .X(_0398_));
 sg13g2_nor2b_1 _3637_ (.A(_0398_),
    .B_N(_0386_),
    .Y(_0399_));
 sg13g2_a21oi_1 _3638_ (.A1(net166),
    .A2(_0399_),
    .Y(_0400_),
    .B1(_0383_));
 sg13g2_mux2_1 _3639_ (.A0(_0391_),
    .A1(_0392_),
    .S(_0393_),
    .X(_0401_));
 sg13g2_buf_1 _3640_ (.A(_0401_),
    .X(_0402_));
 sg13g2_buf_2 _3641_ (.A(\g.g_y[6].g_x[4].t.r_v ),
    .X(_0403_));
 sg13g2_buf_2 _3642_ (.A(\g.g_y[6].g_x[4].t.out_sc ),
    .X(_0404_));
 sg13g2_buf_8 _3643_ (.A(\g.g_y[6].g_x[4].t.r_d ),
    .X(_0405_));
 sg13g2_mux2_1 _3644_ (.A0(\g.g_y[6].g_x[4].t.r_gnl ),
    .A1(_0404_),
    .S(_0405_),
    .X(_0406_));
 sg13g2_buf_2 _3645_ (.A(\g.g_y[6].g_x[4].t.r_ghl ),
    .X(_0407_));
 sg13g2_nor2b_1 _3646_ (.A(_0403_),
    .B_N(_0407_),
    .Y(_0408_));
 sg13g2_a21oi_1 _3647_ (.A1(_0403_),
    .A2(_0406_),
    .Y(_0409_),
    .B1(_0408_));
 sg13g2_nor2_1 _3648_ (.A(_0386_),
    .B(_0409_),
    .Y(_0410_));
 sg13g2_nand3_1 _3649_ (.B(_0402_),
    .C(_0410_),
    .A(_0385_),
    .Y(_0411_));
 sg13g2_inv_1 _3650_ (.Y(_0412_),
    .A(net166));
 sg13g2_nand3_1 _3651_ (.B(net119),
    .C(_0409_),
    .A(_0412_),
    .Y(_0413_));
 sg13g2_nand4_1 _3652_ (.B(_0400_),
    .C(_0411_),
    .A(_0397_),
    .Y(_0414_),
    .D(_0413_));
 sg13g2_inv_1 _3653_ (.Y(_0415_),
    .A(_0378_));
 sg13g2_inv_1 _3654_ (.Y(_0416_),
    .A(_0379_));
 sg13g2_nor2b_1 _3655_ (.A(\g.g_y[1].g_x[3].t.r_h ),
    .B_N(_2770_),
    .Y(_0417_));
 sg13g2_a21o_1 _3656_ (.A2(_2850_),
    .A1(net171),
    .B1(_0417_),
    .X(_0418_));
 sg13g2_mux2_1 _3657_ (.A0(_0336_),
    .A1(\g.g_y[1].g_x[5].t.r_gnl ),
    .S(_0337_),
    .X(_0419_));
 sg13g2_buf_2 _3658_ (.A(\g.g_y[1].g_x[5].t.r_h ),
    .X(_0420_));
 sg13g2_mux2_1 _3659_ (.A0(_0419_),
    .A1(_0340_),
    .S(_0420_),
    .X(_0421_));
 sg13g2_buf_2 _3660_ (.A(_0421_),
    .X(_0422_));
 sg13g2_buf_2 _3661_ (.A(\g.g_y[1].g_x[4].t.r_h ),
    .X(_0423_));
 sg13g2_inv_2 _3662_ (.Y(_0424_),
    .A(_0423_));
 sg13g2_mux2_1 _3663_ (.A0(_0418_),
    .A1(_0422_),
    .S(_0424_),
    .X(_0425_));
 sg13g2_mux2_1 _3664_ (.A0(\g.g_y[0].g_x[4].t.r_gnl ),
    .A1(_2776_),
    .S(_2777_),
    .X(_0426_));
 sg13g2_nor2b_1 _3665_ (.A(_0383_),
    .B_N(_2780_),
    .Y(_0427_));
 sg13g2_a21o_1 _3666_ (.A2(_0426_),
    .A1(_0383_),
    .B1(_0427_),
    .X(_0428_));
 sg13g2_buf_2 _3667_ (.A(\g.g_y[2].g_x[4].t.r_ghl ),
    .X(_0429_));
 sg13g2_buf_2 _3668_ (.A(\g.g_y[2].g_x[4].t.out_sc ),
    .X(_0430_));
 sg13g2_buf_2 _3669_ (.A(\g.g_y[2].g_x[4].t.r_d ),
    .X(_0431_));
 sg13g2_mux2_1 _3670_ (.A0(\g.g_y[2].g_x[4].t.r_gnl ),
    .A1(_0430_),
    .S(_0431_),
    .X(_0432_));
 sg13g2_buf_1 _3671_ (.A(_0432_),
    .X(_0433_));
 sg13g2_buf_2 _3672_ (.A(\g.g_y[2].g_x[4].t.r_v ),
    .X(_0434_));
 sg13g2_inv_2 _3673_ (.Y(_0435_),
    .A(_0434_));
 sg13g2_mux2_1 _3674_ (.A0(_0429_),
    .A1(_0433_),
    .S(_0435_),
    .X(_0436_));
 sg13g2_mux2_1 _3675_ (.A0(_0428_),
    .A1(_0436_),
    .S(_0415_),
    .X(_0437_));
 sg13g2_nand3_1 _3676_ (.B(_0425_),
    .C(_0437_),
    .A(_0416_),
    .Y(_0438_));
 sg13g2_buf_1 _3677_ (.A(_0379_),
    .X(_0439_));
 sg13g2_a21oi_1 _3678_ (.A1(_0383_),
    .A2(_0426_),
    .Y(_0440_),
    .B1(_0427_));
 sg13g2_nand2b_1 _3679_ (.Y(_0441_),
    .B(_0434_),
    .A_N(_0429_));
 sg13g2_o21ai_1 _3680_ (.B1(_0441_),
    .Y(_0442_),
    .A1(_0434_),
    .A2(_0433_));
 sg13g2_mux2_1 _3681_ (.A0(_0440_),
    .A1(_0442_),
    .S(_0378_),
    .X(_0443_));
 sg13g2_buf_1 _3682_ (.A(_0443_),
    .X(_0444_));
 sg13g2_nand2_1 _3683_ (.Y(_0445_),
    .A(net118),
    .B(_0444_));
 sg13g2_inv_1 _3684_ (.Y(_0446_),
    .A(_2770_));
 sg13g2_a21oi_1 _3685_ (.A1(_0446_),
    .A2(_2851_),
    .Y(_0447_),
    .B1(_0423_));
 sg13g2_or2_1 _3686_ (.X(_0448_),
    .B(_2850_),
    .A(_2851_));
 sg13g2_a221oi_1 _3687_ (.B2(_0448_),
    .C1(_0379_),
    .B1(_0447_),
    .A1(_0423_),
    .Y(_0449_),
    .A2(_0422_));
 sg13g2_nor2_1 _3688_ (.A(_0415_),
    .B(_0449_),
    .Y(_0450_));
 sg13g2_inv_1 _3689_ (.Y(_0451_),
    .A(_0383_));
 sg13g2_a221oi_1 _3690_ (.B2(_0450_),
    .C1(_0451_),
    .B1(_0445_),
    .A1(_0415_),
    .Y(_0452_),
    .A2(_0438_));
 sg13g2_a21o_1 _3691_ (.A2(_0414_),
    .A1(_0384_),
    .B1(_0452_),
    .X(_0453_));
 sg13g2_mux2_1 _3692_ (.A0(_0377_),
    .A1(_0453_),
    .S(_2777_),
    .X(_0454_));
 sg13g2_o21ai_1 _3693_ (.B1(_2696_),
    .Y(_0455_),
    .A1(_2780_),
    .A2(net45));
 sg13g2_a21oi_1 _3694_ (.A1(net46),
    .A2(_0454_),
    .Y(_0021_),
    .B1(_0455_));
 sg13g2_nand2_1 _3695_ (.Y(_0456_),
    .A(net182),
    .B(_2596_));
 sg13g2_buf_2 _3696_ (.A(_0456_),
    .X(_0457_));
 sg13g2_mux2_1 _3697_ (.A0(_0376_),
    .A1(_0334_),
    .S(net174),
    .X(_0458_));
 sg13g2_a21oi_1 _3698_ (.A1(_0402_),
    .A2(_0410_),
    .Y(_0459_),
    .B1(_0399_));
 sg13g2_a21oi_1 _3699_ (.A1(net119),
    .A2(_0409_),
    .Y(_0460_),
    .B1(net166));
 sg13g2_or2_1 _3700_ (.X(_0461_),
    .B(_0396_),
    .A(net119));
 sg13g2_a221oi_1 _3701_ (.B2(_0461_),
    .C1(_0451_),
    .B1(_0460_),
    .A1(net166),
    .Y(_0462_),
    .A2(_0459_));
 sg13g2_and2_1 _3702_ (.A(_0415_),
    .B(_0438_),
    .X(_0463_));
 sg13g2_a221oi_1 _3703_ (.B2(_0450_),
    .C1(_0383_),
    .B1(_0445_),
    .A1(_0382_),
    .Y(_0464_),
    .A2(_0463_));
 sg13g2_nor4_1 _3704_ (.A(_0457_),
    .B(_0458_),
    .C(_0462_),
    .D(_0464_),
    .Y(_0465_));
 sg13g2_buf_1 _3705_ (.A(net181),
    .X(_0466_));
 sg13g2_o21ai_1 _3706_ (.B1(_0466_),
    .Y(_0467_),
    .A1(\g.g_y[0].g_x[4].t.r_gnl ),
    .A2(_2689_));
 sg13g2_nor2_1 _3707_ (.A(_0465_),
    .B(_0467_),
    .Y(_0022_));
 sg13g2_nand2_1 _3708_ (.Y(_0468_),
    .A(_2776_),
    .B(net44));
 sg13g2_o21ai_1 _3709_ (.B1(_2781_),
    .Y(_0469_),
    .A1(net65),
    .A2(net98));
 sg13g2_a21oi_1 _3710_ (.A1(_0468_),
    .A2(_0469_),
    .Y(_0023_),
    .B1(net93));
 sg13g2_mux2_1 _3711_ (.A0(_0453_),
    .A1(_0377_),
    .S(_2777_),
    .X(_0470_));
 sg13g2_a22oi_1 _3712_ (.Y(_0471_),
    .B1(_2723_),
    .B2(_2788_),
    .A2(_2720_),
    .A1(_2776_));
 sg13g2_o21ai_1 _3713_ (.B1(_0471_),
    .Y(_0024_),
    .A1(_2716_),
    .A2(_0470_));
 sg13g2_nand2_1 _3714_ (.Y(_0472_),
    .A(_2776_),
    .B(net43));
 sg13g2_o21ai_1 _3715_ (.B1(_0383_),
    .Y(_0473_),
    .A1(net65),
    .A2(net95));
 sg13g2_a21oi_1 _3716_ (.A1(_0472_),
    .A2(_0473_),
    .Y(_0025_),
    .B1(net93));
 sg13g2_mux2_1 _3717_ (.A0(_0364_),
    .A1(net167),
    .S(net47),
    .X(_0474_));
 sg13g2_and2_1 _3718_ (.A(net131),
    .B(_0474_),
    .X(_0026_));
 sg13g2_nand2_1 _3719_ (.Y(_0475_),
    .A(_0364_),
    .B(net44));
 sg13g2_buf_1 _3720_ (.A(net99),
    .X(_0476_));
 sg13g2_o21ai_1 _3721_ (.B1(_0363_),
    .Y(_0477_),
    .A1(net58),
    .A2(net98));
 sg13g2_a21oi_1 _3722_ (.A1(_0475_),
    .A2(_0477_),
    .Y(_0027_),
    .B1(net93));
 sg13g2_nor2_1 _3723_ (.A(_0364_),
    .B(net121),
    .Y(_0478_));
 sg13g2_nor2b_1 _3724_ (.A(net174),
    .B_N(_2780_),
    .Y(_0479_));
 sg13g2_a21oi_1 _3725_ (.A1(net174),
    .A2(_2779_),
    .Y(_0480_),
    .B1(_0479_));
 sg13g2_mux2_1 _3726_ (.A0(_0480_),
    .A1(_0369_),
    .S(_0363_),
    .X(_0481_));
 sg13g2_a221oi_1 _3727_ (.B2(_0373_),
    .C1(net167),
    .B1(_0372_),
    .A1(_0352_),
    .Y(_0482_),
    .A2(_0371_));
 sg13g2_a21oi_1 _3728_ (.A1(net167),
    .A2(_0481_),
    .Y(_0483_),
    .B1(_0482_));
 sg13g2_mux2_1 _3729_ (.A0(_2776_),
    .A1(_0483_),
    .S(net124),
    .X(_0484_));
 sg13g2_nor2_1 _3730_ (.A(net91),
    .B(_0484_),
    .Y(_0485_));
 sg13g2_nor3_1 _3731_ (.A(net92),
    .B(_0478_),
    .C(_0485_),
    .Y(_0028_));
 sg13g2_nand2_1 _3732_ (.Y(_0486_),
    .A(_0364_),
    .B(net43));
 sg13g2_o21ai_1 _3733_ (.B1(_0352_),
    .Y(_0487_),
    .A1(net58),
    .A2(net95));
 sg13g2_a21oi_1 _3734_ (.A1(_0486_),
    .A2(_0487_),
    .Y(_0029_),
    .B1(net93));
 sg13g2_mux2_1 _3735_ (.A0(_0354_),
    .A1(_0355_),
    .S(net47),
    .X(_0488_));
 sg13g2_and2_1 _3736_ (.A(net131),
    .B(_0488_),
    .X(_0030_));
 sg13g2_a21o_1 _3737_ (.A2(_2779_),
    .A1(net174),
    .B1(_0479_),
    .X(_0489_));
 sg13g2_nand3b_1 _3738_ (.B(_0489_),
    .C(_0361_),
    .Y(_0490_),
    .A_N(_0353_));
 sg13g2_nor2b_1 _3739_ (.A(_0365_),
    .B_N(_0363_),
    .Y(_0491_));
 sg13g2_nor2_1 _3740_ (.A(net167),
    .B(_0489_),
    .Y(_0492_));
 sg13g2_nor3_1 _3741_ (.A(_0363_),
    .B(_0374_),
    .C(_0492_),
    .Y(_0493_));
 sg13g2_a21oi_1 _3742_ (.A1(_0490_),
    .A2(_0491_),
    .Y(_0494_),
    .B1(_0493_));
 sg13g2_buf_1 _3743_ (.A(\g.g_y[0].g_x[7].t.out_sc ),
    .X(_0495_));
 sg13g2_inv_1 _3744_ (.Y(_0496_),
    .A(_0495_));
 sg13g2_nand2b_1 _3745_ (.Y(_0497_),
    .B(net180),
    .A_N(_2617_));
 sg13g2_o21ai_1 _3746_ (.B1(_0497_),
    .Y(_0498_),
    .A1(net180),
    .A2(_2618_));
 sg13g2_mux2_1 _3747_ (.A0(_2618_),
    .A1(_2617_),
    .S(net180),
    .X(_0499_));
 sg13g2_nor2b_1 _3748_ (.A(net168),
    .B_N(_0358_),
    .Y(_0500_));
 sg13g2_a21o_1 _3749_ (.A2(_0357_),
    .A1(net168),
    .B1(_0500_),
    .X(_0501_));
 sg13g2_buf_2 _3750_ (.A(\g.g_y[0].g_x[7].t.r_h ),
    .X(_0502_));
 sg13g2_mux2_1 _3751_ (.A0(_0499_),
    .A1(_0501_),
    .S(_0502_),
    .X(_0503_));
 sg13g2_buf_2 _3752_ (.A(\g.g_y[1].g_x[7].t.out_sc ),
    .X(_0504_));
 sg13g2_buf_2 _3753_ (.A(\g.g_y[1].g_x[7].t.r_d ),
    .X(_0505_));
 sg13g2_mux2_1 _3754_ (.A0(\g.g_y[1].g_x[7].t.r_gnl ),
    .A1(_0504_),
    .S(_0505_),
    .X(_0506_));
 sg13g2_buf_1 _3755_ (.A(_0506_),
    .X(_0507_));
 sg13g2_buf_1 _3756_ (.A(\g.g_y[1].g_x[7].t.r_ghl ),
    .X(_0508_));
 sg13g2_buf_1 _3757_ (.A(\g.g_y[1].g_x[7].t.r_v ),
    .X(_0509_));
 sg13g2_mux2_1 _3758_ (.A0(_0507_),
    .A1(_0508_),
    .S(net165),
    .X(_0510_));
 sg13g2_buf_2 _3759_ (.A(\g.g_y[7].g_x[7].t.r_v ),
    .X(_0511_));
 sg13g2_buf_1 _3760_ (.A(\g.g_y[7].g_x[7].t.out_sc ),
    .X(_0512_));
 sg13g2_buf_8 _3761_ (.A(\g.g_y[7].g_x[7].t.r_d ),
    .X(_0513_));
 sg13g2_mux2_1 _3762_ (.A0(\g.g_y[7].g_x[7].t.r_gnl ),
    .A1(_0512_),
    .S(_0513_),
    .X(_0514_));
 sg13g2_buf_1 _3763_ (.A(\g.g_y[7].g_x[7].t.r_ghl ),
    .X(_0515_));
 sg13g2_nor2b_1 _3764_ (.A(_0511_),
    .B_N(_0515_),
    .Y(_0516_));
 sg13g2_a21o_1 _3765_ (.A2(_0514_),
    .A1(_0511_),
    .B1(_0516_),
    .X(_0517_));
 sg13g2_buf_1 _3766_ (.A(\g.g_y[0].g_x[7].t.r_v ),
    .X(_0518_));
 sg13g2_mux2_1 _3767_ (.A0(_0510_),
    .A1(_0517_),
    .S(_0518_),
    .X(_0519_));
 sg13g2_and2_1 _3768_ (.A(_0503_),
    .B(_0519_),
    .X(_0520_));
 sg13g2_nand2_1 _3769_ (.Y(_0521_),
    .A(_0518_),
    .B(_0510_));
 sg13g2_inv_1 _3770_ (.Y(_0522_),
    .A(_0518_));
 sg13g2_nand2_1 _3771_ (.Y(_0523_),
    .A(_0522_),
    .B(_0517_));
 sg13g2_and2_1 _3772_ (.A(_0521_),
    .B(_0523_),
    .X(_0524_));
 sg13g2_buf_2 _3773_ (.A(\g.g_y[0].g_x[7].t.r_d ),
    .X(_0525_));
 sg13g2_mux4_1 _3774_ (.S0(_0502_),
    .A0(_0496_),
    .A1(_0498_),
    .A2(_0520_),
    .A3(_0524_),
    .S1(_0525_),
    .X(_0526_));
 sg13g2_mux2_1 _3775_ (.A0(_0494_),
    .A1(_0526_),
    .S(net168),
    .X(_0527_));
 sg13g2_buf_1 _3776_ (.A(\g.g_y[7].g_x[6].t.r_d ),
    .X(_0528_));
 sg13g2_buf_1 _3777_ (.A(\g.g_y[0].g_x[6].t.r_v ),
    .X(_0529_));
 sg13g2_mux2_1 _3778_ (.A0(\g.g_y[0].g_x[6].t.r_gnl ),
    .A1(_0354_),
    .S(_0355_),
    .X(_0530_));
 sg13g2_buf_1 _3779_ (.A(_0530_),
    .X(_0531_));
 sg13g2_nand2b_1 _3780_ (.Y(_0532_),
    .B(net163),
    .A_N(_0358_));
 sg13g2_o21ai_1 _3781_ (.B1(_0532_),
    .Y(_0533_),
    .A1(net163),
    .A2(_0531_));
 sg13g2_buf_2 _3782_ (.A(\g.g_y[6].g_x[6].t.r_v ),
    .X(_0534_));
 sg13g2_inv_1 _3783_ (.Y(_0535_),
    .A(_0534_));
 sg13g2_buf_2 _3784_ (.A(\g.g_y[6].g_x[6].t.out_sc ),
    .X(_0536_));
 sg13g2_buf_8 _3785_ (.A(\g.g_y[6].g_x[6].t.r_d ),
    .X(_0537_));
 sg13g2_mux2_1 _3786_ (.A0(\g.g_y[6].g_x[6].t.r_gnl ),
    .A1(_0536_),
    .S(_0537_),
    .X(_0538_));
 sg13g2_buf_1 _3787_ (.A(\g.g_y[6].g_x[6].t.r_ghl ),
    .X(_0539_));
 sg13g2_or2_1 _3788_ (.X(_0540_),
    .B(_0534_),
    .A(_0539_));
 sg13g2_o21ai_1 _3789_ (.B1(_0540_),
    .Y(_0541_),
    .A1(_0535_),
    .A2(_0538_));
 sg13g2_buf_1 _3790_ (.A(\g.g_y[7].g_x[6].t.r_v ),
    .X(_0542_));
 sg13g2_mux2_1 _3791_ (.A0(_0533_),
    .A1(_0541_),
    .S(net162),
    .X(_0543_));
 sg13g2_buf_2 _3792_ (.A(\g.g_y[7].g_x[7].t.r_h ),
    .X(_0544_));
 sg13g2_mux2_1 _3793_ (.A0(_0512_),
    .A1(\g.g_y[7].g_x[7].t.r_gnl ),
    .S(_0513_),
    .X(_0545_));
 sg13g2_nand2b_1 _3794_ (.Y(_0546_),
    .B(_0544_),
    .A_N(_0515_));
 sg13g2_o21ai_1 _3795_ (.B1(_0546_),
    .Y(_0547_),
    .A1(_0544_),
    .A2(_0545_));
 sg13g2_nor2b_1 _3796_ (.A(_0389_),
    .B_N(_0349_),
    .Y(_0548_));
 sg13g2_a21oi_1 _3797_ (.A1(_0389_),
    .A2(_0388_),
    .Y(_0549_),
    .B1(_0548_));
 sg13g2_buf_2 _3798_ (.A(\g.g_y[7].g_x[6].t.r_h ),
    .X(_0550_));
 sg13g2_mux2_1 _3799_ (.A0(_0547_),
    .A1(_0549_),
    .S(_0550_),
    .X(_0551_));
 sg13g2_or3_1 _3800_ (.A(net164),
    .B(_0543_),
    .C(_0551_),
    .X(_0552_));
 sg13g2_buf_2 _3801_ (.A(\g.g_y[7].g_x[6].t.out_sc ),
    .X(_0553_));
 sg13g2_nand2b_1 _3802_ (.Y(_0554_),
    .B(net164),
    .A_N(_0553_));
 sg13g2_and2_1 _3803_ (.A(net162),
    .B(_0554_),
    .X(_0555_));
 sg13g2_inv_1 _3804_ (.Y(_0556_),
    .A(net164));
 sg13g2_mux2_1 _3805_ (.A0(_0549_),
    .A1(_0547_),
    .S(_0550_),
    .X(_0557_));
 sg13g2_mux2_1 _3806_ (.A0(_0531_),
    .A1(_0358_),
    .S(net163),
    .X(_0558_));
 sg13g2_or2_1 _3807_ (.X(_0559_),
    .B(_0538_),
    .A(_0535_));
 sg13g2_inv_1 _3808_ (.Y(_0560_),
    .A(net162));
 sg13g2_and2_1 _3809_ (.A(_0560_),
    .B(_0540_),
    .X(_0561_));
 sg13g2_a221oi_1 _3810_ (.B2(_0561_),
    .C1(_0556_),
    .B1(_0559_),
    .A1(net162),
    .Y(_0562_),
    .A2(_0558_));
 sg13g2_a21oi_1 _3811_ (.A1(_0556_),
    .A2(_0557_),
    .Y(_0563_),
    .B1(_0562_));
 sg13g2_a22oi_1 _3812_ (.Y(_0564_),
    .B1(_0563_),
    .B2(_0560_),
    .A2(_0555_),
    .A1(_0552_));
 sg13g2_mux2_1 _3813_ (.A0(_0504_),
    .A1(\g.g_y[1].g_x[7].t.r_gnl ),
    .S(_0505_),
    .X(_0565_));
 sg13g2_buf_2 _3814_ (.A(\g.g_y[1].g_x[7].t.r_h ),
    .X(_0566_));
 sg13g2_mux2_1 _3815_ (.A0(_0565_),
    .A1(_0508_),
    .S(_0566_),
    .X(_0567_));
 sg13g2_nor2b_1 _3816_ (.A(_0420_),
    .B_N(_0340_),
    .Y(_0568_));
 sg13g2_a21o_1 _3817_ (.A2(_0419_),
    .A1(_0420_),
    .B1(_0568_),
    .X(_0569_));
 sg13g2_buf_2 _3818_ (.A(\g.g_y[1].g_x[6].t.r_h ),
    .X(_0570_));
 sg13g2_mux2_1 _3819_ (.A0(_0567_),
    .A1(_0569_),
    .S(_0570_),
    .X(_0571_));
 sg13g2_buf_2 _3820_ (.A(\g.g_y[2].g_x[6].t.out_sc ),
    .X(_0572_));
 sg13g2_buf_2 _3821_ (.A(\g.g_y[2].g_x[6].t.r_d ),
    .X(_0573_));
 sg13g2_mux2_1 _3822_ (.A0(\g.g_y[2].g_x[6].t.r_gnl ),
    .A1(_0572_),
    .S(_0573_),
    .X(_0574_));
 sg13g2_buf_1 _3823_ (.A(\g.g_y[2].g_x[6].t.r_ghl ),
    .X(_0575_));
 sg13g2_buf_2 _3824_ (.A(\g.g_y[2].g_x[6].t.r_v ),
    .X(_0576_));
 sg13g2_mux2_1 _3825_ (.A0(_0574_),
    .A1(_0575_),
    .S(_0576_),
    .X(_0577_));
 sg13g2_nor2b_1 _3826_ (.A(net163),
    .B_N(_0358_),
    .Y(_0578_));
 sg13g2_a21o_1 _3827_ (.A2(_0531_),
    .A1(net163),
    .B1(_0578_),
    .X(_0579_));
 sg13g2_buf_2 _3828_ (.A(\g.g_y[1].g_x[6].t.r_v ),
    .X(_0580_));
 sg13g2_mux2_1 _3829_ (.A0(_0577_),
    .A1(_0579_),
    .S(_0580_),
    .X(_0581_));
 sg13g2_and2_1 _3830_ (.A(_0571_),
    .B(_0581_),
    .X(_0582_));
 sg13g2_a21oi_1 _3831_ (.A1(_0420_),
    .A2(_0419_),
    .Y(_0583_),
    .B1(_0568_));
 sg13g2_nand2b_1 _3832_ (.Y(_0584_),
    .B(_0566_),
    .A_N(_0508_));
 sg13g2_o21ai_1 _3833_ (.B1(_0584_),
    .Y(_0585_),
    .A1(_0566_),
    .A2(_0565_));
 sg13g2_mux2_1 _3834_ (.A0(_0583_),
    .A1(_0585_),
    .S(_0570_),
    .X(_0586_));
 sg13g2_buf_1 _3835_ (.A(\g.g_y[1].g_x[6].t.out_sc ),
    .X(_0587_));
 sg13g2_inv_1 _3836_ (.Y(_0588_),
    .A(_0587_));
 sg13g2_inv_1 _3837_ (.Y(_0589_),
    .A(_0577_));
 sg13g2_buf_2 _3838_ (.A(\g.g_y[1].g_x[6].t.r_d ),
    .X(_0590_));
 sg13g2_mux4_1 _3839_ (.S0(_0580_),
    .A0(_0582_),
    .A1(_0586_),
    .A2(_0588_),
    .A3(_0589_),
    .S1(_0590_),
    .X(_0591_));
 sg13g2_mux2_1 _3840_ (.A0(_0564_),
    .A1(_0591_),
    .S(net163),
    .X(_0592_));
 sg13g2_mux2_1 _3841_ (.A0(_0527_),
    .A1(_0592_),
    .S(_0355_),
    .X(_0593_));
 sg13g2_o21ai_1 _3842_ (.B1(net176),
    .Y(_0594_),
    .A1(_0358_),
    .A2(net59));
 sg13g2_a21oi_1 _3843_ (.A1(net60),
    .A2(_0593_),
    .Y(_0031_),
    .B1(_0594_));
 sg13g2_nand2_1 _3844_ (.Y(_0595_),
    .A(net182),
    .B(_2751_));
 sg13g2_buf_2 _3845_ (.A(_0595_),
    .X(_0596_));
 sg13g2_mux2_1 _3846_ (.A0(_0526_),
    .A1(_0494_),
    .S(net168),
    .X(_0597_));
 sg13g2_mux2_1 _3847_ (.A0(_0591_),
    .A1(_0564_),
    .S(net163),
    .X(_0598_));
 sg13g2_nor3_1 _3848_ (.A(_0596_),
    .B(_0597_),
    .C(_0598_),
    .Y(_0599_));
 sg13g2_o21ai_1 _3849_ (.B1(net117),
    .Y(_0600_),
    .A1(\g.g_y[0].g_x[6].t.r_gnl ),
    .A2(net59));
 sg13g2_nor2_1 _3850_ (.A(_0599_),
    .B(_0600_),
    .Y(_0032_));
 sg13g2_nand2_1 _3851_ (.Y(_0601_),
    .A(_0354_),
    .B(net44));
 sg13g2_o21ai_1 _3852_ (.B1(_0359_),
    .Y(_0602_),
    .A1(net58),
    .A2(net98));
 sg13g2_a21oi_1 _3853_ (.A1(_0601_),
    .A2(_0602_),
    .Y(_0033_),
    .B1(_2889_));
 sg13g2_mux2_1 _3854_ (.A0(_0592_),
    .A1(_0527_),
    .S(_0355_),
    .X(_0603_));
 sg13g2_a22oi_1 _3855_ (.Y(_0604_),
    .B1(net62),
    .B2(_0364_),
    .A2(net63),
    .A1(_0354_));
 sg13g2_o21ai_1 _3856_ (.B1(_0604_),
    .Y(_0034_),
    .A1(net64),
    .A2(_0603_));
 sg13g2_nand2_1 _3857_ (.Y(_0605_),
    .A(_0354_),
    .B(net43));
 sg13g2_o21ai_1 _3858_ (.B1(_0529_),
    .Y(_0606_),
    .A1(_0476_),
    .A2(net95));
 sg13g2_a21oi_1 _3859_ (.A1(_0605_),
    .A2(_0606_),
    .Y(_0035_),
    .B1(_2889_));
 sg13g2_buf_1 _3860_ (.A(_2592_),
    .X(_0607_));
 sg13g2_buf_1 _3861_ (.A(_0607_),
    .X(_0608_));
 sg13g2_buf_1 _3862_ (.A(_2592_),
    .X(_0609_));
 sg13g2_nor2_1 _3863_ (.A(_0496_),
    .B(net41),
    .Y(_0610_));
 sg13g2_a21oi_1 _3864_ (.A1(_0525_),
    .A2(_0608_),
    .Y(_0611_),
    .B1(_0610_));
 sg13g2_nor2_1 _3865_ (.A(net94),
    .B(_0611_),
    .Y(_0036_));
 sg13g2_nand2_1 _3866_ (.Y(_0612_),
    .A(_0495_),
    .B(_2702_));
 sg13g2_o21ai_1 _3867_ (.B1(_0502_),
    .Y(_0613_),
    .A1(_0476_),
    .A2(net98));
 sg13g2_a21oi_1 _3868_ (.A1(_0612_),
    .A2(_0613_),
    .Y(_0037_),
    .B1(net93));
 sg13g2_buf_1 _3869_ (.A(net170),
    .X(_0614_));
 sg13g2_nand2_1 _3870_ (.Y(_0615_),
    .A(_0521_),
    .B(_0523_));
 sg13g2_a21oi_1 _3871_ (.A1(net168),
    .A2(_0357_),
    .Y(_0616_),
    .B1(_0500_));
 sg13g2_mux2_1 _3872_ (.A0(_0616_),
    .A1(_0498_),
    .S(_0502_),
    .X(_0617_));
 sg13g2_nand2_1 _3873_ (.Y(_0618_),
    .A(_0525_),
    .B(_0617_));
 sg13g2_o21ai_1 _3874_ (.B1(_0618_),
    .Y(_0619_),
    .A1(_0525_),
    .A2(_0615_));
 sg13g2_nand2_1 _3875_ (.Y(_0620_),
    .A(net169),
    .B(_0354_));
 sg13g2_o21ai_1 _3876_ (.B1(_0620_),
    .Y(_0621_),
    .A1(net116),
    .A2(_0619_));
 sg13g2_nor2_1 _3877_ (.A(_0496_),
    .B(net123),
    .Y(_0622_));
 sg13g2_a21oi_1 _3878_ (.A1(net125),
    .A2(_0621_),
    .Y(_0623_),
    .B1(_0622_));
 sg13g2_nor2_1 _3879_ (.A(_2738_),
    .B(_0623_),
    .Y(_0038_));
 sg13g2_buf_1 _3880_ (.A(net61),
    .X(_0624_));
 sg13g2_mux2_1 _3881_ (.A0(_0522_),
    .A1(_0496_),
    .S(net40),
    .X(_0625_));
 sg13g2_nor2_1 _3882_ (.A(_2738_),
    .B(_0625_),
    .Y(_0039_));
 sg13g2_inv_1 _3883_ (.Y(_0626_),
    .A(_2682_));
 sg13g2_nor2_1 _3884_ (.A(_0626_),
    .B(net41),
    .Y(_0627_));
 sg13g2_a21oi_1 _3885_ (.A1(_2677_),
    .A2(net22),
    .Y(_0628_),
    .B1(_0627_));
 sg13g2_nor2_1 _3886_ (.A(net94),
    .B(_0628_),
    .Y(_0040_));
 sg13g2_nand2_1 _3887_ (.Y(_0629_),
    .A(_2682_),
    .B(net44));
 sg13g2_o21ai_1 _3888_ (.B1(_2668_),
    .Y(_0630_),
    .A1(net58),
    .A2(net98));
 sg13g2_a21oi_1 _3889_ (.A1(_0629_),
    .A2(_0630_),
    .Y(_0041_),
    .B1(net93));
 sg13g2_buf_8 _3890_ (.A(net170),
    .X(_0631_));
 sg13g2_nand2_1 _3891_ (.Y(_0632_),
    .A(_0631_),
    .B(_0495_));
 sg13g2_mux2_1 _3892_ (.A0(\g.g_y[0].g_x[0].t.r_gnl ),
    .A1(_2584_),
    .S(_2585_),
    .X(_0633_));
 sg13g2_mux2_1 _3893_ (.A0(_2617_),
    .A1(_0633_),
    .S(_2686_),
    .X(_0634_));
 sg13g2_buf_1 _3894_ (.A(_0634_),
    .X(_0635_));
 sg13g2_mux2_1 _3895_ (.A0(_0635_),
    .A1(_2676_),
    .S(_2663_),
    .X(_0636_));
 sg13g2_mux2_1 _3896_ (.A0(_2669_),
    .A1(_0636_),
    .S(_2679_),
    .X(_0637_));
 sg13g2_nand2_1 _3897_ (.Y(_0638_),
    .A(_2743_),
    .B(_0637_));
 sg13g2_nand3_1 _3898_ (.B(_0632_),
    .C(_0638_),
    .A(net123),
    .Y(_0639_));
 sg13g2_o21ai_1 _3899_ (.B1(_0639_),
    .Y(_0640_),
    .A1(_2682_),
    .A2(net125));
 sg13g2_nor2_1 _3900_ (.A(net94),
    .B(_0640_),
    .Y(_0042_));
 sg13g2_nand2_1 _3901_ (.Y(_0641_),
    .A(_2682_),
    .B(net43));
 sg13g2_o21ai_1 _3902_ (.B1(_2663_),
    .Y(_0642_),
    .A1(net58),
    .A2(net95));
 sg13g2_buf_1 _3903_ (.A(net126),
    .X(_0643_));
 sg13g2_a21oi_1 _3904_ (.A1(_0641_),
    .A2(_0642_),
    .Y(_0043_),
    .B1(net90));
 sg13g2_mux2_1 _3905_ (.A0(_2608_),
    .A1(_2609_),
    .S(net47),
    .X(_0644_));
 sg13g2_and2_1 _3906_ (.A(net131),
    .B(_0644_),
    .X(_0044_));
 sg13g2_o21ai_1 _3907_ (.B1(net12),
    .Y(_0645_),
    .A1(net183),
    .A2(_2699_));
 sg13g2_and2_1 _3908_ (.A(net182),
    .B(_0645_),
    .X(_0646_));
 sg13g2_buf_1 _3909_ (.A(_0646_),
    .X(_0647_));
 sg13g2_buf_1 _3910_ (.A(net57),
    .X(_0648_));
 sg13g2_mux2_1 _3911_ (.A0(_2676_),
    .A1(_0635_),
    .S(_2663_),
    .X(_0649_));
 sg13g2_inv_1 _3912_ (.Y(_0650_),
    .A(net2));
 sg13g2_nor2_1 _3913_ (.A(_0650_),
    .B(_2679_),
    .Y(_0651_));
 sg13g2_o21ai_1 _3914_ (.B1(_2668_),
    .Y(_0652_),
    .A1(_2677_),
    .A2(_2682_));
 sg13g2_a21oi_1 _3915_ (.A1(_0649_),
    .A2(_0651_),
    .Y(_0653_),
    .B1(_0652_));
 sg13g2_a21oi_1 _3916_ (.A1(_0650_),
    .A2(_2679_),
    .Y(_0654_),
    .B1(_2668_));
 sg13g2_o21ai_1 _3917_ (.B1(_0654_),
    .Y(_0655_),
    .A1(_2679_),
    .A2(_0636_));
 sg13g2_nor2b_1 _3918_ (.A(_0653_),
    .B_N(_0655_),
    .Y(_0656_));
 sg13g2_nand3_1 _3919_ (.B(_2846_),
    .C(_2855_),
    .A(_2835_),
    .Y(_0657_));
 sg13g2_nor2_1 _3920_ (.A(_2835_),
    .B(_2858_),
    .Y(_0658_));
 sg13g2_nor2_1 _3921_ (.A(_2853_),
    .B(_0658_),
    .Y(_0659_));
 sg13g2_a21oi_1 _3922_ (.A1(net173),
    .A2(_2809_),
    .Y(_0660_),
    .B1(_2836_));
 sg13g2_mux2_1 _3923_ (.A0(_0660_),
    .A1(_2868_),
    .S(_2844_),
    .X(_0661_));
 sg13g2_nor2_1 _3924_ (.A(_2835_),
    .B(_2852_),
    .Y(_0662_));
 sg13g2_a21oi_1 _3925_ (.A1(net122),
    .A2(_0661_),
    .Y(_0663_),
    .B1(_0662_));
 sg13g2_a22oi_1 _3926_ (.Y(_0664_),
    .B1(_0663_),
    .B2(_2853_),
    .A2(_0659_),
    .A1(_0657_));
 sg13g2_mux2_1 _3927_ (.A0(_0656_),
    .A1(_0664_),
    .S(_2665_),
    .X(_0665_));
 sg13g2_nand3b_1 _3928_ (.B(_2616_),
    .C(_2628_),
    .Y(_0666_),
    .A_N(net179));
 sg13g2_nand2b_1 _3929_ (.Y(_0667_),
    .B(net179),
    .A_N(_2630_));
 sg13g2_and2_1 _3930_ (.A(_2614_),
    .B(_0667_),
    .X(_0668_));
 sg13g2_mux2_1 _3931_ (.A0(_2741_),
    .A1(_2633_),
    .S(net179),
    .X(_0669_));
 sg13g2_a22oi_1 _3932_ (.Y(_0670_),
    .B1(_0669_),
    .B2(_2615_),
    .A2(_0668_),
    .A1(_0666_));
 sg13g2_buf_2 _3933_ (.A(\g.g_y[3].g_x[1].t.r_v ),
    .X(_0671_));
 sg13g2_buf_2 _3934_ (.A(\g.g_y[3].g_x[1].t.out_sc ),
    .X(_0672_));
 sg13g2_buf_2 _3935_ (.A(\g.g_y[3].g_x[1].t.r_d ),
    .X(_0673_));
 sg13g2_mux2_1 _3936_ (.A0(\g.g_y[3].g_x[1].t.r_gnl ),
    .A1(_0672_),
    .S(_0673_),
    .X(_0674_));
 sg13g2_buf_1 _3937_ (.A(\g.g_y[3].g_x[1].t.r_ghl ),
    .X(_0675_));
 sg13g2_nand2b_1 _3938_ (.Y(_0676_),
    .B(_0671_),
    .A_N(_0675_));
 sg13g2_o21ai_1 _3939_ (.B1(_0676_),
    .Y(_0677_),
    .A1(_0671_),
    .A2(_0674_));
 sg13g2_mux2_1 _3940_ (.A0(_2670_),
    .A1(\g.g_y[2].g_x[0].t.r_gnl ),
    .S(_2671_),
    .X(_0678_));
 sg13g2_buf_1 _3941_ (.A(\g.g_y[2].g_x[0].t.r_h ),
    .X(_0679_));
 sg13g2_mux2_1 _3942_ (.A0(_2673_),
    .A1(_0678_),
    .S(net161),
    .X(_0680_));
 sg13g2_buf_1 _3943_ (.A(_0680_),
    .X(_0681_));
 sg13g2_buf_1 _3944_ (.A(\g.g_y[2].g_x[1].t.r_d ),
    .X(_0682_));
 sg13g2_buf_2 _3945_ (.A(\g.g_y[2].g_x[1].t.r_h ),
    .X(_0683_));
 sg13g2_nor2b_1 _3946_ (.A(_0682_),
    .B_N(_0683_),
    .Y(_0684_));
 sg13g2_nor2_1 _3947_ (.A(_0683_),
    .B(_0682_),
    .Y(_0685_));
 sg13g2_mux2_1 _3948_ (.A0(_2838_),
    .A1(\g.g_y[2].g_x[2].t.r_gnl ),
    .S(_2839_),
    .X(_0686_));
 sg13g2_buf_2 _3949_ (.A(\g.g_y[2].g_x[2].t.r_h ),
    .X(_0687_));
 sg13g2_mux2_1 _3950_ (.A0(_0686_),
    .A1(_2841_),
    .S(_0687_),
    .X(_0688_));
 sg13g2_buf_1 _3951_ (.A(_0688_),
    .X(_0689_));
 sg13g2_a22oi_1 _3952_ (.Y(_0690_),
    .B1(_0685_),
    .B2(_0689_),
    .A2(_0684_),
    .A1(_0681_));
 sg13g2_buf_2 _3953_ (.A(\g.g_y[2].g_x[1].t.out_sc ),
    .X(_0691_));
 sg13g2_nand2b_1 _3954_ (.Y(_0692_),
    .B(_0682_),
    .A_N(_0691_));
 sg13g2_o21ai_1 _3955_ (.B1(_0692_),
    .Y(_0693_),
    .A1(_0677_),
    .A2(_0690_));
 sg13g2_buf_1 _3956_ (.A(_0682_),
    .X(_0694_));
 sg13g2_mux2_1 _3957_ (.A0(_0681_),
    .A1(_0689_),
    .S(_0683_),
    .X(_0695_));
 sg13g2_nand2_1 _3958_ (.Y(_0696_),
    .A(net114),
    .B(_0677_));
 sg13g2_o21ai_1 _3959_ (.B1(_0696_),
    .Y(_0697_),
    .A1(net114),
    .A2(_0695_));
 sg13g2_buf_1 _3960_ (.A(\g.g_y[2].g_x[1].t.r_v ),
    .X(_0698_));
 sg13g2_mux2_1 _3961_ (.A0(_0693_),
    .A1(_0697_),
    .S(_0698_),
    .X(_0699_));
 sg13g2_mux2_1 _3962_ (.A0(_0670_),
    .A1(_0699_),
    .S(_2612_),
    .X(_0700_));
 sg13g2_mux2_1 _3963_ (.A0(_0665_),
    .A1(_0700_),
    .S(_2609_),
    .X(_0701_));
 sg13g2_buf_1 _3964_ (.A(net57),
    .X(_0702_));
 sg13g2_o21ai_1 _3965_ (.B1(net176),
    .Y(_0703_),
    .A1(_2611_),
    .A2(net38));
 sg13g2_a21oi_1 _3966_ (.A1(_0648_),
    .A2(_0701_),
    .Y(_0045_),
    .B1(_0703_));
 sg13g2_nand2_2 _3967_ (.Y(_0704_),
    .A(_2587_),
    .B(_0645_));
 sg13g2_mux2_1 _3968_ (.A0(_0664_),
    .A1(_0656_),
    .S(_2665_),
    .X(_0705_));
 sg13g2_mux2_1 _3969_ (.A0(_0699_),
    .A1(_0670_),
    .S(_2612_),
    .X(_0706_));
 sg13g2_nor3_1 _3970_ (.A(_0704_),
    .B(_0705_),
    .C(_0706_),
    .Y(_0707_));
 sg13g2_o21ai_1 _3971_ (.B1(net117),
    .Y(_0708_),
    .A1(\g.g_y[1].g_x[1].t.r_gnl ),
    .A2(net38));
 sg13g2_nor2_1 _3972_ (.A(_0707_),
    .B(_0708_),
    .Y(_0046_));
 sg13g2_nand2_1 _3973_ (.Y(_0709_),
    .A(_2608_),
    .B(net44));
 sg13g2_o21ai_1 _3974_ (.B1(_2665_),
    .Y(_0710_),
    .A1(net58),
    .A2(net98));
 sg13g2_a21oi_1 _3975_ (.A1(_0709_),
    .A2(_0710_),
    .Y(_0047_),
    .B1(_0643_));
 sg13g2_mux2_1 _3976_ (.A0(_0700_),
    .A1(_0665_),
    .S(_2609_),
    .X(_0711_));
 sg13g2_a22oi_1 _3977_ (.Y(_0712_),
    .B1(_2723_),
    .B2(_2682_),
    .A2(_2720_),
    .A1(_2608_));
 sg13g2_o21ai_1 _3978_ (.B1(_0712_),
    .Y(_0048_),
    .A1(net64),
    .A2(_0711_));
 sg13g2_nand2_1 _3979_ (.Y(_0713_),
    .A(_2608_),
    .B(net43));
 sg13g2_o21ai_1 _3980_ (.B1(_2612_),
    .Y(_0714_),
    .A1(net58),
    .A2(net95));
 sg13g2_a21oi_1 _3981_ (.A1(_0713_),
    .A2(_0714_),
    .Y(_0049_),
    .B1(net90));
 sg13g2_nor2_1 _3982_ (.A(_2859_),
    .B(net41),
    .Y(_0715_));
 sg13g2_a21oi_1 _3983_ (.A1(_2857_),
    .A2(_0608_),
    .Y(_0716_),
    .B1(_0715_));
 sg13g2_nor2_1 _3984_ (.A(net94),
    .B(_0716_),
    .Y(_0050_));
 sg13g2_buf_1 _3985_ (.A(net66),
    .X(_0717_));
 sg13g2_mux2_1 _3986_ (.A0(_2854_),
    .A1(_2859_),
    .S(net37),
    .X(_0718_));
 sg13g2_nor2_1 _3987_ (.A(net94),
    .B(_0718_),
    .Y(_0051_));
 sg13g2_nor2_1 _3988_ (.A(_2858_),
    .B(net121),
    .Y(_0719_));
 sg13g2_mux2_1 _3989_ (.A0(_0661_),
    .A1(_2865_),
    .S(net122),
    .X(_0720_));
 sg13g2_nand2_1 _3990_ (.Y(_0721_),
    .A(net169),
    .B(_2608_));
 sg13g2_o21ai_1 _3991_ (.B1(_0721_),
    .Y(_0722_),
    .A1(net120),
    .A2(_0720_));
 sg13g2_nor2_1 _3992_ (.A(_2894_),
    .B(_0722_),
    .Y(_0723_));
 sg13g2_nor3_1 _3993_ (.A(_2890_),
    .B(_0719_),
    .C(_0723_),
    .Y(_0052_));
 sg13g2_mux2_1 _3994_ (.A0(_2845_),
    .A1(_2859_),
    .S(net40),
    .X(_0724_));
 sg13g2_nor2_1 _3995_ (.A(net94),
    .B(_0724_),
    .Y(_0053_));
 sg13g2_mux2_1 _3996_ (.A0(_2766_),
    .A1(_2767_),
    .S(net47),
    .X(_0725_));
 sg13g2_and2_1 _3997_ (.A(net131),
    .B(_0725_),
    .X(_0054_));
 sg13g2_buf_1 _3998_ (.A(net184),
    .X(_0726_));
 sg13g2_o21ai_1 _3999_ (.B1(net12),
    .Y(_0727_),
    .A1(net183),
    .A2(_2726_));
 sg13g2_nand2_1 _4000_ (.Y(_0728_),
    .A(net182),
    .B(_0727_));
 sg13g2_buf_1 _4001_ (.A(_0728_),
    .X(_0729_));
 sg13g2_nand3_1 _4002_ (.B(_0726_),
    .C(net56),
    .A(_2770_),
    .Y(_0730_));
 sg13g2_inv_1 _4003_ (.Y(_0731_),
    .A(_2767_));
 sg13g2_nand3b_1 _4004_ (.B(_2853_),
    .C(_0657_),
    .Y(_0732_),
    .A_N(_0658_));
 sg13g2_o21ai_1 _4005_ (.B1(_2854_),
    .Y(_0733_),
    .A1(net122),
    .A2(_2848_));
 sg13g2_a21oi_1 _4006_ (.A1(net122),
    .A2(_0661_),
    .Y(_0734_),
    .B1(_0733_));
 sg13g2_nor2_1 _4007_ (.A(net171),
    .B(_0734_),
    .Y(_0735_));
 sg13g2_and4_1 _4008_ (.A(_0424_),
    .B(_0439_),
    .C(_0422_),
    .D(_0437_),
    .X(_0736_));
 sg13g2_and3_1 _4009_ (.X(_0737_),
    .A(_0423_),
    .B(net118),
    .C(_0444_));
 sg13g2_nor3_1 _4010_ (.A(_0423_),
    .B(net118),
    .C(_0380_),
    .Y(_0738_));
 sg13g2_nor3_1 _4011_ (.A(_0424_),
    .B(_0439_),
    .C(_0422_),
    .Y(_0739_));
 sg13g2_or4_1 _4012_ (.A(_0736_),
    .B(_0737_),
    .C(_0738_),
    .D(_0739_),
    .X(_0740_));
 sg13g2_a22oi_1 _4013_ (.Y(_0741_),
    .B1(_0740_),
    .B2(net171),
    .A2(_0735_),
    .A1(_0732_));
 sg13g2_and2_1 _4014_ (.A(net182),
    .B(_0727_),
    .X(_0742_));
 sg13g2_buf_2 _4015_ (.A(_0742_),
    .X(_0743_));
 sg13g2_nand4_1 _4016_ (.B(net181),
    .C(_0741_),
    .A(_0731_),
    .Y(_0744_),
    .D(_0743_));
 sg13g2_nor2b_1 _4017_ (.A(_0687_),
    .B_N(_2841_),
    .Y(_0745_));
 sg13g2_a21o_1 _4018_ (.A2(_0686_),
    .A1(_0687_),
    .B1(_0745_),
    .X(_0746_));
 sg13g2_buf_1 _4019_ (.A(\g.g_y[2].g_x[3].t.r_h ),
    .X(_0747_));
 sg13g2_inv_1 _4020_ (.Y(_0748_),
    .A(_0747_));
 sg13g2_buf_1 _4021_ (.A(\g.g_y[2].g_x[3].t.r_d ),
    .X(_0749_));
 sg13g2_nor2_1 _4022_ (.A(_0748_),
    .B(net159),
    .Y(_0750_));
 sg13g2_nor2_1 _4023_ (.A(_0747_),
    .B(_0749_),
    .Y(_0751_));
 sg13g2_mux2_1 _4024_ (.A0(_0430_),
    .A1(\g.g_y[2].g_x[4].t.r_gnl ),
    .S(_0431_),
    .X(_0752_));
 sg13g2_buf_2 _4025_ (.A(\g.g_y[2].g_x[4].t.r_h ),
    .X(_0753_));
 sg13g2_mux2_1 _4026_ (.A0(_0752_),
    .A1(_0429_),
    .S(_0753_),
    .X(_0754_));
 sg13g2_a22oi_1 _4027_ (.Y(_0755_),
    .B1(_0751_),
    .B2(_0754_),
    .A2(_0750_),
    .A1(_0746_));
 sg13g2_buf_1 _4028_ (.A(\g.g_y[2].g_x[3].t.r_v ),
    .X(_0756_));
 sg13g2_inv_1 _4029_ (.Y(_0757_),
    .A(_0756_));
 sg13g2_buf_2 _4030_ (.A(\g.g_y[3].g_x[3].t.r_ghl ),
    .X(_0758_));
 sg13g2_buf_2 _4031_ (.A(\g.g_y[3].g_x[3].t.out_sc ),
    .X(_0759_));
 sg13g2_buf_2 _4032_ (.A(\g.g_y[3].g_x[3].t.r_d ),
    .X(_0760_));
 sg13g2_mux2_1 _4033_ (.A0(\g.g_y[3].g_x[3].t.r_gnl ),
    .A1(_0759_),
    .S(_0760_),
    .X(_0761_));
 sg13g2_buf_2 _4034_ (.A(\g.g_y[3].g_x[3].t.r_v ),
    .X(_0762_));
 sg13g2_inv_1 _4035_ (.Y(_0763_),
    .A(_0762_));
 sg13g2_mux2_1 _4036_ (.A0(_0758_),
    .A1(_0761_),
    .S(_0763_),
    .X(_0764_));
 sg13g2_nand2_1 _4037_ (.Y(_0765_),
    .A(_0757_),
    .B(_0764_));
 sg13g2_inv_1 _4038_ (.Y(_0766_),
    .A(net159));
 sg13g2_buf_2 _4039_ (.A(\g.g_y[2].g_x[3].t.out_sc ),
    .X(_0767_));
 sg13g2_nor2_1 _4040_ (.A(_0766_),
    .B(_0767_),
    .Y(_0768_));
 sg13g2_nand2_1 _4041_ (.Y(_0769_),
    .A(_0757_),
    .B(_0768_));
 sg13g2_o21ai_1 _4042_ (.B1(_0769_),
    .Y(_0770_),
    .A1(_0755_),
    .A2(_0765_));
 sg13g2_a21oi_1 _4043_ (.A1(_0687_),
    .A2(_0686_),
    .Y(_0771_),
    .B1(_0745_));
 sg13g2_nand2b_1 _4044_ (.Y(_0772_),
    .B(_0753_),
    .A_N(_0429_));
 sg13g2_o21ai_1 _4045_ (.B1(_0772_),
    .Y(_0773_),
    .A1(_0753_),
    .A2(_0752_));
 sg13g2_mux2_1 _4046_ (.A0(_0771_),
    .A1(_0773_),
    .S(_0747_),
    .X(_0774_));
 sg13g2_a21oi_1 _4047_ (.A1(net159),
    .A2(_0764_),
    .Y(_0775_),
    .B1(_0757_));
 sg13g2_o21ai_1 _4048_ (.B1(_0775_),
    .Y(_0776_),
    .A1(net159),
    .A2(_0774_));
 sg13g2_buf_1 _4049_ (.A(_2771_),
    .X(_0777_));
 sg13g2_nand3b_1 _4050_ (.B(_0776_),
    .C(net113),
    .Y(_0778_),
    .A_N(_0770_));
 sg13g2_nand3_1 _4051_ (.B(_2775_),
    .C(_2786_),
    .A(_0332_),
    .Y(_0779_));
 sg13g2_nor2_1 _4052_ (.A(_2788_),
    .B(_0332_),
    .Y(_0780_));
 sg13g2_nor3_1 _4053_ (.A(net113),
    .B(_2774_),
    .C(_0780_),
    .Y(_0781_));
 sg13g2_nand2_1 _4054_ (.Y(_0782_),
    .A(_0332_),
    .B(_0322_));
 sg13g2_nor2_1 _4055_ (.A(_0332_),
    .B(_2765_),
    .Y(_0783_));
 sg13g2_nor3_1 _4056_ (.A(net113),
    .B(_2773_),
    .C(_0783_),
    .Y(_0784_));
 sg13g2_a22oi_1 _4057_ (.Y(_0785_),
    .B1(_0782_),
    .B2(_0784_),
    .A2(_0781_),
    .A1(_0779_));
 sg13g2_and2_1 _4058_ (.A(_0778_),
    .B(_0785_),
    .X(_0786_));
 sg13g2_or4_1 _4059_ (.A(_0731_),
    .B(_2709_),
    .C(_0728_),
    .D(_0786_),
    .X(_0787_));
 sg13g2_nand3_1 _4060_ (.B(_0744_),
    .C(_0787_),
    .A(_0730_),
    .Y(_0055_));
 sg13g2_nand2b_1 _4061_ (.Y(_0788_),
    .B(net171),
    .A_N(_0734_));
 sg13g2_a21oi_1 _4062_ (.A1(_2853_),
    .A2(_0657_),
    .Y(_0789_),
    .B1(_0788_));
 sg13g2_nand2_1 _4063_ (.Y(_0790_),
    .A(net113),
    .B(_2774_));
 sg13g2_a21oi_1 _4064_ (.A1(_2795_),
    .A2(_0782_),
    .Y(_0791_),
    .B1(_0790_));
 sg13g2_nand3_1 _4065_ (.B(_2853_),
    .C(_0658_),
    .A(_2862_),
    .Y(_0792_));
 sg13g2_nand2_1 _4066_ (.Y(_0793_),
    .A(_2851_),
    .B(_0738_));
 sg13g2_nand3_1 _4067_ (.B(_2773_),
    .C(_0780_),
    .A(_0777_),
    .Y(_0794_));
 sg13g2_nand4_1 _4068_ (.B(_0792_),
    .C(_0793_),
    .A(_0743_),
    .Y(_0795_),
    .D(_0794_));
 sg13g2_nor3_1 _4069_ (.A(_0789_),
    .B(_0791_),
    .C(_0795_),
    .Y(_0796_));
 sg13g2_nor2_1 _4070_ (.A(net118),
    .B(_0422_),
    .Y(_0797_));
 sg13g2_a21o_1 _4071_ (.A2(_0444_),
    .A1(net118),
    .B1(_0797_),
    .X(_0798_));
 sg13g2_a21oi_1 _4072_ (.A1(_0423_),
    .A2(_0798_),
    .Y(_0799_),
    .B1(_0736_));
 sg13g2_nor2_1 _4073_ (.A(net171),
    .B(_0799_),
    .Y(_0800_));
 sg13g2_nand2b_1 _4074_ (.Y(_0801_),
    .B(_0776_),
    .A_N(_0770_));
 sg13g2_o21ai_1 _4075_ (.B1(_0777_),
    .Y(_0802_),
    .A1(_2774_),
    .A2(_0779_));
 sg13g2_o21ai_1 _4076_ (.B1(_0802_),
    .Y(_0803_),
    .A1(net113),
    .A2(_0801_));
 sg13g2_nor2b_1 _4077_ (.A(_0800_),
    .B_N(_0803_),
    .Y(_0804_));
 sg13g2_buf_1 _4078_ (.A(_0743_),
    .X(_0805_));
 sg13g2_o21ai_1 _4079_ (.B1(net176),
    .Y(_0806_),
    .A1(\g.g_y[1].g_x[3].t.r_gnl ),
    .A2(net36));
 sg13g2_a21oi_1 _4080_ (.A1(_0796_),
    .A2(_0804_),
    .Y(_0056_),
    .B1(_0806_));
 sg13g2_buf_1 _4081_ (.A(net66),
    .X(_0807_));
 sg13g2_nand2_1 _4082_ (.Y(_0808_),
    .A(_2766_),
    .B(net35));
 sg13g2_buf_1 _4083_ (.A(net129),
    .X(_0809_));
 sg13g2_o21ai_1 _4084_ (.B1(net171),
    .Y(_0810_),
    .A1(net58),
    .A2(net89));
 sg13g2_a21oi_1 _4085_ (.A1(_0808_),
    .A2(_0810_),
    .Y(_0057_),
    .B1(net90));
 sg13g2_nor2_1 _4086_ (.A(net183),
    .B(_2713_),
    .Y(_0811_));
 sg13g2_buf_1 _4087_ (.A(_0811_),
    .X(_0812_));
 sg13g2_nand3_1 _4088_ (.B(net88),
    .C(_0741_),
    .A(_2767_),
    .Y(_0813_));
 sg13g2_or3_1 _4089_ (.A(_2767_),
    .B(_2715_),
    .C(_0786_),
    .X(_0814_));
 sg13g2_buf_1 _4090_ (.A(_2719_),
    .X(_0815_));
 sg13g2_a22oi_1 _4091_ (.Y(_0816_),
    .B1(net96),
    .B2(_2858_),
    .A2(net55),
    .A1(_2766_));
 sg13g2_nand3_1 _4092_ (.B(_0814_),
    .C(_0816_),
    .A(_0813_),
    .Y(_0058_));
 sg13g2_nand2_1 _4093_ (.Y(_0817_),
    .A(_2766_),
    .B(net43));
 sg13g2_buf_1 _4094_ (.A(net99),
    .X(_0818_));
 sg13g2_o21ai_1 _4095_ (.B1(net113),
    .Y(_0819_),
    .A1(_0818_),
    .A2(net95));
 sg13g2_a21oi_1 _4096_ (.A1(_0817_),
    .A2(_0819_),
    .Y(_0059_),
    .B1(_0643_));
 sg13g2_nor2_1 _4097_ (.A(_0381_),
    .B(_0609_),
    .Y(_0820_));
 sg13g2_a21oi_1 _4098_ (.A1(net118),
    .A2(net22),
    .Y(_0821_),
    .B1(_0820_));
 sg13g2_nor2_1 _4099_ (.A(net94),
    .B(_0821_),
    .Y(_0060_));
 sg13g2_buf_1 _4100_ (.A(net126),
    .X(_0822_));
 sg13g2_mux2_1 _4101_ (.A0(_0424_),
    .A1(_0381_),
    .S(net37),
    .X(_0823_));
 sg13g2_nor2_1 _4102_ (.A(_0822_),
    .B(_0823_),
    .Y(_0061_));
 sg13g2_nor2_1 _4103_ (.A(_0380_),
    .B(_2891_),
    .Y(_0824_));
 sg13g2_a22oi_1 _4104_ (.Y(_0825_),
    .B1(_0447_),
    .B2(_0448_),
    .A2(_0422_),
    .A1(_0423_));
 sg13g2_mux2_1 _4105_ (.A0(_0444_),
    .A1(_0825_),
    .S(net118),
    .X(_0826_));
 sg13g2_nand2_1 _4106_ (.Y(_0827_),
    .A(net169),
    .B(_2766_));
 sg13g2_o21ai_1 _4107_ (.B1(_0827_),
    .Y(_0828_),
    .A1(_2896_),
    .A2(_0826_));
 sg13g2_nor2_1 _4108_ (.A(_2894_),
    .B(_0828_),
    .Y(_0829_));
 sg13g2_nor3_1 _4109_ (.A(_2890_),
    .B(_0824_),
    .C(_0829_),
    .Y(_0062_));
 sg13g2_mux2_1 _4110_ (.A0(_0415_),
    .A1(_0381_),
    .S(net40),
    .X(_0830_));
 sg13g2_nor2_1 _4111_ (.A(_0822_),
    .B(_0830_),
    .Y(_0063_));
 sg13g2_mux2_1 _4112_ (.A0(_0336_),
    .A1(_0337_),
    .S(net47),
    .X(_0831_));
 sg13g2_and2_1 _4113_ (.A(net131),
    .B(_0831_),
    .X(_0064_));
 sg13g2_a21oi_1 _4114_ (.A1(net171),
    .A2(_2850_),
    .Y(_0832_),
    .B1(_0417_));
 sg13g2_and2_1 _4115_ (.A(_0425_),
    .B(_0437_),
    .X(_0833_));
 sg13g2_mux4_1 _4116_ (.S0(_0424_),
    .A0(_0381_),
    .A1(_0832_),
    .A2(_0833_),
    .A3(_0444_),
    .S1(net118),
    .X(_0834_));
 sg13g2_a21oi_1 _4117_ (.A1(net163),
    .A2(_0531_),
    .Y(_0835_),
    .B1(_0578_));
 sg13g2_nor2_1 _4118_ (.A(_0580_),
    .B(_0835_),
    .Y(_0836_));
 sg13g2_nand2_1 _4119_ (.Y(_0837_),
    .A(_0580_),
    .B(_0577_));
 sg13g2_nor2b_1 _4120_ (.A(_0836_),
    .B_N(_0837_),
    .Y(_0838_));
 sg13g2_mux4_1 _4121_ (.S0(_0570_),
    .A0(_0588_),
    .A1(_0585_),
    .A2(_0582_),
    .A3(_0838_),
    .S1(_0590_),
    .X(_0839_));
 sg13g2_mux2_1 _4122_ (.A0(_0834_),
    .A1(_0839_),
    .S(_0420_),
    .X(_0840_));
 sg13g2_buf_2 _4123_ (.A(\g.g_y[2].g_x[5].t.r_h ),
    .X(_0841_));
 sg13g2_inv_2 _4124_ (.Y(_0842_),
    .A(_0841_));
 sg13g2_buf_1 _4125_ (.A(\g.g_y[2].g_x[5].t.r_d ),
    .X(_0843_));
 sg13g2_nor2_1 _4126_ (.A(_0842_),
    .B(net158),
    .Y(_0844_));
 sg13g2_buf_1 _4127_ (.A(\g.g_y[2].g_x[5].t.r_v ),
    .X(_0845_));
 sg13g2_buf_1 _4128_ (.A(\g.g_y[2].g_x[6].t.r_h ),
    .X(_0846_));
 sg13g2_mux2_1 _4129_ (.A0(_0572_),
    .A1(\g.g_y[2].g_x[6].t.r_gnl ),
    .S(_0573_),
    .X(_0847_));
 sg13g2_buf_2 _4130_ (.A(_0847_),
    .X(_0848_));
 sg13g2_nand2b_1 _4131_ (.Y(_0849_),
    .B(net156),
    .A_N(_0575_));
 sg13g2_o21ai_1 _4132_ (.B1(_0849_),
    .Y(_0850_),
    .A1(_0846_),
    .A2(_0848_));
 sg13g2_buf_2 _4133_ (.A(\g.g_y[3].g_x[5].t.r_v ),
    .X(_0851_));
 sg13g2_buf_2 _4134_ (.A(\g.g_y[3].g_x[5].t.out_sc ),
    .X(_0852_));
 sg13g2_buf_2 _4135_ (.A(\g.g_y[3].g_x[5].t.r_d ),
    .X(_0853_));
 sg13g2_mux2_1 _4136_ (.A0(\g.g_y[3].g_x[5].t.r_gnl ),
    .A1(_0852_),
    .S(_0853_),
    .X(_0854_));
 sg13g2_buf_1 _4137_ (.A(\g.g_y[3].g_x[5].t.r_ghl ),
    .X(_0855_));
 sg13g2_nand2b_1 _4138_ (.Y(_0856_),
    .B(_0851_),
    .A_N(_0855_));
 sg13g2_o21ai_1 _4139_ (.B1(_0856_),
    .Y(_0857_),
    .A1(_0851_),
    .A2(_0854_));
 sg13g2_nor2_1 _4140_ (.A(net157),
    .B(_0857_),
    .Y(_0858_));
 sg13g2_mux2_1 _4141_ (.A0(_0429_),
    .A1(_0752_),
    .S(_0753_),
    .X(_0859_));
 sg13g2_buf_2 _4142_ (.A(_0859_),
    .X(_0860_));
 sg13g2_a22oi_1 _4143_ (.Y(_0861_),
    .B1(_0858_),
    .B2(_0860_),
    .A2(_0850_),
    .A1(net157));
 sg13g2_buf_1 _4144_ (.A(\g.g_y[2].g_x[5].t.out_sc ),
    .X(_0862_));
 sg13g2_inv_1 _4145_ (.Y(_0863_),
    .A(_0851_));
 sg13g2_mux2_1 _4146_ (.A0(_0855_),
    .A1(_0854_),
    .S(_0863_),
    .X(_0864_));
 sg13g2_buf_1 _4147_ (.A(_0864_),
    .X(_0865_));
 sg13g2_mux2_1 _4148_ (.A0(net155),
    .A1(_0865_),
    .S(net157),
    .X(_0866_));
 sg13g2_nor3_1 _4149_ (.A(net157),
    .B(_0857_),
    .C(_0850_),
    .Y(_0867_));
 sg13g2_nor2b_1 _4150_ (.A(_0860_),
    .B_N(net157),
    .Y(_0868_));
 sg13g2_nor4_1 _4151_ (.A(_0841_),
    .B(net158),
    .C(_0867_),
    .D(_0868_),
    .Y(_0869_));
 sg13g2_a221oi_1 _4152_ (.B2(net158),
    .C1(_0869_),
    .B1(_0866_),
    .A1(_0844_),
    .Y(_0870_),
    .A2(_0861_));
 sg13g2_a21o_1 _4153_ (.A2(_0481_),
    .A1(_0367_),
    .B1(_0374_),
    .X(_0871_));
 sg13g2_nor2b_1 _4154_ (.A(net167),
    .B_N(_0363_),
    .Y(_0872_));
 sg13g2_nor2_1 _4155_ (.A(_0363_),
    .B(net167),
    .Y(_0873_));
 sg13g2_a22oi_1 _4156_ (.Y(_0874_),
    .B1(_0873_),
    .B2(_0360_),
    .A2(_0872_),
    .A1(_0489_));
 sg13g2_nand2b_1 _4157_ (.Y(_0875_),
    .B(_0361_),
    .A_N(_0364_));
 sg13g2_o21ai_1 _4158_ (.B1(_0875_),
    .Y(_0876_),
    .A1(_0353_),
    .A2(_0874_));
 sg13g2_mux2_1 _4159_ (.A0(_0871_),
    .A1(_0876_),
    .S(_0352_),
    .X(_0877_));
 sg13g2_mux2_1 _4160_ (.A0(_0870_),
    .A1(_0877_),
    .S(_0370_),
    .X(_0878_));
 sg13g2_mux2_1 _4161_ (.A0(_0840_),
    .A1(_0878_),
    .S(_0337_),
    .X(_0879_));
 sg13g2_o21ai_1 _4162_ (.B1(net176),
    .Y(_0880_),
    .A1(_0340_),
    .A2(net38));
 sg13g2_a21oi_1 _4163_ (.A1(_0648_),
    .A2(_0879_),
    .Y(_0065_),
    .B1(_0880_));
 sg13g2_mux2_1 _4164_ (.A0(_0839_),
    .A1(_0834_),
    .S(_0420_),
    .X(_0881_));
 sg13g2_mux2_1 _4165_ (.A0(_0870_),
    .A1(_0877_),
    .S(_0335_),
    .X(_0882_));
 sg13g2_nor3_1 _4166_ (.A(_0704_),
    .B(_0881_),
    .C(_0882_),
    .Y(_0883_));
 sg13g2_o21ai_1 _4167_ (.B1(net117),
    .Y(_0884_),
    .A1(\g.g_y[1].g_x[5].t.r_gnl ),
    .A2(net38));
 sg13g2_nor2_1 _4168_ (.A(_0883_),
    .B(_0884_),
    .Y(_0066_));
 sg13g2_nand2_1 _4169_ (.Y(_0885_),
    .A(_0336_),
    .B(net35));
 sg13g2_o21ai_1 _4170_ (.B1(_0420_),
    .Y(_0886_),
    .A1(_0818_),
    .A2(net89));
 sg13g2_a21oi_1 _4171_ (.A1(_0885_),
    .A2(_0886_),
    .Y(_0067_),
    .B1(net90));
 sg13g2_mux2_1 _4172_ (.A0(_0878_),
    .A1(_0840_),
    .S(_0337_),
    .X(_0887_));
 sg13g2_a22oi_1 _4173_ (.Y(_0888_),
    .B1(net62),
    .B2(_0380_),
    .A2(net63),
    .A1(_0336_));
 sg13g2_o21ai_1 _4174_ (.B1(_0888_),
    .Y(_0068_),
    .A1(net64),
    .A2(_0887_));
 sg13g2_buf_1 _4175_ (.A(net61),
    .X(_0889_));
 sg13g2_nand2_1 _4176_ (.Y(_0890_),
    .A(_0336_),
    .B(net34));
 sg13g2_buf_1 _4177_ (.A(net127),
    .X(_0891_));
 sg13g2_o21ai_1 _4178_ (.B1(_0335_),
    .Y(_0892_),
    .A1(net54),
    .A2(net86));
 sg13g2_a21oi_1 _4179_ (.A1(_0890_),
    .A2(_0892_),
    .Y(_0069_),
    .B1(net90));
 sg13g2_nor2_1 _4180_ (.A(_0588_),
    .B(_0609_),
    .Y(_0893_));
 sg13g2_a21oi_1 _4181_ (.A1(_0590_),
    .A2(net22),
    .Y(_0894_),
    .B1(_0893_));
 sg13g2_nor2_1 _4182_ (.A(net87),
    .B(_0894_),
    .Y(_0070_));
 sg13g2_nand2_1 _4183_ (.Y(_0895_),
    .A(_0587_),
    .B(_0807_));
 sg13g2_o21ai_1 _4184_ (.B1(_0570_),
    .Y(_0896_),
    .A1(net54),
    .A2(net89));
 sg13g2_a21oi_1 _4185_ (.A1(_0895_),
    .A2(_0896_),
    .Y(_0071_),
    .B1(net90));
 sg13g2_nor2_1 _4186_ (.A(_0587_),
    .B(_2891_),
    .Y(_0897_));
 sg13g2_nand2b_1 _4187_ (.Y(_0898_),
    .B(_0837_),
    .A_N(_0836_));
 sg13g2_nand2_1 _4188_ (.Y(_0899_),
    .A(_0590_),
    .B(_0586_));
 sg13g2_o21ai_1 _4189_ (.B1(_0899_),
    .Y(_0900_),
    .A1(_0590_),
    .A2(_0898_));
 sg13g2_nand2_1 _4190_ (.Y(_0901_),
    .A(net169),
    .B(_0336_));
 sg13g2_o21ai_1 _4191_ (.B1(_0901_),
    .Y(_0902_),
    .A1(net120),
    .A2(_0900_));
 sg13g2_nor2_1 _4192_ (.A(net91),
    .B(_0902_),
    .Y(_0903_));
 sg13g2_nor3_1 _4193_ (.A(net92),
    .B(_0897_),
    .C(_0903_),
    .Y(_0072_));
 sg13g2_nand2_1 _4194_ (.Y(_0904_),
    .A(_0587_),
    .B(net34));
 sg13g2_o21ai_1 _4195_ (.B1(_0580_),
    .Y(_0905_),
    .A1(net54),
    .A2(net86));
 sg13g2_a21oi_1 _4196_ (.A1(_0904_),
    .A2(_0905_),
    .Y(_0073_),
    .B1(net90));
 sg13g2_buf_1 _4197_ (.A(net181),
    .X(_0906_));
 sg13g2_buf_2 _4198_ (.A(_2592_),
    .X(_0907_));
 sg13g2_mux2_1 _4199_ (.A0(_0504_),
    .A1(_0505_),
    .S(net33),
    .X(_0908_));
 sg13g2_and2_1 _4200_ (.A(_0906_),
    .B(_0908_),
    .X(_0074_));
 sg13g2_inv_1 _4201_ (.Y(_0909_),
    .A(_0505_));
 sg13g2_buf_1 _4202_ (.A(_0743_),
    .X(_0910_));
 sg13g2_nand2_1 _4203_ (.Y(_0911_),
    .A(_0571_),
    .B(_0581_));
 sg13g2_mux4_1 _4204_ (.S0(_0590_),
    .A0(_0569_),
    .A1(_0898_),
    .A2(_0587_),
    .A3(_0911_),
    .S1(_0570_),
    .X(_0912_));
 sg13g2_and2_1 _4205_ (.A(_2677_),
    .B(_2667_),
    .X(_0913_));
 sg13g2_a22oi_1 _4206_ (.Y(_0914_),
    .B1(_0649_),
    .B2(_0913_),
    .A2(_0626_),
    .A1(_2679_));
 sg13g2_mux2_1 _4207_ (.A0(_2667_),
    .A1(_0636_),
    .S(_2677_),
    .X(_0915_));
 sg13g2_mux2_1 _4208_ (.A0(_0914_),
    .A1(_0915_),
    .S(_2668_),
    .X(_0916_));
 sg13g2_mux2_1 _4209_ (.A0(_0912_),
    .A1(_0916_),
    .S(_0566_),
    .X(_0917_));
 sg13g2_nand4_1 _4210_ (.B(net160),
    .C(net32),
    .A(_0909_),
    .Y(_0918_),
    .D(_0917_));
 sg13g2_a21oi_1 _4211_ (.A1(_0511_),
    .A2(_0514_),
    .Y(_0919_),
    .B1(_0516_));
 sg13g2_mux4_1 _4212_ (.S0(_0522_),
    .A0(_0520_),
    .A1(_0617_),
    .A2(_0496_),
    .A3(_0919_),
    .S1(_0525_),
    .X(_0920_));
 sg13g2_buf_2 _4213_ (.A(\g.g_y[2].g_x[7].t.r_h ),
    .X(_0921_));
 sg13g2_inv_1 _4214_ (.Y(_0922_),
    .A(_0921_));
 sg13g2_buf_1 _4215_ (.A(\g.g_y[2].g_x[7].t.r_d ),
    .X(_0923_));
 sg13g2_nor2_1 _4216_ (.A(_0922_),
    .B(net154),
    .Y(_0924_));
 sg13g2_buf_1 _4217_ (.A(\g.g_y[2].g_x[7].t.r_v ),
    .X(_0925_));
 sg13g2_nand2b_1 _4218_ (.Y(_0926_),
    .B(net161),
    .A_N(_2673_));
 sg13g2_o21ai_1 _4219_ (.B1(_0926_),
    .Y(_0927_),
    .A1(net161),
    .A2(_0678_));
 sg13g2_nor2b_1 _4220_ (.A(\g.g_y[2].g_x[6].t.r_h ),
    .B_N(_0575_),
    .Y(_0928_));
 sg13g2_a21o_1 _4221_ (.A2(_0848_),
    .A1(net156),
    .B1(_0928_),
    .X(_0929_));
 sg13g2_buf_2 _4222_ (.A(_0929_),
    .X(_0930_));
 sg13g2_a21oi_1 _4223_ (.A1(net153),
    .A2(_0927_),
    .Y(_0931_),
    .B1(_0930_));
 sg13g2_nand2_1 _4224_ (.Y(_0932_),
    .A(_0924_),
    .B(_0931_));
 sg13g2_inv_1 _4225_ (.Y(_0933_),
    .A(net153));
 sg13g2_buf_1 _4226_ (.A(\g.g_y[2].g_x[7].t.out_sc ),
    .X(_0934_));
 sg13g2_nand3_1 _4227_ (.B(net154),
    .C(net152),
    .A(_0933_),
    .Y(_0935_));
 sg13g2_mux2_1 _4228_ (.A0(_0678_),
    .A1(_2673_),
    .S(net161),
    .X(_0936_));
 sg13g2_buf_2 _4229_ (.A(_0936_),
    .X(_0937_));
 sg13g2_inv_2 _4230_ (.Y(_0938_),
    .A(\g.g_y[2].g_x[7].t.r_d ));
 sg13g2_nand2_1 _4231_ (.Y(_0939_),
    .A(_0922_),
    .B(_0938_));
 sg13g2_nor2_1 _4232_ (.A(_0937_),
    .B(_0939_),
    .Y(_0940_));
 sg13g2_o21ai_1 _4233_ (.B1(_0940_),
    .Y(_0941_),
    .A1(_0933_),
    .A2(_0930_));
 sg13g2_mux2_1 _4234_ (.A0(_0937_),
    .A1(_0930_),
    .S(_0922_),
    .X(_0942_));
 sg13g2_nand2_1 _4235_ (.Y(_0943_),
    .A(net153),
    .B(_0938_));
 sg13g2_buf_2 _4236_ (.A(\g.g_y[3].g_x[7].t.r_v ),
    .X(_0944_));
 sg13g2_buf_2 _4237_ (.A(\g.g_y[3].g_x[7].t.out_sc ),
    .X(_0945_));
 sg13g2_buf_2 _4238_ (.A(\g.g_y[3].g_x[7].t.r_d ),
    .X(_0946_));
 sg13g2_mux2_1 _4239_ (.A0(\g.g_y[3].g_x[7].t.r_gnl ),
    .A1(_0945_),
    .S(_0946_),
    .X(_0947_));
 sg13g2_buf_1 _4240_ (.A(\g.g_y[3].g_x[7].t.r_ghl ),
    .X(_0948_));
 sg13g2_nand2b_1 _4241_ (.Y(_0949_),
    .B(_0944_),
    .A_N(_0948_));
 sg13g2_o21ai_1 _4242_ (.B1(_0949_),
    .Y(_0950_),
    .A1(_0944_),
    .A2(_0947_));
 sg13g2_mux2_1 _4243_ (.A0(net153),
    .A1(_0938_),
    .S(_0950_),
    .X(_0951_));
 sg13g2_o21ai_1 _4244_ (.B1(_0951_),
    .Y(_0952_),
    .A1(_0942_),
    .A2(_0943_));
 sg13g2_and4_1 _4245_ (.A(_0932_),
    .B(_0935_),
    .C(_0941_),
    .D(_0952_),
    .X(_0953_));
 sg13g2_mux2_1 _4246_ (.A0(_0920_),
    .A1(_0953_),
    .S(net165),
    .X(_0954_));
 sg13g2_or4_1 _4247_ (.A(_0909_),
    .B(net128),
    .C(net56),
    .D(_0954_),
    .X(_0955_));
 sg13g2_nand3_1 _4248_ (.B(net160),
    .C(net56),
    .A(_0508_),
    .Y(_0956_));
 sg13g2_nand3_1 _4249_ (.B(_0955_),
    .C(_0956_),
    .A(_0918_),
    .Y(_0075_));
 sg13g2_mux2_1 _4250_ (.A0(_0916_),
    .A1(_0912_),
    .S(_0566_),
    .X(_0957_));
 sg13g2_mux2_1 _4251_ (.A0(_0953_),
    .A1(_0920_),
    .S(net165),
    .X(_0958_));
 sg13g2_nor2_1 _4252_ (.A(net56),
    .B(_0958_),
    .Y(_0959_));
 sg13g2_o21ai_1 _4253_ (.B1(net176),
    .Y(_0960_),
    .A1(\g.g_y[1].g_x[7].t.r_gnl ),
    .A2(net32));
 sg13g2_a21oi_1 _4254_ (.A1(_0957_),
    .A2(_0959_),
    .Y(_0076_),
    .B1(_0960_));
 sg13g2_nand2_1 _4255_ (.Y(_0961_),
    .A(_0504_),
    .B(net35));
 sg13g2_o21ai_1 _4256_ (.B1(_0566_),
    .Y(_0962_),
    .A1(net54),
    .A2(_0809_));
 sg13g2_a21oi_1 _4257_ (.A1(_0961_),
    .A2(_0962_),
    .Y(_0077_),
    .B1(net90));
 sg13g2_nand3_1 _4258_ (.B(net88),
    .C(_0917_),
    .A(_0505_),
    .Y(_0963_));
 sg13g2_or3_1 _4259_ (.A(_0505_),
    .B(_2715_),
    .C(_0954_),
    .X(_0964_));
 sg13g2_a22oi_1 _4260_ (.Y(_0965_),
    .B1(net96),
    .B2(_0587_),
    .A2(net55),
    .A1(_0504_));
 sg13g2_nand3_1 _4261_ (.B(_0964_),
    .C(_0965_),
    .A(_0963_),
    .Y(_0078_));
 sg13g2_nand2_1 _4262_ (.Y(_0966_),
    .A(_0504_),
    .B(net34));
 sg13g2_o21ai_1 _4263_ (.B1(_0509_),
    .Y(_0967_),
    .A1(net54),
    .A2(net86));
 sg13g2_buf_1 _4264_ (.A(net126),
    .X(_0968_));
 sg13g2_a21oi_1 _4265_ (.A1(_0966_),
    .A2(_0967_),
    .Y(_0079_),
    .B1(net85));
 sg13g2_mux2_1 _4266_ (.A0(_2670_),
    .A1(_2671_),
    .S(_0907_),
    .X(_0969_));
 sg13g2_and2_1 _4267_ (.A(net112),
    .B(_0969_),
    .X(_0080_));
 sg13g2_mux2_1 _4268_ (.A0(_2669_),
    .A1(_0635_),
    .S(_2677_),
    .X(_0970_));
 sg13g2_and2_1 _4269_ (.A(_2679_),
    .B(_0635_),
    .X(_0971_));
 sg13g2_a21oi_1 _4270_ (.A1(_2680_),
    .A2(_0971_),
    .Y(_0972_),
    .B1(_2683_));
 sg13g2_mux2_1 _4271_ (.A0(_0970_),
    .A1(_0972_),
    .S(_2663_),
    .X(_0973_));
 sg13g2_buf_1 _4272_ (.A(\g.g_y[3].g_x[0].t.r_v ),
    .X(_0974_));
 sg13g2_buf_1 _4273_ (.A(\g.g_y[3].g_x[0].t.r_h ),
    .X(_0975_));
 sg13g2_inv_1 _4274_ (.Y(_0976_),
    .A(_0975_));
 sg13g2_mux2_1 _4275_ (.A0(_0672_),
    .A1(\g.g_y[3].g_x[1].t.r_gnl ),
    .S(_0673_),
    .X(_0977_));
 sg13g2_buf_2 _4276_ (.A(\g.g_y[3].g_x[1].t.r_h ),
    .X(_0978_));
 sg13g2_mux2_1 _4277_ (.A0(_0977_),
    .A1(_0675_),
    .S(_0978_),
    .X(_0979_));
 sg13g2_buf_1 _4278_ (.A(_0979_),
    .X(_0980_));
 sg13g2_and2_1 _4279_ (.A(net4),
    .B(_0975_),
    .X(_0981_));
 sg13g2_a21oi_1 _4280_ (.A1(_0976_),
    .A2(_0980_),
    .Y(_0982_),
    .B1(_0981_));
 sg13g2_buf_1 _4281_ (.A(\g.g_y[3].g_x[0].t.r_d ),
    .X(_0983_));
 sg13g2_inv_1 _4282_ (.Y(_0984_),
    .A(_0983_));
 sg13g2_buf_2 _4283_ (.A(\g.g_y[4].g_x[0].t.out_sc ),
    .X(_0985_));
 sg13g2_buf_2 _4284_ (.A(\g.g_y[4].g_x[0].t.r_d ),
    .X(_0986_));
 sg13g2_mux2_1 _4285_ (.A0(\g.g_y[4].g_x[0].t.r_gnl ),
    .A1(_0985_),
    .S(_0986_),
    .X(_0987_));
 sg13g2_buf_1 _4286_ (.A(_0987_),
    .X(_0988_));
 sg13g2_buf_1 _4287_ (.A(\g.g_y[4].g_x[0].t.r_ghl ),
    .X(_0989_));
 sg13g2_buf_1 _4288_ (.A(\g.g_y[4].g_x[0].t.r_v ),
    .X(_0990_));
 sg13g2_mux2_1 _4289_ (.A0(_0988_),
    .A1(_0989_),
    .S(net151),
    .X(_0991_));
 sg13g2_nand2_1 _4290_ (.Y(_0992_),
    .A(_0984_),
    .B(_0991_));
 sg13g2_buf_2 _4291_ (.A(\g.g_y[3].g_x[0].t.out_sc ),
    .X(_0993_));
 sg13g2_nand2b_1 _4292_ (.Y(_0994_),
    .B(_0983_),
    .A_N(_0993_));
 sg13g2_o21ai_1 _4293_ (.B1(_0994_),
    .Y(_0995_),
    .A1(_0982_),
    .A2(_0992_));
 sg13g2_buf_1 _4294_ (.A(_0983_),
    .X(_0996_));
 sg13g2_mux2_1 _4295_ (.A0(net4),
    .A1(_0980_),
    .S(_0975_),
    .X(_0997_));
 sg13g2_nand2b_1 _4296_ (.Y(_0998_),
    .B(net151),
    .A_N(_0989_));
 sg13g2_o21ai_1 _4297_ (.B1(_0998_),
    .Y(_0999_),
    .A1(_0990_),
    .A2(_0988_));
 sg13g2_inv_1 _4298_ (.Y(_1000_),
    .A(_0974_));
 sg13g2_a21oi_1 _4299_ (.A1(_0996_),
    .A2(_0999_),
    .Y(_1001_),
    .B1(_1000_));
 sg13g2_o21ai_1 _4300_ (.B1(_1001_),
    .Y(_1002_),
    .A1(net111),
    .A2(_0997_));
 sg13g2_o21ai_1 _4301_ (.B1(_1002_),
    .Y(_1003_),
    .A1(_0974_),
    .A2(_0995_));
 sg13g2_mux2_1 _4302_ (.A0(_0973_),
    .A1(_1003_),
    .S(_2674_),
    .X(_1004_));
 sg13g2_mux2_1 _4303_ (.A0(_0674_),
    .A1(_0675_),
    .S(_0671_),
    .X(_1005_));
 sg13g2_nor2b_1 _4304_ (.A(_2612_),
    .B_N(_2611_),
    .Y(_1006_));
 sg13g2_a21o_1 _4305_ (.A2(_2610_),
    .A1(_2612_),
    .B1(_1006_),
    .X(_1007_));
 sg13g2_mux2_1 _4306_ (.A0(_1005_),
    .A1(_1007_),
    .S(_0698_),
    .X(_1008_));
 sg13g2_nand3_1 _4307_ (.B(_0689_),
    .C(_1008_),
    .A(net114),
    .Y(_1009_));
 sg13g2_nor2_1 _4308_ (.A(_0682_),
    .B(_0691_),
    .Y(_1010_));
 sg13g2_nor2_1 _4309_ (.A(_0683_),
    .B(_1010_),
    .Y(_1011_));
 sg13g2_a21oi_1 _4310_ (.A1(_2612_),
    .A2(_2610_),
    .Y(_1012_),
    .B1(_1006_));
 sg13g2_inv_1 _4311_ (.Y(_1013_),
    .A(_0698_));
 sg13g2_mux2_1 _4312_ (.A0(_0677_),
    .A1(_1012_),
    .S(_1013_),
    .X(_1014_));
 sg13g2_nand2_1 _4313_ (.Y(_1015_),
    .A(_0694_),
    .B(_1014_));
 sg13g2_o21ai_1 _4314_ (.B1(_0683_),
    .Y(_1016_),
    .A1(net114),
    .A2(_0689_));
 sg13g2_inv_1 _4315_ (.Y(_1017_),
    .A(_1016_));
 sg13g2_a22oi_1 _4316_ (.Y(_1018_),
    .B1(_1015_),
    .B2(_1017_),
    .A2(_1011_),
    .A1(_1009_));
 sg13g2_nand2_1 _4317_ (.Y(_1019_),
    .A(net161),
    .B(_1018_));
 sg13g2_nor2_1 _4318_ (.A(net161),
    .B(net3),
    .Y(_1020_));
 sg13g2_nor2_1 _4319_ (.A(_2671_),
    .B(_1020_),
    .Y(_1021_));
 sg13g2_a22oi_1 _4320_ (.Y(_1022_),
    .B1(_1019_),
    .B2(_1021_),
    .A2(_1004_),
    .A1(_2671_));
 sg13g2_o21ai_1 _4321_ (.B1(net176),
    .Y(_1023_),
    .A1(_2673_),
    .A2(net59));
 sg13g2_a21oi_1 _4322_ (.A1(net60),
    .A2(_1022_),
    .Y(_0081_),
    .B1(_1023_));
 sg13g2_nand2_1 _4323_ (.Y(_1024_),
    .A(net161),
    .B(net3));
 sg13g2_or2_1 _4324_ (.X(_1025_),
    .B(_1018_),
    .A(_0679_));
 sg13g2_nand2_1 _4325_ (.Y(_1026_),
    .A(_2674_),
    .B(_0973_));
 sg13g2_nand2b_1 _4326_ (.Y(_1027_),
    .B(_1003_),
    .A_N(_2674_));
 sg13g2_a22oi_1 _4327_ (.Y(_1028_),
    .B1(_1026_),
    .B2(_1027_),
    .A2(_1025_),
    .A1(_1024_));
 sg13g2_buf_1 _4328_ (.A(net184),
    .X(_1029_));
 sg13g2_o21ai_1 _4329_ (.B1(_1029_),
    .Y(_1030_),
    .A1(\g.g_y[2].g_x[0].t.r_gnl ),
    .A2(net59));
 sg13g2_a21oi_1 _4330_ (.A1(net60),
    .A2(_1028_),
    .Y(_0082_),
    .B1(_1030_));
 sg13g2_nand2_1 _4331_ (.Y(_1031_),
    .A(_2670_),
    .B(_0807_));
 sg13g2_o21ai_1 _4332_ (.B1(net161),
    .Y(_1032_),
    .A1(net54),
    .A2(_0809_));
 sg13g2_a21oi_1 _4333_ (.A1(_1031_),
    .A2(_1032_),
    .Y(_0083_),
    .B1(_0968_));
 sg13g2_nand2b_1 _4334_ (.Y(_1033_),
    .B(_1004_),
    .A_N(_2671_));
 sg13g2_a21oi_1 _4335_ (.A1(_0679_),
    .A2(_1018_),
    .Y(_1034_),
    .B1(_1020_));
 sg13g2_a221oi_1 _4336_ (.B2(_2671_),
    .C1(net120),
    .B1(_1034_),
    .A1(_2670_),
    .Y(_1035_),
    .A2(_2719_));
 sg13g2_nor2_1 _4337_ (.A(net124),
    .B(_0504_),
    .Y(_1036_));
 sg13g2_buf_1 _4338_ (.A(net175),
    .X(_1037_));
 sg13g2_o21ai_1 _4339_ (.B1(net160),
    .Y(_1038_),
    .A1(_2670_),
    .A2(net110));
 sg13g2_a221oi_1 _4340_ (.B2(net125),
    .C1(_1038_),
    .B1(_1036_),
    .A1(_1033_),
    .Y(_0084_),
    .A2(_1035_));
 sg13g2_nand2_1 _4341_ (.Y(_1039_),
    .A(_2670_),
    .B(net34));
 sg13g2_o21ai_1 _4342_ (.B1(_2674_),
    .Y(_1040_),
    .A1(net54),
    .A2(net86));
 sg13g2_a21oi_1 _4343_ (.A1(_1039_),
    .A2(_1040_),
    .Y(_0085_),
    .B1(net85));
 sg13g2_mux2_1 _4344_ (.A0(_0691_),
    .A1(net114),
    .S(net33),
    .X(_1041_));
 sg13g2_and2_1 _4345_ (.A(_0906_),
    .B(_1041_),
    .X(_0086_));
 sg13g2_nand2_1 _4346_ (.Y(_1042_),
    .A(_0691_),
    .B(net35));
 sg13g2_o21ai_1 _4347_ (.B1(_0683_),
    .Y(_1043_),
    .A1(net54),
    .A2(net89));
 sg13g2_a21oi_1 _4348_ (.A1(_1042_),
    .A2(_1043_),
    .Y(_0087_),
    .B1(net85));
 sg13g2_or2_1 _4349_ (.X(_1044_),
    .B(net123),
    .A(_0691_));
 sg13g2_inv_1 _4350_ (.Y(_1045_),
    .A(_0694_));
 sg13g2_nor2_1 _4351_ (.A(_1045_),
    .B(_0695_),
    .Y(_1046_));
 sg13g2_and2_1 _4352_ (.A(_1045_),
    .B(_1014_),
    .X(_1047_));
 sg13g2_nor3_1 _4353_ (.A(net169),
    .B(_1046_),
    .C(_1047_),
    .Y(_1048_));
 sg13g2_buf_1 _4354_ (.A(net175),
    .X(_1049_));
 sg13g2_nand2_1 _4355_ (.Y(_1050_),
    .A(net116),
    .B(_2670_));
 sg13g2_nand3b_1 _4356_ (.B(net109),
    .C(_1050_),
    .Y(_1051_),
    .A_N(_1048_));
 sg13g2_and3_1 _4357_ (.X(_0088_),
    .A(net117),
    .B(_1044_),
    .C(_1051_));
 sg13g2_nand2_1 _4358_ (.Y(_1052_),
    .A(_0691_),
    .B(_0889_));
 sg13g2_buf_1 _4359_ (.A(net99),
    .X(_1053_));
 sg13g2_o21ai_1 _4360_ (.B1(_0698_),
    .Y(_1054_),
    .A1(net53),
    .A2(net86));
 sg13g2_a21oi_1 _4361_ (.A1(_1052_),
    .A2(_1054_),
    .Y(_0089_),
    .B1(net85));
 sg13g2_mux2_1 _4362_ (.A0(_2838_),
    .A1(_2839_),
    .S(net33),
    .X(_1055_));
 sg13g2_and2_1 _4363_ (.A(net112),
    .B(_1055_),
    .X(_0090_));
 sg13g2_and2_1 _4364_ (.A(_0682_),
    .B(_0681_),
    .X(_1056_));
 sg13g2_a21oi_1 _4365_ (.A1(_1008_),
    .A2(_1056_),
    .Y(_1057_),
    .B1(_1010_));
 sg13g2_nor2_1 _4366_ (.A(net114),
    .B(_0681_),
    .Y(_1058_));
 sg13g2_nor2_1 _4367_ (.A(_0683_),
    .B(_1058_),
    .Y(_1059_));
 sg13g2_a22oi_1 _4368_ (.Y(_1060_),
    .B1(_1059_),
    .B2(_1015_),
    .A2(_1057_),
    .A1(_0683_));
 sg13g2_nor2b_1 _4369_ (.A(_2771_),
    .B_N(_2770_),
    .Y(_1061_));
 sg13g2_a21o_1 _4370_ (.A2(_2769_),
    .A1(net113),
    .B1(_1061_),
    .X(_1062_));
 sg13g2_mux2_1 _4371_ (.A0(_0764_),
    .A1(_1062_),
    .S(_0756_),
    .X(_1063_));
 sg13g2_nor2_1 _4372_ (.A(_0766_),
    .B(_0773_),
    .Y(_1064_));
 sg13g2_nor2_1 _4373_ (.A(net159),
    .B(_0767_),
    .Y(_1065_));
 sg13g2_a21oi_1 _4374_ (.A1(_1063_),
    .A2(_1064_),
    .Y(_1066_),
    .B1(_1065_));
 sg13g2_nand2b_1 _4375_ (.Y(_1067_),
    .B(_0762_),
    .A_N(_0758_));
 sg13g2_o21ai_1 _4376_ (.B1(_1067_),
    .Y(_1068_),
    .A1(_0762_),
    .A2(_0761_));
 sg13g2_a21oi_1 _4377_ (.A1(net113),
    .A2(_2769_),
    .Y(_1069_),
    .B1(_1061_));
 sg13g2_mux2_1 _4378_ (.A0(_1068_),
    .A1(_1069_),
    .S(_0757_),
    .X(_1070_));
 sg13g2_nand2_1 _4379_ (.Y(_1071_),
    .A(net159),
    .B(_1070_));
 sg13g2_a21oi_1 _4380_ (.A1(_0766_),
    .A2(_0773_),
    .Y(_1072_),
    .B1(_0748_));
 sg13g2_a22oi_1 _4381_ (.Y(_1073_),
    .B1(_1071_),
    .B2(_1072_),
    .A2(_1066_),
    .A1(_0748_));
 sg13g2_mux2_1 _4382_ (.A0(_1060_),
    .A1(_1073_),
    .S(_0687_),
    .X(_1074_));
 sg13g2_a21oi_1 _4383_ (.A1(net122),
    .A2(_2859_),
    .Y(_1075_),
    .B1(_2845_));
 sg13g2_a21oi_1 _4384_ (.A1(net122),
    .A2(_0660_),
    .Y(_1076_),
    .B1(_2844_));
 sg13g2_a22oi_1 _4385_ (.Y(_1077_),
    .B1(_1076_),
    .B2(_2866_),
    .A2(_1075_),
    .A1(_2856_));
 sg13g2_buf_1 _4386_ (.A(\g.g_y[3].g_x[2].t.r_d ),
    .X(_1078_));
 sg13g2_inv_1 _4387_ (.Y(_1079_),
    .A(net149));
 sg13g2_mux2_1 _4388_ (.A0(_2841_),
    .A1(_2840_),
    .S(_2842_),
    .X(_1080_));
 sg13g2_buf_2 _4389_ (.A(\g.g_y[4].g_x[2].t.out_sc ),
    .X(_1081_));
 sg13g2_buf_2 _4390_ (.A(\g.g_y[4].g_x[2].t.r_d ),
    .X(_1082_));
 sg13g2_mux2_1 _4391_ (.A0(\g.g_y[4].g_x[2].t.r_gnl ),
    .A1(_1081_),
    .S(_1082_),
    .X(_1083_));
 sg13g2_buf_1 _4392_ (.A(\g.g_y[4].g_x[2].t.r_ghl ),
    .X(_1084_));
 sg13g2_buf_2 _4393_ (.A(\g.g_y[4].g_x[2].t.r_v ),
    .X(_1085_));
 sg13g2_mux2_1 _4394_ (.A0(_1083_),
    .A1(_1084_),
    .S(_1085_),
    .X(_1086_));
 sg13g2_buf_1 _4395_ (.A(\g.g_y[3].g_x[2].t.r_v ),
    .X(_1087_));
 sg13g2_inv_1 _4396_ (.Y(_1088_),
    .A(_1087_));
 sg13g2_mux2_1 _4397_ (.A0(_1080_),
    .A1(_1086_),
    .S(_1088_),
    .X(_1089_));
 sg13g2_nor2b_1 _4398_ (.A(_0978_),
    .B_N(_0675_),
    .Y(_1090_));
 sg13g2_a21o_1 _4399_ (.A2(_0977_),
    .A1(_0978_),
    .B1(_1090_),
    .X(_1091_));
 sg13g2_mux2_1 _4400_ (.A0(_0759_),
    .A1(\g.g_y[3].g_x[3].t.r_gnl ),
    .S(_0760_),
    .X(_1092_));
 sg13g2_buf_1 _4401_ (.A(_1092_),
    .X(_1093_));
 sg13g2_buf_2 _4402_ (.A(\g.g_y[3].g_x[3].t.r_h ),
    .X(_1094_));
 sg13g2_inv_1 _4403_ (.Y(_1095_),
    .A(_1094_));
 sg13g2_mux2_1 _4404_ (.A0(_0758_),
    .A1(_1093_),
    .S(_1095_),
    .X(_1096_));
 sg13g2_buf_2 _4405_ (.A(\g.g_y[3].g_x[2].t.r_h ),
    .X(_1097_));
 sg13g2_inv_1 _4406_ (.Y(_1098_),
    .A(_1097_));
 sg13g2_mux2_1 _4407_ (.A0(_1091_),
    .A1(_1096_),
    .S(_1098_),
    .X(_1099_));
 sg13g2_nand3_1 _4408_ (.B(_1089_),
    .C(_1099_),
    .A(_1079_),
    .Y(_1100_));
 sg13g2_inv_2 _4409_ (.Y(_1101_),
    .A(\g.g_y[3].g_x[2].t.out_sc ));
 sg13g2_a21oi_1 _4410_ (.A1(net149),
    .A2(_1101_),
    .Y(_1102_),
    .B1(_1087_));
 sg13g2_a21oi_1 _4411_ (.A1(_0978_),
    .A2(_0977_),
    .Y(_1103_),
    .B1(_1090_));
 sg13g2_nand2b_1 _4412_ (.Y(_1104_),
    .B(_1094_),
    .A_N(_0758_));
 sg13g2_o21ai_1 _4413_ (.B1(_1104_),
    .Y(_1105_),
    .A1(_1094_),
    .A2(_1093_));
 sg13g2_mux2_1 _4414_ (.A0(_1103_),
    .A1(_1105_),
    .S(_1097_),
    .X(_1106_));
 sg13g2_o21ai_1 _4415_ (.B1(_1087_),
    .Y(_1107_),
    .A1(_1079_),
    .A2(_1086_));
 sg13g2_a21oi_1 _4416_ (.A1(_1079_),
    .A2(_1106_),
    .Y(_1108_),
    .B1(_1107_));
 sg13g2_a21oi_1 _4417_ (.A1(_1100_),
    .A2(_1102_),
    .Y(_1109_),
    .B1(_1108_));
 sg13g2_mux2_1 _4418_ (.A0(_1077_),
    .A1(_1109_),
    .S(_2842_),
    .X(_1110_));
 sg13g2_mux2_1 _4419_ (.A0(_1074_),
    .A1(_1110_),
    .S(_2839_),
    .X(_1111_));
 sg13g2_o21ai_1 _4420_ (.B1(net150),
    .Y(_1112_),
    .A1(_2841_),
    .A2(net45));
 sg13g2_a21oi_1 _4421_ (.A1(net46),
    .A2(_1111_),
    .Y(_0091_),
    .B1(_1112_));
 sg13g2_mux2_1 _4422_ (.A0(_1109_),
    .A1(_1077_),
    .S(_2842_),
    .X(_1113_));
 sg13g2_mux2_1 _4423_ (.A0(_1073_),
    .A1(_1060_),
    .S(_0687_),
    .X(_1114_));
 sg13g2_nor3_1 _4424_ (.A(_0457_),
    .B(_1113_),
    .C(_1114_),
    .Y(_1115_));
 sg13g2_o21ai_1 _4425_ (.B1(net117),
    .Y(_1116_),
    .A1(\g.g_y[2].g_x[2].t.r_gnl ),
    .A2(net45));
 sg13g2_nor2_1 _4426_ (.A(_1115_),
    .B(_1116_),
    .Y(_0092_));
 sg13g2_nand2_1 _4427_ (.Y(_1117_),
    .A(_2838_),
    .B(net35));
 sg13g2_o21ai_1 _4428_ (.B1(_0687_),
    .Y(_1118_),
    .A1(net53),
    .A2(net89));
 sg13g2_a21oi_1 _4429_ (.A1(_1117_),
    .A2(_1118_),
    .Y(_0093_),
    .B1(net85));
 sg13g2_mux2_1 _4430_ (.A0(_1110_),
    .A1(_1074_),
    .S(_2839_),
    .X(_1119_));
 sg13g2_a22oi_1 _4431_ (.Y(_1120_),
    .B1(net62),
    .B2(_0691_),
    .A2(net63),
    .A1(_2838_));
 sg13g2_o21ai_1 _4432_ (.B1(_1120_),
    .Y(_0094_),
    .A1(net64),
    .A2(_1119_));
 sg13g2_nand2_1 _4433_ (.Y(_1121_),
    .A(_2838_),
    .B(_0889_));
 sg13g2_o21ai_1 _4434_ (.B1(_2842_),
    .Y(_1122_),
    .A1(net53),
    .A2(_0891_));
 sg13g2_a21oi_1 _4435_ (.A1(_1121_),
    .A2(_1122_),
    .Y(_0095_),
    .B1(_0968_));
 sg13g2_mux2_1 _4436_ (.A0(_0767_),
    .A1(_0749_),
    .S(net33),
    .X(_1123_));
 sg13g2_and2_1 _4437_ (.A(net112),
    .B(_1123_),
    .X(_0096_));
 sg13g2_nand2_1 _4438_ (.Y(_1124_),
    .A(_0767_),
    .B(net35));
 sg13g2_o21ai_1 _4439_ (.B1(_0747_),
    .Y(_1125_),
    .A1(net53),
    .A2(net89));
 sg13g2_a21oi_1 _4440_ (.A1(_1124_),
    .A2(_1125_),
    .Y(_0097_),
    .B1(net85));
 sg13g2_mux2_1 _4441_ (.A0(_0774_),
    .A1(_1070_),
    .S(_0766_),
    .X(_1126_));
 sg13g2_buf_1 _4442_ (.A(net183),
    .X(_1127_));
 sg13g2_nand2_1 _4443_ (.Y(_1128_),
    .A(net148),
    .B(_2838_));
 sg13g2_o21ai_1 _4444_ (.B1(_1128_),
    .Y(_1129_),
    .A1(net116),
    .A2(_1126_));
 sg13g2_nor2b_1 _4445_ (.A(net123),
    .B_N(_0767_),
    .Y(_1130_));
 sg13g2_a21oi_1 _4446_ (.A1(net125),
    .A2(_1129_),
    .Y(_1131_),
    .B1(_1130_));
 sg13g2_nor2_1 _4447_ (.A(net87),
    .B(_1131_),
    .Y(_0098_));
 sg13g2_nand2_1 _4448_ (.Y(_1132_),
    .A(_0767_),
    .B(net34));
 sg13g2_o21ai_1 _4449_ (.B1(_0756_),
    .Y(_1133_),
    .A1(net53),
    .A2(net86));
 sg13g2_a21oi_1 _4450_ (.A1(_1132_),
    .A2(_1133_),
    .Y(_0099_),
    .B1(net85));
 sg13g2_mux2_1 _4451_ (.A0(_0430_),
    .A1(_0431_),
    .S(net33),
    .X(_1134_));
 sg13g2_and2_1 _4452_ (.A(net112),
    .B(_1134_),
    .X(_0100_));
 sg13g2_inv_1 _4453_ (.Y(_1135_),
    .A(\g.g_y[2].g_x[6].t.r_h ));
 sg13g2_mux2_1 _4454_ (.A0(_0575_),
    .A1(_0848_),
    .S(_1135_),
    .X(_1136_));
 sg13g2_mux2_1 _4455_ (.A0(_0860_),
    .A1(_1136_),
    .S(_0842_),
    .X(_1137_));
 sg13g2_mux2_1 _4456_ (.A0(_0340_),
    .A1(_0339_),
    .S(_0335_),
    .X(_1138_));
 sg13g2_mux2_1 _4457_ (.A0(_0865_),
    .A1(_1138_),
    .S(net157),
    .X(_1139_));
 sg13g2_nand3_1 _4458_ (.B(_1137_),
    .C(_1139_),
    .A(_0843_),
    .Y(_1140_));
 sg13g2_nor2_1 _4459_ (.A(net158),
    .B(_0862_),
    .Y(_1141_));
 sg13g2_nor2_1 _4460_ (.A(_0841_),
    .B(_1141_),
    .Y(_1142_));
 sg13g2_inv_1 _4461_ (.Y(_1143_),
    .A(net158));
 sg13g2_nand2b_1 _4462_ (.Y(_1144_),
    .B(_1135_),
    .A_N(_0848_));
 sg13g2_and2_1 _4463_ (.A(_0841_),
    .B(_0849_),
    .X(_1145_));
 sg13g2_a22oi_1 _4464_ (.Y(_1146_),
    .B1(_1144_),
    .B2(_1145_),
    .A2(_0860_),
    .A1(_0842_));
 sg13g2_or2_1 _4465_ (.X(_1147_),
    .B(_0339_),
    .A(_0370_));
 sg13g2_inv_1 _4466_ (.Y(_1148_),
    .A(_0340_));
 sg13g2_a21oi_1 _4467_ (.A1(_1148_),
    .A2(_0370_),
    .Y(_1149_),
    .B1(\g.g_y[2].g_x[5].t.r_v ));
 sg13g2_a221oi_1 _4468_ (.B2(_1149_),
    .C1(_1143_),
    .B1(_1147_),
    .A1(net157),
    .Y(_1150_),
    .A2(_0865_));
 sg13g2_a21oi_1 _4469_ (.A1(_1143_),
    .A2(_1146_),
    .Y(_1151_),
    .B1(_1150_));
 sg13g2_a22oi_1 _4470_ (.Y(_1152_),
    .B1(_1151_),
    .B2(_0841_),
    .A2(_1142_),
    .A1(_1140_));
 sg13g2_nand3_1 _4471_ (.B(_0746_),
    .C(_1063_),
    .A(net159),
    .Y(_1153_));
 sg13g2_nor2_1 _4472_ (.A(_0748_),
    .B(_1065_),
    .Y(_1154_));
 sg13g2_a21oi_1 _4473_ (.A1(_0766_),
    .A2(_0771_),
    .Y(_1155_),
    .B1(_0747_));
 sg13g2_a221oi_1 _4474_ (.B2(_1071_),
    .C1(_0753_),
    .B1(_1155_),
    .A1(_1153_),
    .Y(_1156_),
    .A2(_1154_));
 sg13g2_a21oi_1 _4475_ (.A1(_0753_),
    .A2(_1152_),
    .Y(_1157_),
    .B1(_1156_));
 sg13g2_nor3_1 _4476_ (.A(_0431_),
    .B(_2709_),
    .C(_0596_),
    .Y(_1158_));
 sg13g2_and3_1 _4477_ (.X(_1159_),
    .A(_0431_),
    .B(net184),
    .C(_2753_));
 sg13g2_inv_1 _4478_ (.Y(_1160_),
    .A(\g.g_y[3].g_x[4].t.r_d ));
 sg13g2_mux2_1 _4479_ (.A0(_0758_),
    .A1(_1093_),
    .S(_1094_),
    .X(_1161_));
 sg13g2_mux2_1 _4480_ (.A0(_0852_),
    .A1(\g.g_y[3].g_x[5].t.r_gnl ),
    .S(_0853_),
    .X(_1162_));
 sg13g2_buf_2 _4481_ (.A(\g.g_y[3].g_x[5].t.r_h ),
    .X(_1163_));
 sg13g2_mux2_1 _4482_ (.A0(_1162_),
    .A1(_0855_),
    .S(_1163_),
    .X(_1164_));
 sg13g2_buf_1 _4483_ (.A(_1164_),
    .X(_1165_));
 sg13g2_buf_2 _4484_ (.A(\g.g_y[3].g_x[4].t.r_h ),
    .X(_1166_));
 sg13g2_inv_1 _4485_ (.Y(_1167_),
    .A(_1166_));
 sg13g2_mux2_1 _4486_ (.A0(_1161_),
    .A1(_1165_),
    .S(_1167_),
    .X(_1168_));
 sg13g2_buf_8 _4487_ (.A(\g.g_y[4].g_x[4].t.r_ghl ),
    .X(_1169_));
 sg13g2_buf_8 _4488_ (.A(\g.g_y[4].g_x[4].t.out_sc ),
    .X(_1170_));
 sg13g2_buf_8 _4489_ (.A(\g.g_y[4].g_x[4].t.r_d ),
    .X(_1171_));
 sg13g2_mux2_1 _4490_ (.A0(\g.g_y[4].g_x[4].t.r_gnl ),
    .A1(_1170_),
    .S(_1171_),
    .X(_1172_));
 sg13g2_buf_2 _4491_ (.A(\g.g_y[4].g_x[4].t.r_v ),
    .X(_1173_));
 sg13g2_inv_1 _4492_ (.Y(_1174_),
    .A(_1173_));
 sg13g2_mux2_1 _4493_ (.A0(_1169_),
    .A1(_1172_),
    .S(_1174_),
    .X(_1175_));
 sg13g2_mux2_1 _4494_ (.A0(_0429_),
    .A1(_0433_),
    .S(_0434_),
    .X(_1176_));
 sg13g2_buf_2 _4495_ (.A(\g.g_y[3].g_x[4].t.r_v ),
    .X(_1177_));
 sg13g2_mux2_1 _4496_ (.A0(_1175_),
    .A1(_1176_),
    .S(_1177_),
    .X(_1178_));
 sg13g2_nand3_1 _4497_ (.B(_1168_),
    .C(_1178_),
    .A(_1160_),
    .Y(_1179_));
 sg13g2_buf_1 _4498_ (.A(\g.g_y[3].g_x[4].t.r_d ),
    .X(_1180_));
 sg13g2_buf_1 _4499_ (.A(\g.g_y[3].g_x[4].t.out_sc ),
    .X(_1181_));
 sg13g2_inv_2 _4500_ (.Y(_1182_),
    .A(_1181_));
 sg13g2_a21oi_1 _4501_ (.A1(net147),
    .A2(_1182_),
    .Y(_1183_),
    .B1(_1177_));
 sg13g2_inv_1 _4502_ (.Y(_1184_),
    .A(_1175_));
 sg13g2_inv_1 _4503_ (.Y(_1185_),
    .A(_0758_));
 sg13g2_a21oi_1 _4504_ (.A1(_1185_),
    .A2(_1095_),
    .Y(_1186_),
    .B1(_1166_));
 sg13g2_or2_1 _4505_ (.X(_1187_),
    .B(_1093_),
    .A(_1095_));
 sg13g2_a221oi_1 _4506_ (.B2(_1187_),
    .C1(\g.g_y[3].g_x[4].t.r_d ),
    .B1(_1186_),
    .A1(_1166_),
    .Y(_1188_),
    .A2(_1165_));
 sg13g2_a21oi_1 _4507_ (.A1(net147),
    .A2(_1184_),
    .Y(_1189_),
    .B1(_1188_));
 sg13g2_a22oi_1 _4508_ (.Y(_1190_),
    .B1(_1189_),
    .B2(_1177_),
    .A2(_1183_),
    .A1(_1179_));
 sg13g2_o21ai_1 _4509_ (.B1(_0415_),
    .Y(_1191_),
    .A1(_0416_),
    .A2(_0428_));
 sg13g2_nand2_1 _4510_ (.Y(_1192_),
    .A(_0378_),
    .B(_0382_));
 sg13g2_o21ai_1 _4511_ (.B1(_1192_),
    .Y(_1193_),
    .A1(_0449_),
    .A2(_1191_));
 sg13g2_nand4_1 _4512_ (.B(_0416_),
    .C(_0425_),
    .A(_0378_),
    .Y(_1194_),
    .D(_0428_));
 sg13g2_nand3_1 _4513_ (.B(_1193_),
    .C(_1194_),
    .A(_0435_),
    .Y(_1195_));
 sg13g2_o21ai_1 _4514_ (.B1(_1195_),
    .Y(_1196_),
    .A1(_0435_),
    .A2(_1190_));
 sg13g2_a22oi_1 _4515_ (.Y(_1197_),
    .B1(_1159_),
    .B2(_1196_),
    .A2(_1158_),
    .A1(_1157_));
 sg13g2_nand3_1 _4516_ (.B(net160),
    .C(_0596_),
    .A(_0429_),
    .Y(_1198_));
 sg13g2_nand2_1 _4517_ (.Y(_0101_),
    .A(_1197_),
    .B(_1198_));
 sg13g2_a21oi_1 _4518_ (.A1(_1193_),
    .A2(_1194_),
    .Y(_1199_),
    .B1(_0435_));
 sg13g2_a21o_1 _4519_ (.A2(_1190_),
    .A1(_0435_),
    .B1(_1199_),
    .X(_1200_));
 sg13g2_a22oi_1 _4520_ (.Y(_1201_),
    .B1(_1155_),
    .B2(_1071_),
    .A2(_1154_),
    .A1(_1153_));
 sg13g2_mux2_1 _4521_ (.A0(_1152_),
    .A1(_1201_),
    .S(_0753_),
    .X(_1202_));
 sg13g2_nor3_1 _4522_ (.A(_0596_),
    .B(_1200_),
    .C(_1202_),
    .Y(_1203_));
 sg13g2_o21ai_1 _4523_ (.B1(net117),
    .Y(_1204_),
    .A1(\g.g_y[2].g_x[4].t.r_gnl ),
    .A2(net59));
 sg13g2_nor2_1 _4524_ (.A(_1203_),
    .B(_1204_),
    .Y(_0102_));
 sg13g2_nand2_1 _4525_ (.Y(_1205_),
    .A(_0430_),
    .B(net35));
 sg13g2_o21ai_1 _4526_ (.B1(_0753_),
    .Y(_1206_),
    .A1(net53),
    .A2(net89));
 sg13g2_a21oi_1 _4527_ (.A1(_1205_),
    .A2(_1206_),
    .Y(_0103_),
    .B1(net85));
 sg13g2_a22oi_1 _4528_ (.Y(_1207_),
    .B1(net62),
    .B2(_0767_),
    .A2(net63),
    .A1(_0430_));
 sg13g2_and2_1 _4529_ (.A(_0431_),
    .B(net88),
    .X(_1208_));
 sg13g2_nor2_1 _4530_ (.A(_0431_),
    .B(_2715_),
    .Y(_1209_));
 sg13g2_a22oi_1 _4531_ (.Y(_1210_),
    .B1(_1209_),
    .B2(_1196_),
    .A2(_1208_),
    .A1(_1157_));
 sg13g2_nand2_1 _4532_ (.Y(_0104_),
    .A(_1207_),
    .B(_1210_));
 sg13g2_nand2_1 _4533_ (.Y(_1211_),
    .A(_0430_),
    .B(net34));
 sg13g2_o21ai_1 _4534_ (.B1(_0434_),
    .Y(_1212_),
    .A1(_1053_),
    .A2(_0891_));
 sg13g2_buf_1 _4535_ (.A(net126),
    .X(_1213_));
 sg13g2_a21oi_1 _4536_ (.A1(_1211_),
    .A2(_1212_),
    .Y(_0105_),
    .B1(_1213_));
 sg13g2_mux2_1 _4537_ (.A0(net155),
    .A1(_0843_),
    .S(net33),
    .X(_1214_));
 sg13g2_and2_1 _4538_ (.A(net112),
    .B(_1214_),
    .X(_0106_));
 sg13g2_nand2_1 _4539_ (.Y(_1215_),
    .A(net155),
    .B(net35));
 sg13g2_o21ai_1 _4540_ (.B1(_0841_),
    .Y(_1216_),
    .A1(net53),
    .A2(net89));
 sg13g2_a21oi_1 _4541_ (.A1(_1215_),
    .A2(_1216_),
    .Y(_0107_),
    .B1(net84));
 sg13g2_a221oi_1 _4542_ (.B2(_1149_),
    .C1(net158),
    .B1(_1147_),
    .A1(net157),
    .Y(_1217_),
    .A2(_0865_));
 sg13g2_a21oi_1 _4543_ (.A1(net158),
    .A2(_1146_),
    .Y(_1218_),
    .B1(_1217_));
 sg13g2_and2_1 _4544_ (.A(net170),
    .B(_0430_),
    .X(_1219_));
 sg13g2_a21oi_1 _4545_ (.A1(net124),
    .A2(_1218_),
    .Y(_1220_),
    .B1(_1219_));
 sg13g2_nor2_1 _4546_ (.A(net155),
    .B(net123),
    .Y(_1221_));
 sg13g2_a21oi_1 _4547_ (.A1(net110),
    .A2(_1220_),
    .Y(_1222_),
    .B1(_1221_));
 sg13g2_and2_1 _4548_ (.A(net112),
    .B(_1222_),
    .X(_0108_));
 sg13g2_nand2_1 _4549_ (.Y(_1223_),
    .A(net155),
    .B(net34));
 sg13g2_o21ai_1 _4550_ (.B1(_0845_),
    .Y(_1224_),
    .A1(_1053_),
    .A2(net86));
 sg13g2_a21oi_1 _4551_ (.A1(_1223_),
    .A2(_1224_),
    .Y(_0109_),
    .B1(_1213_));
 sg13g2_mux2_1 _4552_ (.A0(_0572_),
    .A1(_0573_),
    .S(net33),
    .X(_1225_));
 sg13g2_and2_1 _4553_ (.A(net112),
    .B(_1225_),
    .X(_0110_));
 sg13g2_o21ai_1 _4554_ (.B1(_0842_),
    .Y(_1226_),
    .A1(net158),
    .A2(_0860_));
 sg13g2_nor2_1 _4555_ (.A(_1150_),
    .B(_1226_),
    .Y(_1227_));
 sg13g2_a21oi_1 _4556_ (.A1(_0841_),
    .A2(_1140_),
    .Y(_1228_),
    .B1(_1227_));
 sg13g2_nand2_1 _4557_ (.Y(_1229_),
    .A(net156),
    .B(_0923_));
 sg13g2_mux2_1 _4558_ (.A0(_0947_),
    .A1(_0948_),
    .S(_0944_),
    .X(_1230_));
 sg13g2_nor2b_1 _4559_ (.A(net165),
    .B_N(_0508_),
    .Y(_1231_));
 sg13g2_a21o_1 _4560_ (.A2(_0507_),
    .A1(net165),
    .B1(_1231_),
    .X(_1232_));
 sg13g2_mux2_1 _4561_ (.A0(_1230_),
    .A1(_1232_),
    .S(_0925_),
    .X(_1233_));
 sg13g2_nor2_1 _4562_ (.A(_0921_),
    .B(_0927_),
    .Y(_1234_));
 sg13g2_a21oi_1 _4563_ (.A1(net165),
    .A2(_0507_),
    .Y(_1235_),
    .B1(_1231_));
 sg13g2_mux2_1 _4564_ (.A0(_0950_),
    .A1(_1235_),
    .S(_0933_),
    .X(_1236_));
 sg13g2_buf_1 _4565_ (.A(_1236_),
    .X(_1237_));
 sg13g2_a22oi_1 _4566_ (.Y(_1238_),
    .B1(_1237_),
    .B2(_0921_),
    .A2(_1234_),
    .A1(_1233_));
 sg13g2_nor2_1 _4567_ (.A(_0846_),
    .B(net155),
    .Y(_1239_));
 sg13g2_a21o_1 _4568_ (.A2(net152),
    .A1(_0922_),
    .B1(net154),
    .X(_1240_));
 sg13g2_a21oi_1 _4569_ (.A1(_0921_),
    .A2(_0937_),
    .Y(_1241_),
    .B1(_1240_));
 sg13g2_a22oi_1 _4570_ (.Y(_1242_),
    .B1(_1241_),
    .B2(net156),
    .A2(_1239_),
    .A1(_0844_));
 sg13g2_o21ai_1 _4571_ (.B1(_1242_),
    .Y(_1243_),
    .A1(_1229_),
    .A2(_1238_));
 sg13g2_a21o_1 _4572_ (.A2(_1228_),
    .A1(_1135_),
    .B1(_1243_),
    .X(_1244_));
 sg13g2_mux4_1 _4573_ (.S0(_0580_),
    .A0(_0586_),
    .A1(_0582_),
    .A2(_0835_),
    .A3(_0588_),
    .S1(_0590_),
    .X(_1245_));
 sg13g2_buf_1 _4574_ (.A(\g.g_y[3].g_x[6].t.r_d ),
    .X(_1246_));
 sg13g2_mux2_1 _4575_ (.A0(_0945_),
    .A1(\g.g_y[3].g_x[7].t.r_gnl ),
    .S(_0946_),
    .X(_1247_));
 sg13g2_buf_2 _4576_ (.A(\g.g_y[3].g_x[7].t.r_h ),
    .X(_1248_));
 sg13g2_mux2_1 _4577_ (.A0(_1247_),
    .A1(_0948_),
    .S(_1248_),
    .X(_1249_));
 sg13g2_mux2_1 _4578_ (.A0(_0855_),
    .A1(_1162_),
    .S(_1163_),
    .X(_1250_));
 sg13g2_buf_2 _4579_ (.A(\g.g_y[3].g_x[6].t.r_h ),
    .X(_1251_));
 sg13g2_mux2_1 _4580_ (.A0(_1249_),
    .A1(_1250_),
    .S(_1251_),
    .X(_1252_));
 sg13g2_buf_2 _4581_ (.A(\g.g_y[4].g_x[6].t.out_sc ),
    .X(_1253_));
 sg13g2_buf_8 _4582_ (.A(\g.g_y[4].g_x[6].t.r_d ),
    .X(_1254_));
 sg13g2_mux2_1 _4583_ (.A0(\g.g_y[4].g_x[6].t.r_gnl ),
    .A1(_1253_),
    .S(_1254_),
    .X(_1255_));
 sg13g2_buf_1 _4584_ (.A(\g.g_y[4].g_x[6].t.r_ghl ),
    .X(_1256_));
 sg13g2_buf_2 _4585_ (.A(\g.g_y[4].g_x[6].t.r_v ),
    .X(_1257_));
 sg13g2_mux2_1 _4586_ (.A0(_1255_),
    .A1(_1256_),
    .S(_1257_),
    .X(_1258_));
 sg13g2_mux2_1 _4587_ (.A0(_0575_),
    .A1(_0574_),
    .S(_0576_),
    .X(_1259_));
 sg13g2_buf_1 _4588_ (.A(\g.g_y[3].g_x[6].t.r_v ),
    .X(_1260_));
 sg13g2_mux2_1 _4589_ (.A0(_1258_),
    .A1(_1259_),
    .S(_1260_),
    .X(_1261_));
 sg13g2_nand3b_1 _4590_ (.B(_1252_),
    .C(_1261_),
    .Y(_1262_),
    .A_N(net146));
 sg13g2_buf_2 _4591_ (.A(\g.g_y[3].g_x[6].t.out_sc ),
    .X(_1263_));
 sg13g2_inv_1 _4592_ (.Y(_1264_),
    .A(_1263_));
 sg13g2_a21oi_1 _4593_ (.A1(net146),
    .A2(_1264_),
    .Y(_1265_),
    .B1(_1260_));
 sg13g2_mux2_1 _4594_ (.A0(_1250_),
    .A1(_1249_),
    .S(_1251_),
    .X(_1266_));
 sg13g2_inv_1 _4595_ (.Y(_1267_),
    .A(_1260_));
 sg13g2_mux2_1 _4596_ (.A0(_1258_),
    .A1(_1259_),
    .S(_1267_),
    .X(_1268_));
 sg13g2_buf_1 _4597_ (.A(_1268_),
    .X(_1269_));
 sg13g2_mux2_1 _4598_ (.A0(_1266_),
    .A1(_1269_),
    .S(net146),
    .X(_1270_));
 sg13g2_a22oi_1 _4599_ (.Y(_1271_),
    .B1(_1270_),
    .B2(_1260_),
    .A2(_1265_),
    .A1(_1262_));
 sg13g2_mux2_1 _4600_ (.A0(_1245_),
    .A1(_1271_),
    .S(_0576_),
    .X(_1272_));
 sg13g2_mux2_1 _4601_ (.A0(_1244_),
    .A1(_1272_),
    .S(_0573_),
    .X(_1273_));
 sg13g2_o21ai_1 _4602_ (.B1(_1029_),
    .Y(_1274_),
    .A1(_0575_),
    .A2(net45));
 sg13g2_a21oi_1 _4603_ (.A1(net46),
    .A2(_1273_),
    .Y(_0111_),
    .B1(_1274_));
 sg13g2_o21ai_1 _4604_ (.B1(net177),
    .Y(_1275_),
    .A1(\g.g_y[2].g_x[6].t.r_gnl ),
    .A2(net45));
 sg13g2_mux2_1 _4605_ (.A0(_0937_),
    .A1(_0930_),
    .S(_0921_),
    .X(_1276_));
 sg13g2_a21oi_1 _4606_ (.A1(_1233_),
    .A2(_1276_),
    .Y(_1277_),
    .B1(_0938_));
 sg13g2_a21oi_1 _4607_ (.A1(_0938_),
    .A2(net152),
    .Y(_1278_),
    .B1(_1277_));
 sg13g2_o21ai_1 _4608_ (.B1(_0921_),
    .Y(_1279_),
    .A1(net154),
    .A2(_0937_));
 sg13g2_a21oi_1 _4609_ (.A1(net154),
    .A2(_1237_),
    .Y(_1280_),
    .B1(_1279_));
 sg13g2_nor2_1 _4610_ (.A(net156),
    .B(_1280_),
    .Y(_1281_));
 sg13g2_o21ai_1 _4611_ (.B1(_1281_),
    .Y(_1282_),
    .A1(_0921_),
    .A2(_1278_));
 sg13g2_nor2_1 _4612_ (.A(_0842_),
    .B(_1141_),
    .Y(_1283_));
 sg13g2_a21oi_1 _4613_ (.A1(_1140_),
    .A2(_1283_),
    .Y(_1284_),
    .B1(_1227_));
 sg13g2_nand2_1 _4614_ (.Y(_1285_),
    .A(net156),
    .B(_1284_));
 sg13g2_nand2b_1 _4615_ (.Y(_1286_),
    .B(_1271_),
    .A_N(_0576_));
 sg13g2_a21oi_1 _4616_ (.A1(_0576_),
    .A2(_1245_),
    .Y(_1287_),
    .B1(_0457_));
 sg13g2_nand4_1 _4617_ (.B(_1285_),
    .C(_1286_),
    .A(_1282_),
    .Y(_1288_),
    .D(_1287_));
 sg13g2_nor2b_1 _4618_ (.A(_1275_),
    .B_N(_1288_),
    .Y(_0112_));
 sg13g2_buf_1 _4619_ (.A(net66),
    .X(_1289_));
 sg13g2_nand2_1 _4620_ (.Y(_1290_),
    .A(_0572_),
    .B(net31));
 sg13g2_buf_1 _4621_ (.A(_2699_),
    .X(_1291_));
 sg13g2_o21ai_1 _4622_ (.B1(net156),
    .Y(_1292_),
    .A1(net53),
    .A2(net108));
 sg13g2_a21oi_1 _4623_ (.A1(_1290_),
    .A2(_1292_),
    .Y(_0113_),
    .B1(net84));
 sg13g2_mux2_1 _4624_ (.A0(_1272_),
    .A1(_1244_),
    .S(_0573_),
    .X(_1293_));
 sg13g2_a22oi_1 _4625_ (.Y(_1294_),
    .B1(net62),
    .B2(net155),
    .A2(net63),
    .A1(_0572_));
 sg13g2_o21ai_1 _4626_ (.B1(_1294_),
    .Y(_0114_),
    .A1(net64),
    .A2(_1293_));
 sg13g2_nand2_1 _4627_ (.Y(_1295_),
    .A(_0572_),
    .B(net34));
 sg13g2_buf_1 _4628_ (.A(net99),
    .X(_1296_));
 sg13g2_o21ai_1 _4629_ (.B1(_0576_),
    .Y(_1297_),
    .A1(net52),
    .A2(net86));
 sg13g2_a21oi_1 _4630_ (.A1(_1295_),
    .A2(_1297_),
    .Y(_0115_),
    .B1(net84));
 sg13g2_mux2_1 _4631_ (.A0(net152),
    .A1(_0923_),
    .S(net33),
    .X(_1298_));
 sg13g2_and2_1 _4632_ (.A(net112),
    .B(_1298_),
    .X(_0116_));
 sg13g2_nand2_1 _4633_ (.Y(_1299_),
    .A(net152),
    .B(net31));
 sg13g2_o21ai_1 _4634_ (.B1(_0921_),
    .Y(_1300_),
    .A1(net52),
    .A2(net108));
 sg13g2_a21oi_1 _4635_ (.A1(_1299_),
    .A2(_1300_),
    .Y(_0117_),
    .B1(net84));
 sg13g2_buf_1 _4636_ (.A(net181),
    .X(_1301_));
 sg13g2_nor2_1 _4637_ (.A(_0938_),
    .B(_0942_),
    .Y(_1302_));
 sg13g2_and2_1 _4638_ (.A(_0938_),
    .B(_1237_),
    .X(_1303_));
 sg13g2_o21ai_1 _4639_ (.B1(net124),
    .Y(_1304_),
    .A1(_1302_),
    .A2(_1303_));
 sg13g2_o21ai_1 _4640_ (.B1(_1304_),
    .Y(_1305_),
    .A1(net124),
    .A2(_0572_));
 sg13g2_nor2_1 _4641_ (.A(net152),
    .B(net175),
    .Y(_1306_));
 sg13g2_a21oi_1 _4642_ (.A1(net110),
    .A2(_1305_),
    .Y(_1307_),
    .B1(_1306_));
 sg13g2_and2_1 _4643_ (.A(net107),
    .B(_1307_),
    .X(_0118_));
 sg13g2_buf_1 _4644_ (.A(net61),
    .X(_1308_));
 sg13g2_nand2_1 _4645_ (.Y(_1309_),
    .A(net152),
    .B(net30));
 sg13g2_buf_1 _4646_ (.A(net127),
    .X(_1310_));
 sg13g2_o21ai_1 _4647_ (.B1(_0925_),
    .Y(_1311_),
    .A1(net52),
    .A2(net83));
 sg13g2_a21oi_1 _4648_ (.A1(_1309_),
    .A2(_1311_),
    .Y(_0119_),
    .B1(net84));
 sg13g2_mux2_1 _4649_ (.A0(_0993_),
    .A1(_0996_),
    .S(_0907_),
    .X(_1312_));
 sg13g2_and2_1 _4650_ (.A(net107),
    .B(_1312_),
    .X(_0120_));
 sg13g2_nand2_1 _4651_ (.Y(_1313_),
    .A(_0993_),
    .B(_1289_));
 sg13g2_o21ai_1 _4652_ (.B1(_0975_),
    .Y(_1314_),
    .A1(_1296_),
    .A2(_1291_));
 sg13g2_a21oi_1 _4653_ (.A1(_1313_),
    .A2(_1314_),
    .Y(_0121_),
    .B1(net84));
 sg13g2_nor2b_1 _4654_ (.A(_2674_),
    .B_N(_2673_),
    .Y(_1315_));
 sg13g2_a21oi_1 _4655_ (.A1(_2674_),
    .A2(_2672_),
    .Y(_1316_),
    .B1(_1315_));
 sg13g2_mux2_1 _4656_ (.A0(_0999_),
    .A1(_1316_),
    .S(_1000_),
    .X(_1317_));
 sg13g2_nor2_1 _4657_ (.A(_0984_),
    .B(_0997_),
    .Y(_1318_));
 sg13g2_a21oi_1 _4658_ (.A1(_0984_),
    .A2(_1317_),
    .Y(_1319_),
    .B1(_1318_));
 sg13g2_nand2b_1 _4659_ (.Y(_1320_),
    .B(net170),
    .A_N(net152));
 sg13g2_o21ai_1 _4660_ (.B1(_1320_),
    .Y(_1321_),
    .A1(net115),
    .A2(_1319_));
 sg13g2_nor2_1 _4661_ (.A(_0993_),
    .B(net175),
    .Y(_1322_));
 sg13g2_a21oi_1 _4662_ (.A1(_1037_),
    .A2(_1321_),
    .Y(_1323_),
    .B1(_1322_));
 sg13g2_and2_1 _4663_ (.A(net107),
    .B(_1323_),
    .X(_0122_));
 sg13g2_nand2_1 _4664_ (.Y(_1324_),
    .A(_0993_),
    .B(net30));
 sg13g2_o21ai_1 _4665_ (.B1(_0974_),
    .Y(_1325_),
    .A1(_1296_),
    .A2(net83));
 sg13g2_a21oi_1 _4666_ (.A1(_1324_),
    .A2(_1325_),
    .Y(_0123_),
    .B1(net84));
 sg13g2_buf_2 _4667_ (.A(_2592_),
    .X(_1326_));
 sg13g2_mux2_1 _4668_ (.A0(_0672_),
    .A1(_0673_),
    .S(_1326_),
    .X(_1327_));
 sg13g2_and2_1 _4669_ (.A(_1301_),
    .B(_1327_),
    .X(_0124_));
 sg13g2_inv_1 _4670_ (.Y(_1328_),
    .A(_0673_));
 sg13g2_a21o_1 _4671_ (.A2(_2672_),
    .A1(_2674_),
    .B1(_1315_),
    .X(_1329_));
 sg13g2_mux2_1 _4672_ (.A0(_0991_),
    .A1(_1329_),
    .S(_0974_),
    .X(_1330_));
 sg13g2_and2_1 _4673_ (.A(net4),
    .B(_0983_),
    .X(_1331_));
 sg13g2_nor2_1 _4674_ (.A(_0983_),
    .B(_0993_),
    .Y(_1332_));
 sg13g2_a21oi_1 _4675_ (.A1(_1330_),
    .A2(_1331_),
    .Y(_1333_),
    .B1(_1332_));
 sg13g2_nor2_1 _4676_ (.A(net4),
    .B(net111),
    .Y(_1334_));
 sg13g2_a21oi_1 _4677_ (.A1(net111),
    .A2(_1317_),
    .Y(_1335_),
    .B1(_1334_));
 sg13g2_mux2_1 _4678_ (.A0(_1333_),
    .A1(_1335_),
    .S(_0976_),
    .X(_1336_));
 sg13g2_nand2_1 _4679_ (.Y(_1337_),
    .A(_1089_),
    .B(_1099_));
 sg13g2_mux2_1 _4680_ (.A0(_1080_),
    .A1(_1086_),
    .S(_1087_),
    .X(_1338_));
 sg13g2_mux4_1 _4681_ (.S0(_1097_),
    .A0(\g.g_y[3].g_x[2].t.out_sc ),
    .A1(_1096_),
    .A2(_1337_),
    .A3(_1338_),
    .S1(net149),
    .X(_1339_));
 sg13g2_mux2_1 _4682_ (.A0(_1336_),
    .A1(_1339_),
    .S(_0978_),
    .X(_1340_));
 sg13g2_nand4_1 _4683_ (.B(net160),
    .C(_0743_),
    .A(_1328_),
    .Y(_1341_),
    .D(_1340_));
 sg13g2_o21ai_1 _4684_ (.B1(_0692_),
    .Y(_1342_),
    .A1(_0690_),
    .A2(_1012_));
 sg13g2_a21oi_1 _4685_ (.A1(net114),
    .A2(_1012_),
    .Y(_1343_),
    .B1(_0698_));
 sg13g2_o21ai_1 _4686_ (.B1(_1343_),
    .Y(_1344_),
    .A1(net114),
    .A2(_0695_));
 sg13g2_o21ai_1 _4687_ (.B1(_1344_),
    .Y(_1345_),
    .A1(_1013_),
    .A2(_1342_));
 sg13g2_buf_1 _4688_ (.A(\g.g_y[5].g_x[1].t.r_v ),
    .X(_1346_));
 sg13g2_buf_2 _4689_ (.A(\g.g_y[5].g_x[1].t.out_sc ),
    .X(_1347_));
 sg13g2_buf_8 _4690_ (.A(\g.g_y[5].g_x[1].t.r_d ),
    .X(_1348_));
 sg13g2_mux2_1 _4691_ (.A0(\g.g_y[5].g_x[1].t.r_gnl ),
    .A1(_1347_),
    .S(_1348_),
    .X(_1349_));
 sg13g2_buf_1 _4692_ (.A(\g.g_y[5].g_x[1].t.r_ghl ),
    .X(_1350_));
 sg13g2_nand2b_1 _4693_ (.Y(_1351_),
    .B(net145),
    .A_N(_1350_));
 sg13g2_o21ai_1 _4694_ (.B1(_1351_),
    .Y(_1352_),
    .A1(net145),
    .A2(_1349_));
 sg13g2_nor2b_1 _4695_ (.A(_0671_),
    .B_N(_0675_),
    .Y(_1353_));
 sg13g2_a21oi_1 _4696_ (.A1(_0671_),
    .A2(_0674_),
    .Y(_1354_),
    .B1(_1353_));
 sg13g2_buf_2 _4697_ (.A(\g.g_y[4].g_x[1].t.r_v ),
    .X(_1355_));
 sg13g2_mux2_1 _4698_ (.A0(_1352_),
    .A1(_1354_),
    .S(_1355_),
    .X(_1356_));
 sg13g2_buf_2 _4699_ (.A(\g.g_y[4].g_x[2].t.r_h ),
    .X(_1357_));
 sg13g2_mux2_1 _4700_ (.A0(_1081_),
    .A1(\g.g_y[4].g_x[2].t.r_gnl ),
    .S(_1082_),
    .X(_1358_));
 sg13g2_nand2b_1 _4701_ (.Y(_1359_),
    .B(_1357_),
    .A_N(_1084_));
 sg13g2_o21ai_1 _4702_ (.B1(_1359_),
    .Y(_1360_),
    .A1(_1357_),
    .A2(_1358_));
 sg13g2_buf_1 _4703_ (.A(\g.g_y[4].g_x[0].t.r_h ),
    .X(_1361_));
 sg13g2_mux2_1 _4704_ (.A0(_0985_),
    .A1(\g.g_y[4].g_x[0].t.r_gnl ),
    .S(_0986_),
    .X(_1362_));
 sg13g2_nor2b_1 _4705_ (.A(net144),
    .B_N(_0989_),
    .Y(_1363_));
 sg13g2_a21oi_1 _4706_ (.A1(net144),
    .A2(_1362_),
    .Y(_1364_),
    .B1(_1363_));
 sg13g2_buf_2 _4707_ (.A(\g.g_y[4].g_x[1].t.r_h ),
    .X(_1365_));
 sg13g2_mux2_1 _4708_ (.A0(_1360_),
    .A1(_1364_),
    .S(_1365_),
    .X(_1366_));
 sg13g2_nor2_1 _4709_ (.A(_1356_),
    .B(_1366_),
    .Y(_1367_));
 sg13g2_buf_1 _4710_ (.A(\g.g_y[4].g_x[1].t.r_d ),
    .X(_1368_));
 sg13g2_nor2_1 _4711_ (.A(_1355_),
    .B(net143),
    .Y(_1369_));
 sg13g2_nor2b_1 _4712_ (.A(net143),
    .B_N(_1355_),
    .Y(_1370_));
 sg13g2_mux2_1 _4713_ (.A0(_1364_),
    .A1(_1360_),
    .S(_1365_),
    .X(_1371_));
 sg13g2_buf_1 _4714_ (.A(_1371_),
    .X(_1372_));
 sg13g2_buf_1 _4715_ (.A(\g.g_y[4].g_x[1].t.out_sc ),
    .X(_1373_));
 sg13g2_inv_1 _4716_ (.Y(_1374_),
    .A(_1373_));
 sg13g2_nand2_1 _4717_ (.Y(_1375_),
    .A(_1368_),
    .B(_1374_));
 sg13g2_nand3_1 _4718_ (.B(net143),
    .C(_1352_),
    .A(_1355_),
    .Y(_1376_));
 sg13g2_o21ai_1 _4719_ (.B1(_1376_),
    .Y(_1377_),
    .A1(_1355_),
    .A2(_1375_));
 sg13g2_a221oi_1 _4720_ (.B2(_1372_),
    .C1(_1377_),
    .B1(_1370_),
    .A1(_1367_),
    .Y(_1378_),
    .A2(_1369_));
 sg13g2_mux2_1 _4721_ (.A0(_1345_),
    .A1(_1378_),
    .S(_0671_),
    .X(_1379_));
 sg13g2_nand4_1 _4722_ (.B(net181),
    .C(_0743_),
    .A(_0673_),
    .Y(_1380_),
    .D(_1379_));
 sg13g2_nand3_1 _4723_ (.B(net160),
    .C(net56),
    .A(_0675_),
    .Y(_1381_));
 sg13g2_nand3_1 _4724_ (.B(_1380_),
    .C(_1381_),
    .A(_1341_),
    .Y(_0125_));
 sg13g2_o21ai_1 _4725_ (.B1(net177),
    .Y(_1382_),
    .A1(\g.g_y[3].g_x[1].t.r_gnl ),
    .A2(net36));
 sg13g2_mux2_1 _4726_ (.A0(_1339_),
    .A1(_1336_),
    .S(_0978_),
    .X(_1383_));
 sg13g2_mux2_1 _4727_ (.A0(_1378_),
    .A1(_1345_),
    .S(_0671_),
    .X(_1384_));
 sg13g2_nand3_1 _4728_ (.B(_1383_),
    .C(_1384_),
    .A(net32),
    .Y(_1385_));
 sg13g2_nor2b_1 _4729_ (.A(_1382_),
    .B_N(_1385_),
    .Y(_0126_));
 sg13g2_nand2_1 _4730_ (.Y(_1386_),
    .A(_0672_),
    .B(_1289_));
 sg13g2_o21ai_1 _4731_ (.B1(_0978_),
    .Y(_1387_),
    .A1(net52),
    .A2(_1291_));
 sg13g2_a21oi_1 _4732_ (.A1(_1386_),
    .A2(_1387_),
    .Y(_0127_),
    .B1(net84));
 sg13g2_a22oi_1 _4733_ (.Y(_1388_),
    .B1(net96),
    .B2(_0993_),
    .A2(net55),
    .A1(_0672_));
 sg13g2_nand3_1 _4734_ (.B(net88),
    .C(_1340_),
    .A(_0673_),
    .Y(_1389_));
 sg13g2_nand3_1 _4735_ (.B(net88),
    .C(_1379_),
    .A(_1328_),
    .Y(_1390_));
 sg13g2_nand3_1 _4736_ (.B(_1389_),
    .C(_1390_),
    .A(_1388_),
    .Y(_0128_));
 sg13g2_nand2_1 _4737_ (.Y(_1391_),
    .A(_0672_),
    .B(_1308_));
 sg13g2_o21ai_1 _4738_ (.B1(_0671_),
    .Y(_1392_),
    .A1(net52),
    .A2(_1310_));
 sg13g2_buf_1 _4739_ (.A(net128),
    .X(_1393_));
 sg13g2_a21oi_1 _4740_ (.A1(_1391_),
    .A2(_1392_),
    .Y(_0129_),
    .B1(_1393_));
 sg13g2_buf_1 _4741_ (.A(_2592_),
    .X(_1394_));
 sg13g2_nor2_1 _4742_ (.A(_1101_),
    .B(net28),
    .Y(_1395_));
 sg13g2_a21oi_1 _4743_ (.A1(_1078_),
    .A2(net22),
    .Y(_1396_),
    .B1(_1395_));
 sg13g2_nor2_1 _4744_ (.A(net87),
    .B(_1396_),
    .Y(_0130_));
 sg13g2_mux2_1 _4745_ (.A0(_1098_),
    .A1(_1101_),
    .S(net66),
    .X(_1397_));
 sg13g2_nor2_1 _4746_ (.A(net87),
    .B(_1397_),
    .Y(_0131_));
 sg13g2_nand2_1 _4747_ (.Y(_1398_),
    .A(net149),
    .B(_1106_));
 sg13g2_o21ai_1 _4748_ (.B1(_1398_),
    .Y(_1399_),
    .A1(net149),
    .A2(_1338_));
 sg13g2_nand2_1 _4749_ (.Y(_1400_),
    .A(net148),
    .B(_0672_));
 sg13g2_o21ai_1 _4750_ (.B1(_1400_),
    .Y(_1401_),
    .A1(net116),
    .A2(_1399_));
 sg13g2_nor2_1 _4751_ (.A(_1101_),
    .B(net123),
    .Y(_1402_));
 sg13g2_a21oi_1 _4752_ (.A1(net125),
    .A2(_1401_),
    .Y(_1403_),
    .B1(_1402_));
 sg13g2_nor2_1 _4753_ (.A(net87),
    .B(_1403_),
    .Y(_0132_));
 sg13g2_mux2_1 _4754_ (.A0(_1088_),
    .A1(_1101_),
    .S(net40),
    .X(_1404_));
 sg13g2_nor2_1 _4755_ (.A(net87),
    .B(_1404_),
    .Y(_0133_));
 sg13g2_mux2_1 _4756_ (.A0(_0759_),
    .A1(_0760_),
    .S(net29),
    .X(_1405_));
 sg13g2_and2_1 _4757_ (.A(net107),
    .B(_1405_),
    .X(_0134_));
 sg13g2_nand3_1 _4758_ (.B(_1089_),
    .C(_1099_),
    .A(net149),
    .Y(_1406_));
 sg13g2_a21oi_1 _4759_ (.A1(_1079_),
    .A2(_1101_),
    .Y(_1407_),
    .B1(_1098_));
 sg13g2_mux2_1 _4760_ (.A0(_1091_),
    .A1(_1096_),
    .S(_1097_),
    .X(_1408_));
 sg13g2_mux2_1 _4761_ (.A0(_1408_),
    .A1(_1338_),
    .S(net149),
    .X(_1409_));
 sg13g2_a22oi_1 _4762_ (.Y(_1410_),
    .B1(_1409_),
    .B2(_1098_),
    .A2(_1407_),
    .A1(_1406_));
 sg13g2_inv_1 _4763_ (.Y(_1411_),
    .A(_1165_));
 sg13g2_and2_1 _4764_ (.A(_1168_),
    .B(_1178_),
    .X(_1412_));
 sg13g2_or2_1 _4765_ (.X(_1413_),
    .B(_0433_),
    .A(_0435_));
 sg13g2_inv_1 _4766_ (.Y(_1414_),
    .A(_0429_));
 sg13g2_a21oi_1 _4767_ (.A1(_1414_),
    .A2(_0435_),
    .Y(_1415_),
    .B1(_1177_));
 sg13g2_a22oi_1 _4768_ (.Y(_1416_),
    .B1(_1413_),
    .B2(_1415_),
    .A2(_1175_),
    .A1(_1177_));
 sg13g2_mux4_1 _4769_ (.S0(_1166_),
    .A0(_1182_),
    .A1(_1411_),
    .A2(_1412_),
    .A3(_1416_),
    .S1(net147),
    .X(_1417_));
 sg13g2_mux2_1 _4770_ (.A0(_1410_),
    .A1(_1417_),
    .S(_1094_),
    .X(_1418_));
 sg13g2_buf_2 _4771_ (.A(\g.g_y[5].g_x[3].t.r_v ),
    .X(_1419_));
 sg13g2_buf_2 _4772_ (.A(\g.g_y[5].g_x[3].t.out_sc ),
    .X(_1420_));
 sg13g2_buf_8 _4773_ (.A(\g.g_y[5].g_x[3].t.r_d ),
    .X(_1421_));
 sg13g2_mux2_1 _4774_ (.A0(\g.g_y[5].g_x[3].t.r_gnl ),
    .A1(_1420_),
    .S(_1421_),
    .X(_1422_));
 sg13g2_buf_2 _4775_ (.A(\g.g_y[5].g_x[3].t.r_ghl ),
    .X(_1423_));
 sg13g2_nand2b_1 _4776_ (.Y(_1424_),
    .B(_1419_),
    .A_N(_1423_));
 sg13g2_o21ai_1 _4777_ (.B1(_1424_),
    .Y(_1425_),
    .A1(_1419_),
    .A2(_1422_));
 sg13g2_or2_1 _4778_ (.X(_1426_),
    .B(_0762_),
    .A(_0758_));
 sg13g2_o21ai_1 _4779_ (.B1(_1426_),
    .Y(_1427_),
    .A1(_0763_),
    .A2(_0761_));
 sg13g2_buf_1 _4780_ (.A(\g.g_y[4].g_x[3].t.r_v ),
    .X(_1428_));
 sg13g2_mux2_1 _4781_ (.A0(_1425_),
    .A1(_1427_),
    .S(_1428_),
    .X(_1429_));
 sg13g2_inv_1 _4782_ (.Y(_1430_),
    .A(_1357_));
 sg13g2_or2_1 _4783_ (.X(_1431_),
    .B(_1358_),
    .A(_1430_));
 sg13g2_buf_2 _4784_ (.A(\g.g_y[4].g_x[3].t.r_h ),
    .X(_1432_));
 sg13g2_inv_1 _4785_ (.Y(_1433_),
    .A(_1432_));
 sg13g2_buf_2 _4786_ (.A(\g.g_y[4].g_x[3].t.r_d ),
    .X(_1434_));
 sg13g2_nor2_1 _4787_ (.A(_1084_),
    .B(_1357_),
    .Y(_1435_));
 sg13g2_nor3_1 _4788_ (.A(_1433_),
    .B(_1434_),
    .C(_1435_),
    .Y(_1436_));
 sg13g2_buf_8 _4789_ (.A(\g.g_y[4].g_x[4].t.r_h ),
    .X(_1437_));
 sg13g2_nor2b_1 _4790_ (.A(_1169_),
    .B_N(_1437_),
    .Y(_1438_));
 sg13g2_nor3_1 _4791_ (.A(_1432_),
    .B(_1434_),
    .C(_1438_),
    .Y(_1439_));
 sg13g2_mux2_1 _4792_ (.A0(_1170_),
    .A1(\g.g_y[4].g_x[4].t.r_gnl ),
    .S(_1171_),
    .X(_1440_));
 sg13g2_buf_1 _4793_ (.A(_1440_),
    .X(_1441_));
 sg13g2_inv_2 _4794_ (.Y(_1442_),
    .A(_1437_));
 sg13g2_nand2b_1 _4795_ (.Y(_1443_),
    .B(_1442_),
    .A_N(_1441_));
 sg13g2_a22oi_1 _4796_ (.Y(_1444_),
    .B1(_1439_),
    .B2(_1443_),
    .A2(_1436_),
    .A1(_1431_));
 sg13g2_buf_1 _4797_ (.A(\g.g_y[4].g_x[3].t.out_sc ),
    .X(_1445_));
 sg13g2_nand2b_1 _4798_ (.Y(_1446_),
    .B(_1434_),
    .A_N(_1445_));
 sg13g2_o21ai_1 _4799_ (.B1(_1446_),
    .Y(_1447_),
    .A1(_1429_),
    .A2(_1444_));
 sg13g2_buf_1 _4800_ (.A(_1434_),
    .X(_1448_));
 sg13g2_mux2_1 _4801_ (.A0(_1084_),
    .A1(_1358_),
    .S(_1357_),
    .X(_1449_));
 sg13g2_mux2_1 _4802_ (.A0(_1169_),
    .A1(_1441_),
    .S(_1442_),
    .X(_1450_));
 sg13g2_mux2_1 _4803_ (.A0(_1449_),
    .A1(_1450_),
    .S(_1432_),
    .X(_1451_));
 sg13g2_nand2_1 _4804_ (.Y(_1452_),
    .A(net106),
    .B(_1425_));
 sg13g2_o21ai_1 _4805_ (.B1(_1452_),
    .Y(_1453_),
    .A1(net106),
    .A2(_1451_));
 sg13g2_mux2_1 _4806_ (.A0(_1447_),
    .A1(_1453_),
    .S(_1428_),
    .X(_1454_));
 sg13g2_nand2_1 _4807_ (.Y(_1455_),
    .A(_0766_),
    .B(_0774_));
 sg13g2_a21oi_1 _4808_ (.A1(net159),
    .A2(_1069_),
    .Y(_1456_),
    .B1(_0756_));
 sg13g2_nor2_1 _4809_ (.A(_0757_),
    .B(_0768_),
    .Y(_1457_));
 sg13g2_nand2b_1 _4810_ (.Y(_1458_),
    .B(_1062_),
    .A_N(_0755_));
 sg13g2_a22oi_1 _4811_ (.Y(_1459_),
    .B1(_1457_),
    .B2(_1458_),
    .A2(_1456_),
    .A1(_1455_));
 sg13g2_mux2_1 _4812_ (.A0(_1454_),
    .A1(_1459_),
    .S(_0763_),
    .X(_1460_));
 sg13g2_mux2_1 _4813_ (.A0(_1418_),
    .A1(_1460_),
    .S(_0760_),
    .X(_1461_));
 sg13g2_o21ai_1 _4814_ (.B1(net150),
    .Y(_1462_),
    .A1(_0758_),
    .A2(net38));
 sg13g2_a21oi_1 _4815_ (.A1(net39),
    .A2(_1461_),
    .Y(_0135_),
    .B1(_1462_));
 sg13g2_or2_1 _4816_ (.X(_1463_),
    .B(_1417_),
    .A(_1094_));
 sg13g2_nand2b_1 _4817_ (.Y(_1464_),
    .B(_1094_),
    .A_N(_1410_));
 sg13g2_and2_1 _4818_ (.A(_0762_),
    .B(_1459_),
    .X(_1465_));
 sg13g2_a221oi_1 _4819_ (.B2(_1464_),
    .C1(_1465_),
    .B1(_1463_),
    .A1(_0763_),
    .Y(_1466_),
    .A2(_1454_));
 sg13g2_o21ai_1 _4820_ (.B1(net150),
    .Y(_1467_),
    .A1(\g.g_y[3].g_x[3].t.r_gnl ),
    .A2(net38));
 sg13g2_a21oi_1 _4821_ (.A1(net39),
    .A2(_1466_),
    .Y(_0136_),
    .B1(_1467_));
 sg13g2_nand2_1 _4822_ (.Y(_1468_),
    .A(_0759_),
    .B(net31));
 sg13g2_o21ai_1 _4823_ (.B1(_1094_),
    .Y(_1469_),
    .A1(net52),
    .A2(net108));
 sg13g2_a21oi_1 _4824_ (.A1(_1468_),
    .A2(_1469_),
    .Y(_0137_),
    .B1(net82));
 sg13g2_mux2_1 _4825_ (.A0(_1460_),
    .A1(_1418_),
    .S(_0760_),
    .X(_1470_));
 sg13g2_buf_1 _4826_ (.A(_2719_),
    .X(_1471_));
 sg13g2_a22oi_1 _4827_ (.Y(_1472_),
    .B1(net62),
    .B2(\g.g_y[3].g_x[2].t.out_sc ),
    .A2(net51),
    .A1(_0759_));
 sg13g2_o21ai_1 _4828_ (.B1(_1472_),
    .Y(_0138_),
    .A1(net64),
    .A2(_1470_));
 sg13g2_nand2_1 _4829_ (.Y(_1473_),
    .A(_0759_),
    .B(net30));
 sg13g2_o21ai_1 _4830_ (.B1(_0762_),
    .Y(_1474_),
    .A1(net52),
    .A2(net83));
 sg13g2_a21oi_1 _4831_ (.A1(_1473_),
    .A2(_1474_),
    .Y(_0139_),
    .B1(net82));
 sg13g2_nor2_1 _4832_ (.A(_1182_),
    .B(net28),
    .Y(_1475_));
 sg13g2_a21oi_1 _4833_ (.A1(net147),
    .A2(net22),
    .Y(_1476_),
    .B1(_1475_));
 sg13g2_nor2_1 _4834_ (.A(net87),
    .B(_1476_),
    .Y(_0140_));
 sg13g2_mux2_1 _4835_ (.A0(_1167_),
    .A1(_1182_),
    .S(net66),
    .X(_1477_));
 sg13g2_nor2_1 _4836_ (.A(net87),
    .B(_1477_),
    .Y(_0141_));
 sg13g2_buf_1 _4837_ (.A(net126),
    .X(_1478_));
 sg13g2_a221oi_1 _4838_ (.B2(_1187_),
    .C1(_1160_),
    .B1(_1186_),
    .A1(_1166_),
    .Y(_1479_),
    .A2(_1165_));
 sg13g2_a21oi_1 _4839_ (.A1(_1160_),
    .A2(_1416_),
    .Y(_1480_),
    .B1(_1479_));
 sg13g2_nand2b_1 _4840_ (.Y(_1481_),
    .B(net170),
    .A_N(_0759_));
 sg13g2_o21ai_1 _4841_ (.B1(_1481_),
    .Y(_1482_),
    .A1(net148),
    .A2(_1480_));
 sg13g2_nand2_1 _4842_ (.Y(_1483_),
    .A(net109),
    .B(_1482_));
 sg13g2_o21ai_1 _4843_ (.B1(_1483_),
    .Y(_1484_),
    .A1(_1181_),
    .A2(net121));
 sg13g2_nor2_1 _4844_ (.A(net81),
    .B(_1484_),
    .Y(_0142_));
 sg13g2_inv_1 _4845_ (.Y(_1485_),
    .A(_1177_));
 sg13g2_mux2_1 _4846_ (.A0(_1485_),
    .A1(_1182_),
    .S(net40),
    .X(_1486_));
 sg13g2_nor2_1 _4847_ (.A(net81),
    .B(_1486_),
    .Y(_0143_));
 sg13g2_mux2_1 _4848_ (.A0(_0852_),
    .A1(_0853_),
    .S(net29),
    .X(_1487_));
 sg13g2_and2_1 _4849_ (.A(net107),
    .B(_1487_),
    .X(_0144_));
 sg13g2_buf_8 _4850_ (.A(\g.g_y[4].g_x[5].t.r_d ),
    .X(_1488_));
 sg13g2_inv_1 _4851_ (.Y(_1489_),
    .A(_1488_));
 sg13g2_buf_1 _4852_ (.A(\g.g_y[4].g_x[6].t.r_h ),
    .X(_1490_));
 sg13g2_mux2_1 _4853_ (.A0(_1253_),
    .A1(\g.g_y[4].g_x[6].t.r_gnl ),
    .S(_1254_),
    .X(_1491_));
 sg13g2_buf_1 _4854_ (.A(_1491_),
    .X(_1492_));
 sg13g2_nand2b_1 _4855_ (.Y(_1493_),
    .B(net141),
    .A_N(_1256_));
 sg13g2_o21ai_1 _4856_ (.B1(_1493_),
    .Y(_1494_),
    .A1(net141),
    .A2(_1492_));
 sg13g2_or2_1 _4857_ (.X(_1495_),
    .B(_1437_),
    .A(_1169_));
 sg13g2_o21ai_1 _4858_ (.B1(_1495_),
    .Y(_1496_),
    .A1(_1442_),
    .A2(_1441_));
 sg13g2_buf_2 _4859_ (.A(\g.g_y[5].g_x[5].t.r_v ),
    .X(_1497_));
 sg13g2_buf_2 _4860_ (.A(\g.g_y[5].g_x[5].t.out_sc ),
    .X(_1498_));
 sg13g2_buf_8 _4861_ (.A(\g.g_y[5].g_x[5].t.r_d ),
    .X(_1499_));
 sg13g2_mux2_1 _4862_ (.A0(\g.g_y[5].g_x[5].t.r_gnl ),
    .A1(_1498_),
    .S(_1499_),
    .X(_1500_));
 sg13g2_buf_1 _4863_ (.A(\g.g_y[5].g_x[5].t.r_ghl ),
    .X(_1501_));
 sg13g2_nand2b_1 _4864_ (.Y(_1502_),
    .B(_1497_),
    .A_N(_1501_));
 sg13g2_o21ai_1 _4865_ (.B1(_1502_),
    .Y(_1503_),
    .A1(_1497_),
    .A2(_1500_));
 sg13g2_buf_8 _4866_ (.A(_1503_),
    .X(_1504_));
 sg13g2_nor2_1 _4867_ (.A(_1504_),
    .B(_1496_),
    .Y(_1505_));
 sg13g2_nor2_1 _4868_ (.A(_1504_),
    .B(_1494_),
    .Y(_1506_));
 sg13g2_buf_8 _4869_ (.A(\g.g_y[4].g_x[5].t.r_h ),
    .X(_1507_));
 sg13g2_inv_2 _4870_ (.Y(_1508_),
    .A(_1507_));
 sg13g2_buf_2 _4871_ (.A(\g.g_y[4].g_x[5].t.r_v ),
    .X(_1509_));
 sg13g2_inv_2 _4872_ (.Y(_1510_),
    .A(_1509_));
 sg13g2_mux4_1 _4873_ (.S0(_1508_),
    .A0(_1494_),
    .A1(_1496_),
    .A2(_1505_),
    .A3(_1506_),
    .S1(_1510_),
    .X(_1511_));
 sg13g2_nand2_1 _4874_ (.Y(_1512_),
    .A(_1489_),
    .B(_1511_));
 sg13g2_buf_2 _4875_ (.A(\g.g_y[4].g_x[5].t.out_sc ),
    .X(_1513_));
 sg13g2_nor2_1 _4876_ (.A(_1510_),
    .B(_1504_),
    .Y(_1514_));
 sg13g2_a21oi_1 _4877_ (.A1(_1510_),
    .A2(_1513_),
    .Y(_1515_),
    .B1(_1514_));
 sg13g2_a21oi_1 _4878_ (.A1(_1488_),
    .A2(_1515_),
    .Y(_1516_),
    .B1(_0863_));
 sg13g2_nand2_1 _4879_ (.Y(_1517_),
    .A(_0842_),
    .B(_0860_));
 sg13g2_o21ai_1 _4880_ (.B1(_1517_),
    .Y(_1518_),
    .A1(_0842_),
    .A2(_0850_));
 sg13g2_nand2_1 _4881_ (.Y(_1519_),
    .A(_1137_),
    .B(_1139_));
 sg13g2_mux4_1 _4882_ (.S0(_1143_),
    .A0(_1138_),
    .A1(_1518_),
    .A2(net155),
    .A3(_1519_),
    .S1(_0845_),
    .X(_1520_));
 sg13g2_a22oi_1 _4883_ (.Y(_1521_),
    .B1(_1520_),
    .B2(_0863_),
    .A2(_1516_),
    .A1(_1512_));
 sg13g2_nand3_1 _4884_ (.B(net181),
    .C(_0743_),
    .A(_0853_),
    .Y(_1522_));
 sg13g2_nor2_1 _4885_ (.A(_1521_),
    .B(_1522_),
    .Y(_1523_));
 sg13g2_nand3_1 _4886_ (.B(_1168_),
    .C(_1178_),
    .A(net147),
    .Y(_1524_));
 sg13g2_o21ai_1 _4887_ (.B1(_1166_),
    .Y(_1525_),
    .A1(net147),
    .A2(_1181_));
 sg13g2_inv_1 _4888_ (.Y(_1526_),
    .A(_1525_));
 sg13g2_nor2_1 _4889_ (.A(_1180_),
    .B(_1161_),
    .Y(_1527_));
 sg13g2_a21oi_1 _4890_ (.A1(_1180_),
    .A2(_1416_),
    .Y(_1528_),
    .B1(_1527_));
 sg13g2_a22oi_1 _4891_ (.Y(_1529_),
    .B1(_1528_),
    .B2(_1167_),
    .A2(_1526_),
    .A1(_1524_));
 sg13g2_nand2_1 _4892_ (.Y(_1530_),
    .A(_1252_),
    .B(_1261_));
 sg13g2_nor2b_1 _4893_ (.A(_1251_),
    .B_N(net146),
    .Y(_1531_));
 sg13g2_and2_1 _4894_ (.A(_1251_),
    .B(net146),
    .X(_1532_));
 sg13g2_nor2b_1 _4895_ (.A(net146),
    .B_N(_1251_),
    .Y(_1533_));
 sg13g2_nor2_1 _4896_ (.A(_1251_),
    .B(net146),
    .Y(_1534_));
 sg13g2_a22oi_1 _4897_ (.Y(_1535_),
    .B1(_1534_),
    .B2(_1263_),
    .A2(_1533_),
    .A1(_1249_));
 sg13g2_inv_1 _4898_ (.Y(_1536_),
    .A(_1535_));
 sg13g2_a221oi_1 _4899_ (.B2(_1269_),
    .C1(_1536_),
    .B1(_1532_),
    .A1(_1530_),
    .Y(_1537_),
    .A2(_1531_));
 sg13g2_mux2_1 _4900_ (.A0(_1529_),
    .A1(_1537_),
    .S(_1163_),
    .X(_1538_));
 sg13g2_or4_1 _4901_ (.A(_0853_),
    .B(_2709_),
    .C(net56),
    .D(_1538_),
    .X(_1539_));
 sg13g2_nand3_1 _4902_ (.B(net160),
    .C(net56),
    .A(_0855_),
    .Y(_1540_));
 sg13g2_nand3b_1 _4903_ (.B(_1539_),
    .C(_1540_),
    .Y(_0145_),
    .A_N(_1523_));
 sg13g2_mux2_1 _4904_ (.A0(_1537_),
    .A1(_1529_),
    .S(_1163_),
    .X(_1541_));
 sg13g2_nor2_1 _4905_ (.A(_0863_),
    .B(_1520_),
    .Y(_1542_));
 sg13g2_mux2_1 _4906_ (.A0(_1494_),
    .A1(_1496_),
    .S(_1507_),
    .X(_1543_));
 sg13g2_or2_1 _4907_ (.X(_1544_),
    .B(_0851_),
    .A(_0855_));
 sg13g2_o21ai_1 _4908_ (.B1(_1544_),
    .Y(_1545_),
    .A1(_0863_),
    .A2(_0854_));
 sg13g2_mux2_1 _4909_ (.A0(_1504_),
    .A1(_1545_),
    .S(_1509_),
    .X(_1546_));
 sg13g2_nor3_1 _4910_ (.A(net142),
    .B(_1543_),
    .C(_1546_),
    .Y(_1547_));
 sg13g2_inv_1 _4911_ (.Y(_1548_),
    .A(_1547_));
 sg13g2_nand2b_1 _4912_ (.Y(_1549_),
    .B(net142),
    .A_N(_1513_));
 sg13g2_and2_1 _4913_ (.A(_1510_),
    .B(_1549_),
    .X(_1550_));
 sg13g2_mux2_1 _4914_ (.A0(_1169_),
    .A1(_1441_),
    .S(_1437_),
    .X(_1551_));
 sg13g2_and2_1 _4915_ (.A(_1507_),
    .B(_1493_),
    .X(_1552_));
 sg13g2_or2_1 _4916_ (.X(_1553_),
    .B(_1492_),
    .A(net141));
 sg13g2_a221oi_1 _4917_ (.B2(_1553_),
    .C1(\g.g_y[4].g_x[5].t.r_d ),
    .B1(_1552_),
    .A1(_1508_),
    .Y(_1554_),
    .A2(_1551_));
 sg13g2_a21oi_1 _4918_ (.A1(net142),
    .A2(_1504_),
    .Y(_1555_),
    .B1(_1554_));
 sg13g2_a221oi_1 _4919_ (.B2(_1509_),
    .C1(_0851_),
    .B1(_1555_),
    .A1(_1548_),
    .Y(_1556_),
    .A2(_1550_));
 sg13g2_nor3_1 _4920_ (.A(_1541_),
    .B(_1542_),
    .C(_1556_),
    .Y(_1557_));
 sg13g2_o21ai_1 _4921_ (.B1(net150),
    .Y(_1558_),
    .A1(\g.g_y[3].g_x[5].t.r_gnl ),
    .A2(net32));
 sg13g2_a21oi_1 _4922_ (.A1(net36),
    .A2(_1557_),
    .Y(_0146_),
    .B1(_1558_));
 sg13g2_nand2_1 _4923_ (.Y(_1559_),
    .A(_0852_),
    .B(net31));
 sg13g2_o21ai_1 _4924_ (.B1(_1163_),
    .Y(_1560_),
    .A1(net52),
    .A2(net108));
 sg13g2_a21oi_1 _4925_ (.A1(_1559_),
    .A2(_1560_),
    .Y(_0147_),
    .B1(net82));
 sg13g2_mux2_1 _4926_ (.A0(_1521_),
    .A1(_1538_),
    .S(_0853_),
    .X(_1561_));
 sg13g2_buf_1 _4927_ (.A(_2721_),
    .X(_1562_));
 sg13g2_a22oi_1 _4928_ (.Y(_1563_),
    .B1(net80),
    .B2(_1181_),
    .A2(net51),
    .A1(_0852_));
 sg13g2_o21ai_1 _4929_ (.B1(_1563_),
    .Y(_0148_),
    .A1(net64),
    .A2(_1561_));
 sg13g2_nand2_1 _4930_ (.Y(_1564_),
    .A(_0852_),
    .B(net30));
 sg13g2_buf_1 _4931_ (.A(net99),
    .X(_1565_));
 sg13g2_o21ai_1 _4932_ (.B1(_0851_),
    .Y(_1566_),
    .A1(net50),
    .A2(net83));
 sg13g2_a21oi_1 _4933_ (.A1(_1564_),
    .A2(_1566_),
    .Y(_0149_),
    .B1(net82));
 sg13g2_nor2_1 _4934_ (.A(_1264_),
    .B(net28),
    .Y(_1567_));
 sg13g2_a21oi_1 _4935_ (.A1(_1246_),
    .A2(net22),
    .Y(_1568_),
    .B1(_1567_));
 sg13g2_nor2_1 _4936_ (.A(net81),
    .B(_1568_),
    .Y(_0150_));
 sg13g2_nand2_1 _4937_ (.Y(_1569_),
    .A(_1263_),
    .B(net31));
 sg13g2_o21ai_1 _4938_ (.B1(_1251_),
    .Y(_1570_),
    .A1(net50),
    .A2(net108));
 sg13g2_a21oi_1 _4939_ (.A1(_1569_),
    .A2(_1570_),
    .Y(_0151_),
    .B1(net82));
 sg13g2_nand2_1 _4940_ (.Y(_1571_),
    .A(net115),
    .B(_0852_));
 sg13g2_mux2_1 _4941_ (.A0(_1269_),
    .A1(_1266_),
    .S(_1246_),
    .X(_1572_));
 sg13g2_nand2_1 _4942_ (.Y(_1573_),
    .A(net124),
    .B(_1572_));
 sg13g2_a21oi_1 _4943_ (.A1(_1571_),
    .A2(_1573_),
    .Y(_1574_),
    .B1(_2893_));
 sg13g2_a21oi_1 _4944_ (.A1(_1263_),
    .A2(net91),
    .Y(_1575_),
    .B1(_1574_));
 sg13g2_nor2_1 _4945_ (.A(net81),
    .B(_1575_),
    .Y(_0152_));
 sg13g2_mux2_1 _4946_ (.A0(_1267_),
    .A1(_1264_),
    .S(net61),
    .X(_1576_));
 sg13g2_nor2_1 _4947_ (.A(net81),
    .B(_1576_),
    .Y(_0153_));
 sg13g2_mux2_1 _4948_ (.A0(_0945_),
    .A1(_0946_),
    .S(net29),
    .X(_1577_));
 sg13g2_and2_1 _4949_ (.A(net107),
    .B(_1577_),
    .X(_0154_));
 sg13g2_a22oi_1 _4950_ (.Y(_1578_),
    .B1(_1534_),
    .B2(_1250_),
    .A2(_1533_),
    .A1(_1263_));
 sg13g2_inv_1 _4951_ (.Y(_1579_),
    .A(_1578_));
 sg13g2_a221oi_1 _4952_ (.B2(_1530_),
    .C1(_1579_),
    .B1(_1532_),
    .A1(_1269_),
    .Y(_1580_),
    .A2(_1531_));
 sg13g2_nand3_1 _4953_ (.B(_0980_),
    .C(_1330_),
    .A(net111),
    .Y(_1581_));
 sg13g2_nor2_1 _4954_ (.A(_0975_),
    .B(_1332_),
    .Y(_1582_));
 sg13g2_o21ai_1 _4955_ (.B1(_0975_),
    .Y(_1583_),
    .A1(net111),
    .A2(_0980_));
 sg13g2_a21oi_1 _4956_ (.A1(net111),
    .A2(_1317_),
    .Y(_1584_),
    .B1(_1583_));
 sg13g2_a21oi_1 _4957_ (.A1(_1581_),
    .A2(_1582_),
    .Y(_1585_),
    .B1(_1584_));
 sg13g2_mux2_1 _4958_ (.A0(_1580_),
    .A1(_1585_),
    .S(_1248_),
    .X(_1586_));
 sg13g2_nand2_1 _4959_ (.Y(_1587_),
    .A(net153),
    .B(_0934_));
 sg13g2_o21ai_1 _4960_ (.B1(_1587_),
    .Y(_1588_),
    .A1(net153),
    .A2(_1235_));
 sg13g2_nand3_1 _4961_ (.B(_0937_),
    .C(_1232_),
    .A(net153),
    .Y(_1589_));
 sg13g2_a21oi_1 _4962_ (.A1(net156),
    .A2(_0848_),
    .Y(_1590_),
    .B1(_0928_));
 sg13g2_a21oi_1 _4963_ (.A1(_0933_),
    .A2(_1590_),
    .Y(_1591_),
    .B1(_0939_));
 sg13g2_nand2_1 _4964_ (.Y(_1592_),
    .A(_0933_),
    .B(_0927_));
 sg13g2_nand3_1 _4965_ (.B(_0930_),
    .C(_1232_),
    .A(net153),
    .Y(_1593_));
 sg13g2_and3_1 _4966_ (.X(_1594_),
    .A(_0924_),
    .B(_1592_),
    .C(_1593_));
 sg13g2_a221oi_1 _4967_ (.B2(_1591_),
    .C1(_1594_),
    .B1(_1589_),
    .A1(net154),
    .Y(_1595_),
    .A2(_1588_));
 sg13g2_buf_1 _4968_ (.A(\g.g_y[4].g_x[7].t.r_d ),
    .X(_1596_));
 sg13g2_nor2b_1 _4969_ (.A(net141),
    .B_N(_1256_),
    .Y(_1597_));
 sg13g2_a21oi_1 _4970_ (.A1(net141),
    .A2(_1492_),
    .Y(_1598_),
    .B1(_1597_));
 sg13g2_nand2b_1 _4971_ (.Y(_1599_),
    .B(net144),
    .A_N(_0989_));
 sg13g2_o21ai_1 _4972_ (.B1(_1599_),
    .Y(_1600_),
    .A1(net144),
    .A2(_1362_));
 sg13g2_buf_2 _4973_ (.A(\g.g_y[4].g_x[7].t.r_h ),
    .X(_1601_));
 sg13g2_mux2_1 _4974_ (.A0(_1598_),
    .A1(_1600_),
    .S(_1601_),
    .X(_1602_));
 sg13g2_nand2b_1 _4975_ (.Y(_1603_),
    .B(_1602_),
    .A_N(net140));
 sg13g2_buf_2 _4976_ (.A(\g.g_y[5].g_x[7].t.r_v ),
    .X(_1604_));
 sg13g2_buf_2 _4977_ (.A(\g.g_y[5].g_x[7].t.out_sc ),
    .X(_1605_));
 sg13g2_buf_8 _4978_ (.A(\g.g_y[5].g_x[7].t.r_d ),
    .X(_1606_));
 sg13g2_mux2_1 _4979_ (.A0(\g.g_y[5].g_x[7].t.r_gnl ),
    .A1(_1605_),
    .S(_1606_),
    .X(_1607_));
 sg13g2_buf_1 _4980_ (.A(\g.g_y[5].g_x[7].t.r_ghl ),
    .X(_1608_));
 sg13g2_nand2b_1 _4981_ (.Y(_1609_),
    .B(_1604_),
    .A_N(_1608_));
 sg13g2_o21ai_1 _4982_ (.B1(_1609_),
    .Y(_1610_),
    .A1(_1604_),
    .A2(_1607_));
 sg13g2_buf_1 _4983_ (.A(\g.g_y[4].g_x[7].t.r_v ),
    .X(_1611_));
 sg13g2_inv_1 _4984_ (.Y(_1612_),
    .A(_1611_));
 sg13g2_a21oi_1 _4985_ (.A1(net140),
    .A2(_1610_),
    .Y(_1613_),
    .B1(_1612_));
 sg13g2_buf_1 _4986_ (.A(\g.g_y[4].g_x[7].t.out_sc ),
    .X(_1614_));
 sg13g2_inv_1 _4987_ (.Y(_1615_),
    .A(_1614_));
 sg13g2_a21o_1 _4988_ (.A2(_1492_),
    .A1(net141),
    .B1(_1597_),
    .X(_1616_));
 sg13g2_mux2_1 _4989_ (.A0(_1362_),
    .A1(_0989_),
    .S(net144),
    .X(_1617_));
 sg13g2_inv_1 _4990_ (.Y(_1618_),
    .A(_1601_));
 sg13g2_mux2_1 _4991_ (.A0(_1616_),
    .A1(_1617_),
    .S(_1618_),
    .X(_1619_));
 sg13g2_nor2_1 _4992_ (.A(\g.g_y[4].g_x[7].t.r_d ),
    .B(_1610_),
    .Y(_1620_));
 sg13g2_a221oi_1 _4993_ (.B2(_1620_),
    .C1(_1611_),
    .B1(_1619_),
    .A1(_1596_),
    .Y(_1621_),
    .A2(_1615_));
 sg13g2_a21oi_1 _4994_ (.A1(_1603_),
    .A2(_1613_),
    .Y(_1622_),
    .B1(_1621_));
 sg13g2_mux2_1 _4995_ (.A0(_1595_),
    .A1(_1622_),
    .S(_0944_),
    .X(_1623_));
 sg13g2_mux2_1 _4996_ (.A0(_1586_),
    .A1(_1623_),
    .S(_0946_),
    .X(_1624_));
 sg13g2_o21ai_1 _4997_ (.B1(net150),
    .Y(_1625_),
    .A1(_0948_),
    .A2(net57));
 sg13g2_a21oi_1 _4998_ (.A1(net39),
    .A2(_1624_),
    .Y(_0155_),
    .B1(_1625_));
 sg13g2_mux2_1 _4999_ (.A0(_1622_),
    .A1(_1595_),
    .S(_0944_),
    .X(_1626_));
 sg13g2_mux2_1 _5000_ (.A0(_1585_),
    .A1(_1580_),
    .S(_1248_),
    .X(_1627_));
 sg13g2_nor3_1 _5001_ (.A(_0704_),
    .B(_1626_),
    .C(_1627_),
    .Y(_1628_));
 sg13g2_o21ai_1 _5002_ (.B1(net177),
    .Y(_1629_),
    .A1(\g.g_y[3].g_x[7].t.r_gnl ),
    .A2(net38));
 sg13g2_nor2_1 _5003_ (.A(_1628_),
    .B(_1629_),
    .Y(_0156_));
 sg13g2_nand2_1 _5004_ (.Y(_1630_),
    .A(_0945_),
    .B(net31));
 sg13g2_o21ai_1 _5005_ (.B1(_1248_),
    .Y(_1631_),
    .A1(net50),
    .A2(net108));
 sg13g2_a21oi_1 _5006_ (.A1(_1630_),
    .A2(_1631_),
    .Y(_0157_),
    .B1(net82));
 sg13g2_buf_1 _5007_ (.A(_2715_),
    .X(_1632_));
 sg13g2_mux2_1 _5008_ (.A0(_1623_),
    .A1(_1586_),
    .S(_0946_),
    .X(_1633_));
 sg13g2_a22oi_1 _5009_ (.Y(_1634_),
    .B1(net80),
    .B2(_1263_),
    .A2(net51),
    .A1(_0945_));
 sg13g2_o21ai_1 _5010_ (.B1(_1634_),
    .Y(_0158_),
    .A1(net49),
    .A2(_1633_));
 sg13g2_nand2_1 _5011_ (.Y(_1635_),
    .A(_0945_),
    .B(net30));
 sg13g2_o21ai_1 _5012_ (.B1(_0944_),
    .Y(_1636_),
    .A1(net50),
    .A2(net83));
 sg13g2_a21oi_1 _5013_ (.A1(_1635_),
    .A2(_1636_),
    .Y(_0159_),
    .B1(net82));
 sg13g2_mux2_1 _5014_ (.A0(_0985_),
    .A1(_0986_),
    .S(net29),
    .X(_1637_));
 sg13g2_and2_1 _5015_ (.A(_1301_),
    .B(_1637_),
    .X(_0160_));
 sg13g2_inv_1 _5016_ (.Y(_1638_),
    .A(_0986_));
 sg13g2_mux2_1 _5017_ (.A0(_0997_),
    .A1(_1329_),
    .S(net111),
    .X(_1639_));
 sg13g2_or3_1 _5018_ (.A(net111),
    .B(_0982_),
    .C(_1316_),
    .X(_1640_));
 sg13g2_and2_1 _5019_ (.A(_0974_),
    .B(_0994_),
    .X(_1641_));
 sg13g2_a22oi_1 _5020_ (.Y(_1642_),
    .B1(_1640_),
    .B2(_1641_),
    .A2(_1639_),
    .A1(_1000_));
 sg13g2_buf_1 _5021_ (.A(\g.g_y[5].g_x[0].t.r_d ),
    .X(_1643_));
 sg13g2_mux2_1 _5022_ (.A0(_1347_),
    .A1(\g.g_y[5].g_x[1].t.r_gnl ),
    .S(_1348_),
    .X(_1644_));
 sg13g2_buf_2 _5023_ (.A(\g.g_y[5].g_x[1].t.r_h ),
    .X(_1645_));
 sg13g2_mux2_1 _5024_ (.A0(_1644_),
    .A1(_1350_),
    .S(_1645_),
    .X(_1646_));
 sg13g2_buf_1 _5025_ (.A(_1646_),
    .X(_1647_));
 sg13g2_buf_2 _5026_ (.A(\g.g_y[5].g_x[0].t.r_h ),
    .X(_1648_));
 sg13g2_mux2_1 _5027_ (.A0(net6),
    .A1(_1647_),
    .S(_1648_),
    .X(_1649_));
 sg13g2_or2_1 _5028_ (.X(_1650_),
    .B(_1649_),
    .A(_1643_));
 sg13g2_buf_1 _5029_ (.A(_1650_),
    .X(_1651_));
 sg13g2_buf_1 _5030_ (.A(_1643_),
    .X(_1652_));
 sg13g2_nand2b_1 _5031_ (.Y(_1653_),
    .B(net178),
    .A_N(_2652_));
 sg13g2_o21ai_1 _5032_ (.B1(_1653_),
    .Y(_1654_),
    .A1(net178),
    .A2(_2651_));
 sg13g2_buf_1 _5033_ (.A(\g.g_y[5].g_x[0].t.r_v ),
    .X(_1655_));
 sg13g2_inv_1 _5034_ (.Y(_1656_),
    .A(_1655_));
 sg13g2_a21oi_1 _5035_ (.A1(net105),
    .A2(_1654_),
    .Y(_1657_),
    .B1(_1656_));
 sg13g2_buf_1 _5036_ (.A(\g.g_y[5].g_x[0].t.out_sc ),
    .X(_1658_));
 sg13g2_inv_1 _5037_ (.Y(_1659_),
    .A(_1658_));
 sg13g2_mux2_1 _5038_ (.A0(_1647_),
    .A1(net6),
    .S(_1648_),
    .X(_1660_));
 sg13g2_nor2_1 _5039_ (.A(net105),
    .B(_1654_),
    .Y(_1661_));
 sg13g2_a22oi_1 _5040_ (.Y(_1662_),
    .B1(_1660_),
    .B2(_1661_),
    .A2(_1659_),
    .A1(net105));
 sg13g2_a22oi_1 _5041_ (.Y(_1663_),
    .B1(_1662_),
    .B2(_1656_),
    .A2(_1657_),
    .A1(_1651_));
 sg13g2_mux2_1 _5042_ (.A0(_1642_),
    .A1(_1663_),
    .S(net151),
    .X(_1664_));
 sg13g2_or2_1 _5043_ (.X(_1665_),
    .B(_1664_),
    .A(_1638_));
 sg13g2_mux2_1 _5044_ (.A0(_1354_),
    .A1(_1352_),
    .S(_1355_),
    .X(_1666_));
 sg13g2_mux4_1 _5045_ (.S0(net143),
    .A0(_1374_),
    .A1(_1367_),
    .A2(_1372_),
    .A3(_1666_),
    .S1(_1365_),
    .X(_1667_));
 sg13g2_nand2_1 _5046_ (.Y(_1668_),
    .A(net144),
    .B(_1667_));
 sg13g2_nor2_1 _5047_ (.A(net144),
    .B(net5),
    .Y(_1669_));
 sg13g2_nor2_1 _5048_ (.A(_0986_),
    .B(_1669_),
    .Y(_1670_));
 sg13g2_a21oi_1 _5049_ (.A1(_1668_),
    .A2(_1670_),
    .Y(_1671_),
    .B1(_0457_));
 sg13g2_o21ai_1 _5050_ (.B1(net150),
    .Y(_1672_),
    .A1(_0989_),
    .A2(net45));
 sg13g2_a21oi_1 _5051_ (.A1(_1665_),
    .A2(_1671_),
    .Y(_0161_),
    .B1(_1672_));
 sg13g2_nand2_1 _5052_ (.Y(_1673_),
    .A(_1361_),
    .B(net5));
 sg13g2_or2_1 _5053_ (.X(_1674_),
    .B(_1667_),
    .A(net144));
 sg13g2_mux2_1 _5054_ (.A0(_1663_),
    .A1(_1642_),
    .S(net151),
    .X(_1675_));
 sg13g2_a21oi_1 _5055_ (.A1(_1673_),
    .A2(_1674_),
    .Y(_1676_),
    .B1(_1675_));
 sg13g2_o21ai_1 _5056_ (.B1(net150),
    .Y(_1677_),
    .A1(\g.g_y[4].g_x[0].t.r_gnl ),
    .A2(net45));
 sg13g2_a21oi_1 _5057_ (.A1(net46),
    .A2(_1676_),
    .Y(_0162_),
    .B1(_1677_));
 sg13g2_nand2_1 _5058_ (.Y(_1678_),
    .A(_0985_),
    .B(net31));
 sg13g2_o21ai_1 _5059_ (.B1(_1361_),
    .Y(_1679_),
    .A1(net50),
    .A2(net108));
 sg13g2_a21oi_1 _5060_ (.A1(_1678_),
    .A2(_1679_),
    .Y(_0163_),
    .B1(_1393_));
 sg13g2_nor2_1 _5061_ (.A(_1638_),
    .B(_1669_),
    .Y(_1680_));
 sg13g2_nand3_1 _5062_ (.B(_1668_),
    .C(_1680_),
    .A(net88),
    .Y(_1681_));
 sg13g2_nand3b_1 _5063_ (.B(_1638_),
    .C(net88),
    .Y(_1682_),
    .A_N(_1664_));
 sg13g2_a22oi_1 _5064_ (.Y(_1683_),
    .B1(net96),
    .B2(_0945_),
    .A2(net55),
    .A1(_0985_));
 sg13g2_nand3_1 _5065_ (.B(_1682_),
    .C(_1683_),
    .A(_1681_),
    .Y(_0164_));
 sg13g2_nand2_1 _5066_ (.Y(_1684_),
    .A(_0985_),
    .B(_1308_));
 sg13g2_o21ai_1 _5067_ (.B1(net151),
    .Y(_1685_),
    .A1(_1565_),
    .A2(_1310_));
 sg13g2_a21oi_1 _5068_ (.A1(_1684_),
    .A2(_1685_),
    .Y(_0165_),
    .B1(net82));
 sg13g2_nor2_1 _5069_ (.A(_1374_),
    .B(net28),
    .Y(_1686_));
 sg13g2_a21oi_1 _5070_ (.A1(net143),
    .A2(net22),
    .Y(_1687_),
    .B1(_1686_));
 sg13g2_nor2_1 _5071_ (.A(_1478_),
    .B(_1687_),
    .Y(_0166_));
 sg13g2_nand2_1 _5072_ (.Y(_1688_),
    .A(_1373_),
    .B(net31));
 sg13g2_o21ai_1 _5073_ (.B1(_1365_),
    .Y(_1689_),
    .A1(_1565_),
    .A2(net108));
 sg13g2_buf_1 _5074_ (.A(net128),
    .X(_1690_));
 sg13g2_a21oi_1 _5075_ (.A1(_1688_),
    .A2(_1689_),
    .Y(_0167_),
    .B1(net79));
 sg13g2_nor2_1 _5076_ (.A(_1373_),
    .B(net121),
    .Y(_1691_));
 sg13g2_inv_1 _5077_ (.Y(_1692_),
    .A(net143));
 sg13g2_mux2_1 _5078_ (.A0(_1372_),
    .A1(_1666_),
    .S(_1692_),
    .X(_1693_));
 sg13g2_nand2_1 _5079_ (.Y(_1694_),
    .A(net169),
    .B(_0985_));
 sg13g2_o21ai_1 _5080_ (.B1(_1694_),
    .Y(_1695_),
    .A1(net120),
    .A2(_1693_));
 sg13g2_nor2_1 _5081_ (.A(net91),
    .B(_1695_),
    .Y(_1696_));
 sg13g2_nor3_1 _5082_ (.A(net92),
    .B(_1691_),
    .C(_1696_),
    .Y(_0168_));
 sg13g2_nand2_1 _5083_ (.Y(_1697_),
    .A(_1373_),
    .B(net30));
 sg13g2_o21ai_1 _5084_ (.B1(_1355_),
    .Y(_1698_),
    .A1(net50),
    .A2(net83));
 sg13g2_a21oi_1 _5085_ (.A1(_1697_),
    .A2(_1698_),
    .Y(_0169_),
    .B1(_1690_));
 sg13g2_mux2_1 _5086_ (.A0(_1081_),
    .A1(_1082_),
    .S(net29),
    .X(_1699_));
 sg13g2_and2_1 _5087_ (.A(net107),
    .B(_1699_),
    .X(_0170_));
 sg13g2_nand2_1 _5088_ (.Y(_1700_),
    .A(_1434_),
    .B(_1450_));
 sg13g2_or2_1 _5089_ (.X(_1701_),
    .B(_1445_),
    .A(_1434_));
 sg13g2_o21ai_1 _5090_ (.B1(_1701_),
    .Y(_1702_),
    .A1(_1429_),
    .A2(_1700_));
 sg13g2_inv_1 _5091_ (.Y(_1703_),
    .A(_1428_));
 sg13g2_mux2_1 _5092_ (.A0(_1425_),
    .A1(_1427_),
    .S(_1703_),
    .X(_1704_));
 sg13g2_nor2_1 _5093_ (.A(_1434_),
    .B(_1450_),
    .Y(_1705_));
 sg13g2_a21o_1 _5094_ (.A2(_1704_),
    .A1(net106),
    .B1(_1705_),
    .X(_1706_));
 sg13g2_mux2_1 _5095_ (.A0(_1702_),
    .A1(_1706_),
    .S(_1432_),
    .X(_1707_));
 sg13g2_or3_1 _5096_ (.A(_1692_),
    .B(_1356_),
    .C(_1364_),
    .X(_1708_));
 sg13g2_o21ai_1 _5097_ (.B1(_1365_),
    .Y(_1709_),
    .A1(net143),
    .A2(_1373_));
 sg13g2_inv_1 _5098_ (.Y(_1710_),
    .A(_1709_));
 sg13g2_a21oi_1 _5099_ (.A1(_1692_),
    .A2(_1364_),
    .Y(_1711_),
    .B1(_1365_));
 sg13g2_nand2_1 _5100_ (.Y(_1712_),
    .A(net143),
    .B(_1666_));
 sg13g2_a22oi_1 _5101_ (.Y(_1713_),
    .B1(_1711_),
    .B2(_1712_),
    .A2(_1710_),
    .A1(_1708_));
 sg13g2_mux2_1 _5102_ (.A0(_1707_),
    .A1(_1713_),
    .S(_1430_),
    .X(_1714_));
 sg13g2_a21oi_1 _5103_ (.A1(net149),
    .A2(_1101_),
    .Y(_1715_),
    .B1(_1088_));
 sg13g2_o21ai_1 _5104_ (.B1(_1088_),
    .Y(_1716_),
    .A1(_1079_),
    .A2(_1080_));
 sg13g2_a21oi_1 _5105_ (.A1(_1079_),
    .A2(_1106_),
    .Y(_1717_),
    .B1(_1716_));
 sg13g2_a21oi_1 _5106_ (.A1(_1100_),
    .A2(_1715_),
    .Y(_1718_),
    .B1(_1717_));
 sg13g2_buf_1 _5107_ (.A(\g.g_y[5].g_x[2].t.r_d ),
    .X(_1719_));
 sg13g2_buf_1 _5108_ (.A(_1719_),
    .X(_1720_));
 sg13g2_mux2_1 _5109_ (.A0(_1350_),
    .A1(_1644_),
    .S(_1645_),
    .X(_1721_));
 sg13g2_mux2_1 _5110_ (.A0(_1420_),
    .A1(\g.g_y[5].g_x[3].t.r_gnl ),
    .S(_1421_),
    .X(_1722_));
 sg13g2_buf_2 _5111_ (.A(\g.g_y[5].g_x[3].t.r_h ),
    .X(_1723_));
 sg13g2_inv_1 _5112_ (.Y(_1724_),
    .A(_1723_));
 sg13g2_mux2_1 _5113_ (.A0(_1423_),
    .A1(_1722_),
    .S(_1724_),
    .X(_1725_));
 sg13g2_buf_1 _5114_ (.A(\g.g_y[5].g_x[2].t.r_h ),
    .X(_1726_));
 sg13g2_inv_1 _5115_ (.Y(_1727_),
    .A(_1726_));
 sg13g2_mux2_1 _5116_ (.A0(_1721_),
    .A1(_1725_),
    .S(_1727_),
    .X(_1728_));
 sg13g2_mux2_1 _5117_ (.A0(_2803_),
    .A1(_2804_),
    .S(_2800_),
    .X(_1729_));
 sg13g2_buf_1 _5118_ (.A(_1729_),
    .X(_1730_));
 sg13g2_nand3b_1 _5119_ (.B(_1728_),
    .C(_1730_),
    .Y(_1731_),
    .A_N(net104));
 sg13g2_buf_2 _5120_ (.A(\g.g_y[5].g_x[2].t.r_v ),
    .X(_1732_));
 sg13g2_buf_2 _5121_ (.A(\g.g_y[5].g_x[2].t.out_sc ),
    .X(_1733_));
 sg13g2_nor2b_1 _5122_ (.A(_1733_),
    .B_N(_1719_),
    .Y(_1734_));
 sg13g2_nor2_1 _5123_ (.A(_1732_),
    .B(_1734_),
    .Y(_1735_));
 sg13g2_mux2_1 _5124_ (.A0(_1721_),
    .A1(_1725_),
    .S(_1726_),
    .X(_1736_));
 sg13g2_buf_1 _5125_ (.A(_1736_),
    .X(_1737_));
 sg13g2_mux2_1 _5126_ (.A0(_1737_),
    .A1(_1730_),
    .S(net104),
    .X(_1738_));
 sg13g2_a22oi_1 _5127_ (.Y(_1739_),
    .B1(_1738_),
    .B2(_1732_),
    .A2(_1735_),
    .A1(_1731_));
 sg13g2_mux2_1 _5128_ (.A0(_1718_),
    .A1(_1739_),
    .S(_1085_),
    .X(_1740_));
 sg13g2_mux2_1 _5129_ (.A0(_1714_),
    .A1(_1740_),
    .S(_1082_),
    .X(_1741_));
 sg13g2_o21ai_1 _5130_ (.B1(net150),
    .Y(_1742_),
    .A1(_1084_),
    .A2(_2753_));
 sg13g2_a21oi_1 _5131_ (.A1(net60),
    .A2(_1741_),
    .Y(_0171_),
    .B1(_1742_));
 sg13g2_mux2_1 _5132_ (.A0(_1739_),
    .A1(_1718_),
    .S(_1085_),
    .X(_1743_));
 sg13g2_mux2_1 _5133_ (.A0(_1707_),
    .A1(_1713_),
    .S(_1357_),
    .X(_1744_));
 sg13g2_nor3_1 _5134_ (.A(_0596_),
    .B(_1743_),
    .C(_1744_),
    .Y(_1745_));
 sg13g2_o21ai_1 _5135_ (.B1(net177),
    .Y(_1746_),
    .A1(\g.g_y[4].g_x[2].t.r_gnl ),
    .A2(net59));
 sg13g2_nor2_1 _5136_ (.A(_1745_),
    .B(_1746_),
    .Y(_0172_));
 sg13g2_buf_1 _5137_ (.A(net66),
    .X(_1747_));
 sg13g2_nand2_1 _5138_ (.Y(_1748_),
    .A(_1081_),
    .B(net27));
 sg13g2_buf_1 _5139_ (.A(_2699_),
    .X(_1749_));
 sg13g2_o21ai_1 _5140_ (.B1(_1357_),
    .Y(_1750_),
    .A1(net50),
    .A2(net103));
 sg13g2_a21oi_1 _5141_ (.A1(_1748_),
    .A2(_1750_),
    .Y(_0173_),
    .B1(net79));
 sg13g2_mux2_1 _5142_ (.A0(_1740_),
    .A1(_1714_),
    .S(_1082_),
    .X(_1751_));
 sg13g2_a22oi_1 _5143_ (.Y(_1752_),
    .B1(net80),
    .B2(_1373_),
    .A2(net51),
    .A1(_1081_));
 sg13g2_o21ai_1 _5144_ (.B1(_1752_),
    .Y(_0174_),
    .A1(net49),
    .A2(_1751_));
 sg13g2_nand2_1 _5145_ (.Y(_1753_),
    .A(_1081_),
    .B(net30));
 sg13g2_o21ai_1 _5146_ (.B1(_1085_),
    .Y(_1754_),
    .A1(net50),
    .A2(net83));
 sg13g2_a21oi_1 _5147_ (.A1(_1753_),
    .A2(_1754_),
    .Y(_0175_),
    .B1(net79));
 sg13g2_mux2_1 _5148_ (.A0(_1445_),
    .A1(_1448_),
    .S(net29),
    .X(_1755_));
 sg13g2_and2_1 _5149_ (.A(net107),
    .B(_1755_),
    .X(_0176_));
 sg13g2_nand2_1 _5150_ (.Y(_1756_),
    .A(_1445_),
    .B(net27));
 sg13g2_buf_1 _5151_ (.A(net99),
    .X(_1757_));
 sg13g2_o21ai_1 _5152_ (.B1(_1432_),
    .Y(_1758_),
    .A1(net48),
    .A2(net103));
 sg13g2_a21oi_1 _5153_ (.A1(_1756_),
    .A2(_1758_),
    .Y(_0177_),
    .B1(net79));
 sg13g2_nor2_1 _5154_ (.A(_1445_),
    .B(net121),
    .Y(_1759_));
 sg13g2_and2_1 _5155_ (.A(net115),
    .B(_1081_),
    .X(_1760_));
 sg13g2_nor2_1 _5156_ (.A(net106),
    .B(_1704_),
    .Y(_1761_));
 sg13g2_a21oi_1 _5157_ (.A1(net106),
    .A2(_1451_),
    .Y(_1762_),
    .B1(_1761_));
 sg13g2_nor2_1 _5158_ (.A(net120),
    .B(_1762_),
    .Y(_1763_));
 sg13g2_nor3_1 _5159_ (.A(net91),
    .B(_1760_),
    .C(_1763_),
    .Y(_1764_));
 sg13g2_nor3_1 _5160_ (.A(net92),
    .B(_1759_),
    .C(_1764_),
    .Y(_0178_));
 sg13g2_nand2_1 _5161_ (.Y(_1765_),
    .A(_1445_),
    .B(net30));
 sg13g2_o21ai_1 _5162_ (.B1(_1428_),
    .Y(_1766_),
    .A1(net48),
    .A2(net83));
 sg13g2_a21oi_1 _5163_ (.A1(_1765_),
    .A2(_1766_),
    .Y(_0179_),
    .B1(net79));
 sg13g2_buf_1 _5164_ (.A(net181),
    .X(_1767_));
 sg13g2_mux2_1 _5165_ (.A0(_1170_),
    .A1(_1171_),
    .S(net29),
    .X(_1768_));
 sg13g2_and2_1 _5166_ (.A(net102),
    .B(_1768_),
    .X(_0180_));
 sg13g2_or3_1 _5167_ (.A(_1489_),
    .B(_1543_),
    .C(_1546_),
    .X(_1769_));
 sg13g2_nor2_1 _5168_ (.A(net142),
    .B(_1513_),
    .Y(_1770_));
 sg13g2_nor2_1 _5169_ (.A(_1507_),
    .B(_1770_),
    .Y(_1771_));
 sg13g2_mux2_1 _5170_ (.A0(_1504_),
    .A1(_1545_),
    .S(_1510_),
    .X(_1772_));
 sg13g2_a21oi_1 _5171_ (.A1(net142),
    .A2(_1772_),
    .Y(_1773_),
    .B1(_1554_));
 sg13g2_a22oi_1 _5172_ (.Y(_1774_),
    .B1(_1773_),
    .B2(_1507_),
    .A2(_1771_),
    .A1(_1769_));
 sg13g2_nand3b_1 _5173_ (.B(net106),
    .C(_1449_),
    .Y(_1775_),
    .A_N(_1429_));
 sg13g2_nand2_1 _5174_ (.Y(_1776_),
    .A(_1432_),
    .B(_1701_));
 sg13g2_inv_1 _5175_ (.Y(_1777_),
    .A(_1776_));
 sg13g2_nor2_1 _5176_ (.A(_1434_),
    .B(_1449_),
    .Y(_1778_));
 sg13g2_a21oi_1 _5177_ (.A1(net106),
    .A2(_1704_),
    .Y(_1779_),
    .B1(_1778_));
 sg13g2_a22oi_1 _5178_ (.Y(_1780_),
    .B1(_1779_),
    .B2(_1433_),
    .A2(_1777_),
    .A1(_1775_));
 sg13g2_mux2_1 _5179_ (.A0(_1774_),
    .A1(_1780_),
    .S(_1442_),
    .X(_1781_));
 sg13g2_buf_2 _5180_ (.A(\g.g_y[5].g_x[4].t.out_sc ),
    .X(_1782_));
 sg13g2_buf_1 _5181_ (.A(\g.g_y[5].g_x[4].t.r_d ),
    .X(_1783_));
 sg13g2_nand2b_1 _5182_ (.Y(_1784_),
    .B(net139),
    .A_N(_1782_));
 sg13g2_buf_2 _5183_ (.A(\g.g_y[5].g_x[4].t.r_v ),
    .X(_1785_));
 sg13g2_inv_2 _5184_ (.Y(_1786_),
    .A(_1785_));
 sg13g2_nand2b_1 _5185_ (.Y(_1787_),
    .B(_1786_),
    .A_N(_1784_));
 sg13g2_or2_1 _5186_ (.X(_1788_),
    .B(_0406_),
    .A(_0403_));
 sg13g2_buf_1 _5187_ (.A(_1788_),
    .X(_1789_));
 sg13g2_nand2b_1 _5188_ (.Y(_1790_),
    .B(_0403_),
    .A_N(_0407_));
 sg13g2_and2_1 _5189_ (.A(_1785_),
    .B(_1790_),
    .X(_1791_));
 sg13g2_mux2_1 _5190_ (.A0(_1169_),
    .A1(_1172_),
    .S(_1173_),
    .X(_1792_));
 sg13g2_buf_1 _5191_ (.A(_1792_),
    .X(_1793_));
 sg13g2_inv_1 _5192_ (.Y(_1794_),
    .A(\g.g_y[5].g_x[4].t.r_d ));
 sg13g2_a221oi_1 _5193_ (.B2(_1786_),
    .C1(_1794_),
    .B1(_1793_),
    .A1(_1789_),
    .Y(_1795_),
    .A2(_1791_));
 sg13g2_buf_1 _5194_ (.A(_1795_),
    .X(_1796_));
 sg13g2_buf_1 _5195_ (.A(\g.g_y[5].g_x[4].t.r_h ),
    .X(_1797_));
 sg13g2_mux2_1 _5196_ (.A0(_1498_),
    .A1(\g.g_y[5].g_x[5].t.r_gnl ),
    .S(_1499_),
    .X(_1798_));
 sg13g2_buf_2 _5197_ (.A(\g.g_y[5].g_x[5].t.r_h ),
    .X(_1799_));
 sg13g2_mux2_1 _5198_ (.A0(_1798_),
    .A1(_1501_),
    .S(_1799_),
    .X(_1800_));
 sg13g2_buf_2 _5199_ (.A(_1800_),
    .X(_1801_));
 sg13g2_or2_1 _5200_ (.X(_1802_),
    .B(_1722_),
    .A(_1724_));
 sg13g2_buf_1 _5201_ (.A(_1802_),
    .X(_1803_));
 sg13g2_inv_1 _5202_ (.Y(_1804_),
    .A(_1423_));
 sg13g2_a21oi_1 _5203_ (.A1(_1804_),
    .A2(_1724_),
    .Y(_1805_),
    .B1(net138));
 sg13g2_a221oi_1 _5204_ (.B2(_1805_),
    .C1(net139),
    .B1(_1803_),
    .A1(net138),
    .Y(_1806_),
    .A2(_1801_));
 sg13g2_o21ai_1 _5205_ (.B1(_1785_),
    .Y(_1807_),
    .A1(_1796_),
    .A2(_1806_));
 sg13g2_a21oi_1 _5206_ (.A1(_1787_),
    .A2(_1807_),
    .Y(_1808_),
    .B1(_1174_));
 sg13g2_nand2_1 _5207_ (.Y(_1809_),
    .A(net147),
    .B(_1182_));
 sg13g2_nor3_1 _5208_ (.A(_1173_),
    .B(_1485_),
    .C(_1809_),
    .Y(_1810_));
 sg13g2_inv_1 _5209_ (.Y(_1811_),
    .A(net138));
 sg13g2_o21ai_1 _5210_ (.B1(net138),
    .Y(_1812_),
    .A1(_1423_),
    .A2(_1723_));
 sg13g2_inv_1 _5211_ (.Y(_1813_),
    .A(_1812_));
 sg13g2_a22oi_1 _5212_ (.Y(_1814_),
    .B1(_1803_),
    .B2(_1813_),
    .A2(_1801_),
    .A1(_1811_));
 sg13g2_and2_1 _5213_ (.A(_1786_),
    .B(_1790_),
    .X(_1815_));
 sg13g2_a22oi_1 _5214_ (.Y(_1816_),
    .B1(_1815_),
    .B2(_1789_),
    .A2(_1793_),
    .A1(_1785_));
 sg13g2_nor3_1 _5215_ (.A(net139),
    .B(_1814_),
    .C(_1816_),
    .Y(_1817_));
 sg13g2_and3_1 _5216_ (.X(_1818_),
    .A(_1173_),
    .B(_1786_),
    .C(_1817_));
 sg13g2_o21ai_1 _5217_ (.B1(_1485_),
    .Y(_1819_),
    .A1(_1160_),
    .A2(_1176_));
 sg13g2_o21ai_1 _5218_ (.B1(_1174_),
    .Y(_1820_),
    .A1(_1188_),
    .A2(_1819_));
 sg13g2_a21oi_1 _5219_ (.A1(_1177_),
    .A2(_1179_),
    .Y(_1821_),
    .B1(_1820_));
 sg13g2_or4_1 _5220_ (.A(_1808_),
    .B(_1810_),
    .C(_1818_),
    .D(_1821_),
    .X(_1822_));
 sg13g2_mux2_1 _5221_ (.A0(_1781_),
    .A1(_1822_),
    .S(_1171_),
    .X(_1823_));
 sg13g2_buf_1 _5222_ (.A(net184),
    .X(_1824_));
 sg13g2_o21ai_1 _5223_ (.B1(net137),
    .Y(_1825_),
    .A1(_1169_),
    .A2(_2598_));
 sg13g2_a21oi_1 _5224_ (.A1(net46),
    .A2(_1823_),
    .Y(_0181_),
    .B1(_1825_));
 sg13g2_a21oi_1 _5225_ (.A1(net147),
    .A2(_1182_),
    .Y(_1826_),
    .B1(_1485_));
 sg13g2_nor2_1 _5226_ (.A(_1188_),
    .B(_1819_),
    .Y(_1827_));
 sg13g2_a21oi_1 _5227_ (.A1(_1179_),
    .A2(_1826_),
    .Y(_1828_),
    .B1(_1827_));
 sg13g2_nand2b_1 _5228_ (.Y(_1829_),
    .B(_1437_),
    .A_N(_1780_));
 sg13g2_or2_1 _5229_ (.X(_1830_),
    .B(_1774_),
    .A(_1437_));
 sg13g2_nor3_1 _5230_ (.A(_1786_),
    .B(_1796_),
    .C(_1806_),
    .Y(_1831_));
 sg13g2_nand2_1 _5231_ (.Y(_1832_),
    .A(_1786_),
    .B(_1784_));
 sg13g2_nor2_1 _5232_ (.A(_1817_),
    .B(_1832_),
    .Y(_1833_));
 sg13g2_nor3_1 _5233_ (.A(_1173_),
    .B(_1831_),
    .C(_1833_),
    .Y(_1834_));
 sg13g2_a221oi_1 _5234_ (.B2(_1830_),
    .C1(_1834_),
    .B1(_1829_),
    .A1(_1173_),
    .Y(_1835_),
    .A2(_1828_));
 sg13g2_o21ai_1 _5235_ (.B1(net137),
    .Y(_1836_),
    .A1(\g.g_y[4].g_x[4].t.r_gnl ),
    .A2(_2598_));
 sg13g2_a21oi_1 _5236_ (.A1(net46),
    .A2(_1835_),
    .Y(_0182_),
    .B1(_1836_));
 sg13g2_nand2_1 _5237_ (.Y(_1837_),
    .A(_1170_),
    .B(net27));
 sg13g2_o21ai_1 _5238_ (.B1(_1437_),
    .Y(_1838_),
    .A1(net48),
    .A2(net103));
 sg13g2_a21oi_1 _5239_ (.A1(_1837_),
    .A2(_1838_),
    .Y(_0183_),
    .B1(net79));
 sg13g2_nor2b_1 _5240_ (.A(net115),
    .B_N(_1171_),
    .Y(_1839_));
 sg13g2_nor2_1 _5241_ (.A(net115),
    .B(_1171_),
    .Y(_1840_));
 sg13g2_nand2b_1 _5242_ (.Y(_1841_),
    .B(net148),
    .A_N(_1445_));
 sg13g2_nand2b_1 _5243_ (.Y(_1842_),
    .B(_1841_),
    .A_N(_2713_));
 sg13g2_a221oi_1 _5244_ (.B2(_1822_),
    .C1(_1842_),
    .B1(_1840_),
    .A1(_1781_),
    .Y(_1843_),
    .A2(_1839_));
 sg13g2_a21o_1 _5245_ (.A2(net63),
    .A1(_1170_),
    .B1(_1843_),
    .X(_0184_));
 sg13g2_buf_1 _5246_ (.A(net61),
    .X(_1844_));
 sg13g2_nand2_1 _5247_ (.Y(_1845_),
    .A(_1170_),
    .B(net26));
 sg13g2_buf_1 _5248_ (.A(net127),
    .X(_1846_));
 sg13g2_o21ai_1 _5249_ (.B1(_1173_),
    .Y(_1847_),
    .A1(net48),
    .A2(net78));
 sg13g2_a21oi_1 _5250_ (.A1(_1845_),
    .A2(_1847_),
    .Y(_0185_),
    .B1(_1690_));
 sg13g2_mux2_1 _5251_ (.A0(_1513_),
    .A1(net142),
    .S(net29),
    .X(_1848_));
 sg13g2_and2_1 _5252_ (.A(net102),
    .B(_1848_),
    .X(_0186_));
 sg13g2_nand2_1 _5253_ (.Y(_1849_),
    .A(_1513_),
    .B(net27));
 sg13g2_o21ai_1 _5254_ (.B1(_1507_),
    .Y(_1850_),
    .A1(net48),
    .A2(net103));
 sg13g2_a21oi_1 _5255_ (.A1(_1849_),
    .A2(_1850_),
    .Y(_0187_),
    .B1(net79));
 sg13g2_nand2_1 _5256_ (.Y(_1851_),
    .A(_1513_),
    .B(net91));
 sg13g2_and2_1 _5257_ (.A(net115),
    .B(_1170_),
    .X(_1852_));
 sg13g2_and2_1 _5258_ (.A(_1489_),
    .B(_1772_),
    .X(_1853_));
 sg13g2_a221oi_1 _5259_ (.B2(_1553_),
    .C1(_1489_),
    .B1(_1552_),
    .A1(_1508_),
    .Y(_1854_),
    .A2(_1551_));
 sg13g2_nor3_1 _5260_ (.A(net115),
    .B(_1853_),
    .C(_1854_),
    .Y(_1855_));
 sg13g2_o21ai_1 _5261_ (.B1(net110),
    .Y(_1856_),
    .A1(_1852_),
    .A2(_1855_));
 sg13g2_a21oi_1 _5262_ (.A1(_1851_),
    .A2(_1856_),
    .Y(_0188_),
    .B1(net79));
 sg13g2_nand2_1 _5263_ (.Y(_1857_),
    .A(_1513_),
    .B(net26));
 sg13g2_o21ai_1 _5264_ (.B1(_1509_),
    .Y(_1858_),
    .A1(net48),
    .A2(net78));
 sg13g2_buf_1 _5265_ (.A(net128),
    .X(_1859_));
 sg13g2_a21oi_1 _5266_ (.A1(_1857_),
    .A2(_1858_),
    .Y(_0189_),
    .B1(net77));
 sg13g2_mux2_1 _5267_ (.A0(_1253_),
    .A1(_1254_),
    .S(_1326_),
    .X(_1860_));
 sg13g2_and2_1 _5268_ (.A(net102),
    .B(_1860_),
    .X(_0190_));
 sg13g2_nor2_1 _5269_ (.A(_1508_),
    .B(_1770_),
    .Y(_1861_));
 sg13g2_a22oi_1 _5270_ (.Y(_1862_),
    .B1(_1861_),
    .B2(_1769_),
    .A2(_1773_),
    .A1(_1508_));
 sg13g2_nand2_1 _5271_ (.Y(_1863_),
    .A(_1601_),
    .B(_1616_));
 sg13g2_nand2_1 _5272_ (.Y(_1864_),
    .A(_1618_),
    .B(_1617_));
 sg13g2_nor2b_1 _5273_ (.A(_0944_),
    .B_N(_0948_),
    .Y(_1865_));
 sg13g2_a21oi_2 _5274_ (.B1(_1865_),
    .Y(_1866_),
    .A2(_0947_),
    .A1(_0944_));
 sg13g2_mux2_1 _5275_ (.A0(_1610_),
    .A1(_1866_),
    .S(_1611_),
    .X(_1867_));
 sg13g2_a21oi_1 _5276_ (.A1(_1863_),
    .A2(_1864_),
    .Y(_1868_),
    .B1(_1867_));
 sg13g2_mux2_1 _5277_ (.A0(_1610_),
    .A1(_1866_),
    .S(_1612_),
    .X(_1869_));
 sg13g2_mux4_1 _5278_ (.S0(_1601_),
    .A0(_1615_),
    .A1(_1600_),
    .A2(_1868_),
    .A3(_1869_),
    .S1(net140),
    .X(_1870_));
 sg13g2_mux2_1 _5279_ (.A0(_1862_),
    .A1(_1870_),
    .S(_1490_),
    .X(_1871_));
 sg13g2_a21oi_1 _5280_ (.A1(net146),
    .A2(_1264_),
    .Y(_1872_),
    .B1(_1267_));
 sg13g2_a22oi_1 _5281_ (.Y(_1873_),
    .B1(_1872_),
    .B2(_1262_),
    .A2(_1270_),
    .A1(_1267_));
 sg13g2_buf_1 _5282_ (.A(\g.g_y[5].g_x[6].t.out_sc ),
    .X(_1874_));
 sg13g2_inv_1 _5283_ (.Y(_1875_),
    .A(_1874_));
 sg13g2_nand2b_1 _5284_ (.Y(_1876_),
    .B(_0534_),
    .A_N(_0539_));
 sg13g2_o21ai_1 _5285_ (.B1(_1876_),
    .Y(_1877_),
    .A1(_0534_),
    .A2(_0538_));
 sg13g2_buf_2 _5286_ (.A(\g.g_y[5].g_x[7].t.r_h ),
    .X(_1878_));
 sg13g2_mux2_1 _5287_ (.A0(_1605_),
    .A1(\g.g_y[5].g_x[7].t.r_gnl ),
    .S(_1606_),
    .X(_1879_));
 sg13g2_nand2b_1 _5288_ (.Y(_1880_),
    .B(_1878_),
    .A_N(_1608_));
 sg13g2_o21ai_1 _5289_ (.B1(_1880_),
    .Y(_1881_),
    .A1(_1878_),
    .A2(_1879_));
 sg13g2_nor2b_1 _5290_ (.A(_1799_),
    .B_N(_1501_),
    .Y(_1882_));
 sg13g2_a21oi_1 _5291_ (.A1(_1799_),
    .A2(_1798_),
    .Y(_1883_),
    .B1(_1882_));
 sg13g2_buf_2 _5292_ (.A(\g.g_y[5].g_x[6].t.r_h ),
    .X(_1884_));
 sg13g2_mux2_1 _5293_ (.A0(_1881_),
    .A1(_1883_),
    .S(_1884_),
    .X(_1885_));
 sg13g2_nor2b_1 _5294_ (.A(_1257_),
    .B_N(_1256_),
    .Y(_1886_));
 sg13g2_a21oi_1 _5295_ (.A1(_1257_),
    .A2(_1255_),
    .Y(_1887_),
    .B1(_1886_));
 sg13g2_buf_2 _5296_ (.A(\g.g_y[5].g_x[6].t.r_v ),
    .X(_1888_));
 sg13g2_mux2_1 _5297_ (.A0(_1877_),
    .A1(_1887_),
    .S(_1888_),
    .X(_1889_));
 sg13g2_nor2_2 _5298_ (.A(_1885_),
    .B(_1889_),
    .Y(_1890_));
 sg13g2_mux2_1 _5299_ (.A0(_1883_),
    .A1(_1881_),
    .S(_1884_),
    .X(_1891_));
 sg13g2_buf_2 _5300_ (.A(\g.g_y[5].g_x[6].t.r_d ),
    .X(_1892_));
 sg13g2_inv_1 _5301_ (.Y(_1893_),
    .A(_1892_));
 sg13g2_mux4_1 _5302_ (.S0(_1888_),
    .A0(_1875_),
    .A1(_1877_),
    .A2(_1890_),
    .A3(_1891_),
    .S1(_1893_),
    .X(_1894_));
 sg13g2_mux2_1 _5303_ (.A0(_1873_),
    .A1(_1894_),
    .S(_1257_),
    .X(_1895_));
 sg13g2_mux2_1 _5304_ (.A0(_1871_),
    .A1(_1895_),
    .S(_1254_),
    .X(_1896_));
 sg13g2_o21ai_1 _5305_ (.B1(net137),
    .Y(_1897_),
    .A1(_1256_),
    .A2(_2753_));
 sg13g2_a21oi_1 _5306_ (.A1(net60),
    .A2(_1896_),
    .Y(_0191_),
    .B1(_1897_));
 sg13g2_nand2b_1 _5307_ (.Y(_1898_),
    .B(net141),
    .A_N(_1862_));
 sg13g2_or2_1 _5308_ (.X(_1899_),
    .B(_1870_),
    .A(_1490_));
 sg13g2_nor2b_1 _5309_ (.A(_1257_),
    .B_N(_1894_),
    .Y(_1900_));
 sg13g2_a221oi_1 _5310_ (.B2(_1899_),
    .C1(_1900_),
    .B1(_1898_),
    .A1(_1257_),
    .Y(_1901_),
    .A2(_1873_));
 sg13g2_o21ai_1 _5311_ (.B1(net137),
    .Y(_1902_),
    .A1(\g.g_y[4].g_x[6].t.r_gnl ),
    .A2(_2753_));
 sg13g2_a21oi_1 _5312_ (.A1(net60),
    .A2(_1901_),
    .Y(_0192_),
    .B1(_1902_));
 sg13g2_nand2_1 _5313_ (.Y(_1903_),
    .A(_1253_),
    .B(net27));
 sg13g2_o21ai_1 _5314_ (.B1(net141),
    .Y(_1904_),
    .A1(_1757_),
    .A2(net103));
 sg13g2_a21oi_1 _5315_ (.A1(_1903_),
    .A2(_1904_),
    .Y(_0193_),
    .B1(net77));
 sg13g2_mux2_1 _5316_ (.A0(_1895_),
    .A1(_1871_),
    .S(_1254_),
    .X(_1905_));
 sg13g2_a22oi_1 _5317_ (.Y(_1906_),
    .B1(net80),
    .B2(_1513_),
    .A2(net51),
    .A1(_1253_));
 sg13g2_o21ai_1 _5318_ (.B1(_1906_),
    .Y(_0194_),
    .A1(net49),
    .A2(_1905_));
 sg13g2_nand2_1 _5319_ (.Y(_1907_),
    .A(_1253_),
    .B(net26));
 sg13g2_o21ai_1 _5320_ (.B1(_1257_),
    .Y(_1908_),
    .A1(net48),
    .A2(net78));
 sg13g2_a21oi_1 _5321_ (.A1(_1907_),
    .A2(_1908_),
    .Y(_0195_),
    .B1(net77));
 sg13g2_nor2_1 _5322_ (.A(_1615_),
    .B(net28),
    .Y(_1909_));
 sg13g2_a21oi_1 _5323_ (.A1(net140),
    .A2(net22),
    .Y(_1910_),
    .B1(_1909_));
 sg13g2_nor2_1 _5324_ (.A(net81),
    .B(_1910_),
    .Y(_0196_));
 sg13g2_nand2_1 _5325_ (.Y(_1911_),
    .A(_1614_),
    .B(net27));
 sg13g2_o21ai_1 _5326_ (.B1(_1601_),
    .Y(_1912_),
    .A1(_1757_),
    .A2(net103));
 sg13g2_a21oi_1 _5327_ (.A1(_1911_),
    .A2(_1912_),
    .Y(_0197_),
    .B1(_1859_));
 sg13g2_nor2_1 _5328_ (.A(_1614_),
    .B(net110),
    .Y(_1913_));
 sg13g2_mux2_1 _5329_ (.A0(_1869_),
    .A1(_1602_),
    .S(net140),
    .X(_1914_));
 sg13g2_nand2_1 _5330_ (.Y(_1915_),
    .A(net169),
    .B(_1253_));
 sg13g2_o21ai_1 _5331_ (.B1(_1915_),
    .Y(_1916_),
    .A1(net120),
    .A2(_1914_));
 sg13g2_nor2_1 _5332_ (.A(net91),
    .B(_1916_),
    .Y(_1917_));
 sg13g2_nor3_1 _5333_ (.A(net92),
    .B(_1913_),
    .C(_1917_),
    .Y(_0198_));
 sg13g2_mux2_1 _5334_ (.A0(_1612_),
    .A1(_1615_),
    .S(net61),
    .X(_1918_));
 sg13g2_nor2_1 _5335_ (.A(net81),
    .B(_1918_),
    .Y(_0199_));
 sg13g2_nor2_1 _5336_ (.A(_1659_),
    .B(net28),
    .Y(_1919_));
 sg13g2_a21oi_1 _5337_ (.A1(_1652_),
    .A2(net41),
    .Y(_1920_),
    .B1(_1919_));
 sg13g2_nor2_1 _5338_ (.A(net81),
    .B(_1920_),
    .Y(_0200_));
 sg13g2_nand2_1 _5339_ (.Y(_1921_),
    .A(_1658_),
    .B(net27));
 sg13g2_o21ai_1 _5340_ (.B1(_1648_),
    .Y(_1922_),
    .A1(net48),
    .A2(net103));
 sg13g2_a21oi_1 _5341_ (.A1(_1921_),
    .A2(_1922_),
    .Y(_0201_),
    .B1(net77));
 sg13g2_mux2_1 _5342_ (.A0(_2651_),
    .A1(_2652_),
    .S(net178),
    .X(_1923_));
 sg13g2_nand2_1 _5343_ (.Y(_1924_),
    .A(_1655_),
    .B(_1923_));
 sg13g2_nor2b_1 _5344_ (.A(net151),
    .B_N(_0989_),
    .Y(_1925_));
 sg13g2_a21o_1 _5345_ (.A2(_0988_),
    .A1(net151),
    .B1(_1925_),
    .X(_1926_));
 sg13g2_nand2_1 _5346_ (.Y(_1927_),
    .A(_1656_),
    .B(_1926_));
 sg13g2_nand2_1 _5347_ (.Y(_1928_),
    .A(_1924_),
    .B(_1927_));
 sg13g2_mux2_1 _5348_ (.A0(_1928_),
    .A1(_1649_),
    .S(net105),
    .X(_1929_));
 sg13g2_nand2_1 _5349_ (.Y(_1930_),
    .A(net148),
    .B(_1615_));
 sg13g2_o21ai_1 _5350_ (.B1(_1930_),
    .Y(_1931_),
    .A1(net116),
    .A2(_1929_));
 sg13g2_mux2_1 _5351_ (.A0(_1659_),
    .A1(_1931_),
    .S(net109),
    .X(_1932_));
 sg13g2_nor2_1 _5352_ (.A(_1478_),
    .B(_1932_),
    .Y(_0202_));
 sg13g2_buf_1 _5353_ (.A(_2737_),
    .X(_1933_));
 sg13g2_mux2_1 _5354_ (.A0(_1656_),
    .A1(_1659_),
    .S(_2728_),
    .X(_1934_));
 sg13g2_nor2_1 _5355_ (.A(net76),
    .B(_1934_),
    .Y(_0203_));
 sg13g2_buf_1 _5356_ (.A(_2592_),
    .X(_1935_));
 sg13g2_mux2_1 _5357_ (.A0(_1347_),
    .A1(_1348_),
    .S(net25),
    .X(_1936_));
 sg13g2_and2_1 _5358_ (.A(net102),
    .B(_1936_),
    .X(_0204_));
 sg13g2_mux2_1 _5359_ (.A0(_1923_),
    .A1(_1926_),
    .S(_1655_),
    .X(_1937_));
 sg13g2_and2_1 _5360_ (.A(net6),
    .B(_1643_),
    .X(_1938_));
 sg13g2_nor2_1 _5361_ (.A(_1643_),
    .B(_1658_),
    .Y(_1939_));
 sg13g2_a21oi_1 _5362_ (.A1(_1937_),
    .A2(_1938_),
    .Y(_1940_),
    .B1(_1939_));
 sg13g2_nand3_1 _5363_ (.B(_1924_),
    .C(_1927_),
    .A(net105),
    .Y(_1941_));
 sg13g2_nor2_1 _5364_ (.A(net6),
    .B(net105),
    .Y(_1942_));
 sg13g2_nor2_1 _5365_ (.A(_1648_),
    .B(_1942_),
    .Y(_1943_));
 sg13g2_a22oi_1 _5366_ (.Y(_1944_),
    .B1(_1941_),
    .B2(_1943_),
    .A2(_1940_),
    .A1(_1648_));
 sg13g2_nor2b_1 _5367_ (.A(_1085_),
    .B_N(_1084_),
    .Y(_1945_));
 sg13g2_a21o_1 _5368_ (.A2(_1083_),
    .A1(_1085_),
    .B1(_1945_),
    .X(_1946_));
 sg13g2_mux2_1 _5369_ (.A0(_1730_),
    .A1(_1946_),
    .S(_1732_),
    .X(_1947_));
 sg13g2_nand3_1 _5370_ (.B(_1728_),
    .C(_1947_),
    .A(net104),
    .Y(_1948_));
 sg13g2_nor2_1 _5371_ (.A(_1719_),
    .B(_1733_),
    .Y(_1949_));
 sg13g2_nor2_1 _5372_ (.A(_1726_),
    .B(_1949_),
    .Y(_1950_));
 sg13g2_mux2_1 _5373_ (.A0(_1946_),
    .A1(_1730_),
    .S(_1732_),
    .X(_1951_));
 sg13g2_mux2_1 _5374_ (.A0(_1725_),
    .A1(_1951_),
    .S(_1720_),
    .X(_1952_));
 sg13g2_a22oi_1 _5375_ (.Y(_1953_),
    .B1(_1952_),
    .B2(_1726_),
    .A2(_1950_),
    .A1(_1948_));
 sg13g2_mux2_1 _5376_ (.A0(_1944_),
    .A1(_1953_),
    .S(_1645_),
    .X(_1954_));
 sg13g2_mux4_1 _5377_ (.S0(_1692_),
    .A0(_1354_),
    .A1(_1372_),
    .A2(_1374_),
    .A3(_1367_),
    .S1(_1355_),
    .X(_1955_));
 sg13g2_buf_1 _5378_ (.A(\g.g_y[6].g_x[1].t.r_d ),
    .X(_1956_));
 sg13g2_inv_1 _5379_ (.Y(_1957_),
    .A(net136));
 sg13g2_nor2b_1 _5380_ (.A(net145),
    .B_N(_1350_),
    .Y(_1958_));
 sg13g2_a21o_1 _5381_ (.A2(_1349_),
    .A1(net145),
    .B1(_1958_),
    .X(_1959_));
 sg13g2_mux2_1 _5382_ (.A0(_2605_),
    .A1(_2602_),
    .S(_2606_),
    .X(_1960_));
 sg13g2_buf_1 _5383_ (.A(\g.g_y[6].g_x[1].t.r_v ),
    .X(_1961_));
 sg13g2_inv_2 _5384_ (.Y(_1962_),
    .A(_1961_));
 sg13g2_mux2_1 _5385_ (.A0(_1959_),
    .A1(_1960_),
    .S(_1962_),
    .X(_1963_));
 sg13g2_mux2_1 _5386_ (.A0(_2648_),
    .A1(\g.g_y[6].g_x[0].t.r_gnl ),
    .S(_2649_),
    .X(_1964_));
 sg13g2_buf_2 _5387_ (.A(\g.g_y[6].g_x[0].t.r_h ),
    .X(_1965_));
 sg13g2_mux2_1 _5388_ (.A0(_2652_),
    .A1(_1964_),
    .S(_1965_),
    .X(_1966_));
 sg13g2_buf_1 _5389_ (.A(_1966_),
    .X(_1967_));
 sg13g2_mux2_1 _5390_ (.A0(_2801_),
    .A1(\g.g_y[6].g_x[2].t.r_gnl ),
    .S(_2802_),
    .X(_1968_));
 sg13g2_buf_1 _5391_ (.A(\g.g_y[6].g_x[2].t.r_h ),
    .X(_1969_));
 sg13g2_mux2_1 _5392_ (.A0(_1968_),
    .A1(_2804_),
    .S(net135),
    .X(_1970_));
 sg13g2_buf_1 _5393_ (.A(\g.g_y[6].g_x[1].t.r_h ),
    .X(_1971_));
 sg13g2_inv_2 _5394_ (.Y(_1972_),
    .A(_1971_));
 sg13g2_mux2_1 _5395_ (.A0(_1967_),
    .A1(_1970_),
    .S(_1972_),
    .X(_1973_));
 sg13g2_nand3_1 _5396_ (.B(_1963_),
    .C(_1973_),
    .A(_1957_),
    .Y(_1974_));
 sg13g2_buf_1 _5397_ (.A(\g.g_y[6].g_x[1].t.out_sc ),
    .X(_1975_));
 sg13g2_inv_1 _5398_ (.Y(_1976_),
    .A(_1975_));
 sg13g2_a21oi_1 _5399_ (.A1(net136),
    .A2(_1976_),
    .Y(_1977_),
    .B1(_1961_));
 sg13g2_or2_1 _5400_ (.X(_1978_),
    .B(_2605_),
    .A(_2606_));
 sg13g2_inv_1 _5401_ (.Y(_1979_),
    .A(_2602_));
 sg13g2_a21oi_1 _5402_ (.A1(_1979_),
    .A2(_2606_),
    .Y(_1980_),
    .B1(_1962_));
 sg13g2_a22oi_1 _5403_ (.Y(_1981_),
    .B1(_1978_),
    .B2(_1980_),
    .A2(_1959_),
    .A1(_1962_));
 sg13g2_or2_1 _5404_ (.X(_1982_),
    .B(_1968_),
    .A(net135));
 sg13g2_nand2b_1 _5405_ (.Y(_1983_),
    .B(_1969_),
    .A_N(_2804_));
 sg13g2_and2_1 _5406_ (.A(_1971_),
    .B(_1983_),
    .X(_1984_));
 sg13g2_a221oi_1 _5407_ (.B2(_1984_),
    .C1(net136),
    .B1(_1982_),
    .A1(_1972_),
    .Y(_1985_),
    .A2(_1967_));
 sg13g2_a21oi_1 _5408_ (.A1(net136),
    .A2(_1981_),
    .Y(_1986_),
    .B1(_1985_));
 sg13g2_a22oi_1 _5409_ (.Y(_1987_),
    .B1(_1986_),
    .B2(_1961_),
    .A2(_1977_),
    .A1(_1974_));
 sg13g2_mux2_1 _5410_ (.A0(_1955_),
    .A1(_1987_),
    .S(_1346_),
    .X(_1988_));
 sg13g2_mux2_1 _5411_ (.A0(_1954_),
    .A1(_1988_),
    .S(_1348_),
    .X(_1989_));
 sg13g2_o21ai_1 _5412_ (.B1(net137),
    .Y(_1990_),
    .A1(_1350_),
    .A2(net57));
 sg13g2_a21oi_1 _5413_ (.A1(net39),
    .A2(_1989_),
    .Y(_0205_),
    .B1(_1990_));
 sg13g2_nand2b_1 _5414_ (.Y(_1991_),
    .B(net145),
    .A_N(_1955_));
 sg13g2_or2_1 _5415_ (.X(_1992_),
    .B(_1987_),
    .A(net145));
 sg13g2_nor2b_1 _5416_ (.A(_1645_),
    .B_N(_1953_),
    .Y(_1993_));
 sg13g2_a221oi_1 _5417_ (.B2(_1992_),
    .C1(_1993_),
    .B1(_1991_),
    .A1(_1645_),
    .Y(_1994_),
    .A2(_1944_));
 sg13g2_o21ai_1 _5418_ (.B1(net137),
    .Y(_1995_),
    .A1(\g.g_y[5].g_x[1].t.r_gnl ),
    .A2(net57));
 sg13g2_a21oi_1 _5419_ (.A1(net39),
    .A2(_1994_),
    .Y(_0206_),
    .B1(_1995_));
 sg13g2_nand2_1 _5420_ (.Y(_1996_),
    .A(_1347_),
    .B(_1747_));
 sg13g2_buf_1 _5421_ (.A(_2589_),
    .X(_1997_));
 sg13g2_o21ai_1 _5422_ (.B1(_1645_),
    .Y(_1998_),
    .A1(net75),
    .A2(net103));
 sg13g2_a21oi_1 _5423_ (.A1(_1996_),
    .A2(_1998_),
    .Y(_0207_),
    .B1(_1859_));
 sg13g2_mux2_1 _5424_ (.A0(_1988_),
    .A1(_1954_),
    .S(_1348_),
    .X(_1999_));
 sg13g2_a22oi_1 _5425_ (.Y(_2000_),
    .B1(net80),
    .B2(_1658_),
    .A2(net51),
    .A1(_1347_));
 sg13g2_o21ai_1 _5426_ (.B1(_2000_),
    .Y(_0208_),
    .A1(net49),
    .A2(_1999_));
 sg13g2_nand2_1 _5427_ (.Y(_2001_),
    .A(_1347_),
    .B(net26));
 sg13g2_o21ai_1 _5428_ (.B1(net145),
    .Y(_2002_),
    .A1(net75),
    .A2(net78));
 sg13g2_a21oi_1 _5429_ (.A1(_2001_),
    .A2(_2002_),
    .Y(_0209_),
    .B1(net77));
 sg13g2_mux2_1 _5430_ (.A0(_1733_),
    .A1(net104),
    .S(net25),
    .X(_2003_));
 sg13g2_and2_1 _5431_ (.A(net102),
    .B(_2003_),
    .X(_0210_));
 sg13g2_nand2_1 _5432_ (.Y(_2004_),
    .A(_1733_),
    .B(_1747_));
 sg13g2_o21ai_1 _5433_ (.B1(_1726_),
    .Y(_2005_),
    .A1(net75),
    .A2(_1749_));
 sg13g2_a21oi_1 _5434_ (.A1(_2004_),
    .A2(_2005_),
    .Y(_0211_),
    .B1(net77));
 sg13g2_mux2_1 _5435_ (.A0(_1951_),
    .A1(_1737_),
    .S(net104),
    .X(_2006_));
 sg13g2_nand2b_1 _5436_ (.Y(_2007_),
    .B(net170),
    .A_N(_1347_));
 sg13g2_o21ai_1 _5437_ (.B1(_2007_),
    .Y(_2008_),
    .A1(net148),
    .A2(_2006_));
 sg13g2_nand2_1 _5438_ (.Y(_2009_),
    .A(net109),
    .B(_2008_));
 sg13g2_o21ai_1 _5439_ (.B1(_2009_),
    .Y(_2010_),
    .A1(_1733_),
    .A2(net121));
 sg13g2_nor2_1 _5440_ (.A(net76),
    .B(_2010_),
    .Y(_0212_));
 sg13g2_nand2_1 _5441_ (.Y(_2011_),
    .A(_1733_),
    .B(net26));
 sg13g2_o21ai_1 _5442_ (.B1(_1732_),
    .Y(_2012_),
    .A1(net75),
    .A2(net78));
 sg13g2_a21oi_1 _5443_ (.A1(_2011_),
    .A2(_2012_),
    .Y(_0213_),
    .B1(net77));
 sg13g2_mux2_1 _5444_ (.A0(_1420_),
    .A1(_1421_),
    .S(net25),
    .X(_2013_));
 sg13g2_and2_1 _5445_ (.A(net102),
    .B(_2013_),
    .X(_0214_));
 sg13g2_nor2_1 _5446_ (.A(_1727_),
    .B(_1949_),
    .Y(_2014_));
 sg13g2_mux2_1 _5447_ (.A0(_1737_),
    .A1(_1951_),
    .S(net104),
    .X(_2015_));
 sg13g2_a22oi_1 _5448_ (.Y(_2016_),
    .B1(_2015_),
    .B2(_1727_),
    .A2(_2014_),
    .A1(_1948_));
 sg13g2_mux2_1 _5449_ (.A0(_1423_),
    .A1(_1722_),
    .S(_1723_),
    .X(_2017_));
 sg13g2_mux2_1 _5450_ (.A0(_1801_),
    .A1(_2017_),
    .S(net138),
    .X(_2018_));
 sg13g2_nand3b_1 _5451_ (.B(_1783_),
    .C(_2018_),
    .Y(_2019_),
    .A_N(_1816_));
 sg13g2_nor2_1 _5452_ (.A(net139),
    .B(_1782_),
    .Y(_2020_));
 sg13g2_nor2_1 _5453_ (.A(net138),
    .B(_2020_),
    .Y(_2021_));
 sg13g2_nor2_1 _5454_ (.A(net139),
    .B(_1801_),
    .Y(_2022_));
 sg13g2_nor2_1 _5455_ (.A(_1796_),
    .B(_2022_),
    .Y(_2023_));
 sg13g2_a22oi_1 _5456_ (.Y(_2024_),
    .B1(_2023_),
    .B2(net138),
    .A2(_2021_),
    .A1(_2019_));
 sg13g2_mux2_1 _5457_ (.A0(_2016_),
    .A1(_2024_),
    .S(_1723_),
    .X(_2025_));
 sg13g2_nand2_1 _5458_ (.Y(_2026_),
    .A(_1448_),
    .B(_1427_));
 sg13g2_o21ai_1 _5459_ (.B1(_2026_),
    .Y(_2027_),
    .A1(net106),
    .A2(_1451_));
 sg13g2_mux2_1 _5460_ (.A0(_1447_),
    .A1(_2027_),
    .S(_1703_),
    .X(_2028_));
 sg13g2_buf_2 _5461_ (.A(\g.g_y[6].g_x[3].t.r_v ),
    .X(_2029_));
 sg13g2_mux2_1 _5462_ (.A0(_1423_),
    .A1(_1422_),
    .S(_1419_),
    .X(_2030_));
 sg13g2_nand2_1 _5463_ (.Y(_2031_),
    .A(_2029_),
    .B(_2030_));
 sg13g2_mux2_1 _5464_ (.A0(_2762_),
    .A1(_2763_),
    .S(_2759_),
    .X(_2032_));
 sg13g2_nand2b_1 _5465_ (.Y(_2033_),
    .B(_2032_),
    .A_N(_2029_));
 sg13g2_buf_2 _5466_ (.A(\g.g_y[6].g_x[4].t.r_h ),
    .X(_2034_));
 sg13g2_mux2_1 _5467_ (.A0(_0404_),
    .A1(\g.g_y[6].g_x[4].t.r_gnl ),
    .S(_0405_),
    .X(_2035_));
 sg13g2_nand2b_1 _5468_ (.Y(_2036_),
    .B(_2034_),
    .A_N(_0407_));
 sg13g2_o21ai_1 _5469_ (.B1(_2036_),
    .Y(_2037_),
    .A1(_2034_),
    .A2(_2035_));
 sg13g2_nor2b_1 _5470_ (.A(net135),
    .B_N(_2804_),
    .Y(_2038_));
 sg13g2_a21oi_1 _5471_ (.A1(net135),
    .A2(_1968_),
    .Y(_2039_),
    .B1(_2038_));
 sg13g2_buf_2 _5472_ (.A(\g.g_y[6].g_x[3].t.r_h ),
    .X(_2040_));
 sg13g2_mux2_1 _5473_ (.A0(_2037_),
    .A1(_2039_),
    .S(_2040_),
    .X(_2041_));
 sg13g2_a21oi_1 _5474_ (.A1(_2031_),
    .A2(_2033_),
    .Y(_2042_),
    .B1(_2041_));
 sg13g2_mux2_1 _5475_ (.A0(_2039_),
    .A1(_2037_),
    .S(_2040_),
    .X(_2043_));
 sg13g2_buf_1 _5476_ (.A(\g.g_y[6].g_x[3].t.out_sc ),
    .X(_2044_));
 sg13g2_inv_1 _5477_ (.Y(_2045_),
    .A(_2044_));
 sg13g2_inv_1 _5478_ (.Y(_2046_),
    .A(_2032_));
 sg13g2_buf_2 _5479_ (.A(\g.g_y[6].g_x[3].t.r_d ),
    .X(_2047_));
 sg13g2_mux4_1 _5480_ (.S0(_2029_),
    .A0(_2042_),
    .A1(_2043_),
    .A2(_2045_),
    .A3(_2046_),
    .S1(_2047_),
    .X(_2048_));
 sg13g2_mux2_1 _5481_ (.A0(_2028_),
    .A1(_2048_),
    .S(_1419_),
    .X(_2049_));
 sg13g2_mux2_1 _5482_ (.A0(_2025_),
    .A1(_2049_),
    .S(_1421_),
    .X(_2050_));
 sg13g2_o21ai_1 _5483_ (.B1(_1824_),
    .Y(_2051_),
    .A1(_1423_),
    .A2(net32));
 sg13g2_a21oi_1 _5484_ (.A1(net36),
    .A2(_2050_),
    .Y(_0215_),
    .B1(_2051_));
 sg13g2_nand2b_1 _5485_ (.Y(_2052_),
    .B(_1723_),
    .A_N(_2016_));
 sg13g2_or2_1 _5486_ (.X(_2053_),
    .B(_2024_),
    .A(_1723_));
 sg13g2_nor2b_1 _5487_ (.A(_1419_),
    .B_N(_2048_),
    .Y(_2054_));
 sg13g2_a221oi_1 _5488_ (.B2(_2053_),
    .C1(_2054_),
    .B1(_2052_),
    .A1(_1419_),
    .Y(_2055_),
    .A2(_2028_));
 sg13g2_o21ai_1 _5489_ (.B1(net137),
    .Y(_2056_),
    .A1(\g.g_y[5].g_x[3].t.r_gnl ),
    .A2(net32));
 sg13g2_a21oi_1 _5490_ (.A1(net36),
    .A2(_2055_),
    .Y(_0216_),
    .B1(_2056_));
 sg13g2_nand2_1 _5491_ (.Y(_2057_),
    .A(_1420_),
    .B(net27));
 sg13g2_o21ai_1 _5492_ (.B1(_1723_),
    .Y(_2058_),
    .A1(net75),
    .A2(_1749_));
 sg13g2_a21oi_1 _5493_ (.A1(_2057_),
    .A2(_2058_),
    .Y(_0217_),
    .B1(net77));
 sg13g2_mux2_1 _5494_ (.A0(_2049_),
    .A1(_2025_),
    .S(_1421_),
    .X(_2059_));
 sg13g2_a22oi_1 _5495_ (.Y(_2060_),
    .B1(net80),
    .B2(_1733_),
    .A2(net51),
    .A1(_1420_));
 sg13g2_o21ai_1 _5496_ (.B1(_2060_),
    .Y(_0218_),
    .A1(net49),
    .A2(_2059_));
 sg13g2_nand2_1 _5497_ (.Y(_2061_),
    .A(_1420_),
    .B(_1844_));
 sg13g2_o21ai_1 _5498_ (.B1(_1419_),
    .Y(_2062_),
    .A1(net75),
    .A2(_1846_));
 sg13g2_buf_1 _5499_ (.A(_2710_),
    .X(_2063_));
 sg13g2_a21oi_1 _5500_ (.A1(_2061_),
    .A2(_2062_),
    .Y(_0219_),
    .B1(net74));
 sg13g2_mux2_1 _5501_ (.A0(_1782_),
    .A1(net139),
    .S(net25),
    .X(_2064_));
 sg13g2_and2_1 _5502_ (.A(net102),
    .B(_2064_),
    .X(_0220_));
 sg13g2_buf_1 _5503_ (.A(net66),
    .X(_2065_));
 sg13g2_nand2_1 _5504_ (.Y(_2066_),
    .A(_1782_),
    .B(net24));
 sg13g2_buf_1 _5505_ (.A(_2699_),
    .X(_2067_));
 sg13g2_o21ai_1 _5506_ (.B1(_1797_),
    .Y(_2068_),
    .A1(_1997_),
    .A2(net101));
 sg13g2_a21oi_1 _5507_ (.A1(_2066_),
    .A2(_2068_),
    .Y(_0221_),
    .B1(_2063_));
 sg13g2_nor2_1 _5508_ (.A(_1782_),
    .B(net110),
    .Y(_2069_));
 sg13g2_and2_1 _5509_ (.A(net115),
    .B(_1420_),
    .X(_2070_));
 sg13g2_a221oi_1 _5510_ (.B2(_1805_),
    .C1(_1794_),
    .B1(_1803_),
    .A1(net138),
    .Y(_2071_),
    .A2(_1801_));
 sg13g2_a221oi_1 _5511_ (.B2(_1786_),
    .C1(_1783_),
    .B1(_1793_),
    .A1(_1789_),
    .Y(_2072_),
    .A2(_1791_));
 sg13g2_nor3_1 _5512_ (.A(net116),
    .B(_2071_),
    .C(_2072_),
    .Y(_2073_));
 sg13g2_nor3_1 _5513_ (.A(_2893_),
    .B(_2070_),
    .C(_2073_),
    .Y(_2074_));
 sg13g2_nor3_1 _5514_ (.A(net92),
    .B(_2069_),
    .C(_2074_),
    .Y(_0222_));
 sg13g2_nand2_1 _5515_ (.Y(_2075_),
    .A(_1782_),
    .B(net26));
 sg13g2_o21ai_1 _5516_ (.B1(_1785_),
    .Y(_2076_),
    .A1(net75),
    .A2(_1846_));
 sg13g2_a21oi_1 _5517_ (.A1(_2075_),
    .A2(_2076_),
    .Y(_0223_),
    .B1(net74));
 sg13g2_mux2_1 _5518_ (.A0(_1498_),
    .A1(_1499_),
    .S(net25),
    .X(_2077_));
 sg13g2_and2_1 _5519_ (.A(net102),
    .B(_2077_),
    .X(_0224_));
 sg13g2_nor2_1 _5520_ (.A(_1811_),
    .B(_2020_),
    .Y(_2078_));
 sg13g2_nor2_1 _5521_ (.A(net139),
    .B(_2017_),
    .Y(_2079_));
 sg13g2_nor2_1 _5522_ (.A(_1796_),
    .B(_2079_),
    .Y(_2080_));
 sg13g2_a22oi_1 _5523_ (.Y(_2081_),
    .B1(_2080_),
    .B2(_1811_),
    .A2(_2078_),
    .A1(_2019_));
 sg13g2_mux2_1 _5524_ (.A0(_1887_),
    .A1(_1877_),
    .S(_1888_),
    .X(_2082_));
 sg13g2_mux4_1 _5525_ (.S0(_1884_),
    .A0(_1875_),
    .A1(_1881_),
    .A2(_1890_),
    .A3(_2082_),
    .S1(_1892_),
    .X(_2083_));
 sg13g2_mux2_1 _5526_ (.A0(_2081_),
    .A1(_2083_),
    .S(_1799_),
    .X(_2084_));
 sg13g2_a21oi_1 _5527_ (.A1(net142),
    .A2(_1545_),
    .Y(_2085_),
    .B1(_1509_));
 sg13g2_nor2b_1 _5528_ (.A(_1554_),
    .B_N(_2085_),
    .Y(_2086_));
 sg13g2_and2_1 _5529_ (.A(_1509_),
    .B(_1549_),
    .X(_2087_));
 sg13g2_or4_1 _5530_ (.A(_1510_),
    .B(net142),
    .C(_1543_),
    .D(_1545_),
    .X(_2088_));
 sg13g2_o21ai_1 _5531_ (.B1(_2088_),
    .Y(_2089_),
    .A1(_2086_),
    .A2(_2087_));
 sg13g2_buf_1 _5532_ (.A(\g.g_y[6].g_x[5].t.r_v ),
    .X(_2090_));
 sg13g2_buf_1 _5533_ (.A(\g.g_y[6].g_x[5].t.r_d ),
    .X(_2091_));
 sg13g2_inv_1 _5534_ (.Y(_2092_),
    .A(_2091_));
 sg13g2_buf_2 _5535_ (.A(\g.g_y[6].g_x[5].t.out_sc ),
    .X(_2093_));
 sg13g2_nor2_1 _5536_ (.A(_2092_),
    .B(_2093_),
    .Y(_2094_));
 sg13g2_nor2_1 _5537_ (.A(_2090_),
    .B(_2094_),
    .Y(_2095_));
 sg13g2_mux2_1 _5538_ (.A0(_0349_),
    .A1(_0348_),
    .S(_0344_),
    .X(_2096_));
 sg13g2_nor2b_1 _5539_ (.A(_1497_),
    .B_N(_1501_),
    .Y(_2097_));
 sg13g2_a21o_1 _5540_ (.A2(_1500_),
    .A1(_1497_),
    .B1(_2097_),
    .X(_2098_));
 sg13g2_mux2_1 _5541_ (.A0(_2096_),
    .A1(_2098_),
    .S(_2090_),
    .X(_2099_));
 sg13g2_mux2_1 _5542_ (.A0(_0536_),
    .A1(\g.g_y[6].g_x[6].t.r_gnl ),
    .S(_0537_),
    .X(_2100_));
 sg13g2_buf_1 _5543_ (.A(\g.g_y[6].g_x[6].t.r_h ),
    .X(_2101_));
 sg13g2_inv_1 _5544_ (.Y(_2102_),
    .A(net134));
 sg13g2_mux2_1 _5545_ (.A0(_0539_),
    .A1(_2100_),
    .S(_2102_),
    .X(_2103_));
 sg13g2_mux2_1 _5546_ (.A0(_0407_),
    .A1(_2035_),
    .S(_2034_),
    .X(_2104_));
 sg13g2_buf_1 _5547_ (.A(\g.g_y[6].g_x[5].t.r_h ),
    .X(_2105_));
 sg13g2_mux2_1 _5548_ (.A0(_2103_),
    .A1(_2104_),
    .S(net133),
    .X(_2106_));
 sg13g2_nand3_1 _5549_ (.B(_2099_),
    .C(_2106_),
    .A(_2092_),
    .Y(_2107_));
 sg13g2_inv_1 _5550_ (.Y(_2108_),
    .A(_2090_));
 sg13g2_inv_1 _5551_ (.Y(_2109_),
    .A(_2034_));
 sg13g2_or2_1 _5552_ (.X(_2110_),
    .B(_2035_),
    .A(_2109_));
 sg13g2_inv_1 _5553_ (.Y(_2111_),
    .A(_0407_));
 sg13g2_a21oi_1 _5554_ (.A1(_2111_),
    .A2(_2109_),
    .Y(_2112_),
    .B1(net133));
 sg13g2_a221oi_1 _5555_ (.B2(_2112_),
    .C1(_2091_),
    .B1(_2110_),
    .A1(net133),
    .Y(_2113_),
    .A2(_2103_));
 sg13g2_nand2b_1 _5556_ (.Y(_2114_),
    .B(_0344_),
    .A_N(_0348_));
 sg13g2_inv_1 _5557_ (.Y(_2115_),
    .A(_0349_));
 sg13g2_a21oi_1 _5558_ (.A1(_2115_),
    .A2(_0343_),
    .Y(_2116_),
    .B1(_2108_));
 sg13g2_a221oi_1 _5559_ (.B2(_2108_),
    .C1(_2092_),
    .B1(_2098_),
    .A1(_2114_),
    .Y(_2117_),
    .A2(_2116_));
 sg13g2_nor3_1 _5560_ (.A(_2108_),
    .B(_2113_),
    .C(_2117_),
    .Y(_2118_));
 sg13g2_a21oi_1 _5561_ (.A1(_2095_),
    .A2(_2107_),
    .Y(_2119_),
    .B1(_2118_));
 sg13g2_mux2_1 _5562_ (.A0(_2089_),
    .A1(_2119_),
    .S(_1497_),
    .X(_2120_));
 sg13g2_mux2_1 _5563_ (.A0(_2084_),
    .A1(_2120_),
    .S(_1499_),
    .X(_2121_));
 sg13g2_o21ai_1 _5564_ (.B1(net137),
    .Y(_2122_),
    .A1(_1501_),
    .A2(_0647_));
 sg13g2_a21oi_1 _5565_ (.A1(net39),
    .A2(_2121_),
    .Y(_0225_),
    .B1(_2122_));
 sg13g2_inv_1 _5566_ (.Y(_2123_),
    .A(_1497_));
 sg13g2_nand2_1 _5567_ (.Y(_2124_),
    .A(_1548_),
    .B(_2087_));
 sg13g2_nor2_1 _5568_ (.A(_2123_),
    .B(_2086_),
    .Y(_2125_));
 sg13g2_mux2_1 _5569_ (.A0(_2083_),
    .A1(_2081_),
    .S(_1799_),
    .X(_2126_));
 sg13g2_a221oi_1 _5570_ (.B2(_2125_),
    .C1(_2126_),
    .B1(_2124_),
    .A1(_2123_),
    .Y(_2127_),
    .A2(_2119_));
 sg13g2_o21ai_1 _5571_ (.B1(_1824_),
    .Y(_2128_),
    .A1(\g.g_y[5].g_x[5].t.r_gnl ),
    .A2(net57));
 sg13g2_a21oi_1 _5572_ (.A1(net39),
    .A2(_2127_),
    .Y(_0226_),
    .B1(_2128_));
 sg13g2_nand2_1 _5573_ (.Y(_2129_),
    .A(_1498_),
    .B(net24));
 sg13g2_o21ai_1 _5574_ (.B1(_1799_),
    .Y(_2130_),
    .A1(_1997_),
    .A2(net101));
 sg13g2_a21oi_1 _5575_ (.A1(_2129_),
    .A2(_2130_),
    .Y(_0227_),
    .B1(net74));
 sg13g2_mux2_1 _5576_ (.A0(_2120_),
    .A1(_2084_),
    .S(_1499_),
    .X(_2131_));
 sg13g2_a22oi_1 _5577_ (.Y(_2132_),
    .B1(net80),
    .B2(_1782_),
    .A2(net51),
    .A1(_1498_));
 sg13g2_o21ai_1 _5578_ (.B1(_2132_),
    .Y(_0228_),
    .A1(net49),
    .A2(_2131_));
 sg13g2_nand2_1 _5579_ (.Y(_2133_),
    .A(_1498_),
    .B(net26));
 sg13g2_o21ai_1 _5580_ (.B1(_1497_),
    .Y(_2134_),
    .A1(net75),
    .A2(net78));
 sg13g2_a21oi_1 _5581_ (.A1(_2133_),
    .A2(_2134_),
    .Y(_0229_),
    .B1(net74));
 sg13g2_nor2_1 _5582_ (.A(_1875_),
    .B(net28),
    .Y(_2135_));
 sg13g2_a21oi_1 _5583_ (.A1(_1892_),
    .A2(net41),
    .Y(_2136_),
    .B1(_2135_));
 sg13g2_nor2_1 _5584_ (.A(net76),
    .B(_2136_),
    .Y(_0230_));
 sg13g2_nand2_1 _5585_ (.Y(_2137_),
    .A(_1874_),
    .B(net24));
 sg13g2_buf_1 _5586_ (.A(_2589_),
    .X(_2138_));
 sg13g2_o21ai_1 _5587_ (.B1(_1884_),
    .Y(_2139_),
    .A1(net73),
    .A2(net101));
 sg13g2_a21oi_1 _5588_ (.A1(_2137_),
    .A2(_2139_),
    .Y(_0231_),
    .B1(net74));
 sg13g2_nand2b_1 _5589_ (.Y(_2140_),
    .B(_1874_),
    .A_N(_1037_));
 sg13g2_mux2_1 _5590_ (.A0(_1891_),
    .A1(_2082_),
    .S(_1893_),
    .X(_2141_));
 sg13g2_nand2_1 _5591_ (.Y(_2142_),
    .A(net148),
    .B(_1498_));
 sg13g2_o21ai_1 _5592_ (.B1(_2142_),
    .Y(_2143_),
    .A1(net116),
    .A2(_2141_));
 sg13g2_nand2_1 _5593_ (.Y(_2144_),
    .A(net125),
    .B(_2143_));
 sg13g2_a21oi_1 _5594_ (.A1(_2140_),
    .A2(_2144_),
    .Y(_0232_),
    .B1(net74));
 sg13g2_nand2_1 _5595_ (.Y(_2145_),
    .A(_1874_),
    .B(_1844_));
 sg13g2_o21ai_1 _5596_ (.B1(_1888_),
    .Y(_2146_),
    .A1(net73),
    .A2(net78));
 sg13g2_a21oi_1 _5597_ (.A1(_2145_),
    .A2(_2146_),
    .Y(_0233_),
    .B1(net74));
 sg13g2_mux2_1 _5598_ (.A0(_1605_),
    .A1(_1606_),
    .S(net25),
    .X(_2147_));
 sg13g2_and2_1 _5599_ (.A(_1767_),
    .B(_2147_),
    .X(_0234_));
 sg13g2_mux4_1 _5600_ (.S0(_1892_),
    .A0(_1883_),
    .A1(_2082_),
    .A2(_1875_),
    .A3(_1890_),
    .S1(_1884_),
    .X(_2148_));
 sg13g2_nand3_1 _5601_ (.B(_1647_),
    .C(_1937_),
    .A(net105),
    .Y(_2149_));
 sg13g2_nor2_1 _5602_ (.A(_1648_),
    .B(_1939_),
    .Y(_2150_));
 sg13g2_o21ai_1 _5603_ (.B1(_1648_),
    .Y(_2151_),
    .A1(_1643_),
    .A2(_1647_));
 sg13g2_inv_1 _5604_ (.Y(_2152_),
    .A(_2151_));
 sg13g2_a22oi_1 _5605_ (.Y(_2153_),
    .B1(_2152_),
    .B2(_1941_),
    .A2(_2150_),
    .A1(_2149_));
 sg13g2_mux2_1 _5606_ (.A0(_2148_),
    .A1(_2153_),
    .S(_1878_),
    .X(_2154_));
 sg13g2_mux4_1 _5607_ (.S0(net140),
    .A0(_1602_),
    .A1(_1866_),
    .A2(_1868_),
    .A3(_1615_),
    .S1(_1611_),
    .X(_2155_));
 sg13g2_buf_2 _5608_ (.A(\g.g_y[6].g_x[7].t.r_h ),
    .X(_2156_));
 sg13g2_inv_1 _5609_ (.Y(_2157_),
    .A(_2156_));
 sg13g2_inv_1 _5610_ (.Y(_2158_),
    .A(_1965_));
 sg13g2_mux2_1 _5611_ (.A0(_2652_),
    .A1(_1964_),
    .S(_2158_),
    .X(_2159_));
 sg13g2_nand2_1 _5612_ (.Y(_2160_),
    .A(_2157_),
    .B(_2159_));
 sg13g2_or2_1 _5613_ (.X(_2161_),
    .B(net134),
    .A(_0539_));
 sg13g2_o21ai_1 _5614_ (.B1(_2161_),
    .Y(_2162_),
    .A1(_2102_),
    .A2(_2100_));
 sg13g2_or2_1 _5615_ (.X(_2163_),
    .B(_2162_),
    .A(_2157_));
 sg13g2_nor2b_1 _5616_ (.A(_1604_),
    .B_N(_1608_),
    .Y(_2164_));
 sg13g2_a21oi_1 _5617_ (.A1(_1604_),
    .A2(_1607_),
    .Y(_2165_),
    .B1(_2164_));
 sg13g2_buf_2 _5618_ (.A(\g.g_y[6].g_x[7].t.r_v ),
    .X(_2166_));
 sg13g2_nand2b_1 _5619_ (.Y(_2167_),
    .B(_0511_),
    .A_N(_0515_));
 sg13g2_o21ai_1 _5620_ (.B1(_2167_),
    .Y(_2168_),
    .A1(_0511_),
    .A2(_0514_));
 sg13g2_nor2b_1 _5621_ (.A(_2166_),
    .B_N(_2168_),
    .Y(_2169_));
 sg13g2_a221oi_1 _5622_ (.B2(_2166_),
    .C1(_2169_),
    .B1(_2165_),
    .A1(_2160_),
    .Y(_2170_),
    .A2(_2163_));
 sg13g2_and2_1 _5623_ (.A(_2156_),
    .B(_2159_),
    .X(_2171_));
 sg13g2_nor2_1 _5624_ (.A(_2156_),
    .B(_2162_),
    .Y(_2172_));
 sg13g2_nor2_1 _5625_ (.A(_2171_),
    .B(_2172_),
    .Y(_2173_));
 sg13g2_inv_1 _5626_ (.Y(_2174_),
    .A(\g.g_y[6].g_x[7].t.out_sc ));
 sg13g2_buf_2 _5627_ (.A(\g.g_y[6].g_x[7].t.r_d ),
    .X(_2175_));
 sg13g2_mux4_1 _5628_ (.S0(_2166_),
    .A0(_2170_),
    .A1(_2173_),
    .A2(_2174_),
    .A3(_2168_),
    .S1(_2175_),
    .X(_2176_));
 sg13g2_mux2_1 _5629_ (.A0(_2155_),
    .A1(_2176_),
    .S(_1604_),
    .X(_2177_));
 sg13g2_mux2_1 _5630_ (.A0(_2154_),
    .A1(_2177_),
    .S(_1606_),
    .X(_2178_));
 sg13g2_buf_1 _5631_ (.A(_2581_),
    .X(_2179_));
 sg13g2_o21ai_1 _5632_ (.B1(net132),
    .Y(_2180_),
    .A1(_1608_),
    .A2(_0910_));
 sg13g2_a21oi_1 _5633_ (.A1(net36),
    .A2(_2178_),
    .Y(_0235_),
    .B1(_2180_));
 sg13g2_nand2b_1 _5634_ (.Y(_2181_),
    .B(_1604_),
    .A_N(_2155_));
 sg13g2_or2_1 _5635_ (.X(_2182_),
    .B(_2176_),
    .A(_1604_));
 sg13g2_nor2b_1 _5636_ (.A(_1878_),
    .B_N(_2153_),
    .Y(_2183_));
 sg13g2_a221oi_1 _5637_ (.B2(_2182_),
    .C1(_2183_),
    .B1(_2181_),
    .A1(_1878_),
    .Y(_2184_),
    .A2(_2148_));
 sg13g2_o21ai_1 _5638_ (.B1(net132),
    .Y(_2185_),
    .A1(\g.g_y[5].g_x[7].t.r_gnl ),
    .A2(_0910_));
 sg13g2_a21oi_1 _5639_ (.A1(net36),
    .A2(_2184_),
    .Y(_0236_),
    .B1(_2185_));
 sg13g2_nand2_1 _5640_ (.Y(_2186_),
    .A(_1605_),
    .B(net24));
 sg13g2_o21ai_1 _5641_ (.B1(_1878_),
    .Y(_2187_),
    .A1(net73),
    .A2(net101));
 sg13g2_a21oi_1 _5642_ (.A1(_2186_),
    .A2(_2187_),
    .Y(_0237_),
    .B1(_2063_));
 sg13g2_mux2_1 _5643_ (.A0(_2177_),
    .A1(_2154_),
    .S(_1606_),
    .X(_2188_));
 sg13g2_a22oi_1 _5644_ (.Y(_2189_),
    .B1(net80),
    .B2(_1874_),
    .A2(_1471_),
    .A1(_1605_));
 sg13g2_o21ai_1 _5645_ (.B1(_2189_),
    .Y(_0238_),
    .A1(net49),
    .A2(_2188_));
 sg13g2_nand2_1 _5646_ (.Y(_2190_),
    .A(_1605_),
    .B(net26));
 sg13g2_o21ai_1 _5647_ (.B1(_1604_),
    .Y(_2191_),
    .A1(net73),
    .A2(net78));
 sg13g2_a21oi_1 _5648_ (.A1(_2190_),
    .A2(_2191_),
    .Y(_0239_),
    .B1(net74));
 sg13g2_mux2_1 _5649_ (.A0(_2648_),
    .A1(_2649_),
    .S(_1935_),
    .X(_2192_));
 sg13g2_and2_1 _5650_ (.A(_1767_),
    .B(_2192_),
    .X(_0240_));
 sg13g2_mux2_1 _5651_ (.A0(_0633_),
    .A1(_2617_),
    .S(_2686_),
    .X(_2193_));
 sg13g2_buf_1 _5652_ (.A(_2193_),
    .X(_2194_));
 sg13g2_mux2_1 _5653_ (.A0(_2645_),
    .A1(_2194_),
    .S(net130),
    .X(_2195_));
 sg13g2_nand3b_1 _5654_ (.B(_2657_),
    .C(_2194_),
    .Y(_2196_),
    .A_N(net130));
 sg13g2_nor2_1 _5655_ (.A(_2655_),
    .B(_2660_),
    .Y(_2197_));
 sg13g2_a22oi_1 _5656_ (.Y(_2198_),
    .B1(_2196_),
    .B2(_2197_),
    .A2(_2195_),
    .A1(_2655_));
 sg13g2_a21oi_1 _5657_ (.A1(net151),
    .A2(_0988_),
    .Y(_2199_),
    .B1(_1925_));
 sg13g2_a21oi_1 _5658_ (.A1(net105),
    .A2(_2199_),
    .Y(_2200_),
    .B1(_1655_));
 sg13g2_nor2_1 _5659_ (.A(_1643_),
    .B(_2199_),
    .Y(_2201_));
 sg13g2_a22oi_1 _5660_ (.Y(_2202_),
    .B1(_1660_),
    .B2(_2201_),
    .A2(_1659_),
    .A1(_1652_));
 sg13g2_a221oi_1 _5661_ (.B2(_1655_),
    .C1(_2647_),
    .B1(_2202_),
    .A1(_1651_),
    .Y(_2203_),
    .A2(_2200_));
 sg13g2_a21oi_1 _5662_ (.A1(net178),
    .A2(_2198_),
    .Y(_2204_),
    .B1(_2203_));
 sg13g2_nand2_1 _5663_ (.Y(_2205_),
    .A(_1963_),
    .B(_1973_));
 sg13g2_nand2_1 _5664_ (.Y(_2206_),
    .A(_1982_),
    .B(_1983_));
 sg13g2_nand2_1 _5665_ (.Y(_2207_),
    .A(_1972_),
    .B(_1967_));
 sg13g2_o21ai_1 _5666_ (.B1(_2207_),
    .Y(_2208_),
    .A1(_1972_),
    .A2(_2206_));
 sg13g2_a21oi_1 _5667_ (.A1(net145),
    .A2(_1349_),
    .Y(_2209_),
    .B1(_1958_));
 sg13g2_nand2_1 _5668_ (.Y(_2210_),
    .A(_1961_),
    .B(_1960_));
 sg13g2_o21ai_1 _5669_ (.B1(_2210_),
    .Y(_2211_),
    .A1(_1961_),
    .A2(_2209_));
 sg13g2_mux4_1 _5670_ (.S0(net136),
    .A0(_1975_),
    .A1(_2205_),
    .A2(_2208_),
    .A3(_2211_),
    .S1(_1971_),
    .X(_2212_));
 sg13g2_or2_1 _5671_ (.X(_2213_),
    .B(_2212_),
    .A(_2158_));
 sg13g2_nor2_1 _5672_ (.A(_1965_),
    .B(net7),
    .Y(_2214_));
 sg13g2_nor2_1 _5673_ (.A(_2649_),
    .B(_2214_),
    .Y(_2215_));
 sg13g2_a22oi_1 _5674_ (.Y(_2216_),
    .B1(_2213_),
    .B2(_2215_),
    .A2(_2204_),
    .A1(_2649_));
 sg13g2_o21ai_1 _5675_ (.B1(net132),
    .Y(_2217_),
    .A1(_2652_),
    .A2(_2753_));
 sg13g2_a21oi_1 _5676_ (.A1(_2754_),
    .A2(_2216_),
    .Y(_0241_),
    .B1(_2217_));
 sg13g2_nor2_1 _5677_ (.A(_2158_),
    .B(net7),
    .Y(_2218_));
 sg13g2_nor2_1 _5678_ (.A(_1965_),
    .B(_2212_),
    .Y(_2219_));
 sg13g2_a22oi_1 _5679_ (.Y(_2220_),
    .B1(_2202_),
    .B2(_1655_),
    .A2(_2200_),
    .A1(_1651_));
 sg13g2_mux2_1 _5680_ (.A0(_2198_),
    .A1(_2220_),
    .S(net178),
    .X(_2221_));
 sg13g2_nor4_1 _5681_ (.A(_0596_),
    .B(_2218_),
    .C(_2219_),
    .D(_2221_),
    .Y(_2222_));
 sg13g2_o21ai_1 _5682_ (.B1(net177),
    .Y(_2223_),
    .A1(\g.g_y[6].g_x[0].t.r_gnl ),
    .A2(_2873_));
 sg13g2_nor2_1 _5683_ (.A(_2222_),
    .B(_2223_),
    .Y(_0242_));
 sg13g2_nand2_1 _5684_ (.Y(_2224_),
    .A(_2648_),
    .B(net24));
 sg13g2_o21ai_1 _5685_ (.B1(_1965_),
    .Y(_2225_),
    .A1(net73),
    .A2(net101));
 sg13g2_buf_1 _5686_ (.A(_2710_),
    .X(_2226_));
 sg13g2_a21oi_1 _5687_ (.A1(_2224_),
    .A2(_2225_),
    .Y(_0243_),
    .B1(net72));
 sg13g2_inv_1 _5688_ (.Y(_2227_),
    .A(_2649_));
 sg13g2_nor2_1 _5689_ (.A(_2227_),
    .B(_2214_),
    .Y(_2228_));
 sg13g2_a22oi_1 _5690_ (.Y(_2229_),
    .B1(_2213_),
    .B2(_2228_),
    .A2(_2204_),
    .A1(_2227_));
 sg13g2_a22oi_1 _5691_ (.Y(_2230_),
    .B1(_1562_),
    .B2(_1605_),
    .A2(_1471_),
    .A1(_2648_));
 sg13g2_o21ai_1 _5692_ (.B1(_2230_),
    .Y(_0244_),
    .A1(net49),
    .A2(_2229_));
 sg13g2_buf_1 _5693_ (.A(net61),
    .X(_2231_));
 sg13g2_nand2_1 _5694_ (.Y(_2232_),
    .A(_2648_),
    .B(net23));
 sg13g2_buf_1 _5695_ (.A(_2731_),
    .X(_2233_));
 sg13g2_o21ai_1 _5696_ (.B1(net178),
    .Y(_2234_),
    .A1(net73),
    .A2(net71));
 sg13g2_a21oi_1 _5697_ (.A1(_2232_),
    .A2(_2234_),
    .Y(_0245_),
    .B1(net72));
 sg13g2_nor2_1 _5698_ (.A(_1976_),
    .B(net28),
    .Y(_2235_));
 sg13g2_a21oi_1 _5699_ (.A1(net136),
    .A2(net41),
    .Y(_2236_),
    .B1(_2235_));
 sg13g2_nor2_1 _5700_ (.A(net76),
    .B(_2236_),
    .Y(_0246_));
 sg13g2_mux2_1 _5701_ (.A0(_1972_),
    .A1(_1976_),
    .S(_2701_),
    .X(_2237_));
 sg13g2_nor2_1 _5702_ (.A(net76),
    .B(_2237_),
    .Y(_0247_));
 sg13g2_mux2_1 _5703_ (.A0(_2208_),
    .A1(_2211_),
    .S(_1957_),
    .X(_2238_));
 sg13g2_nand2b_1 _5704_ (.Y(_2239_),
    .B(net148),
    .A_N(_2648_));
 sg13g2_o21ai_1 _5705_ (.B1(_2239_),
    .Y(_2240_),
    .A1(_0614_),
    .A2(_2238_));
 sg13g2_mux2_1 _5706_ (.A0(_1976_),
    .A1(_2240_),
    .S(net109),
    .X(_2241_));
 sg13g2_nor2_1 _5707_ (.A(net76),
    .B(_2241_),
    .Y(_0248_));
 sg13g2_mux2_1 _5708_ (.A0(_1962_),
    .A1(_1976_),
    .S(net61),
    .X(_2242_));
 sg13g2_nor2_1 _5709_ (.A(_1933_),
    .B(_2242_),
    .Y(_0249_));
 sg13g2_buf_1 _5710_ (.A(_2582_),
    .X(_2243_));
 sg13g2_mux2_1 _5711_ (.A0(_2801_),
    .A1(_2802_),
    .S(net25),
    .X(_2244_));
 sg13g2_and2_1 _5712_ (.A(net100),
    .B(_2244_),
    .X(_0250_));
 sg13g2_and2_1 _5713_ (.A(_1971_),
    .B(_1967_),
    .X(_2245_));
 sg13g2_a22oi_1 _5714_ (.Y(_2246_),
    .B1(_1981_),
    .B2(_1972_),
    .A2(_2245_),
    .A1(_1963_));
 sg13g2_a21oi_1 _5715_ (.A1(_1971_),
    .A2(_1975_),
    .Y(_2247_),
    .B1(net136));
 sg13g2_nand2_1 _5716_ (.Y(_2248_),
    .A(_2207_),
    .B(_2247_));
 sg13g2_o21ai_1 _5717_ (.B1(_2248_),
    .Y(_2249_),
    .A1(_1957_),
    .A2(_2246_));
 sg13g2_inv_1 _5718_ (.Y(_2250_),
    .A(_2030_));
 sg13g2_mux2_1 _5719_ (.A0(_2250_),
    .A1(_2046_),
    .S(_2029_),
    .X(_2251_));
 sg13g2_mux4_1 _5720_ (.S0(_2040_),
    .A0(_2045_),
    .A1(_2037_),
    .A2(_2042_),
    .A3(_2251_),
    .S1(_2047_),
    .X(_2252_));
 sg13g2_mux2_1 _5721_ (.A0(_2249_),
    .A1(_2252_),
    .S(net135),
    .X(_2253_));
 sg13g2_a21oi_1 _5722_ (.A1(_1085_),
    .A2(_1083_),
    .Y(_2254_),
    .B1(_1945_));
 sg13g2_nor2_1 _5723_ (.A(net104),
    .B(_2254_),
    .Y(_2255_));
 sg13g2_a21oi_1 _5724_ (.A1(_1728_),
    .A2(_2255_),
    .Y(_2256_),
    .B1(_1734_));
 sg13g2_a21oi_1 _5725_ (.A1(net104),
    .A2(_2254_),
    .Y(_2257_),
    .B1(_1732_));
 sg13g2_or2_1 _5726_ (.X(_2258_),
    .B(_1737_),
    .A(_1720_));
 sg13g2_a22oi_1 _5727_ (.Y(_2259_),
    .B1(_2257_),
    .B2(_2258_),
    .A2(_2256_),
    .A1(_1732_));
 sg13g2_mux2_1 _5728_ (.A0(_2833_),
    .A1(_2824_),
    .S(_2812_),
    .X(_2260_));
 sg13g2_mux2_1 _5729_ (.A0(_2259_),
    .A1(_2260_),
    .S(_2800_),
    .X(_2261_));
 sg13g2_mux2_1 _5730_ (.A0(_2253_),
    .A1(_2261_),
    .S(_2802_),
    .X(_2262_));
 sg13g2_o21ai_1 _5731_ (.B1(net132),
    .Y(_2263_),
    .A1(_2804_),
    .A2(_2598_));
 sg13g2_a21oi_1 _5732_ (.A1(_2599_),
    .A2(_2262_),
    .Y(_0251_),
    .B1(_2263_));
 sg13g2_nand2b_1 _5733_ (.Y(_2264_),
    .B(_2800_),
    .A_N(_2259_));
 sg13g2_or2_1 _5734_ (.X(_2265_),
    .B(_2260_),
    .A(_2800_));
 sg13g2_nor2b_1 _5735_ (.A(net135),
    .B_N(_2252_),
    .Y(_2266_));
 sg13g2_a221oi_1 _5736_ (.B2(_2265_),
    .C1(_2266_),
    .B1(_2264_),
    .A1(net135),
    .Y(_2267_),
    .A2(_2249_));
 sg13g2_o21ai_1 _5737_ (.B1(net132),
    .Y(_2268_),
    .A1(\g.g_y[6].g_x[2].t.r_gnl ),
    .A2(_2598_));
 sg13g2_a21oi_1 _5738_ (.A1(_2599_),
    .A2(_2267_),
    .Y(_0252_),
    .B1(_2268_));
 sg13g2_nand2_1 _5739_ (.Y(_2269_),
    .A(_2801_),
    .B(net24));
 sg13g2_o21ai_1 _5740_ (.B1(net135),
    .Y(_2270_),
    .A1(net73),
    .A2(net101));
 sg13g2_a21oi_1 _5741_ (.A1(_2269_),
    .A2(_2270_),
    .Y(_0253_),
    .B1(net72));
 sg13g2_mux2_1 _5742_ (.A0(_2261_),
    .A1(_2253_),
    .S(_2802_),
    .X(_2271_));
 sg13g2_a22oi_1 _5743_ (.Y(_2272_),
    .B1(_1562_),
    .B2(_1975_),
    .A2(_0815_),
    .A1(_2801_));
 sg13g2_o21ai_1 _5744_ (.B1(_2272_),
    .Y(_0254_),
    .A1(_1632_),
    .A2(_2271_));
 sg13g2_nand2_1 _5745_ (.Y(_2273_),
    .A(_2801_),
    .B(net23));
 sg13g2_o21ai_1 _5746_ (.B1(_2800_),
    .Y(_2274_),
    .A1(net73),
    .A2(net71));
 sg13g2_a21oi_1 _5747_ (.A1(_2273_),
    .A2(_2274_),
    .Y(_0255_),
    .B1(net72));
 sg13g2_nor2_1 _5748_ (.A(_2045_),
    .B(_1394_),
    .Y(_2275_));
 sg13g2_a21oi_1 _5749_ (.A1(_2047_),
    .A2(net41),
    .Y(_2276_),
    .B1(_2275_));
 sg13g2_nor2_1 _5750_ (.A(net76),
    .B(_2276_),
    .Y(_0256_));
 sg13g2_nand2_1 _5751_ (.Y(_2277_),
    .A(_2044_),
    .B(net24));
 sg13g2_o21ai_1 _5752_ (.B1(_2040_),
    .Y(_2278_),
    .A1(_2138_),
    .A2(net101));
 sg13g2_a21oi_1 _5753_ (.A1(_2277_),
    .A2(_2278_),
    .Y(_0257_),
    .B1(net72));
 sg13g2_nor2_1 _5754_ (.A(_2044_),
    .B(net110),
    .Y(_2279_));
 sg13g2_mux2_1 _5755_ (.A0(_2251_),
    .A1(_2043_),
    .S(_2047_),
    .X(_2280_));
 sg13g2_nand2_1 _5756_ (.Y(_2281_),
    .A(_0324_),
    .B(_2801_));
 sg13g2_o21ai_1 _5757_ (.B1(_2281_),
    .Y(_2282_),
    .A1(net120),
    .A2(_2280_));
 sg13g2_nor2b_1 _5758_ (.A(_2282_),
    .B_N(net109),
    .Y(_2283_));
 sg13g2_nor3_1 _5759_ (.A(net92),
    .B(_2279_),
    .C(_2283_),
    .Y(_0258_));
 sg13g2_nand2_1 _5760_ (.Y(_2284_),
    .A(_2044_),
    .B(net23));
 sg13g2_o21ai_1 _5761_ (.B1(_2029_),
    .Y(_2285_),
    .A1(_2138_),
    .A2(net71));
 sg13g2_a21oi_1 _5762_ (.A1(_2284_),
    .A2(_2285_),
    .Y(_0259_),
    .B1(net72));
 sg13g2_mux2_1 _5763_ (.A0(_0404_),
    .A1(_0405_),
    .S(net25),
    .X(_2286_));
 sg13g2_and2_1 _5764_ (.A(net100),
    .B(_2286_),
    .X(_0260_));
 sg13g2_nor2_1 _5765_ (.A(_2113_),
    .B(_2117_),
    .Y(_2287_));
 sg13g2_nand3_1 _5766_ (.B(_2099_),
    .C(_2106_),
    .A(_2091_),
    .Y(_2288_));
 sg13g2_nor2_1 _5767_ (.A(_2091_),
    .B(_2093_),
    .Y(_2289_));
 sg13g2_nor2_1 _5768_ (.A(net133),
    .B(_2289_),
    .Y(_2290_));
 sg13g2_a22oi_1 _5769_ (.Y(_2291_),
    .B1(_2288_),
    .B2(_2290_),
    .A2(_2287_),
    .A1(net133));
 sg13g2_mux4_1 _5770_ (.S0(_2047_),
    .A0(_2039_),
    .A1(_2251_),
    .A2(_2045_),
    .A3(_2042_),
    .S1(_2040_),
    .X(_2292_));
 sg13g2_mux2_1 _5771_ (.A0(_2291_),
    .A1(_2292_),
    .S(_2109_),
    .X(_2293_));
 sg13g2_nand3_1 _5772_ (.B(_1793_),
    .C(_2018_),
    .A(_1794_),
    .Y(_2294_));
 sg13g2_and2_1 _5773_ (.A(_1785_),
    .B(_1784_),
    .X(_2295_));
 sg13g2_or2_1 _5774_ (.X(_2296_),
    .B(_1173_),
    .A(_1169_));
 sg13g2_o21ai_1 _5775_ (.B1(_2296_),
    .Y(_2297_),
    .A1(_1174_),
    .A2(_1172_));
 sg13g2_a21oi_1 _5776_ (.A1(net139),
    .A2(_2297_),
    .Y(_2298_),
    .B1(_1806_));
 sg13g2_a22oi_1 _5777_ (.Y(_2299_),
    .B1(_2298_),
    .B2(_1786_),
    .A2(_2295_),
    .A1(_2294_));
 sg13g2_mux2_1 _5778_ (.A0(_2780_),
    .A1(_0426_),
    .S(_0451_),
    .X(_2300_));
 sg13g2_buf_1 _5779_ (.A(_2300_),
    .X(_2301_));
 sg13g2_nand3b_1 _5780_ (.B(_0402_),
    .C(_2301_),
    .Y(_2302_),
    .A_N(net119));
 sg13g2_nor2_1 _5781_ (.A(net166),
    .B(_0399_),
    .Y(_2303_));
 sg13g2_mux2_1 _5782_ (.A0(_0396_),
    .A1(_2301_),
    .S(_0387_),
    .X(_2304_));
 sg13g2_a22oi_1 _5783_ (.Y(_2305_),
    .B1(_2304_),
    .B2(net166),
    .A2(_2303_),
    .A1(_2302_));
 sg13g2_mux2_1 _5784_ (.A0(_2299_),
    .A1(_2305_),
    .S(_0403_),
    .X(_2306_));
 sg13g2_mux2_1 _5785_ (.A0(_2293_),
    .A1(_2306_),
    .S(_0405_),
    .X(_2307_));
 sg13g2_o21ai_1 _5786_ (.B1(net132),
    .Y(_2308_),
    .A1(_0407_),
    .A2(_2753_));
 sg13g2_a21oi_1 _5787_ (.A1(_2754_),
    .A2(_2307_),
    .Y(_0261_),
    .B1(_2308_));
 sg13g2_mux2_1 _5788_ (.A0(_2291_),
    .A1(_2292_),
    .S(_2034_),
    .X(_2309_));
 sg13g2_mux2_1 _5789_ (.A0(_2305_),
    .A1(_2299_),
    .S(_0403_),
    .X(_2310_));
 sg13g2_nor3_1 _5790_ (.A(_0596_),
    .B(_2309_),
    .C(_2310_),
    .Y(_2311_));
 sg13g2_o21ai_1 _5791_ (.B1(net177),
    .Y(_2312_),
    .A1(\g.g_y[6].g_x[4].t.r_gnl ),
    .A2(_2873_));
 sg13g2_nor2_1 _5792_ (.A(_2311_),
    .B(_2312_),
    .Y(_0262_));
 sg13g2_nand2_1 _5793_ (.Y(_2313_),
    .A(_0404_),
    .B(net24));
 sg13g2_buf_1 _5794_ (.A(_2589_),
    .X(_2314_));
 sg13g2_o21ai_1 _5795_ (.B1(_2034_),
    .Y(_2315_),
    .A1(net70),
    .A2(net101));
 sg13g2_a21oi_1 _5796_ (.A1(_2313_),
    .A2(_2315_),
    .Y(_0263_),
    .B1(_2226_));
 sg13g2_mux2_1 _5797_ (.A0(_2306_),
    .A1(_2293_),
    .S(_0405_),
    .X(_2316_));
 sg13g2_a22oi_1 _5798_ (.Y(_2317_),
    .B1(net96),
    .B2(_2044_),
    .A2(net55),
    .A1(_0404_));
 sg13g2_o21ai_1 _5799_ (.B1(_2317_),
    .Y(_0264_),
    .A1(_1632_),
    .A2(_2316_));
 sg13g2_nand2_1 _5800_ (.Y(_2318_),
    .A(_0404_),
    .B(net23));
 sg13g2_o21ai_1 _5801_ (.B1(_0403_),
    .Y(_2319_),
    .A1(net70),
    .A2(net71));
 sg13g2_a21oi_1 _5802_ (.A1(_2318_),
    .A2(_2319_),
    .Y(_0265_),
    .B1(net72));
 sg13g2_mux2_1 _5803_ (.A0(_2093_),
    .A1(_2091_),
    .S(_1935_),
    .X(_2320_));
 sg13g2_and2_1 _5804_ (.A(net100),
    .B(_2320_),
    .X(_0266_));
 sg13g2_nand2_1 _5805_ (.Y(_2321_),
    .A(_2093_),
    .B(_2065_));
 sg13g2_o21ai_1 _5806_ (.B1(_2105_),
    .Y(_2322_),
    .A1(net70),
    .A2(_2067_));
 sg13g2_a21oi_1 _5807_ (.A1(_2321_),
    .A2(_2322_),
    .Y(_0267_),
    .B1(net72));
 sg13g2_a22oi_1 _5808_ (.Y(_2323_),
    .B1(_2098_),
    .B2(_2108_),
    .A2(_2116_),
    .A1(_2114_));
 sg13g2_a221oi_1 _5809_ (.B2(_2112_),
    .C1(_2092_),
    .B1(_2110_),
    .A1(net133),
    .Y(_2324_),
    .A2(_2103_));
 sg13g2_a21oi_1 _5810_ (.A1(_2092_),
    .A2(_2323_),
    .Y(_2325_),
    .B1(_2324_));
 sg13g2_mux2_1 _5811_ (.A0(_0404_),
    .A1(_2325_),
    .S(net124),
    .X(_2326_));
 sg13g2_nor2b_1 _5812_ (.A(net123),
    .B_N(_2093_),
    .Y(_2327_));
 sg13g2_a21oi_1 _5813_ (.A1(_2740_),
    .A2(_2326_),
    .Y(_2328_),
    .B1(_2327_));
 sg13g2_nor2_1 _5814_ (.A(net76),
    .B(_2328_),
    .Y(_0268_));
 sg13g2_nand2_1 _5815_ (.Y(_2329_),
    .A(_2093_),
    .B(net23));
 sg13g2_o21ai_1 _5816_ (.B1(_2090_),
    .Y(_2330_),
    .A1(net70),
    .A2(net71));
 sg13g2_a21oi_1 _5817_ (.A1(_2329_),
    .A2(_2330_),
    .Y(_0269_),
    .B1(_2226_));
 sg13g2_mux2_1 _5818_ (.A0(_0536_),
    .A1(_0537_),
    .S(net42),
    .X(_2331_));
 sg13g2_and2_1 _5819_ (.A(net100),
    .B(_2331_),
    .X(_0270_));
 sg13g2_mux2_1 _5820_ (.A0(_2165_),
    .A1(_2168_),
    .S(_2166_),
    .X(_2332_));
 sg13g2_nor3_1 _5821_ (.A(_2175_),
    .B(_2171_),
    .C(_2172_),
    .Y(_2333_));
 sg13g2_a21oi_1 _5822_ (.A1(_2175_),
    .A2(_2332_),
    .Y(_2334_),
    .B1(_2333_));
 sg13g2_nand3b_1 _5823_ (.B(_2156_),
    .C(net134),
    .Y(_2335_),
    .A_N(_2334_));
 sg13g2_nand2_1 _5824_ (.Y(_2336_),
    .A(_2175_),
    .B(_2170_));
 sg13g2_or2_1 _5825_ (.X(_2337_),
    .B(\g.g_y[6].g_x[7].t.out_sc ),
    .A(_2175_));
 sg13g2_buf_1 _5826_ (.A(_2337_),
    .X(_2338_));
 sg13g2_nand2_1 _5827_ (.Y(_2339_),
    .A(net134),
    .B(_2157_));
 sg13g2_a21o_1 _5828_ (.A2(_2338_),
    .A1(_2336_),
    .B1(_2339_),
    .X(_2340_));
 sg13g2_inv_1 _5829_ (.Y(_2341_),
    .A(net133));
 sg13g2_nor3_1 _5830_ (.A(net134),
    .B(_2341_),
    .C(_2288_),
    .Y(_2342_));
 sg13g2_nor3_1 _5831_ (.A(net134),
    .B(net133),
    .C(_2287_),
    .Y(_2343_));
 sg13g2_nor4_1 _5832_ (.A(net134),
    .B(_2341_),
    .C(_2091_),
    .D(_2093_),
    .Y(_2344_));
 sg13g2_nor3_1 _5833_ (.A(_2342_),
    .B(_2343_),
    .C(_2344_),
    .Y(_2345_));
 sg13g2_nor3_1 _5834_ (.A(_0537_),
    .B(_2709_),
    .C(_0457_),
    .Y(_2346_));
 sg13g2_nand4_1 _5835_ (.B(_2340_),
    .C(_2345_),
    .A(_2335_),
    .Y(_2347_),
    .D(_2346_));
 sg13g2_mux2_1 _5836_ (.A0(_0552_),
    .A1(_0563_),
    .S(net162),
    .X(_2348_));
 sg13g2_nor2_1 _5837_ (.A(net162),
    .B(_0554_),
    .Y(_2349_));
 sg13g2_nor2_1 _5838_ (.A(_0535_),
    .B(_2349_),
    .Y(_2350_));
 sg13g2_nor2b_1 _5839_ (.A(_1892_),
    .B_N(_1888_),
    .Y(_2351_));
 sg13g2_o21ai_1 _5840_ (.B1(_1888_),
    .Y(_2352_),
    .A1(_1893_),
    .A2(_1874_));
 sg13g2_a21o_1 _5841_ (.A2(_1887_),
    .A1(_1892_),
    .B1(_1888_),
    .X(_2353_));
 sg13g2_a21o_1 _5842_ (.A2(_1891_),
    .A1(_1893_),
    .B1(_2353_),
    .X(_2354_));
 sg13g2_a221oi_1 _5843_ (.B2(_2354_),
    .C1(_0534_),
    .B1(_2352_),
    .A1(_1890_),
    .Y(_2355_),
    .A2(_2351_));
 sg13g2_a21o_1 _5844_ (.A2(_2350_),
    .A1(_2348_),
    .B1(_2355_),
    .X(_2356_));
 sg13g2_nand4_1 _5845_ (.B(_2582_),
    .C(_2598_),
    .A(_0537_),
    .Y(_2357_),
    .D(_2356_));
 sg13g2_nand3_1 _5846_ (.B(net160),
    .C(_0457_),
    .A(_0539_),
    .Y(_2358_));
 sg13g2_nand3_1 _5847_ (.B(_2357_),
    .C(_2358_),
    .A(_2347_),
    .Y(_0271_));
 sg13g2_and2_1 _5848_ (.A(_0560_),
    .B(_0554_),
    .X(_2359_));
 sg13g2_a22oi_1 _5849_ (.Y(_2360_),
    .B1(_2359_),
    .B2(_0552_),
    .A2(_0563_),
    .A1(net162));
 sg13g2_a21o_1 _5850_ (.A2(_1890_),
    .A1(_1893_),
    .B1(_2352_),
    .X(_2361_));
 sg13g2_and3_1 _5851_ (.X(_2362_),
    .A(_0534_),
    .B(_2354_),
    .C(_2361_));
 sg13g2_a21oi_1 _5852_ (.A1(_0535_),
    .A2(_2360_),
    .Y(_2363_),
    .B1(_2362_));
 sg13g2_nor2_1 _5853_ (.A(_2341_),
    .B(_2289_),
    .Y(_2364_));
 sg13g2_a221oi_1 _5854_ (.B2(_2364_),
    .C1(_2102_),
    .B1(_2288_),
    .A1(_2341_),
    .Y(_2365_),
    .A2(_2287_));
 sg13g2_and2_1 _5855_ (.A(_2157_),
    .B(_2338_),
    .X(_2366_));
 sg13g2_a221oi_1 _5856_ (.B2(_2366_),
    .C1(net134),
    .B1(_2336_),
    .A1(_2156_),
    .Y(_2367_),
    .A2(_2334_));
 sg13g2_nor3_1 _5857_ (.A(_0457_),
    .B(_2365_),
    .C(_2367_),
    .Y(_2368_));
 sg13g2_o21ai_1 _5858_ (.B1(net132),
    .Y(_2369_),
    .A1(\g.g_y[6].g_x[6].t.r_gnl ),
    .A2(_2598_));
 sg13g2_a21oi_1 _5859_ (.A1(_2363_),
    .A2(_2368_),
    .Y(_0272_),
    .B1(_2369_));
 sg13g2_nand2_1 _5860_ (.Y(_2370_),
    .A(_0536_),
    .B(_2065_));
 sg13g2_o21ai_1 _5861_ (.B1(_2101_),
    .Y(_2371_),
    .A1(net70),
    .A2(_2067_));
 sg13g2_buf_1 _5862_ (.A(net128),
    .X(_2372_));
 sg13g2_a21oi_1 _5863_ (.A1(_2370_),
    .A2(_2371_),
    .Y(_0273_),
    .B1(net69));
 sg13g2_and2_1 _5864_ (.A(_0537_),
    .B(net88),
    .X(_2373_));
 sg13g2_nand4_1 _5865_ (.B(_2340_),
    .C(_2345_),
    .A(_2335_),
    .Y(_2374_),
    .D(_2373_));
 sg13g2_nand3b_1 _5866_ (.B(_0812_),
    .C(_2356_),
    .Y(_2375_),
    .A_N(_0537_));
 sg13g2_a22oi_1 _5867_ (.Y(_2376_),
    .B1(net96),
    .B2(_2093_),
    .A2(_0815_),
    .A1(_0536_));
 sg13g2_nand3_1 _5868_ (.B(_2375_),
    .C(_2376_),
    .A(_2374_),
    .Y(_0274_));
 sg13g2_nand2_1 _5869_ (.Y(_2377_),
    .A(_0536_),
    .B(net23));
 sg13g2_o21ai_1 _5870_ (.B1(_0534_),
    .Y(_2378_),
    .A1(net70),
    .A2(net71));
 sg13g2_a21oi_1 _5871_ (.A1(_2377_),
    .A2(_2378_),
    .Y(_0275_),
    .B1(net69));
 sg13g2_nor2_1 _5872_ (.A(_2174_),
    .B(_1394_),
    .Y(_2379_));
 sg13g2_a21oi_1 _5873_ (.A1(_2175_),
    .A2(net41),
    .Y(_2380_),
    .B1(_2379_));
 sg13g2_nor2_1 _5874_ (.A(_1933_),
    .B(_2380_),
    .Y(_0276_));
 sg13g2_mux2_1 _5875_ (.A0(_2157_),
    .A1(_2174_),
    .S(_2701_),
    .X(_2381_));
 sg13g2_nor2_1 _5876_ (.A(net97),
    .B(_2381_),
    .Y(_0277_));
 sg13g2_mux2_1 _5877_ (.A0(_2332_),
    .A1(_2173_),
    .S(_2175_),
    .X(_2382_));
 sg13g2_nand2_1 _5878_ (.Y(_2383_),
    .A(_1127_),
    .B(_0536_));
 sg13g2_o21ai_1 _5879_ (.B1(_2383_),
    .Y(_2384_),
    .A1(_0614_),
    .A2(_2382_));
 sg13g2_nor2_1 _5880_ (.A(_2174_),
    .B(_2745_),
    .Y(_2385_));
 sg13g2_a21oi_1 _5881_ (.A1(_2740_),
    .A2(_2384_),
    .Y(_2386_),
    .B1(_2385_));
 sg13g2_nor2_1 _5882_ (.A(net97),
    .B(_2386_),
    .Y(_0278_));
 sg13g2_nand2_1 _5883_ (.Y(_2387_),
    .A(\g.g_y[6].g_x[7].t.out_sc ),
    .B(_2231_));
 sg13g2_o21ai_1 _5884_ (.B1(_2166_),
    .Y(_2388_),
    .A1(net70),
    .A2(_2233_));
 sg13g2_a21oi_1 _5885_ (.A1(_2387_),
    .A2(_2388_),
    .Y(_0279_),
    .B1(net69));
 sg13g2_mux2_1 _5886_ (.A0(_2659_),
    .A1(net130),
    .S(net42),
    .X(_2389_));
 sg13g2_and2_1 _5887_ (.A(net100),
    .B(_2389_),
    .X(_0280_));
 sg13g2_nand2_1 _5888_ (.Y(_2390_),
    .A(_2659_),
    .B(net37));
 sg13g2_o21ai_1 _5889_ (.B1(_2644_),
    .Y(_2391_),
    .A1(_2314_),
    .A2(net129));
 sg13g2_a21oi_1 _5890_ (.A1(_2390_),
    .A2(_2391_),
    .Y(_0281_),
    .B1(net69));
 sg13g2_nand2_1 _5891_ (.Y(_2392_),
    .A(_2655_),
    .B(_2194_));
 sg13g2_a21o_1 _5892_ (.A2(_2651_),
    .A1(_2647_),
    .B1(_2653_),
    .X(_2393_));
 sg13g2_nand2b_1 _5893_ (.Y(_2394_),
    .B(_2393_),
    .A_N(_2655_));
 sg13g2_nand2_1 _5894_ (.Y(_2395_),
    .A(_2392_),
    .B(_2394_));
 sg13g2_mux2_1 _5895_ (.A0(_2395_),
    .A1(_2645_),
    .S(net130),
    .X(_2396_));
 sg13g2_nand2_1 _5896_ (.Y(_2397_),
    .A(net170),
    .B(_2174_));
 sg13g2_o21ai_1 _5897_ (.B1(_2397_),
    .Y(_2398_),
    .A1(_0631_),
    .A2(_2396_));
 sg13g2_nor2_1 _5898_ (.A(_2659_),
    .B(_2739_),
    .Y(_2399_));
 sg13g2_a21oi_1 _5899_ (.A1(net109),
    .A2(_2398_),
    .Y(_2400_),
    .B1(_2399_));
 sg13g2_and2_1 _5900_ (.A(net100),
    .B(_2400_),
    .X(_0282_));
 sg13g2_nand2_1 _5901_ (.Y(_2401_),
    .A(_2659_),
    .B(_2231_));
 sg13g2_o21ai_1 _5902_ (.B1(_2655_),
    .Y(_2402_),
    .A1(_2314_),
    .A2(_2233_));
 sg13g2_a21oi_1 _5903_ (.A1(_2401_),
    .A2(_2402_),
    .Y(_0283_),
    .B1(_2372_));
 sg13g2_mux2_1 _5904_ (.A0(_2603_),
    .A1(_2604_),
    .S(net42),
    .X(_2403_));
 sg13g2_and2_1 _5905_ (.A(_2243_),
    .B(_2403_),
    .X(_0284_));
 sg13g2_mux2_1 _5906_ (.A0(_2194_),
    .A1(_2393_),
    .S(_2655_),
    .X(_2404_));
 sg13g2_and2_1 _5907_ (.A(net8),
    .B(_2638_),
    .X(_2405_));
 sg13g2_nor2_1 _5908_ (.A(_2659_),
    .B(_2638_),
    .Y(_2406_));
 sg13g2_a21oi_1 _5909_ (.A1(_2404_),
    .A2(_2405_),
    .Y(_2407_),
    .B1(_2406_));
 sg13g2_nand3_1 _5910_ (.B(_2392_),
    .C(_2394_),
    .A(net130),
    .Y(_2408_));
 sg13g2_nor2_1 _5911_ (.A(net8),
    .B(_2639_),
    .Y(_2409_));
 sg13g2_nor2_1 _5912_ (.A(_2644_),
    .B(_2409_),
    .Y(_2410_));
 sg13g2_a22oi_1 _5913_ (.Y(_2411_),
    .B1(_2408_),
    .B2(_2410_),
    .A2(_2407_),
    .A1(_2644_));
 sg13g2_mux2_1 _5914_ (.A0(_2809_),
    .A1(_2623_),
    .S(net173),
    .X(_2412_));
 sg13g2_a21o_1 _5915_ (.A2(_2803_),
    .A1(_2800_),
    .B1(_2805_),
    .X(_2413_));
 sg13g2_mux2_1 _5916_ (.A0(_2412_),
    .A1(_2413_),
    .S(_2812_),
    .X(_2414_));
 sg13g2_nand3_1 _5917_ (.B(_2414_),
    .C(_2826_),
    .A(net172),
    .Y(_2415_));
 sg13g2_nor2_1 _5918_ (.A(net172),
    .B(_2831_),
    .Y(_2416_));
 sg13g2_nor2_1 _5919_ (.A(_2820_),
    .B(_2416_),
    .Y(_2417_));
 sg13g2_o21ai_1 _5920_ (.B1(_2820_),
    .Y(_2418_),
    .A1(net172),
    .A2(_2826_));
 sg13g2_inv_1 _5921_ (.Y(_2419_),
    .A(_2418_));
 sg13g2_nand2_1 _5922_ (.Y(_2420_),
    .A(net172),
    .B(_2813_));
 sg13g2_a22oi_1 _5923_ (.Y(_2421_),
    .B1(_2419_),
    .B2(_2420_),
    .A2(_2417_),
    .A1(_2415_));
 sg13g2_mux2_1 _5924_ (.A0(_2411_),
    .A1(_2421_),
    .S(_2641_),
    .X(_2422_));
 sg13g2_a21oi_1 _5925_ (.A1(_1956_),
    .A2(_1976_),
    .Y(_2423_),
    .B1(_1962_));
 sg13g2_a21oi_1 _5926_ (.A1(net136),
    .A2(_2209_),
    .Y(_2424_),
    .B1(_1985_));
 sg13g2_a22oi_1 _5927_ (.Y(_2425_),
    .B1(_2424_),
    .B2(_1962_),
    .A2(_2423_),
    .A1(_1974_));
 sg13g2_and2_1 _5928_ (.A(_2615_),
    .B(_0667_),
    .X(_2426_));
 sg13g2_mux2_1 _5929_ (.A0(_2741_),
    .A1(_2613_),
    .S(_2601_),
    .X(_2427_));
 sg13g2_a22oi_1 _5930_ (.Y(_2428_),
    .B1(_2427_),
    .B2(_2614_),
    .A2(_2426_),
    .A1(_0666_));
 sg13g2_mux2_1 _5931_ (.A0(_2425_),
    .A1(_2428_),
    .S(_2606_),
    .X(_2429_));
 sg13g2_mux2_1 _5932_ (.A0(_2422_),
    .A1(_2429_),
    .S(_2604_),
    .X(_2430_));
 sg13g2_o21ai_1 _5933_ (.B1(_2179_),
    .Y(_2431_),
    .A1(_2602_),
    .A2(net32));
 sg13g2_a21oi_1 _5934_ (.A1(_0805_),
    .A2(_2430_),
    .Y(_0285_),
    .B1(_2431_));
 sg13g2_nand2b_1 _5935_ (.Y(_2432_),
    .B(_2606_),
    .A_N(_2425_));
 sg13g2_or2_1 _5936_ (.X(_2433_),
    .B(_2428_),
    .A(_2606_));
 sg13g2_nor2b_1 _5937_ (.A(_2641_),
    .B_N(_2421_),
    .Y(_2434_));
 sg13g2_a221oi_1 _5938_ (.B2(_2433_),
    .C1(_2434_),
    .B1(_2432_),
    .A1(_2641_),
    .Y(_2435_),
    .A2(_2411_));
 sg13g2_o21ai_1 _5939_ (.B1(_2179_),
    .Y(_2436_),
    .A1(\g.g_y[7].g_x[1].t.r_gnl ),
    .A2(net32));
 sg13g2_a21oi_1 _5940_ (.A1(_0805_),
    .A2(_2435_),
    .Y(_0286_),
    .B1(_2436_));
 sg13g2_nand2_1 _5941_ (.Y(_2437_),
    .A(_2603_),
    .B(net37));
 sg13g2_o21ai_1 _5942_ (.B1(_2641_),
    .Y(_2438_),
    .A1(net70),
    .A2(net129));
 sg13g2_a21oi_1 _5943_ (.A1(_2437_),
    .A2(_2438_),
    .Y(_0287_),
    .B1(net69));
 sg13g2_mux2_1 _5944_ (.A0(_2429_),
    .A1(_2422_),
    .S(_2604_),
    .X(_2439_));
 sg13g2_a22oi_1 _5945_ (.Y(_2440_),
    .B1(_2722_),
    .B2(_2659_),
    .A2(net55),
    .A1(_2603_));
 sg13g2_o21ai_1 _5946_ (.B1(_2440_),
    .Y(_0288_),
    .A1(_2715_),
    .A2(_2439_));
 sg13g2_nand2_1 _5947_ (.Y(_2441_),
    .A(_2603_),
    .B(net23));
 sg13g2_buf_1 _5948_ (.A(_2589_),
    .X(_2442_));
 sg13g2_o21ai_1 _5949_ (.B1(_2606_),
    .Y(_2443_),
    .A1(net68),
    .A2(net71));
 sg13g2_a21oi_1 _5950_ (.A1(_2441_),
    .A2(_2443_),
    .Y(_0289_),
    .B1(net69));
 sg13g2_mux2_1 _5951_ (.A0(_2831_),
    .A1(_2822_),
    .S(_0607_),
    .X(_2444_));
 sg13g2_and2_1 _5952_ (.A(_2243_),
    .B(_2444_),
    .X(_0290_));
 sg13g2_nand2_1 _5953_ (.Y(_2445_),
    .A(_2831_),
    .B(net37));
 sg13g2_o21ai_1 _5954_ (.B1(_2820_),
    .Y(_2446_),
    .A1(net68),
    .A2(net129));
 sg13g2_a21oi_1 _5955_ (.A1(_2445_),
    .A2(_2446_),
    .Y(_0291_),
    .B1(net69));
 sg13g2_nor2_1 _5956_ (.A(_2831_),
    .B(net110),
    .Y(_2447_));
 sg13g2_mux2_1 _5957_ (.A0(_2813_),
    .A1(_2821_),
    .S(net172),
    .X(_2448_));
 sg13g2_nand2_1 _5958_ (.Y(_2449_),
    .A(_0324_),
    .B(_2603_));
 sg13g2_o21ai_1 _5959_ (.B1(_2449_),
    .Y(_2450_),
    .A1(net120),
    .A2(_2448_));
 sg13g2_nor2b_1 _5960_ (.A(_2450_),
    .B_N(net109),
    .Y(_2451_));
 sg13g2_nor3_1 _5961_ (.A(net126),
    .B(_2447_),
    .C(_2451_),
    .Y(_0292_));
 sg13g2_nand2_1 _5962_ (.Y(_2452_),
    .A(_2831_),
    .B(net23));
 sg13g2_o21ai_1 _5963_ (.B1(_2812_),
    .Y(_2453_),
    .A1(_2442_),
    .A2(net71));
 sg13g2_a21oi_1 _5964_ (.A1(_2452_),
    .A2(_2453_),
    .Y(_0293_),
    .B1(_2372_));
 sg13g2_mux2_1 _5965_ (.A0(_2760_),
    .A1(_2761_),
    .S(net42),
    .X(_2454_));
 sg13g2_and2_1 _5966_ (.A(net100),
    .B(_2454_),
    .X(_0294_));
 sg13g2_nor2_1 _5967_ (.A(_2823_),
    .B(_2815_),
    .Y(_2455_));
 sg13g2_a21oi_1 _5968_ (.A1(_2414_),
    .A2(_2455_),
    .Y(_2456_),
    .B1(_2416_));
 sg13g2_a21oi_1 _5969_ (.A1(_2823_),
    .A2(_2815_),
    .Y(_2457_),
    .B1(_2820_));
 sg13g2_a22oi_1 _5970_ (.Y(_2458_),
    .B1(_2457_),
    .B2(_2420_),
    .A2(_2456_),
    .A1(_2820_));
 sg13g2_a21o_1 _5971_ (.A2(_0406_),
    .A1(_0403_),
    .B1(_0408_),
    .X(_2459_));
 sg13g2_mux2_1 _5972_ (.A0(_2459_),
    .A1(_2301_),
    .S(_0412_),
    .X(_2460_));
 sg13g2_nand3_1 _5973_ (.B(_0391_),
    .C(_2460_),
    .A(net119),
    .Y(_2461_));
 sg13g2_nor2_1 _5974_ (.A(_0386_),
    .B(_0398_),
    .Y(_2462_));
 sg13g2_nor2_1 _5975_ (.A(_0393_),
    .B(_2462_),
    .Y(_2463_));
 sg13g2_mux2_1 _5976_ (.A0(_2459_),
    .A1(_2301_),
    .S(net166),
    .X(_2464_));
 sg13g2_mux2_1 _5977_ (.A0(_0391_),
    .A1(_2464_),
    .S(_0386_),
    .X(_2465_));
 sg13g2_a22oi_1 _5978_ (.Y(_2466_),
    .B1(_2465_),
    .B2(_0393_),
    .A2(_2463_),
    .A1(_2461_));
 sg13g2_mux2_1 _5979_ (.A0(_2458_),
    .A1(_2466_),
    .S(_2816_),
    .X(_2467_));
 sg13g2_mux4_1 _5980_ (.S0(_2029_),
    .A0(_2043_),
    .A1(_2042_),
    .A2(_2250_),
    .A3(_2045_),
    .S1(_2047_),
    .X(_2468_));
 sg13g2_nor2_1 _5981_ (.A(_2773_),
    .B(_0780_),
    .Y(_2469_));
 sg13g2_a21oi_1 _5982_ (.A1(_2758_),
    .A2(_2793_),
    .Y(_2470_),
    .B1(_2774_));
 sg13g2_a22oi_1 _5983_ (.Y(_2471_),
    .B1(_2470_),
    .B2(_0782_),
    .A2(_2469_),
    .A1(_0779_));
 sg13g2_mux2_1 _5984_ (.A0(_2468_),
    .A1(_2471_),
    .S(_2759_),
    .X(_2472_));
 sg13g2_mux2_1 _5985_ (.A0(_2467_),
    .A1(_2472_),
    .S(_2761_),
    .X(_2473_));
 sg13g2_o21ai_1 _5986_ (.B1(net132),
    .Y(_2474_),
    .A1(_2763_),
    .A2(net57));
 sg13g2_a21oi_1 _5987_ (.A1(net39),
    .A2(_2473_),
    .Y(_0295_),
    .B1(_2474_));
 sg13g2_mux2_1 _5988_ (.A0(_2471_),
    .A1(_2468_),
    .S(_2759_),
    .X(_2475_));
 sg13g2_mux2_1 _5989_ (.A0(_2466_),
    .A1(_2458_),
    .S(_2816_),
    .X(_2476_));
 sg13g2_nor3_1 _5990_ (.A(_0704_),
    .B(_2475_),
    .C(_2476_),
    .Y(_2477_));
 sg13g2_o21ai_1 _5991_ (.B1(net177),
    .Y(_2478_),
    .A1(\g.g_y[7].g_x[3].t.r_gnl ),
    .A2(_0702_));
 sg13g2_nor2_1 _5992_ (.A(_2477_),
    .B(_2478_),
    .Y(_0296_));
 sg13g2_nand2_1 _5993_ (.Y(_2479_),
    .A(_2760_),
    .B(net37));
 sg13g2_o21ai_1 _5994_ (.B1(_2816_),
    .Y(_2480_),
    .A1(net68),
    .A2(net129));
 sg13g2_a21oi_1 _5995_ (.A1(_2479_),
    .A2(_2480_),
    .Y(_0297_),
    .B1(net69));
 sg13g2_mux2_1 _5996_ (.A0(_2472_),
    .A1(_2467_),
    .S(_2761_),
    .X(_2481_));
 sg13g2_a22oi_1 _5997_ (.Y(_2482_),
    .B1(net96),
    .B2(_2831_),
    .A2(net55),
    .A1(_2760_));
 sg13g2_o21ai_1 _5998_ (.B1(_2482_),
    .Y(_0298_),
    .A1(_2715_),
    .A2(_2481_));
 sg13g2_nand2_1 _5999_ (.Y(_2483_),
    .A(_2760_),
    .B(net40));
 sg13g2_o21ai_1 _6000_ (.B1(_2759_),
    .Y(_2484_),
    .A1(net68),
    .A2(net127));
 sg13g2_buf_1 _6001_ (.A(net128),
    .X(_2485_));
 sg13g2_a21oi_1 _6002_ (.A1(_2483_),
    .A2(_2484_),
    .Y(_0299_),
    .B1(net67));
 sg13g2_mux2_1 _6003_ (.A0(_0398_),
    .A1(net119),
    .S(net42),
    .X(_2486_));
 sg13g2_and2_1 _6004_ (.A(net100),
    .B(_2486_),
    .X(_0300_));
 sg13g2_nand2_1 _6005_ (.Y(_2487_),
    .A(_0398_),
    .B(net37));
 sg13g2_o21ai_1 _6006_ (.B1(_0393_),
    .Y(_2488_),
    .A1(net68),
    .A2(net129));
 sg13g2_a21oi_1 _6007_ (.A1(_2487_),
    .A2(_2488_),
    .Y(_0301_),
    .B1(net67));
 sg13g2_mux2_1 _6008_ (.A0(_2464_),
    .A1(_0396_),
    .S(net119),
    .X(_2489_));
 sg13g2_nand2b_1 _6009_ (.Y(_2490_),
    .B(_2895_),
    .A_N(_2760_));
 sg13g2_o21ai_1 _6010_ (.B1(_2490_),
    .Y(_2491_),
    .A1(_1127_),
    .A2(_2489_));
 sg13g2_nand2_1 _6011_ (.Y(_2492_),
    .A(_1049_),
    .B(_2491_));
 sg13g2_o21ai_1 _6012_ (.B1(_2492_),
    .Y(_2493_),
    .A1(_0398_),
    .A2(net121));
 sg13g2_nor2_1 _6013_ (.A(net97),
    .B(_2493_),
    .Y(_0302_));
 sg13g2_nand2_1 _6014_ (.Y(_2494_),
    .A(_0398_),
    .B(net40));
 sg13g2_o21ai_1 _6015_ (.B1(_0385_),
    .Y(_2495_),
    .A1(net68),
    .A2(_2731_));
 sg13g2_a21oi_1 _6016_ (.A1(_2494_),
    .A2(_2495_),
    .Y(_0303_),
    .B1(net67));
 sg13g2_mux2_1 _6017_ (.A0(_0345_),
    .A1(_0346_),
    .S(net42),
    .X(_2496_));
 sg13g2_and2_1 _6018_ (.A(net117),
    .B(_2496_),
    .X(_0304_));
 sg13g2_nand3_1 _6019_ (.B(_0402_),
    .C(_2460_),
    .A(_0387_),
    .Y(_2497_));
 sg13g2_nor2_1 _6020_ (.A(_0394_),
    .B(_2462_),
    .Y(_2498_));
 sg13g2_mux2_1 _6021_ (.A0(_0396_),
    .A1(_2464_),
    .S(_0386_),
    .X(_2499_));
 sg13g2_a22oi_1 _6022_ (.Y(_2500_),
    .B1(_2499_),
    .B2(_0394_),
    .A2(_2498_),
    .A1(_2497_));
 sg13g2_or3_1 _6023_ (.A(_0556_),
    .B(_0543_),
    .C(_0547_),
    .X(_2501_));
 sg13g2_nor2_1 _6024_ (.A(_0528_),
    .B(_0553_),
    .Y(_2502_));
 sg13g2_nor2_1 _6025_ (.A(_0550_),
    .B(_2502_),
    .Y(_2503_));
 sg13g2_a21oi_1 _6026_ (.A1(_0556_),
    .A2(_0547_),
    .Y(_2504_),
    .B1(_0562_));
 sg13g2_a22oi_1 _6027_ (.Y(_2505_),
    .B1(_2504_),
    .B2(_0550_),
    .A2(_2503_),
    .A1(_2501_));
 sg13g2_mux2_1 _6028_ (.A0(_2500_),
    .A1(_2505_),
    .S(_0389_),
    .X(_2506_));
 sg13g2_inv_1 _6029_ (.Y(_2507_),
    .A(_0346_));
 sg13g2_nand2b_1 _6030_ (.Y(_2508_),
    .B(_2507_),
    .A_N(_2506_));
 sg13g2_mux2_1 _6031_ (.A0(_0876_),
    .A1(_0871_),
    .S(_0352_),
    .X(_2509_));
 sg13g2_nand2_1 _6032_ (.Y(_2510_),
    .A(_0343_),
    .B(_2509_));
 sg13g2_a21oi_1 _6033_ (.A1(_1497_),
    .A2(_1500_),
    .Y(_2511_),
    .B1(_2097_));
 sg13g2_a21oi_1 _6034_ (.A1(_2091_),
    .A2(_2511_),
    .Y(_2512_),
    .B1(_2113_));
 sg13g2_nor2_1 _6035_ (.A(_2108_),
    .B(_2094_),
    .Y(_2513_));
 sg13g2_a22oi_1 _6036_ (.Y(_2514_),
    .B1(_2513_),
    .B2(_2107_),
    .A2(_2512_),
    .A1(_2108_));
 sg13g2_a21oi_1 _6037_ (.A1(_0344_),
    .A2(_2514_),
    .Y(_2515_),
    .B1(_2507_));
 sg13g2_a21oi_1 _6038_ (.A1(_2510_),
    .A2(_2515_),
    .Y(_2516_),
    .B1(net56));
 sg13g2_a221oi_1 _6039_ (.B2(_2516_),
    .C1(net67),
    .B1(_2508_),
    .A1(_2115_),
    .Y(_0305_),
    .A2(_0729_));
 sg13g2_mux2_1 _6040_ (.A0(_2505_),
    .A1(_2500_),
    .S(_0389_),
    .X(_2517_));
 sg13g2_mux2_1 _6041_ (.A0(_2509_),
    .A1(_2514_),
    .S(_0343_),
    .X(_2518_));
 sg13g2_nor3_1 _6042_ (.A(_0729_),
    .B(_2517_),
    .C(_2518_),
    .Y(_2519_));
 sg13g2_o21ai_1 _6043_ (.B1(_2690_),
    .Y(_2520_),
    .A1(\g.g_y[7].g_x[5].t.r_gnl ),
    .A2(net36));
 sg13g2_nor2_1 _6044_ (.A(_2519_),
    .B(_2520_),
    .Y(_0306_));
 sg13g2_nand2_1 _6045_ (.Y(_2521_),
    .A(_0345_),
    .B(net37));
 sg13g2_o21ai_1 _6046_ (.B1(_0389_),
    .Y(_2522_),
    .A1(net68),
    .A2(net129));
 sg13g2_a21oi_1 _6047_ (.A1(_2521_),
    .A2(_2522_),
    .Y(_0307_),
    .B1(net67));
 sg13g2_a21oi_1 _6048_ (.A1(_0345_),
    .A2(_2719_),
    .Y(_2523_),
    .B1(net170));
 sg13g2_and3_1 _6049_ (.X(_2524_),
    .A(_0346_),
    .B(_2506_),
    .C(_2523_));
 sg13g2_nand2_1 _6050_ (.Y(_2525_),
    .A(_0344_),
    .B(_2514_));
 sg13g2_nand2_1 _6051_ (.Y(_2526_),
    .A(_2507_),
    .B(_2523_));
 sg13g2_a21oi_1 _6052_ (.A1(_2510_),
    .A2(_2525_),
    .Y(_2527_),
    .B1(_2526_));
 sg13g2_nand3b_1 _6053_ (.B(_2739_),
    .C(net116),
    .Y(_2528_),
    .A_N(_0398_));
 sg13g2_o21ai_1 _6054_ (.B1(_2528_),
    .Y(_2529_),
    .A1(_0345_),
    .A2(_1049_));
 sg13g2_nor4_1 _6055_ (.A(net126),
    .B(_2524_),
    .C(_2527_),
    .D(_2529_),
    .Y(_0308_));
 sg13g2_nand2_1 _6056_ (.Y(_2530_),
    .A(_0345_),
    .B(net40));
 sg13g2_o21ai_1 _6057_ (.B1(_0343_),
    .Y(_2531_),
    .A1(net68),
    .A2(net127));
 sg13g2_a21oi_1 _6058_ (.A1(_2530_),
    .A2(_2531_),
    .Y(_0309_),
    .B1(net67));
 sg13g2_mux2_1 _6059_ (.A0(_0553_),
    .A1(net164),
    .S(net42),
    .X(_2532_));
 sg13g2_and2_1 _6060_ (.A(_0466_),
    .B(_2532_),
    .X(_0310_));
 sg13g2_nand2_1 _6061_ (.Y(_2533_),
    .A(_0553_),
    .B(_0717_));
 sg13g2_o21ai_1 _6062_ (.B1(_0550_),
    .Y(_2534_),
    .A1(_2442_),
    .A2(_2706_));
 sg13g2_a21oi_1 _6063_ (.A1(_2533_),
    .A2(_2534_),
    .Y(_0311_),
    .B1(net67));
 sg13g2_a221oi_1 _6064_ (.B2(_0561_),
    .C1(net164),
    .B1(_0559_),
    .A1(net162),
    .Y(_2535_),
    .A2(_0558_));
 sg13g2_a21oi_1 _6065_ (.A1(net164),
    .A2(_0557_),
    .Y(_2536_),
    .B1(_2535_));
 sg13g2_mux2_1 _6066_ (.A0(_0345_),
    .A1(_2536_),
    .S(_2743_),
    .X(_2537_));
 sg13g2_nor2b_1 _6067_ (.A(_2745_),
    .B_N(_0553_),
    .Y(_2538_));
 sg13g2_a21oi_1 _6068_ (.A1(net125),
    .A2(_2537_),
    .Y(_2539_),
    .B1(_2538_));
 sg13g2_nor2_1 _6069_ (.A(net97),
    .B(_2539_),
    .Y(_0312_));
 sg13g2_nand2_1 _6070_ (.Y(_2540_),
    .A(_0553_),
    .B(_0624_));
 sg13g2_o21ai_1 _6071_ (.B1(_0542_),
    .Y(_2541_),
    .A1(net99),
    .A2(net127));
 sg13g2_a21oi_1 _6072_ (.A1(_2540_),
    .A2(_2541_),
    .Y(_0313_),
    .B1(_2485_));
 sg13g2_mux2_1 _6073_ (.A0(_0512_),
    .A1(_0513_),
    .S(net42),
    .X(_2542_));
 sg13g2_and2_1 _6074_ (.A(net117),
    .B(_2542_),
    .X(_0314_));
 sg13g2_a21o_1 _6075_ (.A2(_0388_),
    .A1(_0389_),
    .B1(_0548_),
    .X(_2543_));
 sg13g2_nand3b_1 _6076_ (.B(_2543_),
    .C(net164),
    .Y(_2544_),
    .A_N(_0543_));
 sg13g2_nor2b_1 _6077_ (.A(_2502_),
    .B_N(_0550_),
    .Y(_2545_));
 sg13g2_nor2_1 _6078_ (.A(net164),
    .B(_2543_),
    .Y(_2546_));
 sg13g2_nor3_1 _6079_ (.A(_0550_),
    .B(_0562_),
    .C(_2546_),
    .Y(_2547_));
 sg13g2_a21oi_1 _6080_ (.A1(_2544_),
    .A2(_2545_),
    .Y(_2548_),
    .B1(_2547_));
 sg13g2_nand3_1 _6081_ (.B(_2643_),
    .C(_2404_),
    .A(net130),
    .Y(_2549_));
 sg13g2_nor2_1 _6082_ (.A(_2644_),
    .B(_2406_),
    .Y(_2550_));
 sg13g2_o21ai_1 _6083_ (.B1(_2644_),
    .Y(_2551_),
    .A1(_2639_),
    .A2(_2643_));
 sg13g2_inv_1 _6084_ (.Y(_2552_),
    .A(_2551_));
 sg13g2_a22oi_1 _6085_ (.Y(_2553_),
    .B1(_2552_),
    .B2(_2408_),
    .A2(_2550_),
    .A1(_2549_));
 sg13g2_mux2_1 _6086_ (.A0(_2548_),
    .A1(_2553_),
    .S(_0544_),
    .X(_2554_));
 sg13g2_mux4_1 _6087_ (.S0(_2166_),
    .A0(_2173_),
    .A1(_2170_),
    .A2(_2165_),
    .A3(_2174_),
    .S1(_2175_),
    .X(_2555_));
 sg13g2_nand2b_1 _6088_ (.Y(_2556_),
    .B(net165),
    .A_N(_0508_));
 sg13g2_o21ai_1 _6089_ (.B1(_2556_),
    .Y(_2557_),
    .A1(net165),
    .A2(_0507_));
 sg13g2_mux4_1 _6090_ (.S0(_0518_),
    .A0(_0520_),
    .A1(_0617_),
    .A2(_0496_),
    .A3(_2557_),
    .S1(_0525_),
    .X(_2558_));
 sg13g2_mux2_1 _6091_ (.A0(_2555_),
    .A1(_2558_),
    .S(_0511_),
    .X(_2559_));
 sg13g2_mux2_1 _6092_ (.A0(_2554_),
    .A1(_2559_),
    .S(_0513_),
    .X(_2560_));
 sg13g2_o21ai_1 _6093_ (.B1(_0726_),
    .Y(_2561_),
    .A1(_0515_),
    .A2(net57));
 sg13g2_a21oi_1 _6094_ (.A1(_0702_),
    .A2(_2560_),
    .Y(_0315_),
    .B1(_2561_));
 sg13g2_mux2_1 _6095_ (.A0(_2558_),
    .A1(_2555_),
    .S(_0511_),
    .X(_2562_));
 sg13g2_mux2_1 _6096_ (.A0(_2553_),
    .A1(_2548_),
    .S(_0544_),
    .X(_2563_));
 sg13g2_nor3_1 _6097_ (.A(_0704_),
    .B(_2562_),
    .C(_2563_),
    .Y(_2564_));
 sg13g2_o21ai_1 _6098_ (.B1(_2690_),
    .Y(_2565_),
    .A1(\g.g_y[7].g_x[7].t.r_gnl ),
    .A2(net38));
 sg13g2_nor2_1 _6099_ (.A(_2564_),
    .B(_2565_),
    .Y(_0316_));
 sg13g2_nand2_1 _6100_ (.Y(_2566_),
    .A(_0512_),
    .B(_0717_));
 sg13g2_o21ai_1 _6101_ (.B1(_0544_),
    .Y(_2567_),
    .A1(_2704_),
    .A2(net129));
 sg13g2_a21oi_1 _6102_ (.A1(_2566_),
    .A2(_2567_),
    .Y(_0317_),
    .B1(_2485_));
 sg13g2_mux2_1 _6103_ (.A0(_2559_),
    .A1(_2554_),
    .S(_0513_),
    .X(_2568_));
 sg13g2_a22oi_1 _6104_ (.Y(_2569_),
    .B1(_2722_),
    .B2(_0553_),
    .A2(net55),
    .A1(_0512_));
 sg13g2_o21ai_1 _6105_ (.B1(_2569_),
    .Y(_0318_),
    .A1(_2715_),
    .A2(_2568_));
 sg13g2_nand2_1 _6106_ (.Y(_2570_),
    .A(_0512_),
    .B(_0624_));
 sg13g2_o21ai_1 _6107_ (.B1(_0511_),
    .Y(_2571_),
    .A1(_2704_),
    .A2(net127));
 sg13g2_a21oi_1 _6108_ (.A1(_2570_),
    .A2(_2571_),
    .Y(_0319_),
    .B1(net67));
 sg13g2_nand2_1 _6109_ (.Y(_2572_),
    .A(_0503_),
    .B(_0519_));
 sg13g2_mux4_1 _6110_ (.S0(_0525_),
    .A0(_0501_),
    .A1(_0615_),
    .A2(_0495_),
    .A3(_2572_),
    .S1(_0502_),
    .X(\g.g_y[0].g_x[7].t.out_r ));
 sg13g2_mux2_1 _6111_ (.A0(_0508_),
    .A1(_0565_),
    .S(_0566_),
    .X(\g.g_y[1].g_x[7].t.out_r ));
 sg13g2_nor2_1 _6112_ (.A(net154),
    .B(_0930_),
    .Y(_2573_));
 sg13g2_a21oi_1 _6113_ (.A1(net154),
    .A2(_1237_),
    .Y(_2574_),
    .B1(_2573_));
 sg13g2_nand2_1 _6114_ (.Y(_2575_),
    .A(_0922_),
    .B(_2574_));
 sg13g2_o21ai_1 _6115_ (.B1(_2575_),
    .Y(\g.g_y[2].g_x[7].t.out_r ),
    .A1(_0922_),
    .A2(_1278_));
 sg13g2_mux2_1 _6116_ (.A0(_0948_),
    .A1(_1247_),
    .S(_1248_),
    .X(\g.g_y[3].g_x[7].t.out_r ));
 sg13g2_nand2_1 _6117_ (.Y(_2576_),
    .A(net140),
    .B(_1868_));
 sg13g2_o21ai_1 _6118_ (.B1(_2576_),
    .Y(_2577_),
    .A1(net140),
    .A2(_1614_));
 sg13g2_nand2_1 _6119_ (.Y(_2578_),
    .A(_1596_),
    .B(_1869_));
 sg13g2_nand3_1 _6120_ (.B(_1603_),
    .C(_2578_),
    .A(_1618_),
    .Y(_2579_));
 sg13g2_o21ai_1 _6121_ (.B1(_2579_),
    .Y(\g.g_y[4].g_x[7].t.out_r ),
    .A1(_1618_),
    .A2(_2577_));
 sg13g2_mux2_1 _6122_ (.A0(_1608_),
    .A1(_1879_),
    .S(_1878_),
    .X(\g.g_y[5].g_x[7].t.out_r ));
 sg13g2_and3_1 _6123_ (.X(_2580_),
    .A(_2156_),
    .B(_2336_),
    .C(_2338_));
 sg13g2_a21o_1 _6124_ (.A2(_2334_),
    .A1(_2157_),
    .B1(_2580_),
    .X(\g.g_y[6].g_x[7].t.out_r ));
 sg13g2_mux2_1 _6125_ (.A0(_0515_),
    .A1(_0545_),
    .S(_0544_),
    .X(\g.g_y[7].g_x[7].t.out_r ));
 sg13g2_buf_2 clkbuf_leaf_0_clk (.A(clknet_3_1__leaf_clk),
    .X(clknet_leaf_0_clk));
 sg13g2_tiehi _6135__199 (.L_HI(net199));
 sg13g2_buf_1 _6128_ (.A(net185),
    .X(uio_oe[0]));
 sg13g2_buf_1 _6129_ (.A(net186),
    .X(uio_oe[1]));
 sg13g2_buf_1 _6130_ (.A(net187),
    .X(uio_oe[2]));
 sg13g2_buf_1 _6131_ (.A(net188),
    .X(uio_oe[3]));
 sg13g2_buf_1 _6132_ (.A(net189),
    .X(uio_oe[4]));
 sg13g2_buf_1 _6133_ (.A(net190),
    .X(uio_oe[5]));
 sg13g2_buf_1 _6134_ (.A(net191),
    .X(uio_oe[6]));
 sg13g2_buf_1 _6135_ (.A(net199),
    .X(uio_oe[7]));
 sg13g2_buf_1 _6136_ (.A(net192),
    .X(uio_out[0]));
 sg13g2_buf_1 _6137_ (.A(net193),
    .X(uio_out[1]));
 sg13g2_buf_1 _6138_ (.A(net194),
    .X(uio_out[2]));
 sg13g2_buf_1 _6139_ (.A(net195),
    .X(uio_out[3]));
 sg13g2_buf_1 _6140_ (.A(net196),
    .X(uio_out[4]));
 sg13g2_buf_1 _6141_ (.A(net197),
    .X(uio_out[5]));
 sg13g2_buf_1 _6142_ (.A(net198),
    .X(uio_out[6]));
 sg13g2_buf_1 _6143_ (.A(\g.g_y[7].g_x[7].t.out_sc ),
    .X(net13));
 sg13g2_buf_1 _6144_ (.A(\g.g_y[0].g_x[7].t.out_r ),
    .X(net14));
 sg13g2_buf_1 _6145_ (.A(\g.g_y[1].g_x[7].t.out_r ),
    .X(net15));
 sg13g2_buf_1 _6146_ (.A(\g.g_y[2].g_x[7].t.out_r ),
    .X(net16));
 sg13g2_buf_1 _6147_ (.A(\g.g_y[3].g_x[7].t.out_r ),
    .X(net17));
 sg13g2_buf_1 _6148_ (.A(\g.g_y[4].g_x[7].t.out_r ),
    .X(net18));
 sg13g2_buf_1 _6149_ (.A(\g.g_y[5].g_x[7].t.out_r ),
    .X(net19));
 sg13g2_buf_1 _6150_ (.A(\g.g_y[6].g_x[7].t.out_r ),
    .X(net20));
 sg13g2_buf_1 _6151_ (.A(\g.g_y[7].g_x[7].t.out_r ),
    .X(net21));
 sg13g2_dfrbp_1 \g.g_y[0].g_x[0].t.r_d$_SDFFE_PN0P_  (.CLK(clknet_leaf_18_clk),
    .RESET_B(net200),
    .D(_0000_),
    .Q_N(_3217_),
    .Q(\g.g_y[0].g_x[0].t.r_d ));
 sg13g2_dfrbp_1 \g.g_y[0].g_x[0].t.r_ghl$_SDFFE_PN0P_  (.CLK(clknet_leaf_18_clk),
    .RESET_B(net201),
    .D(_0001_),
    .Q_N(_3216_),
    .Q(\g.g_y[0].g_x[0].t.r_ghl ));
 sg13g2_dfrbp_1 \g.g_y[0].g_x[0].t.r_gnl$_SDFFE_PN0P_  (.CLK(clknet_leaf_19_clk),
    .RESET_B(net202),
    .D(_0002_),
    .Q_N(_3215_),
    .Q(\g.g_y[0].g_x[0].t.r_gnl ));
 sg13g2_dfrbp_1 \g.g_y[0].g_x[0].t.r_h$_SDFFE_PN0P_  (.CLK(clknet_leaf_18_clk),
    .RESET_B(net203),
    .D(_0003_),
    .Q_N(_3214_),
    .Q(\g.g_y[0].g_x[0].t.r_h ));
 sg13g2_dfrbp_1 \g.g_y[0].g_x[0].t.r_sc$_SDFFE_PN0P_  (.CLK(clknet_leaf_19_clk),
    .RESET_B(net204),
    .D(_0004_),
    .Q_N(_3213_),
    .Q(\g.g_y[0].g_x[0].t.out_sc ));
 sg13g2_dfrbp_1 \g.g_y[0].g_x[0].t.r_v$_SDFFE_PN0P_  (.CLK(clknet_leaf_18_clk),
    .RESET_B(net205),
    .D(_0005_),
    .Q_N(_3212_),
    .Q(\g.g_y[0].g_x[0].t.r_v ));
 sg13g2_dfrbp_1 \g.g_y[0].g_x[1].t.r_d$_SDFFE_PN0P_  (.CLK(clknet_leaf_18_clk),
    .RESET_B(net206),
    .D(_0006_),
    .Q_N(_3211_),
    .Q(\g.g_y[0].g_x[1].t.r_d ));
 sg13g2_dfrbp_1 \g.g_y[0].g_x[1].t.r_h$_SDFFE_PN0P_  (.CLK(clknet_leaf_18_clk),
    .RESET_B(net207),
    .D(_0007_),
    .Q_N(_3210_),
    .Q(\g.g_y[0].g_x[1].t.r_h ));
 sg13g2_dfrbp_1 \g.g_y[0].g_x[1].t.r_sc$_SDFFE_PN0P_  (.CLK(clknet_leaf_19_clk),
    .RESET_B(net208),
    .D(_0008_),
    .Q_N(_3209_),
    .Q(\g.g_y[0].g_x[1].t.out_sc ));
 sg13g2_dfrbp_1 \g.g_y[0].g_x[1].t.r_v$_SDFFE_PN0P_  (.CLK(clknet_leaf_19_clk),
    .RESET_B(net209),
    .D(_0009_),
    .Q_N(_3208_),
    .Q(\g.g_y[0].g_x[1].t.r_v ));
 sg13g2_dfrbp_1 \g.g_y[0].g_x[2].t.r_d$_SDFFE_PN0P_  (.CLK(clknet_leaf_19_clk),
    .RESET_B(net210),
    .D(_0010_),
    .Q_N(_3207_),
    .Q(\g.g_y[0].g_x[2].t.r_d ));
 sg13g2_dfrbp_1 \g.g_y[0].g_x[2].t.r_ghl$_SDFFE_PN0P_  (.CLK(clknet_leaf_19_clk),
    .RESET_B(net211),
    .D(_0011_),
    .Q_N(_3206_),
    .Q(\g.g_y[0].g_x[2].t.r_ghl ));
 sg13g2_dfrbp_1 \g.g_y[0].g_x[2].t.r_gnl$_SDFFE_PN0P_  (.CLK(clknet_leaf_20_clk),
    .RESET_B(net212),
    .D(_0012_),
    .Q_N(_3205_),
    .Q(\g.g_y[0].g_x[2].t.r_gnl ));
 sg13g2_dfrbp_1 \g.g_y[0].g_x[2].t.r_h$_SDFFE_PN0P_  (.CLK(clknet_leaf_20_clk),
    .RESET_B(net213),
    .D(_0013_),
    .Q_N(_3204_),
    .Q(\g.g_y[0].g_x[2].t.r_h ));
 sg13g2_dfrbp_1 \g.g_y[0].g_x[2].t.r_sc$_SDFFE_PN0P_  (.CLK(clknet_leaf_19_clk),
    .RESET_B(net214),
    .D(_0014_),
    .Q_N(_3203_),
    .Q(\g.g_y[0].g_x[2].t.out_sc ));
 sg13g2_dfrbp_1 \g.g_y[0].g_x[2].t.r_v$_SDFFE_PN0P_  (.CLK(clknet_leaf_19_clk),
    .RESET_B(net215),
    .D(_0015_),
    .Q_N(_3202_),
    .Q(\g.g_y[0].g_x[2].t.r_v ));
 sg13g2_dfrbp_1 \g.g_y[0].g_x[3].t.r_d$_SDFFE_PN0P_  (.CLK(clknet_leaf_20_clk),
    .RESET_B(net216),
    .D(_0016_),
    .Q_N(_3201_),
    .Q(\g.g_y[0].g_x[3].t.r_d ));
 sg13g2_dfrbp_1 \g.g_y[0].g_x[3].t.r_h$_SDFFE_PN0P_  (.CLK(clknet_leaf_20_clk),
    .RESET_B(net217),
    .D(_0017_),
    .Q_N(_3200_),
    .Q(\g.g_y[0].g_x[3].t.r_h ));
 sg13g2_dfrbp_1 \g.g_y[0].g_x[3].t.r_sc$_SDFFE_PN0P_  (.CLK(clknet_leaf_21_clk),
    .RESET_B(net218),
    .D(_0018_),
    .Q_N(_3199_),
    .Q(\g.g_y[0].g_x[3].t.out_sc ));
 sg13g2_dfrbp_1 \g.g_y[0].g_x[3].t.r_v$_SDFFE_PN0P_  (.CLK(clknet_leaf_21_clk),
    .RESET_B(net219),
    .D(_0019_),
    .Q_N(_3198_),
    .Q(\g.g_y[0].g_x[3].t.r_v ));
 sg13g2_dfrbp_1 \g.g_y[0].g_x[4].t.r_d$_SDFFE_PN0P_  (.CLK(clknet_leaf_21_clk),
    .RESET_B(net220),
    .D(_0020_),
    .Q_N(_3197_),
    .Q(\g.g_y[0].g_x[4].t.r_d ));
 sg13g2_dfrbp_1 \g.g_y[0].g_x[4].t.r_ghl$_SDFFE_PN0P_  (.CLK(clknet_leaf_21_clk),
    .RESET_B(net221),
    .D(_0021_),
    .Q_N(_3196_),
    .Q(\g.g_y[0].g_x[4].t.r_ghl ));
 sg13g2_dfrbp_1 \g.g_y[0].g_x[4].t.r_gnl$_SDFFE_PN0P_  (.CLK(clknet_leaf_14_clk),
    .RESET_B(net222),
    .D(_0022_),
    .Q_N(_3195_),
    .Q(\g.g_y[0].g_x[4].t.r_gnl ));
 sg13g2_dfrbp_1 \g.g_y[0].g_x[4].t.r_h$_SDFFE_PN0P_  (.CLK(clknet_leaf_20_clk),
    .RESET_B(net223),
    .D(_0023_),
    .Q_N(_3194_),
    .Q(\g.g_y[0].g_x[4].t.r_h ));
 sg13g2_dfrbp_1 \g.g_y[0].g_x[4].t.r_sc$_SDFFE_PN0P_  (.CLK(clknet_leaf_20_clk),
    .RESET_B(net224),
    .D(_0024_),
    .Q_N(_3193_),
    .Q(\g.g_y[0].g_x[4].t.out_sc ));
 sg13g2_dfrbp_1 \g.g_y[0].g_x[4].t.r_v$_SDFFE_PN0P_  (.CLK(clknet_leaf_21_clk),
    .RESET_B(net225),
    .D(_0025_),
    .Q_N(_3192_),
    .Q(\g.g_y[0].g_x[4].t.r_v ));
 sg13g2_dfrbp_1 \g.g_y[0].g_x[5].t.r_d$_SDFFE_PN0P_  (.CLK(clknet_leaf_15_clk),
    .RESET_B(net226),
    .D(_0026_),
    .Q_N(_3191_),
    .Q(\g.g_y[0].g_x[5].t.r_d ));
 sg13g2_dfrbp_1 \g.g_y[0].g_x[5].t.r_h$_SDFFE_PN0P_  (.CLK(clknet_leaf_17_clk),
    .RESET_B(net227),
    .D(_0027_),
    .Q_N(_3190_),
    .Q(\g.g_y[0].g_x[5].t.r_h ));
 sg13g2_dfrbp_1 \g.g_y[0].g_x[5].t.r_sc$_SDFFE_PN0P_  (.CLK(clknet_leaf_23_clk),
    .RESET_B(net228),
    .D(_0028_),
    .Q_N(_3189_),
    .Q(\g.g_y[0].g_x[5].t.out_sc ));
 sg13g2_dfrbp_1 \g.g_y[0].g_x[5].t.r_v$_SDFFE_PN0P_  (.CLK(clknet_leaf_17_clk),
    .RESET_B(net229),
    .D(_0029_),
    .Q_N(_3188_),
    .Q(\g.g_y[0].g_x[5].t.r_v ));
 sg13g2_dfrbp_1 \g.g_y[0].g_x[6].t.r_d$_SDFFE_PN0P_  (.CLK(clknet_leaf_17_clk),
    .RESET_B(net230),
    .D(_0030_),
    .Q_N(_3187_),
    .Q(\g.g_y[0].g_x[6].t.r_d ));
 sg13g2_dfrbp_1 \g.g_y[0].g_x[6].t.r_ghl$_SDFFE_PN0P_  (.CLK(clknet_leaf_17_clk),
    .RESET_B(net231),
    .D(_0031_),
    .Q_N(_3186_),
    .Q(\g.g_y[0].g_x[6].t.r_ghl ));
 sg13g2_dfrbp_1 \g.g_y[0].g_x[6].t.r_gnl$_SDFFE_PN0P_  (.CLK(clknet_leaf_17_clk),
    .RESET_B(net232),
    .D(_0032_),
    .Q_N(_3185_),
    .Q(\g.g_y[0].g_x[6].t.r_gnl ));
 sg13g2_dfrbp_1 \g.g_y[0].g_x[6].t.r_h$_SDFFE_PN0P_  (.CLK(clknet_leaf_18_clk),
    .RESET_B(net233),
    .D(_0033_),
    .Q_N(_3184_),
    .Q(\g.g_y[0].g_x[6].t.r_h ));
 sg13g2_dfrbp_1 \g.g_y[0].g_x[6].t.r_sc$_SDFFE_PN0P_  (.CLK(clknet_leaf_17_clk),
    .RESET_B(net234),
    .D(_0034_),
    .Q_N(_3183_),
    .Q(\g.g_y[0].g_x[6].t.out_sc ));
 sg13g2_dfrbp_1 \g.g_y[0].g_x[6].t.r_v$_SDFFE_PN0P_  (.CLK(clknet_leaf_17_clk),
    .RESET_B(net235),
    .D(_0035_),
    .Q_N(_3182_),
    .Q(\g.g_y[0].g_x[6].t.r_v ));
 sg13g2_dfrbp_1 \g.g_y[0].g_x[7].t.r_d$_SDFFE_PN0P_  (.CLK(clknet_leaf_16_clk),
    .RESET_B(net236),
    .D(_0036_),
    .Q_N(_3181_),
    .Q(\g.g_y[0].g_x[7].t.r_d ));
 sg13g2_dfrbp_1 \g.g_y[0].g_x[7].t.r_h$_SDFFE_PN0P_  (.CLK(clknet_leaf_18_clk),
    .RESET_B(net237),
    .D(_0037_),
    .Q_N(_3180_),
    .Q(\g.g_y[0].g_x[7].t.r_h ));
 sg13g2_dfrbp_1 \g.g_y[0].g_x[7].t.r_sc$_SDFFE_PN0P_  (.CLK(clknet_leaf_16_clk),
    .RESET_B(net238),
    .D(_0038_),
    .Q_N(_3179_),
    .Q(\g.g_y[0].g_x[7].t.out_sc ));
 sg13g2_dfrbp_1 \g.g_y[0].g_x[7].t.r_v$_SDFFE_PN0P_  (.CLK(clknet_leaf_17_clk),
    .RESET_B(net239),
    .D(_0039_),
    .Q_N(_3178_),
    .Q(\g.g_y[0].g_x[7].t.r_v ));
 sg13g2_dfrbp_1 \g.g_y[1].g_x[0].t.r_d$_SDFFE_PN0P_  (.CLK(clknet_leaf_21_clk),
    .RESET_B(net240),
    .D(_0040_),
    .Q_N(_3177_),
    .Q(\g.g_y[1].g_x[0].t.r_d ));
 sg13g2_dfrbp_1 \g.g_y[1].g_x[0].t.r_h$_SDFFE_PN0P_  (.CLK(clknet_leaf_20_clk),
    .RESET_B(net241),
    .D(_0041_),
    .Q_N(_3176_),
    .Q(\g.g_y[1].g_x[0].t.r_h ));
 sg13g2_dfrbp_1 \g.g_y[1].g_x[0].t.r_sc$_SDFFE_PN0P_  (.CLK(clknet_leaf_20_clk),
    .RESET_B(net242),
    .D(_0042_),
    .Q_N(_3175_),
    .Q(\g.g_y[1].g_x[0].t.out_sc ));
 sg13g2_dfrbp_1 \g.g_y[1].g_x[0].t.r_v$_SDFFE_PN0P_  (.CLK(clknet_leaf_21_clk),
    .RESET_B(net243),
    .D(_0043_),
    .Q_N(_3174_),
    .Q(\g.g_y[1].g_x[0].t.r_v ));
 sg13g2_dfrbp_1 \g.g_y[1].g_x[1].t.r_d$_SDFFE_PN0P_  (.CLK(clknet_leaf_26_clk),
    .RESET_B(net244),
    .D(_0044_),
    .Q_N(_3173_),
    .Q(\g.g_y[1].g_x[1].t.r_d ));
 sg13g2_dfrbp_1 \g.g_y[1].g_x[1].t.r_ghl$_SDFFE_PN0P_  (.CLK(clknet_leaf_26_clk),
    .RESET_B(net245),
    .D(_0045_),
    .Q_N(_3172_),
    .Q(\g.g_y[1].g_x[1].t.r_ghl ));
 sg13g2_dfrbp_1 \g.g_y[1].g_x[1].t.r_gnl$_SDFFE_PN0P_  (.CLK(clknet_leaf_22_clk),
    .RESET_B(net246),
    .D(_0046_),
    .Q_N(_3171_),
    .Q(\g.g_y[1].g_x[1].t.r_gnl ));
 sg13g2_dfrbp_1 \g.g_y[1].g_x[1].t.r_h$_SDFFE_PN0P_  (.CLK(clknet_leaf_21_clk),
    .RESET_B(net247),
    .D(_0047_),
    .Q_N(_3170_),
    .Q(\g.g_y[1].g_x[1].t.r_h ));
 sg13g2_dfrbp_1 \g.g_y[1].g_x[1].t.r_sc$_SDFFE_PN0P_  (.CLK(clknet_leaf_22_clk),
    .RESET_B(net248),
    .D(_0048_),
    .Q_N(_3169_),
    .Q(\g.g_y[1].g_x[1].t.out_sc ));
 sg13g2_dfrbp_1 \g.g_y[1].g_x[1].t.r_v$_SDFFE_PN0P_  (.CLK(clknet_leaf_22_clk),
    .RESET_B(net249),
    .D(_0049_),
    .Q_N(_3168_),
    .Q(\g.g_y[1].g_x[1].t.r_v ));
 sg13g2_dfrbp_1 \g.g_y[1].g_x[2].t.r_d$_SDFFE_PN0P_  (.CLK(clknet_leaf_22_clk),
    .RESET_B(net250),
    .D(_0050_),
    .Q_N(_3167_),
    .Q(\g.g_y[1].g_x[2].t.r_d ));
 sg13g2_dfrbp_1 \g.g_y[1].g_x[2].t.r_h$_SDFFE_PN0P_  (.CLK(clknet_leaf_22_clk),
    .RESET_B(net251),
    .D(_0051_),
    .Q_N(_3166_),
    .Q(\g.g_y[1].g_x[2].t.r_h ));
 sg13g2_dfrbp_1 \g.g_y[1].g_x[2].t.r_sc$_SDFFE_PN0P_  (.CLK(clknet_leaf_26_clk),
    .RESET_B(net252),
    .D(_0052_),
    .Q_N(_3165_),
    .Q(\g.g_y[1].g_x[2].t.out_sc ));
 sg13g2_dfrbp_1 \g.g_y[1].g_x[2].t.r_v$_SDFFE_PN0P_  (.CLK(clknet_leaf_22_clk),
    .RESET_B(net253),
    .D(_0053_),
    .Q_N(_3164_),
    .Q(\g.g_y[1].g_x[2].t.r_v ));
 sg13g2_dfrbp_1 \g.g_y[1].g_x[3].t.r_d$_SDFFE_PN0P_  (.CLK(clknet_leaf_23_clk),
    .RESET_B(net254),
    .D(_0054_),
    .Q_N(_3163_),
    .Q(\g.g_y[1].g_x[3].t.r_d ));
 sg13g2_dfrbp_1 \g.g_y[1].g_x[3].t.r_ghl$_SDFFE_PN0P_  (.CLK(clknet_leaf_23_clk),
    .RESET_B(net255),
    .D(_0055_),
    .Q_N(_3162_),
    .Q(\g.g_y[1].g_x[3].t.r_ghl ));
 sg13g2_dfrbp_1 \g.g_y[1].g_x[3].t.r_gnl$_SDFFE_PN0P_  (.CLK(clknet_leaf_22_clk),
    .RESET_B(net256),
    .D(_0056_),
    .Q_N(_3161_),
    .Q(\g.g_y[1].g_x[3].t.r_gnl ));
 sg13g2_dfrbp_1 \g.g_y[1].g_x[3].t.r_h$_SDFFE_PN0P_  (.CLK(clknet_leaf_22_clk),
    .RESET_B(net257),
    .D(_0057_),
    .Q_N(_3160_),
    .Q(\g.g_y[1].g_x[3].t.r_h ));
 sg13g2_dfrbp_1 \g.g_y[1].g_x[3].t.r_sc$_SDFFE_PN0P_  (.CLK(clknet_leaf_23_clk),
    .RESET_B(net258),
    .D(_0058_),
    .Q_N(_3159_),
    .Q(\g.g_y[1].g_x[3].t.out_sc ));
 sg13g2_dfrbp_1 \g.g_y[1].g_x[3].t.r_v$_SDFFE_PN0P_  (.CLK(clknet_leaf_23_clk),
    .RESET_B(net259),
    .D(_0059_),
    .Q_N(_3158_),
    .Q(\g.g_y[1].g_x[3].t.r_v ));
 sg13g2_dfrbp_1 \g.g_y[1].g_x[4].t.r_d$_SDFFE_PN0P_  (.CLK(clknet_leaf_23_clk),
    .RESET_B(net260),
    .D(_0060_),
    .Q_N(_3157_),
    .Q(\g.g_y[1].g_x[4].t.r_d ));
 sg13g2_dfrbp_1 \g.g_y[1].g_x[4].t.r_h$_SDFFE_PN0P_  (.CLK(clknet_leaf_24_clk),
    .RESET_B(net261),
    .D(_0061_),
    .Q_N(_3156_),
    .Q(\g.g_y[1].g_x[4].t.r_h ));
 sg13g2_dfrbp_1 \g.g_y[1].g_x[4].t.r_sc$_SDFFE_PN0P_  (.CLK(clknet_leaf_25_clk),
    .RESET_B(net262),
    .D(_0062_),
    .Q_N(_3155_),
    .Q(\g.g_y[1].g_x[4].t.out_sc ));
 sg13g2_dfrbp_1 \g.g_y[1].g_x[4].t.r_v$_SDFFE_PN0P_  (.CLK(clknet_leaf_24_clk),
    .RESET_B(net263),
    .D(_0063_),
    .Q_N(_3154_),
    .Q(\g.g_y[1].g_x[4].t.r_v ));
 sg13g2_dfrbp_1 \g.g_y[1].g_x[5].t.r_d$_SDFFE_PN0P_  (.CLK(clknet_leaf_26_clk),
    .RESET_B(net264),
    .D(_0064_),
    .Q_N(_3153_),
    .Q(\g.g_y[1].g_x[5].t.r_d ));
 sg13g2_dfrbp_1 \g.g_y[1].g_x[5].t.r_ghl$_SDFFE_PN0P_  (.CLK(clknet_leaf_26_clk),
    .RESET_B(net265),
    .D(_0065_),
    .Q_N(_3152_),
    .Q(\g.g_y[1].g_x[5].t.r_ghl ));
 sg13g2_dfrbp_1 \g.g_y[1].g_x[5].t.r_gnl$_SDFFE_PN0P_  (.CLK(clknet_leaf_26_clk),
    .RESET_B(net266),
    .D(_0066_),
    .Q_N(_3151_),
    .Q(\g.g_y[1].g_x[5].t.r_gnl ));
 sg13g2_dfrbp_1 \g.g_y[1].g_x[5].t.r_h$_SDFFE_PN0P_  (.CLK(clknet_leaf_26_clk),
    .RESET_B(net267),
    .D(_0067_),
    .Q_N(_3150_),
    .Q(\g.g_y[1].g_x[5].t.r_h ));
 sg13g2_dfrbp_1 \g.g_y[1].g_x[5].t.r_sc$_SDFFE_PN0P_  (.CLK(clknet_leaf_26_clk),
    .RESET_B(net268),
    .D(_0068_),
    .Q_N(_3149_),
    .Q(\g.g_y[1].g_x[5].t.out_sc ));
 sg13g2_dfrbp_1 \g.g_y[1].g_x[5].t.r_v$_SDFFE_PN0P_  (.CLK(clknet_leaf_28_clk),
    .RESET_B(net269),
    .D(_0069_),
    .Q_N(_3148_),
    .Q(\g.g_y[1].g_x[5].t.r_v ));
 sg13g2_dfrbp_1 \g.g_y[1].g_x[6].t.r_d$_SDFFE_PN0P_  (.CLK(clknet_leaf_24_clk),
    .RESET_B(net270),
    .D(_0070_),
    .Q_N(_3147_),
    .Q(\g.g_y[1].g_x[6].t.r_d ));
 sg13g2_dfrbp_1 \g.g_y[1].g_x[6].t.r_h$_SDFFE_PN0P_  (.CLK(clknet_leaf_25_clk),
    .RESET_B(net271),
    .D(_0071_),
    .Q_N(_3146_),
    .Q(\g.g_y[1].g_x[6].t.r_h ));
 sg13g2_dfrbp_1 \g.g_y[1].g_x[6].t.r_sc$_SDFFE_PN0P_  (.CLK(clknet_leaf_25_clk),
    .RESET_B(net272),
    .D(_0072_),
    .Q_N(_3145_),
    .Q(\g.g_y[1].g_x[6].t.out_sc ));
 sg13g2_dfrbp_1 \g.g_y[1].g_x[6].t.r_v$_SDFFE_PN0P_  (.CLK(clknet_leaf_25_clk),
    .RESET_B(net273),
    .D(_0073_),
    .Q_N(_3144_),
    .Q(\g.g_y[1].g_x[6].t.r_v ));
 sg13g2_dfrbp_1 \g.g_y[1].g_x[7].t.r_d$_SDFFE_PN0P_  (.CLK(clknet_leaf_25_clk),
    .RESET_B(net274),
    .D(_0074_),
    .Q_N(_3143_),
    .Q(\g.g_y[1].g_x[7].t.r_d ));
 sg13g2_dfrbp_1 \g.g_y[1].g_x[7].t.r_ghl$_SDFFE_PN0P_  (.CLK(clknet_leaf_25_clk),
    .RESET_B(net275),
    .D(_0075_),
    .Q_N(_3142_),
    .Q(\g.g_y[1].g_x[7].t.r_ghl ));
 sg13g2_dfrbp_1 \g.g_y[1].g_x[7].t.r_gnl$_SDFFE_PN0P_  (.CLK(clknet_leaf_24_clk),
    .RESET_B(net276),
    .D(_0076_),
    .Q_N(_3141_),
    .Q(\g.g_y[1].g_x[7].t.r_gnl ));
 sg13g2_dfrbp_1 \g.g_y[1].g_x[7].t.r_h$_SDFFE_PN0P_  (.CLK(clknet_leaf_28_clk),
    .RESET_B(net277),
    .D(_0077_),
    .Q_N(_3140_),
    .Q(\g.g_y[1].g_x[7].t.r_h ));
 sg13g2_dfrbp_1 \g.g_y[1].g_x[7].t.r_sc$_SDFFE_PN0P_  (.CLK(clknet_leaf_25_clk),
    .RESET_B(net278),
    .D(_0078_),
    .Q_N(_3139_),
    .Q(\g.g_y[1].g_x[7].t.out_sc ));
 sg13g2_dfrbp_1 \g.g_y[1].g_x[7].t.r_v$_SDFFE_PN0P_  (.CLK(clknet_leaf_27_clk),
    .RESET_B(net279),
    .D(_0079_),
    .Q_N(_3138_),
    .Q(\g.g_y[1].g_x[7].t.r_v ));
 sg13g2_dfrbp_1 \g.g_y[2].g_x[0].t.r_d$_SDFFE_PN0P_  (.CLK(clknet_leaf_27_clk),
    .RESET_B(net280),
    .D(_0080_),
    .Q_N(_3137_),
    .Q(\g.g_y[2].g_x[0].t.r_d ));
 sg13g2_dfrbp_1 \g.g_y[2].g_x[0].t.r_ghl$_SDFFE_PN0P_  (.CLK(clknet_leaf_27_clk),
    .RESET_B(net281),
    .D(_0081_),
    .Q_N(_3136_),
    .Q(\g.g_y[2].g_x[0].t.r_ghl ));
 sg13g2_dfrbp_1 \g.g_y[2].g_x[0].t.r_gnl$_SDFFE_PN0P_  (.CLK(clknet_leaf_27_clk),
    .RESET_B(net282),
    .D(_0082_),
    .Q_N(_3135_),
    .Q(\g.g_y[2].g_x[0].t.r_gnl ));
 sg13g2_dfrbp_1 \g.g_y[2].g_x[0].t.r_h$_SDFFE_PN0P_  (.CLK(clknet_leaf_28_clk),
    .RESET_B(net283),
    .D(_0083_),
    .Q_N(_3134_),
    .Q(\g.g_y[2].g_x[0].t.r_h ));
 sg13g2_dfrbp_1 \g.g_y[2].g_x[0].t.r_sc$_SDFFE_PN0P_  (.CLK(clknet_leaf_27_clk),
    .RESET_B(net284),
    .D(_0084_),
    .Q_N(_3133_),
    .Q(\g.g_y[2].g_x[0].t.out_sc ));
 sg13g2_dfrbp_1 \g.g_y[2].g_x[0].t.r_v$_SDFFE_PN0P_  (.CLK(clknet_leaf_27_clk),
    .RESET_B(net285),
    .D(_0085_),
    .Q_N(_3132_),
    .Q(\g.g_y[2].g_x[0].t.r_v ));
 sg13g2_dfrbp_1 \g.g_y[2].g_x[1].t.r_d$_SDFFE_PN0P_  (.CLK(clknet_leaf_29_clk),
    .RESET_B(net286),
    .D(_0086_),
    .Q_N(_3131_),
    .Q(\g.g_y[2].g_x[1].t.r_d ));
 sg13g2_dfrbp_1 \g.g_y[2].g_x[1].t.r_h$_SDFFE_PN0P_  (.CLK(clknet_leaf_27_clk),
    .RESET_B(net287),
    .D(_0087_),
    .Q_N(_3130_),
    .Q(\g.g_y[2].g_x[1].t.r_h ));
 sg13g2_dfrbp_1 \g.g_y[2].g_x[1].t.r_sc$_SDFFE_PN0P_  (.CLK(clknet_leaf_28_clk),
    .RESET_B(net288),
    .D(_0088_),
    .Q_N(_3129_),
    .Q(\g.g_y[2].g_x[1].t.out_sc ));
 sg13g2_dfrbp_1 \g.g_y[2].g_x[1].t.r_v$_SDFFE_PN0P_  (.CLK(clknet_leaf_27_clk),
    .RESET_B(net289),
    .D(_0089_),
    .Q_N(_3128_),
    .Q(\g.g_y[2].g_x[1].t.r_v ));
 sg13g2_dfrbp_1 \g.g_y[2].g_x[2].t.r_d$_SDFFE_PN0P_  (.CLK(clknet_leaf_29_clk),
    .RESET_B(net290),
    .D(_0090_),
    .Q_N(_3127_),
    .Q(\g.g_y[2].g_x[2].t.r_d ));
 sg13g2_dfrbp_1 \g.g_y[2].g_x[2].t.r_ghl$_SDFFE_PN0P_  (.CLK(clknet_leaf_29_clk),
    .RESET_B(net291),
    .D(_0091_),
    .Q_N(_3126_),
    .Q(\g.g_y[2].g_x[2].t.r_ghl ));
 sg13g2_dfrbp_1 \g.g_y[2].g_x[2].t.r_gnl$_SDFFE_PN0P_  (.CLK(clknet_leaf_29_clk),
    .RESET_B(net292),
    .D(_0092_),
    .Q_N(_3125_),
    .Q(\g.g_y[2].g_x[2].t.r_gnl ));
 sg13g2_dfrbp_1 \g.g_y[2].g_x[2].t.r_h$_SDFFE_PN0P_  (.CLK(clknet_leaf_29_clk),
    .RESET_B(net293),
    .D(_0093_),
    .Q_N(_3124_),
    .Q(\g.g_y[2].g_x[2].t.r_h ));
 sg13g2_dfrbp_1 \g.g_y[2].g_x[2].t.r_sc$_SDFFE_PN0P_  (.CLK(clknet_leaf_29_clk),
    .RESET_B(net294),
    .D(_0094_),
    .Q_N(_3123_),
    .Q(\g.g_y[2].g_x[2].t.out_sc ));
 sg13g2_dfrbp_1 \g.g_y[2].g_x[2].t.r_v$_SDFFE_PN0P_  (.CLK(clknet_leaf_28_clk),
    .RESET_B(net295),
    .D(_0095_),
    .Q_N(_3122_),
    .Q(\g.g_y[2].g_x[2].t.r_v ));
 sg13g2_dfrbp_1 \g.g_y[2].g_x[3].t.r_d$_SDFFE_PN0P_  (.CLK(clknet_leaf_29_clk),
    .RESET_B(net296),
    .D(_0096_),
    .Q_N(_3121_),
    .Q(\g.g_y[2].g_x[3].t.r_d ));
 sg13g2_dfrbp_1 \g.g_y[2].g_x[3].t.r_h$_SDFFE_PN0P_  (.CLK(clknet_leaf_29_clk),
    .RESET_B(net297),
    .D(_0097_),
    .Q_N(_3120_),
    .Q(\g.g_y[2].g_x[3].t.r_h ));
 sg13g2_dfrbp_1 \g.g_y[2].g_x[3].t.r_sc$_SDFFE_PN0P_  (.CLK(clknet_leaf_28_clk),
    .RESET_B(net298),
    .D(_0098_),
    .Q_N(_3119_),
    .Q(\g.g_y[2].g_x[3].t.out_sc ));
 sg13g2_dfrbp_1 \g.g_y[2].g_x[3].t.r_v$_SDFFE_PN0P_  (.CLK(clknet_leaf_30_clk),
    .RESET_B(net299),
    .D(_0099_),
    .Q_N(_3118_),
    .Q(\g.g_y[2].g_x[3].t.r_v ));
 sg13g2_dfrbp_1 \g.g_y[2].g_x[4].t.r_d$_SDFFE_PN0P_  (.CLK(clknet_leaf_30_clk),
    .RESET_B(net300),
    .D(_0100_),
    .Q_N(_3117_),
    .Q(\g.g_y[2].g_x[4].t.r_d ));
 sg13g2_dfrbp_1 \g.g_y[2].g_x[4].t.r_ghl$_SDFFE_PN0P_  (.CLK(clknet_leaf_25_clk),
    .RESET_B(net301),
    .D(_0101_),
    .Q_N(_3116_),
    .Q(\g.g_y[2].g_x[4].t.r_ghl ));
 sg13g2_dfrbp_1 \g.g_y[2].g_x[4].t.r_gnl$_SDFFE_PN0P_  (.CLK(clknet_leaf_33_clk),
    .RESET_B(net302),
    .D(_0102_),
    .Q_N(_3115_),
    .Q(\g.g_y[2].g_x[4].t.r_gnl ));
 sg13g2_dfrbp_1 \g.g_y[2].g_x[4].t.r_h$_SDFFE_PN0P_  (.CLK(clknet_leaf_30_clk),
    .RESET_B(net303),
    .D(_0103_),
    .Q_N(_3114_),
    .Q(\g.g_y[2].g_x[4].t.r_h ));
 sg13g2_dfrbp_1 \g.g_y[2].g_x[4].t.r_sc$_SDFFE_PN0P_  (.CLK(clknet_leaf_28_clk),
    .RESET_B(net304),
    .D(_0104_),
    .Q_N(_3113_),
    .Q(\g.g_y[2].g_x[4].t.out_sc ));
 sg13g2_dfrbp_1 \g.g_y[2].g_x[4].t.r_v$_SDFFE_PN0P_  (.CLK(clknet_leaf_33_clk),
    .RESET_B(net305),
    .D(_0105_),
    .Q_N(_3112_),
    .Q(\g.g_y[2].g_x[4].t.r_v ));
 sg13g2_dfrbp_1 \g.g_y[2].g_x[5].t.r_d$_SDFFE_PN0P_  (.CLK(clknet_leaf_30_clk),
    .RESET_B(net306),
    .D(_0106_),
    .Q_N(_3111_),
    .Q(\g.g_y[2].g_x[5].t.r_d ));
 sg13g2_dfrbp_1 \g.g_y[2].g_x[5].t.r_h$_SDFFE_PN0P_  (.CLK(clknet_leaf_30_clk),
    .RESET_B(net307),
    .D(_0107_),
    .Q_N(_3110_),
    .Q(\g.g_y[2].g_x[5].t.r_h ));
 sg13g2_dfrbp_1 \g.g_y[2].g_x[5].t.r_sc$_SDFFE_PN0P_  (.CLK(clknet_leaf_30_clk),
    .RESET_B(net308),
    .D(_0108_),
    .Q_N(_3109_),
    .Q(\g.g_y[2].g_x[5].t.out_sc ));
 sg13g2_dfrbp_1 \g.g_y[2].g_x[5].t.r_v$_SDFFE_PN0P_  (.CLK(clknet_leaf_28_clk),
    .RESET_B(net309),
    .D(_0109_),
    .Q_N(_3108_),
    .Q(\g.g_y[2].g_x[5].t.r_v ));
 sg13g2_dfrbp_1 \g.g_y[2].g_x[6].t.r_d$_SDFFE_PN0P_  (.CLK(clknet_leaf_31_clk),
    .RESET_B(net310),
    .D(_0110_),
    .Q_N(_3107_),
    .Q(\g.g_y[2].g_x[6].t.r_d ));
 sg13g2_dfrbp_1 \g.g_y[2].g_x[6].t.r_ghl$_SDFFE_PN0P_  (.CLK(clknet_leaf_30_clk),
    .RESET_B(net311),
    .D(_0111_),
    .Q_N(_3106_),
    .Q(\g.g_y[2].g_x[6].t.r_ghl ));
 sg13g2_dfrbp_1 \g.g_y[2].g_x[6].t.r_gnl$_SDFFE_PN0P_  (.CLK(clknet_leaf_30_clk),
    .RESET_B(net312),
    .D(_0112_),
    .Q_N(_3105_),
    .Q(\g.g_y[2].g_x[6].t.r_gnl ));
 sg13g2_dfrbp_1 \g.g_y[2].g_x[6].t.r_h$_SDFFE_PN0P_  (.CLK(clknet_leaf_31_clk),
    .RESET_B(net313),
    .D(_0113_),
    .Q_N(_3104_),
    .Q(\g.g_y[2].g_x[6].t.r_h ));
 sg13g2_dfrbp_1 \g.g_y[2].g_x[6].t.r_sc$_SDFFE_PN0P_  (.CLK(clknet_leaf_31_clk),
    .RESET_B(net314),
    .D(_0114_),
    .Q_N(_3103_),
    .Q(\g.g_y[2].g_x[6].t.out_sc ));
 sg13g2_dfrbp_1 \g.g_y[2].g_x[6].t.r_v$_SDFFE_PN0P_  (.CLK(clknet_leaf_31_clk),
    .RESET_B(net315),
    .D(_0115_),
    .Q_N(_3102_),
    .Q(\g.g_y[2].g_x[6].t.r_v ));
 sg13g2_dfrbp_1 \g.g_y[2].g_x[7].t.r_d$_SDFFE_PN0P_  (.CLK(clknet_leaf_31_clk),
    .RESET_B(net316),
    .D(_0116_),
    .Q_N(_3101_),
    .Q(\g.g_y[2].g_x[7].t.r_d ));
 sg13g2_dfrbp_1 \g.g_y[2].g_x[7].t.r_h$_SDFFE_PN0P_  (.CLK(clknet_leaf_31_clk),
    .RESET_B(net317),
    .D(_0117_),
    .Q_N(_3100_),
    .Q(\g.g_y[2].g_x[7].t.r_h ));
 sg13g2_dfrbp_1 \g.g_y[2].g_x[7].t.r_sc$_SDFFE_PN0P_  (.CLK(clknet_leaf_32_clk),
    .RESET_B(net318),
    .D(_0118_),
    .Q_N(_3099_),
    .Q(\g.g_y[2].g_x[7].t.out_sc ));
 sg13g2_dfrbp_1 \g.g_y[2].g_x[7].t.r_v$_SDFFE_PN0P_  (.CLK(clknet_leaf_31_clk),
    .RESET_B(net319),
    .D(_0119_),
    .Q_N(_3098_),
    .Q(\g.g_y[2].g_x[7].t.r_v ));
 sg13g2_dfrbp_1 \g.g_y[3].g_x[0].t.r_d$_SDFFE_PN0P_  (.CLK(clknet_leaf_24_clk),
    .RESET_B(net320),
    .D(_0120_),
    .Q_N(_3097_),
    .Q(\g.g_y[3].g_x[0].t.r_d ));
 sg13g2_dfrbp_1 \g.g_y[3].g_x[0].t.r_h$_SDFFE_PN0P_  (.CLK(clknet_leaf_33_clk),
    .RESET_B(net321),
    .D(_0121_),
    .Q_N(_3096_),
    .Q(\g.g_y[3].g_x[0].t.r_h ));
 sg13g2_dfrbp_1 \g.g_y[3].g_x[0].t.r_sc$_SDFFE_PN0P_  (.CLK(clknet_leaf_24_clk),
    .RESET_B(net322),
    .D(_0122_),
    .Q_N(_3095_),
    .Q(\g.g_y[3].g_x[0].t.out_sc ));
 sg13g2_dfrbp_1 \g.g_y[3].g_x[0].t.r_v$_SDFFE_PN0P_  (.CLK(clknet_leaf_33_clk),
    .RESET_B(net323),
    .D(_0123_),
    .Q_N(_3094_),
    .Q(\g.g_y[3].g_x[0].t.r_v ));
 sg13g2_dfrbp_1 \g.g_y[3].g_x[1].t.r_d$_SDFFE_PN0P_  (.CLK(clknet_leaf_34_clk),
    .RESET_B(net324),
    .D(_0124_),
    .Q_N(_3093_),
    .Q(\g.g_y[3].g_x[1].t.r_d ));
 sg13g2_dfrbp_1 \g.g_y[3].g_x[1].t.r_ghl$_SDFFE_PN0P_  (.CLK(clknet_leaf_34_clk),
    .RESET_B(net325),
    .D(_0125_),
    .Q_N(_3092_),
    .Q(\g.g_y[3].g_x[1].t.r_ghl ));
 sg13g2_dfrbp_1 \g.g_y[3].g_x[1].t.r_gnl$_SDFFE_PN0P_  (.CLK(clknet_leaf_34_clk),
    .RESET_B(net326),
    .D(_0126_),
    .Q_N(_3091_),
    .Q(\g.g_y[3].g_x[1].t.r_gnl ));
 sg13g2_dfrbp_1 \g.g_y[3].g_x[1].t.r_h$_SDFFE_PN0P_  (.CLK(clknet_leaf_33_clk),
    .RESET_B(net327),
    .D(_0127_),
    .Q_N(_3090_),
    .Q(\g.g_y[3].g_x[1].t.r_h ));
 sg13g2_dfrbp_1 \g.g_y[3].g_x[1].t.r_sc$_SDFFE_PN0P_  (.CLK(clknet_leaf_34_clk),
    .RESET_B(net328),
    .D(_0128_),
    .Q_N(_3089_),
    .Q(\g.g_y[3].g_x[1].t.out_sc ));
 sg13g2_dfrbp_1 \g.g_y[3].g_x[1].t.r_v$_SDFFE_PN0P_  (.CLK(clknet_leaf_35_clk),
    .RESET_B(net329),
    .D(_0129_),
    .Q_N(_3088_),
    .Q(\g.g_y[3].g_x[1].t.r_v ));
 sg13g2_dfrbp_1 \g.g_y[3].g_x[2].t.r_d$_SDFFE_PN0P_  (.CLK(clknet_leaf_33_clk),
    .RESET_B(net330),
    .D(_0130_),
    .Q_N(_3087_),
    .Q(\g.g_y[3].g_x[2].t.r_d ));
 sg13g2_dfrbp_1 \g.g_y[3].g_x[2].t.r_h$_SDFFE_PN0P_  (.CLK(clknet_leaf_33_clk),
    .RESET_B(net331),
    .D(_0131_),
    .Q_N(_3086_),
    .Q(\g.g_y[3].g_x[2].t.r_h ));
 sg13g2_dfrbp_1 \g.g_y[3].g_x[2].t.r_sc$_SDFFE_PN0P_  (.CLK(clknet_leaf_32_clk),
    .RESET_B(net332),
    .D(_0132_),
    .Q_N(_3085_),
    .Q(\g.g_y[3].g_x[2].t.out_sc ));
 sg13g2_dfrbp_1 \g.g_y[3].g_x[2].t.r_v$_SDFFE_PN0P_  (.CLK(clknet_leaf_33_clk),
    .RESET_B(net333),
    .D(_0133_),
    .Q_N(_3084_),
    .Q(\g.g_y[3].g_x[2].t.r_v ));
 sg13g2_dfrbp_1 \g.g_y[3].g_x[3].t.r_d$_SDFFE_PN0P_  (.CLK(clknet_leaf_32_clk),
    .RESET_B(net334),
    .D(_0134_),
    .Q_N(_3083_),
    .Q(\g.g_y[3].g_x[3].t.r_d ));
 sg13g2_dfrbp_1 \g.g_y[3].g_x[3].t.r_ghl$_SDFFE_PN0P_  (.CLK(clknet_leaf_31_clk),
    .RESET_B(net335),
    .D(_0135_),
    .Q_N(_3082_),
    .Q(\g.g_y[3].g_x[3].t.r_ghl ));
 sg13g2_dfrbp_1 \g.g_y[3].g_x[3].t.r_gnl$_SDFFE_PN0P_  (.CLK(clknet_leaf_32_clk),
    .RESET_B(net336),
    .D(_0136_),
    .Q_N(_3081_),
    .Q(\g.g_y[3].g_x[3].t.r_gnl ));
 sg13g2_dfrbp_1 \g.g_y[3].g_x[3].t.r_h$_SDFFE_PN0P_  (.CLK(clknet_leaf_32_clk),
    .RESET_B(net337),
    .D(_0137_),
    .Q_N(_3080_),
    .Q(\g.g_y[3].g_x[3].t.r_h ));
 sg13g2_dfrbp_1 \g.g_y[3].g_x[3].t.r_sc$_SDFFE_PN0P_  (.CLK(clknet_leaf_32_clk),
    .RESET_B(net338),
    .D(_0138_),
    .Q_N(_3079_),
    .Q(\g.g_y[3].g_x[3].t.out_sc ));
 sg13g2_dfrbp_1 \g.g_y[3].g_x[3].t.r_v$_SDFFE_PN0P_  (.CLK(clknet_leaf_32_clk),
    .RESET_B(net339),
    .D(_0139_),
    .Q_N(_3078_),
    .Q(\g.g_y[3].g_x[3].t.r_v ));
 sg13g2_dfrbp_1 \g.g_y[3].g_x[4].t.r_d$_SDFFE_PN0P_  (.CLK(clknet_leaf_36_clk),
    .RESET_B(net340),
    .D(_0140_),
    .Q_N(_3077_),
    .Q(\g.g_y[3].g_x[4].t.r_d ));
 sg13g2_dfrbp_1 \g.g_y[3].g_x[4].t.r_h$_SDFFE_PN0P_  (.CLK(clknet_leaf_36_clk),
    .RESET_B(net341),
    .D(_0141_),
    .Q_N(_3076_),
    .Q(\g.g_y[3].g_x[4].t.r_h ));
 sg13g2_dfrbp_1 \g.g_y[3].g_x[4].t.r_sc$_SDFFE_PN0P_  (.CLK(clknet_leaf_35_clk),
    .RESET_B(net342),
    .D(_0142_),
    .Q_N(_3075_),
    .Q(\g.g_y[3].g_x[4].t.out_sc ));
 sg13g2_dfrbp_1 \g.g_y[3].g_x[4].t.r_v$_SDFFE_PN0P_  (.CLK(clknet_leaf_34_clk),
    .RESET_B(net343),
    .D(_0143_),
    .Q_N(_3074_),
    .Q(\g.g_y[3].g_x[4].t.r_v ));
 sg13g2_dfrbp_1 \g.g_y[3].g_x[5].t.r_d$_SDFFE_PN0P_  (.CLK(clknet_leaf_37_clk),
    .RESET_B(net344),
    .D(_0144_),
    .Q_N(_3073_),
    .Q(\g.g_y[3].g_x[5].t.r_d ));
 sg13g2_dfrbp_1 \g.g_y[3].g_x[5].t.r_ghl$_SDFFE_PN0P_  (.CLK(clknet_leaf_35_clk),
    .RESET_B(net345),
    .D(_0145_),
    .Q_N(_3072_),
    .Q(\g.g_y[3].g_x[5].t.r_ghl ));
 sg13g2_dfrbp_1 \g.g_y[3].g_x[5].t.r_gnl$_SDFFE_PN0P_  (.CLK(clknet_leaf_36_clk),
    .RESET_B(net346),
    .D(_0146_),
    .Q_N(_3071_),
    .Q(\g.g_y[3].g_x[5].t.r_gnl ));
 sg13g2_dfrbp_1 \g.g_y[3].g_x[5].t.r_h$_SDFFE_PN0P_  (.CLK(clknet_leaf_37_clk),
    .RESET_B(net347),
    .D(_0147_),
    .Q_N(_3070_),
    .Q(\g.g_y[3].g_x[5].t.r_h ));
 sg13g2_dfrbp_1 \g.g_y[3].g_x[5].t.r_sc$_SDFFE_PN0P_  (.CLK(clknet_leaf_36_clk),
    .RESET_B(net348),
    .D(_0148_),
    .Q_N(_3069_),
    .Q(\g.g_y[3].g_x[5].t.out_sc ));
 sg13g2_dfrbp_1 \g.g_y[3].g_x[5].t.r_v$_SDFFE_PN0P_  (.CLK(clknet_leaf_37_clk),
    .RESET_B(net349),
    .D(_0149_),
    .Q_N(_3068_),
    .Q(\g.g_y[3].g_x[5].t.r_v ));
 sg13g2_dfrbp_1 \g.g_y[3].g_x[6].t.r_d$_SDFFE_PN0P_  (.CLK(clknet_leaf_36_clk),
    .RESET_B(net350),
    .D(_0150_),
    .Q_N(_3067_),
    .Q(\g.g_y[3].g_x[6].t.r_d ));
 sg13g2_dfrbp_1 \g.g_y[3].g_x[6].t.r_h$_SDFFE_PN0P_  (.CLK(clknet_leaf_37_clk),
    .RESET_B(net351),
    .D(_0151_),
    .Q_N(_3066_),
    .Q(\g.g_y[3].g_x[6].t.r_h ));
 sg13g2_dfrbp_1 \g.g_y[3].g_x[6].t.r_sc$_SDFFE_PN0P_  (.CLK(clknet_leaf_38_clk),
    .RESET_B(net352),
    .D(_0152_),
    .Q_N(_3065_),
    .Q(\g.g_y[3].g_x[6].t.out_sc ));
 sg13g2_dfrbp_1 \g.g_y[3].g_x[6].t.r_v$_SDFFE_PN0P_  (.CLK(clknet_leaf_38_clk),
    .RESET_B(net353),
    .D(_0153_),
    .Q_N(_3064_),
    .Q(\g.g_y[3].g_x[6].t.r_v ));
 sg13g2_dfrbp_1 \g.g_y[3].g_x[7].t.r_d$_SDFFE_PN0P_  (.CLK(clknet_leaf_36_clk),
    .RESET_B(net354),
    .D(_0154_),
    .Q_N(_3063_),
    .Q(\g.g_y[3].g_x[7].t.r_d ));
 sg13g2_dfrbp_1 \g.g_y[3].g_x[7].t.r_ghl$_SDFFE_PN0P_  (.CLK(clknet_leaf_36_clk),
    .RESET_B(net355),
    .D(_0155_),
    .Q_N(_3062_),
    .Q(\g.g_y[3].g_x[7].t.r_ghl ));
 sg13g2_dfrbp_1 \g.g_y[3].g_x[7].t.r_gnl$_SDFFE_PN0P_  (.CLK(clknet_leaf_32_clk),
    .RESET_B(net356),
    .D(_0156_),
    .Q_N(_3061_),
    .Q(\g.g_y[3].g_x[7].t.r_gnl ));
 sg13g2_dfrbp_1 \g.g_y[3].g_x[7].t.r_h$_SDFFE_PN0P_  (.CLK(clknet_leaf_37_clk),
    .RESET_B(net357),
    .D(_0157_),
    .Q_N(_3060_),
    .Q(\g.g_y[3].g_x[7].t.r_h ));
 sg13g2_dfrbp_1 \g.g_y[3].g_x[7].t.r_sc$_SDFFE_PN0P_  (.CLK(clknet_leaf_37_clk),
    .RESET_B(net358),
    .D(_0158_),
    .Q_N(_3059_),
    .Q(\g.g_y[3].g_x[7].t.out_sc ));
 sg13g2_dfrbp_1 \g.g_y[3].g_x[7].t.r_v$_SDFFE_PN0P_  (.CLK(clknet_leaf_36_clk),
    .RESET_B(net359),
    .D(_0159_),
    .Q_N(_3058_),
    .Q(\g.g_y[3].g_x[7].t.r_v ));
 sg13g2_dfrbp_1 \g.g_y[4].g_x[0].t.r_d$_SDFFE_PN0P_  (.CLK(clknet_leaf_3_clk),
    .RESET_B(net360),
    .D(_0160_),
    .Q_N(_3057_),
    .Q(\g.g_y[4].g_x[0].t.r_d ));
 sg13g2_dfrbp_1 \g.g_y[4].g_x[0].t.r_ghl$_SDFFE_PN0P_  (.CLK(clknet_leaf_34_clk),
    .RESET_B(net361),
    .D(_0161_),
    .Q_N(_3056_),
    .Q(\g.g_y[4].g_x[0].t.r_ghl ));
 sg13g2_dfrbp_1 \g.g_y[4].g_x[0].t.r_gnl$_SDFFE_PN0P_  (.CLK(clknet_leaf_3_clk),
    .RESET_B(net362),
    .D(_0162_),
    .Q_N(_3055_),
    .Q(\g.g_y[4].g_x[0].t.r_gnl ));
 sg13g2_dfrbp_1 \g.g_y[4].g_x[0].t.r_h$_SDFFE_PN0P_  (.CLK(clknet_leaf_34_clk),
    .RESET_B(net363),
    .D(_0163_),
    .Q_N(_3054_),
    .Q(\g.g_y[4].g_x[0].t.r_h ));
 sg13g2_dfrbp_1 \g.g_y[4].g_x[0].t.r_sc$_SDFFE_PN0P_  (.CLK(clknet_leaf_34_clk),
    .RESET_B(net364),
    .D(_0164_),
    .Q_N(_3053_),
    .Q(\g.g_y[4].g_x[0].t.out_sc ));
 sg13g2_dfrbp_1 \g.g_y[4].g_x[0].t.r_v$_SDFFE_PN0P_  (.CLK(clknet_leaf_35_clk),
    .RESET_B(net365),
    .D(_0165_),
    .Q_N(_3052_),
    .Q(\g.g_y[4].g_x[0].t.r_v ));
 sg13g2_dfrbp_1 \g.g_y[4].g_x[1].t.r_d$_SDFFE_PN0P_  (.CLK(clknet_leaf_3_clk),
    .RESET_B(net366),
    .D(_0166_),
    .Q_N(_3051_),
    .Q(\g.g_y[4].g_x[1].t.r_d ));
 sg13g2_dfrbp_1 \g.g_y[4].g_x[1].t.r_h$_SDFFE_PN0P_  (.CLK(clknet_leaf_35_clk),
    .RESET_B(net367),
    .D(_0167_),
    .Q_N(_3050_),
    .Q(\g.g_y[4].g_x[1].t.r_h ));
 sg13g2_dfrbp_1 \g.g_y[4].g_x[1].t.r_sc$_SDFFE_PN0P_  (.CLK(clknet_leaf_35_clk),
    .RESET_B(net368),
    .D(_0168_),
    .Q_N(_3049_),
    .Q(\g.g_y[4].g_x[1].t.out_sc ));
 sg13g2_dfrbp_1 \g.g_y[4].g_x[1].t.r_v$_SDFFE_PN0P_  (.CLK(clknet_leaf_2_clk),
    .RESET_B(net369),
    .D(_0169_),
    .Q_N(_3048_),
    .Q(\g.g_y[4].g_x[1].t.r_v ));
 sg13g2_dfrbp_1 \g.g_y[4].g_x[2].t.r_d$_SDFFE_PN0P_  (.CLK(clknet_leaf_37_clk),
    .RESET_B(net370),
    .D(_0170_),
    .Q_N(_3047_),
    .Q(\g.g_y[4].g_x[2].t.r_d ));
 sg13g2_dfrbp_1 \g.g_y[4].g_x[2].t.r_ghl$_SDFFE_PN0P_  (.CLK(clknet_leaf_35_clk),
    .RESET_B(net371),
    .D(_0171_),
    .Q_N(_3046_),
    .Q(\g.g_y[4].g_x[2].t.r_ghl ));
 sg13g2_dfrbp_1 \g.g_y[4].g_x[2].t.r_gnl$_SDFFE_PN0P_  (.CLK(clknet_leaf_38_clk),
    .RESET_B(net372),
    .D(_0172_),
    .Q_N(_3045_),
    .Q(\g.g_y[4].g_x[2].t.r_gnl ));
 sg13g2_dfrbp_1 \g.g_y[4].g_x[2].t.r_h$_SDFFE_PN0P_  (.CLK(clknet_leaf_38_clk),
    .RESET_B(net373),
    .D(_0173_),
    .Q_N(_3044_),
    .Q(\g.g_y[4].g_x[2].t.r_h ));
 sg13g2_dfrbp_1 \g.g_y[4].g_x[2].t.r_sc$_SDFFE_PN0P_  (.CLK(clknet_leaf_38_clk),
    .RESET_B(net374),
    .D(_0174_),
    .Q_N(_3043_),
    .Q(\g.g_y[4].g_x[2].t.out_sc ));
 sg13g2_dfrbp_1 \g.g_y[4].g_x[2].t.r_v$_SDFFE_PN0P_  (.CLK(clknet_leaf_37_clk),
    .RESET_B(net375),
    .D(_0175_),
    .Q_N(_3042_),
    .Q(\g.g_y[4].g_x[2].t.r_v ));
 sg13g2_dfrbp_1 \g.g_y[4].g_x[3].t.r_d$_SDFFE_PN0P_  (.CLK(clknet_leaf_38_clk),
    .RESET_B(net376),
    .D(_0176_),
    .Q_N(_3041_),
    .Q(\g.g_y[4].g_x[3].t.r_d ));
 sg13g2_dfrbp_1 \g.g_y[4].g_x[3].t.r_h$_SDFFE_PN0P_  (.CLK(clknet_leaf_38_clk),
    .RESET_B(net377),
    .D(_0177_),
    .Q_N(_3040_),
    .Q(\g.g_y[4].g_x[3].t.r_h ));
 sg13g2_dfrbp_1 \g.g_y[4].g_x[3].t.r_sc$_SDFFE_PN0P_  (.CLK(clknet_leaf_35_clk),
    .RESET_B(net378),
    .D(_0178_),
    .Q_N(_3039_),
    .Q(\g.g_y[4].g_x[3].t.out_sc ));
 sg13g2_dfrbp_1 \g.g_y[4].g_x[3].t.r_v$_SDFFE_PN0P_  (.CLK(clknet_leaf_38_clk),
    .RESET_B(net379),
    .D(_0179_),
    .Q_N(_3038_),
    .Q(\g.g_y[4].g_x[3].t.r_v ));
 sg13g2_dfrbp_1 \g.g_y[4].g_x[4].t.r_d$_SDFFE_PN0P_  (.CLK(clknet_leaf_39_clk),
    .RESET_B(net380),
    .D(_0180_),
    .Q_N(_3037_),
    .Q(\g.g_y[4].g_x[4].t.r_d ));
 sg13g2_dfrbp_1 \g.g_y[4].g_x[4].t.r_ghl$_SDFFE_PN0P_  (.CLK(clknet_leaf_39_clk),
    .RESET_B(net381),
    .D(_0181_),
    .Q_N(_3036_),
    .Q(\g.g_y[4].g_x[4].t.r_ghl ));
 sg13g2_dfrbp_1 \g.g_y[4].g_x[4].t.r_gnl$_SDFFE_PN0P_  (.CLK(clknet_leaf_0_clk),
    .RESET_B(net382),
    .D(_0182_),
    .Q_N(_3035_),
    .Q(\g.g_y[4].g_x[4].t.r_gnl ));
 sg13g2_dfrbp_1 \g.g_y[4].g_x[4].t.r_h$_SDFFE_PN0P_  (.CLK(clknet_leaf_39_clk),
    .RESET_B(net383),
    .D(_0183_),
    .Q_N(_3034_),
    .Q(\g.g_y[4].g_x[4].t.r_h ));
 sg13g2_dfrbp_1 \g.g_y[4].g_x[4].t.r_sc$_SDFFE_PN0P_  (.CLK(clknet_leaf_39_clk),
    .RESET_B(net384),
    .D(_0184_),
    .Q_N(_3033_),
    .Q(\g.g_y[4].g_x[4].t.out_sc ));
 sg13g2_dfrbp_1 \g.g_y[4].g_x[4].t.r_v$_SDFFE_PN0P_  (.CLK(clknet_leaf_0_clk),
    .RESET_B(net385),
    .D(_0185_),
    .Q_N(_3032_),
    .Q(\g.g_y[4].g_x[4].t.r_v ));
 sg13g2_dfrbp_1 \g.g_y[4].g_x[5].t.r_d$_SDFFE_PN0P_  (.CLK(clknet_leaf_39_clk),
    .RESET_B(net386),
    .D(_0186_),
    .Q_N(_3031_),
    .Q(\g.g_y[4].g_x[5].t.r_d ));
 sg13g2_dfrbp_1 \g.g_y[4].g_x[5].t.r_h$_SDFFE_PN0P_  (.CLK(clknet_leaf_39_clk),
    .RESET_B(net387),
    .D(_0187_),
    .Q_N(_3030_),
    .Q(\g.g_y[4].g_x[5].t.r_h ));
 sg13g2_dfrbp_1 \g.g_y[4].g_x[5].t.r_sc$_SDFFE_PN0P_  (.CLK(clknet_leaf_39_clk),
    .RESET_B(net388),
    .D(_0188_),
    .Q_N(_3029_),
    .Q(\g.g_y[4].g_x[5].t.out_sc ));
 sg13g2_dfrbp_1 \g.g_y[4].g_x[5].t.r_v$_SDFFE_PN0P_  (.CLK(clknet_leaf_39_clk),
    .RESET_B(net389),
    .D(_0189_),
    .Q_N(_3028_),
    .Q(\g.g_y[4].g_x[5].t.r_v ));
 sg13g2_dfrbp_1 \g.g_y[4].g_x[6].t.r_d$_SDFFE_PN0P_  (.CLK(clknet_leaf_0_clk),
    .RESET_B(net390),
    .D(_0190_),
    .Q_N(_3027_),
    .Q(\g.g_y[4].g_x[6].t.r_d ));
 sg13g2_dfrbp_1 \g.g_y[4].g_x[6].t.r_ghl$_SDFFE_PN0P_  (.CLK(clknet_leaf_0_clk),
    .RESET_B(net391),
    .D(_0191_),
    .Q_N(_3026_),
    .Q(\g.g_y[4].g_x[6].t.r_ghl ));
 sg13g2_dfrbp_1 \g.g_y[4].g_x[6].t.r_gnl$_SDFFE_PN0P_  (.CLK(clknet_leaf_2_clk),
    .RESET_B(net392),
    .D(_0192_),
    .Q_N(_3025_),
    .Q(\g.g_y[4].g_x[6].t.r_gnl ));
 sg13g2_dfrbp_1 \g.g_y[4].g_x[6].t.r_h$_SDFFE_PN0P_  (.CLK(clknet_leaf_2_clk),
    .RESET_B(net393),
    .D(_0193_),
    .Q_N(_3024_),
    .Q(\g.g_y[4].g_x[6].t.r_h ));
 sg13g2_dfrbp_1 \g.g_y[4].g_x[6].t.r_sc$_SDFFE_PN0P_  (.CLK(clknet_leaf_0_clk),
    .RESET_B(net394),
    .D(_0194_),
    .Q_N(_3023_),
    .Q(\g.g_y[4].g_x[6].t.out_sc ));
 sg13g2_dfrbp_1 \g.g_y[4].g_x[6].t.r_v$_SDFFE_PN0P_  (.CLK(clknet_leaf_0_clk),
    .RESET_B(net395),
    .D(_0195_),
    .Q_N(_3022_),
    .Q(\g.g_y[4].g_x[6].t.r_v ));
 sg13g2_dfrbp_1 \g.g_y[4].g_x[7].t.r_d$_SDFFE_PN0P_  (.CLK(clknet_leaf_3_clk),
    .RESET_B(net396),
    .D(_0196_),
    .Q_N(_3021_),
    .Q(\g.g_y[4].g_x[7].t.r_d ));
 sg13g2_dfrbp_1 \g.g_y[4].g_x[7].t.r_h$_SDFFE_PN0P_  (.CLK(clknet_leaf_2_clk),
    .RESET_B(net397),
    .D(_0197_),
    .Q_N(_3020_),
    .Q(\g.g_y[4].g_x[7].t.r_h ));
 sg13g2_dfrbp_1 \g.g_y[4].g_x[7].t.r_sc$_SDFFE_PN0P_  (.CLK(clknet_leaf_2_clk),
    .RESET_B(net398),
    .D(_0198_),
    .Q_N(_3019_),
    .Q(\g.g_y[4].g_x[7].t.out_sc ));
 sg13g2_dfrbp_1 \g.g_y[4].g_x[7].t.r_v$_SDFFE_PN0P_  (.CLK(clknet_leaf_3_clk),
    .RESET_B(net399),
    .D(_0199_),
    .Q_N(_3018_),
    .Q(\g.g_y[4].g_x[7].t.r_v ));
 sg13g2_dfrbp_1 \g.g_y[5].g_x[0].t.r_d$_SDFFE_PN0P_  (.CLK(clknet_leaf_4_clk),
    .RESET_B(net400),
    .D(_0200_),
    .Q_N(_3017_),
    .Q(\g.g_y[5].g_x[0].t.r_d ));
 sg13g2_dfrbp_1 \g.g_y[5].g_x[0].t.r_h$_SDFFE_PN0P_  (.CLK(clknet_leaf_3_clk),
    .RESET_B(net401),
    .D(_0201_),
    .Q_N(_3016_),
    .Q(\g.g_y[5].g_x[0].t.r_h ));
 sg13g2_dfrbp_1 \g.g_y[5].g_x[0].t.r_sc$_SDFFE_PN0P_  (.CLK(clknet_leaf_3_clk),
    .RESET_B(net402),
    .D(_0202_),
    .Q_N(_3015_),
    .Q(\g.g_y[5].g_x[0].t.out_sc ));
 sg13g2_dfrbp_1 \g.g_y[5].g_x[0].t.r_v$_SDFFE_PN0P_  (.CLK(clknet_leaf_4_clk),
    .RESET_B(net403),
    .D(_0203_),
    .Q_N(_3014_),
    .Q(\g.g_y[5].g_x[0].t.r_v ));
 sg13g2_dfrbp_1 \g.g_y[5].g_x[1].t.r_d$_SDFFE_PN0P_  (.CLK(clknet_leaf_6_clk),
    .RESET_B(net404),
    .D(_0204_),
    .Q_N(_3013_),
    .Q(\g.g_y[5].g_x[1].t.r_d ));
 sg13g2_dfrbp_1 \g.g_y[5].g_x[1].t.r_ghl$_SDFFE_PN0P_  (.CLK(clknet_leaf_5_clk),
    .RESET_B(net405),
    .D(_0205_),
    .Q_N(_3012_),
    .Q(\g.g_y[5].g_x[1].t.r_ghl ));
 sg13g2_dfrbp_1 \g.g_y[5].g_x[1].t.r_gnl$_SDFFE_PN0P_  (.CLK(clknet_leaf_5_clk),
    .RESET_B(net406),
    .D(_0206_),
    .Q_N(_3011_),
    .Q(\g.g_y[5].g_x[1].t.r_gnl ));
 sg13g2_dfrbp_1 \g.g_y[5].g_x[1].t.r_h$_SDFFE_PN0P_  (.CLK(clknet_leaf_1_clk),
    .RESET_B(net407),
    .D(_0207_),
    .Q_N(_3010_),
    .Q(\g.g_y[5].g_x[1].t.r_h ));
 sg13g2_dfrbp_1 \g.g_y[5].g_x[1].t.r_sc$_SDFFE_PN0P_  (.CLK(clknet_leaf_5_clk),
    .RESET_B(net408),
    .D(_0208_),
    .Q_N(_3009_),
    .Q(\g.g_y[5].g_x[1].t.out_sc ));
 sg13g2_dfrbp_1 \g.g_y[5].g_x[1].t.r_v$_SDFFE_PN0P_  (.CLK(clknet_leaf_2_clk),
    .RESET_B(net409),
    .D(_0209_),
    .Q_N(_3008_),
    .Q(\g.g_y[5].g_x[1].t.r_v ));
 sg13g2_dfrbp_1 \g.g_y[5].g_x[2].t.r_d$_SDFFE_PN0P_  (.CLK(clknet_leaf_2_clk),
    .RESET_B(net410),
    .D(_0210_),
    .Q_N(_3007_),
    .Q(\g.g_y[5].g_x[2].t.r_d ));
 sg13g2_dfrbp_1 \g.g_y[5].g_x[2].t.r_h$_SDFFE_PN0P_  (.CLK(clknet_leaf_1_clk),
    .RESET_B(net411),
    .D(_0211_),
    .Q_N(_3006_),
    .Q(\g.g_y[5].g_x[2].t.r_h ));
 sg13g2_dfrbp_1 \g.g_y[5].g_x[2].t.r_sc$_SDFFE_PN0P_  (.CLK(clknet_leaf_2_clk),
    .RESET_B(net412),
    .D(_0212_),
    .Q_N(_3005_),
    .Q(\g.g_y[5].g_x[2].t.out_sc ));
 sg13g2_dfrbp_1 \g.g_y[5].g_x[2].t.r_v$_SDFFE_PN0P_  (.CLK(clknet_leaf_1_clk),
    .RESET_B(net413),
    .D(_0213_),
    .Q_N(_3004_),
    .Q(\g.g_y[5].g_x[2].t.r_v ));
 sg13g2_dfrbp_1 \g.g_y[5].g_x[3].t.r_d$_SDFFE_PN0P_  (.CLK(clknet_leaf_1_clk),
    .RESET_B(net414),
    .D(_0214_),
    .Q_N(_3003_),
    .Q(\g.g_y[5].g_x[3].t.r_d ));
 sg13g2_dfrbp_1 \g.g_y[5].g_x[3].t.r_ghl$_SDFFE_PN0P_  (.CLK(clknet_leaf_1_clk),
    .RESET_B(net415),
    .D(_0215_),
    .Q_N(_3002_),
    .Q(\g.g_y[5].g_x[3].t.r_ghl ));
 sg13g2_dfrbp_1 \g.g_y[5].g_x[3].t.r_gnl$_SDFFE_PN0P_  (.CLK(clknet_leaf_1_clk),
    .RESET_B(net416),
    .D(_0216_),
    .Q_N(_3001_),
    .Q(\g.g_y[5].g_x[3].t.r_gnl ));
 sg13g2_dfrbp_1 \g.g_y[5].g_x[3].t.r_h$_SDFFE_PN0P_  (.CLK(clknet_leaf_1_clk),
    .RESET_B(net417),
    .D(_0217_),
    .Q_N(_3000_),
    .Q(\g.g_y[5].g_x[3].t.r_h ));
 sg13g2_dfrbp_1 \g.g_y[5].g_x[3].t.r_sc$_SDFFE_PN0P_  (.CLK(clknet_leaf_1_clk),
    .RESET_B(net418),
    .D(_0218_),
    .Q_N(_2999_),
    .Q(\g.g_y[5].g_x[3].t.out_sc ));
 sg13g2_dfrbp_1 \g.g_y[5].g_x[3].t.r_v$_SDFFE_PN0P_  (.CLK(clknet_leaf_6_clk),
    .RESET_B(net419),
    .D(_0219_),
    .Q_N(_2998_),
    .Q(\g.g_y[5].g_x[3].t.r_v ));
 sg13g2_dfrbp_1 \g.g_y[5].g_x[4].t.r_d$_SDFFE_PN0P_  (.CLK(clknet_leaf_0_clk),
    .RESET_B(net420),
    .D(_0220_),
    .Q_N(_2997_),
    .Q(\g.g_y[5].g_x[4].t.r_d ));
 sg13g2_dfrbp_1 \g.g_y[5].g_x[4].t.r_h$_SDFFE_PN0P_  (.CLK(clknet_leaf_6_clk),
    .RESET_B(net421),
    .D(_0221_),
    .Q_N(_2996_),
    .Q(\g.g_y[5].g_x[4].t.r_h ));
 sg13g2_dfrbp_1 \g.g_y[5].g_x[4].t.r_sc$_SDFFE_PN0P_  (.CLK(clknet_leaf_0_clk),
    .RESET_B(net422),
    .D(_0222_),
    .Q_N(_2995_),
    .Q(\g.g_y[5].g_x[4].t.out_sc ));
 sg13g2_dfrbp_1 \g.g_y[5].g_x[4].t.r_v$_SDFFE_PN0P_  (.CLK(clknet_leaf_6_clk),
    .RESET_B(net423),
    .D(_0223_),
    .Q_N(_2994_),
    .Q(\g.g_y[5].g_x[4].t.r_v ));
 sg13g2_dfrbp_1 \g.g_y[5].g_x[5].t.r_d$_SDFFE_PN0P_  (.CLK(clknet_leaf_6_clk),
    .RESET_B(net424),
    .D(_0224_),
    .Q_N(_2993_),
    .Q(\g.g_y[5].g_x[5].t.r_d ));
 sg13g2_dfrbp_1 \g.g_y[5].g_x[5].t.r_ghl$_SDFFE_PN0P_  (.CLK(clknet_leaf_5_clk),
    .RESET_B(net425),
    .D(_0225_),
    .Q_N(_2992_),
    .Q(\g.g_y[5].g_x[5].t.r_ghl ));
 sg13g2_dfrbp_1 \g.g_y[5].g_x[5].t.r_gnl$_SDFFE_PN0P_  (.CLK(clknet_leaf_5_clk),
    .RESET_B(net426),
    .D(_0226_),
    .Q_N(_2991_),
    .Q(\g.g_y[5].g_x[5].t.r_gnl ));
 sg13g2_dfrbp_1 \g.g_y[5].g_x[5].t.r_h$_SDFFE_PN0P_  (.CLK(clknet_leaf_6_clk),
    .RESET_B(net427),
    .D(_0227_),
    .Q_N(_2990_),
    .Q(\g.g_y[5].g_x[5].t.r_h ));
 sg13g2_dfrbp_1 \g.g_y[5].g_x[5].t.r_sc$_SDFFE_PN0P_  (.CLK(clknet_leaf_6_clk),
    .RESET_B(net428),
    .D(_0228_),
    .Q_N(_2989_),
    .Q(\g.g_y[5].g_x[5].t.out_sc ));
 sg13g2_dfrbp_1 \g.g_y[5].g_x[5].t.r_v$_SDFFE_PN0P_  (.CLK(clknet_leaf_6_clk),
    .RESET_B(net429),
    .D(_0229_),
    .Q_N(_2988_),
    .Q(\g.g_y[5].g_x[5].t.r_v ));
 sg13g2_dfrbp_1 \g.g_y[5].g_x[6].t.r_d$_SDFFE_PN0P_  (.CLK(clknet_leaf_8_clk),
    .RESET_B(net430),
    .D(_0230_),
    .Q_N(_2987_),
    .Q(\g.g_y[5].g_x[6].t.r_d ));
 sg13g2_dfrbp_1 \g.g_y[5].g_x[6].t.r_h$_SDFFE_PN0P_  (.CLK(clknet_leaf_7_clk),
    .RESET_B(net431),
    .D(_0231_),
    .Q_N(_2986_),
    .Q(\g.g_y[5].g_x[6].t.r_h ));
 sg13g2_dfrbp_1 \g.g_y[5].g_x[6].t.r_sc$_SDFFE_PN0P_  (.CLK(clknet_leaf_7_clk),
    .RESET_B(net432),
    .D(_0232_),
    .Q_N(_2985_),
    .Q(\g.g_y[5].g_x[6].t.out_sc ));
 sg13g2_dfrbp_1 \g.g_y[5].g_x[6].t.r_v$_SDFFE_PN0P_  (.CLK(clknet_leaf_7_clk),
    .RESET_B(net433),
    .D(_0233_),
    .Q_N(_2984_),
    .Q(\g.g_y[5].g_x[6].t.r_v ));
 sg13g2_dfrbp_1 \g.g_y[5].g_x[7].t.r_d$_SDFFE_PN0P_  (.CLK(clknet_leaf_8_clk),
    .RESET_B(net434),
    .D(_0234_),
    .Q_N(_2983_),
    .Q(\g.g_y[5].g_x[7].t.r_d ));
 sg13g2_dfrbp_1 \g.g_y[5].g_x[7].t.r_ghl$_SDFFE_PN0P_  (.CLK(clknet_leaf_9_clk),
    .RESET_B(net435),
    .D(_0235_),
    .Q_N(_2982_),
    .Q(\g.g_y[5].g_x[7].t.r_ghl ));
 sg13g2_dfrbp_1 \g.g_y[5].g_x[7].t.r_gnl$_SDFFE_PN0P_  (.CLK(clknet_leaf_8_clk),
    .RESET_B(net436),
    .D(_0236_),
    .Q_N(_2981_),
    .Q(\g.g_y[5].g_x[7].t.r_gnl ));
 sg13g2_dfrbp_1 \g.g_y[5].g_x[7].t.r_h$_SDFFE_PN0P_  (.CLK(clknet_leaf_8_clk),
    .RESET_B(net437),
    .D(_0237_),
    .Q_N(_2980_),
    .Q(\g.g_y[5].g_x[7].t.r_h ));
 sg13g2_dfrbp_1 \g.g_y[5].g_x[7].t.r_sc$_SDFFE_PN0P_  (.CLK(clknet_leaf_8_clk),
    .RESET_B(net438),
    .D(_0238_),
    .Q_N(_2979_),
    .Q(\g.g_y[5].g_x[7].t.out_sc ));
 sg13g2_dfrbp_1 \g.g_y[5].g_x[7].t.r_v$_SDFFE_PN0P_  (.CLK(clknet_leaf_8_clk),
    .RESET_B(net439),
    .D(_0239_),
    .Q_N(_2978_),
    .Q(\g.g_y[5].g_x[7].t.r_v ));
 sg13g2_dfrbp_1 \g.g_y[6].g_x[0].t.r_d$_SDFFE_PN0P_  (.CLK(clknet_leaf_9_clk),
    .RESET_B(net440),
    .D(_0240_),
    .Q_N(_2977_),
    .Q(\g.g_y[6].g_x[0].t.r_d ));
 sg13g2_dfrbp_1 \g.g_y[6].g_x[0].t.r_ghl$_SDFFE_PN0P_  (.CLK(clknet_leaf_10_clk),
    .RESET_B(net441),
    .D(_0241_),
    .Q_N(_2976_),
    .Q(\g.g_y[6].g_x[0].t.r_ghl ));
 sg13g2_dfrbp_1 \g.g_y[6].g_x[0].t.r_gnl$_SDFFE_PN0P_  (.CLK(clknet_leaf_10_clk),
    .RESET_B(net442),
    .D(_0242_),
    .Q_N(_2975_),
    .Q(\g.g_y[6].g_x[0].t.r_gnl ));
 sg13g2_dfrbp_1 \g.g_y[6].g_x[0].t.r_h$_SDFFE_PN0P_  (.CLK(clknet_leaf_10_clk),
    .RESET_B(net443),
    .D(_0243_),
    .Q_N(_2974_),
    .Q(\g.g_y[6].g_x[0].t.r_h ));
 sg13g2_dfrbp_1 \g.g_y[6].g_x[0].t.r_sc$_SDFFE_PN0P_  (.CLK(clknet_leaf_8_clk),
    .RESET_B(net444),
    .D(_0244_),
    .Q_N(_2973_),
    .Q(\g.g_y[6].g_x[0].t.out_sc ));
 sg13g2_dfrbp_1 \g.g_y[6].g_x[0].t.r_v$_SDFFE_PN0P_  (.CLK(clknet_leaf_10_clk),
    .RESET_B(net445),
    .D(_0245_),
    .Q_N(_2972_),
    .Q(\g.g_y[6].g_x[0].t.r_v ));
 sg13g2_dfrbp_1 \g.g_y[6].g_x[1].t.r_d$_SDFFE_PN0P_  (.CLK(clknet_leaf_9_clk),
    .RESET_B(net446),
    .D(_0246_),
    .Q_N(_2971_),
    .Q(\g.g_y[6].g_x[1].t.r_d ));
 sg13g2_dfrbp_1 \g.g_y[6].g_x[1].t.r_h$_SDFFE_PN0P_  (.CLK(clknet_leaf_9_clk),
    .RESET_B(net447),
    .D(_0247_),
    .Q_N(_2970_),
    .Q(\g.g_y[6].g_x[1].t.r_h ));
 sg13g2_dfrbp_1 \g.g_y[6].g_x[1].t.r_sc$_SDFFE_PN0P_  (.CLK(clknet_leaf_9_clk),
    .RESET_B(net448),
    .D(_0248_),
    .Q_N(_2969_),
    .Q(\g.g_y[6].g_x[1].t.out_sc ));
 sg13g2_dfrbp_1 \g.g_y[6].g_x[1].t.r_v$_SDFFE_PN0P_  (.CLK(clknet_leaf_9_clk),
    .RESET_B(net449),
    .D(_0249_),
    .Q_N(_2968_),
    .Q(\g.g_y[6].g_x[1].t.r_v ));
 sg13g2_dfrbp_1 \g.g_y[6].g_x[2].t.r_d$_SDFFE_PN0P_  (.CLK(clknet_leaf_9_clk),
    .RESET_B(net450),
    .D(_0250_),
    .Q_N(_2967_),
    .Q(\g.g_y[6].g_x[2].t.r_d ));
 sg13g2_dfrbp_1 \g.g_y[6].g_x[2].t.r_ghl$_SDFFE_PN0P_  (.CLK(clknet_leaf_9_clk),
    .RESET_B(net451),
    .D(_0251_),
    .Q_N(_2966_),
    .Q(\g.g_y[6].g_x[2].t.r_ghl ));
 sg13g2_dfrbp_1 \g.g_y[6].g_x[2].t.r_gnl$_SDFFE_PN0P_  (.CLK(clknet_leaf_8_clk),
    .RESET_B(net452),
    .D(_0252_),
    .Q_N(_2965_),
    .Q(\g.g_y[6].g_x[2].t.r_gnl ));
 sg13g2_dfrbp_1 \g.g_y[6].g_x[2].t.r_h$_SDFFE_PN0P_  (.CLK(clknet_leaf_7_clk),
    .RESET_B(net453),
    .D(_0253_),
    .Q_N(_2964_),
    .Q(\g.g_y[6].g_x[2].t.r_h ));
 sg13g2_dfrbp_1 \g.g_y[6].g_x[2].t.r_sc$_SDFFE_PN0P_  (.CLK(clknet_leaf_10_clk),
    .RESET_B(net454),
    .D(_0254_),
    .Q_N(_2963_),
    .Q(\g.g_y[6].g_x[2].t.out_sc ));
 sg13g2_dfrbp_1 \g.g_y[6].g_x[2].t.r_v$_SDFFE_PN0P_  (.CLK(clknet_leaf_7_clk),
    .RESET_B(net455),
    .D(_0255_),
    .Q_N(_2962_),
    .Q(\g.g_y[6].g_x[2].t.r_v ));
 sg13g2_dfrbp_1 \g.g_y[6].g_x[3].t.r_d$_SDFFE_PN0P_  (.CLK(clknet_leaf_7_clk),
    .RESET_B(net456),
    .D(_0256_),
    .Q_N(_2961_),
    .Q(\g.g_y[6].g_x[3].t.r_d ));
 sg13g2_dfrbp_1 \g.g_y[6].g_x[3].t.r_h$_SDFFE_PN0P_  (.CLK(clknet_leaf_7_clk),
    .RESET_B(net457),
    .D(_0257_),
    .Q_N(_2960_),
    .Q(\g.g_y[6].g_x[3].t.r_h ));
 sg13g2_dfrbp_1 \g.g_y[6].g_x[3].t.r_sc$_SDFFE_PN0P_  (.CLK(clknet_leaf_4_clk),
    .RESET_B(net458),
    .D(_0258_),
    .Q_N(_2959_),
    .Q(\g.g_y[6].g_x[3].t.out_sc ));
 sg13g2_dfrbp_1 \g.g_y[6].g_x[3].t.r_v$_SDFFE_PN0P_  (.CLK(clknet_leaf_7_clk),
    .RESET_B(net459),
    .D(_0259_),
    .Q_N(_2958_),
    .Q(\g.g_y[6].g_x[3].t.r_v ));
 sg13g2_dfrbp_1 \g.g_y[6].g_x[4].t.r_d$_SDFFE_PN0P_  (.CLK(clknet_leaf_5_clk),
    .RESET_B(net460),
    .D(_0260_),
    .Q_N(_2957_),
    .Q(\g.g_y[6].g_x[4].t.r_d ));
 sg13g2_dfrbp_1 \g.g_y[6].g_x[4].t.r_ghl$_SDFFE_PN0P_  (.CLK(clknet_leaf_4_clk),
    .RESET_B(net461),
    .D(_0261_),
    .Q_N(_2956_),
    .Q(\g.g_y[6].g_x[4].t.r_ghl ));
 sg13g2_dfrbp_1 \g.g_y[6].g_x[4].t.r_gnl$_SDFFE_PN0P_  (.CLK(clknet_leaf_4_clk),
    .RESET_B(net462),
    .D(_0262_),
    .Q_N(_2955_),
    .Q(\g.g_y[6].g_x[4].t.r_gnl ));
 sg13g2_dfrbp_1 \g.g_y[6].g_x[4].t.r_h$_SDFFE_PN0P_  (.CLK(clknet_leaf_5_clk),
    .RESET_B(net463),
    .D(_0263_),
    .Q_N(_2954_),
    .Q(\g.g_y[6].g_x[4].t.r_h ));
 sg13g2_dfrbp_1 \g.g_y[6].g_x[4].t.r_sc$_SDFFE_PN0P_  (.CLK(clknet_leaf_4_clk),
    .RESET_B(net464),
    .D(_0264_),
    .Q_N(_2953_),
    .Q(\g.g_y[6].g_x[4].t.out_sc ));
 sg13g2_dfrbp_1 \g.g_y[6].g_x[4].t.r_v$_SDFFE_PN0P_  (.CLK(clknet_leaf_5_clk),
    .RESET_B(net465),
    .D(_0265_),
    .Q_N(_2952_),
    .Q(\g.g_y[6].g_x[4].t.r_v ));
 sg13g2_dfrbp_1 \g.g_y[6].g_x[5].t.r_d$_SDFFE_PN0P_  (.CLK(clknet_leaf_4_clk),
    .RESET_B(net466),
    .D(_0266_),
    .Q_N(_2951_),
    .Q(\g.g_y[6].g_x[5].t.r_d ));
 sg13g2_dfrbp_1 \g.g_y[6].g_x[5].t.r_h$_SDFFE_PN0P_  (.CLK(clknet_leaf_12_clk),
    .RESET_B(net467),
    .D(_0267_),
    .Q_N(_2950_),
    .Q(\g.g_y[6].g_x[5].t.r_h ));
 sg13g2_dfrbp_1 \g.g_y[6].g_x[5].t.r_sc$_SDFFE_PN0P_  (.CLK(clknet_leaf_13_clk),
    .RESET_B(net468),
    .D(_0268_),
    .Q_N(_2949_),
    .Q(\g.g_y[6].g_x[5].t.out_sc ));
 sg13g2_dfrbp_1 \g.g_y[6].g_x[5].t.r_v$_SDFFE_PN0P_  (.CLK(clknet_leaf_12_clk),
    .RESET_B(net469),
    .D(_0269_),
    .Q_N(_2948_),
    .Q(\g.g_y[6].g_x[5].t.r_v ));
 sg13g2_dfrbp_1 \g.g_y[6].g_x[6].t.r_d$_SDFFE_PN0P_  (.CLK(clknet_leaf_13_clk),
    .RESET_B(net470),
    .D(_0270_),
    .Q_N(_2947_),
    .Q(\g.g_y[6].g_x[6].t.r_d ));
 sg13g2_dfrbp_1 \g.g_y[6].g_x[6].t.r_ghl$_SDFFE_PN0P_  (.CLK(clknet_leaf_13_clk),
    .RESET_B(net471),
    .D(_0271_),
    .Q_N(_2946_),
    .Q(\g.g_y[6].g_x[6].t.r_ghl ));
 sg13g2_dfrbp_1 \g.g_y[6].g_x[6].t.r_gnl$_SDFFE_PN0P_  (.CLK(clknet_leaf_12_clk),
    .RESET_B(net472),
    .D(_0272_),
    .Q_N(_2945_),
    .Q(\g.g_y[6].g_x[6].t.r_gnl ));
 sg13g2_dfrbp_1 \g.g_y[6].g_x[6].t.r_h$_SDFFE_PN0P_  (.CLK(clknet_leaf_12_clk),
    .RESET_B(net473),
    .D(_0273_),
    .Q_N(_2944_),
    .Q(\g.g_y[6].g_x[6].t.r_h ));
 sg13g2_dfrbp_1 \g.g_y[6].g_x[6].t.r_sc$_SDFFE_PN0P_  (.CLK(clknet_leaf_13_clk),
    .RESET_B(net474),
    .D(_0274_),
    .Q_N(_2943_),
    .Q(\g.g_y[6].g_x[6].t.out_sc ));
 sg13g2_dfrbp_1 \g.g_y[6].g_x[6].t.r_v$_SDFFE_PN0P_  (.CLK(clknet_leaf_12_clk),
    .RESET_B(net475),
    .D(_0275_),
    .Q_N(_2942_),
    .Q(\g.g_y[6].g_x[6].t.r_v ));
 sg13g2_dfrbp_1 \g.g_y[6].g_x[7].t.r_d$_SDFFE_PN0P_  (.CLK(clknet_leaf_10_clk),
    .RESET_B(net476),
    .D(_0276_),
    .Q_N(_2941_),
    .Q(\g.g_y[6].g_x[7].t.r_d ));
 sg13g2_dfrbp_1 \g.g_y[6].g_x[7].t.r_h$_SDFFE_PN0P_  (.CLK(clknet_leaf_12_clk),
    .RESET_B(net477),
    .D(_0277_),
    .Q_N(_2940_),
    .Q(\g.g_y[6].g_x[7].t.r_h ));
 sg13g2_dfrbp_1 \g.g_y[6].g_x[7].t.r_sc$_SDFFE_PN0P_  (.CLK(clknet_leaf_10_clk),
    .RESET_B(net478),
    .D(_0278_),
    .Q_N(_2939_),
    .Q(\g.g_y[6].g_x[7].t.out_sc ));
 sg13g2_dfrbp_1 \g.g_y[6].g_x[7].t.r_v$_SDFFE_PN0P_  (.CLK(clknet_leaf_11_clk),
    .RESET_B(net479),
    .D(_0279_),
    .Q_N(_2938_),
    .Q(\g.g_y[6].g_x[7].t.r_v ));
 sg13g2_dfrbp_1 \g.g_y[7].g_x[0].t.r_d$_SDFFE_PN0P_  (.CLK(clknet_leaf_16_clk),
    .RESET_B(net480),
    .D(_0280_),
    .Q_N(_2937_),
    .Q(\g.g_y[7].g_x[0].t.r_d ));
 sg13g2_dfrbp_1 \g.g_y[7].g_x[0].t.r_h$_SDFFE_PN0P_  (.CLK(clknet_leaf_11_clk),
    .RESET_B(net481),
    .D(_0281_),
    .Q_N(_2936_),
    .Q(\g.g_y[7].g_x[0].t.r_h ));
 sg13g2_dfrbp_1 \g.g_y[7].g_x[0].t.r_sc$_SDFFE_PN0P_  (.CLK(clknet_leaf_16_clk),
    .RESET_B(net482),
    .D(_0282_),
    .Q_N(_2935_),
    .Q(\g.g_y[7].g_x[0].t.out_sc ));
 sg13g2_dfrbp_1 \g.g_y[7].g_x[0].t.r_v$_SDFFE_PN0P_  (.CLK(clknet_leaf_11_clk),
    .RESET_B(net483),
    .D(_0283_),
    .Q_N(_2934_),
    .Q(\g.g_y[7].g_x[0].t.r_v ));
 sg13g2_dfrbp_1 \g.g_y[7].g_x[1].t.r_d$_SDFFE_PN0P_  (.CLK(clknet_leaf_11_clk),
    .RESET_B(net484),
    .D(_0284_),
    .Q_N(_2933_),
    .Q(\g.g_y[7].g_x[1].t.r_d ));
 sg13g2_dfrbp_1 \g.g_y[7].g_x[1].t.r_ghl$_SDFFE_PN0P_  (.CLK(clknet_leaf_11_clk),
    .RESET_B(net485),
    .D(_0285_),
    .Q_N(_2932_),
    .Q(\g.g_y[7].g_x[1].t.r_ghl ));
 sg13g2_dfrbp_1 \g.g_y[7].g_x[1].t.r_gnl$_SDFFE_PN0P_  (.CLK(clknet_leaf_11_clk),
    .RESET_B(net486),
    .D(_0286_),
    .Q_N(_2931_),
    .Q(\g.g_y[7].g_x[1].t.r_gnl ));
 sg13g2_dfrbp_1 \g.g_y[7].g_x[1].t.r_h$_SDFFE_PN0P_  (.CLK(clknet_leaf_11_clk),
    .RESET_B(net487),
    .D(_0287_),
    .Q_N(_2930_),
    .Q(\g.g_y[7].g_x[1].t.r_h ));
 sg13g2_dfrbp_1 \g.g_y[7].g_x[1].t.r_sc$_SDFFE_PN0P_  (.CLK(clknet_leaf_11_clk),
    .RESET_B(net488),
    .D(_0288_),
    .Q_N(_2929_),
    .Q(\g.g_y[7].g_x[1].t.out_sc ));
 sg13g2_dfrbp_1 \g.g_y[7].g_x[1].t.r_v$_SDFFE_PN0P_  (.CLK(clknet_leaf_10_clk),
    .RESET_B(net489),
    .D(_0289_),
    .Q_N(_2928_),
    .Q(\g.g_y[7].g_x[1].t.r_v ));
 sg13g2_dfrbp_1 \g.g_y[7].g_x[2].t.r_d$_SDFFE_PN0P_  (.CLK(clknet_leaf_15_clk),
    .RESET_B(net490),
    .D(_0290_),
    .Q_N(_2927_),
    .Q(\g.g_y[7].g_x[2].t.r_d ));
 sg13g2_dfrbp_1 \g.g_y[7].g_x[2].t.r_h$_SDFFE_PN0P_  (.CLK(clknet_leaf_12_clk),
    .RESET_B(net491),
    .D(_0291_),
    .Q_N(_2926_),
    .Q(\g.g_y[7].g_x[2].t.r_h ));
 sg13g2_dfrbp_1 \g.g_y[7].g_x[2].t.r_sc$_SDFFE_PN0P_  (.CLK(clknet_leaf_13_clk),
    .RESET_B(net492),
    .D(_0292_),
    .Q_N(_2925_),
    .Q(\g.g_y[7].g_x[2].t.out_sc ));
 sg13g2_dfrbp_1 \g.g_y[7].g_x[2].t.r_v$_SDFFE_PN0P_  (.CLK(clknet_leaf_12_clk),
    .RESET_B(net493),
    .D(_0293_),
    .Q_N(_2924_),
    .Q(\g.g_y[7].g_x[2].t.r_v ));
 sg13g2_dfrbp_1 \g.g_y[7].g_x[3].t.r_d$_SDFFE_PN0P_  (.CLK(clknet_leaf_3_clk),
    .RESET_B(net494),
    .D(_0294_),
    .Q_N(_2923_),
    .Q(\g.g_y[7].g_x[3].t.r_d ));
 sg13g2_dfrbp_1 \g.g_y[7].g_x[3].t.r_ghl$_SDFFE_PN0P_  (.CLK(clknet_leaf_4_clk),
    .RESET_B(net495),
    .D(_0295_),
    .Q_N(_2922_),
    .Q(\g.g_y[7].g_x[3].t.r_ghl ));
 sg13g2_dfrbp_1 \g.g_y[7].g_x[3].t.r_gnl$_SDFFE_PN0P_  (.CLK(clknet_leaf_13_clk),
    .RESET_B(net496),
    .D(_0296_),
    .Q_N(_2921_),
    .Q(\g.g_y[7].g_x[3].t.r_gnl ));
 sg13g2_dfrbp_1 \g.g_y[7].g_x[3].t.r_h$_SDFFE_PN0P_  (.CLK(clknet_leaf_13_clk),
    .RESET_B(net497),
    .D(_0297_),
    .Q_N(_2920_),
    .Q(\g.g_y[7].g_x[3].t.r_h ));
 sg13g2_dfrbp_1 \g.g_y[7].g_x[3].t.r_sc$_SDFFE_PN0P_  (.CLK(clknet_leaf_13_clk),
    .RESET_B(net498),
    .D(_0298_),
    .Q_N(_2919_),
    .Q(\g.g_y[7].g_x[3].t.out_sc ));
 sg13g2_dfrbp_1 \g.g_y[7].g_x[3].t.r_v$_SDFFE_PN0P_  (.CLK(clknet_leaf_14_clk),
    .RESET_B(net499),
    .D(_0299_),
    .Q_N(_2918_),
    .Q(\g.g_y[7].g_x[3].t.r_v ));
 sg13g2_dfrbp_1 \g.g_y[7].g_x[4].t.r_d$_SDFFE_PN0P_  (.CLK(clknet_leaf_24_clk),
    .RESET_B(net500),
    .D(_0300_),
    .Q_N(_2917_),
    .Q(\g.g_y[7].g_x[4].t.r_d ));
 sg13g2_dfrbp_1 \g.g_y[7].g_x[4].t.r_h$_SDFFE_PN0P_  (.CLK(clknet_leaf_24_clk),
    .RESET_B(net501),
    .D(_0301_),
    .Q_N(_2916_),
    .Q(\g.g_y[7].g_x[4].t.r_h ));
 sg13g2_dfrbp_1 \g.g_y[7].g_x[4].t.r_sc$_SDFFE_PN0P_  (.CLK(clknet_leaf_14_clk),
    .RESET_B(net502),
    .D(_0302_),
    .Q_N(_2915_),
    .Q(\g.g_y[7].g_x[4].t.out_sc ));
 sg13g2_dfrbp_1 \g.g_y[7].g_x[4].t.r_v$_SDFFE_PN0P_  (.CLK(clknet_leaf_23_clk),
    .RESET_B(net503),
    .D(_0303_),
    .Q_N(_2914_),
    .Q(\g.g_y[7].g_x[4].t.r_v ));
 sg13g2_dfrbp_1 \g.g_y[7].g_x[5].t.r_d$_SDFFE_PN0P_  (.CLK(clknet_leaf_14_clk),
    .RESET_B(net504),
    .D(_0304_),
    .Q_N(_2913_),
    .Q(\g.g_y[7].g_x[5].t.r_d ));
 sg13g2_dfrbp_1 \g.g_y[7].g_x[5].t.r_ghl$_SDFFE_PN0P_  (.CLK(clknet_leaf_14_clk),
    .RESET_B(net505),
    .D(_0305_),
    .Q_N(_2912_),
    .Q(\g.g_y[7].g_x[5].t.r_ghl ));
 sg13g2_dfrbp_1 \g.g_y[7].g_x[5].t.r_gnl$_SDFFE_PN0P_  (.CLK(clknet_leaf_14_clk),
    .RESET_B(net506),
    .D(_0306_),
    .Q_N(_2911_),
    .Q(\g.g_y[7].g_x[5].t.r_gnl ));
 sg13g2_dfrbp_1 \g.g_y[7].g_x[5].t.r_h$_SDFFE_PN0P_  (.CLK(clknet_leaf_14_clk),
    .RESET_B(net507),
    .D(_0307_),
    .Q_N(_2910_),
    .Q(\g.g_y[7].g_x[5].t.r_h ));
 sg13g2_dfrbp_1 \g.g_y[7].g_x[5].t.r_sc$_SDFFE_PN0P_  (.CLK(clknet_leaf_23_clk),
    .RESET_B(net508),
    .D(_0308_),
    .Q_N(_2909_),
    .Q(\g.g_y[7].g_x[5].t.out_sc ));
 sg13g2_dfrbp_1 \g.g_y[7].g_x[5].t.r_v$_SDFFE_PN0P_  (.CLK(clknet_leaf_14_clk),
    .RESET_B(net509),
    .D(_0309_),
    .Q_N(_2908_),
    .Q(\g.g_y[7].g_x[5].t.r_v ));
 sg13g2_dfrbp_1 \g.g_y[7].g_x[6].t.r_d$_SDFFE_PN0P_  (.CLK(clknet_leaf_15_clk),
    .RESET_B(net510),
    .D(_0310_),
    .Q_N(_2907_),
    .Q(\g.g_y[7].g_x[6].t.r_d ));
 sg13g2_dfrbp_1 \g.g_y[7].g_x[6].t.r_h$_SDFFE_PN0P_  (.CLK(clknet_leaf_15_clk),
    .RESET_B(net511),
    .D(_0311_),
    .Q_N(_2906_),
    .Q(\g.g_y[7].g_x[6].t.r_h ));
 sg13g2_dfrbp_1 \g.g_y[7].g_x[6].t.r_sc$_SDFFE_PN0P_  (.CLK(clknet_leaf_15_clk),
    .RESET_B(net512),
    .D(_0312_),
    .Q_N(_2905_),
    .Q(\g.g_y[7].g_x[6].t.out_sc ));
 sg13g2_dfrbp_1 \g.g_y[7].g_x[6].t.r_v$_SDFFE_PN0P_  (.CLK(clknet_leaf_15_clk),
    .RESET_B(net513),
    .D(_0313_),
    .Q_N(_2904_),
    .Q(\g.g_y[7].g_x[6].t.r_v ));
 sg13g2_dfrbp_1 \g.g_y[7].g_x[7].t.r_d$_SDFFE_PN0P_  (.CLK(clknet_leaf_16_clk),
    .RESET_B(net514),
    .D(_0314_),
    .Q_N(_2903_),
    .Q(\g.g_y[7].g_x[7].t.r_d ));
 sg13g2_dfrbp_1 \g.g_y[7].g_x[7].t.r_ghl$_SDFFE_PN0P_  (.CLK(clknet_leaf_16_clk),
    .RESET_B(net515),
    .D(_0315_),
    .Q_N(_2902_),
    .Q(\g.g_y[7].g_x[7].t.r_ghl ));
 sg13g2_dfrbp_1 \g.g_y[7].g_x[7].t.r_gnl$_SDFFE_PN0P_  (.CLK(clknet_leaf_16_clk),
    .RESET_B(net516),
    .D(_0316_),
    .Q_N(_2901_),
    .Q(\g.g_y[7].g_x[7].t.r_gnl ));
 sg13g2_dfrbp_1 \g.g_y[7].g_x[7].t.r_h$_SDFFE_PN0P_  (.CLK(clknet_leaf_15_clk),
    .RESET_B(net517),
    .D(_0317_),
    .Q_N(_2900_),
    .Q(\g.g_y[7].g_x[7].t.r_h ));
 sg13g2_dfrbp_1 \g.g_y[7].g_x[7].t.r_sc$_SDFFE_PN0P_  (.CLK(clknet_leaf_16_clk),
    .RESET_B(net518),
    .D(_0318_),
    .Q_N(_2899_),
    .Q(\g.g_y[7].g_x[7].t.out_sc ));
 sg13g2_dfrbp_1 \g.g_y[7].g_x[7].t.r_v$_SDFFE_PN0P_  (.CLK(clknet_leaf_15_clk),
    .RESET_B(net519),
    .D(_0319_),
    .Q_N(_2898_),
    .Q(\g.g_y[7].g_x[7].t.r_v ));
 sg13g2_buf_1 input1 (.A(ui_in[0]),
    .X(net1));
 sg13g2_buf_1 input2 (.A(ui_in[1]),
    .X(net2));
 sg13g2_buf_1 input3 (.A(ui_in[2]),
    .X(net3));
 sg13g2_buf_1 input4 (.A(ui_in[3]),
    .X(net4));
 sg13g2_buf_1 input5 (.A(ui_in[4]),
    .X(net5));
 sg13g2_buf_1 input6 (.A(ui_in[5]),
    .X(net6));
 sg13g2_buf_1 input7 (.A(ui_in[6]),
    .X(net7));
 sg13g2_buf_1 input8 (.A(ui_in[7]),
    .X(net8));
 sg13g2_buf_1 input9 (.A(uio_in[1]),
    .X(net9));
 sg13g2_buf_1 input10 (.A(uio_in[2]),
    .X(net10));
 sg13g2_buf_1 input11 (.A(uio_in[3]),
    .X(net11));
 sg13g2_buf_1 input12 (.A(uio_in[4]),
    .X(net12));
 sg13g2_buf_1 output13 (.A(net13),
    .X(uio_out[7]));
 sg13g2_buf_1 output14 (.A(net14),
    .X(uo_out[0]));
 sg13g2_buf_1 output15 (.A(net15),
    .X(uo_out[1]));
 sg13g2_buf_1 output16 (.A(net16),
    .X(uo_out[2]));
 sg13g2_buf_1 output17 (.A(net17),
    .X(uo_out[3]));
 sg13g2_buf_1 output18 (.A(net18),
    .X(uo_out[4]));
 sg13g2_buf_1 output19 (.A(net19),
    .X(uo_out[5]));
 sg13g2_buf_1 output20 (.A(net20),
    .X(uo_out[6]));
 sg13g2_buf_1 output21 (.A(net21),
    .X(uo_out[7]));
 sg13g2_buf_2 fanout22 (.A(_0608_),
    .X(net22));
 sg13g2_buf_2 fanout23 (.A(_2231_),
    .X(net23));
 sg13g2_buf_2 fanout24 (.A(_2065_),
    .X(net24));
 sg13g2_buf_4 fanout25 (.X(net25),
    .A(_1935_));
 sg13g2_buf_2 fanout26 (.A(_1844_),
    .X(net26));
 sg13g2_buf_2 fanout27 (.A(_1747_),
    .X(net27));
 sg13g2_buf_2 fanout28 (.A(_1394_),
    .X(net28));
 sg13g2_buf_4 fanout29 (.X(net29),
    .A(_1326_));
 sg13g2_buf_2 fanout30 (.A(_1308_),
    .X(net30));
 sg13g2_buf_2 fanout31 (.A(_1289_),
    .X(net31));
 sg13g2_buf_2 fanout32 (.A(_0910_),
    .X(net32));
 sg13g2_buf_4 fanout33 (.X(net33),
    .A(_0907_));
 sg13g2_buf_2 fanout34 (.A(_0889_),
    .X(net34));
 sg13g2_buf_2 fanout35 (.A(_0807_),
    .X(net35));
 sg13g2_buf_2 fanout36 (.A(_0805_),
    .X(net36));
 sg13g2_buf_2 fanout37 (.A(_0717_),
    .X(net37));
 sg13g2_buf_2 fanout38 (.A(_0702_),
    .X(net38));
 sg13g2_buf_2 fanout39 (.A(_0648_),
    .X(net39));
 sg13g2_buf_2 fanout40 (.A(_0624_),
    .X(net40));
 sg13g2_buf_2 fanout41 (.A(_0609_),
    .X(net41));
 sg13g2_buf_4 fanout42 (.X(net42),
    .A(_0607_));
 sg13g2_buf_2 fanout43 (.A(_2729_),
    .X(net43));
 sg13g2_buf_2 fanout44 (.A(_2702_),
    .X(net44));
 sg13g2_buf_2 fanout45 (.A(_2689_),
    .X(net45));
 sg13g2_buf_2 fanout46 (.A(_2599_),
    .X(net46));
 sg13g2_buf_4 fanout47 (.X(net47),
    .A(_2593_));
 sg13g2_buf_2 fanout48 (.A(_1757_),
    .X(net48));
 sg13g2_buf_2 fanout49 (.A(_1632_),
    .X(net49));
 sg13g2_buf_2 fanout50 (.A(_1565_),
    .X(net50));
 sg13g2_buf_2 fanout51 (.A(_1471_),
    .X(net51));
 sg13g2_buf_2 fanout52 (.A(_1296_),
    .X(net52));
 sg13g2_buf_2 fanout53 (.A(_1053_),
    .X(net53));
 sg13g2_buf_2 fanout54 (.A(_0818_),
    .X(net54));
 sg13g2_buf_2 fanout55 (.A(_0815_),
    .X(net55));
 sg13g2_buf_2 fanout56 (.A(_0729_),
    .X(net56));
 sg13g2_buf_2 fanout57 (.A(_0647_),
    .X(net57));
 sg13g2_buf_2 fanout58 (.A(_0476_),
    .X(net58));
 sg13g2_buf_2 fanout59 (.A(_2873_),
    .X(net59));
 sg13g2_buf_2 fanout60 (.A(_2754_),
    .X(net60));
 sg13g2_buf_2 fanout61 (.A(_2728_),
    .X(net61));
 sg13g2_buf_2 fanout62 (.A(_2723_),
    .X(net62));
 sg13g2_buf_2 fanout63 (.A(_2720_),
    .X(net63));
 sg13g2_buf_2 fanout64 (.A(_2716_),
    .X(net64));
 sg13g2_buf_2 fanout65 (.A(_2705_),
    .X(net65));
 sg13g2_buf_2 fanout66 (.A(_2701_),
    .X(net66));
 sg13g2_buf_2 fanout67 (.A(_2485_),
    .X(net67));
 sg13g2_buf_2 fanout68 (.A(_2442_),
    .X(net68));
 sg13g2_buf_2 fanout69 (.A(_2372_),
    .X(net69));
 sg13g2_buf_2 fanout70 (.A(_2314_),
    .X(net70));
 sg13g2_buf_2 fanout71 (.A(_2233_),
    .X(net71));
 sg13g2_buf_2 fanout72 (.A(_2226_),
    .X(net72));
 sg13g2_buf_2 fanout73 (.A(_2138_),
    .X(net73));
 sg13g2_buf_2 fanout74 (.A(_2063_),
    .X(net74));
 sg13g2_buf_2 fanout75 (.A(_1997_),
    .X(net75));
 sg13g2_buf_2 fanout76 (.A(_1933_),
    .X(net76));
 sg13g2_buf_2 fanout77 (.A(_1859_),
    .X(net77));
 sg13g2_buf_2 fanout78 (.A(_1846_),
    .X(net78));
 sg13g2_buf_2 fanout79 (.A(_1690_),
    .X(net79));
 sg13g2_buf_2 fanout80 (.A(_1562_),
    .X(net80));
 sg13g2_buf_2 fanout81 (.A(_1478_),
    .X(net81));
 sg13g2_buf_2 fanout82 (.A(_1393_),
    .X(net82));
 sg13g2_buf_2 fanout83 (.A(_1310_),
    .X(net83));
 sg13g2_buf_2 fanout84 (.A(_1213_),
    .X(net84));
 sg13g2_buf_2 fanout85 (.A(_0968_),
    .X(net85));
 sg13g2_buf_2 fanout86 (.A(_0891_),
    .X(net86));
 sg13g2_buf_2 fanout87 (.A(_0822_),
    .X(net87));
 sg13g2_buf_2 fanout88 (.A(_0812_),
    .X(net88));
 sg13g2_buf_2 fanout89 (.A(_0809_),
    .X(net89));
 sg13g2_buf_2 fanout90 (.A(_0643_),
    .X(net90));
 sg13g2_buf_2 fanout91 (.A(_2894_),
    .X(net91));
 sg13g2_buf_2 fanout92 (.A(_2890_),
    .X(net92));
 sg13g2_buf_2 fanout93 (.A(_2889_),
    .X(net93));
 sg13g2_buf_2 fanout94 (.A(_2738_),
    .X(net94));
 sg13g2_buf_2 fanout95 (.A(_2732_),
    .X(net95));
 sg13g2_buf_2 fanout96 (.A(_2722_),
    .X(net96));
 sg13g2_buf_2 fanout97 (.A(_2711_),
    .X(net97));
 sg13g2_buf_2 fanout98 (.A(_2707_),
    .X(net98));
 sg13g2_buf_2 fanout99 (.A(_2704_),
    .X(net99));
 sg13g2_buf_2 fanout100 (.A(_2243_),
    .X(net100));
 sg13g2_buf_2 fanout101 (.A(_2067_),
    .X(net101));
 sg13g2_buf_2 fanout102 (.A(_1767_),
    .X(net102));
 sg13g2_buf_2 fanout103 (.A(_1749_),
    .X(net103));
 sg13g2_buf_2 fanout104 (.A(_1720_),
    .X(net104));
 sg13g2_buf_2 fanout105 (.A(_1652_),
    .X(net105));
 sg13g2_buf_2 fanout106 (.A(_1448_),
    .X(net106));
 sg13g2_buf_2 fanout107 (.A(_1301_),
    .X(net107));
 sg13g2_buf_2 fanout108 (.A(_1291_),
    .X(net108));
 sg13g2_buf_2 fanout109 (.A(_1049_),
    .X(net109));
 sg13g2_buf_2 fanout110 (.A(_1037_),
    .X(net110));
 sg13g2_buf_2 fanout111 (.A(_0996_),
    .X(net111));
 sg13g2_buf_2 fanout112 (.A(_0906_),
    .X(net112));
 sg13g2_buf_2 fanout113 (.A(_0777_),
    .X(net113));
 sg13g2_buf_2 fanout114 (.A(_0694_),
    .X(net114));
 sg13g2_buf_2 fanout115 (.A(_0631_),
    .X(net115));
 sg13g2_buf_2 fanout116 (.A(_0614_),
    .X(net116));
 sg13g2_buf_2 fanout117 (.A(_0466_),
    .X(net117));
 sg13g2_buf_2 fanout118 (.A(_0439_),
    .X(net118));
 sg13g2_buf_2 fanout119 (.A(_0387_),
    .X(net119));
 sg13g2_buf_2 fanout120 (.A(_2896_),
    .X(net120));
 sg13g2_buf_2 fanout121 (.A(_2891_),
    .X(net121));
 sg13g2_buf_2 fanout122 (.A(_2857_),
    .X(net122));
 sg13g2_buf_2 fanout123 (.A(_2745_),
    .X(net123));
 sg13g2_buf_2 fanout124 (.A(_2743_),
    .X(net124));
 sg13g2_buf_2 fanout125 (.A(_2740_),
    .X(net125));
 sg13g2_buf_2 fanout126 (.A(_2737_),
    .X(net126));
 sg13g2_buf_2 fanout127 (.A(_2731_),
    .X(net127));
 sg13g2_buf_2 fanout128 (.A(_2710_),
    .X(net128));
 sg13g2_buf_2 fanout129 (.A(_2706_),
    .X(net129));
 sg13g2_buf_2 fanout130 (.A(_2639_),
    .X(net130));
 sg13g2_buf_2 fanout131 (.A(_2583_),
    .X(net131));
 sg13g2_buf_2 fanout132 (.A(_2179_),
    .X(net132));
 sg13g2_buf_2 fanout133 (.A(_2105_),
    .X(net133));
 sg13g2_buf_2 fanout134 (.A(_2101_),
    .X(net134));
 sg13g2_buf_2 fanout135 (.A(_1969_),
    .X(net135));
 sg13g2_buf_2 fanout136 (.A(_1956_),
    .X(net136));
 sg13g2_buf_2 fanout137 (.A(_1824_),
    .X(net137));
 sg13g2_buf_2 fanout138 (.A(_1797_),
    .X(net138));
 sg13g2_buf_2 fanout139 (.A(_1783_),
    .X(net139));
 sg13g2_buf_2 fanout140 (.A(_1596_),
    .X(net140));
 sg13g2_buf_2 fanout141 (.A(_1490_),
    .X(net141));
 sg13g2_buf_2 fanout142 (.A(_1488_),
    .X(net142));
 sg13g2_buf_2 fanout143 (.A(_1368_),
    .X(net143));
 sg13g2_buf_2 fanout144 (.A(_1361_),
    .X(net144));
 sg13g2_buf_2 fanout145 (.A(_1346_),
    .X(net145));
 sg13g2_buf_2 fanout146 (.A(_1246_),
    .X(net146));
 sg13g2_buf_2 fanout147 (.A(_1180_),
    .X(net147));
 sg13g2_buf_2 fanout148 (.A(_1127_),
    .X(net148));
 sg13g2_buf_2 fanout149 (.A(_1078_),
    .X(net149));
 sg13g2_buf_2 fanout150 (.A(_1029_),
    .X(net150));
 sg13g2_buf_2 fanout151 (.A(_0990_),
    .X(net151));
 sg13g2_buf_2 fanout152 (.A(_0934_),
    .X(net152));
 sg13g2_buf_2 fanout153 (.A(_0925_),
    .X(net153));
 sg13g2_buf_2 fanout154 (.A(_0923_),
    .X(net154));
 sg13g2_buf_2 fanout155 (.A(_0862_),
    .X(net155));
 sg13g2_buf_2 fanout156 (.A(_0846_),
    .X(net156));
 sg13g2_buf_2 fanout157 (.A(_0845_),
    .X(net157));
 sg13g2_buf_2 fanout158 (.A(_0843_),
    .X(net158));
 sg13g2_buf_2 fanout159 (.A(_0749_),
    .X(net159));
 sg13g2_buf_2 fanout160 (.A(_0726_),
    .X(net160));
 sg13g2_buf_2 fanout161 (.A(_0679_),
    .X(net161));
 sg13g2_buf_2 fanout162 (.A(_0542_),
    .X(net162));
 sg13g2_buf_2 fanout163 (.A(_0529_),
    .X(net163));
 sg13g2_buf_2 fanout164 (.A(_0528_),
    .X(net164));
 sg13g2_buf_2 fanout165 (.A(_0509_),
    .X(net165));
 sg13g2_buf_2 fanout166 (.A(_0385_),
    .X(net166));
 sg13g2_buf_2 fanout167 (.A(_0361_),
    .X(net167));
 sg13g2_buf_2 fanout168 (.A(_0359_),
    .X(net168));
 sg13g2_buf_2 fanout169 (.A(_0324_),
    .X(net169));
 sg13g2_buf_2 fanout170 (.A(_2895_),
    .X(net170));
 sg13g2_buf_2 fanout171 (.A(_2862_),
    .X(net171));
 sg13g2_buf_2 fanout172 (.A(_2822_),
    .X(net172));
 sg13g2_buf_2 fanout173 (.A(_2807_),
    .X(net173));
 sg13g2_buf_2 fanout174 (.A(_2781_),
    .X(net174));
 sg13g2_buf_2 fanout175 (.A(_2739_),
    .X(net175));
 sg13g2_buf_2 fanout176 (.A(_2696_),
    .X(net176));
 sg13g2_buf_2 fanout177 (.A(_2690_),
    .X(net177));
 sg13g2_buf_2 fanout178 (.A(_2647_),
    .X(net178));
 sg13g2_buf_2 fanout179 (.A(_2601_),
    .X(net179));
 sg13g2_buf_2 fanout180 (.A(_2600_),
    .X(net180));
 sg13g2_buf_2 fanout181 (.A(_2582_),
    .X(net181));
 sg13g2_buf_2 fanout182 (.A(_2587_),
    .X(net182));
 sg13g2_buf_2 fanout183 (.A(_2586_),
    .X(net183));
 sg13g2_buf_2 fanout184 (.A(_2581_),
    .X(net184));
 sg13g2_tielo _6128__185 (.L_LO(net185));
 sg13g2_tielo _6129__186 (.L_LO(net186));
 sg13g2_tielo _6130__187 (.L_LO(net187));
 sg13g2_tielo _6131__188 (.L_LO(net188));
 sg13g2_tielo _6132__189 (.L_LO(net189));
 sg13g2_tielo _6133__190 (.L_LO(net190));
 sg13g2_tielo _6134__191 (.L_LO(net191));
 sg13g2_tielo _6136__192 (.L_LO(net192));
 sg13g2_tielo _6137__193 (.L_LO(net193));
 sg13g2_tielo _6138__194 (.L_LO(net194));
 sg13g2_tielo _6139__195 (.L_LO(net195));
 sg13g2_tielo _6140__196 (.L_LO(net196));
 sg13g2_tielo _6141__197 (.L_LO(net197));
 sg13g2_tielo _6142__198 (.L_LO(net198));
 sg13g2_tiehi \g.g_y[0].g_x[0].t.r_d$_SDFFE_PN0P__200  (.L_HI(net200));
 sg13g2_tiehi \g.g_y[0].g_x[0].t.r_ghl$_SDFFE_PN0P__201  (.L_HI(net201));
 sg13g2_tiehi \g.g_y[0].g_x[0].t.r_gnl$_SDFFE_PN0P__202  (.L_HI(net202));
 sg13g2_tiehi \g.g_y[0].g_x[0].t.r_h$_SDFFE_PN0P__203  (.L_HI(net203));
 sg13g2_tiehi \g.g_y[0].g_x[0].t.r_sc$_SDFFE_PN0P__204  (.L_HI(net204));
 sg13g2_tiehi \g.g_y[0].g_x[0].t.r_v$_SDFFE_PN0P__205  (.L_HI(net205));
 sg13g2_tiehi \g.g_y[0].g_x[1].t.r_d$_SDFFE_PN0P__206  (.L_HI(net206));
 sg13g2_tiehi \g.g_y[0].g_x[1].t.r_h$_SDFFE_PN0P__207  (.L_HI(net207));
 sg13g2_tiehi \g.g_y[0].g_x[1].t.r_sc$_SDFFE_PN0P__208  (.L_HI(net208));
 sg13g2_tiehi \g.g_y[0].g_x[1].t.r_v$_SDFFE_PN0P__209  (.L_HI(net209));
 sg13g2_tiehi \g.g_y[0].g_x[2].t.r_d$_SDFFE_PN0P__210  (.L_HI(net210));
 sg13g2_tiehi \g.g_y[0].g_x[2].t.r_ghl$_SDFFE_PN0P__211  (.L_HI(net211));
 sg13g2_tiehi \g.g_y[0].g_x[2].t.r_gnl$_SDFFE_PN0P__212  (.L_HI(net212));
 sg13g2_tiehi \g.g_y[0].g_x[2].t.r_h$_SDFFE_PN0P__213  (.L_HI(net213));
 sg13g2_tiehi \g.g_y[0].g_x[2].t.r_sc$_SDFFE_PN0P__214  (.L_HI(net214));
 sg13g2_tiehi \g.g_y[0].g_x[2].t.r_v$_SDFFE_PN0P__215  (.L_HI(net215));
 sg13g2_tiehi \g.g_y[0].g_x[3].t.r_d$_SDFFE_PN0P__216  (.L_HI(net216));
 sg13g2_tiehi \g.g_y[0].g_x[3].t.r_h$_SDFFE_PN0P__217  (.L_HI(net217));
 sg13g2_tiehi \g.g_y[0].g_x[3].t.r_sc$_SDFFE_PN0P__218  (.L_HI(net218));
 sg13g2_tiehi \g.g_y[0].g_x[3].t.r_v$_SDFFE_PN0P__219  (.L_HI(net219));
 sg13g2_tiehi \g.g_y[0].g_x[4].t.r_d$_SDFFE_PN0P__220  (.L_HI(net220));
 sg13g2_tiehi \g.g_y[0].g_x[4].t.r_ghl$_SDFFE_PN0P__221  (.L_HI(net221));
 sg13g2_tiehi \g.g_y[0].g_x[4].t.r_gnl$_SDFFE_PN0P__222  (.L_HI(net222));
 sg13g2_tiehi \g.g_y[0].g_x[4].t.r_h$_SDFFE_PN0P__223  (.L_HI(net223));
 sg13g2_tiehi \g.g_y[0].g_x[4].t.r_sc$_SDFFE_PN0P__224  (.L_HI(net224));
 sg13g2_tiehi \g.g_y[0].g_x[4].t.r_v$_SDFFE_PN0P__225  (.L_HI(net225));
 sg13g2_tiehi \g.g_y[0].g_x[5].t.r_d$_SDFFE_PN0P__226  (.L_HI(net226));
 sg13g2_tiehi \g.g_y[0].g_x[5].t.r_h$_SDFFE_PN0P__227  (.L_HI(net227));
 sg13g2_tiehi \g.g_y[0].g_x[5].t.r_sc$_SDFFE_PN0P__228  (.L_HI(net228));
 sg13g2_tiehi \g.g_y[0].g_x[5].t.r_v$_SDFFE_PN0P__229  (.L_HI(net229));
 sg13g2_tiehi \g.g_y[0].g_x[6].t.r_d$_SDFFE_PN0P__230  (.L_HI(net230));
 sg13g2_tiehi \g.g_y[0].g_x[6].t.r_ghl$_SDFFE_PN0P__231  (.L_HI(net231));
 sg13g2_tiehi \g.g_y[0].g_x[6].t.r_gnl$_SDFFE_PN0P__232  (.L_HI(net232));
 sg13g2_tiehi \g.g_y[0].g_x[6].t.r_h$_SDFFE_PN0P__233  (.L_HI(net233));
 sg13g2_tiehi \g.g_y[0].g_x[6].t.r_sc$_SDFFE_PN0P__234  (.L_HI(net234));
 sg13g2_tiehi \g.g_y[0].g_x[6].t.r_v$_SDFFE_PN0P__235  (.L_HI(net235));
 sg13g2_tiehi \g.g_y[0].g_x[7].t.r_d$_SDFFE_PN0P__236  (.L_HI(net236));
 sg13g2_tiehi \g.g_y[0].g_x[7].t.r_h$_SDFFE_PN0P__237  (.L_HI(net237));
 sg13g2_tiehi \g.g_y[0].g_x[7].t.r_sc$_SDFFE_PN0P__238  (.L_HI(net238));
 sg13g2_tiehi \g.g_y[0].g_x[7].t.r_v$_SDFFE_PN0P__239  (.L_HI(net239));
 sg13g2_tiehi \g.g_y[1].g_x[0].t.r_d$_SDFFE_PN0P__240  (.L_HI(net240));
 sg13g2_tiehi \g.g_y[1].g_x[0].t.r_h$_SDFFE_PN0P__241  (.L_HI(net241));
 sg13g2_tiehi \g.g_y[1].g_x[0].t.r_sc$_SDFFE_PN0P__242  (.L_HI(net242));
 sg13g2_tiehi \g.g_y[1].g_x[0].t.r_v$_SDFFE_PN0P__243  (.L_HI(net243));
 sg13g2_tiehi \g.g_y[1].g_x[1].t.r_d$_SDFFE_PN0P__244  (.L_HI(net244));
 sg13g2_tiehi \g.g_y[1].g_x[1].t.r_ghl$_SDFFE_PN0P__245  (.L_HI(net245));
 sg13g2_tiehi \g.g_y[1].g_x[1].t.r_gnl$_SDFFE_PN0P__246  (.L_HI(net246));
 sg13g2_tiehi \g.g_y[1].g_x[1].t.r_h$_SDFFE_PN0P__247  (.L_HI(net247));
 sg13g2_tiehi \g.g_y[1].g_x[1].t.r_sc$_SDFFE_PN0P__248  (.L_HI(net248));
 sg13g2_tiehi \g.g_y[1].g_x[1].t.r_v$_SDFFE_PN0P__249  (.L_HI(net249));
 sg13g2_tiehi \g.g_y[1].g_x[2].t.r_d$_SDFFE_PN0P__250  (.L_HI(net250));
 sg13g2_tiehi \g.g_y[1].g_x[2].t.r_h$_SDFFE_PN0P__251  (.L_HI(net251));
 sg13g2_tiehi \g.g_y[1].g_x[2].t.r_sc$_SDFFE_PN0P__252  (.L_HI(net252));
 sg13g2_tiehi \g.g_y[1].g_x[2].t.r_v$_SDFFE_PN0P__253  (.L_HI(net253));
 sg13g2_tiehi \g.g_y[1].g_x[3].t.r_d$_SDFFE_PN0P__254  (.L_HI(net254));
 sg13g2_tiehi \g.g_y[1].g_x[3].t.r_ghl$_SDFFE_PN0P__255  (.L_HI(net255));
 sg13g2_tiehi \g.g_y[1].g_x[3].t.r_gnl$_SDFFE_PN0P__256  (.L_HI(net256));
 sg13g2_tiehi \g.g_y[1].g_x[3].t.r_h$_SDFFE_PN0P__257  (.L_HI(net257));
 sg13g2_tiehi \g.g_y[1].g_x[3].t.r_sc$_SDFFE_PN0P__258  (.L_HI(net258));
 sg13g2_tiehi \g.g_y[1].g_x[3].t.r_v$_SDFFE_PN0P__259  (.L_HI(net259));
 sg13g2_tiehi \g.g_y[1].g_x[4].t.r_d$_SDFFE_PN0P__260  (.L_HI(net260));
 sg13g2_tiehi \g.g_y[1].g_x[4].t.r_h$_SDFFE_PN0P__261  (.L_HI(net261));
 sg13g2_tiehi \g.g_y[1].g_x[4].t.r_sc$_SDFFE_PN0P__262  (.L_HI(net262));
 sg13g2_tiehi \g.g_y[1].g_x[4].t.r_v$_SDFFE_PN0P__263  (.L_HI(net263));
 sg13g2_tiehi \g.g_y[1].g_x[5].t.r_d$_SDFFE_PN0P__264  (.L_HI(net264));
 sg13g2_tiehi \g.g_y[1].g_x[5].t.r_ghl$_SDFFE_PN0P__265  (.L_HI(net265));
 sg13g2_tiehi \g.g_y[1].g_x[5].t.r_gnl$_SDFFE_PN0P__266  (.L_HI(net266));
 sg13g2_tiehi \g.g_y[1].g_x[5].t.r_h$_SDFFE_PN0P__267  (.L_HI(net267));
 sg13g2_tiehi \g.g_y[1].g_x[5].t.r_sc$_SDFFE_PN0P__268  (.L_HI(net268));
 sg13g2_tiehi \g.g_y[1].g_x[5].t.r_v$_SDFFE_PN0P__269  (.L_HI(net269));
 sg13g2_tiehi \g.g_y[1].g_x[6].t.r_d$_SDFFE_PN0P__270  (.L_HI(net270));
 sg13g2_tiehi \g.g_y[1].g_x[6].t.r_h$_SDFFE_PN0P__271  (.L_HI(net271));
 sg13g2_tiehi \g.g_y[1].g_x[6].t.r_sc$_SDFFE_PN0P__272  (.L_HI(net272));
 sg13g2_tiehi \g.g_y[1].g_x[6].t.r_v$_SDFFE_PN0P__273  (.L_HI(net273));
 sg13g2_tiehi \g.g_y[1].g_x[7].t.r_d$_SDFFE_PN0P__274  (.L_HI(net274));
 sg13g2_tiehi \g.g_y[1].g_x[7].t.r_ghl$_SDFFE_PN0P__275  (.L_HI(net275));
 sg13g2_tiehi \g.g_y[1].g_x[7].t.r_gnl$_SDFFE_PN0P__276  (.L_HI(net276));
 sg13g2_tiehi \g.g_y[1].g_x[7].t.r_h$_SDFFE_PN0P__277  (.L_HI(net277));
 sg13g2_tiehi \g.g_y[1].g_x[7].t.r_sc$_SDFFE_PN0P__278  (.L_HI(net278));
 sg13g2_tiehi \g.g_y[1].g_x[7].t.r_v$_SDFFE_PN0P__279  (.L_HI(net279));
 sg13g2_tiehi \g.g_y[2].g_x[0].t.r_d$_SDFFE_PN0P__280  (.L_HI(net280));
 sg13g2_tiehi \g.g_y[2].g_x[0].t.r_ghl$_SDFFE_PN0P__281  (.L_HI(net281));
 sg13g2_tiehi \g.g_y[2].g_x[0].t.r_gnl$_SDFFE_PN0P__282  (.L_HI(net282));
 sg13g2_tiehi \g.g_y[2].g_x[0].t.r_h$_SDFFE_PN0P__283  (.L_HI(net283));
 sg13g2_tiehi \g.g_y[2].g_x[0].t.r_sc$_SDFFE_PN0P__284  (.L_HI(net284));
 sg13g2_tiehi \g.g_y[2].g_x[0].t.r_v$_SDFFE_PN0P__285  (.L_HI(net285));
 sg13g2_tiehi \g.g_y[2].g_x[1].t.r_d$_SDFFE_PN0P__286  (.L_HI(net286));
 sg13g2_tiehi \g.g_y[2].g_x[1].t.r_h$_SDFFE_PN0P__287  (.L_HI(net287));
 sg13g2_tiehi \g.g_y[2].g_x[1].t.r_sc$_SDFFE_PN0P__288  (.L_HI(net288));
 sg13g2_tiehi \g.g_y[2].g_x[1].t.r_v$_SDFFE_PN0P__289  (.L_HI(net289));
 sg13g2_tiehi \g.g_y[2].g_x[2].t.r_d$_SDFFE_PN0P__290  (.L_HI(net290));
 sg13g2_tiehi \g.g_y[2].g_x[2].t.r_ghl$_SDFFE_PN0P__291  (.L_HI(net291));
 sg13g2_tiehi \g.g_y[2].g_x[2].t.r_gnl$_SDFFE_PN0P__292  (.L_HI(net292));
 sg13g2_tiehi \g.g_y[2].g_x[2].t.r_h$_SDFFE_PN0P__293  (.L_HI(net293));
 sg13g2_tiehi \g.g_y[2].g_x[2].t.r_sc$_SDFFE_PN0P__294  (.L_HI(net294));
 sg13g2_tiehi \g.g_y[2].g_x[2].t.r_v$_SDFFE_PN0P__295  (.L_HI(net295));
 sg13g2_tiehi \g.g_y[2].g_x[3].t.r_d$_SDFFE_PN0P__296  (.L_HI(net296));
 sg13g2_tiehi \g.g_y[2].g_x[3].t.r_h$_SDFFE_PN0P__297  (.L_HI(net297));
 sg13g2_tiehi \g.g_y[2].g_x[3].t.r_sc$_SDFFE_PN0P__298  (.L_HI(net298));
 sg13g2_tiehi \g.g_y[2].g_x[3].t.r_v$_SDFFE_PN0P__299  (.L_HI(net299));
 sg13g2_tiehi \g.g_y[2].g_x[4].t.r_d$_SDFFE_PN0P__300  (.L_HI(net300));
 sg13g2_tiehi \g.g_y[2].g_x[4].t.r_ghl$_SDFFE_PN0P__301  (.L_HI(net301));
 sg13g2_tiehi \g.g_y[2].g_x[4].t.r_gnl$_SDFFE_PN0P__302  (.L_HI(net302));
 sg13g2_tiehi \g.g_y[2].g_x[4].t.r_h$_SDFFE_PN0P__303  (.L_HI(net303));
 sg13g2_tiehi \g.g_y[2].g_x[4].t.r_sc$_SDFFE_PN0P__304  (.L_HI(net304));
 sg13g2_tiehi \g.g_y[2].g_x[4].t.r_v$_SDFFE_PN0P__305  (.L_HI(net305));
 sg13g2_tiehi \g.g_y[2].g_x[5].t.r_d$_SDFFE_PN0P__306  (.L_HI(net306));
 sg13g2_tiehi \g.g_y[2].g_x[5].t.r_h$_SDFFE_PN0P__307  (.L_HI(net307));
 sg13g2_tiehi \g.g_y[2].g_x[5].t.r_sc$_SDFFE_PN0P__308  (.L_HI(net308));
 sg13g2_tiehi \g.g_y[2].g_x[5].t.r_v$_SDFFE_PN0P__309  (.L_HI(net309));
 sg13g2_tiehi \g.g_y[2].g_x[6].t.r_d$_SDFFE_PN0P__310  (.L_HI(net310));
 sg13g2_tiehi \g.g_y[2].g_x[6].t.r_ghl$_SDFFE_PN0P__311  (.L_HI(net311));
 sg13g2_tiehi \g.g_y[2].g_x[6].t.r_gnl$_SDFFE_PN0P__312  (.L_HI(net312));
 sg13g2_tiehi \g.g_y[2].g_x[6].t.r_h$_SDFFE_PN0P__313  (.L_HI(net313));
 sg13g2_tiehi \g.g_y[2].g_x[6].t.r_sc$_SDFFE_PN0P__314  (.L_HI(net314));
 sg13g2_tiehi \g.g_y[2].g_x[6].t.r_v$_SDFFE_PN0P__315  (.L_HI(net315));
 sg13g2_tiehi \g.g_y[2].g_x[7].t.r_d$_SDFFE_PN0P__316  (.L_HI(net316));
 sg13g2_tiehi \g.g_y[2].g_x[7].t.r_h$_SDFFE_PN0P__317  (.L_HI(net317));
 sg13g2_tiehi \g.g_y[2].g_x[7].t.r_sc$_SDFFE_PN0P__318  (.L_HI(net318));
 sg13g2_tiehi \g.g_y[2].g_x[7].t.r_v$_SDFFE_PN0P__319  (.L_HI(net319));
 sg13g2_tiehi \g.g_y[3].g_x[0].t.r_d$_SDFFE_PN0P__320  (.L_HI(net320));
 sg13g2_tiehi \g.g_y[3].g_x[0].t.r_h$_SDFFE_PN0P__321  (.L_HI(net321));
 sg13g2_tiehi \g.g_y[3].g_x[0].t.r_sc$_SDFFE_PN0P__322  (.L_HI(net322));
 sg13g2_tiehi \g.g_y[3].g_x[0].t.r_v$_SDFFE_PN0P__323  (.L_HI(net323));
 sg13g2_tiehi \g.g_y[3].g_x[1].t.r_d$_SDFFE_PN0P__324  (.L_HI(net324));
 sg13g2_tiehi \g.g_y[3].g_x[1].t.r_ghl$_SDFFE_PN0P__325  (.L_HI(net325));
 sg13g2_tiehi \g.g_y[3].g_x[1].t.r_gnl$_SDFFE_PN0P__326  (.L_HI(net326));
 sg13g2_tiehi \g.g_y[3].g_x[1].t.r_h$_SDFFE_PN0P__327  (.L_HI(net327));
 sg13g2_tiehi \g.g_y[3].g_x[1].t.r_sc$_SDFFE_PN0P__328  (.L_HI(net328));
 sg13g2_tiehi \g.g_y[3].g_x[1].t.r_v$_SDFFE_PN0P__329  (.L_HI(net329));
 sg13g2_tiehi \g.g_y[3].g_x[2].t.r_d$_SDFFE_PN0P__330  (.L_HI(net330));
 sg13g2_tiehi \g.g_y[3].g_x[2].t.r_h$_SDFFE_PN0P__331  (.L_HI(net331));
 sg13g2_tiehi \g.g_y[3].g_x[2].t.r_sc$_SDFFE_PN0P__332  (.L_HI(net332));
 sg13g2_tiehi \g.g_y[3].g_x[2].t.r_v$_SDFFE_PN0P__333  (.L_HI(net333));
 sg13g2_tiehi \g.g_y[3].g_x[3].t.r_d$_SDFFE_PN0P__334  (.L_HI(net334));
 sg13g2_tiehi \g.g_y[3].g_x[3].t.r_ghl$_SDFFE_PN0P__335  (.L_HI(net335));
 sg13g2_tiehi \g.g_y[3].g_x[3].t.r_gnl$_SDFFE_PN0P__336  (.L_HI(net336));
 sg13g2_tiehi \g.g_y[3].g_x[3].t.r_h$_SDFFE_PN0P__337  (.L_HI(net337));
 sg13g2_tiehi \g.g_y[3].g_x[3].t.r_sc$_SDFFE_PN0P__338  (.L_HI(net338));
 sg13g2_tiehi \g.g_y[3].g_x[3].t.r_v$_SDFFE_PN0P__339  (.L_HI(net339));
 sg13g2_tiehi \g.g_y[3].g_x[4].t.r_d$_SDFFE_PN0P__340  (.L_HI(net340));
 sg13g2_tiehi \g.g_y[3].g_x[4].t.r_h$_SDFFE_PN0P__341  (.L_HI(net341));
 sg13g2_tiehi \g.g_y[3].g_x[4].t.r_sc$_SDFFE_PN0P__342  (.L_HI(net342));
 sg13g2_tiehi \g.g_y[3].g_x[4].t.r_v$_SDFFE_PN0P__343  (.L_HI(net343));
 sg13g2_tiehi \g.g_y[3].g_x[5].t.r_d$_SDFFE_PN0P__344  (.L_HI(net344));
 sg13g2_tiehi \g.g_y[3].g_x[5].t.r_ghl$_SDFFE_PN0P__345  (.L_HI(net345));
 sg13g2_tiehi \g.g_y[3].g_x[5].t.r_gnl$_SDFFE_PN0P__346  (.L_HI(net346));
 sg13g2_tiehi \g.g_y[3].g_x[5].t.r_h$_SDFFE_PN0P__347  (.L_HI(net347));
 sg13g2_tiehi \g.g_y[3].g_x[5].t.r_sc$_SDFFE_PN0P__348  (.L_HI(net348));
 sg13g2_tiehi \g.g_y[3].g_x[5].t.r_v$_SDFFE_PN0P__349  (.L_HI(net349));
 sg13g2_tiehi \g.g_y[3].g_x[6].t.r_d$_SDFFE_PN0P__350  (.L_HI(net350));
 sg13g2_tiehi \g.g_y[3].g_x[6].t.r_h$_SDFFE_PN0P__351  (.L_HI(net351));
 sg13g2_tiehi \g.g_y[3].g_x[6].t.r_sc$_SDFFE_PN0P__352  (.L_HI(net352));
 sg13g2_tiehi \g.g_y[3].g_x[6].t.r_v$_SDFFE_PN0P__353  (.L_HI(net353));
 sg13g2_tiehi \g.g_y[3].g_x[7].t.r_d$_SDFFE_PN0P__354  (.L_HI(net354));
 sg13g2_tiehi \g.g_y[3].g_x[7].t.r_ghl$_SDFFE_PN0P__355  (.L_HI(net355));
 sg13g2_tiehi \g.g_y[3].g_x[7].t.r_gnl$_SDFFE_PN0P__356  (.L_HI(net356));
 sg13g2_tiehi \g.g_y[3].g_x[7].t.r_h$_SDFFE_PN0P__357  (.L_HI(net357));
 sg13g2_tiehi \g.g_y[3].g_x[7].t.r_sc$_SDFFE_PN0P__358  (.L_HI(net358));
 sg13g2_tiehi \g.g_y[3].g_x[7].t.r_v$_SDFFE_PN0P__359  (.L_HI(net359));
 sg13g2_tiehi \g.g_y[4].g_x[0].t.r_d$_SDFFE_PN0P__360  (.L_HI(net360));
 sg13g2_tiehi \g.g_y[4].g_x[0].t.r_ghl$_SDFFE_PN0P__361  (.L_HI(net361));
 sg13g2_tiehi \g.g_y[4].g_x[0].t.r_gnl$_SDFFE_PN0P__362  (.L_HI(net362));
 sg13g2_tiehi \g.g_y[4].g_x[0].t.r_h$_SDFFE_PN0P__363  (.L_HI(net363));
 sg13g2_tiehi \g.g_y[4].g_x[0].t.r_sc$_SDFFE_PN0P__364  (.L_HI(net364));
 sg13g2_tiehi \g.g_y[4].g_x[0].t.r_v$_SDFFE_PN0P__365  (.L_HI(net365));
 sg13g2_tiehi \g.g_y[4].g_x[1].t.r_d$_SDFFE_PN0P__366  (.L_HI(net366));
 sg13g2_tiehi \g.g_y[4].g_x[1].t.r_h$_SDFFE_PN0P__367  (.L_HI(net367));
 sg13g2_tiehi \g.g_y[4].g_x[1].t.r_sc$_SDFFE_PN0P__368  (.L_HI(net368));
 sg13g2_tiehi \g.g_y[4].g_x[1].t.r_v$_SDFFE_PN0P__369  (.L_HI(net369));
 sg13g2_tiehi \g.g_y[4].g_x[2].t.r_d$_SDFFE_PN0P__370  (.L_HI(net370));
 sg13g2_tiehi \g.g_y[4].g_x[2].t.r_ghl$_SDFFE_PN0P__371  (.L_HI(net371));
 sg13g2_tiehi \g.g_y[4].g_x[2].t.r_gnl$_SDFFE_PN0P__372  (.L_HI(net372));
 sg13g2_tiehi \g.g_y[4].g_x[2].t.r_h$_SDFFE_PN0P__373  (.L_HI(net373));
 sg13g2_tiehi \g.g_y[4].g_x[2].t.r_sc$_SDFFE_PN0P__374  (.L_HI(net374));
 sg13g2_tiehi \g.g_y[4].g_x[2].t.r_v$_SDFFE_PN0P__375  (.L_HI(net375));
 sg13g2_tiehi \g.g_y[4].g_x[3].t.r_d$_SDFFE_PN0P__376  (.L_HI(net376));
 sg13g2_tiehi \g.g_y[4].g_x[3].t.r_h$_SDFFE_PN0P__377  (.L_HI(net377));
 sg13g2_tiehi \g.g_y[4].g_x[3].t.r_sc$_SDFFE_PN0P__378  (.L_HI(net378));
 sg13g2_tiehi \g.g_y[4].g_x[3].t.r_v$_SDFFE_PN0P__379  (.L_HI(net379));
 sg13g2_tiehi \g.g_y[4].g_x[4].t.r_d$_SDFFE_PN0P__380  (.L_HI(net380));
 sg13g2_tiehi \g.g_y[4].g_x[4].t.r_ghl$_SDFFE_PN0P__381  (.L_HI(net381));
 sg13g2_tiehi \g.g_y[4].g_x[4].t.r_gnl$_SDFFE_PN0P__382  (.L_HI(net382));
 sg13g2_tiehi \g.g_y[4].g_x[4].t.r_h$_SDFFE_PN0P__383  (.L_HI(net383));
 sg13g2_tiehi \g.g_y[4].g_x[4].t.r_sc$_SDFFE_PN0P__384  (.L_HI(net384));
 sg13g2_tiehi \g.g_y[4].g_x[4].t.r_v$_SDFFE_PN0P__385  (.L_HI(net385));
 sg13g2_tiehi \g.g_y[4].g_x[5].t.r_d$_SDFFE_PN0P__386  (.L_HI(net386));
 sg13g2_tiehi \g.g_y[4].g_x[5].t.r_h$_SDFFE_PN0P__387  (.L_HI(net387));
 sg13g2_tiehi \g.g_y[4].g_x[5].t.r_sc$_SDFFE_PN0P__388  (.L_HI(net388));
 sg13g2_tiehi \g.g_y[4].g_x[5].t.r_v$_SDFFE_PN0P__389  (.L_HI(net389));
 sg13g2_tiehi \g.g_y[4].g_x[6].t.r_d$_SDFFE_PN0P__390  (.L_HI(net390));
 sg13g2_tiehi \g.g_y[4].g_x[6].t.r_ghl$_SDFFE_PN0P__391  (.L_HI(net391));
 sg13g2_tiehi \g.g_y[4].g_x[6].t.r_gnl$_SDFFE_PN0P__392  (.L_HI(net392));
 sg13g2_tiehi \g.g_y[4].g_x[6].t.r_h$_SDFFE_PN0P__393  (.L_HI(net393));
 sg13g2_tiehi \g.g_y[4].g_x[6].t.r_sc$_SDFFE_PN0P__394  (.L_HI(net394));
 sg13g2_tiehi \g.g_y[4].g_x[6].t.r_v$_SDFFE_PN0P__395  (.L_HI(net395));
 sg13g2_tiehi \g.g_y[4].g_x[7].t.r_d$_SDFFE_PN0P__396  (.L_HI(net396));
 sg13g2_tiehi \g.g_y[4].g_x[7].t.r_h$_SDFFE_PN0P__397  (.L_HI(net397));
 sg13g2_tiehi \g.g_y[4].g_x[7].t.r_sc$_SDFFE_PN0P__398  (.L_HI(net398));
 sg13g2_tiehi \g.g_y[4].g_x[7].t.r_v$_SDFFE_PN0P__399  (.L_HI(net399));
 sg13g2_tiehi \g.g_y[5].g_x[0].t.r_d$_SDFFE_PN0P__400  (.L_HI(net400));
 sg13g2_tiehi \g.g_y[5].g_x[0].t.r_h$_SDFFE_PN0P__401  (.L_HI(net401));
 sg13g2_tiehi \g.g_y[5].g_x[0].t.r_sc$_SDFFE_PN0P__402  (.L_HI(net402));
 sg13g2_tiehi \g.g_y[5].g_x[0].t.r_v$_SDFFE_PN0P__403  (.L_HI(net403));
 sg13g2_tiehi \g.g_y[5].g_x[1].t.r_d$_SDFFE_PN0P__404  (.L_HI(net404));
 sg13g2_tiehi \g.g_y[5].g_x[1].t.r_ghl$_SDFFE_PN0P__405  (.L_HI(net405));
 sg13g2_tiehi \g.g_y[5].g_x[1].t.r_gnl$_SDFFE_PN0P__406  (.L_HI(net406));
 sg13g2_tiehi \g.g_y[5].g_x[1].t.r_h$_SDFFE_PN0P__407  (.L_HI(net407));
 sg13g2_tiehi \g.g_y[5].g_x[1].t.r_sc$_SDFFE_PN0P__408  (.L_HI(net408));
 sg13g2_tiehi \g.g_y[5].g_x[1].t.r_v$_SDFFE_PN0P__409  (.L_HI(net409));
 sg13g2_tiehi \g.g_y[5].g_x[2].t.r_d$_SDFFE_PN0P__410  (.L_HI(net410));
 sg13g2_tiehi \g.g_y[5].g_x[2].t.r_h$_SDFFE_PN0P__411  (.L_HI(net411));
 sg13g2_tiehi \g.g_y[5].g_x[2].t.r_sc$_SDFFE_PN0P__412  (.L_HI(net412));
 sg13g2_tiehi \g.g_y[5].g_x[2].t.r_v$_SDFFE_PN0P__413  (.L_HI(net413));
 sg13g2_tiehi \g.g_y[5].g_x[3].t.r_d$_SDFFE_PN0P__414  (.L_HI(net414));
 sg13g2_tiehi \g.g_y[5].g_x[3].t.r_ghl$_SDFFE_PN0P__415  (.L_HI(net415));
 sg13g2_tiehi \g.g_y[5].g_x[3].t.r_gnl$_SDFFE_PN0P__416  (.L_HI(net416));
 sg13g2_tiehi \g.g_y[5].g_x[3].t.r_h$_SDFFE_PN0P__417  (.L_HI(net417));
 sg13g2_tiehi \g.g_y[5].g_x[3].t.r_sc$_SDFFE_PN0P__418  (.L_HI(net418));
 sg13g2_tiehi \g.g_y[5].g_x[3].t.r_v$_SDFFE_PN0P__419  (.L_HI(net419));
 sg13g2_tiehi \g.g_y[5].g_x[4].t.r_d$_SDFFE_PN0P__420  (.L_HI(net420));
 sg13g2_tiehi \g.g_y[5].g_x[4].t.r_h$_SDFFE_PN0P__421  (.L_HI(net421));
 sg13g2_tiehi \g.g_y[5].g_x[4].t.r_sc$_SDFFE_PN0P__422  (.L_HI(net422));
 sg13g2_tiehi \g.g_y[5].g_x[4].t.r_v$_SDFFE_PN0P__423  (.L_HI(net423));
 sg13g2_tiehi \g.g_y[5].g_x[5].t.r_d$_SDFFE_PN0P__424  (.L_HI(net424));
 sg13g2_tiehi \g.g_y[5].g_x[5].t.r_ghl$_SDFFE_PN0P__425  (.L_HI(net425));
 sg13g2_tiehi \g.g_y[5].g_x[5].t.r_gnl$_SDFFE_PN0P__426  (.L_HI(net426));
 sg13g2_tiehi \g.g_y[5].g_x[5].t.r_h$_SDFFE_PN0P__427  (.L_HI(net427));
 sg13g2_tiehi \g.g_y[5].g_x[5].t.r_sc$_SDFFE_PN0P__428  (.L_HI(net428));
 sg13g2_tiehi \g.g_y[5].g_x[5].t.r_v$_SDFFE_PN0P__429  (.L_HI(net429));
 sg13g2_tiehi \g.g_y[5].g_x[6].t.r_d$_SDFFE_PN0P__430  (.L_HI(net430));
 sg13g2_tiehi \g.g_y[5].g_x[6].t.r_h$_SDFFE_PN0P__431  (.L_HI(net431));
 sg13g2_tiehi \g.g_y[5].g_x[6].t.r_sc$_SDFFE_PN0P__432  (.L_HI(net432));
 sg13g2_tiehi \g.g_y[5].g_x[6].t.r_v$_SDFFE_PN0P__433  (.L_HI(net433));
 sg13g2_tiehi \g.g_y[5].g_x[7].t.r_d$_SDFFE_PN0P__434  (.L_HI(net434));
 sg13g2_tiehi \g.g_y[5].g_x[7].t.r_ghl$_SDFFE_PN0P__435  (.L_HI(net435));
 sg13g2_tiehi \g.g_y[5].g_x[7].t.r_gnl$_SDFFE_PN0P__436  (.L_HI(net436));
 sg13g2_tiehi \g.g_y[5].g_x[7].t.r_h$_SDFFE_PN0P__437  (.L_HI(net437));
 sg13g2_tiehi \g.g_y[5].g_x[7].t.r_sc$_SDFFE_PN0P__438  (.L_HI(net438));
 sg13g2_tiehi \g.g_y[5].g_x[7].t.r_v$_SDFFE_PN0P__439  (.L_HI(net439));
 sg13g2_tiehi \g.g_y[6].g_x[0].t.r_d$_SDFFE_PN0P__440  (.L_HI(net440));
 sg13g2_tiehi \g.g_y[6].g_x[0].t.r_ghl$_SDFFE_PN0P__441  (.L_HI(net441));
 sg13g2_tiehi \g.g_y[6].g_x[0].t.r_gnl$_SDFFE_PN0P__442  (.L_HI(net442));
 sg13g2_tiehi \g.g_y[6].g_x[0].t.r_h$_SDFFE_PN0P__443  (.L_HI(net443));
 sg13g2_tiehi \g.g_y[6].g_x[0].t.r_sc$_SDFFE_PN0P__444  (.L_HI(net444));
 sg13g2_tiehi \g.g_y[6].g_x[0].t.r_v$_SDFFE_PN0P__445  (.L_HI(net445));
 sg13g2_tiehi \g.g_y[6].g_x[1].t.r_d$_SDFFE_PN0P__446  (.L_HI(net446));
 sg13g2_tiehi \g.g_y[6].g_x[1].t.r_h$_SDFFE_PN0P__447  (.L_HI(net447));
 sg13g2_tiehi \g.g_y[6].g_x[1].t.r_sc$_SDFFE_PN0P__448  (.L_HI(net448));
 sg13g2_tiehi \g.g_y[6].g_x[1].t.r_v$_SDFFE_PN0P__449  (.L_HI(net449));
 sg13g2_tiehi \g.g_y[6].g_x[2].t.r_d$_SDFFE_PN0P__450  (.L_HI(net450));
 sg13g2_tiehi \g.g_y[6].g_x[2].t.r_ghl$_SDFFE_PN0P__451  (.L_HI(net451));
 sg13g2_tiehi \g.g_y[6].g_x[2].t.r_gnl$_SDFFE_PN0P__452  (.L_HI(net452));
 sg13g2_tiehi \g.g_y[6].g_x[2].t.r_h$_SDFFE_PN0P__453  (.L_HI(net453));
 sg13g2_tiehi \g.g_y[6].g_x[2].t.r_sc$_SDFFE_PN0P__454  (.L_HI(net454));
 sg13g2_tiehi \g.g_y[6].g_x[2].t.r_v$_SDFFE_PN0P__455  (.L_HI(net455));
 sg13g2_tiehi \g.g_y[6].g_x[3].t.r_d$_SDFFE_PN0P__456  (.L_HI(net456));
 sg13g2_tiehi \g.g_y[6].g_x[3].t.r_h$_SDFFE_PN0P__457  (.L_HI(net457));
 sg13g2_tiehi \g.g_y[6].g_x[3].t.r_sc$_SDFFE_PN0P__458  (.L_HI(net458));
 sg13g2_tiehi \g.g_y[6].g_x[3].t.r_v$_SDFFE_PN0P__459  (.L_HI(net459));
 sg13g2_tiehi \g.g_y[6].g_x[4].t.r_d$_SDFFE_PN0P__460  (.L_HI(net460));
 sg13g2_tiehi \g.g_y[6].g_x[4].t.r_ghl$_SDFFE_PN0P__461  (.L_HI(net461));
 sg13g2_tiehi \g.g_y[6].g_x[4].t.r_gnl$_SDFFE_PN0P__462  (.L_HI(net462));
 sg13g2_tiehi \g.g_y[6].g_x[4].t.r_h$_SDFFE_PN0P__463  (.L_HI(net463));
 sg13g2_tiehi \g.g_y[6].g_x[4].t.r_sc$_SDFFE_PN0P__464  (.L_HI(net464));
 sg13g2_tiehi \g.g_y[6].g_x[4].t.r_v$_SDFFE_PN0P__465  (.L_HI(net465));
 sg13g2_tiehi \g.g_y[6].g_x[5].t.r_d$_SDFFE_PN0P__466  (.L_HI(net466));
 sg13g2_tiehi \g.g_y[6].g_x[5].t.r_h$_SDFFE_PN0P__467  (.L_HI(net467));
 sg13g2_tiehi \g.g_y[6].g_x[5].t.r_sc$_SDFFE_PN0P__468  (.L_HI(net468));
 sg13g2_tiehi \g.g_y[6].g_x[5].t.r_v$_SDFFE_PN0P__469  (.L_HI(net469));
 sg13g2_tiehi \g.g_y[6].g_x[6].t.r_d$_SDFFE_PN0P__470  (.L_HI(net470));
 sg13g2_tiehi \g.g_y[6].g_x[6].t.r_ghl$_SDFFE_PN0P__471  (.L_HI(net471));
 sg13g2_tiehi \g.g_y[6].g_x[6].t.r_gnl$_SDFFE_PN0P__472  (.L_HI(net472));
 sg13g2_tiehi \g.g_y[6].g_x[6].t.r_h$_SDFFE_PN0P__473  (.L_HI(net473));
 sg13g2_tiehi \g.g_y[6].g_x[6].t.r_sc$_SDFFE_PN0P__474  (.L_HI(net474));
 sg13g2_tiehi \g.g_y[6].g_x[6].t.r_v$_SDFFE_PN0P__475  (.L_HI(net475));
 sg13g2_tiehi \g.g_y[6].g_x[7].t.r_d$_SDFFE_PN0P__476  (.L_HI(net476));
 sg13g2_tiehi \g.g_y[6].g_x[7].t.r_h$_SDFFE_PN0P__477  (.L_HI(net477));
 sg13g2_tiehi \g.g_y[6].g_x[7].t.r_sc$_SDFFE_PN0P__478  (.L_HI(net478));
 sg13g2_tiehi \g.g_y[6].g_x[7].t.r_v$_SDFFE_PN0P__479  (.L_HI(net479));
 sg13g2_tiehi \g.g_y[7].g_x[0].t.r_d$_SDFFE_PN0P__480  (.L_HI(net480));
 sg13g2_tiehi \g.g_y[7].g_x[0].t.r_h$_SDFFE_PN0P__481  (.L_HI(net481));
 sg13g2_tiehi \g.g_y[7].g_x[0].t.r_sc$_SDFFE_PN0P__482  (.L_HI(net482));
 sg13g2_tiehi \g.g_y[7].g_x[0].t.r_v$_SDFFE_PN0P__483  (.L_HI(net483));
 sg13g2_tiehi \g.g_y[7].g_x[1].t.r_d$_SDFFE_PN0P__484  (.L_HI(net484));
 sg13g2_tiehi \g.g_y[7].g_x[1].t.r_ghl$_SDFFE_PN0P__485  (.L_HI(net485));
 sg13g2_tiehi \g.g_y[7].g_x[1].t.r_gnl$_SDFFE_PN0P__486  (.L_HI(net486));
 sg13g2_tiehi \g.g_y[7].g_x[1].t.r_h$_SDFFE_PN0P__487  (.L_HI(net487));
 sg13g2_tiehi \g.g_y[7].g_x[1].t.r_sc$_SDFFE_PN0P__488  (.L_HI(net488));
 sg13g2_tiehi \g.g_y[7].g_x[1].t.r_v$_SDFFE_PN0P__489  (.L_HI(net489));
 sg13g2_tiehi \g.g_y[7].g_x[2].t.r_d$_SDFFE_PN0P__490  (.L_HI(net490));
 sg13g2_tiehi \g.g_y[7].g_x[2].t.r_h$_SDFFE_PN0P__491  (.L_HI(net491));
 sg13g2_tiehi \g.g_y[7].g_x[2].t.r_sc$_SDFFE_PN0P__492  (.L_HI(net492));
 sg13g2_tiehi \g.g_y[7].g_x[2].t.r_v$_SDFFE_PN0P__493  (.L_HI(net493));
 sg13g2_tiehi \g.g_y[7].g_x[3].t.r_d$_SDFFE_PN0P__494  (.L_HI(net494));
 sg13g2_tiehi \g.g_y[7].g_x[3].t.r_ghl$_SDFFE_PN0P__495  (.L_HI(net495));
 sg13g2_tiehi \g.g_y[7].g_x[3].t.r_gnl$_SDFFE_PN0P__496  (.L_HI(net496));
 sg13g2_tiehi \g.g_y[7].g_x[3].t.r_h$_SDFFE_PN0P__497  (.L_HI(net497));
 sg13g2_tiehi \g.g_y[7].g_x[3].t.r_sc$_SDFFE_PN0P__498  (.L_HI(net498));
 sg13g2_tiehi \g.g_y[7].g_x[3].t.r_v$_SDFFE_PN0P__499  (.L_HI(net499));
 sg13g2_tiehi \g.g_y[7].g_x[4].t.r_d$_SDFFE_PN0P__500  (.L_HI(net500));
 sg13g2_tiehi \g.g_y[7].g_x[4].t.r_h$_SDFFE_PN0P__501  (.L_HI(net501));
 sg13g2_tiehi \g.g_y[7].g_x[4].t.r_sc$_SDFFE_PN0P__502  (.L_HI(net502));
 sg13g2_tiehi \g.g_y[7].g_x[4].t.r_v$_SDFFE_PN0P__503  (.L_HI(net503));
 sg13g2_tiehi \g.g_y[7].g_x[5].t.r_d$_SDFFE_PN0P__504  (.L_HI(net504));
 sg13g2_tiehi \g.g_y[7].g_x[5].t.r_ghl$_SDFFE_PN0P__505  (.L_HI(net505));
 sg13g2_tiehi \g.g_y[7].g_x[5].t.r_gnl$_SDFFE_PN0P__506  (.L_HI(net506));
 sg13g2_tiehi \g.g_y[7].g_x[5].t.r_h$_SDFFE_PN0P__507  (.L_HI(net507));
 sg13g2_tiehi \g.g_y[7].g_x[5].t.r_sc$_SDFFE_PN0P__508  (.L_HI(net508));
 sg13g2_tiehi \g.g_y[7].g_x[5].t.r_v$_SDFFE_PN0P__509  (.L_HI(net509));
 sg13g2_tiehi \g.g_y[7].g_x[6].t.r_d$_SDFFE_PN0P__510  (.L_HI(net510));
 sg13g2_tiehi \g.g_y[7].g_x[6].t.r_h$_SDFFE_PN0P__511  (.L_HI(net511));
 sg13g2_tiehi \g.g_y[7].g_x[6].t.r_sc$_SDFFE_PN0P__512  (.L_HI(net512));
 sg13g2_tiehi \g.g_y[7].g_x[6].t.r_v$_SDFFE_PN0P__513  (.L_HI(net513));
 sg13g2_tiehi \g.g_y[7].g_x[7].t.r_d$_SDFFE_PN0P__514  (.L_HI(net514));
 sg13g2_tiehi \g.g_y[7].g_x[7].t.r_ghl$_SDFFE_PN0P__515  (.L_HI(net515));
 sg13g2_tiehi \g.g_y[7].g_x[7].t.r_gnl$_SDFFE_PN0P__516  (.L_HI(net516));
 sg13g2_tiehi \g.g_y[7].g_x[7].t.r_h$_SDFFE_PN0P__517  (.L_HI(net517));
 sg13g2_tiehi \g.g_y[7].g_x[7].t.r_sc$_SDFFE_PN0P__518  (.L_HI(net518));
 sg13g2_tiehi \g.g_y[7].g_x[7].t.r_v$_SDFFE_PN0P__519  (.L_HI(net519));
 sg13g2_buf_2 clkbuf_leaf_1_clk (.A(clknet_3_1__leaf_clk),
    .X(clknet_leaf_1_clk));
 sg13g2_buf_2 clkbuf_leaf_2_clk (.A(clknet_3_1__leaf_clk),
    .X(clknet_leaf_2_clk));
 sg13g2_buf_2 clkbuf_leaf_3_clk (.A(clknet_3_1__leaf_clk),
    .X(clknet_leaf_3_clk));
 sg13g2_buf_2 clkbuf_leaf_4_clk (.A(clknet_3_4__leaf_clk),
    .X(clknet_leaf_4_clk));
 sg13g2_buf_2 clkbuf_leaf_5_clk (.A(clknet_3_4__leaf_clk),
    .X(clknet_leaf_5_clk));
 sg13g2_buf_2 clkbuf_leaf_6_clk (.A(clknet_3_4__leaf_clk),
    .X(clknet_leaf_6_clk));
 sg13g2_buf_2 clkbuf_leaf_7_clk (.A(clknet_3_4__leaf_clk),
    .X(clknet_leaf_7_clk));
 sg13g2_buf_2 clkbuf_leaf_8_clk (.A(clknet_3_5__leaf_clk),
    .X(clknet_leaf_8_clk));
 sg13g2_buf_2 clkbuf_leaf_9_clk (.A(clknet_3_5__leaf_clk),
    .X(clknet_leaf_9_clk));
 sg13g2_buf_2 clkbuf_leaf_10_clk (.A(clknet_3_5__leaf_clk),
    .X(clknet_leaf_10_clk));
 sg13g2_buf_2 clkbuf_leaf_11_clk (.A(clknet_3_5__leaf_clk),
    .X(clknet_leaf_11_clk));
 sg13g2_buf_2 clkbuf_leaf_12_clk (.A(clknet_3_5__leaf_clk),
    .X(clknet_leaf_12_clk));
 sg13g2_buf_2 clkbuf_leaf_13_clk (.A(clknet_3_4__leaf_clk),
    .X(clknet_leaf_13_clk));
 sg13g2_buf_2 clkbuf_leaf_14_clk (.A(clknet_3_6__leaf_clk),
    .X(clknet_leaf_14_clk));
 sg13g2_buf_2 clkbuf_leaf_15_clk (.A(clknet_3_7__leaf_clk),
    .X(clknet_leaf_15_clk));
 sg13g2_buf_2 clkbuf_leaf_16_clk (.A(clknet_3_7__leaf_clk),
    .X(clknet_leaf_16_clk));
 sg13g2_buf_2 clkbuf_leaf_17_clk (.A(clknet_3_7__leaf_clk),
    .X(clknet_leaf_17_clk));
 sg13g2_buf_2 clkbuf_leaf_18_clk (.A(clknet_3_7__leaf_clk),
    .X(clknet_leaf_18_clk));
 sg13g2_buf_2 clkbuf_leaf_19_clk (.A(clknet_3_7__leaf_clk),
    .X(clknet_leaf_19_clk));
 sg13g2_buf_2 clkbuf_leaf_20_clk (.A(clknet_3_6__leaf_clk),
    .X(clknet_leaf_20_clk));
 sg13g2_buf_2 clkbuf_leaf_21_clk (.A(clknet_3_6__leaf_clk),
    .X(clknet_leaf_21_clk));
 sg13g2_buf_2 clkbuf_leaf_22_clk (.A(clknet_3_6__leaf_clk),
    .X(clknet_leaf_22_clk));
 sg13g2_buf_2 clkbuf_leaf_23_clk (.A(clknet_3_6__leaf_clk),
    .X(clknet_leaf_23_clk));
 sg13g2_buf_2 clkbuf_leaf_24_clk (.A(clknet_3_3__leaf_clk),
    .X(clknet_leaf_24_clk));
 sg13g2_buf_2 clkbuf_leaf_25_clk (.A(clknet_3_3__leaf_clk),
    .X(clknet_leaf_25_clk));
 sg13g2_buf_2 clkbuf_leaf_26_clk (.A(clknet_3_3__leaf_clk),
    .X(clknet_leaf_26_clk));
 sg13g2_buf_2 clkbuf_leaf_27_clk (.A(clknet_3_3__leaf_clk),
    .X(clknet_leaf_27_clk));
 sg13g2_buf_2 clkbuf_leaf_28_clk (.A(clknet_3_3__leaf_clk),
    .X(clknet_leaf_28_clk));
 sg13g2_buf_2 clkbuf_leaf_29_clk (.A(clknet_3_2__leaf_clk),
    .X(clknet_leaf_29_clk));
 sg13g2_buf_2 clkbuf_leaf_30_clk (.A(clknet_3_2__leaf_clk),
    .X(clknet_leaf_30_clk));
 sg13g2_buf_2 clkbuf_leaf_31_clk (.A(clknet_3_2__leaf_clk),
    .X(clknet_leaf_31_clk));
 sg13g2_buf_2 clkbuf_leaf_32_clk (.A(clknet_3_2__leaf_clk),
    .X(clknet_leaf_32_clk));
 sg13g2_buf_2 clkbuf_leaf_33_clk (.A(clknet_3_2__leaf_clk),
    .X(clknet_leaf_33_clk));
 sg13g2_buf_2 clkbuf_leaf_34_clk (.A(clknet_3_1__leaf_clk),
    .X(clknet_leaf_34_clk));
 sg13g2_buf_2 clkbuf_leaf_35_clk (.A(clknet_3_0__leaf_clk),
    .X(clknet_leaf_35_clk));
 sg13g2_buf_2 clkbuf_leaf_36_clk (.A(clknet_3_0__leaf_clk),
    .X(clknet_leaf_36_clk));
 sg13g2_buf_2 clkbuf_leaf_37_clk (.A(clknet_3_0__leaf_clk),
    .X(clknet_leaf_37_clk));
 sg13g2_buf_2 clkbuf_leaf_38_clk (.A(clknet_3_0__leaf_clk),
    .X(clknet_leaf_38_clk));
 sg13g2_buf_2 clkbuf_leaf_39_clk (.A(clknet_3_0__leaf_clk),
    .X(clknet_leaf_39_clk));
 sg13g2_buf_1 clkbuf_0_clk (.A(clk),
    .X(clknet_0_clk));
 sg13g2_buf_1 clkbuf_3_0__f_clk (.A(clknet_0_clk),
    .X(clknet_3_0__leaf_clk));
 sg13g2_buf_1 clkbuf_3_1__f_clk (.A(clknet_0_clk),
    .X(clknet_3_1__leaf_clk));
 sg13g2_buf_1 clkbuf_3_2__f_clk (.A(clknet_0_clk),
    .X(clknet_3_2__leaf_clk));
 sg13g2_buf_1 clkbuf_3_3__f_clk (.A(clknet_0_clk),
    .X(clknet_3_3__leaf_clk));
 sg13g2_buf_1 clkbuf_3_4__f_clk (.A(clknet_0_clk),
    .X(clknet_3_4__leaf_clk));
 sg13g2_buf_1 clkbuf_3_5__f_clk (.A(clknet_0_clk),
    .X(clknet_3_5__leaf_clk));
 sg13g2_buf_1 clkbuf_3_6__f_clk (.A(clknet_0_clk),
    .X(clknet_3_6__leaf_clk));
 sg13g2_buf_1 clkbuf_3_7__f_clk (.A(clknet_0_clk),
    .X(clknet_3_7__leaf_clk));
 sg13g2_antennanp ANTENNA_1 (.A(clk));
 sg13g2_antennanp ANTENNA_2 (.A(clk));
 sg13g2_antennanp ANTENNA_3 (.A(clk));
 sg13g2_antennanp ANTENNA_4 (.A(\g.g_y[1].g_x[7].t.out_r ));
 sg13g2_antennanp ANTENNA_5 (.A(\g.g_y[2].g_x[7].t.out_r ));
 sg13g2_antennanp ANTENNA_6 (.A(\g.g_y[3].g_x[7].t.out_r ));
 sg13g2_antennanp ANTENNA_7 (.A(\g.g_y[1].g_x[7].t.out_r ));
 sg13g2_antennanp ANTENNA_8 (.A(\g.g_y[2].g_x[7].t.out_r ));
 sg13g2_antennanp ANTENNA_9 (.A(\g.g_y[3].g_x[7].t.out_r ));
 sg13g2_antennanp ANTENNA_10 (.A(\g.g_y[1].g_x[7].t.out_r ));
 sg13g2_antennanp ANTENNA_11 (.A(\g.g_y[2].g_x[7].t.out_r ));
 sg13g2_antennanp ANTENNA_12 (.A(\g.g_y[3].g_x[7].t.out_r ));
 sg13g2_antennanp ANTENNA_13 (.A(\g.g_y[1].g_x[7].t.out_r ));
 sg13g2_antennanp ANTENNA_14 (.A(\g.g_y[2].g_x[7].t.out_r ));
 sg13g2_antennanp ANTENNA_15 (.A(\g.g_y[3].g_x[7].t.out_r ));
 sg13g2_antennanp ANTENNA_16 (.A(\g.g_y[1].g_x[7].t.out_r ));
 sg13g2_antennanp ANTENNA_17 (.A(\g.g_y[2].g_x[7].t.out_r ));
 sg13g2_antennanp ANTENNA_18 (.A(\g.g_y[3].g_x[7].t.out_r ));
 sg13g2_decap_8 FILLER_0_0 ();
 sg13g2_decap_8 FILLER_0_7 ();
 sg13g2_decap_8 FILLER_0_14 ();
 sg13g2_decap_8 FILLER_0_21 ();
 sg13g2_decap_8 FILLER_0_28 ();
 sg13g2_decap_8 FILLER_0_35 ();
 sg13g2_decap_8 FILLER_0_42 ();
 sg13g2_decap_8 FILLER_0_49 ();
 sg13g2_decap_8 FILLER_0_56 ();
 sg13g2_decap_8 FILLER_0_63 ();
 sg13g2_decap_8 FILLER_0_70 ();
 sg13g2_decap_8 FILLER_0_77 ();
 sg13g2_decap_8 FILLER_0_84 ();
 sg13g2_decap_8 FILLER_0_91 ();
 sg13g2_decap_8 FILLER_0_102 ();
 sg13g2_decap_8 FILLER_0_114 ();
 sg13g2_fill_2 FILLER_0_121 ();
 sg13g2_fill_1 FILLER_0_123 ();
 sg13g2_decap_4 FILLER_0_128 ();
 sg13g2_fill_1 FILLER_0_132 ();
 sg13g2_decap_8 FILLER_0_138 ();
 sg13g2_decap_4 FILLER_0_145 ();
 sg13g2_fill_2 FILLER_0_149 ();
 sg13g2_decap_8 FILLER_0_169 ();
 sg13g2_decap_4 FILLER_0_176 ();
 sg13g2_fill_2 FILLER_0_180 ();
 sg13g2_fill_2 FILLER_0_190 ();
 sg13g2_fill_1 FILLER_0_192 ();
 sg13g2_decap_4 FILLER_0_245 ();
 sg13g2_fill_2 FILLER_0_249 ();
 sg13g2_decap_8 FILLER_0_255 ();
 sg13g2_fill_1 FILLER_0_262 ();
 sg13g2_fill_1 FILLER_0_268 ();
 sg13g2_decap_4 FILLER_0_273 ();
 sg13g2_fill_1 FILLER_0_277 ();
 sg13g2_decap_4 FILLER_0_282 ();
 sg13g2_decap_4 FILLER_0_299 ();
 sg13g2_fill_1 FILLER_0_303 ();
 sg13g2_decap_4 FILLER_0_308 ();
 sg13g2_fill_2 FILLER_0_312 ();
 sg13g2_decap_8 FILLER_0_319 ();
 sg13g2_fill_1 FILLER_0_326 ();
 sg13g2_decap_4 FILLER_0_337 ();
 sg13g2_fill_1 FILLER_0_341 ();
 sg13g2_decap_8 FILLER_0_346 ();
 sg13g2_decap_8 FILLER_0_353 ();
 sg13g2_decap_8 FILLER_0_360 ();
 sg13g2_decap_8 FILLER_0_367 ();
 sg13g2_decap_8 FILLER_0_374 ();
 sg13g2_decap_8 FILLER_0_381 ();
 sg13g2_decap_8 FILLER_0_388 ();
 sg13g2_decap_8 FILLER_0_395 ();
 sg13g2_decap_8 FILLER_0_402 ();
 sg13g2_decap_8 FILLER_0_409 ();
 sg13g2_decap_8 FILLER_0_416 ();
 sg13g2_decap_8 FILLER_0_423 ();
 sg13g2_decap_8 FILLER_1_0 ();
 sg13g2_decap_8 FILLER_1_7 ();
 sg13g2_decap_8 FILLER_1_14 ();
 sg13g2_decap_8 FILLER_1_21 ();
 sg13g2_decap_8 FILLER_1_28 ();
 sg13g2_decap_8 FILLER_1_35 ();
 sg13g2_decap_8 FILLER_1_42 ();
 sg13g2_decap_8 FILLER_1_49 ();
 sg13g2_decap_8 FILLER_1_56 ();
 sg13g2_decap_8 FILLER_1_63 ();
 sg13g2_decap_8 FILLER_1_70 ();
 sg13g2_decap_8 FILLER_1_77 ();
 sg13g2_decap_8 FILLER_1_84 ();
 sg13g2_fill_1 FILLER_1_143 ();
 sg13g2_fill_1 FILLER_1_185 ();
 sg13g2_fill_1 FILLER_1_212 ();
 sg13g2_fill_1 FILLER_1_244 ();
 sg13g2_fill_2 FILLER_1_333 ();
 sg13g2_decap_8 FILLER_1_361 ();
 sg13g2_decap_8 FILLER_1_368 ();
 sg13g2_decap_8 FILLER_1_375 ();
 sg13g2_decap_8 FILLER_1_382 ();
 sg13g2_decap_8 FILLER_1_389 ();
 sg13g2_decap_8 FILLER_1_396 ();
 sg13g2_decap_8 FILLER_1_403 ();
 sg13g2_decap_8 FILLER_1_410 ();
 sg13g2_decap_8 FILLER_1_417 ();
 sg13g2_decap_4 FILLER_1_424 ();
 sg13g2_fill_2 FILLER_1_428 ();
 sg13g2_decap_8 FILLER_2_0 ();
 sg13g2_decap_8 FILLER_2_7 ();
 sg13g2_decap_8 FILLER_2_14 ();
 sg13g2_decap_8 FILLER_2_21 ();
 sg13g2_decap_8 FILLER_2_28 ();
 sg13g2_decap_8 FILLER_2_35 ();
 sg13g2_decap_8 FILLER_2_42 ();
 sg13g2_decap_8 FILLER_2_49 ();
 sg13g2_decap_8 FILLER_2_56 ();
 sg13g2_decap_8 FILLER_2_63 ();
 sg13g2_decap_8 FILLER_2_70 ();
 sg13g2_decap_8 FILLER_2_77 ();
 sg13g2_decap_4 FILLER_2_84 ();
 sg13g2_fill_1 FILLER_2_102 ();
 sg13g2_fill_1 FILLER_2_118 ();
 sg13g2_fill_1 FILLER_2_124 ();
 sg13g2_fill_2 FILLER_2_197 ();
 sg13g2_fill_1 FILLER_2_209 ();
 sg13g2_fill_2 FILLER_2_251 ();
 sg13g2_fill_1 FILLER_2_253 ();
 sg13g2_fill_1 FILLER_2_331 ();
 sg13g2_decap_8 FILLER_2_362 ();
 sg13g2_decap_8 FILLER_2_369 ();
 sg13g2_decap_8 FILLER_2_376 ();
 sg13g2_decap_8 FILLER_2_383 ();
 sg13g2_decap_8 FILLER_2_390 ();
 sg13g2_decap_8 FILLER_2_397 ();
 sg13g2_decap_8 FILLER_2_404 ();
 sg13g2_decap_8 FILLER_2_411 ();
 sg13g2_decap_8 FILLER_2_418 ();
 sg13g2_decap_4 FILLER_2_425 ();
 sg13g2_fill_1 FILLER_2_429 ();
 sg13g2_decap_8 FILLER_3_0 ();
 sg13g2_decap_8 FILLER_3_7 ();
 sg13g2_decap_8 FILLER_3_14 ();
 sg13g2_decap_8 FILLER_3_21 ();
 sg13g2_decap_8 FILLER_3_28 ();
 sg13g2_decap_8 FILLER_3_35 ();
 sg13g2_decap_8 FILLER_3_42 ();
 sg13g2_decap_4 FILLER_3_49 ();
 sg13g2_fill_2 FILLER_3_53 ();
 sg13g2_decap_8 FILLER_3_59 ();
 sg13g2_decap_8 FILLER_3_66 ();
 sg13g2_decap_8 FILLER_3_73 ();
 sg13g2_decap_4 FILLER_3_80 ();
 sg13g2_fill_1 FILLER_3_198 ();
 sg13g2_decap_8 FILLER_3_203 ();
 sg13g2_fill_1 FILLER_3_210 ();
 sg13g2_fill_1 FILLER_3_216 ();
 sg13g2_fill_1 FILLER_3_231 ();
 sg13g2_decap_4 FILLER_3_236 ();
 sg13g2_fill_2 FILLER_3_245 ();
 sg13g2_fill_1 FILLER_3_273 ();
 sg13g2_fill_2 FILLER_3_310 ();
 sg13g2_decap_8 FILLER_3_359 ();
 sg13g2_decap_8 FILLER_3_366 ();
 sg13g2_decap_8 FILLER_3_373 ();
 sg13g2_decap_8 FILLER_3_380 ();
 sg13g2_decap_8 FILLER_3_387 ();
 sg13g2_decap_8 FILLER_3_394 ();
 sg13g2_decap_8 FILLER_3_401 ();
 sg13g2_decap_8 FILLER_3_408 ();
 sg13g2_decap_8 FILLER_3_415 ();
 sg13g2_decap_8 FILLER_3_422 ();
 sg13g2_fill_1 FILLER_3_429 ();
 sg13g2_decap_8 FILLER_4_0 ();
 sg13g2_decap_8 FILLER_4_7 ();
 sg13g2_decap_8 FILLER_4_14 ();
 sg13g2_decap_8 FILLER_4_21 ();
 sg13g2_decap_8 FILLER_4_28 ();
 sg13g2_decap_8 FILLER_4_35 ();
 sg13g2_decap_4 FILLER_4_42 ();
 sg13g2_fill_1 FILLER_4_46 ();
 sg13g2_fill_1 FILLER_4_103 ();
 sg13g2_fill_1 FILLER_4_109 ();
 sg13g2_fill_1 FILLER_4_132 ();
 sg13g2_fill_1 FILLER_4_160 ();
 sg13g2_fill_1 FILLER_4_184 ();
 sg13g2_fill_1 FILLER_4_228 ();
 sg13g2_fill_1 FILLER_4_234 ();
 sg13g2_decap_4 FILLER_4_240 ();
 sg13g2_fill_2 FILLER_4_244 ();
 sg13g2_fill_1 FILLER_4_259 ();
 sg13g2_fill_1 FILLER_4_264 ();
 sg13g2_fill_2 FILLER_4_270 ();
 sg13g2_fill_1 FILLER_4_272 ();
 sg13g2_fill_1 FILLER_4_318 ();
 sg13g2_fill_1 FILLER_4_324 ();
 sg13g2_fill_2 FILLER_4_343 ();
 sg13g2_decap_8 FILLER_4_375 ();
 sg13g2_decap_8 FILLER_4_382 ();
 sg13g2_decap_8 FILLER_4_389 ();
 sg13g2_decap_8 FILLER_4_396 ();
 sg13g2_decap_8 FILLER_4_403 ();
 sg13g2_decap_8 FILLER_4_410 ();
 sg13g2_decap_8 FILLER_4_417 ();
 sg13g2_decap_4 FILLER_4_424 ();
 sg13g2_fill_2 FILLER_4_428 ();
 sg13g2_decap_8 FILLER_5_0 ();
 sg13g2_decap_8 FILLER_5_7 ();
 sg13g2_decap_8 FILLER_5_14 ();
 sg13g2_decap_8 FILLER_5_21 ();
 sg13g2_decap_8 FILLER_5_28 ();
 sg13g2_decap_8 FILLER_5_35 ();
 sg13g2_decap_8 FILLER_5_42 ();
 sg13g2_fill_2 FILLER_5_49 ();
 sg13g2_decap_8 FILLER_5_60 ();
 sg13g2_fill_2 FILLER_5_67 ();
 sg13g2_fill_2 FILLER_5_74 ();
 sg13g2_fill_1 FILLER_5_76 ();
 sg13g2_fill_2 FILLER_5_104 ();
 sg13g2_fill_1 FILLER_5_119 ();
 sg13g2_fill_1 FILLER_5_124 ();
 sg13g2_fill_1 FILLER_5_130 ();
 sg13g2_fill_1 FILLER_5_135 ();
 sg13g2_decap_8 FILLER_5_141 ();
 sg13g2_decap_4 FILLER_5_148 ();
 sg13g2_fill_1 FILLER_5_156 ();
 sg13g2_fill_1 FILLER_5_162 ();
 sg13g2_fill_1 FILLER_5_172 ();
 sg13g2_fill_1 FILLER_5_178 ();
 sg13g2_fill_1 FILLER_5_189 ();
 sg13g2_fill_2 FILLER_5_194 ();
 sg13g2_fill_2 FILLER_5_201 ();
 sg13g2_decap_4 FILLER_5_207 ();
 sg13g2_fill_1 FILLER_5_211 ();
 sg13g2_fill_1 FILLER_5_217 ();
 sg13g2_decap_8 FILLER_5_226 ();
 sg13g2_decap_4 FILLER_5_233 ();
 sg13g2_fill_2 FILLER_5_237 ();
 sg13g2_fill_2 FILLER_5_244 ();
 sg13g2_fill_2 FILLER_5_249 ();
 sg13g2_fill_2 FILLER_5_256 ();
 sg13g2_fill_1 FILLER_5_258 ();
 sg13g2_fill_2 FILLER_5_268 ();
 sg13g2_fill_1 FILLER_5_274 ();
 sg13g2_fill_2 FILLER_5_284 ();
 sg13g2_fill_1 FILLER_5_286 ();
 sg13g2_decap_4 FILLER_5_295 ();
 sg13g2_fill_2 FILLER_5_299 ();
 sg13g2_decap_4 FILLER_5_306 ();
 sg13g2_decap_4 FILLER_5_314 ();
 sg13g2_fill_1 FILLER_5_318 ();
 sg13g2_fill_2 FILLER_5_328 ();
 sg13g2_decap_8 FILLER_5_396 ();
 sg13g2_fill_2 FILLER_5_403 ();
 sg13g2_fill_1 FILLER_5_405 ();
 sg13g2_decap_8 FILLER_5_410 ();
 sg13g2_decap_8 FILLER_5_417 ();
 sg13g2_decap_4 FILLER_5_424 ();
 sg13g2_fill_2 FILLER_5_428 ();
 sg13g2_decap_8 FILLER_6_0 ();
 sg13g2_decap_8 FILLER_6_7 ();
 sg13g2_decap_8 FILLER_6_14 ();
 sg13g2_decap_8 FILLER_6_21 ();
 sg13g2_decap_8 FILLER_6_28 ();
 sg13g2_decap_4 FILLER_6_35 ();
 sg13g2_decap_8 FILLER_6_69 ();
 sg13g2_decap_4 FILLER_6_76 ();
 sg13g2_decap_4 FILLER_6_84 ();
 sg13g2_fill_2 FILLER_6_93 ();
 sg13g2_fill_1 FILLER_6_103 ();
 sg13g2_fill_1 FILLER_6_122 ();
 sg13g2_decap_8 FILLER_6_180 ();
 sg13g2_decap_4 FILLER_6_187 ();
 sg13g2_fill_1 FILLER_6_191 ();
 sg13g2_fill_2 FILLER_6_218 ();
 sg13g2_fill_1 FILLER_6_220 ();
 sg13g2_fill_1 FILLER_6_251 ();
 sg13g2_fill_2 FILLER_6_257 ();
 sg13g2_fill_2 FILLER_6_264 ();
 sg13g2_fill_2 FILLER_6_292 ();
 sg13g2_fill_1 FILLER_6_294 ();
 sg13g2_decap_8 FILLER_6_400 ();
 sg13g2_decap_8 FILLER_6_407 ();
 sg13g2_decap_8 FILLER_6_414 ();
 sg13g2_decap_8 FILLER_6_421 ();
 sg13g2_fill_2 FILLER_6_428 ();
 sg13g2_decap_8 FILLER_7_0 ();
 sg13g2_decap_8 FILLER_7_7 ();
 sg13g2_decap_8 FILLER_7_14 ();
 sg13g2_decap_8 FILLER_7_21 ();
 sg13g2_decap_8 FILLER_7_28 ();
 sg13g2_decap_8 FILLER_7_35 ();
 sg13g2_decap_4 FILLER_7_42 ();
 sg13g2_fill_2 FILLER_7_50 ();
 sg13g2_fill_1 FILLER_7_52 ();
 sg13g2_fill_1 FILLER_7_92 ();
 sg13g2_fill_2 FILLER_7_180 ();
 sg13g2_fill_1 FILLER_7_182 ();
 sg13g2_fill_1 FILLER_7_274 ();
 sg13g2_fill_2 FILLER_7_289 ();
 sg13g2_fill_2 FILLER_7_378 ();
 sg13g2_fill_2 FILLER_7_384 ();
 sg13g2_decap_8 FILLER_7_412 ();
 sg13g2_decap_8 FILLER_7_419 ();
 sg13g2_decap_4 FILLER_7_426 ();
 sg13g2_decap_8 FILLER_8_0 ();
 sg13g2_decap_8 FILLER_8_7 ();
 sg13g2_decap_8 FILLER_8_14 ();
 sg13g2_decap_8 FILLER_8_21 ();
 sg13g2_decap_8 FILLER_8_28 ();
 sg13g2_decap_8 FILLER_8_35 ();
 sg13g2_decap_8 FILLER_8_42 ();
 sg13g2_fill_1 FILLER_8_49 ();
 sg13g2_fill_2 FILLER_8_148 ();
 sg13g2_fill_1 FILLER_8_155 ();
 sg13g2_fill_2 FILLER_8_179 ();
 sg13g2_fill_2 FILLER_8_211 ();
 sg13g2_fill_2 FILLER_8_297 ();
 sg13g2_fill_1 FILLER_8_304 ();
 sg13g2_fill_2 FILLER_8_329 ();
 sg13g2_fill_2 FILLER_8_336 ();
 sg13g2_decap_4 FILLER_8_342 ();
 sg13g2_fill_2 FILLER_8_346 ();
 sg13g2_fill_2 FILLER_8_372 ();
 sg13g2_fill_1 FILLER_8_404 ();
 sg13g2_decap_8 FILLER_8_409 ();
 sg13g2_decap_8 FILLER_8_416 ();
 sg13g2_decap_8 FILLER_8_423 ();
 sg13g2_decap_8 FILLER_9_0 ();
 sg13g2_decap_8 FILLER_9_7 ();
 sg13g2_decap_8 FILLER_9_14 ();
 sg13g2_decap_8 FILLER_9_21 ();
 sg13g2_decap_4 FILLER_9_28 ();
 sg13g2_decap_8 FILLER_9_36 ();
 sg13g2_fill_1 FILLER_9_43 ();
 sg13g2_fill_2 FILLER_9_57 ();
 sg13g2_fill_1 FILLER_9_59 ();
 sg13g2_fill_1 FILLER_9_107 ();
 sg13g2_fill_2 FILLER_9_118 ();
 sg13g2_fill_2 FILLER_9_125 ();
 sg13g2_fill_2 FILLER_9_153 ();
 sg13g2_fill_1 FILLER_9_155 ();
 sg13g2_fill_1 FILLER_9_176 ();
 sg13g2_fill_1 FILLER_9_217 ();
 sg13g2_fill_1 FILLER_9_228 ();
 sg13g2_fill_1 FILLER_9_234 ();
 sg13g2_fill_1 FILLER_9_255 ();
 sg13g2_fill_1 FILLER_9_276 ();
 sg13g2_fill_2 FILLER_9_296 ();
 sg13g2_fill_1 FILLER_9_298 ();
 sg13g2_decap_4 FILLER_9_329 ();
 sg13g2_fill_1 FILLER_9_333 ();
 sg13g2_fill_2 FILLER_9_339 ();
 sg13g2_fill_2 FILLER_9_399 ();
 sg13g2_decap_8 FILLER_9_406 ();
 sg13g2_decap_8 FILLER_9_413 ();
 sg13g2_decap_8 FILLER_9_420 ();
 sg13g2_fill_2 FILLER_9_427 ();
 sg13g2_fill_1 FILLER_9_429 ();
 sg13g2_decap_8 FILLER_10_0 ();
 sg13g2_decap_8 FILLER_10_7 ();
 sg13g2_decap_8 FILLER_10_14 ();
 sg13g2_decap_4 FILLER_10_21 ();
 sg13g2_fill_1 FILLER_10_51 ();
 sg13g2_fill_1 FILLER_10_64 ();
 sg13g2_fill_2 FILLER_10_85 ();
 sg13g2_fill_1 FILLER_10_97 ();
 sg13g2_fill_1 FILLER_10_105 ();
 sg13g2_fill_2 FILLER_10_109 ();
 sg13g2_fill_2 FILLER_10_116 ();
 sg13g2_decap_8 FILLER_10_122 ();
 sg13g2_decap_4 FILLER_10_129 ();
 sg13g2_fill_1 FILLER_10_133 ();
 sg13g2_fill_1 FILLER_10_142 ();
 sg13g2_fill_2 FILLER_10_161 ();
 sg13g2_fill_1 FILLER_10_217 ();
 sg13g2_decap_4 FILLER_10_223 ();
 sg13g2_fill_2 FILLER_10_242 ();
 sg13g2_fill_1 FILLER_10_244 ();
 sg13g2_decap_8 FILLER_10_250 ();
 sg13g2_fill_1 FILLER_10_257 ();
 sg13g2_fill_1 FILLER_10_268 ();
 sg13g2_fill_2 FILLER_10_285 ();
 sg13g2_fill_1 FILLER_10_337 ();
 sg13g2_fill_2 FILLER_10_342 ();
 sg13g2_decap_8 FILLER_10_402 ();
 sg13g2_decap_8 FILLER_10_409 ();
 sg13g2_decap_8 FILLER_10_416 ();
 sg13g2_decap_8 FILLER_10_423 ();
 sg13g2_decap_8 FILLER_11_0 ();
 sg13g2_decap_8 FILLER_11_7 ();
 sg13g2_decap_8 FILLER_11_14 ();
 sg13g2_decap_8 FILLER_11_21 ();
 sg13g2_decap_8 FILLER_11_28 ();
 sg13g2_decap_4 FILLER_11_35 ();
 sg13g2_fill_2 FILLER_11_39 ();
 sg13g2_fill_1 FILLER_11_51 ();
 sg13g2_decap_4 FILLER_11_82 ();
 sg13g2_fill_2 FILLER_11_86 ();
 sg13g2_decap_8 FILLER_11_92 ();
 sg13g2_fill_1 FILLER_11_105 ();
 sg13g2_decap_8 FILLER_11_121 ();
 sg13g2_fill_1 FILLER_11_183 ();
 sg13g2_fill_2 FILLER_11_189 ();
 sg13g2_fill_1 FILLER_11_205 ();
 sg13g2_decap_4 FILLER_11_232 ();
 sg13g2_fill_2 FILLER_11_241 ();
 sg13g2_fill_1 FILLER_11_243 ();
 sg13g2_fill_2 FILLER_11_248 ();
 sg13g2_decap_8 FILLER_11_255 ();
 sg13g2_fill_1 FILLER_11_270 ();
 sg13g2_fill_1 FILLER_11_284 ();
 sg13g2_fill_2 FILLER_11_290 ();
 sg13g2_fill_1 FILLER_11_341 ();
 sg13g2_fill_1 FILLER_11_347 ();
 sg13g2_fill_1 FILLER_11_353 ();
 sg13g2_fill_1 FILLER_11_374 ();
 sg13g2_fill_2 FILLER_11_382 ();
 sg13g2_fill_1 FILLER_11_384 ();
 sg13g2_decap_8 FILLER_11_415 ();
 sg13g2_decap_8 FILLER_11_422 ();
 sg13g2_fill_1 FILLER_11_429 ();
 sg13g2_decap_8 FILLER_12_0 ();
 sg13g2_decap_8 FILLER_12_7 ();
 sg13g2_decap_4 FILLER_12_14 ();
 sg13g2_fill_2 FILLER_12_18 ();
 sg13g2_fill_2 FILLER_12_91 ();
 sg13g2_decap_8 FILLER_12_97 ();
 sg13g2_decap_4 FILLER_12_104 ();
 sg13g2_fill_1 FILLER_12_108 ();
 sg13g2_fill_1 FILLER_12_148 ();
 sg13g2_fill_2 FILLER_12_155 ();
 sg13g2_fill_2 FILLER_12_168 ();
 sg13g2_decap_8 FILLER_12_190 ();
 sg13g2_fill_2 FILLER_12_197 ();
 sg13g2_fill_1 FILLER_12_199 ();
 sg13g2_decap_8 FILLER_12_205 ();
 sg13g2_fill_2 FILLER_12_212 ();
 sg13g2_fill_2 FILLER_12_218 ();
 sg13g2_fill_1 FILLER_12_220 ();
 sg13g2_fill_1 FILLER_12_230 ();
 sg13g2_fill_1 FILLER_12_283 ();
 sg13g2_fill_2 FILLER_12_289 ();
 sg13g2_fill_1 FILLER_12_295 ();
 sg13g2_fill_2 FILLER_12_302 ();
 sg13g2_fill_2 FILLER_12_309 ();
 sg13g2_fill_2 FILLER_12_318 ();
 sg13g2_fill_1 FILLER_12_320 ();
 sg13g2_decap_8 FILLER_12_383 ();
 sg13g2_fill_2 FILLER_12_390 ();
 sg13g2_decap_8 FILLER_12_412 ();
 sg13g2_decap_8 FILLER_12_419 ();
 sg13g2_decap_4 FILLER_12_426 ();
 sg13g2_decap_8 FILLER_13_0 ();
 sg13g2_decap_8 FILLER_13_7 ();
 sg13g2_decap_8 FILLER_13_14 ();
 sg13g2_decap_8 FILLER_13_21 ();
 sg13g2_decap_4 FILLER_13_28 ();
 sg13g2_fill_1 FILLER_13_32 ();
 sg13g2_decap_8 FILLER_13_37 ();
 sg13g2_decap_8 FILLER_13_44 ();
 sg13g2_decap_4 FILLER_13_51 ();
 sg13g2_fill_1 FILLER_13_65 ();
 sg13g2_fill_2 FILLER_13_75 ();
 sg13g2_fill_1 FILLER_13_83 ();
 sg13g2_decap_8 FILLER_13_98 ();
 sg13g2_fill_2 FILLER_13_125 ();
 sg13g2_decap_4 FILLER_13_168 ();
 sg13g2_decap_8 FILLER_13_202 ();
 sg13g2_fill_1 FILLER_13_214 ();
 sg13g2_fill_1 FILLER_13_220 ();
 sg13g2_fill_2 FILLER_13_224 ();
 sg13g2_fill_1 FILLER_13_226 ();
 sg13g2_decap_4 FILLER_13_253 ();
 sg13g2_fill_2 FILLER_13_261 ();
 sg13g2_decap_4 FILLER_13_273 ();
 sg13g2_fill_1 FILLER_13_287 ();
 sg13g2_fill_2 FILLER_13_397 ();
 sg13g2_decap_8 FILLER_13_403 ();
 sg13g2_decap_8 FILLER_13_414 ();
 sg13g2_decap_8 FILLER_13_421 ();
 sg13g2_fill_2 FILLER_13_428 ();
 sg13g2_decap_8 FILLER_14_0 ();
 sg13g2_decap_8 FILLER_14_7 ();
 sg13g2_decap_8 FILLER_14_14 ();
 sg13g2_decap_8 FILLER_14_21 ();
 sg13g2_decap_8 FILLER_14_28 ();
 sg13g2_fill_2 FILLER_14_40 ();
 sg13g2_decap_4 FILLER_14_52 ();
 sg13g2_fill_2 FILLER_14_56 ();
 sg13g2_fill_1 FILLER_14_67 ();
 sg13g2_fill_1 FILLER_14_75 ();
 sg13g2_fill_2 FILLER_14_94 ();
 sg13g2_fill_1 FILLER_14_96 ();
 sg13g2_decap_8 FILLER_14_136 ();
 sg13g2_decap_8 FILLER_14_143 ();
 sg13g2_decap_8 FILLER_14_160 ();
 sg13g2_fill_1 FILLER_14_177 ();
 sg13g2_fill_1 FILLER_14_236 ();
 sg13g2_decap_8 FILLER_14_241 ();
 sg13g2_decap_8 FILLER_14_248 ();
 sg13g2_decap_8 FILLER_14_255 ();
 sg13g2_fill_2 FILLER_14_262 ();
 sg13g2_fill_1 FILLER_14_273 ();
 sg13g2_fill_2 FILLER_14_279 ();
 sg13g2_fill_1 FILLER_14_290 ();
 sg13g2_fill_1 FILLER_14_295 ();
 sg13g2_fill_1 FILLER_14_302 ();
 sg13g2_fill_2 FILLER_14_308 ();
 sg13g2_fill_1 FILLER_14_348 ();
 sg13g2_fill_1 FILLER_14_354 ();
 sg13g2_fill_1 FILLER_14_360 ();
 sg13g2_fill_1 FILLER_14_365 ();
 sg13g2_fill_1 FILLER_14_380 ();
 sg13g2_fill_1 FILLER_14_385 ();
 sg13g2_decap_8 FILLER_14_412 ();
 sg13g2_decap_8 FILLER_14_419 ();
 sg13g2_decap_4 FILLER_14_426 ();
 sg13g2_decap_8 FILLER_15_0 ();
 sg13g2_decap_8 FILLER_15_7 ();
 sg13g2_decap_8 FILLER_15_14 ();
 sg13g2_decap_8 FILLER_15_21 ();
 sg13g2_fill_2 FILLER_15_28 ();
 sg13g2_fill_1 FILLER_15_136 ();
 sg13g2_fill_1 FILLER_15_142 ();
 sg13g2_fill_1 FILLER_15_148 ();
 sg13g2_fill_2 FILLER_15_159 ();
 sg13g2_fill_2 FILLER_15_165 ();
 sg13g2_fill_1 FILLER_15_167 ();
 sg13g2_fill_2 FILLER_15_178 ();
 sg13g2_fill_2 FILLER_15_195 ();
 sg13g2_fill_1 FILLER_15_197 ();
 sg13g2_decap_4 FILLER_15_211 ();
 sg13g2_fill_2 FILLER_15_215 ();
 sg13g2_decap_4 FILLER_15_232 ();
 sg13g2_decap_4 FILLER_15_255 ();
 sg13g2_fill_1 FILLER_15_259 ();
 sg13g2_fill_1 FILLER_15_270 ();
 sg13g2_decap_4 FILLER_15_274 ();
 sg13g2_fill_1 FILLER_15_278 ();
 sg13g2_fill_2 FILLER_15_286 ();
 sg13g2_decap_4 FILLER_15_293 ();
 sg13g2_decap_8 FILLER_15_306 ();
 sg13g2_decap_8 FILLER_15_361 ();
 sg13g2_decap_4 FILLER_15_368 ();
 sg13g2_fill_2 FILLER_15_372 ();
 sg13g2_fill_1 FILLER_15_384 ();
 sg13g2_decap_8 FILLER_15_405 ();
 sg13g2_decap_8 FILLER_15_412 ();
 sg13g2_decap_8 FILLER_15_419 ();
 sg13g2_decap_4 FILLER_15_426 ();
 sg13g2_decap_8 FILLER_16_0 ();
 sg13g2_decap_8 FILLER_16_7 ();
 sg13g2_decap_8 FILLER_16_14 ();
 sg13g2_decap_8 FILLER_16_21 ();
 sg13g2_decap_8 FILLER_16_28 ();
 sg13g2_decap_4 FILLER_16_35 ();
 sg13g2_fill_1 FILLER_16_39 ();
 sg13g2_fill_1 FILLER_16_44 ();
 sg13g2_fill_2 FILLER_16_99 ();
 sg13g2_fill_2 FILLER_16_137 ();
 sg13g2_fill_1 FILLER_16_139 ();
 sg13g2_fill_1 FILLER_16_189 ();
 sg13g2_fill_2 FILLER_16_194 ();
 sg13g2_fill_1 FILLER_16_201 ();
 sg13g2_fill_2 FILLER_16_222 ();
 sg13g2_fill_1 FILLER_16_224 ();
 sg13g2_fill_2 FILLER_16_234 ();
 sg13g2_fill_1 FILLER_16_236 ();
 sg13g2_fill_1 FILLER_16_251 ();
 sg13g2_decap_8 FILLER_16_277 ();
 sg13g2_fill_1 FILLER_16_284 ();
 sg13g2_fill_1 FILLER_16_308 ();
 sg13g2_fill_1 FILLER_16_314 ();
 sg13g2_decap_8 FILLER_16_356 ();
 sg13g2_fill_2 FILLER_16_363 ();
 sg13g2_fill_1 FILLER_16_365 ();
 sg13g2_fill_2 FILLER_16_371 ();
 sg13g2_fill_2 FILLER_16_393 ();
 sg13g2_fill_2 FILLER_16_400 ();
 sg13g2_fill_1 FILLER_16_402 ();
 sg13g2_decap_4 FILLER_16_407 ();
 sg13g2_fill_1 FILLER_16_411 ();
 sg13g2_decap_8 FILLER_16_417 ();
 sg13g2_decap_4 FILLER_16_424 ();
 sg13g2_fill_2 FILLER_16_428 ();
 sg13g2_decap_8 FILLER_17_0 ();
 sg13g2_decap_8 FILLER_17_7 ();
 sg13g2_decap_8 FILLER_17_14 ();
 sg13g2_decap_8 FILLER_17_21 ();
 sg13g2_decap_8 FILLER_17_28 ();
 sg13g2_decap_4 FILLER_17_35 ();
 sg13g2_decap_4 FILLER_17_43 ();
 sg13g2_fill_2 FILLER_17_60 ();
 sg13g2_fill_1 FILLER_17_85 ();
 sg13g2_fill_2 FILLER_17_106 ();
 sg13g2_fill_1 FILLER_17_123 ();
 sg13g2_fill_2 FILLER_17_165 ();
 sg13g2_fill_1 FILLER_17_177 ();
 sg13g2_fill_2 FILLER_17_188 ();
 sg13g2_fill_1 FILLER_17_190 ();
 sg13g2_fill_1 FILLER_17_196 ();
 sg13g2_fill_1 FILLER_17_203 ();
 sg13g2_fill_1 FILLER_17_228 ();
 sg13g2_decap_4 FILLER_17_310 ();
 sg13g2_fill_1 FILLER_17_344 ();
 sg13g2_decap_4 FILLER_17_350 ();
 sg13g2_fill_2 FILLER_17_367 ();
 sg13g2_decap_4 FILLER_17_426 ();
 sg13g2_decap_8 FILLER_18_0 ();
 sg13g2_decap_8 FILLER_18_7 ();
 sg13g2_decap_8 FILLER_18_14 ();
 sg13g2_decap_8 FILLER_18_21 ();
 sg13g2_decap_4 FILLER_18_28 ();
 sg13g2_fill_1 FILLER_18_63 ();
 sg13g2_fill_1 FILLER_18_68 ();
 sg13g2_fill_1 FILLER_18_73 ();
 sg13g2_decap_4 FILLER_18_79 ();
 sg13g2_fill_2 FILLER_18_83 ();
 sg13g2_fill_2 FILLER_18_90 ();
 sg13g2_fill_2 FILLER_18_107 ();
 sg13g2_fill_1 FILLER_18_109 ();
 sg13g2_fill_2 FILLER_18_115 ();
 sg13g2_fill_2 FILLER_18_127 ();
 sg13g2_fill_1 FILLER_18_149 ();
 sg13g2_fill_2 FILLER_18_155 ();
 sg13g2_fill_1 FILLER_18_157 ();
 sg13g2_decap_8 FILLER_18_163 ();
 sg13g2_decap_4 FILLER_18_170 ();
 sg13g2_fill_2 FILLER_18_227 ();
 sg13g2_fill_1 FILLER_18_257 ();
 sg13g2_fill_1 FILLER_18_268 ();
 sg13g2_fill_1 FILLER_18_272 ();
 sg13g2_fill_2 FILLER_18_282 ();
 sg13g2_fill_1 FILLER_18_293 ();
 sg13g2_fill_1 FILLER_18_299 ();
 sg13g2_fill_2 FILLER_18_305 ();
 sg13g2_fill_1 FILLER_18_307 ();
 sg13g2_decap_4 FILLER_18_312 ();
 sg13g2_fill_1 FILLER_18_316 ();
 sg13g2_fill_2 FILLER_18_321 ();
 sg13g2_fill_1 FILLER_18_323 ();
 sg13g2_fill_2 FILLER_18_339 ();
 sg13g2_fill_1 FILLER_18_341 ();
 sg13g2_fill_1 FILLER_18_346 ();
 sg13g2_fill_2 FILLER_18_357 ();
 sg13g2_fill_1 FILLER_18_359 ();
 sg13g2_fill_1 FILLER_18_386 ();
 sg13g2_fill_1 FILLER_18_392 ();
 sg13g2_fill_2 FILLER_18_423 ();
 sg13g2_fill_1 FILLER_18_425 ();
 sg13g2_decap_8 FILLER_19_0 ();
 sg13g2_decap_8 FILLER_19_7 ();
 sg13g2_decap_8 FILLER_19_14 ();
 sg13g2_fill_2 FILLER_19_21 ();
 sg13g2_fill_2 FILLER_19_77 ();
 sg13g2_fill_2 FILLER_19_84 ();
 sg13g2_fill_1 FILLER_19_86 ();
 sg13g2_fill_2 FILLER_19_92 ();
 sg13g2_fill_1 FILLER_19_94 ();
 sg13g2_decap_4 FILLER_19_99 ();
 sg13g2_fill_2 FILLER_19_103 ();
 sg13g2_decap_4 FILLER_19_126 ();
 sg13g2_fill_2 FILLER_19_130 ();
 sg13g2_decap_8 FILLER_19_136 ();
 sg13g2_fill_2 FILLER_19_143 ();
 sg13g2_fill_1 FILLER_19_200 ();
 sg13g2_fill_2 FILLER_19_204 ();
 sg13g2_fill_1 FILLER_19_206 ();
 sg13g2_decap_4 FILLER_19_212 ();
 sg13g2_decap_8 FILLER_19_221 ();
 sg13g2_fill_1 FILLER_19_228 ();
 sg13g2_fill_1 FILLER_19_237 ();
 sg13g2_decap_4 FILLER_19_286 ();
 sg13g2_fill_2 FILLER_19_294 ();
 sg13g2_decap_4 FILLER_19_332 ();
 sg13g2_fill_2 FILLER_19_336 ();
 sg13g2_fill_1 FILLER_19_373 ();
 sg13g2_decap_8 FILLER_19_393 ();
 sg13g2_decap_8 FILLER_20_0 ();
 sg13g2_decap_8 FILLER_20_7 ();
 sg13g2_decap_8 FILLER_20_14 ();
 sg13g2_fill_2 FILLER_20_21 ();
 sg13g2_fill_1 FILLER_20_23 ();
 sg13g2_fill_2 FILLER_20_55 ();
 sg13g2_fill_2 FILLER_20_62 ();
 sg13g2_fill_2 FILLER_20_69 ();
 sg13g2_fill_1 FILLER_20_71 ();
 sg13g2_fill_1 FILLER_20_80 ();
 sg13g2_fill_1 FILLER_20_86 ();
 sg13g2_fill_1 FILLER_20_113 ();
 sg13g2_fill_2 FILLER_20_140 ();
 sg13g2_fill_2 FILLER_20_150 ();
 sg13g2_fill_1 FILLER_20_152 ();
 sg13g2_fill_2 FILLER_20_157 ();
 sg13g2_fill_2 FILLER_20_163 ();
 sg13g2_fill_2 FILLER_20_169 ();
 sg13g2_fill_1 FILLER_20_171 ();
 sg13g2_fill_2 FILLER_20_176 ();
 sg13g2_fill_1 FILLER_20_178 ();
 sg13g2_fill_1 FILLER_20_183 ();
 sg13g2_fill_1 FILLER_20_189 ();
 sg13g2_fill_1 FILLER_20_194 ();
 sg13g2_fill_1 FILLER_20_205 ();
 sg13g2_fill_2 FILLER_20_225 ();
 sg13g2_fill_1 FILLER_20_227 ();
 sg13g2_fill_1 FILLER_20_238 ();
 sg13g2_fill_2 FILLER_20_249 ();
 sg13g2_fill_1 FILLER_20_309 ();
 sg13g2_decap_4 FILLER_20_367 ();
 sg13g2_decap_4 FILLER_20_375 ();
 sg13g2_fill_2 FILLER_20_379 ();
 sg13g2_fill_1 FILLER_20_419 ();
 sg13g2_fill_1 FILLER_20_424 ();
 sg13g2_decap_8 FILLER_21_0 ();
 sg13g2_decap_8 FILLER_21_7 ();
 sg13g2_decap_8 FILLER_21_14 ();
 sg13g2_decap_4 FILLER_21_21 ();
 sg13g2_fill_2 FILLER_21_25 ();
 sg13g2_fill_2 FILLER_21_41 ();
 sg13g2_fill_1 FILLER_21_48 ();
 sg13g2_fill_1 FILLER_21_54 ();
 sg13g2_fill_2 FILLER_21_103 ();
 sg13g2_fill_2 FILLER_21_166 ();
 sg13g2_fill_1 FILLER_21_292 ();
 sg13g2_fill_2 FILLER_21_298 ();
 sg13g2_fill_2 FILLER_21_304 ();
 sg13g2_fill_1 FILLER_21_306 ();
 sg13g2_decap_4 FILLER_21_313 ();
 sg13g2_fill_1 FILLER_21_317 ();
 sg13g2_decap_4 FILLER_21_322 ();
 sg13g2_fill_1 FILLER_21_326 ();
 sg13g2_fill_2 FILLER_21_331 ();
 sg13g2_fill_1 FILLER_21_333 ();
 sg13g2_fill_1 FILLER_21_338 ();
 sg13g2_fill_1 FILLER_21_349 ();
 sg13g2_decap_4 FILLER_21_355 ();
 sg13g2_fill_2 FILLER_21_367 ();
 sg13g2_fill_1 FILLER_21_369 ();
 sg13g2_fill_2 FILLER_21_405 ();
 sg13g2_fill_1 FILLER_21_411 ();
 sg13g2_fill_2 FILLER_21_427 ();
 sg13g2_fill_1 FILLER_21_429 ();
 sg13g2_decap_8 FILLER_22_0 ();
 sg13g2_decap_8 FILLER_22_7 ();
 sg13g2_fill_1 FILLER_22_55 ();
 sg13g2_decap_4 FILLER_22_62 ();
 sg13g2_fill_2 FILLER_22_94 ();
 sg13g2_fill_2 FILLER_22_101 ();
 sg13g2_decap_4 FILLER_22_107 ();
 sg13g2_fill_1 FILLER_22_116 ();
 sg13g2_fill_2 FILLER_22_122 ();
 sg13g2_fill_2 FILLER_22_128 ();
 sg13g2_fill_2 FILLER_22_135 ();
 sg13g2_fill_1 FILLER_22_137 ();
 sg13g2_fill_1 FILLER_22_192 ();
 sg13g2_fill_2 FILLER_22_239 ();
 sg13g2_fill_1 FILLER_22_241 ();
 sg13g2_fill_2 FILLER_22_247 ();
 sg13g2_fill_1 FILLER_22_249 ();
 sg13g2_fill_2 FILLER_22_260 ();
 sg13g2_fill_1 FILLER_22_305 ();
 sg13g2_fill_1 FILLER_22_342 ();
 sg13g2_fill_2 FILLER_22_347 ();
 sg13g2_fill_2 FILLER_22_363 ();
 sg13g2_fill_1 FILLER_22_370 ();
 sg13g2_fill_2 FILLER_22_397 ();
 sg13g2_fill_2 FILLER_22_404 ();
 sg13g2_fill_1 FILLER_22_406 ();
 sg13g2_fill_1 FILLER_22_423 ();
 sg13g2_fill_1 FILLER_22_429 ();
 sg13g2_decap_4 FILLER_23_0 ();
 sg13g2_fill_1 FILLER_23_48 ();
 sg13g2_fill_1 FILLER_23_54 ();
 sg13g2_fill_1 FILLER_23_73 ();
 sg13g2_fill_1 FILLER_23_97 ();
 sg13g2_fill_1 FILLER_23_134 ();
 sg13g2_fill_1 FILLER_23_165 ();
 sg13g2_fill_1 FILLER_23_191 ();
 sg13g2_fill_1 FILLER_23_204 ();
 sg13g2_fill_1 FILLER_23_209 ();
 sg13g2_fill_2 FILLER_23_280 ();
 sg13g2_fill_1 FILLER_23_296 ();
 sg13g2_fill_2 FILLER_23_302 ();
 sg13g2_fill_1 FILLER_23_308 ();
 sg13g2_fill_2 FILLER_23_314 ();
 sg13g2_fill_2 FILLER_23_320 ();
 sg13g2_fill_2 FILLER_23_325 ();
 sg13g2_fill_2 FILLER_23_375 ();
 sg13g2_fill_1 FILLER_23_377 ();
 sg13g2_decap_4 FILLER_23_425 ();
 sg13g2_fill_1 FILLER_23_429 ();
 sg13g2_decap_8 FILLER_24_0 ();
 sg13g2_decap_8 FILLER_24_7 ();
 sg13g2_decap_4 FILLER_24_14 ();
 sg13g2_fill_2 FILLER_24_73 ();
 sg13g2_fill_2 FILLER_24_120 ();
 sg13g2_fill_1 FILLER_24_127 ();
 sg13g2_fill_1 FILLER_24_133 ();
 sg13g2_fill_1 FILLER_24_156 ();
 sg13g2_fill_1 FILLER_24_161 ();
 sg13g2_fill_2 FILLER_24_171 ();
 sg13g2_decap_8 FILLER_24_203 ();
 sg13g2_decap_8 FILLER_24_210 ();
 sg13g2_fill_1 FILLER_24_217 ();
 sg13g2_decap_4 FILLER_24_222 ();
 sg13g2_fill_2 FILLER_24_230 ();
 sg13g2_fill_1 FILLER_24_232 ();
 sg13g2_decap_8 FILLER_24_261 ();
 sg13g2_fill_2 FILLER_24_268 ();
 sg13g2_fill_1 FILLER_24_270 ();
 sg13g2_decap_4 FILLER_24_288 ();
 sg13g2_fill_1 FILLER_24_292 ();
 sg13g2_fill_1 FILLER_24_301 ();
 sg13g2_fill_1 FILLER_24_309 ();
 sg13g2_fill_1 FILLER_24_314 ();
 sg13g2_fill_1 FILLER_24_320 ();
 sg13g2_fill_1 FILLER_24_325 ();
 sg13g2_fill_1 FILLER_24_384 ();
 sg13g2_fill_1 FILLER_24_390 ();
 sg13g2_fill_2 FILLER_24_410 ();
 sg13g2_fill_2 FILLER_24_422 ();
 sg13g2_fill_1 FILLER_24_424 ();
 sg13g2_decap_8 FILLER_25_0 ();
 sg13g2_decap_8 FILLER_25_7 ();
 sg13g2_decap_8 FILLER_25_14 ();
 sg13g2_decap_8 FILLER_25_21 ();
 sg13g2_decap_4 FILLER_25_28 ();
 sg13g2_fill_1 FILLER_25_32 ();
 sg13g2_decap_8 FILLER_25_37 ();
 sg13g2_fill_2 FILLER_25_44 ();
 sg13g2_fill_1 FILLER_25_55 ();
 sg13g2_decap_4 FILLER_25_60 ();
 sg13g2_fill_2 FILLER_25_68 ();
 sg13g2_fill_1 FILLER_25_70 ();
 sg13g2_decap_4 FILLER_25_80 ();
 sg13g2_fill_1 FILLER_25_84 ();
 sg13g2_fill_1 FILLER_25_99 ();
 sg13g2_fill_1 FILLER_25_110 ();
 sg13g2_fill_2 FILLER_25_158 ();
 sg13g2_fill_1 FILLER_25_165 ();
 sg13g2_fill_2 FILLER_25_170 ();
 sg13g2_fill_1 FILLER_25_220 ();
 sg13g2_fill_2 FILLER_25_236 ();
 sg13g2_fill_2 FILLER_25_248 ();
 sg13g2_fill_1 FILLER_25_250 ();
 sg13g2_decap_8 FILLER_25_266 ();
 sg13g2_decap_8 FILLER_25_273 ();
 sg13g2_fill_1 FILLER_25_280 ();
 sg13g2_fill_2 FILLER_25_338 ();
 sg13g2_fill_2 FILLER_25_428 ();
 sg13g2_decap_8 FILLER_26_0 ();
 sg13g2_decap_8 FILLER_26_7 ();
 sg13g2_decap_8 FILLER_26_14 ();
 sg13g2_decap_8 FILLER_26_21 ();
 sg13g2_decap_4 FILLER_26_28 ();
 sg13g2_fill_1 FILLER_26_32 ();
 sg13g2_decap_4 FILLER_26_72 ();
 sg13g2_fill_1 FILLER_26_76 ();
 sg13g2_fill_2 FILLER_26_81 ();
 sg13g2_decap_4 FILLER_26_88 ();
 sg13g2_fill_1 FILLER_26_116 ();
 sg13g2_fill_1 FILLER_26_121 ();
 sg13g2_fill_1 FILLER_26_127 ();
 sg13g2_fill_2 FILLER_26_206 ();
 sg13g2_fill_2 FILLER_26_239 ();
 sg13g2_fill_2 FILLER_26_281 ();
 sg13g2_fill_1 FILLER_26_293 ();
 sg13g2_fill_1 FILLER_26_300 ();
 sg13g2_fill_1 FILLER_26_363 ();
 sg13g2_fill_1 FILLER_26_369 ();
 sg13g2_fill_2 FILLER_26_375 ();
 sg13g2_fill_1 FILLER_26_384 ();
 sg13g2_fill_2 FILLER_26_399 ();
 sg13g2_decap_4 FILLER_27_0 ();
 sg13g2_fill_1 FILLER_27_4 ();
 sg13g2_fill_1 FILLER_27_36 ();
 sg13g2_fill_1 FILLER_27_45 ();
 sg13g2_fill_1 FILLER_27_61 ();
 sg13g2_decap_4 FILLER_27_72 ();
 sg13g2_fill_1 FILLER_27_86 ();
 sg13g2_fill_1 FILLER_27_101 ();
 sg13g2_fill_1 FILLER_27_109 ();
 sg13g2_fill_1 FILLER_27_142 ();
 sg13g2_fill_1 FILLER_27_153 ();
 sg13g2_fill_1 FILLER_27_225 ();
 sg13g2_fill_1 FILLER_27_251 ();
 sg13g2_fill_1 FILLER_27_278 ();
 sg13g2_fill_2 FILLER_27_331 ();
 sg13g2_fill_2 FILLER_27_361 ();
 sg13g2_fill_1 FILLER_27_363 ();
 sg13g2_fill_1 FILLER_27_429 ();
 sg13g2_decap_8 FILLER_28_0 ();
 sg13g2_fill_1 FILLER_28_7 ();
 sg13g2_fill_1 FILLER_28_42 ();
 sg13g2_fill_1 FILLER_28_72 ();
 sg13g2_fill_2 FILLER_28_107 ();
 sg13g2_fill_1 FILLER_28_109 ();
 sg13g2_fill_1 FILLER_28_170 ();
 sg13g2_fill_2 FILLER_28_176 ();
 sg13g2_fill_2 FILLER_28_229 ();
 sg13g2_fill_2 FILLER_28_265 ();
 sg13g2_fill_1 FILLER_28_276 ();
 sg13g2_fill_1 FILLER_28_281 ();
 sg13g2_fill_1 FILLER_28_292 ();
 sg13g2_fill_2 FILLER_28_297 ();
 sg13g2_fill_2 FILLER_28_309 ();
 sg13g2_fill_1 FILLER_28_311 ();
 sg13g2_fill_1 FILLER_28_387 ();
 sg13g2_fill_2 FILLER_28_393 ();
 sg13g2_fill_1 FILLER_28_395 ();
 sg13g2_fill_2 FILLER_28_401 ();
 sg13g2_fill_1 FILLER_28_429 ();
 sg13g2_decap_8 FILLER_29_0 ();
 sg13g2_decap_4 FILLER_29_7 ();
 sg13g2_fill_1 FILLER_29_11 ();
 sg13g2_decap_8 FILLER_29_16 ();
 sg13g2_fill_2 FILLER_29_23 ();
 sg13g2_fill_1 FILLER_29_25 ();
 sg13g2_fill_2 FILLER_29_102 ();
 sg13g2_decap_8 FILLER_29_138 ();
 sg13g2_fill_2 FILLER_29_167 ();
 sg13g2_fill_1 FILLER_29_195 ();
 sg13g2_fill_2 FILLER_29_230 ();
 sg13g2_decap_4 FILLER_29_246 ();
 sg13g2_fill_1 FILLER_29_250 ();
 sg13g2_fill_2 FILLER_29_255 ();
 sg13g2_decap_8 FILLER_29_266 ();
 sg13g2_fill_2 FILLER_29_273 ();
 sg13g2_fill_1 FILLER_29_275 ();
 sg13g2_fill_2 FILLER_29_286 ();
 sg13g2_fill_1 FILLER_29_288 ();
 sg13g2_fill_2 FILLER_29_293 ();
 sg13g2_fill_1 FILLER_29_295 ();
 sg13g2_fill_1 FILLER_29_310 ();
 sg13g2_fill_1 FILLER_29_316 ();
 sg13g2_fill_1 FILLER_29_322 ();
 sg13g2_fill_1 FILLER_29_349 ();
 sg13g2_fill_1 FILLER_29_376 ();
 sg13g2_fill_1 FILLER_29_382 ();
 sg13g2_fill_1 FILLER_29_392 ();
 sg13g2_fill_1 FILLER_29_407 ();
 sg13g2_decap_4 FILLER_29_413 ();
 sg13g2_decap_4 FILLER_29_426 ();
 sg13g2_decap_8 FILLER_30_0 ();
 sg13g2_decap_8 FILLER_30_7 ();
 sg13g2_decap_8 FILLER_30_14 ();
 sg13g2_fill_2 FILLER_30_21 ();
 sg13g2_fill_2 FILLER_30_54 ();
 sg13g2_fill_2 FILLER_30_75 ();
 sg13g2_fill_2 FILLER_30_130 ();
 sg13g2_fill_1 FILLER_30_136 ();
 sg13g2_decap_8 FILLER_30_140 ();
 sg13g2_fill_2 FILLER_30_147 ();
 sg13g2_fill_2 FILLER_30_179 ();
 sg13g2_fill_1 FILLER_30_211 ();
 sg13g2_fill_1 FILLER_30_218 ();
 sg13g2_fill_1 FILLER_30_245 ();
 sg13g2_fill_1 FILLER_30_255 ();
 sg13g2_fill_1 FILLER_30_266 ();
 sg13g2_fill_1 FILLER_30_272 ();
 sg13g2_fill_2 FILLER_30_338 ();
 sg13g2_fill_1 FILLER_30_340 ();
 sg13g2_fill_1 FILLER_30_351 ();
 sg13g2_fill_1 FILLER_30_357 ();
 sg13g2_fill_1 FILLER_30_362 ();
 sg13g2_decap_4 FILLER_30_408 ();
 sg13g2_fill_2 FILLER_30_412 ();
 sg13g2_decap_8 FILLER_30_418 ();
 sg13g2_fill_1 FILLER_30_429 ();
 sg13g2_decap_8 FILLER_31_0 ();
 sg13g2_decap_8 FILLER_31_7 ();
 sg13g2_decap_8 FILLER_31_14 ();
 sg13g2_decap_4 FILLER_31_21 ();
 sg13g2_fill_2 FILLER_31_33 ();
 sg13g2_fill_1 FILLER_31_48 ();
 sg13g2_decap_4 FILLER_31_57 ();
 sg13g2_fill_2 FILLER_31_61 ();
 sg13g2_decap_8 FILLER_31_78 ();
 sg13g2_decap_8 FILLER_31_85 ();
 sg13g2_fill_2 FILLER_31_92 ();
 sg13g2_decap_4 FILLER_31_98 ();
 sg13g2_fill_1 FILLER_31_102 ();
 sg13g2_fill_1 FILLER_31_126 ();
 sg13g2_fill_2 FILLER_31_153 ();
 sg13g2_fill_1 FILLER_31_155 ();
 sg13g2_fill_1 FILLER_31_172 ();
 sg13g2_fill_1 FILLER_31_197 ();
 sg13g2_decap_8 FILLER_31_202 ();
 sg13g2_fill_1 FILLER_31_209 ();
 sg13g2_fill_2 FILLER_31_218 ();
 sg13g2_fill_1 FILLER_31_228 ();
 sg13g2_fill_1 FILLER_31_233 ();
 sg13g2_fill_1 FILLER_31_239 ();
 sg13g2_fill_1 FILLER_31_246 ();
 sg13g2_fill_1 FILLER_31_272 ();
 sg13g2_fill_2 FILLER_31_277 ();
 sg13g2_fill_1 FILLER_31_284 ();
 sg13g2_fill_2 FILLER_31_289 ();
 sg13g2_fill_1 FILLER_31_296 ();
 sg13g2_fill_2 FILLER_31_303 ();
 sg13g2_fill_2 FILLER_31_347 ();
 sg13g2_decap_8 FILLER_31_354 ();
 sg13g2_fill_1 FILLER_31_374 ();
 sg13g2_fill_1 FILLER_31_383 ();
 sg13g2_fill_2 FILLER_31_394 ();
 sg13g2_fill_2 FILLER_31_402 ();
 sg13g2_decap_8 FILLER_32_0 ();
 sg13g2_decap_8 FILLER_32_7 ();
 sg13g2_decap_8 FILLER_32_14 ();
 sg13g2_decap_4 FILLER_32_21 ();
 sg13g2_fill_2 FILLER_32_25 ();
 sg13g2_fill_1 FILLER_32_52 ();
 sg13g2_fill_1 FILLER_32_62 ();
 sg13g2_fill_2 FILLER_32_111 ();
 sg13g2_decap_4 FILLER_32_118 ();
 sg13g2_fill_1 FILLER_32_147 ();
 sg13g2_fill_2 FILLER_32_153 ();
 sg13g2_fill_1 FILLER_32_155 ();
 sg13g2_fill_2 FILLER_32_176 ();
 sg13g2_fill_1 FILLER_32_178 ();
 sg13g2_decap_8 FILLER_32_205 ();
 sg13g2_fill_1 FILLER_32_212 ();
 sg13g2_fill_1 FILLER_32_248 ();
 sg13g2_fill_1 FILLER_32_280 ();
 sg13g2_decap_8 FILLER_32_284 ();
 sg13g2_fill_2 FILLER_32_291 ();
 sg13g2_fill_1 FILLER_32_301 ();
 sg13g2_fill_2 FILLER_32_306 ();
 sg13g2_fill_2 FILLER_32_329 ();
 sg13g2_fill_2 FILLER_32_336 ();
 sg13g2_fill_1 FILLER_32_338 ();
 sg13g2_decap_4 FILLER_32_370 ();
 sg13g2_fill_1 FILLER_32_374 ();
 sg13g2_fill_2 FILLER_32_399 ();
 sg13g2_fill_2 FILLER_32_427 ();
 sg13g2_fill_1 FILLER_32_429 ();
 sg13g2_decap_8 FILLER_33_0 ();
 sg13g2_fill_1 FILLER_33_33 ();
 sg13g2_fill_1 FILLER_33_39 ();
 sg13g2_fill_1 FILLER_33_55 ();
 sg13g2_fill_1 FILLER_33_97 ();
 sg13g2_fill_1 FILLER_33_108 ();
 sg13g2_fill_1 FILLER_33_157 ();
 sg13g2_fill_1 FILLER_33_162 ();
 sg13g2_fill_1 FILLER_33_183 ();
 sg13g2_fill_1 FILLER_33_206 ();
 sg13g2_fill_2 FILLER_33_211 ();
 sg13g2_decap_4 FILLER_33_228 ();
 sg13g2_fill_1 FILLER_33_232 ();
 sg13g2_decap_4 FILLER_33_238 ();
 sg13g2_fill_1 FILLER_33_242 ();
 sg13g2_decap_4 FILLER_33_248 ();
 sg13g2_fill_1 FILLER_33_252 ();
 sg13g2_fill_1 FILLER_33_288 ();
 sg13g2_fill_1 FILLER_33_311 ();
 sg13g2_fill_1 FILLER_33_316 ();
 sg13g2_fill_1 FILLER_33_327 ();
 sg13g2_decap_4 FILLER_33_332 ();
 sg13g2_decap_4 FILLER_33_341 ();
 sg13g2_fill_2 FILLER_33_345 ();
 sg13g2_fill_1 FILLER_33_351 ();
 sg13g2_decap_8 FILLER_33_362 ();
 sg13g2_fill_1 FILLER_33_369 ();
 sg13g2_fill_2 FILLER_33_395 ();
 sg13g2_decap_8 FILLER_33_411 ();
 sg13g2_decap_8 FILLER_33_418 ();
 sg13g2_decap_4 FILLER_33_425 ();
 sg13g2_fill_1 FILLER_33_429 ();
 sg13g2_decap_8 FILLER_34_0 ();
 sg13g2_decap_8 FILLER_34_7 ();
 sg13g2_fill_2 FILLER_34_14 ();
 sg13g2_decap_8 FILLER_34_20 ();
 sg13g2_decap_4 FILLER_34_27 ();
 sg13g2_fill_2 FILLER_34_51 ();
 sg13g2_fill_2 FILLER_34_193 ();
 sg13g2_fill_1 FILLER_34_225 ();
 sg13g2_fill_1 FILLER_34_235 ();
 sg13g2_fill_1 FILLER_34_241 ();
 sg13g2_fill_1 FILLER_34_247 ();
 sg13g2_fill_2 FILLER_34_253 ();
 sg13g2_fill_1 FILLER_34_321 ();
 sg13g2_fill_1 FILLER_34_332 ();
 sg13g2_fill_1 FILLER_34_347 ();
 sg13g2_fill_1 FILLER_34_382 ();
 sg13g2_fill_1 FILLER_34_388 ();
 sg13g2_fill_1 FILLER_34_394 ();
 sg13g2_fill_2 FILLER_34_405 ();
 sg13g2_decap_4 FILLER_34_424 ();
 sg13g2_fill_2 FILLER_34_428 ();
 sg13g2_decap_8 FILLER_35_0 ();
 sg13g2_decap_4 FILLER_35_7 ();
 sg13g2_fill_2 FILLER_35_11 ();
 sg13g2_fill_2 FILLER_35_17 ();
 sg13g2_decap_4 FILLER_35_39 ();
 sg13g2_fill_1 FILLER_35_70 ();
 sg13g2_decap_8 FILLER_35_114 ();
 sg13g2_fill_2 FILLER_35_149 ();
 sg13g2_fill_1 FILLER_35_151 ();
 sg13g2_fill_1 FILLER_35_156 ();
 sg13g2_fill_2 FILLER_35_166 ();
 sg13g2_decap_4 FILLER_35_173 ();
 sg13g2_fill_2 FILLER_35_252 ();
 sg13g2_fill_2 FILLER_35_279 ();
 sg13g2_decap_4 FILLER_35_363 ();
 sg13g2_fill_2 FILLER_35_397 ();
 sg13g2_decap_4 FILLER_36_0 ();
 sg13g2_fill_2 FILLER_36_4 ();
 sg13g2_fill_2 FILLER_36_32 ();
 sg13g2_fill_1 FILLER_36_34 ();
 sg13g2_fill_1 FILLER_36_65 ();
 sg13g2_fill_2 FILLER_36_70 ();
 sg13g2_fill_1 FILLER_36_72 ();
 sg13g2_fill_2 FILLER_36_102 ();
 sg13g2_fill_1 FILLER_36_109 ();
 sg13g2_decap_4 FILLER_36_115 ();
 sg13g2_fill_2 FILLER_36_119 ();
 sg13g2_fill_1 FILLER_36_139 ();
 sg13g2_fill_1 FILLER_36_149 ();
 sg13g2_fill_2 FILLER_36_162 ();
 sg13g2_fill_1 FILLER_36_164 ();
 sg13g2_fill_2 FILLER_36_216 ();
 sg13g2_fill_1 FILLER_36_223 ();
 sg13g2_fill_1 FILLER_36_250 ();
 sg13g2_fill_1 FILLER_36_265 ();
 sg13g2_decap_4 FILLER_36_271 ();
 sg13g2_fill_2 FILLER_36_279 ();
 sg13g2_fill_1 FILLER_36_281 ();
 sg13g2_decap_4 FILLER_36_286 ();
 sg13g2_fill_1 FILLER_36_290 ();
 sg13g2_decap_4 FILLER_36_295 ();
 sg13g2_fill_1 FILLER_36_299 ();
 sg13g2_decap_4 FILLER_36_305 ();
 sg13g2_fill_1 FILLER_36_314 ();
 sg13g2_fill_1 FILLER_36_320 ();
 sg13g2_fill_1 FILLER_36_328 ();
 sg13g2_fill_1 FILLER_36_339 ();
 sg13g2_fill_2 FILLER_36_366 ();
 sg13g2_fill_2 FILLER_36_394 ();
 sg13g2_decap_8 FILLER_37_0 ();
 sg13g2_fill_2 FILLER_37_7 ();
 sg13g2_fill_1 FILLER_37_9 ();
 sg13g2_fill_2 FILLER_37_49 ();
 sg13g2_decap_8 FILLER_37_83 ();
 sg13g2_fill_2 FILLER_37_90 ();
 sg13g2_fill_2 FILLER_37_127 ();
 sg13g2_fill_1 FILLER_37_129 ();
 sg13g2_fill_2 FILLER_37_160 ();
 sg13g2_fill_1 FILLER_37_167 ();
 sg13g2_fill_1 FILLER_37_172 ();
 sg13g2_fill_2 FILLER_37_188 ();
 sg13g2_fill_2 FILLER_37_194 ();
 sg13g2_fill_1 FILLER_37_196 ();
 sg13g2_fill_2 FILLER_37_202 ();
 sg13g2_fill_1 FILLER_37_204 ();
 sg13g2_fill_1 FILLER_37_209 ();
 sg13g2_fill_2 FILLER_37_215 ();
 sg13g2_fill_2 FILLER_37_222 ();
 sg13g2_fill_2 FILLER_37_229 ();
 sg13g2_fill_2 FILLER_37_235 ();
 sg13g2_fill_2 FILLER_37_242 ();
 sg13g2_fill_1 FILLER_37_244 ();
 sg13g2_fill_1 FILLER_37_249 ();
 sg13g2_fill_2 FILLER_37_258 ();
 sg13g2_fill_2 FILLER_37_269 ();
 sg13g2_decap_4 FILLER_37_276 ();
 sg13g2_fill_2 FILLER_37_280 ();
 sg13g2_decap_4 FILLER_37_308 ();
 sg13g2_decap_4 FILLER_37_322 ();
 sg13g2_fill_1 FILLER_37_381 ();
 sg13g2_decap_4 FILLER_37_397 ();
 sg13g2_fill_1 FILLER_37_401 ();
 sg13g2_fill_2 FILLER_37_407 ();
 sg13g2_fill_1 FILLER_37_413 ();
 sg13g2_fill_2 FILLER_37_427 ();
 sg13g2_fill_1 FILLER_37_429 ();
 sg13g2_decap_4 FILLER_38_0 ();
 sg13g2_fill_2 FILLER_38_43 ();
 sg13g2_fill_2 FILLER_38_54 ();
 sg13g2_fill_2 FILLER_38_61 ();
 sg13g2_fill_1 FILLER_38_63 ();
 sg13g2_fill_1 FILLER_38_69 ();
 sg13g2_fill_2 FILLER_38_96 ();
 sg13g2_fill_1 FILLER_38_98 ();
 sg13g2_fill_1 FILLER_38_108 ();
 sg13g2_fill_1 FILLER_38_140 ();
 sg13g2_fill_2 FILLER_38_145 ();
 sg13g2_decap_8 FILLER_38_211 ();
 sg13g2_fill_2 FILLER_38_218 ();
 sg13g2_fill_1 FILLER_38_220 ();
 sg13g2_decap_4 FILLER_38_225 ();
 sg13g2_fill_1 FILLER_38_229 ();
 sg13g2_decap_4 FILLER_38_298 ();
 sg13g2_fill_1 FILLER_38_302 ();
 sg13g2_decap_8 FILLER_38_307 ();
 sg13g2_fill_2 FILLER_38_314 ();
 sg13g2_fill_1 FILLER_38_316 ();
 sg13g2_decap_8 FILLER_38_322 ();
 sg13g2_fill_2 FILLER_38_329 ();
 sg13g2_fill_1 FILLER_38_331 ();
 sg13g2_fill_2 FILLER_38_337 ();
 sg13g2_fill_1 FILLER_38_339 ();
 sg13g2_fill_2 FILLER_38_354 ();
 sg13g2_fill_2 FILLER_38_361 ();
 sg13g2_fill_2 FILLER_38_367 ();
 sg13g2_fill_1 FILLER_38_369 ();
 sg13g2_decap_4 FILLER_38_375 ();
 sg13g2_fill_1 FILLER_38_379 ();
 sg13g2_fill_2 FILLER_38_389 ();
 sg13g2_decap_8 FILLER_39_0 ();
 sg13g2_fill_1 FILLER_39_7 ();
 sg13g2_fill_2 FILLER_39_98 ();
 sg13g2_fill_1 FILLER_39_100 ();
 sg13g2_fill_1 FILLER_39_142 ();
 sg13g2_fill_1 FILLER_39_148 ();
 sg13g2_fill_2 FILLER_39_159 ();
 sg13g2_fill_1 FILLER_39_182 ();
 sg13g2_decap_8 FILLER_39_216 ();
 sg13g2_decap_8 FILLER_39_287 ();
 sg13g2_fill_2 FILLER_39_294 ();
 sg13g2_fill_2 FILLER_39_322 ();
 sg13g2_fill_1 FILLER_39_324 ();
 sg13g2_decap_4 FILLER_39_328 ();
 sg13g2_fill_1 FILLER_39_332 ();
 sg13g2_fill_1 FILLER_39_341 ();
 sg13g2_fill_1 FILLER_39_368 ();
 sg13g2_fill_1 FILLER_39_395 ();
 sg13g2_fill_1 FILLER_39_411 ();
 sg13g2_fill_2 FILLER_39_427 ();
 sg13g2_fill_1 FILLER_39_429 ();
 sg13g2_decap_8 FILLER_40_0 ();
 sg13g2_decap_8 FILLER_40_7 ();
 sg13g2_fill_2 FILLER_40_14 ();
 sg13g2_decap_8 FILLER_40_20 ();
 sg13g2_decap_4 FILLER_40_27 ();
 sg13g2_fill_1 FILLER_40_31 ();
 sg13g2_decap_8 FILLER_40_36 ();
 sg13g2_fill_1 FILLER_40_43 ();
 sg13g2_fill_2 FILLER_40_48 ();
 sg13g2_fill_2 FILLER_40_55 ();
 sg13g2_decap_8 FILLER_40_62 ();
 sg13g2_decap_4 FILLER_40_69 ();
 sg13g2_fill_1 FILLER_40_73 ();
 sg13g2_decap_8 FILLER_40_101 ();
 sg13g2_decap_8 FILLER_40_114 ();
 sg13g2_fill_1 FILLER_40_121 ();
 sg13g2_fill_1 FILLER_40_126 ();
 sg13g2_fill_2 FILLER_40_131 ();
 sg13g2_fill_1 FILLER_40_137 ();
 sg13g2_fill_2 FILLER_40_142 ();
 sg13g2_fill_1 FILLER_40_217 ();
 sg13g2_decap_8 FILLER_40_252 ();
 sg13g2_decap_4 FILLER_40_259 ();
 sg13g2_fill_1 FILLER_40_263 ();
 sg13g2_fill_2 FILLER_40_268 ();
 sg13g2_fill_1 FILLER_40_270 ();
 sg13g2_fill_2 FILLER_40_275 ();
 sg13g2_fill_2 FILLER_40_281 ();
 sg13g2_fill_1 FILLER_40_283 ();
 sg13g2_fill_1 FILLER_40_294 ();
 sg13g2_fill_1 FILLER_40_309 ();
 sg13g2_fill_2 FILLER_40_330 ();
 sg13g2_fill_1 FILLER_40_380 ();
 sg13g2_decap_8 FILLER_40_390 ();
 sg13g2_fill_2 FILLER_40_397 ();
 sg13g2_decap_8 FILLER_41_0 ();
 sg13g2_decap_8 FILLER_41_7 ();
 sg13g2_decap_4 FILLER_41_14 ();
 sg13g2_fill_1 FILLER_41_54 ();
 sg13g2_fill_2 FILLER_41_60 ();
 sg13g2_fill_2 FILLER_41_66 ();
 sg13g2_fill_2 FILLER_41_73 ();
 sg13g2_fill_1 FILLER_41_75 ();
 sg13g2_fill_2 FILLER_41_106 ();
 sg13g2_fill_2 FILLER_41_112 ();
 sg13g2_fill_1 FILLER_41_114 ();
 sg13g2_fill_2 FILLER_41_120 ();
 sg13g2_fill_1 FILLER_41_122 ();
 sg13g2_decap_4 FILLER_41_170 ();
 sg13g2_fill_1 FILLER_41_174 ();
 sg13g2_fill_2 FILLER_41_184 ();
 sg13g2_fill_1 FILLER_41_186 ();
 sg13g2_decap_8 FILLER_41_199 ();
 sg13g2_fill_2 FILLER_41_211 ();
 sg13g2_decap_4 FILLER_41_220 ();
 sg13g2_fill_2 FILLER_41_224 ();
 sg13g2_decap_8 FILLER_41_238 ();
 sg13g2_fill_1 FILLER_41_245 ();
 sg13g2_fill_2 FILLER_41_250 ();
 sg13g2_fill_1 FILLER_41_257 ();
 sg13g2_decap_4 FILLER_41_262 ();
 sg13g2_fill_1 FILLER_41_266 ();
 sg13g2_fill_1 FILLER_41_336 ();
 sg13g2_fill_2 FILLER_41_370 ();
 sg13g2_fill_1 FILLER_41_372 ();
 sg13g2_fill_2 FILLER_41_387 ();
 sg13g2_fill_1 FILLER_41_389 ();
 sg13g2_decap_4 FILLER_41_395 ();
 sg13g2_fill_2 FILLER_41_399 ();
 sg13g2_fill_1 FILLER_41_429 ();
 sg13g2_decap_8 FILLER_42_0 ();
 sg13g2_decap_8 FILLER_42_7 ();
 sg13g2_decap_4 FILLER_42_14 ();
 sg13g2_fill_1 FILLER_42_18 ();
 sg13g2_fill_1 FILLER_42_49 ();
 sg13g2_fill_2 FILLER_42_55 ();
 sg13g2_fill_2 FILLER_42_83 ();
 sg13g2_fill_2 FILLER_42_132 ();
 sg13g2_fill_1 FILLER_42_134 ();
 sg13g2_fill_1 FILLER_42_166 ();
 sg13g2_fill_1 FILLER_42_172 ();
 sg13g2_fill_2 FILLER_42_179 ();
 sg13g2_decap_4 FILLER_42_190 ();
 sg13g2_fill_2 FILLER_42_194 ();
 sg13g2_decap_4 FILLER_42_235 ();
 sg13g2_fill_2 FILLER_42_239 ();
 sg13g2_fill_1 FILLER_42_259 ();
 sg13g2_decap_4 FILLER_42_269 ();
 sg13g2_fill_1 FILLER_42_273 ();
 sg13g2_fill_2 FILLER_42_347 ();
 sg13g2_fill_2 FILLER_42_374 ();
 sg13g2_fill_1 FILLER_42_401 ();
 sg13g2_fill_2 FILLER_42_427 ();
 sg13g2_fill_1 FILLER_42_429 ();
 sg13g2_decap_8 FILLER_43_0 ();
 sg13g2_decap_8 FILLER_43_7 ();
 sg13g2_decap_8 FILLER_43_14 ();
 sg13g2_decap_8 FILLER_43_21 ();
 sg13g2_fill_1 FILLER_43_37 ();
 sg13g2_fill_2 FILLER_43_42 ();
 sg13g2_fill_1 FILLER_43_49 ();
 sg13g2_fill_1 FILLER_43_124 ();
 sg13g2_fill_1 FILLER_43_190 ();
 sg13g2_fill_2 FILLER_43_201 ();
 sg13g2_fill_1 FILLER_43_203 ();
 sg13g2_fill_2 FILLER_43_218 ();
 sg13g2_fill_1 FILLER_43_220 ();
 sg13g2_fill_2 FILLER_43_248 ();
 sg13g2_fill_2 FILLER_43_300 ();
 sg13g2_fill_2 FILLER_43_312 ();
 sg13g2_fill_1 FILLER_43_314 ();
 sg13g2_fill_2 FILLER_43_331 ();
 sg13g2_fill_1 FILLER_43_348 ();
 sg13g2_fill_2 FILLER_43_395 ();
 sg13g2_decap_4 FILLER_43_424 ();
 sg13g2_fill_2 FILLER_43_428 ();
 sg13g2_decap_8 FILLER_44_0 ();
 sg13g2_decap_8 FILLER_44_7 ();
 sg13g2_decap_8 FILLER_44_14 ();
 sg13g2_decap_8 FILLER_44_21 ();
 sg13g2_decap_8 FILLER_44_28 ();
 sg13g2_fill_2 FILLER_44_35 ();
 sg13g2_decap_4 FILLER_44_47 ();
 sg13g2_fill_2 FILLER_44_51 ();
 sg13g2_decap_4 FILLER_44_58 ();
 sg13g2_fill_1 FILLER_44_66 ();
 sg13g2_fill_1 FILLER_44_77 ();
 sg13g2_fill_1 FILLER_44_88 ();
 sg13g2_fill_2 FILLER_44_99 ();
 sg13g2_fill_1 FILLER_44_106 ();
 sg13g2_fill_2 FILLER_44_111 ();
 sg13g2_fill_1 FILLER_44_113 ();
 sg13g2_fill_2 FILLER_44_141 ();
 sg13g2_fill_1 FILLER_44_148 ();
 sg13g2_fill_2 FILLER_44_176 ();
 sg13g2_fill_2 FILLER_44_181 ();
 sg13g2_fill_1 FILLER_44_183 ();
 sg13g2_fill_1 FILLER_44_194 ();
 sg13g2_fill_2 FILLER_44_200 ();
 sg13g2_fill_1 FILLER_44_202 ();
 sg13g2_decap_4 FILLER_44_229 ();
 sg13g2_fill_2 FILLER_44_233 ();
 sg13g2_fill_1 FILLER_44_312 ();
 sg13g2_fill_1 FILLER_44_318 ();
 sg13g2_fill_2 FILLER_44_338 ();
 sg13g2_decap_4 FILLER_44_344 ();
 sg13g2_fill_2 FILLER_44_354 ();
 sg13g2_fill_1 FILLER_44_356 ();
 sg13g2_fill_2 FILLER_44_367 ();
 sg13g2_fill_2 FILLER_44_404 ();
 sg13g2_decap_4 FILLER_44_426 ();
 sg13g2_decap_8 FILLER_45_0 ();
 sg13g2_decap_8 FILLER_45_7 ();
 sg13g2_fill_2 FILLER_45_14 ();
 sg13g2_fill_1 FILLER_45_16 ();
 sg13g2_decap_4 FILLER_45_47 ();
 sg13g2_decap_8 FILLER_45_71 ();
 sg13g2_decap_4 FILLER_45_78 ();
 sg13g2_fill_2 FILLER_45_86 ();
 sg13g2_decap_4 FILLER_45_93 ();
 sg13g2_fill_1 FILLER_45_116 ();
 sg13g2_fill_2 FILLER_45_127 ();
 sg13g2_fill_2 FILLER_45_133 ();
 sg13g2_decap_8 FILLER_45_140 ();
 sg13g2_fill_2 FILLER_45_163 ();
 sg13g2_fill_1 FILLER_45_170 ();
 sg13g2_fill_2 FILLER_45_203 ();
 sg13g2_fill_2 FILLER_45_215 ();
 sg13g2_fill_1 FILLER_45_217 ();
 sg13g2_fill_2 FILLER_45_281 ();
 sg13g2_fill_1 FILLER_45_283 ();
 sg13g2_decap_8 FILLER_45_314 ();
 sg13g2_decap_8 FILLER_45_321 ();
 sg13g2_fill_2 FILLER_45_328 ();
 sg13g2_decap_4 FILLER_45_335 ();
 sg13g2_fill_2 FILLER_45_344 ();
 sg13g2_fill_1 FILLER_45_346 ();
 sg13g2_decap_4 FILLER_45_361 ();
 sg13g2_fill_2 FILLER_45_365 ();
 sg13g2_fill_2 FILLER_45_373 ();
 sg13g2_decap_4 FILLER_45_425 ();
 sg13g2_fill_1 FILLER_45_429 ();
 sg13g2_decap_8 FILLER_46_0 ();
 sg13g2_decap_8 FILLER_46_7 ();
 sg13g2_decap_8 FILLER_46_14 ();
 sg13g2_fill_1 FILLER_46_21 ();
 sg13g2_decap_4 FILLER_46_32 ();
 sg13g2_fill_2 FILLER_46_46 ();
 sg13g2_fill_2 FILLER_46_58 ();
 sg13g2_fill_1 FILLER_46_60 ();
 sg13g2_fill_1 FILLER_46_64 ();
 sg13g2_decap_8 FILLER_46_73 ();
 sg13g2_fill_2 FILLER_46_106 ();
 sg13g2_fill_2 FILLER_46_115 ();
 sg13g2_fill_1 FILLER_46_117 ();
 sg13g2_fill_2 FILLER_46_138 ();
 sg13g2_fill_1 FILLER_46_140 ();
 sg13g2_fill_2 FILLER_46_146 ();
 sg13g2_fill_1 FILLER_46_148 ();
 sg13g2_fill_2 FILLER_46_154 ();
 sg13g2_decap_8 FILLER_46_160 ();
 sg13g2_fill_1 FILLER_46_167 ();
 sg13g2_fill_2 FILLER_46_172 ();
 sg13g2_fill_1 FILLER_46_224 ();
 sg13g2_fill_1 FILLER_46_229 ();
 sg13g2_fill_1 FILLER_46_253 ();
 sg13g2_fill_2 FILLER_46_259 ();
 sg13g2_fill_1 FILLER_46_275 ();
 sg13g2_fill_1 FILLER_46_286 ();
 sg13g2_fill_1 FILLER_46_296 ();
 sg13g2_fill_1 FILLER_46_343 ();
 sg13g2_fill_1 FILLER_46_351 ();
 sg13g2_fill_1 FILLER_46_362 ();
 sg13g2_fill_1 FILLER_46_423 ();
 sg13g2_fill_1 FILLER_46_429 ();
 sg13g2_decap_8 FILLER_47_0 ();
 sg13g2_fill_1 FILLER_47_7 ();
 sg13g2_decap_4 FILLER_47_34 ();
 sg13g2_fill_1 FILLER_47_48 ();
 sg13g2_fill_1 FILLER_47_79 ();
 sg13g2_fill_1 FILLER_47_85 ();
 sg13g2_fill_2 FILLER_47_112 ();
 sg13g2_fill_2 FILLER_47_180 ();
 sg13g2_decap_4 FILLER_47_186 ();
 sg13g2_decap_4 FILLER_47_209 ();
 sg13g2_fill_2 FILLER_47_213 ();
 sg13g2_fill_2 FILLER_47_219 ();
 sg13g2_fill_1 FILLER_47_221 ();
 sg13g2_fill_2 FILLER_47_241 ();
 sg13g2_fill_1 FILLER_47_247 ();
 sg13g2_fill_1 FILLER_47_253 ();
 sg13g2_decap_4 FILLER_47_262 ();
 sg13g2_decap_8 FILLER_47_271 ();
 sg13g2_fill_2 FILLER_47_283 ();
 sg13g2_fill_2 FILLER_47_292 ();
 sg13g2_fill_1 FILLER_47_294 ();
 sg13g2_fill_2 FILLER_47_300 ();
 sg13g2_fill_1 FILLER_47_302 ();
 sg13g2_decap_4 FILLER_47_308 ();
 sg13g2_fill_1 FILLER_47_312 ();
 sg13g2_decap_4 FILLER_47_317 ();
 sg13g2_fill_1 FILLER_47_321 ();
 sg13g2_fill_1 FILLER_47_332 ();
 sg13g2_fill_1 FILLER_47_373 ();
 sg13g2_fill_1 FILLER_47_394 ();
 sg13g2_fill_2 FILLER_48_0 ();
 sg13g2_fill_1 FILLER_48_2 ();
 sg13g2_decap_4 FILLER_48_51 ();
 sg13g2_fill_1 FILLER_48_55 ();
 sg13g2_fill_2 FILLER_48_91 ();
 sg13g2_fill_1 FILLER_48_93 ();
 sg13g2_fill_1 FILLER_48_137 ();
 sg13g2_fill_1 FILLER_48_148 ();
 sg13g2_fill_1 FILLER_48_184 ();
 sg13g2_fill_1 FILLER_48_190 ();
 sg13g2_fill_2 FILLER_48_195 ();
 sg13g2_fill_2 FILLER_48_212 ();
 sg13g2_fill_2 FILLER_48_219 ();
 sg13g2_fill_2 FILLER_48_226 ();
 sg13g2_fill_2 FILLER_48_277 ();
 sg13g2_fill_1 FILLER_48_285 ();
 sg13g2_fill_1 FILLER_48_293 ();
 sg13g2_fill_1 FILLER_48_299 ();
 sg13g2_fill_1 FILLER_48_336 ();
 sg13g2_fill_1 FILLER_48_342 ();
 sg13g2_fill_1 FILLER_48_360 ();
 sg13g2_fill_1 FILLER_48_365 ();
 sg13g2_fill_1 FILLER_48_397 ();
 sg13g2_fill_1 FILLER_48_402 ();
 sg13g2_fill_2 FILLER_48_408 ();
 sg13g2_fill_1 FILLER_48_410 ();
 sg13g2_decap_8 FILLER_48_415 ();
 sg13g2_fill_1 FILLER_48_422 ();
 sg13g2_fill_2 FILLER_48_428 ();
 sg13g2_decap_8 FILLER_49_0 ();
 sg13g2_decap_4 FILLER_49_7 ();
 sg13g2_fill_1 FILLER_49_11 ();
 sg13g2_fill_1 FILLER_49_31 ();
 sg13g2_fill_1 FILLER_49_42 ();
 sg13g2_fill_1 FILLER_49_63 ();
 sg13g2_fill_1 FILLER_49_69 ();
 sg13g2_fill_2 FILLER_49_75 ();
 sg13g2_fill_1 FILLER_49_102 ();
 sg13g2_fill_1 FILLER_49_108 ();
 sg13g2_fill_1 FILLER_49_119 ();
 sg13g2_fill_1 FILLER_49_130 ();
 sg13g2_fill_2 FILLER_49_135 ();
 sg13g2_fill_1 FILLER_49_142 ();
 sg13g2_fill_2 FILLER_49_157 ();
 sg13g2_fill_1 FILLER_49_159 ();
 sg13g2_fill_2 FILLER_49_192 ();
 sg13g2_fill_2 FILLER_49_199 ();
 sg13g2_fill_1 FILLER_49_201 ();
 sg13g2_fill_2 FILLER_49_207 ();
 sg13g2_fill_1 FILLER_49_209 ();
 sg13g2_fill_2 FILLER_49_236 ();
 sg13g2_fill_1 FILLER_49_238 ();
 sg13g2_fill_2 FILLER_49_244 ();
 sg13g2_fill_1 FILLER_49_246 ();
 sg13g2_fill_2 FILLER_49_252 ();
 sg13g2_decap_4 FILLER_49_261 ();
 sg13g2_fill_1 FILLER_49_265 ();
 sg13g2_decap_4 FILLER_49_270 ();
 sg13g2_fill_1 FILLER_49_279 ();
 sg13g2_fill_1 FILLER_49_297 ();
 sg13g2_fill_1 FILLER_49_340 ();
 sg13g2_fill_2 FILLER_49_366 ();
 sg13g2_fill_1 FILLER_49_368 ();
 sg13g2_decap_8 FILLER_50_0 ();
 sg13g2_decap_8 FILLER_50_7 ();
 sg13g2_decap_8 FILLER_50_14 ();
 sg13g2_fill_2 FILLER_50_21 ();
 sg13g2_decap_8 FILLER_50_31 ();
 sg13g2_decap_8 FILLER_50_53 ();
 sg13g2_fill_2 FILLER_50_60 ();
 sg13g2_fill_1 FILLER_50_62 ();
 sg13g2_fill_2 FILLER_50_111 ();
 sg13g2_decap_4 FILLER_50_117 ();
 sg13g2_fill_1 FILLER_50_126 ();
 sg13g2_fill_1 FILLER_50_153 ();
 sg13g2_fill_2 FILLER_50_157 ();
 sg13g2_fill_1 FILLER_50_164 ();
 sg13g2_fill_1 FILLER_50_170 ();
 sg13g2_decap_4 FILLER_50_176 ();
 sg13g2_fill_2 FILLER_50_180 ();
 sg13g2_fill_1 FILLER_50_218 ();
 sg13g2_fill_1 FILLER_50_254 ();
 sg13g2_fill_2 FILLER_50_338 ();
 sg13g2_fill_1 FILLER_50_340 ();
 sg13g2_decap_4 FILLER_50_351 ();
 sg13g2_fill_1 FILLER_50_355 ();
 sg13g2_fill_2 FILLER_50_366 ();
 sg13g2_fill_1 FILLER_50_372 ();
 sg13g2_fill_1 FILLER_50_377 ();
 sg13g2_fill_1 FILLER_50_382 ();
 sg13g2_fill_2 FILLER_50_402 ();
 sg13g2_decap_8 FILLER_51_0 ();
 sg13g2_decap_4 FILLER_51_7 ();
 sg13g2_fill_2 FILLER_51_11 ();
 sg13g2_fill_2 FILLER_51_39 ();
 sg13g2_fill_1 FILLER_51_71 ();
 sg13g2_decap_4 FILLER_51_139 ();
 sg13g2_fill_1 FILLER_51_143 ();
 sg13g2_fill_2 FILLER_51_227 ();
 sg13g2_fill_1 FILLER_51_233 ();
 sg13g2_decap_4 FILLER_51_239 ();
 sg13g2_fill_1 FILLER_51_243 ();
 sg13g2_fill_1 FILLER_51_282 ();
 sg13g2_fill_1 FILLER_51_287 ();
 sg13g2_fill_1 FILLER_51_293 ();
 sg13g2_fill_1 FILLER_51_299 ();
 sg13g2_fill_2 FILLER_51_304 ();
 sg13g2_fill_2 FILLER_51_310 ();
 sg13g2_fill_2 FILLER_51_316 ();
 sg13g2_decap_8 FILLER_51_322 ();
 sg13g2_fill_1 FILLER_51_329 ();
 sg13g2_fill_2 FILLER_51_335 ();
 sg13g2_fill_2 FILLER_51_350 ();
 sg13g2_decap_4 FILLER_51_366 ();
 sg13g2_fill_2 FILLER_51_370 ();
 sg13g2_decap_8 FILLER_51_376 ();
 sg13g2_decap_8 FILLER_51_383 ();
 sg13g2_decap_4 FILLER_51_390 ();
 sg13g2_decap_8 FILLER_52_0 ();
 sg13g2_decap_8 FILLER_52_7 ();
 sg13g2_decap_4 FILLER_52_14 ();
 sg13g2_fill_2 FILLER_52_18 ();
 sg13g2_fill_1 FILLER_52_25 ();
 sg13g2_fill_1 FILLER_52_52 ();
 sg13g2_fill_1 FILLER_52_57 ();
 sg13g2_fill_1 FILLER_52_105 ();
 sg13g2_fill_1 FILLER_52_132 ();
 sg13g2_fill_1 FILLER_52_137 ();
 sg13g2_fill_1 FILLER_52_165 ();
 sg13g2_fill_2 FILLER_52_169 ();
 sg13g2_fill_2 FILLER_52_176 ();
 sg13g2_fill_2 FILLER_52_184 ();
 sg13g2_fill_1 FILLER_52_200 ();
 sg13g2_fill_2 FILLER_52_211 ();
 sg13g2_fill_1 FILLER_52_213 ();
 sg13g2_fill_2 FILLER_52_224 ();
 sg13g2_fill_2 FILLER_52_230 ();
 sg13g2_fill_1 FILLER_52_290 ();
 sg13g2_decap_8 FILLER_52_295 ();
 sg13g2_fill_2 FILLER_52_337 ();
 sg13g2_fill_1 FILLER_52_339 ();
 sg13g2_fill_2 FILLER_52_396 ();
 sg13g2_fill_1 FILLER_52_398 ();
 sg13g2_fill_1 FILLER_52_404 ();
 sg13g2_fill_2 FILLER_52_409 ();
 sg13g2_fill_1 FILLER_52_429 ();
 sg13g2_decap_8 FILLER_53_0 ();
 sg13g2_fill_2 FILLER_53_7 ();
 sg13g2_decap_4 FILLER_53_17 ();
 sg13g2_fill_1 FILLER_53_35 ();
 sg13g2_fill_1 FILLER_53_40 ();
 sg13g2_fill_1 FILLER_53_45 ();
 sg13g2_fill_2 FILLER_53_61 ();
 sg13g2_fill_1 FILLER_53_68 ();
 sg13g2_fill_1 FILLER_53_73 ();
 sg13g2_fill_1 FILLER_53_104 ();
 sg13g2_fill_2 FILLER_53_110 ();
 sg13g2_fill_2 FILLER_53_144 ();
 sg13g2_fill_2 FILLER_53_169 ();
 sg13g2_fill_1 FILLER_53_179 ();
 sg13g2_fill_2 FILLER_53_184 ();
 sg13g2_decap_8 FILLER_53_191 ();
 sg13g2_decap_4 FILLER_53_198 ();
 sg13g2_decap_8 FILLER_53_282 ();
 sg13g2_decap_4 FILLER_53_289 ();
 sg13g2_fill_2 FILLER_53_293 ();
 sg13g2_fill_1 FILLER_53_300 ();
 sg13g2_fill_2 FILLER_53_309 ();
 sg13g2_fill_2 FILLER_53_335 ();
 sg13g2_fill_2 FILLER_53_359 ();
 sg13g2_fill_2 FILLER_53_370 ();
 sg13g2_decap_4 FILLER_53_410 ();
 sg13g2_fill_2 FILLER_53_414 ();
 sg13g2_decap_4 FILLER_54_0 ();
 sg13g2_fill_2 FILLER_54_4 ();
 sg13g2_fill_1 FILLER_54_32 ();
 sg13g2_decap_4 FILLER_54_47 ();
 sg13g2_fill_2 FILLER_54_51 ();
 sg13g2_fill_1 FILLER_54_58 ();
 sg13g2_fill_1 FILLER_54_64 ();
 sg13g2_fill_1 FILLER_54_69 ();
 sg13g2_fill_1 FILLER_54_75 ();
 sg13g2_decap_8 FILLER_54_94 ();
 sg13g2_decap_4 FILLER_54_101 ();
 sg13g2_fill_2 FILLER_54_127 ();
 sg13g2_fill_1 FILLER_54_129 ();
 sg13g2_fill_1 FILLER_54_135 ();
 sg13g2_fill_1 FILLER_54_140 ();
 sg13g2_fill_1 FILLER_54_162 ();
 sg13g2_fill_1 FILLER_54_167 ();
 sg13g2_fill_1 FILLER_54_212 ();
 sg13g2_fill_2 FILLER_54_218 ();
 sg13g2_fill_1 FILLER_54_225 ();
 sg13g2_fill_2 FILLER_54_230 ();
 sg13g2_fill_2 FILLER_54_244 ();
 sg13g2_fill_1 FILLER_54_251 ();
 sg13g2_fill_1 FILLER_54_296 ();
 sg13g2_fill_2 FILLER_54_302 ();
 sg13g2_fill_1 FILLER_54_304 ();
 sg13g2_fill_2 FILLER_54_318 ();
 sg13g2_decap_4 FILLER_54_338 ();
 sg13g2_fill_2 FILLER_54_342 ();
 sg13g2_fill_2 FILLER_54_391 ();
 sg13g2_fill_1 FILLER_54_422 ();
 sg13g2_fill_2 FILLER_54_428 ();
 sg13g2_decap_8 FILLER_55_0 ();
 sg13g2_decap_8 FILLER_55_7 ();
 sg13g2_decap_8 FILLER_55_14 ();
 sg13g2_decap_8 FILLER_55_21 ();
 sg13g2_fill_2 FILLER_55_28 ();
 sg13g2_decap_8 FILLER_55_35 ();
 sg13g2_decap_4 FILLER_55_42 ();
 sg13g2_fill_2 FILLER_55_56 ();
 sg13g2_decap_8 FILLER_55_64 ();
 sg13g2_fill_2 FILLER_55_71 ();
 sg13g2_fill_1 FILLER_55_73 ();
 sg13g2_decap_8 FILLER_55_78 ();
 sg13g2_decap_4 FILLER_55_85 ();
 sg13g2_fill_1 FILLER_55_89 ();
 sg13g2_fill_1 FILLER_55_105 ();
 sg13g2_fill_1 FILLER_55_110 ();
 sg13g2_fill_1 FILLER_55_115 ();
 sg13g2_fill_1 FILLER_55_121 ();
 sg13g2_fill_2 FILLER_55_126 ();
 sg13g2_fill_2 FILLER_55_141 ();
 sg13g2_fill_1 FILLER_55_143 ();
 sg13g2_fill_2 FILLER_55_149 ();
 sg13g2_fill_1 FILLER_55_151 ();
 sg13g2_fill_1 FILLER_55_156 ();
 sg13g2_decap_8 FILLER_55_161 ();
 sg13g2_fill_1 FILLER_55_168 ();
 sg13g2_fill_2 FILLER_55_255 ();
 sg13g2_fill_1 FILLER_55_261 ();
 sg13g2_fill_1 FILLER_55_267 ();
 sg13g2_fill_1 FILLER_55_290 ();
 sg13g2_fill_2 FILLER_55_296 ();
 sg13g2_fill_2 FILLER_55_308 ();
 sg13g2_fill_2 FILLER_55_314 ();
 sg13g2_fill_1 FILLER_55_316 ();
 sg13g2_fill_1 FILLER_55_322 ();
 sg13g2_fill_1 FILLER_55_386 ();
 sg13g2_fill_2 FILLER_55_427 ();
 sg13g2_fill_1 FILLER_55_429 ();
 sg13g2_decap_8 FILLER_56_0 ();
 sg13g2_fill_2 FILLER_56_7 ();
 sg13g2_fill_1 FILLER_56_40 ();
 sg13g2_fill_2 FILLER_56_72 ();
 sg13g2_fill_1 FILLER_56_74 ();
 sg13g2_fill_1 FILLER_56_106 ();
 sg13g2_decap_4 FILLER_56_194 ();
 sg13g2_fill_1 FILLER_56_198 ();
 sg13g2_fill_2 FILLER_56_214 ();
 sg13g2_fill_1 FILLER_56_216 ();
 sg13g2_fill_2 FILLER_56_248 ();
 sg13g2_fill_1 FILLER_56_286 ();
 sg13g2_fill_2 FILLER_56_313 ();
 sg13g2_fill_1 FILLER_56_315 ();
 sg13g2_fill_2 FILLER_56_335 ();
 sg13g2_fill_1 FILLER_56_347 ();
 sg13g2_fill_1 FILLER_56_353 ();
 sg13g2_fill_1 FILLER_56_358 ();
 sg13g2_fill_1 FILLER_56_364 ();
 sg13g2_fill_1 FILLER_56_370 ();
 sg13g2_fill_1 FILLER_56_375 ();
 sg13g2_fill_2 FILLER_56_381 ();
 sg13g2_fill_1 FILLER_56_424 ();
 sg13g2_decap_8 FILLER_57_0 ();
 sg13g2_fill_2 FILLER_57_7 ();
 sg13g2_fill_2 FILLER_57_75 ();
 sg13g2_fill_1 FILLER_57_183 ();
 sg13g2_fill_2 FILLER_57_234 ();
 sg13g2_fill_1 FILLER_57_248 ();
 sg13g2_fill_2 FILLER_57_283 ();
 sg13g2_fill_2 FILLER_57_289 ();
 sg13g2_fill_1 FILLER_57_291 ();
 sg13g2_fill_2 FILLER_57_296 ();
 sg13g2_fill_1 FILLER_57_298 ();
 sg13g2_fill_2 FILLER_57_303 ();
 sg13g2_fill_2 FILLER_57_315 ();
 sg13g2_fill_2 FILLER_57_332 ();
 sg13g2_fill_2 FILLER_57_362 ();
 sg13g2_fill_2 FILLER_57_394 ();
 sg13g2_fill_1 FILLER_57_423 ();
 sg13g2_fill_1 FILLER_57_429 ();
 sg13g2_decap_8 FILLER_58_0 ();
 sg13g2_decap_8 FILLER_58_7 ();
 sg13g2_decap_8 FILLER_58_14 ();
 sg13g2_fill_1 FILLER_58_21 ();
 sg13g2_fill_1 FILLER_58_31 ();
 sg13g2_fill_2 FILLER_58_104 ();
 sg13g2_fill_1 FILLER_58_156 ();
 sg13g2_fill_2 FILLER_58_172 ();
 sg13g2_fill_1 FILLER_58_186 ();
 sg13g2_fill_1 FILLER_58_192 ();
 sg13g2_fill_1 FILLER_58_198 ();
 sg13g2_fill_1 FILLER_58_203 ();
 sg13g2_fill_1 FILLER_58_209 ();
 sg13g2_fill_1 FILLER_58_218 ();
 sg13g2_fill_1 FILLER_58_227 ();
 sg13g2_fill_2 FILLER_58_263 ();
 sg13g2_fill_2 FILLER_58_270 ();
 sg13g2_fill_1 FILLER_58_272 ();
 sg13g2_decap_8 FILLER_58_278 ();
 sg13g2_fill_1 FILLER_58_285 ();
 sg13g2_fill_1 FILLER_58_290 ();
 sg13g2_fill_2 FILLER_58_296 ();
 sg13g2_fill_2 FILLER_58_341 ();
 sg13g2_decap_4 FILLER_58_402 ();
 sg13g2_fill_2 FILLER_58_406 ();
 sg13g2_decap_4 FILLER_58_412 ();
 sg13g2_decap_4 FILLER_58_426 ();
 sg13g2_decap_8 FILLER_59_0 ();
 sg13g2_decap_8 FILLER_59_7 ();
 sg13g2_decap_8 FILLER_59_14 ();
 sg13g2_decap_8 FILLER_59_21 ();
 sg13g2_fill_1 FILLER_59_28 ();
 sg13g2_fill_1 FILLER_59_37 ();
 sg13g2_fill_1 FILLER_59_46 ();
 sg13g2_fill_2 FILLER_59_62 ();
 sg13g2_fill_2 FILLER_59_95 ();
 sg13g2_fill_2 FILLER_59_102 ();
 sg13g2_fill_2 FILLER_59_120 ();
 sg13g2_fill_1 FILLER_59_126 ();
 sg13g2_fill_1 FILLER_59_132 ();
 sg13g2_fill_2 FILLER_59_146 ();
 sg13g2_fill_1 FILLER_59_148 ();
 sg13g2_fill_2 FILLER_59_152 ();
 sg13g2_fill_1 FILLER_59_158 ();
 sg13g2_fill_1 FILLER_59_162 ();
 sg13g2_fill_1 FILLER_59_168 ();
 sg13g2_fill_1 FILLER_59_179 ();
 sg13g2_fill_1 FILLER_59_200 ();
 sg13g2_fill_1 FILLER_59_208 ();
 sg13g2_fill_1 FILLER_59_213 ();
 sg13g2_fill_1 FILLER_59_219 ();
 sg13g2_fill_1 FILLER_59_226 ();
 sg13g2_fill_1 FILLER_59_233 ();
 sg13g2_fill_1 FILLER_59_239 ();
 sg13g2_fill_1 FILLER_59_244 ();
 sg13g2_fill_2 FILLER_59_256 ();
 sg13g2_fill_1 FILLER_59_289 ();
 sg13g2_fill_1 FILLER_59_395 ();
 sg13g2_decap_4 FILLER_59_426 ();
 sg13g2_decap_8 FILLER_60_0 ();
 sg13g2_decap_8 FILLER_60_7 ();
 sg13g2_decap_8 FILLER_60_14 ();
 sg13g2_decap_4 FILLER_60_21 ();
 sg13g2_fill_1 FILLER_60_25 ();
 sg13g2_decap_4 FILLER_60_30 ();
 sg13g2_fill_2 FILLER_60_48 ();
 sg13g2_decap_8 FILLER_60_67 ();
 sg13g2_decap_4 FILLER_60_74 ();
 sg13g2_fill_1 FILLER_60_87 ();
 sg13g2_fill_1 FILLER_60_127 ();
 sg13g2_fill_1 FILLER_60_132 ();
 sg13g2_fill_1 FILLER_60_141 ();
 sg13g2_fill_1 FILLER_60_151 ();
 sg13g2_fill_1 FILLER_60_156 ();
 sg13g2_fill_1 FILLER_60_162 ();
 sg13g2_fill_1 FILLER_60_172 ();
 sg13g2_decap_4 FILLER_60_178 ();
 sg13g2_fill_2 FILLER_60_182 ();
 sg13g2_decap_8 FILLER_60_189 ();
 sg13g2_fill_2 FILLER_60_196 ();
 sg13g2_fill_1 FILLER_60_198 ();
 sg13g2_decap_4 FILLER_60_202 ();
 sg13g2_fill_2 FILLER_60_206 ();
 sg13g2_fill_1 FILLER_60_266 ();
 sg13g2_fill_2 FILLER_60_271 ();
 sg13g2_fill_2 FILLER_60_278 ();
 sg13g2_fill_1 FILLER_60_285 ();
 sg13g2_decap_4 FILLER_60_290 ();
 sg13g2_fill_1 FILLER_60_294 ();
 sg13g2_fill_2 FILLER_60_315 ();
 sg13g2_fill_1 FILLER_60_359 ();
 sg13g2_fill_1 FILLER_60_369 ();
 sg13g2_fill_2 FILLER_60_396 ();
 sg13g2_fill_1 FILLER_60_403 ();
 sg13g2_decap_8 FILLER_61_0 ();
 sg13g2_decap_8 FILLER_61_7 ();
 sg13g2_decap_8 FILLER_61_14 ();
 sg13g2_fill_2 FILLER_61_21 ();
 sg13g2_fill_1 FILLER_61_23 ();
 sg13g2_fill_1 FILLER_61_61 ();
 sg13g2_decap_8 FILLER_61_67 ();
 sg13g2_fill_2 FILLER_61_74 ();
 sg13g2_decap_4 FILLER_61_116 ();
 sg13g2_fill_2 FILLER_61_120 ();
 sg13g2_decap_4 FILLER_61_127 ();
 sg13g2_fill_2 FILLER_61_150 ();
 sg13g2_fill_1 FILLER_61_157 ();
 sg13g2_fill_2 FILLER_61_193 ();
 sg13g2_fill_1 FILLER_61_200 ();
 sg13g2_fill_2 FILLER_61_211 ();
 sg13g2_fill_1 FILLER_61_217 ();
 sg13g2_fill_2 FILLER_61_223 ();
 sg13g2_fill_2 FILLER_61_230 ();
 sg13g2_fill_1 FILLER_61_291 ();
 sg13g2_fill_1 FILLER_61_296 ();
 sg13g2_fill_2 FILLER_61_304 ();
 sg13g2_decap_8 FILLER_61_311 ();
 sg13g2_fill_2 FILLER_61_342 ();
 sg13g2_fill_2 FILLER_61_350 ();
 sg13g2_fill_1 FILLER_61_352 ();
 sg13g2_decap_4 FILLER_61_366 ();
 sg13g2_fill_1 FILLER_61_370 ();
 sg13g2_fill_1 FILLER_61_376 ();
 sg13g2_fill_2 FILLER_61_381 ();
 sg13g2_fill_2 FILLER_61_388 ();
 sg13g2_fill_2 FILLER_61_395 ();
 sg13g2_fill_2 FILLER_61_428 ();
 sg13g2_decap_8 FILLER_62_0 ();
 sg13g2_decap_8 FILLER_62_7 ();
 sg13g2_fill_1 FILLER_62_14 ();
 sg13g2_decap_4 FILLER_62_41 ();
 sg13g2_fill_2 FILLER_62_80 ();
 sg13g2_fill_1 FILLER_62_82 ();
 sg13g2_fill_2 FILLER_62_93 ();
 sg13g2_fill_1 FILLER_62_95 ();
 sg13g2_fill_1 FILLER_62_108 ();
 sg13g2_fill_1 FILLER_62_114 ();
 sg13g2_fill_1 FILLER_62_120 ();
 sg13g2_fill_2 FILLER_62_126 ();
 sg13g2_fill_1 FILLER_62_138 ();
 sg13g2_fill_2 FILLER_62_144 ();
 sg13g2_decap_4 FILLER_62_181 ();
 sg13g2_fill_1 FILLER_62_185 ();
 sg13g2_fill_1 FILLER_62_194 ();
 sg13g2_fill_1 FILLER_62_201 ();
 sg13g2_fill_2 FILLER_62_206 ();
 sg13g2_fill_1 FILLER_62_208 ();
 sg13g2_fill_1 FILLER_62_219 ();
 sg13g2_decap_8 FILLER_62_223 ();
 sg13g2_fill_2 FILLER_62_230 ();
 sg13g2_decap_4 FILLER_62_273 ();
 sg13g2_fill_2 FILLER_62_277 ();
 sg13g2_fill_2 FILLER_62_284 ();
 sg13g2_decap_8 FILLER_62_311 ();
 sg13g2_fill_1 FILLER_62_318 ();
 sg13g2_fill_1 FILLER_62_332 ();
 sg13g2_fill_2 FILLER_62_365 ();
 sg13g2_fill_1 FILLER_62_367 ();
 sg13g2_fill_2 FILLER_62_373 ();
 sg13g2_fill_1 FILLER_62_379 ();
 sg13g2_fill_1 FILLER_62_392 ();
 sg13g2_fill_2 FILLER_62_398 ();
 sg13g2_fill_2 FILLER_62_417 ();
 sg13g2_fill_1 FILLER_62_429 ();
 sg13g2_decap_4 FILLER_63_0 ();
 sg13g2_fill_2 FILLER_63_4 ();
 sg13g2_decap_8 FILLER_63_51 ();
 sg13g2_fill_2 FILLER_63_58 ();
 sg13g2_fill_1 FILLER_63_166 ();
 sg13g2_fill_2 FILLER_63_171 ();
 sg13g2_fill_1 FILLER_63_173 ();
 sg13g2_fill_1 FILLER_63_191 ();
 sg13g2_fill_2 FILLER_63_206 ();
 sg13g2_fill_1 FILLER_63_218 ();
 sg13g2_decap_8 FILLER_63_223 ();
 sg13g2_fill_2 FILLER_63_230 ();
 sg13g2_fill_1 FILLER_63_232 ();
 sg13g2_fill_1 FILLER_63_243 ();
 sg13g2_fill_2 FILLER_63_249 ();
 sg13g2_fill_2 FILLER_63_256 ();
 sg13g2_fill_2 FILLER_63_262 ();
 sg13g2_fill_1 FILLER_63_264 ();
 sg13g2_fill_2 FILLER_63_275 ();
 sg13g2_fill_2 FILLER_63_307 ();
 sg13g2_fill_2 FILLER_63_313 ();
 sg13g2_fill_1 FILLER_63_319 ();
 sg13g2_fill_1 FILLER_63_346 ();
 sg13g2_fill_2 FILLER_63_417 ();
 sg13g2_decap_4 FILLER_63_424 ();
 sg13g2_fill_2 FILLER_63_428 ();
 sg13g2_decap_8 FILLER_64_0 ();
 sg13g2_decap_8 FILLER_64_7 ();
 sg13g2_fill_2 FILLER_64_14 ();
 sg13g2_fill_1 FILLER_64_16 ();
 sg13g2_decap_8 FILLER_64_21 ();
 sg13g2_fill_1 FILLER_64_28 ();
 sg13g2_decap_8 FILLER_64_39 ();
 sg13g2_decap_8 FILLER_64_51 ();
 sg13g2_fill_2 FILLER_64_58 ();
 sg13g2_fill_1 FILLER_64_109 ();
 sg13g2_fill_1 FILLER_64_119 ();
 sg13g2_fill_2 FILLER_64_135 ();
 sg13g2_fill_1 FILLER_64_151 ();
 sg13g2_fill_1 FILLER_64_157 ();
 sg13g2_fill_1 FILLER_64_166 ();
 sg13g2_fill_2 FILLER_64_174 ();
 sg13g2_fill_1 FILLER_64_180 ();
 sg13g2_fill_2 FILLER_64_186 ();
 sg13g2_fill_2 FILLER_64_198 ();
 sg13g2_fill_1 FILLER_64_200 ();
 sg13g2_fill_2 FILLER_64_236 ();
 sg13g2_fill_1 FILLER_64_243 ();
 sg13g2_fill_1 FILLER_64_248 ();
 sg13g2_fill_2 FILLER_64_267 ();
 sg13g2_fill_1 FILLER_64_278 ();
 sg13g2_fill_1 FILLER_64_303 ();
 sg13g2_fill_1 FILLER_64_335 ();
 sg13g2_fill_1 FILLER_64_341 ();
 sg13g2_fill_1 FILLER_64_385 ();
 sg13g2_decap_4 FILLER_64_390 ();
 sg13g2_decap_8 FILLER_65_0 ();
 sg13g2_decap_8 FILLER_65_7 ();
 sg13g2_decap_8 FILLER_65_14 ();
 sg13g2_decap_4 FILLER_65_21 ();
 sg13g2_fill_2 FILLER_65_35 ();
 sg13g2_fill_1 FILLER_65_47 ();
 sg13g2_fill_1 FILLER_65_56 ();
 sg13g2_fill_2 FILLER_65_62 ();
 sg13g2_fill_2 FILLER_65_70 ();
 sg13g2_fill_2 FILLER_65_107 ();
 sg13g2_fill_1 FILLER_65_113 ();
 sg13g2_fill_1 FILLER_65_118 ();
 sg13g2_fill_1 FILLER_65_149 ();
 sg13g2_fill_1 FILLER_65_155 ();
 sg13g2_fill_1 FILLER_65_161 ();
 sg13g2_fill_2 FILLER_65_167 ();
 sg13g2_fill_2 FILLER_65_200 ();
 sg13g2_fill_2 FILLER_65_304 ();
 sg13g2_fill_1 FILLER_65_310 ();
 sg13g2_fill_1 FILLER_65_334 ();
 sg13g2_fill_1 FILLER_65_365 ();
 sg13g2_decap_4 FILLER_65_371 ();
 sg13g2_fill_1 FILLER_65_403 ();
 sg13g2_decap_4 FILLER_66_0 ();
 sg13g2_fill_2 FILLER_66_30 ();
 sg13g2_fill_1 FILLER_66_32 ();
 sg13g2_fill_1 FILLER_66_38 ();
 sg13g2_fill_1 FILLER_66_73 ();
 sg13g2_fill_2 FILLER_66_104 ();
 sg13g2_decap_8 FILLER_66_112 ();
 sg13g2_fill_2 FILLER_66_144 ();
 sg13g2_fill_1 FILLER_66_146 ();
 sg13g2_fill_1 FILLER_66_161 ();
 sg13g2_fill_1 FILLER_66_166 ();
 sg13g2_fill_1 FILLER_66_178 ();
 sg13g2_fill_1 FILLER_66_188 ();
 sg13g2_fill_2 FILLER_66_193 ();
 sg13g2_fill_1 FILLER_66_195 ();
 sg13g2_decap_4 FILLER_66_211 ();
 sg13g2_fill_1 FILLER_66_215 ();
 sg13g2_fill_1 FILLER_66_235 ();
 sg13g2_fill_1 FILLER_66_241 ();
 sg13g2_fill_2 FILLER_66_246 ();
 sg13g2_fill_1 FILLER_66_248 ();
 sg13g2_fill_2 FILLER_66_259 ();
 sg13g2_fill_1 FILLER_66_261 ();
 sg13g2_fill_1 FILLER_66_267 ();
 sg13g2_fill_1 FILLER_66_277 ();
 sg13g2_fill_2 FILLER_66_322 ();
 sg13g2_fill_1 FILLER_66_328 ();
 sg13g2_fill_1 FILLER_66_334 ();
 sg13g2_decap_4 FILLER_66_339 ();
 sg13g2_fill_1 FILLER_66_343 ();
 sg13g2_fill_1 FILLER_66_348 ();
 sg13g2_fill_2 FILLER_66_362 ();
 sg13g2_decap_4 FILLER_66_369 ();
 sg13g2_fill_1 FILLER_66_398 ();
 sg13g2_decap_8 FILLER_67_0 ();
 sg13g2_fill_2 FILLER_67_7 ();
 sg13g2_fill_1 FILLER_67_9 ();
 sg13g2_fill_1 FILLER_67_65 ();
 sg13g2_fill_1 FILLER_67_76 ();
 sg13g2_fill_2 FILLER_67_82 ();
 sg13g2_fill_1 FILLER_67_94 ();
 sg13g2_fill_1 FILLER_67_121 ();
 sg13g2_fill_1 FILLER_67_128 ();
 sg13g2_fill_1 FILLER_67_160 ();
 sg13g2_fill_1 FILLER_67_165 ();
 sg13g2_fill_1 FILLER_67_169 ();
 sg13g2_fill_1 FILLER_67_177 ();
 sg13g2_fill_1 FILLER_67_182 ();
 sg13g2_fill_1 FILLER_67_188 ();
 sg13g2_fill_1 FILLER_67_194 ();
 sg13g2_fill_2 FILLER_67_200 ();
 sg13g2_fill_2 FILLER_67_207 ();
 sg13g2_fill_2 FILLER_67_219 ();
 sg13g2_fill_2 FILLER_67_295 ();
 sg13g2_fill_2 FILLER_67_301 ();
 sg13g2_fill_1 FILLER_67_303 ();
 sg13g2_fill_2 FILLER_67_334 ();
 sg13g2_fill_1 FILLER_67_336 ();
 sg13g2_decap_4 FILLER_67_347 ();
 sg13g2_fill_1 FILLER_67_351 ();
 sg13g2_decap_4 FILLER_67_356 ();
 sg13g2_fill_2 FILLER_67_360 ();
 sg13g2_fill_1 FILLER_67_372 ();
 sg13g2_fill_1 FILLER_67_377 ();
 sg13g2_fill_1 FILLER_67_388 ();
 sg13g2_fill_2 FILLER_67_422 ();
 sg13g2_fill_2 FILLER_67_428 ();
 sg13g2_decap_8 FILLER_68_0 ();
 sg13g2_decap_8 FILLER_68_7 ();
 sg13g2_fill_2 FILLER_68_14 ();
 sg13g2_fill_1 FILLER_68_16 ();
 sg13g2_fill_2 FILLER_68_39 ();
 sg13g2_fill_2 FILLER_68_51 ();
 sg13g2_fill_1 FILLER_68_112 ();
 sg13g2_fill_2 FILLER_68_169 ();
 sg13g2_decap_8 FILLER_68_285 ();
 sg13g2_fill_1 FILLER_68_292 ();
 sg13g2_fill_1 FILLER_68_298 ();
 sg13g2_fill_1 FILLER_68_309 ();
 sg13g2_fill_1 FILLER_68_320 ();
 sg13g2_fill_2 FILLER_68_326 ();
 sg13g2_fill_2 FILLER_68_354 ();
 sg13g2_fill_1 FILLER_68_401 ();
 sg13g2_fill_1 FILLER_68_412 ();
 sg13g2_fill_2 FILLER_68_417 ();
 sg13g2_fill_1 FILLER_68_419 ();
 sg13g2_decap_4 FILLER_68_425 ();
 sg13g2_fill_1 FILLER_68_429 ();
 sg13g2_decap_8 FILLER_69_0 ();
 sg13g2_decap_8 FILLER_69_7 ();
 sg13g2_decap_8 FILLER_69_14 ();
 sg13g2_decap_8 FILLER_69_21 ();
 sg13g2_decap_8 FILLER_69_28 ();
 sg13g2_fill_2 FILLER_69_35 ();
 sg13g2_fill_2 FILLER_69_93 ();
 sg13g2_decap_8 FILLER_69_100 ();
 sg13g2_fill_1 FILLER_69_107 ();
 sg13g2_fill_1 FILLER_69_142 ();
 sg13g2_fill_1 FILLER_69_158 ();
 sg13g2_fill_1 FILLER_69_173 ();
 sg13g2_decap_4 FILLER_69_223 ();
 sg13g2_fill_2 FILLER_69_227 ();
 sg13g2_decap_4 FILLER_69_233 ();
 sg13g2_fill_1 FILLER_69_237 ();
 sg13g2_fill_2 FILLER_69_272 ();
 sg13g2_fill_1 FILLER_69_300 ();
 sg13g2_fill_1 FILLER_69_327 ();
 sg13g2_fill_1 FILLER_69_386 ();
 sg13g2_fill_1 FILLER_69_397 ();
 sg13g2_fill_1 FILLER_69_403 ();
 sg13g2_decap_8 FILLER_70_0 ();
 sg13g2_decap_8 FILLER_70_7 ();
 sg13g2_decap_8 FILLER_70_14 ();
 sg13g2_decap_8 FILLER_70_21 ();
 sg13g2_decap_8 FILLER_70_28 ();
 sg13g2_fill_2 FILLER_70_35 ();
 sg13g2_decap_4 FILLER_70_47 ();
 sg13g2_fill_2 FILLER_70_60 ();
 sg13g2_fill_2 FILLER_70_66 ();
 sg13g2_fill_1 FILLER_70_68 ();
 sg13g2_fill_2 FILLER_70_73 ();
 sg13g2_fill_1 FILLER_70_75 ();
 sg13g2_fill_2 FILLER_70_80 ();
 sg13g2_fill_1 FILLER_70_82 ();
 sg13g2_fill_1 FILLER_70_92 ();
 sg13g2_fill_1 FILLER_70_98 ();
 sg13g2_fill_1 FILLER_70_145 ();
 sg13g2_fill_2 FILLER_70_158 ();
 sg13g2_fill_1 FILLER_70_181 ();
 sg13g2_fill_1 FILLER_70_189 ();
 sg13g2_fill_1 FILLER_70_194 ();
 sg13g2_fill_1 FILLER_70_201 ();
 sg13g2_fill_2 FILLER_70_206 ();
 sg13g2_fill_1 FILLER_70_208 ();
 sg13g2_fill_2 FILLER_70_240 ();
 sg13g2_fill_1 FILLER_70_242 ();
 sg13g2_fill_2 FILLER_70_263 ();
 sg13g2_fill_1 FILLER_70_316 ();
 sg13g2_fill_2 FILLER_70_332 ();
 sg13g2_fill_2 FILLER_70_339 ();
 sg13g2_fill_1 FILLER_70_345 ();
 sg13g2_fill_2 FILLER_70_351 ();
 sg13g2_fill_2 FILLER_70_359 ();
 sg13g2_fill_1 FILLER_70_361 ();
 sg13g2_fill_2 FILLER_70_366 ();
 sg13g2_fill_2 FILLER_70_372 ();
 sg13g2_fill_1 FILLER_70_374 ();
 sg13g2_fill_1 FILLER_70_380 ();
 sg13g2_fill_2 FILLER_70_386 ();
 sg13g2_fill_1 FILLER_70_388 ();
 sg13g2_decap_8 FILLER_71_0 ();
 sg13g2_decap_8 FILLER_71_7 ();
 sg13g2_decap_8 FILLER_71_14 ();
 sg13g2_decap_8 FILLER_71_21 ();
 sg13g2_decap_8 FILLER_71_28 ();
 sg13g2_decap_8 FILLER_71_35 ();
 sg13g2_fill_2 FILLER_71_42 ();
 sg13g2_fill_1 FILLER_71_93 ();
 sg13g2_fill_1 FILLER_71_107 ();
 sg13g2_fill_1 FILLER_71_112 ();
 sg13g2_fill_1 FILLER_71_123 ();
 sg13g2_fill_2 FILLER_71_134 ();
 sg13g2_fill_2 FILLER_71_189 ();
 sg13g2_decap_8 FILLER_71_195 ();
 sg13g2_fill_2 FILLER_71_202 ();
 sg13g2_fill_1 FILLER_71_209 ();
 sg13g2_decap_8 FILLER_71_215 ();
 sg13g2_fill_1 FILLER_71_222 ();
 sg13g2_decap_4 FILLER_71_227 ();
 sg13g2_fill_2 FILLER_71_231 ();
 sg13g2_decap_8 FILLER_71_238 ();
 sg13g2_decap_4 FILLER_71_245 ();
 sg13g2_fill_2 FILLER_71_249 ();
 sg13g2_fill_2 FILLER_71_261 ();
 sg13g2_fill_1 FILLER_71_263 ();
 sg13g2_fill_1 FILLER_71_287 ();
 sg13g2_fill_1 FILLER_71_292 ();
 sg13g2_fill_1 FILLER_71_297 ();
 sg13g2_fill_1 FILLER_71_303 ();
 sg13g2_fill_1 FILLER_71_309 ();
 sg13g2_fill_1 FILLER_71_325 ();
 sg13g2_fill_2 FILLER_71_351 ();
 sg13g2_fill_2 FILLER_71_363 ();
 sg13g2_fill_1 FILLER_71_365 ();
 sg13g2_fill_1 FILLER_71_376 ();
 sg13g2_fill_1 FILLER_71_381 ();
 sg13g2_fill_1 FILLER_71_392 ();
 sg13g2_fill_2 FILLER_71_402 ();
 sg13g2_decap_8 FILLER_72_0 ();
 sg13g2_decap_8 FILLER_72_7 ();
 sg13g2_decap_8 FILLER_72_14 ();
 sg13g2_decap_8 FILLER_72_21 ();
 sg13g2_decap_4 FILLER_72_28 ();
 sg13g2_fill_1 FILLER_72_58 ();
 sg13g2_fill_1 FILLER_72_90 ();
 sg13g2_fill_2 FILLER_72_101 ();
 sg13g2_fill_1 FILLER_72_113 ();
 sg13g2_fill_2 FILLER_72_118 ();
 sg13g2_fill_2 FILLER_72_124 ();
 sg13g2_decap_4 FILLER_72_159 ();
 sg13g2_decap_8 FILLER_72_166 ();
 sg13g2_fill_2 FILLER_72_177 ();
 sg13g2_fill_1 FILLER_72_219 ();
 sg13g2_fill_2 FILLER_72_269 ();
 sg13g2_fill_1 FILLER_72_317 ();
 sg13g2_fill_1 FILLER_72_344 ();
 sg13g2_fill_1 FILLER_72_375 ();
 sg13g2_fill_1 FILLER_72_381 ();
 sg13g2_fill_1 FILLER_72_412 ();
 sg13g2_fill_1 FILLER_72_417 ();
 sg13g2_fill_2 FILLER_72_422 ();
 sg13g2_fill_2 FILLER_72_428 ();
 sg13g2_decap_8 FILLER_73_0 ();
 sg13g2_decap_8 FILLER_73_7 ();
 sg13g2_decap_8 FILLER_73_14 ();
 sg13g2_decap_8 FILLER_73_21 ();
 sg13g2_decap_8 FILLER_73_28 ();
 sg13g2_fill_1 FILLER_73_35 ();
 sg13g2_decap_8 FILLER_73_40 ();
 sg13g2_decap_4 FILLER_73_47 ();
 sg13g2_fill_1 FILLER_73_55 ();
 sg13g2_fill_2 FILLER_73_86 ();
 sg13g2_fill_1 FILLER_73_96 ();
 sg13g2_fill_2 FILLER_73_107 ();
 sg13g2_decap_8 FILLER_73_113 ();
 sg13g2_decap_8 FILLER_73_120 ();
 sg13g2_fill_2 FILLER_73_127 ();
 sg13g2_decap_4 FILLER_73_160 ();
 sg13g2_fill_1 FILLER_73_164 ();
 sg13g2_fill_1 FILLER_73_169 ();
 sg13g2_fill_1 FILLER_73_175 ();
 sg13g2_fill_1 FILLER_73_211 ();
 sg13g2_fill_1 FILLER_73_303 ();
 sg13g2_fill_2 FILLER_73_314 ();
 sg13g2_fill_1 FILLER_73_316 ();
 sg13g2_fill_2 FILLER_73_332 ();
 sg13g2_fill_1 FILLER_73_334 ();
 sg13g2_fill_1 FILLER_73_413 ();
 sg13g2_fill_1 FILLER_73_423 ();
 sg13g2_fill_1 FILLER_73_429 ();
 sg13g2_decap_8 FILLER_74_0 ();
 sg13g2_decap_8 FILLER_74_7 ();
 sg13g2_decap_8 FILLER_74_14 ();
 sg13g2_decap_8 FILLER_74_21 ();
 sg13g2_decap_8 FILLER_74_28 ();
 sg13g2_decap_8 FILLER_74_35 ();
 sg13g2_decap_8 FILLER_74_42 ();
 sg13g2_decap_8 FILLER_74_49 ();
 sg13g2_decap_4 FILLER_74_56 ();
 sg13g2_fill_1 FILLER_74_60 ();
 sg13g2_fill_1 FILLER_74_74 ();
 sg13g2_fill_1 FILLER_74_116 ();
 sg13g2_fill_1 FILLER_74_143 ();
 sg13g2_fill_2 FILLER_74_149 ();
 sg13g2_fill_2 FILLER_74_155 ();
 sg13g2_fill_2 FILLER_74_162 ();
 sg13g2_fill_1 FILLER_74_164 ();
 sg13g2_fill_2 FILLER_74_170 ();
 sg13g2_fill_1 FILLER_74_172 ();
 sg13g2_fill_2 FILLER_74_177 ();
 sg13g2_fill_1 FILLER_74_179 ();
 sg13g2_fill_2 FILLER_74_195 ();
 sg13g2_fill_2 FILLER_74_202 ();
 sg13g2_fill_1 FILLER_74_204 ();
 sg13g2_decap_4 FILLER_74_210 ();
 sg13g2_decap_4 FILLER_74_219 ();
 sg13g2_fill_2 FILLER_74_223 ();
 sg13g2_decap_4 FILLER_74_240 ();
 sg13g2_fill_1 FILLER_74_244 ();
 sg13g2_fill_1 FILLER_74_278 ();
 sg13g2_fill_1 FILLER_74_336 ();
 sg13g2_fill_2 FILLER_74_341 ();
 sg13g2_fill_2 FILLER_74_387 ();
 sg13g2_fill_2 FILLER_74_393 ();
 sg13g2_fill_2 FILLER_74_403 ();
 sg13g2_decap_8 FILLER_75_0 ();
 sg13g2_decap_8 FILLER_75_7 ();
 sg13g2_decap_8 FILLER_75_14 ();
 sg13g2_decap_8 FILLER_75_21 ();
 sg13g2_decap_8 FILLER_75_28 ();
 sg13g2_decap_8 FILLER_75_35 ();
 sg13g2_decap_8 FILLER_75_42 ();
 sg13g2_decap_8 FILLER_75_49 ();
 sg13g2_decap_4 FILLER_75_56 ();
 sg13g2_fill_1 FILLER_75_60 ();
 sg13g2_decap_4 FILLER_75_65 ();
 sg13g2_fill_2 FILLER_75_69 ();
 sg13g2_fill_1 FILLER_75_85 ();
 sg13g2_fill_1 FILLER_75_91 ();
 sg13g2_fill_1 FILLER_75_112 ();
 sg13g2_fill_2 FILLER_75_119 ();
 sg13g2_fill_1 FILLER_75_126 ();
 sg13g2_fill_2 FILLER_75_131 ();
 sg13g2_fill_1 FILLER_75_137 ();
 sg13g2_fill_2 FILLER_75_164 ();
 sg13g2_fill_1 FILLER_75_180 ();
 sg13g2_fill_1 FILLER_75_186 ();
 sg13g2_fill_1 FILLER_75_196 ();
 sg13g2_fill_1 FILLER_75_202 ();
 sg13g2_decap_8 FILLER_75_207 ();
 sg13g2_fill_2 FILLER_75_214 ();
 sg13g2_fill_1 FILLER_75_216 ();
 sg13g2_fill_1 FILLER_75_232 ();
 sg13g2_fill_2 FILLER_75_243 ();
 sg13g2_fill_2 FILLER_75_255 ();
 sg13g2_fill_1 FILLER_75_257 ();
 sg13g2_fill_1 FILLER_75_292 ();
 sg13g2_fill_2 FILLER_75_297 ();
 sg13g2_fill_2 FILLER_75_304 ();
 sg13g2_fill_2 FILLER_75_310 ();
 sg13g2_fill_2 FILLER_75_341 ();
 sg13g2_fill_1 FILLER_75_348 ();
 sg13g2_fill_1 FILLER_75_354 ();
 sg13g2_fill_1 FILLER_75_365 ();
 sg13g2_fill_1 FILLER_75_376 ();
 sg13g2_fill_1 FILLER_75_429 ();
 sg13g2_decap_8 FILLER_76_0 ();
 sg13g2_decap_8 FILLER_76_7 ();
 sg13g2_decap_8 FILLER_76_14 ();
 sg13g2_decap_8 FILLER_76_21 ();
 sg13g2_decap_8 FILLER_76_28 ();
 sg13g2_decap_8 FILLER_76_35 ();
 sg13g2_decap_8 FILLER_76_42 ();
 sg13g2_decap_8 FILLER_76_49 ();
 sg13g2_fill_1 FILLER_76_56 ();
 sg13g2_fill_2 FILLER_76_83 ();
 sg13g2_fill_2 FILLER_76_99 ();
 sg13g2_decap_8 FILLER_76_129 ();
 sg13g2_fill_2 FILLER_76_136 ();
 sg13g2_fill_1 FILLER_76_138 ();
 sg13g2_fill_1 FILLER_76_191 ();
 sg13g2_fill_2 FILLER_76_214 ();
 sg13g2_fill_2 FILLER_76_226 ();
 sg13g2_fill_1 FILLER_76_240 ();
 sg13g2_fill_1 FILLER_76_245 ();
 sg13g2_fill_1 FILLER_76_256 ();
 sg13g2_fill_2 FILLER_76_276 ();
 sg13g2_decap_4 FILLER_76_291 ();
 sg13g2_fill_1 FILLER_76_317 ();
 sg13g2_fill_1 FILLER_76_333 ();
 sg13g2_fill_1 FILLER_76_356 ();
 sg13g2_fill_2 FILLER_76_366 ();
 sg13g2_fill_2 FILLER_76_393 ();
 sg13g2_decap_8 FILLER_77_0 ();
 sg13g2_decap_8 FILLER_77_7 ();
 sg13g2_decap_8 FILLER_77_14 ();
 sg13g2_decap_8 FILLER_77_21 ();
 sg13g2_decap_8 FILLER_77_28 ();
 sg13g2_decap_8 FILLER_77_35 ();
 sg13g2_decap_8 FILLER_77_42 ();
 sg13g2_decap_8 FILLER_77_49 ();
 sg13g2_decap_4 FILLER_77_56 ();
 sg13g2_fill_1 FILLER_77_60 ();
 sg13g2_decap_8 FILLER_77_65 ();
 sg13g2_decap_8 FILLER_77_72 ();
 sg13g2_fill_2 FILLER_77_79 ();
 sg13g2_fill_1 FILLER_77_81 ();
 sg13g2_fill_1 FILLER_77_115 ();
 sg13g2_fill_1 FILLER_77_183 ();
 sg13g2_fill_1 FILLER_77_194 ();
 sg13g2_fill_1 FILLER_77_209 ();
 sg13g2_fill_2 FILLER_77_259 ();
 sg13g2_fill_2 FILLER_77_287 ();
 sg13g2_fill_1 FILLER_77_310 ();
 sg13g2_fill_1 FILLER_77_364 ();
 sg13g2_fill_2 FILLER_77_399 ();
 sg13g2_fill_1 FILLER_77_421 ();
 sg13g2_fill_1 FILLER_77_429 ();
 sg13g2_decap_8 FILLER_78_0 ();
 sg13g2_decap_8 FILLER_78_7 ();
 sg13g2_decap_8 FILLER_78_14 ();
 sg13g2_decap_8 FILLER_78_21 ();
 sg13g2_decap_8 FILLER_78_28 ();
 sg13g2_decap_8 FILLER_78_35 ();
 sg13g2_decap_8 FILLER_78_42 ();
 sg13g2_decap_8 FILLER_78_49 ();
 sg13g2_decap_8 FILLER_78_56 ();
 sg13g2_decap_8 FILLER_78_63 ();
 sg13g2_fill_2 FILLER_78_70 ();
 sg13g2_decap_4 FILLER_78_80 ();
 sg13g2_fill_1 FILLER_78_149 ();
 sg13g2_fill_2 FILLER_78_241 ();
 sg13g2_fill_1 FILLER_78_309 ();
 sg13g2_fill_2 FILLER_78_318 ();
 sg13g2_fill_2 FILLER_78_428 ();
 sg13g2_decap_8 FILLER_79_0 ();
 sg13g2_decap_8 FILLER_79_7 ();
 sg13g2_decap_8 FILLER_79_14 ();
 sg13g2_decap_8 FILLER_79_21 ();
 sg13g2_decap_8 FILLER_79_28 ();
 sg13g2_decap_8 FILLER_79_35 ();
 sg13g2_decap_8 FILLER_79_42 ();
 sg13g2_decap_8 FILLER_79_49 ();
 sg13g2_decap_8 FILLER_79_56 ();
 sg13g2_fill_1 FILLER_79_127 ();
 sg13g2_fill_1 FILLER_79_168 ();
 sg13g2_fill_1 FILLER_79_179 ();
 sg13g2_fill_2 FILLER_79_185 ();
 sg13g2_fill_1 FILLER_79_221 ();
 sg13g2_fill_2 FILLER_79_278 ();
 sg13g2_fill_1 FILLER_79_403 ();
 sg13g2_decap_8 FILLER_80_0 ();
 sg13g2_decap_8 FILLER_80_7 ();
 sg13g2_decap_8 FILLER_80_14 ();
 sg13g2_decap_8 FILLER_80_21 ();
 sg13g2_decap_8 FILLER_80_28 ();
 sg13g2_decap_8 FILLER_80_35 ();
 sg13g2_decap_8 FILLER_80_42 ();
 sg13g2_decap_8 FILLER_80_49 ();
 sg13g2_decap_8 FILLER_80_56 ();
 sg13g2_decap_8 FILLER_80_63 ();
 sg13g2_fill_2 FILLER_80_70 ();
 sg13g2_fill_1 FILLER_80_72 ();
 sg13g2_decap_4 FILLER_80_77 ();
 sg13g2_fill_1 FILLER_80_161 ();
 sg13g2_fill_1 FILLER_80_166 ();
 sg13g2_fill_1 FILLER_80_171 ();
 sg13g2_fill_1 FILLER_80_180 ();
 sg13g2_fill_1 FILLER_80_185 ();
 sg13g2_fill_2 FILLER_80_214 ();
 sg13g2_fill_2 FILLER_80_233 ();
 sg13g2_fill_1 FILLER_80_247 ();
 sg13g2_fill_2 FILLER_80_252 ();
 sg13g2_fill_2 FILLER_80_258 ();
 sg13g2_fill_1 FILLER_80_334 ();
 sg13g2_fill_1 FILLER_80_340 ();
 sg13g2_fill_2 FILLER_80_399 ();
 sg13g2_fill_1 FILLER_80_401 ();
 sg13g2_fill_2 FILLER_80_415 ();
endmodule
