module tt_um_edwintorok (clk,
    ena,
    rst_n,
    ui_in,
    uio_in,
    uio_oe,
    uio_out,
    uo_out);
 input clk;
 input ena;
 input rst_n;
 input [7:0] ui_in;
 input [7:0] uio_in;
 output [7:0] uio_oe;
 output [7:0] uio_out;
 output [7:0] uo_out;

 wire _0000_;
 wire _0001_;
 wire _0002_;
 wire _0003_;
 wire _0004_;
 wire _0005_;
 wire _0006_;
 wire _0007_;
 wire _0008_;
 wire _0009_;
 wire _0010_;
 wire _0011_;
 wire _0012_;
 wire _0013_;
 wire _0014_;
 wire _0015_;
 wire _0016_;
 wire _0017_;
 wire _0018_;
 wire _0019_;
 wire _0020_;
 wire _0021_;
 wire _0022_;
 wire _0023_;
 wire _0024_;
 wire _0025_;
 wire _0026_;
 wire _0027_;
 wire _0028_;
 wire _0029_;
 wire _0030_;
 wire _0031_;
 wire _0032_;
 wire _0033_;
 wire _0034_;
 wire _0035_;
 wire _0036_;
 wire _0037_;
 wire _0038_;
 wire _0039_;
 wire _0040_;
 wire _0041_;
 wire _0042_;
 wire _0043_;
 wire _0044_;
 wire _0045_;
 wire _0046_;
 wire _0047_;
 wire _0048_;
 wire _0049_;
 wire _0050_;
 wire _0051_;
 wire _0052_;
 wire _0053_;
 wire _0054_;
 wire _0055_;
 wire _0056_;
 wire _0057_;
 wire _0058_;
 wire _0059_;
 wire _0060_;
 wire _0061_;
 wire _0062_;
 wire _0063_;
 wire _0064_;
 wire _0065_;
 wire _0066_;
 wire _0067_;
 wire _0068_;
 wire _0069_;
 wire _0070_;
 wire _0071_;
 wire _0072_;
 wire _0073_;
 wire _0074_;
 wire _0075_;
 wire _0076_;
 wire _0077_;
 wire _0078_;
 wire _0079_;
 wire _0080_;
 wire _0081_;
 wire _0082_;
 wire _0083_;
 wire _0084_;
 wire _0085_;
 wire _0086_;
 wire _0087_;
 wire _0088_;
 wire _0089_;
 wire _0090_;
 wire _0091_;
 wire _0092_;
 wire _0093_;
 wire _0094_;
 wire _0095_;
 wire _0096_;
 wire _0097_;
 wire _0098_;
 wire _0099_;
 wire _0100_;
 wire _0101_;
 wire _0102_;
 wire _0103_;
 wire _0104_;
 wire _0105_;
 wire _0106_;
 wire _0107_;
 wire _0108_;
 wire _0109_;
 wire _0110_;
 wire _0111_;
 wire _0112_;
 wire _0113_;
 wire _0114_;
 wire _0115_;
 wire _0116_;
 wire _0117_;
 wire _0118_;
 wire _0119_;
 wire _0120_;
 wire _0121_;
 wire _0122_;
 wire _0123_;
 wire _0124_;
 wire _0125_;
 wire _0126_;
 wire _0127_;
 wire _0128_;
 wire _0129_;
 wire _0130_;
 wire _0131_;
 wire _0132_;
 wire _0133_;
 wire _0134_;
 wire _0135_;
 wire _0136_;
 wire _0137_;
 wire _0138_;
 wire _0139_;
 wire _0140_;
 wire _0141_;
 wire _0142_;
 wire _0143_;
 wire _0144_;
 wire _0145_;
 wire _0146_;
 wire _0147_;
 wire _0148_;
 wire _0149_;
 wire _0150_;
 wire _0151_;
 wire _0152_;
 wire _0153_;
 wire _0154_;
 wire _0155_;
 wire _0156_;
 wire _0157_;
 wire _0158_;
 wire _0159_;
 wire _0160_;
 wire _0161_;
 wire _0162_;
 wire _0163_;
 wire _0164_;
 wire _0165_;
 wire _0166_;
 wire _0167_;
 wire _0168_;
 wire _0169_;
 wire _0170_;
 wire _0171_;
 wire _0172_;
 wire _0173_;
 wire _0174_;
 wire _0175_;
 wire _0176_;
 wire _0177_;
 wire _0178_;
 wire _0179_;
 wire _0180_;
 wire _0181_;
 wire _0182_;
 wire _0183_;
 wire _0184_;
 wire _0185_;
 wire _0186_;
 wire _0187_;
 wire _0188_;
 wire _0189_;
 wire _0190_;
 wire _0191_;
 wire _0192_;
 wire _0193_;
 wire _0194_;
 wire _0195_;
 wire _0196_;
 wire _0197_;
 wire _0198_;
 wire _0199_;
 wire _0200_;
 wire _0201_;
 wire _0202_;
 wire _0203_;
 wire _0204_;
 wire _0205_;
 wire _0206_;
 wire _0207_;
 wire _0208_;
 wire _0209_;
 wire _0210_;
 wire _0211_;
 wire _0212_;
 wire _0213_;
 wire _0214_;
 wire _0215_;
 wire _0216_;
 wire _0217_;
 wire _0218_;
 wire _0219_;
 wire _0220_;
 wire _0221_;
 wire _0222_;
 wire _0223_;
 wire _0224_;
 wire _0225_;
 wire _0226_;
 wire _0227_;
 wire _0228_;
 wire _0229_;
 wire _0230_;
 wire _0231_;
 wire _0232_;
 wire _0233_;
 wire _0234_;
 wire _0235_;
 wire _0236_;
 wire _0237_;
 wire _0238_;
 wire _0239_;
 wire _0240_;
 wire _0241_;
 wire _0242_;
 wire _0243_;
 wire _0244_;
 wire _0245_;
 wire _0246_;
 wire _0247_;
 wire _0248_;
 wire _0249_;
 wire _0250_;
 wire _0251_;
 wire _0252_;
 wire _0253_;
 wire _0254_;
 wire _0255_;
 wire _0256_;
 wire _0257_;
 wire _0258_;
 wire _0259_;
 wire _0260_;
 wire _0261_;
 wire _0262_;
 wire _0263_;
 wire _0264_;
 wire _0265_;
 wire _0266_;
 wire _0267_;
 wire _0268_;
 wire _0269_;
 wire _0270_;
 wire _0271_;
 wire _0272_;
 wire _0273_;
 wire _0274_;
 wire _0275_;
 wire _0276_;
 wire _0277_;
 wire _0278_;
 wire _0279_;
 wire _0280_;
 wire _0281_;
 wire _0282_;
 wire _0283_;
 wire _0284_;
 wire _0285_;
 wire _0286_;
 wire _0287_;
 wire _0288_;
 wire _0289_;
 wire _0290_;
 wire _0291_;
 wire _0292_;
 wire _0293_;
 wire _0294_;
 wire _0295_;
 wire _0296_;
 wire _0297_;
 wire _0298_;
 wire _0299_;
 wire _0300_;
 wire _0301_;
 wire _0302_;
 wire _0303_;
 wire _0304_;
 wire _0305_;
 wire _0306_;
 wire _0307_;
 wire _0308_;
 wire _0309_;
 wire _0310_;
 wire _0311_;
 wire _0312_;
 wire _0313_;
 wire _0314_;
 wire _0315_;
 wire _0316_;
 wire _0317_;
 wire _0318_;
 wire _0319_;
 wire _0320_;
 wire _0321_;
 wire _0322_;
 wire _0323_;
 wire _0324_;
 wire _0325_;
 wire _0326_;
 wire _0327_;
 wire _0328_;
 wire _0329_;
 wire _0330_;
 wire _0331_;
 wire _0332_;
 wire _0333_;
 wire _0334_;
 wire _0335_;
 wire _0336_;
 wire _0337_;
 wire _0338_;
 wire _0339_;
 wire _0340_;
 wire _0341_;
 wire _0342_;
 wire _0343_;
 wire _0344_;
 wire _0345_;
 wire _0346_;
 wire _0347_;
 wire _0348_;
 wire _0349_;
 wire _0350_;
 wire _0351_;
 wire _0352_;
 wire _0353_;
 wire _0354_;
 wire _0355_;
 wire _0356_;
 wire _0357_;
 wire _0358_;
 wire _0359_;
 wire _0360_;
 wire _0361_;
 wire _0362_;
 wire _0363_;
 wire _0364_;
 wire _0365_;
 wire _0366_;
 wire _0367_;
 wire _0368_;
 wire _0369_;
 wire _0370_;
 wire _0371_;
 wire _0372_;
 wire _0373_;
 wire _0374_;
 wire _0375_;
 wire _0376_;
 wire _0377_;
 wire _0378_;
 wire _0379_;
 wire _0380_;
 wire _0381_;
 wire _0382_;
 wire _0383_;
 wire _0384_;
 wire _0385_;
 wire _0386_;
 wire _0387_;
 wire _0388_;
 wire _0389_;
 wire _0390_;
 wire _0391_;
 wire _0392_;
 wire _0393_;
 wire _0394_;
 wire _0395_;
 wire _0396_;
 wire _0397_;
 wire _0398_;
 wire _0399_;
 wire _0400_;
 wire _0401_;
 wire _0402_;
 wire _0403_;
 wire _0404_;
 wire _0405_;
 wire _0406_;
 wire _0407_;
 wire _0408_;
 wire _0409_;
 wire _0410_;
 wire _0411_;
 wire _0412_;
 wire _0413_;
 wire _0414_;
 wire _0415_;
 wire _0416_;
 wire _0417_;
 wire _0418_;
 wire _0419_;
 wire _0420_;
 wire _0421_;
 wire _0422_;
 wire _0423_;
 wire _0424_;
 wire _0425_;
 wire _0426_;
 wire _0427_;
 wire _0428_;
 wire _0429_;
 wire _0430_;
 wire _0431_;
 wire _0432_;
 wire _0433_;
 wire _0434_;
 wire _0435_;
 wire _0436_;
 wire _0437_;
 wire _0438_;
 wire _0439_;
 wire _0440_;
 wire _0441_;
 wire _0442_;
 wire _0443_;
 wire _0444_;
 wire _0445_;
 wire _0446_;
 wire _0447_;
 wire _0448_;
 wire _0449_;
 wire _0450_;
 wire _0451_;
 wire _0452_;
 wire _0453_;
 wire _0454_;
 wire _0455_;
 wire _0456_;
 wire _0457_;
 wire _0458_;
 wire _0459_;
 wire _0460_;
 wire _0461_;
 wire _0462_;
 wire _0463_;
 wire _0464_;
 wire _0465_;
 wire _0466_;
 wire _0467_;
 wire _0468_;
 wire _0469_;
 wire _0470_;
 wire _0471_;
 wire _0472_;
 wire _0473_;
 wire _0474_;
 wire _0475_;
 wire _0476_;
 wire _0477_;
 wire _0478_;
 wire _0479_;
 wire _0480_;
 wire _0481_;
 wire _0482_;
 wire _0483_;
 wire _0484_;
 wire _0485_;
 wire _0486_;
 wire _0487_;
 wire _0488_;
 wire _0489_;
 wire _0490_;
 wire _0491_;
 wire _0492_;
 wire _0493_;
 wire _0494_;
 wire _0495_;
 wire _0496_;
 wire _0497_;
 wire _0498_;
 wire _0499_;
 wire _0500_;
 wire _0501_;
 wire _0502_;
 wire _0503_;
 wire _0504_;
 wire _0505_;
 wire _0506_;
 wire _0507_;
 wire _0508_;
 wire _0509_;
 wire _0510_;
 wire _0511_;
 wire _0512_;
 wire _0513_;
 wire _0514_;
 wire _0515_;
 wire _0516_;
 wire _0517_;
 wire _0518_;
 wire _0519_;
 wire _0520_;
 wire _0521_;
 wire _0522_;
 wire _0523_;
 wire _0524_;
 wire _0525_;
 wire _0526_;
 wire _0527_;
 wire _0528_;
 wire _0529_;
 wire _0530_;
 wire _0531_;
 wire _0532_;
 wire _0533_;
 wire _0534_;
 wire _0535_;
 wire _0536_;
 wire _0537_;
 wire _0538_;
 wire _0539_;
 wire _0540_;
 wire _0541_;
 wire _0542_;
 wire _0543_;
 wire _0544_;
 wire _0545_;
 wire _0546_;
 wire _0547_;
 wire _0548_;
 wire _0549_;
 wire _0550_;
 wire _0551_;
 wire _0552_;
 wire _0553_;
 wire _0554_;
 wire _0555_;
 wire _0556_;
 wire _0557_;
 wire _0558_;
 wire _0559_;
 wire _0560_;
 wire _0561_;
 wire _0562_;
 wire _0563_;
 wire _0564_;
 wire _0565_;
 wire _0566_;
 wire _0567_;
 wire _0568_;
 wire _0569_;
 wire _0570_;
 wire _0571_;
 wire _0572_;
 wire _0573_;
 wire _0574_;
 wire _0575_;
 wire _0576_;
 wire _0577_;
 wire _0578_;
 wire _0579_;
 wire _0580_;
 wire _0581_;
 wire _0582_;
 wire _0583_;
 wire _0584_;
 wire _0585_;
 wire _0586_;
 wire _0587_;
 wire _0588_;
 wire _0589_;
 wire _0590_;
 wire _0591_;
 wire _0592_;
 wire _0593_;
 wire _0594_;
 wire _0595_;
 wire _0596_;
 wire _0597_;
 wire _0598_;
 wire _0599_;
 wire _0600_;
 wire _0601_;
 wire _0602_;
 wire _0603_;
 wire _0604_;
 wire _0605_;
 wire _0606_;
 wire _0607_;
 wire _0608_;
 wire _0609_;
 wire _0610_;
 wire _0611_;
 wire _0612_;
 wire _0613_;
 wire _0614_;
 wire _0615_;
 wire _0616_;
 wire _0617_;
 wire _0618_;
 wire _0619_;
 wire _0620_;
 wire _0621_;
 wire _0622_;
 wire _0623_;
 wire _0624_;
 wire _0625_;
 wire _0626_;
 wire _0627_;
 wire _0628_;
 wire _0629_;
 wire _0630_;
 wire _0631_;
 wire _0632_;
 wire _0633_;
 wire _0634_;
 wire _0635_;
 wire _0636_;
 wire _0637_;
 wire _0638_;
 wire _0639_;
 wire _0640_;
 wire _0641_;
 wire _0642_;
 wire _0643_;
 wire _0644_;
 wire _0645_;
 wire _0646_;
 wire _0647_;
 wire _0648_;
 wire _0649_;
 wire _0650_;
 wire _0651_;
 wire _0652_;
 wire _0653_;
 wire _0654_;
 wire _0655_;
 wire _0656_;
 wire _0657_;
 wire _0658_;
 wire _0659_;
 wire _0660_;
 wire _0661_;
 wire _0662_;
 wire _0663_;
 wire _0664_;
 wire _0665_;
 wire _0666_;
 wire _0667_;
 wire _0668_;
 wire _0669_;
 wire _0670_;
 wire _0671_;
 wire _0672_;
 wire _0673_;
 wire _0674_;
 wire _0675_;
 wire _0676_;
 wire _0677_;
 wire _0678_;
 wire _0679_;
 wire _0680_;
 wire _0681_;
 wire _0682_;
 wire _0683_;
 wire _0684_;
 wire _0685_;
 wire _0686_;
 wire _0687_;
 wire _0688_;
 wire _0689_;
 wire _0690_;
 wire _0691_;
 wire _0692_;
 wire _0693_;
 wire _0694_;
 wire _0695_;
 wire _0696_;
 wire _0697_;
 wire _0698_;
 wire _0699_;
 wire _0700_;
 wire _0701_;
 wire _0702_;
 wire _0703_;
 wire _0704_;
 wire _0705_;
 wire _0706_;
 wire _0707_;
 wire _0708_;
 wire _0709_;
 wire _0710_;
 wire _0711_;
 wire _0712_;
 wire _0713_;
 wire _0714_;
 wire _0715_;
 wire _0716_;
 wire _0717_;
 wire _0718_;
 wire _0719_;
 wire _0720_;
 wire _0721_;
 wire _0722_;
 wire _0723_;
 wire _0724_;
 wire _0725_;
 wire _0726_;
 wire _0727_;
 wire _0728_;
 wire _0729_;
 wire _0730_;
 wire _0731_;
 wire _0732_;
 wire _0733_;
 wire _0734_;
 wire _0735_;
 wire _0736_;
 wire _0737_;
 wire _0738_;
 wire _0739_;
 wire _0740_;
 wire _0741_;
 wire _0742_;
 wire _0743_;
 wire _0744_;
 wire _0745_;
 wire _0746_;
 wire _0747_;
 wire _0748_;
 wire _0749_;
 wire _0750_;
 wire _0751_;
 wire _0752_;
 wire _0753_;
 wire _0754_;
 wire _0755_;
 wire _0756_;
 wire _0757_;
 wire _0758_;
 wire _0759_;
 wire _0760_;
 wire _0761_;
 wire _0762_;
 wire _0763_;
 wire _0764_;
 wire _0765_;
 wire _0766_;
 wire _0767_;
 wire _0768_;
 wire _0769_;
 wire _0770_;
 wire _0771_;
 wire _0772_;
 wire _0773_;
 wire _0774_;
 wire _0775_;
 wire _0776_;
 wire _0777_;
 wire _0778_;
 wire _0779_;
 wire _0780_;
 wire _0781_;
 wire _0782_;
 wire _0783_;
 wire _0784_;
 wire _0785_;
 wire _0786_;
 wire _0787_;
 wire _0788_;
 wire _0789_;
 wire _0790_;
 wire _0791_;
 wire _0792_;
 wire _0793_;
 wire _0794_;
 wire _0795_;
 wire _0796_;
 wire _0797_;
 wire _0798_;
 wire _0799_;
 wire _0800_;
 wire _0801_;
 wire _0802_;
 wire _0803_;
 wire _0804_;
 wire _0805_;
 wire _0806_;
 wire _0807_;
 wire _0808_;
 wire _0809_;
 wire _0810_;
 wire _0811_;
 wire _0812_;
 wire _0813_;
 wire _0814_;
 wire _0815_;
 wire _0816_;
 wire _0817_;
 wire _0818_;
 wire _0819_;
 wire _0820_;
 wire _0821_;
 wire _0822_;
 wire _0823_;
 wire _0824_;
 wire _0825_;
 wire _0826_;
 wire _0827_;
 wire _0828_;
 wire _0829_;
 wire _0830_;
 wire _0831_;
 wire _0832_;
 wire _0833_;
 wire _0834_;
 wire _0835_;
 wire _0836_;
 wire _0837_;
 wire _0838_;
 wire _0839_;
 wire _0840_;
 wire _0841_;
 wire _0842_;
 wire _0843_;
 wire _0844_;
 wire _0845_;
 wire _0846_;
 wire _0847_;
 wire _0848_;
 wire _0849_;
 wire _0850_;
 wire _0851_;
 wire _0852_;
 wire _0853_;
 wire _0854_;
 wire _0855_;
 wire _0856_;
 wire _0857_;
 wire _0858_;
 wire _0859_;
 wire _0860_;
 wire _0861_;
 wire _0862_;
 wire _0863_;
 wire _0864_;
 wire _0865_;
 wire _0866_;
 wire _0867_;
 wire _0868_;
 wire _0869_;
 wire _0870_;
 wire _0871_;
 wire _0872_;
 wire _0873_;
 wire _0874_;
 wire _0875_;
 wire _0876_;
 wire _0877_;
 wire _0878_;
 wire _0879_;
 wire _0880_;
 wire _0881_;
 wire _0882_;
 wire _0883_;
 wire _0884_;
 wire _0885_;
 wire _0886_;
 wire _0887_;
 wire _0888_;
 wire _0889_;
 wire _0890_;
 wire _0891_;
 wire _0892_;
 wire _0893_;
 wire _0894_;
 wire _0895_;
 wire _0896_;
 wire _0897_;
 wire _0898_;
 wire _0899_;
 wire _0900_;
 wire _0901_;
 wire _0902_;
 wire _0903_;
 wire _0904_;
 wire _0905_;
 wire _0906_;
 wire _0907_;
 wire _0908_;
 wire _0909_;
 wire _0910_;
 wire _0911_;
 wire _0912_;
 wire _0913_;
 wire _0914_;
 wire _0915_;
 wire _0916_;
 wire _0917_;
 wire _0918_;
 wire _0919_;
 wire _0920_;
 wire _0921_;
 wire _0922_;
 wire _0923_;
 wire _0924_;
 wire _0925_;
 wire _0926_;
 wire _0927_;
 wire _0928_;
 wire _0929_;
 wire _0930_;
 wire _0931_;
 wire _0932_;
 wire _0933_;
 wire _0934_;
 wire _0935_;
 wire _0936_;
 wire _0937_;
 wire _0938_;
 wire _0939_;
 wire _0940_;
 wire _0941_;
 wire _0942_;
 wire _0943_;
 wire _0944_;
 wire _0945_;
 wire _0946_;
 wire _0947_;
 wire _0948_;
 wire _0949_;
 wire _0950_;
 wire _0951_;
 wire _0952_;
 wire _0953_;
 wire _0954_;
 wire _0955_;
 wire _0956_;
 wire _0957_;
 wire _0958_;
 wire _0959_;
 wire _0960_;
 wire _0961_;
 wire _0962_;
 wire _0963_;
 wire _0964_;
 wire _0965_;
 wire _0966_;
 wire _0967_;
 wire _0968_;
 wire _0969_;
 wire _0970_;
 wire _0971_;
 wire _0972_;
 wire _0973_;
 wire _0974_;
 wire _0975_;
 wire _0976_;
 wire _0977_;
 wire _0978_;
 wire _0979_;
 wire _0980_;
 wire _0981_;
 wire _0982_;
 wire _0983_;
 wire _0984_;
 wire _0985_;
 wire _0986_;
 wire _0987_;
 wire _0988_;
 wire _0989_;
 wire _0990_;
 wire _0991_;
 wire _0992_;
 wire _0993_;
 wire _0994_;
 wire _0995_;
 wire _0996_;
 wire _0997_;
 wire _0998_;
 wire _0999_;
 wire _1000_;
 wire _1001_;
 wire _1002_;
 wire _1003_;
 wire _1004_;
 wire _1005_;
 wire _1006_;
 wire _1007_;
 wire _1008_;
 wire _1009_;
 wire _1010_;
 wire _1011_;
 wire _1012_;
 wire _1013_;
 wire _1014_;
 wire _1015_;
 wire _1016_;
 wire _1017_;
 wire _1018_;
 wire _1019_;
 wire _1020_;
 wire _1021_;
 wire _1022_;
 wire _1023_;
 wire _1024_;
 wire _1025_;
 wire _1026_;
 wire _1027_;
 wire _1028_;
 wire _1029_;
 wire _1030_;
 wire _1031_;
 wire _1032_;
 wire _1033_;
 wire _1034_;
 wire _1035_;
 wire _1036_;
 wire _1037_;
 wire _1038_;
 wire _1039_;
 wire _1040_;
 wire _1041_;
 wire _1042_;
 wire _1043_;
 wire _1044_;
 wire _1045_;
 wire _1046_;
 wire _1047_;
 wire _1048_;
 wire _1049_;
 wire _1050_;
 wire _1051_;
 wire _1052_;
 wire _1053_;
 wire _1054_;
 wire _1055_;
 wire _1056_;
 wire _1057_;
 wire _1058_;
 wire _1059_;
 wire _1060_;
 wire _1061_;
 wire _1062_;
 wire _1063_;
 wire _1064_;
 wire _1065_;
 wire _1066_;
 wire _1067_;
 wire _1068_;
 wire _1069_;
 wire _1070_;
 wire _1071_;
 wire _1072_;
 wire _1073_;
 wire _1074_;
 wire _1075_;
 wire _1076_;
 wire _1077_;
 wire _1078_;
 wire _1079_;
 wire _1080_;
 wire _1081_;
 wire _1082_;
 wire _1083_;
 wire _1084_;
 wire _1085_;
 wire _1086_;
 wire _1087_;
 wire _1088_;
 wire _1089_;
 wire _1090_;
 wire _1091_;
 wire _1092_;
 wire _1093_;
 wire _1094_;
 wire _1095_;
 wire _1096_;
 wire _1097_;
 wire _1098_;
 wire _1099_;
 wire _1100_;
 wire _1101_;
 wire _1102_;
 wire _1103_;
 wire _1104_;
 wire _1105_;
 wire _1106_;
 wire _1107_;
 wire _1108_;
 wire _1109_;
 wire _1110_;
 wire _1111_;
 wire _1112_;
 wire _1113_;
 wire _1114_;
 wire _1115_;
 wire _1116_;
 wire _1117_;
 wire _1118_;
 wire _1119_;
 wire _1120_;
 wire _1121_;
 wire _1122_;
 wire _1123_;
 wire _1124_;
 wire _1125_;
 wire _1126_;
 wire _1127_;
 wire _1128_;
 wire _1129_;
 wire _1130_;
 wire _1131_;
 wire _1132_;
 wire _1133_;
 wire _1134_;
 wire _1135_;
 wire _1136_;
 wire _1137_;
 wire _1138_;
 wire _1139_;
 wire _1140_;
 wire _1141_;
 wire _1142_;
 wire _1143_;
 wire _1144_;
 wire _1145_;
 wire _1146_;
 wire _1147_;
 wire _1148_;
 wire _1149_;
 wire _1150_;
 wire _1151_;
 wire _1152_;
 wire _1153_;
 wire _1154_;
 wire _1155_;
 wire _1156_;
 wire _1157_;
 wire _1158_;
 wire _1159_;
 wire _1160_;
 wire _1161_;
 wire _1162_;
 wire _1163_;
 wire _1164_;
 wire _1165_;
 wire _1166_;
 wire _1167_;
 wire _1168_;
 wire _1169_;
 wire _1170_;
 wire _1171_;
 wire _1172_;
 wire _1173_;
 wire _1174_;
 wire _1175_;
 wire _1176_;
 wire _1177_;
 wire _1178_;
 wire _1179_;
 wire _1180_;
 wire _1181_;
 wire _1182_;
 wire _1183_;
 wire _1184_;
 wire _1185_;
 wire _1186_;
 wire _1187_;
 wire _1188_;
 wire _1189_;
 wire _1190_;
 wire _1191_;
 wire _1192_;
 wire _1193_;
 wire _1194_;
 wire _1195_;
 wire _1196_;
 wire _1197_;
 wire _1198_;
 wire _1199_;
 wire _1200_;
 wire _1201_;
 wire _1202_;
 wire _1203_;
 wire _1204_;
 wire _1205_;
 wire _1206_;
 wire _1207_;
 wire _1208_;
 wire _1209_;
 wire _1210_;
 wire _1211_;
 wire _1212_;
 wire _1213_;
 wire _1214_;
 wire _1215_;
 wire _1216_;
 wire _1217_;
 wire _1218_;
 wire _1219_;
 wire _1220_;
 wire _1221_;
 wire _1222_;
 wire _1223_;
 wire _1224_;
 wire _1225_;
 wire _1226_;
 wire _1227_;
 wire _1228_;
 wire _1229_;
 wire _1230_;
 wire _1231_;
 wire _1232_;
 wire _1233_;
 wire _1234_;
 wire _1235_;
 wire _1236_;
 wire _1237_;
 wire _1238_;
 wire _1239_;
 wire _1240_;
 wire _1241_;
 wire _1242_;
 wire _1243_;
 wire _1244_;
 wire _1245_;
 wire _1246_;
 wire _1247_;
 wire _1248_;
 wire _1249_;
 wire _1250_;
 wire _1251_;
 wire _1252_;
 wire _1253_;
 wire _1254_;
 wire _1255_;
 wire _1256_;
 wire _1257_;
 wire _1258_;
 wire _1259_;
 wire _1260_;
 wire _1261_;
 wire _1262_;
 wire _1263_;
 wire _1264_;
 wire _1265_;
 wire _1266_;
 wire _1267_;
 wire _1268_;
 wire _1269_;
 wire _1270_;
 wire _1271_;
 wire _1272_;
 wire _1273_;
 wire _1274_;
 wire _1275_;
 wire _1276_;
 wire _1277_;
 wire _1278_;
 wire _1279_;
 wire _1280_;
 wire _1281_;
 wire _1282_;
 wire _1283_;
 wire _1284_;
 wire _1285_;
 wire _1286_;
 wire _1287_;
 wire _1288_;
 wire _1289_;
 wire _1290_;
 wire _1291_;
 wire _1292_;
 wire _1293_;
 wire _1294_;
 wire _1295_;
 wire _1296_;
 wire _1297_;
 wire _1298_;
 wire _1299_;
 wire _1300_;
 wire _1301_;
 wire _1302_;
 wire _1303_;
 wire _1304_;
 wire _1305_;
 wire _1306_;
 wire _1307_;
 wire _1308_;
 wire _1309_;
 wire _1310_;
 wire _1311_;
 wire _1312_;
 wire _1313_;
 wire _1314_;
 wire _1315_;
 wire _1316_;
 wire _1317_;
 wire _1318_;
 wire _1319_;
 wire _1320_;
 wire _1321_;
 wire _1322_;
 wire _1323_;
 wire _1324_;
 wire _1325_;
 wire _1326_;
 wire _1327_;
 wire _1328_;
 wire _1329_;
 wire _1330_;
 wire _1331_;
 wire _1332_;
 wire _1333_;
 wire _1334_;
 wire _1335_;
 wire _1336_;
 wire _1337_;
 wire _1338_;
 wire _1339_;
 wire _1340_;
 wire _1341_;
 wire _1342_;
 wire _1343_;
 wire _1344_;
 wire _1345_;
 wire _1346_;
 wire _1347_;
 wire _1348_;
 wire _1349_;
 wire _1350_;
 wire _1351_;
 wire _1352_;
 wire _1353_;
 wire _1354_;
 wire _1355_;
 wire _1356_;
 wire _1357_;
 wire _1358_;
 wire _1359_;
 wire _1360_;
 wire _1361_;
 wire _1362_;
 wire _1363_;
 wire _1364_;
 wire _1365_;
 wire _1366_;
 wire _1367_;
 wire _1368_;
 wire _1369_;
 wire _1370_;
 wire _1371_;
 wire _1372_;
 wire _1373_;
 wire _1374_;
 wire _1375_;
 wire _1376_;
 wire _1377_;
 wire _1378_;
 wire _1379_;
 wire _1380_;
 wire _1381_;
 wire _1382_;
 wire _1383_;
 wire _1384_;
 wire _1385_;
 wire _1386_;
 wire _1387_;
 wire _1388_;
 wire _1389_;
 wire _1390_;
 wire _1391_;
 wire _1392_;
 wire _1393_;
 wire _1394_;
 wire _1395_;
 wire _1396_;
 wire _1397_;
 wire _1398_;
 wire _1399_;
 wire _1400_;
 wire _1401_;
 wire _1402_;
 wire _1403_;
 wire _1404_;
 wire _1405_;
 wire _1406_;
 wire _1407_;
 wire _1408_;
 wire _1409_;
 wire _1410_;
 wire _1411_;
 wire _1412_;
 wire _1413_;
 wire _1414_;
 wire _1415_;
 wire _1416_;
 wire _1417_;
 wire _1418_;
 wire _1419_;
 wire _1420_;
 wire _1421_;
 wire _1422_;
 wire _1423_;
 wire _1424_;
 wire _1425_;
 wire _1426_;
 wire _1427_;
 wire _1428_;
 wire _1429_;
 wire _1430_;
 wire _1431_;
 wire _1432_;
 wire _1433_;
 wire _1434_;
 wire _1435_;
 wire _1436_;
 wire _1437_;
 wire _1438_;
 wire _1439_;
 wire _1440_;
 wire _1441_;
 wire _1442_;
 wire _1443_;
 wire _1444_;
 wire _1445_;
 wire _1446_;
 wire _1447_;
 wire _1448_;
 wire _1449_;
 wire _1450_;
 wire _1451_;
 wire _1452_;
 wire _1453_;
 wire _1454_;
 wire _1455_;
 wire _1456_;
 wire _1457_;
 wire _1458_;
 wire _1459_;
 wire _1460_;
 wire _1461_;
 wire _1462_;
 wire _1463_;
 wire _1464_;
 wire _1465_;
 wire _1466_;
 wire _1467_;
 wire _1468_;
 wire _1469_;
 wire _1470_;
 wire _1471_;
 wire _1472_;
 wire _1473_;
 wire _1474_;
 wire _1475_;
 wire _1476_;
 wire _1477_;
 wire _1478_;
 wire _1479_;
 wire _1480_;
 wire _1481_;
 wire _1482_;
 wire _1483_;
 wire _1484_;
 wire _1485_;
 wire _1486_;
 wire _1487_;
 wire _1488_;
 wire _1489_;
 wire _1490_;
 wire _1491_;
 wire _1492_;
 wire _1493_;
 wire _1494_;
 wire _1495_;
 wire _1496_;
 wire _1497_;
 wire _1498_;
 wire _1499_;
 wire _1500_;
 wire _1501_;
 wire _1502_;
 wire _1503_;
 wire _1504_;
 wire _1505_;
 wire _1506_;
 wire _1507_;
 wire _1508_;
 wire _1509_;
 wire _1510_;
 wire _1511_;
 wire _1512_;
 wire _1513_;
 wire _1514_;
 wire _1515_;
 wire _1516_;
 wire _1517_;
 wire _1518_;
 wire _1519_;
 wire _1520_;
 wire _1521_;
 wire _1522_;
 wire _1523_;
 wire _1524_;
 wire _1525_;
 wire _1526_;
 wire _1527_;
 wire _1528_;
 wire _1529_;
 wire _1530_;
 wire _1531_;
 wire _1532_;
 wire _1533_;
 wire _1534_;
 wire _1535_;
 wire _1536_;
 wire _1537_;
 wire _1538_;
 wire _1539_;
 wire _1540_;
 wire _1541_;
 wire _1542_;
 wire _1543_;
 wire _1544_;
 wire _1545_;
 wire _1546_;
 wire _1547_;
 wire _1548_;
 wire _1549_;
 wire _1550_;
 wire _1551_;
 wire _1552_;
 wire _1553_;
 wire _1554_;
 wire _1555_;
 wire _1556_;
 wire _1557_;
 wire _1558_;
 wire _1559_;
 wire _1560_;
 wire _1561_;
 wire _1562_;
 wire _1563_;
 wire _1564_;
 wire _1565_;
 wire _1566_;
 wire _1567_;
 wire _1568_;
 wire _1569_;
 wire _1570_;
 wire _1571_;
 wire _1572_;
 wire _1573_;
 wire _1574_;
 wire _1575_;
 wire _1576_;
 wire _1577_;
 wire _1578_;
 wire _1579_;
 wire _1580_;
 wire _1581_;
 wire _1582_;
 wire _1583_;
 wire _1584_;
 wire _1585_;
 wire _1586_;
 wire _1587_;
 wire _1588_;
 wire _1589_;
 wire _1590_;
 wire _1591_;
 wire _1592_;
 wire _1593_;
 wire _1594_;
 wire _1595_;
 wire _1596_;
 wire _1597_;
 wire _1598_;
 wire _1599_;
 wire _1600_;
 wire _1601_;
 wire _1602_;
 wire _1603_;
 wire _1604_;
 wire _1605_;
 wire _1606_;
 wire _1607_;
 wire _1608_;
 wire _1609_;
 wire _1610_;
 wire _1611_;
 wire _1612_;
 wire _1613_;
 wire _1614_;
 wire _1615_;
 wire _1616_;
 wire _1617_;
 wire _1618_;
 wire _1619_;
 wire _1620_;
 wire _1621_;
 wire _1622_;
 wire _1623_;
 wire _1624_;
 wire _1625_;
 wire _1626_;
 wire _1627_;
 wire _1628_;
 wire _1629_;
 wire _1630_;
 wire _1631_;
 wire _1632_;
 wire _1633_;
 wire _1634_;
 wire _1635_;
 wire _1636_;
 wire _1637_;
 wire _1638_;
 wire _1639_;
 wire _1640_;
 wire _1641_;
 wire _1642_;
 wire _1643_;
 wire _1644_;
 wire _1645_;
 wire _1646_;
 wire _1647_;
 wire _1648_;
 wire _1649_;
 wire _1650_;
 wire _1651_;
 wire _1652_;
 wire _1653_;
 wire _1654_;
 wire _1655_;
 wire _1656_;
 wire _1657_;
 wire _1658_;
 wire _1659_;
 wire _1660_;
 wire _1661_;
 wire _1662_;
 wire _1663_;
 wire _1664_;
 wire _1665_;
 wire _1666_;
 wire _1667_;
 wire _1668_;
 wire _1669_;
 wire _1670_;
 wire _1671_;
 wire _1672_;
 wire _1673_;
 wire _1674_;
 wire _1675_;
 wire _1676_;
 wire _1677_;
 wire _1678_;
 wire _1679_;
 wire _1680_;
 wire _1681_;
 wire _1682_;
 wire _1683_;
 wire _1684_;
 wire _1685_;
 wire _1686_;
 wire _1687_;
 wire _1688_;
 wire _1689_;
 wire _1690_;
 wire _1691_;
 wire _1692_;
 wire _1693_;
 wire _1694_;
 wire _1695_;
 wire _1696_;
 wire _1697_;
 wire _1698_;
 wire _1699_;
 wire _1700_;
 wire _1701_;
 wire _1702_;
 wire _1703_;
 wire _1704_;
 wire _1705_;
 wire _1706_;
 wire _1707_;
 wire _1708_;
 wire _1709_;
 wire _1710_;
 wire _1711_;
 wire _1712_;
 wire _1713_;
 wire _1714_;
 wire _1715_;
 wire _1716_;
 wire _1717_;
 wire _1718_;
 wire _1719_;
 wire _1720_;
 wire _1721_;
 wire _1722_;
 wire _1723_;
 wire _1724_;
 wire _1725_;
 wire _1726_;
 wire _1727_;
 wire _1728_;
 wire _1729_;
 wire _1730_;
 wire _1731_;
 wire _1732_;
 wire _1733_;
 wire _1734_;
 wire _1735_;
 wire _1736_;
 wire _1737_;
 wire _1738_;
 wire _1739_;
 wire _1740_;
 wire _1741_;
 wire _1742_;
 wire _1743_;
 wire _1744_;
 wire _1745_;
 wire _1746_;
 wire _1747_;
 wire _1748_;
 wire _1749_;
 wire _1750_;
 wire _1751_;
 wire _1752_;
 wire _1753_;
 wire _1754_;
 wire _1755_;
 wire _1756_;
 wire _1757_;
 wire _1758_;
 wire _1759_;
 wire _1760_;
 wire _1761_;
 wire _1762_;
 wire _1763_;
 wire _1764_;
 wire _1765_;
 wire _1766_;
 wire _1767_;
 wire _1768_;
 wire _1769_;
 wire _1770_;
 wire _1771_;
 wire _1772_;
 wire _1773_;
 wire _1774_;
 wire _1775_;
 wire _1776_;
 wire _1777_;
 wire _1778_;
 wire _1779_;
 wire _1780_;
 wire _1781_;
 wire _1782_;
 wire _1783_;
 wire _1784_;
 wire _1785_;
 wire _1786_;
 wire _1787_;
 wire _1788_;
 wire _1789_;
 wire _1790_;
 wire _1791_;
 wire _1792_;
 wire _1793_;
 wire _1794_;
 wire _1795_;
 wire _1796_;
 wire _1797_;
 wire _1798_;
 wire _1799_;
 wire _1800_;
 wire _1801_;
 wire _1802_;
 wire _1803_;
 wire _1804_;
 wire _1805_;
 wire _1806_;
 wire _1807_;
 wire _1808_;
 wire _1809_;
 wire _1810_;
 wire _1811_;
 wire _1812_;
 wire _1813_;
 wire _1814_;
 wire _1815_;
 wire _1816_;
 wire _1817_;
 wire _1818_;
 wire _1819_;
 wire _1820_;
 wire _1821_;
 wire _1822_;
 wire _1823_;
 wire _1824_;
 wire _1825_;
 wire _1826_;
 wire _1827_;
 wire _1828_;
 wire _1829_;
 wire _1830_;
 wire _1831_;
 wire _1832_;
 wire _1833_;
 wire _1834_;
 wire _1835_;
 wire _1836_;
 wire _1837_;
 wire _1838_;
 wire _1839_;
 wire _1840_;
 wire _1841_;
 wire _1842_;
 wire _1843_;
 wire _1844_;
 wire _1845_;
 wire _1846_;
 wire _1847_;
 wire _1848_;
 wire _1849_;
 wire _1850_;
 wire _1851_;
 wire _1852_;
 wire _1853_;
 wire _1854_;
 wire _1855_;
 wire _1856_;
 wire _1857_;
 wire _1858_;
 wire _1859_;
 wire _1860_;
 wire _1861_;
 wire _1862_;
 wire _1863_;
 wire _1864_;
 wire _1865_;
 wire _1866_;
 wire _1867_;
 wire _1868_;
 wire _1869_;
 wire _1870_;
 wire _1871_;
 wire _1872_;
 wire _1873_;
 wire _1874_;
 wire _1875_;
 wire _1876_;
 wire _1877_;
 wire _1878_;
 wire _1879_;
 wire _1880_;
 wire _1881_;
 wire _1882_;
 wire _1883_;
 wire _1884_;
 wire _1885_;
 wire _1886_;
 wire _1887_;
 wire _1888_;
 wire _1889_;
 wire _1890_;
 wire _1891_;
 wire _1892_;
 wire _1893_;
 wire _1894_;
 wire _1895_;
 wire _1896_;
 wire _1897_;
 wire _1898_;
 wire _1899_;
 wire _1900_;
 wire _1901_;
 wire _1902_;
 wire _1903_;
 wire _1904_;
 wire _1905_;
 wire _1906_;
 wire _1907_;
 wire _1908_;
 wire _1909_;
 wire _1910_;
 wire _1911_;
 wire _1912_;
 wire _1913_;
 wire _1914_;
 wire _1915_;
 wire _1916_;
 wire _1917_;
 wire _1918_;
 wire _1919_;
 wire _1920_;
 wire _1921_;
 wire _1922_;
 wire _1923_;
 wire _1924_;
 wire _1925_;
 wire _1926_;
 wire _1927_;
 wire _1928_;
 wire _1929_;
 wire _1930_;
 wire _1931_;
 wire _1932_;
 wire _1933_;
 wire _1934_;
 wire _1935_;
 wire _1936_;
 wire _1937_;
 wire _1938_;
 wire _1939_;
 wire _1940_;
 wire _1941_;
 wire _1942_;
 wire _1943_;
 wire _1944_;
 wire _1945_;
 wire _1946_;
 wire _1947_;
 wire _1948_;
 wire _1949_;
 wire _1950_;
 wire _1951_;
 wire _1952_;
 wire _1953_;
 wire _1954_;
 wire _1955_;
 wire _1956_;
 wire _1957_;
 wire _1958_;
 wire _1959_;
 wire _1960_;
 wire _1961_;
 wire _1962_;
 wire _1963_;
 wire _1964_;
 wire _1965_;
 wire _1966_;
 wire _1967_;
 wire _1968_;
 wire _1969_;
 wire _1970_;
 wire _1971_;
 wire _1972_;
 wire _1973_;
 wire _1974_;
 wire _1975_;
 wire _1976_;
 wire _1977_;
 wire _1978_;
 wire _1979_;
 wire _1980_;
 wire _1981_;
 wire _1982_;
 wire _1983_;
 wire _1984_;
 wire _1985_;
 wire _1986_;
 wire _1987_;
 wire _1988_;
 wire _1989_;
 wire _1990_;
 wire _1991_;
 wire _1992_;
 wire _1993_;
 wire _1994_;
 wire _1995_;
 wire _1996_;
 wire _1997_;
 wire _1998_;
 wire _1999_;
 wire _2000_;
 wire _2001_;
 wire _2002_;
 wire _2003_;
 wire _2004_;
 wire _2005_;
 wire _2006_;
 wire _2007_;
 wire _2008_;
 wire _2009_;
 wire _2010_;
 wire _2011_;
 wire _2012_;
 wire _2013_;
 wire _2014_;
 wire _2015_;
 wire _2016_;
 wire _2017_;
 wire _2018_;
 wire _2019_;
 wire _2020_;
 wire _2021_;
 wire _2022_;
 wire _2023_;
 wire _2024_;
 wire _2025_;
 wire _2026_;
 wire _2027_;
 wire _2028_;
 wire _2029_;
 wire _2030_;
 wire _2031_;
 wire _2032_;
 wire _2033_;
 wire _2034_;
 wire _2035_;
 wire _2036_;
 wire _2037_;
 wire _2038_;
 wire _2039_;
 wire _2040_;
 wire _2041_;
 wire _2042_;
 wire _2043_;
 wire _2044_;
 wire _2045_;
 wire _2046_;
 wire _2047_;
 wire _2048_;
 wire _2049_;
 wire _2050_;
 wire _2051_;
 wire _2052_;
 wire _2053_;
 wire _2054_;
 wire _2055_;
 wire _2056_;
 wire _2057_;
 wire _2058_;
 wire _2059_;
 wire _2060_;
 wire _2061_;
 wire _2062_;
 wire _2063_;
 wire _2064_;
 wire _2065_;
 wire _2066_;
 wire _2067_;
 wire _2068_;
 wire _2069_;
 wire _2070_;
 wire _2071_;
 wire _2072_;
 wire _2073_;
 wire _2074_;
 wire _2075_;
 wire _2076_;
 wire _2077_;
 wire _2078_;
 wire _2079_;
 wire _2080_;
 wire _2081_;
 wire _2082_;
 wire _2083_;
 wire _2084_;
 wire _2085_;
 wire _2086_;
 wire _2087_;
 wire _2088_;
 wire _2089_;
 wire _2090_;
 wire _2091_;
 wire _2092_;
 wire _2093_;
 wire _2094_;
 wire _2095_;
 wire _2096_;
 wire _2097_;
 wire _2098_;
 wire _2099_;
 wire _2100_;
 wire _2101_;
 wire _2102_;
 wire _2103_;
 wire _2104_;
 wire _2105_;
 wire _2106_;
 wire _2107_;
 wire _2108_;
 wire _2109_;
 wire _2110_;
 wire _2111_;
 wire _2112_;
 wire _2113_;
 wire _2114_;
 wire _2115_;
 wire _2116_;
 wire _2117_;
 wire _2118_;
 wire _2119_;
 wire _2120_;
 wire _2121_;
 wire _2122_;
 wire _2123_;
 wire _2124_;
 wire _2125_;
 wire _2126_;
 wire _2127_;
 wire _2128_;
 wire _2129_;
 wire _2130_;
 wire _2131_;
 wire _2132_;
 wire _2133_;
 wire _2134_;
 wire _2135_;
 wire _2136_;
 wire _2137_;
 wire _2138_;
 wire _2139_;
 wire _2140_;
 wire _2141_;
 wire _2142_;
 wire _2143_;
 wire _2144_;
 wire _2145_;
 wire _2146_;
 wire _2147_;
 wire _2148_;
 wire _2149_;
 wire _2150_;
 wire _2151_;
 wire _2152_;
 wire _2153_;
 wire _2154_;
 wire _2155_;
 wire _2156_;
 wire _2157_;
 wire _2158_;
 wire _2159_;
 wire _2160_;
 wire _2161_;
 wire _2162_;
 wire _2163_;
 wire _2164_;
 wire _2165_;
 wire _2166_;
 wire _2167_;
 wire _2168_;
 wire _2169_;
 wire _2170_;
 wire _2171_;
 wire _2172_;
 wire _2173_;
 wire _2174_;
 wire _2175_;
 wire _2176_;
 wire _2177_;
 wire _2178_;
 wire _2179_;
 wire _2180_;
 wire _2181_;
 wire _2182_;
 wire _2183_;
 wire _2184_;
 wire _2185_;
 wire _2186_;
 wire _2187_;
 wire _2188_;
 wire _2189_;
 wire _2190_;
 wire _2191_;
 wire _2192_;
 wire _2193_;
 wire _2194_;
 wire _2195_;
 wire _2196_;
 wire _2197_;
 wire _2198_;
 wire _2199_;
 wire _2200_;
 wire _2201_;
 wire _2202_;
 wire _2203_;
 wire _2204_;
 wire _2205_;
 wire _2206_;
 wire _2207_;
 wire _2208_;
 wire _2209_;
 wire _2210_;
 wire _2211_;
 wire _2212_;
 wire _2213_;
 wire _2214_;
 wire _2215_;
 wire _2216_;
 wire _2217_;
 wire _2218_;
 wire _2219_;
 wire _2220_;
 wire _2221_;
 wire _2222_;
 wire _2223_;
 wire _2224_;
 wire _2225_;
 wire _2226_;
 wire _2227_;
 wire _2228_;
 wire _2229_;
 wire _2230_;
 wire _2231_;
 wire _2232_;
 wire _2233_;
 wire _2234_;
 wire _2235_;
 wire _2236_;
 wire _2237_;
 wire _2238_;
 wire _2239_;
 wire _2240_;
 wire _2241_;
 wire _2242_;
 wire _2243_;
 wire _2244_;
 wire _2245_;
 wire _2246_;
 wire _2247_;
 wire _2248_;
 wire _2249_;
 wire _2250_;
 wire _2251_;
 wire _2252_;
 wire _2253_;
 wire _2254_;
 wire _2255_;
 wire _2256_;
 wire _2257_;
 wire _2258_;
 wire _2259_;
 wire _2260_;
 wire _2261_;
 wire _2262_;
 wire _2263_;
 wire _2264_;
 wire _2265_;
 wire _2266_;
 wire _2267_;
 wire _2268_;
 wire _2269_;
 wire _2270_;
 wire _2271_;
 wire _2272_;
 wire _2273_;
 wire _2274_;
 wire _2275_;
 wire _2276_;
 wire _2277_;
 wire _2278_;
 wire _2279_;
 wire _2280_;
 wire _2281_;
 wire _2282_;
 wire _2283_;
 wire _2284_;
 wire _2285_;
 wire _2286_;
 wire _2287_;
 wire _2288_;
 wire _2289_;
 wire _2290_;
 wire _2291_;
 wire _2292_;
 wire _2293_;
 wire _2294_;
 wire _2295_;
 wire _2296_;
 wire _2297_;
 wire _2298_;
 wire _2299_;
 wire _2300_;
 wire _2301_;
 wire _2302_;
 wire _2303_;
 wire _2304_;
 wire _2305_;
 wire _2306_;
 wire _2307_;
 wire _2308_;
 wire _2309_;
 wire _2310_;
 wire _2311_;
 wire _2312_;
 wire _2313_;
 wire _2314_;
 wire _2315_;
 wire _2316_;
 wire _2317_;
 wire _2318_;
 wire _2319_;
 wire _2320_;
 wire _2321_;
 wire _2322_;
 wire _2323_;
 wire _2324_;
 wire _2325_;
 wire _2326_;
 wire _2327_;
 wire _2328_;
 wire _2329_;
 wire _2330_;
 wire _2331_;
 wire _2332_;
 wire _2333_;
 wire _2334_;
 wire _2335_;
 wire _2336_;
 wire _2337_;
 wire _2338_;
 wire _2339_;
 wire _2340_;
 wire _2341_;
 wire _2342_;
 wire _2343_;
 wire _2344_;
 wire _2345_;
 wire _2346_;
 wire _2347_;
 wire _2348_;
 wire _2349_;
 wire _2350_;
 wire _2351_;
 wire _2352_;
 wire _2353_;
 wire _2354_;
 wire _2355_;
 wire _2356_;
 wire _2357_;
 wire _2358_;
 wire _2359_;
 wire _2360_;
 wire _2361_;
 wire _2362_;
 wire _2363_;
 wire _2364_;
 wire _2365_;
 wire _2366_;
 wire _2367_;
 wire _2368_;
 wire _2369_;
 wire _2370_;
 wire _2371_;
 wire _2372_;
 wire _2373_;
 wire _2374_;
 wire _2375_;
 wire _2376_;
 wire _2377_;
 wire _2378_;
 wire _2379_;
 wire _2380_;
 wire _2381_;
 wire _2382_;
 wire _2383_;
 wire _2384_;
 wire _2385_;
 wire _2386_;
 wire _2387_;
 wire _2388_;
 wire _2389_;
 wire _2390_;
 wire _2391_;
 wire _2392_;
 wire _2393_;
 wire _2394_;
 wire _2395_;
 wire _2396_;
 wire _2397_;
 wire _2398_;
 wire _2399_;
 wire _2400_;
 wire _2401_;
 wire _2402_;
 wire _2403_;
 wire _2404_;
 wire _2405_;
 wire _2406_;
 wire _2407_;
 wire _2408_;
 wire _2409_;
 wire _2410_;
 wire _2411_;
 wire _2412_;
 wire _2413_;
 wire _2414_;
 wire _2415_;
 wire _2416_;
 wire _2417_;
 wire _2418_;
 wire _2419_;
 wire _2420_;
 wire _2421_;
 wire _2422_;
 wire _2423_;
 wire _2424_;
 wire _2425_;
 wire _2426_;
 wire _2427_;
 wire _2428_;
 wire _2429_;
 wire _2430_;
 wire _2431_;
 wire _2432_;
 wire _2433_;
 wire _2434_;
 wire _2435_;
 wire _2436_;
 wire _2437_;
 wire _2438_;
 wire _2439_;
 wire _2440_;
 wire _2441_;
 wire _2442_;
 wire _2443_;
 wire _2444_;
 wire _2445_;
 wire _2446_;
 wire _2447_;
 wire _2448_;
 wire _2449_;
 wire _2450_;
 wire _2451_;
 wire _2452_;
 wire _2453_;
 wire _2454_;
 wire _2455_;
 wire _2456_;
 wire _2457_;
 wire _2458_;
 wire _2459_;
 wire _2460_;
 wire _2461_;
 wire _2462_;
 wire _2463_;
 wire _2464_;
 wire _2465_;
 wire _2466_;
 wire _2467_;
 wire _2468_;
 wire _2469_;
 wire _2470_;
 wire _2471_;
 wire _2472_;
 wire _2473_;
 wire _2474_;
 wire _2475_;
 wire _2476_;
 wire _2477_;
 wire _2478_;
 wire _2479_;
 wire _2480_;
 wire _2481_;
 wire _2482_;
 wire _2483_;
 wire _2484_;
 wire _2485_;
 wire _2486_;
 wire _2487_;
 wire _2488_;
 wire _2489_;
 wire _2490_;
 wire _2491_;
 wire _2492_;
 wire _2493_;
 wire _2494_;
 wire _2495_;
 wire _2496_;
 wire _2497_;
 wire _2498_;
 wire _2499_;
 wire _2500_;
 wire _2501_;
 wire _2502_;
 wire _2503_;
 wire _2504_;
 wire _2505_;
 wire _2506_;
 wire _2507_;
 wire _2508_;
 wire _2509_;
 wire _2510_;
 wire _2511_;
 wire _2512_;
 wire _2513_;
 wire _2514_;
 wire _2515_;
 wire _2516_;
 wire _2517_;
 wire _2518_;
 wire _2519_;
 wire _2520_;
 wire _2521_;
 wire _2522_;
 wire _2523_;
 wire _2524_;
 wire _2525_;
 wire _2526_;
 wire _2527_;
 wire _2528_;
 wire _2529_;
 wire _2530_;
 wire _2531_;
 wire _2532_;
 wire _2533_;
 wire _2534_;
 wire _2535_;
 wire _2536_;
 wire _2537_;
 wire _2538_;
 wire _2539_;
 wire _2540_;
 wire _2541_;
 wire _2542_;
 wire _2543_;
 wire _2544_;
 wire _2545_;
 wire _2546_;
 wire _2547_;
 wire _2548_;
 wire _2549_;
 wire _2550_;
 wire _2551_;
 wire _2552_;
 wire _2553_;
 wire _2554_;
 wire _2555_;
 wire _2556_;
 wire _2557_;
 wire _2558_;
 wire _2559_;
 wire _2560_;
 wire _2561_;
 wire _2562_;
 wire _2563_;
 wire _2564_;
 wire _2565_;
 wire _2566_;
 wire _2567_;
 wire _2568_;
 wire _2569_;
 wire _2570_;
 wire _2571_;
 wire _2572_;
 wire _2573_;
 wire _2574_;
 wire _2575_;
 wire _2576_;
 wire _2577_;
 wire _2578_;
 wire _2579_;
 wire _2580_;
 wire _2581_;
 wire _2582_;
 wire _2583_;
 wire _2584_;
 wire _2585_;
 wire _2586_;
 wire _2587_;
 wire _2588_;
 wire _2589_;
 wire _2590_;
 wire _2591_;
 wire _2592_;
 wire _2593_;
 wire _2594_;
 wire _2595_;
 wire _2596_;
 wire _2597_;
 wire _2598_;
 wire _2599_;
 wire _2600_;
 wire _2601_;
 wire _2602_;
 wire _2603_;
 wire _2604_;
 wire _2605_;
 wire _2606_;
 wire _2607_;
 wire _2608_;
 wire _2609_;
 wire _2610_;
 wire _2611_;
 wire _2612_;
 wire _2613_;
 wire _2614_;
 wire _2615_;
 wire _2616_;
 wire _2617_;
 wire _2618_;
 wire _2619_;
 wire _2620_;
 wire _2621_;
 wire _2622_;
 wire _2623_;
 wire _2624_;
 wire _2625_;
 wire _2626_;
 wire _2627_;
 wire _2628_;
 wire _2629_;
 wire _2630_;
 wire _2631_;
 wire _2632_;
 wire _2633_;
 wire _2634_;
 wire _2635_;
 wire _2636_;
 wire _2637_;
 wire _2638_;
 wire _2639_;
 wire _2640_;
 wire _2641_;
 wire _2642_;
 wire _2643_;
 wire _2644_;
 wire _2645_;
 wire _2646_;
 wire _2647_;
 wire _2648_;
 wire _2649_;
 wire _2650_;
 wire _2651_;
 wire _2652_;
 wire _2653_;
 wire _2654_;
 wire _2655_;
 wire _2656_;
 wire _2657_;
 wire _2658_;
 wire _2659_;
 wire _2660_;
 wire _2661_;
 wire _2662_;
 wire _2663_;
 wire _2664_;
 wire _2665_;
 wire _2666_;
 wire _2667_;
 wire _2668_;
 wire _2669_;
 wire _2670_;
 wire _2671_;
 wire _2672_;
 wire _2673_;
 wire _2674_;
 wire _2675_;
 wire _2676_;
 wire _2677_;
 wire _2678_;
 wire _2679_;
 wire _2680_;
 wire _2681_;
 wire _2682_;
 wire _2683_;
 wire _2684_;
 wire _2685_;
 wire _2686_;
 wire _2687_;
 wire _2688_;
 wire _2689_;
 wire _2690_;
 wire _2691_;
 wire _2692_;
 wire _2693_;
 wire _2694_;
 wire _2695_;
 wire _2696_;
 wire _2697_;
 wire _2698_;
 wire _2699_;
 wire _2700_;
 wire _2701_;
 wire _2702_;
 wire _2703_;
 wire _2704_;
 wire _2705_;
 wire _2706_;
 wire _2707_;
 wire _2708_;
 wire _2709_;
 wire _2710_;
 wire _2711_;
 wire _2712_;
 wire _2713_;
 wire _2714_;
 wire _2715_;
 wire _2716_;
 wire _2717_;
 wire _2718_;
 wire _2719_;
 wire _2720_;
 wire _2721_;
 wire _2722_;
 wire _2723_;
 wire _2724_;
 wire _2725_;
 wire _2726_;
 wire _2727_;
 wire _2728_;
 wire _2729_;
 wire _2730_;
 wire _2731_;
 wire _2732_;
 wire _2733_;
 wire _2734_;
 wire _2735_;
 wire _2736_;
 wire _2737_;
 wire _2738_;
 wire _2739_;
 wire _2740_;
 wire _2741_;
 wire _2742_;
 wire _2743_;
 wire _2744_;
 wire _2745_;
 wire _2746_;
 wire _2747_;
 wire _2748_;
 wire _2749_;
 wire _2750_;
 wire _2751_;
 wire _2752_;
 wire _2753_;
 wire _2754_;
 wire _2755_;
 wire _2756_;
 wire _2757_;
 wire _2758_;
 wire _2759_;
 wire _2760_;
 wire _2761_;
 wire _2762_;
 wire _2763_;
 wire _2764_;
 wire _2765_;
 wire _2766_;
 wire _2767_;
 wire _2768_;
 wire _2769_;
 wire _2770_;
 wire _2771_;
 wire _2772_;
 wire _2773_;
 wire _2774_;
 wire _2775_;
 wire _2776_;
 wire _2777_;
 wire _2778_;
 wire _2779_;
 wire _2780_;
 wire _2781_;
 wire _2782_;
 wire _2783_;
 wire _2784_;
 wire _2785_;
 wire _2786_;
 wire _2787_;
 wire _2788_;
 wire _2789_;
 wire _2790_;
 wire _2791_;
 wire _2792_;
 wire _2793_;
 wire _2794_;
 wire _2795_;
 wire _2796_;
 wire _2797_;
 wire _2798_;
 wire _2799_;
 wire _2800_;
 wire _2801_;
 wire _2802_;
 wire _2803_;
 wire _2804_;
 wire _2805_;
 wire _2806_;
 wire _2807_;
 wire _2808_;
 wire _2809_;
 wire _2810_;
 wire _2811_;
 wire _2812_;
 wire _2813_;
 wire _2814_;
 wire _2815_;
 wire _2816_;
 wire _2817_;
 wire _2818_;
 wire _2819_;
 wire _2820_;
 wire _2821_;
 wire _2822_;
 wire _2823_;
 wire _2824_;
 wire _2825_;
 wire _2826_;
 wire _2827_;
 wire _2828_;
 wire _2829_;
 wire _2830_;
 wire _2831_;
 wire _2832_;
 wire _2833_;
 wire _2834_;
 wire _2835_;
 wire _2836_;
 wire _2837_;
 wire _2838_;
 wire _2839_;
 wire _2840_;
 wire _2841_;
 wire _2842_;
 wire _2843_;
 wire _2844_;
 wire _2845_;
 wire _2846_;
 wire _2847_;
 wire _2848_;
 wire _2849_;
 wire _2850_;
 wire _2851_;
 wire _2852_;
 wire _2853_;
 wire _2854_;
 wire _2855_;
 wire _2856_;
 wire _2857_;
 wire _2858_;
 wire _2859_;
 wire _2860_;
 wire _2861_;
 wire _2862_;
 wire _2863_;
 wire _2864_;
 wire _2865_;
 wire _2866_;
 wire _2867_;
 wire _2868_;
 wire _2869_;
 wire _2870_;
 wire _2871_;
 wire _2872_;
 wire _2873_;
 wire _2874_;
 wire _2875_;
 wire _2876_;
 wire _2877_;
 wire _2878_;
 wire _2879_;
 wire _2880_;
 wire _2881_;
 wire _2882_;
 wire _2883_;
 wire _2884_;
 wire _2885_;
 wire _2886_;
 wire _2887_;
 wire _2888_;
 wire _2889_;
 wire _2890_;
 wire _2891_;
 wire _2892_;
 wire _2893_;
 wire _2894_;
 wire _2895_;
 wire _2896_;
 wire _2897_;
 wire _2898_;
 wire _2899_;
 wire _2900_;
 wire _2901_;
 wire _2902_;
 wire _2903_;
 wire _2904_;
 wire _2905_;
 wire _2906_;
 wire _2907_;
 wire _2908_;
 wire _2909_;
 wire _2910_;
 wire _2911_;
 wire _2912_;
 wire _2913_;
 wire _2914_;
 wire _2915_;
 wire _2916_;
 wire _2917_;
 wire _2918_;
 wire _2919_;
 wire _2920_;
 wire _2921_;
 wire _2922_;
 wire _2923_;
 wire _2924_;
 wire _2925_;
 wire _2926_;
 wire _2927_;
 wire _2928_;
 wire _2929_;
 wire _2930_;
 wire _2931_;
 wire _2932_;
 wire _2933_;
 wire _2934_;
 wire _2935_;
 wire _2936_;
 wire _2937_;
 wire _2938_;
 wire _2939_;
 wire _2940_;
 wire _2941_;
 wire _2942_;
 wire _2943_;
 wire _2944_;
 wire _2945_;
 wire _2946_;
 wire _2947_;
 wire _2948_;
 wire _2949_;
 wire _2950_;
 wire _2951_;
 wire _2952_;
 wire _2953_;
 wire _2954_;
 wire _2955_;
 wire _2956_;
 wire _2957_;
 wire _2958_;
 wire _2959_;
 wire _2960_;
 wire _2961_;
 wire _2962_;
 wire _2963_;
 wire _2964_;
 wire _2965_;
 wire _2966_;
 wire _2967_;
 wire _2968_;
 wire _2969_;
 wire _2970_;
 wire _2971_;
 wire _2972_;
 wire _2973_;
 wire _2974_;
 wire _2975_;
 wire _2976_;
 wire _2977_;
 wire _2978_;
 wire _2979_;
 wire _2980_;
 wire _2981_;
 wire _2982_;
 wire _2983_;
 wire _2984_;
 wire _2985_;
 wire _2986_;
 wire _2987_;
 wire _2988_;
 wire _2989_;
 wire _2990_;
 wire _2991_;
 wire _2992_;
 wire _2993_;
 wire _2994_;
 wire _2995_;
 wire _2996_;
 wire _2997_;
 wire _2998_;
 wire _2999_;
 wire _3000_;
 wire _3001_;
 wire _3002_;
 wire _3003_;
 wire _3004_;
 wire _3005_;
 wire _3006_;
 wire _3007_;
 wire _3008_;
 wire _3009_;
 wire _3010_;
 wire _3011_;
 wire _3012_;
 wire _3013_;
 wire _3014_;
 wire _3015_;
 wire _3016_;
 wire _3017_;
 wire _3018_;
 wire _3019_;
 wire _3020_;
 wire _3021_;
 wire _3022_;
 wire _3023_;
 wire _3024_;
 wire _3025_;
 wire _3026_;
 wire _3027_;
 wire _3028_;
 wire _3029_;
 wire _3030_;
 wire _3031_;
 wire _3032_;
 wire _3033_;
 wire _3034_;
 wire _3035_;
 wire _3036_;
 wire _3037_;
 wire _3038_;
 wire _3039_;
 wire _3040_;
 wire _3041_;
 wire _3042_;
 wire _3043_;
 wire _3044_;
 wire _3045_;
 wire _3046_;
 wire _3047_;
 wire _3048_;
 wire _3049_;
 wire _3050_;
 wire _3051_;
 wire _3052_;
 wire _3053_;
 wire _3054_;
 wire _3055_;
 wire _3056_;
 wire _3057_;
 wire _3058_;
 wire _3059_;
 wire _3060_;
 wire _3061_;
 wire _3062_;
 wire _3063_;
 wire _3064_;
 wire _3065_;
 wire _3066_;
 wire _3067_;
 wire _3068_;
 wire _3069_;
 wire _3070_;
 wire _3071_;
 wire _3072_;
 wire _3073_;
 wire _3074_;
 wire _3075_;
 wire _3076_;
 wire _3077_;
 wire _3078_;
 wire _3079_;
 wire _3080_;
 wire _3081_;
 wire _3082_;
 wire _3083_;
 wire _3084_;
 wire _3085_;
 wire _3086_;
 wire _3087_;
 wire _3088_;
 wire _3089_;
 wire _3090_;
 wire _3091_;
 wire _3092_;
 wire _3093_;
 wire _3094_;
 wire _3095_;
 wire _3096_;
 wire _3097_;
 wire _3098_;
 wire _3099_;
 wire _3100_;
 wire _3101_;
 wire _3102_;
 wire _3103_;
 wire _3104_;
 wire _3105_;
 wire _3106_;
 wire _3107_;
 wire _3108_;
 wire _3109_;
 wire _3110_;
 wire _3111_;
 wire _3112_;
 wire _3113_;
 wire _3114_;
 wire _3115_;
 wire _3116_;
 wire _3117_;
 wire _3118_;
 wire _3119_;
 wire _3120_;
 wire _3121_;
 wire _3122_;
 wire _3123_;
 wire _3124_;
 wire _3125_;
 wire _3126_;
 wire _3127_;
 wire _3128_;
 wire _3129_;
 wire _3130_;
 wire _3131_;
 wire _3132_;
 wire _3133_;
 wire _3134_;
 wire _3135_;
 wire _3136_;
 wire _3137_;
 wire _3138_;
 wire _3139_;
 wire _3140_;
 wire _3141_;
 wire _3142_;
 wire _3143_;
 wire _3144_;
 wire _3145_;
 wire _3146_;
 wire _3147_;
 wire _3148_;
 wire _3149_;
 wire _3150_;
 wire _3151_;
 wire _3152_;
 wire _3153_;
 wire _3154_;
 wire _3155_;
 wire _3156_;
 wire _3157_;
 wire _3158_;
 wire _3159_;
 wire _3160_;
 wire _3161_;
 wire _3162_;
 wire _3163_;
 wire _3164_;
 wire _3165_;
 wire _3166_;
 wire _3167_;
 wire _3168_;
 wire _3169_;
 wire _3170_;
 wire _3171_;
 wire _3172_;
 wire _3173_;
 wire _3174_;
 wire _3175_;
 wire _3176_;
 wire _3177_;
 wire _3178_;
 wire _3179_;
 wire _3180_;
 wire _3181_;
 wire _3182_;
 wire _3183_;
 wire _3184_;
 wire _3185_;
 wire _3186_;
 wire _3187_;
 wire _3188_;
 wire _3189_;
 wire _3190_;
 wire _3191_;
 wire _3192_;
 wire _3193_;
 wire _3194_;
 wire _3195_;
 wire _3196_;
 wire _3197_;
 wire _3198_;
 wire _3199_;
 wire _3200_;
 wire _3201_;
 wire _3202_;
 wire _3203_;
 wire _3204_;
 wire _3205_;
 wire _3206_;
 wire _3207_;
 wire _3208_;
 wire _3209_;
 wire _3210_;
 wire _3211_;
 wire _3212_;
 wire _3213_;
 wire _3214_;
 wire _3215_;
 wire _3216_;
 wire _3217_;
 wire _3218_;
 wire _3219_;
 wire _3220_;
 wire _3221_;
 wire _3222_;
 wire _3223_;
 wire _3224_;
 wire _3225_;
 wire _3226_;
 wire _3227_;
 wire _3228_;
 wire _3229_;
 wire _3230_;
 wire _3231_;
 wire _3232_;
 wire _3233_;
 wire _3234_;
 wire _3235_;
 wire _3236_;
 wire _3237_;
 wire _3238_;
 wire _3239_;
 wire _3240_;
 wire _3241_;
 wire _3242_;
 wire _3243_;
 wire _3244_;
 wire _3245_;
 wire _3246_;
 wire _3247_;
 wire _3248_;
 wire _3249_;
 wire _3250_;
 wire _3251_;
 wire _3252_;
 wire _3253_;
 wire _3254_;
 wire _3255_;
 wire _3256_;
 wire _3257_;
 wire _3258_;
 wire _3259_;
 wire _3260_;
 wire _3261_;
 wire _3262_;
 wire _3263_;
 wire _3264_;
 wire _3265_;
 wire _3266_;
 wire _3267_;
 wire _3268_;
 wire _3269_;
 wire _3270_;
 wire _3271_;
 wire _3272_;
 wire _3273_;
 wire _3274_;
 wire _3275_;
 wire _3276_;
 wire _3277_;
 wire _3278_;
 wire _3279_;
 wire _3280_;
 wire _3281_;
 wire _3282_;
 wire _3283_;
 wire _3284_;
 wire _3285_;
 wire _3286_;
 wire _3287_;
 wire _3288_;
 wire _3289_;
 wire _3290_;
 wire _3291_;
 wire _3292_;
 wire _3293_;
 wire _3294_;
 wire _3295_;
 wire _3296_;
 wire _3297_;
 wire _3298_;
 wire _3299_;
 wire _3300_;
 wire _3301_;
 wire _3302_;
 wire _3303_;
 wire _3304_;
 wire _3305_;
 wire _3306_;
 wire _3307_;
 wire _3308_;
 wire _3309_;
 wire _3310_;
 wire _3311_;
 wire _3312_;
 wire _3313_;
 wire _3314_;
 wire _3315_;
 wire _3316_;
 wire _3317_;
 wire _3318_;
 wire _3319_;
 wire _3320_;
 wire _3321_;
 wire _3322_;
 wire _3323_;
 wire _3324_;
 wire _3325_;
 wire _3326_;
 wire _3327_;
 wire _3328_;
 wire _3329_;
 wire _3330_;
 wire _3331_;
 wire _3332_;
 wire _3333_;
 wire _3334_;
 wire _3335_;
 wire _3336_;
 wire _3337_;
 wire _3338_;
 wire _3339_;
 wire _3340_;
 wire _3341_;
 wire _3342_;
 wire _3343_;
 wire _3344_;
 wire _3345_;
 wire _3346_;
 wire _3347_;
 wire _3348_;
 wire _3349_;
 wire _3350_;
 wire _3351_;
 wire _3352_;
 wire _3353_;
 wire _3354_;
 wire _3355_;
 wire _3356_;
 wire _3357_;
 wire _3358_;
 wire _3359_;
 wire _3360_;
 wire _3361_;
 wire _3362_;
 wire _3363_;
 wire _3364_;
 wire _3365_;
 wire _3366_;
 wire _3367_;
 wire _3368_;
 wire _3369_;
 wire _3370_;
 wire _3371_;
 wire _3372_;
 wire _3373_;
 wire _3374_;
 wire _3375_;
 wire _3376_;
 wire _3377_;
 wire _3378_;
 wire _3379_;
 wire _3380_;
 wire _3381_;
 wire _3382_;
 wire _3383_;
 wire _3384_;
 wire _3385_;
 wire _3386_;
 wire _3387_;
 wire _3388_;
 wire _3389_;
 wire _3390_;
 wire _3391_;
 wire _3392_;
 wire _3393_;
 wire _3394_;
 wire _3395_;
 wire _3396_;
 wire _3397_;
 wire _3398_;
 wire _3399_;
 wire _3400_;
 wire _3401_;
 wire _3402_;
 wire _3403_;
 wire _3404_;
 wire _3405_;
 wire _3406_;
 wire _3407_;
 wire _3408_;
 wire _3409_;
 wire _3410_;
 wire _3411_;
 wire _3412_;
 wire _3413_;
 wire _3414_;
 wire _3415_;
 wire _3416_;
 wire _3417_;
 wire _3418_;
 wire _3419_;
 wire _3420_;
 wire _3421_;
 wire _3422_;
 wire _3423_;
 wire _3424_;
 wire _3425_;
 wire _3426_;
 wire _3427_;
 wire _3428_;
 wire _3429_;
 wire _3430_;
 wire _3431_;
 wire _3432_;
 wire _3433_;
 wire _3434_;
 wire _3435_;
 wire _3436_;
 wire _3437_;
 wire _3438_;
 wire _3439_;
 wire _3440_;
 wire _3441_;
 wire _3442_;
 wire _3443_;
 wire _3444_;
 wire _3445_;
 wire _3446_;
 wire _3447_;
 wire _3448_;
 wire _3449_;
 wire _3450_;
 wire _3451_;
 wire _3452_;
 wire _3453_;
 wire _3454_;
 wire _3455_;
 wire _3456_;
 wire _3457_;
 wire _3458_;
 wire _3459_;
 wire _3460_;
 wire _3461_;
 wire _3462_;
 wire _3463_;
 wire _3464_;
 wire _3465_;
 wire _3466_;
 wire _3467_;
 wire _3468_;
 wire _3469_;
 wire _3470_;
 wire _3471_;
 wire _3472_;
 wire _3473_;
 wire _3474_;
 wire _3475_;
 wire _3476_;
 wire _3477_;
 wire _3478_;
 wire _3479_;
 wire _3480_;
 wire _3481_;
 wire _3482_;
 wire _3483_;
 wire _3484_;
 wire _3485_;
 wire _3486_;
 wire _3487_;
 wire _3488_;
 wire _3489_;
 wire _3490_;
 wire _3491_;
 wire _3492_;
 wire _3493_;
 wire _3494_;
 wire _3495_;
 wire _3496_;
 wire _3497_;
 wire _3498_;
 wire _3499_;
 wire _3500_;
 wire _3501_;
 wire _3502_;
 wire _3503_;
 wire _3504_;
 wire _3505_;
 wire _3506_;
 wire _3507_;
 wire _3508_;
 wire _3509_;
 wire _3510_;
 wire _3511_;
 wire _3512_;
 wire _3513_;
 wire _3514_;
 wire _3515_;
 wire _3516_;
 wire _3517_;
 wire _3518_;
 wire _3519_;
 wire _3520_;
 wire _3521_;
 wire _3522_;
 wire _3523_;
 wire _3524_;
 wire _3525_;
 wire _3526_;
 wire _3527_;
 wire _3528_;
 wire _3529_;
 wire _3530_;
 wire _3531_;
 wire _3532_;
 wire _3533_;
 wire _3534_;
 wire _3535_;
 wire _3536_;
 wire _3537_;
 wire _3538_;
 wire _3539_;
 wire _3540_;
 wire _3541_;
 wire _3542_;
 wire _3543_;
 wire _3544_;
 wire _3545_;
 wire _3546_;
 wire _3547_;
 wire _3548_;
 wire _3549_;
 wire _3550_;
 wire _3551_;
 wire _3552_;
 wire _3553_;
 wire _3554_;
 wire _3555_;
 wire _3556_;
 wire _3557_;
 wire _3558_;
 wire _3559_;
 wire _3560_;
 wire _3561_;
 wire _3562_;
 wire _3563_;
 wire _3564_;
 wire _3565_;
 wire _3566_;
 wire _3567_;
 wire _3568_;
 wire _3569_;
 wire _3570_;
 wire _3571_;
 wire _3572_;
 wire _3573_;
 wire _3574_;
 wire _3575_;
 wire _3576_;
 wire _3577_;
 wire _3578_;
 wire _3579_;
 wire _3580_;
 wire _3581_;
 wire _3582_;
 wire _3583_;
 wire _3584_;
 wire _3585_;
 wire _3586_;
 wire _3587_;
 wire _3588_;
 wire _3589_;
 wire _3590_;
 wire _3591_;
 wire _3592_;
 wire _3593_;
 wire _3594_;
 wire _3595_;
 wire _3596_;
 wire _3597_;
 wire _3598_;
 wire _3599_;
 wire _3600_;
 wire _3601_;
 wire _3602_;
 wire _3603_;
 wire _3604_;
 wire _3605_;
 wire _3606_;
 wire _3607_;
 wire _3608_;
 wire _3609_;
 wire _3610_;
 wire _3611_;
 wire _3612_;
 wire _3613_;
 wire _3614_;
 wire _3615_;
 wire _3616_;
 wire _3617_;
 wire _3618_;
 wire _3619_;
 wire _3620_;
 wire _3621_;
 wire _3622_;
 wire _3623_;
 wire _3624_;
 wire _3625_;
 wire _3626_;
 wire _3627_;
 wire _3628_;
 wire _3629_;
 wire _3630_;
 wire _3631_;
 wire _3632_;
 wire _3633_;
 wire _3634_;
 wire _3635_;
 wire _3636_;
 wire _3637_;
 wire _3638_;
 wire _3639_;
 wire _3640_;
 wire _3641_;
 wire _3642_;
 wire _3643_;
 wire _3644_;
 wire _3645_;
 wire _3646_;
 wire _3647_;
 wire _3648_;
 wire _3649_;
 wire _3650_;
 wire _3651_;
 wire _3652_;
 wire _3653_;
 wire _3654_;
 wire _3655_;
 wire _3656_;
 wire _3657_;
 wire _3658_;
 wire _3659_;
 wire _3660_;
 wire _3661_;
 wire _3662_;
 wire _3663_;
 wire _3664_;
 wire _3665_;
 wire _3666_;
 wire _3667_;
 wire _3668_;
 wire _3669_;
 wire _3670_;
 wire _3671_;
 wire _3672_;
 wire _3673_;
 wire _3674_;
 wire _3675_;
 wire _3676_;
 wire _3677_;
 wire _3678_;
 wire _3679_;
 wire _3680_;
 wire _3681_;
 wire _3682_;
 wire _3683_;
 wire _3684_;
 wire _3685_;
 wire _3686_;
 wire _3687_;
 wire _3688_;
 wire _3689_;
 wire _3690_;
 wire _3691_;
 wire _3692_;
 wire _3693_;
 wire _3694_;
 wire _3695_;
 wire _3696_;
 wire _3697_;
 wire _3698_;
 wire _3699_;
 wire _3700_;
 wire _3701_;
 wire _3702_;
 wire _3703_;
 wire _3704_;
 wire _3705_;
 wire _3706_;
 wire _3707_;
 wire _3708_;
 wire _3709_;
 wire _3710_;
 wire _3711_;
 wire _3712_;
 wire _3713_;
 wire _3714_;
 wire _3715_;
 wire _3716_;
 wire _3717_;
 wire _3718_;
 wire _3719_;
 wire _3720_;
 wire _3721_;
 wire _3722_;
 wire _3723_;
 wire _3724_;
 wire _3725_;
 wire _3726_;
 wire _3727_;
 wire _3728_;
 wire _3729_;
 wire _3730_;
 wire _3731_;
 wire _3732_;
 wire _3733_;
 wire _3734_;
 wire _3735_;
 wire _3736_;
 wire _3737_;
 wire _3738_;
 wire _3739_;
 wire _3740_;
 wire _3741_;
 wire _3742_;
 wire _3743_;
 wire _3744_;
 wire _3745_;
 wire _3746_;
 wire _3747_;
 wire _3748_;
 wire _3749_;
 wire _3750_;
 wire _3751_;
 wire _3752_;
 wire _3753_;
 wire _3754_;
 wire _3755_;
 wire _3756_;
 wire _3757_;
 wire _3758_;
 wire _3759_;
 wire _3760_;
 wire _3761_;
 wire _3762_;
 wire _3763_;
 wire _3764_;
 wire _3765_;
 wire _3766_;
 wire _3767_;
 wire _3768_;
 wire _3769_;
 wire _3770_;
 wire _3771_;
 wire _3772_;
 wire _3773_;
 wire _3774_;
 wire _3775_;
 wire _3776_;
 wire _3777_;
 wire _3778_;
 wire _3779_;
 wire _3780_;
 wire _3781_;
 wire _3782_;
 wire _3783_;
 wire _3784_;
 wire _3785_;
 wire _3786_;
 wire _3787_;
 wire _3788_;
 wire _3789_;
 wire _3790_;
 wire _3791_;
 wire _3792_;
 wire _3793_;
 wire _3794_;
 wire _3795_;
 wire _3796_;
 wire _3797_;
 wire _3798_;
 wire _3799_;
 wire _3800_;
 wire _3801_;
 wire _3802_;
 wire _3803_;
 wire _3804_;
 wire _3805_;
 wire _3806_;
 wire _3807_;
 wire _3808_;
 wire _3809_;
 wire _3810_;
 wire _3811_;
 wire _3812_;
 wire _3813_;
 wire _3814_;
 wire _3815_;
 wire _3816_;
 wire _3817_;
 wire _3818_;
 wire _3819_;
 wire _3820_;
 wire _3821_;
 wire _3822_;
 wire _3823_;
 wire _3824_;
 wire _3825_;
 wire _3826_;
 wire _3827_;
 wire _3828_;
 wire _3829_;
 wire _3830_;
 wire _3831_;
 wire _3832_;
 wire _3833_;
 wire _3834_;
 wire _3835_;
 wire _3836_;
 wire _3837_;
 wire _3838_;
 wire _3839_;
 wire _3840_;
 wire _3841_;
 wire _3842_;
 wire _3843_;
 wire _3844_;
 wire _3845_;
 wire _3846_;
 wire _3847_;
 wire _3848_;
 wire _3849_;
 wire _3850_;
 wire _3851_;
 wire _3852_;
 wire _3853_;
 wire _3854_;
 wire _3855_;
 wire _3856_;
 wire _3857_;
 wire _3858_;
 wire _3859_;
 wire _3860_;
 wire _3861_;
 wire _3862_;
 wire _3863_;
 wire _3864_;
 wire _3865_;
 wire _3866_;
 wire _3867_;
 wire _3868_;
 wire _3869_;
 wire _3870_;
 wire _3871_;
 wire _3872_;
 wire _3873_;
 wire _3874_;
 wire _3875_;
 wire _3876_;
 wire _3877_;
 wire _3878_;
 wire _3879_;
 wire _3880_;
 wire _3881_;
 wire _3882_;
 wire _3883_;
 wire _3884_;
 wire _3885_;
 wire _3886_;
 wire _3887_;
 wire _3888_;
 wire _3889_;
 wire _3890_;
 wire _3891_;
 wire _3892_;
 wire _3893_;
 wire _3894_;
 wire _3895_;
 wire _3896_;
 wire _3897_;
 wire _3898_;
 wire _3899_;
 wire _3900_;
 wire _3901_;
 wire _3902_;
 wire _3903_;
 wire _3904_;
 wire _3905_;
 wire _3906_;
 wire _3907_;
 wire _3908_;
 wire _3909_;
 wire _3910_;
 wire _3911_;
 wire _3912_;
 wire _3913_;
 wire _3914_;
 wire _3915_;
 wire _3916_;
 wire _3917_;
 wire _3918_;
 wire _3919_;
 wire _3920_;
 wire _3921_;
 wire _3922_;
 wire _3923_;
 wire _3924_;
 wire _3925_;
 wire _3926_;
 wire _3927_;
 wire _3928_;
 wire _3929_;
 wire _3930_;
 wire _3931_;
 wire _3932_;
 wire _3933_;
 wire _3934_;
 wire _3935_;
 wire _3936_;
 wire _3937_;
 wire _3938_;
 wire _3939_;
 wire _3940_;
 wire _3941_;
 wire _3942_;
 wire _3943_;
 wire _3944_;
 wire _3945_;
 wire _3946_;
 wire _3947_;
 wire _3948_;
 wire _3949_;
 wire _3950_;
 wire _3951_;
 wire _3952_;
 wire _3953_;
 wire _3954_;
 wire _3955_;
 wire _3956_;
 wire _3957_;
 wire _3958_;
 wire _3959_;
 wire _3960_;
 wire _3961_;
 wire _3962_;
 wire _3963_;
 wire _3964_;
 wire _3965_;
 wire _3966_;
 wire _3967_;
 wire _3968_;
 wire _3969_;
 wire _3970_;
 wire _3971_;
 wire _3972_;
 wire _3973_;
 wire _3974_;
 wire _3975_;
 wire _3976_;
 wire _3977_;
 wire _3978_;
 wire _3979_;
 wire _3980_;
 wire _3981_;
 wire _3982_;
 wire _3983_;
 wire _3984_;
 wire _3985_;
 wire _3986_;
 wire _3987_;
 wire _3988_;
 wire _3989_;
 wire _3990_;
 wire _3991_;
 wire _3992_;
 wire _3993_;
 wire _3994_;
 wire _3995_;
 wire _3996_;
 wire _3997_;
 wire _3998_;
 wire _3999_;
 wire _4000_;
 wire _4001_;
 wire _4002_;
 wire _4003_;
 wire _4004_;
 wire _4005_;
 wire _4006_;
 wire _4007_;
 wire _4008_;
 wire _4009_;
 wire _4010_;
 wire _4011_;
 wire _4012_;
 wire _4013_;
 wire _4014_;
 wire _4015_;
 wire _4016_;
 wire _4017_;
 wire _4018_;
 wire _4019_;
 wire _4020_;
 wire _4021_;
 wire _4022_;
 wire _4023_;
 wire _4024_;
 wire _4025_;
 wire _4026_;
 wire _4027_;
 wire _4028_;
 wire _4029_;
 wire _4030_;
 wire _4031_;
 wire _4032_;
 wire _4033_;
 wire _4034_;
 wire _4035_;
 wire _4036_;
 wire _4037_;
 wire _4038_;
 wire _4039_;
 wire _4040_;
 wire _4041_;
 wire _4042_;
 wire _4043_;
 wire _4044_;
 wire _4045_;
 wire _4046_;
 wire _4047_;
 wire _4048_;
 wire _4049_;
 wire _4050_;
 wire _4051_;
 wire _4052_;
 wire _4053_;
 wire _4054_;
 wire _4055_;
 wire _4056_;
 wire _4057_;
 wire _4058_;
 wire _4059_;
 wire _4060_;
 wire _4061_;
 wire _4062_;
 wire _4063_;
 wire _4064_;
 wire _4065_;
 wire _4066_;
 wire _4067_;
 wire _4068_;
 wire _4069_;
 wire _4070_;
 wire _4071_;
 wire _4072_;
 wire _4073_;
 wire _4074_;
 wire _4075_;
 wire _4076_;
 wire _4077_;
 wire _4078_;
 wire _4079_;
 wire _4080_;
 wire _4081_;
 wire _4082_;
 wire _4083_;
 wire _4084_;
 wire _4085_;
 wire _4086_;
 wire _4087_;
 wire _4088_;
 wire _4089_;
 wire _4090_;
 wire _4091_;
 wire _4092_;
 wire _4093_;
 wire _4094_;
 wire _4095_;
 wire _4096_;
 wire _4097_;
 wire _4098_;
 wire _4099_;
 wire _4100_;
 wire _4101_;
 wire _4102_;
 wire _4103_;
 wire _4104_;
 wire _4105_;
 wire _4106_;
 wire _4107_;
 wire _4108_;
 wire _4109_;
 wire _4110_;
 wire _4111_;
 wire _4112_;
 wire _4113_;
 wire _4114_;
 wire _4115_;
 wire _4116_;
 wire _4117_;
 wire _4118_;
 wire _4119_;
 wire _4120_;
 wire _4121_;
 wire _4122_;
 wire _4123_;
 wire _4124_;
 wire _4125_;
 wire _4126_;
 wire _4127_;
 wire _4128_;
 wire _4129_;
 wire _4130_;
 wire _4131_;
 wire _4132_;
 wire _4133_;
 wire _4134_;
 wire _4135_;
 wire _4136_;
 wire _4137_;
 wire _4138_;
 wire _4139_;
 wire _4140_;
 wire _4141_;
 wire _4142_;
 wire _4143_;
 wire _4144_;
 wire _4145_;
 wire _4146_;
 wire _4147_;
 wire _4148_;
 wire _4149_;
 wire _4150_;
 wire _4151_;
 wire _4152_;
 wire _4153_;
 wire _4154_;
 wire _4155_;
 wire _4156_;
 wire _4157_;
 wire _4158_;
 wire _4159_;
 wire _4160_;
 wire _4161_;
 wire _4162_;
 wire _4163_;
 wire _4164_;
 wire _4165_;
 wire _4166_;
 wire _4167_;
 wire _4168_;
 wire _4169_;
 wire _4170_;
 wire _4171_;
 wire _4172_;
 wire _4173_;
 wire _4174_;
 wire _4175_;
 wire _4176_;
 wire _4177_;
 wire _4178_;
 wire _4179_;
 wire _4180_;
 wire _4181_;
 wire _4182_;
 wire _4183_;
 wire _4184_;
 wire _4185_;
 wire _4186_;
 wire _4187_;
 wire _4188_;
 wire _4189_;
 wire _4190_;
 wire _4191_;
 wire _4192_;
 wire _4193_;
 wire _4194_;
 wire _4195_;
 wire _4196_;
 wire _4197_;
 wire _4198_;
 wire _4199_;
 wire _4200_;
 wire _4201_;
 wire _4202_;
 wire _4203_;
 wire _4204_;
 wire _4205_;
 wire _4206_;
 wire _4207_;
 wire _4208_;
 wire _4209_;
 wire _4210_;
 wire _4211_;
 wire _4212_;
 wire _4213_;
 wire _4214_;
 wire _4215_;
 wire _4216_;
 wire _4217_;
 wire _4218_;
 wire _4219_;
 wire _4220_;
 wire _4221_;
 wire _4222_;
 wire _4223_;
 wire _4224_;
 wire _4225_;
 wire _4226_;
 wire _4227_;
 wire _4228_;
 wire _4229_;
 wire _4230_;
 wire _4231_;
 wire _4232_;
 wire _4233_;
 wire _4234_;
 wire _4235_;
 wire _4236_;
 wire _4237_;
 wire _4238_;
 wire _4239_;
 wire _4240_;
 wire _4241_;
 wire _4242_;
 wire _4243_;
 wire _4244_;
 wire _4245_;
 wire _4246_;
 wire _4247_;
 wire _4248_;
 wire _4249_;
 wire _4250_;
 wire _4251_;
 wire _4252_;
 wire _4253_;
 wire _4254_;
 wire _4255_;
 wire _4256_;
 wire _4257_;
 wire _4258_;
 wire _4259_;
 wire _4260_;
 wire _4261_;
 wire _4262_;
 wire _4263_;
 wire _4264_;
 wire _4265_;
 wire _4266_;
 wire _4267_;
 wire _4268_;
 wire _4269_;
 wire _4270_;
 wire _4271_;
 wire _4272_;
 wire _4273_;
 wire _4274_;
 wire _4275_;
 wire _4276_;
 wire _4277_;
 wire _4278_;
 wire _4279_;
 wire _4280_;
 wire _4281_;
 wire _4282_;
 wire _4283_;
 wire _4284_;
 wire _4285_;
 wire _4286_;
 wire _4287_;
 wire _4288_;
 wire _4289_;
 wire _4290_;
 wire _4291_;
 wire _4292_;
 wire _4293_;
 wire _4294_;
 wire _4295_;
 wire _4296_;
 wire _4297_;
 wire _4298_;
 wire _4299_;
 wire _4300_;
 wire _4301_;
 wire _4302_;
 wire _4303_;
 wire _4304_;
 wire _4305_;
 wire _4306_;
 wire _4307_;
 wire _4308_;
 wire _4309_;
 wire _4310_;
 wire _4311_;
 wire _4312_;
 wire _4313_;
 wire _4314_;
 wire _4315_;
 wire _4316_;
 wire _4317_;
 wire _4318_;
 wire _4319_;
 wire _4320_;
 wire _4321_;
 wire _4322_;
 wire _4323_;
 wire _4324_;
 wire _4325_;
 wire _4326_;
 wire _4327_;
 wire _4328_;
 wire _4329_;
 wire _4330_;
 wire _4331_;
 wire _4332_;
 wire _4333_;
 wire _4334_;
 wire _4335_;
 wire _4336_;
 wire _4337_;
 wire _4338_;
 wire _4339_;
 wire _4340_;
 wire _4341_;
 wire _4342_;
 wire _4343_;
 wire _4344_;
 wire _4345_;
 wire _4346_;
 wire _4347_;
 wire _4348_;
 wire _4349_;
 wire _4350_;
 wire _4351_;
 wire _4352_;
 wire _4353_;
 wire _4354_;
 wire _4355_;
 wire _4356_;
 wire _4357_;
 wire _4358_;
 wire _4359_;
 wire _4360_;
 wire _4361_;
 wire _4362_;
 wire _4363_;
 wire _4364_;
 wire _4365_;
 wire _4366_;
 wire _4367_;
 wire _4368_;
 wire _4369_;
 wire _4370_;
 wire _4371_;
 wire _4372_;
 wire _4373_;
 wire _4374_;
 wire _4375_;
 wire _4376_;
 wire _4377_;
 wire _4378_;
 wire _4379_;
 wire _4380_;
 wire _4381_;
 wire _4382_;
 wire _4383_;
 wire _4384_;
 wire _4385_;
 wire _4386_;
 wire _4387_;
 wire _4388_;
 wire _4389_;
 wire _4390_;
 wire _4391_;
 wire _4392_;
 wire _4393_;
 wire _4394_;
 wire _4395_;
 wire _4396_;
 wire _4397_;
 wire _4398_;
 wire _4399_;
 wire _4400_;
 wire _4401_;
 wire _4402_;
 wire _4403_;
 wire _4404_;
 wire _4405_;
 wire _4406_;
 wire _4407_;
 wire _4408_;
 wire _4409_;
 wire _4410_;
 wire _4411_;
 wire _4412_;
 wire _4413_;
 wire _4414_;
 wire _4415_;
 wire _4416_;
 wire _4417_;
 wire _4418_;
 wire _4419_;
 wire _4420_;
 wire _4421_;
 wire _4422_;
 wire _4423_;
 wire _4424_;
 wire _4425_;
 wire _4426_;
 wire _4427_;
 wire _4428_;
 wire _4429_;
 wire _4430_;
 wire _4431_;
 wire _4432_;
 wire _4433_;
 wire _4434_;
 wire _4435_;
 wire _4436_;
 wire _4437_;
 wire _4438_;
 wire _4439_;
 wire _4440_;
 wire _4441_;
 wire _4442_;
 wire _4443_;
 wire _4444_;
 wire _4445_;
 wire _4446_;
 wire _4447_;
 wire _4448_;
 wire _4449_;
 wire _4450_;
 wire _4451_;
 wire _4452_;
 wire _4453_;
 wire _4454_;
 wire _4455_;
 wire _4456_;
 wire _4457_;
 wire _4458_;
 wire _4459_;
 wire _4460_;
 wire _4461_;
 wire _4462_;
 wire _4463_;
 wire _4464_;
 wire _4465_;
 wire _4466_;
 wire _4467_;
 wire _4468_;
 wire _4469_;
 wire _4470_;
 wire _4471_;
 wire _4472_;
 wire _4473_;
 wire _4474_;
 wire _4475_;
 wire _4476_;
 wire _4477_;
 wire _4478_;
 wire _4479_;
 wire _4480_;
 wire _4481_;
 wire _4482_;
 wire _4483_;
 wire _4484_;
 wire _4485_;
 wire _4486_;
 wire _4487_;
 wire _4488_;
 wire _4489_;
 wire _4490_;
 wire _4491_;
 wire _4492_;
 wire _4493_;
 wire _4494_;
 wire _4495_;
 wire _4496_;
 wire _4497_;
 wire _4498_;
 wire _4499_;
 wire _4500_;
 wire _4501_;
 wire _4502_;
 wire _4503_;
 wire _4504_;
 wire _4505_;
 wire _4506_;
 wire _4507_;
 wire _4508_;
 wire _4509_;
 wire _4510_;
 wire _4511_;
 wire _4512_;
 wire _4513_;
 wire _4514_;
 wire _4515_;
 wire _4516_;
 wire _4517_;
 wire _4518_;
 wire _4519_;
 wire _4520_;
 wire _4521_;
 wire _4522_;
 wire _4523_;
 wire _4524_;
 wire _4525_;
 wire _4526_;
 wire _4527_;
 wire _4528_;
 wire _4529_;
 wire _4530_;
 wire _4531_;
 wire _4532_;
 wire _4533_;
 wire _4534_;
 wire _4535_;
 wire _4536_;
 wire _4537_;
 wire _4538_;
 wire _4539_;
 wire _4540_;
 wire _4541_;
 wire _4542_;
 wire _4543_;
 wire _4544_;
 wire _4545_;
 wire _4546_;
 wire _4547_;
 wire _4548_;
 wire _4549_;
 wire _4550_;
 wire _4551_;
 wire _4552_;
 wire _4553_;
 wire _4554_;
 wire _4555_;
 wire _4556_;
 wire _4557_;
 wire _4558_;
 wire _4559_;
 wire _4560_;
 wire _4561_;
 wire _4562_;
 wire _4563_;
 wire _4564_;
 wire _4565_;
 wire _4566_;
 wire _4567_;
 wire _4568_;
 wire _4569_;
 wire _4570_;
 wire _4571_;
 wire _4572_;
 wire _4573_;
 wire _4574_;
 wire _4575_;
 wire _4576_;
 wire _4577_;
 wire _4578_;
 wire _4579_;
 wire _4580_;
 wire _4581_;
 wire _4582_;
 wire _4583_;
 wire _4584_;
 wire _4585_;
 wire _4586_;
 wire _4587_;
 wire _4588_;
 wire _4589_;
 wire _4590_;
 wire _4591_;
 wire _4592_;
 wire _4593_;
 wire _4594_;
 wire _4595_;
 wire _4596_;
 wire _4597_;
 wire _4598_;
 wire _4599_;
 wire _4600_;
 wire _4601_;
 wire _4602_;
 wire _4603_;
 wire _4604_;
 wire _4605_;
 wire _4606_;
 wire _4607_;
 wire _4608_;
 wire _4609_;
 wire _4610_;
 wire _4611_;
 wire _4612_;
 wire _4613_;
 wire _4614_;
 wire _4615_;
 wire _4616_;
 wire _4617_;
 wire _4618_;
 wire _4619_;
 wire _4620_;
 wire _4621_;
 wire _4622_;
 wire _4623_;
 wire _4624_;
 wire _4625_;
 wire _4626_;
 wire _4627_;
 wire _4628_;
 wire _4629_;
 wire _4630_;
 wire _4631_;
 wire _4632_;
 wire clknet_leaf_0_clk;
 wire net122;
 wire \generated._1019[3] ;
 wire \generated._1019[4] ;
 wire \generated._1019[5] ;
 wire \generated._1019[6] ;
 wire \generated._1019[7] ;
 wire \generated._1019[8] ;
 wire \generated._1019[9] ;
 wire \generated._1020[0] ;
 wire \generated._1020[1] ;
 wire \generated._1020[2] ;
 wire \generated._1020[3] ;
 wire \generated._1020[4] ;
 wire \generated._1020[5] ;
 wire \generated._1020[6] ;
 wire \generated._1020[7] ;
 wire \generated._1020[8] ;
 wire \generated._1020[9] ;
 wire \generated._1021[0] ;
 wire \generated._1037[0] ;
 wire \generated._1069[3] ;
 wire \generated._1069[4] ;
 wire \generated._1069[5] ;
 wire \generated._1069[6] ;
 wire \generated._1069[7] ;
 wire \generated._1069[8] ;
 wire \generated._1069[9] ;
 wire \generated._1070[0] ;
 wire \generated._1070[1] ;
 wire \generated._1070[2] ;
 wire \generated._1070[3] ;
 wire \generated._1070[4] ;
 wire \generated._1070[5] ;
 wire \generated._1070[6] ;
 wire \generated._1070[7] ;
 wire \generated._1070[8] ;
 wire \generated._1070[9] ;
 wire \generated._1073[0] ;
 wire \generated._1073[1] ;
 wire \generated._1073[2] ;
 wire \generated._1073[3] ;
 wire \generated._1074[0] ;
 wire \generated._1074[1] ;
 wire \generated._1074[2] ;
 wire \generated._1074[3] ;
 wire \generated._108 ;
 wire \generated._1080[0] ;
 wire \generated._1080[1] ;
 wire \generated._1080[2] ;
 wire \generated._1080[3] ;
 wire \generated._1080[4] ;
 wire \generated._1080[5] ;
 wire \generated._1080[6] ;
 wire \generated._1080[7] ;
 wire \generated._1080[8] ;
 wire \generated._1080[9] ;
 wire \generated._1083[0] ;
 wire \generated._111 ;
 wire \generated._1115[0] ;
 wire \generated._1115[1] ;
 wire \generated._1115[2] ;
 wire \generated._1115[3] ;
 wire \generated._1115[4] ;
 wire \generated._1115[5] ;
 wire \generated._1115[6] ;
 wire \generated._1115[7] ;
 wire \generated._1115[8] ;
 wire \generated._1115[9] ;
 wire \generated._1144[0] ;
 wire \generated._1149[0] ;
 wire \generated._1149[1] ;
 wire \generated._118 ;
 wire \generated._119 ;
 wire \generated._14[0] ;
 wire \generated._14[1] ;
 wire \generated._14[2] ;
 wire \generated._14[3] ;
 wire \generated._14[4] ;
 wire \generated._161[4] ;
 wire \generated._19[0] ;
 wire \generated._19[1] ;
 wire \generated._19[2] ;
 wire \generated._19[3] ;
 wire \generated._19[4] ;
 wire \generated._217[0] ;
 wire \generated._217[1] ;
 wire \generated._217[2] ;
 wire \generated._217[3] ;
 wire \generated._231[0] ;
 wire \generated._231[1] ;
 wire \generated._26[0] ;
 wire \generated._26[1] ;
 wire \generated._26[2] ;
 wire \generated._26[3] ;
 wire \generated._284[0] ;
 wire \generated._284[1] ;
 wire \generated._297[0] ;
 wire \generated._31[0] ;
 wire \generated._31[1] ;
 wire \generated._31[2] ;
 wire \generated._31[3] ;
 wire \generated._31[4] ;
 wire \generated._31[5] ;
 wire \generated._31[6] ;
 wire \generated._324[0] ;
 wire \generated._342[0] ;
 wire \generated._342[1] ;
 wire \generated._342[2] ;
 wire \generated._342[3] ;
 wire \generated._342[4] ;
 wire \generated._342[5] ;
 wire \generated._349[0] ;
 wire \generated._353[0] ;
 wire \generated._353[1] ;
 wire \generated._353[2] ;
 wire \generated._353[3] ;
 wire \generated._353[4] ;
 wire \generated._367 ;
 wire \generated._369[0] ;
 wire \generated._369[1] ;
 wire \generated._369[2] ;
 wire \generated._369[3] ;
 wire \generated._369[4] ;
 wire \generated._369[5] ;
 wire \generated._369[6] ;
 wire \generated._369[7] ;
 wire \generated._369[8] ;
 wire \generated._374 ;
 wire \generated._375 ;
 wire \generated._376 ;
 wire \generated._377[0] ;
 wire \generated._377[1] ;
 wire \generated._377[2] ;
 wire \generated._377[3] ;
 wire \generated._377[4] ;
 wire \generated._377[5] ;
 wire \generated._377[6] ;
 wire \generated._377[7] ;
 wire \generated._390[0] ;
 wire \generated._390[1] ;
 wire \generated._390[2] ;
 wire \generated._390[3] ;
 wire \generated._390[4] ;
 wire \generated._390[5] ;
 wire \generated._390[6] ;
 wire \generated._390[7] ;
 wire \generated._390[8] ;
 wire \generated._390[9] ;
 wire \generated._391[0] ;
 wire \generated._402[1] ;
 wire \generated._402[2] ;
 wire \generated._402[3] ;
 wire \generated._402[4] ;
 wire \generated._402[5] ;
 wire \generated._402[6] ;
 wire \generated._402[7] ;
 wire \generated._421[1] ;
 wire \generated._430[10] ;
 wire \generated._430[11] ;
 wire \generated._430[12] ;
 wire \generated._430[13] ;
 wire \generated._430[14] ;
 wire \generated._430[15] ;
 wire \generated._430[16] ;
 wire \generated._430[17] ;
 wire \generated._430[18] ;
 wire \generated._430[19] ;
 wire \generated._477[0] ;
 wire \generated._477[1] ;
 wire \generated._477[2] ;
 wire \generated._477[3] ;
 wire \generated._477[4] ;
 wire \generated._477[5] ;
 wire \generated._477[6] ;
 wire \generated._477[7] ;
 wire \generated._477[8] ;
 wire \generated._477[9] ;
 wire \generated._482[0] ;
 wire \generated._482[1] ;
 wire \generated._482[2] ;
 wire \generated._482[3] ;
 wire \generated._483[0] ;
 wire \generated._483[1] ;
 wire \generated._483[2] ;
 wire \generated._483[3] ;
 wire \generated._497[0] ;
 wire \generated._499 ;
 wire \generated._501[0] ;
 wire \generated._501[1] ;
 wire \generated._501[2] ;
 wire \generated._501[3] ;
 wire \generated._501[4] ;
 wire \generated._501[5] ;
 wire \generated._501[6] ;
 wire \generated._501[7] ;
 wire \generated._501[8] ;
 wire \generated._505 ;
 wire \generated._506 ;
 wire \generated._507 ;
 wire \generated._508[0] ;
 wire \generated._508[1] ;
 wire \generated._508[2] ;
 wire \generated._508[3] ;
 wire \generated._508[4] ;
 wire \generated._508[5] ;
 wire \generated._508[6] ;
 wire \generated._508[7] ;
 wire \generated._557[0] ;
 wire \generated._557[1] ;
 wire \generated._557[2] ;
 wire \generated._557[3] ;
 wire \generated._557[4] ;
 wire \generated._557[5] ;
 wire \generated._557[6] ;
 wire \generated._557[7] ;
 wire \generated._557[8] ;
 wire \generated._557[9] ;
 wire \generated._558[0] ;
 wire \generated._558[1] ;
 wire \generated._558[2] ;
 wire \generated._558[3] ;
 wire \generated._558[4] ;
 wire \generated._558[5] ;
 wire \generated._558[6] ;
 wire \generated._558[7] ;
 wire \generated._558[8] ;
 wire \generated._558[9] ;
 wire \generated._559[0] ;
 wire \generated._568[0] ;
 wire \generated._568[1] ;
 wire \generated._568[2] ;
 wire \generated._568[3] ;
 wire \generated._568[4] ;
 wire \generated._568[5] ;
 wire \generated._568[6] ;
 wire \generated._568[7] ;
 wire \generated._568[8] ;
 wire \generated._568[9] ;
 wire \generated._60[0] ;
 wire \generated._60[1] ;
 wire \generated._60[2] ;
 wire \generated._60[3] ;
 wire \generated._610[0] ;
 wire \generated._610[1] ;
 wire \generated._610[2] ;
 wire \generated._610[3] ;
 wire \generated._610[4] ;
 wire \generated._610[5] ;
 wire \generated._61[0] ;
 wire \generated._61[1] ;
 wire \generated._61[2] ;
 wire \generated._61[3] ;
 wire \generated._62[0] ;
 wire \generated._63[2] ;
 wire \generated._63[3] ;
 wire \generated._63[4] ;
 wire \generated._63[5] ;
 wire \generated._63[6] ;
 wire \generated._64[1] ;
 wire \generated._64[2] ;
 wire \generated._64[3] ;
 wire \generated._64[4] ;
 wire \generated._64[5] ;
 wire \generated._64[6] ;
 wire \generated._64[7] ;
 wire \generated._64[8] ;
 wire \generated._64[9] ;
 wire \generated._67[0] ;
 wire \generated._67[1] ;
 wire \generated._67[2] ;
 wire \generated._67[3] ;
 wire \generated._67[4] ;
 wire \generated._67[5] ;
 wire \generated._67[6] ;
 wire \generated._67[7] ;
 wire \generated._67[8] ;
 wire \generated._67[9] ;
 wire \generated._68[0] ;
 wire \generated._68[1] ;
 wire \generated._68[2] ;
 wire \generated._68[3] ;
 wire \generated._691[0] ;
 wire \generated._691[1] ;
 wire \generated._691[2] ;
 wire \generated._691[3] ;
 wire \generated._691[4] ;
 wire \generated._691[5] ;
 wire \generated._691[6] ;
 wire \generated._691[7] ;
 wire \generated._691[8] ;
 wire \generated._691[9] ;
 wire \generated._69[0] ;
 wire \generated._69[1] ;
 wire \generated._69[2] ;
 wire \generated._69[3] ;
 wire \generated._75[0] ;
 wire \generated._825[2] ;
 wire \generated._825[3] ;
 wire \generated._825[4] ;
 wire \generated._825[5] ;
 wire \generated._825[6] ;
 wire \generated._825[7] ;
 wire \generated._825[8] ;
 wire \generated._839 ;
 wire \generated._840 ;
 wire \generated._885[3] ;
 wire \generated._885[4] ;
 wire \generated._885[5] ;
 wire \generated._885[6] ;
 wire \generated._885[7] ;
 wire \generated._885[8] ;
 wire \generated._885[9] ;
 wire \generated._887[0] ;
 wire \generated._934[3] ;
 wire \generated._934[4] ;
 wire \generated._934[5] ;
 wire \generated._934[6] ;
 wire \generated._934[7] ;
 wire \generated._934[8] ;
 wire \generated._934[9] ;
 wire \generated._965 ;
 wire \generated._966 ;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net120;
 wire net121;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net180;
 wire net181;
 wire net182;
 wire net183;
 wire net184;
 wire net185;
 wire net186;
 wire net187;
 wire net188;
 wire net189;
 wire net190;
 wire net191;
 wire net192;
 wire net193;
 wire net194;
 wire net195;
 wire net196;
 wire net197;
 wire net198;
 wire net199;
 wire net200;
 wire net201;
 wire net202;
 wire net203;
 wire net204;
 wire net205;
 wire net206;
 wire net207;
 wire net208;
 wire net209;
 wire net210;
 wire net211;
 wire net212;
 wire net213;
 wire net214;
 wire net215;
 wire net216;
 wire net217;
 wire net218;
 wire net219;
 wire net220;
 wire net221;
 wire net222;
 wire net223;
 wire net224;
 wire net225;
 wire net226;
 wire net227;
 wire net228;
 wire net229;
 wire net230;
 wire net231;
 wire net232;
 wire net233;
 wire net234;
 wire net235;
 wire net236;
 wire net237;
 wire net238;
 wire net239;
 wire net240;
 wire net241;
 wire net242;
 wire net243;
 wire net244;
 wire net245;
 wire net246;
 wire net247;
 wire net248;
 wire net249;
 wire net250;
 wire net251;
 wire net252;
 wire net253;
 wire net254;
 wire net255;
 wire net256;
 wire net257;
 wire net258;
 wire net259;
 wire net260;
 wire net261;
 wire net262;
 wire net263;
 wire net264;
 wire net265;
 wire net266;
 wire net267;
 wire net268;
 wire net269;
 wire net270;
 wire net271;
 wire net272;
 wire net273;
 wire net274;
 wire net275;
 wire net276;
 wire net277;
 wire net278;
 wire net279;
 wire net280;
 wire net281;
 wire net282;
 wire net283;
 wire net284;
 wire net285;
 wire net286;
 wire net287;
 wire net288;
 wire net289;
 wire net290;
 wire net291;
 wire clknet_leaf_1_clk;
 wire clknet_leaf_2_clk;
 wire clknet_leaf_3_clk;
 wire clknet_leaf_4_clk;
 wire clknet_leaf_5_clk;
 wire clknet_leaf_6_clk;
 wire clknet_leaf_7_clk;
 wire clknet_leaf_8_clk;
 wire clknet_leaf_9_clk;
 wire clknet_leaf_10_clk;
 wire clknet_leaf_11_clk;
 wire clknet_leaf_12_clk;
 wire clknet_leaf_13_clk;
 wire clknet_leaf_14_clk;
 wire clknet_leaf_15_clk;
 wire clknet_leaf_16_clk;
 wire clknet_leaf_17_clk;
 wire clknet_leaf_19_clk;
 wire clknet_leaf_20_clk;
 wire clknet_leaf_21_clk;
 wire clknet_leaf_22_clk;
 wire clknet_leaf_23_clk;
 wire clknet_leaf_24_clk;
 wire clknet_leaf_25_clk;
 wire clknet_leaf_26_clk;
 wire clknet_leaf_27_clk;
 wire clknet_leaf_28_clk;
 wire clknet_leaf_29_clk;
 wire clknet_leaf_30_clk;
 wire clknet_leaf_31_clk;
 wire clknet_leaf_32_clk;
 wire clknet_leaf_33_clk;
 wire clknet_leaf_34_clk;
 wire clknet_0_clk;
 wire clknet_3_0__leaf_clk;
 wire clknet_3_1__leaf_clk;
 wire clknet_3_2__leaf_clk;
 wire clknet_3_3__leaf_clk;
 wire clknet_3_4__leaf_clk;
 wire clknet_3_5__leaf_clk;
 wire clknet_3_6__leaf_clk;
 wire clknet_3_7__leaf_clk;

 sg13g2_inv_1 _4635_ (.Y(_4147_),
    .A(\generated._14[3] ));
 sg13g2_nor2b_1 _4636_ (.A(\generated._19[1] ),
    .B_N(\generated._19[0] ),
    .Y(_4148_));
 sg13g2_inv_1 _4637_ (.Y(_4149_),
    .A(\generated._19[2] ));
 sg13g2_nand4_1 _4638_ (.B(_4149_),
    .C(\generated._19[3] ),
    .A(_4148_),
    .Y(_4150_),
    .D(\generated._19[4] ));
 sg13g2_buf_2 _4639_ (.A(_4150_),
    .X(_4151_));
 sg13g2_inv_1 _4640_ (.Y(_4152_),
    .A(_4151_));
 sg13g2_buf_1 _4641_ (.A(\generated._14[0] ),
    .X(_4153_));
 sg13g2_nand4_1 _4642_ (.B(\generated._14[1] ),
    .C(_4153_),
    .A(_4152_),
    .Y(_4154_),
    .D(\generated._14[2] ));
 sg13g2_buf_2 _4643_ (.A(\generated._568[5] ),
    .X(_4155_));
 sg13g2_buf_8 _4644_ (.A(\generated._568[7] ),
    .X(_4156_));
 sg13g2_buf_8 _4645_ (.A(\generated._568[6] ),
    .X(_4157_));
 sg13g2_nor3_1 _4646_ (.A(_4155_),
    .B(_4156_),
    .C(_4157_),
    .Y(_4158_));
 sg13g2_buf_8 _4647_ (.A(\generated._568[8] ),
    .X(_4159_));
 sg13g2_inv_8 _4648_ (.Y(_4160_),
    .A(_4159_));
 sg13g2_inv_1 _4649_ (.Y(_4161_),
    .A(\generated._568[9] ));
 sg13g2_buf_8 _4650_ (.A(\generated._568[3] ),
    .X(_4162_));
 sg13g2_buf_1 _4651_ (.A(\generated._568[4] ),
    .X(_4163_));
 sg13g2_nor2_1 _4652_ (.A(_4162_),
    .B(net95),
    .Y(_4164_));
 sg13g2_nand4_1 _4653_ (.B(_4160_),
    .C(_4161_),
    .A(_4158_),
    .Y(_4165_),
    .D(_4164_));
 sg13g2_inv_1 _4654_ (.Y(_4166_),
    .A(_4165_));
 sg13g2_inv_1 _4655_ (.Y(_4167_),
    .A(\generated._568[2] ));
 sg13g2_nor2_1 _4656_ (.A(\generated._568[1] ),
    .B(\generated._568[0] ),
    .Y(_4168_));
 sg13g2_nand3_1 _4657_ (.B(_4167_),
    .C(_4168_),
    .A(_4166_),
    .Y(_4169_));
 sg13g2_buf_2 _4658_ (.A(_4169_),
    .X(_4170_));
 sg13g2_inv_1 _4659_ (.Y(_4171_),
    .A(\generated._14[2] ));
 sg13g2_nand2_1 _4660_ (.Y(_4172_),
    .A(\generated._14[1] ),
    .B(_4153_));
 sg13g2_nor3_1 _4661_ (.A(_4171_),
    .B(_4147_),
    .C(_4172_),
    .Y(_4173_));
 sg13g2_nand2_1 _4662_ (.Y(_4174_),
    .A(_4171_),
    .B(\generated._14[3] ));
 sg13g2_nor4_2 _4663_ (.A(\generated._14[1] ),
    .B(_4153_),
    .C(_0111_),
    .Y(_4175_),
    .D(_4174_));
 sg13g2_o21ai_1 _4664_ (.B1(_4152_),
    .Y(_4176_),
    .A1(_4173_),
    .A2(_4175_));
 sg13g2_nand2_1 _4665_ (.Y(_4177_),
    .A(_4170_),
    .B(_4176_));
 sg13g2_a21oi_1 _4666_ (.A1(_4147_),
    .A2(_4154_),
    .Y(_0149_),
    .B1(_4177_));
 sg13g2_inv_2 _4667_ (.Y(_4178_),
    .A(_4170_));
 sg13g2_buf_1 _4668_ (.A(_4178_),
    .X(_4179_));
 sg13g2_xnor2_1 _4669_ (.Y(_4180_),
    .A(_0111_),
    .B(_4173_));
 sg13g2_nor2_1 _4670_ (.A(_4175_),
    .B(_4151_),
    .Y(_4181_));
 sg13g2_a22oi_1 _4671_ (.Y(_4182_),
    .B1(_4180_),
    .B2(_4181_),
    .A2(_4151_),
    .A1(\generated._14[4] ));
 sg13g2_nor2_1 _4672_ (.A(net29),
    .B(_4182_),
    .Y(_0150_));
 sg13g2_nor3_1 _4673_ (.A(_4153_),
    .B(_4175_),
    .C(_4151_),
    .Y(_4183_));
 sg13g2_a21oi_1 _4674_ (.A1(_4153_),
    .A2(_4151_),
    .Y(_4184_),
    .B1(_4183_));
 sg13g2_nor2_1 _4675_ (.A(net29),
    .B(_4184_),
    .Y(_0146_));
 sg13g2_a21oi_1 _4676_ (.A1(_0149_),
    .A2(_0150_),
    .Y(_0003_),
    .B1(_0146_));
 sg13g2_inv_1 _4677_ (.Y(_4185_),
    .A(\generated._342[3] ));
 sg13g2_inv_1 _4678_ (.Y(_4186_),
    .A(\generated._353[4] ));
 sg13g2_nand2_1 _4679_ (.Y(_4187_),
    .A(\generated._353[1] ),
    .B(\generated._353[0] ));
 sg13g2_inv_1 _4680_ (.Y(_4188_),
    .A(_4187_));
 sg13g2_inv_1 _4681_ (.Y(_4189_),
    .A(\generated._353[2] ));
 sg13g2_nand2_1 _4682_ (.Y(_4190_),
    .A(_4188_),
    .B(_4189_));
 sg13g2_nor3_2 _4683_ (.A(\generated._353[3] ),
    .B(_4186_),
    .C(_4190_),
    .Y(_4191_));
 sg13g2_inv_1 _4684_ (.Y(_4192_),
    .A(_4191_));
 sg13g2_buf_1 _4685_ (.A(\generated._342[5] ),
    .X(_4193_));
 sg13g2_inv_1 _4686_ (.Y(_4194_),
    .A(_4193_));
 sg13g2_nor2_1 _4687_ (.A(\generated._342[1] ),
    .B(\generated._342[0] ),
    .Y(_4195_));
 sg13g2_buf_1 _4688_ (.A(\generated._342[2] ),
    .X(_4196_));
 sg13g2_inv_1 _4689_ (.Y(_4197_),
    .A(_4196_));
 sg13g2_nand3_1 _4690_ (.B(_4185_),
    .C(_4197_),
    .A(_4195_),
    .Y(_4198_));
 sg13g2_nor3_1 _4691_ (.A(net91),
    .B(\generated._342[4] ),
    .C(_4198_),
    .Y(_4199_));
 sg13g2_nor2_1 _4692_ (.A(_4192_),
    .B(_4199_),
    .Y(_4200_));
 sg13g2_nand2_1 _4693_ (.Y(_4201_),
    .A(\generated._342[1] ),
    .B(\generated._342[0] ));
 sg13g2_inv_1 _4694_ (.Y(_4202_),
    .A(_4201_));
 sg13g2_nand2_1 _4695_ (.Y(_4203_),
    .A(_4202_),
    .B(_4196_));
 sg13g2_xor2_1 _4696_ (.B(_4203_),
    .A(_0114_),
    .X(_4204_));
 sg13g2_nand2_1 _4697_ (.Y(_4205_),
    .A(_4200_),
    .B(_4204_));
 sg13g2_o21ai_1 _4698_ (.B1(_4205_),
    .Y(_4206_),
    .A1(_4185_),
    .A2(_4191_));
 sg13g2_nand2_2 _4699_ (.Y(_4207_),
    .A(_4206_),
    .B(_4170_));
 sg13g2_a21oi_1 _4700_ (.A1(_4191_),
    .A2(_4199_),
    .Y(_4208_),
    .B1(_4178_));
 sg13g2_inv_1 _4701_ (.Y(_4209_),
    .A(\generated._342[0] ));
 sg13g2_nor2_1 _4702_ (.A(_0112_),
    .B(_4192_),
    .Y(_4210_));
 sg13g2_a21oi_1 _4703_ (.A1(_4209_),
    .A2(_4192_),
    .Y(_4211_),
    .B1(_4210_));
 sg13g2_and2_1 _4704_ (.A(_4208_),
    .B(_4211_),
    .X(_0167_));
 sg13g2_inv_1 _4705_ (.Y(_4212_),
    .A(_0167_));
 sg13g2_nor2_1 _4706_ (.A(_4207_),
    .B(_4212_),
    .Y(_0004_));
 sg13g2_nor3_1 _4707_ (.A(_4185_),
    .B(_4203_),
    .C(_4192_),
    .Y(_4213_));
 sg13g2_xnor2_1 _4708_ (.Y(_4214_),
    .A(\generated._342[4] ),
    .B(_4213_));
 sg13g2_nor2_1 _4709_ (.A(_4178_),
    .B(_4214_),
    .Y(_0171_));
 sg13g2_inv_1 _4710_ (.Y(_4215_),
    .A(_0171_));
 sg13g2_inv_1 _4711_ (.Y(_4216_),
    .A(_4206_));
 sg13g2_nor2_1 _4712_ (.A(_4216_),
    .B(_4215_),
    .Y(_4217_));
 sg13g2_a21oi_1 _4713_ (.A1(_4207_),
    .A2(_4215_),
    .Y(_4218_),
    .B1(_4217_));
 sg13g2_nor2_1 _4714_ (.A(_4212_),
    .B(_4218_),
    .Y(_0000_));
 sg13g2_inv_1 _4715_ (.Y(_4219_),
    .A(_0115_));
 sg13g2_nor2_1 _4716_ (.A(_4191_),
    .B(_4178_),
    .Y(_4220_));
 sg13g2_nor4_1 _4717_ (.A(_4192_),
    .B(_4195_),
    .C(_4202_),
    .D(_4178_),
    .Y(_4221_));
 sg13g2_a21oi_1 _4718_ (.A1(_4219_),
    .A2(_4220_),
    .Y(_4222_),
    .B1(_4221_));
 sg13g2_nor2_1 _4719_ (.A(_4207_),
    .B(_4222_),
    .Y(_0005_));
 sg13g2_nor2_1 _4720_ (.A(_4222_),
    .B(_4218_),
    .Y(_0001_));
 sg13g2_xor2_1 _4721_ (.B(_4201_),
    .A(_0113_),
    .X(_4223_));
 sg13g2_nor2b_1 _4722_ (.A(_4178_),
    .B_N(_4223_),
    .Y(_4224_));
 sg13g2_a22oi_1 _4723_ (.Y(_4225_),
    .B1(_4196_),
    .B2(_4220_),
    .A2(_4200_),
    .A1(_4224_));
 sg13g2_buf_1 _4724_ (.A(_4225_),
    .X(_4226_));
 sg13g2_nor2_1 _4725_ (.A(_4207_),
    .B(_4226_),
    .Y(_0006_));
 sg13g2_inv_1 _4726_ (.Y(_4227_),
    .A(_4217_));
 sg13g2_nand2_1 _4727_ (.Y(_4228_),
    .A(_4215_),
    .B(_4216_));
 sg13g2_a21oi_1 _4728_ (.A1(_4227_),
    .A2(_4228_),
    .Y(_0002_),
    .B1(_4226_));
 sg13g2_inv_1 _4729_ (.Y(_4229_),
    .A(\generated._1037[0] ));
 sg13g2_buf_2 _4730_ (.A(\generated._217[3] ),
    .X(_4230_));
 sg13g2_buf_2 _4731_ (.A(\generated._610[3] ),
    .X(_4231_));
 sg13g2_buf_1 _4732_ (.A(\generated._610[1] ),
    .X(_4232_));
 sg13g2_nor2_1 _4733_ (.A(_4232_),
    .B(\generated._610[0] ),
    .Y(_4233_));
 sg13g2_inv_1 _4734_ (.Y(_4234_),
    .A(\generated._610[2] ));
 sg13g2_nand2_1 _4735_ (.Y(_4235_),
    .A(_4233_),
    .B(_4234_));
 sg13g2_buf_8 _4736_ (.A(\generated._217[0] ),
    .X(_4236_));
 sg13g2_buf_8 _4737_ (.A(\generated._610[5] ),
    .X(_4237_));
 sg13g2_nor2_1 _4738_ (.A(_4236_),
    .B(_4237_),
    .Y(_4238_));
 sg13g2_inv_1 _4739_ (.Y(_4239_),
    .A(\generated._217[2] ));
 sg13g2_inv_1 _4740_ (.Y(_4240_),
    .A(\generated._217[1] ));
 sg13g2_buf_8 _4741_ (.A(\generated._610[4] ),
    .X(_4241_));
 sg13g2_inv_1 _4742_ (.Y(_4242_),
    .A(_4241_));
 sg13g2_nand4_1 _4743_ (.B(_4239_),
    .C(_4240_),
    .A(_4238_),
    .Y(_4243_),
    .D(_4242_));
 sg13g2_nor4_1 _4744_ (.A(_4230_),
    .B(_4231_),
    .C(_4235_),
    .D(_4243_),
    .Y(_4244_));
 sg13g2_nand2_2 _4745_ (.Y(_4245_),
    .A(_4178_),
    .B(_4244_));
 sg13g2_nor2_1 _4746_ (.A(\generated._75[0] ),
    .B(_4245_),
    .Y(_4246_));
 sg13g2_a21oi_1 _4747_ (.A1(_4229_),
    .A2(_4245_),
    .Y(_0234_),
    .B1(_4246_));
 sg13g2_inv_1 _4748_ (.Y(_4247_),
    .A(\generated._402[1] ));
 sg13g2_nor3_2 _4749_ (.A(_4247_),
    .B(_4229_),
    .C(_4245_),
    .Y(_4248_));
 sg13g2_o21ai_1 _4750_ (.B1(_4247_),
    .Y(_4249_),
    .A1(_4229_),
    .A2(_4245_));
 sg13g2_nor2b_1 _4751_ (.A(_4248_),
    .B_N(_4249_),
    .Y(_0235_));
 sg13g2_inv_1 _4752_ (.Y(_4250_),
    .A(\generated._402[2] ));
 sg13g2_xnor2_1 _4753_ (.Y(_0236_),
    .A(_4250_),
    .B(_4248_));
 sg13g2_inv_1 _4754_ (.Y(_4251_),
    .A(\generated._402[3] ));
 sg13g2_nor4_2 _4755_ (.A(_4247_),
    .B(_4250_),
    .C(_4229_),
    .Y(_4252_),
    .D(_4245_));
 sg13g2_xnor2_1 _4756_ (.Y(_0237_),
    .A(_4251_),
    .B(_4252_));
 sg13g2_buf_1 _4757_ (.A(\generated._402[4] ),
    .X(_4253_));
 sg13g2_nand2_1 _4758_ (.Y(_4254_),
    .A(_4252_),
    .B(\generated._402[3] ));
 sg13g2_xnor2_1 _4759_ (.Y(_0238_),
    .A(_4253_),
    .B(_4254_));
 sg13g2_nand4_1 _4760_ (.B(\generated._402[2] ),
    .C(\generated._402[3] ),
    .A(_4248_),
    .Y(_4255_),
    .D(_4253_));
 sg13g2_xnor2_1 _4761_ (.Y(_0239_),
    .A(\generated._402[5] ),
    .B(_4255_));
 sg13g2_inv_1 _4762_ (.Y(_4256_),
    .A(\generated._402[6] ));
 sg13g2_inv_1 _4763_ (.Y(_4257_),
    .A(\generated._402[5] ));
 sg13g2_nor2_1 _4764_ (.A(_4257_),
    .B(_4255_),
    .Y(_4258_));
 sg13g2_xnor2_1 _4765_ (.Y(_0240_),
    .A(_4256_),
    .B(_4258_));
 sg13g2_nand2_1 _4766_ (.Y(_4259_),
    .A(_4258_),
    .B(\generated._402[6] ));
 sg13g2_xnor2_1 _4767_ (.Y(_0241_),
    .A(\generated._402[7] ),
    .B(_4259_));
 sg13g2_inv_2 _4768_ (.Y(_4260_),
    .A(_4162_));
 sg13g2_nand2_1 _4769_ (.Y(_4261_),
    .A(\generated._568[1] ),
    .B(\generated._568[0] ));
 sg13g2_nor2_1 _4770_ (.A(_4167_),
    .B(_4261_),
    .Y(_4262_));
 sg13g2_inv_1 _4771_ (.Y(_4263_),
    .A(_4262_));
 sg13g2_nor2_1 _4772_ (.A(_4260_),
    .B(_4263_),
    .Y(_4264_));
 sg13g2_inv_8 _4773_ (.Y(_4265_),
    .A(_4156_));
 sg13g2_nor2_1 _4774_ (.A(_4159_),
    .B(_4161_),
    .Y(_4266_));
 sg13g2_inv_1 _4775_ (.Y(_4267_),
    .A(_4266_));
 sg13g2_nor2_1 _4776_ (.A(_4265_),
    .B(_4267_),
    .Y(_4268_));
 sg13g2_nor2_1 _4777_ (.A(net95),
    .B(_4155_),
    .Y(_4269_));
 sg13g2_inv_2 _4778_ (.Y(_4270_),
    .A(_4157_));
 sg13g2_nand2_1 _4779_ (.Y(_4271_),
    .A(_4269_),
    .B(_4270_));
 sg13g2_inv_1 _4780_ (.Y(_4272_),
    .A(_4271_));
 sg13g2_nand3_1 _4781_ (.B(_4268_),
    .C(_4272_),
    .A(_4264_),
    .Y(_4273_));
 sg13g2_buf_2 _4782_ (.A(_4273_),
    .X(_4274_));
 sg13g2_nand2_1 _4783_ (.Y(_4275_),
    .A(_4231_),
    .B(\generated._610[2] ));
 sg13g2_nand2_1 _4784_ (.Y(_4276_),
    .A(_4233_),
    .B(_4230_));
 sg13g2_nor3_1 _4785_ (.A(_4275_),
    .B(_4276_),
    .C(_4243_),
    .Y(_4277_));
 sg13g2_nor2_1 _4786_ (.A(_4274_),
    .B(_4277_),
    .Y(_4278_));
 sg13g2_inv_1 _4787_ (.Y(_4279_),
    .A(_4278_));
 sg13g2_inv_1 _4788_ (.Y(_4280_),
    .A(\generated._610[0] ));
 sg13g2_nor2_1 _4789_ (.A(_4280_),
    .B(_4274_),
    .Y(_4281_));
 sg13g2_a21oi_1 _4790_ (.A1(_4279_),
    .A2(_4280_),
    .Y(_0224_),
    .B1(_4281_));
 sg13g2_inv_1 _4791_ (.Y(_4282_),
    .A(_4232_));
 sg13g2_xnor2_1 _4792_ (.Y(_0225_),
    .A(_4282_),
    .B(_4281_));
 sg13g2_nand2_1 _4793_ (.Y(_4283_),
    .A(_4281_),
    .B(_4232_));
 sg13g2_inv_1 _4794_ (.Y(_4284_),
    .A(_4274_));
 sg13g2_nand2_1 _4795_ (.Y(_4285_),
    .A(_4232_),
    .B(\generated._610[0] ));
 sg13g2_nor2_1 _4796_ (.A(_4234_),
    .B(_4285_),
    .Y(_4286_));
 sg13g2_inv_1 _4797_ (.Y(_4287_),
    .A(_4286_));
 sg13g2_nand2b_1 _4798_ (.Y(_4288_),
    .B(_4287_),
    .A_N(_4277_));
 sg13g2_a22oi_1 _4799_ (.Y(_0226_),
    .B1(_4284_),
    .B2(_4288_),
    .A2(_4234_),
    .A1(_4283_));
 sg13g2_inv_1 _4800_ (.Y(_4289_),
    .A(_0116_));
 sg13g2_xnor2_1 _4801_ (.Y(_4290_),
    .A(_4289_),
    .B(_4286_));
 sg13g2_nand2_1 _4802_ (.Y(_4291_),
    .A(_4274_),
    .B(_4231_));
 sg13g2_o21ai_1 _4803_ (.B1(_4291_),
    .Y(_0227_),
    .A1(_4290_),
    .A2(_4279_));
 sg13g2_nor3_1 _4804_ (.A(_4275_),
    .B(_4285_),
    .C(_4274_),
    .Y(_4292_));
 sg13g2_xnor2_1 _4805_ (.Y(_0228_),
    .A(_4242_),
    .B(_4292_));
 sg13g2_buf_1 _4806_ (.A(_0123_),
    .X(_4293_));
 sg13g2_inv_1 _4807_ (.Y(_4294_),
    .A(net94));
 sg13g2_buf_1 _4808_ (.A(_4294_),
    .X(_4295_));
 sg13g2_nand2_2 _4809_ (.Y(_4296_),
    .A(_4241_),
    .B(_4231_));
 sg13g2_nor2_2 _4810_ (.A(_4296_),
    .B(_4287_),
    .Y(_4297_));
 sg13g2_o21ai_1 _4811_ (.B1(_4278_),
    .Y(_4298_),
    .A1(net79),
    .A2(_4297_));
 sg13g2_a21oi_1 _4812_ (.A1(net79),
    .A2(_4297_),
    .Y(_4299_),
    .B1(_4298_));
 sg13g2_a21o_1 _4813_ (.A2(_4274_),
    .A1(_4237_),
    .B1(_4299_),
    .X(_0229_));
 sg13g2_nand2_1 _4814_ (.Y(_4300_),
    .A(_4297_),
    .B(_4237_));
 sg13g2_o21ai_1 _4815_ (.B1(_4278_),
    .Y(_4301_),
    .A1(_0118_),
    .A2(_4300_));
 sg13g2_a21oi_1 _4816_ (.A1(_0118_),
    .A2(_4300_),
    .Y(_4302_),
    .B1(_4301_));
 sg13g2_a21o_1 _4817_ (.A2(_4274_),
    .A1(_4236_),
    .B1(_4302_),
    .X(_0230_));
 sg13g2_nand2_1 _4818_ (.Y(_4303_),
    .A(_4236_),
    .B(_4237_));
 sg13g2_nor2_1 _4819_ (.A(_4296_),
    .B(_4303_),
    .Y(_4304_));
 sg13g2_xnor2_1 _4820_ (.Y(_4305_),
    .A(_0124_),
    .B(_4304_));
 sg13g2_a21oi_1 _4821_ (.A1(_0124_),
    .A2(_4287_),
    .Y(_4306_),
    .B1(_4279_));
 sg13g2_o21ai_1 _4822_ (.B1(_4306_),
    .Y(_4307_),
    .A1(_4287_),
    .A2(_4305_));
 sg13g2_o21ai_1 _4823_ (.B1(_4307_),
    .Y(_0231_),
    .A1(_4240_),
    .A2(_4284_));
 sg13g2_nand3_1 _4824_ (.B(_4286_),
    .C(\generated._217[1] ),
    .A(_4304_),
    .Y(_4308_));
 sg13g2_xnor2_1 _4825_ (.Y(_4309_),
    .A(_0125_),
    .B(_4308_));
 sg13g2_nand2_1 _4826_ (.Y(_4310_),
    .A(_4274_),
    .B(\generated._217[2] ));
 sg13g2_o21ai_1 _4827_ (.B1(_4310_),
    .Y(_0232_),
    .A1(_4309_),
    .A2(_4279_));
 sg13g2_inv_1 _4828_ (.Y(_4311_),
    .A(_4230_));
 sg13g2_nand2_1 _4829_ (.Y(_4312_),
    .A(\generated._217[1] ),
    .B(_4236_));
 sg13g2_nor2_1 _4830_ (.A(_4239_),
    .B(_4312_),
    .Y(_4313_));
 sg13g2_nand2_1 _4831_ (.Y(_4314_),
    .A(_4313_),
    .B(_4237_));
 sg13g2_inv_1 _4832_ (.Y(_4315_),
    .A(_4314_));
 sg13g2_inv_1 _4833_ (.Y(_4316_),
    .A(_0126_));
 sg13g2_nand3_1 _4834_ (.B(_4315_),
    .C(_4316_),
    .A(_4297_),
    .Y(_4317_));
 sg13g2_a21o_1 _4835_ (.A2(_4315_),
    .A1(_4297_),
    .B1(_4316_),
    .X(_4318_));
 sg13g2_nand3_1 _4836_ (.B(_4317_),
    .C(_4318_),
    .A(_4278_),
    .Y(_4319_));
 sg13g2_o21ai_1 _4837_ (.B1(_4319_),
    .Y(_0233_),
    .A1(_4311_),
    .A2(_4284_));
 sg13g2_nor2_1 _4838_ (.A(\generated._1074[1] ),
    .B(\generated._1074[0] ),
    .Y(_4320_));
 sg13g2_inv_1 _4839_ (.Y(_4321_),
    .A(\generated._1074[2] ));
 sg13g2_inv_1 _4840_ (.Y(_4322_),
    .A(\generated._1074[3] ));
 sg13g2_nand3_1 _4841_ (.B(_4321_),
    .C(_4322_),
    .A(_4320_),
    .Y(_4323_));
 sg13g2_buf_2 _4842_ (.A(_4323_),
    .X(_4324_));
 sg13g2_inv_1 _4843_ (.Y(_4325_),
    .A(_4324_));
 sg13g2_buf_1 _4844_ (.A(_4325_),
    .X(_4326_));
 sg13g2_buf_1 _4845_ (.A(net48),
    .X(_4327_));
 sg13g2_buf_1 _4846_ (.A(\generated._966 ),
    .X(_4328_));
 sg13g2_nor2_1 _4847_ (.A(_4328_),
    .B(\generated._965 ),
    .Y(_4329_));
 sg13g2_buf_2 _4848_ (.A(_4329_),
    .X(_4330_));
 sg13g2_buf_1 _4849_ (.A(\generated._965 ),
    .X(_4331_));
 sg13g2_inv_1 _4850_ (.Y(_4332_),
    .A(_4328_));
 sg13g2_nor2_2 _4851_ (.A(_4331_),
    .B(_4332_),
    .Y(_4333_));
 sg13g2_a22oi_1 _4852_ (.Y(_4334_),
    .B1(_0022_),
    .B2(_4333_),
    .A2(_0096_),
    .A1(_4330_));
 sg13g2_buf_1 _4853_ (.A(_4328_),
    .X(_4335_));
 sg13g2_inv_1 _4854_ (.Y(_4336_),
    .A(_0016_));
 sg13g2_nor2_1 _4855_ (.A(net90),
    .B(_0021_),
    .Y(_4337_));
 sg13g2_a21oi_1 _4856_ (.A1(net90),
    .A2(_4336_),
    .Y(_4338_),
    .B1(_4337_));
 sg13g2_nand2_1 _4857_ (.Y(_4339_),
    .A(_4338_),
    .B(net93));
 sg13g2_and2_1 _4858_ (.A(_4334_),
    .B(_4339_),
    .X(_4340_));
 sg13g2_buf_1 _4859_ (.A(_4340_),
    .X(_4341_));
 sg13g2_xor2_1 _4860_ (.B(_4341_),
    .A(_0097_),
    .X(_4342_));
 sg13g2_nor2_1 _4861_ (.A(net36),
    .B(_4342_),
    .Y(_0130_));
 sg13g2_nand2_1 _4862_ (.Y(_4343_),
    .A(_4341_),
    .B(\generated._1020[0] ));
 sg13g2_nand2_1 _4863_ (.Y(_4344_),
    .A(net90),
    .B(_0023_));
 sg13g2_o21ai_1 _4864_ (.B1(_4344_),
    .Y(_4345_),
    .A1(net90),
    .A2(_4336_));
 sg13g2_and2_1 _4865_ (.A(_4330_),
    .B(_0022_),
    .X(_4346_));
 sg13g2_a221oi_1 _4866_ (.B2(net93),
    .C1(_4346_),
    .B1(_4345_),
    .A1(_0021_),
    .Y(_4347_),
    .A2(_4333_));
 sg13g2_nor4_1 _4867_ (.A(\generated._1070[3] ),
    .B(\generated._1070[2] ),
    .C(\generated._1070[1] ),
    .D(\generated._1070[0] ),
    .Y(_4348_));
 sg13g2_nor4_1 _4868_ (.A(\generated._1070[7] ),
    .B(\generated._1070[6] ),
    .C(\generated._1070[5] ),
    .D(\generated._1070[4] ),
    .Y(_4349_));
 sg13g2_nor2_1 _4869_ (.A(\generated._1070[8] ),
    .B(\generated._1070[9] ),
    .Y(_4350_));
 sg13g2_nand3_1 _4870_ (.B(_4349_),
    .C(_4350_),
    .A(_4348_),
    .Y(_4351_));
 sg13g2_inv_1 _4871_ (.Y(_4352_),
    .A(_0020_));
 sg13g2_nand2_1 _4872_ (.Y(_4353_),
    .A(_4351_),
    .B(_4352_));
 sg13g2_buf_1 _4873_ (.A(_4353_),
    .X(_4354_));
 sg13g2_inv_1 _4874_ (.Y(_4355_),
    .A(_4354_));
 sg13g2_nand2_1 _4875_ (.Y(_4356_),
    .A(net47),
    .B(_4341_));
 sg13g2_xor2_1 _4876_ (.B(_4356_),
    .A(_4347_),
    .X(_4357_));
 sg13g2_xor2_1 _4877_ (.B(_4357_),
    .A(\generated._1020[1] ),
    .X(_4358_));
 sg13g2_nor2_1 _4878_ (.A(_4343_),
    .B(_4358_),
    .Y(_4359_));
 sg13g2_a21oi_1 _4879_ (.A1(_4358_),
    .A2(_4343_),
    .Y(_4360_),
    .B1(net48));
 sg13g2_nor2b_1 _4880_ (.A(_4359_),
    .B_N(_4360_),
    .Y(_0131_));
 sg13g2_inv_1 _4881_ (.Y(_4361_),
    .A(net93));
 sg13g2_buf_1 _4882_ (.A(_4361_),
    .X(_4362_));
 sg13g2_buf_1 _4883_ (.A(_4335_),
    .X(_4363_));
 sg13g2_inv_1 _4884_ (.Y(_4364_),
    .A(_0026_));
 sg13g2_nand2_1 _4885_ (.Y(_4365_),
    .A(_4364_),
    .B(net90));
 sg13g2_o21ai_1 _4886_ (.B1(_4365_),
    .Y(_4366_),
    .A1(net77),
    .A2(_0023_));
 sg13g2_nor2_1 _4887_ (.A(_4361_),
    .B(_4366_),
    .Y(_4367_));
 sg13g2_a21oi_1 _4888_ (.A1(net78),
    .A2(_4338_),
    .Y(_4368_),
    .B1(_4367_));
 sg13g2_buf_1 _4889_ (.A(_4354_),
    .X(_4369_));
 sg13g2_nor2_1 _4890_ (.A(_4341_),
    .B(_4347_),
    .Y(_4370_));
 sg13g2_nor2_1 _4891_ (.A(net46),
    .B(_4370_),
    .Y(_4371_));
 sg13g2_xor2_1 _4892_ (.B(_4371_),
    .A(_4368_),
    .X(_4372_));
 sg13g2_xor2_1 _4893_ (.B(_4372_),
    .A(\generated._1020[2] ),
    .X(_4373_));
 sg13g2_nor2_1 _4894_ (.A(_0098_),
    .B(_4357_),
    .Y(_4374_));
 sg13g2_nor2_1 _4895_ (.A(_4374_),
    .B(_4359_),
    .Y(_4375_));
 sg13g2_inv_1 _4896_ (.Y(_4376_),
    .A(_4375_));
 sg13g2_buf_1 _4897_ (.A(_4324_),
    .X(_4377_));
 sg13g2_o21ai_1 _4898_ (.B1(net65),
    .Y(_4378_),
    .A1(_4373_),
    .A2(_4376_));
 sg13g2_nand2_1 _4899_ (.Y(_4379_),
    .A(_4376_),
    .B(_4373_));
 sg13g2_nor2b_1 _4900_ (.A(_4378_),
    .B_N(_4379_),
    .Y(_0132_));
 sg13g2_inv_1 _4901_ (.Y(_4380_),
    .A(_0096_));
 sg13g2_a22oi_1 _4902_ (.Y(_4381_),
    .B1(_0098_),
    .B2(_4333_),
    .A2(_0097_),
    .A1(_4330_));
 sg13g2_inv_1 _4903_ (.Y(_4382_),
    .A(_0099_));
 sg13g2_nand2_1 _4904_ (.Y(_4383_),
    .A(_4328_),
    .B(_0100_));
 sg13g2_o21ai_1 _4905_ (.B1(_4383_),
    .Y(_4384_),
    .A1(_4328_),
    .A2(_4382_));
 sg13g2_nand2_1 _4906_ (.Y(_4385_),
    .A(_4384_),
    .B(net93));
 sg13g2_and2_1 _4907_ (.A(_4381_),
    .B(_4385_),
    .X(_4386_));
 sg13g2_inv_1 _4908_ (.Y(_4387_),
    .A(_4386_));
 sg13g2_nor2_1 _4909_ (.A(_4380_),
    .B(_4387_),
    .Y(_4388_));
 sg13g2_inv_1 _4910_ (.Y(_4389_),
    .A(_4388_));
 sg13g2_nand2_1 _4911_ (.Y(_4390_),
    .A(_4387_),
    .B(_4380_));
 sg13g2_a21oi_1 _4912_ (.A1(_4389_),
    .A2(_4390_),
    .Y(_0133_),
    .B1(net36));
 sg13g2_nand2_1 _4913_ (.Y(_4391_),
    .A(net90),
    .B(_0017_));
 sg13g2_inv_1 _4914_ (.Y(_4392_),
    .A(_4391_));
 sg13g2_a21oi_1 _4915_ (.A1(_4332_),
    .A2(_0100_),
    .Y(_4393_),
    .B1(_4392_));
 sg13g2_nor2_1 _4916_ (.A(_4361_),
    .B(_4393_),
    .Y(_4394_));
 sg13g2_a221oi_1 _4917_ (.B2(_4333_),
    .C1(_4394_),
    .B1(_0099_),
    .A1(_0098_),
    .Y(_4395_),
    .A2(_4330_));
 sg13g2_nor2_1 _4918_ (.A(_4387_),
    .B(_4354_),
    .Y(_4396_));
 sg13g2_xnor2_1 _4919_ (.Y(_4397_),
    .A(_4395_),
    .B(_4396_));
 sg13g2_xor2_1 _4920_ (.B(_4397_),
    .A(_0022_),
    .X(_4398_));
 sg13g2_nor2_1 _4921_ (.A(_4388_),
    .B(_4398_),
    .Y(_4399_));
 sg13g2_inv_1 _4922_ (.Y(_4400_),
    .A(_4399_));
 sg13g2_nand2_1 _4923_ (.Y(_4401_),
    .A(_4400_),
    .B(net65));
 sg13g2_a21oi_1 _4924_ (.A1(_4388_),
    .A2(_4398_),
    .Y(_0134_),
    .B1(_4401_));
 sg13g2_inv_1 _4925_ (.Y(_4402_),
    .A(_0017_));
 sg13g2_nor2_1 _4926_ (.A(net90),
    .B(_4402_),
    .Y(_4403_));
 sg13g2_a21oi_1 _4927_ (.A1(_4335_),
    .A2(_0018_),
    .Y(_4404_),
    .B1(_4403_));
 sg13g2_nor2_1 _4928_ (.A(_4361_),
    .B(_4404_),
    .Y(_4405_));
 sg13g2_a21oi_1 _4929_ (.A1(_4361_),
    .A2(_4384_),
    .Y(_4406_),
    .B1(_4405_));
 sg13g2_nor2_1 _4930_ (.A(_4386_),
    .B(_4395_),
    .Y(_4407_));
 sg13g2_nor2_1 _4931_ (.A(_4354_),
    .B(_4407_),
    .Y(_4408_));
 sg13g2_xnor2_1 _4932_ (.Y(_4409_),
    .A(_4406_),
    .B(_4408_));
 sg13g2_xnor2_1 _4933_ (.Y(_4410_),
    .A(_0021_),
    .B(_4409_));
 sg13g2_a21o_1 _4934_ (.A2(_4397_),
    .A1(\generated._1070[1] ),
    .B1(_4399_),
    .X(_4411_));
 sg13g2_o21ai_1 _4935_ (.B1(net65),
    .Y(_4412_),
    .A1(_4410_),
    .A2(_4411_));
 sg13g2_nand2_1 _4936_ (.Y(_4413_),
    .A(_4411_),
    .B(_4410_));
 sg13g2_nor2b_1 _4937_ (.A(_4412_),
    .B_N(_4413_),
    .Y(_0135_));
 sg13g2_inv_1 _4938_ (.Y(_4414_),
    .A(_0088_));
 sg13g2_nand2_1 _4939_ (.Y(_4415_),
    .A(net77),
    .B(net93));
 sg13g2_xnor2_1 _4940_ (.Y(_4416_),
    .A(_4414_),
    .B(_4415_));
 sg13g2_nor2_1 _4941_ (.A(_4416_),
    .B(net36),
    .Y(_0136_));
 sg13g2_buf_1 _4942_ (.A(\generated._1080[1] ),
    .X(_4417_));
 sg13g2_xnor2_1 _4943_ (.Y(_4418_),
    .A(_4330_),
    .B(_4354_));
 sg13g2_inv_1 _4944_ (.Y(_4419_),
    .A(_4418_));
 sg13g2_nand2_2 _4945_ (.Y(_4420_),
    .A(_4419_),
    .B(_4415_));
 sg13g2_xnor2_1 _4946_ (.Y(_4421_),
    .A(_4417_),
    .B(_4420_));
 sg13g2_nand2_1 _4947_ (.Y(_4422_),
    .A(_4415_),
    .B(\generated._1080[0] ));
 sg13g2_nor2b_1 _4948_ (.A(_4421_),
    .B_N(_4422_),
    .Y(_4423_));
 sg13g2_nor2b_1 _4949_ (.A(_4422_),
    .B_N(_4421_),
    .Y(_4424_));
 sg13g2_nor3_1 _4950_ (.A(net36),
    .B(_4423_),
    .C(_4424_),
    .Y(_0137_));
 sg13g2_buf_1 _4951_ (.A(\generated._1080[2] ),
    .X(_4425_));
 sg13g2_buf_1 _4952_ (.A(_4363_),
    .X(_4426_));
 sg13g2_nor2_1 _4953_ (.A(_4333_),
    .B(net46),
    .Y(_4427_));
 sg13g2_a21oi_1 _4954_ (.A1(net64),
    .A2(net46),
    .Y(_4428_),
    .B1(_4427_));
 sg13g2_nor2_1 _4955_ (.A(_4425_),
    .B(_4428_),
    .Y(_4429_));
 sg13g2_inv_1 _4956_ (.Y(_4430_),
    .A(_4425_));
 sg13g2_nor2b_1 _4957_ (.A(_4430_),
    .B_N(_4428_),
    .Y(_4431_));
 sg13g2_nor2_1 _4958_ (.A(_4429_),
    .B(_4431_),
    .Y(_4432_));
 sg13g2_inv_1 _4959_ (.Y(_4433_),
    .A(_4417_));
 sg13g2_nor2_1 _4960_ (.A(_4433_),
    .B(_4420_),
    .Y(_4434_));
 sg13g2_nor2_1 _4961_ (.A(_4434_),
    .B(_4424_),
    .Y(_4435_));
 sg13g2_xor2_1 _4962_ (.B(_4435_),
    .A(_4432_),
    .X(_4436_));
 sg13g2_nor2_1 _4963_ (.A(net36),
    .B(_4436_),
    .Y(_0138_));
 sg13g2_buf_1 _4964_ (.A(\generated._1080[3] ),
    .X(_4437_));
 sg13g2_xnor2_1 _4965_ (.Y(_4438_),
    .A(_4437_),
    .B(_4420_));
 sg13g2_inv_1 _4966_ (.Y(_4439_),
    .A(_4438_));
 sg13g2_nor2_1 _4967_ (.A(_4429_),
    .B(_4435_),
    .Y(_4440_));
 sg13g2_nor2_1 _4968_ (.A(_4431_),
    .B(_4440_),
    .Y(_4441_));
 sg13g2_o21ai_1 _4969_ (.B1(net65),
    .Y(_4442_),
    .A1(_4439_),
    .A2(_4441_));
 sg13g2_a21oi_1 _4970_ (.A1(_4439_),
    .A2(_4441_),
    .Y(_0139_),
    .B1(_4442_));
 sg13g2_buf_1 _4971_ (.A(\generated._1080[4] ),
    .X(_4443_));
 sg13g2_buf_1 _4972_ (.A(net46),
    .X(_4444_));
 sg13g2_buf_1 _4973_ (.A(_4331_),
    .X(_4445_));
 sg13g2_xnor2_1 _4974_ (.Y(_4446_),
    .A(net64),
    .B(net89));
 sg13g2_nor2_1 _4975_ (.A(_4446_),
    .B(net35),
    .Y(_4447_));
 sg13g2_a21oi_1 _4976_ (.A1(_4330_),
    .A2(net35),
    .Y(_4448_),
    .B1(_4447_));
 sg13g2_nor2_1 _4977_ (.A(_4443_),
    .B(_4448_),
    .Y(_4449_));
 sg13g2_nand2_1 _4978_ (.Y(_4450_),
    .A(_4448_),
    .B(_4443_));
 sg13g2_nor2b_1 _4979_ (.A(_4449_),
    .B_N(_4450_),
    .Y(_4451_));
 sg13g2_inv_1 _4980_ (.Y(_4452_),
    .A(_4441_));
 sg13g2_nor2b_1 _4981_ (.A(_4420_),
    .B_N(_4437_),
    .Y(_4453_));
 sg13g2_a21oi_1 _4982_ (.A1(_4452_),
    .A2(_4438_),
    .Y(_4454_),
    .B1(_4453_));
 sg13g2_xor2_1 _4983_ (.B(_4454_),
    .A(_4451_),
    .X(_4455_));
 sg13g2_nor2_1 _4984_ (.A(_4327_),
    .B(_4455_),
    .Y(_0140_));
 sg13g2_buf_1 _4985_ (.A(\generated._1080[5] ),
    .X(_4456_));
 sg13g2_inv_1 _4986_ (.Y(_4457_),
    .A(_4456_));
 sg13g2_xnor2_1 _4987_ (.Y(_4458_),
    .A(net89),
    .B(net35));
 sg13g2_nor2_1 _4988_ (.A(_4457_),
    .B(_4458_),
    .Y(_4459_));
 sg13g2_inv_1 _4989_ (.Y(_4460_),
    .A(_4459_));
 sg13g2_nand2_1 _4990_ (.Y(_4461_),
    .A(_4458_),
    .B(_4457_));
 sg13g2_o21ai_1 _4991_ (.B1(_4450_),
    .Y(_4462_),
    .A1(_4449_),
    .A2(_4454_));
 sg13g2_a21oi_1 _4992_ (.A1(_4460_),
    .A2(_4461_),
    .Y(_4463_),
    .B1(_4462_));
 sg13g2_nand2_1 _4993_ (.Y(_4464_),
    .A(_4462_),
    .B(_4461_));
 sg13g2_nor2_1 _4994_ (.A(_4459_),
    .B(_4464_),
    .Y(_4465_));
 sg13g2_nor3_1 _4995_ (.A(net36),
    .B(_4463_),
    .C(_4465_),
    .Y(_0141_));
 sg13g2_buf_1 _4996_ (.A(\generated._1080[6] ),
    .X(_4466_));
 sg13g2_nor2_1 _4997_ (.A(_4466_),
    .B(_4418_),
    .Y(_4467_));
 sg13g2_nor2b_1 _4998_ (.A(_4419_),
    .B_N(_4466_),
    .Y(_4468_));
 sg13g2_nor2_1 _4999_ (.A(_4467_),
    .B(_4468_),
    .Y(_4469_));
 sg13g2_nand2_1 _5000_ (.Y(_4470_),
    .A(_4464_),
    .B(_4460_));
 sg13g2_o21ai_1 _5001_ (.B1(_4377_),
    .Y(_4471_),
    .A1(_4469_),
    .A2(_4470_));
 sg13g2_nand2_1 _5002_ (.Y(_4472_),
    .A(_4470_),
    .B(_4469_));
 sg13g2_nor2b_1 _5003_ (.A(_4471_),
    .B_N(_4472_),
    .Y(_0142_));
 sg13g2_buf_1 _5004_ (.A(\generated._1080[7] ),
    .X(_4473_));
 sg13g2_nor2b_1 _5005_ (.A(net35),
    .B_N(_4473_),
    .Y(_4474_));
 sg13g2_nor2_1 _5006_ (.A(_4473_),
    .B(net47),
    .Y(_4475_));
 sg13g2_nor2_1 _5007_ (.A(_4474_),
    .B(_4475_),
    .Y(_4476_));
 sg13g2_inv_1 _5008_ (.Y(_4477_),
    .A(_4467_));
 sg13g2_a21oi_1 _5009_ (.A1(_4470_),
    .A2(_4477_),
    .Y(_4478_),
    .B1(_4468_));
 sg13g2_inv_1 _5010_ (.Y(_4479_),
    .A(_4478_));
 sg13g2_nor2_1 _5011_ (.A(_4476_),
    .B(_4479_),
    .Y(_4480_));
 sg13g2_nand2_1 _5012_ (.Y(_4481_),
    .A(_4479_),
    .B(_4476_));
 sg13g2_inv_1 _5013_ (.Y(_4482_),
    .A(_4481_));
 sg13g2_nor3_1 _5014_ (.A(net48),
    .B(_4480_),
    .C(_4482_),
    .Y(_0143_));
 sg13g2_buf_1 _5015_ (.A(\generated._1080[8] ),
    .X(_4483_));
 sg13g2_xnor2_1 _5016_ (.Y(_4484_),
    .A(_4483_),
    .B(net35));
 sg13g2_nor2_1 _5017_ (.A(_4474_),
    .B(_4468_),
    .Y(_4485_));
 sg13g2_a21oi_1 _5018_ (.A1(_4472_),
    .A2(_4485_),
    .Y(_4486_),
    .B1(_4475_));
 sg13g2_o21ai_1 _5019_ (.B1(net65),
    .Y(_4487_),
    .A1(_4484_),
    .A2(_4486_));
 sg13g2_a21oi_1 _5020_ (.A1(_4484_),
    .A2(_4486_),
    .Y(_0144_),
    .B1(_4487_));
 sg13g2_buf_1 _5021_ (.A(\generated._1080[9] ),
    .X(_4488_));
 sg13g2_buf_1 _5022_ (.A(_4488_),
    .X(_4489_));
 sg13g2_buf_1 _5023_ (.A(_4489_),
    .X(_4490_));
 sg13g2_buf_1 _5024_ (.A(net76),
    .X(_4491_));
 sg13g2_buf_1 _5025_ (.A(net63),
    .X(_4492_));
 sg13g2_xnor2_1 _5026_ (.Y(_4493_),
    .A(net45),
    .B(net35));
 sg13g2_nor2b_1 _5027_ (.A(net35),
    .B_N(_4483_),
    .Y(_4494_));
 sg13g2_a221oi_1 _5028_ (.B2(_4484_),
    .C1(_4494_),
    .B1(_4482_),
    .A1(_4473_),
    .Y(_4495_),
    .A2(_4355_));
 sg13g2_xor2_1 _5029_ (.B(_4495_),
    .A(_4493_),
    .X(_4496_));
 sg13g2_nor2_1 _5030_ (.A(net36),
    .B(_4496_),
    .Y(_0145_));
 sg13g2_a21oi_1 _5031_ (.A1(_4152_),
    .A2(_4153_),
    .Y(_4497_),
    .B1(\generated._14[1] ));
 sg13g2_nor2_1 _5032_ (.A(_4172_),
    .B(_4151_),
    .Y(_4498_));
 sg13g2_nor3_1 _5033_ (.A(_4497_),
    .B(_4498_),
    .C(net29),
    .Y(_0147_));
 sg13g2_o21ai_1 _5034_ (.B1(_4154_),
    .Y(_4499_),
    .A1(\generated._14[2] ),
    .A2(_4498_));
 sg13g2_nor2_1 _5035_ (.A(net29),
    .B(_4499_),
    .Y(_0148_));
 sg13g2_nand2_2 _5036_ (.Y(_4500_),
    .A(_4170_),
    .B(_4151_));
 sg13g2_nor2b_1 _5037_ (.A(_4500_),
    .B_N(\generated._297[0] ),
    .Y(_0151_));
 sg13g2_nand2_1 _5038_ (.Y(_4501_),
    .A(\generated._19[1] ),
    .B(\generated._19[0] ));
 sg13g2_inv_1 _5039_ (.Y(_4502_),
    .A(_4501_));
 sg13g2_nor2_1 _5040_ (.A(\generated._19[1] ),
    .B(\generated._19[0] ),
    .Y(_4503_));
 sg13g2_nor3_1 _5041_ (.A(_4502_),
    .B(_4503_),
    .C(_4500_),
    .Y(_0152_));
 sg13g2_nor2_1 _5042_ (.A(_4149_),
    .B(_4501_),
    .Y(_4504_));
 sg13g2_nor2_1 _5043_ (.A(\generated._19[2] ),
    .B(_4502_),
    .Y(_4505_));
 sg13g2_nor3_1 _5044_ (.A(_4504_),
    .B(_4505_),
    .C(_4500_),
    .Y(_0153_));
 sg13g2_and2_1 _5045_ (.A(_4504_),
    .B(\generated._19[3] ),
    .X(_4506_));
 sg13g2_nor2_1 _5046_ (.A(\generated._19[3] ),
    .B(_4504_),
    .Y(_4507_));
 sg13g2_nor3_1 _5047_ (.A(_4506_),
    .B(_4507_),
    .C(_4500_),
    .Y(_0154_));
 sg13g2_xnor2_1 _5048_ (.Y(_4508_),
    .A(\generated._19[4] ),
    .B(_4506_));
 sg13g2_nor2_1 _5049_ (.A(_4508_),
    .B(_4500_),
    .Y(_0155_));
 sg13g2_buf_1 _5050_ (.A(\generated._26[0] ),
    .X(_4509_));
 sg13g2_inv_1 _5051_ (.Y(_4510_),
    .A(\generated._31[6] ));
 sg13g2_inv_1 _5052_ (.Y(_4511_),
    .A(\generated._31[3] ));
 sg13g2_inv_1 _5053_ (.Y(_4512_),
    .A(\generated._31[2] ));
 sg13g2_nand2_1 _5054_ (.Y(_4513_),
    .A(\generated._31[1] ),
    .B(\generated._31[0] ));
 sg13g2_nor2_1 _5055_ (.A(_4512_),
    .B(_4513_),
    .Y(_4514_));
 sg13g2_inv_1 _5056_ (.Y(_4515_),
    .A(_4514_));
 sg13g2_nor2_1 _5057_ (.A(_4511_),
    .B(_4515_),
    .Y(_4516_));
 sg13g2_inv_1 _5058_ (.Y(_4517_),
    .A(_4516_));
 sg13g2_nor4_2 _5059_ (.A(\generated._31[5] ),
    .B(\generated._31[4] ),
    .C(_4510_),
    .Y(_4518_),
    .D(_4517_));
 sg13g2_xnor2_1 _5060_ (.Y(_4519_),
    .A(_4509_),
    .B(_4518_));
 sg13g2_buf_1 _5061_ (.A(\generated._26[3] ),
    .X(_4520_));
 sg13g2_inv_1 _5062_ (.Y(_4521_),
    .A(_4520_));
 sg13g2_buf_1 _5063_ (.A(\generated._26[2] ),
    .X(_4522_));
 sg13g2_nor4_1 _5064_ (.A(\generated._26[1] ),
    .B(_4509_),
    .C(_4521_),
    .D(_4522_),
    .Y(_0250_));
 sg13g2_a21o_1 _5065_ (.A2(_0250_),
    .A1(_4518_),
    .B1(net29),
    .X(_0251_));
 sg13g2_nor2_1 _5066_ (.A(_4519_),
    .B(_0251_),
    .Y(_0156_));
 sg13g2_nand2_1 _5067_ (.Y(_0252_),
    .A(\generated._26[1] ),
    .B(_4509_));
 sg13g2_inv_1 _5068_ (.Y(_0253_),
    .A(_4518_));
 sg13g2_nor2_1 _5069_ (.A(_0252_),
    .B(_0253_),
    .Y(_0254_));
 sg13g2_a21oi_1 _5070_ (.A1(_4518_),
    .A2(_4509_),
    .Y(_0255_),
    .B1(\generated._26[1] ));
 sg13g2_nor3_1 _5071_ (.A(_4179_),
    .B(_0254_),
    .C(_0255_),
    .Y(_0157_));
 sg13g2_xnor2_1 _5072_ (.Y(_0256_),
    .A(_4522_),
    .B(_0254_));
 sg13g2_nor2_1 _5073_ (.A(_4179_),
    .B(_0256_),
    .Y(_0158_));
 sg13g2_nand2_1 _5074_ (.Y(_0257_),
    .A(_0254_),
    .B(_4522_));
 sg13g2_xnor2_1 _5075_ (.Y(_0258_),
    .A(_4521_),
    .B(_0257_));
 sg13g2_nor2_1 _5076_ (.A(_0251_),
    .B(_0258_),
    .Y(_0159_));
 sg13g2_nand2_2 _5077_ (.Y(_0259_),
    .A(_0253_),
    .B(_4170_));
 sg13g2_nor2b_1 _5078_ (.A(_0259_),
    .B_N(\generated._324[0] ),
    .Y(_0160_));
 sg13g2_inv_1 _5079_ (.Y(_0260_),
    .A(_4513_));
 sg13g2_nor2_1 _5080_ (.A(\generated._31[1] ),
    .B(\generated._31[0] ),
    .Y(_0261_));
 sg13g2_nor3_1 _5081_ (.A(_0260_),
    .B(_0261_),
    .C(_0259_),
    .Y(_0161_));
 sg13g2_nor2_1 _5082_ (.A(\generated._31[2] ),
    .B(_0260_),
    .Y(_0262_));
 sg13g2_nor3_1 _5083_ (.A(_4514_),
    .B(_0262_),
    .C(net29),
    .Y(_0162_));
 sg13g2_nor2_1 _5084_ (.A(\generated._31[3] ),
    .B(_4514_),
    .Y(_0263_));
 sg13g2_nor3_1 _5085_ (.A(_4516_),
    .B(_0263_),
    .C(net29),
    .Y(_0163_));
 sg13g2_nor2_1 _5086_ (.A(\generated._31[4] ),
    .B(_4516_),
    .Y(_0264_));
 sg13g2_nand2_1 _5087_ (.Y(_0265_),
    .A(_4516_),
    .B(\generated._31[4] ));
 sg13g2_inv_1 _5088_ (.Y(_0266_),
    .A(_0265_));
 sg13g2_nor3_1 _5089_ (.A(_0264_),
    .B(_0266_),
    .C(_0259_),
    .Y(_0164_));
 sg13g2_nor2_1 _5090_ (.A(\generated._31[5] ),
    .B(_0266_),
    .Y(_0267_));
 sg13g2_inv_1 _5091_ (.Y(_0268_),
    .A(\generated._31[5] ));
 sg13g2_nor2_1 _5092_ (.A(_0268_),
    .B(_0265_),
    .Y(_0269_));
 sg13g2_nor3_1 _5093_ (.A(_0267_),
    .B(_0269_),
    .C(_0259_),
    .Y(_0165_));
 sg13g2_nand2_1 _5094_ (.Y(_0270_),
    .A(_0269_),
    .B(_4510_));
 sg13g2_o21ai_1 _5095_ (.B1(\generated._31[6] ),
    .Y(_0271_),
    .A1(_0268_),
    .A2(_0265_));
 sg13g2_a21oi_1 _5096_ (.A1(_0270_),
    .A2(_0271_),
    .Y(_0166_),
    .B1(_0259_));
 sg13g2_a21o_1 _5097_ (.A2(_4220_),
    .A1(\generated._342[1] ),
    .B1(_4221_),
    .X(_0168_));
 sg13g2_inv_1 _5098_ (.Y(_0169_),
    .A(_4226_));
 sg13g2_inv_1 _5099_ (.Y(_0170_),
    .A(_4207_));
 sg13g2_nand4_1 _5100_ (.B(\generated._342[3] ),
    .C(_4196_),
    .A(\generated._342[1] ),
    .Y(_0272_),
    .D(\generated._342[4] ));
 sg13g2_nand2b_1 _5101_ (.Y(_0273_),
    .B(_4210_),
    .A_N(_0272_));
 sg13g2_o21ai_1 _5102_ (.B1(_4208_),
    .Y(_0274_),
    .A1(net91),
    .A2(_0273_));
 sg13g2_a21oi_1 _5103_ (.A1(net91),
    .A2(_0273_),
    .Y(_0172_),
    .B1(_0274_));
 sg13g2_inv_1 _5104_ (.Y(_0275_),
    .A(_4220_));
 sg13g2_nor2b_1 _5105_ (.A(_0275_),
    .B_N(\generated._349[0] ),
    .Y(_0173_));
 sg13g2_nor2_1 _5106_ (.A(\generated._353[1] ),
    .B(\generated._353[0] ),
    .Y(_0276_));
 sg13g2_nor3_1 _5107_ (.A(_4188_),
    .B(_0276_),
    .C(net29),
    .Y(_0174_));
 sg13g2_nand2_1 _5108_ (.Y(_0277_),
    .A(_4187_),
    .B(\generated._353[2] ));
 sg13g2_a21oi_1 _5109_ (.A1(_4190_),
    .A2(_0277_),
    .Y(_0175_),
    .B1(_0275_));
 sg13g2_nor2_1 _5110_ (.A(_4189_),
    .B(_4187_),
    .Y(_0278_));
 sg13g2_nor2_1 _5111_ (.A(\generated._353[3] ),
    .B(_0278_),
    .Y(_0279_));
 sg13g2_and2_1 _5112_ (.A(_0278_),
    .B(\generated._353[3] ),
    .X(_0280_));
 sg13g2_nor3_1 _5113_ (.A(_0279_),
    .B(_0280_),
    .C(_0275_),
    .Y(_0176_));
 sg13g2_xnor2_1 _5114_ (.Y(_0281_),
    .A(\generated._353[4] ),
    .B(_0280_));
 sg13g2_nor2_1 _5115_ (.A(_0281_),
    .B(_0275_),
    .Y(_0177_));
 sg13g2_inv_1 _5116_ (.Y(_0282_),
    .A(_0106_));
 sg13g2_buf_1 _5117_ (.A(\generated._375 ),
    .X(_0283_));
 sg13g2_buf_1 _5118_ (.A(\generated._374 ),
    .X(_0284_));
 sg13g2_nor2_2 _5119_ (.A(_0283_),
    .B(_0284_),
    .Y(_0285_));
 sg13g2_buf_1 _5120_ (.A(_0107_),
    .X(_0286_));
 sg13g2_nor2b_1 _5121_ (.A(_0284_),
    .B_N(_0283_),
    .Y(_0287_));
 sg13g2_buf_1 _5122_ (.A(_0287_),
    .X(_0288_));
 sg13g2_a22oi_1 _5123_ (.Y(_0289_),
    .B1(_0108_),
    .B2(_0288_),
    .A2(_0286_),
    .A1(_0285_));
 sg13g2_buf_1 _5124_ (.A(_0283_),
    .X(_0290_));
 sg13g2_inv_1 _5125_ (.Y(_0291_),
    .A(_0109_));
 sg13g2_nand2_1 _5126_ (.Y(_0292_),
    .A(net87),
    .B(_0110_));
 sg13g2_o21ai_1 _5127_ (.B1(_0292_),
    .Y(_0293_),
    .A1(net87),
    .A2(_0291_));
 sg13g2_buf_1 _5128_ (.A(_0284_),
    .X(_0294_));
 sg13g2_nand2_1 _5129_ (.Y(_0295_),
    .A(_0293_),
    .B(net86));
 sg13g2_and2_1 _5130_ (.A(_0289_),
    .B(_0295_),
    .X(_0296_));
 sg13g2_buf_1 _5131_ (.A(_0296_),
    .X(_0297_));
 sg13g2_inv_1 _5132_ (.Y(_0298_),
    .A(_0297_));
 sg13g2_nor2_1 _5133_ (.A(_0282_),
    .B(_0298_),
    .Y(_0299_));
 sg13g2_inv_1 _5134_ (.Y(_0300_),
    .A(_0299_));
 sg13g2_nand2_1 _5135_ (.Y(_0301_),
    .A(_0298_),
    .B(_0282_));
 sg13g2_nor2_1 _5136_ (.A(\generated._483[1] ),
    .B(\generated._483[0] ),
    .Y(_0302_));
 sg13g2_inv_1 _5137_ (.Y(_0303_),
    .A(_0302_));
 sg13g2_nor3_1 _5138_ (.A(\generated._483[3] ),
    .B(\generated._483[2] ),
    .C(_0303_),
    .Y(_0304_));
 sg13g2_buf_1 _5139_ (.A(_0304_),
    .X(_0305_));
 sg13g2_buf_1 _5140_ (.A(net62),
    .X(_0306_));
 sg13g2_a21oi_1 _5141_ (.A1(_0300_),
    .A2(_0301_),
    .Y(_0178_),
    .B1(net44));
 sg13g2_buf_1 _5142_ (.A(\generated._367 ),
    .X(_0307_));
 sg13g2_nand2_1 _5143_ (.Y(_0308_),
    .A(_0297_),
    .B(_0307_));
 sg13g2_inv_1 _5144_ (.Y(_0309_),
    .A(_0110_));
 sg13g2_nand2_1 _5145_ (.Y(_0310_),
    .A(net87),
    .B(_0090_));
 sg13g2_o21ai_1 _5146_ (.B1(_0310_),
    .Y(_0311_),
    .A1(_0290_),
    .A2(_0309_));
 sg13g2_nor2b_1 _5147_ (.A(_0291_),
    .B_N(_0288_),
    .Y(_0312_));
 sg13g2_a221oi_1 _5148_ (.B2(net86),
    .C1(_0312_),
    .B1(_0311_),
    .A1(_0108_),
    .Y(_0313_),
    .A2(_0285_));
 sg13g2_xnor2_1 _5149_ (.Y(_0314_),
    .A(_0308_),
    .B(_0313_));
 sg13g2_xnor2_1 _5150_ (.Y(_0315_),
    .A(_0063_),
    .B(_0314_));
 sg13g2_nor2_1 _5151_ (.A(_0299_),
    .B(_0315_),
    .Y(_0316_));
 sg13g2_inv_1 _5152_ (.Y(_0317_),
    .A(_0316_));
 sg13g2_inv_1 _5153_ (.Y(_0318_),
    .A(net62));
 sg13g2_buf_1 _5154_ (.A(_0318_),
    .X(_0319_));
 sg13g2_nand2_1 _5155_ (.Y(_0320_),
    .A(_0317_),
    .B(net34));
 sg13g2_a21oi_1 _5156_ (.A1(_0299_),
    .A2(_0315_),
    .Y(_0179_),
    .B1(_0320_));
 sg13g2_inv_1 _5157_ (.Y(_0321_),
    .A(net86));
 sg13g2_buf_1 _5158_ (.A(_0321_),
    .X(_0322_));
 sg13g2_buf_1 _5159_ (.A(net87),
    .X(_0323_));
 sg13g2_inv_1 _5160_ (.Y(_0324_),
    .A(_0090_));
 sg13g2_nor2_1 _5161_ (.A(_0290_),
    .B(_0324_),
    .Y(_0325_));
 sg13g2_a21oi_1 _5162_ (.A1(net75),
    .A2(_0091_),
    .Y(_0326_),
    .B1(_0325_));
 sg13g2_nor2_1 _5163_ (.A(_0321_),
    .B(_0326_),
    .Y(_0327_));
 sg13g2_a21oi_1 _5164_ (.A1(net61),
    .A2(_0293_),
    .Y(_0328_),
    .B1(_0327_));
 sg13g2_nor2_1 _5165_ (.A(_0297_),
    .B(_0313_),
    .Y(_0329_));
 sg13g2_inv_1 _5166_ (.Y(_0330_),
    .A(_0329_));
 sg13g2_nand2_1 _5167_ (.Y(_0331_),
    .A(_0330_),
    .B(_0307_));
 sg13g2_xor2_1 _5168_ (.B(_0331_),
    .A(_0328_),
    .X(_0332_));
 sg13g2_xnor2_1 _5169_ (.Y(_0333_),
    .A(_0064_),
    .B(_0332_));
 sg13g2_buf_1 _5170_ (.A(\generated._390[1] ),
    .X(_0334_));
 sg13g2_inv_1 _5171_ (.Y(_0335_),
    .A(_0334_));
 sg13g2_o21ai_1 _5172_ (.B1(_0317_),
    .Y(_0336_),
    .A1(_0335_),
    .A2(_0314_));
 sg13g2_xnor2_1 _5173_ (.Y(_0337_),
    .A(_0333_),
    .B(_0336_));
 sg13g2_nand2_1 _5174_ (.Y(_0180_),
    .A(_0337_),
    .B(net34));
 sg13g2_inv_1 _5175_ (.Y(_0338_),
    .A(_0091_));
 sg13g2_nor2_1 _5176_ (.A(net75),
    .B(_0338_),
    .Y(_0339_));
 sg13g2_a21oi_1 _5177_ (.A1(net75),
    .A2(_0092_),
    .Y(_0340_),
    .B1(_0339_));
 sg13g2_nor2_1 _5178_ (.A(_0322_),
    .B(_0340_),
    .Y(_0341_));
 sg13g2_a21oi_1 _5179_ (.A1(net61),
    .A2(_0311_),
    .Y(_0342_),
    .B1(_0341_));
 sg13g2_inv_2 _5180_ (.Y(_0343_),
    .A(_0307_));
 sg13g2_nor2_1 _5181_ (.A(_0328_),
    .B(_0330_),
    .Y(_0344_));
 sg13g2_nor2_1 _5182_ (.A(_0343_),
    .B(_0344_),
    .Y(_0345_));
 sg13g2_xnor2_1 _5183_ (.Y(_0346_),
    .A(_0342_),
    .B(_0345_));
 sg13g2_xnor2_1 _5184_ (.Y(_0347_),
    .A(_0062_),
    .B(_0346_));
 sg13g2_inv_1 _5185_ (.Y(_0348_),
    .A(\generated._390[2] ));
 sg13g2_inv_1 _5186_ (.Y(_0349_),
    .A(_0332_));
 sg13g2_nand2_1 _5187_ (.Y(_0350_),
    .A(_0336_),
    .B(_0333_));
 sg13g2_o21ai_1 _5188_ (.B1(_0350_),
    .Y(_0351_),
    .A1(_0348_),
    .A2(_0349_));
 sg13g2_xnor2_1 _5189_ (.Y(_0352_),
    .A(_0347_),
    .B(_0351_));
 sg13g2_nand2_1 _5190_ (.Y(_0181_),
    .A(_0352_),
    .B(net34));
 sg13g2_inv_1 _5191_ (.Y(_0353_),
    .A(_0092_));
 sg13g2_buf_1 _5192_ (.A(_0093_),
    .X(_0354_));
 sg13g2_nand2_1 _5193_ (.Y(_0355_),
    .A(_0323_),
    .B(_0354_));
 sg13g2_o21ai_1 _5194_ (.B1(_0355_),
    .Y(_0356_),
    .A1(_0323_),
    .A2(_0353_));
 sg13g2_nor2_1 _5195_ (.A(net86),
    .B(_0326_),
    .Y(_0357_));
 sg13g2_a21oi_1 _5196_ (.A1(_0294_),
    .A2(_0356_),
    .Y(_0358_),
    .B1(_0357_));
 sg13g2_inv_1 _5197_ (.Y(_0359_),
    .A(_0344_));
 sg13g2_nor2_1 _5198_ (.A(_0342_),
    .B(_0359_),
    .Y(_0360_));
 sg13g2_nor2_1 _5199_ (.A(_0343_),
    .B(_0360_),
    .Y(_0361_));
 sg13g2_xnor2_1 _5200_ (.Y(_0362_),
    .A(_0358_),
    .B(_0361_));
 sg13g2_xnor2_1 _5201_ (.Y(_0363_),
    .A(_0061_),
    .B(_0362_));
 sg13g2_inv_1 _5202_ (.Y(_0364_),
    .A(_0363_));
 sg13g2_buf_1 _5203_ (.A(\generated._390[3] ),
    .X(_0365_));
 sg13g2_a22oi_1 _5204_ (.Y(_0366_),
    .B1(_0347_),
    .B2(_0351_),
    .A2(_0346_),
    .A1(_0365_));
 sg13g2_nor2_1 _5205_ (.A(_0364_),
    .B(_0366_),
    .Y(_0367_));
 sg13g2_nor2b_1 _5206_ (.A(_0363_),
    .B_N(_0366_),
    .Y(_0368_));
 sg13g2_o21ai_1 _5207_ (.B1(net34),
    .Y(_0182_),
    .A1(_0367_),
    .A2(_0368_));
 sg13g2_buf_1 _5208_ (.A(\generated._390[4] ),
    .X(_0369_));
 sg13g2_a21o_1 _5209_ (.A2(_0362_),
    .A1(_0369_),
    .B1(_0367_),
    .X(_0370_));
 sg13g2_buf_1 _5210_ (.A(_0060_),
    .X(_0371_));
 sg13g2_buf_1 _5211_ (.A(net86),
    .X(_0372_));
 sg13g2_buf_1 _5212_ (.A(net75),
    .X(_0373_));
 sg13g2_inv_1 _5213_ (.Y(_0374_),
    .A(_0094_));
 sg13g2_nor2_1 _5214_ (.A(net60),
    .B(_0354_),
    .Y(_0375_));
 sg13g2_a21oi_1 _5215_ (.A1(net60),
    .A2(_0374_),
    .Y(_0376_),
    .B1(_0375_));
 sg13g2_nor2_1 _5216_ (.A(net74),
    .B(_0340_),
    .Y(_0377_));
 sg13g2_a21oi_1 _5217_ (.A1(net74),
    .A2(_0376_),
    .Y(_0378_),
    .B1(_0377_));
 sg13g2_buf_1 _5218_ (.A(_0343_),
    .X(_0379_));
 sg13g2_inv_1 _5219_ (.Y(_0380_),
    .A(_0360_));
 sg13g2_nor2_1 _5220_ (.A(_0358_),
    .B(_0380_),
    .Y(_0381_));
 sg13g2_nor2_1 _5221_ (.A(net73),
    .B(_0381_),
    .Y(_0382_));
 sg13g2_xnor2_1 _5222_ (.Y(_0383_),
    .A(_0378_),
    .B(_0382_));
 sg13g2_xnor2_1 _5223_ (.Y(_0384_),
    .A(_0371_),
    .B(_0383_));
 sg13g2_o21ai_1 _5224_ (.B1(net34),
    .Y(_0385_),
    .A1(_0384_),
    .A2(_0370_));
 sg13g2_a21oi_1 _5225_ (.A1(_0370_),
    .A2(_0384_),
    .Y(_0183_),
    .B1(_0385_));
 sg13g2_nand2_1 _5226_ (.Y(_0386_),
    .A(net60),
    .B(_0095_));
 sg13g2_o21ai_1 _5227_ (.B1(_0386_),
    .Y(_0387_),
    .A1(net60),
    .A2(_0374_));
 sg13g2_mux2_1 _5228_ (.A0(_0387_),
    .A1(_0356_),
    .S(net61),
    .X(_0388_));
 sg13g2_inv_1 _5229_ (.Y(_0389_),
    .A(_0381_));
 sg13g2_buf_1 _5230_ (.A(_0307_),
    .X(_0390_));
 sg13g2_o21ai_1 _5231_ (.B1(net85),
    .Y(_0391_),
    .A1(_0378_),
    .A2(_0389_));
 sg13g2_xnor2_1 _5232_ (.Y(_0392_),
    .A(_0388_),
    .B(_0391_));
 sg13g2_xnor2_1 _5233_ (.Y(_0393_),
    .A(_0059_),
    .B(_0392_));
 sg13g2_nand2_1 _5234_ (.Y(_0394_),
    .A(_0370_),
    .B(_0384_));
 sg13g2_nand2_1 _5235_ (.Y(_0395_),
    .A(_0383_),
    .B(\generated._390[5] ));
 sg13g2_nand2_1 _5236_ (.Y(_0396_),
    .A(_0394_),
    .B(_0395_));
 sg13g2_o21ai_1 _5237_ (.B1(net34),
    .Y(_0397_),
    .A1(_0393_),
    .A2(_0396_));
 sg13g2_nand2_1 _5238_ (.Y(_0398_),
    .A(_0396_),
    .B(_0393_));
 sg13g2_nor2b_1 _5239_ (.A(_0397_),
    .B_N(_0398_),
    .Y(_0184_));
 sg13g2_nand2_1 _5240_ (.Y(_0399_),
    .A(net74),
    .B(_0095_));
 sg13g2_inv_1 _5241_ (.Y(_0400_),
    .A(_0399_));
 sg13g2_a21oi_1 _5242_ (.A1(_0376_),
    .A2(net61),
    .Y(_0401_),
    .B1(_0400_));
 sg13g2_inv_1 _5243_ (.Y(_0402_),
    .A(_0401_));
 sg13g2_nand3b_1 _5244_ (.B(_0381_),
    .C(_0388_),
    .Y(_0403_),
    .A_N(_0378_));
 sg13g2_buf_1 _5245_ (.A(_0403_),
    .X(_0404_));
 sg13g2_nand2_1 _5246_ (.Y(_0405_),
    .A(_0404_),
    .B(net85));
 sg13g2_xnor2_1 _5247_ (.Y(_0406_),
    .A(_0402_),
    .B(_0405_));
 sg13g2_xnor2_1 _5248_ (.Y(_0407_),
    .A(_0070_),
    .B(_0406_));
 sg13g2_buf_1 _5249_ (.A(\generated._390[6] ),
    .X(_0408_));
 sg13g2_inv_1 _5250_ (.Y(_0409_),
    .A(_0408_));
 sg13g2_inv_1 _5251_ (.Y(_0410_),
    .A(_0392_));
 sg13g2_o21ai_1 _5252_ (.B1(_0398_),
    .Y(_0411_),
    .A1(_0409_),
    .A2(_0410_));
 sg13g2_xnor2_1 _5253_ (.Y(_0412_),
    .A(_0407_),
    .B(_0411_));
 sg13g2_nand2_1 _5254_ (.Y(_0185_),
    .A(_0412_),
    .B(net34));
 sg13g2_a22oi_1 _5255_ (.Y(_0413_),
    .B1(_0407_),
    .B2(_0411_),
    .A2(_0406_),
    .A1(\generated._390[7] ));
 sg13g2_buf_1 _5256_ (.A(_0073_),
    .X(_0414_));
 sg13g2_a21oi_1 _5257_ (.A1(_0387_),
    .A2(net61),
    .Y(_0415_),
    .B1(_0400_));
 sg13g2_o21ai_1 _5258_ (.B1(net85),
    .Y(_0416_),
    .A1(_0401_),
    .A2(_0404_));
 sg13g2_xnor2_1 _5259_ (.Y(_0417_),
    .A(_0415_),
    .B(_0416_));
 sg13g2_xnor2_1 _5260_ (.Y(_0418_),
    .A(_0414_),
    .B(_0417_));
 sg13g2_nor2_1 _5261_ (.A(_0418_),
    .B(_0413_),
    .Y(_0419_));
 sg13g2_inv_1 _5262_ (.Y(_0420_),
    .A(_0419_));
 sg13g2_nand2_1 _5263_ (.Y(_0421_),
    .A(_0420_),
    .B(net34));
 sg13g2_a21oi_1 _5264_ (.A1(_0413_),
    .A2(_0418_),
    .Y(_0186_),
    .B1(_0421_));
 sg13g2_buf_1 _5265_ (.A(_0076_),
    .X(_0422_));
 sg13g2_nor3_1 _5266_ (.A(_0401_),
    .B(_0415_),
    .C(_0404_),
    .Y(_0423_));
 sg13g2_xnor2_1 _5267_ (.Y(_0424_),
    .A(\generated._376 ),
    .B(_0423_));
 sg13g2_nand2_1 _5268_ (.Y(_0425_),
    .A(net73),
    .B(_0095_));
 sg13g2_o21ai_1 _5269_ (.B1(_0425_),
    .Y(_0426_),
    .A1(net73),
    .A2(_0424_));
 sg13g2_xor2_1 _5270_ (.B(_0426_),
    .A(_0422_),
    .X(_0427_));
 sg13g2_inv_1 _5271_ (.Y(_0428_),
    .A(\generated._390[8] ));
 sg13g2_o21ai_1 _5272_ (.B1(_0420_),
    .Y(_0429_),
    .A1(_0428_),
    .A2(_0417_));
 sg13g2_xor2_1 _5273_ (.B(_0429_),
    .A(_0427_),
    .X(_0430_));
 sg13g2_nor2_1 _5274_ (.A(net44),
    .B(_0430_),
    .Y(_0187_));
 sg13g2_a22oi_1 _5275_ (.Y(_0431_),
    .B1(_0063_),
    .B2(_0288_),
    .A2(_0106_),
    .A1(_0285_));
 sg13g2_inv_1 _5276_ (.Y(_0432_),
    .A(_0064_));
 sg13g2_nand2_1 _5277_ (.Y(_0433_),
    .A(_0283_),
    .B(_0062_));
 sg13g2_o21ai_1 _5278_ (.B1(_0433_),
    .Y(_0434_),
    .A1(_0283_),
    .A2(_0432_));
 sg13g2_nand2_1 _5279_ (.Y(_0435_),
    .A(_0434_),
    .B(_0284_));
 sg13g2_nand2_1 _5280_ (.Y(_0436_),
    .A(_0431_),
    .B(_0435_));
 sg13g2_buf_1 _5281_ (.A(_0318_),
    .X(_0437_));
 sg13g2_o21ai_1 _5282_ (.B1(net33),
    .Y(_0438_),
    .A1(_0286_),
    .A2(_0436_));
 sg13g2_a21oi_1 _5283_ (.A1(_0286_),
    .A2(_0436_),
    .Y(_0188_),
    .B1(_0438_));
 sg13g2_buf_1 _5284_ (.A(\generated._497[0] ),
    .X(_0439_));
 sg13g2_inv_1 _5285_ (.Y(_0440_),
    .A(_0439_));
 sg13g2_nor2_1 _5286_ (.A(_0440_),
    .B(_0436_),
    .Y(_0441_));
 sg13g2_buf_1 _5287_ (.A(\generated._377[0] ),
    .X(_0442_));
 sg13g2_inv_1 _5288_ (.Y(_0443_),
    .A(_0436_));
 sg13g2_nand2_1 _5289_ (.Y(_0444_),
    .A(_0443_),
    .B(_0307_));
 sg13g2_inv_1 _5290_ (.Y(_0445_),
    .A(_0062_));
 sg13g2_nand2_1 _5291_ (.Y(_0446_),
    .A(_0283_),
    .B(_0061_));
 sg13g2_o21ai_1 _5292_ (.B1(_0446_),
    .Y(_0447_),
    .A1(net87),
    .A2(_0445_));
 sg13g2_inv_1 _5293_ (.Y(_0448_),
    .A(_0063_));
 sg13g2_nor3_1 _5294_ (.A(net87),
    .B(_0284_),
    .C(_0448_),
    .Y(_0449_));
 sg13g2_a221oi_1 _5295_ (.B2(net86),
    .C1(_0449_),
    .B1(_0447_),
    .A1(_0064_),
    .Y(_0450_),
    .A2(_0288_));
 sg13g2_xnor2_1 _5296_ (.Y(_0451_),
    .A(_0444_),
    .B(_0450_));
 sg13g2_xnor2_1 _5297_ (.Y(_0452_),
    .A(_0442_),
    .B(_0451_));
 sg13g2_inv_1 _5298_ (.Y(_0453_),
    .A(_0452_));
 sg13g2_nor2_1 _5299_ (.A(_0441_),
    .B(_0453_),
    .Y(_0454_));
 sg13g2_nand2_1 _5300_ (.Y(_0455_),
    .A(_0453_),
    .B(_0441_));
 sg13g2_inv_1 _5301_ (.Y(_0456_),
    .A(_0455_));
 sg13g2_nor3_1 _5302_ (.A(_0306_),
    .B(_0454_),
    .C(_0456_),
    .Y(_0189_));
 sg13g2_buf_1 _5303_ (.A(\generated._377[1] ),
    .X(_0457_));
 sg13g2_inv_1 _5304_ (.Y(_0458_),
    .A(_0061_));
 sg13g2_nor2_1 _5305_ (.A(net87),
    .B(_0458_),
    .Y(_0459_));
 sg13g2_a21oi_1 _5306_ (.A1(net87),
    .A2(_0371_),
    .Y(_0460_),
    .B1(_0459_));
 sg13g2_nor2_1 _5307_ (.A(_0321_),
    .B(_0460_),
    .Y(_0461_));
 sg13g2_a21oi_1 _5308_ (.A1(_0321_),
    .A2(_0434_),
    .Y(_0462_),
    .B1(_0461_));
 sg13g2_nor2_1 _5309_ (.A(_0443_),
    .B(_0450_),
    .Y(_0463_));
 sg13g2_nor2_1 _5310_ (.A(_0343_),
    .B(_0463_),
    .Y(_0464_));
 sg13g2_xor2_1 _5311_ (.B(_0464_),
    .A(_0462_),
    .X(_0465_));
 sg13g2_xor2_1 _5312_ (.B(_0465_),
    .A(_0457_),
    .X(_0466_));
 sg13g2_inv_1 _5313_ (.Y(_0467_),
    .A(_0108_));
 sg13g2_a21oi_1 _5314_ (.A1(_0467_),
    .A2(_0451_),
    .Y(_0468_),
    .B1(_0456_));
 sg13g2_inv_1 _5315_ (.Y(_0469_),
    .A(_0468_));
 sg13g2_o21ai_1 _5316_ (.B1(_0319_),
    .Y(_0470_),
    .A1(_0466_),
    .A2(_0469_));
 sg13g2_nand2_1 _5317_ (.Y(_0471_),
    .A(_0469_),
    .B(_0466_));
 sg13g2_nor2b_1 _5318_ (.A(_0470_),
    .B_N(_0471_),
    .Y(_0190_));
 sg13g2_nand2_1 _5319_ (.Y(_0472_),
    .A(_0465_),
    .B(_0291_));
 sg13g2_nand2_1 _5320_ (.Y(_0473_),
    .A(_0471_),
    .B(_0472_));
 sg13g2_inv_1 _5321_ (.Y(_0474_),
    .A(\generated._377[2] ));
 sg13g2_inv_1 _5322_ (.Y(_0475_),
    .A(_0059_));
 sg13g2_nand2_1 _5323_ (.Y(_0476_),
    .A(_0475_),
    .B(net75));
 sg13g2_o21ai_1 _5324_ (.B1(_0476_),
    .Y(_0477_),
    .A1(net75),
    .A2(_0371_));
 sg13g2_nor2_1 _5325_ (.A(net61),
    .B(_0477_),
    .Y(_0478_));
 sg13g2_a21oi_1 _5326_ (.A1(net61),
    .A2(_0447_),
    .Y(_0479_),
    .B1(_0478_));
 sg13g2_inv_1 _5327_ (.Y(_0480_),
    .A(_0463_));
 sg13g2_nor2_1 _5328_ (.A(_0462_),
    .B(_0480_),
    .Y(_0481_));
 sg13g2_nor2_1 _5329_ (.A(_0343_),
    .B(_0481_),
    .Y(_0482_));
 sg13g2_xor2_1 _5330_ (.B(_0482_),
    .A(_0479_),
    .X(_0483_));
 sg13g2_xnor2_1 _5331_ (.Y(_0484_),
    .A(_0474_),
    .B(_0483_));
 sg13g2_o21ai_1 _5332_ (.B1(net33),
    .Y(_0485_),
    .A1(_0484_),
    .A2(_0473_));
 sg13g2_a21oi_1 _5333_ (.A1(_0473_),
    .A2(_0484_),
    .Y(_0191_),
    .B1(_0485_));
 sg13g2_nand2_1 _5334_ (.Y(_0486_),
    .A(_0473_),
    .B(_0484_));
 sg13g2_nand2_1 _5335_ (.Y(_0487_),
    .A(_0483_),
    .B(_0309_));
 sg13g2_nand2_1 _5336_ (.Y(_0488_),
    .A(_0486_),
    .B(_0487_));
 sg13g2_inv_1 _5337_ (.Y(_0489_),
    .A(\generated._377[3] ));
 sg13g2_nand2_1 _5338_ (.Y(_0490_),
    .A(net75),
    .B(_0070_));
 sg13g2_o21ai_1 _5339_ (.B1(_0490_),
    .Y(_0491_),
    .A1(net75),
    .A2(_0475_));
 sg13g2_nor2_1 _5340_ (.A(net86),
    .B(_0460_),
    .Y(_0492_));
 sg13g2_a21oi_1 _5341_ (.A1(_0294_),
    .A2(_0491_),
    .Y(_0493_),
    .B1(_0492_));
 sg13g2_inv_1 _5342_ (.Y(_0494_),
    .A(_0481_));
 sg13g2_nor2_1 _5343_ (.A(_0479_),
    .B(_0494_),
    .Y(_0495_));
 sg13g2_nor2_1 _5344_ (.A(_0343_),
    .B(_0495_),
    .Y(_0496_));
 sg13g2_xor2_1 _5345_ (.B(_0496_),
    .A(_0493_),
    .X(_0497_));
 sg13g2_xnor2_1 _5346_ (.Y(_0498_),
    .A(_0489_),
    .B(_0497_));
 sg13g2_o21ai_1 _5347_ (.B1(net33),
    .Y(_0499_),
    .A1(_0498_),
    .A2(_0488_));
 sg13g2_a21oi_1 _5348_ (.A1(_0488_),
    .A2(_0498_),
    .Y(_0192_),
    .B1(_0499_));
 sg13g2_nand2_1 _5349_ (.Y(_0500_),
    .A(_0488_),
    .B(_0498_));
 sg13g2_nand2_1 _5350_ (.Y(_0501_),
    .A(_0497_),
    .B(_0324_));
 sg13g2_nand2_1 _5351_ (.Y(_0502_),
    .A(_0500_),
    .B(_0501_));
 sg13g2_inv_1 _5352_ (.Y(_0503_),
    .A(\generated._377[4] ));
 sg13g2_inv_1 _5353_ (.Y(_0504_),
    .A(_0070_));
 sg13g2_nand2_1 _5354_ (.Y(_0505_),
    .A(_0373_),
    .B(_0414_));
 sg13g2_o21ai_1 _5355_ (.B1(_0505_),
    .Y(_0506_),
    .A1(net60),
    .A2(_0504_));
 sg13g2_nor2_1 _5356_ (.A(net74),
    .B(_0477_),
    .Y(_0507_));
 sg13g2_a21oi_2 _5357_ (.B1(_0507_),
    .Y(_0508_),
    .A2(_0506_),
    .A1(net74));
 sg13g2_inv_1 _5358_ (.Y(_0509_),
    .A(_0495_));
 sg13g2_nor2_1 _5359_ (.A(_0493_),
    .B(_0509_),
    .Y(_0510_));
 sg13g2_nor2_1 _5360_ (.A(_0343_),
    .B(_0510_),
    .Y(_0511_));
 sg13g2_xor2_1 _5361_ (.B(_0511_),
    .A(_0508_),
    .X(_0512_));
 sg13g2_xnor2_1 _5362_ (.Y(_0513_),
    .A(_0503_),
    .B(_0512_));
 sg13g2_o21ai_1 _5363_ (.B1(net33),
    .Y(_0514_),
    .A1(_0513_),
    .A2(_0502_));
 sg13g2_a21oi_1 _5364_ (.A1(_0502_),
    .A2(_0513_),
    .Y(_0193_),
    .B1(_0514_));
 sg13g2_nand2_1 _5365_ (.Y(_0515_),
    .A(_0502_),
    .B(_0513_));
 sg13g2_nand2_1 _5366_ (.Y(_0516_),
    .A(_0512_),
    .B(_0338_));
 sg13g2_nand2_1 _5367_ (.Y(_0517_),
    .A(_0515_),
    .B(_0516_));
 sg13g2_buf_1 _5368_ (.A(\generated._377[5] ),
    .X(_0518_));
 sg13g2_inv_1 _5369_ (.Y(_0519_),
    .A(_0414_));
 sg13g2_nand2_1 _5370_ (.Y(_0520_),
    .A(_0373_),
    .B(_0422_));
 sg13g2_o21ai_1 _5371_ (.B1(_0520_),
    .Y(_0521_),
    .A1(net60),
    .A2(_0519_));
 sg13g2_nor2b_1 _5372_ (.A(_0372_),
    .B_N(_0491_),
    .Y(_0522_));
 sg13g2_a21oi_1 _5373_ (.A1(_0372_),
    .A2(_0521_),
    .Y(_0523_),
    .B1(_0522_));
 sg13g2_inv_1 _5374_ (.Y(_0524_),
    .A(_0510_));
 sg13g2_nor2_1 _5375_ (.A(_0508_),
    .B(_0524_),
    .Y(_0525_));
 sg13g2_nor2_1 _5376_ (.A(_0379_),
    .B(_0525_),
    .Y(_0526_));
 sg13g2_xor2_1 _5377_ (.B(_0526_),
    .A(_0523_),
    .X(_0527_));
 sg13g2_xor2_1 _5378_ (.B(_0527_),
    .A(_0518_),
    .X(_0528_));
 sg13g2_o21ai_1 _5379_ (.B1(_0437_),
    .Y(_0529_),
    .A1(_0528_),
    .A2(_0517_));
 sg13g2_a21oi_1 _5380_ (.A1(_0517_),
    .A2(_0528_),
    .Y(_0194_),
    .B1(_0529_));
 sg13g2_buf_1 _5381_ (.A(\generated._377[6] ),
    .X(_0530_));
 sg13g2_nand2_1 _5382_ (.Y(_0531_),
    .A(net74),
    .B(_0422_));
 sg13g2_inv_1 _5383_ (.Y(_0532_),
    .A(_0531_));
 sg13g2_a21oi_1 _5384_ (.A1(_0506_),
    .A2(_0322_),
    .Y(_0533_),
    .B1(_0532_));
 sg13g2_nor3_1 _5385_ (.A(_0508_),
    .B(_0523_),
    .C(_0524_),
    .Y(_0534_));
 sg13g2_nor2_1 _5386_ (.A(net73),
    .B(_0534_),
    .Y(_0535_));
 sg13g2_xnor2_1 _5387_ (.Y(_0536_),
    .A(_0533_),
    .B(_0535_));
 sg13g2_xnor2_1 _5388_ (.Y(_0537_),
    .A(_0530_),
    .B(_0536_));
 sg13g2_nand2_1 _5389_ (.Y(_0538_),
    .A(_0517_),
    .B(_0528_));
 sg13g2_nand2_1 _5390_ (.Y(_0539_),
    .A(_0527_),
    .B(_0353_));
 sg13g2_nand2_1 _5391_ (.Y(_0540_),
    .A(_0538_),
    .B(_0539_));
 sg13g2_nor2_1 _5392_ (.A(_0537_),
    .B(_0540_),
    .Y(_0541_));
 sg13g2_nand2_1 _5393_ (.Y(_0542_),
    .A(_0540_),
    .B(_0537_));
 sg13g2_inv_1 _5394_ (.Y(_0543_),
    .A(_0542_));
 sg13g2_nor3_1 _5395_ (.A(net44),
    .B(_0541_),
    .C(_0543_),
    .Y(_0195_));
 sg13g2_inv_1 _5396_ (.Y(_0544_),
    .A(\generated._377[7] ));
 sg13g2_a21oi_1 _5397_ (.A1(_0521_),
    .A2(net61),
    .Y(_0545_),
    .B1(_0532_));
 sg13g2_inv_1 _5398_ (.Y(_0546_),
    .A(_0534_));
 sg13g2_nor2_1 _5399_ (.A(_0533_),
    .B(_0546_),
    .Y(_0547_));
 sg13g2_nor2_1 _5400_ (.A(_0379_),
    .B(_0547_),
    .Y(_0548_));
 sg13g2_xnor2_1 _5401_ (.Y(_0549_),
    .A(_0545_),
    .B(_0548_));
 sg13g2_xnor2_1 _5402_ (.Y(_0550_),
    .A(_0544_),
    .B(_0549_));
 sg13g2_nor2_1 _5403_ (.A(_0354_),
    .B(_0536_),
    .Y(_0551_));
 sg13g2_nor2_1 _5404_ (.A(_0551_),
    .B(_0543_),
    .Y(_0552_));
 sg13g2_nor2_1 _5405_ (.A(_0550_),
    .B(_0552_),
    .Y(_0553_));
 sg13g2_a21oi_1 _5406_ (.A1(_0552_),
    .A2(_0550_),
    .Y(_0554_),
    .B1(_0305_));
 sg13g2_nor2b_1 _5407_ (.A(_0553_),
    .B_N(_0554_),
    .Y(_0196_));
 sg13g2_nor2_1 _5408_ (.A(_0094_),
    .B(_0549_),
    .Y(_0555_));
 sg13g2_nor2_1 _5409_ (.A(_0555_),
    .B(_0553_),
    .Y(_0556_));
 sg13g2_inv_1 _5410_ (.Y(_0557_),
    .A(_0547_));
 sg13g2_o21ai_1 _5411_ (.B1(\generated._390[9] ),
    .Y(_0558_),
    .A1(_0545_),
    .A2(_0557_));
 sg13g2_inv_1 _5412_ (.Y(_0559_),
    .A(\generated._390[9] ));
 sg13g2_nand3b_1 _5413_ (.B(_0547_),
    .C(_0559_),
    .Y(_0560_),
    .A_N(_0545_));
 sg13g2_nand3_1 _5414_ (.B(_0390_),
    .C(_0560_),
    .A(_0558_),
    .Y(_0561_));
 sg13g2_o21ai_1 _5415_ (.B1(_0561_),
    .Y(_0562_),
    .A1(_0422_),
    .A2(_0390_));
 sg13g2_xnor2_1 _5416_ (.Y(_0563_),
    .A(\generated._376 ),
    .B(_0562_));
 sg13g2_o21ai_1 _5417_ (.B1(_0437_),
    .Y(_0564_),
    .A1(_0563_),
    .A2(_0556_));
 sg13g2_a21oi_1 _5418_ (.A1(_0556_),
    .A2(_0563_),
    .Y(_0197_),
    .B1(_0564_));
 sg13g2_buf_1 _5419_ (.A(\generated._506 ),
    .X(_0565_));
 sg13g2_buf_2 _5420_ (.A(\generated._505 ),
    .X(_0566_));
 sg13g2_nor2_2 _5421_ (.A(_0565_),
    .B(_0566_),
    .Y(_0567_));
 sg13g2_inv_1 _5422_ (.Y(_0568_),
    .A(_0565_));
 sg13g2_nor2_2 _5423_ (.A(_0566_),
    .B(_0568_),
    .Y(_0569_));
 sg13g2_a22oi_1 _5424_ (.Y(_0570_),
    .B1(_0071_),
    .B2(_0569_),
    .A2(_0065_),
    .A1(_0567_));
 sg13g2_inv_1 _5425_ (.Y(_0571_),
    .A(_0077_));
 sg13g2_buf_1 _5426_ (.A(_0074_),
    .X(_0572_));
 sg13g2_nor2_1 _5427_ (.A(_0565_),
    .B(_0572_),
    .Y(_0573_));
 sg13g2_a21oi_1 _5428_ (.A1(_0565_),
    .A2(_0571_),
    .Y(_0574_),
    .B1(_0573_));
 sg13g2_nand2_1 _5429_ (.Y(_0575_),
    .A(_0574_),
    .B(_0566_));
 sg13g2_nand2_1 _5430_ (.Y(_0576_),
    .A(_0570_),
    .B(_0575_));
 sg13g2_nor2_1 _5431_ (.A(\generated._61[1] ),
    .B(\generated._61[0] ),
    .Y(_0577_));
 sg13g2_inv_1 _5432_ (.Y(_0578_),
    .A(\generated._61[2] ));
 sg13g2_inv_1 _5433_ (.Y(_0579_),
    .A(\generated._61[3] ));
 sg13g2_nand3_1 _5434_ (.B(_0578_),
    .C(_0579_),
    .A(_0577_),
    .Y(_0580_));
 sg13g2_buf_1 _5435_ (.A(_0580_),
    .X(_0581_));
 sg13g2_buf_1 _5436_ (.A(net72),
    .X(_0582_));
 sg13g2_o21ai_1 _5437_ (.B1(_0582_),
    .Y(_0583_),
    .A1(_0067_),
    .A2(_0576_));
 sg13g2_a21oi_1 _5438_ (.A1(_0067_),
    .A2(_0576_),
    .Y(_0198_),
    .B1(_0583_));
 sg13g2_inv_2 _5439_ (.Y(_0584_),
    .A(net72));
 sg13g2_buf_1 _5440_ (.A(_0584_),
    .X(_0585_));
 sg13g2_buf_1 _5441_ (.A(\generated._62[0] ),
    .X(_0586_));
 sg13g2_inv_1 _5442_ (.Y(_0587_),
    .A(_0586_));
 sg13g2_nor2_1 _5443_ (.A(_0587_),
    .B(_0576_),
    .Y(_0588_));
 sg13g2_buf_1 _5444_ (.A(\generated._508[0] ),
    .X(_0589_));
 sg13g2_inv_1 _5445_ (.Y(_0590_),
    .A(_0576_));
 sg13g2_buf_1 _5446_ (.A(\generated._499 ),
    .X(_0591_));
 sg13g2_nand2_1 _5447_ (.Y(_0592_),
    .A(_0590_),
    .B(_0591_));
 sg13g2_buf_1 _5448_ (.A(_0565_),
    .X(_0593_));
 sg13g2_buf_1 _5449_ (.A(_0079_),
    .X(_0594_));
 sg13g2_nand2_1 _5450_ (.Y(_0595_),
    .A(net84),
    .B(_0594_));
 sg13g2_o21ai_1 _5451_ (.B1(_0595_),
    .Y(_0596_),
    .A1(_0593_),
    .A2(_0571_));
 sg13g2_inv_1 _5452_ (.Y(_0597_),
    .A(_0071_));
 sg13g2_nor3_1 _5453_ (.A(_0593_),
    .B(_0566_),
    .C(_0597_),
    .Y(_0598_));
 sg13g2_a221oi_1 _5454_ (.B2(_0566_),
    .C1(_0598_),
    .B1(_0596_),
    .A1(_0572_),
    .Y(_0599_),
    .A2(_0569_));
 sg13g2_xnor2_1 _5455_ (.Y(_0600_),
    .A(_0592_),
    .B(_0599_));
 sg13g2_xnor2_1 _5456_ (.Y(_0601_),
    .A(_0589_),
    .B(_0600_));
 sg13g2_inv_1 _5457_ (.Y(_0602_),
    .A(_0601_));
 sg13g2_nor2_1 _5458_ (.A(_0588_),
    .B(_0602_),
    .Y(_0603_));
 sg13g2_nand2_1 _5459_ (.Y(_0604_),
    .A(_0602_),
    .B(_0588_));
 sg13g2_inv_1 _5460_ (.Y(_0605_),
    .A(_0604_));
 sg13g2_nor3_1 _5461_ (.A(net43),
    .B(_0603_),
    .C(_0605_),
    .Y(_0199_));
 sg13g2_inv_1 _5462_ (.Y(_0606_),
    .A(\generated._508[1] ));
 sg13g2_buf_1 _5463_ (.A(_0566_),
    .X(_0607_));
 sg13g2_inv_1 _5464_ (.Y(_0608_),
    .A(net83));
 sg13g2_buf_1 _5465_ (.A(_0608_),
    .X(_0609_));
 sg13g2_buf_1 _5466_ (.A(net84),
    .X(_0610_));
 sg13g2_inv_1 _5467_ (.Y(_0611_),
    .A(_0081_));
 sg13g2_nand2_1 _5468_ (.Y(_0612_),
    .A(_0611_),
    .B(net84));
 sg13g2_o21ai_1 _5469_ (.B1(_0612_),
    .Y(_0613_),
    .A1(net71),
    .A2(_0594_));
 sg13g2_nor2_1 _5470_ (.A(_0608_),
    .B(_0613_),
    .Y(_0614_));
 sg13g2_a21oi_1 _5471_ (.A1(net58),
    .A2(_0574_),
    .Y(_0615_),
    .B1(_0614_));
 sg13g2_buf_1 _5472_ (.A(_0591_),
    .X(_0616_));
 sg13g2_inv_1 _5473_ (.Y(_0617_),
    .A(net82));
 sg13g2_buf_1 _5474_ (.A(_0617_),
    .X(_0618_));
 sg13g2_nor2_1 _5475_ (.A(_0590_),
    .B(_0599_),
    .Y(_0619_));
 sg13g2_nor2_1 _5476_ (.A(net57),
    .B(_0619_),
    .Y(_0620_));
 sg13g2_xor2_1 _5477_ (.B(_0620_),
    .A(_0615_),
    .X(_0621_));
 sg13g2_xnor2_1 _5478_ (.Y(_0622_),
    .A(_0606_),
    .B(_0621_));
 sg13g2_buf_1 _5479_ (.A(_0066_),
    .X(_0623_));
 sg13g2_inv_1 _5480_ (.Y(_0624_),
    .A(_0623_));
 sg13g2_a21oi_1 _5481_ (.A1(_0624_),
    .A2(_0600_),
    .Y(_0625_),
    .B1(_0605_));
 sg13g2_inv_1 _5482_ (.Y(_0626_),
    .A(_0625_));
 sg13g2_buf_1 _5483_ (.A(net72),
    .X(_0627_));
 sg13g2_o21ai_1 _5484_ (.B1(_0627_),
    .Y(_0628_),
    .A1(_0622_),
    .A2(_0626_));
 sg13g2_nand2_1 _5485_ (.Y(_0629_),
    .A(_0626_),
    .B(_0622_));
 sg13g2_nor2b_1 _5486_ (.A(_0628_),
    .B_N(_0629_),
    .Y(_0200_));
 sg13g2_inv_1 _5487_ (.Y(_0630_),
    .A(_0068_));
 sg13g2_nand2_1 _5488_ (.Y(_0631_),
    .A(_0621_),
    .B(_0630_));
 sg13g2_nand2_1 _5489_ (.Y(_0632_),
    .A(_0629_),
    .B(_0631_));
 sg13g2_inv_1 _5490_ (.Y(_0633_),
    .A(\generated._508[2] ));
 sg13g2_buf_1 _5491_ (.A(_0083_),
    .X(_0634_));
 sg13g2_nor2_1 _5492_ (.A(_0610_),
    .B(_0611_),
    .Y(_0635_));
 sg13g2_a21oi_1 _5493_ (.A1(_0610_),
    .A2(_0634_),
    .Y(_0636_),
    .B1(_0635_));
 sg13g2_nor2_1 _5494_ (.A(net58),
    .B(_0636_),
    .Y(_0637_));
 sg13g2_a21oi_1 _5495_ (.A1(net58),
    .A2(_0596_),
    .Y(_0638_),
    .B1(_0637_));
 sg13g2_inv_1 _5496_ (.Y(_0639_),
    .A(_0619_));
 sg13g2_nor2_1 _5497_ (.A(_0615_),
    .B(_0639_),
    .Y(_0640_));
 sg13g2_nor2_1 _5498_ (.A(net57),
    .B(_0640_),
    .Y(_0641_));
 sg13g2_xor2_1 _5499_ (.B(_0641_),
    .A(_0638_),
    .X(_0642_));
 sg13g2_xnor2_1 _5500_ (.Y(_0643_),
    .A(_0633_),
    .B(_0642_));
 sg13g2_o21ai_1 _5501_ (.B1(_0582_),
    .Y(_0644_),
    .A1(_0643_),
    .A2(_0632_));
 sg13g2_a21oi_1 _5502_ (.A1(_0632_),
    .A2(_0643_),
    .Y(_0201_),
    .B1(_0644_));
 sg13g2_inv_1 _5503_ (.Y(_0645_),
    .A(\generated._508[3] ));
 sg13g2_inv_1 _5504_ (.Y(_0646_),
    .A(_0085_));
 sg13g2_nor2_1 _5505_ (.A(net71),
    .B(_0634_),
    .Y(_0647_));
 sg13g2_a21oi_1 _5506_ (.A1(net71),
    .A2(_0646_),
    .Y(_0648_),
    .B1(_0647_));
 sg13g2_nor2_1 _5507_ (.A(net83),
    .B(_0613_),
    .Y(_0649_));
 sg13g2_a21oi_1 _5508_ (.A1(net83),
    .A2(_0648_),
    .Y(_0650_),
    .B1(_0649_));
 sg13g2_inv_1 _5509_ (.Y(_0651_),
    .A(_0640_));
 sg13g2_nor2_1 _5510_ (.A(_0638_),
    .B(_0651_),
    .Y(_0652_));
 sg13g2_nor2_1 _5511_ (.A(_0618_),
    .B(_0652_),
    .Y(_0653_));
 sg13g2_xor2_1 _5512_ (.B(_0653_),
    .A(_0650_),
    .X(_0654_));
 sg13g2_xnor2_1 _5513_ (.Y(_0655_),
    .A(_0645_),
    .B(_0654_));
 sg13g2_nand2_1 _5514_ (.Y(_0656_),
    .A(_0632_),
    .B(_0643_));
 sg13g2_inv_1 _5515_ (.Y(_0657_),
    .A(_0069_));
 sg13g2_nand2_1 _5516_ (.Y(_0658_),
    .A(_0642_),
    .B(_0657_));
 sg13g2_nand2_1 _5517_ (.Y(_0659_),
    .A(_0656_),
    .B(_0658_));
 sg13g2_nor2_1 _5518_ (.A(_0655_),
    .B(_0659_),
    .Y(_0660_));
 sg13g2_nand2_1 _5519_ (.Y(_0661_),
    .A(_0659_),
    .B(_0655_));
 sg13g2_inv_1 _5520_ (.Y(_0662_),
    .A(_0661_));
 sg13g2_nor3_1 _5521_ (.A(net43),
    .B(_0660_),
    .C(_0662_),
    .Y(_0202_));
 sg13g2_inv_1 _5522_ (.Y(_0663_),
    .A(\generated._508[4] ));
 sg13g2_buf_1 _5523_ (.A(net83),
    .X(_0664_));
 sg13g2_buf_1 _5524_ (.A(net71),
    .X(_0665_));
 sg13g2_buf_1 _5525_ (.A(_0086_),
    .X(_0666_));
 sg13g2_nand2_1 _5526_ (.Y(_0667_),
    .A(net55),
    .B(_0666_));
 sg13g2_o21ai_1 _5527_ (.B1(_0667_),
    .Y(_0668_),
    .A1(net55),
    .A2(_0646_));
 sg13g2_nor2_1 _5528_ (.A(net70),
    .B(_0636_),
    .Y(_0669_));
 sg13g2_a21oi_2 _5529_ (.B1(_0669_),
    .Y(_0670_),
    .A2(_0668_),
    .A1(net70));
 sg13g2_inv_1 _5530_ (.Y(_0671_),
    .A(_0652_));
 sg13g2_nor2_1 _5531_ (.A(_0650_),
    .B(_0671_),
    .Y(_0672_));
 sg13g2_nor2_1 _5532_ (.A(net57),
    .B(_0672_),
    .Y(_0673_));
 sg13g2_xor2_1 _5533_ (.B(_0673_),
    .A(_0670_),
    .X(_0674_));
 sg13g2_xnor2_1 _5534_ (.Y(_0675_),
    .A(_0663_),
    .B(_0674_));
 sg13g2_inv_1 _5535_ (.Y(_0676_),
    .A(_0072_));
 sg13g2_a21oi_1 _5536_ (.A1(_0676_),
    .A2(_0654_),
    .Y(_0677_),
    .B1(_0662_));
 sg13g2_inv_1 _5537_ (.Y(_0678_),
    .A(_0677_));
 sg13g2_nor2_1 _5538_ (.A(_0675_),
    .B(_0678_),
    .Y(_0679_));
 sg13g2_nand2_1 _5539_ (.Y(_0680_),
    .A(_0678_),
    .B(_0675_));
 sg13g2_inv_1 _5540_ (.Y(_0681_),
    .A(_0680_));
 sg13g2_nor3_1 _5541_ (.A(_0585_),
    .B(_0679_),
    .C(_0681_),
    .Y(_0203_));
 sg13g2_inv_1 _5542_ (.Y(_0682_),
    .A(_0075_));
 sg13g2_a21oi_1 _5543_ (.A1(_0682_),
    .A2(_0674_),
    .Y(_0683_),
    .B1(_0681_));
 sg13g2_inv_1 _5544_ (.Y(_0684_),
    .A(_0683_));
 sg13g2_buf_1 _5545_ (.A(\generated._508[5] ),
    .X(_0685_));
 sg13g2_inv_1 _5546_ (.Y(_0686_),
    .A(_0666_));
 sg13g2_buf_1 _5547_ (.A(_0087_),
    .X(_0687_));
 sg13g2_nand2_1 _5548_ (.Y(_0688_),
    .A(net55),
    .B(_0687_));
 sg13g2_o21ai_1 _5549_ (.B1(_0688_),
    .Y(_0689_),
    .A1(net55),
    .A2(_0686_));
 sg13g2_nor2b_1 _5550_ (.A(net70),
    .B_N(_0648_),
    .Y(_0690_));
 sg13g2_a21oi_1 _5551_ (.A1(net70),
    .A2(_0689_),
    .Y(_0691_),
    .B1(_0690_));
 sg13g2_buf_1 _5552_ (.A(net57),
    .X(_0692_));
 sg13g2_inv_1 _5553_ (.Y(_0693_),
    .A(_0672_));
 sg13g2_nor2_1 _5554_ (.A(_0670_),
    .B(_0693_),
    .Y(_0694_));
 sg13g2_nor2_1 _5555_ (.A(_0692_),
    .B(_0694_),
    .Y(_0695_));
 sg13g2_xor2_1 _5556_ (.B(_0695_),
    .A(_0691_),
    .X(_0696_));
 sg13g2_xor2_1 _5557_ (.B(_0696_),
    .A(_0685_),
    .X(_0697_));
 sg13g2_o21ai_1 _5558_ (.B1(net59),
    .Y(_0698_),
    .A1(_0697_),
    .A2(_0684_));
 sg13g2_a21oi_1 _5559_ (.A1(_0684_),
    .A2(_0697_),
    .Y(_0204_),
    .B1(_0698_));
 sg13g2_nand2_1 _5560_ (.Y(_0699_),
    .A(net70),
    .B(_0687_));
 sg13g2_inv_1 _5561_ (.Y(_0700_),
    .A(_0699_));
 sg13g2_a21oi_1 _5562_ (.A1(_0668_),
    .A2(net58),
    .Y(_0701_),
    .B1(_0700_));
 sg13g2_nor3_1 _5563_ (.A(_0670_),
    .B(_0691_),
    .C(_0693_),
    .Y(_0702_));
 sg13g2_nor2_1 _5564_ (.A(_0692_),
    .B(_0702_),
    .Y(_0703_));
 sg13g2_xnor2_1 _5565_ (.Y(_0704_),
    .A(_0701_),
    .B(_0703_));
 sg13g2_xnor2_1 _5566_ (.Y(_0705_),
    .A(\generated._508[6] ),
    .B(_0704_));
 sg13g2_nand2_1 _5567_ (.Y(_0706_),
    .A(_0684_),
    .B(_0697_));
 sg13g2_inv_1 _5568_ (.Y(_0707_),
    .A(_0078_));
 sg13g2_nand2_1 _5569_ (.Y(_0708_),
    .A(_0696_),
    .B(_0707_));
 sg13g2_nand2_1 _5570_ (.Y(_0709_),
    .A(_0706_),
    .B(_0708_));
 sg13g2_nor2_1 _5571_ (.A(_0705_),
    .B(_0709_),
    .Y(_0710_));
 sg13g2_nand2_1 _5572_ (.Y(_0711_),
    .A(_0709_),
    .B(_0705_));
 sg13g2_inv_1 _5573_ (.Y(_0712_),
    .A(_0711_));
 sg13g2_nor3_1 _5574_ (.A(net43),
    .B(_0710_),
    .C(_0712_),
    .Y(_0205_));
 sg13g2_inv_1 _5575_ (.Y(_0713_),
    .A(\generated._508[7] ));
 sg13g2_a21oi_2 _5576_ (.B1(_0700_),
    .Y(_0714_),
    .A2(net58),
    .A1(_0689_));
 sg13g2_inv_1 _5577_ (.Y(_0715_),
    .A(_0702_));
 sg13g2_nor2_1 _5578_ (.A(_0701_),
    .B(_0715_),
    .Y(_0716_));
 sg13g2_nor2_1 _5579_ (.A(net42),
    .B(_0716_),
    .Y(_0717_));
 sg13g2_xor2_1 _5580_ (.B(_0717_),
    .A(_0714_),
    .X(_0718_));
 sg13g2_xnor2_1 _5581_ (.Y(_0719_),
    .A(_0713_),
    .B(_0718_));
 sg13g2_buf_1 _5582_ (.A(_0080_),
    .X(_0720_));
 sg13g2_nor2_1 _5583_ (.A(_0720_),
    .B(_0704_),
    .Y(_0721_));
 sg13g2_nor2_1 _5584_ (.A(_0721_),
    .B(_0712_),
    .Y(_0722_));
 sg13g2_inv_1 _5585_ (.Y(_0723_),
    .A(_0722_));
 sg13g2_nor2_1 _5586_ (.A(_0719_),
    .B(_0723_),
    .Y(_0724_));
 sg13g2_nand2_1 _5587_ (.Y(_0725_),
    .A(_0723_),
    .B(_0719_));
 sg13g2_inv_1 _5588_ (.Y(_0726_),
    .A(_0725_));
 sg13g2_nor3_1 _5589_ (.A(net43),
    .B(_0724_),
    .C(_0726_),
    .Y(_0206_));
 sg13g2_inv_1 _5590_ (.Y(_0727_),
    .A(_0082_));
 sg13g2_a21oi_1 _5591_ (.A1(_0727_),
    .A2(_0718_),
    .Y(_0728_),
    .B1(_0726_));
 sg13g2_buf_1 _5592_ (.A(\generated._507 ),
    .X(_0729_));
 sg13g2_inv_1 _5593_ (.Y(_0730_),
    .A(_0716_));
 sg13g2_nor3_1 _5594_ (.A(\generated._558[9] ),
    .B(_0714_),
    .C(_0730_),
    .Y(_0731_));
 sg13g2_o21ai_1 _5595_ (.B1(\generated._558[9] ),
    .Y(_0732_),
    .A1(_0714_),
    .A2(_0730_));
 sg13g2_nand3b_1 _5596_ (.B(_0732_),
    .C(net82),
    .Y(_0733_),
    .A_N(_0731_));
 sg13g2_o21ai_1 _5597_ (.B1(_0733_),
    .Y(_0734_),
    .A1(net82),
    .A2(_0687_));
 sg13g2_xnor2_1 _5598_ (.Y(_0735_),
    .A(_0729_),
    .B(_0734_));
 sg13g2_o21ai_1 _5599_ (.B1(net59),
    .Y(_0736_),
    .A1(_0735_),
    .A2(_0728_));
 sg13g2_a21oi_1 _5600_ (.A1(_0728_),
    .A2(_0735_),
    .Y(_0207_),
    .B1(_0736_));
 sg13g2_buf_2 _5601_ (.A(\generated._840 ),
    .X(_0737_));
 sg13g2_buf_1 _5602_ (.A(\generated._839 ),
    .X(_0738_));
 sg13g2_nor2_1 _5603_ (.A(_0737_),
    .B(_0738_),
    .Y(_0739_));
 sg13g2_buf_1 _5604_ (.A(_0738_),
    .X(_0740_));
 sg13g2_inv_1 _5605_ (.Y(_0741_),
    .A(_0737_));
 sg13g2_nor2_2 _5606_ (.A(net81),
    .B(_0741_),
    .Y(_0742_));
 sg13g2_a22oi_1 _5607_ (.Y(_0743_),
    .B1(_0041_),
    .B2(_0742_),
    .A2(_0101_),
    .A1(_0739_));
 sg13g2_buf_1 _5608_ (.A(_0737_),
    .X(_0744_));
 sg13g2_inv_1 _5609_ (.Y(_0745_),
    .A(_0035_));
 sg13g2_nor2_1 _5610_ (.A(net80),
    .B(_0040_),
    .Y(_0746_));
 sg13g2_a21oi_1 _5611_ (.A1(net80),
    .A2(_0745_),
    .Y(_0747_),
    .B1(_0746_));
 sg13g2_nand2_1 _5612_ (.Y(_0748_),
    .A(_0747_),
    .B(net81));
 sg13g2_and2_1 _5613_ (.A(_0743_),
    .B(_0748_),
    .X(_0749_));
 sg13g2_inv_1 _5614_ (.Y(_0750_),
    .A(_0749_));
 sg13g2_nor2_1 _5615_ (.A(\generated._69[1] ),
    .B(\generated._69[0] ),
    .Y(_0751_));
 sg13g2_inv_1 _5616_ (.Y(_0752_),
    .A(\generated._69[2] ));
 sg13g2_inv_1 _5617_ (.Y(_0753_),
    .A(\generated._69[3] ));
 sg13g2_nand3_1 _5618_ (.B(_0752_),
    .C(_0753_),
    .A(_0751_),
    .Y(_0754_));
 sg13g2_buf_1 _5619_ (.A(_0754_),
    .X(_0755_));
 sg13g2_buf_1 _5620_ (.A(_0755_),
    .X(_0756_));
 sg13g2_o21ai_1 _5621_ (.B1(net54),
    .Y(_0757_),
    .A1(_0102_),
    .A2(_0750_));
 sg13g2_a21oi_1 _5622_ (.A1(_0102_),
    .A2(_0750_),
    .Y(_0208_),
    .B1(_0757_));
 sg13g2_inv_1 _5623_ (.Y(_0758_),
    .A(_0755_));
 sg13g2_buf_1 _5624_ (.A(_0758_),
    .X(_0759_));
 sg13g2_buf_1 _5625_ (.A(\generated._421[1] ),
    .X(_0760_));
 sg13g2_inv_1 _5626_ (.Y(_0761_),
    .A(_0760_));
 sg13g2_nor2_1 _5627_ (.A(_0761_),
    .B(_0750_),
    .Y(_0762_));
 sg13g2_buf_2 _5628_ (.A(\generated._64[1] ),
    .X(_0763_));
 sg13g2_nand2_1 _5629_ (.Y(_0764_),
    .A(net80),
    .B(_0042_));
 sg13g2_o21ai_1 _5630_ (.B1(_0764_),
    .Y(_0765_),
    .A1(net80),
    .A2(_0745_));
 sg13g2_inv_1 _5631_ (.Y(_0766_),
    .A(_0739_));
 sg13g2_nor2b_1 _5632_ (.A(_0766_),
    .B_N(_0041_),
    .Y(_0767_));
 sg13g2_a221oi_1 _5633_ (.B2(net81),
    .C1(_0767_),
    .B1(_0765_),
    .A1(_0040_),
    .Y(_0768_),
    .A2(_0742_));
 sg13g2_nor4_1 _5634_ (.A(\generated._67[3] ),
    .B(\generated._67[2] ),
    .C(\generated._67[1] ),
    .D(\generated._67[0] ),
    .Y(_0769_));
 sg13g2_nor4_1 _5635_ (.A(\generated._67[7] ),
    .B(\generated._67[6] ),
    .C(\generated._67[5] ),
    .D(\generated._67[4] ),
    .Y(_0770_));
 sg13g2_nor2_1 _5636_ (.A(\generated._67[8] ),
    .B(\generated._67[9] ),
    .Y(_0771_));
 sg13g2_nand3_1 _5637_ (.B(_0770_),
    .C(_0771_),
    .A(_0769_),
    .Y(_0772_));
 sg13g2_inv_1 _5638_ (.Y(_0773_),
    .A(_0039_));
 sg13g2_nand2_1 _5639_ (.Y(_0774_),
    .A(_0772_),
    .B(_0773_));
 sg13g2_buf_1 _5640_ (.A(_0774_),
    .X(_0775_));
 sg13g2_nor2_1 _5641_ (.A(_0750_),
    .B(net53),
    .Y(_0776_));
 sg13g2_xor2_1 _5642_ (.B(_0776_),
    .A(_0768_),
    .X(_0777_));
 sg13g2_xnor2_1 _5643_ (.Y(_0778_),
    .A(_0763_),
    .B(_0777_));
 sg13g2_inv_1 _5644_ (.Y(_0779_),
    .A(_0778_));
 sg13g2_nor2_1 _5645_ (.A(_0762_),
    .B(_0779_),
    .Y(_0780_));
 sg13g2_nand2_1 _5646_ (.Y(_0781_),
    .A(_0779_),
    .B(_0762_));
 sg13g2_inv_1 _5647_ (.Y(_0782_),
    .A(_0781_));
 sg13g2_nor3_1 _5648_ (.A(net41),
    .B(_0780_),
    .C(_0782_),
    .Y(_0209_));
 sg13g2_buf_1 _5649_ (.A(\generated._64[2] ),
    .X(_0783_));
 sg13g2_inv_1 _5650_ (.Y(_0784_),
    .A(net92));
 sg13g2_inv_1 _5651_ (.Y(_0785_),
    .A(_0738_));
 sg13g2_buf_1 _5652_ (.A(net80),
    .X(_0786_));
 sg13g2_inv_1 _5653_ (.Y(_0787_),
    .A(_0044_));
 sg13g2_nand2_1 _5654_ (.Y(_0788_),
    .A(_0787_),
    .B(net69));
 sg13g2_o21ai_1 _5655_ (.B1(_0788_),
    .Y(_0789_),
    .A1(net69),
    .A2(_0042_));
 sg13g2_nor2_1 _5656_ (.A(_0785_),
    .B(_0789_),
    .Y(_0790_));
 sg13g2_a21oi_1 _5657_ (.A1(_0785_),
    .A2(_0747_),
    .Y(_0791_),
    .B1(_0790_));
 sg13g2_buf_1 _5658_ (.A(net53),
    .X(_0792_));
 sg13g2_nor2_1 _5659_ (.A(_0749_),
    .B(_0768_),
    .Y(_0793_));
 sg13g2_nor2_1 _5660_ (.A(net40),
    .B(_0793_),
    .Y(_0794_));
 sg13g2_xor2_1 _5661_ (.B(_0794_),
    .A(_0791_),
    .X(_0795_));
 sg13g2_xnor2_1 _5662_ (.Y(_0796_),
    .A(_0784_),
    .B(_0795_));
 sg13g2_inv_1 _5663_ (.Y(_0797_),
    .A(_0103_));
 sg13g2_a21oi_1 _5664_ (.A1(_0797_),
    .A2(_0777_),
    .Y(_0798_),
    .B1(_0782_));
 sg13g2_inv_1 _5665_ (.Y(_0799_),
    .A(_0798_));
 sg13g2_o21ai_1 _5666_ (.B1(net54),
    .Y(_0800_),
    .A1(_0796_),
    .A2(_0799_));
 sg13g2_nand2_1 _5667_ (.Y(_0801_),
    .A(_0799_),
    .B(_0796_));
 sg13g2_nor2b_1 _5668_ (.A(_0800_),
    .B_N(_0801_),
    .Y(_0210_));
 sg13g2_inv_1 _5669_ (.Y(_0802_),
    .A(_0101_));
 sg13g2_a22oi_1 _5670_ (.Y(_0803_),
    .B1(_0103_),
    .B2(_0742_),
    .A2(_0102_),
    .A1(_0739_));
 sg13g2_inv_1 _5671_ (.Y(_0804_),
    .A(_0104_));
 sg13g2_nand2_1 _5672_ (.Y(_0805_),
    .A(_0737_),
    .B(_0105_));
 sg13g2_o21ai_1 _5673_ (.B1(_0805_),
    .Y(_0806_),
    .A1(_0737_),
    .A2(_0804_));
 sg13g2_nand2_1 _5674_ (.Y(_0807_),
    .A(_0806_),
    .B(net81));
 sg13g2_and2_1 _5675_ (.A(_0803_),
    .B(_0807_),
    .X(_0808_));
 sg13g2_inv_1 _5676_ (.Y(_0809_),
    .A(_0808_));
 sg13g2_nor2_1 _5677_ (.A(_0802_),
    .B(_0809_),
    .Y(_0810_));
 sg13g2_inv_1 _5678_ (.Y(_0811_),
    .A(_0810_));
 sg13g2_nand2_1 _5679_ (.Y(_0812_),
    .A(_0809_),
    .B(_0802_));
 sg13g2_a21oi_1 _5680_ (.A1(_0811_),
    .A2(_0812_),
    .Y(_0211_),
    .B1(net41));
 sg13g2_inv_1 _5681_ (.Y(_0813_),
    .A(_0036_));
 sg13g2_nor2_1 _5682_ (.A(net80),
    .B(_0105_),
    .Y(_0814_));
 sg13g2_a21oi_1 _5683_ (.A1(_0744_),
    .A2(_0813_),
    .Y(_0815_),
    .B1(_0814_));
 sg13g2_nor2_1 _5684_ (.A(_0797_),
    .B(_0766_),
    .Y(_0816_));
 sg13g2_a221oi_1 _5685_ (.B2(net81),
    .C1(_0816_),
    .B1(_0815_),
    .A1(_0104_),
    .Y(_0817_),
    .A2(_0742_));
 sg13g2_nor2_1 _5686_ (.A(_0809_),
    .B(net53),
    .Y(_0818_));
 sg13g2_xnor2_1 _5687_ (.Y(_0819_),
    .A(_0817_),
    .B(_0818_));
 sg13g2_xor2_1 _5688_ (.B(_0819_),
    .A(_0041_),
    .X(_0820_));
 sg13g2_nor2_1 _5689_ (.A(_0810_),
    .B(_0820_),
    .Y(_0821_));
 sg13g2_inv_1 _5690_ (.Y(_0822_),
    .A(_0821_));
 sg13g2_nand2_1 _5691_ (.Y(_0823_),
    .A(_0822_),
    .B(net54));
 sg13g2_a21oi_1 _5692_ (.A1(_0810_),
    .A2(_0820_),
    .Y(_0212_),
    .B1(_0823_));
 sg13g2_nor2_1 _5693_ (.A(_0744_),
    .B(_0813_),
    .Y(_0824_));
 sg13g2_a21oi_1 _5694_ (.A1(net69),
    .A2(_0037_),
    .Y(_0825_),
    .B1(_0824_));
 sg13g2_nor2_1 _5695_ (.A(_0785_),
    .B(_0825_),
    .Y(_0826_));
 sg13g2_a21oi_1 _5696_ (.A1(_0785_),
    .A2(_0806_),
    .Y(_0827_),
    .B1(_0826_));
 sg13g2_nor2_1 _5697_ (.A(_0808_),
    .B(_0817_),
    .Y(_0828_));
 sg13g2_nor2_1 _5698_ (.A(_0775_),
    .B(_0828_),
    .Y(_0829_));
 sg13g2_xnor2_1 _5699_ (.Y(_0830_),
    .A(_0827_),
    .B(_0829_));
 sg13g2_xnor2_1 _5700_ (.Y(_0831_),
    .A(_0040_),
    .B(_0830_));
 sg13g2_a21o_1 _5701_ (.A2(_0819_),
    .A1(\generated._67[1] ),
    .B1(_0821_),
    .X(_0832_));
 sg13g2_o21ai_1 _5702_ (.B1(net54),
    .Y(_0833_),
    .A1(_0831_),
    .A2(_0832_));
 sg13g2_nand2_1 _5703_ (.Y(_0834_),
    .A(_0832_),
    .B(_0831_));
 sg13g2_nor2b_1 _5704_ (.A(_0833_),
    .B_N(_0834_),
    .Y(_0213_));
 sg13g2_nand2_1 _5705_ (.Y(_0835_),
    .A(_0737_),
    .B(net81));
 sg13g2_xor2_1 _5706_ (.B(_0835_),
    .A(_0048_),
    .X(_0836_));
 sg13g2_nor2_1 _5707_ (.A(net41),
    .B(_0836_),
    .Y(_0214_));
 sg13g2_buf_1 _5708_ (.A(\generated._430[10] ),
    .X(_0837_));
 sg13g2_nand2_1 _5709_ (.Y(_0838_),
    .A(_0835_),
    .B(_0837_));
 sg13g2_inv_1 _5710_ (.Y(_0839_),
    .A(net53));
 sg13g2_nand2_1 _5711_ (.Y(_0840_),
    .A(_0839_),
    .B(_0785_));
 sg13g2_nand2_1 _5712_ (.Y(_0841_),
    .A(net53),
    .B(_0766_));
 sg13g2_o21ai_1 _5713_ (.B1(_0841_),
    .Y(_0842_),
    .A1(_0737_),
    .A2(_0840_));
 sg13g2_buf_1 _5714_ (.A(_0842_),
    .X(_0843_));
 sg13g2_nand2_2 _5715_ (.Y(_0844_),
    .A(_0843_),
    .B(_0835_));
 sg13g2_xor2_1 _5716_ (.B(_0844_),
    .A(\generated._430[11] ),
    .X(_0845_));
 sg13g2_nor2_1 _5717_ (.A(_0838_),
    .B(_0845_),
    .Y(_0846_));
 sg13g2_inv_1 _5718_ (.Y(_0847_),
    .A(_0846_));
 sg13g2_nand2_1 _5719_ (.Y(_0848_),
    .A(_0847_),
    .B(net54));
 sg13g2_a21oi_1 _5720_ (.A1(_0838_),
    .A2(_0845_),
    .Y(_0215_),
    .B1(_0848_));
 sg13g2_o21ai_1 _5721_ (.B1(_0847_),
    .Y(_0849_),
    .A1(_0056_),
    .A2(_0844_));
 sg13g2_inv_1 _5722_ (.Y(_0850_),
    .A(\generated._430[12] ));
 sg13g2_nor2_1 _5723_ (.A(_0742_),
    .B(net53),
    .Y(_0851_));
 sg13g2_a21oi_1 _5724_ (.A1(net80),
    .A2(net53),
    .Y(_0852_),
    .B1(_0851_));
 sg13g2_xnor2_1 _5725_ (.Y(_0853_),
    .A(_0850_),
    .B(_0852_));
 sg13g2_o21ai_1 _5726_ (.B1(net54),
    .Y(_0854_),
    .A1(_0853_),
    .A2(_0849_));
 sg13g2_a21oi_1 _5727_ (.A1(_0849_),
    .A2(_0853_),
    .Y(_0216_),
    .B1(_0854_));
 sg13g2_inv_1 _5728_ (.Y(_0855_),
    .A(\generated._430[13] ));
 sg13g2_xnor2_1 _5729_ (.Y(_0856_),
    .A(_0855_),
    .B(_0844_));
 sg13g2_inv_1 _5730_ (.Y(_0857_),
    .A(_0856_));
 sg13g2_nand2_1 _5731_ (.Y(_0858_),
    .A(_0849_),
    .B(_0853_));
 sg13g2_inv_1 _5732_ (.Y(_0859_),
    .A(_0055_));
 sg13g2_nand2_1 _5733_ (.Y(_0860_),
    .A(_0852_),
    .B(_0859_));
 sg13g2_nand2_1 _5734_ (.Y(_0861_),
    .A(_0858_),
    .B(_0860_));
 sg13g2_nor2_1 _5735_ (.A(_0857_),
    .B(_0861_),
    .Y(_0862_));
 sg13g2_nand2_1 _5736_ (.Y(_0863_),
    .A(_0861_),
    .B(_0857_));
 sg13g2_inv_1 _5737_ (.Y(_0864_),
    .A(_0863_));
 sg13g2_nor3_1 _5738_ (.A(net41),
    .B(_0862_),
    .C(_0864_),
    .Y(_0217_));
 sg13g2_nor2_1 _5739_ (.A(_0057_),
    .B(_0844_),
    .Y(_0865_));
 sg13g2_nor2_1 _5740_ (.A(_0865_),
    .B(_0864_),
    .Y(_0866_));
 sg13g2_buf_1 _5741_ (.A(\generated._430[14] ),
    .X(_0867_));
 sg13g2_xnor2_1 _5742_ (.Y(_0868_),
    .A(net80),
    .B(net81));
 sg13g2_inv_1 _5743_ (.Y(_0869_),
    .A(_0868_));
 sg13g2_o21ai_1 _5744_ (.B1(_0841_),
    .Y(_0870_),
    .A1(net53),
    .A2(_0869_));
 sg13g2_xnor2_1 _5745_ (.Y(_0871_),
    .A(_0867_),
    .B(_0870_));
 sg13g2_nor2_1 _5746_ (.A(_0871_),
    .B(_0866_),
    .Y(_0872_));
 sg13g2_inv_1 _5747_ (.Y(_0873_),
    .A(_0872_));
 sg13g2_nand2_1 _5748_ (.Y(_0874_),
    .A(_0873_),
    .B(net54));
 sg13g2_a21oi_1 _5749_ (.A1(_0866_),
    .A2(_0871_),
    .Y(_0218_),
    .B1(_0874_));
 sg13g2_xnor2_1 _5750_ (.Y(_0875_),
    .A(_0740_),
    .B(net40));
 sg13g2_xnor2_1 _5751_ (.Y(_0876_),
    .A(\generated._430[15] ),
    .B(_0875_));
 sg13g2_inv_1 _5752_ (.Y(_0877_),
    .A(_0054_));
 sg13g2_a21o_1 _5753_ (.A2(_0870_),
    .A1(_0877_),
    .B1(_0872_),
    .X(_0878_));
 sg13g2_nor2_1 _5754_ (.A(_0876_),
    .B(_0878_),
    .Y(_0879_));
 sg13g2_nand2_1 _5755_ (.Y(_0880_),
    .A(_0878_),
    .B(_0876_));
 sg13g2_inv_1 _5756_ (.Y(_0881_),
    .A(_0880_));
 sg13g2_nor3_1 _5757_ (.A(net41),
    .B(_0879_),
    .C(_0881_),
    .Y(_0219_));
 sg13g2_xor2_1 _5758_ (.B(_0843_),
    .A(\generated._430[16] ),
    .X(_0882_));
 sg13g2_buf_1 _5759_ (.A(_0053_),
    .X(_0883_));
 sg13g2_inv_1 _5760_ (.Y(_0884_),
    .A(_0883_));
 sg13g2_inv_1 _5761_ (.Y(_0885_),
    .A(_0875_));
 sg13g2_a21oi_1 _5762_ (.A1(_0884_),
    .A2(_0885_),
    .Y(_0886_),
    .B1(_0881_));
 sg13g2_nor2_1 _5763_ (.A(_0882_),
    .B(_0886_),
    .Y(_0887_));
 sg13g2_a21oi_1 _5764_ (.A1(_0886_),
    .A2(_0882_),
    .Y(_0888_),
    .B1(_0758_));
 sg13g2_nor2b_1 _5765_ (.A(_0887_),
    .B_N(_0888_),
    .Y(_0220_));
 sg13g2_buf_1 _5766_ (.A(net40),
    .X(_0889_));
 sg13g2_xnor2_1 _5767_ (.Y(_0890_),
    .A(\generated._430[17] ),
    .B(net32));
 sg13g2_inv_1 _5768_ (.Y(_0891_),
    .A(_0052_));
 sg13g2_inv_1 _5769_ (.Y(_0892_),
    .A(_0843_));
 sg13g2_a21oi_1 _5770_ (.A1(_0891_),
    .A2(_0892_),
    .Y(_0893_),
    .B1(_0887_));
 sg13g2_inv_1 _5771_ (.Y(_0894_),
    .A(_0893_));
 sg13g2_nor2_1 _5772_ (.A(_0890_),
    .B(_0894_),
    .Y(_0895_));
 sg13g2_nand2_1 _5773_ (.Y(_0896_),
    .A(_0894_),
    .B(_0890_));
 sg13g2_inv_1 _5774_ (.Y(_0897_),
    .A(_0896_));
 sg13g2_nor3_1 _5775_ (.A(_0759_),
    .B(_0895_),
    .C(_0897_),
    .Y(_0221_));
 sg13g2_xnor2_1 _5776_ (.Y(_0898_),
    .A(\generated._430[18] ),
    .B(net32));
 sg13g2_inv_1 _5777_ (.Y(_0899_),
    .A(_0058_));
 sg13g2_a21oi_1 _5778_ (.A1(_0899_),
    .A2(_0839_),
    .Y(_0900_),
    .B1(_0897_));
 sg13g2_inv_1 _5779_ (.Y(_0901_),
    .A(_0900_));
 sg13g2_nor2_1 _5780_ (.A(_0898_),
    .B(_0901_),
    .Y(_0902_));
 sg13g2_nand2_1 _5781_ (.Y(_0903_),
    .A(_0901_),
    .B(_0898_));
 sg13g2_inv_1 _5782_ (.Y(_0904_),
    .A(_0903_));
 sg13g2_nor3_1 _5783_ (.A(_0759_),
    .B(_0902_),
    .C(_0904_),
    .Y(_0222_));
 sg13g2_inv_1 _5784_ (.Y(_0905_),
    .A(\generated._430[19] ));
 sg13g2_inv_1 _5785_ (.Y(_0906_),
    .A(_0051_));
 sg13g2_nor3_1 _5786_ (.A(_0906_),
    .B(_0889_),
    .C(_0904_),
    .Y(_0907_));
 sg13g2_a21oi_1 _5787_ (.A1(_0889_),
    .A2(_0904_),
    .Y(_0908_),
    .B1(_0907_));
 sg13g2_buf_1 _5788_ (.A(_0755_),
    .X(_0909_));
 sg13g2_o21ai_1 _5789_ (.B1(net52),
    .Y(_0910_),
    .A1(_0905_),
    .A2(_0908_));
 sg13g2_a21oi_1 _5790_ (.A1(_0905_),
    .A2(_0908_),
    .Y(_0223_),
    .B1(_0910_));
 sg13g2_nor2b_1 _5791_ (.A(net44),
    .B_N(\generated._391[0] ),
    .Y(_0242_));
 sg13g2_nand2_1 _5792_ (.Y(_0911_),
    .A(net60),
    .B(net86));
 sg13g2_a21oi_1 _5793_ (.A1(_0911_),
    .A2(net74),
    .Y(_0912_),
    .B1(_0288_));
 sg13g2_nor2_1 _5794_ (.A(_0912_),
    .B(_0306_),
    .Y(_0243_));
 sg13g2_nor2b_1 _5795_ (.A(net43),
    .B_N(\generated._559[0] ),
    .Y(_0244_));
 sg13g2_nand2_2 _5796_ (.Y(_0913_),
    .A(net55),
    .B(net83));
 sg13g2_a21oi_1 _5797_ (.A1(_0913_),
    .A2(net70),
    .Y(_0914_),
    .B1(_0569_));
 sg13g2_nor2_1 _5798_ (.A(_0914_),
    .B(net43),
    .Y(_0245_));
 sg13g2_nor2b_1 _5799_ (.A(net41),
    .B_N(\generated._887[0] ),
    .Y(_0246_));
 sg13g2_nor2_1 _5800_ (.A(_0868_),
    .B(net41),
    .Y(_0247_));
 sg13g2_nor2b_1 _5801_ (.A(net36),
    .B_N(\generated._1021[0] ),
    .Y(_0248_));
 sg13g2_nor2_1 _5802_ (.A(_4446_),
    .B(_4327_),
    .Y(_0249_));
 sg13g2_nor2_1 _5803_ (.A(_4215_),
    .B(_4212_),
    .Y(_0127_));
 sg13g2_nor2_1 _5804_ (.A(_4215_),
    .B(_4222_),
    .Y(_0128_));
 sg13g2_nor2_1 _5805_ (.A(_4215_),
    .B(_4226_),
    .Y(_0129_));
 sg13g2_nor2_1 _5806_ (.A(net77),
    .B(_4364_),
    .Y(_0915_));
 sg13g2_a21oi_1 _5807_ (.A1(net77),
    .A2(_0028_),
    .Y(_0916_),
    .B1(_0915_));
 sg13g2_nor2_1 _5808_ (.A(net78),
    .B(_0916_),
    .Y(_0917_));
 sg13g2_a21oi_1 _5809_ (.A1(net78),
    .A2(_4345_),
    .Y(_0918_),
    .B1(_0917_));
 sg13g2_inv_1 _5810_ (.Y(_0919_),
    .A(_4370_));
 sg13g2_nor2_1 _5811_ (.A(_4368_),
    .B(_0919_),
    .Y(_0920_));
 sg13g2_nor2_1 _5812_ (.A(_4369_),
    .B(_0920_),
    .Y(_0921_));
 sg13g2_xnor2_1 _5813_ (.Y(_0922_),
    .A(_0918_),
    .B(_0921_));
 sg13g2_xor2_1 _5814_ (.B(_0922_),
    .A(\generated._1020[3] ),
    .X(_0923_));
 sg13g2_inv_1 _5815_ (.Y(_0924_),
    .A(_0923_));
 sg13g2_nand2_1 _5816_ (.Y(_0925_),
    .A(_4372_),
    .B(_4382_));
 sg13g2_nand2_1 _5817_ (.Y(_0926_),
    .A(_4379_),
    .B(_0925_));
 sg13g2_xnor2_1 _5818_ (.Y(_0927_),
    .A(_0924_),
    .B(_0926_));
 sg13g2_buf_1 _5819_ (.A(_4324_),
    .X(_0928_));
 sg13g2_nor2_1 _5820_ (.A(\generated._402[1] ),
    .B(\generated._402[2] ),
    .Y(_0929_));
 sg13g2_nor2_1 _5821_ (.A(_4251_),
    .B(_0929_),
    .Y(_0930_));
 sg13g2_inv_1 _5822_ (.Y(_0931_),
    .A(_0930_));
 sg13g2_nand2_1 _5823_ (.Y(_0932_),
    .A(_0929_),
    .B(_4251_));
 sg13g2_a21oi_1 _5824_ (.A1(_0931_),
    .A2(_0932_),
    .Y(_0933_),
    .B1(net65));
 sg13g2_a21oi_1 _5825_ (.A1(_0927_),
    .A2(net51),
    .Y(\generated._1019[3] ),
    .B1(_0933_));
 sg13g2_inv_1 _5826_ (.Y(_0934_),
    .A(_4253_));
 sg13g2_xnor2_1 _5827_ (.Y(_0935_),
    .A(_0934_),
    .B(_0930_));
 sg13g2_nor2_1 _5828_ (.A(_0100_),
    .B(_0922_),
    .Y(_0936_));
 sg13g2_a21oi_1 _5829_ (.A1(_0926_),
    .A2(_0924_),
    .Y(_0937_),
    .B1(_0936_));
 sg13g2_inv_1 _5830_ (.Y(_0938_),
    .A(_0030_));
 sg13g2_nor2_1 _5831_ (.A(net77),
    .B(_0028_),
    .Y(_0939_));
 sg13g2_a21oi_1 _5832_ (.A1(net64),
    .A2(_0938_),
    .Y(_0940_),
    .B1(_0939_));
 sg13g2_nor2_1 _5833_ (.A(net89),
    .B(_4366_),
    .Y(_0941_));
 sg13g2_a21oi_1 _5834_ (.A1(net89),
    .A2(_0940_),
    .Y(_0942_),
    .B1(_0941_));
 sg13g2_inv_1 _5835_ (.Y(_0943_),
    .A(_0920_));
 sg13g2_nor2_1 _5836_ (.A(_0918_),
    .B(_0943_),
    .Y(_0944_));
 sg13g2_nor2_1 _5837_ (.A(_4369_),
    .B(_0944_),
    .Y(_0945_));
 sg13g2_xor2_1 _5838_ (.B(_0945_),
    .A(_0942_),
    .X(_0946_));
 sg13g2_xor2_1 _5839_ (.B(_0946_),
    .A(\generated._1020[4] ),
    .X(_0947_));
 sg13g2_inv_1 _5840_ (.Y(_0948_),
    .A(_0947_));
 sg13g2_a21oi_1 _5841_ (.A1(_0937_),
    .A2(_0948_),
    .Y(_0949_),
    .B1(net48));
 sg13g2_nor2_1 _5842_ (.A(_0948_),
    .B(_0937_),
    .Y(_0950_));
 sg13g2_inv_1 _5843_ (.Y(_0951_),
    .A(_0950_));
 sg13g2_nand2_1 _5844_ (.Y(_0952_),
    .A(_0949_),
    .B(_0951_));
 sg13g2_o21ai_1 _5845_ (.B1(_0952_),
    .Y(\generated._1019[4] ),
    .A1(net51),
    .A2(_0935_));
 sg13g2_nand2_1 _5846_ (.Y(_0953_),
    .A(net64),
    .B(_0031_));
 sg13g2_o21ai_1 _5847_ (.B1(_0953_),
    .Y(_0954_),
    .A1(net64),
    .A2(_0938_));
 sg13g2_nor2_1 _5848_ (.A(net89),
    .B(_0916_),
    .Y(_0955_));
 sg13g2_a21oi_1 _5849_ (.A1(net89),
    .A2(_0954_),
    .Y(_0956_),
    .B1(_0955_));
 sg13g2_inv_1 _5850_ (.Y(_0957_),
    .A(_0944_));
 sg13g2_nor2_1 _5851_ (.A(_0942_),
    .B(_0957_),
    .Y(_0958_));
 sg13g2_nor2_1 _5852_ (.A(_4444_),
    .B(_0958_),
    .Y(_0959_));
 sg13g2_xor2_1 _5853_ (.B(_0959_),
    .A(_0956_),
    .X(_0960_));
 sg13g2_xor2_1 _5854_ (.B(_0960_),
    .A(\generated._1020[5] ),
    .X(_0961_));
 sg13g2_inv_1 _5855_ (.Y(_0962_),
    .A(_0961_));
 sg13g2_a21o_1 _5856_ (.A2(_0946_),
    .A1(_4402_),
    .B1(_0950_),
    .X(_0963_));
 sg13g2_inv_1 _5857_ (.Y(_0964_),
    .A(_0963_));
 sg13g2_nor2_1 _5858_ (.A(_0962_),
    .B(_0964_),
    .Y(_0965_));
 sg13g2_o21ai_1 _5859_ (.B1(_4324_),
    .Y(_0966_),
    .A1(_0961_),
    .A2(_0963_));
 sg13g2_o21ai_1 _5860_ (.B1(_0033_),
    .Y(_0967_),
    .A1(_4253_),
    .A2(_0931_));
 sg13g2_xnor2_1 _5861_ (.Y(_0968_),
    .A(_4257_),
    .B(_0967_));
 sg13g2_nand2_1 _5862_ (.Y(_0969_),
    .A(_0968_),
    .B(_4326_));
 sg13g2_o21ai_1 _5863_ (.B1(_0969_),
    .Y(\generated._1019[5] ),
    .A1(_0965_),
    .A2(_0966_));
 sg13g2_a21oi_1 _5864_ (.A1(_0931_),
    .A2(_0934_),
    .Y(_0970_),
    .B1(_4257_));
 sg13g2_xnor2_1 _5865_ (.Y(_0971_),
    .A(_4256_),
    .B(_0970_));
 sg13g2_inv_1 _5866_ (.Y(_0972_),
    .A(_0971_));
 sg13g2_inv_1 _5867_ (.Y(_0973_),
    .A(_0018_));
 sg13g2_a21oi_1 _5868_ (.A1(_0973_),
    .A2(_0960_),
    .Y(_0974_),
    .B1(_0965_));
 sg13g2_inv_1 _5869_ (.Y(_0975_),
    .A(_0031_));
 sg13g2_nand2_1 _5870_ (.Y(_0976_),
    .A(net64),
    .B(_0020_));
 sg13g2_o21ai_1 _5871_ (.B1(_0976_),
    .Y(_0977_),
    .A1(net64),
    .A2(_0975_));
 sg13g2_mux2_1 _5872_ (.A0(_0977_),
    .A1(_0940_),
    .S(_4362_),
    .X(_0978_));
 sg13g2_inv_1 _5873_ (.Y(_0979_),
    .A(_0956_));
 sg13g2_a21oi_1 _5874_ (.A1(_0958_),
    .A2(_0979_),
    .Y(_0980_),
    .B1(net35));
 sg13g2_xnor2_1 _5875_ (.Y(_0981_),
    .A(_0978_),
    .B(_0980_));
 sg13g2_xor2_1 _5876_ (.B(_0981_),
    .A(\generated._1020[6] ),
    .X(_0982_));
 sg13g2_inv_1 _5877_ (.Y(_0983_),
    .A(_0982_));
 sg13g2_a21oi_1 _5878_ (.A1(_0974_),
    .A2(_0983_),
    .Y(_0984_),
    .B1(_4326_));
 sg13g2_nor2_1 _5879_ (.A(_0983_),
    .B(_0974_),
    .Y(_0985_));
 sg13g2_inv_1 _5880_ (.Y(_0986_),
    .A(_0985_));
 sg13g2_nand2_1 _5881_ (.Y(_0987_),
    .A(_0984_),
    .B(_0986_));
 sg13g2_o21ai_1 _5882_ (.B1(_0987_),
    .Y(\generated._1019[6] ),
    .A1(net51),
    .A2(_0972_));
 sg13g2_nand2_1 _5883_ (.Y(_0988_),
    .A(net89),
    .B(_0020_));
 sg13g2_inv_1 _5884_ (.Y(_0989_),
    .A(_0988_));
 sg13g2_a21oi_2 _5885_ (.B1(_0989_),
    .Y(_0990_),
    .A2(net78),
    .A1(_0954_));
 sg13g2_nand3b_1 _5886_ (.B(_0958_),
    .C(_0978_),
    .Y(_0991_),
    .A_N(_0956_));
 sg13g2_buf_1 _5887_ (.A(_0991_),
    .X(_0992_));
 sg13g2_nand2_1 _5888_ (.Y(_0993_),
    .A(_0992_),
    .B(net47));
 sg13g2_xnor2_1 _5889_ (.Y(_0994_),
    .A(_0990_),
    .B(_0993_));
 sg13g2_xnor2_1 _5890_ (.Y(_0995_),
    .A(\generated._1020[7] ),
    .B(_0994_));
 sg13g2_inv_1 _5891_ (.Y(_0996_),
    .A(_0995_));
 sg13g2_inv_1 _5892_ (.Y(_0997_),
    .A(_0019_));
 sg13g2_a21o_1 _5893_ (.A2(_0981_),
    .A1(_0997_),
    .B1(_0985_),
    .X(_0998_));
 sg13g2_xnor2_1 _5894_ (.Y(_0999_),
    .A(_0996_),
    .B(_0998_));
 sg13g2_nand3_1 _5895_ (.B(\generated._402[5] ),
    .C(\generated._402[6] ),
    .A(_0967_),
    .Y(_1000_));
 sg13g2_xor2_1 _5896_ (.B(_1000_),
    .A(_0034_),
    .X(_1001_));
 sg13g2_nor2_1 _5897_ (.A(net65),
    .B(_1001_),
    .Y(_1002_));
 sg13g2_a21oi_1 _5898_ (.A1(_0999_),
    .A2(net51),
    .Y(\generated._1019[7] ),
    .B1(_1002_));
 sg13g2_nand3_1 _5899_ (.B(\generated._402[6] ),
    .C(\generated._402[7] ),
    .A(_0970_),
    .Y(_1003_));
 sg13g2_inv_1 _5900_ (.Y(_1004_),
    .A(_1003_));
 sg13g2_a21oi_1 _5901_ (.A1(_0977_),
    .A2(_4362_),
    .Y(_1005_),
    .B1(_0989_));
 sg13g2_o21ai_1 _5902_ (.B1(net47),
    .Y(_1006_),
    .A1(_0990_),
    .A2(_0992_));
 sg13g2_xor2_1 _5903_ (.B(_1006_),
    .A(_1005_),
    .X(_1007_));
 sg13g2_xnor2_1 _5904_ (.Y(_1008_),
    .A(\generated._1020[8] ),
    .B(_1007_));
 sg13g2_nand2_1 _5905_ (.Y(_1009_),
    .A(_0998_),
    .B(_0996_));
 sg13g2_inv_1 _5906_ (.Y(_1010_),
    .A(_0024_));
 sg13g2_nand2_1 _5907_ (.Y(_1011_),
    .A(_0994_),
    .B(_1010_));
 sg13g2_nand2_1 _5908_ (.Y(_1012_),
    .A(_1009_),
    .B(_1011_));
 sg13g2_o21ai_1 _5909_ (.B1(_4324_),
    .Y(_1013_),
    .A1(_1008_),
    .A2(_1012_));
 sg13g2_nand2_1 _5910_ (.Y(_1014_),
    .A(_1012_),
    .B(_1008_));
 sg13g2_nand2b_1 _5911_ (.Y(_1015_),
    .B(_1014_),
    .A_N(_1013_));
 sg13g2_o21ai_1 _5912_ (.B1(_1015_),
    .Y(\generated._1019[8] ),
    .A1(_0928_),
    .A2(_1004_));
 sg13g2_nor3_1 _5913_ (.A(_0990_),
    .B(_1005_),
    .C(_0992_),
    .Y(_1016_));
 sg13g2_a21oi_1 _5914_ (.A1(_1016_),
    .A2(\generated._1070[9] ),
    .Y(_1017_),
    .B1(_4444_));
 sg13g2_o21ai_1 _5915_ (.B1(_1017_),
    .Y(_1018_),
    .A1(\generated._1070[9] ),
    .A2(_1016_));
 sg13g2_nand2_1 _5916_ (.Y(_1019_),
    .A(_1018_),
    .B(_4352_));
 sg13g2_xnor2_1 _5917_ (.Y(_1020_),
    .A(\generated._1020[9] ),
    .B(_1019_));
 sg13g2_o21ai_1 _5918_ (.B1(_1014_),
    .Y(_1021_),
    .A1(_0027_),
    .A2(_1007_));
 sg13g2_xnor2_1 _5919_ (.Y(_1022_),
    .A(_1020_),
    .B(_1021_));
 sg13g2_nor2_1 _5920_ (.A(_0034_),
    .B(_1000_),
    .Y(_1023_));
 sg13g2_nor2_1 _5921_ (.A(_4377_),
    .B(_1023_),
    .Y(_1024_));
 sg13g2_a21oi_1 _5922_ (.A1(_1022_),
    .A2(_0928_),
    .Y(\generated._1019[9] ),
    .B1(_1024_));
 sg13g2_buf_2 _5923_ (.A(\generated._64[3] ),
    .X(_1025_));
 sg13g2_inv_2 _5924_ (.Y(_1026_),
    .A(_1025_));
 sg13g2_buf_2 _5925_ (.A(\generated._64[4] ),
    .X(_1027_));
 sg13g2_buf_2 _5926_ (.A(\generated._64[5] ),
    .X(_1028_));
 sg13g2_xnor2_1 _5927_ (.Y(_1029_),
    .A(_1027_),
    .B(_1028_));
 sg13g2_nand2_1 _5928_ (.Y(_1030_),
    .A(_1027_),
    .B(_1028_));
 sg13g2_o21ai_1 _5929_ (.B1(_1030_),
    .Y(_1031_),
    .A1(_1026_),
    .A2(_1029_));
 sg13g2_buf_1 _5930_ (.A(\generated._64[6] ),
    .X(_1032_));
 sg13g2_inv_1 _5931_ (.Y(_1033_),
    .A(_1032_));
 sg13g2_inv_1 _5932_ (.Y(_1034_),
    .A(_1028_));
 sg13g2_nand2_1 _5933_ (.Y(_1035_),
    .A(_1033_),
    .B(_1034_));
 sg13g2_nand2_1 _5934_ (.Y(_1036_),
    .A(_1032_),
    .B(_1028_));
 sg13g2_a21oi_1 _5935_ (.A1(_1035_),
    .A2(_1036_),
    .Y(_1037_),
    .B1(_1027_));
 sg13g2_nand3_1 _5936_ (.B(_1027_),
    .C(_1036_),
    .A(_1035_),
    .Y(_1038_));
 sg13g2_nand2b_1 _5937_ (.Y(_1039_),
    .B(_1038_),
    .A_N(_1037_));
 sg13g2_xnor2_1 _5938_ (.Y(_1040_),
    .A(_1031_),
    .B(_1039_));
 sg13g2_nor2b_1 _5939_ (.A(_1039_),
    .B_N(_1031_),
    .Y(_1041_));
 sg13g2_a21oi_1 _5940_ (.A1(_1040_),
    .A2(_0763_),
    .Y(_1042_),
    .B1(_1041_));
 sg13g2_nand2_1 _5941_ (.Y(_1043_),
    .A(_1038_),
    .B(_1036_));
 sg13g2_buf_2 _5942_ (.A(\generated._64[7] ),
    .X(_1044_));
 sg13g2_inv_1 _5943_ (.Y(_1045_),
    .A(_1044_));
 sg13g2_nand2_1 _5944_ (.Y(_1046_),
    .A(_1045_),
    .B(_1033_));
 sg13g2_nand2_1 _5945_ (.Y(_1047_),
    .A(_1044_),
    .B(_1032_));
 sg13g2_a21oi_1 _5946_ (.A1(_1046_),
    .A2(_1047_),
    .Y(_1048_),
    .B1(_1028_));
 sg13g2_nand3_1 _5947_ (.B(_1028_),
    .C(_1047_),
    .A(_1046_),
    .Y(_1049_));
 sg13g2_nand2b_1 _5948_ (.Y(_1050_),
    .B(_1049_),
    .A_N(_1048_));
 sg13g2_xnor2_1 _5949_ (.Y(_1051_),
    .A(_1043_),
    .B(_1050_));
 sg13g2_xnor2_1 _5950_ (.Y(_1052_),
    .A(net92),
    .B(_1051_));
 sg13g2_or2_1 _5951_ (.X(_1053_),
    .B(_1052_),
    .A(_1042_));
 sg13g2_nand2_1 _5952_ (.Y(_1054_),
    .A(_1049_),
    .B(_1047_));
 sg13g2_buf_2 _5953_ (.A(\generated._64[8] ),
    .X(_1055_));
 sg13g2_xor2_1 _5954_ (.B(_1044_),
    .A(_1055_),
    .X(_1056_));
 sg13g2_xnor2_1 _5955_ (.Y(_1057_),
    .A(_1032_),
    .B(_1056_));
 sg13g2_xnor2_1 _5956_ (.Y(_1058_),
    .A(_1054_),
    .B(_1057_));
 sg13g2_xnor2_1 _5957_ (.Y(_1059_),
    .A(_1025_),
    .B(_1058_));
 sg13g2_nor2b_1 _5958_ (.A(_1050_),
    .B_N(_1043_),
    .Y(_1060_));
 sg13g2_a21oi_1 _5959_ (.A1(_1051_),
    .A2(net92),
    .Y(_1061_),
    .B1(_1060_));
 sg13g2_xor2_1 _5960_ (.B(_1061_),
    .A(_1059_),
    .X(_1062_));
 sg13g2_nand2b_1 _5961_ (.Y(_1063_),
    .B(_1062_),
    .A_N(_1053_));
 sg13g2_nor2_1 _5962_ (.A(_1059_),
    .B(_1061_),
    .Y(_1064_));
 sg13g2_nor2b_1 _5963_ (.A(_1057_),
    .B_N(_1054_),
    .Y(_1065_));
 sg13g2_a21oi_1 _5964_ (.A1(_1058_),
    .A2(_1025_),
    .Y(_1066_),
    .B1(_1065_));
 sg13g2_buf_2 _5965_ (.A(\generated._64[9] ),
    .X(_1067_));
 sg13g2_xnor2_1 _5966_ (.Y(_1068_),
    .A(_1067_),
    .B(_1056_));
 sg13g2_nor2b_1 _5967_ (.A(_1033_),
    .B_N(_1056_),
    .Y(_1069_));
 sg13g2_a21oi_1 _5968_ (.A1(_1055_),
    .A2(_1044_),
    .Y(_1070_),
    .B1(_1069_));
 sg13g2_xor2_1 _5969_ (.B(_1070_),
    .A(_1068_),
    .X(_1071_));
 sg13g2_xnor2_1 _5970_ (.Y(_1072_),
    .A(_1027_),
    .B(_1071_));
 sg13g2_xnor2_1 _5971_ (.Y(_1073_),
    .A(_1066_),
    .B(_1072_));
 sg13g2_xor2_1 _5972_ (.B(_1073_),
    .A(_1064_),
    .X(_1074_));
 sg13g2_nor2_1 _5973_ (.A(_1063_),
    .B(_1074_),
    .Y(_1075_));
 sg13g2_nand2_1 _5974_ (.Y(_1076_),
    .A(_1074_),
    .B(_1063_));
 sg13g2_nand2b_1 _5975_ (.Y(_1077_),
    .B(_1076_),
    .A_N(_1075_));
 sg13g2_xnor2_1 _5976_ (.Y(_1078_),
    .A(_1026_),
    .B(_1029_));
 sg13g2_inv_1 _5977_ (.Y(_1079_),
    .A(_1027_));
 sg13g2_xor2_1 _5978_ (.B(_1025_),
    .A(_1027_),
    .X(_1080_));
 sg13g2_nand2_1 _5979_ (.Y(_1081_),
    .A(_1080_),
    .B(net92));
 sg13g2_o21ai_1 _5980_ (.B1(_1081_),
    .Y(_1082_),
    .A1(_1079_),
    .A2(_1026_));
 sg13g2_inv_1 _5981_ (.Y(_1083_),
    .A(_1082_));
 sg13g2_nor2_1 _5982_ (.A(_1078_),
    .B(_1083_),
    .Y(_1084_));
 sg13g2_nand2_1 _5983_ (.Y(_1085_),
    .A(_1083_),
    .B(_1078_));
 sg13g2_nand2b_1 _5984_ (.Y(_1086_),
    .B(_1085_),
    .A_N(_1084_));
 sg13g2_xnor2_1 _5985_ (.Y(_1087_),
    .A(_0760_),
    .B(_1086_));
 sg13g2_xnor2_1 _5986_ (.Y(_1088_),
    .A(_0783_),
    .B(_1080_));
 sg13g2_inv_1 _5987_ (.Y(_1089_),
    .A(_0763_));
 sg13g2_nor2_1 _5988_ (.A(_1025_),
    .B(net92),
    .Y(_1090_));
 sg13g2_nand2_1 _5989_ (.Y(_1091_),
    .A(_1025_),
    .B(net92));
 sg13g2_o21ai_1 _5990_ (.B1(_1091_),
    .Y(_1092_),
    .A1(_1089_),
    .A2(_1090_));
 sg13g2_nor2b_1 _5991_ (.A(_1088_),
    .B_N(_1092_),
    .Y(_1093_));
 sg13g2_nand2_1 _5992_ (.Y(_1094_),
    .A(_1087_),
    .B(_1093_));
 sg13g2_a21oi_1 _5993_ (.A1(_1085_),
    .A2(_0760_),
    .Y(_1095_),
    .B1(_1084_));
 sg13g2_xnor2_1 _5994_ (.Y(_1096_),
    .A(_0763_),
    .B(_1040_));
 sg13g2_xor2_1 _5995_ (.B(_1096_),
    .A(_1095_),
    .X(_1097_));
 sg13g2_nor2b_1 _5996_ (.A(_1094_),
    .B_N(_1097_),
    .Y(_1098_));
 sg13g2_inv_1 _5997_ (.Y(_1099_),
    .A(_1098_));
 sg13g2_nor2_1 _5998_ (.A(_1095_),
    .B(_1096_),
    .Y(_1100_));
 sg13g2_xnor2_1 _5999_ (.Y(_1101_),
    .A(_1042_),
    .B(_1052_));
 sg13g2_xor2_1 _6000_ (.B(_1101_),
    .A(_1100_),
    .X(_1102_));
 sg13g2_or2_1 _6001_ (.X(_1103_),
    .B(_1087_),
    .A(_1093_));
 sg13g2_xnor2_1 _6002_ (.Y(_1104_),
    .A(_1092_),
    .B(_1088_));
 sg13g2_inv_1 _6003_ (.Y(_1105_),
    .A(_1104_));
 sg13g2_nand2_1 _6004_ (.Y(_1106_),
    .A(net92),
    .B(_0763_));
 sg13g2_nor2_1 _6005_ (.A(net92),
    .B(_0763_),
    .Y(_1107_));
 sg13g2_nor2b_1 _6006_ (.A(_1107_),
    .B_N(_1106_),
    .Y(_1108_));
 sg13g2_nand3_1 _6007_ (.B(_1026_),
    .C(_0760_),
    .A(_1108_),
    .Y(_1109_));
 sg13g2_o21ai_1 _6008_ (.B1(_1109_),
    .Y(_1110_),
    .A1(_1026_),
    .A2(_1106_));
 sg13g2_nor2b_1 _6009_ (.A(_1105_),
    .B_N(_1110_),
    .Y(_1111_));
 sg13g2_nand4_1 _6010_ (.B(_1097_),
    .C(_1094_),
    .A(_1103_),
    .Y(_1112_),
    .D(_1111_));
 sg13g2_nor4_1 _6011_ (.A(_1025_),
    .B(_0761_),
    .C(_1106_),
    .D(_1105_),
    .Y(_1113_));
 sg13g2_nand3_1 _6012_ (.B(_1097_),
    .C(_1113_),
    .A(_1103_),
    .Y(_1114_));
 sg13g2_nand2b_1 _6013_ (.Y(_1115_),
    .B(_1100_),
    .A_N(_1101_));
 sg13g2_xor2_1 _6014_ (.B(_1062_),
    .A(_1053_),
    .X(_1116_));
 sg13g2_xnor2_1 _6015_ (.Y(_1117_),
    .A(_1115_),
    .B(_1116_));
 sg13g2_a221oi_1 _6016_ (.B2(_1114_),
    .C1(_1117_),
    .B1(_1112_),
    .A1(_1099_),
    .Y(_1118_),
    .A2(_1102_));
 sg13g2_nor2_1 _6017_ (.A(_1099_),
    .B(_1102_),
    .Y(_1119_));
 sg13g2_nand2b_1 _6018_ (.Y(_1120_),
    .B(_1119_),
    .A_N(_1117_));
 sg13g2_o21ai_1 _6019_ (.B1(_1120_),
    .Y(_1121_),
    .A1(_1115_),
    .A2(_1116_));
 sg13g2_or2_1 _6020_ (.X(_1122_),
    .B(_1121_),
    .A(_1118_));
 sg13g2_xor2_1 _6021_ (.B(_1122_),
    .A(_1077_),
    .X(_1123_));
 sg13g2_nand2_1 _6022_ (.Y(_1124_),
    .A(_4409_),
    .B(\generated._1070[2] ));
 sg13g2_nand2_1 _6023_ (.Y(_1125_),
    .A(_4413_),
    .B(_1124_));
 sg13g2_nor2_1 _6024_ (.A(net90),
    .B(_0973_),
    .Y(_1126_));
 sg13g2_a21oi_1 _6025_ (.A1(net77),
    .A2(_0019_),
    .Y(_1127_),
    .B1(_1126_));
 sg13g2_mux2_1 _6026_ (.A0(_1127_),
    .A1(_4393_),
    .S(net78),
    .X(_1128_));
 sg13g2_inv_1 _6027_ (.Y(_1129_),
    .A(_4407_));
 sg13g2_nor2_1 _6028_ (.A(_4406_),
    .B(_1129_),
    .Y(_1130_));
 sg13g2_nor2_1 _6029_ (.A(net46),
    .B(_1130_),
    .Y(_1131_));
 sg13g2_xnor2_1 _6030_ (.Y(_1132_),
    .A(_1128_),
    .B(_1131_));
 sg13g2_xnor2_1 _6031_ (.Y(_1133_),
    .A(_0016_),
    .B(_1132_));
 sg13g2_a21oi_1 _6032_ (.A1(_1125_),
    .A2(_1133_),
    .Y(_1134_),
    .B1(_4325_));
 sg13g2_o21ai_1 _6033_ (.B1(_1134_),
    .Y(_1135_),
    .A1(_1125_),
    .A2(_1133_));
 sg13g2_o21ai_1 _6034_ (.B1(_1135_),
    .Y(\generated._1069[3] ),
    .A1(net51),
    .A2(_1123_));
 sg13g2_nand2_1 _6035_ (.Y(_1136_),
    .A(net77),
    .B(_0024_));
 sg13g2_o21ai_1 _6036_ (.B1(_1136_),
    .Y(_1137_),
    .A1(_4363_),
    .A2(_0997_));
 sg13g2_nor2_1 _6037_ (.A(net93),
    .B(_4404_),
    .Y(_1138_));
 sg13g2_a21oi_1 _6038_ (.A1(net93),
    .A2(_1137_),
    .Y(_1139_),
    .B1(_1138_));
 sg13g2_inv_1 _6039_ (.Y(_1140_),
    .A(_1130_));
 sg13g2_nor2_1 _6040_ (.A(_1128_),
    .B(_1140_),
    .Y(_1141_));
 sg13g2_nor2_1 _6041_ (.A(net46),
    .B(_1141_),
    .Y(_1142_));
 sg13g2_xnor2_1 _6042_ (.Y(_1143_),
    .A(_1139_),
    .B(_1142_));
 sg13g2_xnor2_1 _6043_ (.Y(_1144_),
    .A(_0023_),
    .B(_1143_));
 sg13g2_nand2_1 _6044_ (.Y(_1145_),
    .A(_1125_),
    .B(_1133_));
 sg13g2_nand2_1 _6045_ (.Y(_1146_),
    .A(_1132_),
    .B(\generated._1070[3] ));
 sg13g2_nand2_1 _6046_ (.Y(_1147_),
    .A(_1145_),
    .B(_1146_));
 sg13g2_xor2_1 _6047_ (.B(_1147_),
    .A(_1144_),
    .X(_1148_));
 sg13g2_nand2b_1 _6048_ (.Y(_1149_),
    .B(_1064_),
    .A_N(_1073_));
 sg13g2_or2_1 _6049_ (.X(_1150_),
    .B(_1072_),
    .A(_1066_));
 sg13g2_nor2_1 _6050_ (.A(_1067_),
    .B(_1044_),
    .Y(_1151_));
 sg13g2_inv_1 _6051_ (.Y(_1152_),
    .A(_1151_));
 sg13g2_nand2_1 _6052_ (.Y(_1153_),
    .A(_1067_),
    .B(_1044_));
 sg13g2_inv_1 _6053_ (.Y(_1154_),
    .A(_1153_));
 sg13g2_nor2_1 _6054_ (.A(_1055_),
    .B(_1154_),
    .Y(_1155_));
 sg13g2_a21oi_1 _6055_ (.A1(_1055_),
    .A2(_1152_),
    .Y(_1156_),
    .B1(_1155_));
 sg13g2_xnor2_1 _6056_ (.Y(_1157_),
    .A(_1034_),
    .B(_1156_));
 sg13g2_nor2_1 _6057_ (.A(_1068_),
    .B(_1070_),
    .Y(_1158_));
 sg13g2_a21oi_1 _6058_ (.A1(_1071_),
    .A2(_1027_),
    .Y(_1159_),
    .B1(_1158_));
 sg13g2_xnor2_1 _6059_ (.Y(_1160_),
    .A(_1157_),
    .B(_1159_));
 sg13g2_xor2_1 _6060_ (.B(_1160_),
    .A(_1150_),
    .X(_1161_));
 sg13g2_nor2_1 _6061_ (.A(_1149_),
    .B(_1161_),
    .Y(_1162_));
 sg13g2_inv_1 _6062_ (.Y(_1163_),
    .A(_1162_));
 sg13g2_nand2_1 _6063_ (.Y(_1164_),
    .A(_1161_),
    .B(_1149_));
 sg13g2_nand2_1 _6064_ (.Y(_1165_),
    .A(_1163_),
    .B(_1164_));
 sg13g2_o21ai_1 _6065_ (.B1(_1076_),
    .Y(_1166_),
    .A1(_1075_),
    .A2(_1122_));
 sg13g2_o21ai_1 _6066_ (.B1(_4325_),
    .Y(_1167_),
    .A1(_1165_),
    .A2(_1166_));
 sg13g2_a21oi_1 _6067_ (.A1(_1165_),
    .A2(_1166_),
    .Y(_1168_),
    .B1(_1167_));
 sg13g2_a21o_1 _6068_ (.A2(_1148_),
    .A1(net51),
    .B1(_1168_),
    .X(\generated._1069[4] ));
 sg13g2_inv_1 _6069_ (.Y(_1169_),
    .A(_0025_));
 sg13g2_nand2_1 _6070_ (.Y(_1170_),
    .A(_1152_),
    .B(_1169_));
 sg13g2_nand2_1 _6071_ (.Y(_1171_),
    .A(_1156_),
    .B(_1028_));
 sg13g2_o21ai_1 _6072_ (.B1(_1171_),
    .Y(_1172_),
    .A1(_1155_),
    .A2(_1170_));
 sg13g2_xnor2_1 _6073_ (.Y(_1173_),
    .A(_1033_),
    .B(_1172_));
 sg13g2_nor2b_1 _6074_ (.A(_1159_),
    .B_N(_1157_),
    .Y(_1174_));
 sg13g2_nor2b_1 _6075_ (.A(_1150_),
    .B_N(_1160_),
    .Y(_1175_));
 sg13g2_nor2_1 _6076_ (.A(_1174_),
    .B(_1175_),
    .Y(_1176_));
 sg13g2_xor2_1 _6077_ (.B(_1176_),
    .A(_1173_),
    .X(_1177_));
 sg13g2_nor2b_1 _6078_ (.A(_1162_),
    .B_N(_1166_),
    .Y(_1178_));
 sg13g2_nor2b_1 _6079_ (.A(_1178_),
    .B_N(_1164_),
    .Y(_1179_));
 sg13g2_inv_1 _6080_ (.Y(_1180_),
    .A(_1179_));
 sg13g2_nor2_1 _6081_ (.A(_1177_),
    .B(_1180_),
    .Y(_1181_));
 sg13g2_inv_1 _6082_ (.Y(_1182_),
    .A(_1181_));
 sg13g2_nand2_1 _6083_ (.Y(_1183_),
    .A(_1180_),
    .B(_1177_));
 sg13g2_nand3_1 _6084_ (.B(net48),
    .C(_1183_),
    .A(_1182_),
    .Y(_1184_));
 sg13g2_nand2_1 _6085_ (.Y(_1185_),
    .A(net77),
    .B(_0027_));
 sg13g2_o21ai_1 _6086_ (.B1(_1185_),
    .Y(_1186_),
    .A1(net64),
    .A2(_1010_));
 sg13g2_nor2_1 _6087_ (.A(net93),
    .B(_1127_),
    .Y(_1187_));
 sg13g2_a21oi_1 _6088_ (.A1(net89),
    .A2(_1186_),
    .Y(_1188_),
    .B1(_1187_));
 sg13g2_inv_1 _6089_ (.Y(_1189_),
    .A(_1141_));
 sg13g2_nor2_1 _6090_ (.A(_1139_),
    .B(_1189_),
    .Y(_1190_));
 sg13g2_nor2_1 _6091_ (.A(net46),
    .B(_1190_),
    .Y(_1191_));
 sg13g2_xnor2_1 _6092_ (.Y(_1192_),
    .A(_1188_),
    .B(_1191_));
 sg13g2_xnor2_1 _6093_ (.Y(_1193_),
    .A(_0026_),
    .B(_1192_));
 sg13g2_inv_1 _6094_ (.Y(_1194_),
    .A(_1193_));
 sg13g2_a22oi_1 _6095_ (.Y(_1195_),
    .B1(_1144_),
    .B2(_1147_),
    .A2(_1143_),
    .A1(\generated._1070[4] ));
 sg13g2_nor2_1 _6096_ (.A(_1194_),
    .B(_1195_),
    .Y(_1196_));
 sg13g2_inv_1 _6097_ (.Y(_1197_),
    .A(_1196_));
 sg13g2_nand2_1 _6098_ (.Y(_1198_),
    .A(_1195_),
    .B(_1194_));
 sg13g2_nand3_1 _6099_ (.B(net65),
    .C(_1198_),
    .A(_1197_),
    .Y(_1199_));
 sg13g2_nand2_1 _6100_ (.Y(\generated._1069[5] ),
    .A(_1184_),
    .B(_1199_));
 sg13g2_nor2_1 _6101_ (.A(_1151_),
    .B(_1154_),
    .Y(_1200_));
 sg13g2_inv_1 _6102_ (.Y(_1201_),
    .A(_1200_));
 sg13g2_nand2_1 _6103_ (.Y(_1202_),
    .A(_1174_),
    .B(_1173_));
 sg13g2_nand2_1 _6104_ (.Y(_1203_),
    .A(_1172_),
    .B(_1032_));
 sg13g2_nand2_1 _6105_ (.Y(_1204_),
    .A(_1202_),
    .B(_1203_));
 sg13g2_xnor2_1 _6106_ (.Y(_1205_),
    .A(_1201_),
    .B(_1204_));
 sg13g2_inv_1 _6107_ (.Y(_1206_),
    .A(_1205_));
 sg13g2_a21o_1 _6108_ (.A2(_1173_),
    .A1(_1175_),
    .B1(_1181_),
    .X(_1207_));
 sg13g2_inv_1 _6109_ (.Y(_1208_),
    .A(_1207_));
 sg13g2_nor2_1 _6110_ (.A(_1206_),
    .B(_1208_),
    .Y(_1209_));
 sg13g2_o21ai_1 _6111_ (.B1(net48),
    .Y(_1210_),
    .A1(_1205_),
    .A2(_1207_));
 sg13g2_nor2b_1 _6112_ (.A(_4426_),
    .B_N(_0027_),
    .Y(_1211_));
 sg13g2_a21oi_1 _6113_ (.A1(_4426_),
    .A2(_0029_),
    .Y(_1212_),
    .B1(_1211_));
 sg13g2_nor2_1 _6114_ (.A(net78),
    .B(_1212_),
    .Y(_1213_));
 sg13g2_a21oi_2 _6115_ (.B1(_1213_),
    .Y(_1214_),
    .A2(_1137_),
    .A1(net78));
 sg13g2_inv_1 _6116_ (.Y(_1215_),
    .A(_1190_));
 sg13g2_nor2_1 _6117_ (.A(_1188_),
    .B(_1215_),
    .Y(_1216_));
 sg13g2_nor2_1 _6118_ (.A(net46),
    .B(_1216_),
    .Y(_1217_));
 sg13g2_xnor2_1 _6119_ (.Y(_1218_),
    .A(_1214_),
    .B(_1217_));
 sg13g2_xnor2_1 _6120_ (.Y(_1219_),
    .A(_0028_),
    .B(_1218_));
 sg13g2_inv_1 _6121_ (.Y(_1220_),
    .A(_1219_));
 sg13g2_a21o_1 _6122_ (.A2(_1192_),
    .A1(\generated._1070[5] ),
    .B1(_1196_),
    .X(_1221_));
 sg13g2_inv_1 _6123_ (.Y(_1222_),
    .A(_1221_));
 sg13g2_nor2_1 _6124_ (.A(_1220_),
    .B(_1222_),
    .Y(_1223_));
 sg13g2_a21oi_1 _6125_ (.A1(_1222_),
    .A2(_1220_),
    .Y(_1224_),
    .B1(_4325_));
 sg13g2_nand2b_1 _6126_ (.Y(_1225_),
    .B(_1224_),
    .A_N(_1223_));
 sg13g2_o21ai_1 _6127_ (.B1(_1225_),
    .Y(\generated._1069[6] ),
    .A1(_1209_),
    .A2(_1210_));
 sg13g2_nor2_1 _6128_ (.A(_1201_),
    .B(_1202_),
    .Y(_1226_));
 sg13g2_inv_1 _6129_ (.Y(_1227_),
    .A(_1067_));
 sg13g2_nand2_1 _6130_ (.Y(_1228_),
    .A(_1227_),
    .B(_1055_));
 sg13g2_o21ai_1 _6131_ (.B1(_1228_),
    .Y(_1229_),
    .A1(_1227_),
    .A2(_1056_));
 sg13g2_nor2_1 _6132_ (.A(_1201_),
    .B(_1203_),
    .Y(_1230_));
 sg13g2_xor2_1 _6133_ (.B(_1230_),
    .A(_1229_),
    .X(_1231_));
 sg13g2_nor3_1 _6134_ (.A(_1226_),
    .B(_1231_),
    .C(_1209_),
    .Y(_1232_));
 sg13g2_o21ai_1 _6135_ (.B1(_1231_),
    .Y(_1233_),
    .A1(_1226_),
    .A2(_1209_));
 sg13g2_nand2_1 _6136_ (.Y(_1234_),
    .A(_1233_),
    .B(net48));
 sg13g2_a21oi_1 _6137_ (.A1(\generated._1070[6] ),
    .A2(_1218_),
    .Y(_1235_),
    .B1(_1223_));
 sg13g2_nand2_1 _6138_ (.Y(_1236_),
    .A(_4445_),
    .B(_0029_));
 sg13g2_inv_1 _6139_ (.Y(_1237_),
    .A(_1236_));
 sg13g2_a21oi_1 _6140_ (.A1(_1186_),
    .A2(net78),
    .Y(_1238_),
    .B1(_1237_));
 sg13g2_inv_1 _6141_ (.Y(_1239_),
    .A(_1216_));
 sg13g2_o21ai_1 _6142_ (.B1(net47),
    .Y(_1240_),
    .A1(_1214_),
    .A2(_1239_));
 sg13g2_xor2_1 _6143_ (.B(_1240_),
    .A(_1238_),
    .X(_1241_));
 sg13g2_xnor2_1 _6144_ (.Y(_1242_),
    .A(_0030_),
    .B(_1241_));
 sg13g2_inv_1 _6145_ (.Y(_1243_),
    .A(_1242_));
 sg13g2_a21oi_1 _6146_ (.A1(_1235_),
    .A2(_1243_),
    .Y(_1244_),
    .B1(net48));
 sg13g2_nor2_1 _6147_ (.A(_1243_),
    .B(_1235_),
    .Y(_1245_));
 sg13g2_inv_1 _6148_ (.Y(_1246_),
    .A(_1245_));
 sg13g2_nand2_1 _6149_ (.Y(_1247_),
    .A(_1244_),
    .B(_1246_));
 sg13g2_o21ai_1 _6150_ (.B1(_1247_),
    .Y(\generated._1069[7] ),
    .A1(_1232_),
    .A2(_1234_));
 sg13g2_nand2_1 _6151_ (.Y(_1248_),
    .A(_1230_),
    .B(_1229_));
 sg13g2_o21ai_1 _6152_ (.B1(_1067_),
    .Y(_1249_),
    .A1(_1055_),
    .A2(_1044_));
 sg13g2_and3_1 _6153_ (.X(_1250_),
    .A(_1233_),
    .B(_1248_),
    .C(_1249_));
 sg13g2_o21ai_1 _6154_ (.B1(_1236_),
    .Y(_1251_),
    .A1(_4445_),
    .A2(_1212_));
 sg13g2_or3_1 _6155_ (.A(_1214_),
    .B(_1238_),
    .C(_1239_),
    .X(_1252_));
 sg13g2_nand2_1 _6156_ (.Y(_1253_),
    .A(_1252_),
    .B(net47));
 sg13g2_xor2_1 _6157_ (.B(_1253_),
    .A(_1251_),
    .X(_1254_));
 sg13g2_xnor2_1 _6158_ (.Y(_1255_),
    .A(_0031_),
    .B(_1254_));
 sg13g2_a21o_1 _6159_ (.A2(_1241_),
    .A1(\generated._1070[7] ),
    .B1(_1245_),
    .X(_1256_));
 sg13g2_inv_1 _6160_ (.Y(_1257_),
    .A(_1256_));
 sg13g2_nor2_1 _6161_ (.A(_1255_),
    .B(_1257_),
    .Y(_1258_));
 sg13g2_inv_1 _6162_ (.Y(_1259_),
    .A(_1258_));
 sg13g2_nand2_1 _6163_ (.Y(_1260_),
    .A(_1257_),
    .B(_1255_));
 sg13g2_nand3_1 _6164_ (.B(_4324_),
    .C(_1260_),
    .A(_1259_),
    .Y(_1261_));
 sg13g2_o21ai_1 _6165_ (.B1(_1261_),
    .Y(\generated._1069[8] ),
    .A1(net51),
    .A2(_1250_));
 sg13g2_buf_1 _6166_ (.A(_0032_),
    .X(_1262_));
 sg13g2_inv_1 _6167_ (.Y(_1263_),
    .A(\generated._1070[8] ));
 sg13g2_o21ai_1 _6168_ (.B1(_1259_),
    .Y(_1264_),
    .A1(_1263_),
    .A2(_1254_));
 sg13g2_nor2b_1 _6169_ (.A(_1252_),
    .B_N(_1251_),
    .Y(_1265_));
 sg13g2_xnor2_1 _6170_ (.Y(_1266_),
    .A(\generated._1020[9] ),
    .B(_1265_));
 sg13g2_nor2_1 _6171_ (.A(_0029_),
    .B(net47),
    .Y(_1267_));
 sg13g2_a21oi_1 _6172_ (.A1(_1266_),
    .A2(net47),
    .Y(_1268_),
    .B1(_1267_));
 sg13g2_xnor2_1 _6173_ (.Y(_1269_),
    .A(_4352_),
    .B(_1268_));
 sg13g2_nand2b_1 _6174_ (.Y(_1270_),
    .B(_1269_),
    .A_N(_1264_));
 sg13g2_nand2b_1 _6175_ (.Y(_1271_),
    .B(_1264_),
    .A_N(_1269_));
 sg13g2_nand3_1 _6176_ (.B(_4324_),
    .C(_1271_),
    .A(_1270_),
    .Y(_1272_));
 sg13g2_o21ai_1 _6177_ (.B1(_1272_),
    .Y(\generated._1069[9] ),
    .A1(_1262_),
    .A2(net51));
 sg13g2_nand3_1 _6178_ (.B(\generated._1074[2] ),
    .C(_4322_),
    .A(_4320_),
    .Y(_1273_));
 sg13g2_nor2b_1 _6179_ (.A(\generated._1074[0] ),
    .B_N(_1273_),
    .Y(\generated._1073[0] ));
 sg13g2_nand2_1 _6180_ (.Y(_1274_),
    .A(\generated._1074[1] ),
    .B(\generated._1074[0] ));
 sg13g2_inv_1 _6181_ (.Y(_1275_),
    .A(_1274_));
 sg13g2_nor2_1 _6182_ (.A(_4320_),
    .B(_1275_),
    .Y(\generated._1073[1] ));
 sg13g2_nand2_1 _6183_ (.Y(_1276_),
    .A(_1275_),
    .B(\generated._1074[2] ));
 sg13g2_nand2_1 _6184_ (.Y(_1277_),
    .A(_1274_),
    .B(_4321_));
 sg13g2_and3_1 _6185_ (.X(\generated._1073[2] ),
    .A(_1273_),
    .B(_1276_),
    .C(_1277_));
 sg13g2_xnor2_1 _6186_ (.Y(\generated._1073[3] ),
    .A(\generated._1074[3] ),
    .B(_1276_));
 sg13g2_nor3_1 _6187_ (.A(_4230_),
    .B(_4241_),
    .C(_4314_),
    .Y(_1278_));
 sg13g2_nand4_1 _6188_ (.B(_4231_),
    .C(_4234_),
    .A(_1278_),
    .Y(\generated._108 ),
    .D(_4232_));
 sg13g2_inv_1 _6189_ (.Y(\generated._1115[0] ),
    .A(\generated._568[0] ));
 sg13g2_nor2b_1 _6190_ (.A(_4168_),
    .B_N(_4261_),
    .Y(\generated._1115[1] ));
 sg13g2_xnor2_1 _6191_ (.Y(\generated._1115[2] ),
    .A(\generated._568[2] ),
    .B(_4261_));
 sg13g2_inv_1 _6192_ (.Y(_1279_),
    .A(_0120_));
 sg13g2_xnor2_1 _6193_ (.Y(_1280_),
    .A(_1279_),
    .B(_4262_));
 sg13g2_nand3_1 _6194_ (.B(_4159_),
    .C(\generated._568[9] ),
    .A(_4158_),
    .Y(_1281_));
 sg13g2_nand2_1 _6195_ (.Y(_1282_),
    .A(_4264_),
    .B(_4163_));
 sg13g2_nor2_1 _6196_ (.A(_1281_),
    .B(_1282_),
    .Y(_1283_));
 sg13g2_nor2_1 _6197_ (.A(_1280_),
    .B(_1283_),
    .Y(\generated._1115[3] ));
 sg13g2_xor2_1 _6198_ (.B(_4264_),
    .A(net95),
    .X(\generated._1115[4] ));
 sg13g2_buf_1 _6199_ (.A(_0121_),
    .X(_1284_));
 sg13g2_a21oi_1 _6200_ (.A1(_1281_),
    .A2(_1284_),
    .Y(_1285_),
    .B1(_1282_));
 sg13g2_a21oi_1 _6201_ (.A1(_1284_),
    .A2(_1282_),
    .Y(\generated._1115[5] ),
    .B1(_1285_));
 sg13g2_nand3_1 _6202_ (.B(_4155_),
    .C(_4157_),
    .A(net95),
    .Y(_1286_));
 sg13g2_nor3_2 _6203_ (.A(_4260_),
    .B(_1286_),
    .C(_4263_),
    .Y(_1287_));
 sg13g2_inv_1 _6204_ (.Y(_1288_),
    .A(_1287_));
 sg13g2_o21ai_1 _6205_ (.B1(_1288_),
    .Y(_1289_),
    .A1(_4155_),
    .A2(_4157_));
 sg13g2_a21oi_1 _6206_ (.A1(_4270_),
    .A2(_1282_),
    .Y(\generated._1115[6] ),
    .B1(_1289_));
 sg13g2_inv_1 _6207_ (.Y(_1290_),
    .A(_0117_));
 sg13g2_xnor2_1 _6208_ (.Y(_1291_),
    .A(_1290_),
    .B(_1287_));
 sg13g2_nor2_1 _6209_ (.A(_1283_),
    .B(_1291_),
    .Y(\generated._1115[7] ));
 sg13g2_a21oi_1 _6210_ (.A1(_1287_),
    .A2(_4156_),
    .Y(_1292_),
    .B1(_4159_));
 sg13g2_nor3_1 _6211_ (.A(_4265_),
    .B(_4160_),
    .C(_1288_),
    .Y(_1293_));
 sg13g2_nor3_1 _6212_ (.A(_1283_),
    .B(_1292_),
    .C(_1293_),
    .Y(\generated._1115[8] ));
 sg13g2_inv_1 _6213_ (.Y(_1294_),
    .A(_0122_));
 sg13g2_xnor2_1 _6214_ (.Y(_1295_),
    .A(_1294_),
    .B(_1293_));
 sg13g2_nor2_1 _6215_ (.A(_1283_),
    .B(_1295_),
    .Y(\generated._1115[9] ));
 sg13g2_o21ai_1 _6216_ (.B1(\generated._568[9] ),
    .Y(_1296_),
    .A1(_4159_),
    .A2(_1290_));
 sg13g2_inv_1 _6217_ (.Y(_1297_),
    .A(_1296_));
 sg13g2_nor3_2 _6218_ (.A(_4230_),
    .B(_1297_),
    .C(_4315_),
    .Y(_1298_));
 sg13g2_inv_1 _6219_ (.Y(_1299_),
    .A(_1298_));
 sg13g2_nor2_1 _6220_ (.A(\generated._217[2] ),
    .B(_4230_),
    .Y(_1300_));
 sg13g2_inv_1 _6221_ (.Y(_1301_),
    .A(_1300_));
 sg13g2_nand2_1 _6222_ (.Y(_1302_),
    .A(_4237_),
    .B(_4241_));
 sg13g2_nor2_1 _6223_ (.A(_1302_),
    .B(_4312_),
    .Y(_1303_));
 sg13g2_nor2_2 _6224_ (.A(_1301_),
    .B(_1303_),
    .Y(_1304_));
 sg13g2_nor2_1 _6225_ (.A(_4193_),
    .B(_0008_),
    .Y(_1305_));
 sg13g2_inv_1 _6226_ (.Y(_1306_),
    .A(_1304_));
 sg13g2_nor3_1 _6227_ (.A(\generated._26[1] ),
    .B(_4520_),
    .C(net39),
    .Y(_1307_));
 sg13g2_a21oi_1 _6228_ (.A1(_4289_),
    .A2(_4241_),
    .Y(_1308_),
    .B1(_4237_));
 sg13g2_o21ai_1 _6229_ (.B1(_1308_),
    .Y(_1309_),
    .A1(_4296_),
    .A2(_4235_));
 sg13g2_o21ai_1 _6230_ (.B1(_4311_),
    .Y(_1310_),
    .A1(_4231_),
    .A2(_4243_));
 sg13g2_a21oi_1 _6231_ (.A1(_4313_),
    .A2(_1309_),
    .Y(_1311_),
    .B1(_1310_));
 sg13g2_nand2_1 _6232_ (.Y(_1312_),
    .A(_4265_),
    .B(_4157_));
 sg13g2_nand3_1 _6233_ (.B(net95),
    .C(_4155_),
    .A(_4162_),
    .Y(_1313_));
 sg13g2_nor3_1 _6234_ (.A(_1312_),
    .B(_4267_),
    .C(_1313_),
    .Y(_1314_));
 sg13g2_nor3_1 _6235_ (.A(_1297_),
    .B(_1314_),
    .C(_4166_),
    .Y(_1315_));
 sg13g2_nand2_1 _6236_ (.Y(_1316_),
    .A(_1311_),
    .B(_1315_));
 sg13g2_buf_2 _6237_ (.A(_1316_),
    .X(_1317_));
 sg13g2_nor2_1 _6238_ (.A(_1307_),
    .B(_1317_),
    .Y(_1318_));
 sg13g2_o21ai_1 _6239_ (.B1(_1318_),
    .Y(_1319_),
    .A1(_1304_),
    .A2(_1305_));
 sg13g2_buf_2 _6240_ (.A(uio_in[0]),
    .X(_1320_));
 sg13g2_inv_1 _6241_ (.Y(_1321_),
    .A(_1320_));
 sg13g2_inv_1 _6242_ (.Y(_1322_),
    .A(_1317_));
 sg13g2_mux2_1 _6243_ (.A0(\generated._1144[0] ),
    .A1(_0118_),
    .S(_1311_),
    .X(_1323_));
 sg13g2_nor2_1 _6244_ (.A(_1322_),
    .B(_1323_),
    .Y(_1324_));
 sg13g2_nor2_1 _6245_ (.A(_1321_),
    .B(_1324_),
    .Y(_1325_));
 sg13g2_buf_1 _6246_ (.A(\generated._63[3] ),
    .X(_1326_));
 sg13g2_buf_2 _6247_ (.A(\generated._63[2] ),
    .X(_1327_));
 sg13g2_buf_2 _6248_ (.A(\generated._161[4] ),
    .X(_1328_));
 sg13g2_nand2_1 _6249_ (.Y(_1329_),
    .A(_1327_),
    .B(_1328_));
 sg13g2_nor2_1 _6250_ (.A(_1326_),
    .B(_1329_),
    .Y(_1330_));
 sg13g2_inv_1 _6251_ (.Y(_1331_),
    .A(_1330_));
 sg13g2_buf_2 _6252_ (.A(\generated._63[4] ),
    .X(_1332_));
 sg13g2_buf_2 _6253_ (.A(\generated._1083[0] ),
    .X(_1333_));
 sg13g2_xor2_1 _6254_ (.B(_1333_),
    .A(_1332_),
    .X(_1334_));
 sg13g2_inv_1 _6255_ (.Y(_1335_),
    .A(_1334_));
 sg13g2_nor2_1 _6256_ (.A(_1331_),
    .B(_1335_),
    .Y(_1336_));
 sg13g2_nand3_1 _6257_ (.B(_1326_),
    .C(_1327_),
    .A(_1335_),
    .Y(_1337_));
 sg13g2_nor2b_1 _6258_ (.A(_1336_),
    .B_N(_1337_),
    .Y(_1338_));
 sg13g2_inv_1 _6259_ (.Y(_1339_),
    .A(_1332_));
 sg13g2_inv_1 _6260_ (.Y(_1340_),
    .A(_1333_));
 sg13g2_inv_1 _6261_ (.Y(_1341_),
    .A(_1326_));
 sg13g2_nor2_1 _6262_ (.A(_1341_),
    .B(_1335_),
    .Y(_1342_));
 sg13g2_inv_1 _6263_ (.Y(_1343_),
    .A(\generated._63[5] ));
 sg13g2_nand2b_1 _6264_ (.Y(_1344_),
    .B(_1343_),
    .A_N(_1328_));
 sg13g2_nand2_1 _6265_ (.Y(_1345_),
    .A(_1328_),
    .B(\generated._63[5] ));
 sg13g2_nand2_1 _6266_ (.Y(_1346_),
    .A(_1344_),
    .B(_1345_));
 sg13g2_xnor2_1 _6267_ (.Y(_1347_),
    .A(_1333_),
    .B(_1346_));
 sg13g2_xnor2_1 _6268_ (.Y(_1348_),
    .A(_1339_),
    .B(_1347_));
 sg13g2_xnor2_1 _6269_ (.Y(_1349_),
    .A(_1342_),
    .B(_1348_));
 sg13g2_o21ai_1 _6270_ (.B1(_1349_),
    .Y(_1350_),
    .A1(_1339_),
    .A2(_1340_));
 sg13g2_nand4_1 _6271_ (.B(_1345_),
    .C(_1332_),
    .A(_1344_),
    .Y(_1351_),
    .D(_1333_));
 sg13g2_nand2_1 _6272_ (.Y(_1352_),
    .A(_1350_),
    .B(_1351_));
 sg13g2_xnor2_1 _6273_ (.Y(_1353_),
    .A(_1338_),
    .B(_1352_));
 sg13g2_nand2_1 _6274_ (.Y(_1354_),
    .A(_1326_),
    .B(_1328_));
 sg13g2_nor3_1 _6275_ (.A(_1340_),
    .B(_1327_),
    .C(_1354_),
    .Y(_1355_));
 sg13g2_inv_1 _6276_ (.Y(_1356_),
    .A(_1355_));
 sg13g2_inv_1 _6277_ (.Y(_1357_),
    .A(_1327_));
 sg13g2_a21oi_1 _6278_ (.A1(_1326_),
    .A2(_1357_),
    .Y(_1358_),
    .B1(_1330_));
 sg13g2_xnor2_1 _6279_ (.Y(_1359_),
    .A(_1334_),
    .B(_1358_));
 sg13g2_inv_1 _6280_ (.Y(_1360_),
    .A(_1359_));
 sg13g2_nor2_1 _6281_ (.A(_1356_),
    .B(_1360_),
    .Y(_1361_));
 sg13g2_nor2_1 _6282_ (.A(_1326_),
    .B(_1328_),
    .Y(_1362_));
 sg13g2_inv_1 _6283_ (.Y(_1363_),
    .A(_1362_));
 sg13g2_nor2_1 _6284_ (.A(_1333_),
    .B(_1327_),
    .Y(_1364_));
 sg13g2_inv_1 _6285_ (.Y(_1365_),
    .A(_1354_));
 sg13g2_nor2_1 _6286_ (.A(_1362_),
    .B(_1365_),
    .Y(_1366_));
 sg13g2_a21oi_1 _6287_ (.A1(_1341_),
    .A2(_1328_),
    .Y(_1367_),
    .B1(_1357_));
 sg13g2_a221oi_1 _6288_ (.B2(_1333_),
    .C1(_1367_),
    .B1(_1366_),
    .A1(_1363_),
    .Y(_1368_),
    .A2(_1364_));
 sg13g2_xnor2_1 _6289_ (.Y(_1369_),
    .A(_1356_),
    .B(_1359_));
 sg13g2_inv_1 _6290_ (.Y(_1370_),
    .A(_1369_));
 sg13g2_nor2_1 _6291_ (.A(_1368_),
    .B(_1370_),
    .Y(_1371_));
 sg13g2_nor2_1 _6292_ (.A(_1361_),
    .B(_1371_),
    .Y(_1372_));
 sg13g2_a21oi_1 _6293_ (.A1(_1353_),
    .A2(_1372_),
    .Y(_1373_),
    .B1(_1320_));
 sg13g2_inv_1 _6294_ (.Y(_1374_),
    .A(_1361_));
 sg13g2_inv_1 _6295_ (.Y(_1375_),
    .A(_1371_));
 sg13g2_a21o_1 _6296_ (.A2(_1375_),
    .A1(_1374_),
    .B1(_1353_),
    .X(_1376_));
 sg13g2_a22oi_1 _6297_ (.Y(_1377_),
    .B1(_1373_),
    .B2(_1376_),
    .A2(_1325_),
    .A1(_1319_));
 sg13g2_o21ai_1 _6298_ (.B1(net39),
    .Y(_1378_),
    .A1(_4193_),
    .A2(_0007_));
 sg13g2_inv_1 _6299_ (.Y(_1379_),
    .A(_1325_));
 sg13g2_a21o_1 _6300_ (.A2(_1378_),
    .A1(_1318_),
    .B1(_1379_),
    .X(_1380_));
 sg13g2_nand2_1 _6301_ (.Y(_1381_),
    .A(_1370_),
    .B(_1368_));
 sg13g2_nand3_1 _6302_ (.B(_1321_),
    .C(_1381_),
    .A(_1375_),
    .Y(_1382_));
 sg13g2_and3_1 _6303_ (.X(_1383_),
    .A(_1377_),
    .B(_1380_),
    .C(_1382_));
 sg13g2_o21ai_1 _6304_ (.B1(_1306_),
    .Y(_1384_),
    .A1(_4193_),
    .A2(_0009_));
 sg13g2_a21oi_1 _6305_ (.A1(_1318_),
    .A2(_1384_),
    .Y(_1385_),
    .B1(_1379_));
 sg13g2_nor2_1 _6306_ (.A(_1375_),
    .B(_1353_),
    .Y(_1386_));
 sg13g2_nand2_1 _6307_ (.Y(_1387_),
    .A(_1348_),
    .B(_1342_));
 sg13g2_nand2_1 _6308_ (.Y(_1388_),
    .A(_1387_),
    .B(_1351_));
 sg13g2_nor2_1 _6309_ (.A(_1328_),
    .B(_1340_),
    .Y(_1389_));
 sg13g2_inv_1 _6310_ (.Y(_1390_),
    .A(_1345_));
 sg13g2_a22oi_1 _6311_ (.Y(_1391_),
    .B1(_1340_),
    .B2(_1390_),
    .A2(_1343_),
    .A1(_1389_));
 sg13g2_xnor2_1 _6312_ (.Y(_1392_),
    .A(_0119_),
    .B(_1391_));
 sg13g2_xnor2_1 _6313_ (.Y(_1393_),
    .A(\generated._63[5] ),
    .B(\generated._63[6] ));
 sg13g2_xnor2_1 _6314_ (.Y(_1394_),
    .A(_1357_),
    .B(_1393_));
 sg13g2_nand2_1 _6315_ (.Y(_1395_),
    .A(_1347_),
    .B(_1332_));
 sg13g2_xnor2_1 _6316_ (.Y(_1396_),
    .A(_1394_),
    .B(_1395_));
 sg13g2_xnor2_1 _6317_ (.Y(_1397_),
    .A(_1392_),
    .B(_1396_));
 sg13g2_xor2_1 _6318_ (.B(_1397_),
    .A(_1388_),
    .X(_1398_));
 sg13g2_nor2_1 _6319_ (.A(_1337_),
    .B(_1352_),
    .Y(_1399_));
 sg13g2_xnor2_1 _6320_ (.Y(_1400_),
    .A(_1398_),
    .B(_1399_));
 sg13g2_nand3_1 _6321_ (.B(_1351_),
    .C(_1336_),
    .A(_1350_),
    .Y(_1401_));
 sg13g2_o21ai_1 _6322_ (.B1(_1401_),
    .Y(_1402_),
    .A1(_1374_),
    .A2(_1353_));
 sg13g2_xnor2_1 _6323_ (.Y(_1403_),
    .A(_1400_),
    .B(_1402_));
 sg13g2_xor2_1 _6324_ (.B(_1403_),
    .A(_1386_),
    .X(_1404_));
 sg13g2_nor2_1 _6325_ (.A(_1320_),
    .B(_1404_),
    .Y(_1405_));
 sg13g2_nor3_1 _6326_ (.A(_1377_),
    .B(_1385_),
    .C(_1405_),
    .Y(_1406_));
 sg13g2_nor3_1 _6327_ (.A(_1299_),
    .B(_1383_),
    .C(_1406_),
    .Y(\generated._1149[0] ));
 sg13g2_nor2_1 _6328_ (.A(_1385_),
    .B(_1405_),
    .Y(_1407_));
 sg13g2_a21oi_1 _6329_ (.A1(_1407_),
    .A2(_1377_),
    .Y(\generated._1149[1] ),
    .B1(_1299_));
 sg13g2_nand3_1 _6330_ (.B(_4271_),
    .C(_1286_),
    .A(_4268_),
    .Y(\generated._118 ));
 sg13g2_o21ai_1 _6331_ (.B1(_1304_),
    .Y(_1408_),
    .A1(_4509_),
    .A2(_4520_));
 sg13g2_nand3b_1 _6332_ (.B(net39),
    .C(net91),
    .Y(_1409_),
    .A_N(_0014_));
 sg13g2_a21oi_1 _6333_ (.A1(_1408_),
    .A2(_1409_),
    .Y(_1410_),
    .B1(_1317_));
 sg13g2_inv_1 _6334_ (.Y(_1411_),
    .A(_1324_));
 sg13g2_nand2b_1 _6335_ (.Y(_1412_),
    .B(_1411_),
    .A_N(_1410_));
 sg13g2_inv_1 _6336_ (.Y(_1413_),
    .A(_1389_));
 sg13g2_nand2_1 _6337_ (.Y(_1414_),
    .A(_1333_),
    .B(_1327_));
 sg13g2_inv_1 _6338_ (.Y(_1415_),
    .A(_1414_));
 sg13g2_nor2_1 _6339_ (.A(_1364_),
    .B(_1415_),
    .Y(_1416_));
 sg13g2_inv_1 _6340_ (.Y(_1417_),
    .A(_1416_));
 sg13g2_a21oi_1 _6341_ (.A1(_0119_),
    .A2(_1413_),
    .Y(_1418_),
    .B1(_1417_));
 sg13g2_xnor2_1 _6342_ (.Y(_1419_),
    .A(_1414_),
    .B(_1366_));
 sg13g2_xor2_1 _6343_ (.B(_1419_),
    .A(_1418_),
    .X(_1420_));
 sg13g2_nor2_1 _6344_ (.A(_1320_),
    .B(_1420_),
    .Y(_1421_));
 sg13g2_a21oi_1 _6345_ (.A1(_1412_),
    .A2(_1320_),
    .Y(_1422_),
    .B1(_1421_));
 sg13g2_nand3b_1 _6346_ (.B(net39),
    .C(net91),
    .Y(_1423_),
    .A_N(_0015_));
 sg13g2_a21oi_1 _6347_ (.A1(_1408_),
    .A2(_1423_),
    .Y(_1424_),
    .B1(_1317_));
 sg13g2_o21ai_1 _6348_ (.B1(_1320_),
    .Y(_1425_),
    .A1(_1424_),
    .A2(_1324_));
 sg13g2_xor2_1 _6349_ (.B(_1327_),
    .A(_1332_),
    .X(_1426_));
 sg13g2_a21oi_1 _6350_ (.A1(_1354_),
    .A2(_1414_),
    .Y(_1427_),
    .B1(_1362_));
 sg13g2_xnor2_1 _6351_ (.Y(_1428_),
    .A(_1426_),
    .B(_1427_));
 sg13g2_nor2_1 _6352_ (.A(_1333_),
    .B(_1328_),
    .Y(_1429_));
 sg13g2_nor2_1 _6353_ (.A(_1429_),
    .B(_1417_),
    .Y(_1430_));
 sg13g2_nand2_1 _6354_ (.Y(_1431_),
    .A(_1419_),
    .B(_1430_));
 sg13g2_xnor2_1 _6355_ (.Y(_1432_),
    .A(_1428_),
    .B(_1431_));
 sg13g2_nand2_1 _6356_ (.Y(_1433_),
    .A(_1432_),
    .B(_1321_));
 sg13g2_nand2_1 _6357_ (.Y(_1434_),
    .A(_1425_),
    .B(_1433_));
 sg13g2_inv_1 _6358_ (.Y(_1435_),
    .A(_1422_));
 sg13g2_nand3b_1 _6359_ (.B(net39),
    .C(net91),
    .Y(_1436_),
    .A_N(_0013_));
 sg13g2_a21oi_1 _6360_ (.A1(_1408_),
    .A2(_1436_),
    .Y(_1437_),
    .B1(_1317_));
 sg13g2_nand2b_1 _6361_ (.Y(_1438_),
    .B(_1325_),
    .A_N(_1437_));
 sg13g2_a21oi_1 _6362_ (.A1(_1357_),
    .A2(_1429_),
    .Y(_1439_),
    .B1(_1430_));
 sg13g2_nand2_1 _6363_ (.Y(_1440_),
    .A(_1439_),
    .B(_1321_));
 sg13g2_nand3_1 _6364_ (.B(_1438_),
    .C(_1440_),
    .A(_1435_),
    .Y(_1441_));
 sg13g2_nand2_1 _6365_ (.Y(_1442_),
    .A(_1441_),
    .B(_1298_));
 sg13g2_a21oi_1 _6366_ (.A1(_1422_),
    .A2(_1434_),
    .Y(\generated._231[0] ),
    .B1(_1442_));
 sg13g2_a21oi_1 _6367_ (.A1(_1435_),
    .A2(_1434_),
    .Y(\generated._231[1] ),
    .B1(_1299_));
 sg13g2_o21ai_1 _6368_ (.B1(_1304_),
    .Y(_1443_),
    .A1(_4520_),
    .A2(_4522_));
 sg13g2_nand3b_1 _6369_ (.B(net39),
    .C(net91),
    .Y(_1444_),
    .A_N(_0012_));
 sg13g2_a21oi_1 _6370_ (.A1(_1443_),
    .A2(_1444_),
    .Y(_1445_),
    .B1(_1317_));
 sg13g2_o21ai_1 _6371_ (.B1(_1320_),
    .Y(_1446_),
    .A1(_1445_),
    .A2(_1324_));
 sg13g2_nand2_1 _6372_ (.Y(_1447_),
    .A(_1446_),
    .B(_1433_));
 sg13g2_nand3b_1 _6373_ (.B(net39),
    .C(net91),
    .Y(_1448_),
    .A_N(_0011_));
 sg13g2_a21oi_1 _6374_ (.A1(_1443_),
    .A2(_1448_),
    .Y(_1449_),
    .B1(_1317_));
 sg13g2_nand2b_1 _6375_ (.Y(_1450_),
    .B(_1411_),
    .A_N(_1449_));
 sg13g2_a21oi_1 _6376_ (.A1(_1450_),
    .A2(_1320_),
    .Y(_1451_),
    .B1(_1421_));
 sg13g2_nand3b_1 _6377_ (.B(net39),
    .C(_4194_),
    .Y(_1452_),
    .A_N(_0010_));
 sg13g2_a21oi_1 _6378_ (.A1(_1443_),
    .A2(_1452_),
    .Y(_1453_),
    .B1(_1317_));
 sg13g2_o21ai_1 _6379_ (.B1(_1440_),
    .Y(_1454_),
    .A1(_1453_),
    .A2(_1379_));
 sg13g2_o21ai_1 _6380_ (.B1(_1298_),
    .Y(_1455_),
    .A1(_1451_),
    .A2(_1454_));
 sg13g2_a21oi_1 _6381_ (.A1(_1447_),
    .A2(_1451_),
    .Y(\generated._284[0] ),
    .B1(_1455_));
 sg13g2_inv_1 _6382_ (.Y(_1456_),
    .A(_1451_));
 sg13g2_a21oi_1 _6383_ (.A1(_1456_),
    .A2(_1447_),
    .Y(\generated._284[1] ),
    .B1(_1299_));
 sg13g2_nand2_1 _6384_ (.Y(_1457_),
    .A(_0911_),
    .B(_0089_));
 sg13g2_inv_1 _6385_ (.Y(_1458_),
    .A(_1457_));
 sg13g2_nor2_1 _6386_ (.A(_0089_),
    .B(_0911_),
    .Y(_1459_));
 sg13g2_nor3_1 _6387_ (.A(_1458_),
    .B(_1459_),
    .C(net62),
    .Y(_1460_));
 sg13g2_a21oi_1 _6388_ (.A1(_4414_),
    .A2(net44),
    .Y(\generated._477[0] ),
    .B1(_1460_));
 sg13g2_inv_1 _6389_ (.Y(_1461_),
    .A(\generated._369[1] ));
 sg13g2_xnor2_1 _6390_ (.Y(_1462_),
    .A(_0343_),
    .B(_0285_));
 sg13g2_inv_1 _6391_ (.Y(_1463_),
    .A(_1462_));
 sg13g2_nand2_1 _6392_ (.Y(_1464_),
    .A(_1463_),
    .B(_0911_));
 sg13g2_xnor2_1 _6393_ (.Y(_1465_),
    .A(_1461_),
    .B(_1464_));
 sg13g2_inv_1 _6394_ (.Y(_1466_),
    .A(_1465_));
 sg13g2_nor2_1 _6395_ (.A(_1458_),
    .B(_1466_),
    .Y(_1467_));
 sg13g2_o21ai_1 _6396_ (.B1(net33),
    .Y(_1468_),
    .A1(_1457_),
    .A2(_1465_));
 sg13g2_xnor2_1 _6397_ (.Y(_1469_),
    .A(net63),
    .B(_4417_));
 sg13g2_xnor2_1 _6398_ (.Y(_1470_),
    .A(_4414_),
    .B(_1469_));
 sg13g2_nand2b_1 _6399_ (.Y(_1471_),
    .B(net44),
    .A_N(_1470_));
 sg13g2_o21ai_1 _6400_ (.B1(_1471_),
    .Y(\generated._477[1] ),
    .A1(_1467_),
    .A2(_1468_));
 sg13g2_xnor2_1 _6401_ (.Y(_1472_),
    .A(net63),
    .B(_4425_));
 sg13g2_inv_1 _6402_ (.Y(_1473_),
    .A(_1472_));
 sg13g2_nand2_1 _6403_ (.Y(_1474_),
    .A(_1469_),
    .B(\generated._1080[0] ));
 sg13g2_o21ai_1 _6404_ (.B1(_1474_),
    .Y(_1475_),
    .A1(net45),
    .A2(_4433_));
 sg13g2_inv_1 _6405_ (.Y(_1476_),
    .A(_1475_));
 sg13g2_nor2_1 _6406_ (.A(_1473_),
    .B(_1476_),
    .Y(_1477_));
 sg13g2_o21ai_1 _6407_ (.B1(net62),
    .Y(_1478_),
    .A1(_1472_),
    .A2(_1475_));
 sg13g2_inv_1 _6408_ (.Y(_1479_),
    .A(_1464_));
 sg13g2_nor2_1 _6409_ (.A(_1461_),
    .B(_1479_),
    .Y(_1480_));
 sg13g2_nor2_1 _6410_ (.A(_1480_),
    .B(_1467_),
    .Y(_1481_));
 sg13g2_inv_1 _6411_ (.Y(_1482_),
    .A(_1481_));
 sg13g2_inv_1 _6412_ (.Y(_1483_),
    .A(\generated._369[2] ));
 sg13g2_nor2_1 _6413_ (.A(net73),
    .B(_0288_),
    .Y(_1484_));
 sg13g2_a21oi_1 _6414_ (.A1(net60),
    .A2(net73),
    .Y(_1485_),
    .B1(_1484_));
 sg13g2_nor2_1 _6415_ (.A(_1483_),
    .B(_1485_),
    .Y(_1486_));
 sg13g2_nand2_1 _6416_ (.Y(_1487_),
    .A(_1485_),
    .B(_1483_));
 sg13g2_nor2b_1 _6417_ (.A(_1486_),
    .B_N(_1487_),
    .Y(_1488_));
 sg13g2_nand2_1 _6418_ (.Y(_1489_),
    .A(_1482_),
    .B(_1488_));
 sg13g2_nand2b_1 _6419_ (.Y(_1490_),
    .B(_1481_),
    .A_N(_1488_));
 sg13g2_nand3_1 _6420_ (.B(net33),
    .C(_1490_),
    .A(_1489_),
    .Y(_1491_));
 sg13g2_o21ai_1 _6421_ (.B1(_1491_),
    .Y(\generated._477[2] ),
    .A1(_1477_),
    .A2(_1478_));
 sg13g2_inv_2 _6422_ (.Y(_1492_),
    .A(_4488_));
 sg13g2_buf_1 _6423_ (.A(_1492_),
    .X(_1493_));
 sg13g2_o21ai_1 _6424_ (.B1(net68),
    .Y(_1494_),
    .A1(_4417_),
    .A2(_4425_));
 sg13g2_o21ai_1 _6425_ (.B1(_1494_),
    .Y(_1495_),
    .A1(_1473_),
    .A2(_1474_));
 sg13g2_xor2_1 _6426_ (.B(_4437_),
    .A(net63),
    .X(_1496_));
 sg13g2_nand2_1 _6427_ (.Y(_1497_),
    .A(_1495_),
    .B(_1496_));
 sg13g2_inv_1 _6428_ (.Y(_1498_),
    .A(_1497_));
 sg13g2_o21ai_1 _6429_ (.B1(net62),
    .Y(_1499_),
    .A1(_1496_),
    .A2(_1495_));
 sg13g2_a21oi_1 _6430_ (.A1(_1482_),
    .A2(_1487_),
    .Y(_1500_),
    .B1(_1486_));
 sg13g2_inv_1 _6431_ (.Y(_1501_),
    .A(_1500_));
 sg13g2_nor2_1 _6432_ (.A(\generated._369[3] ),
    .B(_1464_),
    .Y(_1502_));
 sg13g2_nor2b_1 _6433_ (.A(_1479_),
    .B_N(\generated._369[3] ),
    .Y(_1503_));
 sg13g2_nor2_1 _6434_ (.A(_1502_),
    .B(_1503_),
    .Y(_1504_));
 sg13g2_a21oi_1 _6435_ (.A1(_1501_),
    .A2(_1504_),
    .Y(_1505_),
    .B1(net62));
 sg13g2_o21ai_1 _6436_ (.B1(_1505_),
    .Y(_1506_),
    .A1(_1501_),
    .A2(_1504_));
 sg13g2_o21ai_1 _6437_ (.B1(_1506_),
    .Y(\generated._477[3] ),
    .A1(_1498_),
    .A2(_1499_));
 sg13g2_o21ai_1 _6438_ (.B1(_4437_),
    .Y(_1507_),
    .A1(net45),
    .A2(_4425_));
 sg13g2_inv_1 _6439_ (.Y(_1508_),
    .A(_1507_));
 sg13g2_a21oi_1 _6440_ (.A1(_1477_),
    .A2(_1496_),
    .Y(_1509_),
    .B1(_1508_));
 sg13g2_xnor2_1 _6441_ (.Y(_1510_),
    .A(net63),
    .B(_4443_));
 sg13g2_nand2b_1 _6442_ (.Y(_1511_),
    .B(_1510_),
    .A_N(_1509_));
 sg13g2_inv_1 _6443_ (.Y(_1512_),
    .A(_1510_));
 sg13g2_a21oi_1 _6444_ (.A1(_1509_),
    .A2(_1512_),
    .Y(_1513_),
    .B1(net33));
 sg13g2_nor2_1 _6445_ (.A(net85),
    .B(_0285_),
    .Y(_1514_));
 sg13g2_a21oi_1 _6446_ (.A1(_0912_),
    .A2(net85),
    .Y(_1515_),
    .B1(_1514_));
 sg13g2_nor2_1 _6447_ (.A(\generated._369[4] ),
    .B(_1515_),
    .Y(_1516_));
 sg13g2_and2_1 _6448_ (.A(_1515_),
    .B(\generated._369[4] ),
    .X(_1517_));
 sg13g2_buf_1 _6449_ (.A(_1517_),
    .X(_1518_));
 sg13g2_nor2_1 _6450_ (.A(_1516_),
    .B(_1518_),
    .Y(_1519_));
 sg13g2_inv_1 _6451_ (.Y(_1520_),
    .A(_1502_));
 sg13g2_a21oi_1 _6452_ (.A1(_1501_),
    .A2(_1520_),
    .Y(_1521_),
    .B1(_1503_));
 sg13g2_inv_1 _6453_ (.Y(_1522_),
    .A(_1521_));
 sg13g2_o21ai_1 _6454_ (.B1(_0318_),
    .Y(_1523_),
    .A1(_1519_),
    .A2(_1522_));
 sg13g2_nand2_1 _6455_ (.Y(_1524_),
    .A(_1522_),
    .B(_1519_));
 sg13g2_nor2b_1 _6456_ (.A(_1523_),
    .B_N(_1524_),
    .Y(_1525_));
 sg13g2_a21o_1 _6457_ (.A2(_1513_),
    .A1(_1511_),
    .B1(_1525_),
    .X(\generated._477[4] ));
 sg13g2_inv_1 _6458_ (.Y(_1526_),
    .A(\generated._369[5] ));
 sg13g2_xnor2_1 _6459_ (.Y(_1527_),
    .A(net74),
    .B(net85));
 sg13g2_xnor2_1 _6460_ (.Y(_1528_),
    .A(_1526_),
    .B(_1527_));
 sg13g2_inv_1 _6461_ (.Y(_1529_),
    .A(_1516_));
 sg13g2_a21oi_1 _6462_ (.A1(_1522_),
    .A2(_1529_),
    .Y(_1530_),
    .B1(_1518_));
 sg13g2_nor2_1 _6463_ (.A(_1528_),
    .B(_1530_),
    .Y(_1531_));
 sg13g2_a21o_1 _6464_ (.A2(_1528_),
    .A1(_1530_),
    .B1(_0305_),
    .X(_1532_));
 sg13g2_o21ai_1 _6465_ (.B1(_4443_),
    .Y(_1533_),
    .A1(_4437_),
    .A2(net68));
 sg13g2_o21ai_1 _6466_ (.B1(_1533_),
    .Y(_1534_),
    .A1(_1512_),
    .A2(_1497_));
 sg13g2_xnor2_1 _6467_ (.Y(_1535_),
    .A(net45),
    .B(_4456_));
 sg13g2_inv_1 _6468_ (.Y(_1536_),
    .A(_1535_));
 sg13g2_inv_1 _6469_ (.Y(_1537_),
    .A(_1534_));
 sg13g2_nor2_1 _6470_ (.A(_1536_),
    .B(_1537_),
    .Y(_1538_));
 sg13g2_nor2_1 _6471_ (.A(_0318_),
    .B(_1538_),
    .Y(_1539_));
 sg13g2_o21ai_1 _6472_ (.B1(_1539_),
    .Y(_1540_),
    .A1(_1534_),
    .A2(_1535_));
 sg13g2_o21ai_1 _6473_ (.B1(_1540_),
    .Y(\generated._477[5] ),
    .A1(_1531_),
    .A2(_1532_));
 sg13g2_inv_1 _6474_ (.Y(_1541_),
    .A(\generated._369[6] ));
 sg13g2_nor2_1 _6475_ (.A(_1541_),
    .B(_1462_),
    .Y(_1542_));
 sg13g2_nor2_1 _6476_ (.A(\generated._369[6] ),
    .B(_1463_),
    .Y(_1543_));
 sg13g2_nor2_1 _6477_ (.A(_1542_),
    .B(_1543_),
    .Y(_1544_));
 sg13g2_nor2_1 _6478_ (.A(_1526_),
    .B(_1527_),
    .Y(_1545_));
 sg13g2_nor2_1 _6479_ (.A(_1545_),
    .B(_1518_),
    .Y(_1546_));
 sg13g2_a22oi_1 _6480_ (.Y(_1547_),
    .B1(_1546_),
    .B2(_1524_),
    .A2(_1527_),
    .A1(_1526_));
 sg13g2_nor2_1 _6481_ (.A(_1544_),
    .B(_1547_),
    .Y(_1548_));
 sg13g2_nand2_1 _6482_ (.Y(_1549_),
    .A(_1547_),
    .B(_1544_));
 sg13g2_nand2_1 _6483_ (.Y(_1550_),
    .A(_1549_),
    .B(net33));
 sg13g2_xor2_1 _6484_ (.B(_4466_),
    .A(net45),
    .X(_1551_));
 sg13g2_o21ai_1 _6485_ (.B1(net68),
    .Y(_1552_),
    .A1(_4443_),
    .A2(_4456_));
 sg13g2_a22oi_1 _6486_ (.Y(_1553_),
    .B1(_1552_),
    .B2(_1511_),
    .A2(_4457_),
    .A1(net45));
 sg13g2_a21oi_1 _6487_ (.A1(_1553_),
    .A2(_1551_),
    .Y(_1554_),
    .B1(_0318_));
 sg13g2_o21ai_1 _6488_ (.B1(_1554_),
    .Y(_1555_),
    .A1(_1551_),
    .A2(_1553_));
 sg13g2_o21ai_1 _6489_ (.B1(_1555_),
    .Y(\generated._477[6] ),
    .A1(_1548_),
    .A2(_1550_));
 sg13g2_nor2_1 _6490_ (.A(\generated._369[7] ),
    .B(net73),
    .Y(_1556_));
 sg13g2_nor2b_1 _6491_ (.A(net85),
    .B_N(\generated._369[7] ),
    .Y(_1557_));
 sg13g2_nor2_1 _6492_ (.A(_1556_),
    .B(_1557_),
    .Y(_1558_));
 sg13g2_nor2_1 _6493_ (.A(_1545_),
    .B(_1542_),
    .Y(_1559_));
 sg13g2_nor2_1 _6494_ (.A(_1543_),
    .B(_1559_),
    .Y(_1560_));
 sg13g2_a21oi_1 _6495_ (.A1(_1531_),
    .A2(_1544_),
    .Y(_1561_),
    .B1(_1560_));
 sg13g2_xor2_1 _6496_ (.B(_1561_),
    .A(_1558_),
    .X(_1562_));
 sg13g2_xor2_1 _6497_ (.B(_4473_),
    .A(net45),
    .X(_1563_));
 sg13g2_inv_1 _6498_ (.Y(_1564_),
    .A(_1563_));
 sg13g2_o21ai_1 _6499_ (.B1(_4466_),
    .Y(_1565_),
    .A1(net45),
    .A2(_4456_));
 sg13g2_inv_1 _6500_ (.Y(_1566_),
    .A(_1565_));
 sg13g2_a21oi_1 _6501_ (.A1(_1538_),
    .A2(_1551_),
    .Y(_1567_),
    .B1(_1566_));
 sg13g2_nor2_1 _6502_ (.A(_1564_),
    .B(_1567_),
    .Y(_1568_));
 sg13g2_a21oi_1 _6503_ (.A1(_1567_),
    .A2(_1564_),
    .Y(_1569_),
    .B1(_0318_));
 sg13g2_nand2b_1 _6504_ (.Y(_1570_),
    .B(_1569_),
    .A_N(_1568_));
 sg13g2_o21ai_1 _6505_ (.B1(_1570_),
    .Y(\generated._477[7] ),
    .A1(net44),
    .A2(_1562_));
 sg13g2_xnor2_1 _6506_ (.Y(_1571_),
    .A(\generated._369[8] ),
    .B(net85));
 sg13g2_nor2_1 _6507_ (.A(_1557_),
    .B(_1542_),
    .Y(_1572_));
 sg13g2_a21oi_1 _6508_ (.A1(_1549_),
    .A2(_1572_),
    .Y(_1573_),
    .B1(_1556_));
 sg13g2_xnor2_1 _6509_ (.Y(_1574_),
    .A(_1571_),
    .B(_1573_));
 sg13g2_nand2_1 _6510_ (.Y(_1575_),
    .A(_4492_),
    .B(_4473_));
 sg13g2_inv_1 _6511_ (.Y(_1576_),
    .A(_1575_));
 sg13g2_xnor2_1 _6512_ (.Y(_1577_),
    .A(_4492_),
    .B(_4483_));
 sg13g2_nor3_1 _6513_ (.A(_1576_),
    .B(_1577_),
    .C(_1568_),
    .Y(_1578_));
 sg13g2_o21ai_1 _6514_ (.B1(_1577_),
    .Y(_1579_),
    .A1(_1576_),
    .A2(_1568_));
 sg13g2_nand3b_1 _6515_ (.B(_1579_),
    .C(net62),
    .Y(_1580_),
    .A_N(_1578_));
 sg13g2_o21ai_1 _6516_ (.B1(_1580_),
    .Y(\generated._477[8] ),
    .A1(net44),
    .A2(_1574_));
 sg13g2_nand3b_1 _6517_ (.B(_1558_),
    .C(_1571_),
    .Y(_1581_),
    .A_N(_1561_));
 sg13g2_o21ai_1 _6518_ (.B1(net73),
    .Y(_1582_),
    .A1(\generated._369[8] ),
    .A2(\generated._369[7] ));
 sg13g2_nand3_1 _6519_ (.B(_0319_),
    .C(_1582_),
    .A(_1581_),
    .Y(_1583_));
 sg13g2_nand2_1 _6520_ (.Y(_1584_),
    .A(net68),
    .B(_4483_));
 sg13g2_nand3_1 _6521_ (.B(net62),
    .C(_1584_),
    .A(_1579_),
    .Y(_1585_));
 sg13g2_nand2_1 _6522_ (.Y(\generated._477[9] ),
    .A(_1583_),
    .B(_1585_));
 sg13g2_inv_1 _6523_ (.Y(_1586_),
    .A(\generated._483[2] ));
 sg13g2_nor3_1 _6524_ (.A(\generated._483[3] ),
    .B(_1586_),
    .C(_0303_),
    .Y(_1587_));
 sg13g2_nor2_1 _6525_ (.A(\generated._483[0] ),
    .B(_1587_),
    .Y(\generated._482[0] ));
 sg13g2_nand2_1 _6526_ (.Y(_1588_),
    .A(\generated._483[1] ),
    .B(\generated._483[0] ));
 sg13g2_inv_1 _6527_ (.Y(_1589_),
    .A(_1588_));
 sg13g2_nor2_1 _6528_ (.A(_0302_),
    .B(_1589_),
    .Y(\generated._482[1] ));
 sg13g2_xnor2_1 _6529_ (.Y(_1590_),
    .A(_1586_),
    .B(_1588_));
 sg13g2_nor2_1 _6530_ (.A(_1590_),
    .B(_1587_),
    .Y(\generated._482[2] ));
 sg13g2_nor2_1 _6531_ (.A(_1586_),
    .B(_1588_),
    .Y(_1591_));
 sg13g2_xor2_1 _6532_ (.B(_1591_),
    .A(\generated._483[3] ),
    .X(\generated._482[3] ));
 sg13g2_buf_1 _6533_ (.A(\generated._390[0] ),
    .X(_1592_));
 sg13g2_nand2_1 _6534_ (.Y(_1593_),
    .A(_1592_),
    .B(_0334_));
 sg13g2_nor2_1 _6535_ (.A(_1592_),
    .B(_0334_),
    .Y(_1594_));
 sg13g2_nor2_1 _6536_ (.A(_1493_),
    .B(_1594_),
    .Y(_1595_));
 sg13g2_a22oi_1 _6537_ (.Y(_1596_),
    .B1(_1593_),
    .B2(_1595_),
    .A2(_0448_),
    .A1(_1493_));
 sg13g2_buf_1 _6538_ (.A(_1596_),
    .X(_1597_));
 sg13g2_nor2_1 _6539_ (.A(net76),
    .B(_0432_),
    .Y(_1598_));
 sg13g2_o21ai_1 _6540_ (.B1(\generated._390[2] ),
    .Y(_1599_),
    .A1(_1592_),
    .A2(_0334_));
 sg13g2_nand2_1 _6541_ (.Y(_1600_),
    .A(_1594_),
    .B(_0348_));
 sg13g2_a21o_1 _6542_ (.A2(_1600_),
    .A1(_1599_),
    .B1(net68),
    .X(_1601_));
 sg13g2_nand2b_1 _6543_ (.Y(_1602_),
    .B(_1601_),
    .A_N(_1598_));
 sg13g2_buf_2 _6544_ (.A(_1602_),
    .X(_1603_));
 sg13g2_nor2_1 _6545_ (.A(_1597_),
    .B(_1603_),
    .Y(_1604_));
 sg13g2_inv_1 _6546_ (.Y(_1605_),
    .A(_1592_));
 sg13g2_inv_1 _6547_ (.Y(_1606_),
    .A(_1597_));
 sg13g2_inv_1 _6548_ (.Y(_1607_),
    .A(_1603_));
 sg13g2_nor2_1 _6549_ (.A(_1606_),
    .B(_1607_),
    .Y(_1608_));
 sg13g2_nor3_1 _6550_ (.A(_1605_),
    .B(_1604_),
    .C(_1608_),
    .Y(_1609_));
 sg13g2_nor2_1 _6551_ (.A(_1604_),
    .B(_1609_),
    .Y(_1610_));
 sg13g2_nor2_1 _6552_ (.A(net76),
    .B(_0445_),
    .Y(_1611_));
 sg13g2_nor3_1 _6553_ (.A(\generated._390[2] ),
    .B(_0334_),
    .C(_0282_),
    .Y(_1612_));
 sg13g2_nor2b_1 _6554_ (.A(_1612_),
    .B_N(_0365_),
    .Y(_1613_));
 sg13g2_inv_1 _6555_ (.Y(_1614_),
    .A(_1612_));
 sg13g2_nor2_1 _6556_ (.A(_0365_),
    .B(_1614_),
    .Y(_1615_));
 sg13g2_o21ai_1 _6557_ (.B1(_4490_),
    .Y(_1616_),
    .A1(_1613_),
    .A2(_1615_));
 sg13g2_nand2b_1 _6558_ (.Y(_1617_),
    .B(_1616_),
    .A_N(_1611_));
 sg13g2_buf_2 _6559_ (.A(_1617_),
    .X(_1618_));
 sg13g2_xnor2_1 _6560_ (.Y(_1619_),
    .A(_1603_),
    .B(_1618_));
 sg13g2_xnor2_1 _6561_ (.Y(_1620_),
    .A(_1606_),
    .B(_1619_));
 sg13g2_inv_1 _6562_ (.Y(_1621_),
    .A(_1620_));
 sg13g2_nor2_1 _6563_ (.A(_1610_),
    .B(_1621_),
    .Y(_1622_));
 sg13g2_a21oi_1 _6564_ (.A1(_1618_),
    .A2(_1603_),
    .Y(_1623_),
    .B1(_1592_));
 sg13g2_nor2_1 _6565_ (.A(_0106_),
    .B(_1597_),
    .Y(_1624_));
 sg13g2_o21ai_1 _6566_ (.B1(_1624_),
    .Y(_1625_),
    .A1(_1605_),
    .A2(_1607_));
 sg13g2_nor2_1 _6567_ (.A(_4490_),
    .B(_0458_),
    .Y(_1626_));
 sg13g2_o21ai_1 _6568_ (.B1(_0369_),
    .Y(_1627_),
    .A1(_0365_),
    .A2(_1600_));
 sg13g2_nor2_1 _6569_ (.A(_0365_),
    .B(_1600_),
    .Y(_1628_));
 sg13g2_nand2b_1 _6570_ (.Y(_1629_),
    .B(_1628_),
    .A_N(_0369_));
 sg13g2_a21o_1 _6571_ (.A2(_1629_),
    .A1(_1627_),
    .B1(net68),
    .X(_1630_));
 sg13g2_nand2b_1 _6572_ (.Y(_1631_),
    .B(_1630_),
    .A_N(_1626_));
 sg13g2_buf_2 _6573_ (.A(_1631_),
    .X(_1632_));
 sg13g2_inv_1 _6574_ (.Y(_1633_),
    .A(_1618_));
 sg13g2_xnor2_1 _6575_ (.Y(_1634_),
    .A(_1633_),
    .B(_1632_));
 sg13g2_nand2_1 _6576_ (.Y(_1635_),
    .A(_1634_),
    .B(_1607_));
 sg13g2_o21ai_1 _6577_ (.B1(_1635_),
    .Y(_1636_),
    .A1(_1618_),
    .A2(_1632_));
 sg13g2_inv_1 _6578_ (.Y(_1637_),
    .A(_1615_));
 sg13g2_o21ai_1 _6579_ (.B1(\generated._390[5] ),
    .Y(_1638_),
    .A1(_0369_),
    .A2(_1637_));
 sg13g2_nor2_1 _6580_ (.A(\generated._390[5] ),
    .B(_0369_),
    .Y(_1639_));
 sg13g2_nand2_1 _6581_ (.Y(_1640_),
    .A(_1615_),
    .B(_1639_));
 sg13g2_nand3_1 _6582_ (.B(net76),
    .C(_1640_),
    .A(_1638_),
    .Y(_1641_));
 sg13g2_o21ai_1 _6583_ (.B1(_1641_),
    .Y(_1642_),
    .A1(net76),
    .A2(_0371_));
 sg13g2_buf_2 _6584_ (.A(_1642_),
    .X(_1643_));
 sg13g2_xnor2_1 _6585_ (.Y(_1644_),
    .A(_1632_),
    .B(_1643_));
 sg13g2_xnor2_1 _6586_ (.Y(_1645_),
    .A(_1633_),
    .B(_1644_));
 sg13g2_xor2_1 _6587_ (.B(_1645_),
    .A(_1636_),
    .X(_1646_));
 sg13g2_xnor2_1 _6588_ (.Y(_1647_),
    .A(_1605_),
    .B(_1646_));
 sg13g2_xnor2_1 _6589_ (.Y(_1648_),
    .A(_1607_),
    .B(_1634_));
 sg13g2_inv_1 _6590_ (.Y(_1649_),
    .A(_1604_));
 sg13g2_o21ai_1 _6591_ (.B1(_1649_),
    .Y(_1650_),
    .A1(_1618_),
    .A2(_1608_));
 sg13g2_nor2b_1 _6592_ (.A(_1648_),
    .B_N(_1650_),
    .Y(_1651_));
 sg13g2_nor2b_1 _6593_ (.A(_1647_),
    .B_N(_1651_),
    .Y(_1652_));
 sg13g2_nor3_1 _6594_ (.A(_1623_),
    .B(_1625_),
    .C(_1652_),
    .Y(_1653_));
 sg13g2_xnor2_1 _6595_ (.Y(_1654_),
    .A(_1650_),
    .B(_1648_));
 sg13g2_nor2b_1 _6596_ (.A(_1647_),
    .B_N(_1654_),
    .Y(_1655_));
 sg13g2_o21ai_1 _6597_ (.B1(_1655_),
    .Y(_1656_),
    .A1(_1622_),
    .A2(_1653_));
 sg13g2_nor2b_1 _6598_ (.A(_1645_),
    .B_N(_1636_),
    .Y(_1657_));
 sg13g2_nor2_1 _6599_ (.A(_1605_),
    .B(_1646_),
    .Y(_1658_));
 sg13g2_nor2_1 _6600_ (.A(_1657_),
    .B(_1658_),
    .Y(_1659_));
 sg13g2_inv_1 _6601_ (.Y(_1660_),
    .A(_1632_));
 sg13g2_a21oi_1 _6602_ (.A1(_1628_),
    .A2(_1639_),
    .Y(_1661_),
    .B1(_0409_));
 sg13g2_nor3_1 _6603_ (.A(\generated._390[5] ),
    .B(_0408_),
    .C(_1629_),
    .Y(_1662_));
 sg13g2_nor2_1 _6604_ (.A(_1661_),
    .B(_1662_),
    .Y(_1663_));
 sg13g2_nor2_1 _6605_ (.A(_0059_),
    .B(net76),
    .Y(_1664_));
 sg13g2_a21oi_2 _6606_ (.B1(_1664_),
    .Y(_1665_),
    .A2(net63),
    .A1(_1663_));
 sg13g2_xnor2_1 _6607_ (.Y(_1666_),
    .A(_1665_),
    .B(_1643_));
 sg13g2_xnor2_1 _6608_ (.Y(_1667_),
    .A(_1660_),
    .B(_1666_));
 sg13g2_inv_1 _6609_ (.Y(_1668_),
    .A(_1644_));
 sg13g2_nand2_1 _6610_ (.Y(_1669_),
    .A(_1643_),
    .B(_1660_));
 sg13g2_o21ai_1 _6611_ (.B1(_1669_),
    .Y(_1670_),
    .A1(_1618_),
    .A2(_1668_));
 sg13g2_xor2_1 _6612_ (.B(_1670_),
    .A(_1667_),
    .X(_1671_));
 sg13g2_xnor2_1 _6613_ (.Y(_1672_),
    .A(_1597_),
    .B(_1671_));
 sg13g2_xnor2_1 _6614_ (.Y(_1673_),
    .A(_1659_),
    .B(_1672_));
 sg13g2_xnor2_1 _6615_ (.Y(_1674_),
    .A(_1652_),
    .B(_1673_));
 sg13g2_inv_1 _6616_ (.Y(_1675_),
    .A(_1674_));
 sg13g2_nor2_1 _6617_ (.A(_1656_),
    .B(_1675_),
    .Y(_1676_));
 sg13g2_inv_1 _6618_ (.Y(_1677_),
    .A(_1676_));
 sg13g2_buf_1 _6619_ (.A(_0584_),
    .X(_1678_));
 sg13g2_nand2_1 _6620_ (.Y(_1679_),
    .A(_1675_),
    .B(_1656_));
 sg13g2_nand3_1 _6621_ (.B(net38),
    .C(_1679_),
    .A(_1677_),
    .Y(_1680_));
 sg13g2_a22oi_1 _6622_ (.Y(_1681_),
    .B1(_0623_),
    .B2(_0569_),
    .A2(_0067_),
    .A1(_0567_));
 sg13g2_nand2_1 _6623_ (.Y(_1682_),
    .A(_0565_),
    .B(_0069_));
 sg13g2_o21ai_1 _6624_ (.B1(_1682_),
    .Y(_1683_),
    .A1(net84),
    .A2(_0630_));
 sg13g2_nand2_1 _6625_ (.Y(_1684_),
    .A(_1683_),
    .B(_0566_));
 sg13g2_and2_1 _6626_ (.A(_1681_),
    .B(_1684_),
    .X(_1685_));
 sg13g2_buf_1 _6627_ (.A(_1685_),
    .X(_1686_));
 sg13g2_nor2_1 _6628_ (.A(_0065_),
    .B(_1686_),
    .Y(_1687_));
 sg13g2_inv_1 _6629_ (.Y(_1688_),
    .A(_0065_));
 sg13g2_nor2b_1 _6630_ (.A(_1688_),
    .B_N(_1686_),
    .Y(_1689_));
 sg13g2_o21ai_1 _6631_ (.B1(net56),
    .Y(_1690_),
    .A1(_1687_),
    .A2(_1689_));
 sg13g2_nand2_1 _6632_ (.Y(\generated._557[0] ),
    .A(_1680_),
    .B(_1690_));
 sg13g2_nor2_1 _6633_ (.A(_1659_),
    .B(_1672_),
    .Y(_1691_));
 sg13g2_nor2b_1 _6634_ (.A(_1667_),
    .B_N(_1670_),
    .Y(_1692_));
 sg13g2_nor2_1 _6635_ (.A(_1597_),
    .B(_1671_),
    .Y(_1693_));
 sg13g2_nor2_1 _6636_ (.A(_1692_),
    .B(_1693_),
    .Y(_1694_));
 sg13g2_inv_1 _6637_ (.Y(_1695_),
    .A(_1666_));
 sg13g2_inv_1 _6638_ (.Y(_1696_),
    .A(_1665_));
 sg13g2_nand2_1 _6639_ (.Y(_1697_),
    .A(_1643_),
    .B(_1696_));
 sg13g2_o21ai_1 _6640_ (.B1(_1697_),
    .Y(_1698_),
    .A1(_1632_),
    .A2(_1695_));
 sg13g2_nor3_1 _6641_ (.A(_0408_),
    .B(\generated._390[7] ),
    .C(_1640_),
    .Y(_1699_));
 sg13g2_o21ai_1 _6642_ (.B1(\generated._390[7] ),
    .Y(_1700_),
    .A1(_0408_),
    .A2(_1640_));
 sg13g2_nand2b_1 _6643_ (.Y(_1701_),
    .B(_1700_),
    .A_N(_1699_));
 sg13g2_nor2_1 _6644_ (.A(net76),
    .B(_0504_),
    .Y(_1702_));
 sg13g2_a21o_1 _6645_ (.A2(net63),
    .A1(_1701_),
    .B1(_1702_),
    .X(_1703_));
 sg13g2_buf_2 _6646_ (.A(_1703_),
    .X(_1704_));
 sg13g2_xnor2_1 _6647_ (.Y(_1705_),
    .A(_1665_),
    .B(_1704_));
 sg13g2_xor2_1 _6648_ (.B(_1705_),
    .A(_1643_),
    .X(_1706_));
 sg13g2_xor2_1 _6649_ (.B(_1706_),
    .A(_1698_),
    .X(_1707_));
 sg13g2_xnor2_1 _6650_ (.Y(_1708_),
    .A(_1603_),
    .B(_1707_));
 sg13g2_xnor2_1 _6651_ (.Y(_1709_),
    .A(_1694_),
    .B(_1708_));
 sg13g2_xnor2_1 _6652_ (.Y(_1710_),
    .A(_1691_),
    .B(_1709_));
 sg13g2_inv_1 _6653_ (.Y(_1711_),
    .A(_1710_));
 sg13g2_nor2_1 _6654_ (.A(_1711_),
    .B(_1677_),
    .Y(_1712_));
 sg13g2_nand2b_1 _6655_ (.Y(_1713_),
    .B(_1652_),
    .A_N(_1673_));
 sg13g2_xor2_1 _6656_ (.B(_1710_),
    .A(_1713_),
    .X(_1714_));
 sg13g2_nand2_1 _6657_ (.Y(_1715_),
    .A(_1714_),
    .B(_1677_));
 sg13g2_nand2_1 _6658_ (.Y(_1716_),
    .A(_1715_),
    .B(net38));
 sg13g2_nand2_1 _6659_ (.Y(_1717_),
    .A(_1686_),
    .B(_0591_));
 sg13g2_nand2_1 _6660_ (.Y(_1718_),
    .A(net84),
    .B(_0072_));
 sg13g2_o21ai_1 _6661_ (.B1(_1718_),
    .Y(_1719_),
    .A1(net84),
    .A2(_0657_));
 sg13g2_nor3_1 _6662_ (.A(_0566_),
    .B(_0568_),
    .C(_0630_),
    .Y(_1720_));
 sg13g2_a221oi_1 _6663_ (.B2(net83),
    .C1(_1720_),
    .B1(_1719_),
    .A1(_0623_),
    .Y(_1721_),
    .A2(_0567_));
 sg13g2_xor2_1 _6664_ (.B(_1721_),
    .A(_1717_),
    .X(_1722_));
 sg13g2_xnor2_1 _6665_ (.Y(_1723_),
    .A(_0597_),
    .B(_1722_));
 sg13g2_or2_1 _6666_ (.X(_1724_),
    .B(_1723_),
    .A(_1689_));
 sg13g2_nand2_1 _6667_ (.Y(_1725_),
    .A(_1723_),
    .B(_1689_));
 sg13g2_nand3_1 _6668_ (.B(net59),
    .C(_1725_),
    .A(_1724_),
    .Y(_1726_));
 sg13g2_o21ai_1 _6669_ (.B1(_1726_),
    .Y(\generated._557[1] ),
    .A1(_1712_),
    .A2(_1716_));
 sg13g2_nor2_1 _6670_ (.A(net84),
    .B(_0676_),
    .Y(_1727_));
 sg13g2_a21oi_1 _6671_ (.A1(net84),
    .A2(_0075_),
    .Y(_1728_),
    .B1(_1727_));
 sg13g2_nor2_1 _6672_ (.A(_0608_),
    .B(_1728_),
    .Y(_1729_));
 sg13g2_a21oi_1 _6673_ (.A1(net58),
    .A2(_1683_),
    .Y(_1730_),
    .B1(_1729_));
 sg13g2_nor2_1 _6674_ (.A(_1686_),
    .B(_1721_),
    .Y(_1731_));
 sg13g2_nor2_1 _6675_ (.A(net57),
    .B(_1731_),
    .Y(_1732_));
 sg13g2_xnor2_1 _6676_ (.Y(_1733_),
    .A(_1730_),
    .B(_1732_));
 sg13g2_xnor2_1 _6677_ (.Y(_1734_),
    .A(_0572_),
    .B(_1733_));
 sg13g2_buf_1 _6678_ (.A(\generated._558[1] ),
    .X(_1735_));
 sg13g2_nand2_1 _6679_ (.Y(_1736_),
    .A(_1722_),
    .B(_1735_));
 sg13g2_nand2_1 _6680_ (.Y(_1737_),
    .A(_1724_),
    .B(_1736_));
 sg13g2_nor2_1 _6681_ (.A(_1734_),
    .B(_1737_),
    .Y(_1738_));
 sg13g2_nand2_1 _6682_ (.Y(_1739_),
    .A(_1737_),
    .B(_1734_));
 sg13g2_nand2_1 _6683_ (.Y(_1740_),
    .A(_1739_),
    .B(net72));
 sg13g2_nor2b_1 _6684_ (.A(_1709_),
    .B_N(_1691_),
    .Y(_1741_));
 sg13g2_inv_1 _6685_ (.Y(_1742_),
    .A(_1741_));
 sg13g2_nor2_1 _6686_ (.A(_1694_),
    .B(_1708_),
    .Y(_1743_));
 sg13g2_nor2b_1 _6687_ (.A(_1706_),
    .B_N(_1698_),
    .Y(_1744_));
 sg13g2_nor2_1 _6688_ (.A(_1603_),
    .B(_1707_),
    .Y(_1745_));
 sg13g2_nor2_1 _6689_ (.A(_1744_),
    .B(_1745_),
    .Y(_1746_));
 sg13g2_nand2b_1 _6690_ (.Y(_1747_),
    .B(_1643_),
    .A_N(_1705_));
 sg13g2_o21ai_1 _6691_ (.B1(_1747_),
    .Y(_1748_),
    .A1(_1665_),
    .A2(_1704_));
 sg13g2_nand2b_1 _6692_ (.Y(_1749_),
    .B(_1662_),
    .A_N(\generated._390[7] ));
 sg13g2_xnor2_1 _6693_ (.Y(_1750_),
    .A(_0428_),
    .B(_1749_));
 sg13g2_nor2_1 _6694_ (.A(net76),
    .B(_0414_),
    .Y(_1751_));
 sg13g2_a21o_1 _6695_ (.A2(net63),
    .A1(_1750_),
    .B1(_1751_),
    .X(_1752_));
 sg13g2_buf_1 _6696_ (.A(_1752_),
    .X(_1753_));
 sg13g2_inv_1 _6697_ (.Y(_1754_),
    .A(_1753_));
 sg13g2_nand2_1 _6698_ (.Y(_1755_),
    .A(_1754_),
    .B(_1704_));
 sg13g2_inv_1 _6699_ (.Y(_1756_),
    .A(_1704_));
 sg13g2_nand2_1 _6700_ (.Y(_1757_),
    .A(_1753_),
    .B(_1756_));
 sg13g2_a21oi_1 _6701_ (.A1(_1755_),
    .A2(_1757_),
    .Y(_1758_),
    .B1(_1696_));
 sg13g2_nand3_1 _6702_ (.B(_1696_),
    .C(_1757_),
    .A(_1755_),
    .Y(_1759_));
 sg13g2_nand2b_1 _6703_ (.Y(_1760_),
    .B(_1759_),
    .A_N(_1758_));
 sg13g2_xor2_1 _6704_ (.B(_1760_),
    .A(_1748_),
    .X(_1761_));
 sg13g2_xnor2_1 _6705_ (.Y(_1762_),
    .A(_1618_),
    .B(_1761_));
 sg13g2_xnor2_1 _6706_ (.Y(_1763_),
    .A(_1746_),
    .B(_1762_));
 sg13g2_xor2_1 _6707_ (.B(_1763_),
    .A(_1743_),
    .X(_1764_));
 sg13g2_xnor2_1 _6708_ (.Y(_1765_),
    .A(_1742_),
    .B(_1764_));
 sg13g2_a21o_1 _6709_ (.A2(_1713_),
    .A1(_1677_),
    .B1(_1711_),
    .X(_1766_));
 sg13g2_nor2_1 _6710_ (.A(_1765_),
    .B(_1766_),
    .Y(_1767_));
 sg13g2_nand2_1 _6711_ (.Y(_1768_),
    .A(_1766_),
    .B(_1765_));
 sg13g2_nand3b_1 _6712_ (.B(net38),
    .C(_1768_),
    .Y(_1769_),
    .A_N(_1767_));
 sg13g2_o21ai_1 _6713_ (.B1(_1769_),
    .Y(\generated._557[2] ),
    .A1(_1738_),
    .A2(_1740_));
 sg13g2_nand2b_1 _6714_ (.Y(_1770_),
    .B(_1743_),
    .A_N(_1763_));
 sg13g2_nor2_1 _6715_ (.A(_1746_),
    .B(_1762_),
    .Y(_1771_));
 sg13g2_nand2_1 _6716_ (.Y(_1772_),
    .A(_1759_),
    .B(_1757_));
 sg13g2_nand2_1 _6717_ (.Y(_1773_),
    .A(_1699_),
    .B(_0428_));
 sg13g2_xnor2_1 _6718_ (.Y(_1774_),
    .A(_0559_),
    .B(_1773_));
 sg13g2_nor2_1 _6719_ (.A(_4491_),
    .B(_0422_),
    .Y(_1775_));
 sg13g2_a21o_1 _6720_ (.A2(_4491_),
    .A1(_1774_),
    .B1(_1775_),
    .X(_1776_));
 sg13g2_buf_1 _6721_ (.A(_1776_),
    .X(_1777_));
 sg13g2_xnor2_1 _6722_ (.Y(_1778_),
    .A(_1753_),
    .B(_1777_));
 sg13g2_xnor2_1 _6723_ (.Y(_1779_),
    .A(_1704_),
    .B(_1778_));
 sg13g2_xor2_1 _6724_ (.B(_1779_),
    .A(_1772_),
    .X(_1780_));
 sg13g2_xnor2_1 _6725_ (.Y(_1781_),
    .A(_1632_),
    .B(_1780_));
 sg13g2_nor2b_1 _6726_ (.A(_1760_),
    .B_N(_1748_),
    .Y(_1782_));
 sg13g2_nor2_1 _6727_ (.A(_1618_),
    .B(_1761_),
    .Y(_1783_));
 sg13g2_nor2_1 _6728_ (.A(_1782_),
    .B(_1783_),
    .Y(_1784_));
 sg13g2_xnor2_1 _6729_ (.Y(_1785_),
    .A(_1781_),
    .B(_1784_));
 sg13g2_xor2_1 _6730_ (.B(_1785_),
    .A(_1771_),
    .X(_1786_));
 sg13g2_xnor2_1 _6731_ (.Y(_1787_),
    .A(_1770_),
    .B(_1786_));
 sg13g2_nor2_1 _6732_ (.A(_1742_),
    .B(_1764_),
    .Y(_1788_));
 sg13g2_nor2_1 _6733_ (.A(_1788_),
    .B(_1767_),
    .Y(_1789_));
 sg13g2_xnor2_1 _6734_ (.Y(_1790_),
    .A(_1787_),
    .B(_1789_));
 sg13g2_nor2_1 _6735_ (.A(net71),
    .B(_0682_),
    .Y(_1791_));
 sg13g2_a21oi_1 _6736_ (.A1(net71),
    .A2(_0078_),
    .Y(_1792_),
    .B1(_1791_));
 sg13g2_nor2_1 _6737_ (.A(_0609_),
    .B(_1792_),
    .Y(_1793_));
 sg13g2_a21oi_1 _6738_ (.A1(_0609_),
    .A2(_1719_),
    .Y(_1794_),
    .B1(_1793_));
 sg13g2_inv_1 _6739_ (.Y(_1795_),
    .A(_1731_));
 sg13g2_nor2_1 _6740_ (.A(_1730_),
    .B(_1795_),
    .Y(_1796_));
 sg13g2_nor2_1 _6741_ (.A(net57),
    .B(_1796_),
    .Y(_1797_));
 sg13g2_xnor2_1 _6742_ (.Y(_1798_),
    .A(_1794_),
    .B(_1797_));
 sg13g2_xnor2_1 _6743_ (.Y(_1799_),
    .A(_0077_),
    .B(_1798_));
 sg13g2_inv_1 _6744_ (.Y(_1800_),
    .A(_1799_));
 sg13g2_inv_1 _6745_ (.Y(_1801_),
    .A(\generated._558[2] ));
 sg13g2_inv_1 _6746_ (.Y(_1802_),
    .A(_1733_));
 sg13g2_o21ai_1 _6747_ (.B1(_1739_),
    .Y(_1803_),
    .A1(_1801_),
    .A2(_1802_));
 sg13g2_inv_1 _6748_ (.Y(_1804_),
    .A(_1803_));
 sg13g2_nor2_1 _6749_ (.A(_1800_),
    .B(_1804_),
    .Y(_1805_));
 sg13g2_inv_1 _6750_ (.Y(_1806_),
    .A(_1805_));
 sg13g2_nand2_1 _6751_ (.Y(_1807_),
    .A(_1804_),
    .B(_1800_));
 sg13g2_nand3_1 _6752_ (.B(net59),
    .C(_1807_),
    .A(_1806_),
    .Y(_1808_));
 sg13g2_o21ai_1 _6753_ (.B1(_1808_),
    .Y(\generated._557[3] ),
    .A1(net56),
    .A2(_1790_));
 sg13g2_nand2_1 _6754_ (.Y(_1809_),
    .A(net71),
    .B(_0720_));
 sg13g2_o21ai_1 _6755_ (.B1(_1809_),
    .Y(_1810_),
    .A1(net71),
    .A2(_0707_));
 sg13g2_nor2_1 _6756_ (.A(net83),
    .B(_1728_),
    .Y(_1811_));
 sg13g2_a21oi_1 _6757_ (.A1(net83),
    .A2(_1810_),
    .Y(_1812_),
    .B1(_1811_));
 sg13g2_inv_1 _6758_ (.Y(_1813_),
    .A(_1796_));
 sg13g2_nor2_1 _6759_ (.A(_1794_),
    .B(_1813_),
    .Y(_1814_));
 sg13g2_nor2_1 _6760_ (.A(_0618_),
    .B(_1814_),
    .Y(_1815_));
 sg13g2_xnor2_1 _6761_ (.Y(_1816_),
    .A(_1812_),
    .B(_1815_));
 sg13g2_xnor2_1 _6762_ (.Y(_1817_),
    .A(_0594_),
    .B(_1816_));
 sg13g2_inv_1 _6763_ (.Y(_1818_),
    .A(_1817_));
 sg13g2_a21o_1 _6764_ (.A2(_1798_),
    .A1(\generated._558[3] ),
    .B1(_1805_),
    .X(_1819_));
 sg13g2_inv_1 _6765_ (.Y(_1820_),
    .A(_1819_));
 sg13g2_nor2_1 _6766_ (.A(_1818_),
    .B(_1820_),
    .Y(_1821_));
 sg13g2_o21ai_1 _6767_ (.B1(net72),
    .Y(_1822_),
    .A1(_1817_),
    .A2(_1819_));
 sg13g2_nor2_1 _6768_ (.A(_1770_),
    .B(_1786_),
    .Y(_1823_));
 sg13g2_nor2_1 _6769_ (.A(_1787_),
    .B(_1789_),
    .Y(_1824_));
 sg13g2_nor2_1 _6770_ (.A(_1823_),
    .B(_1824_),
    .Y(_1825_));
 sg13g2_nand2b_1 _6771_ (.Y(_1826_),
    .B(_1771_),
    .A_N(_1785_));
 sg13g2_or2_1 _6772_ (.X(_1827_),
    .B(_1784_),
    .A(_1781_));
 sg13g2_inv_1 _6773_ (.Y(_1828_),
    .A(_1777_));
 sg13g2_nor2_1 _6774_ (.A(_1704_),
    .B(_1828_),
    .Y(_1829_));
 sg13g2_inv_1 _6775_ (.Y(_1830_),
    .A(_1829_));
 sg13g2_nor2_1 _6776_ (.A(_1756_),
    .B(_1777_),
    .Y(_1831_));
 sg13g2_nor2_1 _6777_ (.A(_1754_),
    .B(_1831_),
    .Y(_1832_));
 sg13g2_a21oi_1 _6778_ (.A1(_1830_),
    .A2(_1754_),
    .Y(_1833_),
    .B1(_1832_));
 sg13g2_xnor2_1 _6779_ (.Y(_1834_),
    .A(_1643_),
    .B(_1833_));
 sg13g2_nor2b_1 _6780_ (.A(_1779_),
    .B_N(_1772_),
    .Y(_1835_));
 sg13g2_nor2_1 _6781_ (.A(_1632_),
    .B(_1780_),
    .Y(_1836_));
 sg13g2_nor2_1 _6782_ (.A(_1835_),
    .B(_1836_),
    .Y(_1837_));
 sg13g2_xor2_1 _6783_ (.B(_1837_),
    .A(_1834_),
    .X(_1838_));
 sg13g2_xor2_1 _6784_ (.B(_1838_),
    .A(_1827_),
    .X(_1839_));
 sg13g2_xnor2_1 _6785_ (.Y(_1840_),
    .A(_1826_),
    .B(_1839_));
 sg13g2_a21oi_1 _6786_ (.A1(_1825_),
    .A2(_1840_),
    .Y(_1841_),
    .B1(net72));
 sg13g2_nor2_1 _6787_ (.A(_1840_),
    .B(_1825_),
    .Y(_1842_));
 sg13g2_inv_1 _6788_ (.Y(_1843_),
    .A(_1842_));
 sg13g2_nand2_1 _6789_ (.Y(_1844_),
    .A(_1841_),
    .B(_1843_));
 sg13g2_o21ai_1 _6790_ (.B1(_1844_),
    .Y(\generated._557[4] ),
    .A1(_1821_),
    .A2(_1822_));
 sg13g2_a21oi_1 _6791_ (.A1(_1833_),
    .A2(_1643_),
    .Y(_1845_),
    .B1(_1832_));
 sg13g2_xnor2_1 _6792_ (.Y(_1846_),
    .A(_1696_),
    .B(_1845_));
 sg13g2_nor2_1 _6793_ (.A(_1834_),
    .B(_1837_),
    .Y(_1847_));
 sg13g2_inv_1 _6794_ (.Y(_1848_),
    .A(_1838_));
 sg13g2_nor2_1 _6795_ (.A(_1827_),
    .B(_1848_),
    .Y(_1849_));
 sg13g2_nor2_1 _6796_ (.A(_1847_),
    .B(_1849_),
    .Y(_1850_));
 sg13g2_xnor2_1 _6797_ (.Y(_1851_),
    .A(_1846_),
    .B(_1850_));
 sg13g2_inv_1 _6798_ (.Y(_1852_),
    .A(_1851_));
 sg13g2_o21ai_1 _6799_ (.B1(_1843_),
    .Y(_1853_),
    .A1(_1826_),
    .A2(_1839_));
 sg13g2_inv_1 _6800_ (.Y(_1854_),
    .A(_1853_));
 sg13g2_nor2_1 _6801_ (.A(_1852_),
    .B(_1854_),
    .Y(_1855_));
 sg13g2_o21ai_1 _6802_ (.B1(net38),
    .Y(_1856_),
    .A1(_1851_),
    .A2(_1853_));
 sg13g2_nand2_1 _6803_ (.Y(_1857_),
    .A(_0727_),
    .B(net55));
 sg13g2_o21ai_1 _6804_ (.B1(_1857_),
    .Y(_1858_),
    .A1(net55),
    .A2(_0720_));
 sg13g2_inv_1 _6805_ (.Y(_1859_),
    .A(_1858_));
 sg13g2_nor2_1 _6806_ (.A(_0607_),
    .B(_1792_),
    .Y(_1860_));
 sg13g2_a21oi_1 _6807_ (.A1(_0607_),
    .A2(_1859_),
    .Y(_1861_),
    .B1(_1860_));
 sg13g2_inv_1 _6808_ (.Y(_1862_),
    .A(_1814_));
 sg13g2_nor2_1 _6809_ (.A(_1812_),
    .B(_1862_),
    .Y(_1863_));
 sg13g2_nor2_1 _6810_ (.A(net57),
    .B(_1863_),
    .Y(_1864_));
 sg13g2_xnor2_1 _6811_ (.Y(_1865_),
    .A(_1861_),
    .B(_1864_));
 sg13g2_xnor2_1 _6812_ (.Y(_1866_),
    .A(_0081_),
    .B(_1865_));
 sg13g2_inv_1 _6813_ (.Y(_1867_),
    .A(_1866_));
 sg13g2_buf_1 _6814_ (.A(\generated._558[4] ),
    .X(_1868_));
 sg13g2_a21oi_1 _6815_ (.A1(_1868_),
    .A2(_1816_),
    .Y(_1869_),
    .B1(_1821_));
 sg13g2_nor2_1 _6816_ (.A(_1867_),
    .B(_1869_),
    .Y(_1870_));
 sg13g2_a21oi_1 _6817_ (.A1(_1869_),
    .A2(_1867_),
    .Y(_1871_),
    .B1(_0584_));
 sg13g2_nand2b_1 _6818_ (.Y(_1872_),
    .B(_1871_),
    .A_N(_1870_));
 sg13g2_o21ai_1 _6819_ (.B1(_1872_),
    .Y(\generated._557[5] ),
    .A1(_1855_),
    .A2(_1856_));
 sg13g2_a21o_1 _6820_ (.A2(_1846_),
    .A1(_1849_),
    .B1(_1855_),
    .X(_1873_));
 sg13g2_nor2_1 _6821_ (.A(_1831_),
    .B(_1829_),
    .Y(_1874_));
 sg13g2_nor2_1 _6822_ (.A(_1665_),
    .B(_1845_),
    .Y(_1875_));
 sg13g2_nand2_1 _6823_ (.Y(_1876_),
    .A(_1847_),
    .B(_1846_));
 sg13g2_inv_1 _6824_ (.Y(_1877_),
    .A(_1876_));
 sg13g2_nor2_1 _6825_ (.A(_1875_),
    .B(_1877_),
    .Y(_1878_));
 sg13g2_xnor2_1 _6826_ (.Y(_1879_),
    .A(_1874_),
    .B(_1878_));
 sg13g2_nand2_1 _6827_ (.Y(_1880_),
    .A(_1873_),
    .B(_1879_));
 sg13g2_inv_1 _6828_ (.Y(_1881_),
    .A(_1880_));
 sg13g2_o21ai_1 _6829_ (.B1(_1678_),
    .Y(_1882_),
    .A1(_1879_),
    .A2(_1873_));
 sg13g2_buf_1 _6830_ (.A(\generated._558[5] ),
    .X(_1883_));
 sg13g2_a21oi_1 _6831_ (.A1(_1883_),
    .A2(_1865_),
    .Y(_1884_),
    .B1(_1870_));
 sg13g2_buf_1 _6832_ (.A(_0084_),
    .X(_1885_));
 sg13g2_nand2_1 _6833_ (.Y(_1886_),
    .A(_0665_),
    .B(_1885_));
 sg13g2_o21ai_1 _6834_ (.B1(_1886_),
    .Y(_1887_),
    .A1(_0665_),
    .A2(_0727_));
 sg13g2_nor2b_1 _6835_ (.A(net70),
    .B_N(_1810_),
    .Y(_1888_));
 sg13g2_a21oi_1 _6836_ (.A1(_0664_),
    .A2(_1887_),
    .Y(_1889_),
    .B1(_1888_));
 sg13g2_inv_1 _6837_ (.Y(_1890_),
    .A(_1863_));
 sg13g2_nor2_1 _6838_ (.A(_1861_),
    .B(_1890_),
    .Y(_1891_));
 sg13g2_nor2_1 _6839_ (.A(net42),
    .B(_1891_),
    .Y(_1892_));
 sg13g2_xnor2_1 _6840_ (.Y(_1893_),
    .A(_1889_),
    .B(_1892_));
 sg13g2_xnor2_1 _6841_ (.Y(_1894_),
    .A(_0634_),
    .B(_1893_));
 sg13g2_inv_1 _6842_ (.Y(_1895_),
    .A(_1894_));
 sg13g2_a21oi_1 _6843_ (.A1(_1884_),
    .A2(_1895_),
    .Y(_1896_),
    .B1(_1678_));
 sg13g2_nor2_1 _6844_ (.A(_1895_),
    .B(_1884_),
    .Y(_1897_));
 sg13g2_inv_1 _6845_ (.Y(_1898_),
    .A(_1897_));
 sg13g2_nand2_1 _6846_ (.Y(_1899_),
    .A(_1896_),
    .B(_1898_));
 sg13g2_o21ai_1 _6847_ (.B1(_1899_),
    .Y(\generated._557[6] ),
    .A1(_1881_),
    .A2(_1882_));
 sg13g2_o21ai_1 _6848_ (.B1(_1757_),
    .Y(_1900_),
    .A1(_1756_),
    .A2(_1778_));
 sg13g2_nand2_1 _6849_ (.Y(_1901_),
    .A(_1875_),
    .B(_1874_));
 sg13g2_inv_1 _6850_ (.Y(_1902_),
    .A(_1901_));
 sg13g2_nor2_1 _6851_ (.A(_1900_),
    .B(_1902_),
    .Y(_1903_));
 sg13g2_nand2_1 _6852_ (.Y(_1904_),
    .A(_1902_),
    .B(_1900_));
 sg13g2_nor2b_1 _6853_ (.A(_1903_),
    .B_N(_1904_),
    .Y(_1905_));
 sg13g2_nand2_1 _6854_ (.Y(_1906_),
    .A(_1877_),
    .B(_1874_));
 sg13g2_nand2_1 _6855_ (.Y(_1907_),
    .A(_1880_),
    .B(_1906_));
 sg13g2_xnor2_1 _6856_ (.Y(_1908_),
    .A(_1905_),
    .B(_1907_));
 sg13g2_buf_1 _6857_ (.A(\generated._558[6] ),
    .X(_1909_));
 sg13g2_a21o_1 _6858_ (.A2(_1893_),
    .A1(_1909_),
    .B1(_1897_),
    .X(_1910_));
 sg13g2_inv_1 _6859_ (.Y(_1911_),
    .A(_1910_));
 sg13g2_nand2_1 _6860_ (.Y(_1912_),
    .A(_0664_),
    .B(_1885_));
 sg13g2_inv_1 _6861_ (.Y(_1913_),
    .A(_1912_));
 sg13g2_a21oi_1 _6862_ (.A1(_1859_),
    .A2(net58),
    .Y(_1914_),
    .B1(_1913_));
 sg13g2_inv_1 _6863_ (.Y(_1915_),
    .A(_1891_));
 sg13g2_nor2_1 _6864_ (.A(_1889_),
    .B(_1915_),
    .Y(_1916_));
 sg13g2_nor2_1 _6865_ (.A(net42),
    .B(_1916_),
    .Y(_1917_));
 sg13g2_xnor2_1 _6866_ (.Y(_1918_),
    .A(_1914_),
    .B(_1917_));
 sg13g2_xnor2_1 _6867_ (.Y(_1919_),
    .A(_0085_),
    .B(_1918_));
 sg13g2_inv_1 _6868_ (.Y(_1920_),
    .A(_1919_));
 sg13g2_a21oi_1 _6869_ (.A1(_1911_),
    .A2(_1920_),
    .Y(_1921_),
    .B1(_0584_));
 sg13g2_nor2_1 _6870_ (.A(_1920_),
    .B(_1911_),
    .Y(_1922_));
 sg13g2_inv_1 _6871_ (.Y(_1923_),
    .A(_1922_));
 sg13g2_nand2_1 _6872_ (.Y(_1924_),
    .A(_1921_),
    .B(_1923_));
 sg13g2_o21ai_1 _6873_ (.B1(_1924_),
    .Y(\generated._557[7] ),
    .A1(net56),
    .A2(_1908_));
 sg13g2_a21oi_2 _6874_ (.B1(_1913_),
    .Y(_1925_),
    .A2(net58),
    .A1(_1887_));
 sg13g2_inv_1 _6875_ (.Y(_1926_),
    .A(_1916_));
 sg13g2_nor2_1 _6876_ (.A(_1914_),
    .B(_1926_),
    .Y(_1927_));
 sg13g2_nor2_1 _6877_ (.A(net42),
    .B(_1927_),
    .Y(_1928_));
 sg13g2_xnor2_1 _6878_ (.Y(_1929_),
    .A(_1925_),
    .B(_1928_));
 sg13g2_xnor2_1 _6879_ (.Y(_1930_),
    .A(_0666_),
    .B(_1929_));
 sg13g2_inv_1 _6880_ (.Y(_1931_),
    .A(_1930_));
 sg13g2_a21o_1 _6881_ (.A2(_1918_),
    .A1(\generated._558[7] ),
    .B1(_1922_),
    .X(_1932_));
 sg13g2_inv_1 _6882_ (.Y(_1933_),
    .A(_1932_));
 sg13g2_nor2_1 _6883_ (.A(_1931_),
    .B(_1933_),
    .Y(_1934_));
 sg13g2_o21ai_1 _6884_ (.B1(_0581_),
    .Y(_1935_),
    .A1(_1930_),
    .A2(_1932_));
 sg13g2_and3_1 _6885_ (.X(_1936_),
    .A(_1880_),
    .B(_1906_),
    .C(_1904_));
 sg13g2_nand2_1 _6886_ (.Y(_1937_),
    .A(_1755_),
    .B(_1777_));
 sg13g2_o21ai_1 _6887_ (.B1(_1937_),
    .Y(_1938_),
    .A1(_1903_),
    .A2(_1936_));
 sg13g2_nand2_1 _6888_ (.Y(_1939_),
    .A(_1938_),
    .B(_0585_));
 sg13g2_o21ai_1 _6889_ (.B1(_1939_),
    .Y(\generated._557[8] ),
    .A1(_1934_),
    .A2(_1935_));
 sg13g2_inv_1 _6890_ (.Y(_1940_),
    .A(_1927_));
 sg13g2_nor3_1 _6891_ (.A(_0729_),
    .B(_1925_),
    .C(_1940_),
    .Y(_1941_));
 sg13g2_o21ai_1 _6892_ (.B1(_0729_),
    .Y(_1942_),
    .A1(_1925_),
    .A2(_1940_));
 sg13g2_nand3b_1 _6893_ (.B(_1942_),
    .C(_0616_),
    .Y(_1943_),
    .A_N(_1941_));
 sg13g2_o21ai_1 _6894_ (.B1(_1943_),
    .Y(_1944_),
    .A1(_0616_),
    .A2(_1885_));
 sg13g2_xnor2_1 _6895_ (.Y(_1945_),
    .A(_0687_),
    .B(_1944_));
 sg13g2_a21oi_1 _6896_ (.A1(\generated._558[8] ),
    .A2(_1929_),
    .Y(_1946_),
    .B1(_1934_));
 sg13g2_a21oi_1 _6897_ (.A1(_1946_),
    .A2(_1945_),
    .Y(_1947_),
    .B1(_0584_));
 sg13g2_o21ai_1 _6898_ (.B1(_1947_),
    .Y(_1948_),
    .A1(_1945_),
    .A2(_1946_));
 sg13g2_o21ai_1 _6899_ (.B1(_1948_),
    .Y(\generated._557[9] ),
    .A1(_0627_),
    .A2(_1828_));
 sg13g2_nand3_1 _6900_ (.B(\generated._61[2] ),
    .C(_0579_),
    .A(_0577_),
    .Y(_1949_));
 sg13g2_nor2b_1 _6901_ (.A(\generated._61[0] ),
    .B_N(_1949_),
    .Y(\generated._60[0] ));
 sg13g2_nand2_1 _6902_ (.Y(_1950_),
    .A(\generated._61[1] ),
    .B(\generated._61[0] ));
 sg13g2_inv_1 _6903_ (.Y(_1951_),
    .A(_1950_));
 sg13g2_nor2_1 _6904_ (.A(_0577_),
    .B(_1951_),
    .Y(\generated._60[1] ));
 sg13g2_nand2_1 _6905_ (.Y(_1952_),
    .A(_1951_),
    .B(\generated._61[2] ));
 sg13g2_nand2_1 _6906_ (.Y(_1953_),
    .A(_1950_),
    .B(_0578_));
 sg13g2_and3_1 _6907_ (.X(\generated._60[2] ),
    .A(_1949_),
    .B(_1952_),
    .C(_1953_));
 sg13g2_xnor2_1 _6908_ (.Y(\generated._60[3] ),
    .A(\generated._61[3] ),
    .B(_1952_));
 sg13g2_nand3_1 _6909_ (.B(\generated._69[2] ),
    .C(_0753_),
    .A(_0751_),
    .Y(_1954_));
 sg13g2_nor2b_1 _6910_ (.A(\generated._69[0] ),
    .B_N(_1954_),
    .Y(\generated._68[0] ));
 sg13g2_nand2_1 _6911_ (.Y(_1955_),
    .A(\generated._69[1] ),
    .B(\generated._69[0] ));
 sg13g2_inv_1 _6912_ (.Y(_1956_),
    .A(_1955_));
 sg13g2_nor2_1 _6913_ (.A(_0751_),
    .B(_1956_),
    .Y(\generated._68[1] ));
 sg13g2_nand2_1 _6914_ (.Y(_1957_),
    .A(_1956_),
    .B(\generated._69[2] ));
 sg13g2_nand2_1 _6915_ (.Y(_1958_),
    .A(_1955_),
    .B(_0752_));
 sg13g2_and3_1 _6916_ (.X(\generated._68[2] ),
    .A(_1954_),
    .B(_1957_),
    .C(_1958_));
 sg13g2_xnor2_1 _6917_ (.Y(\generated._68[3] ),
    .A(\generated._69[3] ),
    .B(_1957_));
 sg13g2_xor2_1 _6918_ (.B(_0913_),
    .A(_0049_),
    .X(_1959_));
 sg13g2_nand2_1 _6919_ (.Y(_1960_),
    .A(_4161_),
    .B(_4159_));
 sg13g2_nor2_1 _6920_ (.A(_1312_),
    .B(_1960_),
    .Y(_1961_));
 sg13g2_nand2_1 _6921_ (.Y(_1962_),
    .A(_4269_),
    .B(_4260_));
 sg13g2_nand2_1 _6922_ (.Y(_1963_),
    .A(_1961_),
    .B(_1962_));
 sg13g2_nor2_1 _6923_ (.A(\generated._568[9] ),
    .B(_4160_),
    .Y(_1964_));
 sg13g2_a21oi_1 _6924_ (.A1(_1964_),
    .A2(_4156_),
    .Y(_1965_),
    .B1(_1294_));
 sg13g2_nand2_1 _6925_ (.Y(_1966_),
    .A(_1963_),
    .B(_1965_));
 sg13g2_buf_8 _6926_ (.A(_1966_),
    .X(_1967_));
 sg13g2_buf_1 _6927_ (.A(_1967_),
    .X(_1968_));
 sg13g2_xnor2_1 _6928_ (.Y(_1969_),
    .A(_0048_),
    .B(net28));
 sg13g2_nor2_1 _6929_ (.A(net59),
    .B(_1969_),
    .Y(_1970_));
 sg13g2_a21oi_1 _6930_ (.A1(net56),
    .A2(_1959_),
    .Y(\generated._691[0] ),
    .B1(_1970_));
 sg13g2_nand2_1 _6931_ (.Y(_1971_),
    .A(_0913_),
    .B(_0049_));
 sg13g2_inv_1 _6932_ (.Y(_1972_),
    .A(\generated._501[1] ));
 sg13g2_xnor2_1 _6933_ (.Y(_1973_),
    .A(net57),
    .B(_0567_));
 sg13g2_inv_1 _6934_ (.Y(_1974_),
    .A(_1973_));
 sg13g2_nand2_2 _6935_ (.Y(_1975_),
    .A(_1974_),
    .B(_0913_));
 sg13g2_xnor2_1 _6936_ (.Y(_1976_),
    .A(_1972_),
    .B(_1975_));
 sg13g2_xnor2_1 _6937_ (.Y(_1977_),
    .A(_1971_),
    .B(_1976_));
 sg13g2_a21oi_1 _6938_ (.A1(_1303_),
    .A2(_4289_),
    .Y(_1978_),
    .B1(_1301_));
 sg13g2_nor2_1 _6939_ (.A(_1978_),
    .B(_1967_),
    .Y(_1979_));
 sg13g2_buf_1 _6940_ (.A(_1979_),
    .X(_1980_));
 sg13g2_xnor2_1 _6941_ (.Y(_1981_),
    .A(\generated._430[11] ),
    .B(net26));
 sg13g2_xnor2_1 _6942_ (.Y(_1982_),
    .A(_0837_),
    .B(_1981_));
 sg13g2_inv_1 _6943_ (.Y(_1983_),
    .A(_0056_));
 sg13g2_nand2_1 _6944_ (.Y(_1984_),
    .A(_1967_),
    .B(_1983_));
 sg13g2_o21ai_1 _6945_ (.B1(_1984_),
    .Y(_1985_),
    .A1(net28),
    .A2(_1982_));
 sg13g2_nand2_1 _6946_ (.Y(_1986_),
    .A(_1964_),
    .B(_4156_));
 sg13g2_nand2_1 _6947_ (.Y(_1987_),
    .A(_1986_),
    .B(_0122_));
 sg13g2_nor3_1 _6948_ (.A(_4162_),
    .B(net95),
    .C(_4155_),
    .Y(_1988_));
 sg13g2_nor2_1 _6949_ (.A(_4156_),
    .B(_4270_),
    .Y(_1989_));
 sg13g2_nand2_1 _6950_ (.Y(_1990_),
    .A(_1989_),
    .B(_1964_));
 sg13g2_nor2_1 _6951_ (.A(_1988_),
    .B(_1990_),
    .Y(_1991_));
 sg13g2_nor2_1 _6952_ (.A(_1987_),
    .B(_1991_),
    .Y(_1992_));
 sg13g2_buf_1 _6953_ (.A(_1992_),
    .X(_1993_));
 sg13g2_nand2_1 _6954_ (.Y(_1994_),
    .A(_1303_),
    .B(_4289_));
 sg13g2_nand2_2 _6955_ (.Y(_1995_),
    .A(_1994_),
    .B(_1300_));
 sg13g2_nand2_1 _6956_ (.Y(_1996_),
    .A(_1993_),
    .B(_1995_));
 sg13g2_inv_1 _6957_ (.Y(_1997_),
    .A(\generated._430[17] ));
 sg13g2_nand2_1 _6958_ (.Y(_1998_),
    .A(_1996_),
    .B(_1997_));
 sg13g2_nand3_1 _6959_ (.B(\generated._430[17] ),
    .C(_1995_),
    .A(_1993_),
    .Y(_1999_));
 sg13g2_nand2_1 _6960_ (.Y(_2000_),
    .A(_1998_),
    .B(_1999_));
 sg13g2_inv_1 _6961_ (.Y(_2001_),
    .A(\generated._430[18] ));
 sg13g2_xnor2_1 _6962_ (.Y(_2002_),
    .A(_2001_),
    .B(net26));
 sg13g2_nor2_1 _6963_ (.A(_2000_),
    .B(_2002_),
    .Y(_2003_));
 sg13g2_nor2_1 _6964_ (.A(_0883_),
    .B(net26),
    .Y(_2004_));
 sg13g2_nand2_1 _6965_ (.Y(_2005_),
    .A(_2004_),
    .B(_0891_));
 sg13g2_buf_8 _6966_ (.A(net26),
    .X(_2006_));
 sg13g2_nand2_1 _6967_ (.Y(_2007_),
    .A(net20),
    .B(\generated._430[16] ));
 sg13g2_nand2_1 _6968_ (.Y(_2008_),
    .A(_2005_),
    .B(_2007_));
 sg13g2_nand2_1 _6969_ (.Y(_2009_),
    .A(_2003_),
    .B(_2008_));
 sg13g2_buf_8 _6970_ (.A(_1996_),
    .X(_2010_));
 sg13g2_nand2_1 _6971_ (.Y(_2011_),
    .A(net25),
    .B(_2001_));
 sg13g2_nand2_1 _6972_ (.Y(_2012_),
    .A(net20),
    .B(\generated._430[18] ));
 sg13g2_nand2_1 _6973_ (.Y(_2013_),
    .A(_2011_),
    .B(_2012_));
 sg13g2_inv_1 _6974_ (.Y(_2014_),
    .A(_1999_));
 sg13g2_nor2_1 _6975_ (.A(_0051_),
    .B(net20),
    .Y(_2015_));
 sg13g2_a21oi_1 _6976_ (.A1(_2013_),
    .A2(_2014_),
    .Y(_2016_),
    .B1(_2015_));
 sg13g2_nand2_1 _6977_ (.Y(_2017_),
    .A(_2009_),
    .B(_2016_));
 sg13g2_nand3_1 _6978_ (.B(_0867_),
    .C(\generated._430[13] ),
    .A(net20),
    .Y(_2018_));
 sg13g2_nand2_1 _6979_ (.Y(_2019_),
    .A(net25),
    .B(_0877_));
 sg13g2_nand2_1 _6980_ (.Y(_2020_),
    .A(_2018_),
    .B(_2019_));
 sg13g2_a21oi_1 _6981_ (.A1(_0850_),
    .A2(_1983_),
    .Y(_2021_),
    .B1(_0859_));
 sg13g2_nor4_1 _6982_ (.A(_0867_),
    .B(_0855_),
    .C(_2021_),
    .D(net20),
    .Y(_2022_));
 sg13g2_nor2_1 _6983_ (.A(_2020_),
    .B(_2022_),
    .Y(_2023_));
 sg13g2_nand2_1 _6984_ (.Y(_2024_),
    .A(net25),
    .B(_0884_));
 sg13g2_nand2_1 _6985_ (.Y(_2025_),
    .A(net26),
    .B(_0883_));
 sg13g2_nand2_1 _6986_ (.Y(_2026_),
    .A(_2024_),
    .B(_2025_));
 sg13g2_xnor2_1 _6987_ (.Y(_2027_),
    .A(_0891_),
    .B(net26));
 sg13g2_nor2_1 _6988_ (.A(_2026_),
    .B(_2027_),
    .Y(_2028_));
 sg13g2_nand2_1 _6989_ (.Y(_2029_),
    .A(_2028_),
    .B(_2003_));
 sg13g2_nor2_1 _6990_ (.A(_2023_),
    .B(_2029_),
    .Y(_2030_));
 sg13g2_nor2_1 _6991_ (.A(_2017_),
    .B(_2030_),
    .Y(_2031_));
 sg13g2_nand2_1 _6992_ (.Y(_2032_),
    .A(net25),
    .B(_0850_));
 sg13g2_nand2_1 _6993_ (.Y(_2033_),
    .A(net26),
    .B(\generated._430[12] ));
 sg13g2_nand2_1 _6994_ (.Y(_2034_),
    .A(_2032_),
    .B(_2033_));
 sg13g2_nand2_1 _6995_ (.Y(_2035_),
    .A(_1981_),
    .B(_2034_));
 sg13g2_xnor2_1 _6996_ (.Y(_2036_),
    .A(_0855_),
    .B(net20));
 sg13g2_xnor2_1 _6997_ (.Y(_2037_),
    .A(_0867_),
    .B(net26));
 sg13g2_nand2_1 _6998_ (.Y(_2038_),
    .A(_2036_),
    .B(_2037_));
 sg13g2_nor2_1 _6999_ (.A(_2035_),
    .B(_2038_),
    .Y(_2039_));
 sg13g2_nand2_1 _7000_ (.Y(_2040_),
    .A(net25),
    .B(_0883_));
 sg13g2_nand2_1 _7001_ (.Y(_2041_),
    .A(_1980_),
    .B(_0884_));
 sg13g2_nand2_1 _7002_ (.Y(_2042_),
    .A(_2040_),
    .B(_2041_));
 sg13g2_nand2_1 _7003_ (.Y(_2043_),
    .A(net25),
    .B(_0891_));
 sg13g2_nand3_1 _7004_ (.B(_0052_),
    .C(_1995_),
    .A(_1993_),
    .Y(_2044_));
 sg13g2_nand2_1 _7005_ (.Y(_2045_),
    .A(_2043_),
    .B(_2044_));
 sg13g2_nand2_1 _7006_ (.Y(_2046_),
    .A(_2042_),
    .B(_2045_));
 sg13g2_xnor2_1 _7007_ (.Y(_2047_),
    .A(_1997_),
    .B(net20));
 sg13g2_nand2_1 _7008_ (.Y(_2048_),
    .A(_2047_),
    .B(_2013_));
 sg13g2_nor2_1 _7009_ (.A(_2046_),
    .B(_2048_),
    .Y(_2049_));
 sg13g2_nand3_1 _7010_ (.B(_2049_),
    .C(_0837_),
    .A(_2039_),
    .Y(_2050_));
 sg13g2_xnor2_1 _7011_ (.Y(_2051_),
    .A(_0050_),
    .B(_2010_));
 sg13g2_nand3_1 _7012_ (.B(_2050_),
    .C(_2051_),
    .A(_2031_),
    .Y(_2052_));
 sg13g2_inv_1 _7013_ (.Y(_2053_),
    .A(_0050_));
 sg13g2_a21oi_1 _7014_ (.A1(_1978_),
    .A2(_2053_),
    .Y(_2054_),
    .B1(_1967_));
 sg13g2_nand2_2 _7015_ (.Y(_2055_),
    .A(_2052_),
    .B(_2054_));
 sg13g2_nand2_1 _7016_ (.Y(_2056_),
    .A(_1967_),
    .B(_0050_));
 sg13g2_nand2_1 _7017_ (.Y(_2057_),
    .A(_2055_),
    .B(_2056_));
 sg13g2_buf_8 _7018_ (.A(_2057_),
    .X(_2058_));
 sg13g2_buf_8 _7019_ (.A(_2058_),
    .X(_2059_));
 sg13g2_xor2_1 _7020_ (.B(net11),
    .A(_1985_),
    .X(_2060_));
 sg13g2_inv_1 _7021_ (.Y(_2061_),
    .A(_2060_));
 sg13g2_a21oi_1 _7022_ (.A1(_2061_),
    .A2(_1969_),
    .Y(_2062_),
    .B1(net72));
 sg13g2_nor2_1 _7023_ (.A(_1969_),
    .B(_2061_),
    .Y(_2063_));
 sg13g2_inv_1 _7024_ (.Y(_2064_),
    .A(_2063_));
 sg13g2_nand2_1 _7025_ (.Y(_2065_),
    .A(_2062_),
    .B(_2064_));
 sg13g2_o21ai_1 _7026_ (.B1(_2065_),
    .Y(\generated._691[1] ),
    .A1(net43),
    .A2(_1977_));
 sg13g2_nand2_1 _7027_ (.Y(_2066_),
    .A(_1981_),
    .B(_0837_));
 sg13g2_o21ai_1 _7028_ (.B1(_2066_),
    .Y(_2067_),
    .A1(_0056_),
    .A2(net20));
 sg13g2_xor2_1 _7029_ (.B(_2067_),
    .A(_2034_),
    .X(_2068_));
 sg13g2_buf_1 _7030_ (.A(_1993_),
    .X(_2069_));
 sg13g2_nor2_1 _7031_ (.A(_0055_),
    .B(net27),
    .Y(_2070_));
 sg13g2_a21oi_1 _7032_ (.A1(_2068_),
    .A2(net27),
    .Y(_2071_),
    .B1(_2070_));
 sg13g2_inv_8 _7033_ (.Y(_2072_),
    .A(_2058_));
 sg13g2_buf_8 _7034_ (.A(_2072_),
    .X(_2073_));
 sg13g2_nor2_1 _7035_ (.A(_2071_),
    .B(net10),
    .Y(_2074_));
 sg13g2_nand2_1 _7036_ (.Y(_2075_),
    .A(net10),
    .B(_2071_));
 sg13g2_nand2b_1 _7037_ (.Y(_2076_),
    .B(_2075_),
    .A_N(_2074_));
 sg13g2_nand2_1 _7038_ (.Y(_2077_),
    .A(_1967_),
    .B(_0905_));
 sg13g2_buf_1 _7039_ (.A(_2077_),
    .X(_2078_));
 sg13g2_nand2_2 _7040_ (.Y(_2079_),
    .A(_2055_),
    .B(net24));
 sg13g2_buf_8 _7041_ (.A(_2079_),
    .X(_2080_));
 sg13g2_a21o_1 _7042_ (.A2(net12),
    .A1(_1985_),
    .B1(_2063_),
    .X(_2081_));
 sg13g2_xor2_1 _7043_ (.B(_2081_),
    .A(_2076_),
    .X(_2082_));
 sg13g2_inv_1 _7044_ (.Y(_2083_),
    .A(_1975_));
 sg13g2_nor2_1 _7045_ (.A(_1972_),
    .B(_2083_),
    .Y(_2084_));
 sg13g2_a21oi_1 _7046_ (.A1(_1976_),
    .A2(_1971_),
    .Y(_2085_),
    .B1(_2084_));
 sg13g2_inv_1 _7047_ (.Y(_2086_),
    .A(_2085_));
 sg13g2_inv_1 _7048_ (.Y(_2087_),
    .A(\generated._501[2] ));
 sg13g2_nor2_1 _7049_ (.A(net42),
    .B(_0569_),
    .Y(_2088_));
 sg13g2_a21oi_1 _7050_ (.A1(net55),
    .A2(net42),
    .Y(_2089_),
    .B1(_2088_));
 sg13g2_nor2_1 _7051_ (.A(_2087_),
    .B(_2089_),
    .Y(_2090_));
 sg13g2_nand2_1 _7052_ (.Y(_2091_),
    .A(_2089_),
    .B(_2087_));
 sg13g2_nor2b_1 _7053_ (.A(_2090_),
    .B_N(_2091_),
    .Y(_2092_));
 sg13g2_nand2_1 _7054_ (.Y(_2093_),
    .A(_2086_),
    .B(_2092_));
 sg13g2_nand2b_1 _7055_ (.Y(_2094_),
    .B(_2085_),
    .A_N(_2092_));
 sg13g2_nand3_1 _7056_ (.B(net59),
    .C(_2094_),
    .A(_2093_),
    .Y(_2095_));
 sg13g2_o21ai_1 _7057_ (.B1(_2095_),
    .Y(\generated._691[2] ),
    .A1(net56),
    .A2(_2082_));
 sg13g2_inv_1 _7058_ (.Y(_2096_),
    .A(_2036_));
 sg13g2_a22oi_1 _7059_ (.Y(_2097_),
    .B1(_2034_),
    .B2(_2067_),
    .A2(net25),
    .A1(_0859_));
 sg13g2_nor2_1 _7060_ (.A(_2096_),
    .B(_2097_),
    .Y(_2098_));
 sg13g2_a21o_1 _7061_ (.A2(_2096_),
    .A1(_2097_),
    .B1(net28),
    .X(_2099_));
 sg13g2_nand2b_1 _7062_ (.Y(_2100_),
    .B(net28),
    .A_N(_0057_));
 sg13g2_o21ai_1 _7063_ (.B1(_2100_),
    .Y(_2101_),
    .A1(_2098_),
    .A2(_2099_));
 sg13g2_xnor2_1 _7064_ (.Y(_2102_),
    .A(net11),
    .B(_2101_));
 sg13g2_a21o_1 _7065_ (.A2(_2075_),
    .A1(_2081_),
    .B1(_2074_),
    .X(_2103_));
 sg13g2_nor2_1 _7066_ (.A(_2102_),
    .B(_2103_),
    .Y(_2104_));
 sg13g2_nand2_1 _7067_ (.Y(_2105_),
    .A(_2103_),
    .B(_2102_));
 sg13g2_nand2_1 _7068_ (.Y(_2106_),
    .A(_2105_),
    .B(net38));
 sg13g2_inv_1 _7069_ (.Y(_2107_),
    .A(\generated._501[3] ));
 sg13g2_xnor2_1 _7070_ (.Y(_2108_),
    .A(_2107_),
    .B(_1975_));
 sg13g2_inv_1 _7071_ (.Y(_2109_),
    .A(_2108_));
 sg13g2_o21ai_1 _7072_ (.B1(_2091_),
    .Y(_2110_),
    .A1(_2090_),
    .A2(_2086_));
 sg13g2_nor2_1 _7073_ (.A(_2109_),
    .B(_2110_),
    .Y(_2111_));
 sg13g2_nand2_1 _7074_ (.Y(_2112_),
    .A(_2110_),
    .B(_2109_));
 sg13g2_nand3b_1 _7075_ (.B(net72),
    .C(_2112_),
    .Y(_2113_),
    .A_N(_2111_));
 sg13g2_o21ai_1 _7076_ (.B1(_2113_),
    .Y(\generated._691[3] ),
    .A1(_2104_),
    .A2(_2106_));
 sg13g2_nor2_1 _7077_ (.A(_0855_),
    .B(net25),
    .Y(_2114_));
 sg13g2_nor2_1 _7078_ (.A(_2114_),
    .B(_2098_),
    .Y(_2115_));
 sg13g2_xor2_1 _7079_ (.B(_2115_),
    .A(_2037_),
    .X(_2116_));
 sg13g2_nor2_1 _7080_ (.A(net28),
    .B(_2116_),
    .Y(_2117_));
 sg13g2_a21oi_1 _7081_ (.A1(_0877_),
    .A2(net28),
    .Y(_2118_),
    .B1(_2117_));
 sg13g2_nor2_1 _7082_ (.A(net10),
    .B(_2118_),
    .Y(_2119_));
 sg13g2_inv_1 _7083_ (.Y(_2120_),
    .A(_2119_));
 sg13g2_nand2_1 _7084_ (.Y(_2121_),
    .A(_2118_),
    .B(net10));
 sg13g2_nand2_1 _7085_ (.Y(_2122_),
    .A(_2120_),
    .B(_2121_));
 sg13g2_nand2_1 _7086_ (.Y(_2123_),
    .A(_2101_),
    .B(net10));
 sg13g2_nand2_1 _7087_ (.Y(_2124_),
    .A(_2105_),
    .B(_2123_));
 sg13g2_xor2_1 _7088_ (.B(_2124_),
    .A(_2122_),
    .X(_2125_));
 sg13g2_a21oi_1 _7089_ (.A1(\generated._501[3] ),
    .A2(_1975_),
    .Y(_2126_),
    .B1(_2111_));
 sg13g2_inv_1 _7090_ (.Y(_2127_),
    .A(_2126_));
 sg13g2_nor2_1 _7091_ (.A(net82),
    .B(_0567_),
    .Y(_2128_));
 sg13g2_a21oi_1 _7092_ (.A1(_0914_),
    .A2(net82),
    .Y(_2129_),
    .B1(_2128_));
 sg13g2_nor2_1 _7093_ (.A(\generated._501[4] ),
    .B(_2129_),
    .Y(_2130_));
 sg13g2_and2_1 _7094_ (.A(_2129_),
    .B(\generated._501[4] ),
    .X(_2131_));
 sg13g2_nor2_1 _7095_ (.A(_2130_),
    .B(_2131_),
    .Y(_2132_));
 sg13g2_a21oi_1 _7096_ (.A1(_2127_),
    .A2(_2132_),
    .Y(_2133_),
    .B1(_0584_));
 sg13g2_o21ai_1 _7097_ (.B1(_2133_),
    .Y(_2134_),
    .A1(_2127_),
    .A2(_2132_));
 sg13g2_o21ai_1 _7098_ (.B1(_2134_),
    .Y(\generated._691[4] ),
    .A1(net56),
    .A2(_2125_));
 sg13g2_inv_1 _7099_ (.Y(_2135_),
    .A(_2115_));
 sg13g2_inv_1 _7100_ (.Y(_2136_),
    .A(_2019_));
 sg13g2_a21oi_1 _7101_ (.A1(_2135_),
    .A2(_2037_),
    .Y(_2137_),
    .B1(_2136_));
 sg13g2_xnor2_1 _7102_ (.Y(_2138_),
    .A(_2042_),
    .B(_2137_));
 sg13g2_nor2_1 _7103_ (.A(_0883_),
    .B(net27),
    .Y(_2139_));
 sg13g2_a21oi_1 _7104_ (.A1(_2138_),
    .A2(net27),
    .Y(_2140_),
    .B1(_2139_));
 sg13g2_xnor2_1 _7105_ (.Y(_2141_),
    .A(net11),
    .B(_2140_));
 sg13g2_inv_1 _7106_ (.Y(_2142_),
    .A(_2141_));
 sg13g2_a21o_1 _7107_ (.A2(_2121_),
    .A1(_2124_),
    .B1(_2119_),
    .X(_2143_));
 sg13g2_inv_1 _7108_ (.Y(_2144_),
    .A(_2143_));
 sg13g2_nor2_1 _7109_ (.A(_2142_),
    .B(_2144_),
    .Y(_2145_));
 sg13g2_o21ai_1 _7110_ (.B1(net38),
    .Y(_2146_),
    .A1(_2141_),
    .A2(_2143_));
 sg13g2_xnor2_1 _7111_ (.Y(_2147_),
    .A(net70),
    .B(net82));
 sg13g2_inv_1 _7112_ (.Y(_2148_),
    .A(_2147_));
 sg13g2_nor2_1 _7113_ (.A(\generated._501[5] ),
    .B(_2148_),
    .Y(_2149_));
 sg13g2_nand2_1 _7114_ (.Y(_2150_),
    .A(_2148_),
    .B(\generated._501[5] ));
 sg13g2_nor2b_1 _7115_ (.A(_2149_),
    .B_N(_2150_),
    .Y(_2151_));
 sg13g2_inv_1 _7116_ (.Y(_2152_),
    .A(_2151_));
 sg13g2_inv_1 _7117_ (.Y(_2153_),
    .A(_2130_));
 sg13g2_a21oi_1 _7118_ (.A1(_2127_),
    .A2(_2153_),
    .Y(_2154_),
    .B1(_2131_));
 sg13g2_nor2_1 _7119_ (.A(_2152_),
    .B(_2154_),
    .Y(_2155_));
 sg13g2_a21oi_1 _7120_ (.A1(_2154_),
    .A2(_2152_),
    .Y(_2156_),
    .B1(_0584_));
 sg13g2_nand2b_1 _7121_ (.Y(_2157_),
    .B(_2156_),
    .A_N(_2155_));
 sg13g2_o21ai_1 _7122_ (.B1(_2157_),
    .Y(\generated._691[5] ),
    .A1(_2145_),
    .A2(_2146_));
 sg13g2_inv_1 _7123_ (.Y(_2158_),
    .A(\generated._501[6] ));
 sg13g2_nor2_1 _7124_ (.A(_2158_),
    .B(_1973_),
    .Y(_2159_));
 sg13g2_inv_1 _7125_ (.Y(_2160_),
    .A(_2159_));
 sg13g2_nand2_1 _7126_ (.Y(_2161_),
    .A(_1973_),
    .B(_2158_));
 sg13g2_nand2_1 _7127_ (.Y(_2162_),
    .A(_2160_),
    .B(_2161_));
 sg13g2_inv_1 _7128_ (.Y(_2163_),
    .A(_2162_));
 sg13g2_o21ai_1 _7129_ (.B1(_2150_),
    .Y(_2164_),
    .A1(_2149_),
    .A2(_2154_));
 sg13g2_xnor2_1 _7130_ (.Y(_2165_),
    .A(_2163_),
    .B(_2164_));
 sg13g2_nor2_1 _7131_ (.A(net10),
    .B(_2140_),
    .Y(_2166_));
 sg13g2_nand2_1 _7132_ (.Y(_2167_),
    .A(_2037_),
    .B(_2042_));
 sg13g2_nor2_1 _7133_ (.A(_2004_),
    .B(_2136_),
    .Y(_2168_));
 sg13g2_o21ai_1 _7134_ (.B1(_2168_),
    .Y(_2169_),
    .A1(_2167_),
    .A2(_2115_));
 sg13g2_nand2b_1 _7135_ (.Y(_2170_),
    .B(_2045_),
    .A_N(_2169_));
 sg13g2_nand2_1 _7136_ (.Y(_2171_),
    .A(_2169_),
    .B(_2027_));
 sg13g2_nand3_1 _7137_ (.B(net27),
    .C(_2171_),
    .A(_2170_),
    .Y(_2172_));
 sg13g2_o21ai_1 _7138_ (.B1(_2172_),
    .Y(_2173_),
    .A1(_0891_),
    .A2(_2069_));
 sg13g2_nor2_1 _7139_ (.A(net11),
    .B(_2173_),
    .Y(_2174_));
 sg13g2_nand2_1 _7140_ (.Y(_2175_),
    .A(_2173_),
    .B(net11));
 sg13g2_inv_1 _7141_ (.Y(_2176_),
    .A(_2175_));
 sg13g2_nor2_1 _7142_ (.A(_2174_),
    .B(_2176_),
    .Y(_2177_));
 sg13g2_o21ai_1 _7143_ (.B1(_2177_),
    .Y(_2178_),
    .A1(_2166_),
    .A2(_2145_));
 sg13g2_nor2_1 _7144_ (.A(_2166_),
    .B(_2145_),
    .Y(_2179_));
 sg13g2_nand2b_1 _7145_ (.Y(_2180_),
    .B(_2179_),
    .A_N(_2177_));
 sg13g2_nand3_1 _7146_ (.B(_2180_),
    .C(net38),
    .A(_2178_),
    .Y(_2181_));
 sg13g2_o21ai_1 _7147_ (.B1(_2181_),
    .Y(\generated._691[6] ),
    .A1(net43),
    .A2(_2165_));
 sg13g2_inv_1 _7148_ (.Y(_2182_),
    .A(_2174_));
 sg13g2_a21oi_1 _7149_ (.A1(_2179_),
    .A2(_2182_),
    .Y(_2183_),
    .B1(_2176_));
 sg13g2_inv_1 _7150_ (.Y(_2184_),
    .A(_2008_));
 sg13g2_o21ai_1 _7151_ (.B1(_2184_),
    .Y(_2185_),
    .A1(_2046_),
    .A2(_2137_));
 sg13g2_nand2b_1 _7152_ (.Y(_2186_),
    .B(_2000_),
    .A_N(_2185_));
 sg13g2_a21oi_1 _7153_ (.A1(_2185_),
    .A2(_2047_),
    .Y(_2187_),
    .B1(net28));
 sg13g2_a22oi_1 _7154_ (.Y(_2188_),
    .B1(_2186_),
    .B2(_2187_),
    .A2(net28),
    .A1(_0899_));
 sg13g2_xor2_1 _7155_ (.B(_2188_),
    .A(net12),
    .X(_2189_));
 sg13g2_inv_1 _7156_ (.Y(_2190_),
    .A(_2189_));
 sg13g2_nand2b_1 _7157_ (.Y(_2191_),
    .B(_2190_),
    .A_N(_2183_));
 sg13g2_nand2_1 _7158_ (.Y(_2192_),
    .A(_2183_),
    .B(_2189_));
 sg13g2_nand3_1 _7159_ (.B(net38),
    .C(_2192_),
    .A(_2191_),
    .Y(_2193_));
 sg13g2_nand2_1 _7160_ (.Y(_2194_),
    .A(_2160_),
    .B(_2150_));
 sg13g2_o21ai_1 _7161_ (.B1(_2161_),
    .Y(_2195_),
    .A1(_2194_),
    .A2(_2155_));
 sg13g2_nor2_1 _7162_ (.A(\generated._501[7] ),
    .B(net42),
    .Y(_2196_));
 sg13g2_nor2b_1 _7163_ (.A(net82),
    .B_N(\generated._501[7] ),
    .Y(_2197_));
 sg13g2_nor2_1 _7164_ (.A(_2196_),
    .B(_2197_),
    .Y(_2198_));
 sg13g2_nand2b_1 _7165_ (.Y(_2199_),
    .B(_2198_),
    .A_N(_2195_));
 sg13g2_nand2b_1 _7166_ (.Y(_2200_),
    .B(_2195_),
    .A_N(_2198_));
 sg13g2_nand3_1 _7167_ (.B(_2200_),
    .C(net59),
    .A(_2199_),
    .Y(_2201_));
 sg13g2_nand2_1 _7168_ (.Y(\generated._691[7] ),
    .A(_2193_),
    .B(_2201_));
 sg13g2_a21oi_1 _7169_ (.A1(_2185_),
    .A2(_1998_),
    .Y(_2202_),
    .B1(_2014_));
 sg13g2_xnor2_1 _7170_ (.Y(_2203_),
    .A(_2002_),
    .B(_2202_));
 sg13g2_nor2_1 _7171_ (.A(_0906_),
    .B(net27),
    .Y(_2204_));
 sg13g2_a21oi_1 _7172_ (.A1(_2203_),
    .A2(net27),
    .Y(_2205_),
    .B1(_2204_));
 sg13g2_xnor2_1 _7173_ (.Y(_2206_),
    .A(net10),
    .B(_2205_));
 sg13g2_nor2_1 _7174_ (.A(net11),
    .B(_2188_),
    .Y(_2207_));
 sg13g2_a21oi_1 _7175_ (.A1(_2189_),
    .A2(_2174_),
    .Y(_2208_),
    .B1(_2207_));
 sg13g2_o21ai_1 _7176_ (.B1(_2208_),
    .Y(_2209_),
    .A1(_2190_),
    .A2(_2178_));
 sg13g2_xnor2_1 _7177_ (.Y(_2210_),
    .A(_2206_),
    .B(_2209_));
 sg13g2_xnor2_1 _7178_ (.Y(_2211_),
    .A(\generated._501[8] ),
    .B(net82));
 sg13g2_nand2_1 _7179_ (.Y(_2212_),
    .A(_2164_),
    .B(_2163_));
 sg13g2_nor2_1 _7180_ (.A(_2197_),
    .B(_2159_),
    .Y(_2213_));
 sg13g2_a21oi_1 _7181_ (.A1(_2212_),
    .A2(_2213_),
    .Y(_2214_),
    .B1(_2196_));
 sg13g2_a21oi_1 _7182_ (.A1(_2214_),
    .A2(_2211_),
    .Y(_2215_),
    .B1(_0584_));
 sg13g2_o21ai_1 _7183_ (.B1(_2215_),
    .Y(_2216_),
    .A1(_2211_),
    .A2(_2214_));
 sg13g2_o21ai_1 _7184_ (.B1(_2216_),
    .Y(\generated._691[8] ),
    .A1(net56),
    .A2(_2210_));
 sg13g2_a21oi_1 _7185_ (.A1(_2031_),
    .A2(_2050_),
    .Y(_2217_),
    .B1(_2051_));
 sg13g2_nand2_1 _7186_ (.Y(_2218_),
    .A(_2052_),
    .B(net27));
 sg13g2_o21ai_1 _7187_ (.B1(_2056_),
    .Y(_2219_),
    .A1(_2217_),
    .A2(_2218_));
 sg13g2_xnor2_1 _7188_ (.Y(_2220_),
    .A(net10),
    .B(_2219_));
 sg13g2_inv_1 _7189_ (.Y(_2221_),
    .A(_2206_));
 sg13g2_o21ai_1 _7190_ (.B1(_2205_),
    .Y(_2222_),
    .A1(net12),
    .A2(_2207_));
 sg13g2_o21ai_1 _7191_ (.B1(_2222_),
    .Y(_2223_),
    .A1(_2221_),
    .A2(_2192_));
 sg13g2_xor2_1 _7192_ (.B(_2223_),
    .A(_2220_),
    .X(_2224_));
 sg13g2_nand2b_1 _7193_ (.Y(_2225_),
    .B(_2211_),
    .A_N(_2199_));
 sg13g2_o21ai_1 _7194_ (.B1(net42),
    .Y(_2226_),
    .A1(\generated._501[8] ),
    .A2(\generated._501[7] ));
 sg13g2_nand3_1 _7195_ (.B(net59),
    .C(_2226_),
    .A(_2225_),
    .Y(_2227_));
 sg13g2_o21ai_1 _7196_ (.B1(_2227_),
    .Y(\generated._691[9] ),
    .A1(net56),
    .A2(_2224_));
 sg13g2_nor2_1 _7197_ (.A(net95),
    .B(_4260_),
    .Y(_2228_));
 sg13g2_nand2_1 _7198_ (.Y(_2229_),
    .A(_2228_),
    .B(_1284_));
 sg13g2_nor2_1 _7199_ (.A(_4270_),
    .B(_1988_),
    .Y(_2230_));
 sg13g2_a21oi_2 _7200_ (.B1(_2230_),
    .Y(_2231_),
    .A2(_4272_),
    .A1(_4260_));
 sg13g2_xor2_1 _7201_ (.B(_2231_),
    .A(_2229_),
    .X(_2232_));
 sg13g2_buf_1 _7202_ (.A(_2232_),
    .X(_2233_));
 sg13g2_inv_1 _7203_ (.Y(_2234_),
    .A(net31));
 sg13g2_nor2_1 _7204_ (.A(_0589_),
    .B(_0586_),
    .Y(_2235_));
 sg13g2_nand3_1 _7205_ (.B(_0606_),
    .C(_0633_),
    .A(_2235_),
    .Y(_2236_));
 sg13g2_nand3b_1 _7206_ (.B(_0645_),
    .C(_0663_),
    .Y(_2237_),
    .A_N(_2236_));
 sg13g2_xnor2_1 _7207_ (.Y(_2238_),
    .A(_0685_),
    .B(_2237_));
 sg13g2_nand2_2 _7208_ (.Y(_2239_),
    .A(net12),
    .B(_2238_));
 sg13g2_buf_8 _7209_ (.A(_2055_),
    .X(_2240_));
 sg13g2_nand3_1 _7210_ (.B(_0078_),
    .C(net24),
    .A(net13),
    .Y(_2241_));
 sg13g2_buf_2 _7211_ (.A(_2241_),
    .X(_2242_));
 sg13g2_nand2_1 _7212_ (.Y(_2243_),
    .A(_2239_),
    .B(_2242_));
 sg13g2_nor2_1 _7213_ (.A(_2234_),
    .B(_2243_),
    .Y(_2244_));
 sg13g2_xor2_1 _7214_ (.B(_4164_),
    .A(_1284_),
    .X(_2245_));
 sg13g2_xor2_1 _7215_ (.B(_2245_),
    .A(_2228_),
    .X(_2246_));
 sg13g2_buf_1 _7216_ (.A(_2246_),
    .X(_2247_));
 sg13g2_inv_1 _7217_ (.Y(_2248_),
    .A(net37));
 sg13g2_inv_1 _7218_ (.Y(_2249_),
    .A(_0067_));
 sg13g2_nor3_1 _7219_ (.A(_0589_),
    .B(\generated._508[1] ),
    .C(_2249_),
    .Y(_2250_));
 sg13g2_nand3_1 _7220_ (.B(_0633_),
    .C(_0645_),
    .A(_2250_),
    .Y(_2251_));
 sg13g2_xnor2_1 _7221_ (.Y(_2252_),
    .A(\generated._508[4] ),
    .B(_2251_));
 sg13g2_nand2_1 _7222_ (.Y(_2253_),
    .A(net12),
    .B(_2252_));
 sg13g2_nand3_1 _7223_ (.B(_0075_),
    .C(net24),
    .A(net13),
    .Y(_2254_));
 sg13g2_nand2_1 _7224_ (.Y(_2255_),
    .A(_2253_),
    .B(_2254_));
 sg13g2_buf_2 _7225_ (.A(_2255_),
    .X(_2256_));
 sg13g2_nor2_1 _7226_ (.A(_2248_),
    .B(_2256_),
    .Y(_2257_));
 sg13g2_nand2_1 _7227_ (.Y(_2258_),
    .A(_2244_),
    .B(_2257_));
 sg13g2_nand3_1 _7228_ (.B(_2242_),
    .C(net37),
    .A(_2239_),
    .Y(_2259_));
 sg13g2_nand3_1 _7229_ (.B(_2254_),
    .C(net31),
    .A(_2253_),
    .Y(_2260_));
 sg13g2_nand2_1 _7230_ (.Y(_2261_),
    .A(_2259_),
    .B(_2260_));
 sg13g2_nand2_1 _7231_ (.Y(_2262_),
    .A(_2258_),
    .B(_2261_));
 sg13g2_xnor2_1 _7232_ (.Y(_2263_),
    .A(_1290_),
    .B(_2230_));
 sg13g2_inv_1 _7233_ (.Y(_2264_),
    .A(_2231_));
 sg13g2_nand2b_1 _7234_ (.Y(_2265_),
    .B(_2264_),
    .A_N(_2229_));
 sg13g2_xor2_1 _7235_ (.B(_2265_),
    .A(_2263_),
    .X(_2266_));
 sg13g2_inv_1 _7236_ (.Y(_2267_),
    .A(_2266_));
 sg13g2_xnor2_1 _7237_ (.Y(_2268_),
    .A(\generated._508[3] ),
    .B(_2236_));
 sg13g2_nand2_1 _7238_ (.Y(_2269_),
    .A(net12),
    .B(_2268_));
 sg13g2_nand3_1 _7239_ (.B(_0072_),
    .C(net24),
    .A(net13),
    .Y(_2270_));
 sg13g2_buf_1 _7240_ (.A(_2270_),
    .X(_2271_));
 sg13g2_nand2_2 _7241_ (.Y(_2272_),
    .A(_2269_),
    .B(_2271_));
 sg13g2_nor2_1 _7242_ (.A(_2267_),
    .B(_2272_),
    .Y(_2273_));
 sg13g2_nand2_1 _7243_ (.Y(_2274_),
    .A(_2262_),
    .B(_2273_));
 sg13g2_nand3_1 _7244_ (.B(_2254_),
    .C(net37),
    .A(_2253_),
    .Y(_2275_));
 sg13g2_nand3_1 _7245_ (.B(_2271_),
    .C(net31),
    .A(_2269_),
    .Y(_2276_));
 sg13g2_nand2_1 _7246_ (.Y(_2277_),
    .A(_2275_),
    .B(_2276_));
 sg13g2_buf_1 _7247_ (.A(_2267_),
    .X(_2278_));
 sg13g2_xnor2_1 _7248_ (.Y(_2279_),
    .A(_0633_),
    .B(_2250_));
 sg13g2_nand2_1 _7249_ (.Y(_2280_),
    .A(net12),
    .B(_2279_));
 sg13g2_nand3_1 _7250_ (.B(_0069_),
    .C(net24),
    .A(net13),
    .Y(_2281_));
 sg13g2_nand2_2 _7251_ (.Y(_2282_),
    .A(_2280_),
    .B(_2281_));
 sg13g2_nor2_1 _7252_ (.A(net19),
    .B(_2282_),
    .Y(_2283_));
 sg13g2_nand3_1 _7253_ (.B(_2271_),
    .C(net37),
    .A(_2269_),
    .Y(_2284_));
 sg13g2_nor2_1 _7254_ (.A(_2260_),
    .B(_2284_),
    .Y(_2285_));
 sg13g2_a21oi_1 _7255_ (.A1(_2277_),
    .A2(_2283_),
    .Y(_2286_),
    .B1(_2285_));
 sg13g2_inv_1 _7256_ (.Y(_2287_),
    .A(_2273_));
 sg13g2_nand3_1 _7257_ (.B(_2261_),
    .C(_2287_),
    .A(_2258_),
    .Y(_2288_));
 sg13g2_nand3_1 _7258_ (.B(_2286_),
    .C(_2288_),
    .A(_2274_),
    .Y(_2289_));
 sg13g2_inv_1 _7259_ (.Y(_2290_),
    .A(_2230_));
 sg13g2_a21oi_1 _7260_ (.A1(_2290_),
    .A2(_4265_),
    .Y(_2291_),
    .B1(_4160_));
 sg13g2_xnor2_1 _7261_ (.Y(_2292_),
    .A(_0122_),
    .B(_2291_));
 sg13g2_inv_1 _7262_ (.Y(_2293_),
    .A(_2292_));
 sg13g2_o21ai_1 _7263_ (.B1(_0117_),
    .Y(_2294_),
    .A1(_1312_),
    .A2(_1988_));
 sg13g2_xnor2_1 _7264_ (.Y(_2295_),
    .A(_4159_),
    .B(_2294_));
 sg13g2_inv_1 _7265_ (.Y(_2296_),
    .A(_2295_));
 sg13g2_nor2_1 _7266_ (.A(_2263_),
    .B(_2265_),
    .Y(_2297_));
 sg13g2_inv_1 _7267_ (.Y(_2298_),
    .A(_2297_));
 sg13g2_nor2_1 _7268_ (.A(_2296_),
    .B(_2298_),
    .Y(_2299_));
 sg13g2_inv_1 _7269_ (.Y(_2300_),
    .A(_2299_));
 sg13g2_nor3_1 _7270_ (.A(_1967_),
    .B(_2293_),
    .C(_2300_),
    .Y(_2301_));
 sg13g2_nor2_1 _7271_ (.A(_2293_),
    .B(_2300_),
    .Y(_2302_));
 sg13g2_nor2_1 _7272_ (.A(_1993_),
    .B(_2302_),
    .Y(_2303_));
 sg13g2_buf_1 _7273_ (.A(_2303_),
    .X(_2304_));
 sg13g2_nor2_1 _7274_ (.A(_2301_),
    .B(net14),
    .Y(_2305_));
 sg13g2_buf_2 _7275_ (.A(_2305_),
    .X(_2306_));
 sg13g2_xnor2_1 _7276_ (.Y(_2307_),
    .A(_0589_),
    .B(_0586_));
 sg13g2_nand2_1 _7277_ (.Y(_2308_),
    .A(net12),
    .B(_2307_));
 sg13g2_nand3_1 _7278_ (.B(_0623_),
    .C(net24),
    .A(net13),
    .Y(_2309_));
 sg13g2_nand2_1 _7279_ (.Y(_2310_),
    .A(_2308_),
    .B(_2309_));
 sg13g2_buf_2 _7280_ (.A(_2310_),
    .X(_2311_));
 sg13g2_nor2_2 _7281_ (.A(_2306_),
    .B(_2311_),
    .Y(_2312_));
 sg13g2_xnor2_1 _7282_ (.Y(_2313_),
    .A(_2296_),
    .B(_2297_));
 sg13g2_buf_2 _7283_ (.A(_2313_),
    .X(_2314_));
 sg13g2_inv_2 _7284_ (.Y(_2315_),
    .A(_2314_));
 sg13g2_nor2_1 _7285_ (.A(_2315_),
    .B(_2282_),
    .Y(_2316_));
 sg13g2_xnor2_1 _7286_ (.Y(_2317_),
    .A(_2293_),
    .B(_2299_));
 sg13g2_inv_2 _7287_ (.Y(_2318_),
    .A(_2317_));
 sg13g2_xnor2_1 _7288_ (.Y(_2319_),
    .A(_0606_),
    .B(_2235_));
 sg13g2_nand2_1 _7289_ (.Y(_2320_),
    .A(_2080_),
    .B(_2319_));
 sg13g2_nand3_1 _7290_ (.B(_0068_),
    .C(net24),
    .A(net13),
    .Y(_2321_));
 sg13g2_nand2_1 _7291_ (.Y(_2322_),
    .A(_2320_),
    .B(_2321_));
 sg13g2_buf_2 _7292_ (.A(_2322_),
    .X(_2323_));
 sg13g2_nor2_1 _7293_ (.A(_2318_),
    .B(_2323_),
    .Y(_2324_));
 sg13g2_nand2b_1 _7294_ (.Y(_2325_),
    .B(_2324_),
    .A_N(_2316_));
 sg13g2_inv_1 _7295_ (.Y(_2326_),
    .A(_2324_));
 sg13g2_nand2_1 _7296_ (.Y(_2327_),
    .A(_2326_),
    .B(_2316_));
 sg13g2_nand2_1 _7297_ (.Y(_2328_),
    .A(_2325_),
    .B(_2327_));
 sg13g2_nand2b_1 _7298_ (.Y(_2329_),
    .B(_2328_),
    .A_N(_2312_));
 sg13g2_nand3_1 _7299_ (.B(_2327_),
    .C(_2312_),
    .A(_2325_),
    .Y(_2330_));
 sg13g2_nand2_1 _7300_ (.Y(_2331_),
    .A(_2329_),
    .B(_2330_));
 sg13g2_a21oi_1 _7301_ (.A1(_2274_),
    .A2(_2288_),
    .Y(_2332_),
    .B1(_2286_));
 sg13g2_a21oi_1 _7302_ (.A1(_2289_),
    .A2(_2331_),
    .Y(_2333_),
    .B1(_2332_));
 sg13g2_nand3_1 _7303_ (.B(_2242_),
    .C(net31),
    .A(_2239_),
    .Y(_2334_));
 sg13g2_nor2_1 _7304_ (.A(_2334_),
    .B(_2275_),
    .Y(_2335_));
 sg13g2_a21oi_1 _7305_ (.A1(_2261_),
    .A2(_2273_),
    .Y(_2336_),
    .B1(_2335_));
 sg13g2_inv_1 _7306_ (.Y(_2337_),
    .A(\generated._508[6] ));
 sg13g2_nor3_1 _7307_ (.A(\generated._508[4] ),
    .B(_0685_),
    .C(_2251_),
    .Y(_2338_));
 sg13g2_xnor2_1 _7308_ (.Y(_2339_),
    .A(_2337_),
    .B(_2338_));
 sg13g2_nand2_2 _7309_ (.Y(_2340_),
    .A(_2079_),
    .B(_2339_));
 sg13g2_nand3_1 _7310_ (.B(_0720_),
    .C(_2078_),
    .A(_2240_),
    .Y(_2341_));
 sg13g2_buf_8 _7311_ (.A(_2341_),
    .X(_2342_));
 sg13g2_nand2_1 _7312_ (.Y(_2343_),
    .A(_2340_),
    .B(_2342_));
 sg13g2_buf_2 _7313_ (.A(_2343_),
    .X(_2344_));
 sg13g2_nor2_1 _7314_ (.A(_2248_),
    .B(_2344_),
    .Y(_2345_));
 sg13g2_nand2_1 _7315_ (.Y(_2346_),
    .A(_2244_),
    .B(_2345_));
 sg13g2_nand3_1 _7316_ (.B(_2342_),
    .C(net37),
    .A(_2340_),
    .Y(_2347_));
 sg13g2_nand2_1 _7317_ (.Y(_2348_),
    .A(_2334_),
    .B(_2347_));
 sg13g2_nand2_1 _7318_ (.Y(_2349_),
    .A(_2346_),
    .B(_2348_));
 sg13g2_nor2_1 _7319_ (.A(_2267_),
    .B(_2256_),
    .Y(_2350_));
 sg13g2_nand2_1 _7320_ (.Y(_2351_),
    .A(_2349_),
    .B(_2350_));
 sg13g2_inv_1 _7321_ (.Y(_2352_),
    .A(_2350_));
 sg13g2_nand3_1 _7322_ (.B(_2348_),
    .C(_2352_),
    .A(_2346_),
    .Y(_2353_));
 sg13g2_nand2_1 _7323_ (.Y(_2354_),
    .A(_2351_),
    .B(_2353_));
 sg13g2_nand2b_1 _7324_ (.Y(_2355_),
    .B(_2354_),
    .A_N(_2336_));
 sg13g2_nand3_1 _7325_ (.B(_2336_),
    .C(_2353_),
    .A(_2351_),
    .Y(_2356_));
 sg13g2_nand2_1 _7326_ (.Y(_2357_),
    .A(_2355_),
    .B(_2356_));
 sg13g2_nor2_1 _7327_ (.A(_2315_),
    .B(_2272_),
    .Y(_2358_));
 sg13g2_nor2_1 _7328_ (.A(_2318_),
    .B(_2282_),
    .Y(_2359_));
 sg13g2_nand2b_1 _7329_ (.Y(_2360_),
    .B(_2359_),
    .A_N(_2358_));
 sg13g2_nand2b_1 _7330_ (.Y(_2361_),
    .B(_2358_),
    .A_N(_2359_));
 sg13g2_nand2_1 _7331_ (.Y(_2362_),
    .A(_2360_),
    .B(_2361_));
 sg13g2_nor2_1 _7332_ (.A(_2306_),
    .B(_2323_),
    .Y(_2363_));
 sg13g2_inv_1 _7333_ (.Y(_2364_),
    .A(_2363_));
 sg13g2_nand2_1 _7334_ (.Y(_2365_),
    .A(_2362_),
    .B(_2364_));
 sg13g2_nand3_1 _7335_ (.B(_2361_),
    .C(_2363_),
    .A(_2360_),
    .Y(_2366_));
 sg13g2_nand2_1 _7336_ (.Y(_2367_),
    .A(_2365_),
    .B(_2366_));
 sg13g2_nand2_1 _7337_ (.Y(_2368_),
    .A(_2357_),
    .B(_2367_));
 sg13g2_nand2_1 _7338_ (.Y(_2369_),
    .A(_2362_),
    .B(_2363_));
 sg13g2_nand3_1 _7339_ (.B(_2361_),
    .C(_2364_),
    .A(_2360_),
    .Y(_2370_));
 sg13g2_nand2_1 _7340_ (.Y(_2371_),
    .A(_2369_),
    .B(_2370_));
 sg13g2_nand3_1 _7341_ (.B(_2356_),
    .C(_2371_),
    .A(_2355_),
    .Y(_2372_));
 sg13g2_nand2_1 _7342_ (.Y(_2373_),
    .A(_2368_),
    .B(_2372_));
 sg13g2_nand2b_1 _7343_ (.Y(_2374_),
    .B(_2373_),
    .A_N(_2333_));
 sg13g2_nand3_1 _7344_ (.B(_2333_),
    .C(_2372_),
    .A(_2368_),
    .Y(_2375_));
 sg13g2_nand2_1 _7345_ (.Y(_2376_),
    .A(_2374_),
    .B(_2375_));
 sg13g2_nor2_1 _7346_ (.A(net14),
    .B(_2311_),
    .Y(_2377_));
 sg13g2_nor2_1 _7347_ (.A(_2315_),
    .B(_2323_),
    .Y(_2378_));
 sg13g2_a22oi_1 _7348_ (.Y(_2379_),
    .B1(_2312_),
    .B2(_2328_),
    .A2(_2378_),
    .A1(_2359_));
 sg13g2_xnor2_1 _7349_ (.Y(_2380_),
    .A(_2377_),
    .B(_2379_));
 sg13g2_nand2_1 _7350_ (.Y(_2381_),
    .A(_2376_),
    .B(_2380_));
 sg13g2_nand2_1 _7351_ (.Y(_2382_),
    .A(_2274_),
    .B(_2288_));
 sg13g2_nand2b_1 _7352_ (.Y(_2383_),
    .B(_2382_),
    .A_N(_2286_));
 sg13g2_nand2_1 _7353_ (.Y(_2384_),
    .A(_2383_),
    .B(_2289_));
 sg13g2_nand2_1 _7354_ (.Y(_2385_),
    .A(_2384_),
    .B(_2331_));
 sg13g2_nor2_1 _7355_ (.A(_2234_),
    .B(_2272_),
    .Y(_2386_));
 sg13g2_nand2_1 _7356_ (.Y(_2387_),
    .A(_2257_),
    .B(_2386_));
 sg13g2_nand2_1 _7357_ (.Y(_2388_),
    .A(_2387_),
    .B(_2277_));
 sg13g2_nand2_1 _7358_ (.Y(_2389_),
    .A(_2388_),
    .B(_2283_));
 sg13g2_nand3_1 _7359_ (.B(_2281_),
    .C(net31),
    .A(_2280_),
    .Y(_2390_));
 sg13g2_nand2_1 _7360_ (.Y(_2391_),
    .A(_2284_),
    .B(_2390_));
 sg13g2_nor2_1 _7361_ (.A(net19),
    .B(_2323_),
    .Y(_2392_));
 sg13g2_nor2_1 _7362_ (.A(_2284_),
    .B(_2390_),
    .Y(_2393_));
 sg13g2_a21oi_1 _7363_ (.A1(_2391_),
    .A2(_2392_),
    .Y(_2394_),
    .B1(_2393_));
 sg13g2_inv_1 _7364_ (.Y(_2395_),
    .A(_2283_));
 sg13g2_nand3_1 _7365_ (.B(_2277_),
    .C(_2395_),
    .A(_2387_),
    .Y(_2396_));
 sg13g2_nand3_1 _7366_ (.B(_2394_),
    .C(_2396_),
    .A(_2389_),
    .Y(_2397_));
 sg13g2_nor2_1 _7367_ (.A(_0587_),
    .B(_2306_),
    .Y(_2398_));
 sg13g2_nor2_1 _7368_ (.A(_2318_),
    .B(_2311_),
    .Y(_2399_));
 sg13g2_nand2b_1 _7369_ (.Y(_2400_),
    .B(_2399_),
    .A_N(_2378_));
 sg13g2_nand2b_1 _7370_ (.Y(_2401_),
    .B(_2378_),
    .A_N(_2399_));
 sg13g2_nand2_1 _7371_ (.Y(_2402_),
    .A(_2400_),
    .B(_2401_));
 sg13g2_nand2b_1 _7372_ (.Y(_2403_),
    .B(_2402_),
    .A_N(_2398_));
 sg13g2_nand3_1 _7373_ (.B(_2401_),
    .C(_2398_),
    .A(_2400_),
    .Y(_2404_));
 sg13g2_nand2_1 _7374_ (.Y(_2405_),
    .A(_2403_),
    .B(_2404_));
 sg13g2_a21oi_1 _7375_ (.A1(_2389_),
    .A2(_2396_),
    .Y(_2406_),
    .B1(_2394_));
 sg13g2_a21oi_1 _7376_ (.A1(_2397_),
    .A2(_2405_),
    .Y(_2407_),
    .B1(_2406_));
 sg13g2_xnor2_1 _7377_ (.Y(_2408_),
    .A(_2312_),
    .B(_2328_));
 sg13g2_nand3_1 _7378_ (.B(_2289_),
    .C(_2408_),
    .A(_2383_),
    .Y(_2409_));
 sg13g2_nand3_1 _7379_ (.B(_2407_),
    .C(_2409_),
    .A(_2385_),
    .Y(_2410_));
 sg13g2_nor2_1 _7380_ (.A(_0587_),
    .B(_2304_),
    .Y(_2411_));
 sg13g2_nor2_1 _7381_ (.A(_2315_),
    .B(_2311_),
    .Y(_2412_));
 sg13g2_a22oi_1 _7382_ (.Y(_2413_),
    .B1(_2398_),
    .B2(_2402_),
    .A2(_2412_),
    .A1(_2324_));
 sg13g2_xnor2_1 _7383_ (.Y(_2414_),
    .A(_2411_),
    .B(_2413_));
 sg13g2_nand2_1 _7384_ (.Y(_2415_),
    .A(_2385_),
    .B(_2409_));
 sg13g2_inv_1 _7385_ (.Y(_2416_),
    .A(_2407_));
 sg13g2_nand2_1 _7386_ (.Y(_2417_),
    .A(_2415_),
    .B(_2416_));
 sg13g2_inv_1 _7387_ (.Y(_2418_),
    .A(_2417_));
 sg13g2_a21oi_1 _7388_ (.A1(_2410_),
    .A2(_2414_),
    .Y(_2419_),
    .B1(_2418_));
 sg13g2_inv_1 _7389_ (.Y(_2420_),
    .A(_2380_));
 sg13g2_nand3_1 _7390_ (.B(_2375_),
    .C(_2420_),
    .A(_2374_),
    .Y(_2421_));
 sg13g2_nand3_1 _7391_ (.B(_2419_),
    .C(_2421_),
    .A(_2381_),
    .Y(_2422_));
 sg13g2_nor2b_2 _7392_ (.A(_2413_),
    .B_N(_2411_),
    .Y(_2423_));
 sg13g2_nand2_1 _7393_ (.Y(_2424_),
    .A(_2381_),
    .B(_2421_));
 sg13g2_inv_1 _7394_ (.Y(_2425_),
    .A(_2419_));
 sg13g2_nand2_1 _7395_ (.Y(_2426_),
    .A(_2424_),
    .B(_2425_));
 sg13g2_inv_1 _7396_ (.Y(_2427_),
    .A(_2426_));
 sg13g2_a21oi_1 _7397_ (.A1(_2422_),
    .A2(_2423_),
    .Y(_2428_),
    .B1(_2427_));
 sg13g2_nor2b_1 _7398_ (.A(_2379_),
    .B_N(_2377_),
    .Y(_2429_));
 sg13g2_inv_1 _7399_ (.Y(_2430_),
    .A(_2374_));
 sg13g2_a21oi_1 _7400_ (.A1(_2375_),
    .A2(_2380_),
    .Y(_2431_),
    .B1(_2430_));
 sg13g2_nand3_1 _7401_ (.B(_2342_),
    .C(net31),
    .A(_2340_),
    .Y(_2432_));
 sg13g2_buf_1 _7402_ (.A(_2432_),
    .X(_2433_));
 sg13g2_nor2_1 _7403_ (.A(_2259_),
    .B(_2433_),
    .Y(_2434_));
 sg13g2_a21oi_1 _7404_ (.A1(_2348_),
    .A2(_2350_),
    .Y(_2435_),
    .B1(_2434_));
 sg13g2_nor3_1 _7405_ (.A(_0685_),
    .B(\generated._508[6] ),
    .C(_2237_),
    .Y(_2436_));
 sg13g2_xnor2_1 _7406_ (.Y(_2437_),
    .A(_0713_),
    .B(_2436_));
 sg13g2_nand2_1 _7407_ (.Y(_2438_),
    .A(_2079_),
    .B(_2437_));
 sg13g2_nand3_1 _7408_ (.B(_0082_),
    .C(_2078_),
    .A(_2240_),
    .Y(_2439_));
 sg13g2_nand2_1 _7409_ (.Y(_2440_),
    .A(_2438_),
    .B(_2439_));
 sg13g2_buf_2 _7410_ (.A(_2440_),
    .X(_2441_));
 sg13g2_nor2_1 _7411_ (.A(_2234_),
    .B(_2441_),
    .Y(_2442_));
 sg13g2_nand2_1 _7412_ (.Y(_2443_),
    .A(_2345_),
    .B(_2442_));
 sg13g2_nand3_1 _7413_ (.B(_2439_),
    .C(net37),
    .A(_2438_),
    .Y(_2444_));
 sg13g2_nand2_1 _7414_ (.Y(_2445_),
    .A(_2433_),
    .B(_2444_));
 sg13g2_nand2_1 _7415_ (.Y(_2446_),
    .A(_2443_),
    .B(_2445_));
 sg13g2_nor2_1 _7416_ (.A(_2267_),
    .B(_2243_),
    .Y(_2447_));
 sg13g2_nand2_1 _7417_ (.Y(_2448_),
    .A(_2446_),
    .B(_2447_));
 sg13g2_inv_1 _7418_ (.Y(_2449_),
    .A(_2447_));
 sg13g2_nand3_1 _7419_ (.B(_2445_),
    .C(_2449_),
    .A(_2443_),
    .Y(_2450_));
 sg13g2_nand2_1 _7420_ (.Y(_2451_),
    .A(_2448_),
    .B(_2450_));
 sg13g2_nand2b_1 _7421_ (.Y(_2452_),
    .B(_2451_),
    .A_N(_2435_));
 sg13g2_nand3_1 _7422_ (.B(_2435_),
    .C(_2450_),
    .A(_2448_),
    .Y(_2453_));
 sg13g2_nand2_1 _7423_ (.Y(_2454_),
    .A(_2452_),
    .B(_2453_));
 sg13g2_nor2_1 _7424_ (.A(_2306_),
    .B(_2282_),
    .Y(_2455_));
 sg13g2_inv_1 _7425_ (.Y(_2456_),
    .A(_2455_));
 sg13g2_nor2_1 _7426_ (.A(_2318_),
    .B(_2272_),
    .Y(_2457_));
 sg13g2_nor2_1 _7427_ (.A(_2315_),
    .B(_2256_),
    .Y(_2458_));
 sg13g2_xnor2_1 _7428_ (.Y(_2459_),
    .A(_2457_),
    .B(_2458_));
 sg13g2_xnor2_1 _7429_ (.Y(_2460_),
    .A(_2456_),
    .B(_2459_));
 sg13g2_inv_1 _7430_ (.Y(_2461_),
    .A(_2460_));
 sg13g2_nand2_1 _7431_ (.Y(_2462_),
    .A(_2454_),
    .B(_2461_));
 sg13g2_nand3_1 _7432_ (.B(_2453_),
    .C(_2460_),
    .A(_2452_),
    .Y(_2463_));
 sg13g2_nand2_1 _7433_ (.Y(_2464_),
    .A(_2462_),
    .B(_2463_));
 sg13g2_a21oi_1 _7434_ (.A1(_2351_),
    .A2(_2353_),
    .Y(_2465_),
    .B1(_2336_));
 sg13g2_a21oi_1 _7435_ (.A1(_2356_),
    .A2(_2367_),
    .Y(_2466_),
    .B1(_2465_));
 sg13g2_inv_1 _7436_ (.Y(_2467_),
    .A(_2466_));
 sg13g2_nand2_1 _7437_ (.Y(_2468_),
    .A(_2464_),
    .B(_2467_));
 sg13g2_nand3_1 _7438_ (.B(_2466_),
    .C(_2463_),
    .A(_2462_),
    .Y(_2469_));
 sg13g2_buf_1 _7439_ (.A(_2469_),
    .X(_2470_));
 sg13g2_nand2_1 _7440_ (.Y(_2471_),
    .A(_2468_),
    .B(_2470_));
 sg13g2_nor2_1 _7441_ (.A(net14),
    .B(_2323_),
    .Y(_2472_));
 sg13g2_a22oi_1 _7442_ (.Y(_2473_),
    .B1(_2363_),
    .B2(_2362_),
    .A2(_2316_),
    .A1(_2457_));
 sg13g2_xnor2_1 _7443_ (.Y(_2474_),
    .A(_2472_),
    .B(_2473_));
 sg13g2_nand2_1 _7444_ (.Y(_2475_),
    .A(_2471_),
    .B(_2474_));
 sg13g2_inv_1 _7445_ (.Y(_2476_),
    .A(_2474_));
 sg13g2_nand3_1 _7446_ (.B(_2470_),
    .C(_2476_),
    .A(_2468_),
    .Y(_2477_));
 sg13g2_nand2_1 _7447_ (.Y(_2478_),
    .A(_2475_),
    .B(_2477_));
 sg13g2_nand2b_1 _7448_ (.Y(_2479_),
    .B(_2478_),
    .A_N(_2431_));
 sg13g2_nand3_1 _7449_ (.B(_2475_),
    .C(_2477_),
    .A(_2431_),
    .Y(_2480_));
 sg13g2_buf_1 _7450_ (.A(_2480_),
    .X(_2481_));
 sg13g2_nand2_1 _7451_ (.Y(_2482_),
    .A(_2479_),
    .B(_2481_));
 sg13g2_nand2b_1 _7452_ (.Y(_2483_),
    .B(_2482_),
    .A_N(_2429_));
 sg13g2_nand3_1 _7453_ (.B(_2481_),
    .C(_2429_),
    .A(_2479_),
    .Y(_2484_));
 sg13g2_nand2_1 _7454_ (.Y(_2485_),
    .A(_2483_),
    .B(_2484_));
 sg13g2_nand2b_1 _7455_ (.Y(_2486_),
    .B(_2485_),
    .A_N(_2428_));
 sg13g2_nand3_1 _7456_ (.B(_2428_),
    .C(_2484_),
    .A(_2483_),
    .Y(_2487_));
 sg13g2_nand2_1 _7457_ (.Y(_2488_),
    .A(_2426_),
    .B(_2422_));
 sg13g2_nand2b_1 _7458_ (.Y(_2489_),
    .B(_2488_),
    .A_N(_2423_));
 sg13g2_nand3_1 _7459_ (.B(_2422_),
    .C(_2423_),
    .A(_2426_),
    .Y(_2490_));
 sg13g2_inv_1 _7460_ (.Y(_2491_),
    .A(_2414_));
 sg13g2_nand2_1 _7461_ (.Y(_2492_),
    .A(_2417_),
    .B(_2410_));
 sg13g2_xnor2_1 _7462_ (.Y(_2493_),
    .A(_2491_),
    .B(_2492_));
 sg13g2_nor2b_1 _7463_ (.A(_2393_),
    .B_N(_2391_),
    .Y(_2494_));
 sg13g2_xnor2_1 _7464_ (.Y(_2495_),
    .A(_2392_),
    .B(_2494_));
 sg13g2_inv_1 _7465_ (.Y(_2496_),
    .A(_2282_));
 sg13g2_nand2_1 _7466_ (.Y(_2497_),
    .A(_2496_),
    .B(net37));
 sg13g2_nand3_1 _7467_ (.B(_2321_),
    .C(net31),
    .A(_2320_),
    .Y(_2498_));
 sg13g2_nand2_1 _7468_ (.Y(_2499_),
    .A(_2497_),
    .B(_2498_));
 sg13g2_nor2_1 _7469_ (.A(net19),
    .B(_2311_),
    .Y(_2500_));
 sg13g2_nor2_1 _7470_ (.A(_2498_),
    .B(_2497_),
    .Y(_2501_));
 sg13g2_a21oi_1 _7471_ (.A1(_2499_),
    .A2(_2500_),
    .Y(_2502_),
    .B1(_2501_));
 sg13g2_nand2_1 _7472_ (.Y(_2503_),
    .A(_2495_),
    .B(_2502_));
 sg13g2_a21oi_1 _7473_ (.A1(_0586_),
    .A2(_2317_),
    .Y(_2504_),
    .B1(_2412_));
 sg13g2_nor2_1 _7474_ (.A(_0587_),
    .B(_2315_),
    .Y(_2505_));
 sg13g2_nand2_1 _7475_ (.Y(_2506_),
    .A(_2399_),
    .B(_2505_));
 sg13g2_nor2b_1 _7476_ (.A(_2504_),
    .B_N(_2506_),
    .Y(_2507_));
 sg13g2_nor2_1 _7477_ (.A(_2502_),
    .B(_2495_),
    .Y(_2508_));
 sg13g2_a21oi_1 _7478_ (.A1(_2503_),
    .A2(_2507_),
    .Y(_2509_),
    .B1(_2508_));
 sg13g2_inv_1 _7479_ (.Y(_2510_),
    .A(_2509_));
 sg13g2_nand2b_1 _7480_ (.Y(_2511_),
    .B(_2397_),
    .A_N(_2406_));
 sg13g2_xnor2_1 _7481_ (.Y(_2512_),
    .A(_2405_),
    .B(_2511_));
 sg13g2_xnor2_1 _7482_ (.Y(_2513_),
    .A(_2510_),
    .B(_2512_));
 sg13g2_nor2_1 _7483_ (.A(_2506_),
    .B(_2513_),
    .Y(_2514_));
 sg13g2_a21oi_1 _7484_ (.A1(_2510_),
    .A2(_2512_),
    .Y(_2515_),
    .B1(_2514_));
 sg13g2_nor2_1 _7485_ (.A(_2493_),
    .B(_2515_),
    .Y(_2516_));
 sg13g2_nand3_1 _7486_ (.B(_2490_),
    .C(_2516_),
    .A(_2489_),
    .Y(_2517_));
 sg13g2_buf_1 _7487_ (.A(_2517_),
    .X(_2518_));
 sg13g2_nand3_1 _7488_ (.B(_2487_),
    .C(_2518_),
    .A(_2486_),
    .Y(_2519_));
 sg13g2_nor2_1 _7489_ (.A(_2304_),
    .B(_2272_),
    .Y(_2520_));
 sg13g2_inv_1 _7490_ (.Y(_2521_),
    .A(net14));
 sg13g2_inv_1 _7491_ (.Y(_2522_),
    .A(_2306_));
 sg13g2_inv_1 _7492_ (.Y(_2523_),
    .A(_2272_));
 sg13g2_a22oi_1 _7493_ (.Y(_2524_),
    .B1(_2522_),
    .B2(_2523_),
    .A2(_2521_),
    .A1(_2496_));
 sg13g2_a21oi_1 _7494_ (.A1(_2455_),
    .A2(_2520_),
    .Y(_2525_),
    .B1(_2524_));
 sg13g2_nor2_1 _7495_ (.A(_2318_),
    .B(_2256_),
    .Y(_2526_));
 sg13g2_inv_1 _7496_ (.Y(_2527_),
    .A(_2459_));
 sg13g2_a22oi_1 _7497_ (.Y(_2528_),
    .B1(_2455_),
    .B2(_2527_),
    .A2(_2526_),
    .A1(_2358_));
 sg13g2_xnor2_1 _7498_ (.Y(_2529_),
    .A(_2525_),
    .B(_2528_));
 sg13g2_inv_1 _7499_ (.Y(_2530_),
    .A(_2452_));
 sg13g2_a21oi_1 _7500_ (.A1(_2453_),
    .A2(_2461_),
    .Y(_2531_),
    .B1(_2530_));
 sg13g2_inv_1 _7501_ (.Y(_2532_),
    .A(_2531_));
 sg13g2_nand3_1 _7502_ (.B(_2242_),
    .C(_2314_),
    .A(_2239_),
    .Y(_2533_));
 sg13g2_inv_2 _7503_ (.Y(_2534_),
    .A(_2533_));
 sg13g2_nand3_1 _7504_ (.B(_2342_),
    .C(_2266_),
    .A(_2340_),
    .Y(_2535_));
 sg13g2_nand2_1 _7505_ (.Y(_2536_),
    .A(_2534_),
    .B(_2535_));
 sg13g2_nor2_1 _7506_ (.A(net19),
    .B(_2344_),
    .Y(_2537_));
 sg13g2_nand2_1 _7507_ (.Y(_2538_),
    .A(_2537_),
    .B(_2533_));
 sg13g2_nand2_1 _7508_ (.Y(_2539_),
    .A(_2536_),
    .B(_2538_));
 sg13g2_inv_1 _7509_ (.Y(_2540_),
    .A(_2526_));
 sg13g2_nand2_1 _7510_ (.Y(_2541_),
    .A(_2539_),
    .B(_2540_));
 sg13g2_nand3_1 _7511_ (.B(_2538_),
    .C(_2526_),
    .A(_2536_),
    .Y(_2542_));
 sg13g2_nand2_1 _7512_ (.Y(_2543_),
    .A(_2541_),
    .B(_2542_));
 sg13g2_nand3_1 _7513_ (.B(_2337_),
    .C(_0713_),
    .A(_2338_),
    .Y(_2544_));
 sg13g2_xnor2_1 _7514_ (.Y(_2545_),
    .A(_0729_),
    .B(_2544_));
 sg13g2_nand2_1 _7515_ (.Y(_2546_),
    .A(_2080_),
    .B(_2545_));
 sg13g2_nand3_1 _7516_ (.B(_1885_),
    .C(net24),
    .A(net13),
    .Y(_2547_));
 sg13g2_nand2_1 _7517_ (.Y(_2548_),
    .A(_2546_),
    .B(_2547_));
 sg13g2_buf_8 _7518_ (.A(_2548_),
    .X(_2549_));
 sg13g2_nor2_1 _7519_ (.A(_2248_),
    .B(_2549_),
    .Y(_2550_));
 sg13g2_xnor2_1 _7520_ (.Y(_2551_),
    .A(_2442_),
    .B(_2550_));
 sg13g2_nor2_1 _7521_ (.A(_2433_),
    .B(_2444_),
    .Y(_2552_));
 sg13g2_a21oi_1 _7522_ (.A1(_2445_),
    .A2(_2447_),
    .Y(_2553_),
    .B1(_2552_));
 sg13g2_xnor2_1 _7523_ (.Y(_2554_),
    .A(_2551_),
    .B(_2553_));
 sg13g2_xnor2_1 _7524_ (.Y(_2555_),
    .A(_2543_),
    .B(_2554_));
 sg13g2_nand2_1 _7525_ (.Y(_2556_),
    .A(_2532_),
    .B(_2555_));
 sg13g2_inv_1 _7526_ (.Y(_2557_),
    .A(_2543_));
 sg13g2_xnor2_1 _7527_ (.Y(_2558_),
    .A(_2557_),
    .B(_2554_));
 sg13g2_nand2_1 _7528_ (.Y(_2559_),
    .A(_2558_),
    .B(_2531_));
 sg13g2_nand2_1 _7529_ (.Y(_2560_),
    .A(_2556_),
    .B(_2559_));
 sg13g2_nand2b_1 _7530_ (.Y(_2561_),
    .B(_2560_),
    .A_N(_2529_));
 sg13g2_nand3_1 _7531_ (.B(_2559_),
    .C(_2529_),
    .A(_2556_),
    .Y(_2562_));
 sg13g2_nand2_1 _7532_ (.Y(_2563_),
    .A(_2561_),
    .B(_2562_));
 sg13g2_inv_1 _7533_ (.Y(_2564_),
    .A(_2468_));
 sg13g2_a21oi_2 _7534_ (.B1(_2564_),
    .Y(_2565_),
    .A2(_2474_),
    .A1(_2470_));
 sg13g2_nand2_2 _7535_ (.Y(_2566_),
    .A(_2563_),
    .B(_2565_));
 sg13g2_nor2b_2 _7536_ (.A(_2473_),
    .B_N(_2472_),
    .Y(_2567_));
 sg13g2_nor2_1 _7537_ (.A(_2565_),
    .B(_2563_),
    .Y(_2568_));
 sg13g2_a21oi_2 _7538_ (.B1(_2568_),
    .Y(_2569_),
    .A2(_2567_),
    .A1(_2566_));
 sg13g2_nand2_1 _7539_ (.Y(_2570_),
    .A(_2456_),
    .B(_2520_));
 sg13g2_nor2_1 _7540_ (.A(_2533_),
    .B(_2535_),
    .Y(_2571_));
 sg13g2_a21oi_1 _7541_ (.A1(_2539_),
    .A2(_2526_),
    .Y(_2572_),
    .B1(_2571_));
 sg13g2_xor2_1 _7542_ (.B(_2572_),
    .A(_2570_),
    .X(_2573_));
 sg13g2_inv_1 _7543_ (.Y(_2574_),
    .A(_2256_));
 sg13g2_nand2_1 _7544_ (.Y(_2575_),
    .A(_2574_),
    .B(_2522_));
 sg13g2_nor2_1 _7545_ (.A(_2318_),
    .B(_2344_),
    .Y(_2576_));
 sg13g2_nand2_1 _7546_ (.Y(_2577_),
    .A(_2534_),
    .B(_2576_));
 sg13g2_nand3_1 _7547_ (.B(_2342_),
    .C(_2314_),
    .A(_2340_),
    .Y(_2578_));
 sg13g2_nand3_1 _7548_ (.B(_2242_),
    .C(_2317_),
    .A(_2239_),
    .Y(_2579_));
 sg13g2_nand2_1 _7549_ (.Y(_2580_),
    .A(_2578_),
    .B(_2579_));
 sg13g2_nand2_1 _7550_ (.Y(_2581_),
    .A(_2577_),
    .B(_2580_));
 sg13g2_xnor2_1 _7551_ (.Y(_2582_),
    .A(_2575_),
    .B(_2581_));
 sg13g2_nand4_1 _7552_ (.B(_2547_),
    .C(_2247_),
    .A(_2546_),
    .Y(_2583_),
    .D(_2233_));
 sg13g2_buf_1 _7553_ (.A(_2583_),
    .X(_2584_));
 sg13g2_a21oi_1 _7554_ (.A1(_2248_),
    .A2(_2234_),
    .Y(_2585_),
    .B1(_2549_));
 sg13g2_nand2_1 _7555_ (.Y(_2586_),
    .A(_2584_),
    .B(_2585_));
 sg13g2_nand2_1 _7556_ (.Y(_2587_),
    .A(_2442_),
    .B(_2550_));
 sg13g2_nor2_1 _7557_ (.A(net19),
    .B(_2441_),
    .Y(_2588_));
 sg13g2_inv_1 _7558_ (.Y(_2589_),
    .A(_2588_));
 sg13g2_nand3_1 _7559_ (.B(_2587_),
    .C(_2589_),
    .A(_2586_),
    .Y(_2590_));
 sg13g2_nand2_1 _7560_ (.Y(_2591_),
    .A(_2585_),
    .B(_2588_));
 sg13g2_nand2_1 _7561_ (.Y(_2592_),
    .A(_2590_),
    .B(_2591_));
 sg13g2_xnor2_1 _7562_ (.Y(_2593_),
    .A(_2582_),
    .B(_2592_));
 sg13g2_nand2_1 _7563_ (.Y(_2594_),
    .A(_2553_),
    .B(_2551_));
 sg13g2_nor2_1 _7564_ (.A(_2551_),
    .B(_2553_),
    .Y(_2595_));
 sg13g2_a21oi_1 _7565_ (.A1(_2543_),
    .A2(_2594_),
    .Y(_2596_),
    .B1(_2595_));
 sg13g2_nand2_1 _7566_ (.Y(_2597_),
    .A(_2593_),
    .B(_2596_));
 sg13g2_inv_1 _7567_ (.Y(_2598_),
    .A(_2575_));
 sg13g2_xnor2_1 _7568_ (.Y(_2599_),
    .A(_2598_),
    .B(_2581_));
 sg13g2_xnor2_1 _7569_ (.Y(_2600_),
    .A(_2599_),
    .B(_2592_));
 sg13g2_inv_1 _7570_ (.Y(_2601_),
    .A(_2596_));
 sg13g2_nand2_1 _7571_ (.Y(_2602_),
    .A(_2600_),
    .B(_2601_));
 sg13g2_nand2_1 _7572_ (.Y(_2603_),
    .A(_2597_),
    .B(_2602_));
 sg13g2_xnor2_1 _7573_ (.Y(_2604_),
    .A(_2573_),
    .B(_2603_));
 sg13g2_nor2_1 _7574_ (.A(_2531_),
    .B(_2558_),
    .Y(_2605_));
 sg13g2_a21oi_1 _7575_ (.A1(_2559_),
    .A2(_2529_),
    .Y(_2606_),
    .B1(_2605_));
 sg13g2_inv_1 _7576_ (.Y(_2607_),
    .A(_2606_));
 sg13g2_nand2_1 _7577_ (.Y(_2608_),
    .A(_2604_),
    .B(_2607_));
 sg13g2_nand2b_1 _7578_ (.Y(_2609_),
    .B(_2603_),
    .A_N(_2573_));
 sg13g2_nand3_1 _7579_ (.B(_2602_),
    .C(_2573_),
    .A(_2597_),
    .Y(_2610_));
 sg13g2_nand2_1 _7580_ (.Y(_2611_),
    .A(_2609_),
    .B(_2610_));
 sg13g2_nand2_1 _7581_ (.Y(_2612_),
    .A(_2611_),
    .B(_2606_));
 sg13g2_nand2_1 _7582_ (.Y(_2613_),
    .A(_2608_),
    .B(_2612_));
 sg13g2_nor2b_1 _7583_ (.A(_2528_),
    .B_N(_2525_),
    .Y(_2614_));
 sg13g2_inv_1 _7584_ (.Y(_2615_),
    .A(_2614_));
 sg13g2_nand2_1 _7585_ (.Y(_2616_),
    .A(_2613_),
    .B(_2615_));
 sg13g2_nand3_1 _7586_ (.B(_2612_),
    .C(_2614_),
    .A(_2608_),
    .Y(_2617_));
 sg13g2_nand2_1 _7587_ (.Y(_2618_),
    .A(_2616_),
    .B(_2617_));
 sg13g2_xnor2_1 _7588_ (.Y(_2619_),
    .A(_2569_),
    .B(_2618_));
 sg13g2_a21oi_1 _7589_ (.A1(_2475_),
    .A2(_2477_),
    .Y(_2620_),
    .B1(_2431_));
 sg13g2_a21oi_2 _7590_ (.B1(_2620_),
    .Y(_2621_),
    .A2(_2429_),
    .A1(_2481_));
 sg13g2_xnor2_1 _7591_ (.Y(_2622_),
    .A(_2529_),
    .B(_2560_));
 sg13g2_inv_1 _7592_ (.Y(_2623_),
    .A(_2565_));
 sg13g2_nand2_1 _7593_ (.Y(_2624_),
    .A(_2622_),
    .B(_2623_));
 sg13g2_nand2_1 _7594_ (.Y(_2625_),
    .A(_2624_),
    .B(_2566_));
 sg13g2_inv_1 _7595_ (.Y(_2626_),
    .A(_2567_));
 sg13g2_nand2_1 _7596_ (.Y(_2627_),
    .A(_2625_),
    .B(_2626_));
 sg13g2_nand3_1 _7597_ (.B(_2566_),
    .C(_2567_),
    .A(_2624_),
    .Y(_2628_));
 sg13g2_nand2_1 _7598_ (.Y(_2629_),
    .A(_2627_),
    .B(_2628_));
 sg13g2_nor2_1 _7599_ (.A(_2621_),
    .B(_2629_),
    .Y(_2630_));
 sg13g2_nand2_1 _7600_ (.Y(_2631_),
    .A(_2619_),
    .B(_2630_));
 sg13g2_inv_1 _7601_ (.Y(_2632_),
    .A(_2569_));
 sg13g2_nand2_1 _7602_ (.Y(_2633_),
    .A(_2618_),
    .B(_2632_));
 sg13g2_nand2_1 _7603_ (.Y(_2634_),
    .A(_2613_),
    .B(_2614_));
 sg13g2_nand3_1 _7604_ (.B(_2612_),
    .C(_2615_),
    .A(_2608_),
    .Y(_2635_));
 sg13g2_nand2_1 _7605_ (.Y(_2636_),
    .A(_2634_),
    .B(_2635_));
 sg13g2_nand2_1 _7606_ (.Y(_2637_),
    .A(_2636_),
    .B(_2569_));
 sg13g2_nand2_1 _7607_ (.Y(_2638_),
    .A(_2633_),
    .B(_2637_));
 sg13g2_nand2_1 _7608_ (.Y(_2639_),
    .A(_2625_),
    .B(_2567_));
 sg13g2_nand3_1 _7609_ (.B(_2566_),
    .C(_2626_),
    .A(_2624_),
    .Y(_2640_));
 sg13g2_nand2_1 _7610_ (.Y(_2641_),
    .A(_2639_),
    .B(_2640_));
 sg13g2_nand2b_1 _7611_ (.Y(_2642_),
    .B(_2641_),
    .A_N(_2621_));
 sg13g2_nand2_1 _7612_ (.Y(_2643_),
    .A(_2638_),
    .B(_2642_));
 sg13g2_nand2_1 _7613_ (.Y(_2644_),
    .A(_2631_),
    .B(_2643_));
 sg13g2_xnor2_1 _7614_ (.Y(_2645_),
    .A(_2621_),
    .B(_2629_));
 sg13g2_nor2_1 _7615_ (.A(_2428_),
    .B(_2485_),
    .Y(_2646_));
 sg13g2_inv_1 _7616_ (.Y(_2647_),
    .A(_2646_));
 sg13g2_nand2_1 _7617_ (.Y(_2648_),
    .A(_2645_),
    .B(_2647_));
 sg13g2_nand3_1 _7618_ (.B(_2644_),
    .C(_2648_),
    .A(_2519_),
    .Y(_2649_));
 sg13g2_nand2_1 _7619_ (.Y(_2650_),
    .A(_2489_),
    .B(_2490_));
 sg13g2_inv_1 _7620_ (.Y(_2651_),
    .A(_2516_));
 sg13g2_nand2_1 _7621_ (.Y(_2652_),
    .A(_2650_),
    .B(_2651_));
 sg13g2_nand2_1 _7622_ (.Y(_2653_),
    .A(_2652_),
    .B(_2518_));
 sg13g2_nand2_1 _7623_ (.Y(_2654_),
    .A(_2515_),
    .B(_2493_));
 sg13g2_inv_1 _7624_ (.Y(_2655_),
    .A(_2654_));
 sg13g2_nor2_1 _7625_ (.A(_2516_),
    .B(_2655_),
    .Y(_2656_));
 sg13g2_nor2b_1 _7626_ (.A(_2508_),
    .B_N(_2503_),
    .Y(_2657_));
 sg13g2_xnor2_1 _7627_ (.Y(_2658_),
    .A(_2507_),
    .B(_2657_));
 sg13g2_nor2b_1 _7628_ (.A(_2501_),
    .B_N(_2499_),
    .Y(_2659_));
 sg13g2_xnor2_1 _7629_ (.Y(_2660_),
    .A(_2500_),
    .B(_2659_));
 sg13g2_nor2_1 _7630_ (.A(_2248_),
    .B(_2323_),
    .Y(_2661_));
 sg13g2_nor2_1 _7631_ (.A(_2234_),
    .B(_2311_),
    .Y(_2662_));
 sg13g2_xor2_1 _7632_ (.B(_2662_),
    .A(_2661_),
    .X(_2663_));
 sg13g2_inv_1 _7633_ (.Y(_2664_),
    .A(_2663_));
 sg13g2_nor3_1 _7634_ (.A(_0587_),
    .B(net19),
    .C(_2664_),
    .Y(_2665_));
 sg13g2_a21oi_1 _7635_ (.A1(_2661_),
    .A2(_2662_),
    .Y(_2666_),
    .B1(_2665_));
 sg13g2_nor2_1 _7636_ (.A(_2660_),
    .B(_2666_),
    .Y(_2667_));
 sg13g2_xnor2_1 _7637_ (.Y(_2668_),
    .A(_2660_),
    .B(_2666_));
 sg13g2_nor2b_1 _7638_ (.A(_2668_),
    .B_N(_2505_),
    .Y(_2669_));
 sg13g2_nor2_1 _7639_ (.A(_2667_),
    .B(_2669_),
    .Y(_2670_));
 sg13g2_xnor2_1 _7640_ (.Y(_2671_),
    .A(_2506_),
    .B(_2513_));
 sg13g2_nor3_2 _7641_ (.A(_2658_),
    .B(_2670_),
    .C(_2671_),
    .Y(_2672_));
 sg13g2_nand2_1 _7642_ (.Y(_2673_),
    .A(_2656_),
    .B(_2672_));
 sg13g2_nand2_1 _7643_ (.Y(_2674_),
    .A(_2653_),
    .B(_2673_));
 sg13g2_and2_1 _7644_ (.A(_2670_),
    .B(_2658_),
    .X(_2675_));
 sg13g2_nand3_1 _7645_ (.B(_2249_),
    .C(net37),
    .A(_2662_),
    .Y(_2676_));
 sg13g2_o21ai_1 _7646_ (.B1(_2664_),
    .Y(_2677_),
    .A1(_0587_),
    .A2(net19));
 sg13g2_nand2b_1 _7647_ (.Y(_2678_),
    .B(_2677_),
    .A_N(_2665_));
 sg13g2_nor2b_1 _7648_ (.A(_2505_),
    .B_N(_2668_),
    .Y(_2679_));
 sg13g2_nor4_1 _7649_ (.A(_2676_),
    .B(_2678_),
    .C(_2669_),
    .D(_2679_),
    .Y(_2680_));
 sg13g2_o21ai_1 _7650_ (.B1(_2680_),
    .Y(_2681_),
    .A1(_2658_),
    .A2(_2670_));
 sg13g2_nor3_1 _7651_ (.A(_2671_),
    .B(_2675_),
    .C(_2681_),
    .Y(_2682_));
 sg13g2_and2_1 _7652_ (.A(_2682_),
    .B(_2656_),
    .X(_2683_));
 sg13g2_nand2_1 _7653_ (.Y(_2684_),
    .A(_2486_),
    .B(_2487_));
 sg13g2_a21oi_1 _7654_ (.A1(_2674_),
    .A2(_2683_),
    .Y(_2685_),
    .B1(_2684_));
 sg13g2_nor2_1 _7655_ (.A(_2649_),
    .B(_2685_),
    .Y(_2686_));
 sg13g2_nand2_1 _7656_ (.Y(_2687_),
    .A(_2674_),
    .B(_2683_));
 sg13g2_xnor2_1 _7657_ (.Y(_2688_),
    .A(_2423_),
    .B(_2488_));
 sg13g2_nand4_1 _7658_ (.B(_2651_),
    .C(_2654_),
    .A(_2688_),
    .Y(_2689_),
    .D(_2672_));
 sg13g2_buf_1 _7659_ (.A(_2689_),
    .X(_2690_));
 sg13g2_nand3_1 _7660_ (.B(_2518_),
    .C(_2690_),
    .A(_2687_),
    .Y(_2691_));
 sg13g2_nand2_1 _7661_ (.Y(_2692_),
    .A(_2686_),
    .B(_2691_));
 sg13g2_xnor2_1 _7662_ (.Y(_2693_),
    .A(_2621_),
    .B(_2641_));
 sg13g2_nand2_1 _7663_ (.Y(_2694_),
    .A(_2693_),
    .B(_2646_));
 sg13g2_inv_2 _7664_ (.Y(_2695_),
    .A(_2644_));
 sg13g2_nor2_1 _7665_ (.A(_2694_),
    .B(_2695_),
    .Y(_2696_));
 sg13g2_nand2_1 _7666_ (.Y(_2697_),
    .A(_2638_),
    .B(_2630_));
 sg13g2_nor2b_1 _7667_ (.A(_2696_),
    .B_N(_2697_),
    .Y(_2698_));
 sg13g2_buf_1 _7668_ (.A(_2698_),
    .X(_2699_));
 sg13g2_nand2_1 _7669_ (.Y(_2700_),
    .A(_2692_),
    .B(_2699_));
 sg13g2_nor2_1 _7670_ (.A(_2569_),
    .B(_2618_),
    .Y(_2701_));
 sg13g2_inv_1 _7671_ (.Y(_2702_),
    .A(_2520_));
 sg13g2_a21oi_1 _7672_ (.A1(_2572_),
    .A2(_2456_),
    .Y(_2703_),
    .B1(_2702_));
 sg13g2_nor2_1 _7673_ (.A(net14),
    .B(_2256_),
    .Y(_2704_));
 sg13g2_a22oi_1 _7674_ (.Y(_2705_),
    .B1(_2598_),
    .B2(_2580_),
    .A2(_2576_),
    .A1(_2534_));
 sg13g2_xnor2_1 _7675_ (.Y(_2706_),
    .A(_2704_),
    .B(_2705_));
 sg13g2_nor2_1 _7676_ (.A(net19),
    .B(_2587_),
    .Y(_2707_));
 sg13g2_nor2_1 _7677_ (.A(_2582_),
    .B(_2592_),
    .Y(_2708_));
 sg13g2_nor2_1 _7678_ (.A(_2707_),
    .B(_2708_),
    .Y(_2709_));
 sg13g2_nand2_1 _7679_ (.Y(_2710_),
    .A(_2591_),
    .B(_2584_));
 sg13g2_nor2_1 _7680_ (.A(_2278_),
    .B(_2549_),
    .Y(_2711_));
 sg13g2_inv_1 _7681_ (.Y(_2712_),
    .A(_2711_));
 sg13g2_xnor2_1 _7682_ (.Y(_2713_),
    .A(_2712_),
    .B(_2586_));
 sg13g2_nand2b_1 _7683_ (.Y(_2714_),
    .B(_2713_),
    .A_N(_2710_));
 sg13g2_nor2_2 _7684_ (.A(_2278_),
    .B(_2584_),
    .Y(_2715_));
 sg13g2_inv_1 _7685_ (.Y(_2716_),
    .A(_2715_));
 sg13g2_nand2_1 _7686_ (.Y(_2717_),
    .A(_2714_),
    .B(_2716_));
 sg13g2_nor2_1 _7687_ (.A(_2306_),
    .B(_2243_),
    .Y(_2718_));
 sg13g2_inv_1 _7688_ (.Y(_2719_),
    .A(_2441_));
 sg13g2_nand2_1 _7689_ (.Y(_2720_),
    .A(_2719_),
    .B(_2314_));
 sg13g2_xnor2_1 _7690_ (.Y(_2721_),
    .A(_2576_),
    .B(_2720_));
 sg13g2_xor2_1 _7691_ (.B(_2721_),
    .A(_2718_),
    .X(_2722_));
 sg13g2_inv_1 _7692_ (.Y(_2723_),
    .A(_2722_));
 sg13g2_nand2_1 _7693_ (.Y(_2724_),
    .A(_2717_),
    .B(_2723_));
 sg13g2_nand3_1 _7694_ (.B(_2722_),
    .C(_2716_),
    .A(_2714_),
    .Y(_2725_));
 sg13g2_nand3b_1 _7695_ (.B(_2724_),
    .C(_2725_),
    .Y(_2726_),
    .A_N(_2709_));
 sg13g2_nand2_1 _7696_ (.Y(_2727_),
    .A(_2724_),
    .B(_2725_));
 sg13g2_nand2_1 _7697_ (.Y(_2728_),
    .A(_2727_),
    .B(_2709_));
 sg13g2_nand2_1 _7698_ (.Y(_2729_),
    .A(_2726_),
    .B(_2728_));
 sg13g2_nand2b_1 _7699_ (.Y(_2730_),
    .B(_2729_),
    .A_N(_2706_));
 sg13g2_nand3_1 _7700_ (.B(_2728_),
    .C(_2706_),
    .A(_2726_),
    .Y(_2731_));
 sg13g2_nand2_1 _7701_ (.Y(_2732_),
    .A(_2730_),
    .B(_2731_));
 sg13g2_nand2_1 _7702_ (.Y(_2733_),
    .A(_2610_),
    .B(_2602_));
 sg13g2_inv_1 _7703_ (.Y(_2734_),
    .A(_2733_));
 sg13g2_nand2_1 _7704_ (.Y(_2735_),
    .A(_2732_),
    .B(_2734_));
 sg13g2_nand3_1 _7705_ (.B(_2731_),
    .C(_2733_),
    .A(_2730_),
    .Y(_2736_));
 sg13g2_nand2_1 _7706_ (.Y(_2737_),
    .A(_2735_),
    .B(_2736_));
 sg13g2_nand2b_1 _7707_ (.Y(_2738_),
    .B(_2737_),
    .A_N(_2703_));
 sg13g2_nand3_1 _7708_ (.B(_2736_),
    .C(_2703_),
    .A(_2735_),
    .Y(_2739_));
 sg13g2_nand2_1 _7709_ (.Y(_2740_),
    .A(_2738_),
    .B(_2739_));
 sg13g2_inv_1 _7710_ (.Y(_2741_),
    .A(_2608_));
 sg13g2_a21oi_1 _7711_ (.A1(_2612_),
    .A2(_2614_),
    .Y(_2742_),
    .B1(_2741_));
 sg13g2_inv_1 _7712_ (.Y(_2743_),
    .A(_2742_));
 sg13g2_nand2_1 _7713_ (.Y(_2744_),
    .A(_2740_),
    .B(_2743_));
 sg13g2_nand3_1 _7714_ (.B(_2739_),
    .C(_2742_),
    .A(_2738_),
    .Y(_2745_));
 sg13g2_nand3b_1 _7715_ (.B(_2744_),
    .C(_2745_),
    .Y(_2746_),
    .A_N(_2701_));
 sg13g2_nand2_1 _7716_ (.Y(_2747_),
    .A(_2744_),
    .B(_2745_));
 sg13g2_nand2_1 _7717_ (.Y(_2748_),
    .A(_2747_),
    .B(_2701_));
 sg13g2_nand2_1 _7718_ (.Y(_2749_),
    .A(_2746_),
    .B(_2748_));
 sg13g2_inv_1 _7719_ (.Y(_2750_),
    .A(_2749_));
 sg13g2_nand2_1 _7720_ (.Y(_2751_),
    .A(_2700_),
    .B(_2750_));
 sg13g2_nand3_1 _7721_ (.B(_2749_),
    .C(_2699_),
    .A(_2692_),
    .Y(_2752_));
 sg13g2_nor2_1 _7722_ (.A(net94),
    .B(_4296_),
    .Y(_2753_));
 sg13g2_inv_1 _7723_ (.Y(_2754_),
    .A(_2753_));
 sg13g2_nor2_1 _7724_ (.A(_0116_),
    .B(_1302_),
    .Y(_2755_));
 sg13g2_xor2_1 _7725_ (.B(_2755_),
    .A(_4236_),
    .X(_2756_));
 sg13g2_buf_2 _7726_ (.A(_2756_),
    .X(_2757_));
 sg13g2_nor3_2 _7727_ (.A(_2754_),
    .B(_2757_),
    .C(_4305_),
    .Y(_2758_));
 sg13g2_xnor2_1 _7728_ (.Y(_2759_),
    .A(_4239_),
    .B(_1994_));
 sg13g2_inv_1 _7729_ (.Y(_2760_),
    .A(_2759_));
 sg13g2_nand2_1 _7730_ (.Y(_2761_),
    .A(_4239_),
    .B(\generated._217[1] ));
 sg13g2_inv_1 _7731_ (.Y(_2762_),
    .A(_4304_));
 sg13g2_o21ai_1 _7732_ (.B1(_0125_),
    .Y(_2763_),
    .A1(_2761_),
    .A2(_2762_));
 sg13g2_xnor2_1 _7733_ (.Y(_2764_),
    .A(_0126_),
    .B(_2763_));
 sg13g2_a21oi_1 _7734_ (.A1(_2758_),
    .A2(_2760_),
    .Y(_2765_),
    .B1(_2764_));
 sg13g2_nand3_1 _7735_ (.B(_2758_),
    .C(_2760_),
    .A(_2764_),
    .Y(_2766_));
 sg13g2_nor2b_1 _7736_ (.A(_2765_),
    .B_N(_2766_),
    .Y(_2767_));
 sg13g2_inv_1 _7737_ (.Y(_2768_),
    .A(_2767_));
 sg13g2_buf_1 _7738_ (.A(\generated._558[0] ),
    .X(_2769_));
 sg13g2_xnor2_1 _7739_ (.Y(_2770_),
    .A(_1735_),
    .B(_2769_));
 sg13g2_nand2_1 _7740_ (.Y(_2771_),
    .A(_2073_),
    .B(_2770_));
 sg13g2_nand2_1 _7741_ (.Y(_2772_),
    .A(net11),
    .B(_0071_));
 sg13g2_nand2_2 _7742_ (.Y(_2773_),
    .A(_2771_),
    .B(_2772_));
 sg13g2_nor2_1 _7743_ (.A(net23),
    .B(_2773_),
    .Y(_2774_));
 sg13g2_inv_1 _7744_ (.Y(_2775_),
    .A(_2774_));
 sg13g2_xnor2_1 _7745_ (.Y(_2776_),
    .A(_2759_),
    .B(_2758_));
 sg13g2_buf_2 _7746_ (.A(_2776_),
    .X(_2777_));
 sg13g2_nand3_1 _7747_ (.B(_2777_),
    .C(_2772_),
    .A(_2771_),
    .Y(_2778_));
 sg13g2_nor2_1 _7748_ (.A(_2754_),
    .B(_2757_),
    .Y(_2779_));
 sg13g2_xnor2_1 _7749_ (.Y(_2780_),
    .A(_4305_),
    .B(_2779_));
 sg13g2_inv_1 _7750_ (.Y(_2781_),
    .A(_2780_));
 sg13g2_buf_1 _7751_ (.A(_2781_),
    .X(_2782_));
 sg13g2_nor2_1 _7752_ (.A(_1735_),
    .B(_2769_),
    .Y(_2783_));
 sg13g2_xnor2_1 _7753_ (.Y(_2784_),
    .A(_1801_),
    .B(_2783_));
 sg13g2_nand2_1 _7754_ (.Y(_2785_),
    .A(_2073_),
    .B(_2784_));
 sg13g2_nand2_1 _7755_ (.Y(_2786_),
    .A(net11),
    .B(_0572_));
 sg13g2_nand2_1 _7756_ (.Y(_2787_),
    .A(_2785_),
    .B(_2786_));
 sg13g2_buf_2 _7757_ (.A(_2787_),
    .X(_2788_));
 sg13g2_nor2_1 _7758_ (.A(net22),
    .B(_2788_),
    .Y(_2789_));
 sg13g2_xnor2_1 _7759_ (.Y(_2790_),
    .A(_2778_),
    .B(_2789_));
 sg13g2_inv_1 _7760_ (.Y(_2791_),
    .A(\generated._558[3] ));
 sg13g2_nand3_1 _7761_ (.B(_1801_),
    .C(_2791_),
    .A(_2783_),
    .Y(_2792_));
 sg13g2_xnor2_1 _7762_ (.Y(_2793_),
    .A(_1868_),
    .B(_2792_));
 sg13g2_nand2_1 _7763_ (.Y(_2794_),
    .A(_2072_),
    .B(_2793_));
 sg13g2_nand2_1 _7764_ (.Y(_2795_),
    .A(_2059_),
    .B(_0594_));
 sg13g2_nand2_1 _7765_ (.Y(_2796_),
    .A(_2794_),
    .B(_2795_));
 sg13g2_buf_2 _7766_ (.A(_2796_),
    .X(_2797_));
 sg13g2_nor2_2 _7767_ (.A(net79),
    .B(_2797_),
    .Y(_2798_));
 sg13g2_xnor2_1 _7768_ (.Y(_2799_),
    .A(_2753_),
    .B(_2757_));
 sg13g2_inv_2 _7769_ (.Y(_2800_),
    .A(_2799_));
 sg13g2_nor3_1 _7770_ (.A(_1735_),
    .B(\generated._558[2] ),
    .C(_1688_),
    .Y(_2801_));
 sg13g2_xnor2_1 _7771_ (.Y(_2802_),
    .A(_2791_),
    .B(_2801_));
 sg13g2_nand2_1 _7772_ (.Y(_2803_),
    .A(_2072_),
    .B(_2802_));
 sg13g2_nand2_1 _7773_ (.Y(_2804_),
    .A(_2059_),
    .B(_0077_));
 sg13g2_nand2_1 _7774_ (.Y(_2805_),
    .A(_2803_),
    .B(_2804_));
 sg13g2_buf_2 _7775_ (.A(_2805_),
    .X(_2806_));
 sg13g2_nor2_2 _7776_ (.A(_2800_),
    .B(_2806_),
    .Y(_2807_));
 sg13g2_xnor2_1 _7777_ (.Y(_2808_),
    .A(_2798_),
    .B(_2807_));
 sg13g2_nor2_1 _7778_ (.A(net79),
    .B(_2788_),
    .Y(_2809_));
 sg13g2_nand2_1 _7779_ (.Y(_2810_),
    .A(_2809_),
    .B(_2807_));
 sg13g2_nand2_1 _7780_ (.Y(_2811_),
    .A(_2808_),
    .B(_2810_));
 sg13g2_inv_1 _7781_ (.Y(_2812_),
    .A(_2788_));
 sg13g2_nand4_1 _7782_ (.B(_2812_),
    .C(net94),
    .A(_2807_),
    .Y(_2813_),
    .D(_2797_));
 sg13g2_nand2_1 _7783_ (.Y(_2814_),
    .A(_2811_),
    .B(_2813_));
 sg13g2_nand2b_1 _7784_ (.Y(_2815_),
    .B(_2814_),
    .A_N(_2790_));
 sg13g2_nand3_1 _7785_ (.B(_2813_),
    .C(_2790_),
    .A(_2811_),
    .Y(_2816_));
 sg13g2_nand2_1 _7786_ (.Y(_2817_),
    .A(_2815_),
    .B(_2816_));
 sg13g2_inv_1 _7787_ (.Y(_2818_),
    .A(_2806_));
 sg13g2_nand2_1 _7788_ (.Y(_2819_),
    .A(_2818_),
    .B(net94));
 sg13g2_nand2_1 _7789_ (.Y(_2820_),
    .A(_2812_),
    .B(_2799_));
 sg13g2_nand2_1 _7790_ (.Y(_2821_),
    .A(_2819_),
    .B(_2820_));
 sg13g2_nand2_1 _7791_ (.Y(_2822_),
    .A(_2821_),
    .B(_2810_));
 sg13g2_nor2_1 _7792_ (.A(_2800_),
    .B(_2773_),
    .Y(_2823_));
 sg13g2_nand2_1 _7793_ (.Y(_2824_),
    .A(_2809_),
    .B(_2823_));
 sg13g2_nand2_1 _7794_ (.Y(_2825_),
    .A(_2822_),
    .B(_2824_));
 sg13g2_nand2_1 _7795_ (.Y(_2826_),
    .A(_2777_),
    .B(_2769_));
 sg13g2_nor2_1 _7796_ (.A(net22),
    .B(_2773_),
    .Y(_2827_));
 sg13g2_xnor2_1 _7797_ (.Y(_2828_),
    .A(_2826_),
    .B(_2827_));
 sg13g2_nor2_1 _7798_ (.A(_2824_),
    .B(_2822_),
    .Y(_2829_));
 sg13g2_a21oi_1 _7799_ (.A1(_2825_),
    .A2(_2828_),
    .Y(_2830_),
    .B1(_2829_));
 sg13g2_nand2_1 _7800_ (.Y(_2831_),
    .A(_2817_),
    .B(_2830_));
 sg13g2_nor3_1 _7801_ (.A(net22),
    .B(_2826_),
    .C(_2773_),
    .Y(_2832_));
 sg13g2_nor2_1 _7802_ (.A(_2830_),
    .B(_2817_),
    .Y(_2833_));
 sg13g2_a21oi_1 _7803_ (.A1(_2831_),
    .A2(_2832_),
    .Y(_2834_),
    .B1(_2833_));
 sg13g2_inv_1 _7804_ (.Y(_2835_),
    .A(_2834_));
 sg13g2_inv_1 _7805_ (.Y(_2836_),
    .A(_2813_));
 sg13g2_a21oi_1 _7806_ (.A1(_2811_),
    .A2(_2790_),
    .Y(_2837_),
    .B1(_2836_));
 sg13g2_nor2_1 _7807_ (.A(net22),
    .B(_2806_),
    .Y(_2838_));
 sg13g2_inv_2 _7808_ (.Y(_2839_),
    .A(_2777_));
 sg13g2_nor2_1 _7809_ (.A(_2839_),
    .B(_2788_),
    .Y(_2840_));
 sg13g2_xor2_1 _7810_ (.B(_2840_),
    .A(_2838_),
    .X(_2841_));
 sg13g2_nand3b_1 _7811_ (.B(_2801_),
    .C(_2791_),
    .Y(_2842_),
    .A_N(_1868_));
 sg13g2_xnor2_1 _7812_ (.Y(_2843_),
    .A(_1883_),
    .B(_2842_));
 sg13g2_nand2_1 _7813_ (.Y(_2844_),
    .A(_2072_),
    .B(_2843_));
 sg13g2_nand2_1 _7814_ (.Y(_2845_),
    .A(_2058_),
    .B(_0081_));
 sg13g2_nand2_1 _7815_ (.Y(_2846_),
    .A(_2844_),
    .B(_2845_));
 sg13g2_buf_2 _7816_ (.A(_2846_),
    .X(_2847_));
 sg13g2_nor2_1 _7817_ (.A(net79),
    .B(_2847_),
    .Y(_2848_));
 sg13g2_nor2_1 _7818_ (.A(_2800_),
    .B(_2797_),
    .Y(_2849_));
 sg13g2_xnor2_1 _7819_ (.Y(_2850_),
    .A(_2848_),
    .B(_2849_));
 sg13g2_nand2_1 _7820_ (.Y(_2851_),
    .A(_2798_),
    .B(_2807_));
 sg13g2_nand2_1 _7821_ (.Y(_2852_),
    .A(_2850_),
    .B(_2851_));
 sg13g2_nand4_1 _7822_ (.B(_2818_),
    .C(net94),
    .A(_2849_),
    .Y(_2853_),
    .D(_2847_));
 sg13g2_nand2_1 _7823_ (.Y(_2854_),
    .A(_2852_),
    .B(_2853_));
 sg13g2_xnor2_1 _7824_ (.Y(_2855_),
    .A(_2841_),
    .B(_2854_));
 sg13g2_nand2b_1 _7825_ (.Y(_2856_),
    .B(_2855_),
    .A_N(_2837_));
 sg13g2_nand2b_1 _7826_ (.Y(_2857_),
    .B(_2854_),
    .A_N(_2841_));
 sg13g2_nand3_1 _7827_ (.B(_2841_),
    .C(_2853_),
    .A(_2852_),
    .Y(_2858_));
 sg13g2_nand2_1 _7828_ (.Y(_2859_),
    .A(_2857_),
    .B(_2858_));
 sg13g2_nand2_1 _7829_ (.Y(_2860_),
    .A(_2859_),
    .B(_2837_));
 sg13g2_nand2_1 _7830_ (.Y(_2861_),
    .A(_2856_),
    .B(_2860_));
 sg13g2_nand2_2 _7831_ (.Y(_2862_),
    .A(_2766_),
    .B(_1995_));
 sg13g2_nor3_1 _7832_ (.A(net22),
    .B(_2788_),
    .C(_2778_),
    .Y(_2863_));
 sg13g2_a21oi_1 _7833_ (.A1(_2769_),
    .A2(_2862_),
    .Y(_2864_),
    .B1(_2863_));
 sg13g2_inv_1 _7834_ (.Y(_2865_),
    .A(_2864_));
 sg13g2_nand2_1 _7835_ (.Y(_2866_),
    .A(_2861_),
    .B(_2865_));
 sg13g2_nand3_1 _7836_ (.B(_2860_),
    .C(_2864_),
    .A(_2856_),
    .Y(_2867_));
 sg13g2_nand2_1 _7837_ (.Y(_2868_),
    .A(_2866_),
    .B(_2867_));
 sg13g2_nor2_1 _7838_ (.A(_2835_),
    .B(_2868_),
    .Y(_2869_));
 sg13g2_nand2_1 _7839_ (.Y(_2870_),
    .A(_2868_),
    .B(_2835_));
 sg13g2_o21ai_1 _7840_ (.B1(_2870_),
    .Y(_2871_),
    .A1(_2775_),
    .A2(_2869_));
 sg13g2_nor2_1 _7841_ (.A(_2837_),
    .B(_2859_),
    .Y(_2872_));
 sg13g2_a21oi_1 _7842_ (.A1(_2860_),
    .A2(_2865_),
    .Y(_2873_),
    .B1(_2872_));
 sg13g2_nor2_1 _7843_ (.A(_2782_),
    .B(_2797_),
    .Y(_2874_));
 sg13g2_nor2_1 _7844_ (.A(_2839_),
    .B(_2806_),
    .Y(_2875_));
 sg13g2_xor2_1 _7845_ (.B(_2875_),
    .A(_2874_),
    .X(_2876_));
 sg13g2_or3_1 _7846_ (.A(_1868_),
    .B(_1883_),
    .C(_2792_),
    .X(_2877_));
 sg13g2_xnor2_1 _7847_ (.Y(_2878_),
    .A(_1909_),
    .B(_2877_));
 sg13g2_nand2_1 _7848_ (.Y(_2879_),
    .A(_2072_),
    .B(_2878_));
 sg13g2_nand2_1 _7849_ (.Y(_2880_),
    .A(_2058_),
    .B(_0634_));
 sg13g2_nand2_2 _7850_ (.Y(_2881_),
    .A(_2879_),
    .B(_2880_));
 sg13g2_nor2_1 _7851_ (.A(_2800_),
    .B(_2881_),
    .Y(_2882_));
 sg13g2_nand2_1 _7852_ (.Y(_2883_),
    .A(_2882_),
    .B(_2848_));
 sg13g2_nand3_1 _7853_ (.B(net94),
    .C(_2880_),
    .A(_2879_),
    .Y(_2884_));
 sg13g2_nand3_1 _7854_ (.B(_2799_),
    .C(_2845_),
    .A(_2844_),
    .Y(_2885_));
 sg13g2_nand2_1 _7855_ (.Y(_2886_),
    .A(_2884_),
    .B(_2885_));
 sg13g2_nand2_1 _7856_ (.Y(_2887_),
    .A(_2883_),
    .B(_2886_));
 sg13g2_nor2_1 _7857_ (.A(_2800_),
    .B(_2847_),
    .Y(_2888_));
 sg13g2_nand2_1 _7858_ (.Y(_2889_),
    .A(_2888_),
    .B(_2798_));
 sg13g2_nand2_1 _7859_ (.Y(_2890_),
    .A(_2887_),
    .B(_2889_));
 sg13g2_nand3_1 _7860_ (.B(_2798_),
    .C(_2884_),
    .A(_2888_),
    .Y(_2891_));
 sg13g2_nand2_1 _7861_ (.Y(_2892_),
    .A(_2890_),
    .B(_2891_));
 sg13g2_xor2_1 _7862_ (.B(_2892_),
    .A(_2876_),
    .X(_2893_));
 sg13g2_inv_1 _7863_ (.Y(_2894_),
    .A(_2853_));
 sg13g2_a21oi_1 _7864_ (.A1(_2852_),
    .A2(_2841_),
    .Y(_2895_),
    .B1(_2894_));
 sg13g2_nand2_1 _7865_ (.Y(_2896_),
    .A(_2893_),
    .B(_2895_));
 sg13g2_xnor2_1 _7866_ (.Y(_2897_),
    .A(_2876_),
    .B(_2892_));
 sg13g2_nand2b_1 _7867_ (.Y(_2898_),
    .B(_2897_),
    .A_N(_2895_));
 sg13g2_nand2_1 _7868_ (.Y(_2899_),
    .A(_2896_),
    .B(_2898_));
 sg13g2_inv_2 _7869_ (.Y(_2900_),
    .A(_2862_));
 sg13g2_nand2_1 _7870_ (.Y(_2901_),
    .A(_2789_),
    .B(_2875_));
 sg13g2_o21ai_1 _7871_ (.B1(_2901_),
    .Y(_2902_),
    .A1(_2900_),
    .A2(_2773_));
 sg13g2_nand2_1 _7872_ (.Y(_2903_),
    .A(_2899_),
    .B(_2902_));
 sg13g2_inv_1 _7873_ (.Y(_2904_),
    .A(_2902_));
 sg13g2_nand3_1 _7874_ (.B(_2898_),
    .C(_2904_),
    .A(_2896_),
    .Y(_2905_));
 sg13g2_nand2_1 _7875_ (.Y(_2906_),
    .A(_2903_),
    .B(_2905_));
 sg13g2_nand2b_1 _7876_ (.Y(_2907_),
    .B(_2906_),
    .A_N(_2873_));
 sg13g2_nand3_1 _7877_ (.B(_2873_),
    .C(_2905_),
    .A(_2903_),
    .Y(_2908_));
 sg13g2_nor2_1 _7878_ (.A(net23),
    .B(_2788_),
    .Y(_2909_));
 sg13g2_nand3_1 _7879_ (.B(_2908_),
    .C(_2909_),
    .A(_2907_),
    .Y(_2910_));
 sg13g2_nand2_1 _7880_ (.Y(_2911_),
    .A(_2907_),
    .B(_2908_));
 sg13g2_nand2b_1 _7881_ (.Y(_2912_),
    .B(_2911_),
    .A_N(_2909_));
 sg13g2_nand3_1 _7882_ (.B(_2910_),
    .C(_2912_),
    .A(_2871_),
    .Y(_2913_));
 sg13g2_a21oi_1 _7883_ (.A1(_2903_),
    .A2(_2905_),
    .Y(_2914_),
    .B1(_2873_));
 sg13g2_a21oi_1 _7884_ (.A1(_2908_),
    .A2(_2909_),
    .Y(_2915_),
    .B1(_2914_));
 sg13g2_inv_1 _7885_ (.Y(_2916_),
    .A(_2898_));
 sg13g2_a21oi_1 _7886_ (.A1(_2896_),
    .A2(_2902_),
    .Y(_2917_),
    .B1(_2916_));
 sg13g2_inv_1 _7887_ (.Y(_2918_),
    .A(_2891_));
 sg13g2_a21oi_1 _7888_ (.A1(_2890_),
    .A2(_2876_),
    .Y(_2919_),
    .B1(_2918_));
 sg13g2_nor2_2 _7889_ (.A(net22),
    .B(_2847_),
    .Y(_2920_));
 sg13g2_nor2_1 _7890_ (.A(_2839_),
    .B(_2797_),
    .Y(_2921_));
 sg13g2_xor2_1 _7891_ (.B(_2921_),
    .A(_2920_),
    .X(_2922_));
 sg13g2_nand2_1 _7892_ (.Y(_2923_),
    .A(_2058_),
    .B(_0085_));
 sg13g2_inv_1 _7893_ (.Y(_2924_),
    .A(\generated._558[7] ));
 sg13g2_nor3_1 _7894_ (.A(_1883_),
    .B(_1909_),
    .C(_2842_),
    .Y(_2925_));
 sg13g2_xnor2_1 _7895_ (.Y(_2926_),
    .A(_2924_),
    .B(_2925_));
 sg13g2_nand3_1 _7896_ (.B(_2056_),
    .C(_2926_),
    .A(net13),
    .Y(_2927_));
 sg13g2_nand2_2 _7897_ (.Y(_2928_),
    .A(_2923_),
    .B(_2927_));
 sg13g2_nor2_2 _7898_ (.A(net79),
    .B(_2928_),
    .Y(_2929_));
 sg13g2_xnor2_1 _7899_ (.Y(_2930_),
    .A(_2929_),
    .B(_2882_));
 sg13g2_nand2_1 _7900_ (.Y(_2931_),
    .A(_2930_),
    .B(_2883_));
 sg13g2_inv_1 _7901_ (.Y(_2932_),
    .A(_2929_));
 sg13g2_nand3_1 _7902_ (.B(_2882_),
    .C(_2848_),
    .A(_2932_),
    .Y(_2933_));
 sg13g2_nand2_1 _7903_ (.Y(_2934_),
    .A(_2931_),
    .B(_2933_));
 sg13g2_xnor2_1 _7904_ (.Y(_2935_),
    .A(_2922_),
    .B(_2934_));
 sg13g2_nand2b_1 _7905_ (.Y(_2936_),
    .B(_2935_),
    .A_N(_2919_));
 sg13g2_inv_1 _7906_ (.Y(_2937_),
    .A(_2922_));
 sg13g2_xnor2_1 _7907_ (.Y(_2938_),
    .A(_2937_),
    .B(_2934_));
 sg13g2_nand2_1 _7908_ (.Y(_2939_),
    .A(_2938_),
    .B(_2919_));
 sg13g2_nand2_1 _7909_ (.Y(_2940_),
    .A(_2936_),
    .B(_2939_));
 sg13g2_nand2_1 _7910_ (.Y(_2941_),
    .A(_2921_),
    .B(_2838_));
 sg13g2_o21ai_1 _7911_ (.B1(_2941_),
    .Y(_2942_),
    .A1(_2900_),
    .A2(_2788_));
 sg13g2_nand2_1 _7912_ (.Y(_2943_),
    .A(_2940_),
    .B(_2942_));
 sg13g2_inv_1 _7913_ (.Y(_2944_),
    .A(_2942_));
 sg13g2_nand3_1 _7914_ (.B(_2939_),
    .C(_2944_),
    .A(_2936_),
    .Y(_2945_));
 sg13g2_nand2_1 _7915_ (.Y(_2946_),
    .A(_2943_),
    .B(_2945_));
 sg13g2_nand2b_1 _7916_ (.Y(_2947_),
    .B(_2946_),
    .A_N(_2917_));
 sg13g2_nand3_1 _7917_ (.B(_2917_),
    .C(_2945_),
    .A(_2943_),
    .Y(_2948_));
 sg13g2_nand2_1 _7918_ (.Y(_2949_),
    .A(_2947_),
    .B(_2948_));
 sg13g2_nor2_1 _7919_ (.A(net23),
    .B(_2806_),
    .Y(_2950_));
 sg13g2_nand2_1 _7920_ (.Y(_2951_),
    .A(_2949_),
    .B(_2950_));
 sg13g2_inv_1 _7921_ (.Y(_2952_),
    .A(_2950_));
 sg13g2_nand3_1 _7922_ (.B(_2948_),
    .C(_2952_),
    .A(_2947_),
    .Y(_2953_));
 sg13g2_nand2_1 _7923_ (.Y(_2954_),
    .A(_2951_),
    .B(_2953_));
 sg13g2_nand2b_1 _7924_ (.Y(_2955_),
    .B(_2954_),
    .A_N(_2915_));
 sg13g2_buf_1 _7925_ (.A(_2955_),
    .X(_2956_));
 sg13g2_nand3_1 _7926_ (.B(_2953_),
    .C(_2915_),
    .A(_2951_),
    .Y(_2957_));
 sg13g2_nand2_1 _7927_ (.Y(_2958_),
    .A(_2956_),
    .B(_2957_));
 sg13g2_nor2_1 _7928_ (.A(_2913_),
    .B(_2958_),
    .Y(_2959_));
 sg13g2_inv_1 _7929_ (.Y(_2960_),
    .A(_2947_));
 sg13g2_a21oi_1 _7930_ (.A1(_2948_),
    .A2(_2950_),
    .Y(_2961_),
    .B1(_2960_));
 sg13g2_nor2_1 _7931_ (.A(net23),
    .B(_2797_),
    .Y(_2962_));
 sg13g2_inv_1 _7932_ (.Y(_2963_),
    .A(_2936_));
 sg13g2_a21oi_1 _7933_ (.A1(_2939_),
    .A2(_2942_),
    .Y(_2964_),
    .B1(_2963_));
 sg13g2_nand2_1 _7934_ (.Y(_2965_),
    .A(_2920_),
    .B(_2921_));
 sg13g2_o21ai_1 _7935_ (.B1(_2965_),
    .Y(_2966_),
    .A1(_2900_),
    .A2(_2806_));
 sg13g2_buf_1 _7936_ (.A(_2966_),
    .X(_2967_));
 sg13g2_inv_1 _7937_ (.Y(_2968_),
    .A(_2933_));
 sg13g2_a21oi_2 _7938_ (.B1(_2968_),
    .Y(_2969_),
    .A2(_2922_),
    .A1(_2931_));
 sg13g2_nand3_1 _7939_ (.B(_2845_),
    .C(_2777_),
    .A(_2844_),
    .Y(_2970_));
 sg13g2_buf_1 _7940_ (.A(_2970_),
    .X(_2971_));
 sg13g2_inv_2 _7941_ (.Y(_2972_),
    .A(_2881_));
 sg13g2_nand2_1 _7942_ (.Y(_2973_),
    .A(_2972_),
    .B(_2780_));
 sg13g2_xnor2_1 _7943_ (.Y(_2974_),
    .A(_2971_),
    .B(_2973_));
 sg13g2_inv_1 _7944_ (.Y(_2975_),
    .A(\generated._558[8] ));
 sg13g2_nor3_1 _7945_ (.A(_1909_),
    .B(\generated._558[7] ),
    .C(_2877_),
    .Y(_2976_));
 sg13g2_xnor2_1 _7946_ (.Y(_2977_),
    .A(_2975_),
    .B(_2976_));
 sg13g2_nand2_1 _7947_ (.Y(_2978_),
    .A(_2072_),
    .B(_2977_));
 sg13g2_nand2_1 _7948_ (.Y(_2979_),
    .A(_2058_),
    .B(_0666_));
 sg13g2_nand2_1 _7949_ (.Y(_2980_),
    .A(_2978_),
    .B(_2979_));
 sg13g2_buf_2 _7950_ (.A(_2980_),
    .X(_2981_));
 sg13g2_nor2_1 _7951_ (.A(_4295_),
    .B(_2981_),
    .Y(_2982_));
 sg13g2_nor2_1 _7952_ (.A(_2800_),
    .B(_2928_),
    .Y(_2983_));
 sg13g2_nand2_1 _7953_ (.Y(_2984_),
    .A(_2884_),
    .B(_2983_));
 sg13g2_xnor2_1 _7954_ (.Y(_2985_),
    .A(_2982_),
    .B(_2984_));
 sg13g2_xor2_1 _7955_ (.B(_2985_),
    .A(_2974_),
    .X(_2986_));
 sg13g2_xnor2_1 _7956_ (.Y(_2987_),
    .A(_2969_),
    .B(_2986_));
 sg13g2_xnor2_1 _7957_ (.Y(_2988_),
    .A(_2967_),
    .B(_2987_));
 sg13g2_nand2b_1 _7958_ (.Y(_2989_),
    .B(_2988_),
    .A_N(_2964_));
 sg13g2_xor2_1 _7959_ (.B(_2987_),
    .A(_2967_),
    .X(_2990_));
 sg13g2_nand2_1 _7960_ (.Y(_2991_),
    .A(_2990_),
    .B(_2964_));
 sg13g2_nand2_1 _7961_ (.Y(_2992_),
    .A(_2989_),
    .B(_2991_));
 sg13g2_xnor2_1 _7962_ (.Y(_2993_),
    .A(_2962_),
    .B(_2992_));
 sg13g2_nand2b_1 _7963_ (.Y(_2994_),
    .B(_2993_),
    .A_N(_2961_));
 sg13g2_buf_1 _7964_ (.A(_2994_),
    .X(_2995_));
 sg13g2_inv_1 _7965_ (.Y(_2996_),
    .A(_2962_));
 sg13g2_xnor2_1 _7966_ (.Y(_2997_),
    .A(_2996_),
    .B(_2992_));
 sg13g2_nand2_1 _7967_ (.Y(_2998_),
    .A(_2997_),
    .B(_2961_));
 sg13g2_nand2_1 _7968_ (.Y(_2999_),
    .A(_2995_),
    .B(_2998_));
 sg13g2_nand2_1 _7969_ (.Y(_3000_),
    .A(_2999_),
    .B(_2956_));
 sg13g2_nor2_1 _7970_ (.A(_2956_),
    .B(_2999_),
    .Y(_3001_));
 sg13g2_a21oi_1 _7971_ (.A1(_2959_),
    .A2(_3000_),
    .Y(_3002_),
    .B1(_3001_));
 sg13g2_a21oi_1 _7972_ (.A1(_2912_),
    .A2(_2910_),
    .Y(_3003_),
    .B1(_2871_));
 sg13g2_nand3_1 _7973_ (.B(_2867_),
    .C(_2834_),
    .A(_2866_),
    .Y(_3004_));
 sg13g2_a21oi_1 _7974_ (.A1(_2870_),
    .A2(_3004_),
    .Y(_3005_),
    .B1(_2774_));
 sg13g2_nand3_1 _7975_ (.B(_3004_),
    .C(_2774_),
    .A(_2870_),
    .Y(_3006_));
 sg13g2_xnor2_1 _7976_ (.Y(_3007_),
    .A(_2790_),
    .B(_2814_));
 sg13g2_nand2b_1 _7977_ (.Y(_3008_),
    .B(_3007_),
    .A_N(_2830_));
 sg13g2_nand2_1 _7978_ (.Y(_3009_),
    .A(_3008_),
    .B(_2831_));
 sg13g2_xor2_1 _7979_ (.B(_3009_),
    .A(_2832_),
    .X(_3010_));
 sg13g2_nand2b_1 _7980_ (.Y(_3011_),
    .B(_2825_),
    .A_N(_2829_));
 sg13g2_nand2b_1 _7981_ (.Y(_3012_),
    .B(_2828_),
    .A_N(_3011_));
 sg13g2_nor2_1 _7982_ (.A(_2809_),
    .B(_2823_),
    .Y(_3013_));
 sg13g2_inv_1 _7983_ (.Y(_3014_),
    .A(_2769_));
 sg13g2_nor2_1 _7984_ (.A(_3014_),
    .B(net22),
    .Y(_3015_));
 sg13g2_nor2_1 _7985_ (.A(_3015_),
    .B(_2824_),
    .Y(_3016_));
 sg13g2_nor2_1 _7986_ (.A(_0065_),
    .B(net79),
    .Y(_3017_));
 sg13g2_a22oi_1 _7987_ (.Y(_3018_),
    .B1(_3015_),
    .B2(_2824_),
    .A2(_3017_),
    .A1(_2823_));
 sg13g2_nor3_1 _7988_ (.A(_3013_),
    .B(_3016_),
    .C(_3018_),
    .Y(_3019_));
 sg13g2_nand2b_1 _7989_ (.Y(_3020_),
    .B(_3011_),
    .A_N(_2828_));
 sg13g2_nand3_1 _7990_ (.B(_3019_),
    .C(_3020_),
    .A(_3012_),
    .Y(_3021_));
 sg13g2_nor2_1 _7991_ (.A(_3014_),
    .B(net23),
    .Y(_3022_));
 sg13g2_nand2b_1 _7992_ (.Y(_3023_),
    .B(_3022_),
    .A_N(_3021_));
 sg13g2_nor2b_1 _7993_ (.A(_3022_),
    .B_N(_3021_),
    .Y(_3024_));
 sg13g2_a21oi_1 _7994_ (.A1(_3010_),
    .A2(_3023_),
    .Y(_3025_),
    .B1(_3024_));
 sg13g2_nand2_1 _7995_ (.Y(_3026_),
    .A(_3006_),
    .B(_3025_));
 sg13g2_nor2_1 _7996_ (.A(_3005_),
    .B(_3026_),
    .Y(_3027_));
 sg13g2_nand2_1 _7997_ (.Y(_3028_),
    .A(_2913_),
    .B(_3027_));
 sg13g2_nor2_1 _7998_ (.A(_3003_),
    .B(_3028_),
    .Y(_3029_));
 sg13g2_inv_1 _7999_ (.Y(_3030_),
    .A(_2958_));
 sg13g2_nand3_1 _8000_ (.B(_3030_),
    .C(_3000_),
    .A(_3029_),
    .Y(_3031_));
 sg13g2_nand2_1 _8001_ (.Y(_3032_),
    .A(_3002_),
    .B(_3031_));
 sg13g2_inv_1 _8002_ (.Y(_3033_),
    .A(_2989_));
 sg13g2_a21oi_1 _8003_ (.A1(_2991_),
    .A2(_2962_),
    .Y(_3034_),
    .B1(_3033_));
 sg13g2_nor2_1 _8004_ (.A(net23),
    .B(_2847_),
    .Y(_3035_));
 sg13g2_nor2_1 _8005_ (.A(_2900_),
    .B(_2797_),
    .Y(_3036_));
 sg13g2_xor2_1 _8006_ (.B(_3036_),
    .A(_3035_),
    .X(_3037_));
 sg13g2_nor3_2 _8007_ (.A(_2881_),
    .B(_2839_),
    .C(_2920_),
    .Y(_3038_));
 sg13g2_nor3_1 _8008_ (.A(_2800_),
    .B(_2981_),
    .C(_2929_),
    .Y(_3039_));
 sg13g2_nor2_1 _8009_ (.A(_2781_),
    .B(_2928_),
    .Y(_3040_));
 sg13g2_nand3_1 _8010_ (.B(_2924_),
    .C(_2975_),
    .A(_2925_),
    .Y(_3041_));
 sg13g2_xnor2_1 _8011_ (.Y(_3042_),
    .A(\generated._558[9] ),
    .B(_3041_));
 sg13g2_nand2_1 _8012_ (.Y(_3043_),
    .A(_2072_),
    .B(_3042_));
 sg13g2_nand2_1 _8013_ (.Y(_3044_),
    .A(_2058_),
    .B(_0687_));
 sg13g2_nand2_2 _8014_ (.Y(_3045_),
    .A(_3043_),
    .B(_3044_));
 sg13g2_nor2_1 _8015_ (.A(_4295_),
    .B(_3045_),
    .Y(_3046_));
 sg13g2_xor2_1 _8016_ (.B(_3046_),
    .A(_3040_),
    .X(_3047_));
 sg13g2_xnor2_1 _8017_ (.Y(_3048_),
    .A(_3039_),
    .B(_3047_));
 sg13g2_nand4_1 _8018_ (.B(_2972_),
    .C(net94),
    .A(_2983_),
    .Y(_3049_),
    .D(_2981_));
 sg13g2_nand2b_1 _8019_ (.Y(_3050_),
    .B(_2985_),
    .A_N(_2974_));
 sg13g2_nand3_1 _8020_ (.B(_3049_),
    .C(_3050_),
    .A(_3048_),
    .Y(_3051_));
 sg13g2_nand2_1 _8021_ (.Y(_3052_),
    .A(_3050_),
    .B(_3049_));
 sg13g2_nand2b_1 _8022_ (.Y(_3053_),
    .B(_3052_),
    .A_N(_3048_));
 sg13g2_nand2_1 _8023_ (.Y(_3054_),
    .A(_3051_),
    .B(_3053_));
 sg13g2_xor2_1 _8024_ (.B(_3054_),
    .A(_3038_),
    .X(_3055_));
 sg13g2_nand2_1 _8025_ (.Y(_3056_),
    .A(_2986_),
    .B(_2969_));
 sg13g2_nor2_1 _8026_ (.A(_2969_),
    .B(_2986_),
    .Y(_3057_));
 sg13g2_a21oi_1 _8027_ (.A1(_3056_),
    .A2(_2967_),
    .Y(_3058_),
    .B1(_3057_));
 sg13g2_nand2_1 _8028_ (.Y(_3059_),
    .A(_3055_),
    .B(_3058_));
 sg13g2_xnor2_1 _8029_ (.Y(_3060_),
    .A(_3038_),
    .B(_3054_));
 sg13g2_nand2b_1 _8030_ (.Y(_3061_),
    .B(_3060_),
    .A_N(_3058_));
 sg13g2_nand2_1 _8031_ (.Y(_3062_),
    .A(_3059_),
    .B(_3061_));
 sg13g2_xnor2_1 _8032_ (.Y(_3063_),
    .A(_3037_),
    .B(_3062_));
 sg13g2_xor2_1 _8033_ (.B(_3063_),
    .A(_3034_),
    .X(_3064_));
 sg13g2_xnor2_1 _8034_ (.Y(_3065_),
    .A(_2995_),
    .B(_3064_));
 sg13g2_inv_1 _8035_ (.Y(_3066_),
    .A(_3036_));
 sg13g2_inv_1 _8036_ (.Y(_3067_),
    .A(_3035_));
 sg13g2_nor2_1 _8037_ (.A(_3066_),
    .B(_3067_),
    .Y(_3068_));
 sg13g2_inv_1 _8038_ (.Y(_3069_),
    .A(_3061_));
 sg13g2_a21oi_1 _8039_ (.A1(_3059_),
    .A2(_3037_),
    .Y(_3070_),
    .B1(_3069_));
 sg13g2_nor2_1 _8040_ (.A(net23),
    .B(_2881_),
    .Y(_3071_));
 sg13g2_inv_1 _8041_ (.Y(_3072_),
    .A(_3071_));
 sg13g2_nor2_1 _8042_ (.A(_2971_),
    .B(_2973_),
    .Y(_3073_));
 sg13g2_xnor2_1 _8043_ (.Y(_3074_),
    .A(_3072_),
    .B(_3073_));
 sg13g2_nor2_1 _8044_ (.A(_2900_),
    .B(_2847_),
    .Y(_3075_));
 sg13g2_nor2_2 _8045_ (.A(net22),
    .B(_3045_),
    .Y(_3076_));
 sg13g2_nand2_1 _8046_ (.Y(_3077_),
    .A(_3076_),
    .B(_2929_));
 sg13g2_xnor2_1 _8047_ (.Y(_3078_),
    .A(_3075_),
    .B(_3077_));
 sg13g2_nand2_1 _8048_ (.Y(_3079_),
    .A(_3047_),
    .B(_3039_));
 sg13g2_nand2_1 _8049_ (.Y(_3080_),
    .A(_2982_),
    .B(_2983_));
 sg13g2_nand2_1 _8050_ (.Y(_3081_),
    .A(_3079_),
    .B(_3080_));
 sg13g2_inv_4 _8051_ (.A(_3045_),
    .Y(_3082_));
 sg13g2_nand2_1 _8052_ (.Y(_3083_),
    .A(_2800_),
    .B(_4294_));
 sg13g2_nand2_1 _8053_ (.Y(_3084_),
    .A(_3082_),
    .B(_3083_));
 sg13g2_nand2b_1 _8054_ (.Y(_3085_),
    .B(_4293_),
    .A_N(_2757_));
 sg13g2_nor2b_1 _8055_ (.A(_3084_),
    .B_N(_3085_),
    .Y(_3086_));
 sg13g2_nand3_1 _8056_ (.B(_2927_),
    .C(_2777_),
    .A(_2923_),
    .Y(_3087_));
 sg13g2_o21ai_1 _8057_ (.B1(_3087_),
    .Y(_3088_),
    .A1(_2781_),
    .A2(_2981_));
 sg13g2_nor2_1 _8058_ (.A(_2839_),
    .B(_2981_),
    .Y(_3089_));
 sg13g2_nand2_1 _8059_ (.Y(_3090_),
    .A(_3089_),
    .B(_3040_));
 sg13g2_nand2_1 _8060_ (.Y(_3091_),
    .A(_3088_),
    .B(_3090_));
 sg13g2_xnor2_1 _8061_ (.Y(_3092_),
    .A(_3086_),
    .B(_3091_));
 sg13g2_inv_1 _8062_ (.Y(_3093_),
    .A(_3092_));
 sg13g2_nand2b_1 _8063_ (.Y(_3094_),
    .B(_3093_),
    .A_N(_3081_));
 sg13g2_nand2_1 _8064_ (.Y(_3095_),
    .A(_3092_),
    .B(_3081_));
 sg13g2_nand2_1 _8065_ (.Y(_3096_),
    .A(_3094_),
    .B(_3095_));
 sg13g2_xor2_1 _8066_ (.B(_3096_),
    .A(_3078_),
    .X(_3097_));
 sg13g2_inv_1 _8067_ (.Y(_3098_),
    .A(_3053_));
 sg13g2_a21oi_1 _8068_ (.A1(_3051_),
    .A2(_3038_),
    .Y(_3099_),
    .B1(_3098_));
 sg13g2_nand2_1 _8069_ (.Y(_3100_),
    .A(_3097_),
    .B(_3099_));
 sg13g2_xnor2_1 _8070_ (.Y(_3101_),
    .A(_3078_),
    .B(_3096_));
 sg13g2_nand2b_1 _8071_ (.Y(_3102_),
    .B(_3101_),
    .A_N(_3099_));
 sg13g2_nand2_1 _8072_ (.Y(_3103_),
    .A(_3100_),
    .B(_3102_));
 sg13g2_xnor2_1 _8073_ (.Y(_3104_),
    .A(_3074_),
    .B(_3103_));
 sg13g2_nand2b_1 _8074_ (.Y(_3105_),
    .B(_3104_),
    .A_N(_3070_));
 sg13g2_inv_1 _8075_ (.Y(_3106_),
    .A(_3074_));
 sg13g2_nand2_1 _8076_ (.Y(_3107_),
    .A(_3103_),
    .B(_3106_));
 sg13g2_nand3_1 _8077_ (.B(_3102_),
    .C(_3074_),
    .A(_3100_),
    .Y(_3108_));
 sg13g2_nand2_1 _8078_ (.Y(_3109_),
    .A(_3107_),
    .B(_3108_));
 sg13g2_nand2_1 _8079_ (.Y(_3110_),
    .A(_3109_),
    .B(_3070_));
 sg13g2_nand2_1 _8080_ (.Y(_3111_),
    .A(_3105_),
    .B(_3110_));
 sg13g2_nand2b_1 _8081_ (.Y(_3112_),
    .B(_3111_),
    .A_N(_3068_));
 sg13g2_nand3_1 _8082_ (.B(_3110_),
    .C(_3068_),
    .A(_3105_),
    .Y(_3113_));
 sg13g2_nand2_1 _8083_ (.Y(_3114_),
    .A(_3112_),
    .B(_3113_));
 sg13g2_nand2b_1 _8084_ (.Y(_3115_),
    .B(_3063_),
    .A_N(_3034_));
 sg13g2_nand2_1 _8085_ (.Y(_3116_),
    .A(_3114_),
    .B(_3115_));
 sg13g2_inv_1 _8086_ (.Y(_3117_),
    .A(_3115_));
 sg13g2_nand3_1 _8087_ (.B(_3113_),
    .C(_3117_),
    .A(_3112_),
    .Y(_3118_));
 sg13g2_nand2_1 _8088_ (.Y(_3119_),
    .A(_3116_),
    .B(_3118_));
 sg13g2_nor2_1 _8089_ (.A(_3065_),
    .B(_3119_),
    .Y(_3120_));
 sg13g2_nand2_1 _8090_ (.Y(_3121_),
    .A(_3032_),
    .B(_3120_));
 sg13g2_nor2_1 _8091_ (.A(_2995_),
    .B(_3064_),
    .Y(_3122_));
 sg13g2_nand2_1 _8092_ (.Y(_3123_),
    .A(_3116_),
    .B(_3122_));
 sg13g2_nand2_1 _8093_ (.Y(_3124_),
    .A(_3123_),
    .B(_3118_));
 sg13g2_inv_1 _8094_ (.Y(_3125_),
    .A(_3124_));
 sg13g2_nand2_1 _8095_ (.Y(_3126_),
    .A(_3121_),
    .B(_3125_));
 sg13g2_inv_1 _8096_ (.Y(_3127_),
    .A(_3105_));
 sg13g2_a21oi_1 _8097_ (.A1(_3110_),
    .A2(_3068_),
    .Y(_3128_),
    .B1(_3127_));
 sg13g2_nor3_2 _8098_ (.A(_2971_),
    .B(_2973_),
    .C(_3072_),
    .Y(_3129_));
 sg13g2_inv_1 _8099_ (.Y(_3130_),
    .A(_3102_));
 sg13g2_a21oi_1 _8100_ (.A1(_3100_),
    .A2(_3074_),
    .Y(_3131_),
    .B1(_3130_));
 sg13g2_nor2_1 _8101_ (.A(net23),
    .B(_2928_),
    .Y(_3132_));
 sg13g2_inv_1 _8102_ (.Y(_3133_),
    .A(_3132_));
 sg13g2_nor2b_1 _8103_ (.A(_3077_),
    .B_N(_3075_),
    .Y(_3134_));
 sg13g2_xnor2_1 _8104_ (.Y(_3135_),
    .A(_3133_),
    .B(_3134_));
 sg13g2_o21ai_1 _8105_ (.B1(_3090_),
    .Y(_3136_),
    .A1(_2881_),
    .A2(_2900_));
 sg13g2_xnor2_1 _8106_ (.Y(_3137_),
    .A(_3076_),
    .B(_3089_));
 sg13g2_buf_2 _8107_ (.A(_3137_),
    .X(_3138_));
 sg13g2_nand3_1 _8108_ (.B(_3088_),
    .C(_3090_),
    .A(_3086_),
    .Y(_3139_));
 sg13g2_inv_1 _8109_ (.Y(_3140_),
    .A(_3084_));
 sg13g2_nand2_1 _8110_ (.Y(_3141_),
    .A(_3139_),
    .B(_3140_));
 sg13g2_xnor2_1 _8111_ (.Y(_3142_),
    .A(_3138_),
    .B(_3141_));
 sg13g2_xnor2_1 _8112_ (.Y(_3143_),
    .A(_3136_),
    .B(_3142_));
 sg13g2_inv_1 _8113_ (.Y(_3144_),
    .A(_3143_));
 sg13g2_inv_1 _8114_ (.Y(_3145_),
    .A(_3095_));
 sg13g2_a21oi_1 _8115_ (.A1(_3094_),
    .A2(_3078_),
    .Y(_3146_),
    .B1(_3145_));
 sg13g2_nand2_1 _8116_ (.Y(_3147_),
    .A(_3144_),
    .B(_3146_));
 sg13g2_nand2b_1 _8117_ (.Y(_3148_),
    .B(_3143_),
    .A_N(_3146_));
 sg13g2_nand2_1 _8118_ (.Y(_3149_),
    .A(_3147_),
    .B(_3148_));
 sg13g2_xnor2_1 _8119_ (.Y(_3150_),
    .A(_3135_),
    .B(_3149_));
 sg13g2_nand2b_1 _8120_ (.Y(_3151_),
    .B(_3150_),
    .A_N(_3131_));
 sg13g2_nand2b_1 _8121_ (.Y(_3152_),
    .B(_3149_),
    .A_N(_3135_));
 sg13g2_nand3_1 _8122_ (.B(_3148_),
    .C(_3135_),
    .A(_3147_),
    .Y(_3153_));
 sg13g2_nand2_1 _8123_ (.Y(_3154_),
    .A(_3152_),
    .B(_3153_));
 sg13g2_nand2_1 _8124_ (.Y(_3155_),
    .A(_3154_),
    .B(_3131_));
 sg13g2_nand2_1 _8125_ (.Y(_3156_),
    .A(_3151_),
    .B(_3155_));
 sg13g2_xnor2_1 _8126_ (.Y(_3157_),
    .A(_3129_),
    .B(_3156_));
 sg13g2_nand2b_1 _8127_ (.Y(_3158_),
    .B(_3157_),
    .A_N(_3128_));
 sg13g2_nand2b_1 _8128_ (.Y(_3159_),
    .B(_3156_),
    .A_N(_3129_));
 sg13g2_nand3_1 _8129_ (.B(_3155_),
    .C(_3129_),
    .A(_3151_),
    .Y(_3160_));
 sg13g2_nand2_1 _8130_ (.Y(_3161_),
    .A(_3159_),
    .B(_3160_));
 sg13g2_nand2_1 _8131_ (.Y(_3162_),
    .A(_3161_),
    .B(_3128_));
 sg13g2_nand2_2 _8132_ (.Y(_3163_),
    .A(_3158_),
    .B(_3162_));
 sg13g2_nand2_1 _8133_ (.Y(_3164_),
    .A(_3126_),
    .B(_3163_));
 sg13g2_inv_1 _8134_ (.Y(_3165_),
    .A(_3163_));
 sg13g2_nand3_1 _8135_ (.B(_3165_),
    .C(_3125_),
    .A(_3121_),
    .Y(_3166_));
 sg13g2_nand2_1 _8136_ (.Y(_3167_),
    .A(_3164_),
    .B(_3166_));
 sg13g2_nand3_1 _8137_ (.B(_2752_),
    .C(_3167_),
    .A(_2751_),
    .Y(_3168_));
 sg13g2_nand2_1 _8138_ (.Y(_3169_),
    .A(_2700_),
    .B(_2749_));
 sg13g2_nand3_1 _8139_ (.B(_2750_),
    .C(_2699_),
    .A(_2692_),
    .Y(_3170_));
 sg13g2_nand2_1 _8140_ (.Y(_3171_),
    .A(_3126_),
    .B(_3165_));
 sg13g2_nand3_1 _8141_ (.B(_3163_),
    .C(_3125_),
    .A(_3121_),
    .Y(_3172_));
 sg13g2_nand2_1 _8142_ (.Y(_3173_),
    .A(_3171_),
    .B(_3172_));
 sg13g2_nand3_1 _8143_ (.B(_3170_),
    .C(_3173_),
    .A(_3169_),
    .Y(_3174_));
 sg13g2_nand2_1 _8144_ (.Y(_3175_),
    .A(_3168_),
    .B(_3174_));
 sg13g2_nand2_1 _8145_ (.Y(_3176_),
    .A(_3029_),
    .B(_3030_));
 sg13g2_nand2b_1 _8146_ (.Y(_3177_),
    .B(_3176_),
    .A_N(_2959_));
 sg13g2_xnor2_1 _8147_ (.Y(_3178_),
    .A(_2956_),
    .B(_2999_));
 sg13g2_nor2_1 _8148_ (.A(_3065_),
    .B(_3178_),
    .Y(_3179_));
 sg13g2_nand2_1 _8149_ (.Y(_3180_),
    .A(_3177_),
    .B(_3179_));
 sg13g2_nand2_1 _8150_ (.Y(_3181_),
    .A(_3064_),
    .B(_2995_));
 sg13g2_a21oi_1 _8151_ (.A1(_3001_),
    .A2(_3181_),
    .Y(_3182_),
    .B1(_3122_));
 sg13g2_nand2_1 _8152_ (.Y(_3183_),
    .A(_3180_),
    .B(_3182_));
 sg13g2_inv_1 _8153_ (.Y(_3184_),
    .A(_3119_));
 sg13g2_nand2_1 _8154_ (.Y(_3185_),
    .A(_3183_),
    .B(_3184_));
 sg13g2_nand3_1 _8155_ (.B(_3182_),
    .C(_3119_),
    .A(_3180_),
    .Y(_3186_));
 sg13g2_nand2_1 _8156_ (.Y(_3187_),
    .A(_3185_),
    .B(_3186_));
 sg13g2_nand2_1 _8157_ (.Y(_3188_),
    .A(_2648_),
    .B(_2694_));
 sg13g2_inv_1 _8158_ (.Y(_3189_),
    .A(_2518_));
 sg13g2_nand2_1 _8159_ (.Y(_3190_),
    .A(_2684_),
    .B(_3189_));
 sg13g2_nand2_1 _8160_ (.Y(_3191_),
    .A(_3190_),
    .B(_2519_));
 sg13g2_nor2_1 _8161_ (.A(_3188_),
    .B(_3191_),
    .Y(_3192_));
 sg13g2_nand2_1 _8162_ (.Y(_3193_),
    .A(_2687_),
    .B(_2690_));
 sg13g2_nand2_1 _8163_ (.Y(_3194_),
    .A(_3192_),
    .B(_3193_));
 sg13g2_inv_1 _8164_ (.Y(_3195_),
    .A(_2648_));
 sg13g2_a21oi_1 _8165_ (.A1(_3190_),
    .A2(_2694_),
    .Y(_3196_),
    .B1(_3195_));
 sg13g2_inv_1 _8166_ (.Y(_3197_),
    .A(_3196_));
 sg13g2_nand2_1 _8167_ (.Y(_3198_),
    .A(_3194_),
    .B(_3197_));
 sg13g2_nand2_1 _8168_ (.Y(_3199_),
    .A(_3198_),
    .B(_2695_));
 sg13g2_nand3_1 _8169_ (.B(_3197_),
    .C(_2644_),
    .A(_3194_),
    .Y(_3200_));
 sg13g2_nand2_1 _8170_ (.Y(_3201_),
    .A(_3199_),
    .B(_3200_));
 sg13g2_nand2b_2 _8171_ (.Y(_3202_),
    .B(_3201_),
    .A_N(_3187_));
 sg13g2_nand2_1 _8172_ (.Y(_3203_),
    .A(_3175_),
    .B(_3202_));
 sg13g2_nand3_1 _8173_ (.B(_3200_),
    .C(_3187_),
    .A(_3199_),
    .Y(_3204_));
 sg13g2_nor3_1 _8174_ (.A(\generated._402[2] ),
    .B(_4247_),
    .C(_4251_),
    .Y(_3205_));
 sg13g2_nand2_1 _8175_ (.Y(_3206_),
    .A(_3205_),
    .B(_4229_));
 sg13g2_nor2_1 _8176_ (.A(_4253_),
    .B(_3206_),
    .Y(_3207_));
 sg13g2_nand2b_1 _8177_ (.Y(_3208_),
    .B(_3207_),
    .A_N(_0968_));
 sg13g2_nor2_1 _8178_ (.A(_0971_),
    .B(_3208_),
    .Y(_3209_));
 sg13g2_inv_1 _8179_ (.Y(_3210_),
    .A(_3209_));
 sg13g2_nor2_1 _8180_ (.A(_1001_),
    .B(_3210_),
    .Y(_3211_));
 sg13g2_inv_1 _8181_ (.Y(_3212_),
    .A(_3211_));
 sg13g2_nand2_1 _8182_ (.Y(_3213_),
    .A(_3212_),
    .B(_1003_));
 sg13g2_nand2_1 _8183_ (.Y(_3214_),
    .A(_3211_),
    .B(_1004_));
 sg13g2_nand2_1 _8184_ (.Y(_3215_),
    .A(_3213_),
    .B(_3214_));
 sg13g2_inv_1 _8185_ (.Y(_3216_),
    .A(_3215_));
 sg13g2_nor2_1 _8186_ (.A(_0442_),
    .B(_0439_),
    .Y(_3217_));
 sg13g2_inv_1 _8187_ (.Y(_3218_),
    .A(_3217_));
 sg13g2_nand2_1 _8188_ (.Y(_3219_),
    .A(_3218_),
    .B(_0457_));
 sg13g2_nor2_1 _8189_ (.A(_0457_),
    .B(_3218_),
    .Y(_3220_));
 sg13g2_nor2_1 _8190_ (.A(net88),
    .B(_3220_),
    .Y(_3221_));
 sg13g2_a22oi_1 _8191_ (.Y(_3222_),
    .B1(_3219_),
    .B2(_3221_),
    .A2(net88),
    .A1(_0291_));
 sg13g2_buf_1 _8192_ (.A(_3222_),
    .X(_3223_));
 sg13g2_inv_1 _8193_ (.Y(_3224_),
    .A(_3223_));
 sg13g2_nand2_1 _8194_ (.Y(_3225_),
    .A(net15),
    .B(_3224_));
 sg13g2_nand2_1 _8195_ (.Y(_3226_),
    .A(_3210_),
    .B(_1001_));
 sg13g2_nand2_1 _8196_ (.Y(_3227_),
    .A(_3212_),
    .B(_3226_));
 sg13g2_buf_2 _8197_ (.A(_3227_),
    .X(_3228_));
 sg13g2_inv_2 _8198_ (.Y(_3229_),
    .A(_3228_));
 sg13g2_inv_1 _8199_ (.Y(_3230_),
    .A(_0286_));
 sg13g2_nor3_1 _8200_ (.A(_0442_),
    .B(_0457_),
    .C(_3230_),
    .Y(_3231_));
 sg13g2_xnor2_1 _8201_ (.Y(_3232_),
    .A(_0474_),
    .B(_3231_));
 sg13g2_nand2_1 _8202_ (.Y(_3233_),
    .A(_0309_),
    .B(net88));
 sg13g2_o21ai_1 _8203_ (.B1(_3233_),
    .Y(_3234_),
    .A1(net88),
    .A2(_3232_));
 sg13g2_buf_2 _8204_ (.A(_3234_),
    .X(_3235_));
 sg13g2_nand2_1 _8205_ (.Y(_3236_),
    .A(_3229_),
    .B(_3235_));
 sg13g2_nand2_1 _8206_ (.Y(_3237_),
    .A(_3225_),
    .B(_3236_));
 sg13g2_nand2_1 _8207_ (.Y(_3238_),
    .A(_0442_),
    .B(_0439_));
 sg13g2_nor2_1 _8208_ (.A(net88),
    .B(_3217_),
    .Y(_3239_));
 sg13g2_a22oi_1 _8209_ (.Y(_3240_),
    .B1(_3238_),
    .B2(_3239_),
    .A2(net88),
    .A1(_0467_));
 sg13g2_buf_1 _8210_ (.A(_3240_),
    .X(_3241_));
 sg13g2_nand3_1 _8211_ (.B(_0934_),
    .C(\generated._75[0] ),
    .A(_3205_),
    .Y(_3242_));
 sg13g2_o21ai_1 _8212_ (.B1(_1023_),
    .Y(_3243_),
    .A1(_1003_),
    .A2(_3242_));
 sg13g2_buf_1 _8213_ (.A(_3243_),
    .X(_3244_));
 sg13g2_inv_2 _8214_ (.Y(_3245_),
    .A(_3244_));
 sg13g2_nor2_1 _8215_ (.A(_3241_),
    .B(_3245_),
    .Y(_3246_));
 sg13g2_nor2_1 _8216_ (.A(_3236_),
    .B(_3225_),
    .Y(_3247_));
 sg13g2_a21oi_1 _8217_ (.A1(_3237_),
    .A2(_3246_),
    .Y(_3248_),
    .B1(_3247_));
 sg13g2_nand2_1 _8218_ (.Y(_3249_),
    .A(_3208_),
    .B(_0971_));
 sg13g2_nand2_1 _8219_ (.Y(_3250_),
    .A(_3210_),
    .B(_3249_));
 sg13g2_buf_1 _8220_ (.A(_3250_),
    .X(_3251_));
 sg13g2_inv_1 _8221_ (.Y(_3252_),
    .A(_3251_));
 sg13g2_inv_1 _8222_ (.Y(_3253_),
    .A(_3220_));
 sg13g2_nor3_1 _8223_ (.A(\generated._377[2] ),
    .B(\generated._377[3] ),
    .C(_3253_),
    .Y(_3254_));
 sg13g2_o21ai_1 _8224_ (.B1(\generated._377[3] ),
    .Y(_3255_),
    .A1(\generated._377[2] ),
    .A2(_3253_));
 sg13g2_nand3b_1 _8225_ (.B(_1492_),
    .C(_3255_),
    .Y(_3256_),
    .A_N(_3254_));
 sg13g2_o21ai_1 _8226_ (.B1(_3256_),
    .Y(_3257_),
    .A1(net68),
    .A2(_0090_));
 sg13g2_buf_2 _8227_ (.A(_3257_),
    .X(_3258_));
 sg13g2_nand2_1 _8228_ (.Y(_3259_),
    .A(net17),
    .B(_3258_));
 sg13g2_nand2_1 _8229_ (.Y(_3260_),
    .A(_3254_),
    .B(_0503_));
 sg13g2_a21oi_1 _8230_ (.A1(_3260_),
    .A2(_0518_),
    .Y(_3261_),
    .B1(_4489_));
 sg13g2_nor2_1 _8231_ (.A(_0518_),
    .B(_3260_),
    .Y(_3262_));
 sg13g2_inv_1 _8232_ (.Y(_3263_),
    .A(_3262_));
 sg13g2_nand2_1 _8233_ (.Y(_3264_),
    .A(_3261_),
    .B(_3263_));
 sg13g2_o21ai_1 _8234_ (.B1(_3264_),
    .Y(_3265_),
    .A1(net68),
    .A2(_0092_));
 sg13g2_buf_2 _8235_ (.A(_3265_),
    .X(_3266_));
 sg13g2_xnor2_1 _8236_ (.Y(_3267_),
    .A(_3206_),
    .B(_0935_));
 sg13g2_buf_2 _8237_ (.A(_3267_),
    .X(_3268_));
 sg13g2_inv_1 _8238_ (.Y(_3269_),
    .A(_3231_));
 sg13g2_nor2_1 _8239_ (.A(\generated._377[2] ),
    .B(_3269_),
    .Y(_3270_));
 sg13g2_a21oi_1 _8240_ (.A1(_3270_),
    .A2(_0489_),
    .Y(_3271_),
    .B1(_0503_));
 sg13g2_nand3_1 _8241_ (.B(_0489_),
    .C(_0503_),
    .A(_3270_),
    .Y(_3272_));
 sg13g2_nand3b_1 _8242_ (.B(_1492_),
    .C(_3272_),
    .Y(_3273_),
    .A_N(_3271_));
 sg13g2_o21ai_1 _8243_ (.B1(_3273_),
    .Y(_3274_),
    .A1(_1492_),
    .A2(_0091_));
 sg13g2_buf_1 _8244_ (.A(_3274_),
    .X(_3275_));
 sg13g2_inv_1 _8245_ (.Y(_3276_),
    .A(_3242_));
 sg13g2_xnor2_1 _8246_ (.Y(_3277_),
    .A(_3276_),
    .B(_0968_));
 sg13g2_buf_1 _8247_ (.A(_3277_),
    .X(_3278_));
 sg13g2_nand2_1 _8248_ (.Y(_3279_),
    .A(_3275_),
    .B(net30));
 sg13g2_inv_1 _8249_ (.Y(_3280_),
    .A(_3279_));
 sg13g2_a21oi_1 _8250_ (.A1(_3266_),
    .A2(_3268_),
    .Y(_3281_),
    .B1(_3280_));
 sg13g2_nand3_1 _8251_ (.B(_3266_),
    .C(_3268_),
    .A(_3280_),
    .Y(_3282_));
 sg13g2_nand2b_1 _8252_ (.Y(_3283_),
    .B(_3282_),
    .A_N(_3281_));
 sg13g2_xnor2_1 _8253_ (.Y(_3284_),
    .A(_3259_),
    .B(_3283_));
 sg13g2_a22oi_1 _8254_ (.Y(_3285_),
    .B1(_3268_),
    .B2(_3275_),
    .A2(_3258_),
    .A1(net30));
 sg13g2_nand2_1 _8255_ (.Y(_3286_),
    .A(_3252_),
    .B(_3235_));
 sg13g2_inv_1 _8256_ (.Y(_3287_),
    .A(_3268_));
 sg13g2_nor2b_1 _8257_ (.A(_3287_),
    .B_N(_3258_),
    .Y(_3288_));
 sg13g2_nand2_1 _8258_ (.Y(_3289_),
    .A(_3280_),
    .B(_3288_));
 sg13g2_o21ai_1 _8259_ (.B1(_3289_),
    .Y(_3290_),
    .A1(_3285_),
    .A2(_3286_));
 sg13g2_nor2b_1 _8260_ (.A(_3284_),
    .B_N(_3290_),
    .Y(_3291_));
 sg13g2_xnor2_1 _8261_ (.Y(_3292_),
    .A(_3236_),
    .B(_3225_));
 sg13g2_xor2_1 _8262_ (.B(_3292_),
    .A(_3246_),
    .X(_3293_));
 sg13g2_xnor2_1 _8263_ (.Y(_3294_),
    .A(_3290_),
    .B(_3284_));
 sg13g2_nor2b_1 _8264_ (.A(_3293_),
    .B_N(_3294_),
    .Y(_3295_));
 sg13g2_nor2_1 _8265_ (.A(_3291_),
    .B(_3295_),
    .Y(_3296_));
 sg13g2_o21ai_1 _8266_ (.B1(_3282_),
    .Y(_3297_),
    .A1(_3259_),
    .A2(_3281_));
 sg13g2_nand2_1 _8267_ (.Y(_3298_),
    .A(net17),
    .B(_3275_));
 sg13g2_nand2_1 _8268_ (.Y(_3299_),
    .A(_3266_),
    .B(net30));
 sg13g2_o21ai_1 _8269_ (.B1(_0530_),
    .Y(_3300_),
    .A1(_0518_),
    .A2(_3272_));
 sg13g2_nor2_1 _8270_ (.A(_0518_),
    .B(_3272_),
    .Y(_3301_));
 sg13g2_nand2b_1 _8271_ (.Y(_3302_),
    .B(_3301_),
    .A_N(_0530_));
 sg13g2_nand3_1 _8272_ (.B(_3302_),
    .C(_1492_),
    .A(_3300_),
    .Y(_3303_));
 sg13g2_o21ai_1 _8273_ (.B1(_3303_),
    .Y(_3304_),
    .A1(_1492_),
    .A2(_0354_));
 sg13g2_buf_2 _8274_ (.A(_3304_),
    .X(_3305_));
 sg13g2_nand2_1 _8275_ (.Y(_3306_),
    .A(_3305_),
    .B(_3268_));
 sg13g2_xnor2_1 _8276_ (.Y(_3307_),
    .A(_3299_),
    .B(_3306_));
 sg13g2_xnor2_1 _8277_ (.Y(_3308_),
    .A(_3298_),
    .B(_3307_));
 sg13g2_xnor2_1 _8278_ (.Y(_3309_),
    .A(_3297_),
    .B(_3308_));
 sg13g2_nor2_1 _8279_ (.A(_3223_),
    .B(_3245_),
    .Y(_3310_));
 sg13g2_nand2_2 _8280_ (.Y(_3311_),
    .A(_3229_),
    .B(_3258_));
 sg13g2_nand2_1 _8281_ (.Y(_3312_),
    .A(net15),
    .B(_3235_));
 sg13g2_xnor2_1 _8282_ (.Y(_3313_),
    .A(_3311_),
    .B(_3312_));
 sg13g2_xor2_1 _8283_ (.B(_3313_),
    .A(_3310_),
    .X(_3314_));
 sg13g2_xor2_1 _8284_ (.B(_3314_),
    .A(_3309_),
    .X(_3315_));
 sg13g2_xnor2_1 _8285_ (.Y(_3316_),
    .A(_3296_),
    .B(_3315_));
 sg13g2_xnor2_1 _8286_ (.Y(_3317_),
    .A(_3248_),
    .B(_3316_));
 sg13g2_nor2_1 _8287_ (.A(_3223_),
    .B(_3228_),
    .Y(_3318_));
 sg13g2_nor2_1 _8288_ (.A(_3241_),
    .B(_3215_),
    .Y(_3319_));
 sg13g2_xnor2_1 _8289_ (.Y(_3320_),
    .A(_3318_),
    .B(_3319_));
 sg13g2_nor2_1 _8290_ (.A(_0440_),
    .B(_3245_),
    .Y(_3321_));
 sg13g2_nor2b_1 _8291_ (.A(_3320_),
    .B_N(_3321_),
    .Y(_3322_));
 sg13g2_a21oi_1 _8292_ (.A1(_3318_),
    .A2(_3319_),
    .Y(_3323_),
    .B1(_3322_));
 sg13g2_xnor2_1 _8293_ (.Y(_3324_),
    .A(_3294_),
    .B(_3293_));
 sg13g2_xor2_1 _8294_ (.B(_3320_),
    .A(_3321_),
    .X(_3325_));
 sg13g2_nand2_1 _8295_ (.Y(_3326_),
    .A(net17),
    .B(_3224_));
 sg13g2_nand2_1 _8296_ (.Y(_3327_),
    .A(net30),
    .B(_3235_));
 sg13g2_xor2_1 _8297_ (.B(_3288_),
    .A(_3327_),
    .X(_3328_));
 sg13g2_nand2b_1 _8298_ (.Y(_3329_),
    .B(_3288_),
    .A_N(_3327_));
 sg13g2_o21ai_1 _8299_ (.B1(_3329_),
    .Y(_3330_),
    .A1(_3326_),
    .A2(_3328_));
 sg13g2_nand2b_1 _8300_ (.Y(_3331_),
    .B(_3289_),
    .A_N(_3285_));
 sg13g2_xnor2_1 _8301_ (.Y(_3332_),
    .A(_3286_),
    .B(_3331_));
 sg13g2_xnor2_1 _8302_ (.Y(_3333_),
    .A(_3330_),
    .B(_3332_));
 sg13g2_nand2b_1 _8303_ (.Y(_3334_),
    .B(_3333_),
    .A_N(_3325_));
 sg13g2_nand2b_1 _8304_ (.Y(_3335_),
    .B(_3330_),
    .A_N(_3332_));
 sg13g2_nand2_1 _8305_ (.Y(_3336_),
    .A(_3334_),
    .B(_3335_));
 sg13g2_xnor2_1 _8306_ (.Y(_3337_),
    .A(_3324_),
    .B(_3336_));
 sg13g2_nand2_1 _8307_ (.Y(_3338_),
    .A(_3336_),
    .B(_3324_));
 sg13g2_o21ai_1 _8308_ (.B1(_3338_),
    .Y(_3339_),
    .A1(_3323_),
    .A2(_3337_));
 sg13g2_nor2b_1 _8309_ (.A(_3317_),
    .B_N(_3339_),
    .Y(_3340_));
 sg13g2_nor2b_1 _8310_ (.A(_3339_),
    .B_N(_3317_),
    .Y(_3341_));
 sg13g2_nand2_1 _8311_ (.Y(_3342_),
    .A(net15),
    .B(_0439_));
 sg13g2_nor2_1 _8312_ (.A(_3241_),
    .B(_3228_),
    .Y(_3343_));
 sg13g2_nor2b_1 _8313_ (.A(_3342_),
    .B_N(_3343_),
    .Y(_3344_));
 sg13g2_a22oi_1 _8314_ (.Y(_3345_),
    .B1(_3224_),
    .B2(net30),
    .A2(_3235_),
    .A1(_3268_));
 sg13g2_nand2b_1 _8315_ (.Y(_3346_),
    .B(net17),
    .A_N(_3241_));
 sg13g2_nor2_1 _8316_ (.A(_3223_),
    .B(_3287_),
    .Y(_3347_));
 sg13g2_nand3_1 _8317_ (.B(_3235_),
    .C(_3347_),
    .A(_3278_),
    .Y(_3348_));
 sg13g2_o21ai_1 _8318_ (.B1(_3348_),
    .Y(_3349_),
    .A1(_3345_),
    .A2(_3346_));
 sg13g2_xnor2_1 _8319_ (.Y(_3350_),
    .A(_3326_),
    .B(_3328_));
 sg13g2_xor2_1 _8320_ (.B(_3350_),
    .A(_3349_),
    .X(_3351_));
 sg13g2_xnor2_1 _8321_ (.Y(_3352_),
    .A(_3343_),
    .B(_3342_));
 sg13g2_nand2b_1 _8322_ (.Y(_3353_),
    .B(_3352_),
    .A_N(_3351_));
 sg13g2_nand2b_1 _8323_ (.Y(_3354_),
    .B(_3349_),
    .A_N(_3350_));
 sg13g2_nand2_1 _8324_ (.Y(_3355_),
    .A(_3353_),
    .B(_3354_));
 sg13g2_xor2_1 _8325_ (.B(_3325_),
    .A(_3333_),
    .X(_3356_));
 sg13g2_xor2_1 _8326_ (.B(_3356_),
    .A(_3355_),
    .X(_3357_));
 sg13g2_xor2_1 _8327_ (.B(_3357_),
    .A(_3344_),
    .X(_3358_));
 sg13g2_nor2b_1 _8328_ (.A(_3345_),
    .B_N(_3348_),
    .Y(_3359_));
 sg13g2_xnor2_1 _8329_ (.Y(_3360_),
    .A(_3346_),
    .B(_3359_));
 sg13g2_inv_1 _8330_ (.Y(_3361_),
    .A(net30));
 sg13g2_nor2_1 _8331_ (.A(_3241_),
    .B(_3361_),
    .Y(_3362_));
 sg13g2_xor2_1 _8332_ (.B(_3362_),
    .A(_3347_),
    .X(_3363_));
 sg13g2_nand3_1 _8333_ (.B(_0439_),
    .C(net17),
    .A(_3363_),
    .Y(_3364_));
 sg13g2_nand2_1 _8334_ (.Y(_3365_),
    .A(_3362_),
    .B(_3347_));
 sg13g2_nand2_1 _8335_ (.Y(_3366_),
    .A(_3364_),
    .B(_3365_));
 sg13g2_xnor2_1 _8336_ (.Y(_3367_),
    .A(_3360_),
    .B(_3366_));
 sg13g2_nor3_1 _8337_ (.A(_0440_),
    .B(_3228_),
    .C(_3367_),
    .Y(_3368_));
 sg13g2_o21ai_1 _8338_ (.B1(_3367_),
    .Y(_3369_),
    .A1(_0440_),
    .A2(_3228_));
 sg13g2_nor2b_1 _8339_ (.A(_3368_),
    .B_N(_3369_),
    .Y(_3370_));
 sg13g2_a21o_1 _8340_ (.A2(net17),
    .A1(_0439_),
    .B1(_3363_),
    .X(_3371_));
 sg13g2_nor4_1 _8341_ (.A(_0286_),
    .B(_3287_),
    .C(_3241_),
    .D(_3361_),
    .Y(_3372_));
 sg13g2_nand4_1 _8342_ (.B(_3364_),
    .C(_3371_),
    .A(_3370_),
    .Y(_3373_),
    .D(_3372_));
 sg13g2_a21oi_1 _8343_ (.A1(_3366_),
    .A2(_3360_),
    .Y(_3374_),
    .B1(_3368_));
 sg13g2_nand2_1 _8344_ (.Y(_3375_),
    .A(_3373_),
    .B(_3374_));
 sg13g2_xnor2_1 _8345_ (.Y(_3376_),
    .A(_3352_),
    .B(_3351_));
 sg13g2_nor2_1 _8346_ (.A(_3374_),
    .B(_3373_),
    .Y(_3377_));
 sg13g2_a21oi_1 _8347_ (.A1(_3375_),
    .A2(_3376_),
    .Y(_3378_),
    .B1(_3377_));
 sg13g2_nor2_1 _8348_ (.A(_3358_),
    .B(_3378_),
    .Y(_3379_));
 sg13g2_xnor2_1 _8349_ (.Y(_3380_),
    .A(_3323_),
    .B(_3337_));
 sg13g2_nor2b_1 _8350_ (.A(_3356_),
    .B_N(_3355_),
    .Y(_3381_));
 sg13g2_nor2b_1 _8351_ (.A(_3357_),
    .B_N(_3344_),
    .Y(_3382_));
 sg13g2_nor2_1 _8352_ (.A(_3381_),
    .B(_3382_),
    .Y(_3383_));
 sg13g2_nand2_1 _8353_ (.Y(_3384_),
    .A(_3380_),
    .B(_3383_));
 sg13g2_nor2_1 _8354_ (.A(_3383_),
    .B(_3380_),
    .Y(_3385_));
 sg13g2_a21oi_1 _8355_ (.A1(_3379_),
    .A2(_3384_),
    .Y(_3386_),
    .B1(_3385_));
 sg13g2_nor2_1 _8356_ (.A(_3296_),
    .B(_3315_),
    .Y(_3387_));
 sg13g2_nor2_1 _8357_ (.A(_3248_),
    .B(_3316_),
    .Y(_3388_));
 sg13g2_nor2_1 _8358_ (.A(_3387_),
    .B(_3388_),
    .Y(_3389_));
 sg13g2_nand2_1 _8359_ (.Y(_3390_),
    .A(_3312_),
    .B(_3311_));
 sg13g2_nor2_1 _8360_ (.A(_3311_),
    .B(_3312_),
    .Y(_3391_));
 sg13g2_a21oi_1 _8361_ (.A1(_3390_),
    .A2(_3310_),
    .Y(_3392_),
    .B1(_3391_));
 sg13g2_nor2b_1 _8362_ (.A(_3308_),
    .B_N(_3297_),
    .Y(_3393_));
 sg13g2_nor2b_1 _8363_ (.A(_3314_),
    .B_N(_3309_),
    .Y(_3394_));
 sg13g2_nor2_1 _8364_ (.A(_3393_),
    .B(_3394_),
    .Y(_3395_));
 sg13g2_nor2b_1 _8365_ (.A(_3245_),
    .B_N(_3235_),
    .Y(_3396_));
 sg13g2_nand2_1 _8366_ (.Y(_3397_),
    .A(net15),
    .B(_3275_));
 sg13g2_nor2_1 _8367_ (.A(_3311_),
    .B(_3397_),
    .Y(_3398_));
 sg13g2_a22oi_1 _8368_ (.Y(_3399_),
    .B1(_3258_),
    .B2(_3216_),
    .A2(_3229_),
    .A1(_3275_));
 sg13g2_nor2_1 _8369_ (.A(_3398_),
    .B(_3399_),
    .Y(_3400_));
 sg13g2_xnor2_1 _8370_ (.Y(_3401_),
    .A(_3396_),
    .B(_3400_));
 sg13g2_inv_1 _8371_ (.Y(_3402_),
    .A(_3306_));
 sg13g2_nand2b_1 _8372_ (.Y(_3403_),
    .B(_3402_),
    .A_N(_3299_));
 sg13g2_o21ai_1 _8373_ (.B1(_3403_),
    .Y(_3404_),
    .A1(_3298_),
    .A2(_3307_));
 sg13g2_nor2b_1 _8374_ (.A(_3251_),
    .B_N(_3266_),
    .Y(_3405_));
 sg13g2_o21ai_1 _8375_ (.B1(_0544_),
    .Y(_3406_),
    .A1(_0530_),
    .A2(_3263_));
 sg13g2_inv_1 _8376_ (.Y(_3407_),
    .A(_0530_));
 sg13g2_nand3_1 _8377_ (.B(_3407_),
    .C(\generated._377[7] ),
    .A(_3262_),
    .Y(_3408_));
 sg13g2_nand3_1 _8378_ (.B(_1492_),
    .C(_3408_),
    .A(_3406_),
    .Y(_3409_));
 sg13g2_nand2_1 _8379_ (.Y(_3410_),
    .A(net88),
    .B(_0094_));
 sg13g2_nand2_2 _8380_ (.Y(_3411_),
    .A(_3409_),
    .B(_3410_));
 sg13g2_inv_1 _8381_ (.Y(_3412_),
    .A(_3411_));
 sg13g2_a22oi_1 _8382_ (.Y(_3413_),
    .B1(_3268_),
    .B2(_3412_),
    .A2(_3305_),
    .A1(net30));
 sg13g2_nor2_1 _8383_ (.A(_3361_),
    .B(_3411_),
    .Y(_3414_));
 sg13g2_nand2_1 _8384_ (.Y(_3415_),
    .A(_3414_),
    .B(_3402_));
 sg13g2_nand2b_1 _8385_ (.Y(_3416_),
    .B(_3415_),
    .A_N(_3413_));
 sg13g2_xor2_1 _8386_ (.B(_3416_),
    .A(_3405_),
    .X(_3417_));
 sg13g2_xnor2_1 _8387_ (.Y(_3418_),
    .A(_3404_),
    .B(_3417_));
 sg13g2_xor2_1 _8388_ (.B(_3418_),
    .A(_3401_),
    .X(_3419_));
 sg13g2_xnor2_1 _8389_ (.Y(_3420_),
    .A(_3395_),
    .B(_3419_));
 sg13g2_xnor2_1 _8390_ (.Y(_3421_),
    .A(_3392_),
    .B(_3420_));
 sg13g2_xnor2_1 _8391_ (.Y(_3422_),
    .A(_3389_),
    .B(_3421_));
 sg13g2_nor4_1 _8392_ (.A(_3340_),
    .B(_3341_),
    .C(_3386_),
    .D(_3422_),
    .Y(_3423_));
 sg13g2_nand2b_1 _8393_ (.Y(_3424_),
    .B(_3340_),
    .A_N(_3422_));
 sg13g2_nand2b_1 _8394_ (.Y(_3425_),
    .B(_3424_),
    .A_N(_3423_));
 sg13g2_nor2_1 _8395_ (.A(_3395_),
    .B(_3419_),
    .Y(_3426_));
 sg13g2_nor2_1 _8396_ (.A(_3392_),
    .B(_3420_),
    .Y(_3427_));
 sg13g2_nor2_1 _8397_ (.A(_3426_),
    .B(_3427_),
    .Y(_3428_));
 sg13g2_nand2_1 _8398_ (.Y(_3429_),
    .A(_3244_),
    .B(_3258_));
 sg13g2_a21oi_1 _8399_ (.A1(_3400_),
    .A2(_3396_),
    .Y(_3430_),
    .B1(_3398_));
 sg13g2_xor2_1 _8400_ (.B(_3430_),
    .A(_3429_),
    .X(_3431_));
 sg13g2_a22oi_1 _8401_ (.Y(_3432_),
    .B1(_3266_),
    .B2(_3229_),
    .A2(net17),
    .A1(_3305_));
 sg13g2_nand3_1 _8402_ (.B(_3229_),
    .C(_3305_),
    .A(_3405_),
    .Y(_3433_));
 sg13g2_nor2b_1 _8403_ (.A(_3432_),
    .B_N(_3433_),
    .Y(_3434_));
 sg13g2_xor2_1 _8404_ (.B(_3434_),
    .A(_3397_),
    .X(_3435_));
 sg13g2_nand2_1 _8405_ (.Y(_3436_),
    .A(net17),
    .B(_3266_));
 sg13g2_o21ai_1 _8406_ (.B1(_3415_),
    .Y(_3437_),
    .A1(_3436_),
    .A2(_3413_));
 sg13g2_nor2_1 _8407_ (.A(\generated._377[7] ),
    .B(_3302_),
    .Y(_3438_));
 sg13g2_xnor2_1 _8408_ (.Y(_3439_),
    .A(\generated._376 ),
    .B(_3438_));
 sg13g2_nor2_1 _8409_ (.A(_4488_),
    .B(_3439_),
    .Y(_3440_));
 sg13g2_a21o_1 _8410_ (.A2(_0095_),
    .A1(net88),
    .B1(_3440_),
    .X(_3441_));
 sg13g2_buf_8 _8411_ (.A(_3441_),
    .X(_3442_));
 sg13g2_nor2_1 _8412_ (.A(_3287_),
    .B(_3442_),
    .Y(_3443_));
 sg13g2_xor2_1 _8413_ (.B(_3443_),
    .A(_3414_),
    .X(_3444_));
 sg13g2_xor2_1 _8414_ (.B(_3444_),
    .A(_3437_),
    .X(_3445_));
 sg13g2_xnor2_1 _8415_ (.Y(_3446_),
    .A(_3435_),
    .B(_3445_));
 sg13g2_nor2b_1 _8416_ (.A(_3417_),
    .B_N(_3404_),
    .Y(_3447_));
 sg13g2_nor2b_1 _8417_ (.A(_3401_),
    .B_N(_3418_),
    .Y(_3448_));
 sg13g2_nor2_1 _8418_ (.A(_3447_),
    .B(_3448_),
    .Y(_3449_));
 sg13g2_xor2_1 _8419_ (.B(_3449_),
    .A(_3446_),
    .X(_3450_));
 sg13g2_xor2_1 _8420_ (.B(_3450_),
    .A(_3431_),
    .X(_3451_));
 sg13g2_xnor2_1 _8421_ (.Y(_3452_),
    .A(_3428_),
    .B(_3451_));
 sg13g2_nor2_1 _8422_ (.A(_3389_),
    .B(_3421_),
    .Y(_3453_));
 sg13g2_nand2b_1 _8423_ (.Y(_3454_),
    .B(_3453_),
    .A_N(_3452_));
 sg13g2_nand2b_1 _8424_ (.Y(_3455_),
    .B(_3452_),
    .A_N(_3453_));
 sg13g2_nand3_1 _8425_ (.B(_3454_),
    .C(_3455_),
    .A(_3425_),
    .Y(_3456_));
 sg13g2_nor2_1 _8426_ (.A(_3428_),
    .B(_3451_),
    .Y(_3457_));
 sg13g2_nor2_1 _8427_ (.A(_3429_),
    .B(_3430_),
    .Y(_3458_));
 sg13g2_nor2b_1 _8428_ (.A(_3449_),
    .B_N(_3446_),
    .Y(_3459_));
 sg13g2_nor2b_1 _8429_ (.A(_3450_),
    .B_N(_3431_),
    .Y(_3460_));
 sg13g2_nor2_1 _8430_ (.A(_3459_),
    .B(_3460_),
    .Y(_3461_));
 sg13g2_o21ai_1 _8431_ (.B1(_3433_),
    .Y(_3462_),
    .A1(_3397_),
    .A2(_3432_));
 sg13g2_nor2b_1 _8432_ (.A(_3245_),
    .B_N(_3275_),
    .Y(_3463_));
 sg13g2_nand2_2 _8433_ (.Y(_3464_),
    .A(_3229_),
    .B(_3305_));
 sg13g2_nand2_1 _8434_ (.Y(_3465_),
    .A(net15),
    .B(_3266_));
 sg13g2_xnor2_1 _8435_ (.Y(_3466_),
    .A(_3464_),
    .B(_3465_));
 sg13g2_xor2_1 _8436_ (.B(_3466_),
    .A(_3463_),
    .X(_3467_));
 sg13g2_nor2_1 _8437_ (.A(_3251_),
    .B(_3411_),
    .Y(_3468_));
 sg13g2_inv_2 _8438_ (.Y(_3469_),
    .A(_3442_));
 sg13g2_o21ai_1 _8439_ (.B1(_3469_),
    .Y(_3470_),
    .A1(net30),
    .A2(_3268_));
 sg13g2_inv_1 _8440_ (.Y(_3471_),
    .A(_3443_));
 sg13g2_nor2_1 _8441_ (.A(_3361_),
    .B(_3471_),
    .Y(_3472_));
 sg13g2_nor2_1 _8442_ (.A(_3470_),
    .B(_3472_),
    .Y(_3473_));
 sg13g2_a21oi_1 _8443_ (.A1(_3414_),
    .A2(_3443_),
    .Y(_3474_),
    .B1(_3473_));
 sg13g2_xnor2_1 _8444_ (.Y(_3475_),
    .A(_3468_),
    .B(_3474_));
 sg13g2_xor2_1 _8445_ (.B(_3475_),
    .A(_3467_),
    .X(_3476_));
 sg13g2_nor2b_1 _8446_ (.A(_3435_),
    .B_N(_3445_),
    .Y(_3477_));
 sg13g2_a21o_1 _8447_ (.A2(_3444_),
    .A1(_3437_),
    .B1(_3477_),
    .X(_3478_));
 sg13g2_xor2_1 _8448_ (.B(_3478_),
    .A(_3476_),
    .X(_3479_));
 sg13g2_xor2_1 _8449_ (.B(_3479_),
    .A(_3462_),
    .X(_3480_));
 sg13g2_nor2_1 _8450_ (.A(_3461_),
    .B(_3480_),
    .Y(_3481_));
 sg13g2_nand2_1 _8451_ (.Y(_3482_),
    .A(_3480_),
    .B(_3461_));
 sg13g2_nor2b_1 _8452_ (.A(_3481_),
    .B_N(_3482_),
    .Y(_3483_));
 sg13g2_xnor2_1 _8453_ (.Y(_3484_),
    .A(_3458_),
    .B(_3483_));
 sg13g2_xnor2_1 _8454_ (.Y(_3485_),
    .A(_3457_),
    .B(_3484_));
 sg13g2_xnor2_1 _8455_ (.Y(_3486_),
    .A(_3454_),
    .B(_3485_));
 sg13g2_xnor2_1 _8456_ (.Y(_3487_),
    .A(_3456_),
    .B(_3486_));
 sg13g2_nand3_1 _8457_ (.B(_3204_),
    .C(_3487_),
    .A(_3202_),
    .Y(_3488_));
 sg13g2_nor2b_1 _8458_ (.A(_3476_),
    .B_N(_3478_),
    .Y(_3489_));
 sg13g2_nor2b_1 _8459_ (.A(_3479_),
    .B_N(_3462_),
    .Y(_3490_));
 sg13g2_nor2_1 _8460_ (.A(_3489_),
    .B(_3490_),
    .Y(_3491_));
 sg13g2_nand2_1 _8461_ (.Y(_3492_),
    .A(_3465_),
    .B(_3464_));
 sg13g2_nor2_1 _8462_ (.A(_3464_),
    .B(_3465_),
    .Y(_3493_));
 sg13g2_a21oi_1 _8463_ (.A1(_3492_),
    .A2(_3463_),
    .Y(_3494_),
    .B1(_3493_));
 sg13g2_nor2b_1 _8464_ (.A(_3245_),
    .B_N(_3266_),
    .Y(_3495_));
 sg13g2_nand2_1 _8465_ (.Y(_3496_),
    .A(net15),
    .B(_3412_));
 sg13g2_nor2_1 _8466_ (.A(_3464_),
    .B(_3496_),
    .Y(_3497_));
 sg13g2_nand2_1 _8467_ (.Y(_3498_),
    .A(net15),
    .B(_3305_));
 sg13g2_nand2_1 _8468_ (.Y(_3499_),
    .A(_3229_),
    .B(_3412_));
 sg13g2_nand2_1 _8469_ (.Y(_3500_),
    .A(_3498_),
    .B(_3499_));
 sg13g2_nor2b_1 _8470_ (.A(_3497_),
    .B_N(_3500_),
    .Y(_3501_));
 sg13g2_xnor2_1 _8471_ (.Y(_3502_),
    .A(_3495_),
    .B(_3501_));
 sg13g2_a21oi_1 _8472_ (.A1(_3473_),
    .A2(_3468_),
    .Y(_3503_),
    .B1(_3472_));
 sg13g2_nor2_1 _8473_ (.A(_3251_),
    .B(_3442_),
    .Y(_3504_));
 sg13g2_inv_1 _8474_ (.Y(_3505_),
    .A(_3504_));
 sg13g2_xnor2_1 _8475_ (.Y(_3506_),
    .A(_3505_),
    .B(_3473_));
 sg13g2_xnor2_1 _8476_ (.Y(_3507_),
    .A(_3503_),
    .B(_3506_));
 sg13g2_xnor2_1 _8477_ (.Y(_3508_),
    .A(_3502_),
    .B(_3507_));
 sg13g2_inv_1 _8478_ (.Y(_3509_),
    .A(_3472_));
 sg13g2_nor2_1 _8479_ (.A(_3251_),
    .B(_3509_),
    .Y(_3510_));
 sg13g2_inv_1 _8480_ (.Y(_3511_),
    .A(_3510_));
 sg13g2_nand2b_1 _8481_ (.Y(_3512_),
    .B(_3475_),
    .A_N(_3467_));
 sg13g2_o21ai_1 _8482_ (.B1(_3512_),
    .Y(_3513_),
    .A1(_3411_),
    .A2(_3511_));
 sg13g2_xnor2_1 _8483_ (.Y(_3514_),
    .A(_3508_),
    .B(_3513_));
 sg13g2_xnor2_1 _8484_ (.Y(_3515_),
    .A(_3494_),
    .B(_3514_));
 sg13g2_xor2_1 _8485_ (.B(_3515_),
    .A(_3491_),
    .X(_3516_));
 sg13g2_a21oi_1 _8486_ (.A1(_3482_),
    .A2(_3458_),
    .Y(_3517_),
    .B1(_3481_));
 sg13g2_xnor2_1 _8487_ (.Y(_3518_),
    .A(_3516_),
    .B(_3517_));
 sg13g2_nand2b_1 _8488_ (.Y(_3519_),
    .B(_3457_),
    .A_N(_3484_));
 sg13g2_xor2_1 _8489_ (.B(_3519_),
    .A(_3518_),
    .X(_3520_));
 sg13g2_nand2_1 _8490_ (.Y(_3521_),
    .A(_3456_),
    .B(_3454_));
 sg13g2_nand2_1 _8491_ (.Y(_3522_),
    .A(_3521_),
    .B(_3485_));
 sg13g2_xor2_1 _8492_ (.B(_3522_),
    .A(_3520_),
    .X(_3523_));
 sg13g2_inv_1 _8493_ (.Y(_3524_),
    .A(_3523_));
 sg13g2_nand2_1 _8494_ (.Y(_3525_),
    .A(_3488_),
    .B(_3524_));
 sg13g2_inv_4 _8495_ (.A(_3202_),
    .Y(_3526_));
 sg13g2_nand3_1 _8496_ (.B(_3174_),
    .C(_3526_),
    .A(_3168_),
    .Y(_3527_));
 sg13g2_nand3_1 _8497_ (.B(_3525_),
    .C(_3527_),
    .A(_3203_),
    .Y(_3528_));
 sg13g2_nand2b_1 _8498_ (.Y(_3529_),
    .B(_3523_),
    .A_N(_3488_));
 sg13g2_nand2_1 _8499_ (.Y(_3530_),
    .A(_3528_),
    .B(_3529_));
 sg13g2_inv_1 _8500_ (.Y(_3531_),
    .A(_3516_));
 sg13g2_nor2_1 _8501_ (.A(_3491_),
    .B(_3515_),
    .Y(_3532_));
 sg13g2_nand2_1 _8502_ (.Y(_3533_),
    .A(_3513_),
    .B(_3508_));
 sg13g2_o21ai_1 _8503_ (.B1(_3533_),
    .Y(_3534_),
    .A1(_3494_),
    .A2(_3514_));
 sg13g2_a21oi_1 _8504_ (.A1(_3500_),
    .A2(_3495_),
    .Y(_3535_),
    .B1(_3497_));
 sg13g2_a21oi_2 _8505_ (.B1(_3510_),
    .Y(_3536_),
    .A2(_3505_),
    .A1(_3470_));
 sg13g2_nor2b_1 _8506_ (.A(_3245_),
    .B_N(_3305_),
    .Y(_3537_));
 sg13g2_nand2_1 _8507_ (.Y(_3538_),
    .A(_3469_),
    .B(net15));
 sg13g2_o21ai_1 _8508_ (.B1(_3496_),
    .Y(_3539_),
    .A1(_3228_),
    .A2(_3442_));
 sg13g2_o21ai_1 _8509_ (.B1(_3539_),
    .Y(_3540_),
    .A1(_3499_),
    .A2(_3538_));
 sg13g2_xor2_1 _8510_ (.B(_3540_),
    .A(_3537_),
    .X(_3541_));
 sg13g2_xor2_1 _8511_ (.B(_3541_),
    .A(_3536_),
    .X(_3542_));
 sg13g2_nor2b_1 _8512_ (.A(_3502_),
    .B_N(_3507_),
    .Y(_3543_));
 sg13g2_nor2_1 _8513_ (.A(_3510_),
    .B(_3543_),
    .Y(_3544_));
 sg13g2_xnor2_1 _8514_ (.Y(_3545_),
    .A(_3542_),
    .B(_3544_));
 sg13g2_xnor2_1 _8515_ (.Y(_3546_),
    .A(_3535_),
    .B(_3545_));
 sg13g2_xor2_1 _8516_ (.B(_3546_),
    .A(_3534_),
    .X(_3547_));
 sg13g2_xor2_1 _8517_ (.B(_3547_),
    .A(_3532_),
    .X(_3548_));
 sg13g2_or3_1 _8518_ (.A(_3517_),
    .B(_3531_),
    .C(_3548_),
    .X(_3549_));
 sg13g2_o21ai_1 _8519_ (.B1(_3548_),
    .Y(_3550_),
    .A1(_3531_),
    .A2(_3517_));
 sg13g2_nand2_1 _8520_ (.Y(_3551_),
    .A(_3549_),
    .B(_3550_));
 sg13g2_nand2b_1 _8521_ (.Y(_3552_),
    .B(_3518_),
    .A_N(_3519_));
 sg13g2_o21ai_1 _8522_ (.B1(_3552_),
    .Y(_3553_),
    .A1(_3520_),
    .A2(_3522_));
 sg13g2_xnor2_1 _8523_ (.Y(_3554_),
    .A(_3551_),
    .B(_3553_));
 sg13g2_inv_1 _8524_ (.Y(_3555_),
    .A(_3554_));
 sg13g2_nor2_1 _8525_ (.A(_3163_),
    .B(_3119_),
    .Y(_3556_));
 sg13g2_nand2_1 _8526_ (.Y(_3557_),
    .A(_3183_),
    .B(_3556_));
 sg13g2_nor2b_2 _8527_ (.A(_3133_),
    .B_N(_3134_),
    .Y(_3558_));
 sg13g2_nor2_2 _8528_ (.A(_2768_),
    .B(_2981_),
    .Y(_3559_));
 sg13g2_nand2_1 _8529_ (.Y(_3560_),
    .A(_3076_),
    .B(_3089_));
 sg13g2_o21ai_1 _8530_ (.B1(_3560_),
    .Y(_3561_),
    .A1(_2928_),
    .A2(_2900_));
 sg13g2_nand2_1 _8531_ (.Y(_3562_),
    .A(_3082_),
    .B(_2777_));
 sg13g2_xnor2_1 _8532_ (.Y(_3563_),
    .A(_3076_),
    .B(_3562_));
 sg13g2_a21oi_1 _8533_ (.A1(_3138_),
    .A2(_3140_),
    .Y(_3564_),
    .B1(_3563_));
 sg13g2_nand3_1 _8534_ (.B(_3138_),
    .C(_3140_),
    .A(_3563_),
    .Y(_3565_));
 sg13g2_nor2b_1 _8535_ (.A(_3564_),
    .B_N(_3565_),
    .Y(_3566_));
 sg13g2_xnor2_1 _8536_ (.Y(_3567_),
    .A(_3561_),
    .B(_3566_));
 sg13g2_inv_1 _8537_ (.Y(_3568_),
    .A(_3567_));
 sg13g2_nor2_1 _8538_ (.A(_3084_),
    .B(_3138_),
    .Y(_3569_));
 sg13g2_inv_1 _8539_ (.Y(_3570_),
    .A(_3138_));
 sg13g2_nor2_1 _8540_ (.A(_3140_),
    .B(_3570_),
    .Y(_3571_));
 sg13g2_o21ai_1 _8541_ (.B1(_3139_),
    .Y(_3572_),
    .A1(_3569_),
    .A2(_3571_));
 sg13g2_nor2_1 _8542_ (.A(_3570_),
    .B(_3139_),
    .Y(_3573_));
 sg13g2_a21oi_1 _8543_ (.A1(_3572_),
    .A2(_3136_),
    .Y(_3574_),
    .B1(_3573_));
 sg13g2_inv_1 _8544_ (.Y(_3575_),
    .A(_3574_));
 sg13g2_nand2_1 _8545_ (.Y(_3576_),
    .A(_3568_),
    .B(_3575_));
 sg13g2_nand2_1 _8546_ (.Y(_3577_),
    .A(_3567_),
    .B(_3574_));
 sg13g2_nand2_1 _8547_ (.Y(_3578_),
    .A(_3576_),
    .B(_3577_));
 sg13g2_xor2_1 _8548_ (.B(_3578_),
    .A(_3559_),
    .X(_3579_));
 sg13g2_inv_1 _8549_ (.Y(_3580_),
    .A(_3148_));
 sg13g2_a21oi_1 _8550_ (.A1(_3147_),
    .A2(_3135_),
    .Y(_3581_),
    .B1(_3580_));
 sg13g2_nand2_1 _8551_ (.Y(_3582_),
    .A(_3579_),
    .B(_3581_));
 sg13g2_xnor2_1 _8552_ (.Y(_3583_),
    .A(_3559_),
    .B(_3578_));
 sg13g2_nand2b_1 _8553_ (.Y(_3584_),
    .B(_3583_),
    .A_N(_3581_));
 sg13g2_nand2_1 _8554_ (.Y(_3585_),
    .A(_3582_),
    .B(_3584_));
 sg13g2_xor2_1 _8555_ (.B(_3585_),
    .A(_3558_),
    .X(_3586_));
 sg13g2_inv_1 _8556_ (.Y(_3587_),
    .A(_3151_));
 sg13g2_a21oi_1 _8557_ (.A1(_3155_),
    .A2(_3129_),
    .Y(_3588_),
    .B1(_3587_));
 sg13g2_nand2_1 _8558_ (.Y(_3589_),
    .A(_3586_),
    .B(_3588_));
 sg13g2_xnor2_1 _8559_ (.Y(_3590_),
    .A(_3558_),
    .B(_3585_));
 sg13g2_inv_1 _8560_ (.Y(_3591_),
    .A(_3588_));
 sg13g2_nand2_1 _8561_ (.Y(_3592_),
    .A(_3590_),
    .B(_3591_));
 sg13g2_nand2_1 _8562_ (.Y(_3593_),
    .A(_3589_),
    .B(_3592_));
 sg13g2_inv_1 _8563_ (.Y(_3594_),
    .A(_3593_));
 sg13g2_nor2_1 _8564_ (.A(_3115_),
    .B(_3114_),
    .Y(_3595_));
 sg13g2_inv_1 _8565_ (.Y(_3596_),
    .A(_3158_));
 sg13g2_a21oi_1 _8566_ (.A1(_3595_),
    .A2(_3162_),
    .Y(_3597_),
    .B1(_3596_));
 sg13g2_nand3_1 _8567_ (.B(_3594_),
    .C(_3597_),
    .A(_3557_),
    .Y(_3598_));
 sg13g2_inv_1 _8568_ (.Y(_3599_),
    .A(_3182_));
 sg13g2_nand2_1 _8569_ (.Y(_3600_),
    .A(_3595_),
    .B(_3162_));
 sg13g2_nand2_1 _8570_ (.Y(_3601_),
    .A(_3600_),
    .B(_3158_));
 sg13g2_nor2_1 _8571_ (.A(_3599_),
    .B(_3601_),
    .Y(_3602_));
 sg13g2_nand2_1 _8572_ (.Y(_3603_),
    .A(_3602_),
    .B(_3180_));
 sg13g2_inv_1 _8573_ (.Y(_3604_),
    .A(_3556_));
 sg13g2_nand2b_1 _8574_ (.Y(_3605_),
    .B(_3604_),
    .A_N(_3601_));
 sg13g2_nand3_1 _8575_ (.B(_3605_),
    .C(_3593_),
    .A(_3603_),
    .Y(_3606_));
 sg13g2_nand2_1 _8576_ (.Y(_3607_),
    .A(_3598_),
    .B(_3606_));
 sg13g2_nor2_1 _8577_ (.A(_2695_),
    .B(_2749_),
    .Y(_3608_));
 sg13g2_inv_1 _8578_ (.Y(_3609_),
    .A(_2746_));
 sg13g2_a21oi_1 _8579_ (.A1(_2748_),
    .A2(_2697_),
    .Y(_3610_),
    .B1(_3609_));
 sg13g2_a21oi_1 _8580_ (.A1(_3196_),
    .A2(_3608_),
    .Y(_3611_),
    .B1(_3610_));
 sg13g2_nand3_1 _8581_ (.B(_3193_),
    .C(_3608_),
    .A(_3192_),
    .Y(_3612_));
 sg13g2_nand2_1 _8582_ (.Y(_3613_),
    .A(_3611_),
    .B(_3612_));
 sg13g2_nor2b_1 _8583_ (.A(_2705_),
    .B_N(_2704_),
    .Y(_3614_));
 sg13g2_nor2_1 _8584_ (.A(net14),
    .B(_2243_),
    .Y(_3615_));
 sg13g2_nor2_1 _8585_ (.A(_2315_),
    .B(_2344_),
    .Y(_3616_));
 sg13g2_nor2_1 _8586_ (.A(_2318_),
    .B(_2441_),
    .Y(_3617_));
 sg13g2_a22oi_1 _8587_ (.Y(_3618_),
    .B1(_2718_),
    .B2(_2721_),
    .A2(_3617_),
    .A1(_3616_));
 sg13g2_xnor2_1 _8588_ (.Y(_3619_),
    .A(_3615_),
    .B(_3618_));
 sg13g2_a21oi_1 _8589_ (.A1(_2714_),
    .A2(_2722_),
    .Y(_3620_),
    .B1(_2715_));
 sg13g2_inv_1 _8590_ (.Y(_3621_),
    .A(_2585_));
 sg13g2_a21oi_2 _8591_ (.B1(_2715_),
    .Y(_3622_),
    .A2(_2712_),
    .A1(_3621_));
 sg13g2_inv_1 _8592_ (.Y(_3623_),
    .A(_3622_));
 sg13g2_nor2_1 _8593_ (.A(_2306_),
    .B(_2344_),
    .Y(_3624_));
 sg13g2_inv_4 _8594_ (.A(_2549_),
    .Y(_3625_));
 sg13g2_nand2_1 _8595_ (.Y(_3626_),
    .A(_3625_),
    .B(_2314_));
 sg13g2_xor2_1 _8596_ (.B(_3626_),
    .A(_3617_),
    .X(_3627_));
 sg13g2_xor2_1 _8597_ (.B(_3627_),
    .A(_3624_),
    .X(_3628_));
 sg13g2_xnor2_1 _8598_ (.Y(_3629_),
    .A(_3623_),
    .B(_3628_));
 sg13g2_nor2_1 _8599_ (.A(_3620_),
    .B(_3629_),
    .Y(_3630_));
 sg13g2_nand2_1 _8600_ (.Y(_3631_),
    .A(_3629_),
    .B(_3620_));
 sg13g2_nand2b_1 _8601_ (.Y(_3632_),
    .B(_3631_),
    .A_N(_3630_));
 sg13g2_xnor2_1 _8602_ (.Y(_3633_),
    .A(_3619_),
    .B(_3632_));
 sg13g2_inv_1 _8603_ (.Y(_3634_),
    .A(_3633_));
 sg13g2_inv_1 _8604_ (.Y(_3635_),
    .A(_2726_));
 sg13g2_a21oi_1 _8605_ (.A1(_2728_),
    .A2(_2706_),
    .Y(_3636_),
    .B1(_3635_));
 sg13g2_nand2_1 _8606_ (.Y(_3637_),
    .A(_3634_),
    .B(_3636_));
 sg13g2_nand2b_1 _8607_ (.Y(_3638_),
    .B(_3633_),
    .A_N(_3636_));
 sg13g2_nand2_1 _8608_ (.Y(_3639_),
    .A(_3637_),
    .B(_3638_));
 sg13g2_nand2b_1 _8609_ (.Y(_3640_),
    .B(_3639_),
    .A_N(_3614_));
 sg13g2_nand3_1 _8610_ (.B(_3638_),
    .C(_3614_),
    .A(_3637_),
    .Y(_3641_));
 sg13g2_nand2_1 _8611_ (.Y(_3642_),
    .A(_3640_),
    .B(_3641_));
 sg13g2_inv_2 _8612_ (.Y(_3643_),
    .A(_2736_));
 sg13g2_a21oi_1 _8613_ (.A1(_2735_),
    .A2(_2703_),
    .Y(_3644_),
    .B1(_3643_));
 sg13g2_nand2_1 _8614_ (.Y(_3645_),
    .A(_3642_),
    .B(_3644_));
 sg13g2_inv_1 _8615_ (.Y(_3646_),
    .A(_3644_));
 sg13g2_nand3_1 _8616_ (.B(_3646_),
    .C(_3641_),
    .A(_3640_),
    .Y(_3647_));
 sg13g2_nand2_1 _8617_ (.Y(_3648_),
    .A(_3645_),
    .B(_3647_));
 sg13g2_nand3_1 _8618_ (.B(_2739_),
    .C(_2743_),
    .A(_2738_),
    .Y(_3649_));
 sg13g2_nand2_1 _8619_ (.Y(_3650_),
    .A(_3648_),
    .B(_3649_));
 sg13g2_inv_1 _8620_ (.Y(_3651_),
    .A(_3649_));
 sg13g2_nand3_1 _8621_ (.B(_3647_),
    .C(_3651_),
    .A(_3645_),
    .Y(_3652_));
 sg13g2_nand2_1 _8622_ (.Y(_3653_),
    .A(_3650_),
    .B(_3652_));
 sg13g2_inv_2 _8623_ (.Y(_3654_),
    .A(_3653_));
 sg13g2_nand2_1 _8624_ (.Y(_3655_),
    .A(_3613_),
    .B(_3654_));
 sg13g2_nand3_1 _8625_ (.B(_3612_),
    .C(_3653_),
    .A(_3611_),
    .Y(_3656_));
 sg13g2_nand2_1 _8626_ (.Y(_3657_),
    .A(_3655_),
    .B(_3656_));
 sg13g2_xor2_1 _8627_ (.B(_3657_),
    .A(_3607_),
    .X(_3658_));
 sg13g2_inv_2 _8628_ (.Y(_3659_),
    .A(_3168_));
 sg13g2_a21oi_1 _8629_ (.A1(_3174_),
    .A2(_3526_),
    .Y(_3660_),
    .B1(_3659_));
 sg13g2_xnor2_1 _8630_ (.Y(_3661_),
    .A(_3658_),
    .B(_3660_));
 sg13g2_nor2_1 _8631_ (.A(_3555_),
    .B(_3661_),
    .Y(_3662_));
 sg13g2_nand2_1 _8632_ (.Y(_3663_),
    .A(_3661_),
    .B(_3555_));
 sg13g2_nand2b_1 _8633_ (.Y(_3664_),
    .B(_3663_),
    .A_N(_3662_));
 sg13g2_xnor2_1 _8634_ (.Y(\generated._825[2] ),
    .A(_3530_),
    .B(_3664_));
 sg13g2_a21oi_1 _8635_ (.A1(_3663_),
    .A2(_3530_),
    .Y(_3665_),
    .B1(_3662_));
 sg13g2_nor2_1 _8636_ (.A(_3202_),
    .B(_3175_),
    .Y(_3666_));
 sg13g2_nand2b_1 _8637_ (.Y(_3667_),
    .B(_3666_),
    .A_N(_3658_));
 sg13g2_nand2_1 _8638_ (.Y(_3668_),
    .A(_2674_),
    .B(_2690_));
 sg13g2_nor2_1 _8639_ (.A(_3668_),
    .B(_3191_),
    .Y(_3669_));
 sg13g2_xnor2_1 _8640_ (.Y(_3670_),
    .A(_2672_),
    .B(_2656_));
 sg13g2_nor2b_1 _8641_ (.A(_3670_),
    .B_N(_2682_),
    .Y(_3671_));
 sg13g2_nand2_1 _8642_ (.Y(_3672_),
    .A(_3669_),
    .B(_3671_));
 sg13g2_inv_1 _8643_ (.Y(_3673_),
    .A(_2684_));
 sg13g2_a21oi_1 _8644_ (.A1(_2690_),
    .A2(_2518_),
    .Y(_3674_),
    .B1(_3673_));
 sg13g2_inv_1 _8645_ (.Y(_3675_),
    .A(_3674_));
 sg13g2_nand2_1 _8646_ (.Y(_3676_),
    .A(_3672_),
    .B(_3675_));
 sg13g2_nand2_1 _8647_ (.Y(_3677_),
    .A(_3654_),
    .B(_2750_));
 sg13g2_nor2_1 _8648_ (.A(_2695_),
    .B(_3188_),
    .Y(_3678_));
 sg13g2_nor2b_1 _8649_ (.A(_3677_),
    .B_N(_3678_),
    .Y(_3679_));
 sg13g2_nand2_1 _8650_ (.Y(_3680_),
    .A(_3676_),
    .B(_3679_));
 sg13g2_inv_1 _8651_ (.Y(_3681_),
    .A(_3650_));
 sg13g2_a21oi_1 _8652_ (.A1(_3652_),
    .A2(_2748_),
    .Y(_3682_),
    .B1(_3681_));
 sg13g2_nor2_1 _8653_ (.A(_2699_),
    .B(_3677_),
    .Y(_3683_));
 sg13g2_nor2_1 _8654_ (.A(_3682_),
    .B(_3683_),
    .Y(_3684_));
 sg13g2_nand2_1 _8655_ (.Y(_3685_),
    .A(_3680_),
    .B(_3684_));
 sg13g2_inv_2 _8656_ (.Y(_3686_),
    .A(_3647_));
 sg13g2_inv_1 _8657_ (.Y(_3687_),
    .A(_3638_));
 sg13g2_a21oi_1 _8658_ (.A1(_3637_),
    .A2(_3614_),
    .Y(_3688_),
    .B1(_3687_));
 sg13g2_nor2_1 _8659_ (.A(net14),
    .B(_2344_),
    .Y(_3689_));
 sg13g2_nand3_1 _8660_ (.B(_2292_),
    .C(_2314_),
    .A(_3625_),
    .Y(_3690_));
 sg13g2_buf_1 _8661_ (.A(_3690_),
    .X(_3691_));
 sg13g2_inv_1 _8662_ (.Y(_3692_),
    .A(_3691_));
 sg13g2_nor2b_1 _8663_ (.A(_3627_),
    .B_N(_3624_),
    .Y(_3693_));
 sg13g2_a21oi_1 _8664_ (.A1(_2719_),
    .A2(_3692_),
    .Y(_3694_),
    .B1(_3693_));
 sg13g2_xnor2_1 _8665_ (.Y(_3695_),
    .A(_3689_),
    .B(_3694_));
 sg13g2_nor2_1 _8666_ (.A(_2306_),
    .B(_2441_),
    .Y(_3696_));
 sg13g2_a21oi_1 _8667_ (.A1(_2315_),
    .A2(_2318_),
    .Y(_3697_),
    .B1(_2549_));
 sg13g2_nand2_1 _8668_ (.Y(_3698_),
    .A(_3691_),
    .B(_3697_));
 sg13g2_xor2_1 _8669_ (.B(_3698_),
    .A(_3696_),
    .X(_3699_));
 sg13g2_xnor2_1 _8670_ (.Y(_3700_),
    .A(_3622_),
    .B(_3699_));
 sg13g2_inv_1 _8671_ (.Y(_3701_),
    .A(_3628_));
 sg13g2_a21oi_1 _8672_ (.A1(_3701_),
    .A2(_3622_),
    .Y(_3702_),
    .B1(_2715_));
 sg13g2_xnor2_1 _8673_ (.Y(_3703_),
    .A(_3700_),
    .B(_3702_));
 sg13g2_xor2_1 _8674_ (.B(_3703_),
    .A(_3695_),
    .X(_3704_));
 sg13g2_a21oi_1 _8675_ (.A1(_3631_),
    .A2(_3619_),
    .Y(_3705_),
    .B1(_3630_));
 sg13g2_inv_1 _8676_ (.Y(_3706_),
    .A(_3705_));
 sg13g2_nand2_1 _8677_ (.Y(_3707_),
    .A(_3704_),
    .B(_3706_));
 sg13g2_xnor2_1 _8678_ (.Y(_3708_),
    .A(_3695_),
    .B(_3703_));
 sg13g2_nand2_1 _8679_ (.Y(_3709_),
    .A(_3708_),
    .B(_3705_));
 sg13g2_nand2_1 _8680_ (.Y(_3710_),
    .A(_3707_),
    .B(_3709_));
 sg13g2_nor2b_1 _8681_ (.A(_3618_),
    .B_N(_3615_),
    .Y(_3711_));
 sg13g2_nand2_1 _8682_ (.Y(_3712_),
    .A(_3710_),
    .B(_3711_));
 sg13g2_inv_1 _8683_ (.Y(_3713_),
    .A(_3711_));
 sg13g2_nand3_1 _8684_ (.B(_3709_),
    .C(_3713_),
    .A(_3707_),
    .Y(_3714_));
 sg13g2_nand2_1 _8685_ (.Y(_3715_),
    .A(_3712_),
    .B(_3714_));
 sg13g2_xnor2_1 _8686_ (.Y(_3716_),
    .A(_3688_),
    .B(_3715_));
 sg13g2_nor2_1 _8687_ (.A(_3686_),
    .B(_3716_),
    .Y(_3717_));
 sg13g2_nand2_1 _8688_ (.Y(_3718_),
    .A(_3716_),
    .B(_3686_));
 sg13g2_nor2b_1 _8689_ (.A(_3717_),
    .B_N(_3718_),
    .Y(_3719_));
 sg13g2_nand2_1 _8690_ (.Y(_3720_),
    .A(_3685_),
    .B(_3719_));
 sg13g2_nand2b_1 _8691_ (.Y(_3721_),
    .B(_3718_),
    .A_N(_3717_));
 sg13g2_nand3_1 _8692_ (.B(_3684_),
    .C(_3721_),
    .A(_3680_),
    .Y(_3722_));
 sg13g2_nand2_1 _8693_ (.Y(_3723_),
    .A(_3720_),
    .B(_3722_));
 sg13g2_nor2_1 _8694_ (.A(_3593_),
    .B(_3163_),
    .Y(_3724_));
 sg13g2_nand2_1 _8695_ (.Y(_3725_),
    .A(_3596_),
    .B(_3589_));
 sg13g2_nand2_1 _8696_ (.Y(_3726_),
    .A(_3725_),
    .B(_3592_));
 sg13g2_a21oi_1 _8697_ (.A1(_3724_),
    .A2(_3124_),
    .Y(_3727_),
    .B1(_3726_));
 sg13g2_nand3_1 _8698_ (.B(_3120_),
    .C(_3724_),
    .A(_3032_),
    .Y(_3728_));
 sg13g2_nand2_1 _8699_ (.Y(_3729_),
    .A(_3727_),
    .B(_3728_));
 sg13g2_inv_1 _8700_ (.Y(_3730_),
    .A(_3576_));
 sg13g2_a21oi_1 _8701_ (.A1(_3577_),
    .A2(_3559_),
    .Y(_3731_),
    .B1(_3730_));
 sg13g2_nor2_1 _8702_ (.A(_2768_),
    .B(_3045_),
    .Y(_3732_));
 sg13g2_inv_1 _8703_ (.Y(_3733_),
    .A(_3732_));
 sg13g2_inv_1 _8704_ (.Y(_3734_),
    .A(_2981_));
 sg13g2_nor3_1 _8705_ (.A(_2782_),
    .B(_2839_),
    .C(_3045_),
    .Y(_3735_));
 sg13g2_a21oi_1 _8706_ (.A1(_3734_),
    .A2(_2862_),
    .Y(_3736_),
    .B1(_3735_));
 sg13g2_nor2_1 _8707_ (.A(_3140_),
    .B(_3563_),
    .Y(_3737_));
 sg13g2_xor2_1 _8708_ (.B(_3737_),
    .A(_3736_),
    .X(_3738_));
 sg13g2_nor3_1 _8709_ (.A(_3084_),
    .B(_3138_),
    .C(_3563_),
    .Y(_3739_));
 sg13g2_a21o_1 _8710_ (.A2(_3561_),
    .A1(_3566_),
    .B1(_3739_),
    .X(_3740_));
 sg13g2_xnor2_1 _8711_ (.Y(_3741_),
    .A(_3738_),
    .B(_3740_));
 sg13g2_xnor2_1 _8712_ (.Y(_3742_),
    .A(_3733_),
    .B(_3741_));
 sg13g2_xor2_1 _8713_ (.B(_3742_),
    .A(_3731_),
    .X(_3743_));
 sg13g2_inv_1 _8714_ (.Y(_3744_),
    .A(_3584_));
 sg13g2_a21oi_1 _8715_ (.A1(_3582_),
    .A2(_3558_),
    .Y(_3745_),
    .B1(_3744_));
 sg13g2_xor2_1 _8716_ (.B(_3745_),
    .A(_3743_),
    .X(_3746_));
 sg13g2_nand2_1 _8717_ (.Y(_3747_),
    .A(_3729_),
    .B(_3746_));
 sg13g2_inv_1 _8718_ (.Y(_3748_),
    .A(_3746_));
 sg13g2_nand3_1 _8719_ (.B(_3728_),
    .C(_3748_),
    .A(_3727_),
    .Y(_3749_));
 sg13g2_nand2_1 _8720_ (.Y(_3750_),
    .A(_3747_),
    .B(_3749_));
 sg13g2_inv_1 _8721_ (.Y(_3751_),
    .A(_3750_));
 sg13g2_nand2_1 _8722_ (.Y(_3752_),
    .A(_3723_),
    .B(_3751_));
 sg13g2_nand3_1 _8723_ (.B(_3722_),
    .C(_3750_),
    .A(_3720_),
    .Y(_3753_));
 sg13g2_nand2_1 _8724_ (.Y(_3754_),
    .A(_3752_),
    .B(_3753_));
 sg13g2_nand2b_1 _8725_ (.Y(_3755_),
    .B(_3657_),
    .A_N(_3607_));
 sg13g2_nor2b_1 _8726_ (.A(_3657_),
    .B_N(_3607_),
    .Y(_3756_));
 sg13g2_a21oi_1 _8727_ (.A1(_3755_),
    .A2(_3659_),
    .Y(_3757_),
    .B1(_3756_));
 sg13g2_nand3_1 _8728_ (.B(_3754_),
    .C(_3757_),
    .A(_3667_),
    .Y(_3758_));
 sg13g2_nor2_1 _8729_ (.A(_3659_),
    .B(_3756_),
    .Y(_3759_));
 sg13g2_nand2_1 _8730_ (.Y(_3760_),
    .A(_3527_),
    .B(_3759_));
 sg13g2_inv_1 _8731_ (.Y(_3761_),
    .A(_3754_));
 sg13g2_nand3_1 _8732_ (.B(_3761_),
    .C(_3755_),
    .A(_3760_),
    .Y(_3762_));
 sg13g2_nand2b_1 _8733_ (.Y(_3763_),
    .B(_3532_),
    .A_N(_3547_));
 sg13g2_nor2b_1 _8734_ (.A(_3546_),
    .B_N(_3534_),
    .Y(_3764_));
 sg13g2_nor2_1 _8735_ (.A(_3228_),
    .B(_3538_),
    .Y(_3765_));
 sg13g2_a22oi_1 _8736_ (.Y(_3766_),
    .B1(_3412_),
    .B2(_3765_),
    .A2(_3537_),
    .A1(_3539_));
 sg13g2_nor2_1 _8737_ (.A(_3245_),
    .B(_3411_),
    .Y(_3767_));
 sg13g2_a21oi_1 _8738_ (.A1(_3215_),
    .A2(_3228_),
    .Y(_3768_),
    .B1(_3442_));
 sg13g2_nor2b_1 _8739_ (.A(_3765_),
    .B_N(_3768_),
    .Y(_3769_));
 sg13g2_xnor2_1 _8740_ (.Y(_3770_),
    .A(_3767_),
    .B(_3769_));
 sg13g2_xnor2_1 _8741_ (.Y(_3771_),
    .A(_3536_),
    .B(_3770_));
 sg13g2_nand2b_1 _8742_ (.Y(_3772_),
    .B(_3536_),
    .A_N(_3541_));
 sg13g2_nand2_1 _8743_ (.Y(_3773_),
    .A(_3772_),
    .B(_3511_));
 sg13g2_xnor2_1 _8744_ (.Y(_3774_),
    .A(_3771_),
    .B(_3773_));
 sg13g2_xnor2_1 _8745_ (.Y(_3775_),
    .A(_3766_),
    .B(_3774_));
 sg13g2_nor2_1 _8746_ (.A(_3542_),
    .B(_3544_),
    .Y(_3776_));
 sg13g2_nor2_1 _8747_ (.A(_3535_),
    .B(_3545_),
    .Y(_3777_));
 sg13g2_nor2_1 _8748_ (.A(_3776_),
    .B(_3777_),
    .Y(_3778_));
 sg13g2_xnor2_1 _8749_ (.Y(_3779_),
    .A(_3775_),
    .B(_3778_));
 sg13g2_xor2_1 _8750_ (.B(_3779_),
    .A(_3764_),
    .X(_3780_));
 sg13g2_nor2_1 _8751_ (.A(_3763_),
    .B(_3780_),
    .Y(_3781_));
 sg13g2_nand2_1 _8752_ (.Y(_3782_),
    .A(_3780_),
    .B(_3763_));
 sg13g2_nand2b_1 _8753_ (.Y(_3783_),
    .B(_3782_),
    .A_N(_3781_));
 sg13g2_nand2_1 _8754_ (.Y(_3784_),
    .A(_3553_),
    .B(_3550_));
 sg13g2_nand2_1 _8755_ (.Y(_3785_),
    .A(_3784_),
    .B(_3549_));
 sg13g2_xnor2_1 _8756_ (.Y(_3786_),
    .A(_3783_),
    .B(_3785_));
 sg13g2_a21oi_1 _8757_ (.A1(_3758_),
    .A2(_3762_),
    .Y(_3787_),
    .B1(_3786_));
 sg13g2_nand3_1 _8758_ (.B(_3762_),
    .C(_3786_),
    .A(_3758_),
    .Y(_3788_));
 sg13g2_inv_1 _8759_ (.Y(_3789_),
    .A(_3788_));
 sg13g2_nor2_1 _8760_ (.A(_3787_),
    .B(_3789_),
    .Y(_3790_));
 sg13g2_xnor2_1 _8761_ (.Y(\generated._825[3] ),
    .A(_3665_),
    .B(_3790_));
 sg13g2_a21oi_1 _8762_ (.A1(_3785_),
    .A2(_3782_),
    .Y(_3791_),
    .B1(_3781_));
 sg13g2_or2_1 _8763_ (.X(_3792_),
    .B(_3778_),
    .A(_3775_));
 sg13g2_nand2b_1 _8764_ (.Y(_3793_),
    .B(_3764_),
    .A_N(_3779_));
 sg13g2_a21oi_1 _8765_ (.A1(_3767_),
    .A2(_3768_),
    .Y(_3794_),
    .B1(_3765_));
 sg13g2_nand2_1 _8766_ (.Y(_3795_),
    .A(_3469_),
    .B(_3244_));
 sg13g2_xnor2_1 _8767_ (.Y(_3796_),
    .A(_3795_),
    .B(_3769_));
 sg13g2_xnor2_1 _8768_ (.Y(_3797_),
    .A(_3536_),
    .B(_3796_));
 sg13g2_nand2b_1 _8769_ (.Y(_3798_),
    .B(_3536_),
    .A_N(_3770_));
 sg13g2_nand2_1 _8770_ (.Y(_3799_),
    .A(_3798_),
    .B(_3511_));
 sg13g2_xnor2_1 _8771_ (.Y(_3800_),
    .A(_3797_),
    .B(_3799_));
 sg13g2_xnor2_1 _8772_ (.Y(_3801_),
    .A(_3794_),
    .B(_3800_));
 sg13g2_nand2_1 _8773_ (.Y(_3802_),
    .A(_3773_),
    .B(_3771_));
 sg13g2_o21ai_1 _8774_ (.B1(_3802_),
    .Y(_3803_),
    .A1(_3766_),
    .A2(_3774_));
 sg13g2_xnor2_1 _8775_ (.Y(_3804_),
    .A(_3801_),
    .B(_3803_));
 sg13g2_nand4_1 _8776_ (.B(_3792_),
    .C(_3793_),
    .A(_3791_),
    .Y(_3805_),
    .D(_3804_));
 sg13g2_nor2_1 _8777_ (.A(_3746_),
    .B(_3593_),
    .Y(_3806_));
 sg13g2_nand3_1 _8778_ (.B(_3556_),
    .C(_3806_),
    .A(_3183_),
    .Y(_3807_));
 sg13g2_nor2_1 _8779_ (.A(_3731_),
    .B(_3742_),
    .Y(_3808_));
 sg13g2_a21oi_1 _8780_ (.A1(_3082_),
    .A2(_2862_),
    .Y(_3809_),
    .B1(_3735_));
 sg13g2_nor2b_1 _8781_ (.A(_3737_),
    .B_N(_3736_),
    .Y(_3810_));
 sg13g2_xnor2_1 _8782_ (.Y(_3811_),
    .A(_3809_),
    .B(_3810_));
 sg13g2_xnor2_1 _8783_ (.Y(_3812_),
    .A(_3733_),
    .B(_3811_));
 sg13g2_nor2_1 _8784_ (.A(_3733_),
    .B(_3741_),
    .Y(_3813_));
 sg13g2_a21oi_1 _8785_ (.A1(_3740_),
    .A2(_3738_),
    .Y(_3814_),
    .B1(_3813_));
 sg13g2_xnor2_1 _8786_ (.Y(_3815_),
    .A(_3812_),
    .B(_3814_));
 sg13g2_nor2_1 _8787_ (.A(_3808_),
    .B(_3815_),
    .Y(_3816_));
 sg13g2_nand2b_1 _8788_ (.Y(_3817_),
    .B(_3743_),
    .A_N(_3745_));
 sg13g2_o21ai_1 _8789_ (.B1(_3817_),
    .Y(_3818_),
    .A1(_3592_),
    .A2(_3746_));
 sg13g2_a21oi_1 _8790_ (.A1(_3601_),
    .A2(_3806_),
    .Y(_3819_),
    .B1(_3818_));
 sg13g2_nand3_1 _8791_ (.B(_3816_),
    .C(_3819_),
    .A(_3807_),
    .Y(_3820_));
 sg13g2_nor2_1 _8792_ (.A(_3653_),
    .B(_3721_),
    .Y(_3821_));
 sg13g2_inv_1 _8793_ (.Y(_3822_),
    .A(_3821_));
 sg13g2_nor2b_1 _8794_ (.A(_3822_),
    .B_N(_3608_),
    .Y(_3823_));
 sg13g2_nand2_1 _8795_ (.Y(_3824_),
    .A(_3198_),
    .B(_3823_));
 sg13g2_a21oi_1 _8796_ (.A1(_3652_),
    .A2(_3718_),
    .Y(_3825_),
    .B1(_3717_));
 sg13g2_a21oi_1 _8797_ (.A1(_3821_),
    .A2(_3610_),
    .Y(_3826_),
    .B1(_3825_));
 sg13g2_nand2_1 _8798_ (.Y(_3827_),
    .A(_3824_),
    .B(_3826_));
 sg13g2_a21oi_1 _8799_ (.A1(_3712_),
    .A2(_3714_),
    .Y(_3828_),
    .B1(_3688_));
 sg13g2_inv_1 _8800_ (.Y(_3829_),
    .A(_3707_));
 sg13g2_a21oi_1 _8801_ (.A1(_3709_),
    .A2(_3711_),
    .Y(_3830_),
    .B1(_3829_));
 sg13g2_inv_1 _8802_ (.Y(_3831_),
    .A(_3689_));
 sg13g2_nor2_1 _8803_ (.A(_3831_),
    .B(_3694_),
    .Y(_3832_));
 sg13g2_nor2_1 _8804_ (.A(net14),
    .B(_2441_),
    .Y(_3833_));
 sg13g2_a21oi_1 _8805_ (.A1(_3697_),
    .A2(_3696_),
    .Y(_3834_),
    .B1(_3692_));
 sg13g2_xnor2_1 _8806_ (.Y(_3835_),
    .A(_3833_),
    .B(_3834_));
 sg13g2_nand2_1 _8807_ (.Y(_3836_),
    .A(_3625_),
    .B(_2522_));
 sg13g2_xnor2_1 _8808_ (.Y(_3837_),
    .A(_3836_),
    .B(_3698_));
 sg13g2_xnor2_1 _8809_ (.Y(_3838_),
    .A(_3622_),
    .B(_3837_));
 sg13g2_inv_1 _8810_ (.Y(_3839_),
    .A(_3699_));
 sg13g2_a21oi_1 _8811_ (.A1(_3839_),
    .A2(_3622_),
    .Y(_3840_),
    .B1(_2715_));
 sg13g2_xnor2_1 _8812_ (.Y(_3841_),
    .A(_3838_),
    .B(_3840_));
 sg13g2_xor2_1 _8813_ (.B(_3841_),
    .A(_3835_),
    .X(_3842_));
 sg13g2_inv_1 _8814_ (.Y(_3843_),
    .A(_3842_));
 sg13g2_inv_1 _8815_ (.Y(_3844_),
    .A(_3700_));
 sg13g2_nand2_1 _8816_ (.Y(_3845_),
    .A(_3702_),
    .B(_3844_));
 sg13g2_nor2_1 _8817_ (.A(_3844_),
    .B(_3702_),
    .Y(_3846_));
 sg13g2_a21oi_1 _8818_ (.A1(_3845_),
    .A2(_3695_),
    .Y(_3847_),
    .B1(_3846_));
 sg13g2_nand2_1 _8819_ (.Y(_3848_),
    .A(_3843_),
    .B(_3847_));
 sg13g2_nand2b_1 _8820_ (.Y(_3849_),
    .B(_3842_),
    .A_N(_3847_));
 sg13g2_nand2_1 _8821_ (.Y(_3850_),
    .A(_3848_),
    .B(_3849_));
 sg13g2_nand2b_1 _8822_ (.Y(_3851_),
    .B(_3850_),
    .A_N(_3832_));
 sg13g2_nand3_1 _8823_ (.B(_3832_),
    .C(_3849_),
    .A(_3848_),
    .Y(_3852_));
 sg13g2_nand2_1 _8824_ (.Y(_3853_),
    .A(_3851_),
    .B(_3852_));
 sg13g2_xnor2_1 _8825_ (.Y(_3854_),
    .A(_3830_),
    .B(_3853_));
 sg13g2_xnor2_1 _8826_ (.Y(_3855_),
    .A(_3828_),
    .B(_3854_));
 sg13g2_nand2_1 _8827_ (.Y(_3856_),
    .A(_3827_),
    .B(_3855_));
 sg13g2_inv_1 _8828_ (.Y(_3857_),
    .A(_3855_));
 sg13g2_nand3_1 _8829_ (.B(_3857_),
    .C(_3826_),
    .A(_3824_),
    .Y(_3858_));
 sg13g2_nand2_1 _8830_ (.Y(_3859_),
    .A(_3856_),
    .B(_3858_));
 sg13g2_nand2b_1 _8831_ (.Y(_3860_),
    .B(_3859_),
    .A_N(_3820_));
 sg13g2_nand3_1 _8832_ (.B(_3858_),
    .C(_3820_),
    .A(_3856_),
    .Y(_3861_));
 sg13g2_buf_8 _8833_ (.A(_3861_),
    .X(_3862_));
 sg13g2_nand2_1 _8834_ (.Y(_3863_),
    .A(_3860_),
    .B(_3862_));
 sg13g2_nor2_1 _8835_ (.A(_3658_),
    .B(_3754_),
    .Y(_3864_));
 sg13g2_inv_1 _8836_ (.Y(_3865_),
    .A(_3660_));
 sg13g2_nand2_1 _8837_ (.Y(_3866_),
    .A(_3864_),
    .B(_3865_));
 sg13g2_inv_1 _8838_ (.Y(_3867_),
    .A(_3753_));
 sg13g2_a21oi_1 _8839_ (.A1(_3752_),
    .A2(_3756_),
    .Y(_3868_),
    .B1(_3867_));
 sg13g2_nand2_1 _8840_ (.Y(_3869_),
    .A(_3866_),
    .B(_3868_));
 sg13g2_nand2b_1 _8841_ (.Y(_3870_),
    .B(_3869_),
    .A_N(_3863_));
 sg13g2_nand3_1 _8842_ (.B(_3868_),
    .C(_3863_),
    .A(_3866_),
    .Y(_3871_));
 sg13g2_nand2_1 _8843_ (.Y(_3872_),
    .A(_3870_),
    .B(_3871_));
 sg13g2_xnor2_1 _8844_ (.Y(_3873_),
    .A(_3805_),
    .B(_3872_));
 sg13g2_o21ai_1 _8845_ (.B1(_3788_),
    .Y(_3874_),
    .A1(_3787_),
    .A2(_3665_));
 sg13g2_xor2_1 _8846_ (.B(_3874_),
    .A(_3873_),
    .X(\generated._825[4] ));
 sg13g2_nor2_1 _8847_ (.A(_3754_),
    .B(_3863_),
    .Y(_3875_));
 sg13g2_nand3_1 _8848_ (.B(_3755_),
    .C(_3760_),
    .A(_3875_),
    .Y(_3876_));
 sg13g2_inv_1 _8849_ (.Y(_3877_),
    .A(_3862_));
 sg13g2_o21ai_1 _8850_ (.B1(_3860_),
    .Y(_3878_),
    .A1(_3867_),
    .A2(_3877_));
 sg13g2_nand2_1 _8851_ (.Y(_3879_),
    .A(_3876_),
    .B(_3878_));
 sg13g2_nand2_1 _8852_ (.Y(_3880_),
    .A(_3737_),
    .B(_3809_));
 sg13g2_nor2_1 _8853_ (.A(_3732_),
    .B(_3880_),
    .Y(_3881_));
 sg13g2_inv_1 _8854_ (.Y(_3882_),
    .A(_3830_));
 sg13g2_nand3_1 _8855_ (.B(_3851_),
    .C(_3852_),
    .A(_3882_),
    .Y(_3883_));
 sg13g2_nand2b_1 _8856_ (.Y(_3884_),
    .B(_3833_),
    .A_N(_3834_));
 sg13g2_nand2_1 _8857_ (.Y(_3885_),
    .A(_3625_),
    .B(_2521_));
 sg13g2_o21ai_1 _8858_ (.B1(_3691_),
    .Y(_3886_),
    .A1(_3836_),
    .A2(_3698_));
 sg13g2_xnor2_1 _8859_ (.Y(_3887_),
    .A(_3885_),
    .B(_3886_));
 sg13g2_nand3_1 _8860_ (.B(_2716_),
    .C(_3623_),
    .A(_3837_),
    .Y(_3888_));
 sg13g2_o21ai_1 _8861_ (.B1(_3888_),
    .Y(_3889_),
    .A1(_2716_),
    .A2(_3837_));
 sg13g2_xor2_1 _8862_ (.B(_3889_),
    .A(_3887_),
    .X(_3890_));
 sg13g2_nor2b_1 _8863_ (.A(_3840_),
    .B_N(_3838_),
    .Y(_3891_));
 sg13g2_a21oi_1 _8864_ (.A1(_3841_),
    .A2(_3835_),
    .Y(_3892_),
    .B1(_3891_));
 sg13g2_xnor2_1 _8865_ (.Y(_3893_),
    .A(_3890_),
    .B(_3892_));
 sg13g2_xnor2_1 _8866_ (.Y(_3894_),
    .A(_3884_),
    .B(_3893_));
 sg13g2_nand4_1 _8867_ (.B(_3849_),
    .C(_3852_),
    .A(_3883_),
    .Y(_3895_),
    .D(_3894_));
 sg13g2_nand2_1 _8868_ (.Y(_3896_),
    .A(_3674_),
    .B(_3678_));
 sg13g2_nand2_1 _8869_ (.Y(_3897_),
    .A(_3896_),
    .B(_2699_));
 sg13g2_nand2_1 _8870_ (.Y(_3898_),
    .A(_3719_),
    .B(_3855_));
 sg13g2_nor2_1 _8871_ (.A(_3898_),
    .B(_3677_),
    .Y(_3899_));
 sg13g2_nand2_1 _8872_ (.Y(_3900_),
    .A(_3897_),
    .B(_3899_));
 sg13g2_nor2_1 _8873_ (.A(_3857_),
    .B(_3721_),
    .Y(_3901_));
 sg13g2_nand2b_1 _8874_ (.Y(_3902_),
    .B(_3855_),
    .A_N(_3718_));
 sg13g2_nand2b_1 _8875_ (.Y(_3903_),
    .B(_3828_),
    .A_N(_3854_));
 sg13g2_nand2_1 _8876_ (.Y(_3904_),
    .A(_3902_),
    .B(_3903_));
 sg13g2_a21oi_1 _8877_ (.A1(_3901_),
    .A2(_3682_),
    .Y(_3905_),
    .B1(_3904_));
 sg13g2_nand3b_1 _8878_ (.B(_3900_),
    .C(_3905_),
    .Y(_3906_),
    .A_N(_3895_));
 sg13g2_xnor2_1 _8879_ (.Y(_3907_),
    .A(_3881_),
    .B(_3906_));
 sg13g2_nand2_1 _8880_ (.Y(_3908_),
    .A(_3879_),
    .B(_3907_));
 sg13g2_inv_2 _8881_ (.Y(_3909_),
    .A(_3907_));
 sg13g2_nand3_1 _8882_ (.B(_3878_),
    .C(_3909_),
    .A(_3876_),
    .Y(_3910_));
 sg13g2_nand2_1 _8883_ (.Y(_3911_),
    .A(_3908_),
    .B(_3910_));
 sg13g2_nand2_1 _8884_ (.Y(_3912_),
    .A(_3911_),
    .B(_3442_));
 sg13g2_nand3_1 _8885_ (.B(_3910_),
    .C(_3469_),
    .A(_3908_),
    .Y(_3913_));
 sg13g2_buf_1 _8886_ (.A(_3913_),
    .X(_3914_));
 sg13g2_nand2_1 _8887_ (.Y(_3915_),
    .A(_3912_),
    .B(_3914_));
 sg13g2_nand2_1 _8888_ (.Y(_3916_),
    .A(_3874_),
    .B(_3873_));
 sg13g2_nand3_1 _8889_ (.B(_3871_),
    .C(_3805_),
    .A(_3870_),
    .Y(_3917_));
 sg13g2_nand2_1 _8890_ (.Y(_3918_),
    .A(_3916_),
    .B(_3917_));
 sg13g2_xnor2_1 _8891_ (.Y(\generated._825[5] ),
    .A(_3915_),
    .B(_3918_));
 sg13g2_nand4_1 _8892_ (.B(_3873_),
    .C(_3912_),
    .A(_3874_),
    .Y(_3919_),
    .D(_3914_));
 sg13g2_inv_1 _8893_ (.Y(_3920_),
    .A(_3914_));
 sg13g2_nor2_1 _8894_ (.A(_3917_),
    .B(_3915_),
    .Y(_3921_));
 sg13g2_nor2_1 _8895_ (.A(_3920_),
    .B(_3921_),
    .Y(_3922_));
 sg13g2_nand2_1 _8896_ (.Y(_3923_),
    .A(_3919_),
    .B(_3922_));
 sg13g2_inv_1 _8897_ (.Y(_3924_),
    .A(_3881_));
 sg13g2_nand2_1 _8898_ (.Y(_3925_),
    .A(_3906_),
    .B(_3924_));
 sg13g2_o21ai_1 _8899_ (.B1(_3925_),
    .Y(_3926_),
    .A1(_3862_),
    .A2(_3909_));
 sg13g2_nand3_1 _8900_ (.B(_3907_),
    .C(_3862_),
    .A(_3860_),
    .Y(_3927_));
 sg13g2_nor2_1 _8901_ (.A(_3927_),
    .B(_3868_),
    .Y(_3928_));
 sg13g2_nor2_1 _8902_ (.A(_3926_),
    .B(_3928_),
    .Y(_3929_));
 sg13g2_nor2_1 _8903_ (.A(_3909_),
    .B(_3863_),
    .Y(_3930_));
 sg13g2_nand3_1 _8904_ (.B(_3864_),
    .C(_3865_),
    .A(_3930_),
    .Y(_3931_));
 sg13g2_nand2_1 _8905_ (.Y(_3932_),
    .A(_3929_),
    .B(_3931_));
 sg13g2_nor2_1 _8906_ (.A(_2549_),
    .B(_3881_),
    .Y(_3933_));
 sg13g2_nor2_1 _8907_ (.A(_3625_),
    .B(_3924_),
    .Y(_3934_));
 sg13g2_nor2_1 _8908_ (.A(_3933_),
    .B(_3934_),
    .Y(_3935_));
 sg13g2_nand2_1 _8909_ (.Y(_3936_),
    .A(_3932_),
    .B(_3935_));
 sg13g2_inv_1 _8910_ (.Y(_3937_),
    .A(_3935_));
 sg13g2_nand3_1 _8911_ (.B(_3931_),
    .C(_3937_),
    .A(_3929_),
    .Y(_3938_));
 sg13g2_nand2_1 _8912_ (.Y(_3939_),
    .A(_3936_),
    .B(_3938_));
 sg13g2_nand2_1 _8913_ (.Y(_3940_),
    .A(_3939_),
    .B(_3442_));
 sg13g2_nand3_1 _8914_ (.B(_3938_),
    .C(_3469_),
    .A(_3936_),
    .Y(_3941_));
 sg13g2_nand2_1 _8915_ (.Y(_3942_),
    .A(_3940_),
    .B(_3941_));
 sg13g2_nand2_1 _8916_ (.Y(_3943_),
    .A(_3923_),
    .B(_3942_));
 sg13g2_inv_1 _8917_ (.Y(_3944_),
    .A(_3942_));
 sg13g2_nand3_1 _8918_ (.B(_3922_),
    .C(_3944_),
    .A(_3919_),
    .Y(_3945_));
 sg13g2_nand2_1 _8919_ (.Y(\generated._825[6] ),
    .A(_3943_),
    .B(_3945_));
 sg13g2_nor2_1 _8920_ (.A(_3915_),
    .B(_3942_),
    .Y(_3946_));
 sg13g2_nand2_1 _8921_ (.Y(_3947_),
    .A(_3918_),
    .B(_3946_));
 sg13g2_nand2b_1 _8922_ (.Y(_3948_),
    .B(_3936_),
    .A_N(_3934_));
 sg13g2_xnor2_1 _8923_ (.Y(_3949_),
    .A(_3469_),
    .B(_3948_));
 sg13g2_nor2b_1 _8924_ (.A(_3920_),
    .B_N(_3941_),
    .Y(_3950_));
 sg13g2_nand3_1 _8925_ (.B(_3949_),
    .C(_3950_),
    .A(_3947_),
    .Y(_3951_));
 sg13g2_nand2b_1 _8926_ (.Y(_3952_),
    .B(_3469_),
    .A_N(_3948_));
 sg13g2_nand2_1 _8927_ (.Y(\generated._825[7] ),
    .A(_3951_),
    .B(_3952_));
 sg13g2_nand2_1 _8928_ (.Y(\generated._825[8] ),
    .A(_3951_),
    .B(_3952_));
 sg13g2_nor2_1 _8929_ (.A(_1995_),
    .B(_1968_),
    .Y(_3953_));
 sg13g2_buf_1 _8930_ (.A(_3953_),
    .X(_3954_));
 sg13g2_nand2_1 _8931_ (.Y(_3955_),
    .A(net18),
    .B(_4242_));
 sg13g2_buf_1 _8932_ (.A(_1968_),
    .X(_3956_));
 sg13g2_xnor2_1 _8933_ (.Y(_3957_),
    .A(_4162_),
    .B(net95));
 sg13g2_buf_1 _8934_ (.A(_2006_),
    .X(_3958_));
 sg13g2_xor2_1 _8935_ (.B(_4231_),
    .A(_4241_),
    .X(_3959_));
 sg13g2_a221oi_1 _8936_ (.B2(_3959_),
    .C1(_0909_),
    .B1(net16),
    .A1(net21),
    .Y(_3960_),
    .A2(_3957_));
 sg13g2_buf_1 _8937_ (.A(_0755_),
    .X(_3961_));
 sg13g2_buf_1 _8938_ (.A(_0785_),
    .X(_3962_));
 sg13g2_nor2_1 _8939_ (.A(net69),
    .B(_0787_),
    .Y(_3963_));
 sg13g2_a21oi_1 _8940_ (.A1(net69),
    .A2(_0045_),
    .Y(_3964_),
    .B1(_3963_));
 sg13g2_nor2_1 _8941_ (.A(net67),
    .B(_3964_),
    .Y(_3965_));
 sg13g2_a21oi_1 _8942_ (.A1(net67),
    .A2(_0765_),
    .Y(_3966_),
    .B1(_3965_));
 sg13g2_inv_1 _8943_ (.Y(_3967_),
    .A(_0793_));
 sg13g2_nor2_1 _8944_ (.A(_0791_),
    .B(_3967_),
    .Y(_3968_));
 sg13g2_nor2_1 _8945_ (.A(net40),
    .B(_3968_),
    .Y(_3969_));
 sg13g2_xor2_1 _8946_ (.B(_3969_),
    .A(_3966_),
    .X(_3970_));
 sg13g2_xnor2_1 _8947_ (.Y(_3971_),
    .A(_1026_),
    .B(_3970_));
 sg13g2_nand2_1 _8948_ (.Y(_3972_),
    .A(_0795_),
    .B(_0804_));
 sg13g2_nand2_1 _8949_ (.Y(_3973_),
    .A(_0801_),
    .B(_3972_));
 sg13g2_xnor2_1 _8950_ (.Y(_3974_),
    .A(_3971_),
    .B(_3973_));
 sg13g2_a22oi_1 _8951_ (.Y(\generated._885[3] ),
    .B1(net50),
    .B2(_3974_),
    .A2(_3960_),
    .A1(_3955_));
 sg13g2_buf_1 _8952_ (.A(_0740_),
    .X(_3975_));
 sg13g2_buf_1 _8953_ (.A(net69),
    .X(_3976_));
 sg13g2_inv_1 _8954_ (.Y(_3977_),
    .A(_0046_));
 sg13g2_nor2_1 _8955_ (.A(net69),
    .B(_0045_),
    .Y(_3978_));
 sg13g2_a21oi_1 _8956_ (.A1(net49),
    .A2(_3977_),
    .Y(_3979_),
    .B1(_3978_));
 sg13g2_nor2_1 _8957_ (.A(net66),
    .B(_0789_),
    .Y(_3980_));
 sg13g2_a21oi_1 _8958_ (.A1(net66),
    .A2(_3979_),
    .Y(_3981_),
    .B1(_3980_));
 sg13g2_inv_1 _8959_ (.Y(_3982_),
    .A(_3968_));
 sg13g2_nor2_1 _8960_ (.A(_3966_),
    .B(_3982_),
    .Y(_3983_));
 sg13g2_nor2_1 _8961_ (.A(net40),
    .B(_3983_),
    .Y(_3984_));
 sg13g2_xor2_1 _8962_ (.B(_3984_),
    .A(_3981_),
    .X(_3985_));
 sg13g2_xnor2_1 _8963_ (.Y(_3986_),
    .A(_1079_),
    .B(_3985_));
 sg13g2_nor2b_1 _8964_ (.A(_0105_),
    .B_N(_3970_),
    .Y(_3987_));
 sg13g2_a21o_1 _8965_ (.A2(_3971_),
    .A1(_3973_),
    .B1(_3987_),
    .X(_3988_));
 sg13g2_xnor2_1 _8966_ (.Y(_3989_),
    .A(_3986_),
    .B(_3988_));
 sg13g2_xnor2_1 _8967_ (.Y(_3990_),
    .A(net79),
    .B(_4296_));
 sg13g2_o21ai_1 _8968_ (.B1(_0758_),
    .Y(_3991_),
    .A1(_2245_),
    .A2(_2069_));
 sg13g2_a221oi_1 _8969_ (.B2(net18),
    .C1(_3991_),
    .B1(net94),
    .A1(net16),
    .Y(_3992_),
    .A2(_3990_));
 sg13g2_a21oi_1 _8970_ (.A1(_3989_),
    .A2(_3961_),
    .Y(\generated._885[4] ),
    .B1(_3992_));
 sg13g2_nand2_1 _8971_ (.Y(_3993_),
    .A(_2799_),
    .B(net18));
 sg13g2_a221oi_1 _8972_ (.B2(_2757_),
    .C1(net52),
    .B1(net16),
    .A1(_2231_),
    .Y(_3994_),
    .A2(net21));
 sg13g2_nand2_1 _8973_ (.Y(_3995_),
    .A(net49),
    .B(_0047_));
 sg13g2_o21ai_1 _8974_ (.B1(_3995_),
    .Y(_3996_),
    .A1(net49),
    .A2(_3977_));
 sg13g2_nor2_1 _8975_ (.A(net66),
    .B(_3964_),
    .Y(_3997_));
 sg13g2_a21oi_2 _8976_ (.B1(_3997_),
    .Y(_3998_),
    .A2(_3996_),
    .A1(net66));
 sg13g2_inv_1 _8977_ (.Y(_3999_),
    .A(_3983_));
 sg13g2_nor2_1 _8978_ (.A(_3981_),
    .B(_3999_),
    .Y(_4000_));
 sg13g2_nor2_1 _8979_ (.A(net40),
    .B(_4000_),
    .Y(_4001_));
 sg13g2_xor2_1 _8980_ (.B(_4001_),
    .A(_3998_),
    .X(_4002_));
 sg13g2_xnor2_1 _8981_ (.Y(_4003_),
    .A(_1034_),
    .B(_4002_));
 sg13g2_nor2b_1 _8982_ (.A(_0036_),
    .B_N(_3985_),
    .Y(_4004_));
 sg13g2_a21o_1 _8983_ (.A2(_3986_),
    .A1(_3988_),
    .B1(_4004_),
    .X(_4005_));
 sg13g2_xnor2_1 _8984_ (.Y(_4006_),
    .A(_4003_),
    .B(_4005_));
 sg13g2_a22oi_1 _8985_ (.Y(\generated._885[5] ),
    .B1(net50),
    .B2(_4006_),
    .A2(_3994_),
    .A1(_3993_));
 sg13g2_nand2_1 _8986_ (.Y(_4007_),
    .A(_2780_),
    .B(net18));
 sg13g2_a221oi_1 _8987_ (.B2(_4305_),
    .C1(net52),
    .B1(net16),
    .A1(_2263_),
    .Y(_4008_),
    .A2(net21));
 sg13g2_nand2_1 _8988_ (.Y(_4009_),
    .A(_0773_),
    .B(net49));
 sg13g2_o21ai_1 _8989_ (.B1(_4009_),
    .Y(_4010_),
    .A1(net49),
    .A2(_0047_));
 sg13g2_nor2_1 _8990_ (.A(net67),
    .B(_4010_),
    .Y(_4011_));
 sg13g2_a21oi_1 _8991_ (.A1(net67),
    .A2(_3979_),
    .Y(_4012_),
    .B1(_4011_));
 sg13g2_inv_1 _8992_ (.Y(_4013_),
    .A(_4000_));
 sg13g2_nor2_1 _8993_ (.A(_3998_),
    .B(_4013_),
    .Y(_4014_));
 sg13g2_nor2_1 _8994_ (.A(net32),
    .B(_4014_),
    .Y(_4015_));
 sg13g2_xor2_1 _8995_ (.B(_4015_),
    .A(_4012_),
    .X(_4016_));
 sg13g2_xnor2_1 _8996_ (.Y(_4017_),
    .A(_1033_),
    .B(_4016_));
 sg13g2_nor2b_1 _8997_ (.A(_0037_),
    .B_N(_4002_),
    .Y(_4018_));
 sg13g2_a21o_1 _8998_ (.A2(_4003_),
    .A1(_4005_),
    .B1(_4018_),
    .X(_4019_));
 sg13g2_xnor2_1 _8999_ (.Y(_4020_),
    .A(_4017_),
    .B(_4019_));
 sg13g2_a22oi_1 _9000_ (.Y(\generated._885[6] ),
    .B1(net50),
    .B2(_4020_),
    .A2(_4008_),
    .A1(_4007_));
 sg13g2_nand2_1 _9001_ (.Y(_4021_),
    .A(_2777_),
    .B(net18));
 sg13g2_a221oi_1 _9002_ (.B2(net21),
    .C1(net52),
    .B1(_2296_),
    .A1(net16),
    .Y(_4022_),
    .A2(_2759_));
 sg13g2_nand2_1 _9003_ (.Y(_4023_),
    .A(net66),
    .B(_0039_));
 sg13g2_inv_1 _9004_ (.Y(_4024_),
    .A(_4023_));
 sg13g2_a21oi_1 _9005_ (.A1(_3996_),
    .A2(net67),
    .Y(_4025_),
    .B1(_4024_));
 sg13g2_nor3_1 _9006_ (.A(_3998_),
    .B(_4012_),
    .C(_4013_),
    .Y(_4026_));
 sg13g2_inv_1 _9007_ (.Y(_4027_),
    .A(_4026_));
 sg13g2_o21ai_1 _9008_ (.B1(_0839_),
    .Y(_4028_),
    .A1(_4025_),
    .A2(_4027_));
 sg13g2_a21oi_1 _9009_ (.A1(_4027_),
    .A2(_4025_),
    .Y(_4029_),
    .B1(_4028_));
 sg13g2_a21o_1 _9010_ (.A2(_4025_),
    .A1(net32),
    .B1(_4029_),
    .X(_4030_));
 sg13g2_xnor2_1 _9011_ (.Y(_4031_),
    .A(_1045_),
    .B(_4030_));
 sg13g2_nor2b_1 _9012_ (.A(_0038_),
    .B_N(_4016_),
    .Y(_4032_));
 sg13g2_a21o_1 _9013_ (.A2(_4017_),
    .A1(_4019_),
    .B1(_4032_),
    .X(_4033_));
 sg13g2_xnor2_1 _9014_ (.Y(_4034_),
    .A(_4031_),
    .B(_4033_));
 sg13g2_a22oi_1 _9015_ (.Y(\generated._885[7] ),
    .B1(net50),
    .B2(_4034_),
    .A2(_4022_),
    .A1(_4021_));
 sg13g2_nand2_1 _9016_ (.Y(_4035_),
    .A(_2767_),
    .B(net18));
 sg13g2_inv_1 _9017_ (.Y(_4036_),
    .A(_2764_));
 sg13g2_a221oi_1 _9018_ (.B2(_3958_),
    .C1(net52),
    .B1(_4036_),
    .A1(_1294_),
    .Y(_4037_),
    .A2(_2291_));
 sg13g2_o21ai_1 _9019_ (.B1(_4023_),
    .Y(_4038_),
    .A1(_3975_),
    .A2(_4010_));
 sg13g2_xnor2_1 _9020_ (.Y(_4039_),
    .A(_4038_),
    .B(_4028_));
 sg13g2_xnor2_1 _9021_ (.Y(_4040_),
    .A(_1055_),
    .B(_4039_));
 sg13g2_nor2b_1 _9022_ (.A(_0043_),
    .B_N(_4030_),
    .Y(_4041_));
 sg13g2_a21o_1 _9023_ (.A2(_4031_),
    .A1(_4033_),
    .B1(_4041_),
    .X(_4042_));
 sg13g2_xnor2_1 _9024_ (.Y(_4043_),
    .A(_4040_),
    .B(_4042_));
 sg13g2_a22oi_1 _9025_ (.Y(\generated._885[8] ),
    .B1(net50),
    .B2(_4043_),
    .A2(_4037_),
    .A1(_4035_));
 sg13g2_inv_1 _9026_ (.Y(_4044_),
    .A(_4039_));
 sg13g2_a22oi_1 _9027_ (.Y(_4045_),
    .B1(_4040_),
    .B2(_4042_),
    .A2(_4044_),
    .A1(_1169_));
 sg13g2_nand3b_1 _9028_ (.B(_4026_),
    .C(_4038_),
    .Y(_4046_),
    .A_N(_4025_));
 sg13g2_xor2_1 _9029_ (.B(_4046_),
    .A(\generated._67[9] ),
    .X(_4047_));
 sg13g2_o21ai_1 _9030_ (.B1(_0773_),
    .Y(_4048_),
    .A1(net32),
    .A2(_4047_));
 sg13g2_xnor2_1 _9031_ (.Y(_4049_),
    .A(_1227_),
    .B(_4048_));
 sg13g2_o21ai_1 _9032_ (.B1(_0909_),
    .Y(_4050_),
    .A1(_4049_),
    .A2(_4045_));
 sg13g2_a21oi_1 _9033_ (.A1(_4045_),
    .A2(_4049_),
    .Y(\generated._885[9] ),
    .B1(_4050_));
 sg13g2_xnor2_1 _9034_ (.Y(_4051_),
    .A(_0120_),
    .B(_3957_));
 sg13g2_nor2_1 _9035_ (.A(_4051_),
    .B(_2010_),
    .Y(_4052_));
 sg13g2_a221oi_1 _9036_ (.B2(_3957_),
    .C1(_4052_),
    .B1(net18),
    .A1(net21),
    .Y(_4053_),
    .A2(_3959_));
 sg13g2_nand2_1 _9037_ (.Y(_4054_),
    .A(_0830_),
    .B(\generated._67[2] ));
 sg13g2_nand2_1 _9038_ (.Y(_4055_),
    .A(_0834_),
    .B(_4054_));
 sg13g2_inv_1 _9039_ (.Y(_4056_),
    .A(_0038_));
 sg13g2_nand2_1 _9040_ (.Y(_4057_),
    .A(_4056_),
    .B(net69));
 sg13g2_o21ai_1 _9041_ (.B1(_4057_),
    .Y(_4058_),
    .A1(_0786_),
    .A2(_0037_));
 sg13g2_nor2_1 _9042_ (.A(net67),
    .B(_4058_),
    .Y(_4059_));
 sg13g2_a21oi_1 _9043_ (.A1(net67),
    .A2(_0815_),
    .Y(_4060_),
    .B1(_4059_));
 sg13g2_inv_1 _9044_ (.Y(_4061_),
    .A(_0828_));
 sg13g2_nor2_1 _9045_ (.A(_0827_),
    .B(_4061_),
    .Y(_4062_));
 sg13g2_nor2_1 _9046_ (.A(net40),
    .B(_4062_),
    .Y(_4063_));
 sg13g2_xnor2_1 _9047_ (.Y(_4064_),
    .A(_4060_),
    .B(_4063_));
 sg13g2_xnor2_1 _9048_ (.Y(_4065_),
    .A(_0035_),
    .B(_4064_));
 sg13g2_a21oi_1 _9049_ (.A1(_4055_),
    .A2(_4065_),
    .Y(_4066_),
    .B1(_0758_));
 sg13g2_o21ai_1 _9050_ (.B1(_4066_),
    .Y(_4067_),
    .A1(_4055_),
    .A2(_4065_));
 sg13g2_o21ai_1 _9051_ (.B1(_4067_),
    .Y(\generated._934[3] ),
    .A1(net54),
    .A2(_4053_));
 sg13g2_nand2_1 _9052_ (.Y(_4068_),
    .A(_0786_),
    .B(_0043_));
 sg13g2_o21ai_1 _9053_ (.B1(_4068_),
    .Y(_4069_),
    .A1(net49),
    .A2(_4056_));
 sg13g2_nor2_1 _9054_ (.A(net81),
    .B(_0825_),
    .Y(_4070_));
 sg13g2_a21oi_1 _9055_ (.A1(net66),
    .A2(_4069_),
    .Y(_4071_),
    .B1(_4070_));
 sg13g2_inv_1 _9056_ (.Y(_4072_),
    .A(_4062_));
 sg13g2_nor2_1 _9057_ (.A(_4060_),
    .B(_4072_),
    .Y(_4073_));
 sg13g2_nor2_1 _9058_ (.A(net40),
    .B(_4073_),
    .Y(_4074_));
 sg13g2_xnor2_1 _9059_ (.Y(_4075_),
    .A(_4071_),
    .B(_4074_));
 sg13g2_xnor2_1 _9060_ (.Y(_4076_),
    .A(_0042_),
    .B(_4075_));
 sg13g2_nand2_1 _9061_ (.Y(_4077_),
    .A(_4055_),
    .B(_4065_));
 sg13g2_nand2_1 _9062_ (.Y(_4078_),
    .A(_4064_),
    .B(\generated._67[3] ));
 sg13g2_nand2_1 _9063_ (.Y(_4079_),
    .A(_4077_),
    .B(_4078_));
 sg13g2_xnor2_1 _9064_ (.Y(_4080_),
    .A(_4076_),
    .B(_4079_));
 sg13g2_inv_1 _9065_ (.Y(_4081_),
    .A(_3953_));
 sg13g2_a22oi_1 _9066_ (.Y(_4082_),
    .B1(_2006_),
    .B2(_2247_),
    .A2(_3990_),
    .A1(_3956_));
 sg13g2_o21ai_1 _9067_ (.B1(_4082_),
    .Y(_4083_),
    .A1(_2245_),
    .A2(_4081_));
 sg13g2_nor2_1 _9068_ (.A(_0756_),
    .B(_4083_),
    .Y(_4084_));
 sg13g2_a21oi_1 _9069_ (.A1(_4080_),
    .A2(_0756_),
    .Y(\generated._934[4] ),
    .B1(_4084_));
 sg13g2_nand2_1 _9070_ (.Y(_4085_),
    .A(net31),
    .B(net16));
 sg13g2_a221oi_1 _9071_ (.B2(_2231_),
    .C1(net52),
    .B1(net18),
    .A1(net21),
    .Y(_4086_),
    .A2(_2757_));
 sg13g2_nand2_1 _9072_ (.Y(_4087_),
    .A(_1169_),
    .B(net49));
 sg13g2_o21ai_1 _9073_ (.B1(_4087_),
    .Y(_4088_),
    .A1(net49),
    .A2(_0043_));
 sg13g2_inv_1 _9074_ (.Y(_4089_),
    .A(_4088_));
 sg13g2_nor2_1 _9075_ (.A(net66),
    .B(_4058_),
    .Y(_4090_));
 sg13g2_a21oi_1 _9076_ (.A1(net66),
    .A2(_4089_),
    .Y(_4091_),
    .B1(_4090_));
 sg13g2_inv_1 _9077_ (.Y(_4092_),
    .A(_4073_));
 sg13g2_nor2_1 _9078_ (.A(_4071_),
    .B(_4092_),
    .Y(_4093_));
 sg13g2_nor2_1 _9079_ (.A(_0792_),
    .B(_4093_),
    .Y(_4094_));
 sg13g2_xnor2_1 _9080_ (.Y(_4095_),
    .A(_4091_),
    .B(_4094_));
 sg13g2_xnor2_1 _9081_ (.Y(_4096_),
    .A(_0044_),
    .B(_4095_));
 sg13g2_nand2_1 _9082_ (.Y(_4097_),
    .A(_4079_),
    .B(_4076_));
 sg13g2_nand2_1 _9083_ (.Y(_4098_),
    .A(_4075_),
    .B(\generated._67[4] ));
 sg13g2_nand2_1 _9084_ (.Y(_4099_),
    .A(_4097_),
    .B(_4098_));
 sg13g2_xnor2_1 _9085_ (.Y(_4100_),
    .A(_4096_),
    .B(_4099_));
 sg13g2_a22oi_1 _9086_ (.Y(\generated._934[5] ),
    .B1(net50),
    .B2(_4100_),
    .A2(_4086_),
    .A1(_4085_));
 sg13g2_nand2_1 _9087_ (.Y(_4101_),
    .A(_2266_),
    .B(net16));
 sg13g2_a221oi_1 _9088_ (.B2(_2263_),
    .C1(net52),
    .B1(_3954_),
    .A1(_4305_),
    .Y(_4102_),
    .A2(net21));
 sg13g2_nand2_1 _9089_ (.Y(_4103_),
    .A(_3976_),
    .B(_1262_));
 sg13g2_o21ai_1 _9090_ (.B1(_4103_),
    .Y(_4104_),
    .A1(_3976_),
    .A2(_1169_));
 sg13g2_mux2_1 _9091_ (.A0(_4104_),
    .A1(_4069_),
    .S(net67),
    .X(_4105_));
 sg13g2_inv_1 _9092_ (.Y(_4106_),
    .A(_4091_));
 sg13g2_a21oi_1 _9093_ (.A1(_4093_),
    .A2(_4106_),
    .Y(_4107_),
    .B1(_0792_));
 sg13g2_xor2_1 _9094_ (.B(_4107_),
    .A(_4105_),
    .X(_4108_));
 sg13g2_xnor2_1 _9095_ (.Y(_4109_),
    .A(_0045_),
    .B(_4108_));
 sg13g2_nand2_1 _9096_ (.Y(_4110_),
    .A(_4099_),
    .B(_4096_));
 sg13g2_nand2_1 _9097_ (.Y(_4111_),
    .A(_4095_),
    .B(\generated._67[5] ));
 sg13g2_nand2_1 _9098_ (.Y(_4112_),
    .A(_4110_),
    .B(_4111_));
 sg13g2_xnor2_1 _9099_ (.Y(_4113_),
    .A(_4109_),
    .B(_4112_));
 sg13g2_a22oi_1 _9100_ (.Y(\generated._934[6] ),
    .B1(net50),
    .B2(_4113_),
    .A2(_4102_),
    .A1(_4101_));
 sg13g2_nand2_1 _9101_ (.Y(_4114_),
    .A(_2314_),
    .B(_3958_));
 sg13g2_a221oi_1 _9102_ (.B2(_3954_),
    .C1(net52),
    .B1(_2296_),
    .A1(net21),
    .Y(_4115_),
    .A2(_2759_));
 sg13g2_nand2_1 _9103_ (.Y(_4116_),
    .A(_3975_),
    .B(_1262_));
 sg13g2_inv_1 _9104_ (.Y(_4117_),
    .A(_4116_));
 sg13g2_a21oi_1 _9105_ (.A1(_4089_),
    .A2(_3962_),
    .Y(_4118_),
    .B1(_4117_));
 sg13g2_inv_1 _9106_ (.Y(_4119_),
    .A(_4118_));
 sg13g2_nand3b_1 _9107_ (.B(_4093_),
    .C(_4105_),
    .Y(_4120_),
    .A_N(_4091_));
 sg13g2_nand2_1 _9108_ (.Y(_4121_),
    .A(_4120_),
    .B(_0839_));
 sg13g2_xnor2_1 _9109_ (.Y(_4122_),
    .A(_4119_),
    .B(_4121_));
 sg13g2_xnor2_1 _9110_ (.Y(_4123_),
    .A(_0046_),
    .B(_4122_));
 sg13g2_nand2_1 _9111_ (.Y(_4124_),
    .A(_4112_),
    .B(_4109_));
 sg13g2_nand2_1 _9112_ (.Y(_4125_),
    .A(_4108_),
    .B(\generated._67[6] ));
 sg13g2_nand2_1 _9113_ (.Y(_4126_),
    .A(_4124_),
    .B(_4125_));
 sg13g2_xnor2_1 _9114_ (.Y(_4127_),
    .A(_4123_),
    .B(_4126_));
 sg13g2_a22oi_1 _9115_ (.Y(\generated._934[7] ),
    .B1(_3961_),
    .B2(_4127_),
    .A2(_4115_),
    .A1(_4114_));
 sg13g2_nand2_1 _9116_ (.Y(_4128_),
    .A(_2317_),
    .B(net16));
 sg13g2_a221oi_1 _9117_ (.B2(_3953_),
    .C1(_0755_),
    .B1(_2293_),
    .A1(_3956_),
    .Y(_4129_),
    .A2(_4036_));
 sg13g2_a21oi_1 _9118_ (.A1(_4104_),
    .A2(_3962_),
    .Y(_4130_),
    .B1(_4117_));
 sg13g2_o21ai_1 _9119_ (.B1(_4121_),
    .Y(_4131_),
    .A1(net32),
    .A2(_4119_));
 sg13g2_xor2_1 _9120_ (.B(_4131_),
    .A(_4130_),
    .X(_4132_));
 sg13g2_xor2_1 _9121_ (.B(_4132_),
    .A(_0047_),
    .X(_4133_));
 sg13g2_nand2_1 _9122_ (.Y(_4134_),
    .A(_4126_),
    .B(_4123_));
 sg13g2_nand2_1 _9123_ (.Y(_4135_),
    .A(_4122_),
    .B(\generated._67[7] ));
 sg13g2_nand2_1 _9124_ (.Y(_4136_),
    .A(_4134_),
    .B(_4135_));
 sg13g2_xnor2_1 _9125_ (.Y(_4137_),
    .A(_4133_),
    .B(_4136_));
 sg13g2_a22oi_1 _9126_ (.Y(\generated._934[8] ),
    .B1(net50),
    .B2(_4137_),
    .A2(_4129_),
    .A1(_4128_));
 sg13g2_nor3_1 _9127_ (.A(_4118_),
    .B(_4130_),
    .C(_4120_),
    .Y(_4138_));
 sg13g2_xnor2_1 _9128_ (.Y(_4139_),
    .A(_1067_),
    .B(_4138_));
 sg13g2_nand2_1 _9129_ (.Y(_4140_),
    .A(net32),
    .B(_1262_));
 sg13g2_o21ai_1 _9130_ (.B1(_4140_),
    .Y(_4141_),
    .A1(net32),
    .A2(_4139_));
 sg13g2_xnor2_1 _9131_ (.Y(_4142_),
    .A(_0039_),
    .B(_4141_));
 sg13g2_inv_1 _9132_ (.Y(_4143_),
    .A(_4132_));
 sg13g2_a22oi_1 _9133_ (.Y(_4144_),
    .B1(_4133_),
    .B2(_4136_),
    .A2(_4143_),
    .A1(\generated._67[8] ));
 sg13g2_xor2_1 _9134_ (.B(_4144_),
    .A(_4142_),
    .X(_4145_));
 sg13g2_o21ai_1 _9135_ (.B1(_0758_),
    .Y(_4146_),
    .A1(_1978_),
    .A2(_2301_));
 sg13g2_o21ai_1 _9136_ (.B1(_4146_),
    .Y(\generated._934[9] ),
    .A1(net41),
    .A2(_4145_));
 sg13g2_dfrbp_1 _9137_ (.CLK(clknet_leaf_14_clk),
    .RESET_B(net122),
    .D(_0004_),
    .Q_N(_4578_),
    .Q(_0010_));
 sg13g2_dfrbp_1 _9138_ (.CLK(clknet_leaf_14_clk),
    .RESET_B(net123),
    .D(_0005_),
    .Q_N(_4579_),
    .Q(_0011_));
 sg13g2_dfrbp_1 _9139_ (.CLK(clknet_leaf_14_clk),
    .RESET_B(net124),
    .D(_0006_),
    .Q_N(_4577_),
    .Q(_0012_));
 sg13g2_dfrbp_1 _9140_ (.CLK(clknet_leaf_14_clk),
    .RESET_B(net125),
    .D(_0127_),
    .Q_N(_4576_),
    .Q(_0013_));
 sg13g2_dfrbp_1 _9141_ (.CLK(clknet_leaf_13_clk),
    .RESET_B(net126),
    .D(_0128_),
    .Q_N(_4575_),
    .Q(_0014_));
 sg13g2_dfrbp_1 _9142_ (.CLK(clknet_leaf_14_clk),
    .RESET_B(net127),
    .D(_0129_),
    .Q_N(_4580_),
    .Q(_0015_));
 sg13g2_dfrbp_1 _9143_ (.CLK(clknet_leaf_14_clk),
    .RESET_B(net128),
    .D(_0000_),
    .Q_N(_4581_),
    .Q(_0007_));
 sg13g2_dfrbp_1 _9144_ (.CLK(clknet_leaf_17_clk),
    .RESET_B(net129),
    .D(_0001_),
    .Q_N(_4582_),
    .Q(_0008_));
 sg13g2_dfrbp_1 _9145_ (.CLK(clknet_leaf_13_clk),
    .RESET_B(net130),
    .D(_0002_),
    .Q_N(_4574_),
    .Q(_0009_));
 sg13g2_buf_2 clkbuf_leaf_0_clk (.A(clknet_3_0__leaf_clk),
    .X(clknet_leaf_0_clk));
 sg13g2_tiehi _9137__122 (.L_HI(net122));
 sg13g2_buf_1 _9148_ (.A(net106),
    .X(uio_oe[0]));
 sg13g2_buf_1 _9149_ (.A(net107),
    .X(uio_oe[1]));
 sg13g2_buf_1 _9150_ (.A(net108),
    .X(uio_oe[2]));
 sg13g2_buf_1 _9151_ (.A(net109),
    .X(uio_oe[3]));
 sg13g2_buf_1 _9152_ (.A(net110),
    .X(uio_oe[4]));
 sg13g2_buf_1 _9153_ (.A(net111),
    .X(uio_oe[5]));
 sg13g2_buf_1 _9154_ (.A(net112),
    .X(uio_oe[6]));
 sg13g2_buf_1 _9155_ (.A(net113),
    .X(uio_oe[7]));
 sg13g2_buf_1 _9156_ (.A(net114),
    .X(uio_out[0]));
 sg13g2_buf_1 _9157_ (.A(net115),
    .X(uio_out[1]));
 sg13g2_buf_1 _9158_ (.A(net116),
    .X(uio_out[2]));
 sg13g2_buf_1 _9159_ (.A(net117),
    .X(uio_out[3]));
 sg13g2_buf_1 _9160_ (.A(net118),
    .X(uio_out[4]));
 sg13g2_buf_1 _9161_ (.A(net119),
    .X(uio_out[5]));
 sg13g2_buf_1 _9162_ (.A(net120),
    .X(uio_out[6]));
 sg13g2_buf_1 _9163_ (.A(net121),
    .X(uio_out[7]));
 sg13g2_buf_1 _9164_ (.A(\generated._111 ),
    .X(net5));
 sg13g2_buf_1 _9165_ (.A(\generated._119 ),
    .X(net9));
 sg13g2_dfrbp_1 \generated._1020[0]$_SDFF_PP0_  (.CLK(clknet_leaf_0_clk),
    .RESET_B(net131),
    .D(_0130_),
    .Q_N(_0097_),
    .Q(\generated._1020[0] ));
 sg13g2_dfrbp_1 \generated._1020[1]$_SDFF_PP0_  (.CLK(clknet_leaf_0_clk),
    .RESET_B(net132),
    .D(_0131_),
    .Q_N(_0098_),
    .Q(\generated._1020[1] ));
 sg13g2_dfrbp_1 \generated._1020[2]$_SDFF_PP0_  (.CLK(clknet_leaf_0_clk),
    .RESET_B(net133),
    .D(_0132_),
    .Q_N(_0099_),
    .Q(\generated._1020[2] ));
 sg13g2_dfrbp_1 \generated._1020[3]$_DFF_P_  (.CLK(clknet_leaf_0_clk),
    .RESET_B(net134),
    .D(\generated._1019[3] ),
    .Q_N(_0100_),
    .Q(\generated._1020[3] ));
 sg13g2_dfrbp_1 \generated._1020[4]$_DFF_P_  (.CLK(clknet_leaf_3_clk),
    .RESET_B(net135),
    .D(\generated._1019[4] ),
    .Q_N(_0017_),
    .Q(\generated._1020[4] ));
 sg13g2_dfrbp_1 \generated._1020[5]$_DFF_P_  (.CLK(clknet_leaf_3_clk),
    .RESET_B(net136),
    .D(\generated._1019[5] ),
    .Q_N(_0018_),
    .Q(\generated._1020[5] ));
 sg13g2_dfrbp_1 \generated._1020[6]$_DFF_P_  (.CLK(clknet_leaf_3_clk),
    .RESET_B(net137),
    .D(\generated._1019[6] ),
    .Q_N(_0019_),
    .Q(\generated._1020[6] ));
 sg13g2_dfrbp_1 \generated._1020[7]$_DFF_P_  (.CLK(clknet_leaf_3_clk),
    .RESET_B(net138),
    .D(\generated._1019[7] ),
    .Q_N(_0024_),
    .Q(\generated._1020[7] ));
 sg13g2_dfrbp_1 \generated._1020[8]$_DFF_P_  (.CLK(clknet_leaf_31_clk),
    .RESET_B(net139),
    .D(\generated._1019[8] ),
    .Q_N(_0027_),
    .Q(\generated._1020[8] ));
 sg13g2_dfrbp_1 \generated._1020[9]$_DFF_P_  (.CLK(clknet_leaf_31_clk),
    .RESET_B(net140),
    .D(\generated._1019[9] ),
    .Q_N(_0029_),
    .Q(\generated._1020[9] ));
 sg13g2_dfrbp_1 \generated._1070[0]$_SDFF_PP0_  (.CLK(clknet_leaf_34_clk),
    .RESET_B(net141),
    .D(_0133_),
    .Q_N(_0096_),
    .Q(\generated._1070[0] ));
 sg13g2_dfrbp_1 \generated._1070[1]$_SDFF_PP0_  (.CLK(clknet_leaf_34_clk),
    .RESET_B(net142),
    .D(_0134_),
    .Q_N(_0022_),
    .Q(\generated._1070[1] ));
 sg13g2_dfrbp_1 \generated._1070[2]$_SDFF_PP0_  (.CLK(clknet_leaf_34_clk),
    .RESET_B(net143),
    .D(_0135_),
    .Q_N(_0021_),
    .Q(\generated._1070[2] ));
 sg13g2_dfrbp_1 \generated._1070[3]$_DFF_P_  (.CLK(clknet_leaf_34_clk),
    .RESET_B(net144),
    .D(\generated._1069[3] ),
    .Q_N(_0016_),
    .Q(\generated._1070[3] ));
 sg13g2_dfrbp_1 \generated._1070[4]$_DFF_P_  (.CLK(clknet_leaf_34_clk),
    .RESET_B(net145),
    .D(\generated._1069[4] ),
    .Q_N(_0023_),
    .Q(\generated._1070[4] ));
 sg13g2_dfrbp_1 \generated._1070[5]$_DFF_P_  (.CLK(clknet_leaf_34_clk),
    .RESET_B(net146),
    .D(\generated._1069[5] ),
    .Q_N(_0026_),
    .Q(\generated._1070[5] ));
 sg13g2_dfrbp_1 \generated._1070[6]$_DFF_P_  (.CLK(clknet_leaf_34_clk),
    .RESET_B(net147),
    .D(\generated._1069[6] ),
    .Q_N(_0028_),
    .Q(\generated._1070[6] ));
 sg13g2_dfrbp_1 \generated._1070[7]$_DFF_P_  (.CLK(clknet_leaf_34_clk),
    .RESET_B(net148),
    .D(\generated._1069[7] ),
    .Q_N(_0030_),
    .Q(\generated._1070[7] ));
 sg13g2_dfrbp_1 \generated._1070[8]$_DFF_P_  (.CLK(clknet_leaf_32_clk),
    .RESET_B(net149),
    .D(\generated._1069[8] ),
    .Q_N(_0031_),
    .Q(\generated._1070[8] ));
 sg13g2_dfrbp_1 \generated._1070[9]$_DFF_P_  (.CLK(clknet_leaf_0_clk),
    .RESET_B(net150),
    .D(\generated._1069[9] ),
    .Q_N(_0020_),
    .Q(\generated._1070[9] ));
 sg13g2_dfrbp_1 \generated._1074[0]$_DFF_PN0_  (.CLK(clknet_leaf_3_clk),
    .RESET_B(net96),
    .D(\generated._1073[0] ),
    .Q_N(_4583_),
    .Q(\generated._1074[0] ));
 sg13g2_dfrbp_1 \generated._1074[1]$_DFF_PN0_  (.CLK(clknet_leaf_4_clk),
    .RESET_B(net97),
    .D(\generated._1073[1] ),
    .Q_N(_4584_),
    .Q(\generated._1074[1] ));
 sg13g2_dfrbp_1 \generated._1074[2]$_DFF_PN0_  (.CLK(clknet_leaf_4_clk),
    .RESET_B(net97),
    .D(\generated._1073[2] ),
    .Q_N(_4585_),
    .Q(\generated._1074[2] ));
 sg13g2_dfrbp_1 \generated._1074[3]$_DFF_PN0_  (.CLK(clknet_leaf_31_clk),
    .RESET_B(net96),
    .D(\generated._1073[3] ),
    .Q_N(_4573_),
    .Q(\generated._1074[3] ));
 sg13g2_dfrbp_1 \generated._1080[0]$_SDFF_PP0_  (.CLK(clknet_leaf_1_clk),
    .RESET_B(net151),
    .D(_0136_),
    .Q_N(_0088_),
    .Q(\generated._1080[0] ));
 sg13g2_dfrbp_1 \generated._1080[1]$_SDFF_PP0_  (.CLK(clknet_leaf_1_clk),
    .RESET_B(net152),
    .D(_0137_),
    .Q_N(_4572_),
    .Q(\generated._1080[1] ));
 sg13g2_dfrbp_1 \generated._1080[2]$_SDFF_PP0_  (.CLK(clknet_leaf_1_clk),
    .RESET_B(net153),
    .D(_0138_),
    .Q_N(_4571_),
    .Q(\generated._1080[2] ));
 sg13g2_dfrbp_1 \generated._1080[3]$_SDFF_PP0_  (.CLK(clknet_leaf_1_clk),
    .RESET_B(net154),
    .D(_0139_),
    .Q_N(_4570_),
    .Q(\generated._1080[3] ));
 sg13g2_dfrbp_1 \generated._1080[4]$_SDFF_PP0_  (.CLK(clknet_leaf_1_clk),
    .RESET_B(net155),
    .D(_0140_),
    .Q_N(_4569_),
    .Q(\generated._1080[4] ));
 sg13g2_dfrbp_1 \generated._1080[5]$_SDFF_PP0_  (.CLK(clknet_leaf_1_clk),
    .RESET_B(net156),
    .D(_0141_),
    .Q_N(_4568_),
    .Q(\generated._1080[5] ));
 sg13g2_dfrbp_1 \generated._1080[6]$_SDFF_PP0_  (.CLK(clknet_leaf_0_clk),
    .RESET_B(net157),
    .D(_0142_),
    .Q_N(_4567_),
    .Q(\generated._1080[6] ));
 sg13g2_dfrbp_1 \generated._1080[7]$_SDFF_PP0_  (.CLK(clknet_leaf_1_clk),
    .RESET_B(net158),
    .D(_0143_),
    .Q_N(_4566_),
    .Q(\generated._1080[7] ));
 sg13g2_dfrbp_1 \generated._1080[8]$_SDFF_PP0_  (.CLK(clknet_leaf_2_clk),
    .RESET_B(net159),
    .D(_0144_),
    .Q_N(_4565_),
    .Q(\generated._1080[8] ));
 sg13g2_dfrbp_1 \generated._1080[9]$_SDFF_PP0_  (.CLK(clknet_leaf_2_clk),
    .RESET_B(net160),
    .D(_0145_),
    .Q_N(_4586_),
    .Q(\generated._1080[9] ));
 sg13g2_dfrbp_1 \generated._111$_DFF_PN0_  (.CLK(clknet_leaf_16_clk),
    .RESET_B(net102),
    .D(\generated._108 ),
    .Q_N(_4587_),
    .Q(\generated._111 ));
 sg13g2_dfrbp_1 \generated._1150[0]$_DFF_PN0_  (.CLK(clknet_leaf_17_clk),
    .RESET_B(net102),
    .D(\generated._1149[0] ),
    .Q_N(_4588_),
    .Q(net6));
 sg13g2_dfrbp_1 \generated._1150[1]$_DFF_PN0_  (.CLK(clknet_leaf_17_clk),
    .RESET_B(net102),
    .D(\generated._1149[1] ),
    .Q_N(_4589_),
    .Q(net2));
 sg13g2_dfrbp_1 \generated._119$_DFF_PN0_  (.CLK(clknet_leaf_16_clk),
    .RESET_B(net104),
    .D(\generated._118 ),
    .Q_N(_4590_),
    .Q(\generated._119 ));
 sg13g2_dfrbp_1 \generated._222[1]$_DFF_P_  (.CLK(clknet_leaf_16_clk),
    .RESET_B(net161),
    .D(_0003_),
    .Q_N(_4591_),
    .Q(\generated._1144[0] ));
 sg13g2_dfrbp_1 \generated._232[0]$_DFF_PN0_  (.CLK(clknet_leaf_17_clk),
    .RESET_B(net102),
    .D(\generated._231[0] ),
    .Q_N(_4592_),
    .Q(net8));
 sg13g2_dfrbp_1 \generated._232[1]$_DFF_PN0_  (.CLK(clknet_leaf_17_clk),
    .RESET_B(net102),
    .D(\generated._231[1] ),
    .Q_N(_4593_),
    .Q(net4));
 sg13g2_dfrbp_1 \generated._285[0]$_DFF_PN0_  (.CLK(clknet_leaf_17_clk),
    .RESET_B(net102),
    .D(\generated._284[0] ),
    .Q_N(_4594_),
    .Q(net7));
 sg13g2_dfrbp_1 \generated._285[1]$_DFF_PN0_  (.CLK(clknet_leaf_17_clk),
    .RESET_B(net102),
    .D(\generated._284[1] ),
    .Q_N(_4564_),
    .Q(net3));
 sg13g2_dfrbp_1 \generated._287[0]$_SDFFE_PP0N_  (.CLK(clknet_leaf_10_clk),
    .RESET_B(net162),
    .D(_0146_),
    .Q_N(_4563_),
    .Q(\generated._14[0] ));
 sg13g2_dfrbp_1 \generated._287[1]$_SDFFE_PP0N_  (.CLK(clknet_leaf_10_clk),
    .RESET_B(net163),
    .D(_0147_),
    .Q_N(_4562_),
    .Q(\generated._14[1] ));
 sg13g2_dfrbp_1 \generated._287[2]$_SDFFE_PP0N_  (.CLK(clknet_leaf_10_clk),
    .RESET_B(net164),
    .D(_0148_),
    .Q_N(_4561_),
    .Q(\generated._14[2] ));
 sg13g2_dfrbp_1 \generated._287[3]$_SDFFE_PP0N_  (.CLK(clknet_leaf_10_clk),
    .RESET_B(net165),
    .D(_0149_),
    .Q_N(_4560_),
    .Q(\generated._14[3] ));
 sg13g2_dfrbp_1 \generated._287[4]$_SDFFE_PP0N_  (.CLK(clknet_leaf_10_clk),
    .RESET_B(net166),
    .D(_0150_),
    .Q_N(_0111_),
    .Q(\generated._14[4] ));
 sg13g2_dfrbp_1 \generated._301[0]$_SDFF_PP0_  (.CLK(clknet_leaf_9_clk),
    .RESET_B(net167),
    .D(_0151_),
    .Q_N(\generated._297[0] ),
    .Q(\generated._19[0] ));
 sg13g2_dfrbp_1 \generated._301[1]$_SDFF_PP0_  (.CLK(clknet_leaf_8_clk),
    .RESET_B(net168),
    .D(_0152_),
    .Q_N(_4559_),
    .Q(\generated._19[1] ));
 sg13g2_dfrbp_1 \generated._301[2]$_SDFF_PP0_  (.CLK(clknet_leaf_9_clk),
    .RESET_B(net169),
    .D(_0153_),
    .Q_N(_4558_),
    .Q(\generated._19[2] ));
 sg13g2_dfrbp_1 \generated._301[3]$_SDFF_PP0_  (.CLK(clknet_leaf_10_clk),
    .RESET_B(net170),
    .D(_0154_),
    .Q_N(_4557_),
    .Q(\generated._19[3] ));
 sg13g2_dfrbp_1 \generated._301[4]$_SDFF_PP0_  (.CLK(clknet_leaf_10_clk),
    .RESET_B(net171),
    .D(_0155_),
    .Q_N(_4556_),
    .Q(\generated._19[4] ));
 sg13g2_dfrbp_1 \generated._315[0]$_SDFFE_PP0P_  (.CLK(clknet_leaf_12_clk),
    .RESET_B(net172),
    .D(_0156_),
    .Q_N(_4555_),
    .Q(\generated._26[0] ));
 sg13g2_dfrbp_1 \generated._315[1]$_SDFFE_PP0P_  (.CLK(clknet_leaf_12_clk),
    .RESET_B(net173),
    .D(_0157_),
    .Q_N(_4554_),
    .Q(\generated._26[1] ));
 sg13g2_dfrbp_1 \generated._315[2]$_SDFFE_PP0P_  (.CLK(clknet_leaf_12_clk),
    .RESET_B(net174),
    .D(_0158_),
    .Q_N(_4553_),
    .Q(\generated._26[2] ));
 sg13g2_dfrbp_1 \generated._315[3]$_SDFFE_PP0P_  (.CLK(clknet_leaf_12_clk),
    .RESET_B(net175),
    .D(_0159_),
    .Q_N(_4552_),
    .Q(\generated._26[3] ));
 sg13g2_dfrbp_1 \generated._328[0]$_SDFF_PP0_  (.CLK(clknet_leaf_11_clk),
    .RESET_B(net176),
    .D(_0160_),
    .Q_N(\generated._324[0] ),
    .Q(\generated._31[0] ));
 sg13g2_dfrbp_1 \generated._328[1]$_SDFF_PP0_  (.CLK(clknet_leaf_11_clk),
    .RESET_B(net177),
    .D(_0161_),
    .Q_N(_4551_),
    .Q(\generated._31[1] ));
 sg13g2_dfrbp_1 \generated._328[2]$_SDFF_PP0_  (.CLK(clknet_leaf_10_clk),
    .RESET_B(net178),
    .D(_0162_),
    .Q_N(_4550_),
    .Q(\generated._31[2] ));
 sg13g2_dfrbp_1 \generated._328[3]$_SDFF_PP0_  (.CLK(clknet_leaf_11_clk),
    .RESET_B(net179),
    .D(_0163_),
    .Q_N(_4549_),
    .Q(\generated._31[3] ));
 sg13g2_dfrbp_1 \generated._328[4]$_SDFF_PP0_  (.CLK(clknet_leaf_11_clk),
    .RESET_B(net180),
    .D(_0164_),
    .Q_N(_4548_),
    .Q(\generated._31[4] ));
 sg13g2_dfrbp_1 \generated._328[5]$_SDFF_PP0_  (.CLK(clknet_leaf_11_clk),
    .RESET_B(net181),
    .D(_0165_),
    .Q_N(_4547_),
    .Q(\generated._31[5] ));
 sg13g2_dfrbp_1 \generated._328[6]$_SDFF_PP0_  (.CLK(clknet_leaf_11_clk),
    .RESET_B(net182),
    .D(_0166_),
    .Q_N(_4546_),
    .Q(\generated._31[6] ));
 sg13g2_dfrbp_1 \generated._342[0]$_SDFFE_PP0N_  (.CLK(clknet_leaf_13_clk),
    .RESET_B(net183),
    .D(_0167_),
    .Q_N(_0112_),
    .Q(\generated._342[0] ));
 sg13g2_dfrbp_1 \generated._342[1]$_SDFFE_PP0N_  (.CLK(clknet_leaf_13_clk),
    .RESET_B(net184),
    .D(_0168_),
    .Q_N(_0115_),
    .Q(\generated._342[1] ));
 sg13g2_dfrbp_1 \generated._342[2]$_SDFFE_PP0N_  (.CLK(clknet_leaf_13_clk),
    .RESET_B(net185),
    .D(_0169_),
    .Q_N(_0113_),
    .Q(\generated._342[2] ));
 sg13g2_dfrbp_1 \generated._342[3]$_SDFFE_PP0N_  (.CLK(clknet_leaf_13_clk),
    .RESET_B(net186),
    .D(_0170_),
    .Q_N(_0114_),
    .Q(\generated._342[3] ));
 sg13g2_dfrbp_1 \generated._342[4]$_SDFFE_PP0N_  (.CLK(clknet_leaf_14_clk),
    .RESET_B(net187),
    .D(_0171_),
    .Q_N(_4545_),
    .Q(\generated._342[4] ));
 sg13g2_dfrbp_1 \generated._342[5]$_SDFFE_PP0N_  (.CLK(clknet_leaf_14_clk),
    .RESET_B(net188),
    .D(_0172_),
    .Q_N(_4544_),
    .Q(\generated._342[5] ));
 sg13g2_dfrbp_1 \generated._353[0]$_SDFF_PP0_  (.CLK(clknet_leaf_12_clk),
    .RESET_B(net189),
    .D(_0173_),
    .Q_N(\generated._349[0] ),
    .Q(\generated._353[0] ));
 sg13g2_dfrbp_1 \generated._353[1]$_SDFF_PP0_  (.CLK(clknet_leaf_11_clk),
    .RESET_B(net190),
    .D(_0174_),
    .Q_N(_4543_),
    .Q(\generated._353[1] ));
 sg13g2_dfrbp_1 \generated._353[2]$_SDFF_PP0_  (.CLK(clknet_leaf_11_clk),
    .RESET_B(net191),
    .D(_0175_),
    .Q_N(_4542_),
    .Q(\generated._353[2] ));
 sg13g2_dfrbp_1 \generated._353[3]$_SDFF_PP0_  (.CLK(clknet_leaf_13_clk),
    .RESET_B(net192),
    .D(_0176_),
    .Q_N(_4541_),
    .Q(\generated._353[3] ));
 sg13g2_dfrbp_1 \generated._353[4]$_SDFF_PP0_  (.CLK(clknet_leaf_13_clk),
    .RESET_B(net193),
    .D(_0177_),
    .Q_N(_4540_),
    .Q(\generated._353[4] ));
 sg13g2_dfrbp_1 \generated._390[0]$_SDFF_PP0_  (.CLK(clknet_leaf_5_clk),
    .RESET_B(net194),
    .D(_0178_),
    .Q_N(_0106_),
    .Q(\generated._390[0] ));
 sg13g2_dfrbp_1 \generated._390[1]$_SDFF_PP0_  (.CLK(clknet_leaf_5_clk),
    .RESET_B(net195),
    .D(_0179_),
    .Q_N(_0063_),
    .Q(\generated._390[1] ));
 sg13g2_dfrbp_1 \generated._390[2]$_SDFF_PP1_  (.CLK(clknet_leaf_5_clk),
    .RESET_B(net196),
    .D(_0180_),
    .Q_N(_0064_),
    .Q(\generated._390[2] ));
 sg13g2_dfrbp_1 \generated._390[3]$_SDFF_PP1_  (.CLK(clknet_leaf_5_clk),
    .RESET_B(net197),
    .D(_0181_),
    .Q_N(_0062_),
    .Q(\generated._390[3] ));
 sg13g2_dfrbp_1 \generated._390[4]$_SDFF_PP1_  (.CLK(clknet_leaf_5_clk),
    .RESET_B(net198),
    .D(_0182_),
    .Q_N(_0061_),
    .Q(\generated._390[4] ));
 sg13g2_dfrbp_1 \generated._390[5]$_SDFF_PP0_  (.CLK(clknet_leaf_5_clk),
    .RESET_B(net199),
    .D(_0183_),
    .Q_N(_0060_),
    .Q(\generated._390[5] ));
 sg13g2_dfrbp_1 \generated._390[6]$_SDFF_PP0_  (.CLK(clknet_leaf_2_clk),
    .RESET_B(net200),
    .D(_0184_),
    .Q_N(_0059_),
    .Q(\generated._390[6] ));
 sg13g2_dfrbp_1 \generated._390[7]$_SDFF_PP1_  (.CLK(clknet_leaf_2_clk),
    .RESET_B(net201),
    .D(_0185_),
    .Q_N(_0070_),
    .Q(\generated._390[7] ));
 sg13g2_dfrbp_1 \generated._390[8]$_SDFF_PP0_  (.CLK(clknet_leaf_2_clk),
    .RESET_B(net202),
    .D(_0186_),
    .Q_N(_0073_),
    .Q(\generated._390[8] ));
 sg13g2_dfrbp_1 \generated._390[9]$_SDFF_PP0_  (.CLK(clknet_leaf_6_clk),
    .RESET_B(net203),
    .D(_0187_),
    .Q_N(_0076_),
    .Q(\generated._390[9] ));
 sg13g2_dfrbp_1 \generated._478[0]$_DFF_P_  (.CLK(clknet_leaf_1_clk),
    .RESET_B(net204),
    .D(\generated._477[0] ),
    .Q_N(_0089_),
    .Q(\generated._369[0] ));
 sg13g2_dfrbp_1 \generated._478[1]$_DFF_P_  (.CLK(clknet_leaf_2_clk),
    .RESET_B(net205),
    .D(\generated._477[1] ),
    .Q_N(_4595_),
    .Q(\generated._369[1] ));
 sg13g2_dfrbp_1 \generated._478[2]$_DFF_P_  (.CLK(clknet_leaf_2_clk),
    .RESET_B(net206),
    .D(\generated._477[2] ),
    .Q_N(_4596_),
    .Q(\generated._369[2] ));
 sg13g2_dfrbp_1 \generated._478[3]$_DFF_P_  (.CLK(clknet_leaf_6_clk),
    .RESET_B(net207),
    .D(\generated._477[3] ),
    .Q_N(_4597_),
    .Q(\generated._369[3] ));
 sg13g2_dfrbp_1 \generated._478[4]$_DFF_P_  (.CLK(clknet_leaf_6_clk),
    .RESET_B(net208),
    .D(\generated._477[4] ),
    .Q_N(_4598_),
    .Q(\generated._369[4] ));
 sg13g2_dfrbp_1 \generated._478[5]$_DFF_P_  (.CLK(clknet_leaf_6_clk),
    .RESET_B(net209),
    .D(\generated._477[5] ),
    .Q_N(_4599_),
    .Q(\generated._369[5] ));
 sg13g2_dfrbp_1 \generated._478[6]$_DFF_P_  (.CLK(clknet_leaf_6_clk),
    .RESET_B(net210),
    .D(\generated._477[6] ),
    .Q_N(_4600_),
    .Q(\generated._369[6] ));
 sg13g2_dfrbp_1 \generated._478[7]$_DFF_P_  (.CLK(clknet_leaf_6_clk),
    .RESET_B(net211),
    .D(\generated._477[7] ),
    .Q_N(_4601_),
    .Q(\generated._369[7] ));
 sg13g2_dfrbp_1 \generated._478[8]$_DFF_P_  (.CLK(clknet_leaf_6_clk),
    .RESET_B(net212),
    .D(\generated._477[8] ),
    .Q_N(_4602_),
    .Q(\generated._369[8] ));
 sg13g2_dfrbp_1 \generated._478[9]$_DFF_P_  (.CLK(clknet_leaf_7_clk),
    .RESET_B(net213),
    .D(\generated._477[9] ),
    .Q_N(_4603_),
    .Q(\generated._367 ));
 sg13g2_dfrbp_1 \generated._483[0]$_DFF_PN0_  (.CLK(clknet_leaf_9_clk),
    .RESET_B(net105),
    .D(\generated._482[0] ),
    .Q_N(_4604_),
    .Q(\generated._483[0] ));
 sg13g2_dfrbp_1 \generated._483[1]$_DFF_PN0_  (.CLK(clknet_leaf_9_clk),
    .RESET_B(net105),
    .D(\generated._482[1] ),
    .Q_N(_4605_),
    .Q(\generated._483[1] ));
 sg13g2_dfrbp_1 \generated._483[2]$_DFF_PN0_  (.CLK(clknet_leaf_9_clk),
    .RESET_B(net105),
    .D(\generated._482[2] ),
    .Q_N(_4606_),
    .Q(\generated._483[2] ));
 sg13g2_dfrbp_1 \generated._483[3]$_DFF_PN0_  (.CLK(clknet_leaf_7_clk),
    .RESET_B(net105),
    .D(\generated._482[3] ),
    .Q_N(_4539_),
    .Q(\generated._483[3] ));
 sg13g2_dfrbp_1 \generated._497[0]$_SDFF_PP0_  (.CLK(clknet_leaf_12_clk),
    .RESET_B(net214),
    .D(_0188_),
    .Q_N(_0107_),
    .Q(\generated._497[0] ));
 sg13g2_dfrbp_1 \generated._497[1]$_SDFF_PP0_  (.CLK(clknet_leaf_8_clk),
    .RESET_B(net215),
    .D(_0189_),
    .Q_N(_0108_),
    .Q(\generated._377[0] ));
 sg13g2_dfrbp_1 \generated._497[2]$_SDFF_PP0_  (.CLK(clknet_leaf_8_clk),
    .RESET_B(net216),
    .D(_0190_),
    .Q_N(_0109_),
    .Q(\generated._377[1] ));
 sg13g2_dfrbp_1 \generated._497[3]$_SDFF_PP0_  (.CLK(clknet_leaf_12_clk),
    .RESET_B(net217),
    .D(_0191_),
    .Q_N(_0110_),
    .Q(\generated._377[2] ));
 sg13g2_dfrbp_1 \generated._497[4]$_SDFF_PP0_  (.CLK(clknet_leaf_12_clk),
    .RESET_B(net218),
    .D(_0192_),
    .Q_N(_0090_),
    .Q(\generated._377[3] ));
 sg13g2_dfrbp_1 \generated._497[5]$_SDFF_PP0_  (.CLK(clknet_leaf_9_clk),
    .RESET_B(net219),
    .D(_0193_),
    .Q_N(_0091_),
    .Q(\generated._377[4] ));
 sg13g2_dfrbp_1 \generated._497[6]$_SDFF_PP0_  (.CLK(clknet_leaf_9_clk),
    .RESET_B(net220),
    .D(_0194_),
    .Q_N(_0092_),
    .Q(\generated._377[5] ));
 sg13g2_dfrbp_1 \generated._497[7]$_SDFF_PP0_  (.CLK(clknet_leaf_9_clk),
    .RESET_B(net221),
    .D(_0195_),
    .Q_N(_0093_),
    .Q(\generated._377[6] ));
 sg13g2_dfrbp_1 \generated._497[8]$_SDFF_PP0_  (.CLK(clknet_leaf_8_clk),
    .RESET_B(net222),
    .D(_0196_),
    .Q_N(_0094_),
    .Q(\generated._377[7] ));
 sg13g2_dfrbp_1 \generated._497[9]$_SDFF_PP0_  (.CLK(clknet_leaf_7_clk),
    .RESET_B(net223),
    .D(_0197_),
    .Q_N(_0095_),
    .Q(\generated._376 ));
 sg13g2_dfrbp_1 \generated._558[0]$_DFF_P_  (.CLK(clknet_leaf_20_clk),
    .RESET_B(net224),
    .D(\generated._557[0] ),
    .Q_N(_0065_),
    .Q(\generated._558[0] ));
 sg13g2_dfrbp_1 \generated._558[1]$_DFF_P_  (.CLK(clknet_leaf_21_clk),
    .RESET_B(net225),
    .D(\generated._557[1] ),
    .Q_N(_0071_),
    .Q(\generated._558[1] ));
 sg13g2_dfrbp_1 \generated._558[2]$_DFF_P_  (.CLK(clknet_leaf_20_clk),
    .RESET_B(net226),
    .D(\generated._557[2] ),
    .Q_N(_0074_),
    .Q(\generated._558[2] ));
 sg13g2_dfrbp_1 \generated._558[3]$_DFF_P_  (.CLK(clknet_leaf_22_clk),
    .RESET_B(net227),
    .D(\generated._557[3] ),
    .Q_N(_0077_),
    .Q(\generated._558[3] ));
 sg13g2_dfrbp_1 \generated._558[4]$_DFF_P_  (.CLK(clknet_leaf_22_clk),
    .RESET_B(net228),
    .D(\generated._557[4] ),
    .Q_N(_0079_),
    .Q(\generated._558[4] ));
 sg13g2_dfrbp_1 \generated._558[5]$_DFF_P_  (.CLK(clknet_leaf_21_clk),
    .RESET_B(net229),
    .D(\generated._557[5] ),
    .Q_N(_0081_),
    .Q(\generated._558[5] ));
 sg13g2_dfrbp_1 \generated._558[6]$_DFF_P_  (.CLK(clknet_leaf_21_clk),
    .RESET_B(net230),
    .D(\generated._557[6] ),
    .Q_N(_0083_),
    .Q(\generated._558[6] ));
 sg13g2_dfrbp_1 \generated._558[7]$_DFF_P_  (.CLK(clknet_leaf_22_clk),
    .RESET_B(net231),
    .D(\generated._557[7] ),
    .Q_N(_0085_),
    .Q(\generated._558[7] ));
 sg13g2_dfrbp_1 \generated._558[8]$_DFF_P_  (.CLK(clknet_leaf_22_clk),
    .RESET_B(net232),
    .D(\generated._557[8] ),
    .Q_N(_0086_),
    .Q(\generated._558[8] ));
 sg13g2_dfrbp_1 \generated._558[9]$_DFF_P_  (.CLK(clknet_leaf_22_clk),
    .RESET_B(net233),
    .D(\generated._557[9] ),
    .Q_N(_0087_),
    .Q(\generated._558[9] ));
 sg13g2_dfrbp_1 \generated._692[0]$_DFF_P_  (.CLK(clknet_leaf_25_clk),
    .RESET_B(net234),
    .D(\generated._691[0] ),
    .Q_N(_0049_),
    .Q(\generated._501[0] ));
 sg13g2_dfrbp_1 \generated._692[1]$_DFF_P_  (.CLK(clknet_leaf_25_clk),
    .RESET_B(net235),
    .D(\generated._691[1] ),
    .Q_N(_4607_),
    .Q(\generated._501[1] ));
 sg13g2_dfrbp_1 \generated._692[2]$_DFF_P_  (.CLK(clknet_leaf_25_clk),
    .RESET_B(net236),
    .D(\generated._691[2] ),
    .Q_N(_4608_),
    .Q(\generated._501[2] ));
 sg13g2_dfrbp_1 \generated._692[3]$_DFF_P_  (.CLK(clknet_leaf_25_clk),
    .RESET_B(net237),
    .D(\generated._691[3] ),
    .Q_N(_4609_),
    .Q(\generated._501[3] ));
 sg13g2_dfrbp_1 \generated._692[4]$_DFF_P_  (.CLK(clknet_leaf_25_clk),
    .RESET_B(net238),
    .D(\generated._691[4] ),
    .Q_N(_4610_),
    .Q(\generated._501[4] ));
 sg13g2_dfrbp_1 \generated._692[5]$_DFF_P_  (.CLK(clknet_leaf_25_clk),
    .RESET_B(net239),
    .D(\generated._691[5] ),
    .Q_N(_4611_),
    .Q(\generated._501[5] ));
 sg13g2_dfrbp_1 \generated._692[6]$_DFF_P_  (.CLK(clknet_leaf_24_clk),
    .RESET_B(net240),
    .D(\generated._691[6] ),
    .Q_N(_4612_),
    .Q(\generated._501[6] ));
 sg13g2_dfrbp_1 \generated._692[7]$_DFF_P_  (.CLK(clknet_leaf_24_clk),
    .RESET_B(net241),
    .D(\generated._691[7] ),
    .Q_N(_4613_),
    .Q(\generated._501[7] ));
 sg13g2_dfrbp_1 \generated._692[8]$_DFF_P_  (.CLK(clknet_leaf_24_clk),
    .RESET_B(net242),
    .D(\generated._691[8] ),
    .Q_N(_4614_),
    .Q(\generated._501[8] ));
 sg13g2_dfrbp_1 \generated._692[9]$_DFF_P_  (.CLK(clknet_leaf_24_clk),
    .RESET_B(net243),
    .D(\generated._691[9] ),
    .Q_N(_4615_),
    .Q(\generated._499 ));
 sg13g2_dfrbp_1 \generated._696[0]$_DFF_PN0_  (.CLK(clknet_leaf_30_clk),
    .RESET_B(net96),
    .D(\generated._60[0] ),
    .Q_N(_4616_),
    .Q(\generated._61[0] ));
 sg13g2_dfrbp_1 \generated._696[1]$_DFF_PN0_  (.CLK(clknet_leaf_30_clk),
    .RESET_B(net96),
    .D(\generated._60[1] ),
    .Q_N(_4617_),
    .Q(\generated._61[1] ));
 sg13g2_dfrbp_1 \generated._696[2]$_DFF_PN0_  (.CLK(clknet_leaf_30_clk),
    .RESET_B(net97),
    .D(\generated._60[2] ),
    .Q_N(_4618_),
    .Q(\generated._61[2] ));
 sg13g2_dfrbp_1 \generated._696[3]$_DFF_PN0_  (.CLK(clknet_leaf_4_clk),
    .RESET_B(net97),
    .D(\generated._60[3] ),
    .Q_N(_4538_),
    .Q(\generated._61[3] ));
 sg13g2_dfrbp_1 \generated._710[0]$_SDFF_PP0_  (.CLK(clknet_leaf_23_clk),
    .RESET_B(net244),
    .D(_0198_),
    .Q_N(_0067_),
    .Q(\generated._62[0] ));
 sg13g2_dfrbp_1 \generated._710[1]$_SDFF_PP0_  (.CLK(clknet_leaf_23_clk),
    .RESET_B(net245),
    .D(_0199_),
    .Q_N(_0066_),
    .Q(\generated._508[0] ));
 sg13g2_dfrbp_1 \generated._710[2]$_SDFF_PP0_  (.CLK(clknet_leaf_23_clk),
    .RESET_B(net246),
    .D(_0200_),
    .Q_N(_0068_),
    .Q(\generated._508[1] ));
 sg13g2_dfrbp_1 \generated._710[3]$_SDFF_PP0_  (.CLK(clknet_leaf_23_clk),
    .RESET_B(net247),
    .D(_0201_),
    .Q_N(_0069_),
    .Q(\generated._508[2] ));
 sg13g2_dfrbp_1 \generated._710[4]$_SDFF_PP0_  (.CLK(clknet_leaf_23_clk),
    .RESET_B(net248),
    .D(_0202_),
    .Q_N(_0072_),
    .Q(\generated._508[3] ));
 sg13g2_dfrbp_1 \generated._710[5]$_SDFF_PP0_  (.CLK(clknet_leaf_23_clk),
    .RESET_B(net249),
    .D(_0203_),
    .Q_N(_0075_),
    .Q(\generated._508[4] ));
 sg13g2_dfrbp_1 \generated._710[6]$_SDFF_PP0_  (.CLK(clknet_leaf_23_clk),
    .RESET_B(net250),
    .D(_0204_),
    .Q_N(_0078_),
    .Q(\generated._508[5] ));
 sg13g2_dfrbp_1 \generated._710[7]$_SDFF_PP0_  (.CLK(clknet_leaf_23_clk),
    .RESET_B(net251),
    .D(_0205_),
    .Q_N(_0080_),
    .Q(\generated._508[6] ));
 sg13g2_dfrbp_1 \generated._710[8]$_SDFF_PP0_  (.CLK(clknet_leaf_24_clk),
    .RESET_B(net252),
    .D(_0206_),
    .Q_N(_0082_),
    .Q(\generated._508[7] ));
 sg13g2_dfrbp_1 \generated._710[9]$_SDFF_PP0_  (.CLK(clknet_leaf_24_clk),
    .RESET_B(net253),
    .D(_0207_),
    .Q_N(_0084_),
    .Q(\generated._507 ));
 sg13g2_dfrbp_1 \generated._830[0]$_DFF_PN0_  (.CLK(clknet_3_7__leaf_clk),
    .RESET_B(net102),
    .D(\generated._825[2] ),
    .Q_N(_4619_),
    .Q(\generated._1083[0] ));
 sg13g2_dfrbp_1 \generated._830[1]$_DFF_PN0_  (.CLK(clknet_leaf_17_clk),
    .RESET_B(net103),
    .D(\generated._825[3] ),
    .Q_N(_0119_),
    .Q(\generated._161[4] ));
 sg13g2_dfrbp_1 \generated._830[2]$_DFF_PN0_  (.CLK(clknet_leaf_19_clk),
    .RESET_B(net103),
    .D(\generated._825[4] ),
    .Q_N(_4620_),
    .Q(\generated._63[2] ));
 sg13g2_dfrbp_1 \generated._830[3]$_DFF_PN0_  (.CLK(clknet_leaf_19_clk),
    .RESET_B(net103),
    .D(\generated._825[5] ),
    .Q_N(_4621_),
    .Q(\generated._63[3] ));
 sg13g2_dfrbp_1 \generated._830[4]$_DFF_PN0_  (.CLK(clknet_leaf_19_clk),
    .RESET_B(net103),
    .D(\generated._825[6] ),
    .Q_N(_4622_),
    .Q(\generated._63[4] ));
 sg13g2_dfrbp_1 \generated._830[5]$_DFF_PN0_  (.CLK(clknet_leaf_19_clk),
    .RESET_B(net103),
    .D(\generated._825[7] ),
    .Q_N(_4623_),
    .Q(\generated._63[5] ));
 sg13g2_dfrbp_1 \generated._830[6]$_DFF_PN0_  (.CLK(clknet_leaf_19_clk),
    .RESET_B(net103),
    .D(\generated._825[8] ),
    .Q_N(_4537_),
    .Q(\generated._63[6] ));
 sg13g2_dfrbp_1 \generated._886[0]$_SDFF_PP0_  (.CLK(clknet_leaf_33_clk),
    .RESET_B(net254),
    .D(_0208_),
    .Q_N(_0102_),
    .Q(\generated._421[1] ));
 sg13g2_dfrbp_1 \generated._886[1]$_SDFF_PP0_  (.CLK(clknet_leaf_27_clk),
    .RESET_B(net255),
    .D(_0209_),
    .Q_N(_0103_),
    .Q(\generated._64[1] ));
 sg13g2_dfrbp_1 \generated._886[2]$_SDFF_PP0_  (.CLK(clknet_leaf_33_clk),
    .RESET_B(net256),
    .D(_0210_),
    .Q_N(_0104_),
    .Q(\generated._64[2] ));
 sg13g2_dfrbp_1 \generated._886[3]$_DFF_P_  (.CLK(clknet_leaf_33_clk),
    .RESET_B(net257),
    .D(\generated._885[3] ),
    .Q_N(_0105_),
    .Q(\generated._64[3] ));
 sg13g2_dfrbp_1 \generated._886[4]$_DFF_P_  (.CLK(clknet_leaf_33_clk),
    .RESET_B(net258),
    .D(\generated._885[4] ),
    .Q_N(_0036_),
    .Q(\generated._64[4] ));
 sg13g2_dfrbp_1 \generated._886[5]$_DFF_P_  (.CLK(clknet_leaf_32_clk),
    .RESET_B(net259),
    .D(\generated._885[5] ),
    .Q_N(_0037_),
    .Q(\generated._64[5] ));
 sg13g2_dfrbp_1 \generated._886[6]$_DFF_P_  (.CLK(clknet_leaf_32_clk),
    .RESET_B(net260),
    .D(\generated._885[6] ),
    .Q_N(_0038_),
    .Q(\generated._64[6] ));
 sg13g2_dfrbp_1 \generated._886[7]$_DFF_P_  (.CLK(clknet_leaf_30_clk),
    .RESET_B(net261),
    .D(\generated._885[7] ),
    .Q_N(_0043_),
    .Q(\generated._64[7] ));
 sg13g2_dfrbp_1 \generated._886[8]$_DFF_P_  (.CLK(clknet_leaf_30_clk),
    .RESET_B(net262),
    .D(\generated._885[8] ),
    .Q_N(_0025_),
    .Q(\generated._64[8] ));
 sg13g2_dfrbp_1 \generated._886[9]$_DFF_P_  (.CLK(clknet_leaf_31_clk),
    .RESET_B(net263),
    .D(\generated._885[9] ),
    .Q_N(_0032_),
    .Q(\generated._64[9] ));
 sg13g2_dfrbp_1 \generated._935[0]$_SDFF_PP0_  (.CLK(clknet_leaf_26_clk),
    .RESET_B(net264),
    .D(_0211_),
    .Q_N(_0101_),
    .Q(\generated._67[0] ));
 sg13g2_dfrbp_1 \generated._935[1]$_SDFF_PP0_  (.CLK(clknet_leaf_26_clk),
    .RESET_B(net265),
    .D(_0212_),
    .Q_N(_0041_),
    .Q(\generated._67[1] ));
 sg13g2_dfrbp_1 \generated._935[2]$_SDFF_PP0_  (.CLK(clknet_leaf_27_clk),
    .RESET_B(net266),
    .D(_0213_),
    .Q_N(_0040_),
    .Q(\generated._67[2] ));
 sg13g2_dfrbp_1 \generated._935[3]$_DFF_P_  (.CLK(clknet_leaf_27_clk),
    .RESET_B(net267),
    .D(\generated._934[3] ),
    .Q_N(_0035_),
    .Q(\generated._67[3] ));
 sg13g2_dfrbp_1 \generated._935[4]$_DFF_P_  (.CLK(clknet_leaf_28_clk),
    .RESET_B(net268),
    .D(\generated._934[4] ),
    .Q_N(_0042_),
    .Q(\generated._67[4] ));
 sg13g2_dfrbp_1 \generated._935[5]$_DFF_P_  (.CLK(clknet_leaf_28_clk),
    .RESET_B(net269),
    .D(\generated._934[5] ),
    .Q_N(_0044_),
    .Q(\generated._67[5] ));
 sg13g2_dfrbp_1 \generated._935[6]$_DFF_P_  (.CLK(clknet_leaf_29_clk),
    .RESET_B(net270),
    .D(\generated._934[6] ),
    .Q_N(_0045_),
    .Q(\generated._67[6] ));
 sg13g2_dfrbp_1 \generated._935[7]$_DFF_P_  (.CLK(clknet_leaf_28_clk),
    .RESET_B(net271),
    .D(\generated._934[7] ),
    .Q_N(_0046_),
    .Q(\generated._67[7] ));
 sg13g2_dfrbp_1 \generated._935[8]$_DFF_P_  (.CLK(clknet_leaf_30_clk),
    .RESET_B(net272),
    .D(\generated._934[8] ),
    .Q_N(_0047_),
    .Q(\generated._67[8] ));
 sg13g2_dfrbp_1 \generated._935[9]$_DFF_P_  (.CLK(clknet_leaf_30_clk),
    .RESET_B(net273),
    .D(\generated._934[9] ),
    .Q_N(_0039_),
    .Q(\generated._67[9] ));
 sg13g2_dfrbp_1 \generated._939[0]$_DFF_PN0_  (.CLK(clknet_leaf_31_clk),
    .RESET_B(net96),
    .D(\generated._68[0] ),
    .Q_N(_4624_),
    .Q(\generated._69[0] ));
 sg13g2_dfrbp_1 \generated._939[1]$_DFF_PN0_  (.CLK(clknet_leaf_31_clk),
    .RESET_B(net96),
    .D(\generated._68[1] ),
    .Q_N(_4625_),
    .Q(\generated._69[1] ));
 sg13g2_dfrbp_1 \generated._939[2]$_DFF_PN0_  (.CLK(clknet_leaf_31_clk),
    .RESET_B(net96),
    .D(\generated._68[2] ),
    .Q_N(_4626_),
    .Q(\generated._69[2] ));
 sg13g2_dfrbp_1 \generated._939[3]$_DFF_PN0_  (.CLK(clknet_leaf_31_clk),
    .RESET_B(net96),
    .D(\generated._68[3] ),
    .Q_N(_4536_),
    .Q(\generated._69[3] ));
 sg13g2_dfrbp_1 \generated._945[0]$_SDFF_PP0_  (.CLK(clknet_leaf_26_clk),
    .RESET_B(net274),
    .D(_0214_),
    .Q_N(_0048_),
    .Q(\generated._430[10] ));
 sg13g2_dfrbp_1 \generated._945[1]$_SDFF_PP0_  (.CLK(clknet_leaf_26_clk),
    .RESET_B(net275),
    .D(_0215_),
    .Q_N(_0056_),
    .Q(\generated._430[11] ));
 sg13g2_dfrbp_1 \generated._945[2]$_SDFF_PP0_  (.CLK(clknet_leaf_26_clk),
    .RESET_B(net276),
    .D(_0216_),
    .Q_N(_0055_),
    .Q(\generated._430[12] ));
 sg13g2_dfrbp_1 \generated._945[3]$_SDFF_PP0_  (.CLK(clknet_leaf_26_clk),
    .RESET_B(net277),
    .D(_0217_),
    .Q_N(_0057_),
    .Q(\generated._430[13] ));
 sg13g2_dfrbp_1 \generated._945[4]$_SDFF_PP0_  (.CLK(clknet_leaf_26_clk),
    .RESET_B(net278),
    .D(_0218_),
    .Q_N(_0054_),
    .Q(\generated._430[14] ));
 sg13g2_dfrbp_1 \generated._945[5]$_SDFF_PP0_  (.CLK(clknet_leaf_28_clk),
    .RESET_B(net279),
    .D(_0219_),
    .Q_N(_0053_),
    .Q(\generated._430[15] ));
 sg13g2_dfrbp_1 \generated._945[6]$_SDFF_PP0_  (.CLK(clknet_leaf_28_clk),
    .RESET_B(net280),
    .D(_0220_),
    .Q_N(_0052_),
    .Q(\generated._430[16] ));
 sg13g2_dfrbp_1 \generated._945[7]$_SDFF_PP0_  (.CLK(clknet_leaf_28_clk),
    .RESET_B(net281),
    .D(_0221_),
    .Q_N(_0058_),
    .Q(\generated._430[17] ));
 sg13g2_dfrbp_1 \generated._945[8]$_SDFF_PP0_  (.CLK(clknet_leaf_28_clk),
    .RESET_B(net282),
    .D(_0222_),
    .Q_N(_0051_),
    .Q(\generated._430[18] ));
 sg13g2_dfrbp_1 \generated._945[9]$_SDFF_PP0_  (.CLK(clknet_leaf_28_clk),
    .RESET_B(net283),
    .D(_0223_),
    .Q_N(_0050_),
    .Q(\generated._430[19] ));
 sg13g2_dfrbp_1 \generated._946[0]$_DFF_PN0_  (.CLK(clknet_leaf_15_clk),
    .RESET_B(net100),
    .D(\generated._1115[0] ),
    .Q_N(_4627_),
    .Q(\generated._568[0] ));
 sg13g2_dfrbp_1 \generated._946[1]$_DFF_PN0_  (.CLK(clknet_leaf_15_clk),
    .RESET_B(net100),
    .D(\generated._1115[1] ),
    .Q_N(_4628_),
    .Q(\generated._568[1] ));
 sg13g2_dfrbp_1 \generated._946[2]$_DFF_PN0_  (.CLK(clknet_leaf_15_clk),
    .RESET_B(net100),
    .D(\generated._1115[2] ),
    .Q_N(_4629_),
    .Q(\generated._568[2] ));
 sg13g2_dfrbp_1 \generated._946[3]$_DFF_PN0_  (.CLK(clknet_leaf_30_clk),
    .RESET_B(net98),
    .D(\generated._1115[3] ),
    .Q_N(_0120_),
    .Q(\generated._568[3] ));
 sg13g2_dfrbp_1 \generated._946[4]$_DFF_PN0_  (.CLK(clknet_leaf_29_clk),
    .RESET_B(net97),
    .D(\generated._1115[4] ),
    .Q_N(_4630_),
    .Q(\generated._568[4] ));
 sg13g2_dfrbp_1 \generated._946[5]$_DFF_PN0_  (.CLK(clknet_leaf_29_clk),
    .RESET_B(net98),
    .D(\generated._1115[5] ),
    .Q_N(_0121_),
    .Q(\generated._568[5] ));
 sg13g2_dfrbp_1 \generated._946[6]$_DFF_PN0_  (.CLK(clknet_leaf_4_clk),
    .RESET_B(net98),
    .D(\generated._1115[6] ),
    .Q_N(_4631_),
    .Q(\generated._568[6] ));
 sg13g2_dfrbp_1 \generated._946[7]$_DFF_PN0_  (.CLK(clknet_leaf_21_clk),
    .RESET_B(net101),
    .D(\generated._1115[7] ),
    .Q_N(_0117_),
    .Q(\generated._568[7] ));
 sg13g2_dfrbp_1 \generated._946[8]$_DFF_PN0_  (.CLK(clknet_leaf_20_clk),
    .RESET_B(net101),
    .D(\generated._1115[8] ),
    .Q_N(_4632_),
    .Q(\generated._568[8] ));
 sg13g2_dfrbp_1 \generated._946[9]$_DFF_PN0_  (.CLK(clknet_leaf_21_clk),
    .RESET_B(net101),
    .D(\generated._1115[9] ),
    .Q_N(_0122_),
    .Q(\generated._568[9] ));
 sg13g2_dfrbp_1 \generated._949[0]$_DFFE_PN0N_  (.CLK(clknet_leaf_16_clk),
    .RESET_B(net105),
    .D(_0224_),
    .Q_N(_4535_),
    .Q(\generated._610[0] ));
 sg13g2_dfrbp_1 \generated._949[1]$_DFFE_PN0N_  (.CLK(clknet_leaf_16_clk),
    .RESET_B(net104),
    .D(_0225_),
    .Q_N(_4534_),
    .Q(\generated._610[1] ));
 sg13g2_dfrbp_1 \generated._949[2]$_DFFE_PN0N_  (.CLK(clknet_leaf_15_clk),
    .RESET_B(net105),
    .D(_0226_),
    .Q_N(_4533_),
    .Q(\generated._610[2] ));
 sg13g2_dfrbp_1 \generated._949[3]$_DFFE_PN0N_  (.CLK(clknet_leaf_15_clk),
    .RESET_B(net101),
    .D(_0227_),
    .Q_N(_0116_),
    .Q(\generated._610[3] ));
 sg13g2_dfrbp_1 \generated._949[4]$_DFFE_PN0N_  (.CLK(clknet_leaf_15_clk),
    .RESET_B(net100),
    .D(_0228_),
    .Q_N(_4532_),
    .Q(\generated._610[4] ));
 sg13g2_dfrbp_1 \generated._949[5]$_DFFE_PN0N_  (.CLK(clknet_leaf_16_clk),
    .RESET_B(net104),
    .D(_0229_),
    .Q_N(_0123_),
    .Q(\generated._610[5] ));
 sg13g2_dfrbp_1 \generated._949[6]$_DFFE_PN0N_  (.CLK(clknet_leaf_16_clk),
    .RESET_B(net104),
    .D(_0230_),
    .Q_N(_0118_),
    .Q(\generated._217[0] ));
 sg13g2_dfrbp_1 \generated._949[7]$_DFFE_PN0N_  (.CLK(clknet_leaf_15_clk),
    .RESET_B(net101),
    .D(_0231_),
    .Q_N(_0124_),
    .Q(\generated._217[1] ));
 sg13g2_dfrbp_1 \generated._949[8]$_DFFE_PN0N_  (.CLK(clknet_leaf_15_clk),
    .RESET_B(net101),
    .D(_0232_),
    .Q_N(_0125_),
    .Q(\generated._217[2] ));
 sg13g2_dfrbp_1 \generated._949[9]$_DFFE_PN0N_  (.CLK(clknet_leaf_16_clk),
    .RESET_B(net104),
    .D(_0233_),
    .Q_N(_0126_),
    .Q(\generated._217[3] ));
 sg13g2_dfrbp_1 \generated._956[0]$_DFFE_PN0P_  (.CLK(clknet_leaf_4_clk),
    .RESET_B(net100),
    .D(_0234_),
    .Q_N(\generated._75[0] ),
    .Q(\generated._1037[0] ));
 sg13g2_dfrbp_1 \generated._956[1]$_DFFE_PN0P_  (.CLK(clknet_leaf_4_clk),
    .RESET_B(net97),
    .D(_0235_),
    .Q_N(_4531_),
    .Q(\generated._402[1] ));
 sg13g2_dfrbp_1 \generated._956[2]$_DFFE_PN0P_  (.CLK(clknet_leaf_4_clk),
    .RESET_B(net97),
    .D(_0236_),
    .Q_N(_4530_),
    .Q(\generated._402[2] ));
 sg13g2_dfrbp_1 \generated._956[3]$_DFFE_PN0P_  (.CLK(clknet_leaf_4_clk),
    .RESET_B(net97),
    .D(_0237_),
    .Q_N(_4529_),
    .Q(\generated._402[3] ));
 sg13g2_dfrbp_1 \generated._956[4]$_DFFE_PN0P_  (.CLK(clknet_leaf_3_clk),
    .RESET_B(net99),
    .D(_0238_),
    .Q_N(_0033_),
    .Q(\generated._402[4] ));
 sg13g2_dfrbp_1 \generated._956[5]$_DFFE_PN0P_  (.CLK(clknet_leaf_2_clk),
    .RESET_B(net99),
    .D(_0239_),
    .Q_N(_4528_),
    .Q(\generated._402[5] ));
 sg13g2_dfrbp_1 \generated._956[6]$_DFFE_PN0P_  (.CLK(clknet_leaf_3_clk),
    .RESET_B(net99),
    .D(_0240_),
    .Q_N(_4527_),
    .Q(\generated._402[6] ));
 sg13g2_dfrbp_1 \generated._956[7]$_DFFE_PN0P_  (.CLK(clknet_leaf_3_clk),
    .RESET_B(net100),
    .D(_0241_),
    .Q_N(_0034_),
    .Q(\generated._402[7] ));
 sg13g2_dfrbp_1 \generated.iter_sel[0]$_SDFF_PP0_  (.CLK(clknet_leaf_6_clk),
    .RESET_B(net284),
    .D(_0242_),
    .Q_N(\generated._391[0] ),
    .Q(\generated._375 ));
 sg13g2_dfrbp_1 \generated.iter_sel[1]$_SDFF_PP0_  (.CLK(clknet_leaf_7_clk),
    .RESET_B(net285),
    .D(_0243_),
    .Q_N(_4526_),
    .Q(\generated._374 ));
 sg13g2_dfrbp_1 \generated.iter_sel_0[0]$_SDFF_PP0_  (.CLK(clknet_leaf_24_clk),
    .RESET_B(net286),
    .D(_0244_),
    .Q_N(\generated._559[0] ),
    .Q(\generated._506 ));
 sg13g2_dfrbp_1 \generated.iter_sel_0[1]$_SDFF_PP0_  (.CLK(clknet_leaf_24_clk),
    .RESET_B(net287),
    .D(_0245_),
    .Q_N(_4525_),
    .Q(\generated._505 ));
 sg13g2_dfrbp_1 \generated.iter_sel_1[0]$_SDFF_PP0_  (.CLK(clknet_leaf_33_clk),
    .RESET_B(net288),
    .D(_0246_),
    .Q_N(\generated._887[0] ),
    .Q(\generated._840 ));
 sg13g2_dfrbp_1 \generated.iter_sel_1[1]$_SDFF_PP0_  (.CLK(clknet_leaf_26_clk),
    .RESET_B(net289),
    .D(_0247_),
    .Q_N(_4524_),
    .Q(\generated._839 ));
 sg13g2_dfrbp_1 \generated.iter_sel_2[0]$_SDFF_PP0_  (.CLK(clknet_leaf_0_clk),
    .RESET_B(net290),
    .D(_0248_),
    .Q_N(\generated._1021[0] ),
    .Q(\generated._966 ));
 sg13g2_dfrbp_1 \generated.iter_sel_2[1]$_SDFF_PP0_  (.CLK(clknet_leaf_0_clk),
    .RESET_B(net291),
    .D(_0249_),
    .Q_N(_4523_),
    .Q(\generated._965 ));
 sg13g2_buf_1 input1 (.A(rst_n),
    .X(net1));
 sg13g2_buf_1 output2 (.A(net2),
    .X(uo_out[0]));
 sg13g2_buf_1 output3 (.A(net3),
    .X(uo_out[1]));
 sg13g2_buf_1 output4 (.A(net4),
    .X(uo_out[2]));
 sg13g2_buf_1 output5 (.A(net5),
    .X(uo_out[3]));
 sg13g2_buf_1 output6 (.A(net6),
    .X(uo_out[4]));
 sg13g2_buf_1 output7 (.A(net7),
    .X(uo_out[5]));
 sg13g2_buf_1 output8 (.A(net8),
    .X(uo_out[6]));
 sg13g2_buf_1 output9 (.A(net9),
    .X(uo_out[7]));
 sg13g2_buf_2 fanout10 (.A(_2073_),
    .X(net10));
 sg13g2_buf_2 fanout11 (.A(_2059_),
    .X(net11));
 sg13g2_buf_2 fanout12 (.A(_2080_),
    .X(net12));
 sg13g2_buf_2 fanout13 (.A(_2240_),
    .X(net13));
 sg13g2_buf_2 fanout14 (.A(_2304_),
    .X(net14));
 sg13g2_buf_2 fanout15 (.A(_3216_),
    .X(net15));
 sg13g2_buf_2 fanout16 (.A(_3958_),
    .X(net16));
 sg13g2_buf_2 fanout17 (.A(_3252_),
    .X(net17));
 sg13g2_buf_2 fanout18 (.A(_3954_),
    .X(net18));
 sg13g2_buf_2 fanout19 (.A(_2278_),
    .X(net19));
 sg13g2_buf_2 fanout20 (.A(_2006_),
    .X(net20));
 sg13g2_buf_2 fanout21 (.A(_3956_),
    .X(net21));
 sg13g2_buf_2 fanout22 (.A(_2782_),
    .X(net22));
 sg13g2_buf_2 fanout23 (.A(_2768_),
    .X(net23));
 sg13g2_buf_2 fanout24 (.A(_2078_),
    .X(net24));
 sg13g2_buf_2 fanout25 (.A(_2010_),
    .X(net25));
 sg13g2_buf_2 fanout26 (.A(_1980_),
    .X(net26));
 sg13g2_buf_2 fanout27 (.A(_2069_),
    .X(net27));
 sg13g2_buf_2 fanout28 (.A(_1968_),
    .X(net28));
 sg13g2_buf_2 fanout29 (.A(_4179_),
    .X(net29));
 sg13g2_buf_2 fanout30 (.A(_3278_),
    .X(net30));
 sg13g2_buf_2 fanout31 (.A(_2233_),
    .X(net31));
 sg13g2_buf_2 fanout32 (.A(_0889_),
    .X(net32));
 sg13g2_buf_2 fanout33 (.A(_0437_),
    .X(net33));
 sg13g2_buf_2 fanout34 (.A(_0319_),
    .X(net34));
 sg13g2_buf_2 fanout35 (.A(_4444_),
    .X(net35));
 sg13g2_buf_2 fanout36 (.A(_4327_),
    .X(net36));
 sg13g2_buf_2 fanout37 (.A(_2247_),
    .X(net37));
 sg13g2_buf_2 fanout38 (.A(_1678_),
    .X(net38));
 sg13g2_buf_2 fanout39 (.A(_1306_),
    .X(net39));
 sg13g2_buf_2 fanout40 (.A(_0792_),
    .X(net40));
 sg13g2_buf_2 fanout41 (.A(_0759_),
    .X(net41));
 sg13g2_buf_2 fanout42 (.A(_0692_),
    .X(net42));
 sg13g2_buf_2 fanout43 (.A(_0585_),
    .X(net43));
 sg13g2_buf_2 fanout44 (.A(_0306_),
    .X(net44));
 sg13g2_buf_2 fanout45 (.A(_4492_),
    .X(net45));
 sg13g2_buf_2 fanout46 (.A(_4369_),
    .X(net46));
 sg13g2_buf_2 fanout47 (.A(_4355_),
    .X(net47));
 sg13g2_buf_2 fanout48 (.A(_4326_),
    .X(net48));
 sg13g2_buf_2 fanout49 (.A(_3976_),
    .X(net49));
 sg13g2_buf_2 fanout50 (.A(_3961_),
    .X(net50));
 sg13g2_buf_2 fanout51 (.A(_0928_),
    .X(net51));
 sg13g2_buf_2 fanout52 (.A(_0909_),
    .X(net52));
 sg13g2_buf_2 fanout53 (.A(_0775_),
    .X(net53));
 sg13g2_buf_2 fanout54 (.A(_0756_),
    .X(net54));
 sg13g2_buf_2 fanout55 (.A(_0665_),
    .X(net55));
 sg13g2_buf_2 fanout56 (.A(_0627_),
    .X(net56));
 sg13g2_buf_2 fanout57 (.A(_0618_),
    .X(net57));
 sg13g2_buf_2 fanout58 (.A(_0609_),
    .X(net58));
 sg13g2_buf_2 fanout59 (.A(_0582_),
    .X(net59));
 sg13g2_buf_2 fanout60 (.A(_0373_),
    .X(net60));
 sg13g2_buf_2 fanout61 (.A(_0322_),
    .X(net61));
 sg13g2_buf_2 fanout62 (.A(_0305_),
    .X(net62));
 sg13g2_buf_2 fanout63 (.A(_4491_),
    .X(net63));
 sg13g2_buf_2 fanout64 (.A(_4426_),
    .X(net64));
 sg13g2_buf_2 fanout65 (.A(_4377_),
    .X(net65));
 sg13g2_buf_2 fanout66 (.A(_3975_),
    .X(net66));
 sg13g2_buf_2 fanout67 (.A(_3962_),
    .X(net67));
 sg13g2_buf_2 fanout68 (.A(_1493_),
    .X(net68));
 sg13g2_buf_2 fanout69 (.A(_0786_),
    .X(net69));
 sg13g2_buf_2 fanout70 (.A(_0664_),
    .X(net70));
 sg13g2_buf_2 fanout71 (.A(_0610_),
    .X(net71));
 sg13g2_buf_2 fanout72 (.A(_0581_),
    .X(net72));
 sg13g2_buf_2 fanout73 (.A(_0379_),
    .X(net73));
 sg13g2_buf_2 fanout74 (.A(_0372_),
    .X(net74));
 sg13g2_buf_2 fanout75 (.A(_0323_),
    .X(net75));
 sg13g2_buf_2 fanout76 (.A(_4490_),
    .X(net76));
 sg13g2_buf_2 fanout77 (.A(_4363_),
    .X(net77));
 sg13g2_buf_2 fanout78 (.A(_4362_),
    .X(net78));
 sg13g2_buf_2 fanout79 (.A(_4295_),
    .X(net79));
 sg13g2_buf_2 fanout80 (.A(_0744_),
    .X(net80));
 sg13g2_buf_2 fanout81 (.A(_0740_),
    .X(net81));
 sg13g2_buf_2 fanout82 (.A(_0616_),
    .X(net82));
 sg13g2_buf_2 fanout83 (.A(_0607_),
    .X(net83));
 sg13g2_buf_2 fanout84 (.A(_0593_),
    .X(net84));
 sg13g2_buf_2 fanout85 (.A(_0390_),
    .X(net85));
 sg13g2_buf_2 fanout86 (.A(_0294_),
    .X(net86));
 sg13g2_buf_2 fanout87 (.A(_0290_),
    .X(net87));
 sg13g2_buf_2 fanout88 (.A(_4489_),
    .X(net88));
 sg13g2_buf_2 fanout89 (.A(_4445_),
    .X(net89));
 sg13g2_buf_2 fanout90 (.A(_4335_),
    .X(net90));
 sg13g2_buf_2 fanout91 (.A(_4194_),
    .X(net91));
 sg13g2_buf_2 fanout92 (.A(_0783_),
    .X(net92));
 sg13g2_buf_2 fanout93 (.A(_4331_),
    .X(net93));
 sg13g2_buf_2 fanout94 (.A(_4293_),
    .X(net94));
 sg13g2_buf_2 fanout95 (.A(_4163_),
    .X(net95));
 sg13g2_buf_4 fanout96 (.X(net96),
    .A(net98));
 sg13g2_buf_4 fanout97 (.X(net97),
    .A(net98));
 sg13g2_buf_2 fanout98 (.A(net99),
    .X(net98));
 sg13g2_buf_2 fanout99 (.A(net100),
    .X(net99));
 sg13g2_buf_4 fanout100 (.X(net100),
    .A(net101));
 sg13g2_buf_4 fanout101 (.X(net101),
    .A(net1));
 sg13g2_buf_4 fanout102 (.X(net102),
    .A(net104));
 sg13g2_buf_2 fanout103 (.A(net104),
    .X(net103));
 sg13g2_buf_4 fanout104 (.X(net104),
    .A(net105));
 sg13g2_buf_4 fanout105 (.X(net105),
    .A(net1));
 sg13g2_tielo _9148__106 (.L_LO(net106));
 sg13g2_tielo _9149__107 (.L_LO(net107));
 sg13g2_tielo _9150__108 (.L_LO(net108));
 sg13g2_tielo _9151__109 (.L_LO(net109));
 sg13g2_tielo _9152__110 (.L_LO(net110));
 sg13g2_tielo _9153__111 (.L_LO(net111));
 sg13g2_tielo _9154__112 (.L_LO(net112));
 sg13g2_tielo _9155__113 (.L_LO(net113));
 sg13g2_tielo _9156__114 (.L_LO(net114));
 sg13g2_tielo _9157__115 (.L_LO(net115));
 sg13g2_tielo _9158__116 (.L_LO(net116));
 sg13g2_tielo _9159__117 (.L_LO(net117));
 sg13g2_tielo _9160__118 (.L_LO(net118));
 sg13g2_tielo _9161__119 (.L_LO(net119));
 sg13g2_tielo _9162__120 (.L_LO(net120));
 sg13g2_tielo _9163__121 (.L_LO(net121));
 sg13g2_tiehi _9138__123 (.L_HI(net123));
 sg13g2_tiehi _9139__124 (.L_HI(net124));
 sg13g2_tiehi _9140__125 (.L_HI(net125));
 sg13g2_tiehi _9141__126 (.L_HI(net126));
 sg13g2_tiehi _9142__127 (.L_HI(net127));
 sg13g2_tiehi _9143__128 (.L_HI(net128));
 sg13g2_tiehi _9144__129 (.L_HI(net129));
 sg13g2_tiehi _9145__130 (.L_HI(net130));
 sg13g2_tiehi \generated._1020[0]$_SDFF_PP0__131  (.L_HI(net131));
 sg13g2_tiehi \generated._1020[1]$_SDFF_PP0__132  (.L_HI(net132));
 sg13g2_tiehi \generated._1020[2]$_SDFF_PP0__133  (.L_HI(net133));
 sg13g2_tiehi \generated._1020[3]$_DFF_P__134  (.L_HI(net134));
 sg13g2_tiehi \generated._1020[4]$_DFF_P__135  (.L_HI(net135));
 sg13g2_tiehi \generated._1020[5]$_DFF_P__136  (.L_HI(net136));
 sg13g2_tiehi \generated._1020[6]$_DFF_P__137  (.L_HI(net137));
 sg13g2_tiehi \generated._1020[7]$_DFF_P__138  (.L_HI(net138));
 sg13g2_tiehi \generated._1020[8]$_DFF_P__139  (.L_HI(net139));
 sg13g2_tiehi \generated._1020[9]$_DFF_P__140  (.L_HI(net140));
 sg13g2_tiehi \generated._1070[0]$_SDFF_PP0__141  (.L_HI(net141));
 sg13g2_tiehi \generated._1070[1]$_SDFF_PP0__142  (.L_HI(net142));
 sg13g2_tiehi \generated._1070[2]$_SDFF_PP0__143  (.L_HI(net143));
 sg13g2_tiehi \generated._1070[3]$_DFF_P__144  (.L_HI(net144));
 sg13g2_tiehi \generated._1070[4]$_DFF_P__145  (.L_HI(net145));
 sg13g2_tiehi \generated._1070[5]$_DFF_P__146  (.L_HI(net146));
 sg13g2_tiehi \generated._1070[6]$_DFF_P__147  (.L_HI(net147));
 sg13g2_tiehi \generated._1070[7]$_DFF_P__148  (.L_HI(net148));
 sg13g2_tiehi \generated._1070[8]$_DFF_P__149  (.L_HI(net149));
 sg13g2_tiehi \generated._1070[9]$_DFF_P__150  (.L_HI(net150));
 sg13g2_tiehi \generated._1080[0]$_SDFF_PP0__151  (.L_HI(net151));
 sg13g2_tiehi \generated._1080[1]$_SDFF_PP0__152  (.L_HI(net152));
 sg13g2_tiehi \generated._1080[2]$_SDFF_PP0__153  (.L_HI(net153));
 sg13g2_tiehi \generated._1080[3]$_SDFF_PP0__154  (.L_HI(net154));
 sg13g2_tiehi \generated._1080[4]$_SDFF_PP0__155  (.L_HI(net155));
 sg13g2_tiehi \generated._1080[5]$_SDFF_PP0__156  (.L_HI(net156));
 sg13g2_tiehi \generated._1080[6]$_SDFF_PP0__157  (.L_HI(net157));
 sg13g2_tiehi \generated._1080[7]$_SDFF_PP0__158  (.L_HI(net158));
 sg13g2_tiehi \generated._1080[8]$_SDFF_PP0__159  (.L_HI(net159));
 sg13g2_tiehi \generated._1080[9]$_SDFF_PP0__160  (.L_HI(net160));
 sg13g2_tiehi \generated._222[1]$_DFF_P__161  (.L_HI(net161));
 sg13g2_tiehi \generated._287[0]$_SDFFE_PP0N__162  (.L_HI(net162));
 sg13g2_tiehi \generated._287[1]$_SDFFE_PP0N__163  (.L_HI(net163));
 sg13g2_tiehi \generated._287[2]$_SDFFE_PP0N__164  (.L_HI(net164));
 sg13g2_tiehi \generated._287[3]$_SDFFE_PP0N__165  (.L_HI(net165));
 sg13g2_tiehi \generated._287[4]$_SDFFE_PP0N__166  (.L_HI(net166));
 sg13g2_tiehi \generated._301[0]$_SDFF_PP0__167  (.L_HI(net167));
 sg13g2_tiehi \generated._301[1]$_SDFF_PP0__168  (.L_HI(net168));
 sg13g2_tiehi \generated._301[2]$_SDFF_PP0__169  (.L_HI(net169));
 sg13g2_tiehi \generated._301[3]$_SDFF_PP0__170  (.L_HI(net170));
 sg13g2_tiehi \generated._301[4]$_SDFF_PP0__171  (.L_HI(net171));
 sg13g2_tiehi \generated._315[0]$_SDFFE_PP0P__172  (.L_HI(net172));
 sg13g2_tiehi \generated._315[1]$_SDFFE_PP0P__173  (.L_HI(net173));
 sg13g2_tiehi \generated._315[2]$_SDFFE_PP0P__174  (.L_HI(net174));
 sg13g2_tiehi \generated._315[3]$_SDFFE_PP0P__175  (.L_HI(net175));
 sg13g2_tiehi \generated._328[0]$_SDFF_PP0__176  (.L_HI(net176));
 sg13g2_tiehi \generated._328[1]$_SDFF_PP0__177  (.L_HI(net177));
 sg13g2_tiehi \generated._328[2]$_SDFF_PP0__178  (.L_HI(net178));
 sg13g2_tiehi \generated._328[3]$_SDFF_PP0__179  (.L_HI(net179));
 sg13g2_tiehi \generated._328[4]$_SDFF_PP0__180  (.L_HI(net180));
 sg13g2_tiehi \generated._328[5]$_SDFF_PP0__181  (.L_HI(net181));
 sg13g2_tiehi \generated._328[6]$_SDFF_PP0__182  (.L_HI(net182));
 sg13g2_tiehi \generated._342[0]$_SDFFE_PP0N__183  (.L_HI(net183));
 sg13g2_tiehi \generated._342[1]$_SDFFE_PP0N__184  (.L_HI(net184));
 sg13g2_tiehi \generated._342[2]$_SDFFE_PP0N__185  (.L_HI(net185));
 sg13g2_tiehi \generated._342[3]$_SDFFE_PP0N__186  (.L_HI(net186));
 sg13g2_tiehi \generated._342[4]$_SDFFE_PP0N__187  (.L_HI(net187));
 sg13g2_tiehi \generated._342[5]$_SDFFE_PP0N__188  (.L_HI(net188));
 sg13g2_tiehi \generated._353[0]$_SDFF_PP0__189  (.L_HI(net189));
 sg13g2_tiehi \generated._353[1]$_SDFF_PP0__190  (.L_HI(net190));
 sg13g2_tiehi \generated._353[2]$_SDFF_PP0__191  (.L_HI(net191));
 sg13g2_tiehi \generated._353[3]$_SDFF_PP0__192  (.L_HI(net192));
 sg13g2_tiehi \generated._353[4]$_SDFF_PP0__193  (.L_HI(net193));
 sg13g2_tiehi \generated._390[0]$_SDFF_PP0__194  (.L_HI(net194));
 sg13g2_tiehi \generated._390[1]$_SDFF_PP0__195  (.L_HI(net195));
 sg13g2_tiehi \generated._390[2]$_SDFF_PP1__196  (.L_HI(net196));
 sg13g2_tiehi \generated._390[3]$_SDFF_PP1__197  (.L_HI(net197));
 sg13g2_tiehi \generated._390[4]$_SDFF_PP1__198  (.L_HI(net198));
 sg13g2_tiehi \generated._390[5]$_SDFF_PP0__199  (.L_HI(net199));
 sg13g2_tiehi \generated._390[6]$_SDFF_PP0__200  (.L_HI(net200));
 sg13g2_tiehi \generated._390[7]$_SDFF_PP1__201  (.L_HI(net201));
 sg13g2_tiehi \generated._390[8]$_SDFF_PP0__202  (.L_HI(net202));
 sg13g2_tiehi \generated._390[9]$_SDFF_PP0__203  (.L_HI(net203));
 sg13g2_tiehi \generated._478[0]$_DFF_P__204  (.L_HI(net204));
 sg13g2_tiehi \generated._478[1]$_DFF_P__205  (.L_HI(net205));
 sg13g2_tiehi \generated._478[2]$_DFF_P__206  (.L_HI(net206));
 sg13g2_tiehi \generated._478[3]$_DFF_P__207  (.L_HI(net207));
 sg13g2_tiehi \generated._478[4]$_DFF_P__208  (.L_HI(net208));
 sg13g2_tiehi \generated._478[5]$_DFF_P__209  (.L_HI(net209));
 sg13g2_tiehi \generated._478[6]$_DFF_P__210  (.L_HI(net210));
 sg13g2_tiehi \generated._478[7]$_DFF_P__211  (.L_HI(net211));
 sg13g2_tiehi \generated._478[8]$_DFF_P__212  (.L_HI(net212));
 sg13g2_tiehi \generated._478[9]$_DFF_P__213  (.L_HI(net213));
 sg13g2_tiehi \generated._497[0]$_SDFF_PP0__214  (.L_HI(net214));
 sg13g2_tiehi \generated._497[1]$_SDFF_PP0__215  (.L_HI(net215));
 sg13g2_tiehi \generated._497[2]$_SDFF_PP0__216  (.L_HI(net216));
 sg13g2_tiehi \generated._497[3]$_SDFF_PP0__217  (.L_HI(net217));
 sg13g2_tiehi \generated._497[4]$_SDFF_PP0__218  (.L_HI(net218));
 sg13g2_tiehi \generated._497[5]$_SDFF_PP0__219  (.L_HI(net219));
 sg13g2_tiehi \generated._497[6]$_SDFF_PP0__220  (.L_HI(net220));
 sg13g2_tiehi \generated._497[7]$_SDFF_PP0__221  (.L_HI(net221));
 sg13g2_tiehi \generated._497[8]$_SDFF_PP0__222  (.L_HI(net222));
 sg13g2_tiehi \generated._497[9]$_SDFF_PP0__223  (.L_HI(net223));
 sg13g2_tiehi \generated._558[0]$_DFF_P__224  (.L_HI(net224));
 sg13g2_tiehi \generated._558[1]$_DFF_P__225  (.L_HI(net225));
 sg13g2_tiehi \generated._558[2]$_DFF_P__226  (.L_HI(net226));
 sg13g2_tiehi \generated._558[3]$_DFF_P__227  (.L_HI(net227));
 sg13g2_tiehi \generated._558[4]$_DFF_P__228  (.L_HI(net228));
 sg13g2_tiehi \generated._558[5]$_DFF_P__229  (.L_HI(net229));
 sg13g2_tiehi \generated._558[6]$_DFF_P__230  (.L_HI(net230));
 sg13g2_tiehi \generated._558[7]$_DFF_P__231  (.L_HI(net231));
 sg13g2_tiehi \generated._558[8]$_DFF_P__232  (.L_HI(net232));
 sg13g2_tiehi \generated._558[9]$_DFF_P__233  (.L_HI(net233));
 sg13g2_tiehi \generated._692[0]$_DFF_P__234  (.L_HI(net234));
 sg13g2_tiehi \generated._692[1]$_DFF_P__235  (.L_HI(net235));
 sg13g2_tiehi \generated._692[2]$_DFF_P__236  (.L_HI(net236));
 sg13g2_tiehi \generated._692[3]$_DFF_P__237  (.L_HI(net237));
 sg13g2_tiehi \generated._692[4]$_DFF_P__238  (.L_HI(net238));
 sg13g2_tiehi \generated._692[5]$_DFF_P__239  (.L_HI(net239));
 sg13g2_tiehi \generated._692[6]$_DFF_P__240  (.L_HI(net240));
 sg13g2_tiehi \generated._692[7]$_DFF_P__241  (.L_HI(net241));
 sg13g2_tiehi \generated._692[8]$_DFF_P__242  (.L_HI(net242));
 sg13g2_tiehi \generated._692[9]$_DFF_P__243  (.L_HI(net243));
 sg13g2_tiehi \generated._710[0]$_SDFF_PP0__244  (.L_HI(net244));
 sg13g2_tiehi \generated._710[1]$_SDFF_PP0__245  (.L_HI(net245));
 sg13g2_tiehi \generated._710[2]$_SDFF_PP0__246  (.L_HI(net246));
 sg13g2_tiehi \generated._710[3]$_SDFF_PP0__247  (.L_HI(net247));
 sg13g2_tiehi \generated._710[4]$_SDFF_PP0__248  (.L_HI(net248));
 sg13g2_tiehi \generated._710[5]$_SDFF_PP0__249  (.L_HI(net249));
 sg13g2_tiehi \generated._710[6]$_SDFF_PP0__250  (.L_HI(net250));
 sg13g2_tiehi \generated._710[7]$_SDFF_PP0__251  (.L_HI(net251));
 sg13g2_tiehi \generated._710[8]$_SDFF_PP0__252  (.L_HI(net252));
 sg13g2_tiehi \generated._710[9]$_SDFF_PP0__253  (.L_HI(net253));
 sg13g2_tiehi \generated._886[0]$_SDFF_PP0__254  (.L_HI(net254));
 sg13g2_tiehi \generated._886[1]$_SDFF_PP0__255  (.L_HI(net255));
 sg13g2_tiehi \generated._886[2]$_SDFF_PP0__256  (.L_HI(net256));
 sg13g2_tiehi \generated._886[3]$_DFF_P__257  (.L_HI(net257));
 sg13g2_tiehi \generated._886[4]$_DFF_P__258  (.L_HI(net258));
 sg13g2_tiehi \generated._886[5]$_DFF_P__259  (.L_HI(net259));
 sg13g2_tiehi \generated._886[6]$_DFF_P__260  (.L_HI(net260));
 sg13g2_tiehi \generated._886[7]$_DFF_P__261  (.L_HI(net261));
 sg13g2_tiehi \generated._886[8]$_DFF_P__262  (.L_HI(net262));
 sg13g2_tiehi \generated._886[9]$_DFF_P__263  (.L_HI(net263));
 sg13g2_tiehi \generated._935[0]$_SDFF_PP0__264  (.L_HI(net264));
 sg13g2_tiehi \generated._935[1]$_SDFF_PP0__265  (.L_HI(net265));
 sg13g2_tiehi \generated._935[2]$_SDFF_PP0__266  (.L_HI(net266));
 sg13g2_tiehi \generated._935[3]$_DFF_P__267  (.L_HI(net267));
 sg13g2_tiehi \generated._935[4]$_DFF_P__268  (.L_HI(net268));
 sg13g2_tiehi \generated._935[5]$_DFF_P__269  (.L_HI(net269));
 sg13g2_tiehi \generated._935[6]$_DFF_P__270  (.L_HI(net270));
 sg13g2_tiehi \generated._935[7]$_DFF_P__271  (.L_HI(net271));
 sg13g2_tiehi \generated._935[8]$_DFF_P__272  (.L_HI(net272));
 sg13g2_tiehi \generated._935[9]$_DFF_P__273  (.L_HI(net273));
 sg13g2_tiehi \generated._945[0]$_SDFF_PP0__274  (.L_HI(net274));
 sg13g2_tiehi \generated._945[1]$_SDFF_PP0__275  (.L_HI(net275));
 sg13g2_tiehi \generated._945[2]$_SDFF_PP0__276  (.L_HI(net276));
 sg13g2_tiehi \generated._945[3]$_SDFF_PP0__277  (.L_HI(net277));
 sg13g2_tiehi \generated._945[4]$_SDFF_PP0__278  (.L_HI(net278));
 sg13g2_tiehi \generated._945[5]$_SDFF_PP0__279  (.L_HI(net279));
 sg13g2_tiehi \generated._945[6]$_SDFF_PP0__280  (.L_HI(net280));
 sg13g2_tiehi \generated._945[7]$_SDFF_PP0__281  (.L_HI(net281));
 sg13g2_tiehi \generated._945[8]$_SDFF_PP0__282  (.L_HI(net282));
 sg13g2_tiehi \generated._945[9]$_SDFF_PP0__283  (.L_HI(net283));
 sg13g2_tiehi \generated.iter_sel[0]$_SDFF_PP0__284  (.L_HI(net284));
 sg13g2_tiehi \generated.iter_sel[1]$_SDFF_PP0__285  (.L_HI(net285));
 sg13g2_tiehi \generated.iter_sel_0[0]$_SDFF_PP0__286  (.L_HI(net286));
 sg13g2_tiehi \generated.iter_sel_0[1]$_SDFF_PP0__287  (.L_HI(net287));
 sg13g2_tiehi \generated.iter_sel_1[0]$_SDFF_PP0__288  (.L_HI(net288));
 sg13g2_tiehi \generated.iter_sel_1[1]$_SDFF_PP0__289  (.L_HI(net289));
 sg13g2_tiehi \generated.iter_sel_2[0]$_SDFF_PP0__290  (.L_HI(net290));
 sg13g2_tiehi \generated.iter_sel_2[1]$_SDFF_PP0__291  (.L_HI(net291));
 sg13g2_buf_2 clkbuf_leaf_1_clk (.A(clknet_3_0__leaf_clk),
    .X(clknet_leaf_1_clk));
 sg13g2_buf_2 clkbuf_leaf_2_clk (.A(clknet_3_0__leaf_clk),
    .X(clknet_leaf_2_clk));
 sg13g2_buf_2 clkbuf_leaf_3_clk (.A(clknet_3_1__leaf_clk),
    .X(clknet_leaf_3_clk));
 sg13g2_buf_2 clkbuf_leaf_4_clk (.A(clknet_3_1__leaf_clk),
    .X(clknet_leaf_4_clk));
 sg13g2_buf_2 clkbuf_leaf_5_clk (.A(clknet_3_4__leaf_clk),
    .X(clknet_leaf_5_clk));
 sg13g2_buf_2 clkbuf_leaf_6_clk (.A(clknet_3_4__leaf_clk),
    .X(clknet_leaf_6_clk));
 sg13g2_buf_2 clkbuf_leaf_7_clk (.A(clknet_3_4__leaf_clk),
    .X(clknet_leaf_7_clk));
 sg13g2_buf_2 clkbuf_leaf_8_clk (.A(clknet_3_4__leaf_clk),
    .X(clknet_leaf_8_clk));
 sg13g2_buf_2 clkbuf_leaf_9_clk (.A(clknet_3_4__leaf_clk),
    .X(clknet_leaf_9_clk));
 sg13g2_buf_2 clkbuf_leaf_10_clk (.A(clknet_3_5__leaf_clk),
    .X(clknet_leaf_10_clk));
 sg13g2_buf_2 clkbuf_leaf_11_clk (.A(clknet_3_5__leaf_clk),
    .X(clknet_leaf_11_clk));
 sg13g2_buf_2 clkbuf_leaf_12_clk (.A(clknet_3_5__leaf_clk),
    .X(clknet_leaf_12_clk));
 sg13g2_buf_2 clkbuf_leaf_13_clk (.A(clknet_3_5__leaf_clk),
    .X(clknet_leaf_13_clk));
 sg13g2_buf_2 clkbuf_leaf_14_clk (.A(clknet_3_7__leaf_clk),
    .X(clknet_leaf_14_clk));
 sg13g2_buf_2 clkbuf_leaf_15_clk (.A(clknet_3_6__leaf_clk),
    .X(clknet_leaf_15_clk));
 sg13g2_buf_2 clkbuf_leaf_16_clk (.A(clknet_3_6__leaf_clk),
    .X(clknet_leaf_16_clk));
 sg13g2_buf_2 clkbuf_leaf_17_clk (.A(clknet_3_7__leaf_clk),
    .X(clknet_leaf_17_clk));
 sg13g2_buf_2 clkbuf_leaf_19_clk (.A(clknet_3_7__leaf_clk),
    .X(clknet_leaf_19_clk));
 sg13g2_buf_2 clkbuf_leaf_20_clk (.A(clknet_3_6__leaf_clk),
    .X(clknet_leaf_20_clk));
 sg13g2_buf_2 clkbuf_leaf_21_clk (.A(clknet_3_6__leaf_clk),
    .X(clknet_leaf_21_clk));
 sg13g2_buf_2 clkbuf_leaf_22_clk (.A(clknet_3_3__leaf_clk),
    .X(clknet_leaf_22_clk));
 sg13g2_buf_2 clkbuf_leaf_23_clk (.A(clknet_3_3__leaf_clk),
    .X(clknet_leaf_23_clk));
 sg13g2_buf_2 clkbuf_leaf_24_clk (.A(clknet_3_3__leaf_clk),
    .X(clknet_leaf_24_clk));
 sg13g2_buf_2 clkbuf_leaf_25_clk (.A(clknet_3_2__leaf_clk),
    .X(clknet_leaf_25_clk));
 sg13g2_buf_2 clkbuf_leaf_26_clk (.A(clknet_3_2__leaf_clk),
    .X(clknet_leaf_26_clk));
 sg13g2_buf_2 clkbuf_leaf_27_clk (.A(clknet_3_2__leaf_clk),
    .X(clknet_leaf_27_clk));
 sg13g2_buf_2 clkbuf_leaf_28_clk (.A(clknet_3_3__leaf_clk),
    .X(clknet_leaf_28_clk));
 sg13g2_buf_2 clkbuf_leaf_29_clk (.A(clknet_3_1__leaf_clk),
    .X(clknet_leaf_29_clk));
 sg13g2_buf_2 clkbuf_leaf_30_clk (.A(clknet_3_1__leaf_clk),
    .X(clknet_leaf_30_clk));
 sg13g2_buf_2 clkbuf_leaf_31_clk (.A(clknet_3_0__leaf_clk),
    .X(clknet_leaf_31_clk));
 sg13g2_buf_2 clkbuf_leaf_32_clk (.A(clknet_3_2__leaf_clk),
    .X(clknet_leaf_32_clk));
 sg13g2_buf_2 clkbuf_leaf_33_clk (.A(clknet_3_2__leaf_clk),
    .X(clknet_leaf_33_clk));
 sg13g2_buf_2 clkbuf_leaf_34_clk (.A(clknet_3_0__leaf_clk),
    .X(clknet_leaf_34_clk));
 sg13g2_buf_1 clkbuf_0_clk (.A(clk),
    .X(clknet_0_clk));
 sg13g2_buf_1 clkbuf_3_0__f_clk (.A(clknet_0_clk),
    .X(clknet_3_0__leaf_clk));
 sg13g2_buf_1 clkbuf_3_1__f_clk (.A(clknet_0_clk),
    .X(clknet_3_1__leaf_clk));
 sg13g2_buf_1 clkbuf_3_2__f_clk (.A(clknet_0_clk),
    .X(clknet_3_2__leaf_clk));
 sg13g2_buf_1 clkbuf_3_3__f_clk (.A(clknet_0_clk),
    .X(clknet_3_3__leaf_clk));
 sg13g2_buf_1 clkbuf_3_4__f_clk (.A(clknet_0_clk),
    .X(clknet_3_4__leaf_clk));
 sg13g2_buf_1 clkbuf_3_5__f_clk (.A(clknet_0_clk),
    .X(clknet_3_5__leaf_clk));
 sg13g2_buf_1 clkbuf_3_6__f_clk (.A(clknet_0_clk),
    .X(clknet_3_6__leaf_clk));
 sg13g2_buf_1 clkbuf_3_7__f_clk (.A(clknet_0_clk),
    .X(clknet_3_7__leaf_clk));
 sg13g2_buf_2 clkload0 (.A(clknet_3_1__leaf_clk));
 sg13g2_buf_2 clkload1 (.A(clknet_3_3__leaf_clk));
 sg13g2_buf_2 clkload2 (.A(clknet_3_5__leaf_clk));
 sg13g2_buf_2 clkload3 (.A(clknet_3_6__leaf_clk));
 sg13g2_buf_1 clkload4 (.A(clknet_3_7__leaf_clk));
 sg13g2_buf_16 clkload5 (.A(clknet_leaf_29_clk));
 sg13g2_inv_2 clkload6 (.A(clknet_leaf_25_clk));
 sg13g2_buf_16 clkload7 (.A(clknet_leaf_27_clk));
 sg13g2_buf_16 clkload8 (.A(clknet_leaf_32_clk));
 sg13g2_buf_8 clkload9 (.A(clknet_leaf_33_clk));
 sg13g2_buf_8 clkload10 (.A(clknet_leaf_22_clk));
 sg13g2_inv_2 clkload11 (.A(clknet_leaf_5_clk));
 sg13g2_inv_4 clkload12 (.A(clknet_leaf_7_clk));
 sg13g2_inv_4 clkload13 (.A(clknet_leaf_8_clk));
 sg13g2_buf_16 clkload14 (.A(clknet_leaf_20_clk));
 sg13g2_buf_8 clkload15 (.A(clknet_leaf_21_clk));
 sg13g2_buf_8 clkload16 (.A(clknet_leaf_19_clk));
 sg13g2_antennanp ANTENNA_1 (.A(clk));
 sg13g2_antennanp ANTENNA_2 (.A(clk));
 sg13g2_antennanp ANTENNA_3 (.A(clk));
 sg13g2_antennanp ANTENNA_4 (.A(clk));
 sg13g2_antennanp ANTENNA_5 (.A(clk));
 sg13g2_antennanp ANTENNA_6 (.A(clk));
 sg13g2_decap_8 FILLER_0_0 ();
 sg13g2_decap_8 FILLER_0_7 ();
 sg13g2_decap_8 FILLER_0_14 ();
 sg13g2_decap_8 FILLER_0_21 ();
 sg13g2_decap_8 FILLER_0_28 ();
 sg13g2_decap_8 FILLER_0_35 ();
 sg13g2_decap_8 FILLER_0_42 ();
 sg13g2_decap_8 FILLER_0_49 ();
 sg13g2_decap_8 FILLER_0_56 ();
 sg13g2_decap_8 FILLER_0_63 ();
 sg13g2_decap_8 FILLER_0_70 ();
 sg13g2_decap_8 FILLER_0_77 ();
 sg13g2_decap_8 FILLER_0_84 ();
 sg13g2_decap_8 FILLER_0_91 ();
 sg13g2_decap_8 FILLER_0_98 ();
 sg13g2_decap_8 FILLER_0_105 ();
 sg13g2_decap_8 FILLER_0_112 ();
 sg13g2_decap_8 FILLER_0_119 ();
 sg13g2_decap_8 FILLER_0_126 ();
 sg13g2_decap_8 FILLER_0_133 ();
 sg13g2_decap_8 FILLER_0_140 ();
 sg13g2_decap_8 FILLER_0_147 ();
 sg13g2_decap_8 FILLER_0_154 ();
 sg13g2_fill_1 FILLER_0_161 ();
 sg13g2_fill_1 FILLER_0_188 ();
 sg13g2_fill_1 FILLER_0_215 ();
 sg13g2_fill_1 FILLER_0_221 ();
 sg13g2_fill_1 FILLER_0_230 ();
 sg13g2_fill_1 FILLER_0_248 ();
 sg13g2_fill_1 FILLER_0_281 ();
 sg13g2_fill_2 FILLER_0_286 ();
 sg13g2_decap_8 FILLER_0_296 ();
 sg13g2_decap_8 FILLER_0_303 ();
 sg13g2_decap_8 FILLER_0_310 ();
 sg13g2_decap_8 FILLER_0_317 ();
 sg13g2_decap_8 FILLER_0_324 ();
 sg13g2_decap_8 FILLER_0_331 ();
 sg13g2_decap_8 FILLER_0_338 ();
 sg13g2_decap_8 FILLER_0_345 ();
 sg13g2_decap_8 FILLER_0_352 ();
 sg13g2_decap_8 FILLER_0_359 ();
 sg13g2_decap_8 FILLER_0_366 ();
 sg13g2_decap_8 FILLER_0_373 ();
 sg13g2_decap_8 FILLER_0_380 ();
 sg13g2_decap_8 FILLER_0_387 ();
 sg13g2_decap_8 FILLER_0_394 ();
 sg13g2_decap_8 FILLER_0_401 ();
 sg13g2_decap_8 FILLER_0_408 ();
 sg13g2_decap_8 FILLER_0_415 ();
 sg13g2_decap_8 FILLER_0_422 ();
 sg13g2_fill_1 FILLER_0_429 ();
 sg13g2_decap_8 FILLER_1_0 ();
 sg13g2_decap_8 FILLER_1_7 ();
 sg13g2_decap_8 FILLER_1_14 ();
 sg13g2_decap_8 FILLER_1_21 ();
 sg13g2_decap_8 FILLER_1_28 ();
 sg13g2_decap_8 FILLER_1_35 ();
 sg13g2_decap_8 FILLER_1_42 ();
 sg13g2_decap_8 FILLER_1_49 ();
 sg13g2_decap_8 FILLER_1_56 ();
 sg13g2_decap_8 FILLER_1_63 ();
 sg13g2_decap_8 FILLER_1_70 ();
 sg13g2_decap_8 FILLER_1_77 ();
 sg13g2_decap_8 FILLER_1_84 ();
 sg13g2_decap_8 FILLER_1_91 ();
 sg13g2_decap_8 FILLER_1_98 ();
 sg13g2_decap_8 FILLER_1_105 ();
 sg13g2_decap_8 FILLER_1_112 ();
 sg13g2_decap_8 FILLER_1_119 ();
 sg13g2_decap_8 FILLER_1_126 ();
 sg13g2_decap_8 FILLER_1_133 ();
 sg13g2_decap_8 FILLER_1_140 ();
 sg13g2_decap_8 FILLER_1_147 ();
 sg13g2_fill_2 FILLER_1_154 ();
 sg13g2_fill_1 FILLER_1_156 ();
 sg13g2_fill_2 FILLER_1_164 ();
 sg13g2_fill_2 FILLER_1_173 ();
 sg13g2_fill_1 FILLER_1_202 ();
 sg13g2_fill_1 FILLER_1_309 ();
 sg13g2_decap_8 FILLER_1_314 ();
 sg13g2_decap_8 FILLER_1_321 ();
 sg13g2_decap_8 FILLER_1_328 ();
 sg13g2_decap_8 FILLER_1_335 ();
 sg13g2_decap_8 FILLER_1_342 ();
 sg13g2_decap_8 FILLER_1_349 ();
 sg13g2_decap_8 FILLER_1_356 ();
 sg13g2_decap_8 FILLER_1_363 ();
 sg13g2_decap_8 FILLER_1_370 ();
 sg13g2_decap_8 FILLER_1_377 ();
 sg13g2_decap_8 FILLER_1_384 ();
 sg13g2_decap_8 FILLER_1_391 ();
 sg13g2_decap_8 FILLER_1_398 ();
 sg13g2_decap_8 FILLER_1_405 ();
 sg13g2_decap_8 FILLER_1_412 ();
 sg13g2_decap_8 FILLER_1_419 ();
 sg13g2_decap_4 FILLER_1_426 ();
 sg13g2_decap_8 FILLER_2_0 ();
 sg13g2_decap_8 FILLER_2_7 ();
 sg13g2_decap_8 FILLER_2_14 ();
 sg13g2_decap_8 FILLER_2_21 ();
 sg13g2_decap_8 FILLER_2_28 ();
 sg13g2_decap_8 FILLER_2_35 ();
 sg13g2_decap_8 FILLER_2_42 ();
 sg13g2_decap_8 FILLER_2_49 ();
 sg13g2_decap_8 FILLER_2_56 ();
 sg13g2_decap_8 FILLER_2_63 ();
 sg13g2_decap_8 FILLER_2_70 ();
 sg13g2_decap_8 FILLER_2_77 ();
 sg13g2_decap_8 FILLER_2_84 ();
 sg13g2_decap_8 FILLER_2_91 ();
 sg13g2_decap_8 FILLER_2_98 ();
 sg13g2_decap_8 FILLER_2_105 ();
 sg13g2_decap_8 FILLER_2_112 ();
 sg13g2_decap_8 FILLER_2_119 ();
 sg13g2_decap_8 FILLER_2_126 ();
 sg13g2_decap_8 FILLER_2_133 ();
 sg13g2_decap_8 FILLER_2_140 ();
 sg13g2_fill_2 FILLER_2_147 ();
 sg13g2_fill_1 FILLER_2_149 ();
 sg13g2_fill_1 FILLER_2_179 ();
 sg13g2_fill_1 FILLER_2_288 ();
 sg13g2_decap_8 FILLER_2_303 ();
 sg13g2_decap_8 FILLER_2_310 ();
 sg13g2_decap_8 FILLER_2_317 ();
 sg13g2_decap_8 FILLER_2_324 ();
 sg13g2_decap_8 FILLER_2_331 ();
 sg13g2_decap_8 FILLER_2_338 ();
 sg13g2_decap_8 FILLER_2_345 ();
 sg13g2_decap_8 FILLER_2_352 ();
 sg13g2_decap_8 FILLER_2_359 ();
 sg13g2_decap_8 FILLER_2_366 ();
 sg13g2_decap_8 FILLER_2_373 ();
 sg13g2_decap_8 FILLER_2_380 ();
 sg13g2_decap_8 FILLER_2_387 ();
 sg13g2_decap_8 FILLER_2_394 ();
 sg13g2_decap_8 FILLER_2_401 ();
 sg13g2_decap_8 FILLER_2_408 ();
 sg13g2_decap_8 FILLER_2_415 ();
 sg13g2_decap_8 FILLER_2_422 ();
 sg13g2_fill_1 FILLER_2_429 ();
 sg13g2_decap_8 FILLER_3_0 ();
 sg13g2_decap_8 FILLER_3_7 ();
 sg13g2_decap_8 FILLER_3_14 ();
 sg13g2_decap_8 FILLER_3_21 ();
 sg13g2_decap_8 FILLER_3_28 ();
 sg13g2_decap_8 FILLER_3_35 ();
 sg13g2_decap_8 FILLER_3_42 ();
 sg13g2_decap_8 FILLER_3_49 ();
 sg13g2_decap_8 FILLER_3_56 ();
 sg13g2_decap_8 FILLER_3_63 ();
 sg13g2_decap_8 FILLER_3_70 ();
 sg13g2_decap_8 FILLER_3_77 ();
 sg13g2_decap_8 FILLER_3_84 ();
 sg13g2_decap_8 FILLER_3_91 ();
 sg13g2_decap_8 FILLER_3_98 ();
 sg13g2_decap_8 FILLER_3_105 ();
 sg13g2_decap_8 FILLER_3_112 ();
 sg13g2_decap_8 FILLER_3_119 ();
 sg13g2_decap_8 FILLER_3_126 ();
 sg13g2_decap_8 FILLER_3_133 ();
 sg13g2_decap_8 FILLER_3_140 ();
 sg13g2_decap_4 FILLER_3_147 ();
 sg13g2_fill_1 FILLER_3_151 ();
 sg13g2_fill_2 FILLER_3_157 ();
 sg13g2_fill_1 FILLER_3_206 ();
 sg13g2_fill_2 FILLER_3_269 ();
 sg13g2_decap_8 FILLER_3_310 ();
 sg13g2_decap_8 FILLER_3_317 ();
 sg13g2_decap_4 FILLER_3_324 ();
 sg13g2_decap_8 FILLER_3_354 ();
 sg13g2_decap_8 FILLER_3_361 ();
 sg13g2_decap_8 FILLER_3_368 ();
 sg13g2_decap_8 FILLER_3_375 ();
 sg13g2_decap_8 FILLER_3_382 ();
 sg13g2_decap_8 FILLER_3_389 ();
 sg13g2_decap_8 FILLER_3_396 ();
 sg13g2_decap_8 FILLER_3_403 ();
 sg13g2_decap_8 FILLER_3_410 ();
 sg13g2_decap_8 FILLER_3_417 ();
 sg13g2_decap_4 FILLER_3_424 ();
 sg13g2_fill_2 FILLER_3_428 ();
 sg13g2_decap_8 FILLER_4_0 ();
 sg13g2_decap_8 FILLER_4_7 ();
 sg13g2_decap_8 FILLER_4_14 ();
 sg13g2_decap_8 FILLER_4_21 ();
 sg13g2_decap_8 FILLER_4_28 ();
 sg13g2_decap_8 FILLER_4_35 ();
 sg13g2_decap_8 FILLER_4_42 ();
 sg13g2_decap_8 FILLER_4_49 ();
 sg13g2_decap_8 FILLER_4_56 ();
 sg13g2_decap_8 FILLER_4_63 ();
 sg13g2_decap_8 FILLER_4_70 ();
 sg13g2_decap_8 FILLER_4_77 ();
 sg13g2_decap_8 FILLER_4_84 ();
 sg13g2_decap_8 FILLER_4_91 ();
 sg13g2_decap_8 FILLER_4_98 ();
 sg13g2_decap_8 FILLER_4_105 ();
 sg13g2_decap_8 FILLER_4_112 ();
 sg13g2_decap_8 FILLER_4_119 ();
 sg13g2_decap_8 FILLER_4_126 ();
 sg13g2_fill_2 FILLER_4_133 ();
 sg13g2_fill_1 FILLER_4_135 ();
 sg13g2_fill_1 FILLER_4_202 ();
 sg13g2_fill_1 FILLER_4_249 ();
 sg13g2_fill_1 FILLER_4_277 ();
 sg13g2_fill_2 FILLER_4_286 ();
 sg13g2_fill_1 FILLER_4_317 ();
 sg13g2_decap_8 FILLER_4_354 ();
 sg13g2_decap_8 FILLER_4_361 ();
 sg13g2_decap_8 FILLER_4_368 ();
 sg13g2_decap_8 FILLER_4_375 ();
 sg13g2_decap_8 FILLER_4_382 ();
 sg13g2_decap_8 FILLER_4_389 ();
 sg13g2_decap_8 FILLER_4_396 ();
 sg13g2_decap_8 FILLER_4_403 ();
 sg13g2_decap_8 FILLER_4_410 ();
 sg13g2_decap_8 FILLER_4_417 ();
 sg13g2_decap_4 FILLER_4_424 ();
 sg13g2_fill_2 FILLER_4_428 ();
 sg13g2_decap_8 FILLER_5_0 ();
 sg13g2_decap_8 FILLER_5_7 ();
 sg13g2_decap_8 FILLER_5_14 ();
 sg13g2_decap_8 FILLER_5_21 ();
 sg13g2_decap_8 FILLER_5_28 ();
 sg13g2_decap_8 FILLER_5_35 ();
 sg13g2_decap_8 FILLER_5_42 ();
 sg13g2_decap_8 FILLER_5_49 ();
 sg13g2_decap_8 FILLER_5_56 ();
 sg13g2_decap_8 FILLER_5_63 ();
 sg13g2_decap_8 FILLER_5_70 ();
 sg13g2_decap_8 FILLER_5_77 ();
 sg13g2_decap_8 FILLER_5_84 ();
 sg13g2_decap_8 FILLER_5_91 ();
 sg13g2_decap_8 FILLER_5_98 ();
 sg13g2_decap_8 FILLER_5_105 ();
 sg13g2_decap_8 FILLER_5_112 ();
 sg13g2_decap_4 FILLER_5_119 ();
 sg13g2_decap_4 FILLER_5_133 ();
 sg13g2_fill_2 FILLER_5_137 ();
 sg13g2_fill_1 FILLER_5_147 ();
 sg13g2_fill_2 FILLER_5_179 ();
 sg13g2_fill_2 FILLER_5_210 ();
 sg13g2_fill_1 FILLER_5_281 ();
 sg13g2_fill_1 FILLER_5_286 ();
 sg13g2_decap_8 FILLER_5_360 ();
 sg13g2_decap_8 FILLER_5_367 ();
 sg13g2_decap_8 FILLER_5_374 ();
 sg13g2_decap_8 FILLER_5_381 ();
 sg13g2_decap_8 FILLER_5_388 ();
 sg13g2_decap_8 FILLER_5_395 ();
 sg13g2_decap_8 FILLER_5_402 ();
 sg13g2_decap_8 FILLER_5_409 ();
 sg13g2_decap_8 FILLER_5_416 ();
 sg13g2_decap_8 FILLER_5_423 ();
 sg13g2_decap_8 FILLER_6_0 ();
 sg13g2_decap_8 FILLER_6_7 ();
 sg13g2_decap_8 FILLER_6_14 ();
 sg13g2_decap_8 FILLER_6_21 ();
 sg13g2_decap_8 FILLER_6_28 ();
 sg13g2_decap_8 FILLER_6_35 ();
 sg13g2_decap_8 FILLER_6_42 ();
 sg13g2_decap_8 FILLER_6_49 ();
 sg13g2_decap_8 FILLER_6_56 ();
 sg13g2_decap_4 FILLER_6_63 ();
 sg13g2_fill_1 FILLER_6_67 ();
 sg13g2_decap_8 FILLER_6_79 ();
 sg13g2_decap_8 FILLER_6_86 ();
 sg13g2_decap_8 FILLER_6_93 ();
 sg13g2_decap_8 FILLER_6_100 ();
 sg13g2_decap_8 FILLER_6_107 ();
 sg13g2_decap_8 FILLER_6_114 ();
 sg13g2_fill_2 FILLER_6_121 ();
 sg13g2_fill_1 FILLER_6_131 ();
 sg13g2_fill_1 FILLER_6_140 ();
 sg13g2_fill_1 FILLER_6_146 ();
 sg13g2_fill_1 FILLER_6_152 ();
 sg13g2_fill_2 FILLER_6_171 ();
 sg13g2_fill_2 FILLER_6_259 ();
 sg13g2_fill_2 FILLER_6_286 ();
 sg13g2_fill_2 FILLER_6_306 ();
 sg13g2_fill_1 FILLER_6_362 ();
 sg13g2_decap_8 FILLER_6_366 ();
 sg13g2_decap_8 FILLER_6_373 ();
 sg13g2_decap_8 FILLER_6_380 ();
 sg13g2_decap_8 FILLER_6_387 ();
 sg13g2_decap_8 FILLER_6_394 ();
 sg13g2_decap_8 FILLER_6_401 ();
 sg13g2_decap_8 FILLER_6_408 ();
 sg13g2_decap_8 FILLER_6_415 ();
 sg13g2_decap_8 FILLER_6_422 ();
 sg13g2_fill_1 FILLER_6_429 ();
 sg13g2_decap_8 FILLER_7_0 ();
 sg13g2_decap_8 FILLER_7_7 ();
 sg13g2_decap_8 FILLER_7_14 ();
 sg13g2_decap_8 FILLER_7_21 ();
 sg13g2_decap_8 FILLER_7_28 ();
 sg13g2_decap_8 FILLER_7_35 ();
 sg13g2_decap_8 FILLER_7_42 ();
 sg13g2_decap_4 FILLER_7_49 ();
 sg13g2_fill_2 FILLER_7_92 ();
 sg13g2_fill_1 FILLER_7_94 ();
 sg13g2_decap_4 FILLER_7_112 ();
 sg13g2_fill_1 FILLER_7_116 ();
 sg13g2_fill_2 FILLER_7_122 ();
 sg13g2_fill_1 FILLER_7_124 ();
 sg13g2_fill_2 FILLER_7_134 ();
 sg13g2_fill_1 FILLER_7_220 ();
 sg13g2_fill_2 FILLER_7_255 ();
 sg13g2_decap_8 FILLER_7_373 ();
 sg13g2_decap_8 FILLER_7_380 ();
 sg13g2_decap_8 FILLER_7_387 ();
 sg13g2_decap_8 FILLER_7_394 ();
 sg13g2_decap_8 FILLER_7_401 ();
 sg13g2_decap_8 FILLER_7_408 ();
 sg13g2_decap_8 FILLER_7_415 ();
 sg13g2_decap_8 FILLER_7_422 ();
 sg13g2_fill_1 FILLER_7_429 ();
 sg13g2_decap_8 FILLER_8_0 ();
 sg13g2_decap_8 FILLER_8_7 ();
 sg13g2_decap_8 FILLER_8_14 ();
 sg13g2_decap_8 FILLER_8_21 ();
 sg13g2_decap_8 FILLER_8_28 ();
 sg13g2_decap_8 FILLER_8_35 ();
 sg13g2_decap_8 FILLER_8_42 ();
 sg13g2_fill_2 FILLER_8_49 ();
 sg13g2_fill_2 FILLER_8_165 ();
 sg13g2_fill_2 FILLER_8_258 ();
 sg13g2_fill_1 FILLER_8_291 ();
 sg13g2_fill_1 FILLER_8_319 ();
 sg13g2_fill_1 FILLER_8_324 ();
 sg13g2_fill_1 FILLER_8_351 ();
 sg13g2_fill_1 FILLER_8_357 ();
 sg13g2_decap_8 FILLER_8_377 ();
 sg13g2_decap_8 FILLER_8_384 ();
 sg13g2_decap_8 FILLER_8_391 ();
 sg13g2_decap_8 FILLER_8_398 ();
 sg13g2_decap_8 FILLER_8_405 ();
 sg13g2_decap_8 FILLER_8_412 ();
 sg13g2_decap_8 FILLER_8_419 ();
 sg13g2_decap_4 FILLER_8_426 ();
 sg13g2_decap_8 FILLER_9_0 ();
 sg13g2_decap_8 FILLER_9_7 ();
 sg13g2_decap_8 FILLER_9_14 ();
 sg13g2_decap_8 FILLER_9_21 ();
 sg13g2_decap_4 FILLER_9_31 ();
 sg13g2_fill_1 FILLER_9_107 ();
 sg13g2_fill_1 FILLER_9_127 ();
 sg13g2_fill_1 FILLER_9_136 ();
 sg13g2_fill_2 FILLER_9_141 ();
 sg13g2_fill_2 FILLER_9_151 ();
 sg13g2_fill_2 FILLER_9_161 ();
 sg13g2_fill_1 FILLER_9_184 ();
 sg13g2_fill_1 FILLER_9_198 ();
 sg13g2_fill_1 FILLER_9_249 ();
 sg13g2_fill_1 FILLER_9_301 ();
 sg13g2_fill_1 FILLER_9_307 ();
 sg13g2_decap_8 FILLER_9_384 ();
 sg13g2_decap_8 FILLER_9_391 ();
 sg13g2_decap_8 FILLER_9_398 ();
 sg13g2_decap_8 FILLER_9_405 ();
 sg13g2_decap_8 FILLER_9_412 ();
 sg13g2_decap_8 FILLER_9_419 ();
 sg13g2_decap_4 FILLER_9_426 ();
 sg13g2_decap_8 FILLER_10_0 ();
 sg13g2_decap_8 FILLER_10_7 ();
 sg13g2_decap_8 FILLER_10_14 ();
 sg13g2_decap_8 FILLER_10_21 ();
 sg13g2_fill_2 FILLER_10_28 ();
 sg13g2_fill_1 FILLER_10_30 ();
 sg13g2_fill_1 FILLER_10_40 ();
 sg13g2_fill_1 FILLER_10_45 ();
 sg13g2_fill_1 FILLER_10_54 ();
 sg13g2_fill_1 FILLER_10_62 ();
 sg13g2_fill_1 FILLER_10_75 ();
 sg13g2_fill_1 FILLER_10_86 ();
 sg13g2_fill_1 FILLER_10_95 ();
 sg13g2_fill_1 FILLER_10_100 ();
 sg13g2_fill_1 FILLER_10_139 ();
 sg13g2_fill_1 FILLER_10_153 ();
 sg13g2_fill_1 FILLER_10_159 ();
 sg13g2_fill_1 FILLER_10_165 ();
 sg13g2_fill_2 FILLER_10_171 ();
 sg13g2_fill_1 FILLER_10_203 ();
 sg13g2_fill_1 FILLER_10_220 ();
 sg13g2_fill_2 FILLER_10_229 ();
 sg13g2_fill_1 FILLER_10_324 ();
 sg13g2_fill_1 FILLER_10_359 ();
 sg13g2_decap_8 FILLER_10_372 ();
 sg13g2_decap_8 FILLER_10_379 ();
 sg13g2_decap_8 FILLER_10_386 ();
 sg13g2_decap_8 FILLER_10_393 ();
 sg13g2_decap_8 FILLER_10_400 ();
 sg13g2_decap_8 FILLER_10_407 ();
 sg13g2_decap_8 FILLER_10_414 ();
 sg13g2_decap_8 FILLER_10_421 ();
 sg13g2_fill_2 FILLER_10_428 ();
 sg13g2_decap_8 FILLER_11_0 ();
 sg13g2_decap_8 FILLER_11_7 ();
 sg13g2_decap_8 FILLER_11_14 ();
 sg13g2_decap_8 FILLER_11_21 ();
 sg13g2_fill_2 FILLER_11_28 ();
 sg13g2_fill_1 FILLER_11_30 ();
 sg13g2_fill_1 FILLER_11_38 ();
 sg13g2_fill_1 FILLER_11_69 ();
 sg13g2_fill_1 FILLER_11_112 ();
 sg13g2_fill_1 FILLER_11_118 ();
 sg13g2_fill_1 FILLER_11_129 ();
 sg13g2_fill_2 FILLER_11_156 ();
 sg13g2_fill_2 FILLER_11_162 ();
 sg13g2_fill_1 FILLER_11_198 ();
 sg13g2_fill_2 FILLER_11_264 ();
 sg13g2_fill_1 FILLER_11_279 ();
 sg13g2_fill_1 FILLER_11_332 ();
 sg13g2_fill_2 FILLER_11_341 ();
 sg13g2_fill_1 FILLER_11_348 ();
 sg13g2_decap_8 FILLER_11_379 ();
 sg13g2_decap_8 FILLER_11_386 ();
 sg13g2_decap_8 FILLER_11_393 ();
 sg13g2_decap_8 FILLER_11_400 ();
 sg13g2_decap_8 FILLER_11_407 ();
 sg13g2_decap_8 FILLER_11_414 ();
 sg13g2_decap_8 FILLER_11_421 ();
 sg13g2_fill_2 FILLER_11_428 ();
 sg13g2_decap_8 FILLER_12_0 ();
 sg13g2_decap_8 FILLER_12_7 ();
 sg13g2_decap_8 FILLER_12_14 ();
 sg13g2_decap_8 FILLER_12_21 ();
 sg13g2_fill_1 FILLER_12_28 ();
 sg13g2_fill_1 FILLER_12_37 ();
 sg13g2_fill_1 FILLER_12_61 ();
 sg13g2_fill_2 FILLER_12_66 ();
 sg13g2_fill_1 FILLER_12_80 ();
 sg13g2_fill_1 FILLER_12_89 ();
 sg13g2_fill_1 FILLER_12_94 ();
 sg13g2_fill_1 FILLER_12_99 ();
 sg13g2_fill_2 FILLER_12_130 ();
 sg13g2_fill_2 FILLER_12_143 ();
 sg13g2_fill_2 FILLER_12_149 ();
 sg13g2_fill_1 FILLER_12_165 ();
 sg13g2_fill_1 FILLER_12_196 ();
 sg13g2_fill_1 FILLER_12_204 ();
 sg13g2_fill_1 FILLER_12_214 ();
 sg13g2_fill_1 FILLER_12_220 ();
 sg13g2_fill_1 FILLER_12_283 ();
 sg13g2_fill_1 FILLER_12_321 ();
 sg13g2_fill_1 FILLER_12_327 ();
 sg13g2_fill_1 FILLER_12_363 ();
 sg13g2_decap_8 FILLER_12_376 ();
 sg13g2_decap_8 FILLER_12_383 ();
 sg13g2_decap_8 FILLER_12_390 ();
 sg13g2_decap_8 FILLER_12_397 ();
 sg13g2_decap_8 FILLER_12_404 ();
 sg13g2_decap_8 FILLER_12_411 ();
 sg13g2_decap_8 FILLER_12_418 ();
 sg13g2_decap_4 FILLER_12_425 ();
 sg13g2_fill_1 FILLER_12_429 ();
 sg13g2_decap_8 FILLER_13_0 ();
 sg13g2_decap_8 FILLER_13_7 ();
 sg13g2_decap_8 FILLER_13_14 ();
 sg13g2_decap_8 FILLER_13_21 ();
 sg13g2_fill_1 FILLER_13_28 ();
 sg13g2_fill_1 FILLER_13_49 ();
 sg13g2_fill_2 FILLER_13_67 ();
 sg13g2_fill_1 FILLER_13_76 ();
 sg13g2_fill_1 FILLER_13_132 ();
 sg13g2_fill_1 FILLER_13_141 ();
 sg13g2_fill_1 FILLER_13_198 ();
 sg13g2_fill_2 FILLER_13_207 ();
 sg13g2_fill_1 FILLER_13_246 ();
 sg13g2_fill_2 FILLER_13_275 ();
 sg13g2_fill_2 FILLER_13_306 ();
 sg13g2_fill_1 FILLER_13_316 ();
 sg13g2_fill_1 FILLER_13_343 ();
 sg13g2_fill_1 FILLER_13_352 ();
 sg13g2_fill_2 FILLER_13_380 ();
 sg13g2_decap_8 FILLER_13_385 ();
 sg13g2_decap_8 FILLER_13_392 ();
 sg13g2_decap_8 FILLER_13_399 ();
 sg13g2_decap_8 FILLER_13_406 ();
 sg13g2_decap_8 FILLER_13_413 ();
 sg13g2_decap_8 FILLER_13_420 ();
 sg13g2_fill_2 FILLER_13_427 ();
 sg13g2_fill_1 FILLER_13_429 ();
 sg13g2_decap_8 FILLER_14_0 ();
 sg13g2_decap_8 FILLER_14_7 ();
 sg13g2_fill_2 FILLER_14_14 ();
 sg13g2_fill_1 FILLER_14_16 ();
 sg13g2_decap_4 FILLER_14_22 ();
 sg13g2_fill_2 FILLER_14_30 ();
 sg13g2_fill_2 FILLER_14_46 ();
 sg13g2_fill_2 FILLER_14_93 ();
 sg13g2_fill_2 FILLER_14_103 ();
 sg13g2_fill_2 FILLER_14_118 ();
 sg13g2_fill_1 FILLER_14_159 ();
 sg13g2_fill_1 FILLER_14_167 ();
 sg13g2_fill_1 FILLER_14_188 ();
 sg13g2_fill_2 FILLER_14_249 ();
 sg13g2_fill_1 FILLER_14_303 ();
 sg13g2_decap_8 FILLER_14_387 ();
 sg13g2_decap_8 FILLER_14_394 ();
 sg13g2_decap_8 FILLER_14_401 ();
 sg13g2_decap_8 FILLER_14_408 ();
 sg13g2_decap_8 FILLER_14_415 ();
 sg13g2_decap_8 FILLER_14_422 ();
 sg13g2_fill_1 FILLER_14_429 ();
 sg13g2_decap_8 FILLER_15_0 ();
 sg13g2_decap_8 FILLER_15_7 ();
 sg13g2_decap_4 FILLER_15_14 ();
 sg13g2_fill_1 FILLER_15_18 ();
 sg13g2_fill_2 FILLER_15_132 ();
 sg13g2_fill_1 FILLER_15_146 ();
 sg13g2_fill_1 FILLER_15_170 ();
 sg13g2_fill_2 FILLER_15_176 ();
 sg13g2_fill_1 FILLER_15_203 ();
 sg13g2_fill_2 FILLER_15_227 ();
 sg13g2_fill_1 FILLER_15_237 ();
 sg13g2_fill_1 FILLER_15_246 ();
 sg13g2_fill_1 FILLER_15_291 ();
 sg13g2_fill_1 FILLER_15_299 ();
 sg13g2_fill_2 FILLER_15_318 ();
 sg13g2_fill_1 FILLER_15_350 ();
 sg13g2_fill_1 FILLER_15_371 ();
 sg13g2_decap_8 FILLER_15_377 ();
 sg13g2_decap_8 FILLER_15_384 ();
 sg13g2_decap_8 FILLER_15_391 ();
 sg13g2_decap_8 FILLER_15_398 ();
 sg13g2_decap_8 FILLER_15_405 ();
 sg13g2_decap_8 FILLER_15_412 ();
 sg13g2_decap_8 FILLER_15_419 ();
 sg13g2_decap_4 FILLER_15_426 ();
 sg13g2_decap_8 FILLER_16_0 ();
 sg13g2_decap_8 FILLER_16_7 ();
 sg13g2_decap_8 FILLER_16_14 ();
 sg13g2_decap_4 FILLER_16_21 ();
 sg13g2_fill_2 FILLER_16_25 ();
 sg13g2_fill_1 FILLER_16_52 ();
 sg13g2_fill_1 FILLER_16_75 ();
 sg13g2_fill_1 FILLER_16_80 ();
 sg13g2_fill_1 FILLER_16_86 ();
 sg13g2_fill_2 FILLER_16_96 ();
 sg13g2_fill_1 FILLER_16_129 ();
 sg13g2_fill_1 FILLER_16_142 ();
 sg13g2_fill_1 FILLER_16_155 ();
 sg13g2_fill_2 FILLER_16_199 ();
 sg13g2_fill_1 FILLER_16_209 ();
 sg13g2_fill_2 FILLER_16_215 ();
 sg13g2_fill_1 FILLER_16_301 ();
 sg13g2_fill_2 FILLER_16_311 ();
 sg13g2_decap_8 FILLER_16_388 ();
 sg13g2_decap_8 FILLER_16_395 ();
 sg13g2_decap_8 FILLER_16_402 ();
 sg13g2_decap_8 FILLER_16_409 ();
 sg13g2_decap_8 FILLER_16_416 ();
 sg13g2_decap_8 FILLER_16_423 ();
 sg13g2_decap_8 FILLER_17_0 ();
 sg13g2_decap_8 FILLER_17_7 ();
 sg13g2_decap_4 FILLER_17_14 ();
 sg13g2_fill_1 FILLER_17_122 ();
 sg13g2_fill_2 FILLER_17_163 ();
 sg13g2_fill_1 FILLER_17_169 ();
 sg13g2_fill_1 FILLER_17_183 ();
 sg13g2_fill_2 FILLER_17_198 ();
 sg13g2_fill_2 FILLER_17_226 ();
 sg13g2_fill_1 FILLER_17_244 ();
 sg13g2_fill_1 FILLER_17_249 ();
 sg13g2_fill_1 FILLER_17_258 ();
 sg13g2_fill_2 FILLER_17_263 ();
 sg13g2_fill_1 FILLER_17_283 ();
 sg13g2_fill_1 FILLER_17_309 ();
 sg13g2_fill_1 FILLER_17_355 ();
 sg13g2_decap_8 FILLER_17_391 ();
 sg13g2_decap_8 FILLER_17_398 ();
 sg13g2_decap_8 FILLER_17_405 ();
 sg13g2_decap_8 FILLER_17_412 ();
 sg13g2_decap_8 FILLER_17_419 ();
 sg13g2_decap_4 FILLER_17_426 ();
 sg13g2_decap_4 FILLER_18_3 ();
 sg13g2_fill_2 FILLER_18_10 ();
 sg13g2_fill_1 FILLER_18_21 ();
 sg13g2_fill_1 FILLER_18_52 ();
 sg13g2_fill_1 FILLER_18_61 ();
 sg13g2_fill_1 FILLER_18_82 ();
 sg13g2_fill_1 FILLER_18_96 ();
 sg13g2_fill_2 FILLER_18_132 ();
 sg13g2_fill_1 FILLER_18_178 ();
 sg13g2_fill_1 FILLER_18_191 ();
 sg13g2_fill_1 FILLER_18_204 ();
 sg13g2_fill_2 FILLER_18_276 ();
 sg13g2_fill_1 FILLER_18_304 ();
 sg13g2_fill_1 FILLER_18_335 ();
 sg13g2_fill_1 FILLER_18_344 ();
 sg13g2_fill_1 FILLER_18_355 ();
 sg13g2_decap_8 FILLER_18_394 ();
 sg13g2_decap_8 FILLER_18_401 ();
 sg13g2_decap_8 FILLER_18_408 ();
 sg13g2_decap_8 FILLER_18_415 ();
 sg13g2_decap_8 FILLER_18_422 ();
 sg13g2_fill_1 FILLER_18_429 ();
 sg13g2_fill_2 FILLER_19_8 ();
 sg13g2_fill_1 FILLER_19_14 ();
 sg13g2_fill_1 FILLER_19_25 ();
 sg13g2_fill_2 FILLER_19_49 ();
 sg13g2_fill_1 FILLER_19_59 ();
 sg13g2_fill_1 FILLER_19_72 ();
 sg13g2_fill_2 FILLER_19_81 ();
 sg13g2_fill_1 FILLER_19_87 ();
 sg13g2_fill_1 FILLER_19_93 ();
 sg13g2_fill_1 FILLER_19_104 ();
 sg13g2_fill_1 FILLER_19_126 ();
 sg13g2_fill_1 FILLER_19_168 ();
 sg13g2_fill_1 FILLER_19_189 ();
 sg13g2_fill_1 FILLER_19_236 ();
 sg13g2_fill_2 FILLER_19_241 ();
 sg13g2_fill_1 FILLER_19_278 ();
 sg13g2_fill_2 FILLER_19_283 ();
 sg13g2_fill_1 FILLER_19_299 ();
 sg13g2_fill_1 FILLER_19_321 ();
 sg13g2_fill_1 FILLER_19_327 ();
 sg13g2_fill_1 FILLER_19_333 ();
 sg13g2_fill_2 FILLER_19_351 ();
 sg13g2_decap_8 FILLER_19_396 ();
 sg13g2_decap_8 FILLER_19_403 ();
 sg13g2_decap_8 FILLER_19_410 ();
 sg13g2_decap_8 FILLER_19_417 ();
 sg13g2_decap_4 FILLER_19_424 ();
 sg13g2_fill_2 FILLER_19_428 ();
 sg13g2_fill_2 FILLER_20_0 ();
 sg13g2_fill_2 FILLER_20_14 ();
 sg13g2_fill_1 FILLER_20_30 ();
 sg13g2_fill_1 FILLER_20_90 ();
 sg13g2_fill_1 FILLER_20_95 ();
 sg13g2_fill_2 FILLER_20_103 ();
 sg13g2_fill_1 FILLER_20_127 ();
 sg13g2_fill_1 FILLER_20_133 ();
 sg13g2_fill_1 FILLER_20_177 ();
 sg13g2_fill_1 FILLER_20_257 ();
 sg13g2_fill_1 FILLER_20_262 ();
 sg13g2_fill_2 FILLER_20_270 ();
 sg13g2_fill_1 FILLER_20_277 ();
 sg13g2_fill_2 FILLER_20_316 ();
 sg13g2_fill_1 FILLER_20_332 ();
 sg13g2_fill_1 FILLER_20_371 ();
 sg13g2_decap_8 FILLER_20_403 ();
 sg13g2_decap_8 FILLER_20_410 ();
 sg13g2_decap_8 FILLER_20_417 ();
 sg13g2_decap_4 FILLER_20_424 ();
 sg13g2_fill_2 FILLER_20_428 ();
 sg13g2_fill_2 FILLER_21_31 ();
 sg13g2_fill_1 FILLER_21_57 ();
 sg13g2_fill_1 FILLER_21_187 ();
 sg13g2_fill_2 FILLER_21_221 ();
 sg13g2_fill_1 FILLER_21_223 ();
 sg13g2_fill_1 FILLER_21_228 ();
 sg13g2_fill_2 FILLER_21_252 ();
 sg13g2_fill_2 FILLER_21_263 ();
 sg13g2_fill_1 FILLER_21_273 ();
 sg13g2_fill_1 FILLER_21_294 ();
 sg13g2_fill_2 FILLER_21_307 ();
 sg13g2_fill_1 FILLER_21_369 ();
 sg13g2_decap_8 FILLER_21_400 ();
 sg13g2_decap_8 FILLER_21_407 ();
 sg13g2_decap_8 FILLER_21_414 ();
 sg13g2_decap_8 FILLER_21_421 ();
 sg13g2_fill_2 FILLER_21_428 ();
 sg13g2_fill_2 FILLER_22_9 ();
 sg13g2_fill_1 FILLER_22_19 ();
 sg13g2_fill_1 FILLER_22_24 ();
 sg13g2_fill_2 FILLER_22_77 ();
 sg13g2_fill_1 FILLER_22_84 ();
 sg13g2_fill_1 FILLER_22_143 ();
 sg13g2_fill_1 FILLER_22_159 ();
 sg13g2_fill_1 FILLER_22_173 ();
 sg13g2_fill_1 FILLER_22_183 ();
 sg13g2_fill_1 FILLER_22_192 ();
 sg13g2_fill_1 FILLER_22_201 ();
 sg13g2_fill_1 FILLER_22_211 ();
 sg13g2_fill_2 FILLER_22_252 ();
 sg13g2_fill_1 FILLER_22_297 ();
 sg13g2_fill_1 FILLER_22_303 ();
 sg13g2_fill_1 FILLER_22_320 ();
 sg13g2_fill_1 FILLER_22_361 ();
 sg13g2_fill_2 FILLER_22_398 ();
 sg13g2_decap_8 FILLER_22_407 ();
 sg13g2_decap_8 FILLER_22_414 ();
 sg13g2_decap_8 FILLER_22_421 ();
 sg13g2_fill_2 FILLER_22_428 ();
 sg13g2_fill_1 FILLER_23_39 ();
 sg13g2_fill_1 FILLER_23_48 ();
 sg13g2_fill_1 FILLER_23_59 ();
 sg13g2_fill_1 FILLER_23_91 ();
 sg13g2_fill_1 FILLER_23_109 ();
 sg13g2_fill_2 FILLER_23_184 ();
 sg13g2_fill_1 FILLER_23_211 ();
 sg13g2_fill_2 FILLER_23_233 ();
 sg13g2_fill_2 FILLER_23_259 ();
 sg13g2_fill_1 FILLER_23_309 ();
 sg13g2_fill_1 FILLER_23_315 ();
 sg13g2_fill_2 FILLER_23_340 ();
 sg13g2_fill_2 FILLER_23_365 ();
 sg13g2_fill_1 FILLER_23_371 ();
 sg13g2_fill_1 FILLER_23_376 ();
 sg13g2_decap_8 FILLER_23_406 ();
 sg13g2_decap_8 FILLER_23_413 ();
 sg13g2_decap_8 FILLER_23_420 ();
 sg13g2_fill_2 FILLER_23_427 ();
 sg13g2_fill_1 FILLER_23_429 ();
 sg13g2_fill_1 FILLER_24_25 ();
 sg13g2_fill_1 FILLER_24_56 ();
 sg13g2_fill_2 FILLER_24_69 ();
 sg13g2_fill_2 FILLER_24_101 ();
 sg13g2_fill_2 FILLER_24_111 ();
 sg13g2_fill_1 FILLER_24_117 ();
 sg13g2_fill_2 FILLER_24_126 ();
 sg13g2_fill_1 FILLER_24_154 ();
 sg13g2_fill_1 FILLER_24_159 ();
 sg13g2_fill_1 FILLER_24_186 ();
 sg13g2_fill_1 FILLER_24_235 ();
 sg13g2_fill_1 FILLER_24_288 ();
 sg13g2_fill_2 FILLER_24_340 ();
 sg13g2_fill_1 FILLER_24_347 ();
 sg13g2_fill_2 FILLER_24_368 ();
 sg13g2_decap_8 FILLER_24_404 ();
 sg13g2_decap_8 FILLER_24_411 ();
 sg13g2_decap_8 FILLER_24_418 ();
 sg13g2_decap_4 FILLER_24_425 ();
 sg13g2_fill_1 FILLER_24_429 ();
 sg13g2_fill_1 FILLER_25_10 ();
 sg13g2_fill_2 FILLER_25_43 ();
 sg13g2_fill_1 FILLER_25_76 ();
 sg13g2_fill_1 FILLER_25_117 ();
 sg13g2_fill_1 FILLER_25_144 ();
 sg13g2_fill_1 FILLER_25_150 ();
 sg13g2_fill_1 FILLER_25_183 ();
 sg13g2_fill_1 FILLER_25_213 ();
 sg13g2_fill_1 FILLER_25_225 ();
 sg13g2_fill_1 FILLER_25_230 ();
 sg13g2_fill_1 FILLER_25_235 ();
 sg13g2_fill_1 FILLER_25_244 ();
 sg13g2_fill_1 FILLER_25_249 ();
 sg13g2_fill_1 FILLER_25_253 ();
 sg13g2_fill_1 FILLER_25_259 ();
 sg13g2_fill_1 FILLER_25_282 ();
 sg13g2_fill_2 FILLER_25_315 ();
 sg13g2_fill_1 FILLER_25_317 ();
 sg13g2_decap_8 FILLER_25_411 ();
 sg13g2_decap_8 FILLER_25_418 ();
 sg13g2_decap_4 FILLER_25_425 ();
 sg13g2_fill_1 FILLER_25_429 ();
 sg13g2_fill_1 FILLER_26_34 ();
 sg13g2_fill_2 FILLER_26_66 ();
 sg13g2_fill_2 FILLER_26_132 ();
 sg13g2_fill_1 FILLER_26_219 ();
 sg13g2_decap_4 FILLER_26_234 ();
 sg13g2_fill_1 FILLER_26_238 ();
 sg13g2_fill_1 FILLER_26_245 ();
 sg13g2_fill_1 FILLER_26_259 ();
 sg13g2_decap_4 FILLER_26_264 ();
 sg13g2_fill_2 FILLER_26_268 ();
 sg13g2_fill_1 FILLER_26_277 ();
 sg13g2_fill_2 FILLER_26_301 ();
 sg13g2_fill_2 FILLER_26_332 ();
 sg13g2_decap_8 FILLER_26_406 ();
 sg13g2_decap_8 FILLER_26_413 ();
 sg13g2_decap_8 FILLER_26_420 ();
 sg13g2_fill_2 FILLER_26_427 ();
 sg13g2_fill_1 FILLER_26_429 ();
 sg13g2_fill_1 FILLER_27_10 ();
 sg13g2_fill_1 FILLER_27_29 ();
 sg13g2_fill_1 FILLER_27_38 ();
 sg13g2_fill_1 FILLER_27_96 ();
 sg13g2_fill_2 FILLER_27_100 ();
 sg13g2_fill_1 FILLER_27_102 ();
 sg13g2_fill_1 FILLER_27_118 ();
 sg13g2_fill_2 FILLER_27_123 ();
 sg13g2_fill_1 FILLER_27_125 ();
 sg13g2_fill_2 FILLER_27_152 ();
 sg13g2_fill_1 FILLER_27_200 ();
 sg13g2_fill_2 FILLER_27_223 ();
 sg13g2_fill_1 FILLER_27_225 ();
 sg13g2_fill_1 FILLER_27_244 ();
 sg13g2_fill_1 FILLER_27_304 ();
 sg13g2_fill_1 FILLER_27_318 ();
 sg13g2_fill_1 FILLER_27_329 ();
 sg13g2_fill_2 FILLER_27_343 ();
 sg13g2_fill_2 FILLER_27_366 ();
 sg13g2_fill_2 FILLER_27_399 ();
 sg13g2_fill_1 FILLER_27_409 ();
 sg13g2_decap_8 FILLER_27_418 ();
 sg13g2_decap_4 FILLER_27_425 ();
 sg13g2_fill_1 FILLER_27_429 ();
 sg13g2_fill_2 FILLER_28_15 ();
 sg13g2_fill_2 FILLER_28_22 ();
 sg13g2_fill_2 FILLER_28_47 ();
 sg13g2_fill_2 FILLER_28_56 ();
 sg13g2_fill_1 FILLER_28_65 ();
 sg13g2_fill_1 FILLER_28_94 ();
 sg13g2_fill_1 FILLER_28_129 ();
 sg13g2_fill_2 FILLER_28_175 ();
 sg13g2_fill_1 FILLER_28_232 ();
 sg13g2_fill_1 FILLER_28_241 ();
 sg13g2_fill_1 FILLER_28_267 ();
 sg13g2_fill_2 FILLER_28_294 ();
 sg13g2_fill_1 FILLER_28_296 ();
 sg13g2_fill_1 FILLER_28_343 ();
 sg13g2_fill_1 FILLER_28_349 ();
 sg13g2_fill_1 FILLER_28_367 ();
 sg13g2_fill_2 FILLER_28_412 ();
 sg13g2_fill_1 FILLER_28_414 ();
 sg13g2_decap_8 FILLER_28_419 ();
 sg13g2_decap_4 FILLER_28_426 ();
 sg13g2_fill_1 FILLER_29_52 ();
 sg13g2_fill_1 FILLER_29_57 ();
 sg13g2_fill_1 FILLER_29_124 ();
 sg13g2_fill_1 FILLER_29_273 ();
 sg13g2_fill_1 FILLER_29_306 ();
 sg13g2_fill_1 FILLER_29_370 ();
 sg13g2_fill_1 FILLER_29_403 ();
 sg13g2_decap_8 FILLER_29_419 ();
 sg13g2_decap_4 FILLER_29_426 ();
 sg13g2_fill_2 FILLER_30_0 ();
 sg13g2_fill_1 FILLER_30_41 ();
 sg13g2_fill_1 FILLER_30_77 ();
 sg13g2_fill_2 FILLER_30_136 ();
 sg13g2_fill_2 FILLER_30_164 ();
 sg13g2_fill_1 FILLER_30_183 ();
 sg13g2_fill_2 FILLER_30_227 ();
 sg13g2_fill_2 FILLER_30_258 ();
 sg13g2_fill_1 FILLER_30_260 ();
 sg13g2_fill_1 FILLER_30_295 ();
 sg13g2_fill_1 FILLER_30_306 ();
 sg13g2_fill_2 FILLER_30_331 ();
 sg13g2_fill_1 FILLER_30_362 ();
 sg13g2_fill_1 FILLER_30_418 ();
 sg13g2_decap_4 FILLER_30_424 ();
 sg13g2_fill_2 FILLER_30_428 ();
 sg13g2_fill_1 FILLER_31_0 ();
 sg13g2_fill_2 FILLER_31_50 ();
 sg13g2_fill_1 FILLER_31_59 ();
 sg13g2_fill_1 FILLER_31_64 ();
 sg13g2_fill_1 FILLER_31_80 ();
 sg13g2_fill_2 FILLER_31_85 ();
 sg13g2_fill_1 FILLER_31_91 ();
 sg13g2_fill_2 FILLER_31_123 ();
 sg13g2_fill_1 FILLER_31_128 ();
 sg13g2_fill_1 FILLER_31_186 ();
 sg13g2_fill_1 FILLER_31_199 ();
 sg13g2_fill_1 FILLER_31_204 ();
 sg13g2_fill_2 FILLER_31_209 ();
 sg13g2_fill_1 FILLER_31_216 ();
 sg13g2_fill_1 FILLER_31_267 ();
 sg13g2_fill_1 FILLER_31_272 ();
 sg13g2_fill_1 FILLER_31_357 ();
 sg13g2_fill_1 FILLER_31_391 ();
 sg13g2_fill_2 FILLER_31_400 ();
 sg13g2_fill_1 FILLER_31_410 ();
 sg13g2_decap_8 FILLER_31_420 ();
 sg13g2_fill_2 FILLER_31_427 ();
 sg13g2_fill_1 FILLER_31_429 ();
 sg13g2_fill_1 FILLER_32_34 ();
 sg13g2_fill_1 FILLER_32_50 ();
 sg13g2_fill_1 FILLER_32_77 ();
 sg13g2_fill_1 FILLER_32_98 ();
 sg13g2_fill_2 FILLER_32_148 ();
 sg13g2_fill_1 FILLER_32_162 ();
 sg13g2_fill_1 FILLER_32_171 ();
 sg13g2_fill_1 FILLER_32_180 ();
 sg13g2_fill_2 FILLER_32_207 ();
 sg13g2_fill_1 FILLER_32_209 ();
 sg13g2_fill_1 FILLER_32_218 ();
 sg13g2_fill_1 FILLER_32_223 ();
 sg13g2_fill_1 FILLER_32_228 ();
 sg13g2_fill_1 FILLER_32_233 ();
 sg13g2_fill_2 FILLER_32_239 ();
 sg13g2_fill_1 FILLER_32_245 ();
 sg13g2_fill_1 FILLER_32_259 ();
 sg13g2_fill_2 FILLER_32_265 ();
 sg13g2_fill_1 FILLER_32_340 ();
 sg13g2_decap_4 FILLER_32_360 ();
 sg13g2_fill_2 FILLER_32_369 ();
 sg13g2_fill_2 FILLER_32_412 ();
 sg13g2_fill_1 FILLER_32_414 ();
 sg13g2_decap_8 FILLER_32_423 ();
 sg13g2_fill_1 FILLER_33_64 ();
 sg13g2_fill_1 FILLER_33_91 ();
 sg13g2_fill_1 FILLER_33_125 ();
 sg13g2_fill_1 FILLER_33_185 ();
 sg13g2_fill_2 FILLER_33_237 ();
 sg13g2_fill_1 FILLER_33_247 ();
 sg13g2_fill_1 FILLER_33_251 ();
 sg13g2_fill_1 FILLER_33_256 ();
 sg13g2_fill_2 FILLER_33_362 ();
 sg13g2_fill_2 FILLER_33_393 ();
 sg13g2_fill_2 FILLER_33_409 ();
 sg13g2_decap_4 FILLER_33_426 ();
 sg13g2_fill_2 FILLER_34_0 ();
 sg13g2_fill_2 FILLER_34_22 ();
 sg13g2_fill_1 FILLER_34_54 ();
 sg13g2_fill_2 FILLER_34_73 ();
 sg13g2_fill_2 FILLER_34_79 ();
 sg13g2_fill_2 FILLER_34_88 ();
 sg13g2_fill_2 FILLER_34_154 ();
 sg13g2_fill_1 FILLER_34_165 ();
 sg13g2_fill_1 FILLER_34_181 ();
 sg13g2_fill_1 FILLER_34_199 ();
 sg13g2_fill_1 FILLER_34_205 ();
 sg13g2_fill_1 FILLER_34_210 ();
 sg13g2_fill_1 FILLER_34_216 ();
 sg13g2_fill_2 FILLER_34_279 ();
 sg13g2_fill_2 FILLER_34_290 ();
 sg13g2_fill_2 FILLER_34_334 ();
 sg13g2_fill_2 FILLER_34_343 ();
 sg13g2_fill_2 FILLER_34_411 ();
 sg13g2_fill_1 FILLER_34_421 ();
 sg13g2_fill_2 FILLER_35_42 ();
 sg13g2_fill_1 FILLER_35_70 ();
 sg13g2_fill_1 FILLER_35_109 ();
 sg13g2_fill_1 FILLER_35_138 ();
 sg13g2_fill_1 FILLER_35_157 ();
 sg13g2_fill_2 FILLER_35_187 ();
 sg13g2_fill_2 FILLER_35_211 ();
 sg13g2_fill_2 FILLER_35_243 ();
 sg13g2_fill_1 FILLER_35_249 ();
 sg13g2_fill_2 FILLER_35_254 ();
 sg13g2_fill_1 FILLER_35_260 ();
 sg13g2_fill_1 FILLER_35_265 ();
 sg13g2_fill_1 FILLER_35_270 ();
 sg13g2_fill_1 FILLER_35_275 ();
 sg13g2_fill_1 FILLER_35_280 ();
 sg13g2_fill_2 FILLER_35_311 ();
 sg13g2_fill_1 FILLER_35_321 ();
 sg13g2_fill_2 FILLER_35_359 ();
 sg13g2_fill_1 FILLER_35_429 ();
 sg13g2_fill_2 FILLER_36_0 ();
 sg13g2_fill_1 FILLER_36_21 ();
 sg13g2_fill_1 FILLER_36_70 ();
 sg13g2_fill_1 FILLER_36_118 ();
 sg13g2_fill_1 FILLER_36_208 ();
 sg13g2_fill_1 FILLER_36_218 ();
 sg13g2_fill_1 FILLER_36_223 ();
 sg13g2_fill_1 FILLER_36_231 ();
 sg13g2_fill_2 FILLER_36_236 ();
 sg13g2_fill_1 FILLER_36_246 ();
 sg13g2_fill_2 FILLER_36_277 ();
 sg13g2_fill_1 FILLER_36_279 ();
 sg13g2_fill_1 FILLER_36_290 ();
 sg13g2_fill_1 FILLER_36_324 ();
 sg13g2_fill_2 FILLER_36_328 ();
 sg13g2_fill_1 FILLER_36_382 ();
 sg13g2_fill_2 FILLER_36_387 ();
 sg13g2_fill_1 FILLER_36_397 ();
 sg13g2_fill_2 FILLER_37_0 ();
 sg13g2_fill_2 FILLER_37_75 ();
 sg13g2_fill_1 FILLER_37_84 ();
 sg13g2_fill_1 FILLER_37_90 ();
 sg13g2_fill_1 FILLER_37_99 ();
 sg13g2_fill_2 FILLER_37_113 ();
 sg13g2_fill_1 FILLER_37_146 ();
 sg13g2_fill_2 FILLER_37_179 ();
 sg13g2_fill_1 FILLER_37_211 ();
 sg13g2_decap_4 FILLER_37_265 ();
 sg13g2_fill_1 FILLER_37_269 ();
 sg13g2_fill_1 FILLER_37_274 ();
 sg13g2_fill_2 FILLER_37_287 ();
 sg13g2_fill_1 FILLER_37_309 ();
 sg13g2_fill_1 FILLER_37_338 ();
 sg13g2_fill_1 FILLER_37_343 ();
 sg13g2_fill_1 FILLER_37_374 ();
 sg13g2_fill_1 FILLER_37_379 ();
 sg13g2_fill_2 FILLER_37_385 ();
 sg13g2_fill_1 FILLER_37_406 ();
 sg13g2_fill_1 FILLER_37_417 ();
 sg13g2_fill_2 FILLER_37_428 ();
 sg13g2_fill_1 FILLER_38_0 ();
 sg13g2_fill_1 FILLER_38_9 ();
 sg13g2_fill_1 FILLER_38_20 ();
 sg13g2_fill_1 FILLER_38_26 ();
 sg13g2_fill_1 FILLER_38_37 ();
 sg13g2_fill_1 FILLER_38_103 ();
 sg13g2_fill_1 FILLER_38_198 ();
 sg13g2_fill_1 FILLER_38_217 ();
 sg13g2_fill_1 FILLER_38_223 ();
 sg13g2_fill_1 FILLER_38_244 ();
 sg13g2_fill_2 FILLER_38_296 ();
 sg13g2_fill_1 FILLER_38_316 ();
 sg13g2_fill_1 FILLER_38_321 ();
 sg13g2_fill_2 FILLER_38_356 ();
 sg13g2_decap_4 FILLER_38_363 ();
 sg13g2_fill_1 FILLER_38_367 ();
 sg13g2_decap_4 FILLER_38_424 ();
 sg13g2_fill_2 FILLER_38_428 ();
 sg13g2_fill_2 FILLER_39_0 ();
 sg13g2_fill_2 FILLER_39_24 ();
 sg13g2_fill_1 FILLER_39_136 ();
 sg13g2_fill_2 FILLER_39_193 ();
 sg13g2_fill_1 FILLER_39_209 ();
 sg13g2_fill_1 FILLER_39_219 ();
 sg13g2_fill_1 FILLER_39_237 ();
 sg13g2_fill_1 FILLER_39_248 ();
 sg13g2_fill_1 FILLER_39_257 ();
 sg13g2_fill_1 FILLER_39_274 ();
 sg13g2_fill_2 FILLER_39_280 ();
 sg13g2_fill_2 FILLER_39_289 ();
 sg13g2_fill_2 FILLER_39_299 ();
 sg13g2_fill_1 FILLER_39_301 ();
 sg13g2_fill_1 FILLER_39_341 ();
 sg13g2_fill_1 FILLER_39_345 ();
 sg13g2_fill_1 FILLER_39_350 ();
 sg13g2_fill_1 FILLER_39_368 ();
 sg13g2_fill_1 FILLER_39_374 ();
 sg13g2_fill_1 FILLER_39_416 ();
 sg13g2_fill_2 FILLER_40_22 ();
 sg13g2_fill_1 FILLER_40_39 ();
 sg13g2_fill_1 FILLER_40_44 ();
 sg13g2_fill_1 FILLER_40_71 ();
 sg13g2_fill_1 FILLER_40_76 ();
 sg13g2_decap_4 FILLER_40_98 ();
 sg13g2_fill_2 FILLER_40_102 ();
 sg13g2_fill_1 FILLER_40_116 ();
 sg13g2_fill_2 FILLER_40_128 ();
 sg13g2_fill_1 FILLER_40_130 ();
 sg13g2_decap_4 FILLER_40_139 ();
 sg13g2_fill_1 FILLER_40_151 ();
 sg13g2_fill_1 FILLER_40_157 ();
 sg13g2_fill_1 FILLER_40_163 ();
 sg13g2_fill_1 FILLER_40_189 ();
 sg13g2_fill_2 FILLER_40_207 ();
 sg13g2_fill_1 FILLER_40_302 ();
 sg13g2_fill_1 FILLER_40_307 ();
 sg13g2_fill_1 FILLER_40_331 ();
 sg13g2_fill_2 FILLER_40_359 ();
 sg13g2_fill_1 FILLER_40_361 ();
 sg13g2_decap_4 FILLER_40_370 ();
 sg13g2_fill_2 FILLER_40_379 ();
 sg13g2_fill_1 FILLER_40_381 ();
 sg13g2_fill_2 FILLER_40_397 ();
 sg13g2_fill_1 FILLER_40_399 ();
 sg13g2_fill_2 FILLER_40_408 ();
 sg13g2_fill_1 FILLER_40_410 ();
 sg13g2_fill_2 FILLER_41_59 ();
 sg13g2_fill_1 FILLER_41_65 ();
 sg13g2_fill_1 FILLER_41_122 ();
 sg13g2_fill_1 FILLER_41_128 ();
 sg13g2_fill_1 FILLER_41_132 ();
 sg13g2_fill_1 FILLER_41_145 ();
 sg13g2_fill_2 FILLER_41_154 ();
 sg13g2_fill_1 FILLER_41_156 ();
 sg13g2_fill_2 FILLER_41_169 ();
 sg13g2_fill_1 FILLER_41_171 ();
 sg13g2_fill_1 FILLER_41_205 ();
 sg13g2_fill_2 FILLER_41_210 ();
 sg13g2_fill_1 FILLER_41_234 ();
 sg13g2_fill_1 FILLER_41_261 ();
 sg13g2_fill_1 FILLER_41_292 ();
 sg13g2_fill_1 FILLER_41_306 ();
 sg13g2_fill_1 FILLER_41_327 ();
 sg13g2_fill_1 FILLER_41_332 ();
 sg13g2_decap_4 FILLER_41_342 ();
 sg13g2_fill_2 FILLER_41_346 ();
 sg13g2_decap_4 FILLER_41_352 ();
 sg13g2_fill_2 FILLER_41_356 ();
 sg13g2_fill_1 FILLER_41_387 ();
 sg13g2_fill_2 FILLER_41_396 ();
 sg13g2_fill_2 FILLER_41_406 ();
 sg13g2_fill_1 FILLER_41_408 ();
 sg13g2_fill_1 FILLER_41_414 ();
 sg13g2_fill_2 FILLER_41_419 ();
 sg13g2_fill_1 FILLER_41_429 ();
 sg13g2_fill_1 FILLER_42_38 ();
 sg13g2_fill_1 FILLER_42_119 ();
 sg13g2_fill_1 FILLER_42_124 ();
 sg13g2_fill_1 FILLER_42_136 ();
 sg13g2_fill_2 FILLER_42_206 ();
 sg13g2_fill_1 FILLER_42_208 ();
 sg13g2_fill_1 FILLER_42_261 ();
 sg13g2_fill_2 FILLER_42_266 ();
 sg13g2_fill_2 FILLER_42_344 ();
 sg13g2_decap_4 FILLER_42_384 ();
 sg13g2_decap_4 FILLER_42_396 ();
 sg13g2_fill_1 FILLER_42_400 ();
 sg13g2_fill_1 FILLER_42_429 ();
 sg13g2_fill_1 FILLER_43_0 ();
 sg13g2_fill_2 FILLER_43_29 ();
 sg13g2_fill_1 FILLER_43_75 ();
 sg13g2_fill_1 FILLER_43_80 ();
 sg13g2_fill_1 FILLER_43_107 ();
 sg13g2_fill_2 FILLER_43_117 ();
 sg13g2_fill_1 FILLER_43_119 ();
 sg13g2_fill_1 FILLER_43_127 ();
 sg13g2_fill_1 FILLER_43_132 ();
 sg13g2_fill_1 FILLER_43_143 ();
 sg13g2_fill_2 FILLER_43_156 ();
 sg13g2_fill_1 FILLER_43_158 ();
 sg13g2_fill_1 FILLER_43_163 ();
 sg13g2_fill_1 FILLER_43_172 ();
 sg13g2_fill_2 FILLER_43_210 ();
 sg13g2_decap_4 FILLER_43_221 ();
 sg13g2_fill_2 FILLER_43_225 ();
 sg13g2_fill_1 FILLER_43_230 ();
 sg13g2_decap_8 FILLER_43_234 ();
 sg13g2_fill_1 FILLER_43_241 ();
 sg13g2_fill_1 FILLER_43_287 ();
 sg13g2_fill_1 FILLER_43_309 ();
 sg13g2_fill_2 FILLER_43_345 ();
 sg13g2_decap_8 FILLER_43_351 ();
 sg13g2_fill_1 FILLER_43_358 ();
 sg13g2_fill_1 FILLER_43_368 ();
 sg13g2_decap_4 FILLER_43_377 ();
 sg13g2_fill_2 FILLER_43_420 ();
 sg13g2_fill_1 FILLER_43_422 ();
 sg13g2_fill_2 FILLER_43_428 ();
 sg13g2_decap_4 FILLER_44_33 ();
 sg13g2_fill_1 FILLER_44_69 ();
 sg13g2_fill_1 FILLER_44_88 ();
 sg13g2_fill_2 FILLER_44_100 ();
 sg13g2_fill_1 FILLER_44_102 ();
 sg13g2_fill_1 FILLER_44_107 ();
 sg13g2_fill_2 FILLER_44_124 ();
 sg13g2_fill_1 FILLER_44_129 ();
 sg13g2_fill_1 FILLER_44_138 ();
 sg13g2_fill_1 FILLER_44_184 ();
 sg13g2_fill_1 FILLER_44_193 ();
 sg13g2_fill_1 FILLER_44_198 ();
 sg13g2_fill_2 FILLER_44_203 ();
 sg13g2_decap_4 FILLER_44_209 ();
 sg13g2_fill_1 FILLER_44_213 ();
 sg13g2_decap_4 FILLER_44_222 ();
 sg13g2_fill_1 FILLER_44_226 ();
 sg13g2_fill_2 FILLER_44_255 ();
 sg13g2_fill_1 FILLER_44_262 ();
 sg13g2_fill_2 FILLER_44_272 ();
 sg13g2_fill_1 FILLER_44_283 ();
 sg13g2_fill_1 FILLER_44_324 ();
 sg13g2_fill_2 FILLER_44_338 ();
 sg13g2_fill_1 FILLER_44_340 ();
 sg13g2_decap_4 FILLER_44_348 ();
 sg13g2_fill_2 FILLER_44_365 ();
 sg13g2_fill_1 FILLER_44_367 ();
 sg13g2_fill_2 FILLER_44_403 ();
 sg13g2_fill_2 FILLER_44_408 ();
 sg13g2_fill_1 FILLER_44_414 ();
 sg13g2_fill_2 FILLER_44_428 ();
 sg13g2_fill_1 FILLER_45_66 ();
 sg13g2_fill_1 FILLER_45_74 ();
 sg13g2_fill_1 FILLER_45_79 ();
 sg13g2_fill_1 FILLER_45_87 ();
 sg13g2_fill_2 FILLER_45_102 ();
 sg13g2_fill_2 FILLER_45_119 ();
 sg13g2_fill_1 FILLER_45_134 ();
 sg13g2_fill_1 FILLER_45_140 ();
 sg13g2_fill_1 FILLER_45_146 ();
 sg13g2_fill_1 FILLER_45_151 ();
 sg13g2_fill_2 FILLER_45_160 ();
 sg13g2_fill_2 FILLER_45_170 ();
 sg13g2_fill_2 FILLER_45_252 ();
 sg13g2_fill_1 FILLER_45_257 ();
 sg13g2_fill_1 FILLER_45_262 ();
 sg13g2_fill_1 FILLER_45_271 ();
 sg13g2_fill_1 FILLER_45_287 ();
 sg13g2_fill_1 FILLER_45_293 ();
 sg13g2_fill_1 FILLER_45_299 ();
 sg13g2_fill_1 FILLER_45_318 ();
 sg13g2_decap_4 FILLER_45_329 ();
 sg13g2_fill_1 FILLER_45_349 ();
 sg13g2_fill_1 FILLER_45_360 ();
 sg13g2_fill_1 FILLER_45_365 ();
 sg13g2_fill_1 FILLER_45_378 ();
 sg13g2_fill_1 FILLER_45_383 ();
 sg13g2_fill_1 FILLER_45_389 ();
 sg13g2_fill_1 FILLER_45_406 ();
 sg13g2_fill_1 FILLER_45_411 ();
 sg13g2_fill_2 FILLER_45_416 ();
 sg13g2_fill_1 FILLER_45_423 ();
 sg13g2_fill_2 FILLER_45_428 ();
 sg13g2_fill_1 FILLER_46_33 ();
 sg13g2_fill_1 FILLER_46_98 ();
 sg13g2_fill_2 FILLER_46_129 ();
 sg13g2_fill_1 FILLER_46_135 ();
 sg13g2_fill_1 FILLER_46_144 ();
 sg13g2_fill_2 FILLER_46_168 ();
 sg13g2_fill_2 FILLER_46_178 ();
 sg13g2_fill_1 FILLER_46_222 ();
 sg13g2_fill_1 FILLER_46_239 ();
 sg13g2_fill_2 FILLER_46_281 ();
 sg13g2_fill_1 FILLER_46_283 ();
 sg13g2_fill_2 FILLER_46_314 ();
 sg13g2_fill_1 FILLER_46_338 ();
 sg13g2_fill_1 FILLER_46_359 ();
 sg13g2_fill_1 FILLER_46_363 ();
 sg13g2_fill_1 FILLER_46_369 ();
 sg13g2_fill_2 FILLER_46_427 ();
 sg13g2_fill_1 FILLER_46_429 ();
 sg13g2_fill_1 FILLER_47_33 ();
 sg13g2_fill_2 FILLER_47_43 ();
 sg13g2_fill_1 FILLER_47_73 ();
 sg13g2_fill_1 FILLER_47_87 ();
 sg13g2_fill_1 FILLER_47_104 ();
 sg13g2_fill_2 FILLER_47_127 ();
 sg13g2_fill_1 FILLER_47_129 ();
 sg13g2_fill_2 FILLER_47_133 ();
 sg13g2_fill_1 FILLER_47_135 ();
 sg13g2_fill_2 FILLER_47_165 ();
 sg13g2_fill_1 FILLER_47_249 ();
 sg13g2_fill_2 FILLER_47_256 ();
 sg13g2_fill_1 FILLER_47_262 ();
 sg13g2_fill_1 FILLER_47_270 ();
 sg13g2_fill_1 FILLER_47_309 ();
 sg13g2_fill_2 FILLER_47_314 ();
 sg13g2_fill_1 FILLER_47_343 ();
 sg13g2_decap_4 FILLER_47_353 ();
 sg13g2_fill_2 FILLER_47_357 ();
 sg13g2_fill_1 FILLER_47_363 ();
 sg13g2_fill_1 FILLER_47_372 ();
 sg13g2_fill_1 FILLER_47_391 ();
 sg13g2_fill_1 FILLER_47_424 ();
 sg13g2_fill_1 FILLER_47_429 ();
 sg13g2_fill_2 FILLER_48_15 ();
 sg13g2_fill_1 FILLER_48_38 ();
 sg13g2_fill_1 FILLER_48_87 ();
 sg13g2_fill_1 FILLER_48_92 ();
 sg13g2_fill_1 FILLER_48_97 ();
 sg13g2_fill_1 FILLER_48_161 ();
 sg13g2_fill_1 FILLER_48_188 ();
 sg13g2_fill_1 FILLER_48_198 ();
 sg13g2_fill_2 FILLER_48_203 ();
 sg13g2_fill_1 FILLER_48_210 ();
 sg13g2_fill_1 FILLER_48_216 ();
 sg13g2_fill_2 FILLER_48_222 ();
 sg13g2_fill_1 FILLER_48_228 ();
 sg13g2_fill_1 FILLER_48_232 ();
 sg13g2_fill_1 FILLER_48_251 ();
 sg13g2_fill_1 FILLER_48_257 ();
 sg13g2_fill_1 FILLER_48_266 ();
 sg13g2_fill_1 FILLER_48_273 ();
 sg13g2_fill_1 FILLER_48_282 ();
 sg13g2_fill_2 FILLER_48_287 ();
 sg13g2_fill_1 FILLER_48_292 ();
 sg13g2_fill_1 FILLER_48_298 ();
 sg13g2_fill_1 FILLER_48_304 ();
 sg13g2_fill_1 FILLER_48_310 ();
 sg13g2_fill_2 FILLER_48_366 ();
 sg13g2_decap_4 FILLER_48_389 ();
 sg13g2_fill_1 FILLER_48_393 ();
 sg13g2_fill_1 FILLER_48_421 ();
 sg13g2_fill_1 FILLER_48_426 ();
 sg13g2_fill_1 FILLER_49_30 ();
 sg13g2_fill_2 FILLER_49_47 ();
 sg13g2_fill_1 FILLER_49_67 ();
 sg13g2_fill_1 FILLER_49_72 ();
 sg13g2_fill_1 FILLER_49_124 ();
 sg13g2_fill_2 FILLER_49_148 ();
 sg13g2_fill_1 FILLER_49_163 ();
 sg13g2_fill_2 FILLER_49_168 ();
 sg13g2_fill_2 FILLER_49_173 ();
 sg13g2_fill_2 FILLER_49_206 ();
 sg13g2_fill_2 FILLER_49_228 ();
 sg13g2_fill_2 FILLER_49_262 ();
 sg13g2_fill_1 FILLER_49_268 ();
 sg13g2_fill_2 FILLER_49_273 ();
 sg13g2_fill_1 FILLER_49_284 ();
 sg13g2_fill_1 FILLER_49_297 ();
 sg13g2_fill_1 FILLER_49_326 ();
 sg13g2_fill_1 FILLER_49_356 ();
 sg13g2_decap_4 FILLER_49_369 ();
 sg13g2_fill_1 FILLER_49_377 ();
 sg13g2_fill_1 FILLER_49_383 ();
 sg13g2_fill_1 FILLER_49_392 ();
 sg13g2_fill_2 FILLER_49_406 ();
 sg13g2_fill_1 FILLER_49_408 ();
 sg13g2_fill_2 FILLER_49_428 ();
 sg13g2_fill_1 FILLER_50_5 ();
 sg13g2_fill_1 FILLER_50_10 ();
 sg13g2_fill_1 FILLER_50_33 ();
 sg13g2_fill_1 FILLER_50_43 ();
 sg13g2_fill_1 FILLER_50_110 ();
 sg13g2_fill_1 FILLER_50_131 ();
 sg13g2_fill_1 FILLER_50_136 ();
 sg13g2_fill_1 FILLER_50_145 ();
 sg13g2_fill_1 FILLER_50_178 ();
 sg13g2_fill_2 FILLER_50_271 ();
 sg13g2_fill_1 FILLER_50_295 ();
 sg13g2_fill_1 FILLER_50_309 ();
 sg13g2_fill_1 FILLER_50_318 ();
 sg13g2_fill_1 FILLER_50_328 ();
 sg13g2_fill_1 FILLER_50_334 ();
 sg13g2_fill_2 FILLER_50_339 ();
 sg13g2_fill_1 FILLER_50_350 ();
 sg13g2_fill_1 FILLER_50_359 ();
 sg13g2_fill_1 FILLER_50_364 ();
 sg13g2_fill_2 FILLER_50_371 ();
 sg13g2_fill_2 FILLER_50_385 ();
 sg13g2_fill_1 FILLER_50_399 ();
 sg13g2_fill_1 FILLER_50_405 ();
 sg13g2_fill_2 FILLER_50_427 ();
 sg13g2_fill_1 FILLER_50_429 ();
 sg13g2_fill_2 FILLER_51_138 ();
 sg13g2_fill_1 FILLER_51_171 ();
 sg13g2_decap_4 FILLER_51_176 ();
 sg13g2_fill_1 FILLER_51_194 ();
 sg13g2_fill_1 FILLER_51_203 ();
 sg13g2_fill_1 FILLER_51_268 ();
 sg13g2_fill_1 FILLER_51_273 ();
 sg13g2_fill_1 FILLER_51_278 ();
 sg13g2_fill_2 FILLER_51_292 ();
 sg13g2_fill_1 FILLER_51_310 ();
 sg13g2_fill_1 FILLER_51_315 ();
 sg13g2_fill_1 FILLER_51_321 ();
 sg13g2_fill_1 FILLER_51_326 ();
 sg13g2_fill_2 FILLER_51_335 ();
 sg13g2_fill_1 FILLER_51_337 ();
 sg13g2_fill_1 FILLER_51_364 ();
 sg13g2_fill_1 FILLER_51_429 ();
 sg13g2_fill_2 FILLER_52_12 ();
 sg13g2_fill_1 FILLER_52_19 ();
 sg13g2_fill_1 FILLER_52_48 ();
 sg13g2_fill_2 FILLER_52_71 ();
 sg13g2_fill_1 FILLER_52_78 ();
 sg13g2_fill_1 FILLER_52_84 ();
 sg13g2_fill_1 FILLER_52_89 ();
 sg13g2_fill_1 FILLER_52_98 ();
 sg13g2_fill_1 FILLER_52_113 ();
 sg13g2_fill_2 FILLER_52_131 ();
 sg13g2_fill_1 FILLER_52_133 ();
 sg13g2_fill_1 FILLER_52_150 ();
 sg13g2_fill_1 FILLER_52_157 ();
 sg13g2_fill_1 FILLER_52_162 ();
 sg13g2_fill_1 FILLER_52_168 ();
 sg13g2_fill_2 FILLER_52_195 ();
 sg13g2_fill_1 FILLER_52_225 ();
 sg13g2_fill_1 FILLER_52_231 ();
 sg13g2_fill_1 FILLER_52_237 ();
 sg13g2_fill_2 FILLER_52_246 ();
 sg13g2_fill_2 FILLER_52_253 ();
 sg13g2_fill_2 FILLER_52_273 ();
 sg13g2_decap_8 FILLER_52_330 ();
 sg13g2_decap_4 FILLER_52_345 ();
 sg13g2_fill_2 FILLER_52_349 ();
 sg13g2_fill_2 FILLER_52_391 ();
 sg13g2_fill_2 FILLER_52_396 ();
 sg13g2_fill_2 FILLER_52_414 ();
 sg13g2_fill_1 FILLER_53_15 ();
 sg13g2_fill_1 FILLER_53_24 ();
 sg13g2_fill_1 FILLER_53_33 ();
 sg13g2_fill_2 FILLER_53_65 ();
 sg13g2_fill_2 FILLER_53_94 ();
 sg13g2_fill_1 FILLER_53_119 ();
 sg13g2_fill_1 FILLER_53_133 ();
 sg13g2_fill_1 FILLER_53_146 ();
 sg13g2_fill_1 FILLER_53_152 ();
 sg13g2_fill_2 FILLER_53_161 ();
 sg13g2_fill_1 FILLER_53_163 ();
 sg13g2_fill_1 FILLER_53_221 ();
 sg13g2_fill_1 FILLER_53_228 ();
 sg13g2_fill_1 FILLER_53_239 ();
 sg13g2_fill_1 FILLER_53_247 ();
 sg13g2_fill_1 FILLER_53_284 ();
 sg13g2_fill_2 FILLER_53_303 ();
 sg13g2_fill_1 FILLER_53_315 ();
 sg13g2_fill_1 FILLER_53_321 ();
 sg13g2_fill_2 FILLER_53_351 ();
 sg13g2_decap_4 FILLER_53_357 ();
 sg13g2_fill_2 FILLER_53_365 ();
 sg13g2_fill_1 FILLER_53_367 ();
 sg13g2_fill_2 FILLER_53_395 ();
 sg13g2_fill_2 FILLER_53_421 ();
 sg13g2_fill_1 FILLER_53_423 ();
 sg13g2_fill_2 FILLER_53_427 ();
 sg13g2_fill_1 FILLER_53_429 ();
 sg13g2_fill_1 FILLER_54_33 ();
 sg13g2_fill_2 FILLER_54_66 ();
 sg13g2_fill_1 FILLER_54_79 ();
 sg13g2_fill_1 FILLER_54_121 ();
 sg13g2_fill_1 FILLER_54_129 ();
 sg13g2_fill_1 FILLER_54_179 ();
 sg13g2_fill_1 FILLER_54_184 ();
 sg13g2_fill_1 FILLER_54_198 ();
 sg13g2_fill_2 FILLER_54_234 ();
 sg13g2_fill_1 FILLER_54_241 ();
 sg13g2_fill_2 FILLER_54_246 ();
 sg13g2_fill_1 FILLER_54_248 ();
 sg13g2_fill_2 FILLER_54_275 ();
 sg13g2_fill_1 FILLER_54_300 ();
 sg13g2_fill_1 FILLER_54_309 ();
 sg13g2_fill_2 FILLER_54_324 ();
 sg13g2_fill_1 FILLER_54_326 ();
 sg13g2_fill_1 FILLER_54_343 ();
 sg13g2_fill_2 FILLER_54_383 ();
 sg13g2_fill_1 FILLER_54_394 ();
 sg13g2_fill_2 FILLER_54_398 ();
 sg13g2_fill_1 FILLER_54_400 ();
 sg13g2_fill_2 FILLER_54_420 ();
 sg13g2_fill_1 FILLER_55_82 ();
 sg13g2_fill_1 FILLER_55_92 ();
 sg13g2_fill_2 FILLER_55_97 ();
 sg13g2_fill_1 FILLER_55_145 ();
 sg13g2_fill_1 FILLER_55_150 ();
 sg13g2_decap_4 FILLER_55_177 ();
 sg13g2_fill_2 FILLER_55_233 ();
 sg13g2_fill_2 FILLER_55_238 ();
 sg13g2_fill_2 FILLER_55_244 ();
 sg13g2_fill_2 FILLER_55_302 ();
 sg13g2_decap_4 FILLER_55_320 ();
 sg13g2_fill_2 FILLER_55_324 ();
 sg13g2_fill_2 FILLER_55_339 ();
 sg13g2_fill_2 FILLER_55_349 ();
 sg13g2_fill_2 FILLER_55_354 ();
 sg13g2_fill_1 FILLER_55_380 ();
 sg13g2_fill_2 FILLER_55_422 ();
 sg13g2_fill_2 FILLER_55_428 ();
 sg13g2_fill_1 FILLER_56_0 ();
 sg13g2_fill_1 FILLER_56_50 ();
 sg13g2_fill_2 FILLER_56_56 ();
 sg13g2_fill_1 FILLER_56_62 ();
 sg13g2_fill_1 FILLER_56_71 ();
 sg13g2_fill_2 FILLER_56_119 ();
 sg13g2_fill_1 FILLER_56_160 ();
 sg13g2_fill_2 FILLER_56_166 ();
 sg13g2_fill_1 FILLER_56_176 ();
 sg13g2_fill_2 FILLER_56_195 ();
 sg13g2_fill_1 FILLER_56_197 ();
 sg13g2_fill_1 FILLER_56_214 ();
 sg13g2_fill_1 FILLER_56_244 ();
 sg13g2_fill_1 FILLER_56_250 ();
 sg13g2_fill_2 FILLER_56_256 ();
 sg13g2_fill_2 FILLER_56_271 ();
 sg13g2_fill_1 FILLER_56_273 ();
 sg13g2_fill_1 FILLER_56_284 ();
 sg13g2_fill_1 FILLER_56_290 ();
 sg13g2_fill_2 FILLER_56_299 ();
 sg13g2_fill_2 FILLER_56_327 ();
 sg13g2_fill_1 FILLER_56_334 ();
 sg13g2_fill_1 FILLER_56_362 ();
 sg13g2_fill_1 FILLER_56_423 ();
 sg13g2_fill_1 FILLER_56_429 ();
 sg13g2_fill_2 FILLER_57_64 ();
 sg13g2_fill_1 FILLER_57_79 ();
 sg13g2_fill_1 FILLER_57_85 ();
 sg13g2_fill_1 FILLER_57_95 ();
 sg13g2_fill_1 FILLER_57_101 ();
 sg13g2_fill_1 FILLER_57_114 ();
 sg13g2_fill_2 FILLER_57_146 ();
 sg13g2_fill_1 FILLER_57_157 ();
 sg13g2_fill_2 FILLER_57_205 ();
 sg13g2_fill_2 FILLER_57_211 ();
 sg13g2_fill_1 FILLER_57_213 ();
 sg13g2_fill_2 FILLER_57_240 ();
 sg13g2_decap_4 FILLER_57_258 ();
 sg13g2_fill_1 FILLER_57_262 ();
 sg13g2_fill_2 FILLER_57_278 ();
 sg13g2_fill_1 FILLER_57_295 ();
 sg13g2_fill_2 FILLER_57_357 ();
 sg13g2_decap_4 FILLER_57_376 ();
 sg13g2_fill_2 FILLER_57_393 ();
 sg13g2_fill_2 FILLER_58_44 ();
 sg13g2_fill_1 FILLER_58_132 ();
 sg13g2_fill_2 FILLER_58_159 ();
 sg13g2_fill_2 FILLER_58_176 ();
 sg13g2_fill_1 FILLER_58_178 ();
 sg13g2_fill_1 FILLER_58_184 ();
 sg13g2_fill_2 FILLER_58_193 ();
 sg13g2_fill_1 FILLER_58_195 ();
 sg13g2_fill_1 FILLER_58_199 ();
 sg13g2_fill_1 FILLER_58_226 ();
 sg13g2_decap_8 FILLER_58_232 ();
 sg13g2_fill_1 FILLER_58_244 ();
 sg13g2_fill_2 FILLER_58_253 ();
 sg13g2_fill_1 FILLER_58_261 ();
 sg13g2_fill_2 FILLER_58_265 ();
 sg13g2_decap_4 FILLER_58_271 ();
 sg13g2_fill_2 FILLER_58_315 ();
 sg13g2_fill_1 FILLER_58_366 ();
 sg13g2_fill_1 FILLER_58_389 ();
 sg13g2_fill_1 FILLER_58_395 ();
 sg13g2_fill_1 FILLER_58_400 ();
 sg13g2_fill_1 FILLER_58_404 ();
 sg13g2_fill_1 FILLER_58_429 ();
 sg13g2_fill_1 FILLER_59_72 ();
 sg13g2_fill_2 FILLER_59_77 ();
 sg13g2_fill_1 FILLER_59_87 ();
 sg13g2_fill_1 FILLER_59_112 ();
 sg13g2_fill_2 FILLER_59_133 ();
 sg13g2_fill_2 FILLER_59_153 ();
 sg13g2_fill_2 FILLER_59_185 ();
 sg13g2_fill_2 FILLER_59_200 ();
 sg13g2_fill_1 FILLER_59_202 ();
 sg13g2_fill_2 FILLER_59_208 ();
 sg13g2_fill_1 FILLER_59_210 ();
 sg13g2_fill_1 FILLER_59_215 ();
 sg13g2_fill_2 FILLER_59_227 ();
 sg13g2_fill_1 FILLER_59_297 ();
 sg13g2_fill_1 FILLER_59_325 ();
 sg13g2_fill_2 FILLER_59_330 ();
 sg13g2_fill_1 FILLER_59_332 ();
 sg13g2_fill_2 FILLER_59_336 ();
 sg13g2_fill_2 FILLER_59_353 ();
 sg13g2_fill_1 FILLER_59_355 ();
 sg13g2_fill_2 FILLER_59_394 ();
 sg13g2_fill_2 FILLER_59_404 ();
 sg13g2_fill_2 FILLER_60_26 ();
 sg13g2_fill_2 FILLER_60_41 ();
 sg13g2_fill_1 FILLER_60_51 ();
 sg13g2_fill_1 FILLER_60_66 ();
 sg13g2_fill_1 FILLER_60_72 ();
 sg13g2_fill_1 FILLER_60_146 ();
 sg13g2_fill_1 FILLER_60_152 ();
 sg13g2_fill_1 FILLER_60_161 ();
 sg13g2_fill_1 FILLER_60_170 ();
 sg13g2_fill_1 FILLER_60_176 ();
 sg13g2_fill_2 FILLER_60_185 ();
 sg13g2_fill_2 FILLER_60_255 ();
 sg13g2_fill_1 FILLER_60_265 ();
 sg13g2_fill_1 FILLER_60_305 ();
 sg13g2_fill_2 FILLER_60_332 ();
 sg13g2_fill_1 FILLER_60_339 ();
 sg13g2_fill_1 FILLER_60_348 ();
 sg13g2_fill_2 FILLER_60_357 ();
 sg13g2_fill_2 FILLER_60_371 ();
 sg13g2_fill_1 FILLER_60_373 ();
 sg13g2_fill_1 FILLER_60_378 ();
 sg13g2_fill_2 FILLER_60_395 ();
 sg13g2_fill_2 FILLER_60_406 ();
 sg13g2_fill_2 FILLER_60_411 ();
 sg13g2_fill_2 FILLER_60_428 ();
 sg13g2_fill_1 FILLER_61_4 ();
 sg13g2_fill_1 FILLER_61_56 ();
 sg13g2_fill_2 FILLER_61_146 ();
 sg13g2_fill_1 FILLER_61_153 ();
 sg13g2_fill_1 FILLER_61_162 ();
 sg13g2_fill_1 FILLER_61_168 ();
 sg13g2_fill_1 FILLER_61_174 ();
 sg13g2_fill_1 FILLER_61_179 ();
 sg13g2_fill_1 FILLER_61_185 ();
 sg13g2_fill_1 FILLER_61_194 ();
 sg13g2_fill_1 FILLER_61_215 ();
 sg13g2_decap_4 FILLER_61_233 ();
 sg13g2_fill_2 FILLER_61_237 ();
 sg13g2_fill_1 FILLER_61_256 ();
 sg13g2_fill_1 FILLER_61_312 ();
 sg13g2_fill_2 FILLER_61_330 ();
 sg13g2_decap_4 FILLER_61_343 ();
 sg13g2_fill_1 FILLER_61_347 ();
 sg13g2_fill_1 FILLER_61_355 ();
 sg13g2_fill_1 FILLER_61_368 ();
 sg13g2_decap_4 FILLER_61_379 ();
 sg13g2_fill_1 FILLER_61_389 ();
 sg13g2_fill_2 FILLER_61_412 ();
 sg13g2_fill_1 FILLER_62_0 ();
 sg13g2_fill_1 FILLER_62_9 ();
 sg13g2_fill_1 FILLER_62_20 ();
 sg13g2_fill_2 FILLER_62_45 ();
 sg13g2_fill_2 FILLER_62_114 ();
 sg13g2_fill_2 FILLER_62_133 ();
 sg13g2_fill_2 FILLER_62_182 ();
 sg13g2_fill_1 FILLER_62_246 ();
 sg13g2_fill_1 FILLER_62_250 ();
 sg13g2_fill_1 FILLER_62_256 ();
 sg13g2_fill_1 FILLER_62_261 ();
 sg13g2_fill_1 FILLER_62_267 ();
 sg13g2_fill_1 FILLER_62_309 ();
 sg13g2_decap_4 FILLER_62_319 ();
 sg13g2_fill_1 FILLER_62_340 ();
 sg13g2_fill_1 FILLER_62_368 ();
 sg13g2_fill_1 FILLER_62_396 ();
 sg13g2_decap_4 FILLER_62_409 ();
 sg13g2_fill_1 FILLER_62_413 ();
 sg13g2_fill_1 FILLER_62_423 ();
 sg13g2_fill_2 FILLER_62_427 ();
 sg13g2_fill_1 FILLER_62_429 ();
 sg13g2_fill_2 FILLER_63_31 ();
 sg13g2_fill_1 FILLER_63_104 ();
 sg13g2_fill_1 FILLER_63_118 ();
 sg13g2_fill_2 FILLER_63_154 ();
 sg13g2_fill_2 FILLER_63_161 ();
 sg13g2_fill_1 FILLER_63_186 ();
 sg13g2_fill_2 FILLER_63_222 ();
 sg13g2_fill_1 FILLER_63_224 ();
 sg13g2_fill_1 FILLER_63_259 ();
 sg13g2_fill_1 FILLER_63_296 ();
 sg13g2_fill_1 FILLER_63_306 ();
 sg13g2_fill_1 FILLER_63_310 ();
 sg13g2_fill_2 FILLER_63_323 ();
 sg13g2_fill_1 FILLER_63_325 ();
 sg13g2_fill_2 FILLER_63_330 ();
 sg13g2_fill_1 FILLER_63_341 ();
 sg13g2_fill_2 FILLER_63_359 ();
 sg13g2_fill_2 FILLER_63_370 ();
 sg13g2_fill_2 FILLER_63_377 ();
 sg13g2_fill_2 FILLER_63_382 ();
 sg13g2_fill_1 FILLER_63_384 ();
 sg13g2_fill_1 FILLER_63_393 ();
 sg13g2_fill_1 FILLER_63_398 ();
 sg13g2_fill_1 FILLER_63_404 ();
 sg13g2_fill_1 FILLER_63_409 ();
 sg13g2_fill_1 FILLER_64_0 ();
 sg13g2_fill_2 FILLER_64_9 ();
 sg13g2_fill_2 FILLER_64_66 ();
 sg13g2_fill_1 FILLER_64_75 ();
 sg13g2_fill_1 FILLER_64_95 ();
 sg13g2_fill_2 FILLER_64_188 ();
 sg13g2_fill_2 FILLER_64_208 ();
 sg13g2_decap_4 FILLER_64_267 ();
 sg13g2_fill_1 FILLER_64_271 ();
 sg13g2_decap_4 FILLER_64_284 ();
 sg13g2_fill_1 FILLER_64_292 ();
 sg13g2_decap_4 FILLER_64_332 ();
 sg13g2_fill_2 FILLER_64_336 ();
 sg13g2_fill_1 FILLER_64_348 ();
 sg13g2_fill_1 FILLER_64_373 ();
 sg13g2_decap_4 FILLER_64_383 ();
 sg13g2_fill_2 FILLER_64_387 ();
 sg13g2_fill_1 FILLER_64_393 ();
 sg13g2_fill_1 FILLER_64_414 ();
 sg13g2_fill_2 FILLER_64_428 ();
 sg13g2_fill_1 FILLER_65_26 ();
 sg13g2_fill_1 FILLER_65_77 ();
 sg13g2_fill_2 FILLER_65_115 ();
 sg13g2_fill_1 FILLER_65_159 ();
 sg13g2_fill_2 FILLER_65_225 ();
 sg13g2_fill_1 FILLER_65_227 ();
 sg13g2_fill_1 FILLER_65_232 ();
 sg13g2_decap_4 FILLER_65_253 ();
 sg13g2_fill_1 FILLER_65_275 ();
 sg13g2_fill_1 FILLER_65_281 ();
 sg13g2_fill_2 FILLER_65_291 ();
 sg13g2_fill_1 FILLER_65_298 ();
 sg13g2_fill_2 FILLER_65_303 ();
 sg13g2_fill_2 FILLER_65_309 ();
 sg13g2_fill_2 FILLER_65_315 ();
 sg13g2_fill_1 FILLER_65_317 ();
 sg13g2_fill_1 FILLER_65_323 ();
 sg13g2_fill_2 FILLER_65_336 ();
 sg13g2_fill_1 FILLER_65_344 ();
 sg13g2_fill_2 FILLER_65_353 ();
 sg13g2_fill_2 FILLER_65_367 ();
 sg13g2_fill_2 FILLER_65_397 ();
 sg13g2_fill_1 FILLER_65_403 ();
 sg13g2_fill_2 FILLER_65_428 ();
 sg13g2_fill_2 FILLER_66_0 ();
 sg13g2_fill_2 FILLER_66_32 ();
 sg13g2_fill_1 FILLER_66_42 ();
 sg13g2_fill_1 FILLER_66_55 ();
 sg13g2_fill_2 FILLER_66_116 ();
 sg13g2_fill_2 FILLER_66_152 ();
 sg13g2_fill_2 FILLER_66_175 ();
 sg13g2_fill_1 FILLER_66_195 ();
 sg13g2_fill_2 FILLER_66_200 ();
 sg13g2_fill_1 FILLER_66_238 ();
 sg13g2_fill_1 FILLER_66_246 ();
 sg13g2_fill_1 FILLER_66_255 ();
 sg13g2_fill_2 FILLER_66_284 ();
 sg13g2_fill_1 FILLER_66_306 ();
 sg13g2_fill_1 FILLER_66_313 ();
 sg13g2_fill_1 FILLER_66_318 ();
 sg13g2_fill_2 FILLER_66_324 ();
 sg13g2_decap_4 FILLER_66_342 ();
 sg13g2_fill_1 FILLER_66_346 ();
 sg13g2_fill_2 FILLER_66_372 ();
 sg13g2_fill_2 FILLER_66_417 ();
 sg13g2_fill_1 FILLER_66_419 ();
 sg13g2_fill_2 FILLER_66_428 ();
 sg13g2_fill_1 FILLER_67_21 ();
 sg13g2_fill_1 FILLER_67_75 ();
 sg13g2_fill_2 FILLER_67_108 ();
 sg13g2_fill_2 FILLER_67_163 ();
 sg13g2_fill_2 FILLER_67_210 ();
 sg13g2_fill_1 FILLER_67_248 ();
 sg13g2_fill_2 FILLER_67_261 ();
 sg13g2_fill_1 FILLER_67_281 ();
 sg13g2_fill_1 FILLER_67_287 ();
 sg13g2_fill_1 FILLER_67_293 ();
 sg13g2_fill_2 FILLER_67_298 ();
 sg13g2_fill_1 FILLER_67_305 ();
 sg13g2_fill_1 FILLER_67_313 ();
 sg13g2_fill_2 FILLER_67_337 ();
 sg13g2_fill_2 FILLER_67_343 ();
 sg13g2_decap_4 FILLER_67_352 ();
 sg13g2_fill_1 FILLER_67_361 ();
 sg13g2_fill_2 FILLER_67_379 ();
 sg13g2_fill_1 FILLER_67_400 ();
 sg13g2_fill_2 FILLER_67_404 ();
 sg13g2_fill_1 FILLER_67_410 ();
 sg13g2_fill_2 FILLER_67_415 ();
 sg13g2_decap_4 FILLER_67_426 ();
 sg13g2_fill_2 FILLER_68_56 ();
 sg13g2_fill_1 FILLER_68_117 ();
 sg13g2_fill_2 FILLER_68_138 ();
 sg13g2_fill_1 FILLER_68_178 ();
 sg13g2_fill_2 FILLER_68_190 ();
 sg13g2_fill_1 FILLER_68_230 ();
 sg13g2_fill_1 FILLER_68_235 ();
 sg13g2_fill_1 FILLER_68_303 ();
 sg13g2_fill_1 FILLER_68_312 ();
 sg13g2_fill_1 FILLER_68_318 ();
 sg13g2_fill_1 FILLER_68_337 ();
 sg13g2_fill_1 FILLER_68_345 ();
 sg13g2_fill_1 FILLER_68_350 ();
 sg13g2_decap_4 FILLER_68_355 ();
 sg13g2_fill_1 FILLER_68_367 ();
 sg13g2_fill_2 FILLER_68_390 ();
 sg13g2_fill_1 FILLER_68_392 ();
 sg13g2_decap_4 FILLER_68_397 ();
 sg13g2_fill_2 FILLER_68_401 ();
 sg13g2_decap_4 FILLER_68_407 ();
 sg13g2_fill_2 FILLER_68_421 ();
 sg13g2_fill_1 FILLER_68_423 ();
 sg13g2_fill_2 FILLER_68_428 ();
 sg13g2_fill_1 FILLER_69_16 ();
 sg13g2_fill_1 FILLER_69_229 ();
 sg13g2_fill_2 FILLER_69_235 ();
 sg13g2_fill_1 FILLER_69_252 ();
 sg13g2_fill_1 FILLER_69_301 ();
 sg13g2_fill_1 FILLER_69_310 ();
 sg13g2_fill_1 FILLER_69_330 ();
 sg13g2_fill_1 FILLER_69_335 ();
 sg13g2_fill_2 FILLER_69_366 ();
 sg13g2_fill_1 FILLER_69_377 ();
 sg13g2_decap_4 FILLER_69_406 ();
 sg13g2_fill_1 FILLER_69_410 ();
 sg13g2_fill_2 FILLER_69_427 ();
 sg13g2_fill_1 FILLER_69_429 ();
 sg13g2_fill_2 FILLER_70_47 ();
 sg13g2_fill_2 FILLER_70_78 ();
 sg13g2_fill_2 FILLER_70_128 ();
 sg13g2_fill_2 FILLER_70_211 ();
 sg13g2_fill_2 FILLER_70_236 ();
 sg13g2_fill_1 FILLER_70_261 ();
 sg13g2_fill_2 FILLER_70_288 ();
 sg13g2_fill_1 FILLER_70_300 ();
 sg13g2_fill_2 FILLER_70_354 ();
 sg13g2_fill_2 FILLER_70_360 ();
 sg13g2_fill_1 FILLER_70_362 ();
 sg13g2_fill_1 FILLER_70_367 ();
 sg13g2_fill_1 FILLER_70_372 ();
 sg13g2_fill_1 FILLER_70_376 ();
 sg13g2_fill_1 FILLER_70_381 ();
 sg13g2_fill_2 FILLER_70_387 ();
 sg13g2_fill_1 FILLER_70_389 ();
 sg13g2_fill_2 FILLER_70_415 ();
 sg13g2_fill_1 FILLER_71_17 ();
 sg13g2_fill_2 FILLER_71_60 ();
 sg13g2_fill_1 FILLER_71_106 ();
 sg13g2_fill_1 FILLER_71_179 ();
 sg13g2_fill_1 FILLER_71_188 ();
 sg13g2_fill_1 FILLER_71_215 ();
 sg13g2_fill_1 FILLER_71_223 ();
 sg13g2_fill_2 FILLER_71_285 ();
 sg13g2_decap_4 FILLER_71_290 ();
 sg13g2_fill_2 FILLER_71_294 ();
 sg13g2_fill_1 FILLER_71_306 ();
 sg13g2_fill_1 FILLER_71_310 ();
 sg13g2_fill_1 FILLER_71_320 ();
 sg13g2_fill_2 FILLER_71_326 ();
 sg13g2_fill_2 FILLER_71_391 ();
 sg13g2_fill_1 FILLER_71_416 ();
 sg13g2_fill_2 FILLER_71_421 ();
 sg13g2_fill_2 FILLER_71_427 ();
 sg13g2_fill_1 FILLER_71_429 ();
 sg13g2_fill_2 FILLER_72_138 ();
 sg13g2_fill_2 FILLER_72_165 ();
 sg13g2_fill_2 FILLER_72_179 ();
 sg13g2_fill_2 FILLER_72_225 ();
 sg13g2_fill_1 FILLER_72_251 ();
 sg13g2_fill_2 FILLER_72_265 ();
 sg13g2_fill_1 FILLER_72_317 ();
 sg13g2_fill_1 FILLER_72_322 ();
 sg13g2_fill_1 FILLER_72_331 ();
 sg13g2_fill_1 FILLER_72_336 ();
 sg13g2_decap_4 FILLER_72_357 ();
 sg13g2_fill_2 FILLER_72_361 ();
 sg13g2_fill_2 FILLER_72_376 ();
 sg13g2_fill_1 FILLER_72_378 ();
 sg13g2_fill_2 FILLER_72_384 ();
 sg13g2_fill_1 FILLER_72_386 ();
 sg13g2_fill_1 FILLER_72_396 ();
 sg13g2_fill_1 FILLER_72_401 ();
 sg13g2_fill_1 FILLER_72_411 ();
 sg13g2_fill_1 FILLER_73_8 ();
 sg13g2_fill_1 FILLER_73_21 ();
 sg13g2_fill_2 FILLER_73_27 ();
 sg13g2_fill_1 FILLER_73_105 ();
 sg13g2_fill_1 FILLER_73_123 ();
 sg13g2_fill_1 FILLER_73_128 ();
 sg13g2_fill_2 FILLER_73_189 ();
 sg13g2_fill_1 FILLER_73_196 ();
 sg13g2_fill_1 FILLER_73_219 ();
 sg13g2_fill_2 FILLER_73_293 ();
 sg13g2_fill_2 FILLER_73_313 ();
 sg13g2_fill_1 FILLER_73_337 ();
 sg13g2_fill_1 FILLER_73_343 ();
 sg13g2_fill_2 FILLER_73_349 ();
 sg13g2_fill_1 FILLER_73_356 ();
 sg13g2_fill_2 FILLER_73_362 ();
 sg13g2_fill_1 FILLER_73_364 ();
 sg13g2_fill_2 FILLER_73_427 ();
 sg13g2_fill_1 FILLER_73_429 ();
 sg13g2_fill_1 FILLER_74_31 ();
 sg13g2_fill_1 FILLER_74_38 ();
 sg13g2_fill_1 FILLER_74_220 ();
 sg13g2_fill_2 FILLER_74_307 ();
 sg13g2_fill_2 FILLER_74_313 ();
 sg13g2_fill_1 FILLER_74_327 ();
 sg13g2_fill_1 FILLER_74_336 ();
 sg13g2_fill_2 FILLER_74_354 ();
 sg13g2_fill_1 FILLER_74_356 ();
 sg13g2_decap_8 FILLER_74_361 ();
 sg13g2_decap_8 FILLER_74_368 ();
 sg13g2_fill_2 FILLER_74_375 ();
 sg13g2_fill_1 FILLER_74_377 ();
 sg13g2_fill_1 FILLER_74_390 ();
 sg13g2_fill_2 FILLER_74_395 ();
 sg13g2_fill_1 FILLER_74_397 ();
 sg13g2_decap_4 FILLER_74_410 ();
 sg13g2_fill_1 FILLER_74_414 ();
 sg13g2_fill_2 FILLER_74_427 ();
 sg13g2_fill_1 FILLER_74_429 ();
 sg13g2_fill_1 FILLER_75_17 ();
 sg13g2_fill_2 FILLER_75_52 ();
 sg13g2_fill_2 FILLER_75_74 ();
 sg13g2_fill_1 FILLER_75_104 ();
 sg13g2_fill_1 FILLER_75_237 ();
 sg13g2_fill_1 FILLER_75_241 ();
 sg13g2_fill_2 FILLER_75_298 ();
 sg13g2_fill_1 FILLER_75_344 ();
 sg13g2_fill_1 FILLER_75_354 ();
 sg13g2_decap_8 FILLER_75_401 ();
 sg13g2_decap_8 FILLER_75_408 ();
 sg13g2_decap_8 FILLER_75_415 ();
 sg13g2_decap_8 FILLER_75_422 ();
 sg13g2_fill_1 FILLER_75_429 ();
 sg13g2_fill_1 FILLER_76_100 ();
 sg13g2_fill_2 FILLER_76_127 ();
 sg13g2_fill_2 FILLER_76_237 ();
 sg13g2_fill_1 FILLER_76_246 ();
 sg13g2_fill_1 FILLER_76_252 ();
 sg13g2_fill_1 FILLER_76_257 ();
 sg13g2_fill_1 FILLER_76_266 ();
 sg13g2_fill_1 FILLER_76_340 ();
 sg13g2_fill_1 FILLER_76_358 ();
 sg13g2_decap_8 FILLER_76_401 ();
 sg13g2_decap_8 FILLER_76_408 ();
 sg13g2_decap_8 FILLER_76_415 ();
 sg13g2_decap_8 FILLER_76_422 ();
 sg13g2_fill_1 FILLER_76_429 ();
 sg13g2_fill_1 FILLER_77_0 ();
 sg13g2_fill_1 FILLER_77_14 ();
 sg13g2_fill_1 FILLER_77_191 ();
 sg13g2_fill_2 FILLER_77_196 ();
 sg13g2_fill_1 FILLER_77_232 ();
 sg13g2_fill_1 FILLER_77_273 ();
 sg13g2_fill_1 FILLER_77_316 ();
 sg13g2_fill_2 FILLER_77_350 ();
 sg13g2_fill_1 FILLER_77_378 ();
 sg13g2_decap_8 FILLER_77_405 ();
 sg13g2_decap_8 FILLER_77_412 ();
 sg13g2_decap_8 FILLER_77_419 ();
 sg13g2_decap_4 FILLER_77_426 ();
 sg13g2_fill_2 FILLER_78_34 ();
 sg13g2_fill_1 FILLER_78_44 ();
 sg13g2_fill_2 FILLER_78_113 ();
 sg13g2_fill_1 FILLER_78_174 ();
 sg13g2_fill_1 FILLER_78_299 ();
 sg13g2_fill_2 FILLER_78_319 ();
 sg13g2_fill_1 FILLER_78_329 ();
 sg13g2_fill_2 FILLER_78_334 ();
 sg13g2_fill_2 FILLER_78_357 ();
 sg13g2_fill_2 FILLER_78_363 ();
 sg13g2_fill_2 FILLER_78_369 ();
 sg13g2_decap_8 FILLER_78_410 ();
 sg13g2_decap_8 FILLER_78_417 ();
 sg13g2_decap_4 FILLER_78_424 ();
 sg13g2_fill_2 FILLER_78_428 ();
 sg13g2_fill_1 FILLER_79_0 ();
 sg13g2_fill_1 FILLER_79_9 ();
 sg13g2_fill_1 FILLER_79_217 ();
 sg13g2_fill_2 FILLER_79_230 ();
 sg13g2_fill_2 FILLER_79_248 ();
 sg13g2_fill_2 FILLER_79_262 ();
 sg13g2_fill_2 FILLER_79_333 ();
 sg13g2_fill_1 FILLER_79_376 ();
 sg13g2_decap_8 FILLER_79_411 ();
 sg13g2_decap_8 FILLER_79_418 ();
 sg13g2_decap_4 FILLER_79_425 ();
 sg13g2_fill_1 FILLER_79_429 ();
 sg13g2_fill_1 FILLER_80_146 ();
 sg13g2_fill_1 FILLER_80_151 ();
 sg13g2_fill_2 FILLER_80_184 ();
 sg13g2_fill_1 FILLER_80_301 ();
 sg13g2_fill_1 FILLER_80_310 ();
 sg13g2_fill_1 FILLER_80_319 ();
 sg13g2_fill_2 FILLER_80_328 ();
 sg13g2_fill_2 FILLER_80_342 ();
 sg13g2_fill_1 FILLER_80_348 ();
 sg13g2_decap_8 FILLER_80_407 ();
 sg13g2_decap_8 FILLER_80_414 ();
 sg13g2_decap_8 FILLER_80_421 ();
 sg13g2_fill_2 FILLER_80_428 ();
endmodule
