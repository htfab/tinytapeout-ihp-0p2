module tt_um_MichaelBell_mandelbrot (clk,
    ena,
    rst_n,
    ui_in,
    uio_in,
    uio_oe,
    uio_out,
    uo_out);
 input clk;
 input ena;
 input rst_n;
 input [7:0] ui_in;
 input [7:0] uio_in;
 output [7:0] uio_oe;
 output [7:0] uio_out;
 output [7:0] uo_out;

 wire _00000_;
 wire _00001_;
 wire _00002_;
 wire _00003_;
 wire _00004_;
 wire _00005_;
 wire _00006_;
 wire _00007_;
 wire _00008_;
 wire _00009_;
 wire _00010_;
 wire _00011_;
 wire _00012_;
 wire _00013_;
 wire _00014_;
 wire _00015_;
 wire _00016_;
 wire _00017_;
 wire _00018_;
 wire _00019_;
 wire _00020_;
 wire _00021_;
 wire _00022_;
 wire _00023_;
 wire _00024_;
 wire _00025_;
 wire _00026_;
 wire _00027_;
 wire _00028_;
 wire _00029_;
 wire _00030_;
 wire _00031_;
 wire _00032_;
 wire _00033_;
 wire _00034_;
 wire _00035_;
 wire _00036_;
 wire _00037_;
 wire _00038_;
 wire _00039_;
 wire _00040_;
 wire _00041_;
 wire _00042_;
 wire _00043_;
 wire _00044_;
 wire _00045_;
 wire _00046_;
 wire _00047_;
 wire _00048_;
 wire _00049_;
 wire _00050_;
 wire _00051_;
 wire _00052_;
 wire _00053_;
 wire _00054_;
 wire _00055_;
 wire _00056_;
 wire _00057_;
 wire _00058_;
 wire _00059_;
 wire _00060_;
 wire _00061_;
 wire _00062_;
 wire _00063_;
 wire _00064_;
 wire _00065_;
 wire _00066_;
 wire _00067_;
 wire _00068_;
 wire _00069_;
 wire _00070_;
 wire _00071_;
 wire _00072_;
 wire _00073_;
 wire _00074_;
 wire _00075_;
 wire _00076_;
 wire _00077_;
 wire _00078_;
 wire _00079_;
 wire _00080_;
 wire _00081_;
 wire _00082_;
 wire _00083_;
 wire _00084_;
 wire _00085_;
 wire _00086_;
 wire _00087_;
 wire _00088_;
 wire _00089_;
 wire _00090_;
 wire _00091_;
 wire _00092_;
 wire _00093_;
 wire _00094_;
 wire _00095_;
 wire _00096_;
 wire _00097_;
 wire _00098_;
 wire _00099_;
 wire _00100_;
 wire _00101_;
 wire _00102_;
 wire _00103_;
 wire _00104_;
 wire _00105_;
 wire _00106_;
 wire _00107_;
 wire _00108_;
 wire _00109_;
 wire _00110_;
 wire _00111_;
 wire _00112_;
 wire _00113_;
 wire _00114_;
 wire _00115_;
 wire _00116_;
 wire _00117_;
 wire _00118_;
 wire _00119_;
 wire _00120_;
 wire _00121_;
 wire _00122_;
 wire _00123_;
 wire _00124_;
 wire _00125_;
 wire _00126_;
 wire _00127_;
 wire _00128_;
 wire _00129_;
 wire _00130_;
 wire _00131_;
 wire _00132_;
 wire _00133_;
 wire _00134_;
 wire _00135_;
 wire _00136_;
 wire _00137_;
 wire _00138_;
 wire _00139_;
 wire _00140_;
 wire _00141_;
 wire _00142_;
 wire _00143_;
 wire _00144_;
 wire _00145_;
 wire _00146_;
 wire _00147_;
 wire _00148_;
 wire _00149_;
 wire _00150_;
 wire _00151_;
 wire _00152_;
 wire _00153_;
 wire _00154_;
 wire _00155_;
 wire _00156_;
 wire _00157_;
 wire _00158_;
 wire _00159_;
 wire _00160_;
 wire _00161_;
 wire _00162_;
 wire _00163_;
 wire _00164_;
 wire _00165_;
 wire _00166_;
 wire _00167_;
 wire _00168_;
 wire _00169_;
 wire _00170_;
 wire _00171_;
 wire _00172_;
 wire _00173_;
 wire _00174_;
 wire _00175_;
 wire _00176_;
 wire _00177_;
 wire _00178_;
 wire _00179_;
 wire _00180_;
 wire _00181_;
 wire _00182_;
 wire _00183_;
 wire _00184_;
 wire _00185_;
 wire _00186_;
 wire _00187_;
 wire _00188_;
 wire _00189_;
 wire _00190_;
 wire _00191_;
 wire _00192_;
 wire _00193_;
 wire _00194_;
 wire _00195_;
 wire _00196_;
 wire _00197_;
 wire _00198_;
 wire _00199_;
 wire _00200_;
 wire _00201_;
 wire _00202_;
 wire _00203_;
 wire _00204_;
 wire _00205_;
 wire _00206_;
 wire _00207_;
 wire _00208_;
 wire _00209_;
 wire _00210_;
 wire _00211_;
 wire _00212_;
 wire _00213_;
 wire _00214_;
 wire _00215_;
 wire _00216_;
 wire _00217_;
 wire _00218_;
 wire _00219_;
 wire _00220_;
 wire _00221_;
 wire _00222_;
 wire _00223_;
 wire _00224_;
 wire _00225_;
 wire _00226_;
 wire _00227_;
 wire _00228_;
 wire _00229_;
 wire _00230_;
 wire _00231_;
 wire _00232_;
 wire _00233_;
 wire _00234_;
 wire _00235_;
 wire _00236_;
 wire _00237_;
 wire _00238_;
 wire _00239_;
 wire _00240_;
 wire _00241_;
 wire _00242_;
 wire _00243_;
 wire _00244_;
 wire _00245_;
 wire _00246_;
 wire _00247_;
 wire _00248_;
 wire _00249_;
 wire _00250_;
 wire _00251_;
 wire _00252_;
 wire _00253_;
 wire _00254_;
 wire _00255_;
 wire _00256_;
 wire _00257_;
 wire _00258_;
 wire _00259_;
 wire _00260_;
 wire _00261_;
 wire _00262_;
 wire _00263_;
 wire _00264_;
 wire _00265_;
 wire _00266_;
 wire _00267_;
 wire _00268_;
 wire _00269_;
 wire _00270_;
 wire _00271_;
 wire _00272_;
 wire _00273_;
 wire _00274_;
 wire _00275_;
 wire _00276_;
 wire _00277_;
 wire _00278_;
 wire _00279_;
 wire _00280_;
 wire _00281_;
 wire _00282_;
 wire _00283_;
 wire _00284_;
 wire _00285_;
 wire _00286_;
 wire _00287_;
 wire _00288_;
 wire _00289_;
 wire _00290_;
 wire _00291_;
 wire _00292_;
 wire _00293_;
 wire _00294_;
 wire _00295_;
 wire _00296_;
 wire _00297_;
 wire _00298_;
 wire _00299_;
 wire _00300_;
 wire _00301_;
 wire _00302_;
 wire _00303_;
 wire _00304_;
 wire _00305_;
 wire _00306_;
 wire _00307_;
 wire _00308_;
 wire _00309_;
 wire _00310_;
 wire _00311_;
 wire _00312_;
 wire _00313_;
 wire _00314_;
 wire _00315_;
 wire _00316_;
 wire _00317_;
 wire _00318_;
 wire _00319_;
 wire _00320_;
 wire _00321_;
 wire _00322_;
 wire _00323_;
 wire _00324_;
 wire _00325_;
 wire _00326_;
 wire _00327_;
 wire _00328_;
 wire _00329_;
 wire _00330_;
 wire _00331_;
 wire _00332_;
 wire _00333_;
 wire _00334_;
 wire _00335_;
 wire _00336_;
 wire _00337_;
 wire _00338_;
 wire _00339_;
 wire _00340_;
 wire _00341_;
 wire _00342_;
 wire _00343_;
 wire _00344_;
 wire _00345_;
 wire _00346_;
 wire _00347_;
 wire _00348_;
 wire _00349_;
 wire _00350_;
 wire _00351_;
 wire _00352_;
 wire _00353_;
 wire _00354_;
 wire _00355_;
 wire _00356_;
 wire _00357_;
 wire _00358_;
 wire _00359_;
 wire _00360_;
 wire _00361_;
 wire _00362_;
 wire _00363_;
 wire _00364_;
 wire _00365_;
 wire _00366_;
 wire _00367_;
 wire _00368_;
 wire _00369_;
 wire _00370_;
 wire _00371_;
 wire _00372_;
 wire _00373_;
 wire _00374_;
 wire _00375_;
 wire _00376_;
 wire _00377_;
 wire _00378_;
 wire _00379_;
 wire _00380_;
 wire _00381_;
 wire _00382_;
 wire _00383_;
 wire _00384_;
 wire _00385_;
 wire _00386_;
 wire _00387_;
 wire _00388_;
 wire _00389_;
 wire _00390_;
 wire _00391_;
 wire _00392_;
 wire _00393_;
 wire _00394_;
 wire _00395_;
 wire _00396_;
 wire _00397_;
 wire _00398_;
 wire _00399_;
 wire _00400_;
 wire _00401_;
 wire _00402_;
 wire _00403_;
 wire _00404_;
 wire _00405_;
 wire _00406_;
 wire _00407_;
 wire _00408_;
 wire _00409_;
 wire _00410_;
 wire _00411_;
 wire _00412_;
 wire _00413_;
 wire _00414_;
 wire _00415_;
 wire _00416_;
 wire _00417_;
 wire _00418_;
 wire _00419_;
 wire _00420_;
 wire _00421_;
 wire _00422_;
 wire _00423_;
 wire _00424_;
 wire _00425_;
 wire _00426_;
 wire _00427_;
 wire _00428_;
 wire _00429_;
 wire _00430_;
 wire _00431_;
 wire _00432_;
 wire _00433_;
 wire _00434_;
 wire _00435_;
 wire _00436_;
 wire _00437_;
 wire _00438_;
 wire _00439_;
 wire _00440_;
 wire _00441_;
 wire _00442_;
 wire _00443_;
 wire _00444_;
 wire _00445_;
 wire _00446_;
 wire _00447_;
 wire _00448_;
 wire _00449_;
 wire _00450_;
 wire _00451_;
 wire _00452_;
 wire _00453_;
 wire _00454_;
 wire _00455_;
 wire _00456_;
 wire _00457_;
 wire _00458_;
 wire _00459_;
 wire _00460_;
 wire _00461_;
 wire _00462_;
 wire _00463_;
 wire _00464_;
 wire _00465_;
 wire _00466_;
 wire _00467_;
 wire _00468_;
 wire _00469_;
 wire _00470_;
 wire _00471_;
 wire _00472_;
 wire _00473_;
 wire _00474_;
 wire _00475_;
 wire _00476_;
 wire _00477_;
 wire _00478_;
 wire _00479_;
 wire _00480_;
 wire _00481_;
 wire _00482_;
 wire _00483_;
 wire _00484_;
 wire _00485_;
 wire _00486_;
 wire _00487_;
 wire _00488_;
 wire _00489_;
 wire _00490_;
 wire _00491_;
 wire _00492_;
 wire _00493_;
 wire _00494_;
 wire _00495_;
 wire _00496_;
 wire _00497_;
 wire _00498_;
 wire _00499_;
 wire _00500_;
 wire _00501_;
 wire _00502_;
 wire _00503_;
 wire _00504_;
 wire _00505_;
 wire _00506_;
 wire _00507_;
 wire _00508_;
 wire _00509_;
 wire _00510_;
 wire _00511_;
 wire _00512_;
 wire _00513_;
 wire _00514_;
 wire _00515_;
 wire _00516_;
 wire _00517_;
 wire _00518_;
 wire _00519_;
 wire _00520_;
 wire _00521_;
 wire _00522_;
 wire _00523_;
 wire _00524_;
 wire _00525_;
 wire _00526_;
 wire _00527_;
 wire _00528_;
 wire _00529_;
 wire _00530_;
 wire _00531_;
 wire _00532_;
 wire _00533_;
 wire _00534_;
 wire _00535_;
 wire _00536_;
 wire _00537_;
 wire _00538_;
 wire _00539_;
 wire _00540_;
 wire _00541_;
 wire _00542_;
 wire _00543_;
 wire _00544_;
 wire _00545_;
 wire _00546_;
 wire _00547_;
 wire _00548_;
 wire _00549_;
 wire _00550_;
 wire _00551_;
 wire _00552_;
 wire _00553_;
 wire _00554_;
 wire _00555_;
 wire _00556_;
 wire _00557_;
 wire _00558_;
 wire _00559_;
 wire _00560_;
 wire _00561_;
 wire _00562_;
 wire _00563_;
 wire _00564_;
 wire _00565_;
 wire _00566_;
 wire _00567_;
 wire _00568_;
 wire _00569_;
 wire _00570_;
 wire _00571_;
 wire _00572_;
 wire _00573_;
 wire _00574_;
 wire _00575_;
 wire _00576_;
 wire _00577_;
 wire _00578_;
 wire _00579_;
 wire _00580_;
 wire _00581_;
 wire _00582_;
 wire _00583_;
 wire _00584_;
 wire _00585_;
 wire _00586_;
 wire _00587_;
 wire _00588_;
 wire _00589_;
 wire _00590_;
 wire _00591_;
 wire _00592_;
 wire _00593_;
 wire _00594_;
 wire _00595_;
 wire _00596_;
 wire _00597_;
 wire _00598_;
 wire _00599_;
 wire _00600_;
 wire _00601_;
 wire _00602_;
 wire _00603_;
 wire _00604_;
 wire _00605_;
 wire _00606_;
 wire _00607_;
 wire _00608_;
 wire _00609_;
 wire _00610_;
 wire _00611_;
 wire _00612_;
 wire _00613_;
 wire _00614_;
 wire _00615_;
 wire _00616_;
 wire _00617_;
 wire _00618_;
 wire _00619_;
 wire _00620_;
 wire _00621_;
 wire _00622_;
 wire _00623_;
 wire _00624_;
 wire _00625_;
 wire _00626_;
 wire _00627_;
 wire _00628_;
 wire _00629_;
 wire _00630_;
 wire _00631_;
 wire _00632_;
 wire _00633_;
 wire _00634_;
 wire _00635_;
 wire _00636_;
 wire _00637_;
 wire _00638_;
 wire _00639_;
 wire _00640_;
 wire _00641_;
 wire _00642_;
 wire _00643_;
 wire _00644_;
 wire _00645_;
 wire _00646_;
 wire _00647_;
 wire _00648_;
 wire _00649_;
 wire _00650_;
 wire _00651_;
 wire _00652_;
 wire _00653_;
 wire _00654_;
 wire _00655_;
 wire _00656_;
 wire _00657_;
 wire _00658_;
 wire _00659_;
 wire _00660_;
 wire _00661_;
 wire _00662_;
 wire _00663_;
 wire _00664_;
 wire _00665_;
 wire _00666_;
 wire _00667_;
 wire _00668_;
 wire _00669_;
 wire _00670_;
 wire _00671_;
 wire _00672_;
 wire _00673_;
 wire _00674_;
 wire _00675_;
 wire _00676_;
 wire _00677_;
 wire _00678_;
 wire _00679_;
 wire _00680_;
 wire _00681_;
 wire _00682_;
 wire _00683_;
 wire _00684_;
 wire _00685_;
 wire _00686_;
 wire _00687_;
 wire _00688_;
 wire _00689_;
 wire _00690_;
 wire _00691_;
 wire _00692_;
 wire _00693_;
 wire _00694_;
 wire _00695_;
 wire _00696_;
 wire _00697_;
 wire _00698_;
 wire _00699_;
 wire _00700_;
 wire _00701_;
 wire _00702_;
 wire _00703_;
 wire _00704_;
 wire _00705_;
 wire _00706_;
 wire _00707_;
 wire _00708_;
 wire _00709_;
 wire _00710_;
 wire _00711_;
 wire _00712_;
 wire _00713_;
 wire _00714_;
 wire _00715_;
 wire _00716_;
 wire _00717_;
 wire _00718_;
 wire _00719_;
 wire _00720_;
 wire _00721_;
 wire _00722_;
 wire _00723_;
 wire _00724_;
 wire _00725_;
 wire _00726_;
 wire _00727_;
 wire _00728_;
 wire _00729_;
 wire _00730_;
 wire _00731_;
 wire _00732_;
 wire _00733_;
 wire _00734_;
 wire _00735_;
 wire _00736_;
 wire _00737_;
 wire _00738_;
 wire _00739_;
 wire _00740_;
 wire _00741_;
 wire _00742_;
 wire _00743_;
 wire _00744_;
 wire _00745_;
 wire _00746_;
 wire _00747_;
 wire _00748_;
 wire _00749_;
 wire _00750_;
 wire _00751_;
 wire _00752_;
 wire _00753_;
 wire _00754_;
 wire _00755_;
 wire _00756_;
 wire _00757_;
 wire _00758_;
 wire _00759_;
 wire _00760_;
 wire _00761_;
 wire _00762_;
 wire _00763_;
 wire _00764_;
 wire _00765_;
 wire _00766_;
 wire _00767_;
 wire _00768_;
 wire _00769_;
 wire _00770_;
 wire _00771_;
 wire _00772_;
 wire _00773_;
 wire _00774_;
 wire _00775_;
 wire _00776_;
 wire _00777_;
 wire _00778_;
 wire _00779_;
 wire _00780_;
 wire _00781_;
 wire _00782_;
 wire _00783_;
 wire _00784_;
 wire _00785_;
 wire _00786_;
 wire _00787_;
 wire _00788_;
 wire _00789_;
 wire _00790_;
 wire _00791_;
 wire _00792_;
 wire _00793_;
 wire _00794_;
 wire _00795_;
 wire _00796_;
 wire _00797_;
 wire _00798_;
 wire _00799_;
 wire _00800_;
 wire _00801_;
 wire _00802_;
 wire _00803_;
 wire _00804_;
 wire _00805_;
 wire _00806_;
 wire _00807_;
 wire _00808_;
 wire _00809_;
 wire _00810_;
 wire _00811_;
 wire _00812_;
 wire _00813_;
 wire _00814_;
 wire _00815_;
 wire _00816_;
 wire _00817_;
 wire _00818_;
 wire _00819_;
 wire _00820_;
 wire _00821_;
 wire _00822_;
 wire _00823_;
 wire _00824_;
 wire _00825_;
 wire _00826_;
 wire _00827_;
 wire _00828_;
 wire _00829_;
 wire _00830_;
 wire _00831_;
 wire _00832_;
 wire _00833_;
 wire _00834_;
 wire _00835_;
 wire _00836_;
 wire _00837_;
 wire _00838_;
 wire _00839_;
 wire _00840_;
 wire _00841_;
 wire _00842_;
 wire _00843_;
 wire _00844_;
 wire _00845_;
 wire _00846_;
 wire _00847_;
 wire _00848_;
 wire _00849_;
 wire _00850_;
 wire _00851_;
 wire _00852_;
 wire _00853_;
 wire _00854_;
 wire _00855_;
 wire _00856_;
 wire _00857_;
 wire _00858_;
 wire _00859_;
 wire _00860_;
 wire _00861_;
 wire _00862_;
 wire _00863_;
 wire _00864_;
 wire _00865_;
 wire _00866_;
 wire _00867_;
 wire _00868_;
 wire _00869_;
 wire _00870_;
 wire _00871_;
 wire _00872_;
 wire _00873_;
 wire _00874_;
 wire _00875_;
 wire _00876_;
 wire _00877_;
 wire _00878_;
 wire _00879_;
 wire _00880_;
 wire _00881_;
 wire _00882_;
 wire _00883_;
 wire _00884_;
 wire _00885_;
 wire _00886_;
 wire _00887_;
 wire _00888_;
 wire _00889_;
 wire _00890_;
 wire _00891_;
 wire _00892_;
 wire _00893_;
 wire _00894_;
 wire _00895_;
 wire _00896_;
 wire _00897_;
 wire _00898_;
 wire _00899_;
 wire _00900_;
 wire _00901_;
 wire _00902_;
 wire _00903_;
 wire _00904_;
 wire _00905_;
 wire _00906_;
 wire _00907_;
 wire _00908_;
 wire _00909_;
 wire _00910_;
 wire _00911_;
 wire _00912_;
 wire _00913_;
 wire _00914_;
 wire _00915_;
 wire _00916_;
 wire _00917_;
 wire _00918_;
 wire _00919_;
 wire _00920_;
 wire _00921_;
 wire _00922_;
 wire _00923_;
 wire _00924_;
 wire _00925_;
 wire _00926_;
 wire _00927_;
 wire _00928_;
 wire _00929_;
 wire _00930_;
 wire _00931_;
 wire _00932_;
 wire _00933_;
 wire _00934_;
 wire _00935_;
 wire _00936_;
 wire _00937_;
 wire _00938_;
 wire _00939_;
 wire _00940_;
 wire _00941_;
 wire _00942_;
 wire _00943_;
 wire _00944_;
 wire _00945_;
 wire _00946_;
 wire _00947_;
 wire _00948_;
 wire _00949_;
 wire _00950_;
 wire _00951_;
 wire _00952_;
 wire _00953_;
 wire _00954_;
 wire _00955_;
 wire _00956_;
 wire _00957_;
 wire _00958_;
 wire _00959_;
 wire _00960_;
 wire _00961_;
 wire _00962_;
 wire _00963_;
 wire _00964_;
 wire _00965_;
 wire _00966_;
 wire _00967_;
 wire _00968_;
 wire _00969_;
 wire _00970_;
 wire _00971_;
 wire _00972_;
 wire _00973_;
 wire _00974_;
 wire _00975_;
 wire _00976_;
 wire _00977_;
 wire _00978_;
 wire _00979_;
 wire _00980_;
 wire _00981_;
 wire _00982_;
 wire _00983_;
 wire _00984_;
 wire _00985_;
 wire _00986_;
 wire _00987_;
 wire _00988_;
 wire _00989_;
 wire _00990_;
 wire _00991_;
 wire _00992_;
 wire _00993_;
 wire _00994_;
 wire _00995_;
 wire _00996_;
 wire _00997_;
 wire _00998_;
 wire _00999_;
 wire _01000_;
 wire _01001_;
 wire _01002_;
 wire _01003_;
 wire _01004_;
 wire _01005_;
 wire _01006_;
 wire _01007_;
 wire _01008_;
 wire _01009_;
 wire _01010_;
 wire _01011_;
 wire _01012_;
 wire _01013_;
 wire _01014_;
 wire _01015_;
 wire _01016_;
 wire _01017_;
 wire _01018_;
 wire _01019_;
 wire _01020_;
 wire _01021_;
 wire _01022_;
 wire _01023_;
 wire _01024_;
 wire _01025_;
 wire _01026_;
 wire _01027_;
 wire _01028_;
 wire _01029_;
 wire _01030_;
 wire _01031_;
 wire _01032_;
 wire _01033_;
 wire _01034_;
 wire _01035_;
 wire _01036_;
 wire _01037_;
 wire _01038_;
 wire _01039_;
 wire _01040_;
 wire _01041_;
 wire _01042_;
 wire _01043_;
 wire _01044_;
 wire _01045_;
 wire _01046_;
 wire _01047_;
 wire _01048_;
 wire _01049_;
 wire _01050_;
 wire _01051_;
 wire _01052_;
 wire _01053_;
 wire _01054_;
 wire _01055_;
 wire _01056_;
 wire _01057_;
 wire _01058_;
 wire _01059_;
 wire _01060_;
 wire _01061_;
 wire _01062_;
 wire _01063_;
 wire _01064_;
 wire _01065_;
 wire _01066_;
 wire _01067_;
 wire _01068_;
 wire _01069_;
 wire _01070_;
 wire _01071_;
 wire _01072_;
 wire _01073_;
 wire _01074_;
 wire _01075_;
 wire _01076_;
 wire _01077_;
 wire _01078_;
 wire _01079_;
 wire _01080_;
 wire _01081_;
 wire _01082_;
 wire _01083_;
 wire _01084_;
 wire _01085_;
 wire _01086_;
 wire _01087_;
 wire _01088_;
 wire _01089_;
 wire _01090_;
 wire _01091_;
 wire _01092_;
 wire _01093_;
 wire _01094_;
 wire _01095_;
 wire _01096_;
 wire _01097_;
 wire _01098_;
 wire _01099_;
 wire _01100_;
 wire _01101_;
 wire _01102_;
 wire _01103_;
 wire _01104_;
 wire _01105_;
 wire _01106_;
 wire _01107_;
 wire _01108_;
 wire _01109_;
 wire _01110_;
 wire _01111_;
 wire _01112_;
 wire _01113_;
 wire _01114_;
 wire _01115_;
 wire _01116_;
 wire _01117_;
 wire _01118_;
 wire _01119_;
 wire _01120_;
 wire _01121_;
 wire _01122_;
 wire _01123_;
 wire _01124_;
 wire _01125_;
 wire _01126_;
 wire _01127_;
 wire _01128_;
 wire _01129_;
 wire _01130_;
 wire _01131_;
 wire _01132_;
 wire _01133_;
 wire _01134_;
 wire _01135_;
 wire _01136_;
 wire _01137_;
 wire _01138_;
 wire _01139_;
 wire _01140_;
 wire _01141_;
 wire _01142_;
 wire _01143_;
 wire _01144_;
 wire _01145_;
 wire _01146_;
 wire _01147_;
 wire _01148_;
 wire _01149_;
 wire _01150_;
 wire _01151_;
 wire _01152_;
 wire _01153_;
 wire _01154_;
 wire _01155_;
 wire _01156_;
 wire _01157_;
 wire _01158_;
 wire _01159_;
 wire _01160_;
 wire _01161_;
 wire _01162_;
 wire _01163_;
 wire _01164_;
 wire _01165_;
 wire _01166_;
 wire _01167_;
 wire _01168_;
 wire _01169_;
 wire _01170_;
 wire _01171_;
 wire _01172_;
 wire _01173_;
 wire _01174_;
 wire _01175_;
 wire _01176_;
 wire _01177_;
 wire _01178_;
 wire _01179_;
 wire _01180_;
 wire _01181_;
 wire _01182_;
 wire _01183_;
 wire _01184_;
 wire _01185_;
 wire _01186_;
 wire _01187_;
 wire _01188_;
 wire _01189_;
 wire _01190_;
 wire _01191_;
 wire _01192_;
 wire _01193_;
 wire _01194_;
 wire _01195_;
 wire _01196_;
 wire _01197_;
 wire _01198_;
 wire _01199_;
 wire _01200_;
 wire _01201_;
 wire _01202_;
 wire _01203_;
 wire _01204_;
 wire _01205_;
 wire _01206_;
 wire _01207_;
 wire _01208_;
 wire _01209_;
 wire _01210_;
 wire _01211_;
 wire _01212_;
 wire _01213_;
 wire _01214_;
 wire _01215_;
 wire _01216_;
 wire _01217_;
 wire _01218_;
 wire _01219_;
 wire _01220_;
 wire _01221_;
 wire _01222_;
 wire _01223_;
 wire _01224_;
 wire _01225_;
 wire _01226_;
 wire _01227_;
 wire _01228_;
 wire _01229_;
 wire _01230_;
 wire _01231_;
 wire _01232_;
 wire _01233_;
 wire _01234_;
 wire _01235_;
 wire _01236_;
 wire _01237_;
 wire _01238_;
 wire _01239_;
 wire _01240_;
 wire _01241_;
 wire _01242_;
 wire _01243_;
 wire _01244_;
 wire _01245_;
 wire _01246_;
 wire _01247_;
 wire _01248_;
 wire _01249_;
 wire _01250_;
 wire _01251_;
 wire _01252_;
 wire _01253_;
 wire _01254_;
 wire _01255_;
 wire _01256_;
 wire _01257_;
 wire _01258_;
 wire _01259_;
 wire _01260_;
 wire _01261_;
 wire _01262_;
 wire _01263_;
 wire _01264_;
 wire _01265_;
 wire _01266_;
 wire _01267_;
 wire _01268_;
 wire _01269_;
 wire _01270_;
 wire _01271_;
 wire _01272_;
 wire _01273_;
 wire _01274_;
 wire _01275_;
 wire _01276_;
 wire _01277_;
 wire _01278_;
 wire _01279_;
 wire _01280_;
 wire _01281_;
 wire _01282_;
 wire _01283_;
 wire _01284_;
 wire _01285_;
 wire _01286_;
 wire _01287_;
 wire _01288_;
 wire _01289_;
 wire _01290_;
 wire _01291_;
 wire _01292_;
 wire _01293_;
 wire _01294_;
 wire _01295_;
 wire _01296_;
 wire _01297_;
 wire _01298_;
 wire _01299_;
 wire _01300_;
 wire _01301_;
 wire _01302_;
 wire _01303_;
 wire _01304_;
 wire _01305_;
 wire _01306_;
 wire _01307_;
 wire _01308_;
 wire _01309_;
 wire _01310_;
 wire _01311_;
 wire _01312_;
 wire _01313_;
 wire _01314_;
 wire _01315_;
 wire _01316_;
 wire _01317_;
 wire _01318_;
 wire _01319_;
 wire _01320_;
 wire _01321_;
 wire _01322_;
 wire _01323_;
 wire _01324_;
 wire _01325_;
 wire _01326_;
 wire _01327_;
 wire _01328_;
 wire _01329_;
 wire _01330_;
 wire _01331_;
 wire _01332_;
 wire _01333_;
 wire _01334_;
 wire _01335_;
 wire _01336_;
 wire _01337_;
 wire _01338_;
 wire _01339_;
 wire _01340_;
 wire _01341_;
 wire _01342_;
 wire _01343_;
 wire _01344_;
 wire _01345_;
 wire _01346_;
 wire _01347_;
 wire _01348_;
 wire _01349_;
 wire _01350_;
 wire _01351_;
 wire _01352_;
 wire _01353_;
 wire _01354_;
 wire _01355_;
 wire _01356_;
 wire _01357_;
 wire _01358_;
 wire _01359_;
 wire _01360_;
 wire _01361_;
 wire _01362_;
 wire _01363_;
 wire _01364_;
 wire _01365_;
 wire _01366_;
 wire _01367_;
 wire _01368_;
 wire _01369_;
 wire _01370_;
 wire _01371_;
 wire _01372_;
 wire _01373_;
 wire _01374_;
 wire _01375_;
 wire _01376_;
 wire _01377_;
 wire _01378_;
 wire _01379_;
 wire _01380_;
 wire _01381_;
 wire _01382_;
 wire _01383_;
 wire _01384_;
 wire _01385_;
 wire _01386_;
 wire _01387_;
 wire _01388_;
 wire _01389_;
 wire _01390_;
 wire _01391_;
 wire _01392_;
 wire _01393_;
 wire _01394_;
 wire _01395_;
 wire _01396_;
 wire _01397_;
 wire _01398_;
 wire _01399_;
 wire _01400_;
 wire _01401_;
 wire _01402_;
 wire _01403_;
 wire _01404_;
 wire _01405_;
 wire _01406_;
 wire _01407_;
 wire _01408_;
 wire _01409_;
 wire _01410_;
 wire _01411_;
 wire _01412_;
 wire _01413_;
 wire _01414_;
 wire _01415_;
 wire _01416_;
 wire _01417_;
 wire _01418_;
 wire _01419_;
 wire _01420_;
 wire _01421_;
 wire _01422_;
 wire _01423_;
 wire _01424_;
 wire _01425_;
 wire _01426_;
 wire _01427_;
 wire _01428_;
 wire _01429_;
 wire _01430_;
 wire _01431_;
 wire _01432_;
 wire _01433_;
 wire _01434_;
 wire _01435_;
 wire _01436_;
 wire _01437_;
 wire _01438_;
 wire _01439_;
 wire _01440_;
 wire _01441_;
 wire _01442_;
 wire _01443_;
 wire _01444_;
 wire _01445_;
 wire _01446_;
 wire _01447_;
 wire _01448_;
 wire _01449_;
 wire _01450_;
 wire _01451_;
 wire _01452_;
 wire _01453_;
 wire _01454_;
 wire _01455_;
 wire _01456_;
 wire _01457_;
 wire _01458_;
 wire _01459_;
 wire _01460_;
 wire _01461_;
 wire _01462_;
 wire _01463_;
 wire _01464_;
 wire _01465_;
 wire _01466_;
 wire _01467_;
 wire _01468_;
 wire _01469_;
 wire _01470_;
 wire _01471_;
 wire _01472_;
 wire _01473_;
 wire _01474_;
 wire _01475_;
 wire _01476_;
 wire _01477_;
 wire _01478_;
 wire _01479_;
 wire _01480_;
 wire _01481_;
 wire _01482_;
 wire _01483_;
 wire _01484_;
 wire _01485_;
 wire _01486_;
 wire _01487_;
 wire _01488_;
 wire _01489_;
 wire _01490_;
 wire _01491_;
 wire _01492_;
 wire _01493_;
 wire _01494_;
 wire _01495_;
 wire _01496_;
 wire _01497_;
 wire _01498_;
 wire _01499_;
 wire _01500_;
 wire _01501_;
 wire _01502_;
 wire _01503_;
 wire _01504_;
 wire _01505_;
 wire _01506_;
 wire _01507_;
 wire _01508_;
 wire _01509_;
 wire _01510_;
 wire _01511_;
 wire _01512_;
 wire _01513_;
 wire _01514_;
 wire _01515_;
 wire _01516_;
 wire _01517_;
 wire _01518_;
 wire _01519_;
 wire _01520_;
 wire _01521_;
 wire _01522_;
 wire _01523_;
 wire _01524_;
 wire _01525_;
 wire _01526_;
 wire _01527_;
 wire _01528_;
 wire _01529_;
 wire _01530_;
 wire _01531_;
 wire _01532_;
 wire _01533_;
 wire _01534_;
 wire _01535_;
 wire _01536_;
 wire _01537_;
 wire _01538_;
 wire _01539_;
 wire _01540_;
 wire _01541_;
 wire _01542_;
 wire _01543_;
 wire _01544_;
 wire _01545_;
 wire _01546_;
 wire _01547_;
 wire _01548_;
 wire _01549_;
 wire _01550_;
 wire _01551_;
 wire _01552_;
 wire _01553_;
 wire _01554_;
 wire _01555_;
 wire _01556_;
 wire _01557_;
 wire _01558_;
 wire _01559_;
 wire _01560_;
 wire _01561_;
 wire _01562_;
 wire _01563_;
 wire _01564_;
 wire _01565_;
 wire _01566_;
 wire _01567_;
 wire _01568_;
 wire _01569_;
 wire _01570_;
 wire _01571_;
 wire _01572_;
 wire _01573_;
 wire _01574_;
 wire _01575_;
 wire _01576_;
 wire _01577_;
 wire _01578_;
 wire _01579_;
 wire _01580_;
 wire _01581_;
 wire _01582_;
 wire _01583_;
 wire _01584_;
 wire _01585_;
 wire _01586_;
 wire _01587_;
 wire _01588_;
 wire _01589_;
 wire _01590_;
 wire _01591_;
 wire _01592_;
 wire _01593_;
 wire _01594_;
 wire _01595_;
 wire _01596_;
 wire _01597_;
 wire _01598_;
 wire _01599_;
 wire _01600_;
 wire _01601_;
 wire _01602_;
 wire _01603_;
 wire _01604_;
 wire _01605_;
 wire _01606_;
 wire _01607_;
 wire _01608_;
 wire _01609_;
 wire _01610_;
 wire _01611_;
 wire _01612_;
 wire _01613_;
 wire _01614_;
 wire _01615_;
 wire _01616_;
 wire _01617_;
 wire _01618_;
 wire _01619_;
 wire _01620_;
 wire _01621_;
 wire _01622_;
 wire _01623_;
 wire _01624_;
 wire _01625_;
 wire _01626_;
 wire _01627_;
 wire _01628_;
 wire _01629_;
 wire _01630_;
 wire _01631_;
 wire _01632_;
 wire _01633_;
 wire _01634_;
 wire _01635_;
 wire _01636_;
 wire _01637_;
 wire _01638_;
 wire _01639_;
 wire _01640_;
 wire _01641_;
 wire _01642_;
 wire _01643_;
 wire _01644_;
 wire _01645_;
 wire _01646_;
 wire _01647_;
 wire _01648_;
 wire _01649_;
 wire _01650_;
 wire _01651_;
 wire _01652_;
 wire _01653_;
 wire _01654_;
 wire _01655_;
 wire _01656_;
 wire _01657_;
 wire _01658_;
 wire _01659_;
 wire _01660_;
 wire _01661_;
 wire _01662_;
 wire _01663_;
 wire _01664_;
 wire _01665_;
 wire _01666_;
 wire _01667_;
 wire _01668_;
 wire _01669_;
 wire _01670_;
 wire _01671_;
 wire _01672_;
 wire _01673_;
 wire _01674_;
 wire _01675_;
 wire _01676_;
 wire _01677_;
 wire _01678_;
 wire _01679_;
 wire _01680_;
 wire _01681_;
 wire _01682_;
 wire _01683_;
 wire _01684_;
 wire _01685_;
 wire _01686_;
 wire _01687_;
 wire _01688_;
 wire _01689_;
 wire _01690_;
 wire _01691_;
 wire _01692_;
 wire _01693_;
 wire _01694_;
 wire _01695_;
 wire _01696_;
 wire _01697_;
 wire _01698_;
 wire _01699_;
 wire _01700_;
 wire _01701_;
 wire _01702_;
 wire _01703_;
 wire _01704_;
 wire _01705_;
 wire _01706_;
 wire _01707_;
 wire _01708_;
 wire _01709_;
 wire _01710_;
 wire _01711_;
 wire _01712_;
 wire _01713_;
 wire _01714_;
 wire _01715_;
 wire _01716_;
 wire _01717_;
 wire _01718_;
 wire _01719_;
 wire _01720_;
 wire _01721_;
 wire _01722_;
 wire _01723_;
 wire _01724_;
 wire _01725_;
 wire _01726_;
 wire _01727_;
 wire _01728_;
 wire _01729_;
 wire _01730_;
 wire _01731_;
 wire _01732_;
 wire _01733_;
 wire _01734_;
 wire _01735_;
 wire _01736_;
 wire _01737_;
 wire _01738_;
 wire _01739_;
 wire _01740_;
 wire _01741_;
 wire _01742_;
 wire _01743_;
 wire _01744_;
 wire _01745_;
 wire _01746_;
 wire _01747_;
 wire _01748_;
 wire _01749_;
 wire _01750_;
 wire _01751_;
 wire _01752_;
 wire _01753_;
 wire _01754_;
 wire _01755_;
 wire _01756_;
 wire _01757_;
 wire _01758_;
 wire _01759_;
 wire _01760_;
 wire _01761_;
 wire _01762_;
 wire _01763_;
 wire _01764_;
 wire _01765_;
 wire _01766_;
 wire _01767_;
 wire _01768_;
 wire _01769_;
 wire _01770_;
 wire _01771_;
 wire _01772_;
 wire _01773_;
 wire _01774_;
 wire _01775_;
 wire _01776_;
 wire _01777_;
 wire _01778_;
 wire _01779_;
 wire _01780_;
 wire _01781_;
 wire _01782_;
 wire _01783_;
 wire _01784_;
 wire _01785_;
 wire _01786_;
 wire _01787_;
 wire _01788_;
 wire _01789_;
 wire _01790_;
 wire _01791_;
 wire _01792_;
 wire _01793_;
 wire _01794_;
 wire _01795_;
 wire _01796_;
 wire _01797_;
 wire _01798_;
 wire _01799_;
 wire _01800_;
 wire _01801_;
 wire _01802_;
 wire _01803_;
 wire _01804_;
 wire _01805_;
 wire _01806_;
 wire _01807_;
 wire _01808_;
 wire _01809_;
 wire _01810_;
 wire _01811_;
 wire _01812_;
 wire _01813_;
 wire _01814_;
 wire _01815_;
 wire _01816_;
 wire _01817_;
 wire _01818_;
 wire _01819_;
 wire _01820_;
 wire _01821_;
 wire _01822_;
 wire _01823_;
 wire _01824_;
 wire _01825_;
 wire _01826_;
 wire _01827_;
 wire _01828_;
 wire _01829_;
 wire _01830_;
 wire _01831_;
 wire _01832_;
 wire _01833_;
 wire _01834_;
 wire _01835_;
 wire _01836_;
 wire _01837_;
 wire _01838_;
 wire _01839_;
 wire _01840_;
 wire _01841_;
 wire _01842_;
 wire _01843_;
 wire _01844_;
 wire _01845_;
 wire _01846_;
 wire _01847_;
 wire _01848_;
 wire _01849_;
 wire _01850_;
 wire _01851_;
 wire _01852_;
 wire _01853_;
 wire _01854_;
 wire _01855_;
 wire _01856_;
 wire _01857_;
 wire _01858_;
 wire _01859_;
 wire _01860_;
 wire _01861_;
 wire _01862_;
 wire _01863_;
 wire _01864_;
 wire _01865_;
 wire _01866_;
 wire _01867_;
 wire _01868_;
 wire _01869_;
 wire _01870_;
 wire _01871_;
 wire _01872_;
 wire _01873_;
 wire _01874_;
 wire _01875_;
 wire _01876_;
 wire _01877_;
 wire _01878_;
 wire _01879_;
 wire _01880_;
 wire _01881_;
 wire _01882_;
 wire _01883_;
 wire _01884_;
 wire _01885_;
 wire _01886_;
 wire _01887_;
 wire _01888_;
 wire _01889_;
 wire _01890_;
 wire _01891_;
 wire _01892_;
 wire _01893_;
 wire _01894_;
 wire _01895_;
 wire _01896_;
 wire _01897_;
 wire _01898_;
 wire _01899_;
 wire _01900_;
 wire _01901_;
 wire _01902_;
 wire _01903_;
 wire _01904_;
 wire _01905_;
 wire _01906_;
 wire _01907_;
 wire _01908_;
 wire _01909_;
 wire _01910_;
 wire _01911_;
 wire _01912_;
 wire _01913_;
 wire _01914_;
 wire _01915_;
 wire _01916_;
 wire _01917_;
 wire _01918_;
 wire _01919_;
 wire _01920_;
 wire _01921_;
 wire _01922_;
 wire _01923_;
 wire _01924_;
 wire _01925_;
 wire _01926_;
 wire _01927_;
 wire _01928_;
 wire _01929_;
 wire _01930_;
 wire _01931_;
 wire _01932_;
 wire _01933_;
 wire _01934_;
 wire _01935_;
 wire _01936_;
 wire _01937_;
 wire _01938_;
 wire _01939_;
 wire _01940_;
 wire _01941_;
 wire _01942_;
 wire _01943_;
 wire _01944_;
 wire _01945_;
 wire _01946_;
 wire _01947_;
 wire _01948_;
 wire _01949_;
 wire _01950_;
 wire _01951_;
 wire _01952_;
 wire _01953_;
 wire _01954_;
 wire _01955_;
 wire _01956_;
 wire _01957_;
 wire _01958_;
 wire _01959_;
 wire _01960_;
 wire _01961_;
 wire _01962_;
 wire _01963_;
 wire _01964_;
 wire _01965_;
 wire _01966_;
 wire _01967_;
 wire _01968_;
 wire _01969_;
 wire _01970_;
 wire _01971_;
 wire _01972_;
 wire _01973_;
 wire _01974_;
 wire _01975_;
 wire _01976_;
 wire _01977_;
 wire _01978_;
 wire _01979_;
 wire _01980_;
 wire _01981_;
 wire _01982_;
 wire _01983_;
 wire _01984_;
 wire _01985_;
 wire _01986_;
 wire _01987_;
 wire _01988_;
 wire _01989_;
 wire _01990_;
 wire _01991_;
 wire _01992_;
 wire _01993_;
 wire _01994_;
 wire _01995_;
 wire _01996_;
 wire _01997_;
 wire _01998_;
 wire _01999_;
 wire _02000_;
 wire _02001_;
 wire _02002_;
 wire _02003_;
 wire _02004_;
 wire _02005_;
 wire _02006_;
 wire _02007_;
 wire _02008_;
 wire _02009_;
 wire _02010_;
 wire _02011_;
 wire _02012_;
 wire _02013_;
 wire _02014_;
 wire _02015_;
 wire _02016_;
 wire _02017_;
 wire _02018_;
 wire _02019_;
 wire _02020_;
 wire _02021_;
 wire _02022_;
 wire _02023_;
 wire _02024_;
 wire _02025_;
 wire _02026_;
 wire _02027_;
 wire _02028_;
 wire _02029_;
 wire _02030_;
 wire _02031_;
 wire _02032_;
 wire _02033_;
 wire _02034_;
 wire _02035_;
 wire _02036_;
 wire _02037_;
 wire _02038_;
 wire _02039_;
 wire _02040_;
 wire _02041_;
 wire _02042_;
 wire _02043_;
 wire _02044_;
 wire _02045_;
 wire _02046_;
 wire _02047_;
 wire _02048_;
 wire _02049_;
 wire _02050_;
 wire _02051_;
 wire _02052_;
 wire _02053_;
 wire _02054_;
 wire _02055_;
 wire _02056_;
 wire _02057_;
 wire _02058_;
 wire _02059_;
 wire _02060_;
 wire _02061_;
 wire _02062_;
 wire _02063_;
 wire _02064_;
 wire _02065_;
 wire _02066_;
 wire _02067_;
 wire _02068_;
 wire _02069_;
 wire _02070_;
 wire _02071_;
 wire _02072_;
 wire _02073_;
 wire _02074_;
 wire _02075_;
 wire _02076_;
 wire _02077_;
 wire _02078_;
 wire _02079_;
 wire _02080_;
 wire _02081_;
 wire _02082_;
 wire _02083_;
 wire _02084_;
 wire _02085_;
 wire _02086_;
 wire _02087_;
 wire _02088_;
 wire _02089_;
 wire _02090_;
 wire _02091_;
 wire _02092_;
 wire _02093_;
 wire _02094_;
 wire _02095_;
 wire _02096_;
 wire _02097_;
 wire _02098_;
 wire _02099_;
 wire _02100_;
 wire _02101_;
 wire _02102_;
 wire _02103_;
 wire _02104_;
 wire _02105_;
 wire _02106_;
 wire _02107_;
 wire _02108_;
 wire _02109_;
 wire _02110_;
 wire _02111_;
 wire _02112_;
 wire _02113_;
 wire _02114_;
 wire _02115_;
 wire _02116_;
 wire _02117_;
 wire _02118_;
 wire _02119_;
 wire _02120_;
 wire _02121_;
 wire _02122_;
 wire _02123_;
 wire _02124_;
 wire _02125_;
 wire _02126_;
 wire _02127_;
 wire _02128_;
 wire _02129_;
 wire _02130_;
 wire _02131_;
 wire _02132_;
 wire _02133_;
 wire _02134_;
 wire _02135_;
 wire _02136_;
 wire _02137_;
 wire _02138_;
 wire _02139_;
 wire _02140_;
 wire _02141_;
 wire _02142_;
 wire _02143_;
 wire _02144_;
 wire _02145_;
 wire _02146_;
 wire _02147_;
 wire _02148_;
 wire _02149_;
 wire _02150_;
 wire _02151_;
 wire _02152_;
 wire _02153_;
 wire _02154_;
 wire _02155_;
 wire _02156_;
 wire _02157_;
 wire _02158_;
 wire _02159_;
 wire _02160_;
 wire _02161_;
 wire _02162_;
 wire _02163_;
 wire _02164_;
 wire _02165_;
 wire _02166_;
 wire _02167_;
 wire _02168_;
 wire _02169_;
 wire _02170_;
 wire _02171_;
 wire _02172_;
 wire _02173_;
 wire _02174_;
 wire _02175_;
 wire _02176_;
 wire _02177_;
 wire _02178_;
 wire _02179_;
 wire _02180_;
 wire _02181_;
 wire _02182_;
 wire _02183_;
 wire _02184_;
 wire _02185_;
 wire _02186_;
 wire _02187_;
 wire _02188_;
 wire _02189_;
 wire _02190_;
 wire _02191_;
 wire _02192_;
 wire _02193_;
 wire _02194_;
 wire _02195_;
 wire _02196_;
 wire _02197_;
 wire _02198_;
 wire _02199_;
 wire _02200_;
 wire _02201_;
 wire _02202_;
 wire _02203_;
 wire _02204_;
 wire _02205_;
 wire _02206_;
 wire _02207_;
 wire _02208_;
 wire _02209_;
 wire _02210_;
 wire _02211_;
 wire _02212_;
 wire _02213_;
 wire _02214_;
 wire _02215_;
 wire _02216_;
 wire _02217_;
 wire _02218_;
 wire _02219_;
 wire _02220_;
 wire _02221_;
 wire _02222_;
 wire _02223_;
 wire _02224_;
 wire _02225_;
 wire _02226_;
 wire _02227_;
 wire _02228_;
 wire _02229_;
 wire _02230_;
 wire _02231_;
 wire _02232_;
 wire _02233_;
 wire _02234_;
 wire _02235_;
 wire _02236_;
 wire _02237_;
 wire _02238_;
 wire _02239_;
 wire _02240_;
 wire _02241_;
 wire _02242_;
 wire _02243_;
 wire _02244_;
 wire _02245_;
 wire _02246_;
 wire _02247_;
 wire _02248_;
 wire _02249_;
 wire _02250_;
 wire _02251_;
 wire _02252_;
 wire _02253_;
 wire _02254_;
 wire _02255_;
 wire _02256_;
 wire _02257_;
 wire _02258_;
 wire _02259_;
 wire _02260_;
 wire _02261_;
 wire _02262_;
 wire _02263_;
 wire _02264_;
 wire _02265_;
 wire _02266_;
 wire _02267_;
 wire _02268_;
 wire _02269_;
 wire _02270_;
 wire _02271_;
 wire _02272_;
 wire _02273_;
 wire _02274_;
 wire _02275_;
 wire _02276_;
 wire _02277_;
 wire _02278_;
 wire _02279_;
 wire _02280_;
 wire _02281_;
 wire _02282_;
 wire _02283_;
 wire _02284_;
 wire _02285_;
 wire _02286_;
 wire _02287_;
 wire _02288_;
 wire _02289_;
 wire _02290_;
 wire _02291_;
 wire _02292_;
 wire _02293_;
 wire _02294_;
 wire _02295_;
 wire _02296_;
 wire _02297_;
 wire _02298_;
 wire _02299_;
 wire _02300_;
 wire _02301_;
 wire _02302_;
 wire _02303_;
 wire _02304_;
 wire _02305_;
 wire _02306_;
 wire _02307_;
 wire _02308_;
 wire _02309_;
 wire _02310_;
 wire _02311_;
 wire _02312_;
 wire _02313_;
 wire _02314_;
 wire _02315_;
 wire _02316_;
 wire _02317_;
 wire _02318_;
 wire _02319_;
 wire _02320_;
 wire _02321_;
 wire _02322_;
 wire _02323_;
 wire _02324_;
 wire _02325_;
 wire _02326_;
 wire _02327_;
 wire _02328_;
 wire _02329_;
 wire _02330_;
 wire _02331_;
 wire _02332_;
 wire _02333_;
 wire _02334_;
 wire _02335_;
 wire _02336_;
 wire _02337_;
 wire _02338_;
 wire _02339_;
 wire _02340_;
 wire _02341_;
 wire _02342_;
 wire _02343_;
 wire _02344_;
 wire _02345_;
 wire _02346_;
 wire _02347_;
 wire _02348_;
 wire _02349_;
 wire _02350_;
 wire _02351_;
 wire _02352_;
 wire _02353_;
 wire _02354_;
 wire _02355_;
 wire _02356_;
 wire _02357_;
 wire _02358_;
 wire _02359_;
 wire _02360_;
 wire _02361_;
 wire _02362_;
 wire _02363_;
 wire _02364_;
 wire _02365_;
 wire _02366_;
 wire _02367_;
 wire _02368_;
 wire _02369_;
 wire _02370_;
 wire _02371_;
 wire _02372_;
 wire _02373_;
 wire _02374_;
 wire _02375_;
 wire _02376_;
 wire _02377_;
 wire _02378_;
 wire _02379_;
 wire _02380_;
 wire _02381_;
 wire _02382_;
 wire _02383_;
 wire _02384_;
 wire _02385_;
 wire _02386_;
 wire _02387_;
 wire _02388_;
 wire _02389_;
 wire _02390_;
 wire _02391_;
 wire _02392_;
 wire _02393_;
 wire _02394_;
 wire _02395_;
 wire _02396_;
 wire _02397_;
 wire _02398_;
 wire _02399_;
 wire _02400_;
 wire _02401_;
 wire _02402_;
 wire _02403_;
 wire _02404_;
 wire _02405_;
 wire _02406_;
 wire _02407_;
 wire _02408_;
 wire _02409_;
 wire _02410_;
 wire _02411_;
 wire _02412_;
 wire _02413_;
 wire _02414_;
 wire _02415_;
 wire _02416_;
 wire _02417_;
 wire _02418_;
 wire _02419_;
 wire _02420_;
 wire _02421_;
 wire _02422_;
 wire _02423_;
 wire _02424_;
 wire _02425_;
 wire _02426_;
 wire _02427_;
 wire _02428_;
 wire _02429_;
 wire _02430_;
 wire _02431_;
 wire _02432_;
 wire _02433_;
 wire _02434_;
 wire _02435_;
 wire _02436_;
 wire _02437_;
 wire _02438_;
 wire _02439_;
 wire _02440_;
 wire _02441_;
 wire _02442_;
 wire _02443_;
 wire _02444_;
 wire _02445_;
 wire _02446_;
 wire _02447_;
 wire _02448_;
 wire _02449_;
 wire _02450_;
 wire _02451_;
 wire _02452_;
 wire _02453_;
 wire _02454_;
 wire _02455_;
 wire _02456_;
 wire _02457_;
 wire _02458_;
 wire _02459_;
 wire _02460_;
 wire _02461_;
 wire _02462_;
 wire _02463_;
 wire _02464_;
 wire _02465_;
 wire _02466_;
 wire _02467_;
 wire _02468_;
 wire _02469_;
 wire _02470_;
 wire _02471_;
 wire _02472_;
 wire _02473_;
 wire _02474_;
 wire _02475_;
 wire _02476_;
 wire _02477_;
 wire _02478_;
 wire _02479_;
 wire _02480_;
 wire _02481_;
 wire _02482_;
 wire _02483_;
 wire _02484_;
 wire _02485_;
 wire _02486_;
 wire _02487_;
 wire _02488_;
 wire _02489_;
 wire _02490_;
 wire _02491_;
 wire _02492_;
 wire _02493_;
 wire _02494_;
 wire _02495_;
 wire _02496_;
 wire _02497_;
 wire _02498_;
 wire _02499_;
 wire _02500_;
 wire _02501_;
 wire _02502_;
 wire _02503_;
 wire _02504_;
 wire _02505_;
 wire _02506_;
 wire _02507_;
 wire _02508_;
 wire _02509_;
 wire _02510_;
 wire _02511_;
 wire _02512_;
 wire _02513_;
 wire _02514_;
 wire _02515_;
 wire _02516_;
 wire _02517_;
 wire _02518_;
 wire _02519_;
 wire _02520_;
 wire _02521_;
 wire _02522_;
 wire _02523_;
 wire _02524_;
 wire _02525_;
 wire _02526_;
 wire _02527_;
 wire _02528_;
 wire _02529_;
 wire _02530_;
 wire _02531_;
 wire _02532_;
 wire _02533_;
 wire _02534_;
 wire _02535_;
 wire _02536_;
 wire _02537_;
 wire _02538_;
 wire _02539_;
 wire _02540_;
 wire _02541_;
 wire _02542_;
 wire _02543_;
 wire _02544_;
 wire _02545_;
 wire _02546_;
 wire _02547_;
 wire _02548_;
 wire _02549_;
 wire _02550_;
 wire _02551_;
 wire _02552_;
 wire _02553_;
 wire _02554_;
 wire _02555_;
 wire _02556_;
 wire _02557_;
 wire _02558_;
 wire _02559_;
 wire _02560_;
 wire _02561_;
 wire _02562_;
 wire _02563_;
 wire _02564_;
 wire _02565_;
 wire _02566_;
 wire _02567_;
 wire _02568_;
 wire _02569_;
 wire _02570_;
 wire _02571_;
 wire _02572_;
 wire _02573_;
 wire _02574_;
 wire _02575_;
 wire _02576_;
 wire _02577_;
 wire _02578_;
 wire _02579_;
 wire _02580_;
 wire _02581_;
 wire _02582_;
 wire _02583_;
 wire _02584_;
 wire _02585_;
 wire _02586_;
 wire _02587_;
 wire _02588_;
 wire _02589_;
 wire _02590_;
 wire _02591_;
 wire _02592_;
 wire _02593_;
 wire _02594_;
 wire _02595_;
 wire _02596_;
 wire _02597_;
 wire _02598_;
 wire _02599_;
 wire _02600_;
 wire _02601_;
 wire _02602_;
 wire _02603_;
 wire _02604_;
 wire _02605_;
 wire _02606_;
 wire _02607_;
 wire _02608_;
 wire _02609_;
 wire _02610_;
 wire _02611_;
 wire _02612_;
 wire _02613_;
 wire _02614_;
 wire _02615_;
 wire _02616_;
 wire _02617_;
 wire _02618_;
 wire _02619_;
 wire _02620_;
 wire _02621_;
 wire _02622_;
 wire _02623_;
 wire _02624_;
 wire _02625_;
 wire _02626_;
 wire _02627_;
 wire _02628_;
 wire _02629_;
 wire _02630_;
 wire _02631_;
 wire _02632_;
 wire _02633_;
 wire _02634_;
 wire _02635_;
 wire _02636_;
 wire _02637_;
 wire _02638_;
 wire _02639_;
 wire _02640_;
 wire _02641_;
 wire _02642_;
 wire _02643_;
 wire _02644_;
 wire _02645_;
 wire _02646_;
 wire _02647_;
 wire _02648_;
 wire _02649_;
 wire _02650_;
 wire _02651_;
 wire _02652_;
 wire _02653_;
 wire _02654_;
 wire _02655_;
 wire _02656_;
 wire _02657_;
 wire _02658_;
 wire _02659_;
 wire _02660_;
 wire _02661_;
 wire _02662_;
 wire _02663_;
 wire _02664_;
 wire _02665_;
 wire _02666_;
 wire _02667_;
 wire _02668_;
 wire _02669_;
 wire _02670_;
 wire _02671_;
 wire _02672_;
 wire _02673_;
 wire _02674_;
 wire _02675_;
 wire _02676_;
 wire _02677_;
 wire _02678_;
 wire _02679_;
 wire _02680_;
 wire _02681_;
 wire _02682_;
 wire _02683_;
 wire _02684_;
 wire _02685_;
 wire _02686_;
 wire _02687_;
 wire _02688_;
 wire _02689_;
 wire _02690_;
 wire _02691_;
 wire _02692_;
 wire _02693_;
 wire _02694_;
 wire _02695_;
 wire _02696_;
 wire _02697_;
 wire _02698_;
 wire _02699_;
 wire _02700_;
 wire _02701_;
 wire _02702_;
 wire _02703_;
 wire _02704_;
 wire _02705_;
 wire _02706_;
 wire _02707_;
 wire _02708_;
 wire _02709_;
 wire _02710_;
 wire _02711_;
 wire _02712_;
 wire _02713_;
 wire _02714_;
 wire _02715_;
 wire _02716_;
 wire _02717_;
 wire _02718_;
 wire _02719_;
 wire _02720_;
 wire _02721_;
 wire _02722_;
 wire _02723_;
 wire _02724_;
 wire _02725_;
 wire _02726_;
 wire _02727_;
 wire _02728_;
 wire _02729_;
 wire _02730_;
 wire _02731_;
 wire _02732_;
 wire _02733_;
 wire _02734_;
 wire _02735_;
 wire _02736_;
 wire _02737_;
 wire _02738_;
 wire _02739_;
 wire _02740_;
 wire _02741_;
 wire _02742_;
 wire _02743_;
 wire _02744_;
 wire _02745_;
 wire _02746_;
 wire _02747_;
 wire _02748_;
 wire _02749_;
 wire _02750_;
 wire _02751_;
 wire _02752_;
 wire _02753_;
 wire _02754_;
 wire _02755_;
 wire _02756_;
 wire _02757_;
 wire _02758_;
 wire _02759_;
 wire _02760_;
 wire _02761_;
 wire _02762_;
 wire _02763_;
 wire _02764_;
 wire _02765_;
 wire _02766_;
 wire _02767_;
 wire _02768_;
 wire _02769_;
 wire _02770_;
 wire _02771_;
 wire _02772_;
 wire _02773_;
 wire _02774_;
 wire _02775_;
 wire _02776_;
 wire _02777_;
 wire _02778_;
 wire _02779_;
 wire _02780_;
 wire _02781_;
 wire _02782_;
 wire _02783_;
 wire _02784_;
 wire _02785_;
 wire _02786_;
 wire _02787_;
 wire _02788_;
 wire _02789_;
 wire _02790_;
 wire _02791_;
 wire _02792_;
 wire _02793_;
 wire _02794_;
 wire _02795_;
 wire _02796_;
 wire _02797_;
 wire _02798_;
 wire _02799_;
 wire _02800_;
 wire _02801_;
 wire _02802_;
 wire _02803_;
 wire _02804_;
 wire _02805_;
 wire _02806_;
 wire _02807_;
 wire _02808_;
 wire _02809_;
 wire _02810_;
 wire _02811_;
 wire _02812_;
 wire _02813_;
 wire _02814_;
 wire _02815_;
 wire _02816_;
 wire _02817_;
 wire _02818_;
 wire _02819_;
 wire _02820_;
 wire _02821_;
 wire _02822_;
 wire _02823_;
 wire _02824_;
 wire _02825_;
 wire _02826_;
 wire _02827_;
 wire _02828_;
 wire _02829_;
 wire _02830_;
 wire _02831_;
 wire _02832_;
 wire _02833_;
 wire _02834_;
 wire _02835_;
 wire _02836_;
 wire _02837_;
 wire _02838_;
 wire _02839_;
 wire _02840_;
 wire _02841_;
 wire _02842_;
 wire _02843_;
 wire _02844_;
 wire _02845_;
 wire _02846_;
 wire _02847_;
 wire _02848_;
 wire _02849_;
 wire _02850_;
 wire _02851_;
 wire _02852_;
 wire _02853_;
 wire _02854_;
 wire _02855_;
 wire _02856_;
 wire _02857_;
 wire _02858_;
 wire _02859_;
 wire _02860_;
 wire _02861_;
 wire _02862_;
 wire _02863_;
 wire _02864_;
 wire _02865_;
 wire _02866_;
 wire _02867_;
 wire _02868_;
 wire _02869_;
 wire _02870_;
 wire _02871_;
 wire _02872_;
 wire _02873_;
 wire _02874_;
 wire _02875_;
 wire _02876_;
 wire _02877_;
 wire _02878_;
 wire _02879_;
 wire _02880_;
 wire _02881_;
 wire _02882_;
 wire _02883_;
 wire _02884_;
 wire _02885_;
 wire _02886_;
 wire _02887_;
 wire _02888_;
 wire _02889_;
 wire _02890_;
 wire _02891_;
 wire _02892_;
 wire _02893_;
 wire _02894_;
 wire _02895_;
 wire _02896_;
 wire _02897_;
 wire _02898_;
 wire _02899_;
 wire _02900_;
 wire _02901_;
 wire _02902_;
 wire _02903_;
 wire _02904_;
 wire _02905_;
 wire _02906_;
 wire _02907_;
 wire _02908_;
 wire _02909_;
 wire _02910_;
 wire _02911_;
 wire _02912_;
 wire _02913_;
 wire _02914_;
 wire _02915_;
 wire _02916_;
 wire _02917_;
 wire _02918_;
 wire _02919_;
 wire _02920_;
 wire _02921_;
 wire _02922_;
 wire _02923_;
 wire _02924_;
 wire _02925_;
 wire _02926_;
 wire _02927_;
 wire _02928_;
 wire _02929_;
 wire _02930_;
 wire _02931_;
 wire _02932_;
 wire _02933_;
 wire _02934_;
 wire _02935_;
 wire _02936_;
 wire _02937_;
 wire _02938_;
 wire _02939_;
 wire _02940_;
 wire _02941_;
 wire _02942_;
 wire _02943_;
 wire _02944_;
 wire _02945_;
 wire _02946_;
 wire _02947_;
 wire _02948_;
 wire _02949_;
 wire _02950_;
 wire _02951_;
 wire _02952_;
 wire _02953_;
 wire _02954_;
 wire _02955_;
 wire _02956_;
 wire _02957_;
 wire _02958_;
 wire _02959_;
 wire _02960_;
 wire _02961_;
 wire _02962_;
 wire _02963_;
 wire _02964_;
 wire _02965_;
 wire _02966_;
 wire _02967_;
 wire _02968_;
 wire _02969_;
 wire _02970_;
 wire _02971_;
 wire _02972_;
 wire _02973_;
 wire _02974_;
 wire _02975_;
 wire _02976_;
 wire _02977_;
 wire _02978_;
 wire _02979_;
 wire _02980_;
 wire _02981_;
 wire _02982_;
 wire _02983_;
 wire _02984_;
 wire _02985_;
 wire _02986_;
 wire _02987_;
 wire _02988_;
 wire _02989_;
 wire _02990_;
 wire _02991_;
 wire _02992_;
 wire _02993_;
 wire _02994_;
 wire _02995_;
 wire _02996_;
 wire _02997_;
 wire _02998_;
 wire _02999_;
 wire _03000_;
 wire _03001_;
 wire _03002_;
 wire _03003_;
 wire _03004_;
 wire _03005_;
 wire _03006_;
 wire _03007_;
 wire _03008_;
 wire _03009_;
 wire _03010_;
 wire _03011_;
 wire _03012_;
 wire _03013_;
 wire _03014_;
 wire _03015_;
 wire _03016_;
 wire _03017_;
 wire _03018_;
 wire _03019_;
 wire _03020_;
 wire _03021_;
 wire _03022_;
 wire _03023_;
 wire _03024_;
 wire _03025_;
 wire _03026_;
 wire _03027_;
 wire _03028_;
 wire _03029_;
 wire _03030_;
 wire _03031_;
 wire _03032_;
 wire _03033_;
 wire _03034_;
 wire _03035_;
 wire _03036_;
 wire _03037_;
 wire _03038_;
 wire _03039_;
 wire _03040_;
 wire _03041_;
 wire _03042_;
 wire _03043_;
 wire _03044_;
 wire _03045_;
 wire _03046_;
 wire _03047_;
 wire _03048_;
 wire _03049_;
 wire _03050_;
 wire _03051_;
 wire _03052_;
 wire _03053_;
 wire _03054_;
 wire _03055_;
 wire _03056_;
 wire _03057_;
 wire _03058_;
 wire _03059_;
 wire _03060_;
 wire _03061_;
 wire _03062_;
 wire _03063_;
 wire _03064_;
 wire _03065_;
 wire _03066_;
 wire _03067_;
 wire _03068_;
 wire _03069_;
 wire _03070_;
 wire _03071_;
 wire _03072_;
 wire _03073_;
 wire _03074_;
 wire _03075_;
 wire _03076_;
 wire _03077_;
 wire _03078_;
 wire _03079_;
 wire _03080_;
 wire _03081_;
 wire _03082_;
 wire _03083_;
 wire _03084_;
 wire _03085_;
 wire _03086_;
 wire _03087_;
 wire _03088_;
 wire _03089_;
 wire _03090_;
 wire _03091_;
 wire _03092_;
 wire _03093_;
 wire _03094_;
 wire _03095_;
 wire _03096_;
 wire _03097_;
 wire _03098_;
 wire _03099_;
 wire _03100_;
 wire _03101_;
 wire _03102_;
 wire _03103_;
 wire _03104_;
 wire _03105_;
 wire _03106_;
 wire _03107_;
 wire _03108_;
 wire _03109_;
 wire _03110_;
 wire _03111_;
 wire _03112_;
 wire _03113_;
 wire _03114_;
 wire _03115_;
 wire _03116_;
 wire _03117_;
 wire _03118_;
 wire _03119_;
 wire _03120_;
 wire _03121_;
 wire _03122_;
 wire _03123_;
 wire _03124_;
 wire _03125_;
 wire _03126_;
 wire _03127_;
 wire _03128_;
 wire _03129_;
 wire _03130_;
 wire _03131_;
 wire _03132_;
 wire _03133_;
 wire _03134_;
 wire _03135_;
 wire _03136_;
 wire _03137_;
 wire _03138_;
 wire _03139_;
 wire _03140_;
 wire _03141_;
 wire _03142_;
 wire _03143_;
 wire _03144_;
 wire _03145_;
 wire _03146_;
 wire _03147_;
 wire _03148_;
 wire _03149_;
 wire _03150_;
 wire _03151_;
 wire _03152_;
 wire _03153_;
 wire _03154_;
 wire _03155_;
 wire _03156_;
 wire _03157_;
 wire _03158_;
 wire _03159_;
 wire _03160_;
 wire _03161_;
 wire _03162_;
 wire _03163_;
 wire _03164_;
 wire _03165_;
 wire _03166_;
 wire _03167_;
 wire _03168_;
 wire _03169_;
 wire _03170_;
 wire _03171_;
 wire _03172_;
 wire _03173_;
 wire _03174_;
 wire _03175_;
 wire _03176_;
 wire _03177_;
 wire _03178_;
 wire _03179_;
 wire _03180_;
 wire _03181_;
 wire _03182_;
 wire _03183_;
 wire _03184_;
 wire _03185_;
 wire _03186_;
 wire _03187_;
 wire _03188_;
 wire _03189_;
 wire _03190_;
 wire _03191_;
 wire _03192_;
 wire _03193_;
 wire _03194_;
 wire _03195_;
 wire _03196_;
 wire _03197_;
 wire _03198_;
 wire _03199_;
 wire _03200_;
 wire _03201_;
 wire _03202_;
 wire _03203_;
 wire _03204_;
 wire _03205_;
 wire _03206_;
 wire _03207_;
 wire _03208_;
 wire _03209_;
 wire _03210_;
 wire _03211_;
 wire _03212_;
 wire _03213_;
 wire _03214_;
 wire _03215_;
 wire _03216_;
 wire _03217_;
 wire _03218_;
 wire _03219_;
 wire _03220_;
 wire _03221_;
 wire _03222_;
 wire _03223_;
 wire _03224_;
 wire _03225_;
 wire _03226_;
 wire _03227_;
 wire _03228_;
 wire _03229_;
 wire _03230_;
 wire _03231_;
 wire _03232_;
 wire _03233_;
 wire _03234_;
 wire _03235_;
 wire _03236_;
 wire _03237_;
 wire _03238_;
 wire _03239_;
 wire _03240_;
 wire _03241_;
 wire _03242_;
 wire _03243_;
 wire _03244_;
 wire _03245_;
 wire _03246_;
 wire _03247_;
 wire _03248_;
 wire _03249_;
 wire _03250_;
 wire _03251_;
 wire _03252_;
 wire _03253_;
 wire _03254_;
 wire _03255_;
 wire _03256_;
 wire _03257_;
 wire _03258_;
 wire _03259_;
 wire _03260_;
 wire _03261_;
 wire _03262_;
 wire _03263_;
 wire _03264_;
 wire _03265_;
 wire _03266_;
 wire _03267_;
 wire _03268_;
 wire _03269_;
 wire _03270_;
 wire _03271_;
 wire _03272_;
 wire _03273_;
 wire _03274_;
 wire _03275_;
 wire _03276_;
 wire _03277_;
 wire _03278_;
 wire _03279_;
 wire _03280_;
 wire _03281_;
 wire _03282_;
 wire _03283_;
 wire _03284_;
 wire _03285_;
 wire _03286_;
 wire _03287_;
 wire _03288_;
 wire _03289_;
 wire _03290_;
 wire _03291_;
 wire _03292_;
 wire _03293_;
 wire _03294_;
 wire _03295_;
 wire _03296_;
 wire _03297_;
 wire _03298_;
 wire _03299_;
 wire _03300_;
 wire _03301_;
 wire _03302_;
 wire _03303_;
 wire _03304_;
 wire _03305_;
 wire _03306_;
 wire _03307_;
 wire _03308_;
 wire _03309_;
 wire _03310_;
 wire _03311_;
 wire _03312_;
 wire _03313_;
 wire _03314_;
 wire _03315_;
 wire _03316_;
 wire _03317_;
 wire _03318_;
 wire _03319_;
 wire _03320_;
 wire _03321_;
 wire _03322_;
 wire _03323_;
 wire _03324_;
 wire _03325_;
 wire _03326_;
 wire _03327_;
 wire _03328_;
 wire _03329_;
 wire _03330_;
 wire _03331_;
 wire _03332_;
 wire _03333_;
 wire _03334_;
 wire _03335_;
 wire _03336_;
 wire _03337_;
 wire _03338_;
 wire _03339_;
 wire _03340_;
 wire _03341_;
 wire _03342_;
 wire _03343_;
 wire _03344_;
 wire _03345_;
 wire _03346_;
 wire _03347_;
 wire _03348_;
 wire _03349_;
 wire _03350_;
 wire _03351_;
 wire _03352_;
 wire _03353_;
 wire _03354_;
 wire _03355_;
 wire _03356_;
 wire _03357_;
 wire _03358_;
 wire _03359_;
 wire _03360_;
 wire _03361_;
 wire _03362_;
 wire _03363_;
 wire _03364_;
 wire _03365_;
 wire _03366_;
 wire _03367_;
 wire _03368_;
 wire _03369_;
 wire _03370_;
 wire _03371_;
 wire _03372_;
 wire _03373_;
 wire _03374_;
 wire _03375_;
 wire _03376_;
 wire _03377_;
 wire _03378_;
 wire _03379_;
 wire _03380_;
 wire _03381_;
 wire _03382_;
 wire _03383_;
 wire _03384_;
 wire _03385_;
 wire _03386_;
 wire _03387_;
 wire _03388_;
 wire _03389_;
 wire _03390_;
 wire _03391_;
 wire _03392_;
 wire _03393_;
 wire _03394_;
 wire _03395_;
 wire _03396_;
 wire _03397_;
 wire _03398_;
 wire _03399_;
 wire _03400_;
 wire _03401_;
 wire _03402_;
 wire _03403_;
 wire _03404_;
 wire _03405_;
 wire _03406_;
 wire _03407_;
 wire _03408_;
 wire _03409_;
 wire _03410_;
 wire _03411_;
 wire _03412_;
 wire _03413_;
 wire _03414_;
 wire _03415_;
 wire _03416_;
 wire _03417_;
 wire _03418_;
 wire _03419_;
 wire _03420_;
 wire _03421_;
 wire _03422_;
 wire _03423_;
 wire _03424_;
 wire _03425_;
 wire _03426_;
 wire _03427_;
 wire _03428_;
 wire _03429_;
 wire _03430_;
 wire _03431_;
 wire _03432_;
 wire _03433_;
 wire _03434_;
 wire _03435_;
 wire _03436_;
 wire _03437_;
 wire _03438_;
 wire _03439_;
 wire _03440_;
 wire _03441_;
 wire _03442_;
 wire _03443_;
 wire _03444_;
 wire _03445_;
 wire _03446_;
 wire _03447_;
 wire _03448_;
 wire _03449_;
 wire _03450_;
 wire _03451_;
 wire _03452_;
 wire _03453_;
 wire _03454_;
 wire _03455_;
 wire _03456_;
 wire _03457_;
 wire _03458_;
 wire _03459_;
 wire _03460_;
 wire _03461_;
 wire _03462_;
 wire _03463_;
 wire _03464_;
 wire _03465_;
 wire _03466_;
 wire _03467_;
 wire _03468_;
 wire _03469_;
 wire _03470_;
 wire _03471_;
 wire _03472_;
 wire _03473_;
 wire _03474_;
 wire _03475_;
 wire _03476_;
 wire _03477_;
 wire _03478_;
 wire _03479_;
 wire _03480_;
 wire _03481_;
 wire _03482_;
 wire _03483_;
 wire _03484_;
 wire _03485_;
 wire _03486_;
 wire _03487_;
 wire _03488_;
 wire _03489_;
 wire _03490_;
 wire _03491_;
 wire _03492_;
 wire _03493_;
 wire _03494_;
 wire _03495_;
 wire _03496_;
 wire _03497_;
 wire _03498_;
 wire _03499_;
 wire _03500_;
 wire _03501_;
 wire _03502_;
 wire _03503_;
 wire _03504_;
 wire _03505_;
 wire _03506_;
 wire _03507_;
 wire _03508_;
 wire _03509_;
 wire _03510_;
 wire _03511_;
 wire _03512_;
 wire _03513_;
 wire _03514_;
 wire _03515_;
 wire _03516_;
 wire _03517_;
 wire _03518_;
 wire _03519_;
 wire _03520_;
 wire _03521_;
 wire _03522_;
 wire _03523_;
 wire _03524_;
 wire _03525_;
 wire _03526_;
 wire _03527_;
 wire _03528_;
 wire _03529_;
 wire _03530_;
 wire _03531_;
 wire _03532_;
 wire _03533_;
 wire _03534_;
 wire _03535_;
 wire _03536_;
 wire _03537_;
 wire _03538_;
 wire _03539_;
 wire _03540_;
 wire _03541_;
 wire _03542_;
 wire _03543_;
 wire _03544_;
 wire _03545_;
 wire _03546_;
 wire _03547_;
 wire _03548_;
 wire _03549_;
 wire _03550_;
 wire _03551_;
 wire _03552_;
 wire _03553_;
 wire _03554_;
 wire _03555_;
 wire _03556_;
 wire _03557_;
 wire _03558_;
 wire _03559_;
 wire _03560_;
 wire _03561_;
 wire _03562_;
 wire _03563_;
 wire _03564_;
 wire _03565_;
 wire _03566_;
 wire _03567_;
 wire _03568_;
 wire _03569_;
 wire _03570_;
 wire _03571_;
 wire _03572_;
 wire _03573_;
 wire _03574_;
 wire _03575_;
 wire _03576_;
 wire _03577_;
 wire _03578_;
 wire _03579_;
 wire _03580_;
 wire _03581_;
 wire _03582_;
 wire _03583_;
 wire _03584_;
 wire _03585_;
 wire _03586_;
 wire _03587_;
 wire _03588_;
 wire _03589_;
 wire _03590_;
 wire _03591_;
 wire _03592_;
 wire _03593_;
 wire _03594_;
 wire _03595_;
 wire _03596_;
 wire _03597_;
 wire _03598_;
 wire _03599_;
 wire _03600_;
 wire _03601_;
 wire _03602_;
 wire _03603_;
 wire _03604_;
 wire _03605_;
 wire _03606_;
 wire _03607_;
 wire _03608_;
 wire _03609_;
 wire _03610_;
 wire _03611_;
 wire _03612_;
 wire _03613_;
 wire _03614_;
 wire _03615_;
 wire _03616_;
 wire _03617_;
 wire _03618_;
 wire _03619_;
 wire _03620_;
 wire _03621_;
 wire _03622_;
 wire _03623_;
 wire _03624_;
 wire _03625_;
 wire _03626_;
 wire _03627_;
 wire _03628_;
 wire _03629_;
 wire _03630_;
 wire _03631_;
 wire _03632_;
 wire _03633_;
 wire _03634_;
 wire _03635_;
 wire _03636_;
 wire _03637_;
 wire _03638_;
 wire _03639_;
 wire _03640_;
 wire _03641_;
 wire _03642_;
 wire _03643_;
 wire _03644_;
 wire _03645_;
 wire _03646_;
 wire _03647_;
 wire _03648_;
 wire _03649_;
 wire _03650_;
 wire _03651_;
 wire _03652_;
 wire _03653_;
 wire _03654_;
 wire _03655_;
 wire _03656_;
 wire _03657_;
 wire _03658_;
 wire _03659_;
 wire _03660_;
 wire _03661_;
 wire _03662_;
 wire _03663_;
 wire _03664_;
 wire _03665_;
 wire _03666_;
 wire _03667_;
 wire _03668_;
 wire _03669_;
 wire _03670_;
 wire _03671_;
 wire _03672_;
 wire _03673_;
 wire _03674_;
 wire _03675_;
 wire _03676_;
 wire _03677_;
 wire _03678_;
 wire _03679_;
 wire _03680_;
 wire _03681_;
 wire _03682_;
 wire _03683_;
 wire _03684_;
 wire _03685_;
 wire _03686_;
 wire _03687_;
 wire _03688_;
 wire _03689_;
 wire _03690_;
 wire _03691_;
 wire _03692_;
 wire _03693_;
 wire _03694_;
 wire _03695_;
 wire _03696_;
 wire _03697_;
 wire _03698_;
 wire _03699_;
 wire _03700_;
 wire _03701_;
 wire _03702_;
 wire _03703_;
 wire _03704_;
 wire _03705_;
 wire _03706_;
 wire _03707_;
 wire _03708_;
 wire _03709_;
 wire _03710_;
 wire _03711_;
 wire _03712_;
 wire _03713_;
 wire _03714_;
 wire _03715_;
 wire _03716_;
 wire _03717_;
 wire _03718_;
 wire _03719_;
 wire _03720_;
 wire _03721_;
 wire _03722_;
 wire _03723_;
 wire _03724_;
 wire _03725_;
 wire _03726_;
 wire _03727_;
 wire _03728_;
 wire _03729_;
 wire _03730_;
 wire _03731_;
 wire _03732_;
 wire _03733_;
 wire _03734_;
 wire _03735_;
 wire _03736_;
 wire _03737_;
 wire _03738_;
 wire _03739_;
 wire _03740_;
 wire _03741_;
 wire _03742_;
 wire _03743_;
 wire _03744_;
 wire _03745_;
 wire _03746_;
 wire _03747_;
 wire _03748_;
 wire _03749_;
 wire _03750_;
 wire _03751_;
 wire _03752_;
 wire _03753_;
 wire _03754_;
 wire _03755_;
 wire _03756_;
 wire _03757_;
 wire _03758_;
 wire _03759_;
 wire _03760_;
 wire _03761_;
 wire _03762_;
 wire _03763_;
 wire _03764_;
 wire _03765_;
 wire _03766_;
 wire _03767_;
 wire _03768_;
 wire _03769_;
 wire _03770_;
 wire _03771_;
 wire _03772_;
 wire _03773_;
 wire _03774_;
 wire _03775_;
 wire _03776_;
 wire _03777_;
 wire _03778_;
 wire _03779_;
 wire _03780_;
 wire _03781_;
 wire _03782_;
 wire _03783_;
 wire _03784_;
 wire _03785_;
 wire _03786_;
 wire _03787_;
 wire _03788_;
 wire _03789_;
 wire _03790_;
 wire _03791_;
 wire _03792_;
 wire _03793_;
 wire _03794_;
 wire _03795_;
 wire _03796_;
 wire _03797_;
 wire _03798_;
 wire _03799_;
 wire _03800_;
 wire _03801_;
 wire _03802_;
 wire _03803_;
 wire _03804_;
 wire _03805_;
 wire _03806_;
 wire _03807_;
 wire _03808_;
 wire _03809_;
 wire _03810_;
 wire _03811_;
 wire _03812_;
 wire _03813_;
 wire _03814_;
 wire _03815_;
 wire _03816_;
 wire _03817_;
 wire _03818_;
 wire _03819_;
 wire _03820_;
 wire _03821_;
 wire _03822_;
 wire _03823_;
 wire _03824_;
 wire _03825_;
 wire _03826_;
 wire _03827_;
 wire _03828_;
 wire _03829_;
 wire _03830_;
 wire _03831_;
 wire _03832_;
 wire _03833_;
 wire _03834_;
 wire _03835_;
 wire _03836_;
 wire _03837_;
 wire _03838_;
 wire _03839_;
 wire _03840_;
 wire _03841_;
 wire _03842_;
 wire _03843_;
 wire _03844_;
 wire _03845_;
 wire _03846_;
 wire _03847_;
 wire _03848_;
 wire _03849_;
 wire _03850_;
 wire _03851_;
 wire _03852_;
 wire _03853_;
 wire _03854_;
 wire _03855_;
 wire _03856_;
 wire _03857_;
 wire _03858_;
 wire _03859_;
 wire _03860_;
 wire _03861_;
 wire _03862_;
 wire _03863_;
 wire _03864_;
 wire _03865_;
 wire _03866_;
 wire _03867_;
 wire _03868_;
 wire _03869_;
 wire _03870_;
 wire _03871_;
 wire _03872_;
 wire _03873_;
 wire _03874_;
 wire _03875_;
 wire _03876_;
 wire _03877_;
 wire _03878_;
 wire _03879_;
 wire _03880_;
 wire _03881_;
 wire _03882_;
 wire _03883_;
 wire _03884_;
 wire _03885_;
 wire _03886_;
 wire _03887_;
 wire _03888_;
 wire _03889_;
 wire _03890_;
 wire _03891_;
 wire _03892_;
 wire _03893_;
 wire _03894_;
 wire _03895_;
 wire _03896_;
 wire _03897_;
 wire _03898_;
 wire _03899_;
 wire _03900_;
 wire _03901_;
 wire _03902_;
 wire _03903_;
 wire _03904_;
 wire _03905_;
 wire _03906_;
 wire _03907_;
 wire _03908_;
 wire _03909_;
 wire _03910_;
 wire _03911_;
 wire _03912_;
 wire _03913_;
 wire _03914_;
 wire _03915_;
 wire _03916_;
 wire _03917_;
 wire _03918_;
 wire _03919_;
 wire _03920_;
 wire _03921_;
 wire _03922_;
 wire _03923_;
 wire _03924_;
 wire _03925_;
 wire _03926_;
 wire _03927_;
 wire _03928_;
 wire _03929_;
 wire _03930_;
 wire _03931_;
 wire _03932_;
 wire _03933_;
 wire _03934_;
 wire _03935_;
 wire _03936_;
 wire _03937_;
 wire _03938_;
 wire _03939_;
 wire _03940_;
 wire _03941_;
 wire _03942_;
 wire _03943_;
 wire _03944_;
 wire _03945_;
 wire _03946_;
 wire _03947_;
 wire _03948_;
 wire _03949_;
 wire _03950_;
 wire _03951_;
 wire _03952_;
 wire _03953_;
 wire _03954_;
 wire _03955_;
 wire _03956_;
 wire _03957_;
 wire _03958_;
 wire _03959_;
 wire _03960_;
 wire _03961_;
 wire _03962_;
 wire _03963_;
 wire _03964_;
 wire _03965_;
 wire _03966_;
 wire _03967_;
 wire _03968_;
 wire _03969_;
 wire _03970_;
 wire _03971_;
 wire _03972_;
 wire _03973_;
 wire _03974_;
 wire _03975_;
 wire _03976_;
 wire _03977_;
 wire _03978_;
 wire _03979_;
 wire _03980_;
 wire _03981_;
 wire _03982_;
 wire _03983_;
 wire _03984_;
 wire _03985_;
 wire _03986_;
 wire _03987_;
 wire _03988_;
 wire _03989_;
 wire _03990_;
 wire _03991_;
 wire _03992_;
 wire _03993_;
 wire _03994_;
 wire _03995_;
 wire _03996_;
 wire _03997_;
 wire _03998_;
 wire _03999_;
 wire _04000_;
 wire _04001_;
 wire _04002_;
 wire _04003_;
 wire _04004_;
 wire _04005_;
 wire _04006_;
 wire _04007_;
 wire _04008_;
 wire _04009_;
 wire _04010_;
 wire _04011_;
 wire _04012_;
 wire _04013_;
 wire _04014_;
 wire _04015_;
 wire _04016_;
 wire _04017_;
 wire _04018_;
 wire _04019_;
 wire _04020_;
 wire _04021_;
 wire _04022_;
 wire _04023_;
 wire _04024_;
 wire _04025_;
 wire _04026_;
 wire _04027_;
 wire _04028_;
 wire _04029_;
 wire _04030_;
 wire _04031_;
 wire _04032_;
 wire _04033_;
 wire _04034_;
 wire _04035_;
 wire _04036_;
 wire _04037_;
 wire _04038_;
 wire _04039_;
 wire _04040_;
 wire _04041_;
 wire _04042_;
 wire _04043_;
 wire _04044_;
 wire _04045_;
 wire _04046_;
 wire _04047_;
 wire _04048_;
 wire _04049_;
 wire _04050_;
 wire _04051_;
 wire _04052_;
 wire _04053_;
 wire _04054_;
 wire _04055_;
 wire _04056_;
 wire _04057_;
 wire _04058_;
 wire _04059_;
 wire _04060_;
 wire _04061_;
 wire _04062_;
 wire _04063_;
 wire _04064_;
 wire _04065_;
 wire _04066_;
 wire _04067_;
 wire _04068_;
 wire _04069_;
 wire _04070_;
 wire _04071_;
 wire _04072_;
 wire _04073_;
 wire _04074_;
 wire _04075_;
 wire _04076_;
 wire _04077_;
 wire _04078_;
 wire _04079_;
 wire _04080_;
 wire _04081_;
 wire _04082_;
 wire _04083_;
 wire _04084_;
 wire _04085_;
 wire _04086_;
 wire _04087_;
 wire _04088_;
 wire _04089_;
 wire _04090_;
 wire _04091_;
 wire _04092_;
 wire _04093_;
 wire _04094_;
 wire _04095_;
 wire _04096_;
 wire _04097_;
 wire _04098_;
 wire _04099_;
 wire _04100_;
 wire _04101_;
 wire _04102_;
 wire _04103_;
 wire _04104_;
 wire _04105_;
 wire _04106_;
 wire _04107_;
 wire _04108_;
 wire _04109_;
 wire _04110_;
 wire _04111_;
 wire _04112_;
 wire _04113_;
 wire _04114_;
 wire _04115_;
 wire _04116_;
 wire _04117_;
 wire _04118_;
 wire _04119_;
 wire _04120_;
 wire _04121_;
 wire _04122_;
 wire _04123_;
 wire _04124_;
 wire _04125_;
 wire _04126_;
 wire _04127_;
 wire _04128_;
 wire _04129_;
 wire _04130_;
 wire _04131_;
 wire _04132_;
 wire _04133_;
 wire _04134_;
 wire _04135_;
 wire _04136_;
 wire _04137_;
 wire _04138_;
 wire _04139_;
 wire _04140_;
 wire _04141_;
 wire _04142_;
 wire _04143_;
 wire _04144_;
 wire _04145_;
 wire _04146_;
 wire _04147_;
 wire _04148_;
 wire _04149_;
 wire _04150_;
 wire _04151_;
 wire _04152_;
 wire _04153_;
 wire _04154_;
 wire _04155_;
 wire _04156_;
 wire _04157_;
 wire _04158_;
 wire _04159_;
 wire _04160_;
 wire _04161_;
 wire _04162_;
 wire _04163_;
 wire _04164_;
 wire _04165_;
 wire _04166_;
 wire _04167_;
 wire _04168_;
 wire _04169_;
 wire _04170_;
 wire _04171_;
 wire _04172_;
 wire _04173_;
 wire _04174_;
 wire _04175_;
 wire _04176_;
 wire _04177_;
 wire _04178_;
 wire _04179_;
 wire _04180_;
 wire _04181_;
 wire _04182_;
 wire _04183_;
 wire _04184_;
 wire _04185_;
 wire _04186_;
 wire _04187_;
 wire _04188_;
 wire _04189_;
 wire _04190_;
 wire _04191_;
 wire _04192_;
 wire _04193_;
 wire _04194_;
 wire _04195_;
 wire _04196_;
 wire _04197_;
 wire _04198_;
 wire _04199_;
 wire _04200_;
 wire _04201_;
 wire _04202_;
 wire _04203_;
 wire _04204_;
 wire _04205_;
 wire _04206_;
 wire _04207_;
 wire _04208_;
 wire _04209_;
 wire _04210_;
 wire _04211_;
 wire _04212_;
 wire _04213_;
 wire _04214_;
 wire _04215_;
 wire _04216_;
 wire _04217_;
 wire _04218_;
 wire _04219_;
 wire _04220_;
 wire _04221_;
 wire _04222_;
 wire _04223_;
 wire _04224_;
 wire _04225_;
 wire _04226_;
 wire _04227_;
 wire _04228_;
 wire _04229_;
 wire _04230_;
 wire _04231_;
 wire _04232_;
 wire _04233_;
 wire _04234_;
 wire _04235_;
 wire _04236_;
 wire _04237_;
 wire _04238_;
 wire _04239_;
 wire _04240_;
 wire _04241_;
 wire _04242_;
 wire _04243_;
 wire _04244_;
 wire _04245_;
 wire _04246_;
 wire _04247_;
 wire _04248_;
 wire _04249_;
 wire _04250_;
 wire _04251_;
 wire _04252_;
 wire _04253_;
 wire _04254_;
 wire _04255_;
 wire _04256_;
 wire _04257_;
 wire _04258_;
 wire _04259_;
 wire _04260_;
 wire _04261_;
 wire _04262_;
 wire _04263_;
 wire _04264_;
 wire _04265_;
 wire _04266_;
 wire _04267_;
 wire _04268_;
 wire _04269_;
 wire _04270_;
 wire _04271_;
 wire _04272_;
 wire _04273_;
 wire _04274_;
 wire _04275_;
 wire _04276_;
 wire _04277_;
 wire _04278_;
 wire _04279_;
 wire _04280_;
 wire _04281_;
 wire _04282_;
 wire _04283_;
 wire _04284_;
 wire _04285_;
 wire _04286_;
 wire _04287_;
 wire _04288_;
 wire _04289_;
 wire _04290_;
 wire _04291_;
 wire _04292_;
 wire _04293_;
 wire _04294_;
 wire _04295_;
 wire _04296_;
 wire _04297_;
 wire _04298_;
 wire _04299_;
 wire _04300_;
 wire _04301_;
 wire _04302_;
 wire _04303_;
 wire _04304_;
 wire _04305_;
 wire _04306_;
 wire _04307_;
 wire _04308_;
 wire _04309_;
 wire _04310_;
 wire _04311_;
 wire _04312_;
 wire _04313_;
 wire _04314_;
 wire _04315_;
 wire _04316_;
 wire _04317_;
 wire _04318_;
 wire _04319_;
 wire _04320_;
 wire _04321_;
 wire _04322_;
 wire _04323_;
 wire _04324_;
 wire _04325_;
 wire _04326_;
 wire _04327_;
 wire _04328_;
 wire _04329_;
 wire _04330_;
 wire _04331_;
 wire _04332_;
 wire _04333_;
 wire _04334_;
 wire _04335_;
 wire _04336_;
 wire _04337_;
 wire _04338_;
 wire _04339_;
 wire _04340_;
 wire _04341_;
 wire _04342_;
 wire _04343_;
 wire _04344_;
 wire _04345_;
 wire _04346_;
 wire _04347_;
 wire _04348_;
 wire _04349_;
 wire _04350_;
 wire _04351_;
 wire _04352_;
 wire _04353_;
 wire _04354_;
 wire _04355_;
 wire _04356_;
 wire _04357_;
 wire _04358_;
 wire _04359_;
 wire _04360_;
 wire _04361_;
 wire _04362_;
 wire _04363_;
 wire _04364_;
 wire _04365_;
 wire _04366_;
 wire _04367_;
 wire _04368_;
 wire _04369_;
 wire _04370_;
 wire _04371_;
 wire _04372_;
 wire _04373_;
 wire _04374_;
 wire _04375_;
 wire _04376_;
 wire _04377_;
 wire _04378_;
 wire _04379_;
 wire _04380_;
 wire _04381_;
 wire _04382_;
 wire _04383_;
 wire _04384_;
 wire _04385_;
 wire _04386_;
 wire _04387_;
 wire _04388_;
 wire _04389_;
 wire _04390_;
 wire _04391_;
 wire _04392_;
 wire _04393_;
 wire _04394_;
 wire _04395_;
 wire _04396_;
 wire _04397_;
 wire _04398_;
 wire _04399_;
 wire _04400_;
 wire _04401_;
 wire _04402_;
 wire _04403_;
 wire _04404_;
 wire _04405_;
 wire _04406_;
 wire _04407_;
 wire _04408_;
 wire _04409_;
 wire _04410_;
 wire _04411_;
 wire _04412_;
 wire _04413_;
 wire _04414_;
 wire _04415_;
 wire _04416_;
 wire _04417_;
 wire _04418_;
 wire _04419_;
 wire _04420_;
 wire _04421_;
 wire _04422_;
 wire _04423_;
 wire _04424_;
 wire _04425_;
 wire _04426_;
 wire _04427_;
 wire _04428_;
 wire _04429_;
 wire _04430_;
 wire _04431_;
 wire _04432_;
 wire _04433_;
 wire _04434_;
 wire _04435_;
 wire _04436_;
 wire _04437_;
 wire _04438_;
 wire _04439_;
 wire _04440_;
 wire _04441_;
 wire _04442_;
 wire _04443_;
 wire _04444_;
 wire _04445_;
 wire _04446_;
 wire _04447_;
 wire _04448_;
 wire _04449_;
 wire _04450_;
 wire _04451_;
 wire _04452_;
 wire _04453_;
 wire _04454_;
 wire _04455_;
 wire _04456_;
 wire _04457_;
 wire _04458_;
 wire _04459_;
 wire _04460_;
 wire _04461_;
 wire _04462_;
 wire _04463_;
 wire _04464_;
 wire _04465_;
 wire _04466_;
 wire _04467_;
 wire _04468_;
 wire _04469_;
 wire _04470_;
 wire _04471_;
 wire _04472_;
 wire _04473_;
 wire _04474_;
 wire _04475_;
 wire _04476_;
 wire _04477_;
 wire _04478_;
 wire _04479_;
 wire _04480_;
 wire _04481_;
 wire _04482_;
 wire _04483_;
 wire _04484_;
 wire _04485_;
 wire _04486_;
 wire _04487_;
 wire _04488_;
 wire _04489_;
 wire _04490_;
 wire _04491_;
 wire _04492_;
 wire _04493_;
 wire _04494_;
 wire _04495_;
 wire _04496_;
 wire _04497_;
 wire _04498_;
 wire _04499_;
 wire _04500_;
 wire _04501_;
 wire _04502_;
 wire _04503_;
 wire _04504_;
 wire _04505_;
 wire _04506_;
 wire _04507_;
 wire _04508_;
 wire _04509_;
 wire _04510_;
 wire _04511_;
 wire _04512_;
 wire _04513_;
 wire _04514_;
 wire _04515_;
 wire _04516_;
 wire _04517_;
 wire _04518_;
 wire _04519_;
 wire _04520_;
 wire _04521_;
 wire _04522_;
 wire _04523_;
 wire _04524_;
 wire _04525_;
 wire _04526_;
 wire _04527_;
 wire _04528_;
 wire _04529_;
 wire _04530_;
 wire _04531_;
 wire _04532_;
 wire _04533_;
 wire _04534_;
 wire _04535_;
 wire _04536_;
 wire _04537_;
 wire _04538_;
 wire _04539_;
 wire _04540_;
 wire _04541_;
 wire _04542_;
 wire _04543_;
 wire _04544_;
 wire _04545_;
 wire _04546_;
 wire _04547_;
 wire _04548_;
 wire _04549_;
 wire _04550_;
 wire _04551_;
 wire _04552_;
 wire _04553_;
 wire _04554_;
 wire _04555_;
 wire _04556_;
 wire _04557_;
 wire _04558_;
 wire _04559_;
 wire _04560_;
 wire _04561_;
 wire _04562_;
 wire _04563_;
 wire _04564_;
 wire _04565_;
 wire _04566_;
 wire _04567_;
 wire _04568_;
 wire _04569_;
 wire _04570_;
 wire _04571_;
 wire _04572_;
 wire _04573_;
 wire _04574_;
 wire _04575_;
 wire _04576_;
 wire _04577_;
 wire _04578_;
 wire _04579_;
 wire _04580_;
 wire _04581_;
 wire _04582_;
 wire _04583_;
 wire _04584_;
 wire _04585_;
 wire _04586_;
 wire _04587_;
 wire _04588_;
 wire _04589_;
 wire _04590_;
 wire _04591_;
 wire _04592_;
 wire _04593_;
 wire _04594_;
 wire _04595_;
 wire _04596_;
 wire _04597_;
 wire _04598_;
 wire _04599_;
 wire _04600_;
 wire _04601_;
 wire _04602_;
 wire _04603_;
 wire _04604_;
 wire _04605_;
 wire _04606_;
 wire _04607_;
 wire _04608_;
 wire _04609_;
 wire _04610_;
 wire _04611_;
 wire _04612_;
 wire _04613_;
 wire _04614_;
 wire _04615_;
 wire _04616_;
 wire _04617_;
 wire _04618_;
 wire _04619_;
 wire _04620_;
 wire _04621_;
 wire _04622_;
 wire _04623_;
 wire _04624_;
 wire _04625_;
 wire _04626_;
 wire _04627_;
 wire _04628_;
 wire _04629_;
 wire _04630_;
 wire _04631_;
 wire _04632_;
 wire _04633_;
 wire _04634_;
 wire _04635_;
 wire _04636_;
 wire _04637_;
 wire _04638_;
 wire _04639_;
 wire _04640_;
 wire _04641_;
 wire _04642_;
 wire _04643_;
 wire _04644_;
 wire _04645_;
 wire _04646_;
 wire _04647_;
 wire _04648_;
 wire _04649_;
 wire _04650_;
 wire _04651_;
 wire _04652_;
 wire _04653_;
 wire _04654_;
 wire _04655_;
 wire _04656_;
 wire _04657_;
 wire _04658_;
 wire _04659_;
 wire _04660_;
 wire _04661_;
 wire _04662_;
 wire _04663_;
 wire _04664_;
 wire _04665_;
 wire _04666_;
 wire _04667_;
 wire _04668_;
 wire _04669_;
 wire _04670_;
 wire _04671_;
 wire _04672_;
 wire _04673_;
 wire _04674_;
 wire _04675_;
 wire _04676_;
 wire _04677_;
 wire _04678_;
 wire _04679_;
 wire _04680_;
 wire _04681_;
 wire _04682_;
 wire _04683_;
 wire _04684_;
 wire _04685_;
 wire _04686_;
 wire _04687_;
 wire _04688_;
 wire _04689_;
 wire _04690_;
 wire _04691_;
 wire _04692_;
 wire _04693_;
 wire _04694_;
 wire _04695_;
 wire _04696_;
 wire _04697_;
 wire _04698_;
 wire _04699_;
 wire _04700_;
 wire _04701_;
 wire _04702_;
 wire _04703_;
 wire _04704_;
 wire _04705_;
 wire _04706_;
 wire _04707_;
 wire _04708_;
 wire _04709_;
 wire _04710_;
 wire _04711_;
 wire _04712_;
 wire _04713_;
 wire _04714_;
 wire _04715_;
 wire _04716_;
 wire _04717_;
 wire _04718_;
 wire _04719_;
 wire _04720_;
 wire _04721_;
 wire _04722_;
 wire _04723_;
 wire _04724_;
 wire _04725_;
 wire _04726_;
 wire _04727_;
 wire _04728_;
 wire _04729_;
 wire _04730_;
 wire _04731_;
 wire _04732_;
 wire _04733_;
 wire _04734_;
 wire _04735_;
 wire _04736_;
 wire _04737_;
 wire _04738_;
 wire _04739_;
 wire _04740_;
 wire _04741_;
 wire _04742_;
 wire _04743_;
 wire _04744_;
 wire _04745_;
 wire _04746_;
 wire _04747_;
 wire _04748_;
 wire _04749_;
 wire _04750_;
 wire _04751_;
 wire _04752_;
 wire _04753_;
 wire _04754_;
 wire _04755_;
 wire _04756_;
 wire _04757_;
 wire _04758_;
 wire _04759_;
 wire _04760_;
 wire _04761_;
 wire _04762_;
 wire _04763_;
 wire _04764_;
 wire _04765_;
 wire _04766_;
 wire _04767_;
 wire _04768_;
 wire _04769_;
 wire _04770_;
 wire _04771_;
 wire _04772_;
 wire _04773_;
 wire _04774_;
 wire _04775_;
 wire _04776_;
 wire _04777_;
 wire _04778_;
 wire _04779_;
 wire _04780_;
 wire _04781_;
 wire _04782_;
 wire _04783_;
 wire _04784_;
 wire _04785_;
 wire _04786_;
 wire _04787_;
 wire _04788_;
 wire _04789_;
 wire _04790_;
 wire _04791_;
 wire _04792_;
 wire _04793_;
 wire _04794_;
 wire _04795_;
 wire _04796_;
 wire _04797_;
 wire _04798_;
 wire _04799_;
 wire _04800_;
 wire _04801_;
 wire _04802_;
 wire _04803_;
 wire _04804_;
 wire _04805_;
 wire _04806_;
 wire _04807_;
 wire _04808_;
 wire _04809_;
 wire _04810_;
 wire _04811_;
 wire _04812_;
 wire _04813_;
 wire _04814_;
 wire _04815_;
 wire _04816_;
 wire _04817_;
 wire _04818_;
 wire _04819_;
 wire _04820_;
 wire _04821_;
 wire _04822_;
 wire _04823_;
 wire _04824_;
 wire _04825_;
 wire _04826_;
 wire _04827_;
 wire _04828_;
 wire _04829_;
 wire _04830_;
 wire _04831_;
 wire _04832_;
 wire _04833_;
 wire _04834_;
 wire _04835_;
 wire _04836_;
 wire _04837_;
 wire _04838_;
 wire _04839_;
 wire _04840_;
 wire _04841_;
 wire _04842_;
 wire _04843_;
 wire _04844_;
 wire _04845_;
 wire _04846_;
 wire _04847_;
 wire _04848_;
 wire _04849_;
 wire _04850_;
 wire _04851_;
 wire _04852_;
 wire _04853_;
 wire _04854_;
 wire _04855_;
 wire _04856_;
 wire _04857_;
 wire _04858_;
 wire _04859_;
 wire _04860_;
 wire _04861_;
 wire _04862_;
 wire _04863_;
 wire _04864_;
 wire _04865_;
 wire _04866_;
 wire _04867_;
 wire _04868_;
 wire _04869_;
 wire _04870_;
 wire _04871_;
 wire _04872_;
 wire _04873_;
 wire _04874_;
 wire _04875_;
 wire _04876_;
 wire _04877_;
 wire _04878_;
 wire _04879_;
 wire _04880_;
 wire _04881_;
 wire _04882_;
 wire _04883_;
 wire _04884_;
 wire _04885_;
 wire _04886_;
 wire _04887_;
 wire _04888_;
 wire _04889_;
 wire _04890_;
 wire _04891_;
 wire _04892_;
 wire _04893_;
 wire _04894_;
 wire _04895_;
 wire _04896_;
 wire _04897_;
 wire _04898_;
 wire _04899_;
 wire _04900_;
 wire _04901_;
 wire _04902_;
 wire _04903_;
 wire _04904_;
 wire _04905_;
 wire _04906_;
 wire _04907_;
 wire _04908_;
 wire _04909_;
 wire _04910_;
 wire _04911_;
 wire _04912_;
 wire _04913_;
 wire _04914_;
 wire _04915_;
 wire _04916_;
 wire _04917_;
 wire _04918_;
 wire _04919_;
 wire _04920_;
 wire _04921_;
 wire _04922_;
 wire _04923_;
 wire _04924_;
 wire _04925_;
 wire _04926_;
 wire _04927_;
 wire _04928_;
 wire _04929_;
 wire _04930_;
 wire _04931_;
 wire _04932_;
 wire _04933_;
 wire _04934_;
 wire _04935_;
 wire _04936_;
 wire _04937_;
 wire _04938_;
 wire _04939_;
 wire _04940_;
 wire _04941_;
 wire _04942_;
 wire _04943_;
 wire _04944_;
 wire _04945_;
 wire _04946_;
 wire _04947_;
 wire _04948_;
 wire _04949_;
 wire _04950_;
 wire _04951_;
 wire _04952_;
 wire _04953_;
 wire _04954_;
 wire _04955_;
 wire _04956_;
 wire _04957_;
 wire _04958_;
 wire _04959_;
 wire _04960_;
 wire _04961_;
 wire _04962_;
 wire _04963_;
 wire _04964_;
 wire _04965_;
 wire _04966_;
 wire _04967_;
 wire _04968_;
 wire _04969_;
 wire _04970_;
 wire _04971_;
 wire _04972_;
 wire _04973_;
 wire _04974_;
 wire _04975_;
 wire _04976_;
 wire _04977_;
 wire _04978_;
 wire _04979_;
 wire _04980_;
 wire _04981_;
 wire _04982_;
 wire _04983_;
 wire _04984_;
 wire _04985_;
 wire _04986_;
 wire _04987_;
 wire _04988_;
 wire _04989_;
 wire _04990_;
 wire _04991_;
 wire _04992_;
 wire _04993_;
 wire _04994_;
 wire _04995_;
 wire _04996_;
 wire _04997_;
 wire _04998_;
 wire _04999_;
 wire _05000_;
 wire _05001_;
 wire _05002_;
 wire _05003_;
 wire _05004_;
 wire _05005_;
 wire _05006_;
 wire _05007_;
 wire _05008_;
 wire _05009_;
 wire _05010_;
 wire _05011_;
 wire _05012_;
 wire _05013_;
 wire _05014_;
 wire _05015_;
 wire _05016_;
 wire _05017_;
 wire _05018_;
 wire _05019_;
 wire _05020_;
 wire _05021_;
 wire _05022_;
 wire _05023_;
 wire _05024_;
 wire _05025_;
 wire _05026_;
 wire _05027_;
 wire _05028_;
 wire _05029_;
 wire _05030_;
 wire _05031_;
 wire _05032_;
 wire _05033_;
 wire _05034_;
 wire _05035_;
 wire _05036_;
 wire _05037_;
 wire _05038_;
 wire _05039_;
 wire _05040_;
 wire _05041_;
 wire _05042_;
 wire _05043_;
 wire _05044_;
 wire _05045_;
 wire _05046_;
 wire _05047_;
 wire _05048_;
 wire _05049_;
 wire _05050_;
 wire _05051_;
 wire _05052_;
 wire _05053_;
 wire _05054_;
 wire _05055_;
 wire _05056_;
 wire _05057_;
 wire _05058_;
 wire _05059_;
 wire _05060_;
 wire _05061_;
 wire _05062_;
 wire _05063_;
 wire _05064_;
 wire _05065_;
 wire _05066_;
 wire _05067_;
 wire _05068_;
 wire _05069_;
 wire _05070_;
 wire _05071_;
 wire _05072_;
 wire _05073_;
 wire _05074_;
 wire _05075_;
 wire _05076_;
 wire _05077_;
 wire _05078_;
 wire _05079_;
 wire _05080_;
 wire _05081_;
 wire _05082_;
 wire _05083_;
 wire _05084_;
 wire _05085_;
 wire _05086_;
 wire _05087_;
 wire _05088_;
 wire _05089_;
 wire _05090_;
 wire _05091_;
 wire _05092_;
 wire _05093_;
 wire _05094_;
 wire _05095_;
 wire _05096_;
 wire _05097_;
 wire _05098_;
 wire _05099_;
 wire _05100_;
 wire _05101_;
 wire _05102_;
 wire _05103_;
 wire _05104_;
 wire _05105_;
 wire _05106_;
 wire _05107_;
 wire _05108_;
 wire _05109_;
 wire _05110_;
 wire _05111_;
 wire _05112_;
 wire _05113_;
 wire _05114_;
 wire _05115_;
 wire _05116_;
 wire _05117_;
 wire _05118_;
 wire _05119_;
 wire _05120_;
 wire _05121_;
 wire _05122_;
 wire _05123_;
 wire _05124_;
 wire _05125_;
 wire _05126_;
 wire _05127_;
 wire _05128_;
 wire _05129_;
 wire _05130_;
 wire _05131_;
 wire _05132_;
 wire _05133_;
 wire _05134_;
 wire _05135_;
 wire _05136_;
 wire _05137_;
 wire _05138_;
 wire _05139_;
 wire _05140_;
 wire _05141_;
 wire _05142_;
 wire _05143_;
 wire _05144_;
 wire _05145_;
 wire _05146_;
 wire _05147_;
 wire _05148_;
 wire _05149_;
 wire _05150_;
 wire _05151_;
 wire _05152_;
 wire _05153_;
 wire _05154_;
 wire _05155_;
 wire _05156_;
 wire _05157_;
 wire _05158_;
 wire _05159_;
 wire _05160_;
 wire _05161_;
 wire _05162_;
 wire _05163_;
 wire _05164_;
 wire _05165_;
 wire _05166_;
 wire _05167_;
 wire _05168_;
 wire _05169_;
 wire _05170_;
 wire _05171_;
 wire _05172_;
 wire _05173_;
 wire _05174_;
 wire _05175_;
 wire _05176_;
 wire _05177_;
 wire _05178_;
 wire _05179_;
 wire _05180_;
 wire _05181_;
 wire _05182_;
 wire _05183_;
 wire _05184_;
 wire _05185_;
 wire _05186_;
 wire _05187_;
 wire _05188_;
 wire _05189_;
 wire _05190_;
 wire _05191_;
 wire _05192_;
 wire _05193_;
 wire _05194_;
 wire _05195_;
 wire _05196_;
 wire _05197_;
 wire _05198_;
 wire _05199_;
 wire _05200_;
 wire _05201_;
 wire _05202_;
 wire _05203_;
 wire _05204_;
 wire _05205_;
 wire _05206_;
 wire _05207_;
 wire _05208_;
 wire _05209_;
 wire _05210_;
 wire _05211_;
 wire _05212_;
 wire _05213_;
 wire _05214_;
 wire _05215_;
 wire _05216_;
 wire _05217_;
 wire _05218_;
 wire _05219_;
 wire _05220_;
 wire _05221_;
 wire _05222_;
 wire _05223_;
 wire _05224_;
 wire _05225_;
 wire _05226_;
 wire _05227_;
 wire _05228_;
 wire _05229_;
 wire _05230_;
 wire _05231_;
 wire _05232_;
 wire _05233_;
 wire _05234_;
 wire _05235_;
 wire _05236_;
 wire _05237_;
 wire _05238_;
 wire _05239_;
 wire _05240_;
 wire _05241_;
 wire _05242_;
 wire _05243_;
 wire _05244_;
 wire _05245_;
 wire _05246_;
 wire _05247_;
 wire _05248_;
 wire _05249_;
 wire _05250_;
 wire _05251_;
 wire _05252_;
 wire _05253_;
 wire _05254_;
 wire _05255_;
 wire _05256_;
 wire _05257_;
 wire _05258_;
 wire _05259_;
 wire _05260_;
 wire _05261_;
 wire _05262_;
 wire _05263_;
 wire _05264_;
 wire _05265_;
 wire _05266_;
 wire _05267_;
 wire _05268_;
 wire _05269_;
 wire _05270_;
 wire _05271_;
 wire _05272_;
 wire _05273_;
 wire _05274_;
 wire _05275_;
 wire _05276_;
 wire _05277_;
 wire _05278_;
 wire _05279_;
 wire _05280_;
 wire _05281_;
 wire _05282_;
 wire _05283_;
 wire _05284_;
 wire _05285_;
 wire _05286_;
 wire _05287_;
 wire _05288_;
 wire _05289_;
 wire _05290_;
 wire _05291_;
 wire _05292_;
 wire _05293_;
 wire _05294_;
 wire _05295_;
 wire _05296_;
 wire _05297_;
 wire _05298_;
 wire _05299_;
 wire _05300_;
 wire _05301_;
 wire _05302_;
 wire _05303_;
 wire _05304_;
 wire _05305_;
 wire _05306_;
 wire _05307_;
 wire _05308_;
 wire _05309_;
 wire _05310_;
 wire _05311_;
 wire _05312_;
 wire _05313_;
 wire _05314_;
 wire _05315_;
 wire _05316_;
 wire _05317_;
 wire _05318_;
 wire _05319_;
 wire _05320_;
 wire _05321_;
 wire _05322_;
 wire _05323_;
 wire _05324_;
 wire _05325_;
 wire _05326_;
 wire _05327_;
 wire _05328_;
 wire _05329_;
 wire _05330_;
 wire _05331_;
 wire _05332_;
 wire _05333_;
 wire _05334_;
 wire _05335_;
 wire _05336_;
 wire _05337_;
 wire _05338_;
 wire _05339_;
 wire _05340_;
 wire _05341_;
 wire _05342_;
 wire _05343_;
 wire _05344_;
 wire _05345_;
 wire _05346_;
 wire _05347_;
 wire _05348_;
 wire _05349_;
 wire _05350_;
 wire _05351_;
 wire _05352_;
 wire _05353_;
 wire _05354_;
 wire _05355_;
 wire _05356_;
 wire _05357_;
 wire _05358_;
 wire _05359_;
 wire _05360_;
 wire _05361_;
 wire _05362_;
 wire _05363_;
 wire _05364_;
 wire _05365_;
 wire _05366_;
 wire _05367_;
 wire _05368_;
 wire _05369_;
 wire _05370_;
 wire _05371_;
 wire _05372_;
 wire _05373_;
 wire _05374_;
 wire _05375_;
 wire _05376_;
 wire _05377_;
 wire _05378_;
 wire _05379_;
 wire _05380_;
 wire _05381_;
 wire _05382_;
 wire _05383_;
 wire _05384_;
 wire _05385_;
 wire _05386_;
 wire _05387_;
 wire _05388_;
 wire _05389_;
 wire _05390_;
 wire _05391_;
 wire _05392_;
 wire _05393_;
 wire _05394_;
 wire _05395_;
 wire _05396_;
 wire _05397_;
 wire _05398_;
 wire _05399_;
 wire _05400_;
 wire _05401_;
 wire _05402_;
 wire _05403_;
 wire _05404_;
 wire _05405_;
 wire _05406_;
 wire _05407_;
 wire _05408_;
 wire _05409_;
 wire _05410_;
 wire _05411_;
 wire _05412_;
 wire _05413_;
 wire _05414_;
 wire _05415_;
 wire _05416_;
 wire _05417_;
 wire _05418_;
 wire _05419_;
 wire _05420_;
 wire _05421_;
 wire _05422_;
 wire _05423_;
 wire _05424_;
 wire _05425_;
 wire _05426_;
 wire _05427_;
 wire _05428_;
 wire _05429_;
 wire _05430_;
 wire _05431_;
 wire _05432_;
 wire _05433_;
 wire _05434_;
 wire _05435_;
 wire _05436_;
 wire _05437_;
 wire _05438_;
 wire _05439_;
 wire _05440_;
 wire _05441_;
 wire _05442_;
 wire _05443_;
 wire _05444_;
 wire _05445_;
 wire _05446_;
 wire _05447_;
 wire _05448_;
 wire _05449_;
 wire _05450_;
 wire _05451_;
 wire _05452_;
 wire _05453_;
 wire _05454_;
 wire _05455_;
 wire _05456_;
 wire _05457_;
 wire _05458_;
 wire _05459_;
 wire _05460_;
 wire _05461_;
 wire _05462_;
 wire _05463_;
 wire _05464_;
 wire _05465_;
 wire _05466_;
 wire _05467_;
 wire _05468_;
 wire _05469_;
 wire _05470_;
 wire _05471_;
 wire _05472_;
 wire _05473_;
 wire _05474_;
 wire _05475_;
 wire _05476_;
 wire _05477_;
 wire _05478_;
 wire _05479_;
 wire _05480_;
 wire _05481_;
 wire _05482_;
 wire _05483_;
 wire _05484_;
 wire _05485_;
 wire _05486_;
 wire _05487_;
 wire _05488_;
 wire _05489_;
 wire _05490_;
 wire _05491_;
 wire _05492_;
 wire _05493_;
 wire _05494_;
 wire _05495_;
 wire _05496_;
 wire _05497_;
 wire _05498_;
 wire _05499_;
 wire _05500_;
 wire _05501_;
 wire _05502_;
 wire _05503_;
 wire _05504_;
 wire _05505_;
 wire _05506_;
 wire _05507_;
 wire _05508_;
 wire _05509_;
 wire _05510_;
 wire _05511_;
 wire _05512_;
 wire _05513_;
 wire _05514_;
 wire _05515_;
 wire _05516_;
 wire _05517_;
 wire _05518_;
 wire _05519_;
 wire _05520_;
 wire _05521_;
 wire _05522_;
 wire _05523_;
 wire _05524_;
 wire _05525_;
 wire _05526_;
 wire _05527_;
 wire _05528_;
 wire _05529_;
 wire _05530_;
 wire _05531_;
 wire _05532_;
 wire _05533_;
 wire _05534_;
 wire _05535_;
 wire _05536_;
 wire _05537_;
 wire _05538_;
 wire _05539_;
 wire _05540_;
 wire _05541_;
 wire _05542_;
 wire _05543_;
 wire _05544_;
 wire _05545_;
 wire _05546_;
 wire _05547_;
 wire _05548_;
 wire _05549_;
 wire _05550_;
 wire _05551_;
 wire _05552_;
 wire _05553_;
 wire _05554_;
 wire _05555_;
 wire _05556_;
 wire _05557_;
 wire _05558_;
 wire _05559_;
 wire _05560_;
 wire _05561_;
 wire _05562_;
 wire _05563_;
 wire _05564_;
 wire _05565_;
 wire _05566_;
 wire _05567_;
 wire _05568_;
 wire _05569_;
 wire _05570_;
 wire _05571_;
 wire _05572_;
 wire _05573_;
 wire _05574_;
 wire _05575_;
 wire _05576_;
 wire _05577_;
 wire _05578_;
 wire _05579_;
 wire _05580_;
 wire _05581_;
 wire _05582_;
 wire _05583_;
 wire _05584_;
 wire _05585_;
 wire _05586_;
 wire _05587_;
 wire _05588_;
 wire _05589_;
 wire _05590_;
 wire _05591_;
 wire _05592_;
 wire _05593_;
 wire _05594_;
 wire _05595_;
 wire _05596_;
 wire _05597_;
 wire _05598_;
 wire _05599_;
 wire _05600_;
 wire _05601_;
 wire _05602_;
 wire _05603_;
 wire _05604_;
 wire _05605_;
 wire _05606_;
 wire _05607_;
 wire _05608_;
 wire _05609_;
 wire _05610_;
 wire _05611_;
 wire _05612_;
 wire _05613_;
 wire _05614_;
 wire _05615_;
 wire _05616_;
 wire _05617_;
 wire _05618_;
 wire _05619_;
 wire _05620_;
 wire _05621_;
 wire _05622_;
 wire _05623_;
 wire _05624_;
 wire _05625_;
 wire _05626_;
 wire _05627_;
 wire _05628_;
 wire _05629_;
 wire _05630_;
 wire _05631_;
 wire _05632_;
 wire _05633_;
 wire _05634_;
 wire _05635_;
 wire _05636_;
 wire _05637_;
 wire _05638_;
 wire _05639_;
 wire _05640_;
 wire _05641_;
 wire _05642_;
 wire _05643_;
 wire _05644_;
 wire _05645_;
 wire _05646_;
 wire _05647_;
 wire _05648_;
 wire _05649_;
 wire _05650_;
 wire _05651_;
 wire _05652_;
 wire _05653_;
 wire _05654_;
 wire _05655_;
 wire _05656_;
 wire _05657_;
 wire _05658_;
 wire _05659_;
 wire _05660_;
 wire _05661_;
 wire _05662_;
 wire _05663_;
 wire _05664_;
 wire _05665_;
 wire _05666_;
 wire _05667_;
 wire _05668_;
 wire _05669_;
 wire _05670_;
 wire _05671_;
 wire _05672_;
 wire _05673_;
 wire _05674_;
 wire _05675_;
 wire _05676_;
 wire _05677_;
 wire _05678_;
 wire _05679_;
 wire _05680_;
 wire _05681_;
 wire _05682_;
 wire _05683_;
 wire _05684_;
 wire _05685_;
 wire _05686_;
 wire _05687_;
 wire _05688_;
 wire _05689_;
 wire _05690_;
 wire _05691_;
 wire _05692_;
 wire _05693_;
 wire _05694_;
 wire _05695_;
 wire _05696_;
 wire _05697_;
 wire _05698_;
 wire _05699_;
 wire _05700_;
 wire _05701_;
 wire _05702_;
 wire _05703_;
 wire _05704_;
 wire _05705_;
 wire _05706_;
 wire _05707_;
 wire _05708_;
 wire _05709_;
 wire _05710_;
 wire _05711_;
 wire _05712_;
 wire _05713_;
 wire _05714_;
 wire _05715_;
 wire _05716_;
 wire _05717_;
 wire _05718_;
 wire _05719_;
 wire _05720_;
 wire _05721_;
 wire _05722_;
 wire _05723_;
 wire _05724_;
 wire _05725_;
 wire _05726_;
 wire _05727_;
 wire _05728_;
 wire _05729_;
 wire _05730_;
 wire _05731_;
 wire _05732_;
 wire _05733_;
 wire _05734_;
 wire _05735_;
 wire _05736_;
 wire _05737_;
 wire _05738_;
 wire _05739_;
 wire _05740_;
 wire _05741_;
 wire _05742_;
 wire _05743_;
 wire _05744_;
 wire _05745_;
 wire _05746_;
 wire _05747_;
 wire _05748_;
 wire _05749_;
 wire _05750_;
 wire _05751_;
 wire _05752_;
 wire _05753_;
 wire _05754_;
 wire _05755_;
 wire _05756_;
 wire _05757_;
 wire _05758_;
 wire _05759_;
 wire _05760_;
 wire _05761_;
 wire _05762_;
 wire _05763_;
 wire _05764_;
 wire _05765_;
 wire _05766_;
 wire _05767_;
 wire _05768_;
 wire _05769_;
 wire _05770_;
 wire _05771_;
 wire _05772_;
 wire _05773_;
 wire _05774_;
 wire _05775_;
 wire _05776_;
 wire _05777_;
 wire _05778_;
 wire _05779_;
 wire _05780_;
 wire _05781_;
 wire _05782_;
 wire _05783_;
 wire _05784_;
 wire _05785_;
 wire _05786_;
 wire _05787_;
 wire _05788_;
 wire _05789_;
 wire _05790_;
 wire _05791_;
 wire _05792_;
 wire _05793_;
 wire _05794_;
 wire _05795_;
 wire _05796_;
 wire _05797_;
 wire _05798_;
 wire _05799_;
 wire _05800_;
 wire _05801_;
 wire _05802_;
 wire _05803_;
 wire _05804_;
 wire _05805_;
 wire _05806_;
 wire _05807_;
 wire _05808_;
 wire _05809_;
 wire _05810_;
 wire _05811_;
 wire _05812_;
 wire _05813_;
 wire _05814_;
 wire _05815_;
 wire _05816_;
 wire _05817_;
 wire _05818_;
 wire _05819_;
 wire _05820_;
 wire _05821_;
 wire _05822_;
 wire _05823_;
 wire _05824_;
 wire _05825_;
 wire _05826_;
 wire _05827_;
 wire _05828_;
 wire _05829_;
 wire _05830_;
 wire _05831_;
 wire _05832_;
 wire _05833_;
 wire _05834_;
 wire _05835_;
 wire _05836_;
 wire _05837_;
 wire _05838_;
 wire _05839_;
 wire _05840_;
 wire _05841_;
 wire _05842_;
 wire _05843_;
 wire _05844_;
 wire _05845_;
 wire _05846_;
 wire _05847_;
 wire _05848_;
 wire _05849_;
 wire _05850_;
 wire _05851_;
 wire _05852_;
 wire _05853_;
 wire _05854_;
 wire _05855_;
 wire _05856_;
 wire _05857_;
 wire _05858_;
 wire _05859_;
 wire _05860_;
 wire _05861_;
 wire _05862_;
 wire _05863_;
 wire _05864_;
 wire _05865_;
 wire _05866_;
 wire _05867_;
 wire _05868_;
 wire _05869_;
 wire _05870_;
 wire _05871_;
 wire _05872_;
 wire _05873_;
 wire _05874_;
 wire _05875_;
 wire _05876_;
 wire _05877_;
 wire _05878_;
 wire _05879_;
 wire _05880_;
 wire _05881_;
 wire _05882_;
 wire _05883_;
 wire _05884_;
 wire _05885_;
 wire _05886_;
 wire _05887_;
 wire _05888_;
 wire _05889_;
 wire _05890_;
 wire _05891_;
 wire _05892_;
 wire _05893_;
 wire _05894_;
 wire _05895_;
 wire _05896_;
 wire _05897_;
 wire _05898_;
 wire _05899_;
 wire _05900_;
 wire _05901_;
 wire _05902_;
 wire _05903_;
 wire _05904_;
 wire _05905_;
 wire _05906_;
 wire _05907_;
 wire _05908_;
 wire _05909_;
 wire _05910_;
 wire _05911_;
 wire _05912_;
 wire _05913_;
 wire _05914_;
 wire _05915_;
 wire _05916_;
 wire _05917_;
 wire _05918_;
 wire _05919_;
 wire _05920_;
 wire _05921_;
 wire _05922_;
 wire _05923_;
 wire _05924_;
 wire _05925_;
 wire _05926_;
 wire _05927_;
 wire _05928_;
 wire _05929_;
 wire _05930_;
 wire _05931_;
 wire _05932_;
 wire _05933_;
 wire _05934_;
 wire _05935_;
 wire _05936_;
 wire _05937_;
 wire _05938_;
 wire _05939_;
 wire _05940_;
 wire _05941_;
 wire _05942_;
 wire _05943_;
 wire _05944_;
 wire _05945_;
 wire _05946_;
 wire _05947_;
 wire _05948_;
 wire _05949_;
 wire _05950_;
 wire _05951_;
 wire _05952_;
 wire _05953_;
 wire _05954_;
 wire _05955_;
 wire _05956_;
 wire _05957_;
 wire _05958_;
 wire _05959_;
 wire _05960_;
 wire _05961_;
 wire _05962_;
 wire _05963_;
 wire _05964_;
 wire _05965_;
 wire _05966_;
 wire _05967_;
 wire _05968_;
 wire _05969_;
 wire _05970_;
 wire _05971_;
 wire _05972_;
 wire _05973_;
 wire _05974_;
 wire _05975_;
 wire _05976_;
 wire _05977_;
 wire _05978_;
 wire _05979_;
 wire _05980_;
 wire _05981_;
 wire _05982_;
 wire _05983_;
 wire _05984_;
 wire _05985_;
 wire _05986_;
 wire _05987_;
 wire _05988_;
 wire _05989_;
 wire _05990_;
 wire _05991_;
 wire _05992_;
 wire _05993_;
 wire _05994_;
 wire _05995_;
 wire _05996_;
 wire _05997_;
 wire _05998_;
 wire _05999_;
 wire _06000_;
 wire _06001_;
 wire _06002_;
 wire _06003_;
 wire _06004_;
 wire _06005_;
 wire _06006_;
 wire _06007_;
 wire _06008_;
 wire _06009_;
 wire _06010_;
 wire _06011_;
 wire _06012_;
 wire _06013_;
 wire _06014_;
 wire _06015_;
 wire _06016_;
 wire _06017_;
 wire _06018_;
 wire _06019_;
 wire _06020_;
 wire _06021_;
 wire _06022_;
 wire _06023_;
 wire _06024_;
 wire _06025_;
 wire _06026_;
 wire _06027_;
 wire _06028_;
 wire _06029_;
 wire _06030_;
 wire _06031_;
 wire _06032_;
 wire _06033_;
 wire _06034_;
 wire _06035_;
 wire _06036_;
 wire _06037_;
 wire _06038_;
 wire _06039_;
 wire _06040_;
 wire _06041_;
 wire _06042_;
 wire _06043_;
 wire _06044_;
 wire _06045_;
 wire _06046_;
 wire _06047_;
 wire _06048_;
 wire _06049_;
 wire _06050_;
 wire _06051_;
 wire _06052_;
 wire _06053_;
 wire _06054_;
 wire _06055_;
 wire _06056_;
 wire _06057_;
 wire _06058_;
 wire _06059_;
 wire _06060_;
 wire _06061_;
 wire _06062_;
 wire _06063_;
 wire _06064_;
 wire _06065_;
 wire _06066_;
 wire _06067_;
 wire _06068_;
 wire _06069_;
 wire _06070_;
 wire _06071_;
 wire _06072_;
 wire _06073_;
 wire _06074_;
 wire _06075_;
 wire _06076_;
 wire _06077_;
 wire _06078_;
 wire _06079_;
 wire _06080_;
 wire _06081_;
 wire _06082_;
 wire _06083_;
 wire _06084_;
 wire _06085_;
 wire _06086_;
 wire _06087_;
 wire _06088_;
 wire _06089_;
 wire _06090_;
 wire _06091_;
 wire _06092_;
 wire _06093_;
 wire _06094_;
 wire _06095_;
 wire _06096_;
 wire _06097_;
 wire _06098_;
 wire _06099_;
 wire _06100_;
 wire _06101_;
 wire _06102_;
 wire _06103_;
 wire _06104_;
 wire _06105_;
 wire _06106_;
 wire _06107_;
 wire _06108_;
 wire _06109_;
 wire _06110_;
 wire _06111_;
 wire _06112_;
 wire _06113_;
 wire _06114_;
 wire _06115_;
 wire _06116_;
 wire _06117_;
 wire _06118_;
 wire _06119_;
 wire _06120_;
 wire _06121_;
 wire _06122_;
 wire _06123_;
 wire _06124_;
 wire _06125_;
 wire _06126_;
 wire _06127_;
 wire _06128_;
 wire _06129_;
 wire _06130_;
 wire _06131_;
 wire _06132_;
 wire _06133_;
 wire _06134_;
 wire _06135_;
 wire _06136_;
 wire _06137_;
 wire _06138_;
 wire _06139_;
 wire _06140_;
 wire _06141_;
 wire _06142_;
 wire _06143_;
 wire _06144_;
 wire _06145_;
 wire _06146_;
 wire _06147_;
 wire _06148_;
 wire _06149_;
 wire _06150_;
 wire _06151_;
 wire _06152_;
 wire _06153_;
 wire _06154_;
 wire _06155_;
 wire _06156_;
 wire _06157_;
 wire _06158_;
 wire _06159_;
 wire _06160_;
 wire _06161_;
 wire _06162_;
 wire _06163_;
 wire _06164_;
 wire _06165_;
 wire _06166_;
 wire _06167_;
 wire _06168_;
 wire _06169_;
 wire _06170_;
 wire _06171_;
 wire _06172_;
 wire _06173_;
 wire _06174_;
 wire _06175_;
 wire _06176_;
 wire _06177_;
 wire _06178_;
 wire _06179_;
 wire _06180_;
 wire _06181_;
 wire _06182_;
 wire _06183_;
 wire _06184_;
 wire _06185_;
 wire _06186_;
 wire _06187_;
 wire _06188_;
 wire _06189_;
 wire _06190_;
 wire _06191_;
 wire _06192_;
 wire _06193_;
 wire _06194_;
 wire _06195_;
 wire _06196_;
 wire _06197_;
 wire _06198_;
 wire _06199_;
 wire _06200_;
 wire _06201_;
 wire _06202_;
 wire _06203_;
 wire _06204_;
 wire _06205_;
 wire _06206_;
 wire _06207_;
 wire _06208_;
 wire _06209_;
 wire _06210_;
 wire _06211_;
 wire _06212_;
 wire _06213_;
 wire _06214_;
 wire _06215_;
 wire _06216_;
 wire _06217_;
 wire _06218_;
 wire _06219_;
 wire _06220_;
 wire _06221_;
 wire _06222_;
 wire _06223_;
 wire _06224_;
 wire _06225_;
 wire _06226_;
 wire _06227_;
 wire _06228_;
 wire _06229_;
 wire _06230_;
 wire _06231_;
 wire _06232_;
 wire _06233_;
 wire _06234_;
 wire _06235_;
 wire _06236_;
 wire _06237_;
 wire _06238_;
 wire _06239_;
 wire _06240_;
 wire _06241_;
 wire _06242_;
 wire _06243_;
 wire _06244_;
 wire _06245_;
 wire _06246_;
 wire _06247_;
 wire _06248_;
 wire _06249_;
 wire _06250_;
 wire _06251_;
 wire _06252_;
 wire _06253_;
 wire _06254_;
 wire _06255_;
 wire _06256_;
 wire _06257_;
 wire _06258_;
 wire _06259_;
 wire _06260_;
 wire _06261_;
 wire _06262_;
 wire _06263_;
 wire _06264_;
 wire _06265_;
 wire _06266_;
 wire _06267_;
 wire _06268_;
 wire _06269_;
 wire _06270_;
 wire _06271_;
 wire _06272_;
 wire _06273_;
 wire _06274_;
 wire _06275_;
 wire _06276_;
 wire _06277_;
 wire _06278_;
 wire _06279_;
 wire _06280_;
 wire _06281_;
 wire _06282_;
 wire _06283_;
 wire _06284_;
 wire _06285_;
 wire _06286_;
 wire _06287_;
 wire _06288_;
 wire _06289_;
 wire _06290_;
 wire _06291_;
 wire _06292_;
 wire _06293_;
 wire _06294_;
 wire _06295_;
 wire _06296_;
 wire _06297_;
 wire _06298_;
 wire _06299_;
 wire _06300_;
 wire _06301_;
 wire _06302_;
 wire _06303_;
 wire _06304_;
 wire _06305_;
 wire _06306_;
 wire _06307_;
 wire _06308_;
 wire _06309_;
 wire _06310_;
 wire _06311_;
 wire _06312_;
 wire _06313_;
 wire _06314_;
 wire _06315_;
 wire _06316_;
 wire _06317_;
 wire _06318_;
 wire _06319_;
 wire _06320_;
 wire _06321_;
 wire _06322_;
 wire _06323_;
 wire _06324_;
 wire _06325_;
 wire _06326_;
 wire _06327_;
 wire _06328_;
 wire _06329_;
 wire _06330_;
 wire _06331_;
 wire _06332_;
 wire _06333_;
 wire _06334_;
 wire _06335_;
 wire _06336_;
 wire _06337_;
 wire _06338_;
 wire _06339_;
 wire _06340_;
 wire _06341_;
 wire _06342_;
 wire _06343_;
 wire _06344_;
 wire _06345_;
 wire _06346_;
 wire _06347_;
 wire _06348_;
 wire _06349_;
 wire _06350_;
 wire _06351_;
 wire _06352_;
 wire _06353_;
 wire _06354_;
 wire _06355_;
 wire _06356_;
 wire _06357_;
 wire _06358_;
 wire _06359_;
 wire _06360_;
 wire _06361_;
 wire _06362_;
 wire _06363_;
 wire _06364_;
 wire _06365_;
 wire _06366_;
 wire _06367_;
 wire _06368_;
 wire _06369_;
 wire _06370_;
 wire _06371_;
 wire _06372_;
 wire _06373_;
 wire _06374_;
 wire _06375_;
 wire _06376_;
 wire _06377_;
 wire _06378_;
 wire _06379_;
 wire _06380_;
 wire _06381_;
 wire _06382_;
 wire _06383_;
 wire _06384_;
 wire _06385_;
 wire _06386_;
 wire _06387_;
 wire _06388_;
 wire _06389_;
 wire _06390_;
 wire _06391_;
 wire _06392_;
 wire _06393_;
 wire _06394_;
 wire _06395_;
 wire _06396_;
 wire _06397_;
 wire _06398_;
 wire _06399_;
 wire _06400_;
 wire _06401_;
 wire _06402_;
 wire _06403_;
 wire _06404_;
 wire _06405_;
 wire _06406_;
 wire _06407_;
 wire _06408_;
 wire _06409_;
 wire _06410_;
 wire _06411_;
 wire _06412_;
 wire _06413_;
 wire _06414_;
 wire _06415_;
 wire _06416_;
 wire _06417_;
 wire _06418_;
 wire _06419_;
 wire _06420_;
 wire _06421_;
 wire _06422_;
 wire _06423_;
 wire _06424_;
 wire _06425_;
 wire _06426_;
 wire _06427_;
 wire _06428_;
 wire _06429_;
 wire _06430_;
 wire _06431_;
 wire _06432_;
 wire _06433_;
 wire _06434_;
 wire _06435_;
 wire _06436_;
 wire _06437_;
 wire _06438_;
 wire _06439_;
 wire _06440_;
 wire _06441_;
 wire _06442_;
 wire _06443_;
 wire _06444_;
 wire _06445_;
 wire _06446_;
 wire _06447_;
 wire _06448_;
 wire _06449_;
 wire _06450_;
 wire _06451_;
 wire _06452_;
 wire _06453_;
 wire _06454_;
 wire _06455_;
 wire _06456_;
 wire _06457_;
 wire _06458_;
 wire _06459_;
 wire _06460_;
 wire _06461_;
 wire _06462_;
 wire _06463_;
 wire _06464_;
 wire _06465_;
 wire _06466_;
 wire _06467_;
 wire _06468_;
 wire _06469_;
 wire _06470_;
 wire _06471_;
 wire _06472_;
 wire _06473_;
 wire _06474_;
 wire _06475_;
 wire _06476_;
 wire _06477_;
 wire _06478_;
 wire _06479_;
 wire _06480_;
 wire _06481_;
 wire _06482_;
 wire _06483_;
 wire _06484_;
 wire _06485_;
 wire _06486_;
 wire _06487_;
 wire _06488_;
 wire _06489_;
 wire _06490_;
 wire _06491_;
 wire _06492_;
 wire _06493_;
 wire _06494_;
 wire _06495_;
 wire _06496_;
 wire _06497_;
 wire _06498_;
 wire _06499_;
 wire _06500_;
 wire _06501_;
 wire _06502_;
 wire _06503_;
 wire _06504_;
 wire _06505_;
 wire _06506_;
 wire _06507_;
 wire _06508_;
 wire _06509_;
 wire _06510_;
 wire _06511_;
 wire _06512_;
 wire _06513_;
 wire _06514_;
 wire _06515_;
 wire _06516_;
 wire _06517_;
 wire _06518_;
 wire _06519_;
 wire _06520_;
 wire _06521_;
 wire _06522_;
 wire _06523_;
 wire _06524_;
 wire _06525_;
 wire _06526_;
 wire _06527_;
 wire _06528_;
 wire _06529_;
 wire _06530_;
 wire _06531_;
 wire _06532_;
 wire _06533_;
 wire _06534_;
 wire _06535_;
 wire _06536_;
 wire _06537_;
 wire _06538_;
 wire _06539_;
 wire _06540_;
 wire _06541_;
 wire _06542_;
 wire _06543_;
 wire _06544_;
 wire _06545_;
 wire _06546_;
 wire _06547_;
 wire _06548_;
 wire _06549_;
 wire _06550_;
 wire _06551_;
 wire _06552_;
 wire _06553_;
 wire _06554_;
 wire _06555_;
 wire _06556_;
 wire _06557_;
 wire _06558_;
 wire _06559_;
 wire _06560_;
 wire _06561_;
 wire _06562_;
 wire _06563_;
 wire _06564_;
 wire _06565_;
 wire _06566_;
 wire _06567_;
 wire _06568_;
 wire _06569_;
 wire _06570_;
 wire _06571_;
 wire _06572_;
 wire _06573_;
 wire _06574_;
 wire _06575_;
 wire _06576_;
 wire _06577_;
 wire _06578_;
 wire _06579_;
 wire _06580_;
 wire _06581_;
 wire _06582_;
 wire _06583_;
 wire _06584_;
 wire _06585_;
 wire _06586_;
 wire _06587_;
 wire _06588_;
 wire _06589_;
 wire _06590_;
 wire _06591_;
 wire _06592_;
 wire _06593_;
 wire _06594_;
 wire _06595_;
 wire _06596_;
 wire _06597_;
 wire _06598_;
 wire _06599_;
 wire _06600_;
 wire _06601_;
 wire _06602_;
 wire _06603_;
 wire _06604_;
 wire _06605_;
 wire _06606_;
 wire _06607_;
 wire _06608_;
 wire _06609_;
 wire _06610_;
 wire _06611_;
 wire _06612_;
 wire _06613_;
 wire _06614_;
 wire _06615_;
 wire _06616_;
 wire _06617_;
 wire _06618_;
 wire _06619_;
 wire _06620_;
 wire _06621_;
 wire _06622_;
 wire _06623_;
 wire _06624_;
 wire _06625_;
 wire _06626_;
 wire _06627_;
 wire _06628_;
 wire _06629_;
 wire _06630_;
 wire _06631_;
 wire _06632_;
 wire _06633_;
 wire _06634_;
 wire _06635_;
 wire _06636_;
 wire _06637_;
 wire _06638_;
 wire _06639_;
 wire _06640_;
 wire _06641_;
 wire _06642_;
 wire _06643_;
 wire _06644_;
 wire _06645_;
 wire _06646_;
 wire _06647_;
 wire _06648_;
 wire _06649_;
 wire _06650_;
 wire _06651_;
 wire _06652_;
 wire _06653_;
 wire _06654_;
 wire _06655_;
 wire _06656_;
 wire _06657_;
 wire _06658_;
 wire _06659_;
 wire _06660_;
 wire _06661_;
 wire _06662_;
 wire _06663_;
 wire _06664_;
 wire _06665_;
 wire _06666_;
 wire _06667_;
 wire _06668_;
 wire _06669_;
 wire _06670_;
 wire _06671_;
 wire _06672_;
 wire _06673_;
 wire _06674_;
 wire _06675_;
 wire _06676_;
 wire _06677_;
 wire _06678_;
 wire _06679_;
 wire _06680_;
 wire _06681_;
 wire _06682_;
 wire _06683_;
 wire _06684_;
 wire _06685_;
 wire _06686_;
 wire _06687_;
 wire _06688_;
 wire _06689_;
 wire _06690_;
 wire _06691_;
 wire _06692_;
 wire _06693_;
 wire _06694_;
 wire _06695_;
 wire _06696_;
 wire _06697_;
 wire _06698_;
 wire _06699_;
 wire _06700_;
 wire _06701_;
 wire _06702_;
 wire _06703_;
 wire _06704_;
 wire _06705_;
 wire _06706_;
 wire _06707_;
 wire _06708_;
 wire _06709_;
 wire _06710_;
 wire _06711_;
 wire _06712_;
 wire _06713_;
 wire _06714_;
 wire _06715_;
 wire _06716_;
 wire _06717_;
 wire _06718_;
 wire _06719_;
 wire _06720_;
 wire _06721_;
 wire _06722_;
 wire _06723_;
 wire _06724_;
 wire _06725_;
 wire _06726_;
 wire _06727_;
 wire _06728_;
 wire _06729_;
 wire _06730_;
 wire _06731_;
 wire _06732_;
 wire _06733_;
 wire _06734_;
 wire _06735_;
 wire _06736_;
 wire _06737_;
 wire _06738_;
 wire _06739_;
 wire _06740_;
 wire _06741_;
 wire _06742_;
 wire _06743_;
 wire _06744_;
 wire _06745_;
 wire _06746_;
 wire _06747_;
 wire _06748_;
 wire _06749_;
 wire _06750_;
 wire _06751_;
 wire _06752_;
 wire _06753_;
 wire _06754_;
 wire _06755_;
 wire _06756_;
 wire _06757_;
 wire _06758_;
 wire _06759_;
 wire _06760_;
 wire _06761_;
 wire _06762_;
 wire _06763_;
 wire _06764_;
 wire _06765_;
 wire _06766_;
 wire _06767_;
 wire _06768_;
 wire _06769_;
 wire _06770_;
 wire _06771_;
 wire _06772_;
 wire _06773_;
 wire _06774_;
 wire _06775_;
 wire _06776_;
 wire _06777_;
 wire _06778_;
 wire _06779_;
 wire _06780_;
 wire _06781_;
 wire _06782_;
 wire _06783_;
 wire _06784_;
 wire _06785_;
 wire _06786_;
 wire _06787_;
 wire _06788_;
 wire _06789_;
 wire _06790_;
 wire _06791_;
 wire _06792_;
 wire _06793_;
 wire _06794_;
 wire _06795_;
 wire _06796_;
 wire _06797_;
 wire _06798_;
 wire _06799_;
 wire _06800_;
 wire _06801_;
 wire _06802_;
 wire _06803_;
 wire _06804_;
 wire _06805_;
 wire _06806_;
 wire _06807_;
 wire _06808_;
 wire _06809_;
 wire _06810_;
 wire _06811_;
 wire _06812_;
 wire _06813_;
 wire _06814_;
 wire _06815_;
 wire _06816_;
 wire _06817_;
 wire _06818_;
 wire _06819_;
 wire _06820_;
 wire _06821_;
 wire _06822_;
 wire _06823_;
 wire _06824_;
 wire _06825_;
 wire _06826_;
 wire _06827_;
 wire _06828_;
 wire _06829_;
 wire _06830_;
 wire _06831_;
 wire _06832_;
 wire _06833_;
 wire _06834_;
 wire _06835_;
 wire _06836_;
 wire _06837_;
 wire _06838_;
 wire _06839_;
 wire _06840_;
 wire _06841_;
 wire _06842_;
 wire _06843_;
 wire _06844_;
 wire _06845_;
 wire _06846_;
 wire _06847_;
 wire _06848_;
 wire _06849_;
 wire _06850_;
 wire _06851_;
 wire _06852_;
 wire _06853_;
 wire _06854_;
 wire _06855_;
 wire _06856_;
 wire _06857_;
 wire _06858_;
 wire _06859_;
 wire _06860_;
 wire _06861_;
 wire _06862_;
 wire _06863_;
 wire _06864_;
 wire _06865_;
 wire _06866_;
 wire _06867_;
 wire _06868_;
 wire _06869_;
 wire _06870_;
 wire _06871_;
 wire _06872_;
 wire _06873_;
 wire _06874_;
 wire _06875_;
 wire _06876_;
 wire _06877_;
 wire _06878_;
 wire _06879_;
 wire _06880_;
 wire _06881_;
 wire _06882_;
 wire _06883_;
 wire _06884_;
 wire _06885_;
 wire _06886_;
 wire _06887_;
 wire _06888_;
 wire _06889_;
 wire _06890_;
 wire _06891_;
 wire _06892_;
 wire _06893_;
 wire _06894_;
 wire _06895_;
 wire _06896_;
 wire _06897_;
 wire _06898_;
 wire _06899_;
 wire _06900_;
 wire _06901_;
 wire _06902_;
 wire _06903_;
 wire _06904_;
 wire _06905_;
 wire _06906_;
 wire _06907_;
 wire _06908_;
 wire _06909_;
 wire _06910_;
 wire _06911_;
 wire _06912_;
 wire _06913_;
 wire _06914_;
 wire _06915_;
 wire _06916_;
 wire _06917_;
 wire _06918_;
 wire _06919_;
 wire _06920_;
 wire _06921_;
 wire _06922_;
 wire _06923_;
 wire _06924_;
 wire _06925_;
 wire _06926_;
 wire _06927_;
 wire _06928_;
 wire _06929_;
 wire _06930_;
 wire _06931_;
 wire _06932_;
 wire _06933_;
 wire _06934_;
 wire _06935_;
 wire _06936_;
 wire _06937_;
 wire _06938_;
 wire _06939_;
 wire _06940_;
 wire _06941_;
 wire _06942_;
 wire _06943_;
 wire _06944_;
 wire _06945_;
 wire _06946_;
 wire _06947_;
 wire _06948_;
 wire _06949_;
 wire _06950_;
 wire _06951_;
 wire _06952_;
 wire _06953_;
 wire _06954_;
 wire _06955_;
 wire _06956_;
 wire _06957_;
 wire _06958_;
 wire _06959_;
 wire _06960_;
 wire _06961_;
 wire _06962_;
 wire _06963_;
 wire _06964_;
 wire _06965_;
 wire _06966_;
 wire _06967_;
 wire _06968_;
 wire _06969_;
 wire _06970_;
 wire _06971_;
 wire _06972_;
 wire _06973_;
 wire _06974_;
 wire _06975_;
 wire _06976_;
 wire _06977_;
 wire _06978_;
 wire _06979_;
 wire _06980_;
 wire _06981_;
 wire _06982_;
 wire _06983_;
 wire _06984_;
 wire _06985_;
 wire _06986_;
 wire _06987_;
 wire _06988_;
 wire _06989_;
 wire _06990_;
 wire _06991_;
 wire _06992_;
 wire _06993_;
 wire _06994_;
 wire _06995_;
 wire _06996_;
 wire _06997_;
 wire _06998_;
 wire _06999_;
 wire _07000_;
 wire _07001_;
 wire _07002_;
 wire _07003_;
 wire _07004_;
 wire _07005_;
 wire _07006_;
 wire _07007_;
 wire _07008_;
 wire _07009_;
 wire _07010_;
 wire _07011_;
 wire _07012_;
 wire _07013_;
 wire _07014_;
 wire _07015_;
 wire _07016_;
 wire _07017_;
 wire _07018_;
 wire _07019_;
 wire _07020_;
 wire _07021_;
 wire _07022_;
 wire _07023_;
 wire _07024_;
 wire _07025_;
 wire _07026_;
 wire _07027_;
 wire _07028_;
 wire _07029_;
 wire _07030_;
 wire _07031_;
 wire _07032_;
 wire _07033_;
 wire _07034_;
 wire _07035_;
 wire _07036_;
 wire _07037_;
 wire _07038_;
 wire _07039_;
 wire _07040_;
 wire _07041_;
 wire _07042_;
 wire _07043_;
 wire _07044_;
 wire _07045_;
 wire _07046_;
 wire _07047_;
 wire _07048_;
 wire _07049_;
 wire _07050_;
 wire _07051_;
 wire _07052_;
 wire _07053_;
 wire _07054_;
 wire _07055_;
 wire _07056_;
 wire _07057_;
 wire _07058_;
 wire _07059_;
 wire _07060_;
 wire _07061_;
 wire _07062_;
 wire _07063_;
 wire _07064_;
 wire _07065_;
 wire _07066_;
 wire _07067_;
 wire _07068_;
 wire _07069_;
 wire _07070_;
 wire _07071_;
 wire _07072_;
 wire _07073_;
 wire _07074_;
 wire _07075_;
 wire _07076_;
 wire _07077_;
 wire _07078_;
 wire _07079_;
 wire _07080_;
 wire _07081_;
 wire _07082_;
 wire _07083_;
 wire _07084_;
 wire _07085_;
 wire _07086_;
 wire _07087_;
 wire _07088_;
 wire _07089_;
 wire _07090_;
 wire _07091_;
 wire _07092_;
 wire _07093_;
 wire _07094_;
 wire _07095_;
 wire _07096_;
 wire _07097_;
 wire _07098_;
 wire _07099_;
 wire _07100_;
 wire _07101_;
 wire _07102_;
 wire _07103_;
 wire _07104_;
 wire _07105_;
 wire _07106_;
 wire _07107_;
 wire _07108_;
 wire _07109_;
 wire _07110_;
 wire _07111_;
 wire _07112_;
 wire _07113_;
 wire _07114_;
 wire _07115_;
 wire _07116_;
 wire _07117_;
 wire _07118_;
 wire _07119_;
 wire _07120_;
 wire _07121_;
 wire _07122_;
 wire _07123_;
 wire _07124_;
 wire _07125_;
 wire _07126_;
 wire _07127_;
 wire _07128_;
 wire _07129_;
 wire _07130_;
 wire _07131_;
 wire _07132_;
 wire _07133_;
 wire _07134_;
 wire _07135_;
 wire _07136_;
 wire _07137_;
 wire _07138_;
 wire _07139_;
 wire _07140_;
 wire _07141_;
 wire _07142_;
 wire _07143_;
 wire _07144_;
 wire _07145_;
 wire _07146_;
 wire _07147_;
 wire _07148_;
 wire _07149_;
 wire _07150_;
 wire _07151_;
 wire _07152_;
 wire _07153_;
 wire _07154_;
 wire _07155_;
 wire _07156_;
 wire _07157_;
 wire _07158_;
 wire _07159_;
 wire _07160_;
 wire _07161_;
 wire _07162_;
 wire _07163_;
 wire _07164_;
 wire _07165_;
 wire _07166_;
 wire _07167_;
 wire _07168_;
 wire _07169_;
 wire _07170_;
 wire _07171_;
 wire _07172_;
 wire _07173_;
 wire _07174_;
 wire _07175_;
 wire _07176_;
 wire _07177_;
 wire _07178_;
 wire _07179_;
 wire _07180_;
 wire _07181_;
 wire _07182_;
 wire _07183_;
 wire _07184_;
 wire _07185_;
 wire _07186_;
 wire _07187_;
 wire _07188_;
 wire _07189_;
 wire _07190_;
 wire _07191_;
 wire _07192_;
 wire _07193_;
 wire _07194_;
 wire _07195_;
 wire _07196_;
 wire _07197_;
 wire _07198_;
 wire _07199_;
 wire _07200_;
 wire _07201_;
 wire _07202_;
 wire _07203_;
 wire _07204_;
 wire _07205_;
 wire _07206_;
 wire _07207_;
 wire _07208_;
 wire _07209_;
 wire _07210_;
 wire _07211_;
 wire _07212_;
 wire _07213_;
 wire _07214_;
 wire _07215_;
 wire _07216_;
 wire _07217_;
 wire _07218_;
 wire _07219_;
 wire _07220_;
 wire _07221_;
 wire _07222_;
 wire _07223_;
 wire _07224_;
 wire _07225_;
 wire _07226_;
 wire _07227_;
 wire _07228_;
 wire _07229_;
 wire _07230_;
 wire _07231_;
 wire _07232_;
 wire _07233_;
 wire _07234_;
 wire _07235_;
 wire _07236_;
 wire _07237_;
 wire _07238_;
 wire _07239_;
 wire _07240_;
 wire _07241_;
 wire _07242_;
 wire _07243_;
 wire _07244_;
 wire _07245_;
 wire _07246_;
 wire _07247_;
 wire _07248_;
 wire _07249_;
 wire _07250_;
 wire _07251_;
 wire _07252_;
 wire _07253_;
 wire _07254_;
 wire _07255_;
 wire _07256_;
 wire _07257_;
 wire _07258_;
 wire _07259_;
 wire _07260_;
 wire _07261_;
 wire _07262_;
 wire _07263_;
 wire _07264_;
 wire _07265_;
 wire _07266_;
 wire _07267_;
 wire _07268_;
 wire _07269_;
 wire _07270_;
 wire _07271_;
 wire _07272_;
 wire _07273_;
 wire _07274_;
 wire _07275_;
 wire _07276_;
 wire _07277_;
 wire _07278_;
 wire _07279_;
 wire _07280_;
 wire _07281_;
 wire _07282_;
 wire _07283_;
 wire _07284_;
 wire _07285_;
 wire _07286_;
 wire _07287_;
 wire _07288_;
 wire _07289_;
 wire _07290_;
 wire _07291_;
 wire _07292_;
 wire _07293_;
 wire _07294_;
 wire _07295_;
 wire _07296_;
 wire _07297_;
 wire _07298_;
 wire _07299_;
 wire _07300_;
 wire _07301_;
 wire _07302_;
 wire _07303_;
 wire _07304_;
 wire _07305_;
 wire _07306_;
 wire _07307_;
 wire _07308_;
 wire _07309_;
 wire _07310_;
 wire _07311_;
 wire _07312_;
 wire _07313_;
 wire _07314_;
 wire _07315_;
 wire _07316_;
 wire _07317_;
 wire _07318_;
 wire _07319_;
 wire _07320_;
 wire _07321_;
 wire _07322_;
 wire _07323_;
 wire _07324_;
 wire _07325_;
 wire _07326_;
 wire _07327_;
 wire _07328_;
 wire _07329_;
 wire _07330_;
 wire _07331_;
 wire _07332_;
 wire _07333_;
 wire _07334_;
 wire _07335_;
 wire _07336_;
 wire _07337_;
 wire _07338_;
 wire _07339_;
 wire _07340_;
 wire _07341_;
 wire _07342_;
 wire _07343_;
 wire _07344_;
 wire _07345_;
 wire _07346_;
 wire _07347_;
 wire _07348_;
 wire _07349_;
 wire _07350_;
 wire _07351_;
 wire _07352_;
 wire _07353_;
 wire _07354_;
 wire _07355_;
 wire _07356_;
 wire _07357_;
 wire _07358_;
 wire _07359_;
 wire _07360_;
 wire _07361_;
 wire _07362_;
 wire _07363_;
 wire _07364_;
 wire _07365_;
 wire _07366_;
 wire _07367_;
 wire _07368_;
 wire _07369_;
 wire _07370_;
 wire _07371_;
 wire _07372_;
 wire _07373_;
 wire _07374_;
 wire _07375_;
 wire _07376_;
 wire _07377_;
 wire _07378_;
 wire _07379_;
 wire _07380_;
 wire _07381_;
 wire _07382_;
 wire _07383_;
 wire _07384_;
 wire _07385_;
 wire _07386_;
 wire _07387_;
 wire _07388_;
 wire _07389_;
 wire _07390_;
 wire _07391_;
 wire _07392_;
 wire _07393_;
 wire _07394_;
 wire _07395_;
 wire _07396_;
 wire _07397_;
 wire _07398_;
 wire _07399_;
 wire _07400_;
 wire _07401_;
 wire _07402_;
 wire _07403_;
 wire _07404_;
 wire _07405_;
 wire _07406_;
 wire _07407_;
 wire _07408_;
 wire _07409_;
 wire _07410_;
 wire _07411_;
 wire _07412_;
 wire _07413_;
 wire _07414_;
 wire _07415_;
 wire _07416_;
 wire _07417_;
 wire _07418_;
 wire _07419_;
 wire _07420_;
 wire _07421_;
 wire _07422_;
 wire _07423_;
 wire _07424_;
 wire _07425_;
 wire _07426_;
 wire _07427_;
 wire _07428_;
 wire _07429_;
 wire _07430_;
 wire _07431_;
 wire _07432_;
 wire _07433_;
 wire _07434_;
 wire _07435_;
 wire _07436_;
 wire _07437_;
 wire _07438_;
 wire _07439_;
 wire _07440_;
 wire _07441_;
 wire _07442_;
 wire _07443_;
 wire _07444_;
 wire _07445_;
 wire _07446_;
 wire _07447_;
 wire _07448_;
 wire _07449_;
 wire _07450_;
 wire _07451_;
 wire _07452_;
 wire _07453_;
 wire _07454_;
 wire _07455_;
 wire _07456_;
 wire _07457_;
 wire _07458_;
 wire _07459_;
 wire _07460_;
 wire _07461_;
 wire _07462_;
 wire _07463_;
 wire _07464_;
 wire _07465_;
 wire _07466_;
 wire _07467_;
 wire _07468_;
 wire _07469_;
 wire _07470_;
 wire _07471_;
 wire _07472_;
 wire _07473_;
 wire _07474_;
 wire _07475_;
 wire _07476_;
 wire _07477_;
 wire _07478_;
 wire _07479_;
 wire _07480_;
 wire _07481_;
 wire _07482_;
 wire _07483_;
 wire _07484_;
 wire _07485_;
 wire _07486_;
 wire _07487_;
 wire _07488_;
 wire _07489_;
 wire _07490_;
 wire _07491_;
 wire _07492_;
 wire _07493_;
 wire _07494_;
 wire _07495_;
 wire _07496_;
 wire _07497_;
 wire _07498_;
 wire _07499_;
 wire _07500_;
 wire _07501_;
 wire _07502_;
 wire _07503_;
 wire _07504_;
 wire _07505_;
 wire _07506_;
 wire _07507_;
 wire _07508_;
 wire _07509_;
 wire _07510_;
 wire _07511_;
 wire _07512_;
 wire _07513_;
 wire _07514_;
 wire _07515_;
 wire _07516_;
 wire _07517_;
 wire _07518_;
 wire _07519_;
 wire _07520_;
 wire _07521_;
 wire _07522_;
 wire _07523_;
 wire _07524_;
 wire _07525_;
 wire _07526_;
 wire _07527_;
 wire _07528_;
 wire _07529_;
 wire _07530_;
 wire _07531_;
 wire _07532_;
 wire _07533_;
 wire _07534_;
 wire _07535_;
 wire _07536_;
 wire _07537_;
 wire _07538_;
 wire _07539_;
 wire _07540_;
 wire _07541_;
 wire _07542_;
 wire _07543_;
 wire _07544_;
 wire _07545_;
 wire _07546_;
 wire _07547_;
 wire _07548_;
 wire _07549_;
 wire _07550_;
 wire _07551_;
 wire _07552_;
 wire _07553_;
 wire _07554_;
 wire _07555_;
 wire _07556_;
 wire _07557_;
 wire _07558_;
 wire _07559_;
 wire _07560_;
 wire _07561_;
 wire _07562_;
 wire _07563_;
 wire _07564_;
 wire _07565_;
 wire _07566_;
 wire _07567_;
 wire _07568_;
 wire _07569_;
 wire _07570_;
 wire _07571_;
 wire _07572_;
 wire _07573_;
 wire _07574_;
 wire _07575_;
 wire _07576_;
 wire _07577_;
 wire _07578_;
 wire _07579_;
 wire _07580_;
 wire _07581_;
 wire _07582_;
 wire _07583_;
 wire _07584_;
 wire _07585_;
 wire _07586_;
 wire _07587_;
 wire _07588_;
 wire _07589_;
 wire _07590_;
 wire _07591_;
 wire _07592_;
 wire _07593_;
 wire _07594_;
 wire _07595_;
 wire _07596_;
 wire _07597_;
 wire _07598_;
 wire _07599_;
 wire _07600_;
 wire _07601_;
 wire _07602_;
 wire _07603_;
 wire _07604_;
 wire _07605_;
 wire _07606_;
 wire _07607_;
 wire _07608_;
 wire _07609_;
 wire _07610_;
 wire _07611_;
 wire _07612_;
 wire _07613_;
 wire _07614_;
 wire _07615_;
 wire _07616_;
 wire _07617_;
 wire _07618_;
 wire _07619_;
 wire _07620_;
 wire _07621_;
 wire _07622_;
 wire _07623_;
 wire _07624_;
 wire _07625_;
 wire _07626_;
 wire _07627_;
 wire _07628_;
 wire _07629_;
 wire _07630_;
 wire _07631_;
 wire _07632_;
 wire _07633_;
 wire _07634_;
 wire _07635_;
 wire _07636_;
 wire _07637_;
 wire _07638_;
 wire _07639_;
 wire _07640_;
 wire _07641_;
 wire _07642_;
 wire _07643_;
 wire _07644_;
 wire _07645_;
 wire _07646_;
 wire _07647_;
 wire _07648_;
 wire _07649_;
 wire _07650_;
 wire _07651_;
 wire _07652_;
 wire _07653_;
 wire _07654_;
 wire _07655_;
 wire _07656_;
 wire _07657_;
 wire _07658_;
 wire _07659_;
 wire _07660_;
 wire _07661_;
 wire _07662_;
 wire _07663_;
 wire _07664_;
 wire _07665_;
 wire _07666_;
 wire _07667_;
 wire _07668_;
 wire _07669_;
 wire _07670_;
 wire clknet_leaf_0_clk;
 wire net353;
 wire \i_coord.demo_update ;
 wire \i_coord.demo_update_delay ;
 wire \i_coord.l_xip.data_out[0] ;
 wire \i_coord.l_xip.data_out[1] ;
 wire \i_coord.l_xip.data_out[2] ;
 wire \i_coord.l_xip.data_out[3] ;
 wire \i_coord.l_xip.data_out[4] ;
 wire \i_coord.l_xip.data_out[5] ;
 wire \i_coord.l_xip.data_out[6] ;
 wire \i_coord.l_xip.data_out[7] ;
 wire \i_coord.l_xip.data_out[8] ;
 wire \i_coord.l_xip.data_out[9] ;
 wire \i_coord.l_xir.data_out[0] ;
 wire \i_coord.l_xir.data_out[1] ;
 wire \i_coord.l_xir.data_out[2] ;
 wire \i_coord.l_xir.data_out[3] ;
 wire \i_coord.l_xir.data_out[4] ;
 wire \i_coord.l_xir.data_out[5] ;
 wire \i_coord.l_xir.data_out[6] ;
 wire \i_coord.l_xir.data_out[7] ;
 wire \i_coord.l_xl.data_out[10] ;
 wire \i_coord.l_xl.data_out[11] ;
 wire \i_coord.l_xl.data_out[12] ;
 wire \i_coord.l_xl.data_out[13] ;
 wire \i_coord.l_xl.data_out[14] ;
 wire \i_coord.l_xl.data_out[15] ;
 wire \i_coord.l_xl.data_out[3] ;
 wire \i_coord.l_xl.data_out[4] ;
 wire \i_coord.l_xl.data_out[5] ;
 wire \i_coord.l_xl.data_out[6] ;
 wire \i_coord.l_xl.data_out[7] ;
 wire \i_coord.l_xl.data_out[8] ;
 wire \i_coord.l_xl.data_out[9] ;
 wire \i_coord.l_yip.data_out[0] ;
 wire \i_coord.l_yip.data_out[1] ;
 wire \i_coord.l_yip.data_out[2] ;
 wire \i_coord.l_yip.data_out[3] ;
 wire \i_coord.l_yip.data_out[4] ;
 wire \i_coord.l_yip.data_out[5] ;
 wire \i_coord.l_yip.data_out[6] ;
 wire \i_coord.l_yip.data_out[7] ;
 wire \i_coord.l_yip.data_out[8] ;
 wire \i_coord.l_yip.data_out[9] ;
 wire \i_coord.l_yt.data_out[0] ;
 wire \i_coord.l_yt.data_out[10] ;
 wire \i_coord.l_yt.data_out[11] ;
 wire \i_coord.l_yt.data_out[12] ;
 wire \i_coord.l_yt.data_out[13] ;
 wire \i_coord.l_yt.data_out[14] ;
 wire \i_coord.l_yt.data_out[1] ;
 wire \i_coord.l_yt.data_out[2] ;
 wire \i_coord.l_yt.data_out[3] ;
 wire \i_coord.l_yt.data_out[4] ;
 wire \i_coord.l_yt.data_out[5] ;
 wire \i_coord.l_yt.data_out[6] ;
 wire \i_coord.l_yt.data_out[7] ;
 wire \i_coord.l_yt.data_out[8] ;
 wire \i_coord.l_yt.data_out[9] ;
 wire \i_coord.x0[-10] ;
 wire \i_coord.x0[-11] ;
 wire \i_coord.x0[-12] ;
 wire \i_coord.x0[-13] ;
 wire \i_coord.x0[-1] ;
 wire \i_coord.x0[-2] ;
 wire \i_coord.x0[-3] ;
 wire \i_coord.x0[-4] ;
 wire \i_coord.x0[-5] ;
 wire \i_coord.x0[-6] ;
 wire \i_coord.x0[-7] ;
 wire \i_coord.x0[-8] ;
 wire \i_coord.x0[-9] ;
 wire \i_coord.x0[0] ;
 wire \i_coord.x0[1] ;
 wire \i_coord.x0[2] ;
 wire \i_coord.x_row_start[-10] ;
 wire \i_coord.x_row_start[-11] ;
 wire \i_coord.x_row_start[-12] ;
 wire \i_coord.x_row_start[-13] ;
 wire \i_coord.x_row_start[-1] ;
 wire \i_coord.x_row_start[-2] ;
 wire \i_coord.x_row_start[-3] ;
 wire \i_coord.x_row_start[-4] ;
 wire \i_coord.x_row_start[-5] ;
 wire \i_coord.x_row_start[-6] ;
 wire \i_coord.x_row_start[-7] ;
 wire \i_coord.x_row_start[-8] ;
 wire \i_coord.x_row_start[-9] ;
 wire \i_coord.x_row_start[0] ;
 wire \i_coord.x_row_start[1] ;
 wire \i_coord.x_row_start[2] ;
 wire \i_coord.y0[-10] ;
 wire \i_coord.y0[-11] ;
 wire \i_coord.y0[-12] ;
 wire \i_coord.y0[-13] ;
 wire \i_coord.y0[-1] ;
 wire \i_coord.y0[-2] ;
 wire \i_coord.y0[-3] ;
 wire \i_coord.y0[-4] ;
 wire \i_coord.y0[-5] ;
 wire \i_coord.y0[-6] ;
 wire \i_coord.y0[-7] ;
 wire \i_coord.y0[-8] ;
 wire \i_coord.y0[-9] ;
 wire \i_coord.y0[0] ;
 wire \i_coord.y0[1] ;
 wire \i_coord.y_inc_row[-10] ;
 wire \i_coord.y_inc_row[-11] ;
 wire \i_coord.y_inc_row[-12] ;
 wire \i_coord.y_inc_row[-13] ;
 wire \i_coord.y_inc_row[-6] ;
 wire \i_coord.y_inc_row[-7] ;
 wire \i_coord.y_inc_row[-8] ;
 wire \i_coord.y_inc_row[-9] ;
 wire \i_coord.y_row_start[-10] ;
 wire \i_coord.y_row_start[-11] ;
 wire \i_coord.y_row_start[-12] ;
 wire \i_coord.y_row_start[-13] ;
 wire \i_coord.y_row_start[-1] ;
 wire \i_coord.y_row_start[-2] ;
 wire \i_coord.y_row_start[-3] ;
 wire \i_coord.y_row_start[-4] ;
 wire \i_coord.y_row_start[-5] ;
 wire \i_coord.y_row_start[-6] ;
 wire \i_coord.y_row_start[-7] ;
 wire \i_coord.y_row_start[-8] ;
 wire \i_coord.y_row_start[-9] ;
 wire \i_coord.y_row_start[0] ;
 wire \i_coord.y_row_start[1] ;
 wire \i_mandel.i_sq_x.x[-10] ;
 wire \i_mandel.i_sq_x.x[-11] ;
 wire \i_mandel.i_sq_x.x[-12] ;
 wire \i_mandel.i_sq_x.x[-13] ;
 wire \i_mandel.i_sq_x.x[-1] ;
 wire \i_mandel.i_sq_x.x[-2] ;
 wire \i_mandel.i_sq_x.x[-3] ;
 wire \i_mandel.i_sq_x.x[-4] ;
 wire \i_mandel.i_sq_x.x[-5] ;
 wire \i_mandel.i_sq_x.x[-6] ;
 wire \i_mandel.i_sq_x.x[-7] ;
 wire \i_mandel.i_sq_x.x[-8] ;
 wire \i_mandel.i_sq_x.x[-9] ;
 wire \i_mandel.i_sq_x.x[0] ;
 wire \i_mandel.i_sq_x.x[1] ;
 wire \i_mandel.i_sq_x.x[2] ;
 wire \i_mandel.i_sq_y.x[-10] ;
 wire \i_mandel.i_sq_y.x[-11] ;
 wire \i_mandel.i_sq_y.x[-12] ;
 wire \i_mandel.i_sq_y.x[-13] ;
 wire \i_mandel.i_sq_y.x[-1] ;
 wire \i_mandel.i_sq_y.x[-2] ;
 wire \i_mandel.i_sq_y.x[-3] ;
 wire \i_mandel.i_sq_y.x[-4] ;
 wire \i_mandel.i_sq_y.x[-5] ;
 wire \i_mandel.i_sq_y.x[-6] ;
 wire \i_mandel.i_sq_y.x[-7] ;
 wire \i_mandel.i_sq_y.x[-8] ;
 wire \i_mandel.i_sq_y.x[-9] ;
 wire \i_mandel.i_sq_y.x[0] ;
 wire \i_mandel.i_sq_y.x[1] ;
 wire \i_mandel.i_sq_y.x[2] ;
 wire \i_vga.hsync ;
 wire \i_vga.timing_hor.counter[0] ;
 wire \i_vga.timing_hor.counter[10] ;
 wire \i_vga.timing_hor.counter[1] ;
 wire \i_vga.timing_hor.counter[2] ;
 wire \i_vga.timing_hor.counter[3] ;
 wire \i_vga.timing_hor.counter[4] ;
 wire \i_vga.timing_hor.counter[5] ;
 wire \i_vga.timing_hor.counter[6] ;
 wire \i_vga.timing_hor.counter[7] ;
 wire \i_vga.timing_hor.counter[8] ;
 wire \i_vga.timing_hor.counter[9] ;
 wire \i_vga.timing_ver.blank ;
 wire \i_vga.timing_ver.counter[0] ;
 wire \i_vga.timing_ver.counter[1] ;
 wire \i_vga.timing_ver.counter[2] ;
 wire \i_vga.timing_ver.counter[3] ;
 wire \i_vga.timing_ver.counter[4] ;
 wire \i_vga.timing_ver.counter[5] ;
 wire \i_vga.timing_ver.counter[6] ;
 wire \i_vga.timing_ver.counter[7] ;
 wire \i_vga.timing_ver.counter[8] ;
 wire \i_vga.timing_ver.counter[9] ;
 wire \i_vga.timing_ver.sync ;
 wire \i_vga.timing_ver.sync_tmp ;
 wire \i_vga.vblank ;
 wire \iter[0] ;
 wire \iter[1] ;
 wire \iter[2] ;
 wire \iter[3] ;
 wire \last_iter[0] ;
 wire \last_iter[1] ;
 wire \last_iter[2] ;
 wire \last_iter[3] ;
 wire \last_iter[4] ;
 wire \step[0] ;
 wire \step[1] ;
 wire \step[2] ;
 wire \step[3] ;
 wire \video_colour[0] ;
 wire \video_colour[1] ;
 wire \video_colour[2] ;
 wire \video_colour[3] ;
 wire \video_colour[4] ;
 wire \video_colour[5] ;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net180;
 wire net181;
 wire net182;
 wire net183;
 wire net184;
 wire net185;
 wire net186;
 wire net187;
 wire net188;
 wire net189;
 wire net190;
 wire net191;
 wire net192;
 wire net193;
 wire net194;
 wire net195;
 wire net196;
 wire net197;
 wire net198;
 wire net199;
 wire net200;
 wire net201;
 wire net202;
 wire net203;
 wire net204;
 wire net205;
 wire net206;
 wire net207;
 wire net208;
 wire net209;
 wire net210;
 wire net211;
 wire net212;
 wire net213;
 wire net214;
 wire net215;
 wire net216;
 wire net217;
 wire net218;
 wire net219;
 wire net220;
 wire net221;
 wire net222;
 wire net223;
 wire net224;
 wire net225;
 wire net226;
 wire net227;
 wire net228;
 wire net229;
 wire net230;
 wire net231;
 wire net232;
 wire net233;
 wire net234;
 wire net235;
 wire net236;
 wire net237;
 wire net238;
 wire net239;
 wire net240;
 wire net241;
 wire net242;
 wire net243;
 wire net244;
 wire net245;
 wire net246;
 wire net247;
 wire net248;
 wire net249;
 wire net250;
 wire net251;
 wire net252;
 wire net253;
 wire net254;
 wire net255;
 wire net256;
 wire net257;
 wire net258;
 wire net259;
 wire net260;
 wire net261;
 wire net262;
 wire net263;
 wire net264;
 wire net265;
 wire net266;
 wire net267;
 wire net268;
 wire net269;
 wire net270;
 wire net271;
 wire net272;
 wire net273;
 wire net274;
 wire net275;
 wire net276;
 wire net277;
 wire net278;
 wire net279;
 wire net280;
 wire net281;
 wire net282;
 wire net283;
 wire net284;
 wire net285;
 wire net286;
 wire net287;
 wire net288;
 wire net289;
 wire net290;
 wire net291;
 wire net292;
 wire net293;
 wire net294;
 wire net295;
 wire net296;
 wire net297;
 wire net298;
 wire net299;
 wire net300;
 wire net301;
 wire net302;
 wire net303;
 wire net304;
 wire net305;
 wire net306;
 wire net307;
 wire net308;
 wire net309;
 wire net310;
 wire net311;
 wire net312;
 wire net313;
 wire net314;
 wire net315;
 wire net316;
 wire net317;
 wire net318;
 wire net319;
 wire net320;
 wire net321;
 wire net322;
 wire net323;
 wire net324;
 wire net325;
 wire net326;
 wire net327;
 wire net328;
 wire net329;
 wire net330;
 wire net331;
 wire net332;
 wire net333;
 wire net334;
 wire net335;
 wire net336;
 wire net337;
 wire net338;
 wire net339;
 wire net340;
 wire net341;
 wire net342;
 wire net343;
 wire net344;
 wire net345;
 wire net346;
 wire net347;
 wire net348;
 wire net349;
 wire net350;
 wire net351;
 wire net352;
 wire net354;
 wire net355;
 wire net356;
 wire net357;
 wire net358;
 wire net359;
 wire net360;
 wire net361;
 wire net362;
 wire net363;
 wire net364;
 wire net365;
 wire net366;
 wire net367;
 wire net368;
 wire net369;
 wire net370;
 wire net371;
 wire net372;
 wire net373;
 wire net374;
 wire net375;
 wire net376;
 wire net377;
 wire net378;
 wire net379;
 wire net380;
 wire net381;
 wire net382;
 wire net383;
 wire net384;
 wire net385;
 wire net386;
 wire net387;
 wire net388;
 wire net389;
 wire net390;
 wire net391;
 wire net392;
 wire net393;
 wire net394;
 wire net395;
 wire net396;
 wire net397;
 wire net398;
 wire net399;
 wire net400;
 wire net401;
 wire net402;
 wire net403;
 wire net404;
 wire net405;
 wire net406;
 wire net407;
 wire net408;
 wire net409;
 wire net410;
 wire net411;
 wire net412;
 wire net413;
 wire net414;
 wire net415;
 wire net416;
 wire net417;
 wire net418;
 wire net419;
 wire net420;
 wire net421;
 wire net422;
 wire net423;
 wire net424;
 wire net425;
 wire net426;
 wire net427;
 wire net428;
 wire net429;
 wire net430;
 wire net431;
 wire net432;
 wire net433;
 wire net434;
 wire net435;
 wire net436;
 wire net437;
 wire net438;
 wire net439;
 wire net440;
 wire net441;
 wire net442;
 wire net443;
 wire net444;
 wire net445;
 wire net446;
 wire net447;
 wire net448;
 wire net449;
 wire net450;
 wire net451;
 wire net452;
 wire net453;
 wire net454;
 wire net455;
 wire net456;
 wire net457;
 wire net458;
 wire net459;
 wire net460;
 wire net461;
 wire net462;
 wire net463;
 wire net464;
 wire net465;
 wire net466;
 wire net467;
 wire net468;
 wire net469;
 wire net470;
 wire net471;
 wire net472;
 wire net473;
 wire net474;
 wire net475;
 wire net476;
 wire net477;
 wire net478;
 wire net479;
 wire net480;
 wire net481;
 wire net482;
 wire net483;
 wire net484;
 wire net485;
 wire net486;
 wire net487;
 wire net488;
 wire net489;
 wire net490;
 wire net491;
 wire net492;
 wire net493;
 wire net494;
 wire net495;
 wire net496;
 wire net497;
 wire net498;
 wire net499;
 wire net500;
 wire net501;
 wire net502;
 wire net503;
 wire net504;
 wire net505;
 wire net506;
 wire net507;
 wire net508;
 wire net509;
 wire net510;
 wire net511;
 wire net512;
 wire net513;
 wire net514;
 wire net515;
 wire net516;
 wire net517;
 wire net518;
 wire net519;
 wire net520;
 wire net521;
 wire net522;
 wire net523;
 wire net524;
 wire net525;
 wire net526;
 wire net527;
 wire net528;
 wire net529;
 wire net530;
 wire net531;
 wire net532;
 wire net533;
 wire net534;
 wire net535;
 wire net536;
 wire net537;
 wire net538;
 wire net539;
 wire net540;
 wire net541;
 wire net542;
 wire net543;
 wire net544;
 wire net545;
 wire net546;
 wire net547;
 wire net548;
 wire net549;
 wire net550;
 wire net551;
 wire net552;
 wire net553;
 wire net554;
 wire net555;
 wire clknet_leaf_1_clk;
 wire clknet_leaf_2_clk;
 wire clknet_leaf_3_clk;
 wire clknet_leaf_4_clk;
 wire clknet_leaf_5_clk;
 wire clknet_leaf_6_clk;
 wire clknet_leaf_7_clk;
 wire clknet_leaf_8_clk;
 wire clknet_leaf_9_clk;
 wire clknet_leaf_10_clk;
 wire clknet_leaf_11_clk;
 wire clknet_leaf_12_clk;
 wire clknet_leaf_13_clk;
 wire clknet_leaf_14_clk;
 wire clknet_leaf_15_clk;
 wire clknet_leaf_16_clk;
 wire clknet_leaf_17_clk;
 wire clknet_leaf_18_clk;
 wire clknet_leaf_19_clk;
 wire clknet_leaf_20_clk;
 wire clknet_leaf_21_clk;
 wire clknet_leaf_22_clk;
 wire clknet_leaf_23_clk;
 wire clknet_leaf_24_clk;
 wire clknet_leaf_25_clk;
 wire clknet_0_clk;
 wire clknet_2_0__leaf_clk;
 wire clknet_2_1__leaf_clk;
 wire clknet_2_2__leaf_clk;
 wire clknet_2_3__leaf_clk;

 sg13g2_buf_1 _07673_ (.A(\step[2] ),
    .X(_03903_));
 sg13g2_and2_1 _07674_ (.A(\step[1] ),
    .B(\step[0] ),
    .X(_03914_));
 sg13g2_buf_2 _07675_ (.A(_03914_),
    .X(_03924_));
 sg13g2_and3_1 _07676_ (.X(_03935_),
    .A(_03903_),
    .B(\step[3] ),
    .C(_03924_));
 sg13g2_buf_2 _07677_ (.A(_03935_),
    .X(_03945_));
 sg13g2_buf_1 _07678_ (.A(\i_vga.timing_hor.counter[1] ),
    .X(_03954_));
 sg13g2_buf_2 _07679_ (.A(\i_vga.timing_hor.counter[0] ),
    .X(_03964_));
 sg13g2_buf_1 _07680_ (.A(\i_vga.timing_hor.counter[2] ),
    .X(_03974_));
 sg13g2_nand3_1 _07681_ (.B(_03964_),
    .C(_03974_),
    .A(_03954_),
    .Y(_03983_));
 sg13g2_buf_1 _07682_ (.A(_03983_),
    .X(_03992_));
 sg13g2_buf_1 _07683_ (.A(\i_vga.timing_hor.counter[3] ),
    .X(_03998_));
 sg13g2_nand2_1 _07684_ (.Y(_04007_),
    .A(_03998_),
    .B(_03924_));
 sg13g2_nor2_1 _07685_ (.A(_03992_),
    .B(_04007_),
    .Y(_04014_));
 sg13g2_buf_1 _07686_ (.A(\i_vga.timing_hor.counter[5] ),
    .X(_04021_));
 sg13g2_buf_1 _07687_ (.A(\i_vga.timing_hor.counter[8] ),
    .X(_04027_));
 sg13g2_buf_1 _07688_ (.A(\i_vga.timing_hor.counter[10] ),
    .X(_04034_));
 sg13g2_buf_1 _07689_ (.A(\i_vga.timing_hor.counter[4] ),
    .X(_04041_));
 sg13g2_inv_1 _07690_ (.Y(_04050_),
    .A(_04041_));
 sg13g2_buf_1 _07691_ (.A(\i_vga.timing_hor.counter[7] ),
    .X(_04060_));
 sg13g2_buf_2 _07692_ (.A(\i_vga.timing_hor.counter[6] ),
    .X(_04071_));
 sg13g2_buf_1 _07693_ (.A(\i_vga.timing_hor.counter[9] ),
    .X(_04081_));
 sg13g2_nand4_1 _07694_ (.B(_04060_),
    .C(_04071_),
    .A(_04050_),
    .Y(_04090_),
    .D(_04081_));
 sg13g2_nor4_1 _07695_ (.A(net336),
    .B(_04027_),
    .C(_04034_),
    .D(_04090_),
    .Y(_04100_));
 sg13g2_and2_1 _07696_ (.A(_04014_),
    .B(_04100_),
    .X(_04109_));
 sg13g2_buf_1 _07697_ (.A(_04109_),
    .X(_04118_));
 sg13g2_buf_1 _07698_ (.A(\i_vga.timing_ver.counter[0] ),
    .X(_04127_));
 sg13g2_buf_1 _07699_ (.A(\i_vga.timing_ver.counter[1] ),
    .X(_04136_));
 sg13g2_inv_1 _07700_ (.Y(_04145_),
    .A(_04136_));
 sg13g2_buf_1 _07701_ (.A(\i_vga.timing_ver.counter[5] ),
    .X(_04155_));
 sg13g2_buf_1 _07702_ (.A(\i_vga.timing_ver.counter[9] ),
    .X(_04166_));
 sg13g2_buf_1 _07703_ (.A(\i_vga.timing_ver.counter[6] ),
    .X(_04177_));
 sg13g2_nand3_1 _07704_ (.B(_04177_),
    .C(\i_vga.timing_ver.counter[8] ),
    .A(\i_vga.timing_ver.counter[7] ),
    .Y(_04188_));
 sg13g2_buf_1 _07705_ (.A(_04188_),
    .X(_04199_));
 sg13g2_inv_1 _07706_ (.Y(_04210_),
    .A(_04199_));
 sg13g2_nand4_1 _07707_ (.B(_04155_),
    .C(_04166_),
    .A(\i_vga.timing_ver.counter[4] ),
    .Y(_04220_),
    .D(_04210_));
 sg13g2_buf_1 _07708_ (.A(_04220_),
    .X(_04231_));
 sg13g2_buf_1 _07709_ (.A(\i_vga.timing_ver.counter[2] ),
    .X(_04241_));
 sg13g2_nand2_1 _07710_ (.Y(_04251_),
    .A(\i_vga.timing_ver.counter[3] ),
    .B(_04241_));
 sg13g2_nor4_1 _07711_ (.A(_04127_),
    .B(_04145_),
    .C(_04231_),
    .D(_04251_),
    .Y(_04261_));
 sg13g2_and2_1 _07712_ (.A(_04118_),
    .B(_04261_),
    .X(_04270_));
 sg13g2_buf_1 _07713_ (.A(_04270_),
    .X(_04280_));
 sg13g2_nand3_1 _07714_ (.B(_04027_),
    .C(_04034_),
    .A(_04081_),
    .Y(_04289_));
 sg13g2_buf_1 _07715_ (.A(_04289_),
    .X(_04298_));
 sg13g2_nand2_1 _07716_ (.Y(_04308_),
    .A(_03964_),
    .B(_03924_));
 sg13g2_inv_1 _07717_ (.Y(_04317_),
    .A(_04060_));
 sg13g2_nor2_1 _07718_ (.A(_03954_),
    .B(_03974_),
    .Y(_04327_));
 sg13g2_nand3_1 _07719_ (.B(_04317_),
    .C(_04327_),
    .A(_04050_),
    .Y(_04338_));
 sg13g2_buf_1 _07720_ (.A(_04338_),
    .X(_04348_));
 sg13g2_inv_1 _07721_ (.Y(_04359_),
    .A(\i_vga.vblank ));
 sg13g2_nand4_1 _07722_ (.B(_03998_),
    .C(net336),
    .A(_04359_),
    .Y(_04370_),
    .D(_04071_));
 sg13g2_buf_1 _07723_ (.A(_04370_),
    .X(_04381_));
 sg13g2_nor4_1 _07724_ (.A(_04298_),
    .B(_04308_),
    .C(_04348_),
    .D(_04381_),
    .Y(_04391_));
 sg13g2_buf_1 _07725_ (.A(_04391_),
    .X(_04401_));
 sg13g2_nor2_1 _07726_ (.A(_04280_),
    .B(net131),
    .Y(_04411_));
 sg13g2_buf_1 _07727_ (.A(_04411_),
    .X(_04420_));
 sg13g2_nand2_1 _07728_ (.Y(_04430_),
    .A(_03945_),
    .B(_04420_));
 sg13g2_buf_2 _07729_ (.A(_04430_),
    .X(_04439_));
 sg13g2_buf_1 _07730_ (.A(\iter[3] ),
    .X(_04449_));
 sg13g2_inv_1 _07731_ (.Y(_04458_),
    .A(_04449_));
 sg13g2_buf_2 _07732_ (.A(\i_mandel.i_sq_y.x[0] ),
    .X(_04468_));
 sg13g2_buf_1 _07733_ (.A(\i_mandel.i_sq_y.x[-1] ),
    .X(_04477_));
 sg13g2_buf_8 _07734_ (.A(_04477_),
    .X(_04488_));
 sg13g2_buf_2 _07735_ (.A(\i_mandel.i_sq_y.x[-2] ),
    .X(_04499_));
 sg13g2_buf_8 _07736_ (.A(\i_mandel.i_sq_y.x[-3] ),
    .X(_04509_));
 sg13g2_and4_1 _07737_ (.A(_04468_),
    .B(net310),
    .C(_04499_),
    .D(_04509_),
    .X(_04520_));
 sg13g2_buf_2 _07738_ (.A(_04520_),
    .X(_04531_));
 sg13g2_buf_1 _07739_ (.A(_04499_),
    .X(_04542_));
 sg13g2_nand2_1 _07740_ (.Y(_04553_),
    .A(net310),
    .B(net309));
 sg13g2_buf_2 _07741_ (.A(_04553_),
    .X(_04563_));
 sg13g2_buf_1 _07742_ (.A(_04468_),
    .X(_04574_));
 sg13g2_buf_8 _07743_ (.A(_04509_),
    .X(_04584_));
 sg13g2_buf_1 _07744_ (.A(net307),
    .X(_04595_));
 sg13g2_nand2_1 _07745_ (.Y(_04605_),
    .A(net308),
    .B(net270));
 sg13g2_buf_2 _07746_ (.A(\i_mandel.i_sq_y.x[1] ),
    .X(_04615_));
 sg13g2_buf_1 _07747_ (.A(_04615_),
    .X(_04626_));
 sg13g2_buf_8 _07748_ (.A(\i_mandel.i_sq_y.x[-4] ),
    .X(_04635_));
 sg13g2_buf_1 _07749_ (.A(_04635_),
    .X(_04645_));
 sg13g2_nand2_1 _07750_ (.Y(_04655_),
    .A(net306),
    .B(net305));
 sg13g2_a21oi_1 _07751_ (.A1(_04563_),
    .A2(_04605_),
    .Y(_04665_),
    .B1(_04655_));
 sg13g2_or2_1 _07752_ (.X(_04675_),
    .B(_04665_),
    .A(_04531_));
 sg13g2_buf_1 _07753_ (.A(_04675_),
    .X(_04685_));
 sg13g2_buf_2 _07754_ (.A(_00039_),
    .X(_04694_));
 sg13g2_inv_1 _07755_ (.Y(_04705_),
    .A(_04694_));
 sg13g2_nand2_1 _07756_ (.Y(_04714_),
    .A(net306),
    .B(net270));
 sg13g2_buf_1 _07757_ (.A(_04714_),
    .X(_04725_));
 sg13g2_xnor2_1 _07758_ (.Y(_04736_),
    .A(_04705_),
    .B(_04725_));
 sg13g2_buf_1 _07759_ (.A(net309),
    .X(_04746_));
 sg13g2_nand2_1 _07760_ (.Y(_04757_),
    .A(net308),
    .B(net269));
 sg13g2_buf_2 _07761_ (.A(_04757_),
    .X(_04768_));
 sg13g2_xnor2_1 _07762_ (.Y(_04779_),
    .A(_04736_),
    .B(_04768_));
 sg13g2_buf_1 _07763_ (.A(net305),
    .X(_04790_));
 sg13g2_buf_1 _07764_ (.A(net268),
    .X(_04801_));
 sg13g2_buf_8 _07765_ (.A(\i_mandel.i_sq_y.x[2] ),
    .X(_04812_));
 sg13g2_inv_1 _07766_ (.Y(_04823_),
    .A(_04812_));
 sg13g2_buf_1 _07767_ (.A(_04823_),
    .X(_04834_));
 sg13g2_nor2_1 _07768_ (.A(net217),
    .B(net267),
    .Y(_04845_));
 sg13g2_a21oi_1 _07769_ (.A1(_04685_),
    .A2(_04779_),
    .Y(_04856_),
    .B1(_04845_));
 sg13g2_nor2_1 _07770_ (.A(_04685_),
    .B(_04779_),
    .Y(_04866_));
 sg13g2_nor2_1 _07771_ (.A(_04856_),
    .B(_04866_),
    .Y(_04877_));
 sg13g2_buf_8 _07772_ (.A(\i_mandel.i_sq_y.x[-6] ),
    .X(_04887_));
 sg13g2_buf_1 _07773_ (.A(net333),
    .X(_04897_));
 sg13g2_buf_1 _07774_ (.A(net304),
    .X(_04907_));
 sg13g2_buf_1 _07775_ (.A(\i_mandel.i_sq_y.x[-7] ),
    .X(_04918_));
 sg13g2_buf_1 _07776_ (.A(_04918_),
    .X(_04928_));
 sg13g2_nand2_1 _07777_ (.Y(_04939_),
    .A(net266),
    .B(net303));
 sg13g2_buf_2 _07778_ (.A(_04939_),
    .X(_04949_));
 sg13g2_buf_1 _07779_ (.A(net266),
    .X(_04959_));
 sg13g2_buf_1 _07780_ (.A(net216),
    .X(_04968_));
 sg13g2_buf_1 _07781_ (.A(net303),
    .X(_04978_));
 sg13g2_buf_1 _07782_ (.A(net265),
    .X(_04988_));
 sg13g2_buf_8 _07783_ (.A(\i_mandel.i_sq_y.x[-5] ),
    .X(_04998_));
 sg13g2_buf_1 _07784_ (.A(_04998_),
    .X(_05008_));
 sg13g2_buf_1 _07785_ (.A(net302),
    .X(_05017_));
 sg13g2_buf_1 _07786_ (.A(net264),
    .X(_05027_));
 sg13g2_o21ai_1 _07787_ (.B1(net214),
    .Y(_05038_),
    .A1(_04968_),
    .A2(net215));
 sg13g2_a21oi_1 _07788_ (.A1(_04949_),
    .A2(_05038_),
    .Y(_05049_),
    .B1(_04834_));
 sg13g2_buf_1 _07789_ (.A(_05049_),
    .X(_05060_));
 sg13g2_buf_1 _07790_ (.A(net334),
    .X(_05070_));
 sg13g2_buf_1 _07791_ (.A(net301),
    .X(_05080_));
 sg13g2_nand2_1 _07792_ (.Y(_05090_),
    .A(_04790_),
    .B(net263));
 sg13g2_xor2_1 _07793_ (.B(_05090_),
    .A(_04725_),
    .X(_05100_));
 sg13g2_xnor2_1 _07794_ (.Y(_05110_),
    .A(_05100_),
    .B(_04768_));
 sg13g2_a21oi_1 _07795_ (.A1(net95),
    .A2(_04685_),
    .Y(_05120_),
    .B1(_05110_));
 sg13g2_nor2_1 _07796_ (.A(net95),
    .B(_04685_),
    .Y(_05130_));
 sg13g2_nor2_1 _07797_ (.A(_05120_),
    .B(_05130_),
    .Y(_05140_));
 sg13g2_nand2_1 _07798_ (.Y(_05150_),
    .A(_04877_),
    .B(_05140_));
 sg13g2_xnor2_1 _07799_ (.Y(_05159_),
    .A(_04694_),
    .B(_04768_));
 sg13g2_buf_1 _07800_ (.A(net310),
    .X(_05169_));
 sg13g2_buf_1 _07801_ (.A(net262),
    .X(_05179_));
 sg13g2_nand3_1 _07802_ (.B(net213),
    .C(net269),
    .A(net308),
    .Y(_05189_));
 sg13g2_o21ai_1 _07803_ (.B1(_05189_),
    .Y(_05200_),
    .A1(_04725_),
    .A2(_05159_));
 sg13g2_buf_1 _07804_ (.A(_05200_),
    .X(_05211_));
 sg13g2_nand2_1 _07805_ (.Y(_05222_),
    .A(net306),
    .B(_04746_));
 sg13g2_buf_1 _07806_ (.A(net270),
    .X(_05233_));
 sg13g2_nor2_1 _07807_ (.A(net212),
    .B(net267),
    .Y(_05244_));
 sg13g2_xnor2_1 _07808_ (.Y(_05255_),
    .A(_05222_),
    .B(_05244_));
 sg13g2_xnor2_1 _07809_ (.Y(_05266_),
    .A(_05211_),
    .B(_05255_));
 sg13g2_nor2_1 _07810_ (.A(_04877_),
    .B(_05140_),
    .Y(_05277_));
 sg13g2_a21oi_1 _07811_ (.A1(_05150_),
    .A2(_05266_),
    .Y(_05288_),
    .B1(_05277_));
 sg13g2_buf_1 _07812_ (.A(_00035_),
    .X(_05299_));
 sg13g2_buf_1 _07813_ (.A(_05299_),
    .X(_05310_));
 sg13g2_and4_1 _07814_ (.A(_04509_),
    .B(net335),
    .C(_04998_),
    .D(net333),
    .X(_05321_));
 sg13g2_buf_1 _07815_ (.A(_05321_),
    .X(_05332_));
 sg13g2_buf_2 _07816_ (.A(_00040_),
    .X(_05343_));
 sg13g2_inv_1 _07817_ (.Y(_05354_),
    .A(_05343_));
 sg13g2_a21oi_1 _07818_ (.A1(net301),
    .A2(net261),
    .Y(_05365_),
    .B1(_05354_));
 sg13g2_buf_2 _07819_ (.A(_05365_),
    .X(_05376_));
 sg13g2_nand4_1 _07820_ (.B(net335),
    .C(_04998_),
    .A(_04509_),
    .Y(_05387_),
    .D(net333));
 sg13g2_buf_2 _07821_ (.A(_05387_),
    .X(_05398_));
 sg13g2_nor3_1 _07822_ (.A(_04823_),
    .B(_05343_),
    .C(_05398_),
    .Y(_05409_));
 sg13g2_buf_2 _07823_ (.A(_05409_),
    .X(_05420_));
 sg13g2_nor3_2 _07824_ (.A(net300),
    .B(_05376_),
    .C(_05420_),
    .Y(_05431_));
 sg13g2_buf_2 _07825_ (.A(_00041_),
    .X(_05442_));
 sg13g2_buf_1 _07826_ (.A(\i_mandel.i_sq_y.x[-12] ),
    .X(_05453_));
 sg13g2_nor2b_1 _07827_ (.A(_05442_),
    .B_N(net332),
    .Y(_05464_));
 sg13g2_and2_1 _07828_ (.A(net332),
    .B(_05442_),
    .X(_05475_));
 sg13g2_and4_1 _07829_ (.A(net335),
    .B(_04998_),
    .C(_04887_),
    .D(\i_mandel.i_sq_y.x[2] ),
    .X(_05486_));
 sg13g2_buf_1 _07830_ (.A(_05486_),
    .X(_05497_));
 sg13g2_buf_8 _07831_ (.A(_05497_),
    .X(_05507_));
 sg13g2_mux2_1 _07832_ (.A0(_05464_),
    .A1(_05475_),
    .S(_05507_),
    .X(_05518_));
 sg13g2_buf_2 _07833_ (.A(_05518_),
    .X(_05529_));
 sg13g2_buf_2 _07834_ (.A(\i_mandel.i_sq_y.x[-11] ),
    .X(_05540_));
 sg13g2_inv_1 _07835_ (.Y(_05551_),
    .A(_05540_));
 sg13g2_buf_1 _07836_ (.A(_05551_),
    .X(_05562_));
 sg13g2_buf_2 _07837_ (.A(_00042_),
    .X(_05573_));
 sg13g2_and3_1 _07838_ (.X(_05584_),
    .A(_04998_),
    .B(net333),
    .C(net334));
 sg13g2_xor2_1 _07839_ (.B(_05584_),
    .A(_05573_),
    .X(_05595_));
 sg13g2_buf_1 _07840_ (.A(_05595_),
    .X(_05606_));
 sg13g2_nor2_1 _07841_ (.A(net260),
    .B(_05606_),
    .Y(_05617_));
 sg13g2_xnor2_1 _07842_ (.Y(_05628_),
    .A(_05529_),
    .B(_05617_));
 sg13g2_xnor2_1 _07843_ (.Y(_05639_),
    .A(_05431_),
    .B(_05628_));
 sg13g2_buf_1 _07844_ (.A(\i_mandel.i_sq_y.x[-10] ),
    .X(_05650_));
 sg13g2_xnor2_1 _07845_ (.Y(_05661_),
    .A(_04998_),
    .B(net333));
 sg13g2_nor2b_1 _07846_ (.A(net334),
    .B_N(_00043_),
    .Y(_05672_));
 sg13g2_a21oi_1 _07847_ (.A1(net334),
    .A2(_05661_),
    .Y(_05683_),
    .B1(_05672_));
 sg13g2_buf_1 _07848_ (.A(_05683_),
    .X(_05694_));
 sg13g2_nand2_1 _07849_ (.Y(_05705_),
    .A(net331),
    .B(net210));
 sg13g2_or2_1 _07850_ (.X(_05716_),
    .B(_05442_),
    .A(_05299_));
 sg13g2_nand2b_1 _07851_ (.Y(_05727_),
    .B(_05442_),
    .A_N(_05299_));
 sg13g2_mux2_1 _07852_ (.A0(_05716_),
    .A1(_05727_),
    .S(_05507_),
    .X(_05738_));
 sg13g2_xnor2_1 _07853_ (.Y(_05749_),
    .A(_05573_),
    .B(_05584_));
 sg13g2_a22oi_1 _07854_ (.Y(_05760_),
    .B1(_05694_),
    .B2(_05540_),
    .A2(_05749_),
    .A1(net332));
 sg13g2_buf_1 _07855_ (.A(net332),
    .X(_05771_));
 sg13g2_buf_1 _07856_ (.A(_05540_),
    .X(_05782_));
 sg13g2_buf_8 _07857_ (.A(_05749_),
    .X(_05793_));
 sg13g2_nand4_1 _07858_ (.B(net298),
    .C(net209),
    .A(net299),
    .Y(_05804_),
    .D(net210));
 sg13g2_o21ai_1 _07859_ (.B1(_05804_),
    .Y(_05815_),
    .A1(_05738_),
    .A2(_05760_));
 sg13g2_nor2b_1 _07860_ (.A(_05705_),
    .B_N(_05815_),
    .Y(_05826_));
 sg13g2_nand2b_1 _07861_ (.Y(_05837_),
    .B(_05705_),
    .A_N(_05815_));
 sg13g2_o21ai_1 _07862_ (.B1(_05837_),
    .Y(_05848_),
    .A1(_05639_),
    .A2(_05826_));
 sg13g2_xnor2_1 _07863_ (.Y(_05859_),
    .A(_05442_),
    .B(_05497_));
 sg13g2_nor2b_1 _07864_ (.A(_05343_),
    .B_N(net332),
    .Y(_05870_));
 sg13g2_o21ai_1 _07865_ (.B1(_05870_),
    .Y(_05881_),
    .A1(_04823_),
    .A2(_05398_));
 sg13g2_nand4_1 _07866_ (.B(net334),
    .C(_05343_),
    .A(net332),
    .Y(_05892_),
    .D(net261));
 sg13g2_buf_1 _07867_ (.A(_05892_),
    .X(_05903_));
 sg13g2_and4_1 _07868_ (.A(net298),
    .B(_05859_),
    .C(_05881_),
    .D(_05903_),
    .X(_05914_));
 sg13g2_buf_8 _07869_ (.A(_05859_),
    .X(_05925_));
 sg13g2_a22oi_1 _07870_ (.Y(_05936_),
    .B1(_05881_),
    .B2(_05903_),
    .A2(net161),
    .A1(net298));
 sg13g2_and2_1 _07871_ (.A(_04499_),
    .B(_04509_),
    .X(_05947_));
 sg13g2_buf_1 _07872_ (.A(_05947_),
    .X(_05958_));
 sg13g2_a21oi_1 _07873_ (.A1(net211),
    .A2(_05958_),
    .Y(_05969_),
    .B1(_04705_));
 sg13g2_buf_2 _07874_ (.A(_05969_),
    .X(_05980_));
 sg13g2_nand4_1 _07875_ (.B(_04998_),
    .C(_04887_),
    .A(net335),
    .Y(_05991_),
    .D(_04812_));
 sg13g2_buf_2 _07876_ (.A(_05991_),
    .X(_06002_));
 sg13g2_nand3b_1 _07877_ (.B(_04509_),
    .C(_04499_),
    .Y(_06013_),
    .A_N(_04694_));
 sg13g2_buf_1 _07878_ (.A(_06013_),
    .X(_06024_));
 sg13g2_nor2_2 _07879_ (.A(_06002_),
    .B(_06024_),
    .Y(_06035_));
 sg13g2_nor3_2 _07880_ (.A(net300),
    .B(_05980_),
    .C(_06035_),
    .Y(_06046_));
 sg13g2_o21ai_1 _07881_ (.B1(_06046_),
    .Y(_06057_),
    .A1(_05914_),
    .A2(_05936_));
 sg13g2_buf_1 _07882_ (.A(_06057_),
    .X(_06068_));
 sg13g2_or3_1 _07883_ (.A(_06046_),
    .B(_05914_),
    .C(_05936_),
    .X(_06079_));
 sg13g2_buf_1 _07884_ (.A(_06079_),
    .X(_06090_));
 sg13g2_nand2_2 _07885_ (.Y(_06101_),
    .A(_06068_),
    .B(_06090_));
 sg13g2_nor2_1 _07886_ (.A(net298),
    .B(_05529_),
    .Y(_06112_));
 sg13g2_nor2_1 _07887_ (.A(_05310_),
    .B(_05354_),
    .Y(_06123_));
 sg13g2_nor2_1 _07888_ (.A(_04823_),
    .B(_05398_),
    .Y(_06134_));
 sg13g2_or2_1 _07889_ (.X(_06145_),
    .B(_05343_),
    .A(_05299_));
 sg13g2_a21oi_1 _07890_ (.A1(net301),
    .A2(net261),
    .Y(_06156_),
    .B1(_06145_));
 sg13g2_a221oi_1 _07891_ (.B2(_06134_),
    .C1(_06156_),
    .B1(_06123_),
    .A1(net298),
    .Y(_06167_),
    .A2(_05529_));
 sg13g2_inv_1 _07892_ (.Y(_06178_),
    .A(net331));
 sg13g2_buf_1 _07893_ (.A(_05606_),
    .X(_06189_));
 sg13g2_nor2_1 _07894_ (.A(_06178_),
    .B(net160),
    .Y(_06200_));
 sg13g2_o21ai_1 _07895_ (.B1(_06200_),
    .Y(_06211_),
    .A1(_06112_),
    .A2(_06167_));
 sg13g2_nand2_1 _07896_ (.Y(_06222_),
    .A(_05540_),
    .B(_06178_));
 sg13g2_buf_2 _07897_ (.A(_06222_),
    .X(_06233_));
 sg13g2_nor2_1 _07898_ (.A(_06233_),
    .B(net160),
    .Y(_06244_));
 sg13g2_buf_8 _07899_ (.A(_06002_),
    .X(_06255_));
 sg13g2_nand2_1 _07900_ (.Y(_06266_),
    .A(_06255_),
    .B(_05464_));
 sg13g2_nand2_1 _07901_ (.Y(_06277_),
    .A(net211),
    .B(_05475_));
 sg13g2_a22oi_1 _07902_ (.Y(_06288_),
    .B1(net209),
    .B2(net331),
    .A2(_06277_),
    .A1(_06266_));
 sg13g2_o21ai_1 _07903_ (.B1(_05431_),
    .Y(_06299_),
    .A1(_06244_),
    .A2(_06288_));
 sg13g2_nand2_1 _07904_ (.Y(_06310_),
    .A(_05529_),
    .B(_06244_));
 sg13g2_nand3_1 _07905_ (.B(_06299_),
    .C(_06310_),
    .A(_06211_),
    .Y(_06321_));
 sg13g2_xnor2_1 _07906_ (.Y(_06332_),
    .A(_06101_),
    .B(_06321_));
 sg13g2_nor2b_1 _07907_ (.A(_05848_),
    .B_N(_06332_),
    .Y(_06343_));
 sg13g2_inv_1 _07908_ (.Y(_06354_),
    .A(_06343_));
 sg13g2_nor2b_1 _07909_ (.A(_06332_),
    .B_N(_05848_),
    .Y(_06365_));
 sg13g2_xnor2_1 _07910_ (.Y(_06376_),
    .A(_05705_),
    .B(_05815_));
 sg13g2_xor2_1 _07911_ (.B(_06376_),
    .A(_05639_),
    .X(_06387_));
 sg13g2_buf_8 _07912_ (.A(_06387_),
    .X(_06398_));
 sg13g2_xor2_1 _07913_ (.B(net334),
    .A(net333),
    .X(_06409_));
 sg13g2_buf_2 _07914_ (.A(_06409_),
    .X(_06420_));
 sg13g2_nand2_1 _07915_ (.Y(_06431_),
    .A(net331),
    .B(_06420_));
 sg13g2_nand2_1 _07916_ (.Y(_06442_),
    .A(net332),
    .B(_05749_));
 sg13g2_a21o_1 _07917_ (.A2(_05683_),
    .A1(_05540_),
    .B1(_05738_),
    .X(_06453_));
 sg13g2_nand3_1 _07918_ (.B(_05683_),
    .C(_05738_),
    .A(_05540_),
    .Y(_06464_));
 sg13g2_nand3_1 _07919_ (.B(_06453_),
    .C(_06464_),
    .A(_06442_),
    .Y(_06475_));
 sg13g2_a21o_1 _07920_ (.A2(_06464_),
    .A1(_06453_),
    .B1(_06442_),
    .X(_06486_));
 sg13g2_buf_1 _07921_ (.A(_06486_),
    .X(_06497_));
 sg13g2_and2_1 _07922_ (.A(net332),
    .B(_05683_),
    .X(_06508_));
 sg13g2_buf_1 _07923_ (.A(_06508_),
    .X(_06519_));
 sg13g2_nand2_1 _07924_ (.Y(_06530_),
    .A(_05540_),
    .B(_06420_));
 sg13g2_o21ai_1 _07925_ (.B1(_06530_),
    .Y(_06541_),
    .A1(net300),
    .A2(net160));
 sg13g2_buf_1 _07926_ (.A(net300),
    .X(_06552_));
 sg13g2_nor3_1 _07927_ (.A(net259),
    .B(_05573_),
    .C(_06530_),
    .Y(_06563_));
 sg13g2_a21o_1 _07928_ (.A2(_06541_),
    .A1(_06519_),
    .B1(_06563_),
    .X(_06574_));
 sg13g2_nand3_1 _07929_ (.B(_06497_),
    .C(_06574_),
    .A(_06475_),
    .Y(_06585_));
 sg13g2_a21oi_1 _07930_ (.A1(_06475_),
    .A2(_06497_),
    .Y(_06596_),
    .B1(_06574_));
 sg13g2_a21oi_1 _07931_ (.A1(_06431_),
    .A2(_06585_),
    .Y(_06607_),
    .B1(_06596_));
 sg13g2_buf_2 _07932_ (.A(_06607_),
    .X(_06618_));
 sg13g2_nor2_2 _07933_ (.A(_06398_),
    .B(_06618_),
    .Y(_06629_));
 sg13g2_o21ai_1 _07934_ (.B1(net260),
    .Y(_06640_),
    .A1(net300),
    .A2(_05606_));
 sg13g2_buf_1 _07935_ (.A(net298),
    .X(_06651_));
 sg13g2_nor2_2 _07936_ (.A(net300),
    .B(_05606_),
    .Y(_06662_));
 sg13g2_nand2_1 _07937_ (.Y(_06673_),
    .A(net258),
    .B(_06662_));
 sg13g2_buf_1 _07938_ (.A(\i_mandel.i_sq_y.x[-13] ),
    .X(_06684_));
 sg13g2_nand3_1 _07939_ (.B(_06420_),
    .C(_06519_),
    .A(_06684_),
    .Y(_06695_));
 sg13g2_a21oi_1 _07940_ (.A1(_06640_),
    .A2(_06673_),
    .Y(_06706_),
    .B1(_06695_));
 sg13g2_and2_1 _07941_ (.A(_06475_),
    .B(_06497_),
    .X(_06717_));
 sg13g2_inv_1 _07942_ (.Y(_06728_),
    .A(_06431_));
 sg13g2_nor3_1 _07943_ (.A(net300),
    .B(net260),
    .C(net160),
    .Y(_06738_));
 sg13g2_o21ai_1 _07944_ (.B1(_06640_),
    .Y(_06749_),
    .A1(_06519_),
    .A2(_06738_));
 sg13g2_or2_1 _07945_ (.X(_06760_),
    .B(_06662_),
    .A(_06519_));
 sg13g2_xnor2_1 _07946_ (.Y(_06771_),
    .A(net333),
    .B(net301));
 sg13g2_nor2_1 _07947_ (.A(_06233_),
    .B(_06771_),
    .Y(_06782_));
 sg13g2_and3_1 _07948_ (.X(_06793_),
    .A(_06431_),
    .B(_06519_),
    .C(_06662_));
 sg13g2_a221oi_1 _07949_ (.B2(_06782_),
    .C1(_06793_),
    .B1(_06760_),
    .A1(_06728_),
    .Y(_06804_),
    .A2(_06749_));
 sg13g2_xnor2_1 _07950_ (.Y(_06815_),
    .A(_06717_),
    .B(_06804_));
 sg13g2_buf_1 _07951_ (.A(_06815_),
    .X(_06826_));
 sg13g2_a22oi_1 _07952_ (.Y(_06836_),
    .B1(_06706_),
    .B2(net69),
    .A2(_06618_),
    .A1(_06398_));
 sg13g2_buf_1 _07953_ (.A(_06836_),
    .X(_06847_));
 sg13g2_or3_1 _07954_ (.A(_06365_),
    .B(_06629_),
    .C(_06847_),
    .X(_06858_));
 sg13g2_buf_1 _07955_ (.A(_06858_),
    .X(_06869_));
 sg13g2_and3_1 _07956_ (.X(_06880_),
    .A(_04477_),
    .B(_04499_),
    .C(net334));
 sg13g2_buf_1 _07957_ (.A(_06880_),
    .X(_06891_));
 sg13g2_buf_2 _07958_ (.A(_00038_),
    .X(_06902_));
 sg13g2_inv_1 _07959_ (.Y(_06912_),
    .A(_06902_));
 sg13g2_a21oi_1 _07960_ (.A1(net261),
    .A2(_06891_),
    .Y(_06923_),
    .B1(_06912_));
 sg13g2_nand3_1 _07961_ (.B(_04499_),
    .C(net334),
    .A(_04477_),
    .Y(_06934_));
 sg13g2_buf_1 _07962_ (.A(_06934_),
    .X(_06945_));
 sg13g2_nor3_1 _07963_ (.A(_06902_),
    .B(_05398_),
    .C(_06945_),
    .Y(_06956_));
 sg13g2_nor3_1 _07964_ (.A(_05310_),
    .B(_06923_),
    .C(_06956_),
    .Y(_06967_));
 sg13g2_buf_2 _07965_ (.A(_06967_),
    .X(_06978_));
 sg13g2_o21ai_1 _07966_ (.B1(net299),
    .Y(_06989_),
    .A1(net208),
    .A2(_06024_));
 sg13g2_nand2_1 _07967_ (.Y(_06999_),
    .A(_04499_),
    .B(net307));
 sg13g2_o21ai_1 _07968_ (.B1(_04694_),
    .Y(_07010_),
    .A1(net208),
    .A2(_06999_));
 sg13g2_buf_2 _07969_ (.A(_07010_),
    .X(_07021_));
 sg13g2_nand2b_1 _07970_ (.Y(_07032_),
    .B(_07021_),
    .A_N(_06989_));
 sg13g2_or3_1 _07971_ (.A(net260),
    .B(_05376_),
    .C(_05420_),
    .X(_07043_));
 sg13g2_xnor2_1 _07972_ (.Y(_07054_),
    .A(_07032_),
    .B(_07043_));
 sg13g2_xnor2_1 _07973_ (.Y(_07065_),
    .A(_06978_),
    .B(_07054_));
 sg13g2_buf_1 _07974_ (.A(_07065_),
    .X(_07075_));
 sg13g2_nand2_1 _07975_ (.Y(_07086_),
    .A(net258),
    .B(net161));
 sg13g2_and2_1 _07976_ (.A(_05881_),
    .B(_05903_),
    .X(_07097_));
 sg13g2_nand2_1 _07977_ (.Y(_07108_),
    .A(_07086_),
    .B(_07097_));
 sg13g2_nor2_1 _07978_ (.A(_07086_),
    .B(_07097_),
    .Y(_07119_));
 sg13g2_a21o_1 _07979_ (.A2(_06046_),
    .A1(_07108_),
    .B1(_07119_),
    .X(_07128_));
 sg13g2_buf_2 _07980_ (.A(_07128_),
    .X(_07137_));
 sg13g2_xnor2_1 _07981_ (.Y(_07146_),
    .A(net80),
    .B(_07137_));
 sg13g2_nor2_1 _07982_ (.A(_06112_),
    .B(_06167_),
    .Y(_07154_));
 sg13g2_nand2_1 _07983_ (.Y(_07163_),
    .A(_07154_),
    .B(_05793_));
 sg13g2_and2_1 _07984_ (.A(_05529_),
    .B(_05431_),
    .X(_07171_));
 sg13g2_nor2_1 _07985_ (.A(_05793_),
    .B(_07171_),
    .Y(_07178_));
 sg13g2_a21o_1 _07986_ (.A2(_07163_),
    .A1(_06101_),
    .B1(_07178_),
    .X(_07187_));
 sg13g2_buf_1 _07987_ (.A(_07187_),
    .X(_07196_));
 sg13g2_nand3_1 _07988_ (.B(_06090_),
    .C(_07154_),
    .A(_06068_),
    .Y(_07203_));
 sg13g2_buf_1 _07989_ (.A(_06178_),
    .X(_07213_));
 sg13g2_a221oi_1 _07990_ (.B2(_07213_),
    .C1(_07178_),
    .B1(_07203_),
    .A1(_06101_),
    .Y(_07221_),
    .A2(_07163_));
 sg13g2_buf_2 _07991_ (.A(_07221_),
    .X(_07230_));
 sg13g2_nand2_1 _07992_ (.Y(_07239_),
    .A(net331),
    .B(net161));
 sg13g2_mux2_1 _07993_ (.A0(_07196_),
    .A1(_07230_),
    .S(_07239_),
    .X(_07248_));
 sg13g2_xor2_1 _07994_ (.B(_07248_),
    .A(_07146_),
    .X(_07256_));
 sg13g2_a21o_1 _07995_ (.A2(_06869_),
    .A1(_06354_),
    .B1(_07256_),
    .X(_07264_));
 sg13g2_buf_8 _07996_ (.A(_07264_),
    .X(_07272_));
 sg13g2_buf_8 _07997_ (.A(_07272_),
    .X(_07282_));
 sg13g2_xor2_1 _07998_ (.B(_07054_),
    .A(_06978_),
    .X(_07289_));
 sg13g2_xnor2_1 _07999_ (.Y(_07296_),
    .A(_05442_),
    .B(net208));
 sg13g2_nor2_1 _08000_ (.A(_06178_),
    .B(_07296_),
    .Y(_07301_));
 sg13g2_buf_1 _08001_ (.A(_07301_),
    .X(_07302_));
 sg13g2_and2_1 _08002_ (.A(_07302_),
    .B(_06046_),
    .X(_07303_));
 sg13g2_a22oi_1 _08003_ (.Y(_07304_),
    .B1(_07303_),
    .B2(_07108_),
    .A2(_07119_),
    .A1(_07302_));
 sg13g2_buf_1 _08004_ (.A(_07304_),
    .X(_07305_));
 sg13g2_nor2_1 _08005_ (.A(_07302_),
    .B(_07137_),
    .Y(_07306_));
 sg13g2_a21oi_2 _08006_ (.B1(_07306_),
    .Y(_07307_),
    .A2(_07305_),
    .A1(_07289_));
 sg13g2_nor2_1 _08007_ (.A(_06923_),
    .B(_06956_),
    .Y(_07308_));
 sg13g2_buf_1 _08008_ (.A(_07308_),
    .X(_07309_));
 sg13g2_nand2_1 _08009_ (.Y(_07310_),
    .A(_05771_),
    .B(net130));
 sg13g2_o21ai_1 _08010_ (.B1(_04705_),
    .Y(_07311_),
    .A1(_06255_),
    .A2(_06999_));
 sg13g2_nand2_1 _08011_ (.Y(_07312_),
    .A(_04468_),
    .B(net310));
 sg13g2_buf_2 _08012_ (.A(_07312_),
    .X(_07313_));
 sg13g2_nand4_1 _08013_ (.B(net211),
    .C(_05958_),
    .A(_04694_),
    .Y(_07314_),
    .D(_07313_));
 sg13g2_buf_1 _08014_ (.A(_00037_),
    .X(_07315_));
 sg13g2_inv_1 _08015_ (.Y(_07316_),
    .A(net330));
 sg13g2_a21oi_1 _08016_ (.A1(_07311_),
    .A2(_07314_),
    .Y(_07317_),
    .B1(_07316_));
 sg13g2_inv_1 _08017_ (.Y(_07318_),
    .A(_05299_));
 sg13g2_buf_1 _08018_ (.A(_07318_),
    .X(_07319_));
 sg13g2_nor3_1 _08019_ (.A(net256),
    .B(_05980_),
    .C(_06035_),
    .Y(_07320_));
 sg13g2_xnor2_1 _08020_ (.Y(_07321_),
    .A(net330),
    .B(_04694_));
 sg13g2_nor3_1 _08021_ (.A(net259),
    .B(_07313_),
    .C(_07321_),
    .Y(_07322_));
 sg13g2_nor3_1 _08022_ (.A(_07317_),
    .B(_07320_),
    .C(_07322_),
    .Y(_07323_));
 sg13g2_nand4_1 _08023_ (.B(net310),
    .C(_04499_),
    .A(_04468_),
    .Y(_07324_),
    .D(net307));
 sg13g2_buf_2 _08024_ (.A(_07324_),
    .X(_07325_));
 sg13g2_nor2_1 _08025_ (.A(net298),
    .B(net330),
    .Y(_07326_));
 sg13g2_o21ai_1 _08026_ (.B1(_07326_),
    .Y(_07327_),
    .A1(net208),
    .A2(_07325_));
 sg13g2_nand4_1 _08027_ (.B(net330),
    .C(net211),
    .A(net260),
    .Y(_07328_),
    .D(_04531_));
 sg13g2_nand2_1 _08028_ (.Y(_07329_),
    .A(_07327_),
    .B(_07328_));
 sg13g2_nand4_1 _08029_ (.B(net211),
    .C(_05958_),
    .A(_04705_),
    .Y(_07330_),
    .D(_07313_));
 sg13g2_a21oi_1 _08030_ (.A1(_07021_),
    .A2(_07330_),
    .Y(_07331_),
    .B1(net330));
 sg13g2_o21ai_1 _08031_ (.B1(net256),
    .Y(_07332_),
    .A1(_07329_),
    .A2(_07331_));
 sg13g2_o21ai_1 _08032_ (.B1(_07332_),
    .Y(_07333_),
    .A1(net260),
    .A2(_07323_));
 sg13g2_xor2_1 _08033_ (.B(_07333_),
    .A(_07310_),
    .X(_07334_));
 sg13g2_or2_1 _08034_ (.X(_07335_),
    .B(_05420_),
    .A(_05376_));
 sg13g2_buf_1 _08035_ (.A(_07335_),
    .X(_07336_));
 sg13g2_nor2_1 _08036_ (.A(_06178_),
    .B(_07336_),
    .Y(_07337_));
 sg13g2_nor2_1 _08037_ (.A(_05980_),
    .B(_06989_),
    .Y(_07338_));
 sg13g2_a21o_1 _08038_ (.A2(_07338_),
    .A1(net298),
    .B1(_06978_),
    .X(_07339_));
 sg13g2_o21ai_1 _08039_ (.B1(_07339_),
    .Y(_07340_),
    .A1(net258),
    .A2(_07338_));
 sg13g2_nor2_1 _08040_ (.A(_07336_),
    .B(_06233_),
    .Y(_07341_));
 sg13g2_nand2b_1 _08041_ (.Y(_07342_),
    .B(_07032_),
    .A_N(_06978_));
 sg13g2_nand2_1 _08042_ (.Y(_07343_),
    .A(_06978_),
    .B(_07338_));
 sg13g2_nor2_1 _08043_ (.A(_07343_),
    .B(_07337_),
    .Y(_07344_));
 sg13g2_a221oi_1 _08044_ (.B2(_07342_),
    .C1(_07344_),
    .B1(_07341_),
    .A1(_07337_),
    .Y(_07345_),
    .A2(_07340_));
 sg13g2_xor2_1 _08045_ (.B(_07345_),
    .A(_07334_),
    .X(_07346_));
 sg13g2_buf_2 _08046_ (.A(_07346_),
    .X(_07347_));
 sg13g2_nor2_1 _08047_ (.A(_07289_),
    .B(_07305_),
    .Y(_07348_));
 sg13g2_nand2b_1 _08048_ (.Y(_07349_),
    .B(_07348_),
    .A_N(_07196_));
 sg13g2_nand3_1 _08049_ (.B(_07347_),
    .C(_07349_),
    .A(_07307_),
    .Y(_07350_));
 sg13g2_buf_1 _08050_ (.A(_07350_),
    .X(_07351_));
 sg13g2_xnor2_1 _08051_ (.Y(_07352_),
    .A(_07334_),
    .B(_07345_));
 sg13g2_and2_1 _08052_ (.A(_06068_),
    .B(_06090_),
    .X(_07353_));
 sg13g2_buf_1 _08053_ (.A(_07353_),
    .X(_07354_));
 sg13g2_buf_1 _08054_ (.A(net331),
    .X(_07355_));
 sg13g2_o21ai_1 _08055_ (.B1(net297),
    .Y(_07356_),
    .A1(_07354_),
    .A2(_07154_));
 sg13g2_buf_1 _08056_ (.A(_06651_),
    .X(_07357_));
 sg13g2_or2_1 _08057_ (.X(_07358_),
    .B(_05431_),
    .A(_05529_));
 sg13g2_nand3_1 _08058_ (.B(_07354_),
    .C(_07358_),
    .A(net207),
    .Y(_07359_));
 sg13g2_a21o_1 _08059_ (.A2(_07359_),
    .A1(_07356_),
    .B1(_06189_),
    .X(_07360_));
 sg13g2_a221oi_1 _08060_ (.B2(_07171_),
    .C1(net80),
    .B1(_07354_),
    .A1(net297),
    .Y(_07361_),
    .A2(net161));
 sg13g2_nand3_1 _08061_ (.B(_07360_),
    .C(_07361_),
    .A(_07352_),
    .Y(_07362_));
 sg13g2_buf_1 _08062_ (.A(_07362_),
    .X(_07363_));
 sg13g2_nand2_1 _08063_ (.Y(_07364_),
    .A(net80),
    .B(_07302_));
 sg13g2_nand2b_1 _08064_ (.Y(_07365_),
    .B(net80),
    .A_N(_07203_));
 sg13g2_o21ai_1 _08065_ (.B1(net297),
    .Y(_07366_),
    .A1(net80),
    .A2(_05925_));
 sg13g2_a22oi_1 _08066_ (.Y(_07367_),
    .B1(_07365_),
    .B2(_07366_),
    .A2(_07196_),
    .A1(_07364_));
 sg13g2_or3_1 _08067_ (.A(_07137_),
    .B(_07347_),
    .C(_07367_),
    .X(_07368_));
 sg13g2_buf_1 _08068_ (.A(_07368_),
    .X(_07369_));
 sg13g2_nand3_1 _08069_ (.B(_07363_),
    .C(_07369_),
    .A(_07351_),
    .Y(_07370_));
 sg13g2_buf_1 _08070_ (.A(_07370_),
    .X(_07371_));
 sg13g2_nor4_1 _08071_ (.A(_07075_),
    .B(_07239_),
    .C(_07137_),
    .D(_07352_),
    .Y(_07372_));
 sg13g2_nor2_1 _08072_ (.A(_07302_),
    .B(_07146_),
    .Y(_07373_));
 sg13g2_mux2_1 _08073_ (.A0(_07348_),
    .A1(_07373_),
    .S(_07347_),
    .X(_07374_));
 sg13g2_o21ai_1 _08074_ (.B1(_07230_),
    .Y(_07375_),
    .A1(_07372_),
    .A2(_07374_));
 sg13g2_o21ai_1 _08075_ (.B1(_07375_),
    .Y(_07376_),
    .A1(net34),
    .A2(_07371_));
 sg13g2_buf_8 _08076_ (.A(_07376_),
    .X(_07377_));
 sg13g2_nand2_1 _08077_ (.Y(_07378_),
    .A(_07307_),
    .B(_07347_));
 sg13g2_nor2_1 _08078_ (.A(_06978_),
    .B(_07338_),
    .Y(_07379_));
 sg13g2_a21oi_1 _08079_ (.A1(_07043_),
    .A2(_07343_),
    .Y(_07380_),
    .B1(_07379_));
 sg13g2_nor2_1 _08080_ (.A(_07337_),
    .B(_07380_),
    .Y(_07381_));
 sg13g2_nand2_1 _08081_ (.Y(_07382_),
    .A(_07337_),
    .B(_07380_));
 sg13g2_o21ai_1 _08082_ (.B1(_07382_),
    .Y(_07383_),
    .A1(_07334_),
    .A2(_07381_));
 sg13g2_buf_2 _08083_ (.A(_07383_),
    .X(_07384_));
 sg13g2_and4_1 _08084_ (.A(_04615_),
    .B(_04468_),
    .C(net310),
    .D(net309),
    .X(_07385_));
 sg13g2_a21oi_1 _08085_ (.A1(_05332_),
    .A2(_07385_),
    .Y(_07386_),
    .B1(_00036_));
 sg13g2_buf_2 _08086_ (.A(_07386_),
    .X(_07387_));
 sg13g2_nor2b_1 _08087_ (.A(_06902_),
    .B_N(_05782_),
    .Y(_07388_));
 sg13g2_o21ai_1 _08088_ (.B1(_07388_),
    .Y(_07389_),
    .A1(_05398_),
    .A2(_06945_));
 sg13g2_nand4_1 _08089_ (.B(_06902_),
    .C(net261),
    .A(_05782_),
    .Y(_07390_),
    .D(_06891_));
 sg13g2_and4_1 _08090_ (.A(net256),
    .B(_07387_),
    .C(_07389_),
    .D(_07390_),
    .X(_07391_));
 sg13g2_a22oi_1 _08091_ (.Y(_07392_),
    .B1(_07389_),
    .B2(_07390_),
    .A2(_07387_),
    .A1(net256));
 sg13g2_o21ai_1 _08092_ (.B1(net330),
    .Y(_07393_),
    .A1(net208),
    .A2(_07325_));
 sg13g2_nand3_1 _08093_ (.B(net211),
    .C(_04531_),
    .A(_07316_),
    .Y(_07394_));
 sg13g2_and3_1 _08094_ (.X(_07395_),
    .A(_05771_),
    .B(_07393_),
    .C(_07394_));
 sg13g2_buf_1 _08095_ (.A(_07395_),
    .X(_07396_));
 sg13g2_o21ai_1 _08096_ (.B1(_07396_),
    .Y(_07397_),
    .A1(_07391_),
    .A2(_07392_));
 sg13g2_buf_1 _08097_ (.A(_07397_),
    .X(_07398_));
 sg13g2_or3_1 _08098_ (.A(_07396_),
    .B(_07391_),
    .C(_07392_),
    .X(_07399_));
 sg13g2_buf_1 _08099_ (.A(_07399_),
    .X(_07400_));
 sg13g2_nand2_1 _08100_ (.Y(_07401_),
    .A(_07398_),
    .B(_07400_));
 sg13g2_nor2b_1 _08101_ (.A(_06902_),
    .B_N(_05453_),
    .Y(_07402_));
 sg13g2_o21ai_1 _08102_ (.B1(_07402_),
    .Y(_07403_),
    .A1(_05398_),
    .A2(_06945_));
 sg13g2_nand4_1 _08103_ (.B(_06902_),
    .C(net261),
    .A(_05453_),
    .Y(_07404_),
    .D(_06891_));
 sg13g2_nor2_1 _08104_ (.A(net300),
    .B(net330),
    .Y(_07405_));
 sg13g2_o21ai_1 _08105_ (.B1(_07405_),
    .Y(_07406_),
    .A1(net208),
    .A2(_07325_));
 sg13g2_nand4_1 _08106_ (.B(_07315_),
    .C(net211),
    .A(net256),
    .Y(_07407_),
    .D(_04531_));
 sg13g2_a22oi_1 _08107_ (.Y(_07408_),
    .B1(_07406_),
    .B2(_07407_),
    .A2(_07404_),
    .A1(_07403_));
 sg13g2_buf_1 _08108_ (.A(_07408_),
    .X(_07409_));
 sg13g2_nor2_1 _08109_ (.A(_05980_),
    .B(_06035_),
    .Y(_07410_));
 sg13g2_buf_2 _08110_ (.A(_07410_),
    .X(_07411_));
 sg13g2_nand2_1 _08111_ (.Y(_07412_),
    .A(net331),
    .B(_07411_));
 sg13g2_nand4_1 _08112_ (.B(_07404_),
    .C(_07406_),
    .A(_07403_),
    .Y(_07413_),
    .D(_07407_));
 sg13g2_buf_1 _08113_ (.A(_07413_),
    .X(_07414_));
 sg13g2_a21oi_1 _08114_ (.A1(net258),
    .A2(_07414_),
    .Y(_07415_),
    .B1(_07409_));
 sg13g2_nor2_1 _08115_ (.A(_05562_),
    .B(net331),
    .Y(_07416_));
 sg13g2_and2_1 _08116_ (.A(_07416_),
    .B(_07414_),
    .X(_07417_));
 sg13g2_a21o_1 _08117_ (.A2(_07415_),
    .A1(_05650_),
    .B1(_07417_),
    .X(_07418_));
 sg13g2_a22oi_1 _08118_ (.Y(_07419_),
    .B1(_07418_),
    .B2(_07411_),
    .A2(_07412_),
    .A1(_07409_));
 sg13g2_xnor2_1 _08119_ (.Y(_07420_),
    .A(_07401_),
    .B(_07419_));
 sg13g2_xor2_1 _08120_ (.B(_07420_),
    .A(_07384_),
    .X(_07421_));
 sg13g2_xnor2_1 _08121_ (.Y(_07422_),
    .A(_07378_),
    .B(_07421_));
 sg13g2_buf_2 _08122_ (.A(_07422_),
    .X(_07423_));
 sg13g2_nand2_1 _08123_ (.Y(_07424_),
    .A(_07319_),
    .B(_07387_));
 sg13g2_nand3_1 _08124_ (.B(_07309_),
    .C(_07396_),
    .A(net258),
    .Y(_07425_));
 sg13g2_a21oi_1 _08125_ (.A1(_06651_),
    .A2(net130),
    .Y(_07426_),
    .B1(_07396_));
 sg13g2_a21o_1 _08126_ (.A2(_07425_),
    .A1(_07424_),
    .B1(_07426_),
    .X(_07427_));
 sg13g2_nand2_1 _08127_ (.Y(_07428_),
    .A(net297),
    .B(_07309_));
 sg13g2_nand3_1 _08128_ (.B(_07393_),
    .C(_07394_),
    .A(net258),
    .Y(_07429_));
 sg13g2_xnor2_1 _08129_ (.Y(_07430_),
    .A(net259),
    .B(net299));
 sg13g2_nand2_1 _08130_ (.Y(_07431_),
    .A(_07387_),
    .B(_07430_));
 sg13g2_xor2_1 _08131_ (.B(_07431_),
    .A(_07429_),
    .X(_07432_));
 sg13g2_xnor2_1 _08132_ (.Y(_07433_),
    .A(_07428_),
    .B(_07432_));
 sg13g2_xnor2_1 _08133_ (.Y(_07434_),
    .A(_07427_),
    .B(_07433_));
 sg13g2_buf_2 _08134_ (.A(_07434_),
    .X(_07435_));
 sg13g2_a221oi_1 _08135_ (.B2(_07357_),
    .C1(_07409_),
    .B1(_07414_),
    .A1(_07398_),
    .Y(_07436_),
    .A2(_07400_));
 sg13g2_a21oi_1 _08136_ (.A1(_07398_),
    .A2(_07400_),
    .Y(_07437_),
    .B1(_07411_));
 sg13g2_nand2_1 _08137_ (.Y(_07438_),
    .A(_07357_),
    .B(_07414_));
 sg13g2_nor2_1 _08138_ (.A(_07355_),
    .B(_07409_),
    .Y(_07439_));
 sg13g2_nor2_1 _08139_ (.A(_07411_),
    .B(_07409_),
    .Y(_07440_));
 sg13g2_a21o_1 _08140_ (.A2(_07439_),
    .A1(_07438_),
    .B1(_07440_),
    .X(_07441_));
 sg13g2_a21oi_1 _08141_ (.A1(_07398_),
    .A2(_07400_),
    .Y(_07442_),
    .B1(net297));
 sg13g2_nor4_2 _08142_ (.A(_07436_),
    .B(_07437_),
    .C(_07441_),
    .Y(_07443_),
    .D(_07442_));
 sg13g2_xnor2_1 _08143_ (.Y(_07444_),
    .A(_07401_),
    .B(_07441_));
 sg13g2_nand2_1 _08144_ (.Y(_07445_),
    .A(_07419_),
    .B(_07444_));
 sg13g2_mux2_1 _08145_ (.A0(_07443_),
    .A1(_07445_),
    .S(_07384_),
    .X(_07446_));
 sg13g2_buf_1 _08146_ (.A(_07446_),
    .X(_07447_));
 sg13g2_xnor2_1 _08147_ (.Y(_07448_),
    .A(_07435_),
    .B(_07447_));
 sg13g2_nor2b_1 _08148_ (.A(_07432_),
    .B_N(_07428_),
    .Y(_07449_));
 sg13g2_nand2b_1 _08149_ (.Y(_07450_),
    .B(_07432_),
    .A_N(_07428_));
 sg13g2_o21ai_1 _08150_ (.B1(_07450_),
    .Y(_07451_),
    .A1(_07449_),
    .A2(_07427_));
 sg13g2_buf_1 _08151_ (.A(_07387_),
    .X(_07452_));
 sg13g2_buf_1 _08152_ (.A(net260),
    .X(_07453_));
 sg13g2_nor2_1 _08153_ (.A(net299),
    .B(net206),
    .Y(_07454_));
 sg13g2_and3_1 _08154_ (.X(_07455_),
    .A(net259),
    .B(net129),
    .C(_07454_));
 sg13g2_inv_1 _08155_ (.Y(_07456_),
    .A(net299));
 sg13g2_and2_1 _08156_ (.A(_07393_),
    .B(_07394_),
    .X(_07457_));
 sg13g2_buf_1 _08157_ (.A(_07457_),
    .X(_07458_));
 sg13g2_nand4_1 _08158_ (.B(net255),
    .C(_07458_),
    .A(net256),
    .Y(_07459_),
    .D(_07387_));
 sg13g2_nand4_1 _08159_ (.B(net299),
    .C(_07458_),
    .A(net259),
    .Y(_07460_),
    .D(_07387_));
 sg13g2_nand2_1 _08160_ (.Y(_07461_),
    .A(net297),
    .B(_07458_));
 sg13g2_nor2_1 _08161_ (.A(net255),
    .B(net258),
    .Y(_07462_));
 sg13g2_nor2_1 _08162_ (.A(net259),
    .B(net258),
    .Y(_07463_));
 sg13g2_o21ai_1 _08163_ (.B1(net129),
    .Y(_07464_),
    .A1(_07462_),
    .A2(_07463_));
 sg13g2_nand4_1 _08164_ (.B(_07460_),
    .C(_07461_),
    .A(_07459_),
    .Y(_07465_),
    .D(_07464_));
 sg13g2_buf_1 _08165_ (.A(net256),
    .X(_07466_));
 sg13g2_nor2_1 _08166_ (.A(net255),
    .B(net206),
    .Y(_07467_));
 sg13g2_nand2_1 _08167_ (.Y(_07468_),
    .A(net255),
    .B(net260));
 sg13g2_nor2_1 _08168_ (.A(net256),
    .B(_07468_),
    .Y(_07469_));
 sg13g2_a21oi_1 _08169_ (.A1(_07466_),
    .A2(_07467_),
    .Y(_07470_),
    .B1(_07469_));
 sg13g2_nand4_1 _08170_ (.B(_07458_),
    .C(_07452_),
    .A(net297),
    .Y(_07471_),
    .D(_07470_));
 sg13g2_o21ai_1 _08171_ (.B1(_07471_),
    .Y(_07472_),
    .A1(_07455_),
    .A2(_07465_));
 sg13g2_xor2_1 _08172_ (.B(_07472_),
    .A(_07451_),
    .X(_07473_));
 sg13g2_buf_1 _08173_ (.A(_07473_),
    .X(_07474_));
 sg13g2_nand2_1 _08174_ (.Y(_07475_),
    .A(_07443_),
    .B(_07435_));
 sg13g2_xor2_1 _08175_ (.B(_07475_),
    .A(_07474_),
    .X(_07476_));
 sg13g2_inv_1 _08176_ (.Y(_07477_),
    .A(_07476_));
 sg13g2_inv_1 _08177_ (.Y(_07478_),
    .A(_07472_));
 sg13g2_buf_1 _08178_ (.A(_07355_),
    .X(_07479_));
 sg13g2_buf_1 _08179_ (.A(net299),
    .X(_07480_));
 sg13g2_nand2_1 _08180_ (.Y(_07481_),
    .A(net253),
    .B(net207));
 sg13g2_a21oi_1 _08181_ (.A1(_07481_),
    .A2(_07458_),
    .Y(_07482_),
    .B1(_06552_));
 sg13g2_buf_1 _08182_ (.A(_07458_),
    .X(_07483_));
 sg13g2_nand2b_1 _08183_ (.Y(_07484_),
    .B(_07468_),
    .A_N(net94));
 sg13g2_nand2b_1 _08184_ (.Y(_07485_),
    .B(_07484_),
    .A_N(_07482_));
 sg13g2_nand2_1 _08185_ (.Y(_07486_),
    .A(_06552_),
    .B(_07213_));
 sg13g2_o21ai_1 _08186_ (.B1(_07452_),
    .Y(_07487_),
    .A1(_07486_),
    .A2(_07468_));
 sg13g2_a21oi_1 _08187_ (.A1(net254),
    .A2(_07485_),
    .Y(_07488_),
    .B1(_07487_));
 sg13g2_a21oi_1 _08188_ (.A1(_07451_),
    .A2(_07478_),
    .Y(_07489_),
    .B1(_07488_));
 sg13g2_buf_2 _08189_ (.A(_07489_),
    .X(_07490_));
 sg13g2_nor4_1 _08190_ (.A(_07423_),
    .B(_07448_),
    .C(_07477_),
    .D(_07490_),
    .Y(_07491_));
 sg13g2_a21oi_1 _08191_ (.A1(_07377_),
    .A2(_07491_),
    .Y(_07492_),
    .B1(_07487_));
 sg13g2_buf_8 _08192_ (.A(_07492_),
    .X(_07493_));
 sg13g2_buf_2 _08193_ (.A(\i_mandel.i_sq_y.x[-9] ),
    .X(_07494_));
 sg13g2_inv_1 _08194_ (.Y(_07495_),
    .A(_07494_));
 sg13g2_buf_1 _08195_ (.A(_07495_),
    .X(_07496_));
 sg13g2_buf_1 _08196_ (.A(\i_mandel.i_sq_y.x[-8] ),
    .X(_07497_));
 sg13g2_buf_1 _08197_ (.A(net329),
    .X(_07498_));
 sg13g2_inv_1 _08198_ (.Y(_07499_),
    .A(net296));
 sg13g2_buf_1 _08199_ (.A(_07499_),
    .X(_07500_));
 sg13g2_nor3_1 _08200_ (.A(net267),
    .B(net252),
    .C(net204),
    .Y(_07501_));
 sg13g2_nand2_1 _08201_ (.Y(_07502_),
    .A(_07493_),
    .B(_07501_));
 sg13g2_buf_1 _08202_ (.A(_07502_),
    .X(_07503_));
 sg13g2_buf_1 _08203_ (.A(_07494_),
    .X(_07504_));
 sg13g2_buf_1 _08204_ (.A(_07504_),
    .X(_07505_));
 sg13g2_buf_1 _08205_ (.A(net296),
    .X(_07506_));
 sg13g2_o21ai_1 _08206_ (.B1(net263),
    .Y(_00240_),
    .A1(net251),
    .A2(net250));
 sg13g2_buf_2 _08207_ (.A(_00240_),
    .X(_00241_));
 sg13g2_inv_1 _08208_ (.Y(_00242_),
    .A(_00241_));
 sg13g2_nor2_1 _08209_ (.A(_07493_),
    .B(_00242_),
    .Y(_00243_));
 sg13g2_buf_2 _08210_ (.A(_00243_),
    .X(_00244_));
 sg13g2_buf_1 _08211_ (.A(net263),
    .X(_00245_));
 sg13g2_xnor2_1 _08212_ (.Y(_00246_),
    .A(net216),
    .B(net215));
 sg13g2_xnor2_1 _08213_ (.Y(_00247_),
    .A(net214),
    .B(_00246_));
 sg13g2_nand2_1 _08214_ (.Y(_00248_),
    .A(net203),
    .B(_00247_));
 sg13g2_buf_2 _08215_ (.A(_00248_),
    .X(_00249_));
 sg13g2_nand2_2 _08216_ (.Y(_00250_),
    .A(_00244_),
    .B(_00249_));
 sg13g2_xnor2_1 _08217_ (.Y(_00251_),
    .A(net270),
    .B(_04790_));
 sg13g2_nor2_1 _08218_ (.A(_04834_),
    .B(_00251_),
    .Y(_00252_));
 sg13g2_xnor2_1 _08219_ (.Y(_00253_),
    .A(_05222_),
    .B(_00252_));
 sg13g2_nand2_1 _08220_ (.Y(_00254_),
    .A(_04725_),
    .B(_04768_));
 sg13g2_o21ai_1 _08221_ (.B1(_05090_),
    .Y(_00255_),
    .A1(_04725_),
    .A2(_04768_));
 sg13g2_and2_1 _08222_ (.A(_00254_),
    .B(_00255_),
    .X(_00256_));
 sg13g2_buf_1 _08223_ (.A(_00256_),
    .X(_00257_));
 sg13g2_xnor2_1 _08224_ (.Y(_00258_),
    .A(_05049_),
    .B(_00257_));
 sg13g2_xnor2_1 _08225_ (.Y(_00259_),
    .A(_00253_),
    .B(_00258_));
 sg13g2_buf_1 _08226_ (.A(_00259_),
    .X(_00260_));
 sg13g2_xor2_1 _08227_ (.B(_05100_),
    .A(_05060_),
    .X(_00261_));
 sg13g2_xor2_1 _08228_ (.B(_04768_),
    .A(_04685_),
    .X(_00262_));
 sg13g2_xnor2_1 _08229_ (.Y(_00263_),
    .A(_00261_),
    .B(_00262_));
 sg13g2_nor2b_1 _08230_ (.A(_00263_),
    .B_N(net68),
    .Y(_00264_));
 sg13g2_nand2_1 _08231_ (.Y(_00265_),
    .A(_00250_),
    .B(_00264_));
 sg13g2_o21ai_1 _08232_ (.B1(_00265_),
    .Y(_00266_),
    .A1(_00250_),
    .A2(net68));
 sg13g2_buf_1 _08233_ (.A(_00249_),
    .X(_00267_));
 sg13g2_nor2_1 _08234_ (.A(_00249_),
    .B(net68),
    .Y(_00268_));
 sg13g2_xnor2_1 _08235_ (.Y(_00269_),
    .A(_05140_),
    .B(_05266_));
 sg13g2_xnor2_1 _08236_ (.Y(_00270_),
    .A(_04877_),
    .B(_00269_));
 sg13g2_a22oi_1 _08237_ (.Y(_00271_),
    .B1(_00268_),
    .B2(_00270_),
    .A2(_00264_),
    .A1(net85));
 sg13g2_or2_1 _08238_ (.X(_00272_),
    .B(_00249_),
    .A(net30));
 sg13g2_buf_1 _08239_ (.A(_00272_),
    .X(_00273_));
 sg13g2_nand2b_1 _08240_ (.Y(_00274_),
    .B(_00263_),
    .A_N(net68));
 sg13g2_nand3_1 _08241_ (.B(_00270_),
    .C(_00274_),
    .A(_00273_),
    .Y(_00275_));
 sg13g2_o21ai_1 _08242_ (.B1(_00275_),
    .Y(_00276_),
    .A1(net30),
    .A2(_00271_));
 sg13g2_a21oi_1 _08243_ (.A1(_07503_),
    .A2(_00266_),
    .Y(_00277_),
    .B1(_00276_));
 sg13g2_nor2_1 _08244_ (.A(_05288_),
    .B(_00277_),
    .Y(_00278_));
 sg13g2_a21o_1 _08245_ (.A2(net85),
    .A1(_00244_),
    .B1(net68),
    .X(_00279_));
 sg13g2_a22oi_1 _08246_ (.Y(_00280_),
    .B1(_00279_),
    .B2(net30),
    .A2(_00260_),
    .A1(net85));
 sg13g2_buf_1 _08247_ (.A(net203),
    .X(_00281_));
 sg13g2_inv_1 _08248_ (.Y(_00282_),
    .A(net309));
 sg13g2_buf_1 _08249_ (.A(_00282_),
    .X(_00283_));
 sg13g2_nor2_1 _08250_ (.A(net270),
    .B(net268),
    .Y(_00284_));
 sg13g2_nand2_1 _08251_ (.Y(_00285_),
    .A(net202),
    .B(_00284_));
 sg13g2_and2_1 _08252_ (.A(_04584_),
    .B(net305),
    .X(_00286_));
 sg13g2_buf_2 _08253_ (.A(_00286_),
    .X(_00287_));
 sg13g2_nor2_1 _08254_ (.A(net306),
    .B(_00284_),
    .Y(_00288_));
 sg13g2_buf_1 _08255_ (.A(net269),
    .X(_00289_));
 sg13g2_o21ai_1 _08256_ (.B1(net201),
    .Y(_00290_),
    .A1(_00287_),
    .A2(_00288_));
 sg13g2_and3_1 _08257_ (.X(_00291_),
    .A(net159),
    .B(_00285_),
    .C(_00290_));
 sg13g2_xnor2_1 _08258_ (.Y(_00292_),
    .A(net95),
    .B(_00291_));
 sg13g2_buf_2 _08259_ (.A(_00292_),
    .X(_00293_));
 sg13g2_nor2_1 _08260_ (.A(_00253_),
    .B(_00257_),
    .Y(_00294_));
 sg13g2_a21oi_1 _08261_ (.A1(_00253_),
    .A2(_00257_),
    .Y(_00295_),
    .B1(_05060_));
 sg13g2_nor2_1 _08262_ (.A(_00294_),
    .B(_00295_),
    .Y(_00296_));
 sg13g2_nand2_1 _08263_ (.Y(_00297_),
    .A(net202),
    .B(net203));
 sg13g2_buf_1 _08264_ (.A(net308),
    .X(_00298_));
 sg13g2_nor2b_1 _08265_ (.A(net213),
    .B_N(_00298_),
    .Y(_00299_));
 sg13g2_xnor2_1 _08266_ (.Y(_00300_),
    .A(_00297_),
    .B(_00299_));
 sg13g2_nor2_1 _08267_ (.A(_05211_),
    .B(_05244_),
    .Y(_00301_));
 sg13g2_nor2_1 _08268_ (.A(_05222_),
    .B(_00301_),
    .Y(_00302_));
 sg13g2_a21oi_1 _08269_ (.A1(_05211_),
    .A2(_05244_),
    .Y(_00303_),
    .B1(_00302_));
 sg13g2_xor2_1 _08270_ (.B(_00303_),
    .A(_00300_),
    .X(_00304_));
 sg13g2_xnor2_1 _08271_ (.Y(_00305_),
    .A(_00296_),
    .B(_00304_));
 sg13g2_xnor2_1 _08272_ (.Y(_00306_),
    .A(_00293_),
    .B(_00305_));
 sg13g2_xnor2_1 _08273_ (.Y(_00307_),
    .A(_00280_),
    .B(_00306_));
 sg13g2_nand2_1 _08274_ (.Y(_00308_),
    .A(_05288_),
    .B(_00277_));
 sg13g2_o21ai_1 _08275_ (.B1(_00308_),
    .Y(_00309_),
    .A1(_00278_),
    .A2(_00307_));
 sg13g2_nand2_1 _08276_ (.Y(_00310_),
    .A(net68),
    .B(_00293_));
 sg13g2_xor2_1 _08277_ (.B(_00291_),
    .A(net95),
    .X(_00311_));
 sg13g2_nand3_1 _08278_ (.B(_00311_),
    .C(_00305_),
    .A(_00244_),
    .Y(_00312_));
 sg13g2_o21ai_1 _08279_ (.B1(_00312_),
    .Y(_00313_),
    .A1(_00244_),
    .A2(_00310_));
 sg13g2_o21ai_1 _08280_ (.B1(_00305_),
    .Y(_00314_),
    .A1(net68),
    .A2(_00293_));
 sg13g2_inv_1 _08281_ (.Y(_00315_),
    .A(_00314_));
 sg13g2_mux2_1 _08282_ (.A0(_00293_),
    .A1(_00310_),
    .S(net30),
    .X(_00316_));
 sg13g2_nor2_1 _08283_ (.A(net85),
    .B(_00316_),
    .Y(_00317_));
 sg13g2_a221oi_1 _08284_ (.B2(_00250_),
    .C1(_00317_),
    .B1(_00315_),
    .A1(net85),
    .Y(_00318_),
    .A2(_00313_));
 sg13g2_buf_1 _08285_ (.A(_00318_),
    .X(_00319_));
 sg13g2_inv_1 _08286_ (.Y(_00320_),
    .A(net30));
 sg13g2_o21ai_1 _08287_ (.B1(_00249_),
    .Y(_00321_),
    .A1(_00244_),
    .A2(_00311_));
 sg13g2_o21ai_1 _08288_ (.B1(_00321_),
    .Y(_00322_),
    .A1(_00320_),
    .A2(_00293_));
 sg13g2_nand2_1 _08289_ (.Y(_00323_),
    .A(_00289_),
    .B(_00287_));
 sg13g2_nand3_1 _08290_ (.B(_00285_),
    .C(_00323_),
    .A(net159),
    .Y(_00324_));
 sg13g2_xnor2_1 _08291_ (.Y(_00325_),
    .A(net95),
    .B(_00324_));
 sg13g2_buf_2 _08292_ (.A(_00325_),
    .X(_00326_));
 sg13g2_nor3_1 _08293_ (.A(net306),
    .B(net202),
    .C(_00284_),
    .Y(_00327_));
 sg13g2_nand3b_1 _08294_ (.B(net95),
    .C(_00285_),
    .Y(_00328_),
    .A_N(_00327_));
 sg13g2_and2_1 _08295_ (.A(_00323_),
    .B(_00328_),
    .X(_00329_));
 sg13g2_nand2b_1 _08296_ (.Y(_00330_),
    .B(net159),
    .A_N(_00329_));
 sg13g2_buf_1 _08297_ (.A(net213),
    .X(_00331_));
 sg13g2_a21oi_1 _08298_ (.A1(_00298_),
    .A2(net202),
    .Y(_00332_),
    .B1(net267));
 sg13g2_buf_1 _08299_ (.A(net306),
    .X(_00333_));
 sg13g2_xor2_1 _08300_ (.B(net249),
    .A(net248),
    .X(_00334_));
 sg13g2_nand2_1 _08301_ (.Y(_00335_),
    .A(net213),
    .B(net203));
 sg13g2_nand2_1 _08302_ (.Y(_00336_),
    .A(_00335_),
    .B(_00334_));
 sg13g2_o21ai_1 _08303_ (.B1(_00336_),
    .Y(_00337_),
    .A1(net267),
    .A2(_00334_));
 sg13g2_o21ai_1 _08304_ (.B1(_00337_),
    .Y(_00338_),
    .A1(net158),
    .A2(_00332_));
 sg13g2_xor2_1 _08305_ (.B(_00338_),
    .A(_00330_),
    .X(_00339_));
 sg13g2_xor2_1 _08306_ (.B(_00339_),
    .A(_00326_),
    .X(_00340_));
 sg13g2_xnor2_1 _08307_ (.Y(_00341_),
    .A(_00322_),
    .B(_00340_));
 sg13g2_o21ai_1 _08308_ (.B1(_00303_),
    .Y(_00342_),
    .A1(_00294_),
    .A2(_00295_));
 sg13g2_nor3_1 _08309_ (.A(_00294_),
    .B(_00295_),
    .C(_00303_),
    .Y(_00343_));
 sg13g2_a21oi_1 _08310_ (.A1(_00300_),
    .A2(_00342_),
    .Y(_00344_),
    .B1(_00343_));
 sg13g2_xnor2_1 _08311_ (.Y(_00345_),
    .A(_00341_),
    .B(_00344_));
 sg13g2_xnor2_1 _08312_ (.Y(_00346_),
    .A(_00319_),
    .B(_00345_));
 sg13g2_nand2_2 _08313_ (.Y(_00347_),
    .A(_00309_),
    .B(_00346_));
 sg13g2_nor2_1 _08314_ (.A(_00319_),
    .B(_00344_),
    .Y(_00348_));
 sg13g2_nand2_1 _08315_ (.Y(_00349_),
    .A(_00319_),
    .B(_00344_));
 sg13g2_o21ai_1 _08316_ (.B1(_00349_),
    .Y(_00350_),
    .A1(_00341_),
    .A2(_00348_));
 sg13g2_buf_1 _08317_ (.A(_00350_),
    .X(_00351_));
 sg13g2_nor2_1 _08318_ (.A(_00293_),
    .B(_00326_),
    .Y(_00352_));
 sg13g2_nor2_1 _08319_ (.A(_00339_),
    .B(_00352_),
    .Y(_00353_));
 sg13g2_nand2_1 _08320_ (.Y(_00354_),
    .A(_00293_),
    .B(_00326_));
 sg13g2_mux2_1 _08321_ (.A0(_00354_),
    .A1(_00326_),
    .S(_00244_),
    .X(_00355_));
 sg13g2_nor2_1 _08322_ (.A(_00320_),
    .B(_00354_),
    .Y(_00356_));
 sg13g2_nor3_1 _08323_ (.A(net30),
    .B(_00326_),
    .C(_00339_),
    .Y(_00357_));
 sg13g2_nor3_1 _08324_ (.A(net85),
    .B(_00356_),
    .C(_00357_),
    .Y(_00358_));
 sg13g2_a21oi_1 _08325_ (.A1(net85),
    .A2(_00355_),
    .Y(_00359_),
    .B1(_00358_));
 sg13g2_a21oi_2 _08326_ (.B1(_00359_),
    .Y(_00360_),
    .A2(_00353_),
    .A1(_00273_));
 sg13g2_buf_1 _08327_ (.A(net158),
    .X(_00361_));
 sg13g2_buf_1 _08328_ (.A(net201),
    .X(_00362_));
 sg13g2_buf_1 _08329_ (.A(net267),
    .X(_00363_));
 sg13g2_a21oi_1 _08330_ (.A1(_00362_),
    .A2(_00329_),
    .Y(_00364_),
    .B1(net200));
 sg13g2_nor2_1 _08331_ (.A(net128),
    .B(_00364_),
    .Y(_00365_));
 sg13g2_buf_1 _08332_ (.A(net249),
    .X(_00366_));
 sg13g2_inv_1 _08333_ (.Y(_00367_),
    .A(_00330_));
 sg13g2_buf_1 _08334_ (.A(net248),
    .X(_00368_));
 sg13g2_nor2_1 _08335_ (.A(net198),
    .B(net200),
    .Y(_00369_));
 sg13g2_a221oi_1 _08336_ (.B2(net198),
    .C1(_00369_),
    .B1(_00335_),
    .A1(net199),
    .Y(_00370_),
    .A2(_00367_));
 sg13g2_buf_1 _08337_ (.A(_00366_),
    .X(_00371_));
 sg13g2_nor2_1 _08338_ (.A(net156),
    .B(_00367_),
    .Y(_00372_));
 sg13g2_nor3_2 _08339_ (.A(_00365_),
    .B(_00370_),
    .C(_00372_),
    .Y(_00373_));
 sg13g2_nor2b_1 _08340_ (.A(_00273_),
    .B_N(_00326_),
    .Y(_00374_));
 sg13g2_nor3_1 _08341_ (.A(_00320_),
    .B(_00250_),
    .C(_00326_),
    .Y(_00375_));
 sg13g2_nor2_1 _08342_ (.A(_00374_),
    .B(_00375_),
    .Y(_00376_));
 sg13g2_buf_1 _08343_ (.A(_00376_),
    .X(_00377_));
 sg13g2_o21ai_1 _08344_ (.B1(_00362_),
    .Y(_00378_),
    .A1(_00287_),
    .A2(net95));
 sg13g2_nand2b_1 _08345_ (.Y(_00379_),
    .B(net95),
    .A_N(_00284_));
 sg13g2_a21oi_1 _08346_ (.A1(_00378_),
    .A2(_00379_),
    .Y(_00380_),
    .B1(net200));
 sg13g2_buf_1 _08347_ (.A(_00380_),
    .X(_00381_));
 sg13g2_buf_1 _08348_ (.A(net159),
    .X(_00382_));
 sg13g2_nor2_1 _08349_ (.A(_00333_),
    .B(_00331_),
    .Y(_00383_));
 sg13g2_xnor2_1 _08350_ (.Y(_00384_),
    .A(_00366_),
    .B(net159));
 sg13g2_a22oi_1 _08351_ (.Y(_00385_),
    .B1(_00384_),
    .B2(net248),
    .A2(_00383_),
    .A1(_00382_));
 sg13g2_xnor2_1 _08352_ (.Y(_00386_),
    .A(net67),
    .B(_00385_));
 sg13g2_xnor2_1 _08353_ (.Y(_00387_),
    .A(_00377_),
    .B(_00386_));
 sg13g2_xnor2_1 _08354_ (.Y(_00388_),
    .A(_00373_),
    .B(_00387_));
 sg13g2_xnor2_1 _08355_ (.Y(_00389_),
    .A(_00360_),
    .B(_00388_));
 sg13g2_nand2_1 _08356_ (.Y(_00390_),
    .A(_00351_),
    .B(_00389_));
 sg13g2_nand2_1 _08357_ (.Y(_00391_),
    .A(_00360_),
    .B(_00373_));
 sg13g2_nor2_1 _08358_ (.A(_00360_),
    .B(_00373_),
    .Y(_00392_));
 sg13g2_a21oi_1 _08359_ (.A1(_00387_),
    .A2(_00391_),
    .Y(_00393_),
    .B1(_00392_));
 sg13g2_nand2b_1 _08360_ (.Y(_00394_),
    .B(_00326_),
    .A_N(_00273_));
 sg13g2_buf_1 _08361_ (.A(_00394_),
    .X(_00395_));
 sg13g2_a21o_1 _08362_ (.A2(_00379_),
    .A1(_00378_),
    .B1(net200),
    .X(_00396_));
 sg13g2_buf_1 _08363_ (.A(_00396_),
    .X(_00397_));
 sg13g2_nor2_1 _08364_ (.A(net27),
    .B(net67),
    .Y(_00398_));
 sg13g2_inv_2 _08365_ (.Y(_00399_),
    .A(_00377_));
 sg13g2_nor2_1 _08366_ (.A(_00399_),
    .B(_00385_),
    .Y(_00400_));
 sg13g2_o21ai_1 _08367_ (.B1(_00395_),
    .Y(_00401_),
    .A1(_00398_),
    .A2(_00400_));
 sg13g2_o21ai_1 _08368_ (.B1(_00401_),
    .Y(_00402_),
    .A1(_00395_),
    .A2(_00397_));
 sg13g2_nand2b_1 _08369_ (.Y(_00403_),
    .B(net67),
    .A_N(net158));
 sg13g2_nand2_1 _08370_ (.Y(_00404_),
    .A(_00369_),
    .B(_00403_));
 sg13g2_nor2_1 _08371_ (.A(net198),
    .B(_00403_),
    .Y(_00405_));
 sg13g2_inv_2 _08372_ (.Y(_00406_),
    .A(net198));
 sg13g2_nor2_1 _08373_ (.A(_00406_),
    .B(_00381_),
    .Y(_00407_));
 sg13g2_o21ai_1 _08374_ (.B1(net156),
    .Y(_00408_),
    .A1(_00405_),
    .A2(_00407_));
 sg13g2_o21ai_1 _08375_ (.B1(_00408_),
    .Y(_00409_),
    .A1(net156),
    .A2(_00404_));
 sg13g2_xnor2_1 _08376_ (.Y(_00410_),
    .A(_00402_),
    .B(_00409_));
 sg13g2_xor2_1 _08377_ (.B(_00410_),
    .A(_00393_),
    .X(_00411_));
 sg13g2_nor2_1 _08378_ (.A(_00351_),
    .B(_00389_),
    .Y(_00412_));
 sg13g2_or2_1 _08379_ (.X(_00413_),
    .B(_00412_),
    .A(_00411_));
 sg13g2_nand2_1 _08380_ (.Y(_00414_),
    .A(_04574_),
    .B(_04645_));
 sg13g2_buf_1 _08381_ (.A(_00414_),
    .X(_00415_));
 sg13g2_nand2_1 _08382_ (.Y(_00416_),
    .A(net262),
    .B(net270));
 sg13g2_and2_1 _08383_ (.A(net197),
    .B(_00416_),
    .X(_00417_));
 sg13g2_or2_1 _08384_ (.X(_00418_),
    .B(_00416_),
    .A(net197));
 sg13g2_o21ai_1 _08385_ (.B1(_00418_),
    .Y(_00419_),
    .A1(net202),
    .A2(_00417_));
 sg13g2_nand2_2 _08386_ (.Y(_00420_),
    .A(_04626_),
    .B(net264));
 sg13g2_nor2_1 _08387_ (.A(_04959_),
    .B(_04988_),
    .Y(_00421_));
 sg13g2_o21ai_1 _08388_ (.B1(_04949_),
    .Y(_00422_),
    .A1(_00420_),
    .A2(_00421_));
 sg13g2_nand2_1 _08389_ (.Y(_00423_),
    .A(net203),
    .B(_00422_));
 sg13g2_xor2_1 _08390_ (.B(_00423_),
    .A(_00419_),
    .X(_00424_));
 sg13g2_xnor2_1 _08391_ (.Y(_00425_),
    .A(_04605_),
    .B(_04655_));
 sg13g2_xnor2_1 _08392_ (.Y(_00426_),
    .A(_04563_),
    .B(_00425_));
 sg13g2_buf_2 _08393_ (.A(_00426_),
    .X(_00427_));
 sg13g2_xnor2_1 _08394_ (.Y(_00428_),
    .A(_00424_),
    .B(_00427_));
 sg13g2_buf_1 _08395_ (.A(net251),
    .X(_00429_));
 sg13g2_nand3_1 _08396_ (.B(net196),
    .C(net250),
    .A(net203),
    .Y(_00430_));
 sg13g2_buf_1 _08397_ (.A(_00430_),
    .X(_00431_));
 sg13g2_nand2b_1 _08398_ (.Y(_00432_),
    .B(net263),
    .A_N(_00246_));
 sg13g2_xor2_1 _08399_ (.B(_00420_),
    .A(_00432_),
    .X(_00433_));
 sg13g2_buf_2 _08400_ (.A(_00433_),
    .X(_00434_));
 sg13g2_nand2_1 _08401_ (.Y(_00435_),
    .A(_00431_),
    .B(_00434_));
 sg13g2_inv_1 _08402_ (.Y(_00436_),
    .A(_07493_));
 sg13g2_a21o_1 _08403_ (.A2(_00428_),
    .A1(_00435_),
    .B1(_00436_),
    .X(_00437_));
 sg13g2_o21ai_1 _08404_ (.B1(_00437_),
    .Y(_00438_),
    .A1(_00241_),
    .A2(_00428_));
 sg13g2_nand3_1 _08405_ (.B(_00241_),
    .C(_00247_),
    .A(_00281_),
    .Y(_00439_));
 sg13g2_nand3_1 _08406_ (.B(_00434_),
    .C(_00249_),
    .A(_00242_),
    .Y(_00440_));
 sg13g2_o21ai_1 _08407_ (.B1(_00440_),
    .Y(_00441_),
    .A1(_00428_),
    .A2(_00439_));
 sg13g2_nand2b_1 _08408_ (.Y(_00442_),
    .B(_00434_),
    .A_N(_00428_));
 sg13g2_a21oi_1 _08409_ (.A1(net30),
    .A2(_00442_),
    .Y(_00443_),
    .B1(net85));
 sg13g2_a221oi_1 _08410_ (.B2(_00436_),
    .C1(_00443_),
    .B1(_00441_),
    .A1(_00267_),
    .Y(_00444_),
    .A2(_00438_));
 sg13g2_xnor2_1 _08411_ (.Y(_00445_),
    .A(_04845_),
    .B(_04736_));
 sg13g2_nand2_1 _08412_ (.Y(_00446_),
    .A(_00423_),
    .B(_00427_));
 sg13g2_nor2_1 _08413_ (.A(_00423_),
    .B(_00427_),
    .Y(_00447_));
 sg13g2_a21oi_1 _08414_ (.A1(_00419_),
    .A2(_00446_),
    .Y(_00448_),
    .B1(_00447_));
 sg13g2_inv_2 _08415_ (.Y(_00449_),
    .A(net302));
 sg13g2_buf_1 _08416_ (.A(_00449_),
    .X(_00450_));
 sg13g2_nand2_1 _08417_ (.Y(_00451_),
    .A(net195),
    .B(_00245_));
 sg13g2_o21ai_1 _08418_ (.B1(_00418_),
    .Y(_00452_),
    .A1(_00420_),
    .A2(_00417_));
 sg13g2_buf_1 _08419_ (.A(_00452_),
    .X(_00453_));
 sg13g2_nor2b_1 _08420_ (.A(_00453_),
    .B_N(_00427_),
    .Y(_00454_));
 sg13g2_nand2b_1 _08421_ (.Y(_00455_),
    .B(_00453_),
    .A_N(_00427_));
 sg13g2_o21ai_1 _08422_ (.B1(_00455_),
    .Y(_00456_),
    .A1(_00451_),
    .A2(_00454_));
 sg13g2_buf_1 _08423_ (.A(_00456_),
    .X(_00457_));
 sg13g2_xnor2_1 _08424_ (.Y(_00458_),
    .A(_00448_),
    .B(_00457_));
 sg13g2_xnor2_1 _08425_ (.Y(_00459_),
    .A(_00445_),
    .B(_00458_));
 sg13g2_nand2_1 _08426_ (.Y(_00460_),
    .A(_00273_),
    .B(_00250_));
 sg13g2_xor2_1 _08427_ (.B(_00460_),
    .A(_00261_),
    .X(_00461_));
 sg13g2_xor2_1 _08428_ (.B(_00461_),
    .A(_00459_),
    .X(_00462_));
 sg13g2_xnor2_1 _08429_ (.Y(_00463_),
    .A(_00444_),
    .B(_00462_));
 sg13g2_nand2_1 _08430_ (.Y(_00464_),
    .A(net263),
    .B(_04978_));
 sg13g2_nand2_1 _08431_ (.Y(_00465_),
    .A(_04615_),
    .B(net266));
 sg13g2_nand2_2 _08432_ (.Y(_00466_),
    .A(net308),
    .B(net302));
 sg13g2_xor2_1 _08433_ (.B(_00466_),
    .A(_00465_),
    .X(_00467_));
 sg13g2_xnor2_1 _08434_ (.Y(_00468_),
    .A(_00464_),
    .B(_00467_));
 sg13g2_buf_1 _08435_ (.A(_00468_),
    .X(_00469_));
 sg13g2_and2_1 _08436_ (.A(_00469_),
    .B(_00434_),
    .X(_00470_));
 sg13g2_nor2_1 _08437_ (.A(_00241_),
    .B(_00434_),
    .Y(_00471_));
 sg13g2_and2_1 _08438_ (.A(_00464_),
    .B(_00466_),
    .X(_00472_));
 sg13g2_or2_1 _08439_ (.X(_00473_),
    .B(_00466_),
    .A(_00464_));
 sg13g2_o21ai_1 _08440_ (.B1(_00473_),
    .Y(_00474_),
    .A1(_00465_),
    .A2(_00472_));
 sg13g2_buf_1 _08441_ (.A(_00474_),
    .X(_00475_));
 sg13g2_nor2_1 _08442_ (.A(net202),
    .B(net270),
    .Y(_00476_));
 sg13g2_nor2b_1 _08443_ (.A(_00476_),
    .B_N(_00416_),
    .Y(_00477_));
 sg13g2_xnor2_1 _08444_ (.Y(_00478_),
    .A(net197),
    .B(_00477_));
 sg13g2_xnor2_1 _08445_ (.Y(_00479_),
    .A(_00475_),
    .B(_00478_));
 sg13g2_o21ai_1 _08446_ (.B1(_00479_),
    .Y(_00480_),
    .A1(_00470_),
    .A2(_00471_));
 sg13g2_nand2_1 _08447_ (.Y(_00481_),
    .A(_00469_),
    .B(_00242_));
 sg13g2_a21oi_1 _08448_ (.A1(_00469_),
    .A2(_00431_),
    .Y(_00482_),
    .B1(_00479_));
 sg13g2_nand2_1 _08449_ (.Y(_00483_),
    .A(_00241_),
    .B(_00479_));
 sg13g2_mux4_1 _08450_ (.S0(_07493_),
    .A0(_00481_),
    .A1(_00482_),
    .A2(_00483_),
    .A3(_00431_),
    .S1(_00434_),
    .X(_00484_));
 sg13g2_nand2_1 _08451_ (.Y(_00485_),
    .A(_00480_),
    .B(_00484_));
 sg13g2_a21oi_1 _08452_ (.A1(_00283_),
    .A2(_04595_),
    .Y(_00486_),
    .B1(net197));
 sg13g2_a21oi_1 _08453_ (.A1(_00475_),
    .A2(net197),
    .Y(_00487_),
    .B1(_00486_));
 sg13g2_nor2_1 _08454_ (.A(_00475_),
    .B(net197),
    .Y(_00488_));
 sg13g2_a21oi_1 _08455_ (.A1(_00283_),
    .A2(net197),
    .Y(_00489_),
    .B1(_00488_));
 sg13g2_xnor2_1 _08456_ (.Y(_00490_),
    .A(net269),
    .B(net197));
 sg13g2_a21o_1 _08457_ (.A2(_00490_),
    .A1(_00475_),
    .B1(_05233_),
    .X(_00491_));
 sg13g2_o21ai_1 _08458_ (.B1(_00491_),
    .Y(_00492_),
    .A1(_05179_),
    .A2(_00489_));
 sg13g2_a21o_1 _08459_ (.A2(_00487_),
    .A1(_05179_),
    .B1(_00492_),
    .X(_00493_));
 sg13g2_nand2_1 _08460_ (.Y(_00494_),
    .A(net262),
    .B(net305));
 sg13g2_and2_1 _08461_ (.A(_00466_),
    .B(_00494_),
    .X(_00495_));
 sg13g2_or2_1 _08462_ (.X(_00496_),
    .B(_00494_),
    .A(_00466_));
 sg13g2_o21ai_1 _08463_ (.B1(_00496_),
    .Y(_00497_),
    .A1(_00465_),
    .A2(_00495_));
 sg13g2_inv_1 _08464_ (.Y(_00498_),
    .A(_00497_));
 sg13g2_xor2_1 _08465_ (.B(_00416_),
    .A(_00420_),
    .X(_00499_));
 sg13g2_xor2_1 _08466_ (.B(_00499_),
    .A(_00415_),
    .X(_00500_));
 sg13g2_xnor2_1 _08467_ (.Y(_00501_),
    .A(_00415_),
    .B(_00499_));
 sg13g2_nor2b_1 _08468_ (.A(net304),
    .B_N(net301),
    .Y(_00502_));
 sg13g2_a21oi_1 _08469_ (.A1(_00497_),
    .A2(_00501_),
    .Y(_00503_),
    .B1(_00502_));
 sg13g2_a21oi_2 _08470_ (.B1(_00503_),
    .Y(_00504_),
    .A2(_00500_),
    .A1(_00498_));
 sg13g2_xor2_1 _08471_ (.B(_00453_),
    .A(_00451_),
    .X(_00505_));
 sg13g2_xnor2_1 _08472_ (.Y(_00506_),
    .A(_00504_),
    .B(_00505_));
 sg13g2_xnor2_1 _08473_ (.Y(_00507_),
    .A(_00493_),
    .B(_00506_));
 sg13g2_o21ai_1 _08474_ (.B1(_07503_),
    .Y(_00508_),
    .A1(_00244_),
    .A2(_00434_));
 sg13g2_xnor2_1 _08475_ (.Y(_00509_),
    .A(_00249_),
    .B(_00424_));
 sg13g2_xnor2_1 _08476_ (.Y(_00510_),
    .A(_00508_),
    .B(_00509_));
 sg13g2_xor2_1 _08477_ (.B(_00510_),
    .A(_00507_),
    .X(_00511_));
 sg13g2_nand2_1 _08478_ (.Y(_00512_),
    .A(_00485_),
    .B(_00511_));
 sg13g2_or3_1 _08479_ (.A(_00507_),
    .B(_00510_),
    .C(_00427_),
    .X(_00513_));
 sg13g2_nand3_1 _08480_ (.B(_00510_),
    .C(_00427_),
    .A(_00507_),
    .Y(_00514_));
 sg13g2_nand3_1 _08481_ (.B(_00513_),
    .C(_00514_),
    .A(_00512_),
    .Y(_00515_));
 sg13g2_xor2_1 _08482_ (.B(_00427_),
    .A(_00505_),
    .X(_00516_));
 sg13g2_nand2_1 _08483_ (.Y(_00517_),
    .A(_00504_),
    .B(_00516_));
 sg13g2_nor2_1 _08484_ (.A(_00504_),
    .B(_00516_),
    .Y(_00518_));
 sg13g2_a21o_1 _08485_ (.A2(_00517_),
    .A1(_00493_),
    .B1(_00518_),
    .X(_00519_));
 sg13g2_buf_1 _08486_ (.A(_00519_),
    .X(_00520_));
 sg13g2_xnor2_1 _08487_ (.Y(_00521_),
    .A(_00515_),
    .B(_00520_));
 sg13g2_xnor2_1 _08488_ (.Y(_00522_),
    .A(_00463_),
    .B(_00521_));
 sg13g2_buf_1 _08489_ (.A(_00522_),
    .X(_00523_));
 sg13g2_nand2_1 _08490_ (.Y(_00524_),
    .A(net308),
    .B(_04897_));
 sg13g2_nand2_1 _08491_ (.Y(_00525_),
    .A(net262),
    .B(net302));
 sg13g2_nand2_1 _08492_ (.Y(_00526_),
    .A(_04615_),
    .B(net303));
 sg13g2_a21o_1 _08493_ (.A2(_00525_),
    .A1(_00524_),
    .B1(_00526_),
    .X(_00527_));
 sg13g2_o21ai_1 _08494_ (.B1(_00527_),
    .Y(_00528_),
    .A1(_00524_),
    .A2(_00525_));
 sg13g2_buf_2 _08495_ (.A(_00528_),
    .X(_00529_));
 sg13g2_o21ai_1 _08496_ (.B1(_05169_),
    .Y(_00530_),
    .A1(net269),
    .A2(_00529_));
 sg13g2_nand2_1 _08497_ (.Y(_00531_),
    .A(_04746_),
    .B(_00529_));
 sg13g2_inv_2 _08498_ (.Y(_00532_),
    .A(_04635_));
 sg13g2_a21oi_2 _08499_ (.B1(_00532_),
    .Y(_00533_),
    .A2(_00531_),
    .A1(_00530_));
 sg13g2_xor2_1 _08500_ (.B(_00494_),
    .A(_00467_),
    .X(_00534_));
 sg13g2_inv_1 _08501_ (.Y(_00535_),
    .A(_00529_));
 sg13g2_inv_1 _08502_ (.Y(_00536_),
    .A(_04918_));
 sg13g2_buf_1 _08503_ (.A(_00536_),
    .X(_00537_));
 sg13g2_nand2_1 _08504_ (.Y(_00538_),
    .A(net263),
    .B(_00537_));
 sg13g2_a21o_1 _08505_ (.A2(_00535_),
    .A1(_00534_),
    .B1(_00538_),
    .X(_00539_));
 sg13g2_o21ai_1 _08506_ (.B1(_00539_),
    .Y(_00540_),
    .A1(_00534_),
    .A2(_00535_));
 sg13g2_buf_1 _08507_ (.A(_00540_),
    .X(_00541_));
 sg13g2_xnor2_1 _08508_ (.Y(_00542_),
    .A(_00502_),
    .B(_00497_));
 sg13g2_xnor2_1 _08509_ (.Y(_00543_),
    .A(_00542_),
    .B(_00501_));
 sg13g2_o21ai_1 _08510_ (.B1(_00543_),
    .Y(_00544_),
    .A1(_00533_),
    .A2(_00541_));
 sg13g2_nand2_1 _08511_ (.Y(_00545_),
    .A(_00533_),
    .B(_00541_));
 sg13g2_nand2_2 _08512_ (.Y(_00546_),
    .A(_00544_),
    .B(_00545_));
 sg13g2_xor2_1 _08513_ (.B(_00525_),
    .A(_00524_),
    .X(_00547_));
 sg13g2_or2_1 _08514_ (.X(_00548_),
    .B(_00547_),
    .A(_00526_));
 sg13g2_nand2_1 _08515_ (.Y(_00549_),
    .A(_00526_),
    .B(_00547_));
 sg13g2_nand2_1 _08516_ (.Y(_00550_),
    .A(_00548_),
    .B(_00549_));
 sg13g2_buf_1 _08517_ (.A(_00550_),
    .X(_00551_));
 sg13g2_nand2_1 _08518_ (.Y(_00552_),
    .A(net262),
    .B(net266));
 sg13g2_nand2_2 _08519_ (.Y(_00553_),
    .A(net309),
    .B(net302));
 sg13g2_and2_1 _08520_ (.A(_04488_),
    .B(net304),
    .X(_00554_));
 sg13g2_buf_1 _08521_ (.A(_00554_),
    .X(_00555_));
 sg13g2_nor2_1 _08522_ (.A(_00282_),
    .B(_00449_),
    .Y(_00556_));
 sg13g2_and2_1 _08523_ (.A(net308),
    .B(net303),
    .X(_00557_));
 sg13g2_a21oi_1 _08524_ (.A1(_00555_),
    .A2(_00556_),
    .Y(_00558_),
    .B1(_00557_));
 sg13g2_a21oi_2 _08525_ (.B1(_00558_),
    .Y(_00559_),
    .A2(_00553_),
    .A1(_00552_));
 sg13g2_nor2_1 _08526_ (.A(net93),
    .B(_00559_),
    .Y(_00560_));
 sg13g2_nand2_1 _08527_ (.Y(_00561_),
    .A(net263),
    .B(_07499_));
 sg13g2_nand2_1 _08528_ (.Y(_00562_),
    .A(net93),
    .B(_00559_));
 sg13g2_o21ai_1 _08529_ (.B1(_00562_),
    .Y(_00563_),
    .A1(_00560_),
    .A2(_00561_));
 sg13g2_buf_1 _08530_ (.A(_00563_),
    .X(_00564_));
 sg13g2_nand2_1 _08531_ (.Y(_00565_),
    .A(_04468_),
    .B(_04918_));
 sg13g2_a22oi_1 _08532_ (.Y(_00566_),
    .B1(_00557_),
    .B2(_00555_),
    .A2(net296),
    .A1(_04615_));
 sg13g2_a21oi_2 _08533_ (.B1(_00566_),
    .Y(_00567_),
    .A2(_00552_),
    .A1(_00565_));
 sg13g2_nand2_1 _08534_ (.Y(_00568_),
    .A(_00567_),
    .B(_00287_));
 sg13g2_nor2_1 _08535_ (.A(_00567_),
    .B(_00287_),
    .Y(_00569_));
 sg13g2_a21oi_1 _08536_ (.A1(_05442_),
    .A2(_00568_),
    .Y(_00570_),
    .B1(_00569_));
 sg13g2_xnor2_1 _08537_ (.Y(_00571_),
    .A(_00538_),
    .B(_00534_));
 sg13g2_xnor2_1 _08538_ (.Y(_00572_),
    .A(_00571_),
    .B(_00529_));
 sg13g2_a21o_1 _08539_ (.A2(_00570_),
    .A1(_00564_),
    .B1(_00572_),
    .X(_00573_));
 sg13g2_o21ai_1 _08540_ (.B1(_00573_),
    .Y(_00574_),
    .A1(_00564_),
    .A2(_00570_));
 sg13g2_buf_1 _08541_ (.A(_00574_),
    .X(_00575_));
 sg13g2_mux2_1 _08542_ (.A0(_00241_),
    .A1(_07501_),
    .S(_07493_),
    .X(_00576_));
 sg13g2_xnor2_1 _08543_ (.Y(_00577_),
    .A(_00469_),
    .B(_00576_));
 sg13g2_xor2_1 _08544_ (.B(net309),
    .A(net262),
    .X(_00578_));
 sg13g2_nand2_1 _08545_ (.Y(_00579_),
    .A(net268),
    .B(_00578_));
 sg13g2_xnor2_1 _08546_ (.Y(_00580_),
    .A(_00579_),
    .B(_00529_));
 sg13g2_nand2_1 _08547_ (.Y(_00581_),
    .A(_00577_),
    .B(_00580_));
 sg13g2_nand2_1 _08548_ (.Y(_00582_),
    .A(net80),
    .B(_07230_));
 sg13g2_a21o_1 _08549_ (.A2(_00582_),
    .A1(_07352_),
    .B1(_07305_),
    .X(_00583_));
 sg13g2_or2_1 _08550_ (.X(_00584_),
    .B(_07137_),
    .A(_07302_));
 sg13g2_nand2_1 _08551_ (.Y(_00585_),
    .A(net80),
    .B(_00584_));
 sg13g2_o21ai_1 _08552_ (.B1(_07230_),
    .Y(_00586_),
    .A1(net80),
    .A2(_00584_));
 sg13g2_a21o_1 _08553_ (.A2(_00586_),
    .A1(_00585_),
    .B1(_07352_),
    .X(_00587_));
 sg13g2_a21o_1 _08554_ (.A2(_00587_),
    .A1(_00583_),
    .B1(_07421_),
    .X(_00588_));
 sg13g2_buf_1 _08555_ (.A(_00588_),
    .X(_00589_));
 sg13g2_or3_1 _08556_ (.A(_07272_),
    .B(_07371_),
    .C(_07423_),
    .X(_00590_));
 sg13g2_buf_1 _08557_ (.A(_00590_),
    .X(_00591_));
 sg13g2_nor2_1 _08558_ (.A(_00036_),
    .B(_07490_),
    .Y(_00592_));
 sg13g2_nand3_1 _08559_ (.B(_00591_),
    .C(_00592_),
    .A(_00589_),
    .Y(_00593_));
 sg13g2_a21oi_1 _08560_ (.A1(_07384_),
    .A2(_07445_),
    .Y(_00594_),
    .B1(_07443_));
 sg13g2_nor3_1 _08561_ (.A(_07401_),
    .B(_07412_),
    .C(_07415_),
    .Y(_00595_));
 sg13g2_a21oi_1 _08562_ (.A1(_07384_),
    .A2(_00595_),
    .Y(_00596_),
    .B1(_07435_));
 sg13g2_or3_1 _08563_ (.A(_07474_),
    .B(_00594_),
    .C(_00596_),
    .X(_00597_));
 sg13g2_nor2b_1 _08564_ (.A(_07474_),
    .B_N(_07435_),
    .Y(_00598_));
 sg13g2_nor2_1 _08565_ (.A(_07474_),
    .B(_07435_),
    .Y(_00599_));
 sg13g2_and4_1 _08566_ (.A(_07384_),
    .B(_07474_),
    .C(_07435_),
    .D(_00595_),
    .X(_00600_));
 sg13g2_a221oi_1 _08567_ (.B2(_07447_),
    .C1(_00600_),
    .B1(_00599_),
    .A1(_00598_),
    .Y(_00601_),
    .A2(_00594_));
 sg13g2_buf_1 _08568_ (.A(_00601_),
    .X(_00602_));
 sg13g2_nand3_1 _08569_ (.B(net295),
    .C(_07490_),
    .A(_05070_),
    .Y(_00603_));
 sg13g2_nand2b_1 _08570_ (.Y(_00604_),
    .B(_00603_),
    .A_N(_00592_));
 sg13g2_nand3_1 _08571_ (.B(_00602_),
    .C(_00604_),
    .A(_00597_),
    .Y(_00605_));
 sg13g2_nand2b_1 _08572_ (.Y(_00606_),
    .B(_07490_),
    .A_N(_00036_));
 sg13g2_or3_1 _08573_ (.A(_00602_),
    .B(_00591_),
    .C(_00606_),
    .X(_00607_));
 sg13g2_nand3b_1 _08574_ (.B(net295),
    .C(_05070_),
    .Y(_00608_),
    .A_N(_07490_));
 sg13g2_nor2_1 _08575_ (.A(_00602_),
    .B(_00608_),
    .Y(_00609_));
 sg13g2_nor3_1 _08576_ (.A(_07474_),
    .B(_00594_),
    .C(_00596_),
    .Y(_00610_));
 sg13g2_a21oi_1 _08577_ (.A1(_00583_),
    .A2(_00587_),
    .Y(_00611_),
    .B1(_07421_));
 sg13g2_nor3_1 _08578_ (.A(_00610_),
    .B(_00611_),
    .C(_00603_),
    .Y(_00612_));
 sg13g2_mux2_1 _08579_ (.A0(_00609_),
    .A1(_00612_),
    .S(_00591_),
    .X(_00613_));
 sg13g2_nand2b_1 _08580_ (.Y(_00614_),
    .B(_00611_),
    .A_N(_00602_));
 sg13g2_a22oi_1 _08581_ (.Y(_00615_),
    .B1(_00614_),
    .B2(_00597_),
    .A2(_00608_),
    .A1(_00606_));
 sg13g2_nor2_1 _08582_ (.A(_00613_),
    .B(_00615_),
    .Y(_00616_));
 sg13g2_and4_1 _08583_ (.A(_00593_),
    .B(_00605_),
    .C(_00607_),
    .D(_00616_),
    .X(_00617_));
 sg13g2_xor2_1 _08584_ (.B(net296),
    .A(_07505_),
    .X(_00618_));
 sg13g2_nand2_1 _08585_ (.Y(_00619_),
    .A(_05080_),
    .B(_00618_));
 sg13g2_xnor2_1 _08586_ (.Y(_00620_),
    .A(_00619_),
    .B(_07493_));
 sg13g2_nand2_1 _08587_ (.Y(_00621_),
    .A(net93),
    .B(_00620_));
 sg13g2_nor2_1 _08588_ (.A(net93),
    .B(_00620_),
    .Y(_00622_));
 sg13g2_a21oi_1 _08589_ (.A1(_00617_),
    .A2(_00621_),
    .Y(_00623_),
    .B1(_00622_));
 sg13g2_o21ai_1 _08590_ (.B1(_00623_),
    .Y(_00624_),
    .A1(_00577_),
    .A2(_00580_));
 sg13g2_nand2_1 _08591_ (.Y(_00625_),
    .A(_00581_),
    .B(_00624_));
 sg13g2_nand2_1 _08592_ (.Y(_00626_),
    .A(_00469_),
    .B(_00431_));
 sg13g2_nor2_1 _08593_ (.A(_00469_),
    .B(_00241_),
    .Y(_00627_));
 sg13g2_a21oi_1 _08594_ (.A1(_07493_),
    .A2(_00626_),
    .Y(_00628_),
    .B1(_00627_));
 sg13g2_xnor2_1 _08595_ (.Y(_00629_),
    .A(_00541_),
    .B(_00542_));
 sg13g2_xnor2_1 _08596_ (.Y(_00630_),
    .A(_00533_),
    .B(_00629_));
 sg13g2_xor2_1 _08597_ (.B(_00476_),
    .A(_00432_),
    .X(_00631_));
 sg13g2_xnor2_1 _08598_ (.Y(_00632_),
    .A(_00475_),
    .B(_00631_));
 sg13g2_xnor2_1 _08599_ (.Y(_00633_),
    .A(_00630_),
    .B(_00632_));
 sg13g2_xnor2_1 _08600_ (.Y(_00634_),
    .A(_00628_),
    .B(_00633_));
 sg13g2_xnor2_1 _08601_ (.Y(_00635_),
    .A(_00625_),
    .B(_00634_));
 sg13g2_buf_2 _08602_ (.A(_00635_),
    .X(_00636_));
 sg13g2_xnor2_1 _08603_ (.Y(_00637_),
    .A(_00579_),
    .B(_00577_));
 sg13g2_xnor2_1 _08604_ (.Y(_00638_),
    .A(_00623_),
    .B(_00637_));
 sg13g2_buf_2 _08605_ (.A(_00638_),
    .X(_00639_));
 sg13g2_xor2_1 _08606_ (.B(_00570_),
    .A(_00571_),
    .X(_00640_));
 sg13g2_xnor2_1 _08607_ (.Y(_00641_),
    .A(_00564_),
    .B(_00640_));
 sg13g2_nand2_1 _08608_ (.Y(_00642_),
    .A(_00639_),
    .B(_00641_));
 sg13g2_inv_1 _08609_ (.Y(_00643_),
    .A(_00641_));
 sg13g2_nand2b_1 _08610_ (.Y(_00644_),
    .B(_00643_),
    .A_N(_00639_));
 sg13g2_xor2_1 _08611_ (.B(_00287_),
    .A(_05442_),
    .X(_00645_));
 sg13g2_xnor2_1 _08612_ (.Y(_00646_),
    .A(_00567_),
    .B(_00645_));
 sg13g2_a21oi_1 _08613_ (.A1(_00589_),
    .A2(_00591_),
    .Y(_00647_),
    .B1(_00602_));
 sg13g2_o21ai_1 _08614_ (.B1(_07490_),
    .Y(_00648_),
    .A1(_00610_),
    .A2(_00647_));
 sg13g2_buf_2 _08615_ (.A(_00648_),
    .X(_00649_));
 sg13g2_or3_1 _08616_ (.A(_07490_),
    .B(_00610_),
    .C(_00647_),
    .X(_00650_));
 sg13g2_buf_1 _08617_ (.A(_00650_),
    .X(_00651_));
 sg13g2_nand2_1 _08618_ (.Y(_00652_),
    .A(_05080_),
    .B(net252));
 sg13g2_buf_1 _08619_ (.A(_00652_),
    .X(_00653_));
 sg13g2_a21oi_1 _08620_ (.A1(_00649_),
    .A2(_00651_),
    .Y(_00654_),
    .B1(_00653_));
 sg13g2_and3_1 _08621_ (.X(_00655_),
    .A(_00653_),
    .B(_00649_),
    .C(_00651_));
 sg13g2_nand3_1 _08622_ (.B(_07347_),
    .C(_07384_),
    .A(_07307_),
    .Y(_00656_));
 sg13g2_a21oi_1 _08623_ (.A1(_07307_),
    .A2(_07347_),
    .Y(_00657_),
    .B1(_07384_));
 sg13g2_a21oi_1 _08624_ (.A1(_07420_),
    .A2(_00656_),
    .Y(_00658_),
    .B1(_00657_));
 sg13g2_xor2_1 _08625_ (.B(_07435_),
    .A(_07443_),
    .X(_00659_));
 sg13g2_nor2_1 _08626_ (.A(_07423_),
    .B(_07448_),
    .Y(_00660_));
 sg13g2_nand2_1 _08627_ (.Y(_00661_),
    .A(_04468_),
    .B(net329));
 sg13g2_nand2_2 _08628_ (.Y(_00662_),
    .A(_04615_),
    .B(_07494_));
 sg13g2_or2_1 _08629_ (.X(_00663_),
    .B(_00662_),
    .A(_00661_));
 sg13g2_nand2_1 _08630_ (.Y(_00664_),
    .A(_00663_),
    .B(_07477_));
 sg13g2_a221oi_1 _08631_ (.B2(_07377_),
    .C1(_00664_),
    .B1(_00660_),
    .A1(_00658_),
    .Y(_00665_),
    .A2(_00659_));
 sg13g2_and2_1 _08632_ (.A(_00663_),
    .B(_07476_),
    .X(_00666_));
 sg13g2_nand3_1 _08633_ (.B(_00660_),
    .C(_00666_),
    .A(_07377_),
    .Y(_00667_));
 sg13g2_and2_1 _08634_ (.A(_00658_),
    .B(_00659_),
    .X(_00668_));
 sg13g2_a22oi_1 _08635_ (.Y(_00669_),
    .B1(_00668_),
    .B2(_00666_),
    .A2(_00662_),
    .A1(_00661_));
 sg13g2_nand3b_1 _08636_ (.B(_00667_),
    .C(_00669_),
    .Y(_00670_),
    .A_N(_00665_));
 sg13g2_buf_8 _08637_ (.A(_00670_),
    .X(_00671_));
 sg13g2_nand2_2 _08638_ (.Y(_00672_),
    .A(_04615_),
    .B(net329));
 sg13g2_xnor2_1 _08639_ (.Y(_00673_),
    .A(_00565_),
    .B(_00555_));
 sg13g2_xor2_1 _08640_ (.B(_00673_),
    .A(_00672_),
    .X(_00674_));
 sg13g2_inv_1 _08641_ (.Y(_00675_),
    .A(_00674_));
 sg13g2_nand2b_1 _08642_ (.Y(_00676_),
    .B(_00675_),
    .A_N(_00671_));
 sg13g2_o21ai_1 _08643_ (.B1(_00676_),
    .Y(_00677_),
    .A1(_00654_),
    .A2(_00655_));
 sg13g2_nand2_1 _08644_ (.Y(_00678_),
    .A(_00671_),
    .B(_00674_));
 sg13g2_and3_1 _08645_ (.X(_00679_),
    .A(_00646_),
    .B(_00677_),
    .C(_00678_));
 sg13g2_xnor2_1 _08646_ (.Y(_00680_),
    .A(_00617_),
    .B(_00620_));
 sg13g2_buf_2 _08647_ (.A(_00680_),
    .X(_00681_));
 sg13g2_xor2_1 _08648_ (.B(_00681_),
    .A(net93),
    .X(_00682_));
 sg13g2_a21o_1 _08649_ (.A2(_00678_),
    .A1(_00677_),
    .B1(_00646_),
    .X(_00683_));
 sg13g2_buf_1 _08650_ (.A(_00683_),
    .X(_00684_));
 sg13g2_o21ai_1 _08651_ (.B1(_00684_),
    .Y(_00685_),
    .A1(_00679_),
    .A2(_00682_));
 sg13g2_a21oi_1 _08652_ (.A1(_00642_),
    .A2(_00644_),
    .Y(_00686_),
    .B1(_00685_));
 sg13g2_and3_1 _08653_ (.X(_00687_),
    .A(_00639_),
    .B(_00643_),
    .C(_00529_));
 sg13g2_nor3_1 _08654_ (.A(_00639_),
    .B(_00643_),
    .C(_00529_),
    .Y(_00688_));
 sg13g2_nor3_1 _08655_ (.A(_00686_),
    .B(_00687_),
    .C(_00688_),
    .Y(_00689_));
 sg13g2_buf_2 _08656_ (.A(_00689_),
    .X(_00690_));
 sg13g2_o21ai_1 _08657_ (.B1(_00690_),
    .Y(_00691_),
    .A1(_00575_),
    .A2(_00636_));
 sg13g2_inv_1 _08658_ (.Y(_00692_),
    .A(_00691_));
 sg13g2_a21oi_2 _08659_ (.B1(_00692_),
    .Y(_00693_),
    .A2(_00636_),
    .A1(_00575_));
 sg13g2_inv_1 _08660_ (.Y(_00694_),
    .A(_00693_));
 sg13g2_xnor2_1 _08661_ (.Y(_00695_),
    .A(_00628_),
    .B(_00632_));
 sg13g2_nand2_1 _08662_ (.Y(_00696_),
    .A(_00630_),
    .B(_00501_));
 sg13g2_nand3b_1 _08663_ (.B(_00695_),
    .C(_00500_),
    .Y(_00697_),
    .A_N(_00630_));
 sg13g2_o21ai_1 _08664_ (.B1(_00697_),
    .Y(_00698_),
    .A1(_00695_),
    .A2(_00696_));
 sg13g2_a21oi_2 _08665_ (.B1(_00698_),
    .Y(_00699_),
    .A2(_00634_),
    .A1(_00625_));
 sg13g2_nand2_1 _08666_ (.Y(_00700_),
    .A(_00694_),
    .B(_00699_));
 sg13g2_nor2_1 _08667_ (.A(_00694_),
    .B(_00699_),
    .Y(_00701_));
 sg13g2_a21o_1 _08668_ (.A2(_00700_),
    .A1(_00546_),
    .B1(_00701_),
    .X(_00702_));
 sg13g2_xnor2_1 _08669_ (.Y(_00703_),
    .A(_00485_),
    .B(_00511_));
 sg13g2_xnor2_1 _08670_ (.Y(_00704_),
    .A(_00703_),
    .B(_00546_));
 sg13g2_xnor2_1 _08671_ (.Y(_00705_),
    .A(_00699_),
    .B(_00704_));
 sg13g2_buf_1 _08672_ (.A(_00705_),
    .X(_00706_));
 sg13g2_and2_1 _08673_ (.A(_00693_),
    .B(_00706_),
    .X(_00707_));
 sg13g2_buf_2 _08674_ (.A(_00707_),
    .X(_00708_));
 sg13g2_inv_1 _08675_ (.Y(_00709_),
    .A(_00703_));
 sg13g2_nand2_1 _08676_ (.Y(_00710_),
    .A(_00709_),
    .B(_00546_));
 sg13g2_nor2_1 _08677_ (.A(_00709_),
    .B(_00546_),
    .Y(_00711_));
 sg13g2_a21oi_1 _08678_ (.A1(_00699_),
    .A2(_00710_),
    .Y(_00712_),
    .B1(_00711_));
 sg13g2_xnor2_1 _08679_ (.Y(_00713_),
    .A(_00523_),
    .B(_00712_));
 sg13g2_buf_1 _08680_ (.A(_00713_),
    .X(_00714_));
 sg13g2_nand2b_1 _08681_ (.Y(_00715_),
    .B(_00714_),
    .A_N(_00708_));
 sg13g2_xnor2_1 _08682_ (.Y(_00716_),
    .A(_00575_),
    .B(_00636_));
 sg13g2_xor2_1 _08683_ (.B(_00716_),
    .A(_00690_),
    .X(_00717_));
 sg13g2_buf_1 _08684_ (.A(_00717_),
    .X(_00718_));
 sg13g2_nand2b_1 _08685_ (.Y(_00719_),
    .B(_00526_),
    .A_N(_00547_));
 sg13g2_nand2b_1 _08686_ (.Y(_00720_),
    .B(_00547_),
    .A_N(_00526_));
 sg13g2_nor2_1 _08687_ (.A(net267),
    .B(_07505_),
    .Y(_00721_));
 sg13g2_buf_1 _08688_ (.A(_00721_),
    .X(_00722_));
 sg13g2_and3_1 _08689_ (.X(_00723_),
    .A(_00671_),
    .B(_00649_),
    .C(_00651_));
 sg13g2_a21oi_1 _08690_ (.A1(_00649_),
    .A2(_00651_),
    .Y(_00724_),
    .B1(_00671_));
 sg13g2_nor3_1 _08691_ (.A(_00674_),
    .B(_00723_),
    .C(_00724_),
    .Y(_00725_));
 sg13g2_nand3_1 _08692_ (.B(_00649_),
    .C(_00651_),
    .A(_00671_),
    .Y(_00726_));
 sg13g2_a21o_1 _08693_ (.A2(_00651_),
    .A1(_00649_),
    .B1(_00671_),
    .X(_00727_));
 sg13g2_a21oi_1 _08694_ (.A1(_00726_),
    .A2(_00727_),
    .Y(_00728_),
    .B1(_00675_));
 sg13g2_nor2_1 _08695_ (.A(_00725_),
    .B(_00728_),
    .Y(_00729_));
 sg13g2_xnor2_1 _08696_ (.Y(_00730_),
    .A(_00722_),
    .B(_00729_));
 sg13g2_a21oi_1 _08697_ (.A1(_07377_),
    .A2(_00660_),
    .Y(_00731_),
    .B1(_00668_));
 sg13g2_and2_1 _08698_ (.A(_04574_),
    .B(net296),
    .X(_00732_));
 sg13g2_buf_1 _08699_ (.A(_00732_),
    .X(_00733_));
 sg13g2_xnor2_1 _08700_ (.Y(_00734_),
    .A(_00733_),
    .B(_07476_));
 sg13g2_xnor2_1 _08701_ (.Y(_00735_),
    .A(_00731_),
    .B(_00734_));
 sg13g2_xnor2_1 _08702_ (.Y(_00736_),
    .A(_00662_),
    .B(_00735_));
 sg13g2_and2_1 _08703_ (.A(_04468_),
    .B(net310),
    .X(_00737_));
 sg13g2_nor2_1 _08704_ (.A(net252),
    .B(net204),
    .Y(_00738_));
 sg13g2_nand2_1 _08705_ (.Y(_00739_),
    .A(net310),
    .B(net329));
 sg13g2_nand2_1 _08706_ (.Y(_00740_),
    .A(net308),
    .B(net295));
 sg13g2_nand2_1 _08707_ (.Y(_00741_),
    .A(_00739_),
    .B(_00740_));
 sg13g2_nor2_1 _08708_ (.A(net34),
    .B(_07371_),
    .Y(_00742_));
 sg13g2_xor2_1 _08709_ (.B(_07447_),
    .A(_07435_),
    .X(_00743_));
 sg13g2_nor2_1 _08710_ (.A(_00743_),
    .B(_00611_),
    .Y(_00744_));
 sg13g2_nor2_1 _08711_ (.A(_07448_),
    .B(_00589_),
    .Y(_00745_));
 sg13g2_a221oi_1 _08712_ (.B2(_00744_),
    .C1(_00745_),
    .B1(_00591_),
    .A1(_00742_),
    .Y(_00746_),
    .A2(_00660_));
 sg13g2_buf_2 _08713_ (.A(_00746_),
    .X(_00747_));
 sg13g2_a22oi_1 _08714_ (.Y(_00748_),
    .B1(_00741_),
    .B2(_00747_),
    .A2(_00738_),
    .A1(_00737_));
 sg13g2_buf_1 _08715_ (.A(_00748_),
    .X(_00749_));
 sg13g2_and2_1 _08716_ (.A(net262),
    .B(net303),
    .X(_00750_));
 sg13g2_buf_1 _08717_ (.A(_00750_),
    .X(_00751_));
 sg13g2_nand2_1 _08718_ (.Y(_00752_),
    .A(net309),
    .B(_04897_));
 sg13g2_buf_1 _08719_ (.A(_00752_),
    .X(_00753_));
 sg13g2_xnor2_1 _08720_ (.Y(_00754_),
    .A(_00751_),
    .B(net194));
 sg13g2_nand2_1 _08721_ (.Y(_00755_),
    .A(net307),
    .B(_05008_));
 sg13g2_buf_2 _08722_ (.A(_00755_),
    .X(_00756_));
 sg13g2_xnor2_1 _08723_ (.Y(_00757_),
    .A(_00754_),
    .B(_00756_));
 sg13g2_nand2b_1 _08724_ (.Y(_00758_),
    .B(_00757_),
    .A_N(_00749_));
 sg13g2_nor2b_1 _08725_ (.A(_00757_),
    .B_N(_00749_),
    .Y(_00759_));
 sg13g2_a21oi_2 _08726_ (.B1(_00759_),
    .Y(_00760_),
    .A2(_00758_),
    .A1(_00736_));
 sg13g2_and2_1 _08727_ (.A(net307),
    .B(net302),
    .X(_00761_));
 sg13g2_buf_1 _08728_ (.A(_00761_),
    .X(_00762_));
 sg13g2_nor2_1 _08729_ (.A(_05573_),
    .B(net194),
    .Y(_00763_));
 sg13g2_a21oi_1 _08730_ (.A1(_00751_),
    .A2(net194),
    .Y(_00764_),
    .B1(_00763_));
 sg13g2_nand2_2 _08731_ (.Y(_00765_),
    .A(_05169_),
    .B(_04928_));
 sg13g2_a21oi_1 _08732_ (.A1(_00765_),
    .A2(net194),
    .Y(_00766_),
    .B1(_00532_));
 sg13g2_a21oi_1 _08733_ (.A1(_00532_),
    .A2(_00764_),
    .Y(_00767_),
    .B1(_00766_));
 sg13g2_xnor2_1 _08734_ (.Y(_00768_),
    .A(_05573_),
    .B(_00751_));
 sg13g2_nor2_1 _08735_ (.A(net194),
    .B(_00762_),
    .Y(_00769_));
 sg13g2_a22oi_1 _08736_ (.Y(_00770_),
    .B1(_00768_),
    .B2(_00769_),
    .A2(_00767_),
    .A1(_00762_));
 sg13g2_xnor2_1 _08737_ (.Y(_00771_),
    .A(_00553_),
    .B(_00770_));
 sg13g2_inv_1 _08738_ (.Y(_00772_),
    .A(_00771_));
 sg13g2_nand2_1 _08739_ (.Y(_00773_),
    .A(_00760_),
    .B(_00772_));
 sg13g2_nor2_1 _08740_ (.A(_00760_),
    .B(_00772_),
    .Y(_00774_));
 sg13g2_a21o_1 _08741_ (.A2(_00773_),
    .A1(_00730_),
    .B1(_00774_),
    .X(_00775_));
 sg13g2_buf_2 _08742_ (.A(_00775_),
    .X(_00776_));
 sg13g2_xnor2_1 _08743_ (.Y(_00777_),
    .A(_00673_),
    .B(_00556_));
 sg13g2_a21o_1 _08744_ (.A2(_00765_),
    .A1(_00661_),
    .B1(_00662_),
    .X(_00778_));
 sg13g2_o21ai_1 _08745_ (.B1(_00778_),
    .Y(_00779_),
    .A1(_00661_),
    .A2(_00765_));
 sg13g2_nor2_1 _08746_ (.A(_00672_),
    .B(_00777_),
    .Y(_00780_));
 sg13g2_nor2_1 _08747_ (.A(_00779_),
    .B(_00780_),
    .Y(_00781_));
 sg13g2_a21oi_2 _08748_ (.B1(_00781_),
    .Y(_00782_),
    .A2(_00777_),
    .A1(_00672_));
 sg13g2_xor2_1 _08749_ (.B(_00561_),
    .A(_00559_),
    .X(_00783_));
 sg13g2_nor3_1 _08750_ (.A(net305),
    .B(_05573_),
    .C(_00756_),
    .Y(_00784_));
 sg13g2_o21ai_1 _08751_ (.B1(_00765_),
    .Y(_00785_),
    .A1(net194),
    .A2(_00756_));
 sg13g2_nand2b_1 _08752_ (.Y(_00786_),
    .B(_00785_),
    .A_N(_00784_));
 sg13g2_a22oi_1 _08753_ (.Y(_00787_),
    .B1(_00756_),
    .B2(_05573_),
    .A2(net194),
    .A1(_00532_));
 sg13g2_a21oi_1 _08754_ (.A1(_00556_),
    .A2(_00751_),
    .Y(_00788_),
    .B1(_00787_));
 sg13g2_a221oi_1 _08755_ (.B2(_00553_),
    .C1(_00788_),
    .B1(_00786_),
    .A1(net194),
    .Y(_00789_),
    .A2(_00756_));
 sg13g2_buf_1 _08756_ (.A(_00789_),
    .X(_00790_));
 sg13g2_xnor2_1 _08757_ (.Y(_00791_),
    .A(_00783_),
    .B(_00790_));
 sg13g2_xnor2_1 _08758_ (.Y(_00792_),
    .A(_00782_),
    .B(_00791_));
 sg13g2_inv_1 _08759_ (.Y(_00793_),
    .A(_00792_));
 sg13g2_nand3_1 _08760_ (.B(_00677_),
    .C(_00678_),
    .A(_00646_),
    .Y(_00794_));
 sg13g2_buf_1 _08761_ (.A(_00794_),
    .X(_00795_));
 sg13g2_a21o_1 _08762_ (.A2(_00684_),
    .A1(_00795_),
    .B1(_00681_),
    .X(_00796_));
 sg13g2_nand3_1 _08763_ (.B(_00681_),
    .C(_00684_),
    .A(_00795_),
    .Y(_00797_));
 sg13g2_nand3_1 _08764_ (.B(_00796_),
    .C(_00797_),
    .A(_00793_),
    .Y(_00798_));
 sg13g2_buf_1 _08765_ (.A(_00798_),
    .X(_00799_));
 sg13g2_a21oi_1 _08766_ (.A1(_00796_),
    .A2(_00797_),
    .Y(_00800_),
    .B1(_00793_));
 sg13g2_a221oi_1 _08767_ (.B2(_00799_),
    .C1(_00800_),
    .B1(_00776_),
    .A1(_00719_),
    .Y(_00801_),
    .A2(_00720_));
 sg13g2_buf_1 _08768_ (.A(_00801_),
    .X(_00802_));
 sg13g2_a21oi_1 _08769_ (.A1(_00795_),
    .A2(_00684_),
    .Y(_00803_),
    .B1(_00681_));
 sg13g2_and3_1 _08770_ (.X(_00804_),
    .A(_00795_),
    .B(_00681_),
    .C(_00684_));
 sg13g2_o21ai_1 _08771_ (.B1(_00792_),
    .Y(_00805_),
    .A1(_00803_),
    .A2(_00804_));
 sg13g2_nor3_1 _08772_ (.A(_00792_),
    .B(_00803_),
    .C(_00804_),
    .Y(_00806_));
 sg13g2_a221oi_1 _08773_ (.B2(_00805_),
    .C1(_00806_),
    .B1(_00776_),
    .A1(_00548_),
    .Y(_00807_),
    .A2(_00549_));
 sg13g2_buf_1 _08774_ (.A(_00807_),
    .X(_00808_));
 sg13g2_nor2_1 _08775_ (.A(_00802_),
    .B(_00808_),
    .Y(_00809_));
 sg13g2_buf_8 _08776_ (.A(_00809_),
    .X(_00810_));
 sg13g2_xor2_1 _08777_ (.B(_00754_),
    .A(_00749_),
    .X(_00811_));
 sg13g2_xnor2_1 _08778_ (.Y(_00812_),
    .A(_00736_),
    .B(_00811_));
 sg13g2_nor2_1 _08779_ (.A(_00532_),
    .B(_00449_),
    .Y(_00813_));
 sg13g2_buf_2 _08780_ (.A(_00813_),
    .X(_00814_));
 sg13g2_nand2_1 _08781_ (.Y(_00815_),
    .A(_04584_),
    .B(net304));
 sg13g2_nand2_1 _08782_ (.Y(_00816_),
    .A(net309),
    .B(_04918_));
 sg13g2_xor2_1 _08783_ (.B(_00816_),
    .A(_00815_),
    .X(_00817_));
 sg13g2_xnor2_1 _08784_ (.Y(_00818_),
    .A(_00814_),
    .B(_00817_));
 sg13g2_buf_1 _08785_ (.A(_00818_),
    .X(_00819_));
 sg13g2_xnor2_1 _08786_ (.Y(_00820_),
    .A(_00739_),
    .B(_00740_));
 sg13g2_nand2_1 _08787_ (.Y(_00821_),
    .A(net111),
    .B(_00820_));
 sg13g2_xor2_1 _08788_ (.B(_00740_),
    .A(_00739_),
    .X(_00822_));
 sg13g2_buf_2 _08789_ (.A(_00822_),
    .X(_00823_));
 sg13g2_nand2_1 _08790_ (.Y(_00824_),
    .A(net111),
    .B(_00823_));
 sg13g2_mux2_1 _08791_ (.A0(_00821_),
    .A1(_00824_),
    .S(_00747_),
    .X(_00825_));
 sg13g2_xor2_1 _08792_ (.B(_07423_),
    .A(_07377_),
    .X(_00826_));
 sg13g2_nand2_1 _08793_ (.Y(_00827_),
    .A(_04488_),
    .B(net295));
 sg13g2_buf_2 _08794_ (.A(_00827_),
    .X(_00828_));
 sg13g2_nand2_1 _08795_ (.Y(_00829_),
    .A(_04542_),
    .B(net329));
 sg13g2_buf_1 _08796_ (.A(_00829_),
    .X(_00830_));
 sg13g2_or2_1 _08797_ (.X(_00831_),
    .B(net193),
    .A(_00828_));
 sg13g2_and2_1 _08798_ (.A(_00828_),
    .B(net193),
    .X(_00832_));
 sg13g2_a21oi_1 _08799_ (.A1(_00826_),
    .A2(_00831_),
    .Y(_00833_),
    .B1(_00832_));
 sg13g2_nor2_1 _08800_ (.A(net111),
    .B(_00823_),
    .Y(_00834_));
 sg13g2_nor3_1 _08801_ (.A(_00747_),
    .B(_00819_),
    .C(_00820_),
    .Y(_00835_));
 sg13g2_a221oi_1 _08802_ (.B2(_00747_),
    .C1(_00835_),
    .B1(_00834_),
    .A1(_00825_),
    .Y(_00836_),
    .A2(_00833_));
 sg13g2_buf_1 _08803_ (.A(_00836_),
    .X(_00837_));
 sg13g2_xor2_1 _08804_ (.B(_00753_),
    .A(_05573_),
    .X(_00838_));
 sg13g2_mux2_1 _08805_ (.A0(_00837_),
    .A1(_00762_),
    .S(_00838_),
    .X(_00839_));
 sg13g2_nand2b_1 _08806_ (.Y(_00840_),
    .B(_00839_),
    .A_N(_00812_));
 sg13g2_mux2_1 _08807_ (.A0(_00756_),
    .A1(_00837_),
    .S(_00838_),
    .X(_00841_));
 sg13g2_nand2_1 _08808_ (.Y(_00842_),
    .A(_00812_),
    .B(_00841_));
 sg13g2_xnor2_1 _08809_ (.Y(_00843_),
    .A(_00672_),
    .B(_00779_));
 sg13g2_xnor2_1 _08810_ (.Y(_00844_),
    .A(_00777_),
    .B(_00843_));
 sg13g2_xor2_1 _08811_ (.B(net265),
    .A(_04626_),
    .X(_00845_));
 sg13g2_nor4_2 _08812_ (.A(net252),
    .B(net204),
    .C(_07313_),
    .Y(_00846_),
    .D(_00845_));
 sg13g2_nor2b_1 _08813_ (.A(_00814_),
    .B_N(_00815_),
    .Y(_00847_));
 sg13g2_o21ai_1 _08814_ (.B1(_05398_),
    .Y(_00848_),
    .A1(_00847_),
    .A2(_00816_));
 sg13g2_buf_1 _08815_ (.A(_00848_),
    .X(_00849_));
 sg13g2_xnor2_1 _08816_ (.Y(_00850_),
    .A(_00846_),
    .B(_00849_));
 sg13g2_xnor2_1 _08817_ (.Y(_00851_),
    .A(_00844_),
    .B(_00850_));
 sg13g2_a21oi_2 _08818_ (.B1(_00851_),
    .Y(_00852_),
    .A2(_00842_),
    .A1(_00840_));
 sg13g2_inv_1 _08819_ (.Y(_00853_),
    .A(_00852_));
 sg13g2_nand3_1 _08820_ (.B(_00726_),
    .C(_00727_),
    .A(_00675_),
    .Y(_00854_));
 sg13g2_o21ai_1 _08821_ (.B1(_00674_),
    .Y(_00855_),
    .A1(_00723_),
    .A2(_00724_));
 sg13g2_nand3_1 _08822_ (.B(_00854_),
    .C(_00855_),
    .A(_00772_),
    .Y(_00856_));
 sg13g2_o21ai_1 _08823_ (.B1(_00771_),
    .Y(_00857_),
    .A1(_00725_),
    .A2(_00728_));
 sg13g2_a21oi_1 _08824_ (.A1(_00856_),
    .A2(_00857_),
    .Y(_00858_),
    .B1(_00760_));
 sg13g2_inv_2 _08825_ (.Y(_00859_),
    .A(_00760_));
 sg13g2_nor3_1 _08826_ (.A(_00771_),
    .B(_00725_),
    .C(_00728_),
    .Y(_00860_));
 sg13g2_a21oi_1 _08827_ (.A1(_00854_),
    .A2(_00855_),
    .Y(_00861_),
    .B1(_00772_));
 sg13g2_nor3_1 _08828_ (.A(_00859_),
    .B(_00860_),
    .C(_00861_),
    .Y(_00862_));
 sg13g2_nor3_1 _08829_ (.A(_00653_),
    .B(_00858_),
    .C(_00862_),
    .Y(_00863_));
 sg13g2_o21ai_1 _08830_ (.B1(_00859_),
    .Y(_00864_),
    .A1(_00860_),
    .A2(_00861_));
 sg13g2_nand3_1 _08831_ (.B(_00856_),
    .C(_00857_),
    .A(_00760_),
    .Y(_00865_));
 sg13g2_buf_1 _08832_ (.A(_00865_),
    .X(_00866_));
 sg13g2_a21oi_1 _08833_ (.A1(_00864_),
    .A2(_00866_),
    .Y(_00867_),
    .B1(_00722_));
 sg13g2_nand3_1 _08834_ (.B(_00840_),
    .C(_00842_),
    .A(_00851_),
    .Y(_00868_));
 sg13g2_buf_1 _08835_ (.A(_00868_),
    .X(_00869_));
 sg13g2_o21ai_1 _08836_ (.B1(_00869_),
    .Y(_00870_),
    .A1(_00863_),
    .A2(_00867_));
 sg13g2_nand2_1 _08837_ (.Y(_00871_),
    .A(_00846_),
    .B(_00849_));
 sg13g2_o21ai_1 _08838_ (.B1(_00844_),
    .Y(_00872_),
    .A1(_00846_),
    .A2(_00849_));
 sg13g2_nand2_1 _08839_ (.Y(_00873_),
    .A(_00871_),
    .B(_00872_));
 sg13g2_buf_2 _08840_ (.A(_00873_),
    .X(_00874_));
 sg13g2_nand2_1 _08841_ (.Y(_00875_),
    .A(_00795_),
    .B(_00684_));
 sg13g2_xnor2_1 _08842_ (.Y(_00876_),
    .A(_00681_),
    .B(_00792_));
 sg13g2_xnor2_1 _08843_ (.Y(_00877_),
    .A(_00875_),
    .B(_00876_));
 sg13g2_xnor2_1 _08844_ (.Y(_00878_),
    .A(_00776_),
    .B(_00877_));
 sg13g2_a22oi_1 _08845_ (.Y(_00879_),
    .B1(_00874_),
    .B2(_00878_),
    .A2(_00870_),
    .A1(_00853_));
 sg13g2_buf_1 _08846_ (.A(_00879_),
    .X(_00880_));
 sg13g2_nor2_1 _08847_ (.A(_00874_),
    .B(_00878_),
    .Y(_00881_));
 sg13g2_nor2_1 _08848_ (.A(_00880_),
    .B(_00881_),
    .Y(_00882_));
 sg13g2_buf_2 _08849_ (.A(_00882_),
    .X(_00883_));
 sg13g2_xnor2_1 _08850_ (.Y(_00884_),
    .A(net93),
    .B(_00783_));
 sg13g2_a21o_1 _08851_ (.A2(_00790_),
    .A1(_00782_),
    .B1(_00884_),
    .X(_00885_));
 sg13g2_o21ai_1 _08852_ (.B1(_00885_),
    .Y(_00886_),
    .A1(_00782_),
    .A2(_00790_));
 sg13g2_buf_1 _08853_ (.A(_00886_),
    .X(_00887_));
 sg13g2_xnor2_1 _08854_ (.Y(_00888_),
    .A(_00639_),
    .B(_00643_));
 sg13g2_xnor2_1 _08855_ (.Y(_00889_),
    .A(_00685_),
    .B(_00888_));
 sg13g2_buf_2 _08856_ (.A(_00889_),
    .X(_00890_));
 sg13g2_nor2_1 _08857_ (.A(_00887_),
    .B(_00890_),
    .Y(_00891_));
 sg13g2_buf_2 _08858_ (.A(_00891_),
    .X(_00892_));
 sg13g2_buf_1 _08859_ (.A(_00887_),
    .X(_00893_));
 sg13g2_nand2_1 _08860_ (.Y(_00894_),
    .A(_00893_),
    .B(_00890_));
 sg13g2_buf_1 _08861_ (.A(_00894_),
    .X(_00895_));
 sg13g2_o21ai_1 _08862_ (.B1(_00895_),
    .Y(_00896_),
    .A1(_00883_),
    .A2(_00892_));
 sg13g2_nor2_1 _08863_ (.A(_00883_),
    .B(_00895_),
    .Y(_00897_));
 sg13g2_a21oi_1 _08864_ (.A1(net22),
    .A2(_00896_),
    .Y(_00898_),
    .B1(_00897_));
 sg13g2_nor2_1 _08865_ (.A(net93),
    .B(_00799_),
    .Y(_00899_));
 sg13g2_a21oi_1 _08866_ (.A1(net93),
    .A2(_00800_),
    .Y(_00900_),
    .B1(_00899_));
 sg13g2_nor2_1 _08867_ (.A(_00776_),
    .B(_00900_),
    .Y(_00901_));
 sg13g2_o21ai_1 _08868_ (.B1(_00799_),
    .Y(_00902_),
    .A1(_00776_),
    .A2(_00800_));
 sg13g2_o21ai_1 _08869_ (.B1(_00805_),
    .Y(_00903_),
    .A1(_00776_),
    .A2(_00806_));
 sg13g2_mux2_1 _08870_ (.A0(_00902_),
    .A1(_00903_),
    .S(_00551_),
    .X(_00904_));
 sg13g2_a21o_1 _08871_ (.A2(_00904_),
    .A1(_00874_),
    .B1(_00901_),
    .X(_00905_));
 sg13g2_and2_1 _08872_ (.A(_00853_),
    .B(_00870_),
    .X(_00906_));
 sg13g2_a22oi_1 _08873_ (.Y(_00907_),
    .B1(_00905_),
    .B2(_00906_),
    .A2(_00901_),
    .A1(_00874_));
 sg13g2_nand2_1 _08874_ (.Y(_00908_),
    .A(_00718_),
    .B(_00892_));
 sg13g2_xnor2_1 _08875_ (.Y(_00909_),
    .A(_00693_),
    .B(_00706_));
 sg13g2_o21ai_1 _08876_ (.B1(_00909_),
    .Y(_00910_),
    .A1(_00907_),
    .A2(_00908_));
 sg13g2_o21ai_1 _08877_ (.B1(_00910_),
    .Y(_00911_),
    .A1(_00718_),
    .A2(_00898_));
 sg13g2_buf_1 _08878_ (.A(_00911_),
    .X(_00912_));
 sg13g2_xor2_1 _08879_ (.B(_00877_),
    .A(_00776_),
    .X(_00913_));
 sg13g2_nand2b_1 _08880_ (.Y(_00914_),
    .B(_00913_),
    .A_N(_00874_));
 sg13g2_or2_1 _08881_ (.X(_00915_),
    .B(_00808_),
    .A(_00802_));
 sg13g2_buf_1 _08882_ (.A(_00915_),
    .X(_00916_));
 sg13g2_nand3b_1 _08883_ (.B(_00914_),
    .C(_00916_),
    .Y(_00917_),
    .A_N(_00880_));
 sg13g2_buf_1 _08884_ (.A(_00917_),
    .X(_00918_));
 sg13g2_o21ai_1 _08885_ (.B1(_00810_),
    .Y(_00919_),
    .A1(_00880_),
    .A2(_00881_));
 sg13g2_buf_1 _08886_ (.A(_00919_),
    .X(_00920_));
 sg13g2_and2_1 _08887_ (.A(net52),
    .B(_00890_),
    .X(_00921_));
 sg13g2_nor2_1 _08888_ (.A(_00921_),
    .B(_00892_),
    .Y(_00922_));
 sg13g2_nand3_1 _08889_ (.B(_00920_),
    .C(_00922_),
    .A(_00918_),
    .Y(_00923_));
 sg13g2_a21o_1 _08890_ (.A2(_00920_),
    .A1(_00918_),
    .B1(_00922_),
    .X(_00924_));
 sg13g2_buf_1 _08891_ (.A(_00924_),
    .X(_00925_));
 sg13g2_nand2_1 _08892_ (.Y(_00926_),
    .A(_00923_),
    .B(_00925_));
 sg13g2_inv_1 _08893_ (.Y(_00927_),
    .A(_00926_));
 sg13g2_xor2_1 _08894_ (.B(_00768_),
    .A(_00749_),
    .X(_00928_));
 sg13g2_xnor2_1 _08895_ (.Y(_00929_),
    .A(_00837_),
    .B(_00928_));
 sg13g2_xnor2_1 _08896_ (.Y(_00930_),
    .A(_00736_),
    .B(_00929_));
 sg13g2_buf_8 _08897_ (.A(_00930_),
    .X(_00931_));
 sg13g2_inv_1 _08898_ (.Y(_00932_),
    .A(net304));
 sg13g2_nor2_1 _08899_ (.A(_00932_),
    .B(net247),
    .Y(_00933_));
 sg13g2_nand2_1 _08900_ (.Y(_00934_),
    .A(_04595_),
    .B(_04928_));
 sg13g2_nand2_1 _08901_ (.Y(_00935_),
    .A(net305),
    .B(net266));
 sg13g2_xor2_1 _08902_ (.B(_00935_),
    .A(_00934_),
    .X(_00936_));
 sg13g2_buf_1 _08903_ (.A(_00936_),
    .X(_00937_));
 sg13g2_a21o_1 _08904_ (.A2(net193),
    .A1(net111),
    .B1(_00449_),
    .X(_00938_));
 sg13g2_o21ai_1 _08905_ (.B1(_00938_),
    .Y(_00939_),
    .A1(net111),
    .A2(net193));
 sg13g2_a22oi_1 _08906_ (.Y(_00940_),
    .B1(_00937_),
    .B2(_00939_),
    .A2(_00933_),
    .A1(_00287_));
 sg13g2_buf_2 _08907_ (.A(_00940_),
    .X(_00941_));
 sg13g2_nor2b_1 _08908_ (.A(_00852_),
    .B_N(_00869_),
    .Y(_00942_));
 sg13g2_nor3_2 _08909_ (.A(_00863_),
    .B(_00867_),
    .C(_00942_),
    .Y(_00943_));
 sg13g2_nand3_1 _08910_ (.B(_00864_),
    .C(_00866_),
    .A(_00722_),
    .Y(_00944_));
 sg13g2_o21ai_1 _08911_ (.B1(_00653_),
    .Y(_00945_),
    .A1(_00858_),
    .A2(_00862_));
 sg13g2_nand2b_1 _08912_ (.Y(_00946_),
    .B(_00869_),
    .A_N(_00852_));
 sg13g2_a21oi_2 _08913_ (.B1(_00946_),
    .Y(_00947_),
    .A2(_00945_),
    .A1(_00944_));
 sg13g2_o21ai_1 _08914_ (.B1(net262),
    .Y(_00948_),
    .A1(net196),
    .A2(_04988_));
 sg13g2_a21oi_1 _08915_ (.A1(_07496_),
    .A2(_00733_),
    .Y(_00949_),
    .B1(_00765_));
 sg13g2_a21oi_1 _08916_ (.A1(_00733_),
    .A2(_00948_),
    .Y(_00950_),
    .B1(_00949_));
 sg13g2_xnor2_1 _08917_ (.Y(_00951_),
    .A(_00662_),
    .B(_00950_));
 sg13g2_nor2_1 _08918_ (.A(_00282_),
    .B(net204),
    .Y(_00952_));
 sg13g2_buf_2 _08919_ (.A(_00952_),
    .X(_00953_));
 sg13g2_a21oi_1 _08920_ (.A1(_06354_),
    .A2(_06869_),
    .Y(_00954_),
    .B1(_07256_));
 sg13g2_nor2_2 _08921_ (.A(_00282_),
    .B(_07496_),
    .Y(_00955_));
 sg13g2_nor2_1 _08922_ (.A(_07479_),
    .B(_07154_),
    .Y(_00956_));
 sg13g2_nor2_1 _08923_ (.A(_07479_),
    .B(_07137_),
    .Y(_00957_));
 sg13g2_a22oi_1 _08924_ (.Y(_00958_),
    .B1(_00957_),
    .B2(_06101_),
    .A2(_00956_),
    .A1(_07306_));
 sg13g2_o21ai_1 _08925_ (.B1(_07306_),
    .Y(_00959_),
    .A1(_07289_),
    .A2(_07196_));
 sg13g2_nand3b_1 _08926_ (.B(_07289_),
    .C(_07305_),
    .Y(_00960_),
    .A_N(_07230_));
 sg13g2_nand4_1 _08927_ (.B(_00958_),
    .C(_00959_),
    .A(_07349_),
    .Y(_00961_),
    .D(_00960_));
 sg13g2_xnor2_1 _08928_ (.Y(_00962_),
    .A(_07347_),
    .B(_00961_));
 sg13g2_nor3_1 _08929_ (.A(_00954_),
    .B(_00955_),
    .C(_00962_),
    .Y(_00963_));
 sg13g2_and2_1 _08930_ (.A(net307),
    .B(_07498_),
    .X(_00964_));
 sg13g2_buf_1 _08931_ (.A(_00964_),
    .X(_00965_));
 sg13g2_nor3_1 _08932_ (.A(_00954_),
    .B(_00962_),
    .C(_00965_),
    .Y(_00966_));
 sg13g2_nor2_1 _08933_ (.A(_00955_),
    .B(_00965_),
    .Y(_00967_));
 sg13g2_nand2_2 _08934_ (.Y(_00968_),
    .A(_04542_),
    .B(_07504_));
 sg13g2_nand4_1 _08935_ (.B(_07363_),
    .C(_07369_),
    .A(_07351_),
    .Y(_00969_),
    .D(_00968_));
 sg13g2_nand2_1 _08936_ (.Y(_00970_),
    .A(net307),
    .B(_07498_));
 sg13g2_nand4_1 _08937_ (.B(_07363_),
    .C(_07369_),
    .A(_07351_),
    .Y(_00971_),
    .D(_00970_));
 sg13g2_a21oi_1 _08938_ (.A1(_00969_),
    .A2(_00971_),
    .Y(_00972_),
    .B1(_07282_));
 sg13g2_or4_1 _08939_ (.A(_00963_),
    .B(_00966_),
    .C(_00967_),
    .D(_00972_),
    .X(_00973_));
 sg13g2_buf_1 _08940_ (.A(_00973_),
    .X(_00974_));
 sg13g2_xor2_1 _08941_ (.B(net193),
    .A(_00828_),
    .X(_00975_));
 sg13g2_nand2b_1 _08942_ (.Y(_00976_),
    .B(_00975_),
    .A_N(_07423_));
 sg13g2_nand2_1 _08943_ (.Y(_00977_),
    .A(_07423_),
    .B(_00975_));
 sg13g2_mux2_1 _08944_ (.A0(_00976_),
    .A1(_00977_),
    .S(_07377_),
    .X(_00978_));
 sg13g2_nand2b_1 _08945_ (.Y(_00979_),
    .B(_07423_),
    .A_N(_00975_));
 sg13g2_or2_1 _08946_ (.X(_00980_),
    .B(_00975_),
    .A(_07423_));
 sg13g2_mux2_1 _08947_ (.A0(_00979_),
    .A1(_00980_),
    .S(_07377_),
    .X(_00981_));
 sg13g2_nand3b_1 _08948_ (.B(_00978_),
    .C(_00981_),
    .Y(_00982_),
    .A_N(_00974_));
 sg13g2_buf_1 _08949_ (.A(_00982_),
    .X(_00983_));
 sg13g2_and3_1 _08950_ (.X(_00984_),
    .A(net264),
    .B(_00953_),
    .C(_00983_));
 sg13g2_xnor2_1 _08951_ (.Y(_00985_),
    .A(net195),
    .B(net193));
 sg13g2_nor2_1 _08952_ (.A(net111),
    .B(_00985_),
    .Y(_00986_));
 sg13g2_o21ai_1 _08953_ (.B1(_00937_),
    .Y(_00987_),
    .A1(_00984_),
    .A2(_00986_));
 sg13g2_xnor2_1 _08954_ (.Y(_00988_),
    .A(_00747_),
    .B(_00823_));
 sg13g2_xnor2_1 _08955_ (.Y(_00989_),
    .A(_00988_),
    .B(_00833_));
 sg13g2_xnor2_1 _08956_ (.Y(_00990_),
    .A(_00934_),
    .B(_00935_));
 sg13g2_buf_2 _08957_ (.A(_00990_),
    .X(_00991_));
 sg13g2_nand2_2 _08958_ (.Y(_00992_),
    .A(_00981_),
    .B(_00978_));
 sg13g2_nand3_1 _08959_ (.B(_00992_),
    .C(net33),
    .A(_00991_),
    .Y(_00993_));
 sg13g2_nor2_1 _08960_ (.A(net264),
    .B(_00937_),
    .Y(_00994_));
 sg13g2_nand2_1 _08961_ (.Y(_00995_),
    .A(net33),
    .B(_00994_));
 sg13g2_and3_1 _08962_ (.X(_00996_),
    .A(_00449_),
    .B(net193),
    .C(net33));
 sg13g2_o21ai_1 _08963_ (.B1(_00992_),
    .Y(_00997_),
    .A1(_00994_),
    .A2(_00996_));
 sg13g2_and4_1 _08964_ (.A(_00989_),
    .B(_00993_),
    .C(_00995_),
    .D(_00997_),
    .X(_00998_));
 sg13g2_nand4_1 _08965_ (.B(_00937_),
    .C(_00992_),
    .A(_00953_),
    .Y(_00999_),
    .D(_00974_));
 sg13g2_o21ai_1 _08966_ (.B1(net111),
    .Y(_01000_),
    .A1(net193),
    .A2(_00991_));
 sg13g2_and2_1 _08967_ (.A(net195),
    .B(_01000_),
    .X(_01001_));
 sg13g2_nor2_1 _08968_ (.A(_00953_),
    .B(_00991_),
    .Y(_01002_));
 sg13g2_o21ai_1 _08969_ (.B1(net111),
    .Y(_01003_),
    .A1(_00953_),
    .A2(_00991_));
 sg13g2_nand2_1 _08970_ (.Y(_01004_),
    .A(net264),
    .B(_01003_));
 sg13g2_a21oi_1 _08971_ (.A1(_00983_),
    .A2(_01002_),
    .Y(_01005_),
    .B1(_01004_));
 sg13g2_a21o_1 _08972_ (.A2(_01001_),
    .A1(_00999_),
    .B1(_01005_),
    .X(_01006_));
 sg13g2_inv_1 _08973_ (.Y(_01007_),
    .A(_00989_));
 sg13g2_a22oi_1 _08974_ (.Y(_01008_),
    .B1(_01006_),
    .B2(_01007_),
    .A2(_00998_),
    .A1(_00987_));
 sg13g2_buf_2 _08975_ (.A(_01008_),
    .X(_01009_));
 sg13g2_or2_1 _08976_ (.X(_01010_),
    .B(_01009_),
    .A(_00951_));
 sg13g2_buf_1 _08977_ (.A(_01010_),
    .X(_01011_));
 sg13g2_inv_1 _08978_ (.Y(_01012_),
    .A(_01011_));
 sg13g2_nor3_1 _08979_ (.A(_00943_),
    .B(_00947_),
    .C(_01012_),
    .Y(_01013_));
 sg13g2_or3_1 _08980_ (.A(_00931_),
    .B(_00941_),
    .C(_01013_),
    .X(_01014_));
 sg13g2_buf_1 _08981_ (.A(_01014_),
    .X(_01015_));
 sg13g2_nand2_1 _08982_ (.Y(_01016_),
    .A(_00951_),
    .B(_01009_));
 sg13g2_nand2b_1 _08983_ (.Y(_01017_),
    .B(_01016_),
    .A_N(_00931_));
 sg13g2_nand2_1 _08984_ (.Y(_01018_),
    .A(_00941_),
    .B(_01011_));
 sg13g2_nand2_1 _08985_ (.Y(_01019_),
    .A(_01016_),
    .B(_01018_));
 sg13g2_nor2_1 _08986_ (.A(_00943_),
    .B(_00947_),
    .Y(_01020_));
 sg13g2_a21o_1 _08987_ (.A2(_01019_),
    .A1(_01017_),
    .B1(_01020_),
    .X(_01021_));
 sg13g2_buf_1 _08988_ (.A(_01021_),
    .X(_01022_));
 sg13g2_nand2_1 _08989_ (.Y(_01023_),
    .A(_01015_),
    .B(_01022_));
 sg13g2_inv_1 _08990_ (.Y(_01024_),
    .A(_01023_));
 sg13g2_xnor2_1 _08991_ (.Y(_01025_),
    .A(_00941_),
    .B(_00950_));
 sg13g2_xnor2_1 _08992_ (.Y(_01026_),
    .A(_00735_),
    .B(_01025_));
 sg13g2_xnor2_1 _08993_ (.Y(_01027_),
    .A(_00929_),
    .B(_01026_));
 sg13g2_xnor2_1 _08994_ (.Y(_01028_),
    .A(_01009_),
    .B(_01027_));
 sg13g2_or4_1 _08995_ (.A(_00449_),
    .B(_00953_),
    .C(_00991_),
    .D(net33),
    .X(_01029_));
 sg13g2_nand3_1 _08996_ (.B(_00830_),
    .C(net33),
    .A(net195),
    .Y(_01030_));
 sg13g2_mux2_1 _08997_ (.A0(_01029_),
    .A1(_01030_),
    .S(_00992_),
    .X(_01031_));
 sg13g2_nor3_1 _08998_ (.A(net195),
    .B(_00830_),
    .C(_00991_),
    .Y(_01032_));
 sg13g2_o21ai_1 _08999_ (.B1(_00983_),
    .Y(_01033_),
    .A1(_00994_),
    .A2(_01032_));
 sg13g2_nand3_1 _09000_ (.B(_00953_),
    .C(_00937_),
    .A(_00450_),
    .Y(_01034_));
 sg13g2_a21o_1 _09001_ (.A2(net33),
    .A1(_00992_),
    .B1(_01034_),
    .X(_01035_));
 sg13g2_nand4_1 _09002_ (.B(_01031_),
    .C(_01033_),
    .A(_00993_),
    .Y(_01036_),
    .D(_01035_));
 sg13g2_xnor2_1 _09003_ (.Y(_01037_),
    .A(_00989_),
    .B(_01036_));
 sg13g2_buf_2 _09004_ (.A(_01037_),
    .X(_01038_));
 sg13g2_nand2_1 _09005_ (.Y(_01039_),
    .A(net264),
    .B(_04907_));
 sg13g2_nand2_1 _09006_ (.Y(_01040_),
    .A(net305),
    .B(net265));
 sg13g2_nor2_1 _09007_ (.A(_00532_),
    .B(_00537_),
    .Y(_01041_));
 sg13g2_a21oi_1 _09008_ (.A1(_00955_),
    .A2(_01041_),
    .Y(_01042_),
    .B1(_00965_));
 sg13g2_a21oi_1 _09009_ (.A1(_00968_),
    .A2(_01040_),
    .Y(_01043_),
    .B1(_01042_));
 sg13g2_xnor2_1 _09010_ (.Y(_01044_),
    .A(_00953_),
    .B(_00991_));
 sg13g2_nor2_1 _09011_ (.A(_01043_),
    .B(_01044_),
    .Y(_01045_));
 sg13g2_nand2_1 _09012_ (.Y(_01046_),
    .A(_01043_),
    .B(_01044_));
 sg13g2_o21ai_1 _09013_ (.B1(_01046_),
    .Y(_01047_),
    .A1(_01039_),
    .A2(_01045_));
 sg13g2_buf_1 _09014_ (.A(_01047_),
    .X(_01048_));
 sg13g2_nand2_1 _09015_ (.Y(_01049_),
    .A(_01038_),
    .B(_01048_));
 sg13g2_xnor2_1 _09016_ (.Y(_01050_),
    .A(_01039_),
    .B(_01043_));
 sg13g2_mux2_1 _09017_ (.A0(_07371_),
    .A1(_00962_),
    .S(_07282_),
    .X(_01051_));
 sg13g2_buf_1 _09018_ (.A(_01051_),
    .X(_01052_));
 sg13g2_xnor2_1 _09019_ (.Y(_01053_),
    .A(_00968_),
    .B(_00965_));
 sg13g2_xnor2_1 _09020_ (.Y(_01054_),
    .A(_01052_),
    .B(_01053_));
 sg13g2_nand2_1 _09021_ (.Y(_01055_),
    .A(net307),
    .B(_07494_));
 sg13g2_buf_1 _09022_ (.A(_01055_),
    .X(_01056_));
 sg13g2_nor2_1 _09023_ (.A(_07500_),
    .B(_01056_),
    .Y(_01057_));
 sg13g2_a21oi_1 _09024_ (.A1(_07500_),
    .A2(_01056_),
    .Y(_01058_),
    .B1(_01040_));
 sg13g2_nand3_1 _09025_ (.B(_06869_),
    .C(_07256_),
    .A(_06354_),
    .Y(_01059_));
 sg13g2_buf_2 _09026_ (.A(_01059_),
    .X(_01060_));
 sg13g2_and2_1 _09027_ (.A(net34),
    .B(_01060_),
    .X(_01061_));
 sg13g2_buf_2 _09028_ (.A(_01061_),
    .X(_01062_));
 sg13g2_a22oi_1 _09029_ (.Y(_01063_),
    .B1(_01058_),
    .B2(_01062_),
    .A2(_01057_),
    .A1(_01041_));
 sg13g2_nand2_1 _09030_ (.Y(_01064_),
    .A(net335),
    .B(net329));
 sg13g2_nand2_1 _09031_ (.Y(_01065_),
    .A(_01056_),
    .B(_01064_));
 sg13g2_nor2_1 _09032_ (.A(_01056_),
    .B(_01064_),
    .Y(_01066_));
 sg13g2_a221oi_1 _09033_ (.B2(_01062_),
    .C1(_01066_),
    .B1(_01065_),
    .A1(_04645_),
    .Y(_01067_),
    .A2(net265));
 sg13g2_a21o_1 _09034_ (.A2(_01063_),
    .A1(_01054_),
    .B1(_01067_),
    .X(_01068_));
 sg13g2_buf_1 _09035_ (.A(_01068_),
    .X(_01069_));
 sg13g2_nor2_1 _09036_ (.A(_01050_),
    .B(_01044_),
    .Y(_01070_));
 sg13g2_a21oi_1 _09037_ (.A1(_01050_),
    .A2(_01069_),
    .Y(_01071_),
    .B1(_01070_));
 sg13g2_inv_1 _09038_ (.Y(_01072_),
    .A(_01050_));
 sg13g2_and2_1 _09039_ (.A(_01050_),
    .B(_01044_),
    .X(_01073_));
 sg13g2_a21oi_1 _09040_ (.A1(_01072_),
    .A2(_01069_),
    .Y(_01074_),
    .B1(_01073_));
 sg13g2_xnor2_1 _09041_ (.Y(_01075_),
    .A(_05017_),
    .B(_00828_));
 sg13g2_xnor2_1 _09042_ (.Y(_01076_),
    .A(_00826_),
    .B(_01075_));
 sg13g2_xnor2_1 _09043_ (.Y(_01077_),
    .A(net33),
    .B(_01076_));
 sg13g2_mux2_1 _09044_ (.A0(_01071_),
    .A1(_01074_),
    .S(_01077_),
    .X(_01078_));
 sg13g2_buf_8 _09045_ (.A(_01078_),
    .X(_01079_));
 sg13g2_inv_1 _09046_ (.Y(_01080_),
    .A(_01079_));
 sg13g2_a21oi_1 _09047_ (.A1(_01028_),
    .A2(_01049_),
    .Y(_01081_),
    .B1(_01080_));
 sg13g2_and2_1 _09048_ (.A(_01079_),
    .B(_01048_),
    .X(_01082_));
 sg13g2_or2_1 _09049_ (.X(_01083_),
    .B(_01048_),
    .A(_01079_));
 sg13g2_o21ai_1 _09050_ (.B1(_01083_),
    .Y(_01084_),
    .A1(_01038_),
    .A2(_01082_));
 sg13g2_o21ai_1 _09051_ (.B1(_00823_),
    .Y(_01085_),
    .A1(_01038_),
    .A2(_01048_));
 sg13g2_a21oi_1 _09052_ (.A1(_01084_),
    .A2(_01085_),
    .Y(_01086_),
    .B1(_01028_));
 sg13g2_a21oi_2 _09053_ (.B1(_01086_),
    .Y(_01087_),
    .A2(_01081_),
    .A1(_00823_));
 sg13g2_nor2_1 _09054_ (.A(_00941_),
    .B(_00951_),
    .Y(_01088_));
 sg13g2_nor2_1 _09055_ (.A(_00931_),
    .B(_01009_),
    .Y(_01089_));
 sg13g2_and2_1 _09056_ (.A(_00931_),
    .B(_00941_),
    .X(_01090_));
 sg13g2_nor2_1 _09057_ (.A(_00931_),
    .B(_00941_),
    .Y(_01091_));
 sg13g2_nor2_1 _09058_ (.A(_01016_),
    .B(_01091_),
    .Y(_01092_));
 sg13g2_a221oi_1 _09059_ (.B2(_01011_),
    .C1(_01092_),
    .B1(_01090_),
    .A1(_01088_),
    .Y(_01093_),
    .A2(_01089_));
 sg13g2_nand2_1 _09060_ (.Y(_01094_),
    .A(_00864_),
    .B(_00866_));
 sg13g2_xnor2_1 _09061_ (.Y(_01095_),
    .A(_01094_),
    .B(_00942_));
 sg13g2_xor2_1 _09062_ (.B(_01095_),
    .A(_01093_),
    .X(_01096_));
 sg13g2_mux2_1 _09063_ (.A0(_00653_),
    .A1(_01087_),
    .S(_01096_),
    .X(_01097_));
 sg13g2_buf_1 _09064_ (.A(_01097_),
    .X(_01098_));
 sg13g2_inv_2 _09065_ (.Y(_01099_),
    .A(_01098_));
 sg13g2_xnor2_1 _09066_ (.Y(_01100_),
    .A(_00859_),
    .B(_00730_));
 sg13g2_xnor2_1 _09067_ (.Y(_01101_),
    .A(_00771_),
    .B(_01100_));
 sg13g2_o21ai_1 _09068_ (.B1(_00869_),
    .Y(_01102_),
    .A1(_00852_),
    .A2(_01101_));
 sg13g2_xnor2_1 _09069_ (.Y(_01103_),
    .A(_00874_),
    .B(_00913_));
 sg13g2_xor2_1 _09070_ (.B(_01103_),
    .A(_01102_),
    .X(_01104_));
 sg13g2_o21ai_1 _09071_ (.B1(_01104_),
    .Y(_01105_),
    .A1(_01023_),
    .A2(_01099_));
 sg13g2_o21ai_1 _09072_ (.B1(_01105_),
    .Y(_01106_),
    .A1(_01024_),
    .A2(_01098_));
 sg13g2_xnor2_1 _09073_ (.Y(_01107_),
    .A(_00941_),
    .B(_00951_));
 sg13g2_a21oi_1 _09074_ (.A1(_01009_),
    .A2(_01107_),
    .Y(_01108_),
    .B1(_00931_));
 sg13g2_nor2_1 _09075_ (.A(_01009_),
    .B(_01107_),
    .Y(_01109_));
 sg13g2_nor4_1 _09076_ (.A(_00943_),
    .B(_00947_),
    .C(_01108_),
    .D(_01109_),
    .Y(_01110_));
 sg13g2_nand2_1 _09077_ (.Y(_01111_),
    .A(_00722_),
    .B(_01088_));
 sg13g2_nor2_1 _09078_ (.A(_00722_),
    .B(_01088_),
    .Y(_01112_));
 sg13g2_nor2_1 _09079_ (.A(_01108_),
    .B(_01109_),
    .Y(_01113_));
 sg13g2_or2_1 _09080_ (.X(_01114_),
    .B(_01113_),
    .A(_01020_));
 sg13g2_inv_1 _09081_ (.Y(_01115_),
    .A(_01087_));
 sg13g2_a221oi_1 _09082_ (.B2(_01114_),
    .C1(_01115_),
    .B1(_01112_),
    .A1(_01110_),
    .Y(_01116_),
    .A2(_01111_));
 sg13g2_nor2_1 _09083_ (.A(_01020_),
    .B(_01113_),
    .Y(_01117_));
 sg13g2_nor3_1 _09084_ (.A(_00943_),
    .B(_00947_),
    .C(_01089_),
    .Y(_01118_));
 sg13g2_o21ai_1 _09085_ (.B1(_01089_),
    .Y(_01119_),
    .A1(_00943_),
    .A2(_00947_));
 sg13g2_o21ai_1 _09086_ (.B1(_01119_),
    .Y(_01120_),
    .A1(_00653_),
    .A2(_01118_));
 sg13g2_a221oi_1 _09087_ (.B2(_01088_),
    .C1(_01087_),
    .B1(_01120_),
    .A1(_00722_),
    .Y(_01121_),
    .A2(_01117_));
 sg13g2_nor2_1 _09088_ (.A(_01111_),
    .B(_01119_),
    .Y(_01122_));
 sg13g2_a21oi_1 _09089_ (.A1(_01110_),
    .A2(_01112_),
    .Y(_01123_),
    .B1(_01122_));
 sg13g2_o21ai_1 _09090_ (.B1(_01123_),
    .Y(_01124_),
    .A1(_01116_),
    .A2(_01121_));
 sg13g2_xnor2_1 _09091_ (.Y(_01125_),
    .A(_01104_),
    .B(_01124_));
 sg13g2_xnor2_1 _09092_ (.Y(_01126_),
    .A(_01093_),
    .B(_01087_));
 sg13g2_xnor2_1 _09093_ (.Y(_01127_),
    .A(_01095_),
    .B(_01126_));
 sg13g2_xnor2_1 _09094_ (.Y(_01128_),
    .A(_00823_),
    .B(_01048_));
 sg13g2_xnor2_1 _09095_ (.Y(_01129_),
    .A(_01079_),
    .B(_01128_));
 sg13g2_xnor2_1 _09096_ (.Y(_01130_),
    .A(_01038_),
    .B(_01129_));
 sg13g2_xnor2_1 _09097_ (.Y(_01131_),
    .A(_00450_),
    .B(_00826_));
 sg13g2_xnor2_1 _09098_ (.Y(_01132_),
    .A(net33),
    .B(_01131_));
 sg13g2_xnor2_1 _09099_ (.Y(_01133_),
    .A(_01072_),
    .B(_01069_));
 sg13g2_xnor2_1 _09100_ (.Y(_01134_),
    .A(_01132_),
    .B(_01133_));
 sg13g2_nand2_1 _09101_ (.Y(_01135_),
    .A(_07506_),
    .B(_00287_));
 sg13g2_xnor2_1 _09102_ (.Y(_01136_),
    .A(_00965_),
    .B(_01040_));
 sg13g2_buf_1 _09103_ (.A(_00003_),
    .X(_01137_));
 sg13g2_nand2_1 _09104_ (.Y(_01138_),
    .A(_04907_),
    .B(_01137_));
 sg13g2_and3_1 _09105_ (.X(_01139_),
    .A(_05017_),
    .B(net265),
    .C(_01138_));
 sg13g2_a21oi_1 _09106_ (.A1(_00282_),
    .A2(_01136_),
    .Y(_01140_),
    .B1(_01139_));
 sg13g2_nand3_1 _09107_ (.B(_04978_),
    .C(_01138_),
    .A(_05008_),
    .Y(_01141_));
 sg13g2_buf_1 _09108_ (.A(_01141_),
    .X(_01142_));
 sg13g2_nand2_1 _09109_ (.Y(_01143_),
    .A(_01142_),
    .B(_01135_));
 sg13g2_inv_1 _09110_ (.Y(_01144_),
    .A(_01136_));
 sg13g2_nand3_1 _09111_ (.B(_01143_),
    .C(_01144_),
    .A(net269),
    .Y(_01145_));
 sg13g2_o21ai_1 _09112_ (.B1(_01145_),
    .Y(_01146_),
    .A1(_01135_),
    .A2(_01140_));
 sg13g2_nor3_1 _09113_ (.A(_00955_),
    .B(_01142_),
    .C(_01144_),
    .Y(_01147_));
 sg13g2_a21o_1 _09114_ (.A2(_01146_),
    .A1(_00429_),
    .B1(_01147_),
    .X(_01148_));
 sg13g2_xor2_1 _09115_ (.B(_05848_),
    .A(_06332_),
    .X(_01149_));
 sg13g2_buf_2 _09116_ (.A(_01149_),
    .X(_01150_));
 sg13g2_buf_1 _09117_ (.A(_01150_),
    .X(_01151_));
 sg13g2_nor2_2 _09118_ (.A(_06629_),
    .B(_06847_),
    .Y(_01152_));
 sg13g2_nand2_1 _09119_ (.Y(_01153_),
    .A(net302),
    .B(_07497_));
 sg13g2_buf_1 _09120_ (.A(_01153_),
    .X(_01154_));
 sg13g2_inv_1 _09121_ (.Y(_01155_),
    .A(_01154_));
 sg13g2_nor2_2 _09122_ (.A(_00532_),
    .B(_07495_),
    .Y(_01156_));
 sg13g2_a21oi_1 _09123_ (.A1(_01152_),
    .A2(_01155_),
    .Y(_01157_),
    .B1(_01156_));
 sg13g2_nand2_1 _09124_ (.Y(_01158_),
    .A(net335),
    .B(_07494_));
 sg13g2_nand2_1 _09125_ (.Y(_01159_),
    .A(_01158_),
    .B(_01154_));
 sg13g2_nand2_1 _09126_ (.Y(_01160_),
    .A(net44),
    .B(_01154_));
 sg13g2_a21oi_1 _09127_ (.A1(_01159_),
    .A2(_01160_),
    .Y(_01161_),
    .B1(_01152_));
 sg13g2_a21oi_1 _09128_ (.A1(net44),
    .A2(_01157_),
    .Y(_01162_),
    .B1(_01161_));
 sg13g2_nor2_1 _09129_ (.A(_01158_),
    .B(_01154_),
    .Y(_01163_));
 sg13g2_or2_1 _09130_ (.X(_01164_),
    .B(_06847_),
    .A(_06629_));
 sg13g2_buf_1 _09131_ (.A(_01164_),
    .X(_01165_));
 sg13g2_nor2_1 _09132_ (.A(_01165_),
    .B(_01151_),
    .Y(_01166_));
 sg13g2_nand2b_1 _09133_ (.Y(_01167_),
    .B(_01166_),
    .A_N(_01163_));
 sg13g2_xor2_1 _09134_ (.B(_01064_),
    .A(_01056_),
    .X(_01168_));
 sg13g2_inv_1 _09135_ (.Y(_01169_),
    .A(_01168_));
 sg13g2_xnor2_1 _09136_ (.Y(_01170_),
    .A(_06343_),
    .B(_01169_));
 sg13g2_xnor2_1 _09137_ (.Y(_01171_),
    .A(_07256_),
    .B(_01170_));
 sg13g2_mux2_1 _09138_ (.A0(_01162_),
    .A1(_01167_),
    .S(_01171_),
    .X(_01172_));
 sg13g2_xnor2_1 _09139_ (.Y(_01173_),
    .A(_01171_),
    .B(_01166_));
 sg13g2_xnor2_1 _09140_ (.Y(_01174_),
    .A(_01152_),
    .B(_01151_));
 sg13g2_o21ai_1 _09141_ (.B1(_01159_),
    .Y(_01175_),
    .A1(_01163_),
    .A2(_01174_));
 sg13g2_o21ai_1 _09142_ (.B1(_01137_),
    .Y(_01176_),
    .A1(_01173_),
    .A2(_01175_));
 sg13g2_nand2_1 _09143_ (.Y(_01177_),
    .A(_01172_),
    .B(_01176_));
 sg13g2_nand3_1 _09144_ (.B(_01060_),
    .C(_01168_),
    .A(net34),
    .Y(_01178_));
 sg13g2_xnor2_1 _09145_ (.Y(_01179_),
    .A(_01142_),
    .B(_01178_));
 sg13g2_xnor2_1 _09146_ (.Y(_01180_),
    .A(_01052_),
    .B(_01179_));
 sg13g2_nand2_1 _09147_ (.Y(_01181_),
    .A(_01177_),
    .B(_01180_));
 sg13g2_xnor2_1 _09148_ (.Y(_01182_),
    .A(_01066_),
    .B(_01139_));
 sg13g2_xnor2_1 _09149_ (.Y(_01183_),
    .A(_01136_),
    .B(_01182_));
 sg13g2_nand2_1 _09150_ (.Y(_01184_),
    .A(_00955_),
    .B(_01183_));
 sg13g2_nand2b_1 _09151_ (.Y(_01185_),
    .B(_00968_),
    .A_N(_01183_));
 sg13g2_a21oi_1 _09152_ (.A1(_01065_),
    .A2(_01062_),
    .Y(_01186_),
    .B1(_01066_));
 sg13g2_xnor2_1 _09153_ (.Y(_01187_),
    .A(_01052_),
    .B(_01136_));
 sg13g2_xnor2_1 _09154_ (.Y(_01188_),
    .A(_01186_),
    .B(_01187_));
 sg13g2_mux2_1 _09155_ (.A0(_01184_),
    .A1(_01185_),
    .S(_01188_),
    .X(_01189_));
 sg13g2_and3_1 _09156_ (.X(_01190_),
    .A(_01148_),
    .B(_01181_),
    .C(_01189_));
 sg13g2_buf_1 _09157_ (.A(_01190_),
    .X(_01191_));
 sg13g2_xnor2_1 _09158_ (.Y(_01192_),
    .A(_00828_),
    .B(_01191_));
 sg13g2_a21oi_1 _09159_ (.A1(_00429_),
    .A2(_01146_),
    .Y(_01193_),
    .B1(_01147_));
 sg13g2_nand2_1 _09160_ (.Y(_01194_),
    .A(_01181_),
    .B(_01189_));
 sg13g2_a21oi_1 _09161_ (.A1(_01193_),
    .A2(_01194_),
    .Y(_01195_),
    .B1(_01134_));
 sg13g2_a21oi_1 _09162_ (.A1(_01134_),
    .A2(_01192_),
    .Y(_01196_),
    .B1(_01195_));
 sg13g2_xor2_1 _09163_ (.B(_01196_),
    .A(_01130_),
    .X(_01197_));
 sg13g2_xnor2_1 _09164_ (.Y(_01198_),
    .A(_01193_),
    .B(_01194_));
 sg13g2_xnor2_1 _09165_ (.Y(_01199_),
    .A(_01134_),
    .B(_01198_));
 sg13g2_xor2_1 _09166_ (.B(_01180_),
    .A(_01177_),
    .X(_01200_));
 sg13g2_xnor2_1 _09167_ (.Y(_01201_),
    .A(net44),
    .B(_01156_));
 sg13g2_buf_1 _09168_ (.A(_06706_),
    .X(_01202_));
 sg13g2_a21oi_1 _09169_ (.A1(net92),
    .A2(net69),
    .Y(_01203_),
    .B1(_06618_));
 sg13g2_and3_1 _09170_ (.X(_01204_),
    .A(_06618_),
    .B(net92),
    .C(net69));
 sg13g2_nor3_1 _09171_ (.A(_06398_),
    .B(_01203_),
    .C(_01204_),
    .Y(_01205_));
 sg13g2_a21o_1 _09172_ (.A2(_01203_),
    .A1(_06398_),
    .B1(_01205_),
    .X(_01206_));
 sg13g2_nand2_1 _09173_ (.Y(_01207_),
    .A(_06398_),
    .B(_06618_));
 sg13g2_nand2_1 _09174_ (.Y(_01208_),
    .A(net92),
    .B(net69));
 sg13g2_nor3_1 _09175_ (.A(_01207_),
    .B(_01208_),
    .C(_01201_),
    .Y(_01209_));
 sg13g2_a21o_1 _09176_ (.A2(_01206_),
    .A1(_01201_),
    .B1(_01209_),
    .X(_01210_));
 sg13g2_nand2_1 _09177_ (.Y(_01211_),
    .A(_04998_),
    .B(_07494_));
 sg13g2_buf_1 _09178_ (.A(_01211_),
    .X(_01212_));
 sg13g2_nand2_1 _09179_ (.Y(_01213_),
    .A(net333),
    .B(net329));
 sg13g2_buf_1 _09180_ (.A(_01213_),
    .X(_01214_));
 sg13g2_nand2_2 _09181_ (.Y(_01215_),
    .A(_01212_),
    .B(_01214_));
 sg13g2_nand3_1 _09182_ (.B(_00932_),
    .C(_07494_),
    .A(net335),
    .Y(_01216_));
 sg13g2_nor2b_1 _09183_ (.A(_01216_),
    .B_N(_01150_),
    .Y(_01217_));
 sg13g2_and2_1 _09184_ (.A(_07495_),
    .B(_01150_),
    .X(_01218_));
 sg13g2_mux2_1 _09185_ (.A0(_01217_),
    .A1(_01218_),
    .S(_01152_),
    .X(_01219_));
 sg13g2_nor2_1 _09186_ (.A(net335),
    .B(net304),
    .Y(_01220_));
 sg13g2_and2_1 _09187_ (.A(_01150_),
    .B(_01220_),
    .X(_01221_));
 sg13g2_nor2_1 _09188_ (.A(net295),
    .B(net44),
    .Y(_01222_));
 sg13g2_mux2_1 _09189_ (.A0(_01221_),
    .A1(_01222_),
    .S(_01165_),
    .X(_01223_));
 sg13g2_nor2b_1 _09190_ (.A(net44),
    .B_N(_01220_),
    .Y(_01224_));
 sg13g2_nor4_1 _09191_ (.A(_06629_),
    .B(_06847_),
    .C(net44),
    .D(_01216_),
    .Y(_01225_));
 sg13g2_a21o_1 _09192_ (.A2(_01224_),
    .A1(_01165_),
    .B1(_01225_),
    .X(_01226_));
 sg13g2_nor4_1 _09193_ (.A(_01154_),
    .B(_01219_),
    .C(_01223_),
    .D(_01226_),
    .Y(_01227_));
 sg13g2_a21o_1 _09194_ (.A2(_01215_),
    .A1(_01210_),
    .B1(_01227_),
    .X(_01228_));
 sg13g2_buf_2 _09195_ (.A(_01228_),
    .X(_01229_));
 sg13g2_nor2_1 _09196_ (.A(_04949_),
    .B(_01168_),
    .Y(_01230_));
 sg13g2_nand2_1 _09197_ (.Y(_01231_),
    .A(_01137_),
    .B(_01159_));
 sg13g2_nand2b_1 _09198_ (.Y(_01232_),
    .B(_01150_),
    .A_N(_01231_));
 sg13g2_nor2_1 _09199_ (.A(_01137_),
    .B(_01163_),
    .Y(_01233_));
 sg13g2_nand2b_1 _09200_ (.Y(_01234_),
    .B(_01233_),
    .A_N(_01150_));
 sg13g2_a21oi_1 _09201_ (.A1(_01232_),
    .A2(_01234_),
    .Y(_01235_),
    .B1(_01165_));
 sg13g2_or2_1 _09202_ (.X(_01236_),
    .B(_01231_),
    .A(_01150_));
 sg13g2_nand2_1 _09203_ (.Y(_01237_),
    .A(_01150_),
    .B(_01233_));
 sg13g2_a21oi_1 _09204_ (.A1(_01236_),
    .A2(_01237_),
    .Y(_01238_),
    .B1(_01152_));
 sg13g2_nand2_1 _09205_ (.Y(_01239_),
    .A(_01137_),
    .B(_01163_));
 sg13g2_o21ai_1 _09206_ (.B1(_01239_),
    .Y(_01240_),
    .A1(_01137_),
    .A2(_01159_));
 sg13g2_nor3_1 _09207_ (.A(_01235_),
    .B(_01238_),
    .C(_01240_),
    .Y(_01241_));
 sg13g2_xnor2_1 _09208_ (.Y(_01242_),
    .A(_01062_),
    .B(_01241_));
 sg13g2_a21oi_1 _09209_ (.A1(_00933_),
    .A2(_01229_),
    .Y(_01243_),
    .B1(_01242_));
 sg13g2_a21oi_2 _09210_ (.B1(_01227_),
    .Y(_01244_),
    .A2(_01215_),
    .A1(_01210_));
 sg13g2_or3_1 _09211_ (.A(_01235_),
    .B(_01238_),
    .C(_01240_),
    .X(_01245_));
 sg13g2_buf_1 _09212_ (.A(_01245_),
    .X(_01246_));
 sg13g2_xnor2_1 _09213_ (.Y(_01247_),
    .A(_01062_),
    .B(_01246_));
 sg13g2_a21oi_1 _09214_ (.A1(_04949_),
    .A2(_01244_),
    .Y(_01248_),
    .B1(_01247_));
 sg13g2_a221oi_1 _09215_ (.B2(_01168_),
    .C1(_01248_),
    .B1(_01243_),
    .A1(_01229_),
    .Y(_01249_),
    .A2(_01230_));
 sg13g2_xnor2_1 _09216_ (.Y(_01250_),
    .A(_01200_),
    .B(_01249_));
 sg13g2_nor2_1 _09217_ (.A(_01212_),
    .B(_01214_),
    .Y(_01251_));
 sg13g2_and2_1 _09218_ (.A(net92),
    .B(_01251_),
    .X(_01252_));
 sg13g2_a22oi_1 _09219_ (.Y(_01253_),
    .B1(_01252_),
    .B2(_06826_),
    .A2(_01251_),
    .A1(_06618_));
 sg13g2_nand4_1 _09220_ (.B(_01202_),
    .C(net69),
    .A(_06618_),
    .Y(_01254_),
    .D(_01215_));
 sg13g2_xnor2_1 _09221_ (.Y(_01255_),
    .A(_05639_),
    .B(_06376_));
 sg13g2_a21o_1 _09222_ (.A2(_01254_),
    .A1(_01253_),
    .B1(_01255_),
    .X(_01256_));
 sg13g2_and2_1 _09223_ (.A(_01212_),
    .B(_01214_),
    .X(_01257_));
 sg13g2_buf_1 _09224_ (.A(_01257_),
    .X(_01258_));
 sg13g2_a22oi_1 _09225_ (.Y(_01259_),
    .B1(_01251_),
    .B2(_01204_),
    .A2(_01258_),
    .A1(_01203_));
 sg13g2_a21oi_1 _09226_ (.A1(_01202_),
    .A2(_06826_),
    .Y(_01260_),
    .B1(_01251_));
 sg13g2_o21ai_1 _09227_ (.B1(_06629_),
    .Y(_01261_),
    .A1(_01258_),
    .A2(_01260_));
 sg13g2_nand3_1 _09228_ (.B(_01208_),
    .C(_01258_),
    .A(_01255_),
    .Y(_01262_));
 sg13g2_nand4_1 _09229_ (.B(_01259_),
    .C(_01261_),
    .A(_01256_),
    .Y(_01263_),
    .D(_01262_));
 sg13g2_xor2_1 _09230_ (.B(_01263_),
    .A(net44),
    .X(_01264_));
 sg13g2_o21ai_1 _09231_ (.B1(net247),
    .Y(_01265_),
    .A1(_01212_),
    .A2(_01214_));
 sg13g2_nand2_1 _09232_ (.Y(_01266_),
    .A(net329),
    .B(_04918_));
 sg13g2_buf_2 _09233_ (.A(_01266_),
    .X(_01267_));
 sg13g2_nand2_1 _09234_ (.Y(_01268_),
    .A(net304),
    .B(_07494_));
 sg13g2_or2_1 _09235_ (.X(_01269_),
    .B(_01268_),
    .A(_01267_));
 sg13g2_nand2b_1 _09236_ (.Y(_01270_),
    .B(_01269_),
    .A_N(net92));
 sg13g2_nand2_1 _09237_ (.Y(_01271_),
    .A(net92),
    .B(_01269_));
 sg13g2_mux2_1 _09238_ (.A0(_01270_),
    .A1(_01271_),
    .S(net69),
    .X(_01272_));
 sg13g2_nand2_1 _09239_ (.Y(_01273_),
    .A(_01267_),
    .B(_01268_));
 sg13g2_and2_1 _09240_ (.A(_01272_),
    .B(_01273_),
    .X(_01274_));
 sg13g2_buf_1 _09241_ (.A(_01274_),
    .X(_01275_));
 sg13g2_xor2_1 _09242_ (.B(_01214_),
    .A(_01212_),
    .X(_01276_));
 sg13g2_xnor2_1 _09243_ (.Y(_01277_),
    .A(_06398_),
    .B(_06618_));
 sg13g2_xnor2_1 _09244_ (.Y(_01278_),
    .A(_01208_),
    .B(_01277_));
 sg13g2_buf_2 _09245_ (.A(_01278_),
    .X(_01279_));
 sg13g2_mux2_1 _09246_ (.A0(_01275_),
    .A1(_01276_),
    .S(_01279_),
    .X(_01280_));
 sg13g2_nor2_1 _09247_ (.A(net247),
    .B(_01276_),
    .Y(_01281_));
 sg13g2_and3_1 _09248_ (.X(_01282_),
    .A(net303),
    .B(_01272_),
    .C(_01273_));
 sg13g2_mux2_1 _09249_ (.A0(_01281_),
    .A1(_01282_),
    .S(_01279_),
    .X(_01283_));
 sg13g2_a221oi_1 _09250_ (.B2(net247),
    .C1(_01283_),
    .B1(_01280_),
    .A1(_01215_),
    .Y(_01284_),
    .A2(_01265_));
 sg13g2_buf_1 _09251_ (.A(_01284_),
    .X(_01285_));
 sg13g2_and2_1 _09252_ (.A(_01264_),
    .B(_01285_),
    .X(_01286_));
 sg13g2_or2_1 _09253_ (.X(_01287_),
    .B(_01276_),
    .A(net247));
 sg13g2_nand3_1 _09254_ (.B(_01272_),
    .C(_01273_),
    .A(net303),
    .Y(_01288_));
 sg13g2_mux2_1 _09255_ (.A0(_01287_),
    .A1(_01288_),
    .S(_01279_),
    .X(_01289_));
 sg13g2_nand3b_1 _09256_ (.B(_01275_),
    .C(net247),
    .Y(_01290_),
    .A_N(_01279_));
 sg13g2_nand2_1 _09257_ (.Y(_01291_),
    .A(_01215_),
    .B(_01265_));
 sg13g2_a21o_1 _09258_ (.A2(_01290_),
    .A1(_01289_),
    .B1(_01291_),
    .X(_01292_));
 sg13g2_buf_1 _09259_ (.A(_01292_),
    .X(_01293_));
 sg13g2_xnor2_1 _09260_ (.Y(_01294_),
    .A(net44),
    .B(_01263_));
 sg13g2_nand3_1 _09261_ (.B(_01293_),
    .C(_01294_),
    .A(_01158_),
    .Y(_01295_));
 sg13g2_nand2b_1 _09262_ (.Y(_01296_),
    .B(_01295_),
    .A_N(_01286_));
 sg13g2_a21o_1 _09263_ (.A2(_01060_),
    .A1(net34),
    .B1(_04949_),
    .X(_01297_));
 sg13g2_nand3_1 _09264_ (.B(_04949_),
    .C(_01060_),
    .A(net34),
    .Y(_01298_));
 sg13g2_a21oi_1 _09265_ (.A1(_01297_),
    .A2(_01298_),
    .Y(_01299_),
    .B1(_01246_));
 sg13g2_a21o_1 _09266_ (.A2(_01060_),
    .A1(net34),
    .B1(_00933_),
    .X(_01300_));
 sg13g2_nand3_1 _09267_ (.B(_00933_),
    .C(_01060_),
    .A(net34),
    .Y(_01301_));
 sg13g2_a21oi_1 _09268_ (.A1(_01300_),
    .A2(_01301_),
    .Y(_01302_),
    .B1(_01241_));
 sg13g2_nor3_1 _09269_ (.A(_01158_),
    .B(_01293_),
    .C(_01264_),
    .Y(_01303_));
 sg13g2_nor4_1 _09270_ (.A(_01229_),
    .B(_01299_),
    .C(_01302_),
    .D(_01303_),
    .Y(_01304_));
 sg13g2_a21o_1 _09271_ (.A2(_01298_),
    .A1(_01297_),
    .B1(_01246_),
    .X(_01305_));
 sg13g2_a21o_1 _09272_ (.A2(_01301_),
    .A1(_01300_),
    .B1(_01241_),
    .X(_01306_));
 sg13g2_nor2_1 _09273_ (.A(_01293_),
    .B(_01264_),
    .Y(_01307_));
 sg13g2_a221oi_1 _09274_ (.B2(_01156_),
    .C1(_01244_),
    .B1(_01307_),
    .A1(_01305_),
    .Y(_01308_),
    .A2(_01306_));
 sg13g2_or3_1 _09275_ (.A(_01296_),
    .B(_01304_),
    .C(_01308_),
    .X(_01309_));
 sg13g2_buf_1 _09276_ (.A(_01309_),
    .X(_01310_));
 sg13g2_nand3_1 _09277_ (.B(_01305_),
    .C(_01306_),
    .A(_01229_),
    .Y(_01311_));
 sg13g2_buf_1 _09278_ (.A(_01311_),
    .X(_01312_));
 sg13g2_o21ai_1 _09279_ (.B1(_01244_),
    .Y(_01313_),
    .A1(_01299_),
    .A2(_01302_));
 sg13g2_buf_1 _09280_ (.A(_01313_),
    .X(_01314_));
 sg13g2_a21oi_1 _09281_ (.A1(_01289_),
    .A2(_01290_),
    .Y(_01315_),
    .B1(_01291_));
 sg13g2_xnor2_1 _09282_ (.Y(_01316_),
    .A(_01156_),
    .B(_01315_));
 sg13g2_a21o_1 _09283_ (.A2(_01316_),
    .A1(_01294_),
    .B1(_01286_),
    .X(_01317_));
 sg13g2_buf_1 _09284_ (.A(_01317_),
    .X(_01318_));
 sg13g2_and3_1 _09285_ (.X(_01319_),
    .A(_01312_),
    .B(_01314_),
    .C(_01318_));
 sg13g2_buf_1 _09286_ (.A(_01319_),
    .X(_01320_));
 sg13g2_a21oi_1 _09287_ (.A1(_01312_),
    .A2(_01314_),
    .Y(_01321_),
    .B1(_01318_));
 sg13g2_o21ai_1 _09288_ (.B1(_01264_),
    .Y(_01322_),
    .A1(_01315_),
    .A2(_01285_));
 sg13g2_or3_1 _09289_ (.A(_01315_),
    .B(_01264_),
    .C(_01285_),
    .X(_01323_));
 sg13g2_buf_1 _09290_ (.A(_01323_),
    .X(_01324_));
 sg13g2_nor2_1 _09291_ (.A(net204),
    .B(_01268_),
    .Y(_01325_));
 sg13g2_xor2_1 _09292_ (.B(net69),
    .A(net92),
    .X(_01326_));
 sg13g2_buf_1 _09293_ (.A(_01326_),
    .X(_01327_));
 sg13g2_buf_1 _09294_ (.A(_06684_),
    .X(_01328_));
 sg13g2_nor2_1 _09295_ (.A(net206),
    .B(_01328_),
    .Y(_01329_));
 sg13g2_buf_1 _09296_ (.A(net207),
    .X(_01330_));
 sg13g2_inv_2 _09297_ (.Y(_01331_),
    .A(net294));
 sg13g2_nor2_1 _09298_ (.A(net155),
    .B(_01331_),
    .Y(_01332_));
 sg13g2_a21oi_1 _09299_ (.A1(_06519_),
    .A2(_01329_),
    .Y(_01333_),
    .B1(_01332_));
 sg13g2_a21o_1 _09300_ (.A2(_06420_),
    .A1(_01330_),
    .B1(_06519_),
    .X(_01334_));
 sg13g2_o21ai_1 _09301_ (.B1(_01334_),
    .Y(_01335_),
    .A1(_06771_),
    .A2(_01333_));
 sg13g2_xnor2_1 _09302_ (.Y(_01336_),
    .A(_06662_),
    .B(_01335_));
 sg13g2_nand2_1 _09303_ (.Y(_01337_),
    .A(_01327_),
    .B(_01336_));
 sg13g2_o21ai_1 _09304_ (.B1(net296),
    .Y(_01338_),
    .A1(_00932_),
    .A2(_01327_));
 sg13g2_nand2_1 _09305_ (.Y(_01339_),
    .A(net295),
    .B(net265));
 sg13g2_a21o_1 _09306_ (.A2(_01338_),
    .A1(_01337_),
    .B1(_01339_),
    .X(_01340_));
 sg13g2_nor2_1 _09307_ (.A(net295),
    .B(net247),
    .Y(_01341_));
 sg13g2_mux2_1 _09308_ (.A0(_01341_),
    .A1(_01336_),
    .S(_01327_),
    .X(_01342_));
 sg13g2_xnor2_1 _09309_ (.Y(_01343_),
    .A(net92),
    .B(net69));
 sg13g2_and4_1 _09310_ (.A(net266),
    .B(net295),
    .C(_01267_),
    .D(_01343_),
    .X(_01344_));
 sg13g2_a21oi_1 _09311_ (.A1(net296),
    .A2(_01342_),
    .Y(_01345_),
    .B1(_01344_));
 sg13g2_xnor2_1 _09312_ (.Y(_01346_),
    .A(_01279_),
    .B(_01275_));
 sg13g2_buf_1 _09313_ (.A(_01346_),
    .X(_01347_));
 sg13g2_a22oi_1 _09314_ (.Y(_01348_),
    .B1(_01347_),
    .B2(net215),
    .A2(_01345_),
    .A1(_01340_));
 sg13g2_or2_1 _09315_ (.X(_01349_),
    .B(_01348_),
    .A(_01325_));
 sg13g2_nand2_1 _09316_ (.Y(_01350_),
    .A(_01340_),
    .B(_01345_));
 sg13g2_nor2_1 _09317_ (.A(net247),
    .B(_01347_),
    .Y(_01351_));
 sg13g2_a21o_1 _09318_ (.A2(_01347_),
    .A1(_01350_),
    .B1(_01351_),
    .X(_01352_));
 sg13g2_and4_1 _09319_ (.A(_01322_),
    .B(_01324_),
    .C(_01349_),
    .D(_01352_),
    .X(_01353_));
 sg13g2_a22oi_1 _09320_ (.Y(_01354_),
    .B1(_01349_),
    .B2(_01352_),
    .A2(_01324_),
    .A1(_01322_));
 sg13g2_xnor2_1 _09321_ (.Y(_01355_),
    .A(net255),
    .B(_05694_));
 sg13g2_nor3_1 _09322_ (.A(_01331_),
    .B(_07495_),
    .C(_06771_),
    .Y(_01356_));
 sg13g2_nand3_1 _09323_ (.B(_01355_),
    .C(_01356_),
    .A(_01336_),
    .Y(_01357_));
 sg13g2_buf_1 _09324_ (.A(_01357_),
    .X(_01358_));
 sg13g2_nor2_1 _09325_ (.A(_01327_),
    .B(_01358_),
    .Y(_01359_));
 sg13g2_nand2_1 _09326_ (.Y(_01360_),
    .A(net204),
    .B(_01339_));
 sg13g2_inv_1 _09327_ (.Y(_01361_),
    .A(_01336_));
 sg13g2_xor2_1 _09328_ (.B(net303),
    .A(net296),
    .X(_01362_));
 sg13g2_nand3_1 _09329_ (.B(_01361_),
    .C(_01362_),
    .A(net251),
    .Y(_01363_));
 sg13g2_o21ai_1 _09330_ (.B1(_01363_),
    .Y(_01364_),
    .A1(_01358_),
    .A2(_01360_));
 sg13g2_a21oi_1 _09331_ (.A1(_01327_),
    .A2(_01358_),
    .Y(_01365_),
    .B1(_07499_));
 sg13g2_nor2_1 _09332_ (.A(_01359_),
    .B(_01365_),
    .Y(_01366_));
 sg13g2_nor2_1 _09333_ (.A(_01339_),
    .B(_01366_),
    .Y(_01367_));
 sg13g2_a221oi_1 _09334_ (.B2(_01327_),
    .C1(_01367_),
    .B1(_01364_),
    .A1(_07506_),
    .Y(_01368_),
    .A2(_01359_));
 sg13g2_buf_1 _09335_ (.A(_01368_),
    .X(_01369_));
 sg13g2_o21ai_1 _09336_ (.B1(net265),
    .Y(_01370_),
    .A1(_07499_),
    .A2(_01268_));
 sg13g2_xnor2_1 _09337_ (.Y(_01371_),
    .A(_01347_),
    .B(_01370_));
 sg13g2_xnor2_1 _09338_ (.Y(_01372_),
    .A(_01350_),
    .B(_01371_));
 sg13g2_nor2_1 _09339_ (.A(_01369_),
    .B(_01372_),
    .Y(_01373_));
 sg13g2_o21ai_1 _09340_ (.B1(_01373_),
    .Y(_01374_),
    .A1(_01353_),
    .A2(_01354_));
 sg13g2_or4_1 _09341_ (.A(_01310_),
    .B(_01320_),
    .C(_01321_),
    .D(_01374_),
    .X(_01375_));
 sg13g2_nor2_1 _09342_ (.A(_01325_),
    .B(_01348_),
    .Y(_01376_));
 sg13g2_a21oi_1 _09343_ (.A1(_01350_),
    .A2(_01347_),
    .Y(_01377_),
    .B1(_01351_));
 sg13g2_nor2_1 _09344_ (.A(_01376_),
    .B(_01377_),
    .Y(_01378_));
 sg13g2_nor2_1 _09345_ (.A(_01373_),
    .B(_01378_),
    .Y(_01379_));
 sg13g2_nor4_1 _09346_ (.A(_01369_),
    .B(_01372_),
    .C(_01376_),
    .D(_01377_),
    .Y(_01380_));
 sg13g2_and2_1 _09347_ (.A(_01322_),
    .B(_01324_),
    .X(_01381_));
 sg13g2_buf_1 _09348_ (.A(_01381_),
    .X(_01382_));
 sg13g2_nor2b_1 _09349_ (.A(_01380_),
    .B_N(_01382_),
    .Y(_01383_));
 sg13g2_or4_1 _09350_ (.A(_01320_),
    .B(_01321_),
    .C(_01379_),
    .D(_01383_),
    .X(_01384_));
 sg13g2_a22oi_1 _09351_ (.Y(_01385_),
    .B1(_01384_),
    .B2(_01310_),
    .A2(_01375_),
    .A1(_01250_));
 sg13g2_buf_1 _09352_ (.A(_01385_),
    .X(_01386_));
 sg13g2_o21ai_1 _09353_ (.B1(_01200_),
    .Y(_01387_),
    .A1(_04949_),
    .A2(_01244_));
 sg13g2_nor2_1 _09354_ (.A(_01169_),
    .B(_01242_),
    .Y(_01388_));
 sg13g2_a21oi_1 _09355_ (.A1(_01244_),
    .A2(_01247_),
    .Y(_01389_),
    .B1(_04949_));
 sg13g2_a21oi_1 _09356_ (.A1(_01229_),
    .A2(_01242_),
    .Y(_01390_),
    .B1(_01389_));
 sg13g2_nor2_1 _09357_ (.A(_01200_),
    .B(_01390_),
    .Y(_01391_));
 sg13g2_a21o_1 _09358_ (.A2(_01388_),
    .A1(_01387_),
    .B1(_01391_),
    .X(_01392_));
 sg13g2_buf_1 _09359_ (.A(_01392_),
    .X(_01393_));
 sg13g2_nor2_1 _09360_ (.A(_01386_),
    .B(_01393_),
    .Y(_01394_));
 sg13g2_nand2_1 _09361_ (.Y(_01395_),
    .A(_01386_),
    .B(_01393_));
 sg13g2_o21ai_1 _09362_ (.B1(_01395_),
    .Y(_01396_),
    .A1(_01199_),
    .A2(_01394_));
 sg13g2_and2_1 _09363_ (.A(_01197_),
    .B(_01396_),
    .X(_01397_));
 sg13g2_buf_1 _09364_ (.A(_01397_),
    .X(_01398_));
 sg13g2_nand2b_1 _09365_ (.Y(_01399_),
    .B(_01134_),
    .A_N(_00828_));
 sg13g2_nor2b_1 _09366_ (.A(_01191_),
    .B_N(_01130_),
    .Y(_01400_));
 sg13g2_nor2_1 _09367_ (.A(_01195_),
    .B(_01191_),
    .Y(_01401_));
 sg13g2_or2_1 _09368_ (.X(_01402_),
    .B(_01401_),
    .A(_01130_));
 sg13g2_o21ai_1 _09369_ (.B1(_01402_),
    .Y(_01403_),
    .A1(_01399_),
    .A2(_01400_));
 sg13g2_buf_1 _09370_ (.A(_01403_),
    .X(_01404_));
 sg13g2_nor2_1 _09371_ (.A(_01398_),
    .B(_01404_),
    .Y(_01405_));
 sg13g2_and2_1 _09372_ (.A(_00823_),
    .B(_01082_),
    .X(_01406_));
 sg13g2_nor2_1 _09373_ (.A(_01038_),
    .B(_01083_),
    .Y(_01407_));
 sg13g2_a221oi_1 _09374_ (.B2(_01038_),
    .C1(_01407_),
    .B1(_01406_),
    .A1(_00820_),
    .Y(_01408_),
    .A2(_01084_));
 sg13g2_xor2_1 _09375_ (.B(_01408_),
    .A(_01028_),
    .X(_01409_));
 sg13g2_nand2_1 _09376_ (.Y(_01410_),
    .A(_01398_),
    .B(_01404_));
 sg13g2_o21ai_1 _09377_ (.B1(_01410_),
    .Y(_01411_),
    .A1(_01405_),
    .A2(_01409_));
 sg13g2_buf_1 _09378_ (.A(_01411_),
    .X(_01412_));
 sg13g2_nand2b_1 _09379_ (.Y(_01413_),
    .B(_01412_),
    .A_N(_01127_));
 sg13g2_xnor2_1 _09380_ (.Y(_01414_),
    .A(_01102_),
    .B(_01103_));
 sg13g2_a21oi_1 _09381_ (.A1(_01015_),
    .A2(_01022_),
    .Y(_01415_),
    .B1(_01414_));
 sg13g2_buf_8 _09382_ (.A(_01415_),
    .X(_01416_));
 sg13g2_a21oi_1 _09383_ (.A1(_00923_),
    .A2(_00925_),
    .Y(_01417_),
    .B1(_01416_));
 sg13g2_and3_1 _09384_ (.X(_01418_),
    .A(_00923_),
    .B(_00925_),
    .C(_01416_));
 sg13g2_nor3_1 _09385_ (.A(_01413_),
    .B(_01417_),
    .C(_01418_),
    .Y(_01419_));
 sg13g2_nand2b_1 _09386_ (.Y(_01420_),
    .B(_00914_),
    .A_N(_00880_));
 sg13g2_buf_2 _09387_ (.A(_01420_),
    .X(_01421_));
 sg13g2_nor2_1 _09388_ (.A(_01421_),
    .B(net22),
    .Y(_01422_));
 sg13g2_nor2b_1 _09389_ (.A(net52),
    .B_N(_00920_),
    .Y(_01423_));
 sg13g2_o21ai_1 _09390_ (.B1(net23),
    .Y(_01424_),
    .A1(_01422_),
    .A2(_01423_));
 sg13g2_xnor2_1 _09391_ (.Y(_01425_),
    .A(_00690_),
    .B(_00716_));
 sg13g2_buf_1 _09392_ (.A(_01425_),
    .X(_01426_));
 sg13g2_a21o_1 _09393_ (.A2(_00918_),
    .A1(_01426_),
    .B1(net52),
    .X(_01427_));
 sg13g2_nand2_1 _09394_ (.Y(_01428_),
    .A(_00717_),
    .B(_00920_));
 sg13g2_a21o_1 _09395_ (.A2(_01428_),
    .A1(_01427_),
    .B1(_00890_),
    .X(_01429_));
 sg13g2_a21oi_1 _09396_ (.A1(_01424_),
    .A2(_01429_),
    .Y(_01430_),
    .B1(_00909_));
 sg13g2_a221oi_1 _09397_ (.B2(_01419_),
    .C1(_01430_),
    .B1(_01125_),
    .A1(_00927_),
    .Y(_01431_),
    .A2(_01106_));
 sg13g2_buf_1 _09398_ (.A(_01431_),
    .X(_01432_));
 sg13g2_nor2_2 _09399_ (.A(_00912_),
    .B(_01432_),
    .Y(_01433_));
 sg13g2_o21ai_1 _09400_ (.B1(_00546_),
    .Y(_01434_),
    .A1(_00523_),
    .A2(_00701_));
 sg13g2_nand2_1 _09401_ (.Y(_01435_),
    .A(_00523_),
    .B(_00700_));
 sg13g2_a21oi_1 _09402_ (.A1(_01434_),
    .A2(_01435_),
    .Y(_01436_),
    .B1(_00703_));
 sg13g2_a221oi_1 _09403_ (.B2(_01433_),
    .C1(_01436_),
    .B1(_00715_),
    .A1(_00523_),
    .Y(_01437_),
    .A2(_00702_));
 sg13g2_inv_1 _09404_ (.Y(_01438_),
    .A(_00347_));
 sg13g2_nor2_2 _09405_ (.A(_00309_),
    .B(_00346_),
    .Y(_01439_));
 sg13g2_nand2b_1 _09406_ (.Y(_01440_),
    .B(_00308_),
    .A_N(_00278_));
 sg13g2_xor2_1 _09407_ (.B(_01440_),
    .A(_00307_),
    .X(_01441_));
 sg13g2_xor2_1 _09408_ (.B(_00262_),
    .A(_00445_),
    .X(_01442_));
 sg13g2_nand2_1 _09409_ (.Y(_01443_),
    .A(_00457_),
    .B(_01442_));
 sg13g2_nand2_1 _09410_ (.Y(_01444_),
    .A(_00448_),
    .B(_01443_));
 sg13g2_o21ai_1 _09411_ (.B1(_01444_),
    .Y(_01445_),
    .A1(_00457_),
    .A2(_01442_));
 sg13g2_a21o_1 _09412_ (.A2(_00249_),
    .A1(_00244_),
    .B1(_00263_),
    .X(_01446_));
 sg13g2_a22oi_1 _09413_ (.Y(_01447_),
    .B1(_01446_),
    .B2(net30),
    .A2(_00263_),
    .A1(_00267_));
 sg13g2_xnor2_1 _09414_ (.Y(_01448_),
    .A(_00270_),
    .B(net68));
 sg13g2_xnor2_1 _09415_ (.Y(_01449_),
    .A(_01447_),
    .B(_01448_));
 sg13g2_nor2_1 _09416_ (.A(_01445_),
    .B(_01449_),
    .Y(_01450_));
 sg13g2_nor2_1 _09417_ (.A(_00459_),
    .B(_00262_),
    .Y(_01451_));
 sg13g2_nand2_1 _09418_ (.Y(_01452_),
    .A(_00459_),
    .B(_00262_));
 sg13g2_nor2_1 _09419_ (.A(_00461_),
    .B(_01452_),
    .Y(_01453_));
 sg13g2_a21oi_1 _09420_ (.A1(_00461_),
    .A2(_01451_),
    .Y(_01454_),
    .B1(_01453_));
 sg13g2_o21ai_1 _09421_ (.B1(_01454_),
    .Y(_01455_),
    .A1(_00444_),
    .A2(_00462_));
 sg13g2_nand2_1 _09422_ (.Y(_01456_),
    .A(_01445_),
    .B(_01449_));
 sg13g2_o21ai_1 _09423_ (.B1(_01456_),
    .Y(_01457_),
    .A1(_01450_),
    .A2(_01455_));
 sg13g2_nor2b_1 _09424_ (.A(_01441_),
    .B_N(_01457_),
    .Y(_01458_));
 sg13g2_nor3_1 _09425_ (.A(_01438_),
    .B(_01439_),
    .C(_01458_),
    .Y(_01459_));
 sg13g2_nor2b_1 _09426_ (.A(_01450_),
    .B_N(_01456_),
    .Y(_01460_));
 sg13g2_xnor2_1 _09427_ (.Y(_01461_),
    .A(_01455_),
    .B(_01460_));
 sg13g2_nor2_1 _09428_ (.A(_00463_),
    .B(_00520_),
    .Y(_01462_));
 sg13g2_nor2_1 _09429_ (.A(_00515_),
    .B(_01462_),
    .Y(_01463_));
 sg13g2_a21oi_1 _09430_ (.A1(_00463_),
    .A2(_00520_),
    .Y(_01464_),
    .B1(_01463_));
 sg13g2_xnor2_1 _09431_ (.Y(_01465_),
    .A(_01461_),
    .B(_01464_));
 sg13g2_buf_2 _09432_ (.A(_01465_),
    .X(_01466_));
 sg13g2_nand2_1 _09433_ (.Y(_01467_),
    .A(_01459_),
    .B(_01466_));
 sg13g2_nor2b_1 _09434_ (.A(_01461_),
    .B_N(_01464_),
    .Y(_01468_));
 sg13g2_buf_2 _09435_ (.A(_01468_),
    .X(_01469_));
 sg13g2_and2_1 _09436_ (.A(_00523_),
    .B(_00712_),
    .X(_01470_));
 sg13g2_buf_1 _09437_ (.A(_01470_),
    .X(_01471_));
 sg13g2_nand2_1 _09438_ (.Y(_01472_),
    .A(_00708_),
    .B(_01471_));
 sg13g2_nand2b_1 _09439_ (.Y(_01473_),
    .B(_01441_),
    .A_N(_01457_));
 sg13g2_buf_1 _09440_ (.A(_01473_),
    .X(_01474_));
 sg13g2_o21ai_1 _09441_ (.B1(_01474_),
    .Y(_01475_),
    .A1(_01438_),
    .A2(_01439_));
 sg13g2_a21oi_1 _09442_ (.A1(_01469_),
    .A2(_01475_),
    .Y(_01476_),
    .B1(_01459_));
 sg13g2_nor2_1 _09443_ (.A(_01472_),
    .B(_01476_),
    .Y(_01477_));
 sg13g2_nor3_1 _09444_ (.A(_01438_),
    .B(_01439_),
    .C(_01474_),
    .Y(_01478_));
 sg13g2_a221oi_1 _09445_ (.B2(_01433_),
    .C1(_01478_),
    .B1(_01477_),
    .A1(_01459_),
    .Y(_01479_),
    .A2(_01469_));
 sg13g2_o21ai_1 _09446_ (.B1(_01479_),
    .Y(_01480_),
    .A1(_01437_),
    .A2(_01467_));
 sg13g2_buf_1 _09447_ (.A(_01480_),
    .X(_01481_));
 sg13g2_a22oi_1 _09448_ (.Y(_01482_),
    .B1(_00413_),
    .B2(_01481_),
    .A2(_00411_),
    .A1(_00390_));
 sg13g2_a21oi_1 _09449_ (.A1(_01481_),
    .A2(_00390_),
    .Y(_01483_),
    .B1(_00412_));
 sg13g2_nand2b_1 _09450_ (.Y(_01484_),
    .B(_00411_),
    .A_N(_01483_));
 sg13g2_o21ai_1 _09451_ (.B1(_01484_),
    .Y(_01485_),
    .A1(_00347_),
    .A2(_01482_));
 sg13g2_buf_1 _09452_ (.A(\i_mandel.i_sq_x.x[1] ),
    .X(_01486_));
 sg13g2_buf_1 _09453_ (.A(_01486_),
    .X(_01487_));
 sg13g2_buf_1 _09454_ (.A(_01487_),
    .X(_01488_));
 sg13g2_buf_1 _09455_ (.A(_01488_),
    .X(_01489_));
 sg13g2_buf_1 _09456_ (.A(net192),
    .X(_01490_));
 sg13g2_buf_1 _09457_ (.A(\i_mandel.i_sq_x.x[-1] ),
    .X(_01491_));
 sg13g2_inv_1 _09458_ (.Y(_01492_),
    .A(net328));
 sg13g2_buf_1 _09459_ (.A(_01492_),
    .X(_01493_));
 sg13g2_buf_8 _09460_ (.A(\i_mandel.i_sq_x.x[2] ),
    .X(_01494_));
 sg13g2_inv_2 _09461_ (.Y(_01495_),
    .A(net327));
 sg13g2_buf_1 _09462_ (.A(_01495_),
    .X(_01496_));
 sg13g2_buf_1 _09463_ (.A(net244),
    .X(_01497_));
 sg13g2_a21oi_1 _09464_ (.A1(net154),
    .A2(net245),
    .Y(_01498_),
    .B1(net191));
 sg13g2_buf_8 _09465_ (.A(\i_mandel.i_sq_x.x[0] ),
    .X(_01499_));
 sg13g2_buf_1 _09466_ (.A(net326),
    .X(_01500_));
 sg13g2_inv_1 _09467_ (.Y(_01501_),
    .A(net292));
 sg13g2_mux2_1 _09468_ (.A0(net154),
    .A1(_01498_),
    .S(_01501_),
    .X(_01502_));
 sg13g2_buf_2 _09469_ (.A(_01502_),
    .X(_01503_));
 sg13g2_buf_8 _09470_ (.A(\i_mandel.i_sq_x.x[-2] ),
    .X(_01504_));
 sg13g2_buf_8 _09471_ (.A(\i_mandel.i_sq_x.x[-3] ),
    .X(_01505_));
 sg13g2_nand2_2 _09472_ (.Y(_01506_),
    .A(_01504_),
    .B(_01505_));
 sg13g2_buf_1 _09473_ (.A(\i_mandel.i_sq_x.x[-4] ),
    .X(_01507_));
 sg13g2_buf_8 _09474_ (.A(\i_mandel.i_sq_x.x[-5] ),
    .X(_01508_));
 sg13g2_buf_8 _09475_ (.A(\i_mandel.i_sq_x.x[-6] ),
    .X(_01509_));
 sg13g2_nand4_1 _09476_ (.B(net324),
    .C(_01509_),
    .A(net325),
    .Y(_01510_),
    .D(net327));
 sg13g2_buf_2 _09477_ (.A(_01510_),
    .X(_01511_));
 sg13g2_buf_8 _09478_ (.A(_01511_),
    .X(_01512_));
 sg13g2_buf_2 _09479_ (.A(_00006_),
    .X(_01513_));
 sg13g2_buf_1 _09480_ (.A(_01513_),
    .X(_01514_));
 sg13g2_buf_1 _09481_ (.A(_00008_),
    .X(_01515_));
 sg13g2_buf_1 _09482_ (.A(_01515_),
    .X(_01516_));
 sg13g2_or2_1 _09483_ (.X(_01517_),
    .B(net290),
    .A(net291));
 sg13g2_o21ai_1 _09484_ (.B1(_01517_),
    .Y(_01518_),
    .A1(_01506_),
    .A2(net190));
 sg13g2_and2_1 _09485_ (.A(_01504_),
    .B(_01505_),
    .X(_01519_));
 sg13g2_buf_1 _09486_ (.A(_01519_),
    .X(_01520_));
 sg13g2_and4_1 _09487_ (.A(net325),
    .B(net324),
    .C(_01509_),
    .D(net327),
    .X(_01521_));
 sg13g2_buf_8 _09488_ (.A(_01521_),
    .X(_01522_));
 sg13g2_buf_8 _09489_ (.A(net243),
    .X(_01523_));
 sg13g2_nand2b_1 _09490_ (.Y(_01524_),
    .B(net290),
    .A_N(net291));
 sg13g2_nand4_1 _09491_ (.B(_01520_),
    .C(net189),
    .A(_01492_),
    .Y(_01525_),
    .D(_01524_));
 sg13g2_buf_1 _09492_ (.A(_00007_),
    .X(_01526_));
 sg13g2_buf_1 _09493_ (.A(_01526_),
    .X(_01527_));
 sg13g2_a21o_1 _09494_ (.A2(_01525_),
    .A1(_01518_),
    .B1(net289),
    .X(_01528_));
 sg13g2_buf_8 _09495_ (.A(_01504_),
    .X(_01529_));
 sg13g2_buf_8 _09496_ (.A(_01505_),
    .X(_01530_));
 sg13g2_nand3_1 _09497_ (.B(_01529_),
    .C(_01530_),
    .A(net328),
    .Y(_01531_));
 sg13g2_buf_1 _09498_ (.A(_01531_),
    .X(_01532_));
 sg13g2_nor2_2 _09499_ (.A(net190),
    .B(_01532_),
    .Y(_01533_));
 sg13g2_nand3_1 _09500_ (.B(net291),
    .C(_01533_),
    .A(net289),
    .Y(_01534_));
 sg13g2_nand2_1 _09501_ (.Y(_01535_),
    .A(_01528_),
    .B(_01534_));
 sg13g2_buf_2 _09502_ (.A(\i_mandel.i_sq_x.x[-11] ),
    .X(_01536_));
 sg13g2_buf_1 _09503_ (.A(_01536_),
    .X(_01537_));
 sg13g2_inv_2 _09504_ (.Y(_01538_),
    .A(_01537_));
 sg13g2_buf_1 _09505_ (.A(\i_mandel.i_sq_x.x[-12] ),
    .X(_01539_));
 sg13g2_buf_1 _09506_ (.A(_01539_),
    .X(_01540_));
 sg13g2_inv_1 _09507_ (.Y(_01541_),
    .A(_01540_));
 sg13g2_buf_1 _09508_ (.A(_01541_),
    .X(_01542_));
 sg13g2_nand4_1 _09509_ (.B(_01491_),
    .C(_01504_),
    .A(net326),
    .Y(_01543_),
    .D(_01505_));
 sg13g2_buf_1 _09510_ (.A(_01543_),
    .X(_01544_));
 sg13g2_buf_1 _09511_ (.A(_00005_),
    .X(_01545_));
 sg13g2_o21ai_1 _09512_ (.B1(_01545_),
    .Y(_01546_),
    .A1(_01544_),
    .A2(_01511_));
 sg13g2_buf_2 _09513_ (.A(_01546_),
    .X(_01547_));
 sg13g2_and4_1 _09514_ (.A(_01499_),
    .B(net328),
    .C(_01504_),
    .D(_01505_),
    .X(_01548_));
 sg13g2_buf_2 _09515_ (.A(_01548_),
    .X(_01549_));
 sg13g2_nand3b_1 _09516_ (.B(_01549_),
    .C(net243),
    .Y(_01550_),
    .A_N(_01545_));
 sg13g2_buf_2 _09517_ (.A(_01550_),
    .X(_01551_));
 sg13g2_nand2_1 _09518_ (.Y(_01552_),
    .A(_01547_),
    .B(_01551_));
 sg13g2_buf_2 _09519_ (.A(_01552_),
    .X(_01553_));
 sg13g2_nor3_1 _09520_ (.A(_01538_),
    .B(net188),
    .C(_01553_),
    .Y(_01554_));
 sg13g2_buf_1 _09521_ (.A(net285),
    .X(_01555_));
 sg13g2_and2_1 _09522_ (.A(_01547_),
    .B(_01551_),
    .X(_01556_));
 sg13g2_buf_1 _09523_ (.A(_01556_),
    .X(_01557_));
 sg13g2_a21oi_1 _09524_ (.A1(_01518_),
    .A2(_01525_),
    .Y(_01558_),
    .B1(net289));
 sg13g2_buf_8 _09525_ (.A(net286),
    .X(_01559_));
 sg13g2_buf_1 _09526_ (.A(_01559_),
    .X(_01560_));
 sg13g2_and4_1 _09527_ (.A(net241),
    .B(net289),
    .C(_01514_),
    .D(_01533_),
    .X(_01561_));
 sg13g2_a221oi_1 _09528_ (.B2(net187),
    .C1(_01561_),
    .B1(_01558_),
    .A1(net242),
    .Y(_01562_),
    .A2(net110));
 sg13g2_buf_1 _09529_ (.A(_01562_),
    .X(_01563_));
 sg13g2_a21oi_1 _09530_ (.A1(_01520_),
    .A2(net243),
    .Y(_01564_),
    .B1(net290));
 sg13g2_nand3_1 _09531_ (.B(net287),
    .C(_01515_),
    .A(_01504_),
    .Y(_01565_));
 sg13g2_buf_1 _09532_ (.A(_01565_),
    .X(_01566_));
 sg13g2_nor3_1 _09533_ (.A(net328),
    .B(_01511_),
    .C(_01566_),
    .Y(_01567_));
 sg13g2_o21ai_1 _09534_ (.B1(net289),
    .Y(_01568_),
    .A1(_01564_),
    .A2(_01567_));
 sg13g2_xor2_1 _09535_ (.B(_01515_),
    .A(_01526_),
    .X(_01569_));
 sg13g2_nand3_1 _09536_ (.B(net241),
    .C(_01569_),
    .A(net328),
    .Y(_01570_));
 sg13g2_nand4_1 _09537_ (.B(net290),
    .C(_01520_),
    .A(_01538_),
    .Y(_01571_),
    .D(net189));
 sg13g2_nor2_1 _09538_ (.A(net286),
    .B(net290),
    .Y(_01572_));
 sg13g2_o21ai_1 _09539_ (.B1(_01572_),
    .Y(_01573_),
    .A1(_01506_),
    .A2(net190));
 sg13g2_and3_1 _09540_ (.X(_01574_),
    .A(_01570_),
    .B(_01571_),
    .C(_01573_));
 sg13g2_a21o_1 _09541_ (.A2(_01574_),
    .A1(_01568_),
    .B1(net291),
    .X(_01575_));
 sg13g2_buf_1 _09542_ (.A(_01575_),
    .X(_01576_));
 sg13g2_inv_2 _09543_ (.Y(_01577_),
    .A(net291));
 sg13g2_nand4_1 _09544_ (.B(_01577_),
    .C(_01547_),
    .A(net242),
    .Y(_01578_),
    .D(_01551_));
 sg13g2_a21oi_1 _09545_ (.A1(_01568_),
    .A2(_01574_),
    .Y(_01579_),
    .B1(_01578_));
 sg13g2_buf_1 _09546_ (.A(_01579_),
    .X(_01580_));
 sg13g2_a221oi_1 _09547_ (.B2(_01576_),
    .C1(_01580_),
    .B1(_01563_),
    .A1(_01535_),
    .Y(_01581_),
    .A2(_01554_));
 sg13g2_buf_2 _09548_ (.A(_01581_),
    .X(_01582_));
 sg13g2_nor2b_1 _09549_ (.A(_01526_),
    .B_N(net285),
    .Y(_01583_));
 sg13g2_o21ai_1 _09550_ (.B1(_01583_),
    .Y(_01584_),
    .A1(net190),
    .A2(_01532_));
 sg13g2_and3_1 _09551_ (.X(_01585_),
    .A(net328),
    .B(_01504_),
    .C(net287));
 sg13g2_buf_1 _09552_ (.A(_01585_),
    .X(_01586_));
 sg13g2_nand4_1 _09553_ (.B(_01526_),
    .C(net189),
    .A(_01540_),
    .Y(_01587_),
    .D(_01586_));
 sg13g2_buf_1 _09554_ (.A(_01587_),
    .X(_01588_));
 sg13g2_nand4_1 _09555_ (.B(net325),
    .C(net324),
    .A(_01530_),
    .Y(_01589_),
    .D(_01509_));
 sg13g2_buf_1 _09556_ (.A(_01589_),
    .X(_01590_));
 sg13g2_buf_2 _09557_ (.A(_00009_),
    .X(_01591_));
 sg13g2_nor2_1 _09558_ (.A(net291),
    .B(_01591_),
    .Y(_01592_));
 sg13g2_o21ai_1 _09559_ (.B1(_01592_),
    .Y(_01593_),
    .A1(_01495_),
    .A2(_01590_));
 sg13g2_buf_1 _09560_ (.A(net327),
    .X(_01594_));
 sg13g2_and4_1 _09561_ (.A(_01505_),
    .B(net325),
    .C(net324),
    .D(_01509_),
    .X(_01595_));
 sg13g2_buf_2 _09562_ (.A(_01595_),
    .X(_01596_));
 sg13g2_nand4_1 _09563_ (.B(_01577_),
    .C(_01591_),
    .A(net284),
    .Y(_01597_),
    .D(_01596_));
 sg13g2_buf_1 _09564_ (.A(_01597_),
    .X(_01598_));
 sg13g2_nand4_1 _09565_ (.B(_01588_),
    .C(_01593_),
    .A(_01584_),
    .Y(_01599_),
    .D(_01598_));
 sg13g2_inv_1 _09566_ (.Y(_01600_),
    .A(_01515_));
 sg13g2_nand3_1 _09567_ (.B(_01520_),
    .C(_01522_),
    .A(_01600_),
    .Y(_01601_));
 sg13g2_buf_2 _09568_ (.A(_01601_),
    .X(_01602_));
 sg13g2_o21ai_1 _09569_ (.B1(net290),
    .Y(_01603_),
    .A1(_01506_),
    .A2(_01511_));
 sg13g2_buf_2 _09570_ (.A(_01603_),
    .X(_01604_));
 sg13g2_and3_1 _09571_ (.X(_01605_),
    .A(_01559_),
    .B(_01602_),
    .C(_01604_));
 sg13g2_buf_1 _09572_ (.A(_01605_),
    .X(_01606_));
 sg13g2_a22oi_1 _09573_ (.Y(_01607_),
    .B1(_01593_),
    .B2(_01598_),
    .A2(_01588_),
    .A1(_01584_));
 sg13g2_a21o_1 _09574_ (.A2(_01606_),
    .A1(_01599_),
    .B1(_01607_),
    .X(_01608_));
 sg13g2_buf_1 _09575_ (.A(_01608_),
    .X(_01609_));
 sg13g2_buf_1 _09576_ (.A(\i_mandel.i_sq_x.x[-13] ),
    .X(_01610_));
 sg13g2_buf_1 _09577_ (.A(_01610_),
    .X(_01611_));
 sg13g2_and4_1 _09578_ (.A(_01486_),
    .B(_01499_),
    .C(net328),
    .D(_01529_),
    .X(_01612_));
 sg13g2_buf_1 _09579_ (.A(_00004_),
    .X(_01613_));
 sg13g2_a21oi_1 _09580_ (.A1(_01596_),
    .A2(_01612_),
    .Y(_01614_),
    .B1(_01613_));
 sg13g2_buf_1 _09581_ (.A(_01614_),
    .X(_01615_));
 sg13g2_and2_1 _09582_ (.A(net283),
    .B(_01615_),
    .X(_01616_));
 sg13g2_buf_1 _09583_ (.A(_01616_),
    .X(_01617_));
 sg13g2_o21ai_1 _09584_ (.B1(_01617_),
    .Y(_01618_),
    .A1(_01582_),
    .A2(net84));
 sg13g2_buf_2 _09585_ (.A(_01618_),
    .X(_01619_));
 sg13g2_buf_8 _09586_ (.A(_01582_),
    .X(_01620_));
 sg13g2_nand2_2 _09587_ (.Y(_01621_),
    .A(net63),
    .B(net84));
 sg13g2_nand4_1 _09588_ (.B(net242),
    .C(_01547_),
    .A(net241),
    .Y(_01622_),
    .D(_01551_));
 sg13g2_a21oi_2 _09589_ (.B1(_01622_),
    .Y(_01623_),
    .A2(_01534_),
    .A1(_01528_));
 sg13g2_buf_1 _09590_ (.A(_01577_),
    .X(_01624_));
 sg13g2_nand2_1 _09591_ (.Y(_01625_),
    .A(net187),
    .B(net186));
 sg13g2_inv_1 _09592_ (.Y(_01626_),
    .A(net289));
 sg13g2_nor2_1 _09593_ (.A(net190),
    .B(_01566_),
    .Y(_01627_));
 sg13g2_buf_1 _09594_ (.A(net328),
    .X(_01628_));
 sg13g2_and2_1 _09595_ (.A(net282),
    .B(net289),
    .X(_01629_));
 sg13g2_nor4_1 _09596_ (.A(net282),
    .B(_01527_),
    .C(net190),
    .D(_01566_),
    .Y(_01630_));
 sg13g2_a221oi_1 _09597_ (.B2(_01629_),
    .C1(_01630_),
    .B1(_01627_),
    .A1(_01626_),
    .Y(_01631_),
    .A2(_01564_));
 sg13g2_nor2_1 _09598_ (.A(_01625_),
    .B(_01631_),
    .Y(_01632_));
 sg13g2_nor3_1 _09599_ (.A(_01580_),
    .B(_01623_),
    .C(_01632_),
    .Y(_01633_));
 sg13g2_buf_2 _09600_ (.A(_01633_),
    .X(_01634_));
 sg13g2_or2_1 _09601_ (.X(_01635_),
    .B(net291),
    .A(_01526_));
 sg13g2_a21o_1 _09602_ (.A2(_01586_),
    .A1(net243),
    .B1(_01635_),
    .X(_01636_));
 sg13g2_nor2b_1 _09603_ (.A(net291),
    .B_N(_01526_),
    .Y(_01637_));
 sg13g2_nand3_1 _09604_ (.B(_01586_),
    .C(_01637_),
    .A(net243),
    .Y(_01638_));
 sg13g2_nand2_1 _09605_ (.Y(_01639_),
    .A(_01549_),
    .B(net189));
 sg13g2_buf_1 _09606_ (.A(_01545_),
    .X(_01640_));
 sg13g2_nor2b_1 _09607_ (.A(net281),
    .B_N(_01536_),
    .Y(_01641_));
 sg13g2_and4_1 _09608_ (.A(net286),
    .B(net281),
    .C(_01549_),
    .D(net189),
    .X(_01642_));
 sg13g2_a221oi_1 _09609_ (.B2(_01641_),
    .C1(_01642_),
    .B1(_01639_),
    .A1(_01636_),
    .Y(_01643_),
    .A2(_01638_));
 sg13g2_buf_1 _09610_ (.A(_01643_),
    .X(_01644_));
 sg13g2_o21ai_1 _09611_ (.B1(_01641_),
    .Y(_01645_),
    .A1(_01544_),
    .A2(net190));
 sg13g2_nand4_1 _09612_ (.B(net281),
    .C(_01549_),
    .A(net286),
    .Y(_01646_),
    .D(net243));
 sg13g2_a21oi_1 _09613_ (.A1(net189),
    .A2(_01586_),
    .Y(_01647_),
    .B1(_01635_));
 sg13g2_a221oi_1 _09614_ (.B2(_01646_),
    .C1(_01647_),
    .B1(_01645_),
    .A1(_01533_),
    .Y(_01648_),
    .A2(_01637_));
 sg13g2_buf_1 _09615_ (.A(_01648_),
    .X(_01649_));
 sg13g2_nor2_1 _09616_ (.A(_01644_),
    .B(_01649_),
    .Y(_01650_));
 sg13g2_xor2_1 _09617_ (.B(_01610_),
    .A(net242),
    .X(_01651_));
 sg13g2_nand2_1 _09618_ (.Y(_01652_),
    .A(_01615_),
    .B(_01651_));
 sg13g2_xnor2_1 _09619_ (.Y(_01653_),
    .A(_01650_),
    .B(_01652_));
 sg13g2_xnor2_1 _09620_ (.Y(_01654_),
    .A(_01634_),
    .B(_01653_));
 sg13g2_a21oi_2 _09621_ (.B1(_01654_),
    .Y(_01655_),
    .A2(_01621_),
    .A1(_01619_));
 sg13g2_and3_1 _09622_ (.X(_01656_),
    .A(_01619_),
    .B(_01621_),
    .C(_01654_));
 sg13g2_buf_2 _09623_ (.A(_01656_),
    .X(_01657_));
 sg13g2_nor2_1 _09624_ (.A(_01655_),
    .B(_01657_),
    .Y(_01658_));
 sg13g2_buf_1 _09625_ (.A(_01658_),
    .X(_01659_));
 sg13g2_nand3_1 _09626_ (.B(_01547_),
    .C(_01551_),
    .A(_01610_),
    .Y(_01660_));
 sg13g2_buf_1 _09627_ (.A(_01660_),
    .X(_01661_));
 sg13g2_buf_2 _09628_ (.A(_00010_),
    .X(_01662_));
 sg13g2_xnor2_1 _09629_ (.Y(_01663_),
    .A(_01662_),
    .B(_01522_));
 sg13g2_buf_8 _09630_ (.A(_01663_),
    .X(_01664_));
 sg13g2_nor2b_1 _09631_ (.A(_01591_),
    .B_N(_01537_),
    .Y(_01665_));
 sg13g2_o21ai_1 _09632_ (.B1(_01665_),
    .Y(_01666_),
    .A1(_01495_),
    .A2(_01590_));
 sg13g2_nand4_1 _09633_ (.B(net284),
    .C(_01591_),
    .A(net241),
    .Y(_01667_),
    .D(_01596_));
 sg13g2_and4_1 _09634_ (.A(net186),
    .B(_01664_),
    .C(_01666_),
    .D(_01667_),
    .X(_01668_));
 sg13g2_a22oi_1 _09635_ (.Y(_01669_),
    .B1(_01666_),
    .B2(_01667_),
    .A2(_01664_),
    .A1(net186));
 sg13g2_and3_1 _09636_ (.X(_01670_),
    .A(net242),
    .B(_01602_),
    .C(_01604_));
 sg13g2_o21ai_1 _09637_ (.B1(_01670_),
    .Y(_01671_),
    .A1(_01668_),
    .A2(_01669_));
 sg13g2_buf_2 _09638_ (.A(_01671_),
    .X(_01672_));
 sg13g2_nor2_1 _09639_ (.A(_01538_),
    .B(_01514_),
    .Y(_01673_));
 sg13g2_inv_1 _09640_ (.Y(_01674_),
    .A(_01591_));
 sg13g2_a21oi_2 _09641_ (.B1(_01674_),
    .Y(_01675_),
    .A2(_01596_),
    .A1(net327));
 sg13g2_nor3_2 _09642_ (.A(_01495_),
    .B(_01591_),
    .C(_01590_),
    .Y(_01676_));
 sg13g2_nor2_1 _09643_ (.A(_01675_),
    .B(_01676_),
    .Y(_01677_));
 sg13g2_buf_1 _09644_ (.A(_01677_),
    .X(_01678_));
 sg13g2_buf_8 _09645_ (.A(_01664_),
    .X(_01679_));
 sg13g2_nand3_1 _09646_ (.B(net108),
    .C(net126),
    .A(_01673_),
    .Y(_01680_));
 sg13g2_buf_1 _09647_ (.A(_01680_),
    .X(_01681_));
 sg13g2_nand3_1 _09648_ (.B(_01672_),
    .C(_01681_),
    .A(_01661_),
    .Y(_01682_));
 sg13g2_and2_1 _09649_ (.A(_01584_),
    .B(_01588_),
    .X(_01683_));
 sg13g2_buf_1 _09650_ (.A(_01683_),
    .X(_01684_));
 sg13g2_nand2_1 _09651_ (.Y(_01685_),
    .A(_01593_),
    .B(_01598_));
 sg13g2_xnor2_1 _09652_ (.Y(_01686_),
    .A(_01685_),
    .B(_01606_));
 sg13g2_buf_2 _09653_ (.A(_01686_),
    .X(_01687_));
 sg13g2_xor2_1 _09654_ (.B(_01687_),
    .A(_01684_),
    .X(_01688_));
 sg13g2_a21oi_1 _09655_ (.A1(_01672_),
    .A2(_01681_),
    .Y(_01689_),
    .B1(_01661_));
 sg13g2_a21o_1 _09656_ (.A2(_01688_),
    .A1(_01682_),
    .B1(_01689_),
    .X(_01690_));
 sg13g2_buf_1 _09657_ (.A(_01690_),
    .X(_01691_));
 sg13g2_nand2_2 _09658_ (.Y(_01692_),
    .A(net283),
    .B(_01615_));
 sg13g2_xnor2_1 _09659_ (.Y(_01693_),
    .A(_01692_),
    .B(net84));
 sg13g2_xor2_1 _09660_ (.B(_01693_),
    .A(_01582_),
    .X(_01694_));
 sg13g2_buf_2 _09661_ (.A(_01694_),
    .X(_01695_));
 sg13g2_nor2_2 _09662_ (.A(net62),
    .B(_01695_),
    .Y(_01696_));
 sg13g2_nand2b_1 _09663_ (.Y(_01697_),
    .B(net109),
    .A_N(net91));
 sg13g2_nand2_1 _09664_ (.Y(_01698_),
    .A(net91),
    .B(net109));
 sg13g2_mux2_1 _09665_ (.A0(_01697_),
    .A1(_01698_),
    .S(_01687_),
    .X(_01699_));
 sg13g2_buf_1 _09666_ (.A(_01699_),
    .X(_01700_));
 sg13g2_nand2b_1 _09667_ (.Y(_01701_),
    .B(net91),
    .A_N(net109));
 sg13g2_or2_1 _09668_ (.X(_01702_),
    .B(net109),
    .A(net91));
 sg13g2_mux2_1 _09669_ (.A0(_01701_),
    .A1(_01702_),
    .S(_01687_),
    .X(_01703_));
 sg13g2_buf_1 _09670_ (.A(_01703_),
    .X(_01704_));
 sg13g2_and2_1 _09671_ (.A(_01672_),
    .B(_01681_),
    .X(_01705_));
 sg13g2_buf_1 _09672_ (.A(_01705_),
    .X(_01706_));
 sg13g2_a21oi_2 _09673_ (.B1(_01706_),
    .Y(_01707_),
    .A2(_01704_),
    .A1(_01700_));
 sg13g2_nand2_1 _09674_ (.Y(_01708_),
    .A(_01672_),
    .B(_01681_));
 sg13g2_nor2b_1 _09675_ (.A(net91),
    .B_N(net109),
    .Y(_01709_));
 sg13g2_and2_1 _09676_ (.A(net91),
    .B(net109),
    .X(_01710_));
 sg13g2_mux2_1 _09677_ (.A0(_01709_),
    .A1(_01710_),
    .S(_01687_),
    .X(_01711_));
 sg13g2_buf_1 _09678_ (.A(_01711_),
    .X(_01712_));
 sg13g2_nor2b_1 _09679_ (.A(net109),
    .B_N(net91),
    .Y(_01713_));
 sg13g2_nor2_1 _09680_ (.A(net91),
    .B(net109),
    .Y(_01714_));
 sg13g2_mux2_1 _09681_ (.A0(_01713_),
    .A1(_01714_),
    .S(_01687_),
    .X(_01715_));
 sg13g2_buf_1 _09682_ (.A(_01715_),
    .X(_01716_));
 sg13g2_nor3_2 _09683_ (.A(_01708_),
    .B(_01712_),
    .C(_01716_),
    .Y(_01717_));
 sg13g2_or3_1 _09684_ (.A(_01668_),
    .B(_01669_),
    .C(_01670_),
    .X(_01718_));
 sg13g2_nand2_1 _09685_ (.Y(_01719_),
    .A(_01672_),
    .B(_01718_));
 sg13g2_buf_2 _09686_ (.A(_01719_),
    .X(_01720_));
 sg13g2_xnor2_1 _09687_ (.Y(_01721_),
    .A(net289),
    .B(_01533_));
 sg13g2_nand2_1 _09688_ (.Y(_01722_),
    .A(net283),
    .B(_01721_));
 sg13g2_or3_1 _09689_ (.A(_01542_),
    .B(_01675_),
    .C(_01676_),
    .X(_01723_));
 sg13g2_buf_2 _09690_ (.A(_01723_),
    .X(_01724_));
 sg13g2_buf_2 _09691_ (.A(_00011_),
    .X(_01725_));
 sg13g2_nor2b_1 _09692_ (.A(_01507_),
    .B_N(net327),
    .Y(_01726_));
 sg13g2_buf_2 _09693_ (.A(_01726_),
    .X(_01727_));
 sg13g2_nand2_1 _09694_ (.Y(_01728_),
    .A(net324),
    .B(_01509_));
 sg13g2_buf_2 _09695_ (.A(_01728_),
    .X(_01729_));
 sg13g2_a221oi_1 _09696_ (.B2(_01729_),
    .C1(net243),
    .B1(_01727_),
    .A1(_01495_),
    .Y(_01730_),
    .A2(_01725_));
 sg13g2_buf_2 _09697_ (.A(_01730_),
    .X(_01731_));
 sg13g2_buf_8 _09698_ (.A(_01731_),
    .X(_01732_));
 sg13g2_nand4_1 _09699_ (.B(net186),
    .C(_01664_),
    .A(net187),
    .Y(_01733_),
    .D(net125));
 sg13g2_a22oi_1 _09700_ (.Y(_01734_),
    .B1(net125),
    .B2(net186),
    .A2(net126),
    .A1(net187));
 sg13g2_a21oi_2 _09701_ (.B1(_01734_),
    .Y(_01735_),
    .A2(_01733_),
    .A1(_01724_));
 sg13g2_nand2b_1 _09702_ (.Y(_01736_),
    .B(_01735_),
    .A_N(_01722_));
 sg13g2_buf_8 _09703_ (.A(_01721_),
    .X(_01737_));
 sg13g2_a21oi_2 _09704_ (.B1(_01735_),
    .Y(_01738_),
    .A2(_01737_),
    .A1(net283));
 sg13g2_a21oi_2 _09705_ (.B1(_01738_),
    .Y(_01739_),
    .A2(_01736_),
    .A1(_01720_));
 sg13g2_o21ai_1 _09706_ (.B1(_01739_),
    .Y(_01740_),
    .A1(_01707_),
    .A2(_01717_));
 sg13g2_buf_2 _09707_ (.A(_01740_),
    .X(_01741_));
 sg13g2_nand2_2 _09708_ (.Y(_01742_),
    .A(net62),
    .B(_01695_));
 sg13g2_o21ai_1 _09709_ (.B1(_01742_),
    .Y(_01743_),
    .A1(_01696_),
    .A2(_01741_));
 sg13g2_buf_1 _09710_ (.A(_01743_),
    .X(_01744_));
 sg13g2_nor3_2 _09711_ (.A(_01696_),
    .B(_01655_),
    .C(_01657_),
    .Y(_01745_));
 sg13g2_nand2b_1 _09712_ (.Y(_01746_),
    .B(net286),
    .A_N(_01662_));
 sg13g2_nand2_1 _09713_ (.Y(_01747_),
    .A(net241),
    .B(_01662_));
 sg13g2_mux2_1 _09714_ (.A0(_01746_),
    .A1(_01747_),
    .S(_01523_),
    .X(_01748_));
 sg13g2_a21o_1 _09715_ (.A2(_01732_),
    .A1(_01624_),
    .B1(_01748_),
    .X(_01749_));
 sg13g2_buf_1 _09716_ (.A(_01749_),
    .X(_01750_));
 sg13g2_nand3_1 _09717_ (.B(_01748_),
    .C(_01732_),
    .A(_01624_),
    .Y(_01751_));
 sg13g2_buf_1 _09718_ (.A(_01751_),
    .X(_01752_));
 sg13g2_nand2_1 _09719_ (.Y(_01753_),
    .A(_01750_),
    .B(_01752_));
 sg13g2_xor2_1 _09720_ (.B(_01753_),
    .A(_01724_),
    .X(_01754_));
 sg13g2_nand3_1 _09721_ (.B(_01602_),
    .C(_01604_),
    .A(net283),
    .Y(_01755_));
 sg13g2_buf_1 _09722_ (.A(_01755_),
    .X(_01756_));
 sg13g2_xnor2_1 _09723_ (.Y(_01757_),
    .A(_01508_),
    .B(_01509_));
 sg13g2_buf_2 _09724_ (.A(_00012_),
    .X(_01758_));
 sg13g2_nor2b_1 _09725_ (.A(net327),
    .B_N(_01758_),
    .Y(_01759_));
 sg13g2_a21oi_1 _09726_ (.A1(net327),
    .A2(_01757_),
    .Y(_01760_),
    .B1(_01759_));
 sg13g2_buf_1 _09727_ (.A(_01760_),
    .X(_01761_));
 sg13g2_a22oi_1 _09728_ (.Y(_01762_),
    .B1(_01761_),
    .B2(net186),
    .A2(_01664_),
    .A1(_01555_));
 sg13g2_nand2_1 _09729_ (.Y(_01763_),
    .A(net241),
    .B(_01731_));
 sg13g2_buf_1 _09730_ (.A(_01555_),
    .X(_01764_));
 sg13g2_nand4_1 _09731_ (.B(net186),
    .C(_01664_),
    .A(net184),
    .Y(_01765_),
    .D(_01761_));
 sg13g2_o21ai_1 _09732_ (.B1(_01765_),
    .Y(_01766_),
    .A1(_01762_),
    .A2(_01763_));
 sg13g2_xor2_1 _09733_ (.B(_01766_),
    .A(_01756_),
    .X(_01767_));
 sg13g2_xnor2_1 _09734_ (.Y(_01768_),
    .A(_01754_),
    .B(_01767_));
 sg13g2_nand2b_1 _09735_ (.Y(_01769_),
    .B(_01539_),
    .A_N(_01662_));
 sg13g2_nand2_1 _09736_ (.Y(_01770_),
    .A(_01539_),
    .B(_01662_));
 sg13g2_mux2_1 _09737_ (.A0(_01769_),
    .A1(_01770_),
    .S(net243),
    .X(_01771_));
 sg13g2_a21o_1 _09738_ (.A2(_01760_),
    .A1(_01577_),
    .B1(_01771_),
    .X(_01772_));
 sg13g2_nand3_1 _09739_ (.B(_01771_),
    .C(net185),
    .A(_01577_),
    .Y(_01773_));
 sg13g2_and3_1 _09740_ (.X(_01774_),
    .A(_01763_),
    .B(_01772_),
    .C(_01773_));
 sg13g2_buf_1 _09741_ (.A(_01774_),
    .X(_01775_));
 sg13g2_a21oi_1 _09742_ (.A1(_01772_),
    .A2(_01773_),
    .Y(_01776_),
    .B1(_01763_));
 sg13g2_or2_1 _09743_ (.X(_01777_),
    .B(_01776_),
    .A(_01775_));
 sg13g2_buf_1 _09744_ (.A(_01777_),
    .X(_01778_));
 sg13g2_buf_1 _09745_ (.A(_01509_),
    .X(_01779_));
 sg13g2_nand2b_1 _09746_ (.Y(_01780_),
    .B(net280),
    .A_N(_01494_));
 sg13g2_nand3b_1 _09747_ (.B(_01494_),
    .C(net324),
    .Y(_01781_),
    .A_N(_01509_));
 sg13g2_o21ai_1 _09748_ (.B1(_01781_),
    .Y(_01782_),
    .A1(_01758_),
    .A2(_01780_));
 sg13g2_buf_1 _09749_ (.A(_01782_),
    .X(_01783_));
 sg13g2_nand2_1 _09750_ (.Y(_01784_),
    .A(_01673_),
    .B(_01783_));
 sg13g2_nand3_1 _09751_ (.B(_01536_),
    .C(_01513_),
    .A(net324),
    .Y(_01785_));
 sg13g2_or2_1 _09752_ (.X(_01786_),
    .B(_01513_),
    .A(_01536_));
 sg13g2_a21oi_1 _09753_ (.A1(_01785_),
    .A2(_01786_),
    .Y(_01787_),
    .B1(net280));
 sg13g2_nand2_1 _09754_ (.Y(_01788_),
    .A(net280),
    .B(_01536_));
 sg13g2_or2_1 _09755_ (.X(_01789_),
    .B(_01513_),
    .A(net280));
 sg13g2_buf_1 _09756_ (.A(net324),
    .X(_01790_));
 sg13g2_a21oi_1 _09757_ (.A1(_01788_),
    .A2(_01789_),
    .Y(_01791_),
    .B1(_01790_));
 sg13g2_or3_1 _09758_ (.A(_01495_),
    .B(_01787_),
    .C(_01791_),
    .X(_01792_));
 sg13g2_nor2b_1 _09759_ (.A(_01513_),
    .B_N(_01779_),
    .Y(_01793_));
 sg13g2_nor2b_1 _09760_ (.A(_01758_),
    .B_N(_01536_),
    .Y(_01794_));
 sg13g2_xnor2_1 _09761_ (.Y(_01795_),
    .A(_01793_),
    .B(_01794_));
 sg13g2_nand2_1 _09762_ (.Y(_01796_),
    .A(net244),
    .B(_01795_));
 sg13g2_nand4_1 _09763_ (.B(net125),
    .C(_01792_),
    .A(net242),
    .Y(_01797_),
    .D(_01796_));
 sg13g2_buf_1 _09764_ (.A(_01797_),
    .X(_01798_));
 sg13g2_nand2_1 _09765_ (.Y(_01799_),
    .A(net283),
    .B(net108));
 sg13g2_a21o_1 _09766_ (.A2(_01798_),
    .A1(_01784_),
    .B1(_01799_),
    .X(_01800_));
 sg13g2_buf_1 _09767_ (.A(_01800_),
    .X(_01801_));
 sg13g2_and3_1 _09768_ (.X(_01802_),
    .A(_01784_),
    .B(_01798_),
    .C(_01799_));
 sg13g2_a21o_1 _09769_ (.A2(_01801_),
    .A1(_01778_),
    .B1(_01802_),
    .X(_01803_));
 sg13g2_buf_1 _09770_ (.A(_01803_),
    .X(_01804_));
 sg13g2_nand2_1 _09771_ (.Y(_01805_),
    .A(_01768_),
    .B(_01804_));
 sg13g2_buf_2 _09772_ (.A(_01805_),
    .X(_01806_));
 sg13g2_nor2_1 _09773_ (.A(_01787_),
    .B(_01791_),
    .Y(_01807_));
 sg13g2_and2_1 _09774_ (.A(_01727_),
    .B(_01729_),
    .X(_01808_));
 sg13g2_nor4_1 _09775_ (.A(net188),
    .B(_01495_),
    .C(net189),
    .D(_01808_),
    .Y(_01809_));
 sg13g2_a22oi_1 _09776_ (.Y(_01810_),
    .B1(_01795_),
    .B2(net244),
    .A2(net125),
    .A1(net285));
 sg13g2_and4_1 _09777_ (.A(net285),
    .B(net244),
    .C(_01731_),
    .D(_01795_),
    .X(_01811_));
 sg13g2_a221oi_1 _09778_ (.B2(_01792_),
    .C1(_01811_),
    .B1(_01810_),
    .A1(_01807_),
    .Y(_01812_),
    .A2(_01809_));
 sg13g2_buf_2 _09779_ (.A(_01812_),
    .X(_01813_));
 sg13g2_nand3_1 _09780_ (.B(net242),
    .C(_01783_),
    .A(net241),
    .Y(_01814_));
 sg13g2_buf_2 _09781_ (.A(_01814_),
    .X(_01815_));
 sg13g2_nand2_1 _09782_ (.Y(_01816_),
    .A(_01610_),
    .B(_01664_));
 sg13g2_xor2_1 _09783_ (.B(_01816_),
    .A(_01815_),
    .X(_01817_));
 sg13g2_xnor2_1 _09784_ (.Y(_01818_),
    .A(_01813_),
    .B(_01817_));
 sg13g2_buf_2 _09785_ (.A(_01818_),
    .X(_01819_));
 sg13g2_nand3b_1 _09786_ (.B(net285),
    .C(_01790_),
    .Y(_01820_),
    .A_N(net286));
 sg13g2_nand2b_1 _09787_ (.Y(_01821_),
    .B(net286),
    .A_N(net285));
 sg13g2_a21o_1 _09788_ (.A2(_01821_),
    .A1(_01820_),
    .B1(net280),
    .X(_01822_));
 sg13g2_inv_2 _09789_ (.Y(_01823_),
    .A(net279));
 sg13g2_mux2_1 _09790_ (.A0(net286),
    .A1(net285),
    .S(net280),
    .X(_01824_));
 sg13g2_a21oi_1 _09791_ (.A1(_01823_),
    .A2(_01824_),
    .Y(_01825_),
    .B1(_01495_));
 sg13g2_nand2b_1 _09792_ (.Y(_01826_),
    .B(net285),
    .A_N(_01758_));
 sg13g2_xnor2_1 _09793_ (.Y(_01827_),
    .A(_01788_),
    .B(_01826_));
 sg13g2_a22oi_1 _09794_ (.Y(_01828_),
    .B1(_01827_),
    .B2(_01496_),
    .A2(_01825_),
    .A1(_01822_));
 sg13g2_buf_1 _09795_ (.A(_01828_),
    .X(_01829_));
 sg13g2_and2_1 _09796_ (.A(net242),
    .B(_01783_),
    .X(_01830_));
 sg13g2_o21ai_1 _09797_ (.B1(_01830_),
    .Y(_01831_),
    .A1(net125),
    .A2(_01829_));
 sg13g2_nand2_1 _09798_ (.Y(_01832_),
    .A(net125),
    .B(_01829_));
 sg13g2_inv_1 _09799_ (.Y(_01833_),
    .A(net283));
 sg13g2_a21oi_1 _09800_ (.A1(_01831_),
    .A2(_01832_),
    .Y(_01834_),
    .B1(net240));
 sg13g2_buf_1 _09801_ (.A(_01834_),
    .X(_01835_));
 sg13g2_nand2_1 _09802_ (.Y(_01836_),
    .A(_01819_),
    .B(_01835_));
 sg13g2_or2_1 _09803_ (.X(_01837_),
    .B(_01815_),
    .A(_01813_));
 sg13g2_buf_1 _09804_ (.A(_01837_),
    .X(_01838_));
 sg13g2_a21o_1 _09805_ (.A2(_01815_),
    .A1(_01813_),
    .B1(_01816_),
    .X(_01839_));
 sg13g2_buf_1 _09806_ (.A(_01839_),
    .X(_01840_));
 sg13g2_nand3_1 _09807_ (.B(_01838_),
    .C(_01840_),
    .A(_01836_),
    .Y(_01841_));
 sg13g2_buf_1 _09808_ (.A(_01841_),
    .X(_01842_));
 sg13g2_nand2_1 _09809_ (.Y(_01843_),
    .A(_01813_),
    .B(_01815_));
 sg13g2_o21ai_1 _09810_ (.B1(_01816_),
    .Y(_01844_),
    .A1(_01813_),
    .A2(_01815_));
 sg13g2_and4_1 _09811_ (.A(_01819_),
    .B(_01835_),
    .C(_01843_),
    .D(_01844_),
    .X(_01845_));
 sg13g2_nand3_1 _09812_ (.B(_01798_),
    .C(_01799_),
    .A(_01784_),
    .Y(_01846_));
 sg13g2_and3_1 _09813_ (.X(_01847_),
    .A(_01778_),
    .B(_01801_),
    .C(_01846_));
 sg13g2_a21oi_1 _09814_ (.A1(_01801_),
    .A2(_01846_),
    .Y(_01848_),
    .B1(_01778_));
 sg13g2_or3_1 _09815_ (.A(_01845_),
    .B(_01847_),
    .C(_01848_),
    .X(_01849_));
 sg13g2_buf_2 _09816_ (.A(_01849_),
    .X(_01850_));
 sg13g2_nand3_1 _09817_ (.B(_01842_),
    .C(_01850_),
    .A(_01806_),
    .Y(_01851_));
 sg13g2_buf_2 _09818_ (.A(_01851_),
    .X(_01852_));
 sg13g2_and2_1 _09819_ (.A(_01602_),
    .B(_01604_),
    .X(_01853_));
 sg13g2_buf_1 _09820_ (.A(_01853_),
    .X(_01854_));
 sg13g2_a221oi_1 _09821_ (.B2(_01752_),
    .C1(_01724_),
    .B1(_01750_),
    .A1(net283),
    .Y(_01855_),
    .A2(_01854_));
 sg13g2_nand4_1 _09822_ (.B(_01756_),
    .C(_01750_),
    .A(_01724_),
    .Y(_01856_),
    .D(_01752_));
 sg13g2_nand3b_1 _09823_ (.B(_01856_),
    .C(_01766_),
    .Y(_01857_),
    .A_N(_01855_));
 sg13g2_o21ai_1 _09824_ (.B1(_01857_),
    .Y(_01858_),
    .A1(_01756_),
    .A2(_01754_));
 sg13g2_buf_1 _09825_ (.A(_01858_),
    .X(_01859_));
 sg13g2_xnor2_1 _09826_ (.Y(_01860_),
    .A(_01722_),
    .B(_01735_));
 sg13g2_xnor2_1 _09827_ (.Y(_01861_),
    .A(_01720_),
    .B(_01860_));
 sg13g2_buf_1 _09828_ (.A(_01861_),
    .X(_01862_));
 sg13g2_and2_1 _09829_ (.A(_01859_),
    .B(_01862_),
    .X(_01863_));
 sg13g2_buf_2 _09830_ (.A(_01863_),
    .X(_01864_));
 sg13g2_nor2_1 _09831_ (.A(_01768_),
    .B(_01804_),
    .Y(_01865_));
 sg13g2_buf_2 _09832_ (.A(_01865_),
    .X(_01866_));
 sg13g2_nor2_1 _09833_ (.A(_01864_),
    .B(_01866_),
    .Y(_01867_));
 sg13g2_nand3_1 _09834_ (.B(_01700_),
    .C(_01704_),
    .A(_01708_),
    .Y(_01868_));
 sg13g2_buf_1 _09835_ (.A(_01868_),
    .X(_01869_));
 sg13g2_o21ai_1 _09836_ (.B1(_01706_),
    .Y(_01870_),
    .A1(_01712_),
    .A2(_01716_));
 sg13g2_buf_1 _09837_ (.A(_01859_),
    .X(_01871_));
 sg13g2_nor2_1 _09838_ (.A(_01738_),
    .B(_01720_),
    .Y(_01872_));
 sg13g2_a22oi_1 _09839_ (.Y(_01873_),
    .B1(net51),
    .B2(_01872_),
    .A2(_01870_),
    .A1(_01869_));
 sg13g2_inv_1 _09840_ (.Y(_01874_),
    .A(_01720_));
 sg13g2_inv_1 _09841_ (.Y(_01875_),
    .A(_01736_));
 sg13g2_o21ai_1 _09842_ (.B1(_01875_),
    .Y(_01876_),
    .A1(_01874_),
    .A2(net51));
 sg13g2_o21ai_1 _09843_ (.B1(_01708_),
    .Y(_01877_),
    .A1(_01712_),
    .A2(_01716_));
 sg13g2_buf_1 _09844_ (.A(_01877_),
    .X(_01878_));
 sg13g2_nand3_1 _09845_ (.B(_01700_),
    .C(_01704_),
    .A(_01706_),
    .Y(_01879_));
 sg13g2_buf_1 _09846_ (.A(_01879_),
    .X(_01880_));
 sg13g2_mux2_1 _09847_ (.A0(_01738_),
    .A1(_01860_),
    .S(_01720_),
    .X(_01881_));
 sg13g2_a221oi_1 _09848_ (.B2(_01859_),
    .C1(_01881_),
    .B1(_01738_),
    .A1(_01878_),
    .Y(_01882_),
    .A2(_01880_));
 sg13g2_a21o_1 _09849_ (.A2(_01876_),
    .A1(_01873_),
    .B1(_01882_),
    .X(_01883_));
 sg13g2_a21oi_1 _09850_ (.A1(_01852_),
    .A2(_01867_),
    .Y(_01884_),
    .B1(_01883_));
 sg13g2_buf_2 _09851_ (.A(_01884_),
    .X(_01885_));
 sg13g2_and2_1 _09852_ (.A(net184),
    .B(_01615_),
    .X(_01886_));
 sg13g2_buf_1 _09853_ (.A(_01886_),
    .X(_01887_));
 sg13g2_o21ai_1 _09854_ (.B1(_01887_),
    .Y(_01888_),
    .A1(_01644_),
    .A2(_01649_));
 sg13g2_buf_1 _09855_ (.A(_01888_),
    .X(_01889_));
 sg13g2_or3_1 _09856_ (.A(_01644_),
    .B(_01649_),
    .C(_01887_),
    .X(_01890_));
 sg13g2_buf_1 _09857_ (.A(_01890_),
    .X(_01891_));
 sg13g2_nand2_1 _09858_ (.Y(_01892_),
    .A(_01889_),
    .B(_01891_));
 sg13g2_a21oi_1 _09859_ (.A1(_01692_),
    .A2(_01634_),
    .Y(_01893_),
    .B1(_01892_));
 sg13g2_nand3_1 _09860_ (.B(net63),
    .C(net84),
    .A(_01634_),
    .Y(_01894_));
 sg13g2_a21oi_1 _09861_ (.A1(_01619_),
    .A2(_01894_),
    .Y(_01895_),
    .B1(_01653_));
 sg13g2_nand3_1 _09862_ (.B(_01620_),
    .C(_01609_),
    .A(_01653_),
    .Y(_01896_));
 sg13g2_a21oi_1 _09863_ (.A1(_01692_),
    .A2(_01896_),
    .Y(_01897_),
    .B1(_01634_));
 sg13g2_or3_1 _09864_ (.A(_01893_),
    .B(_01895_),
    .C(_01897_),
    .X(_01898_));
 sg13g2_and2_1 _09865_ (.A(_01889_),
    .B(_01891_),
    .X(_01899_));
 sg13g2_or3_1 _09866_ (.A(_01580_),
    .B(_01623_),
    .C(_01632_),
    .X(_01900_));
 sg13g2_buf_1 _09867_ (.A(_01900_),
    .X(_01901_));
 sg13g2_nand2_1 _09868_ (.Y(_01902_),
    .A(_01899_),
    .B(_01901_));
 sg13g2_nand4_1 _09869_ (.B(net186),
    .C(_01721_),
    .A(net187),
    .Y(_01903_),
    .D(net110));
 sg13g2_nand2_1 _09870_ (.Y(_01904_),
    .A(net184),
    .B(_01615_));
 sg13g2_nand4_1 _09871_ (.B(_01638_),
    .C(_01645_),
    .A(_01636_),
    .Y(_01905_),
    .D(_01646_));
 sg13g2_or2_1 _09872_ (.X(_01906_),
    .B(_01905_),
    .A(_01904_));
 sg13g2_o21ai_1 _09873_ (.B1(_01906_),
    .Y(_01907_),
    .A1(_01887_),
    .A2(_01903_));
 sg13g2_buf_1 _09874_ (.A(\i_mandel.i_sq_x.x[-10] ),
    .X(_01908_));
 sg13g2_nand2b_1 _09875_ (.Y(_01909_),
    .B(net323),
    .A_N(net281));
 sg13g2_a21oi_1 _09876_ (.A1(_01549_),
    .A2(_01523_),
    .Y(_01910_),
    .B1(_01909_));
 sg13g2_and4_1 _09877_ (.A(net323),
    .B(net281),
    .C(_01549_),
    .D(net189),
    .X(_01911_));
 sg13g2_nand2b_1 _09878_ (.Y(_01912_),
    .B(net241),
    .A_N(_01613_));
 sg13g2_a21o_1 _09879_ (.A2(_01612_),
    .A1(_01596_),
    .B1(_01912_),
    .X(_01913_));
 sg13g2_nor3_1 _09880_ (.A(_01910_),
    .B(_01911_),
    .C(_01913_),
    .Y(_01914_));
 sg13g2_and4_1 _09881_ (.A(net323),
    .B(_01547_),
    .C(_01551_),
    .D(_01913_),
    .X(_01915_));
 sg13g2_buf_1 _09882_ (.A(_01915_),
    .X(_01916_));
 sg13g2_or2_1 _09883_ (.X(_01917_),
    .B(_01916_),
    .A(_01914_));
 sg13g2_xnor2_1 _09884_ (.Y(_01918_),
    .A(_01617_),
    .B(_01917_));
 sg13g2_xor2_1 _09885_ (.B(_01918_),
    .A(_01907_),
    .X(_01919_));
 sg13g2_o21ai_1 _09886_ (.B1(_01919_),
    .Y(_01920_),
    .A1(_01619_),
    .A2(_01902_));
 sg13g2_buf_1 _09887_ (.A(_01615_),
    .X(_01921_));
 sg13g2_inv_2 _09888_ (.Y(_01922_),
    .A(net323));
 sg13g2_nor2_1 _09889_ (.A(net187),
    .B(net184),
    .Y(_01923_));
 sg13g2_nand3_1 _09890_ (.B(net240),
    .C(_01923_),
    .A(_01922_),
    .Y(_01924_));
 sg13g2_buf_1 _09891_ (.A(_01611_),
    .X(_01925_));
 sg13g2_buf_1 _09892_ (.A(net239),
    .X(_01926_));
 sg13g2_buf_1 _09893_ (.A(_01617_),
    .X(_01927_));
 sg13g2_o21ai_1 _09894_ (.B1(net90),
    .Y(_01928_),
    .A1(_01914_),
    .A2(_01916_));
 sg13g2_nor3_1 _09895_ (.A(net90),
    .B(_01914_),
    .C(_01916_),
    .Y(_01929_));
 sg13g2_a21oi_1 _09896_ (.A1(_01903_),
    .A2(_01928_),
    .Y(_01930_),
    .B1(_01929_));
 sg13g2_a21oi_1 _09897_ (.A1(net90),
    .A2(_01905_),
    .Y(_01931_),
    .B1(_01904_));
 sg13g2_nor2_1 _09898_ (.A(net90),
    .B(_01905_),
    .Y(_01932_));
 sg13g2_a21oi_1 _09899_ (.A1(_01917_),
    .A2(_01931_),
    .Y(_01933_),
    .B1(_01932_));
 sg13g2_o21ai_1 _09900_ (.B1(_01933_),
    .Y(_01934_),
    .A1(_01887_),
    .A2(_01930_));
 sg13g2_buf_1 _09901_ (.A(_01934_),
    .X(_01935_));
 sg13g2_nor2_1 _09902_ (.A(_01538_),
    .B(net188),
    .Y(_01936_));
 sg13g2_a21oi_1 _09903_ (.A1(_01547_),
    .A2(_01551_),
    .Y(_01937_),
    .B1(_01923_));
 sg13g2_nor2_1 _09904_ (.A(_01936_),
    .B(_01937_),
    .Y(_01938_));
 sg13g2_nor2_1 _09905_ (.A(_01922_),
    .B(_01938_),
    .Y(_01939_));
 sg13g2_nand3_1 _09906_ (.B(_01935_),
    .C(_01939_),
    .A(net183),
    .Y(_01940_));
 sg13g2_o21ai_1 _09907_ (.B1(net323),
    .Y(_01941_),
    .A1(_01936_),
    .A2(_01937_));
 sg13g2_nand3b_1 _09908_ (.B(_01941_),
    .C(_01833_),
    .Y(_01942_),
    .A_N(_01935_));
 sg13g2_nand4_1 _09909_ (.B(_01924_),
    .C(_01940_),
    .A(net124),
    .Y(_01943_),
    .D(_01942_));
 sg13g2_a21o_1 _09910_ (.A2(_01920_),
    .A1(_01898_),
    .B1(_01943_),
    .X(_01944_));
 sg13g2_a221oi_1 _09911_ (.B2(_01885_),
    .C1(_01944_),
    .B1(_01745_),
    .A1(net35),
    .Y(_01945_),
    .A2(_01744_));
 sg13g2_buf_1 _09912_ (.A(_01945_),
    .X(_01946_));
 sg13g2_and3_1 _09913_ (.X(_01947_),
    .A(_01889_),
    .B(_01891_),
    .C(_01927_));
 sg13g2_o21ai_1 _09914_ (.B1(_01947_),
    .Y(_01948_),
    .A1(net63),
    .A2(net84));
 sg13g2_a21o_1 _09915_ (.A2(_01891_),
    .A1(_01889_),
    .B1(_01927_),
    .X(_01949_));
 sg13g2_a21o_1 _09916_ (.A2(net84),
    .A1(_01620_),
    .B1(_01949_),
    .X(_01950_));
 sg13g2_and2_1 _09917_ (.A(_01948_),
    .B(_01950_),
    .X(_01951_));
 sg13g2_nor2_1 _09918_ (.A(_01634_),
    .B(_01919_),
    .Y(_01952_));
 sg13g2_xnor2_1 _09919_ (.Y(_01953_),
    .A(_01907_),
    .B(_01918_));
 sg13g2_and3_1 _09920_ (.X(_01954_),
    .A(_01889_),
    .B(_01891_),
    .C(_01692_));
 sg13g2_o21ai_1 _09921_ (.B1(net90),
    .Y(_01955_),
    .A1(_01625_),
    .A2(_01631_));
 sg13g2_nor3_1 _09922_ (.A(_01580_),
    .B(_01623_),
    .C(_01955_),
    .Y(_01956_));
 sg13g2_a21o_1 _09923_ (.A2(_01954_),
    .A1(net63),
    .B1(_01956_),
    .X(_01957_));
 sg13g2_inv_1 _09924_ (.Y(_01958_),
    .A(_01609_));
 sg13g2_or3_1 _09925_ (.A(_01580_),
    .B(_01623_),
    .C(_01955_),
    .X(_01959_));
 sg13g2_nand2b_1 _09926_ (.Y(_01960_),
    .B(_01685_),
    .A_N(_01684_));
 sg13g2_nand2_1 _09927_ (.Y(_01961_),
    .A(_01599_),
    .B(_01606_));
 sg13g2_and4_1 _09928_ (.A(_01576_),
    .B(_01563_),
    .C(_01960_),
    .D(_01961_),
    .X(_01962_));
 sg13g2_a22oi_1 _09929_ (.Y(_01963_),
    .B1(_01962_),
    .B2(_01892_),
    .A2(_01959_),
    .A1(_01958_));
 sg13g2_and3_1 _09930_ (.X(_01964_),
    .A(_01953_),
    .B(_01957_),
    .C(_01963_));
 sg13g2_a21oi_1 _09931_ (.A1(_01951_),
    .A2(_01952_),
    .Y(_01965_),
    .B1(_01964_));
 sg13g2_nand3_1 _09932_ (.B(_01948_),
    .C(_01950_),
    .A(_01901_),
    .Y(_01966_));
 sg13g2_a21oi_1 _09933_ (.A1(_01957_),
    .A2(_01963_),
    .Y(_01967_),
    .B1(_01953_));
 sg13g2_nand2_1 _09934_ (.Y(_01968_),
    .A(_01966_),
    .B(_01967_));
 sg13g2_a221oi_1 _09935_ (.B2(_01968_),
    .C1(_01943_),
    .B1(_01965_),
    .A1(_01898_),
    .Y(_01969_),
    .A2(_01920_));
 sg13g2_nand2_1 _09936_ (.Y(_01970_),
    .A(_01922_),
    .B(_01923_));
 sg13g2_a21oi_1 _09937_ (.A1(_01970_),
    .A2(_01941_),
    .Y(_01971_),
    .B1(net240));
 sg13g2_and3_1 _09938_ (.X(_01972_),
    .A(net240),
    .B(_01970_),
    .C(_01941_));
 sg13g2_o21ai_1 _09939_ (.B1(net124),
    .Y(_01973_),
    .A1(_01971_),
    .A2(_01972_));
 sg13g2_xor2_1 _09940_ (.B(_01973_),
    .A(_01935_),
    .X(_01974_));
 sg13g2_nor2_1 _09941_ (.A(_01943_),
    .B(_01974_),
    .Y(_01975_));
 sg13g2_and4_1 _09942_ (.A(net183),
    .B(net124),
    .C(_01935_),
    .D(_01939_),
    .X(_01976_));
 sg13g2_or3_1 _09943_ (.A(_01969_),
    .B(_01975_),
    .C(_01976_),
    .X(_01977_));
 sg13g2_buf_1 _09944_ (.A(_01977_),
    .X(_01978_));
 sg13g2_nor2_1 _09945_ (.A(_01946_),
    .B(_01978_),
    .Y(_01979_));
 sg13g2_buf_1 _09946_ (.A(_01979_),
    .X(_01980_));
 sg13g2_buf_1 _09947_ (.A(net284),
    .X(_01981_));
 sg13g2_buf_1 _09948_ (.A(net238),
    .X(_01982_));
 sg13g2_buf_1 _09949_ (.A(_01823_),
    .X(_01983_));
 sg13g2_buf_2 _09950_ (.A(\i_mandel.i_sq_x.x[-8] ),
    .X(_01984_));
 sg13g2_buf_1 _09951_ (.A(\i_mandel.i_sq_x.x[-9] ),
    .X(_01985_));
 sg13g2_buf_1 _09952_ (.A(_01985_),
    .X(_01986_));
 sg13g2_xor2_1 _09953_ (.B(net278),
    .A(_01984_),
    .X(_01987_));
 sg13g2_buf_2 _09954_ (.A(_01987_),
    .X(_01988_));
 sg13g2_xnor2_1 _09955_ (.Y(_01989_),
    .A(net181),
    .B(_01988_));
 sg13g2_buf_1 _09956_ (.A(net280),
    .X(_01990_));
 sg13g2_inv_1 _09957_ (.Y(_01991_),
    .A(net237));
 sg13g2_buf_2 _09958_ (.A(\i_mandel.i_sq_x.x[-7] ),
    .X(_01992_));
 sg13g2_inv_1 _09959_ (.Y(_01993_),
    .A(_01992_));
 sg13g2_nor2_2 _09960_ (.A(_01991_),
    .B(_01993_),
    .Y(_01994_));
 sg13g2_nand3_1 _09961_ (.B(_01989_),
    .C(_01994_),
    .A(net182),
    .Y(_01995_));
 sg13g2_buf_1 _09962_ (.A(_01995_),
    .X(_01996_));
 sg13g2_nor2_1 _09963_ (.A(net32),
    .B(_01996_),
    .Y(_01997_));
 sg13g2_buf_1 _09964_ (.A(_01997_),
    .X(_01998_));
 sg13g2_nand2_1 _09965_ (.Y(_01999_),
    .A(_01984_),
    .B(net278));
 sg13g2_buf_1 _09966_ (.A(_01999_),
    .X(_02000_));
 sg13g2_buf_1 _09967_ (.A(_01984_),
    .X(_02001_));
 sg13g2_buf_1 _09968_ (.A(net279),
    .X(_02002_));
 sg13g2_o21ai_1 _09969_ (.B1(net236),
    .Y(_02003_),
    .A1(net277),
    .A2(net278));
 sg13g2_a21oi_1 _09970_ (.A1(_02000_),
    .A2(_02003_),
    .Y(_02004_),
    .B1(net244));
 sg13g2_buf_1 _09971_ (.A(_02004_),
    .X(_02005_));
 sg13g2_buf_1 _09972_ (.A(net288),
    .X(_02006_));
 sg13g2_buf_1 _09973_ (.A(net235),
    .X(_02007_));
 sg13g2_buf_1 _09974_ (.A(net180),
    .X(_02008_));
 sg13g2_buf_1 _09975_ (.A(net287),
    .X(_02009_));
 sg13g2_buf_1 _09976_ (.A(net325),
    .X(_02010_));
 sg13g2_and2_1 _09977_ (.A(net234),
    .B(net276),
    .X(_02011_));
 sg13g2_buf_1 _09978_ (.A(_02011_),
    .X(_02012_));
 sg13g2_buf_1 _09979_ (.A(net234),
    .X(_02013_));
 sg13g2_buf_1 _09980_ (.A(net179),
    .X(_02014_));
 sg13g2_buf_1 _09981_ (.A(net276),
    .X(_02015_));
 sg13g2_buf_1 _09982_ (.A(_02015_),
    .X(_02016_));
 sg13g2_buf_1 _09983_ (.A(net178),
    .X(_02017_));
 sg13g2_or2_1 _09984_ (.X(_02018_),
    .B(net151),
    .A(net152));
 sg13g2_buf_1 _09985_ (.A(net182),
    .X(_02019_));
 sg13g2_o21ai_1 _09986_ (.B1(net150),
    .Y(_02020_),
    .A1(net180),
    .A2(_02018_));
 sg13g2_a21o_1 _09987_ (.A2(_02012_),
    .A1(net153),
    .B1(_02020_),
    .X(_02021_));
 sg13g2_xor2_1 _09988_ (.B(_02021_),
    .A(net123),
    .X(_02022_));
 sg13g2_buf_1 _09989_ (.A(_02022_),
    .X(_02023_));
 sg13g2_nand2_2 _09990_ (.Y(_02024_),
    .A(net234),
    .B(net233));
 sg13g2_nand2b_1 _09991_ (.Y(_02025_),
    .B(_02024_),
    .A_N(_02005_));
 sg13g2_a22oi_1 _09992_ (.Y(_02026_),
    .B1(_02025_),
    .B2(net153),
    .A2(_02018_),
    .A1(net123));
 sg13g2_nor2_1 _09993_ (.A(net191),
    .B(_02026_),
    .Y(_02027_));
 sg13g2_buf_1 _09994_ (.A(_02027_),
    .X(_02028_));
 sg13g2_buf_1 _09995_ (.A(net150),
    .X(_02029_));
 sg13g2_buf_1 _09996_ (.A(net282),
    .X(_02030_));
 sg13g2_buf_1 _09997_ (.A(net232),
    .X(_02031_));
 sg13g2_buf_1 _09998_ (.A(net177),
    .X(_02032_));
 sg13g2_nor2_1 _09999_ (.A(net154),
    .B(net149),
    .Y(_02033_));
 sg13g2_buf_1 _10000_ (.A(net292),
    .X(_02034_));
 sg13g2_xnor2_1 _10001_ (.Y(_02035_),
    .A(_02034_),
    .B(net122));
 sg13g2_a22oi_1 _10002_ (.Y(_02036_),
    .B1(_02035_),
    .B2(net154),
    .A2(_02033_),
    .A1(net122));
 sg13g2_buf_1 _10003_ (.A(_02036_),
    .X(_02037_));
 sg13g2_nand2_1 _10004_ (.Y(_02038_),
    .A(net79),
    .B(_02037_));
 sg13g2_o21ai_1 _10005_ (.B1(_02038_),
    .Y(_02039_),
    .A1(net79),
    .A2(net78));
 sg13g2_buf_1 _10006_ (.A(_01991_),
    .X(_02040_));
 sg13g2_buf_1 _10007_ (.A(_01993_),
    .X(_02041_));
 sg13g2_nand2_1 _10008_ (.Y(_02042_),
    .A(net148),
    .B(net230));
 sg13g2_o21ai_1 _10009_ (.B1(net182),
    .Y(_02043_),
    .A1(_01989_),
    .A2(_02042_));
 sg13g2_buf_1 _10010_ (.A(_02043_),
    .X(_02044_));
 sg13g2_and2_1 _10011_ (.A(net32),
    .B(_02044_),
    .X(_02045_));
 sg13g2_buf_1 _10012_ (.A(_02045_),
    .X(_02046_));
 sg13g2_and2_1 _10013_ (.A(_02046_),
    .B(net79),
    .X(_02047_));
 sg13g2_buf_1 _10014_ (.A(_02047_),
    .X(_02048_));
 sg13g2_nand2_1 _10015_ (.Y(_02049_),
    .A(_02048_),
    .B(net78));
 sg13g2_nand2b_1 _10016_ (.Y(_02050_),
    .B(_02037_),
    .A_N(_02048_));
 sg13g2_a21oi_1 _10017_ (.A1(_02049_),
    .A2(_02050_),
    .Y(_02051_),
    .B1(net29));
 sg13g2_a21oi_1 _10018_ (.A1(net29),
    .A2(_02039_),
    .Y(_02052_),
    .B1(_02051_));
 sg13g2_xor2_1 _10019_ (.B(_02052_),
    .A(_01503_),
    .X(_02053_));
 sg13g2_buf_1 _10020_ (.A(net231),
    .X(_02054_));
 sg13g2_nand2_1 _10021_ (.Y(_02055_),
    .A(net176),
    .B(net78));
 sg13g2_o21ai_1 _10022_ (.B1(_02055_),
    .Y(_02056_),
    .A1(net176),
    .A2(net245));
 sg13g2_buf_1 _10023_ (.A(_01490_),
    .X(_02057_));
 sg13g2_a22oi_1 _10024_ (.Y(_02058_),
    .B1(_02056_),
    .B2(net121),
    .A2(_02033_),
    .A1(_02028_));
 sg13g2_buf_1 _10025_ (.A(net122),
    .X(_02059_));
 sg13g2_nand2b_1 _10026_ (.Y(_02060_),
    .B(net106),
    .A_N(_02058_));
 sg13g2_inv_1 _10027_ (.Y(_02061_),
    .A(net29));
 sg13g2_nor2_1 _10028_ (.A(_02061_),
    .B(_02023_),
    .Y(_02062_));
 sg13g2_nor2_1 _10029_ (.A(_02048_),
    .B(_02062_),
    .Y(_02063_));
 sg13g2_or2_1 _10030_ (.X(_02064_),
    .B(_01503_),
    .A(_02037_));
 sg13g2_nand3_1 _10031_ (.B(_02037_),
    .C(_01503_),
    .A(net78),
    .Y(_02065_));
 sg13g2_o21ai_1 _10032_ (.B1(_02065_),
    .Y(_02066_),
    .A1(net78),
    .A2(_02064_));
 sg13g2_xor2_1 _10033_ (.B(_01503_),
    .A(net78),
    .X(_02067_));
 sg13g2_a22oi_1 _10034_ (.Y(_02068_),
    .B1(_02067_),
    .B2(_02062_),
    .A2(_02066_),
    .A1(_02063_));
 sg13g2_inv_2 _10035_ (.Y(_02069_),
    .A(net288));
 sg13g2_nor2_1 _10036_ (.A(net152),
    .B(net151),
    .Y(_02070_));
 sg13g2_nor3_1 _10037_ (.A(net192),
    .B(_02069_),
    .C(_02070_),
    .Y(_02071_));
 sg13g2_a21oi_1 _10038_ (.A1(_02069_),
    .A2(_02070_),
    .Y(_02072_),
    .B1(_02071_));
 sg13g2_a22oi_1 _10039_ (.Y(_02073_),
    .B1(_02072_),
    .B2(_02005_),
    .A2(_02012_),
    .A1(net153));
 sg13g2_nand2b_1 _10040_ (.Y(_02074_),
    .B(net122),
    .A_N(_02073_));
 sg13g2_inv_1 _10041_ (.Y(_02075_),
    .A(_02074_));
 sg13g2_o21ai_1 _10042_ (.B1(net106),
    .Y(_02076_),
    .A1(_02069_),
    .A2(_02075_));
 sg13g2_or2_1 _10043_ (.X(_02077_),
    .B(_02029_),
    .A(net154));
 sg13g2_nand3_1 _10044_ (.B(net149),
    .C(_02029_),
    .A(net154),
    .Y(_02078_));
 sg13g2_a22oi_1 _10045_ (.Y(_02079_),
    .B1(_02077_),
    .B2(_02078_),
    .A2(_02075_),
    .A1(net176));
 sg13g2_a221oi_1 _10046_ (.B2(net245),
    .C1(_02079_),
    .B1(_02076_),
    .A1(_01501_),
    .Y(_02080_),
    .A2(_02074_));
 sg13g2_o21ai_1 _10047_ (.B1(_02019_),
    .Y(_02081_),
    .A1(_01501_),
    .A2(net153));
 sg13g2_xnor2_1 _10048_ (.Y(_02082_),
    .A(net192),
    .B(_02034_));
 sg13g2_a21o_1 _10049_ (.A2(_02019_),
    .A1(net149),
    .B1(_02082_),
    .X(_02083_));
 sg13g2_nand2_1 _10050_ (.Y(_02084_),
    .A(net122),
    .B(_02082_));
 sg13g2_a22oi_1 _10051_ (.Y(_02085_),
    .B1(_02083_),
    .B2(_02084_),
    .A2(_02081_),
    .A1(_01493_));
 sg13g2_xnor2_1 _10052_ (.Y(_02086_),
    .A(_02074_),
    .B(_02085_));
 sg13g2_o21ai_1 _10053_ (.B1(_02086_),
    .Y(_02087_),
    .A1(_02046_),
    .A2(net79));
 sg13g2_o21ai_1 _10054_ (.B1(_02024_),
    .Y(_02088_),
    .A1(net192),
    .A2(_02070_));
 sg13g2_a21oi_1 _10055_ (.A1(net180),
    .A2(_02088_),
    .Y(_02089_),
    .B1(_02020_));
 sg13g2_xnor2_1 _10056_ (.Y(_02090_),
    .A(net123),
    .B(_02089_));
 sg13g2_buf_1 _10057_ (.A(_02090_),
    .X(_02091_));
 sg13g2_nor2_1 _10058_ (.A(net79),
    .B(_02086_),
    .Y(_02092_));
 sg13g2_a221oi_1 _10059_ (.B2(_02091_),
    .C1(_02092_),
    .B1(_02087_),
    .A1(_02046_),
    .Y(_02093_),
    .A2(net79));
 sg13g2_inv_1 _10060_ (.Y(_02094_),
    .A(_02086_));
 sg13g2_nand3_1 _10061_ (.B(net79),
    .C(_02094_),
    .A(net29),
    .Y(_02095_));
 sg13g2_o21ai_1 _10062_ (.B1(_02095_),
    .Y(_02096_),
    .A1(net29),
    .A2(_02093_));
 sg13g2_buf_1 _10063_ (.A(_02096_),
    .X(_02097_));
 sg13g2_xnor2_1 _10064_ (.Y(_02098_),
    .A(net78),
    .B(_02037_));
 sg13g2_xnor2_1 _10065_ (.Y(_02099_),
    .A(_02063_),
    .B(_02098_));
 sg13g2_nand2_1 _10066_ (.Y(_02100_),
    .A(_02097_),
    .B(_02099_));
 sg13g2_nor2_1 _10067_ (.A(_02097_),
    .B(_02099_),
    .Y(_02101_));
 sg13g2_a21oi_1 _10068_ (.A1(_02080_),
    .A2(_02100_),
    .Y(_02102_),
    .B1(_02101_));
 sg13g2_a21oi_1 _10069_ (.A1(_02053_),
    .A2(_02060_),
    .Y(_02103_),
    .B1(_02102_));
 sg13g2_xor2_1 _10070_ (.B(_02103_),
    .A(_02068_),
    .X(_02104_));
 sg13g2_o21ai_1 _10071_ (.B1(_02104_),
    .Y(_02105_),
    .A1(_02053_),
    .A2(_02060_));
 sg13g2_nor2_1 _10072_ (.A(net198),
    .B(_00399_),
    .Y(_02106_));
 sg13g2_nand2_1 _10073_ (.Y(_02107_),
    .A(net127),
    .B(_07313_));
 sg13g2_and2_1 _10074_ (.A(_02106_),
    .B(_02107_),
    .X(_02108_));
 sg13g2_buf_1 _10075_ (.A(net156),
    .X(_02109_));
 sg13g2_nor2_1 _10076_ (.A(net127),
    .B(net27),
    .Y(_02110_));
 sg13g2_nor2_1 _10077_ (.A(net156),
    .B(net128),
    .Y(_02111_));
 sg13g2_a22oi_1 _10078_ (.Y(_02112_),
    .B1(_02111_),
    .B2(net27),
    .A2(_02110_),
    .A1(net120));
 sg13g2_nor2_1 _10079_ (.A(_00406_),
    .B(_02112_),
    .Y(_02113_));
 sg13g2_nand2_1 _10080_ (.Y(_02114_),
    .A(net200),
    .B(net27));
 sg13g2_nand3_1 _10081_ (.B(_00369_),
    .C(_00399_),
    .A(net128),
    .Y(_02115_));
 sg13g2_a21oi_1 _10082_ (.A1(_02114_),
    .A2(_02115_),
    .Y(_02116_),
    .B1(net120));
 sg13g2_nor4_1 _10083_ (.A(_00397_),
    .B(_02108_),
    .C(_02113_),
    .D(_02116_),
    .Y(_02117_));
 sg13g2_nor2b_1 _10084_ (.A(net27),
    .B_N(_02111_),
    .Y(_02118_));
 sg13g2_a21oi_1 _10085_ (.A1(net120),
    .A2(net27),
    .Y(_02119_),
    .B1(_02118_));
 sg13g2_nor2_1 _10086_ (.A(_02109_),
    .B(_00382_),
    .Y(_02120_));
 sg13g2_nor2_1 _10087_ (.A(_00371_),
    .B(net200),
    .Y(_02121_));
 sg13g2_mux2_1 _10088_ (.A0(net156),
    .A1(_02121_),
    .S(net27),
    .X(_02122_));
 sg13g2_a22oi_1 _10089_ (.Y(_02123_),
    .B1(_02122_),
    .B2(_00406_),
    .A2(_00399_),
    .A1(_02120_));
 sg13g2_o21ai_1 _10090_ (.B1(_02123_),
    .Y(_02124_),
    .A1(_00406_),
    .A2(_02119_));
 sg13g2_nor2_1 _10091_ (.A(net67),
    .B(_02124_),
    .Y(_02125_));
 sg13g2_a21oi_1 _10092_ (.A1(net120),
    .A2(net67),
    .Y(_02126_),
    .B1(net128));
 sg13g2_nor2_1 _10093_ (.A(_00406_),
    .B(_00399_),
    .Y(_02127_));
 sg13g2_a21o_1 _10094_ (.A2(_00405_),
    .A1(_00399_),
    .B1(_02127_),
    .X(_02128_));
 sg13g2_a22oi_1 _10095_ (.Y(_02129_),
    .B1(_02128_),
    .B2(net120),
    .A2(_02126_),
    .A1(_02106_));
 sg13g2_nand2_1 _10096_ (.Y(_02130_),
    .A(net198),
    .B(net127));
 sg13g2_buf_1 _10097_ (.A(_02130_),
    .X(_02131_));
 sg13g2_nor4_1 _10098_ (.A(net156),
    .B(net27),
    .C(net67),
    .D(_02131_),
    .Y(_02132_));
 sg13g2_a21o_1 _10099_ (.A2(_02106_),
    .A1(net67),
    .B1(_02132_),
    .X(_02133_));
 sg13g2_a21oi_1 _10100_ (.A1(net127),
    .A2(_00397_),
    .Y(_02134_),
    .B1(net120));
 sg13g2_a221oi_1 _10101_ (.B2(_02127_),
    .C1(_00374_),
    .B1(_02134_),
    .A1(net128),
    .Y(_02135_),
    .A2(_02133_));
 sg13g2_o21ai_1 _10102_ (.B1(_02135_),
    .Y(_02136_),
    .A1(_00363_),
    .A2(_02129_));
 sg13g2_o21ai_1 _10103_ (.B1(_02136_),
    .Y(_02137_),
    .A1(_02117_),
    .A2(_02125_));
 sg13g2_nand2_1 _10104_ (.Y(_02138_),
    .A(_00393_),
    .B(_00410_));
 sg13g2_nand2_1 _10105_ (.Y(_02139_),
    .A(_00368_),
    .B(_00371_));
 sg13g2_o21ai_1 _10106_ (.B1(_02121_),
    .Y(_02140_),
    .A1(_00406_),
    .A2(_00361_));
 sg13g2_a21oi_1 _10107_ (.A1(_02139_),
    .A2(_02140_),
    .Y(_02141_),
    .B1(_00399_));
 sg13g2_o21ai_1 _10108_ (.B1(_00395_),
    .Y(_02142_),
    .A1(_00398_),
    .A2(_02141_));
 sg13g2_o21ai_1 _10109_ (.B1(_02142_),
    .Y(_02143_),
    .A1(_00395_),
    .A2(_00397_));
 sg13g2_o21ai_1 _10110_ (.B1(_02049_),
    .Y(_02144_),
    .A1(_02048_),
    .A2(_01503_));
 sg13g2_mux2_1 _10111_ (.A0(net78),
    .A1(_01503_),
    .S(_02023_),
    .X(_02145_));
 sg13g2_nand2_1 _10112_ (.Y(_02146_),
    .A(_01998_),
    .B(_02145_));
 sg13g2_o21ai_1 _10113_ (.B1(_02146_),
    .Y(_02147_),
    .A1(_01998_),
    .A2(_02144_));
 sg13g2_nor3_1 _10114_ (.A(_00368_),
    .B(net156),
    .C(_00397_),
    .Y(_02148_));
 sg13g2_nor3_1 _10115_ (.A(_00406_),
    .B(net67),
    .C(_02111_),
    .Y(_02149_));
 sg13g2_o21ai_1 _10116_ (.B1(net127),
    .Y(_02150_),
    .A1(_02148_),
    .A2(_02149_));
 sg13g2_nor4_1 _10117_ (.A(net121),
    .B(net176),
    .C(net191),
    .D(_02026_),
    .Y(_02151_));
 sg13g2_o21ai_1 _10118_ (.B1(net154),
    .Y(_02152_),
    .A1(net176),
    .A2(net149));
 sg13g2_nor2_1 _10119_ (.A(_02028_),
    .B(_02152_),
    .Y(_02153_));
 sg13g2_o21ai_1 _10120_ (.B1(net106),
    .Y(_02154_),
    .A1(_02151_),
    .A2(_02153_));
 sg13g2_xnor2_1 _10121_ (.Y(_02155_),
    .A(_02150_),
    .B(_02154_));
 sg13g2_xnor2_1 _10122_ (.Y(_02156_),
    .A(_02147_),
    .B(_02155_));
 sg13g2_xnor2_1 _10123_ (.Y(_02157_),
    .A(_02143_),
    .B(_02156_));
 sg13g2_xnor2_1 _10124_ (.Y(_02158_),
    .A(_02138_),
    .B(_02157_));
 sg13g2_xnor2_1 _10125_ (.Y(_02159_),
    .A(_02137_),
    .B(_02158_));
 sg13g2_xnor2_1 _10126_ (.Y(_02160_),
    .A(_02105_),
    .B(_02159_));
 sg13g2_xnor2_1 _10127_ (.Y(_02161_),
    .A(_01485_),
    .B(_02160_));
 sg13g2_xnor2_1 _10128_ (.Y(_02162_),
    .A(_02053_),
    .B(_02060_));
 sg13g2_xnor2_1 _10129_ (.Y(_02163_),
    .A(_02102_),
    .B(_02162_));
 sg13g2_nand2_2 _10130_ (.Y(_02164_),
    .A(net232),
    .B(net288));
 sg13g2_nand2_1 _10131_ (.Y(_02165_),
    .A(net292),
    .B(net234));
 sg13g2_nand2_1 _10132_ (.Y(_02166_),
    .A(net293),
    .B(net233));
 sg13g2_a21oi_1 _10133_ (.A1(_02164_),
    .A2(_02165_),
    .Y(_02167_),
    .B1(_02166_));
 sg13g2_or2_1 _10134_ (.X(_02168_),
    .B(_02167_),
    .A(_01549_));
 sg13g2_buf_1 _10135_ (.A(_02168_),
    .X(_02169_));
 sg13g2_nand2_1 _10136_ (.Y(_02170_),
    .A(net292),
    .B(_02006_));
 sg13g2_buf_2 _10137_ (.A(_02170_),
    .X(_02171_));
 sg13g2_nand2_1 _10138_ (.Y(_02172_),
    .A(net178),
    .B(_01982_));
 sg13g2_nand2_1 _10139_ (.Y(_02173_),
    .A(_01488_),
    .B(net179));
 sg13g2_buf_2 _10140_ (.A(_02173_),
    .X(_02174_));
 sg13g2_xor2_1 _10141_ (.B(_02174_),
    .A(_02172_),
    .X(_02175_));
 sg13g2_xnor2_1 _10142_ (.Y(_02176_),
    .A(_02171_),
    .B(_02175_));
 sg13g2_a21oi_1 _10143_ (.A1(net123),
    .A2(_02169_),
    .Y(_02177_),
    .B1(_02176_));
 sg13g2_nor2_1 _10144_ (.A(net123),
    .B(_02169_),
    .Y(_02178_));
 sg13g2_nor2_1 _10145_ (.A(_02177_),
    .B(_02178_),
    .Y(_02179_));
 sg13g2_xnor2_1 _10146_ (.Y(_02180_),
    .A(net290),
    .B(_02171_));
 sg13g2_xor2_1 _10147_ (.B(_02180_),
    .A(_02174_),
    .X(_02181_));
 sg13g2_a21oi_1 _10148_ (.A1(_02169_),
    .A2(_02181_),
    .Y(_02182_),
    .B1(_01727_));
 sg13g2_nor2_1 _10149_ (.A(_02169_),
    .B(_02181_),
    .Y(_02183_));
 sg13g2_nor2_1 _10150_ (.A(_02182_),
    .B(_02183_),
    .Y(_02184_));
 sg13g2_nand2_1 _10151_ (.Y(_02185_),
    .A(_02179_),
    .B(_02184_));
 sg13g2_nand3_1 _10152_ (.B(net177),
    .C(net180),
    .A(net292),
    .Y(_02186_));
 sg13g2_o21ai_1 _10153_ (.B1(_02186_),
    .Y(_02187_),
    .A1(_02174_),
    .A2(_02180_));
 sg13g2_inv_1 _10154_ (.Y(_02188_),
    .A(net287));
 sg13g2_nand2_1 _10155_ (.Y(_02189_),
    .A(_02188_),
    .B(net150));
 sg13g2_and2_1 _10156_ (.A(net246),
    .B(_02006_),
    .X(_02190_));
 sg13g2_buf_1 _10157_ (.A(_02190_),
    .X(_02191_));
 sg13g2_xnor2_1 _10158_ (.Y(_02192_),
    .A(_02189_),
    .B(_02191_));
 sg13g2_xnor2_1 _10159_ (.Y(_02193_),
    .A(_02187_),
    .B(_02192_));
 sg13g2_nor2_1 _10160_ (.A(_02179_),
    .B(_02184_),
    .Y(_02194_));
 sg13g2_a21oi_1 _10161_ (.A1(_02185_),
    .A2(_02193_),
    .Y(_02195_),
    .B1(_02194_));
 sg13g2_xor2_1 _10162_ (.B(net178),
    .A(net179),
    .X(_02196_));
 sg13g2_nand2_1 _10163_ (.Y(_02197_),
    .A(_01982_),
    .B(_02196_));
 sg13g2_xnor2_1 _10164_ (.Y(_02198_),
    .A(_02191_),
    .B(_02197_));
 sg13g2_nand2_1 _10165_ (.Y(_02199_),
    .A(_02171_),
    .B(_02174_));
 sg13g2_o21ai_1 _10166_ (.B1(_02172_),
    .Y(_02200_),
    .A1(_02171_),
    .A2(_02174_));
 sg13g2_and2_1 _10167_ (.A(_02199_),
    .B(_02200_),
    .X(_02201_));
 sg13g2_buf_1 _10168_ (.A(_02201_),
    .X(_02202_));
 sg13g2_xor2_1 _10169_ (.B(_02202_),
    .A(net123),
    .X(_02203_));
 sg13g2_xnor2_1 _10170_ (.Y(_02204_),
    .A(_02198_),
    .B(_02203_));
 sg13g2_buf_2 _10171_ (.A(_02204_),
    .X(_02205_));
 sg13g2_nand2_1 _10172_ (.Y(_02206_),
    .A(net32),
    .B(_02044_));
 sg13g2_o21ai_1 _10173_ (.B1(_02206_),
    .Y(_02207_),
    .A1(net29),
    .A2(_02205_));
 sg13g2_nor2_1 _10174_ (.A(_02198_),
    .B(_02202_),
    .Y(_02208_));
 sg13g2_a21oi_1 _10175_ (.A1(_02198_),
    .A2(_02202_),
    .Y(_02209_),
    .B1(net123));
 sg13g2_nor2_1 _10176_ (.A(_02208_),
    .B(_02209_),
    .Y(_02210_));
 sg13g2_nand2_1 _10177_ (.Y(_02211_),
    .A(_02069_),
    .B(net150));
 sg13g2_nor2_1 _10178_ (.A(_01501_),
    .B(net177),
    .Y(_02212_));
 sg13g2_xnor2_1 _10179_ (.Y(_02213_),
    .A(_02211_),
    .B(_02212_));
 sg13g2_nand2b_1 _10180_ (.Y(_02214_),
    .B(_02189_),
    .A_N(_02187_));
 sg13g2_nor3_1 _10181_ (.A(net152),
    .B(net191),
    .C(_02186_),
    .Y(_02215_));
 sg13g2_a21oi_1 _10182_ (.A1(_02191_),
    .A2(_02214_),
    .Y(_02216_),
    .B1(_02215_));
 sg13g2_xnor2_1 _10183_ (.Y(_02217_),
    .A(_02213_),
    .B(_02216_));
 sg13g2_xnor2_1 _10184_ (.Y(_02218_),
    .A(_02210_),
    .B(_02217_));
 sg13g2_xor2_1 _10185_ (.B(_02218_),
    .A(_02091_),
    .X(_02219_));
 sg13g2_xnor2_1 _10186_ (.Y(_02220_),
    .A(_02207_),
    .B(_02219_));
 sg13g2_or2_1 _10187_ (.X(_02221_),
    .B(_02220_),
    .A(_02195_));
 sg13g2_nand2_1 _10188_ (.Y(_02222_),
    .A(_02195_),
    .B(_02220_));
 sg13g2_xnor2_1 _10189_ (.Y(_02223_),
    .A(_02175_),
    .B(net123));
 sg13g2_xnor2_1 _10190_ (.Y(_02224_),
    .A(_02171_),
    .B(_02169_));
 sg13g2_xnor2_1 _10191_ (.Y(_02225_),
    .A(_02223_),
    .B(_02224_));
 sg13g2_xor2_1 _10192_ (.B(_02184_),
    .A(_02179_),
    .X(_02226_));
 sg13g2_xnor2_1 _10193_ (.Y(_02227_),
    .A(_02193_),
    .B(_02226_));
 sg13g2_o21ai_1 _10194_ (.B1(_02227_),
    .Y(_02228_),
    .A1(_02205_),
    .A2(_02225_));
 sg13g2_inv_1 _10195_ (.Y(_02229_),
    .A(_02228_));
 sg13g2_nand2_1 _10196_ (.Y(_02230_),
    .A(_02205_),
    .B(_02225_));
 sg13g2_nand3b_1 _10197_ (.B(_02227_),
    .C(_02044_),
    .Y(_02231_),
    .A_N(_02205_));
 sg13g2_o21ai_1 _10198_ (.B1(_02231_),
    .Y(_02232_),
    .A1(_02044_),
    .A2(_02230_));
 sg13g2_mux2_1 _10199_ (.A0(_02205_),
    .A1(_02230_),
    .S(_01996_),
    .X(_02233_));
 sg13g2_nor2_1 _10200_ (.A(net32),
    .B(_02233_),
    .Y(_02234_));
 sg13g2_a221oi_1 _10201_ (.B2(_01980_),
    .C1(_02234_),
    .B1(_02232_),
    .A1(_02206_),
    .Y(_02235_),
    .A2(_02229_));
 sg13g2_nand2_1 _10202_ (.Y(_02236_),
    .A(_02222_),
    .B(_02235_));
 sg13g2_nand2_1 _10203_ (.Y(_02237_),
    .A(_02221_),
    .B(_02236_));
 sg13g2_a21o_1 _10204_ (.A2(_02218_),
    .A1(net29),
    .B1(_02046_),
    .X(_02238_));
 sg13g2_a21oi_1 _10205_ (.A1(_02206_),
    .A2(_02205_),
    .Y(_02239_),
    .B1(_02218_));
 sg13g2_nand2_1 _10206_ (.Y(_02240_),
    .A(_02205_),
    .B(_02218_));
 sg13g2_o21ai_1 _10207_ (.B1(_02240_),
    .Y(_02241_),
    .A1(_02091_),
    .A2(_02239_));
 sg13g2_a22oi_1 _10208_ (.Y(_02242_),
    .B1(_02241_),
    .B2(_02061_),
    .A2(_02238_),
    .A1(_02091_));
 sg13g2_a21oi_1 _10209_ (.A1(_02206_),
    .A2(_02091_),
    .Y(_02243_),
    .B1(net29));
 sg13g2_xor2_1 _10210_ (.B(_02086_),
    .A(net79),
    .X(_02244_));
 sg13g2_xnor2_1 _10211_ (.Y(_02245_),
    .A(_02243_),
    .B(_02244_));
 sg13g2_o21ai_1 _10212_ (.B1(_02216_),
    .Y(_02246_),
    .A1(_02208_),
    .A2(_02209_));
 sg13g2_nor3_1 _10213_ (.A(_02208_),
    .B(_02209_),
    .C(_02216_),
    .Y(_02247_));
 sg13g2_a21oi_2 _10214_ (.B1(_02247_),
    .Y(_02248_),
    .A2(_02246_),
    .A1(_02213_));
 sg13g2_xnor2_1 _10215_ (.Y(_02249_),
    .A(_02245_),
    .B(_02248_));
 sg13g2_xnor2_1 _10216_ (.Y(_02250_),
    .A(_02242_),
    .B(_02249_));
 sg13g2_nor2b_1 _10217_ (.A(_02237_),
    .B_N(_02250_),
    .Y(_02251_));
 sg13g2_xnor2_1 _10218_ (.Y(_02252_),
    .A(_02080_),
    .B(_02099_));
 sg13g2_xnor2_1 _10219_ (.Y(_02253_),
    .A(_02097_),
    .B(_02252_));
 sg13g2_or2_1 _10220_ (.X(_02254_),
    .B(_02253_),
    .A(_02251_));
 sg13g2_buf_1 _10221_ (.A(_02254_),
    .X(_02255_));
 sg13g2_nor2_1 _10222_ (.A(_02245_),
    .B(_02248_),
    .Y(_02256_));
 sg13g2_nand2_1 _10223_ (.Y(_02257_),
    .A(_02245_),
    .B(_02248_));
 sg13g2_o21ai_1 _10224_ (.B1(_02257_),
    .Y(_02258_),
    .A1(_02242_),
    .A2(_02256_));
 sg13g2_buf_1 _10225_ (.A(_02258_),
    .X(_02259_));
 sg13g2_nand2b_1 _10226_ (.Y(_02260_),
    .B(_02259_),
    .A_N(_02253_));
 sg13g2_nand2_1 _10227_ (.Y(_02261_),
    .A(_02221_),
    .B(_02222_));
 sg13g2_xnor2_1 _10228_ (.Y(_02262_),
    .A(_02235_),
    .B(_02261_));
 sg13g2_or2_1 _10229_ (.X(_02263_),
    .B(_02225_),
    .A(_02044_));
 sg13g2_a22oi_1 _10230_ (.Y(_02264_),
    .B1(_02263_),
    .B2(_01980_),
    .A2(_02225_),
    .A1(_01996_));
 sg13g2_xor2_1 _10231_ (.B(_02227_),
    .A(_02205_),
    .X(_02265_));
 sg13g2_xnor2_1 _10232_ (.Y(_02266_),
    .A(_02264_),
    .B(_02265_));
 sg13g2_nor2_1 _10233_ (.A(_02046_),
    .B(_01997_),
    .Y(_02267_));
 sg13g2_xnor2_1 _10234_ (.Y(_02268_),
    .A(_02223_),
    .B(_02267_));
 sg13g2_nand2_1 _10235_ (.Y(_02269_),
    .A(_02030_),
    .B(net234));
 sg13g2_nand2_1 _10236_ (.Y(_02270_),
    .A(net293),
    .B(net236));
 sg13g2_buf_2 _10237_ (.A(_02270_),
    .X(_02271_));
 sg13g2_nand2_1 _10238_ (.Y(_02272_),
    .A(_02269_),
    .B(_02271_));
 sg13g2_nand2_1 _10239_ (.Y(_02273_),
    .A(net292),
    .B(net233));
 sg13g2_buf_2 _10240_ (.A(_02273_),
    .X(_02274_));
 sg13g2_o21ai_1 _10241_ (.B1(_02274_),
    .Y(_02275_),
    .A1(_02269_),
    .A2(_02271_));
 sg13g2_and2_1 _10242_ (.A(_02272_),
    .B(_02275_),
    .X(_02276_));
 sg13g2_buf_1 _10243_ (.A(_02276_),
    .X(_02277_));
 sg13g2_inv_1 _10244_ (.Y(_02278_),
    .A(_02277_));
 sg13g2_xnor2_1 _10245_ (.Y(_02279_),
    .A(_02165_),
    .B(_02166_));
 sg13g2_xnor2_1 _10246_ (.Y(_02280_),
    .A(_02164_),
    .B(_02279_));
 sg13g2_inv_1 _10247_ (.Y(_02281_),
    .A(_02280_));
 sg13g2_buf_1 _10248_ (.A(net236),
    .X(_02282_));
 sg13g2_nor2_2 _10249_ (.A(net175),
    .B(_01496_),
    .Y(_02283_));
 sg13g2_a21oi_1 _10250_ (.A1(_02277_),
    .A2(_02281_),
    .Y(_02284_),
    .B1(_02283_));
 sg13g2_a21oi_2 _10251_ (.B1(_02284_),
    .Y(_02285_),
    .A2(_02280_),
    .A1(_02278_));
 sg13g2_xor2_1 _10252_ (.B(_01727_),
    .A(_02174_),
    .X(_02286_));
 sg13g2_xnor2_1 _10253_ (.Y(_02287_),
    .A(net290),
    .B(_02286_));
 sg13g2_buf_1 _10254_ (.A(net277),
    .X(_02288_));
 sg13g2_buf_1 _10255_ (.A(net278),
    .X(_02289_));
 sg13g2_buf_1 _10256_ (.A(_02289_),
    .X(_02290_));
 sg13g2_nor2_1 _10257_ (.A(net229),
    .B(net174),
    .Y(_02291_));
 sg13g2_buf_1 _10258_ (.A(_02000_),
    .X(_02292_));
 sg13g2_o21ai_1 _10259_ (.B1(net147),
    .Y(_02293_),
    .A1(_02291_),
    .A2(_02271_));
 sg13g2_nand2_1 _10260_ (.Y(_02294_),
    .A(net182),
    .B(_02293_));
 sg13g2_a21oi_1 _10261_ (.A1(_02030_),
    .A2(_02009_),
    .Y(_02295_),
    .B1(net235));
 sg13g2_a21oi_1 _10262_ (.A1(_01532_),
    .A2(_02274_),
    .Y(_02296_),
    .B1(_02295_));
 sg13g2_nor2_1 _10263_ (.A(_02281_),
    .B(_02296_),
    .Y(_02297_));
 sg13g2_nand2_1 _10264_ (.Y(_02298_),
    .A(_02281_),
    .B(_02296_));
 sg13g2_o21ai_1 _10265_ (.B1(_02298_),
    .Y(_02299_),
    .A1(_02294_),
    .A2(_02297_));
 sg13g2_buf_1 _10266_ (.A(_02299_),
    .X(_02300_));
 sg13g2_xor2_1 _10267_ (.B(_02300_),
    .A(_02287_),
    .X(_02301_));
 sg13g2_xnor2_1 _10268_ (.Y(_02302_),
    .A(_02285_),
    .B(_02301_));
 sg13g2_buf_1 _10269_ (.A(net237),
    .X(_02303_));
 sg13g2_buf_1 _10270_ (.A(net173),
    .X(_02304_));
 sg13g2_nor2_1 _10271_ (.A(net293),
    .B(net146),
    .Y(_02305_));
 sg13g2_a21oi_1 _10272_ (.A1(_01988_),
    .A2(_02305_),
    .Y(_02306_),
    .B1(_01994_));
 sg13g2_nor2_1 _10273_ (.A(net148),
    .B(net238),
    .Y(_02307_));
 sg13g2_nand2_1 _10274_ (.Y(_02308_),
    .A(net284),
    .B(_01988_));
 sg13g2_buf_2 _10275_ (.A(_02308_),
    .X(_02309_));
 sg13g2_xnor2_1 _10276_ (.Y(_02310_),
    .A(net175),
    .B(_02309_));
 sg13g2_o21ai_1 _10277_ (.B1(net246),
    .Y(_02311_),
    .A1(_02307_),
    .A2(_02310_));
 sg13g2_o21ai_1 _10278_ (.B1(_02311_),
    .Y(_02312_),
    .A1(net191),
    .A2(_02306_));
 sg13g2_buf_1 _10279_ (.A(_01992_),
    .X(_02313_));
 sg13g2_nand2_1 _10280_ (.Y(_02314_),
    .A(net173),
    .B(net275));
 sg13g2_a21oi_1 _10281_ (.A1(_01988_),
    .A2(_02314_),
    .Y(_02315_),
    .B1(net293));
 sg13g2_nand2_1 _10282_ (.Y(_02316_),
    .A(net238),
    .B(_02042_));
 sg13g2_nor2_1 _10283_ (.A(net181),
    .B(_01988_),
    .Y(_02317_));
 sg13g2_a21oi_1 _10284_ (.A1(_01988_),
    .A2(_02271_),
    .Y(_02318_),
    .B1(_02317_));
 sg13g2_nor3_1 _10285_ (.A(_02315_),
    .B(_02316_),
    .C(_02318_),
    .Y(_02319_));
 sg13g2_mux2_1 _10286_ (.A0(_02312_),
    .A1(_02319_),
    .S(_01979_),
    .X(_02320_));
 sg13g2_buf_1 _10287_ (.A(_02320_),
    .X(_02321_));
 sg13g2_xnor2_1 _10288_ (.Y(_02322_),
    .A(_02294_),
    .B(_02296_));
 sg13g2_xnor2_1 _10289_ (.Y(_02323_),
    .A(_02280_),
    .B(_02322_));
 sg13g2_nor2_1 _10290_ (.A(_02321_),
    .B(_02323_),
    .Y(_02324_));
 sg13g2_nand2_1 _10291_ (.Y(_02325_),
    .A(net182),
    .B(_01989_));
 sg13g2_nand2_1 _10292_ (.Y(_02326_),
    .A(net238),
    .B(_01994_));
 sg13g2_nor3_1 _10293_ (.A(_01969_),
    .B(_01975_),
    .C(_01976_),
    .Y(_02327_));
 sg13g2_nand2b_1 _10294_ (.Y(_02328_),
    .B(_02327_),
    .A_N(_01946_));
 sg13g2_buf_1 _10295_ (.A(_02328_),
    .X(_02329_));
 sg13g2_mux2_1 _10296_ (.A0(_02042_),
    .A1(_02326_),
    .S(net31),
    .X(_02330_));
 sg13g2_nand3_1 _10297_ (.B(_02325_),
    .C(_02330_),
    .A(net182),
    .Y(_02331_));
 sg13g2_buf_1 _10298_ (.A(net275),
    .X(_02332_));
 sg13g2_buf_1 _10299_ (.A(_02332_),
    .X(_02333_));
 sg13g2_nand2b_1 _10300_ (.Y(_02334_),
    .B(_01594_),
    .A_N(_01779_));
 sg13g2_buf_1 _10301_ (.A(_02334_),
    .X(_02335_));
 sg13g2_nor2_1 _10302_ (.A(net172),
    .B(_02335_),
    .Y(_02336_));
 sg13g2_a21oi_1 _10303_ (.A1(_01989_),
    .A2(_02336_),
    .Y(_02337_),
    .B1(net31));
 sg13g2_a221oi_1 _10304_ (.B2(_02325_),
    .C1(net32),
    .B1(_02326_),
    .A1(_01989_),
    .Y(_02338_),
    .A2(_01994_));
 sg13g2_a21o_1 _10305_ (.A2(_02337_),
    .A1(_02331_),
    .B1(_02338_),
    .X(_02339_));
 sg13g2_nand2_1 _10306_ (.Y(_02340_),
    .A(_02321_),
    .B(_02323_));
 sg13g2_o21ai_1 _10307_ (.B1(_02340_),
    .Y(_02341_),
    .A1(_02324_),
    .A2(_02339_));
 sg13g2_buf_1 _10308_ (.A(_02341_),
    .X(_02342_));
 sg13g2_nand2_1 _10309_ (.Y(_02343_),
    .A(_02224_),
    .B(_02302_));
 sg13g2_o21ai_1 _10310_ (.B1(_02343_),
    .Y(_02344_),
    .A1(_02302_),
    .A2(_02342_));
 sg13g2_mux2_1 _10311_ (.A0(_02224_),
    .A1(_02342_),
    .S(_02302_),
    .X(_02345_));
 sg13g2_nor2_1 _10312_ (.A(_02268_),
    .B(_02345_),
    .Y(_02346_));
 sg13g2_a21oi_2 _10313_ (.B1(_02346_),
    .Y(_02347_),
    .A2(_02344_),
    .A1(_02268_));
 sg13g2_nand2_1 _10314_ (.Y(_02348_),
    .A(_02285_),
    .B(_02300_));
 sg13g2_xnor2_1 _10315_ (.Y(_02349_),
    .A(_02224_),
    .B(_02287_));
 sg13g2_o21ai_1 _10316_ (.B1(_02349_),
    .Y(_02350_),
    .A1(_02285_),
    .A2(_02300_));
 sg13g2_nand2_1 _10317_ (.Y(_02351_),
    .A(_02348_),
    .B(_02350_));
 sg13g2_a21o_1 _10318_ (.A2(_02347_),
    .A1(_02266_),
    .B1(_02351_),
    .X(_02352_));
 sg13g2_o21ai_1 _10319_ (.B1(_02352_),
    .Y(_02353_),
    .A1(_02266_),
    .A2(_02347_));
 sg13g2_nand2_1 _10320_ (.Y(_02354_),
    .A(_02262_),
    .B(_02353_));
 sg13g2_xnor2_1 _10321_ (.Y(_02355_),
    .A(_02266_),
    .B(_02351_));
 sg13g2_xnor2_1 _10322_ (.Y(_02356_),
    .A(_02347_),
    .B(_02355_));
 sg13g2_buf_2 _10323_ (.A(_02356_),
    .X(_02357_));
 sg13g2_inv_1 _10324_ (.Y(_02358_),
    .A(net278));
 sg13g2_nand2_1 _10325_ (.Y(_02359_),
    .A(net282),
    .B(net275));
 sg13g2_buf_1 _10326_ (.A(_02359_),
    .X(_02360_));
 sg13g2_nor2_1 _10327_ (.A(_01492_),
    .B(_01993_),
    .Y(_02361_));
 sg13g2_a21oi_1 _10328_ (.A1(net228),
    .A2(_02361_),
    .Y(_02362_),
    .B1(_01500_));
 sg13g2_a21oi_1 _10329_ (.A1(_02358_),
    .A2(net171),
    .Y(_02363_),
    .B1(_02362_));
 sg13g2_nand2_1 _10330_ (.Y(_02364_),
    .A(net282),
    .B(net237));
 sg13g2_buf_2 _10331_ (.A(_02364_),
    .X(_02365_));
 sg13g2_nand2_1 _10332_ (.Y(_02366_),
    .A(net326),
    .B(_01992_));
 sg13g2_buf_2 _10333_ (.A(_02366_),
    .X(_02367_));
 sg13g2_nand2_1 _10334_ (.Y(_02368_),
    .A(net288),
    .B(net279));
 sg13g2_buf_1 _10335_ (.A(_02368_),
    .X(_02369_));
 sg13g2_xnor2_1 _10336_ (.Y(_02370_),
    .A(_02367_),
    .B(_02369_));
 sg13g2_xnor2_1 _10337_ (.Y(_02371_),
    .A(_02365_),
    .B(_02370_));
 sg13g2_nand2b_1 _10338_ (.Y(_02372_),
    .B(_02371_),
    .A_N(_02363_));
 sg13g2_nor2_1 _10339_ (.A(net171),
    .B(_02371_),
    .Y(_02373_));
 sg13g2_a22oi_1 _10340_ (.Y(_02374_),
    .B1(_02373_),
    .B2(net174),
    .A2(_02372_),
    .A1(net229));
 sg13g2_inv_1 _10341_ (.Y(_02375_),
    .A(_02374_));
 sg13g2_nand2_1 _10342_ (.Y(_02376_),
    .A(net326),
    .B(_01984_));
 sg13g2_buf_2 _10343_ (.A(_02376_),
    .X(_02377_));
 sg13g2_nor3_1 _10344_ (.A(net171),
    .B(_02377_),
    .C(_02371_),
    .Y(_02378_));
 sg13g2_a21oi_2 _10345_ (.B1(_02378_),
    .Y(_02379_),
    .A2(_02375_),
    .A1(net246));
 sg13g2_nand2_1 _10346_ (.Y(_02380_),
    .A(net288),
    .B(net237));
 sg13g2_buf_2 _10347_ (.A(_02380_),
    .X(_02381_));
 sg13g2_nand2_1 _10348_ (.Y(_02382_),
    .A(net234),
    .B(net279));
 sg13g2_buf_2 _10349_ (.A(_02382_),
    .X(_02383_));
 sg13g2_xnor2_1 _10350_ (.Y(_02384_),
    .A(_01725_),
    .B(_02383_));
 sg13g2_nand3_1 _10351_ (.B(net276),
    .C(net236),
    .A(net234),
    .Y(_02385_));
 sg13g2_o21ai_1 _10352_ (.B1(_02385_),
    .Y(_02386_),
    .A1(_02381_),
    .A2(_02384_));
 sg13g2_buf_1 _10353_ (.A(_02386_),
    .X(_02387_));
 sg13g2_nand2_1 _10354_ (.Y(_02388_),
    .A(_02377_),
    .B(_02383_));
 sg13g2_nand2_1 _10355_ (.Y(_02389_),
    .A(net293),
    .B(net278));
 sg13g2_o21ai_1 _10356_ (.B1(_02389_),
    .Y(_02390_),
    .A1(_02377_),
    .A2(_02383_));
 sg13g2_and2_1 _10357_ (.A(_02388_),
    .B(_02390_),
    .X(_02391_));
 sg13g2_buf_1 _10358_ (.A(_02391_),
    .X(_02392_));
 sg13g2_nor2_1 _10359_ (.A(_02387_),
    .B(_02392_),
    .Y(_02393_));
 sg13g2_nand2_1 _10360_ (.Y(_02394_),
    .A(_02387_),
    .B(_02392_));
 sg13g2_o21ai_1 _10361_ (.B1(_02394_),
    .Y(_02395_),
    .A1(_02369_),
    .A2(_02393_));
 sg13g2_nor2b_1 _10362_ (.A(_02379_),
    .B_N(_02395_),
    .Y(_02396_));
 sg13g2_and2_1 _10363_ (.A(net293),
    .B(net227),
    .X(_02397_));
 sg13g2_buf_2 _10364_ (.A(_02397_),
    .X(_02398_));
 sg13g2_a21o_1 _10365_ (.A2(_02369_),
    .A1(_02367_),
    .B1(_02365_),
    .X(_02399_));
 sg13g2_o21ai_1 _10366_ (.B1(_02399_),
    .Y(_02400_),
    .A1(_02367_),
    .A2(_02369_));
 sg13g2_buf_1 _10367_ (.A(_02400_),
    .X(_02401_));
 sg13g2_nand2_1 _10368_ (.Y(_02402_),
    .A(net326),
    .B(net237));
 sg13g2_buf_2 _10369_ (.A(_02402_),
    .X(_02403_));
 sg13g2_nand2_2 _10370_ (.Y(_02404_),
    .A(net232),
    .B(net236));
 sg13g2_xor2_1 _10371_ (.B(_02404_),
    .A(_02403_),
    .X(_02405_));
 sg13g2_nor2_1 _10372_ (.A(net244),
    .B(net277),
    .Y(_02406_));
 sg13g2_xor2_1 _10373_ (.B(_02406_),
    .A(_02405_),
    .X(_02407_));
 sg13g2_xnor2_1 _10374_ (.Y(_02408_),
    .A(_02401_),
    .B(_02407_));
 sg13g2_xnor2_1 _10375_ (.Y(_02409_),
    .A(_02398_),
    .B(_02408_));
 sg13g2_nand2b_1 _10376_ (.Y(_02410_),
    .B(_02379_),
    .A_N(_02395_));
 sg13g2_o21ai_1 _10377_ (.B1(_02410_),
    .Y(_02411_),
    .A1(_02396_),
    .A2(_02409_));
 sg13g2_buf_1 _10378_ (.A(_02411_),
    .X(_02412_));
 sg13g2_nand2_1 _10379_ (.Y(_02413_),
    .A(net293),
    .B(net227));
 sg13g2_buf_2 _10380_ (.A(_02413_),
    .X(_02414_));
 sg13g2_xnor2_1 _10381_ (.Y(_02415_),
    .A(_02369_),
    .B(_02392_));
 sg13g2_xor2_1 _10382_ (.B(_02415_),
    .A(_02387_),
    .X(_02416_));
 sg13g2_nand2_1 _10383_ (.Y(_02417_),
    .A(_01965_),
    .B(_01968_));
 sg13g2_a221oi_1 _10384_ (.B2(_01885_),
    .C1(_02417_),
    .B1(_01745_),
    .A1(net35),
    .Y(_02418_),
    .A2(_01744_));
 sg13g2_nand2_1 _10385_ (.Y(_02419_),
    .A(net171),
    .B(_02381_));
 sg13g2_a221oi_1 _10386_ (.B2(_01966_),
    .C1(_01964_),
    .B1(_01967_),
    .A1(_01951_),
    .Y(_02420_),
    .A2(_01952_));
 sg13g2_buf_1 _10387_ (.A(_02420_),
    .X(_02421_));
 sg13g2_nor2b_1 _10388_ (.A(_02421_),
    .B_N(_02419_),
    .Y(_02422_));
 sg13g2_nand2b_1 _10389_ (.Y(_02423_),
    .B(net35),
    .A_N(_01696_));
 sg13g2_a21oi_1 _10390_ (.A1(_01873_),
    .A2(_01876_),
    .Y(_02424_),
    .B1(_01882_));
 sg13g2_nand2_1 _10391_ (.Y(_02425_),
    .A(_01742_),
    .B(_01741_));
 sg13g2_o21ai_1 _10392_ (.B1(_01742_),
    .Y(_02426_),
    .A1(_01655_),
    .A2(_01657_));
 sg13g2_o21ai_1 _10393_ (.B1(_02426_),
    .Y(_02427_),
    .A1(_02424_),
    .A2(_02425_));
 sg13g2_buf_1 _10394_ (.A(_02427_),
    .X(_02428_));
 sg13g2_and3_1 _10395_ (.X(_02429_),
    .A(_01806_),
    .B(_01842_),
    .C(_01850_));
 sg13g2_buf_2 _10396_ (.A(_02429_),
    .X(_02430_));
 sg13g2_nand2_2 _10397_ (.Y(_02431_),
    .A(net51),
    .B(net61));
 sg13g2_or2_1 _10398_ (.X(_02432_),
    .B(_01804_),
    .A(_01768_));
 sg13g2_buf_2 _10399_ (.A(_02432_),
    .X(_02433_));
 sg13g2_nand2_1 _10400_ (.Y(_02434_),
    .A(_02431_),
    .B(_02433_));
 sg13g2_nor3_2 _10401_ (.A(_02430_),
    .B(_02434_),
    .C(_02425_),
    .Y(_02435_));
 sg13g2_nor3_2 _10402_ (.A(_02423_),
    .B(_02428_),
    .C(_02435_),
    .Y(_02436_));
 sg13g2_nor2_1 _10403_ (.A(net171),
    .B(_02381_),
    .Y(_02437_));
 sg13g2_a221oi_1 _10404_ (.B2(_02436_),
    .C1(_02437_),
    .B1(_02422_),
    .A1(_02418_),
    .Y(_02438_),
    .A2(_02419_));
 sg13g2_buf_1 _10405_ (.A(_02438_),
    .X(_02439_));
 sg13g2_a21o_1 _10406_ (.A2(_01850_),
    .A1(_01842_),
    .B1(_01866_),
    .X(_02440_));
 sg13g2_buf_2 _10407_ (.A(_02440_),
    .X(_02441_));
 sg13g2_a21o_1 _10408_ (.A2(_01736_),
    .A1(_01720_),
    .B1(_01738_),
    .X(_02442_));
 sg13g2_buf_1 _10409_ (.A(_02442_),
    .X(_02443_));
 sg13g2_a21oi_1 _10410_ (.A1(_01878_),
    .A2(_01880_),
    .Y(_02444_),
    .B1(_02443_));
 sg13g2_buf_2 _10411_ (.A(_02444_),
    .X(_02445_));
 sg13g2_nor3_2 _10412_ (.A(_01707_),
    .B(_01717_),
    .C(_01739_),
    .Y(_02446_));
 sg13g2_xnor2_1 _10413_ (.Y(_02447_),
    .A(_01859_),
    .B(_01862_));
 sg13g2_buf_2 _10414_ (.A(_02447_),
    .X(_02448_));
 sg13g2_xnor2_1 _10415_ (.Y(_02449_),
    .A(net62),
    .B(_01695_));
 sg13g2_buf_2 _10416_ (.A(_02449_),
    .X(_02450_));
 sg13g2_nor4_2 _10417_ (.A(_02445_),
    .B(_02446_),
    .C(_02448_),
    .Y(_02451_),
    .D(_02450_));
 sg13g2_o21ai_1 _10418_ (.B1(net90),
    .Y(_02452_),
    .A1(_01899_),
    .A2(_01901_));
 sg13g2_a21oi_2 _10419_ (.B1(_01919_),
    .Y(_02453_),
    .A2(_02452_),
    .A1(_01902_));
 sg13g2_and3_1 _10420_ (.X(_02454_),
    .A(_01919_),
    .B(_01902_),
    .C(_02452_));
 sg13g2_buf_1 _10421_ (.A(_02454_),
    .X(_02455_));
 sg13g2_nor3_1 _10422_ (.A(_01657_),
    .B(_02453_),
    .C(_02455_),
    .Y(_02456_));
 sg13g2_and4_1 _10423_ (.A(_01806_),
    .B(_02441_),
    .C(_02451_),
    .D(_02456_),
    .X(_02457_));
 sg13g2_buf_1 _10424_ (.A(_02457_),
    .X(_02458_));
 sg13g2_a22oi_1 _10425_ (.Y(_02459_),
    .B1(net51),
    .B2(net61),
    .A2(_01695_),
    .A1(net62));
 sg13g2_a22oi_1 _10426_ (.Y(_02460_),
    .B1(_02459_),
    .B2(_01741_),
    .A2(_02446_),
    .A1(_01742_));
 sg13g2_nor4_1 _10427_ (.A(_01696_),
    .B(_01657_),
    .C(_02453_),
    .D(_02455_),
    .Y(_02461_));
 sg13g2_a21o_1 _10428_ (.A2(_01621_),
    .A1(_01619_),
    .B1(_01654_),
    .X(_02462_));
 sg13g2_buf_1 _10429_ (.A(_02462_),
    .X(_02463_));
 sg13g2_nor3_1 _10430_ (.A(_02463_),
    .B(_02453_),
    .C(_02455_),
    .Y(_02464_));
 sg13g2_a21o_1 _10431_ (.A2(_02461_),
    .A1(_02460_),
    .B1(_02464_),
    .X(_02465_));
 sg13g2_buf_1 _10432_ (.A(_02465_),
    .X(_02466_));
 sg13g2_xor2_1 _10433_ (.B(_02453_),
    .A(_01974_),
    .X(_02467_));
 sg13g2_buf_1 _10434_ (.A(_02467_),
    .X(_02468_));
 sg13g2_nand2_1 _10435_ (.Y(_02469_),
    .A(net284),
    .B(net278));
 sg13g2_nand2_1 _10436_ (.Y(_02470_),
    .A(_01486_),
    .B(_01984_));
 sg13g2_xor2_1 _10437_ (.B(_02470_),
    .A(_02367_),
    .X(_02471_));
 sg13g2_xnor2_1 _10438_ (.Y(_02472_),
    .A(_02469_),
    .B(_02471_));
 sg13g2_xnor2_1 _10439_ (.Y(_02473_),
    .A(net284),
    .B(_02365_));
 sg13g2_nand2_1 _10440_ (.Y(_02474_),
    .A(_02472_),
    .B(_02473_));
 sg13g2_nor2_1 _10441_ (.A(net40),
    .B(_02474_),
    .Y(_02475_));
 sg13g2_o21ai_1 _10442_ (.B1(_02475_),
    .Y(_02476_),
    .A1(_02458_),
    .A2(_02466_));
 sg13g2_nand4_1 _10443_ (.B(_02441_),
    .C(_02451_),
    .A(_01806_),
    .Y(_02477_),
    .D(_02456_));
 sg13g2_buf_2 _10444_ (.A(_02477_),
    .X(_02478_));
 sg13g2_a21oi_1 _10445_ (.A1(_02460_),
    .A2(_02461_),
    .Y(_02479_),
    .B1(_02464_));
 sg13g2_buf_1 _10446_ (.A(_02479_),
    .X(_02480_));
 sg13g2_xnor2_1 _10447_ (.Y(_02481_),
    .A(_01974_),
    .B(_02453_));
 sg13g2_buf_1 _10448_ (.A(_02481_),
    .X(_02482_));
 sg13g2_xnor2_1 _10449_ (.Y(_02483_),
    .A(net244),
    .B(_02365_));
 sg13g2_nor2_1 _10450_ (.A(_02472_),
    .B(_02483_),
    .Y(_02484_));
 sg13g2_nand4_1 _10451_ (.B(_02480_),
    .C(_02482_),
    .A(_02478_),
    .Y(_02485_),
    .D(_02484_));
 sg13g2_and2_1 _10452_ (.A(net40),
    .B(_02484_),
    .X(_02486_));
 sg13g2_o21ai_1 _10453_ (.B1(_02486_),
    .Y(_02487_),
    .A1(_02458_),
    .A2(_02466_));
 sg13g2_or4_1 _10454_ (.A(_02458_),
    .B(_02466_),
    .C(_02482_),
    .D(_02474_),
    .X(_02488_));
 sg13g2_and4_1 _10455_ (.A(_02476_),
    .B(_02485_),
    .C(_02487_),
    .D(_02488_),
    .X(_02489_));
 sg13g2_buf_1 _10456_ (.A(_02489_),
    .X(_02490_));
 sg13g2_nor2_1 _10457_ (.A(_02472_),
    .B(_02473_),
    .Y(_02491_));
 sg13g2_nand2_1 _10458_ (.Y(_02492_),
    .A(_02482_),
    .B(_02491_));
 sg13g2_a21oi_1 _10459_ (.A1(_02478_),
    .A2(_02480_),
    .Y(_02493_),
    .B1(_02492_));
 sg13g2_and2_1 _10460_ (.A(_02472_),
    .B(_02483_),
    .X(_02494_));
 sg13g2_and4_1 _10461_ (.A(_02478_),
    .B(_02480_),
    .C(_02482_),
    .D(_02494_),
    .X(_02495_));
 sg13g2_nand2_1 _10462_ (.Y(_02496_),
    .A(net40),
    .B(_02494_));
 sg13g2_a21oi_1 _10463_ (.A1(_02478_),
    .A2(_02480_),
    .Y(_02497_),
    .B1(_02496_));
 sg13g2_and4_1 _10464_ (.A(_02478_),
    .B(_02480_),
    .C(net40),
    .D(_02491_),
    .X(_02498_));
 sg13g2_nor4_2 _10465_ (.A(_02493_),
    .B(_02495_),
    .C(_02497_),
    .Y(_02499_),
    .D(_02498_));
 sg13g2_nand2_1 _10466_ (.Y(_02500_),
    .A(_02490_),
    .B(_02499_));
 sg13g2_xnor2_1 _10467_ (.Y(_02501_),
    .A(_02439_),
    .B(_02500_));
 sg13g2_nor2_1 _10468_ (.A(_02069_),
    .B(_01993_),
    .Y(_02502_));
 sg13g2_buf_2 _10469_ (.A(_02502_),
    .X(_02503_));
 sg13g2_nand2_1 _10470_ (.Y(_02504_),
    .A(_01852_),
    .B(_02433_));
 sg13g2_xor2_1 _10471_ (.B(net61),
    .A(net51),
    .X(_02505_));
 sg13g2_buf_2 _10472_ (.A(_02505_),
    .X(_02506_));
 sg13g2_buf_1 _10473_ (.A(_02506_),
    .X(_02507_));
 sg13g2_nand2b_1 _10474_ (.Y(_02508_),
    .B(_01901_),
    .A_N(_01653_));
 sg13g2_nand2_1 _10475_ (.Y(_02509_),
    .A(_01634_),
    .B(_01653_));
 sg13g2_xor2_1 _10476_ (.B(_01691_),
    .A(net63),
    .X(_02510_));
 sg13g2_and2_1 _10477_ (.A(net90),
    .B(net84),
    .X(_02511_));
 sg13g2_nor2b_1 _10478_ (.A(net63),
    .B_N(_02511_),
    .Y(_02512_));
 sg13g2_nor2_1 _10479_ (.A(net90),
    .B(net84),
    .Y(_02513_));
 sg13g2_and2_1 _10480_ (.A(net63),
    .B(_02513_),
    .X(_02514_));
 sg13g2_mux2_1 _10481_ (.A0(_02512_),
    .A1(_02514_),
    .S(net62),
    .X(_02515_));
 sg13g2_a221oi_1 _10482_ (.B2(_01693_),
    .C1(_02515_),
    .B1(_02510_),
    .A1(_02508_),
    .Y(_02516_),
    .A2(_02509_));
 sg13g2_nor2_1 _10483_ (.A(_01580_),
    .B(_01623_),
    .Y(_02517_));
 sg13g2_nand2_1 _10484_ (.Y(_02518_),
    .A(_01576_),
    .B(_01563_));
 sg13g2_a221oi_1 _10485_ (.B2(_01688_),
    .C1(_01689_),
    .B1(_01682_),
    .A1(_02517_),
    .Y(_02519_),
    .A2(_02518_));
 sg13g2_and2_1 _10486_ (.A(net63),
    .B(_02511_),
    .X(_02520_));
 sg13g2_a221oi_1 _10487_ (.B2(net62),
    .C1(_01654_),
    .B1(_02520_),
    .A1(_02513_),
    .Y(_02521_),
    .A2(_02519_));
 sg13g2_or2_1 _10488_ (.X(_02522_),
    .B(_02521_),
    .A(_02516_));
 sg13g2_nand2b_1 _10489_ (.Y(_02523_),
    .B(net35),
    .A_N(_02460_));
 sg13g2_a22oi_1 _10490_ (.Y(_02524_),
    .B1(_02522_),
    .B2(_02523_),
    .A2(net36),
    .A1(_02504_));
 sg13g2_a21oi_1 _10491_ (.A1(_02445_),
    .A2(_01864_),
    .Y(_02525_),
    .B1(_02521_));
 sg13g2_nand2b_1 _10492_ (.Y(_02526_),
    .B(_02525_),
    .A_N(_02516_));
 sg13g2_a22oi_1 _10493_ (.Y(_02527_),
    .B1(_01871_),
    .B2(net61),
    .A2(_01870_),
    .A1(_01869_));
 sg13g2_nand4_1 _10494_ (.B(_01870_),
    .C(_01871_),
    .A(_01869_),
    .Y(_02528_),
    .D(net61));
 sg13g2_o21ai_1 _10495_ (.B1(_02528_),
    .Y(_02529_),
    .A1(_02443_),
    .A2(_02527_));
 sg13g2_nand3_1 _10496_ (.B(_01621_),
    .C(_01654_),
    .A(_01619_),
    .Y(_02530_));
 sg13g2_a21oi_1 _10497_ (.A1(_02463_),
    .A2(_02530_),
    .Y(_02531_),
    .B1(_02450_));
 sg13g2_and2_1 _10498_ (.A(_02446_),
    .B(_02459_),
    .X(_02532_));
 sg13g2_a22oi_1 _10499_ (.Y(_02533_),
    .B1(_02532_),
    .B2(_01659_),
    .A2(_02531_),
    .A1(_02529_));
 sg13g2_nand2_1 _10500_ (.Y(_02534_),
    .A(_02526_),
    .B(_02533_));
 sg13g2_o21ai_1 _10501_ (.B1(_02451_),
    .Y(_02535_),
    .A1(_02430_),
    .A2(_01866_));
 sg13g2_nor2_1 _10502_ (.A(_02535_),
    .B(net35),
    .Y(_02536_));
 sg13g2_or4_1 _10503_ (.A(_02503_),
    .B(_02524_),
    .C(_02534_),
    .D(_02536_),
    .X(_02537_));
 sg13g2_buf_1 _10504_ (.A(_02537_),
    .X(_02538_));
 sg13g2_nor2_2 _10505_ (.A(_02188_),
    .B(_01991_),
    .Y(_02539_));
 sg13g2_nand2_1 _10506_ (.Y(_02540_),
    .A(net288),
    .B(net275));
 sg13g2_buf_1 _10507_ (.A(_02540_),
    .X(_02541_));
 sg13g2_a21oi_1 _10508_ (.A1(_02526_),
    .A2(_02533_),
    .Y(_02542_),
    .B1(_02541_));
 sg13g2_a221oi_1 _10509_ (.B2(_02523_),
    .C1(_02541_),
    .B1(_02522_),
    .A1(_02504_),
    .Y(_02543_),
    .A2(_02506_));
 sg13g2_nor3_1 _10510_ (.A(_02535_),
    .B(net35),
    .C(_02541_),
    .Y(_02544_));
 sg13g2_or4_1 _10511_ (.A(_02539_),
    .B(_02542_),
    .C(_02543_),
    .D(_02544_),
    .X(_02545_));
 sg13g2_buf_1 _10512_ (.A(_02545_),
    .X(_02546_));
 sg13g2_xor2_1 _10513_ (.B(_02389_),
    .A(_02377_),
    .X(_02547_));
 sg13g2_xnor2_1 _10514_ (.Y(_02548_),
    .A(_02547_),
    .B(_02383_));
 sg13g2_xnor2_1 _10515_ (.Y(_02549_),
    .A(net171),
    .B(_02381_));
 sg13g2_nand3_1 _10516_ (.B(_01745_),
    .C(_02549_),
    .A(_02421_),
    .Y(_02550_));
 sg13g2_nor3_1 _10517_ (.A(_02428_),
    .B(_02435_),
    .C(_02550_),
    .Y(_02551_));
 sg13g2_nand2b_1 _10518_ (.Y(_02552_),
    .B(_02549_),
    .A_N(_02421_));
 sg13g2_a221oi_1 _10519_ (.B2(_01885_),
    .C1(_02552_),
    .B1(_01745_),
    .A1(net35),
    .Y(_02553_),
    .A2(_01744_));
 sg13g2_xor2_1 _10520_ (.B(_02381_),
    .A(net171),
    .X(_02554_));
 sg13g2_nand2_1 _10521_ (.Y(_02555_),
    .A(_02421_),
    .B(_02554_));
 sg13g2_a221oi_1 _10522_ (.B2(_01885_),
    .C1(_02555_),
    .B1(_01745_),
    .A1(net35),
    .Y(_02556_),
    .A2(_01744_));
 sg13g2_nand2b_1 _10523_ (.Y(_02557_),
    .B(_02554_),
    .A_N(_02421_));
 sg13g2_nor4_1 _10524_ (.A(_02423_),
    .B(_02428_),
    .C(_02435_),
    .D(_02557_),
    .Y(_02558_));
 sg13g2_nor4_1 _10525_ (.A(_02551_),
    .B(_02553_),
    .C(_02556_),
    .D(_02558_),
    .Y(_02559_));
 sg13g2_a22oi_1 _10526_ (.Y(_02560_),
    .B1(_02548_),
    .B2(_02559_),
    .A2(_02546_),
    .A1(_02538_));
 sg13g2_nor2_1 _10527_ (.A(_02548_),
    .B(_02559_),
    .Y(_02561_));
 sg13g2_nand2_1 _10528_ (.Y(_02562_),
    .A(_02418_),
    .B(_02419_));
 sg13g2_a21oi_1 _10529_ (.A1(_02436_),
    .A2(_02422_),
    .Y(_02563_),
    .B1(_02437_));
 sg13g2_a221oi_1 _10530_ (.B2(_02499_),
    .C1(_02416_),
    .B1(_02490_),
    .A1(_02562_),
    .Y(_02564_),
    .A2(_02563_));
 sg13g2_inv_1 _10531_ (.Y(_02565_),
    .A(_02416_));
 sg13g2_and4_1 _10532_ (.A(_02565_),
    .B(_02439_),
    .C(_02490_),
    .D(_02499_),
    .X(_02566_));
 sg13g2_nor4_1 _10533_ (.A(_02560_),
    .B(_02561_),
    .C(_02564_),
    .D(_02566_),
    .Y(_02567_));
 sg13g2_a21o_1 _10534_ (.A2(_02501_),
    .A1(_02416_),
    .B1(_02567_),
    .X(_02568_));
 sg13g2_buf_1 _10535_ (.A(_02568_),
    .X(_02569_));
 sg13g2_xor2_1 _10536_ (.B(_02408_),
    .A(_02395_),
    .X(_02570_));
 sg13g2_xnor2_1 _10537_ (.Y(_02571_),
    .A(_02379_),
    .B(_02570_));
 sg13g2_nand3_1 _10538_ (.B(net173),
    .C(net238),
    .A(net232),
    .Y(_02572_));
 sg13g2_xor2_1 _10539_ (.B(_02404_),
    .A(_02309_),
    .X(_02573_));
 sg13g2_nand3_1 _10540_ (.B(_02572_),
    .C(_02573_),
    .A(_02482_),
    .Y(_02574_));
 sg13g2_nand3_1 _10541_ (.B(_02572_),
    .C(_02573_),
    .A(net40),
    .Y(_02575_));
 sg13g2_nand2_1 _10542_ (.Y(_02576_),
    .A(_02478_),
    .B(_02480_));
 sg13g2_buf_8 _10543_ (.A(_02576_),
    .X(_02577_));
 sg13g2_mux2_1 _10544_ (.A0(_02574_),
    .A1(_02575_),
    .S(_02577_),
    .X(_02578_));
 sg13g2_nor2_1 _10545_ (.A(net191),
    .B(_02365_),
    .Y(_02579_));
 sg13g2_xnor2_1 _10546_ (.Y(_02580_),
    .A(_02309_),
    .B(_02404_));
 sg13g2_buf_2 _10547_ (.A(_02580_),
    .X(_02581_));
 sg13g2_nand3_1 _10548_ (.B(_02579_),
    .C(_02581_),
    .A(_02482_),
    .Y(_02582_));
 sg13g2_nand3_1 _10549_ (.B(_02579_),
    .C(_02581_),
    .A(net40),
    .Y(_02583_));
 sg13g2_mux2_1 _10550_ (.A0(_02582_),
    .A1(_02583_),
    .S(_02577_),
    .X(_02584_));
 sg13g2_o21ai_1 _10551_ (.B1(_01613_),
    .Y(_02585_),
    .A1(net284),
    .A2(_02365_));
 sg13g2_nand3_1 _10552_ (.B(_02585_),
    .C(_02581_),
    .A(net40),
    .Y(_02586_));
 sg13g2_nand3_1 _10553_ (.B(_02585_),
    .C(_02581_),
    .A(_02482_),
    .Y(_02587_));
 sg13g2_mux2_1 _10554_ (.A0(_02586_),
    .A1(_02587_),
    .S(_02577_),
    .X(_02588_));
 sg13g2_nor2_1 _10555_ (.A(_02585_),
    .B(_02581_),
    .Y(_02589_));
 sg13g2_o21ai_1 _10556_ (.B1(_02589_),
    .Y(_02590_),
    .A1(_02577_),
    .A2(_02468_));
 sg13g2_nand4_1 _10557_ (.B(_02584_),
    .C(_02588_),
    .A(_02578_),
    .Y(_02591_),
    .D(_02590_));
 sg13g2_a21o_1 _10558_ (.A2(_02469_),
    .A1(_02367_),
    .B1(_02470_),
    .X(_02592_));
 sg13g2_o21ai_1 _10559_ (.B1(_02592_),
    .Y(_02593_),
    .A1(_02367_),
    .A2(_02469_));
 sg13g2_buf_1 _10560_ (.A(_02593_),
    .X(_02594_));
 sg13g2_xnor2_1 _10561_ (.Y(_02595_),
    .A(_01662_),
    .B(_02012_));
 sg13g2_xnor2_1 _10562_ (.Y(_02596_),
    .A(_02594_),
    .B(_02595_));
 sg13g2_xor2_1 _10563_ (.B(_02596_),
    .A(_02403_),
    .X(_02597_));
 sg13g2_xnor2_1 _10564_ (.Y(_02598_),
    .A(net32),
    .B(_02597_));
 sg13g2_xnor2_1 _10565_ (.Y(_02599_),
    .A(_02591_),
    .B(_02598_));
 sg13g2_xnor2_1 _10566_ (.Y(_02600_),
    .A(_02468_),
    .B(_02483_));
 sg13g2_xnor2_1 _10567_ (.Y(_02601_),
    .A(_02577_),
    .B(_02600_));
 sg13g2_nand2_1 _10568_ (.Y(_02602_),
    .A(_02439_),
    .B(_02601_));
 sg13g2_nor2_1 _10569_ (.A(_02439_),
    .B(_02601_),
    .Y(_02603_));
 sg13g2_a21oi_1 _10570_ (.A1(_02472_),
    .A2(_02602_),
    .Y(_02604_),
    .B1(_02603_));
 sg13g2_xnor2_1 _10571_ (.Y(_02605_),
    .A(_02599_),
    .B(_02604_));
 sg13g2_nand2_1 _10572_ (.Y(_02606_),
    .A(_02571_),
    .B(_02605_));
 sg13g2_nor2_1 _10573_ (.A(_02571_),
    .B(_02605_),
    .Y(_02607_));
 sg13g2_a21oi_1 _10574_ (.A1(_02569_),
    .A2(_02606_),
    .Y(_02608_),
    .B1(_02607_));
 sg13g2_o21ai_1 _10575_ (.B1(_02569_),
    .Y(_02609_),
    .A1(_02571_),
    .A2(_02605_));
 sg13g2_and3_1 _10576_ (.X(_02610_),
    .A(_02398_),
    .B(_02606_),
    .C(_02609_));
 sg13g2_a21o_1 _10577_ (.A2(_02608_),
    .A1(_02414_),
    .B1(_02610_),
    .X(_02611_));
 sg13g2_nand2b_1 _10578_ (.Y(_02612_),
    .B(_02398_),
    .A_N(_02412_));
 sg13g2_inv_1 _10579_ (.Y(_02613_),
    .A(_02612_));
 sg13g2_and2_1 _10580_ (.A(_02569_),
    .B(_02613_),
    .X(_02614_));
 sg13g2_nor2_1 _10581_ (.A(_02398_),
    .B(_02412_),
    .Y(_02615_));
 sg13g2_mux2_1 _10582_ (.A0(_02614_),
    .A1(_02615_),
    .S(_02607_),
    .X(_02616_));
 sg13g2_and3_1 _10583_ (.X(_02617_),
    .A(_02569_),
    .B(_02606_),
    .C(_02615_));
 sg13g2_nor2_1 _10584_ (.A(_02606_),
    .B(_02612_),
    .Y(_02618_));
 sg13g2_xnor2_1 _10585_ (.Y(_02619_),
    .A(_02403_),
    .B(_02414_));
 sg13g2_xnor2_1 _10586_ (.Y(_02620_),
    .A(net31),
    .B(_02619_));
 sg13g2_xnor2_1 _10587_ (.Y(_02621_),
    .A(_02591_),
    .B(_02620_));
 sg13g2_nand2_1 _10588_ (.Y(_02622_),
    .A(_02596_),
    .B(_02621_));
 sg13g2_o21ai_1 _10589_ (.B1(_02604_),
    .Y(_02623_),
    .A1(_02596_),
    .A2(_02621_));
 sg13g2_nand2_1 _10590_ (.Y(_02624_),
    .A(_02622_),
    .B(_02623_));
 sg13g2_nor2_1 _10591_ (.A(net238),
    .B(_02365_),
    .Y(_02625_));
 sg13g2_nor2b_1 _10592_ (.A(_02625_),
    .B_N(_01613_),
    .Y(_02626_));
 sg13g2_xnor2_1 _10593_ (.Y(_02627_),
    .A(_02577_),
    .B(net40));
 sg13g2_mux2_1 _10594_ (.A0(_02626_),
    .A1(_02572_),
    .S(_02627_),
    .X(_02628_));
 sg13g2_nand2_1 _10595_ (.Y(_02629_),
    .A(_02628_),
    .B(_02581_));
 sg13g2_nor2_1 _10596_ (.A(_02628_),
    .B(_02581_),
    .Y(_02630_));
 sg13g2_a21oi_2 _10597_ (.B1(_02630_),
    .Y(_02631_),
    .A2(_02620_),
    .A1(_02629_));
 sg13g2_inv_1 _10598_ (.Y(_02632_),
    .A(_02594_));
 sg13g2_a21oi_1 _10599_ (.A1(_02024_),
    .A2(_02632_),
    .Y(_02633_),
    .B1(_01662_));
 sg13g2_a21oi_2 _10600_ (.B1(_02633_),
    .Y(_02634_),
    .A2(_02594_),
    .A1(_02012_));
 sg13g2_xnor2_1 _10601_ (.Y(_02635_),
    .A(_02414_),
    .B(_02405_));
 sg13g2_a21oi_1 _10602_ (.A1(_02401_),
    .A2(_02635_),
    .Y(_02636_),
    .B1(_02406_));
 sg13g2_nor2_1 _10603_ (.A(_02401_),
    .B(_02635_),
    .Y(_02637_));
 sg13g2_nor2_1 _10604_ (.A(_02636_),
    .B(_02637_),
    .Y(_02638_));
 sg13g2_xor2_1 _10605_ (.B(_02638_),
    .A(_02634_),
    .X(_02639_));
 sg13g2_nand2_1 _10606_ (.Y(_02640_),
    .A(net292),
    .B(net236));
 sg13g2_buf_2 _10607_ (.A(_02640_),
    .X(_02641_));
 sg13g2_nand2_1 _10608_ (.Y(_02642_),
    .A(net232),
    .B(net233));
 sg13g2_xor2_1 _10609_ (.B(_02642_),
    .A(_02641_),
    .X(_02643_));
 sg13g2_nand2_1 _10610_ (.Y(_02644_),
    .A(_01981_),
    .B(net230));
 sg13g2_nand2_1 _10611_ (.Y(_02645_),
    .A(net326),
    .B(net232));
 sg13g2_nand2_1 _10612_ (.Y(_02646_),
    .A(_02398_),
    .B(_02405_));
 sg13g2_o21ai_1 _10613_ (.B1(_02646_),
    .Y(_02647_),
    .A1(_02645_),
    .A2(_01729_));
 sg13g2_buf_1 _10614_ (.A(_02647_),
    .X(_02648_));
 sg13g2_xnor2_1 _10615_ (.Y(_02649_),
    .A(_02644_),
    .B(_02648_));
 sg13g2_xnor2_1 _10616_ (.Y(_02650_),
    .A(_02643_),
    .B(_02649_));
 sg13g2_xnor2_1 _10617_ (.Y(_02651_),
    .A(_02639_),
    .B(_02650_));
 sg13g2_nand2_1 _10618_ (.Y(_02652_),
    .A(_02403_),
    .B(_02414_));
 sg13g2_nand2b_1 _10619_ (.Y(_02653_),
    .B(_02398_),
    .A_N(_02403_));
 sg13g2_mux2_1 _10620_ (.A0(_02652_),
    .A1(_02653_),
    .S(_01979_),
    .X(_02654_));
 sg13g2_nor2_1 _10621_ (.A(net244),
    .B(_02003_),
    .Y(_02655_));
 sg13g2_nand2_1 _10622_ (.Y(_02656_),
    .A(net233),
    .B(_02004_));
 sg13g2_o21ai_1 _10623_ (.B1(_02656_),
    .Y(_02657_),
    .A1(net233),
    .A2(_02655_));
 sg13g2_nand4_1 _10624_ (.B(net229),
    .C(net174),
    .A(net238),
    .Y(_02658_),
    .D(_02642_));
 sg13g2_o21ai_1 _10625_ (.B1(_02658_),
    .Y(_02659_),
    .A1(net245),
    .A2(_02657_));
 sg13g2_nand2_1 _10626_ (.Y(_02660_),
    .A(net235),
    .B(net233));
 sg13g2_xnor2_1 _10627_ (.Y(_02661_),
    .A(_02659_),
    .B(_02660_));
 sg13g2_nand2_1 _10628_ (.Y(_02662_),
    .A(net284),
    .B(net227));
 sg13g2_xnor2_1 _10629_ (.Y(_02663_),
    .A(_02309_),
    .B(_02641_));
 sg13g2_xnor2_1 _10630_ (.Y(_02664_),
    .A(_02662_),
    .B(_02663_));
 sg13g2_xnor2_1 _10631_ (.Y(_02665_),
    .A(_02661_),
    .B(_02664_));
 sg13g2_xnor2_1 _10632_ (.Y(_02666_),
    .A(_02654_),
    .B(_02665_));
 sg13g2_xnor2_1 _10633_ (.Y(_02667_),
    .A(_02651_),
    .B(_02666_));
 sg13g2_xnor2_1 _10634_ (.Y(_02668_),
    .A(_02631_),
    .B(_02667_));
 sg13g2_xnor2_1 _10635_ (.Y(_02669_),
    .A(_02624_),
    .B(_02668_));
 sg13g2_nor4_1 _10636_ (.A(_02616_),
    .B(_02617_),
    .C(_02618_),
    .D(_02669_),
    .Y(_02670_));
 sg13g2_a21o_1 _10637_ (.A2(_02611_),
    .A1(_02412_),
    .B1(_02670_),
    .X(_02671_));
 sg13g2_buf_2 _10638_ (.A(_02671_),
    .X(_02672_));
 sg13g2_xnor2_1 _10639_ (.Y(_02673_),
    .A(_02412_),
    .B(_02669_));
 sg13g2_xnor2_1 _10640_ (.Y(_02674_),
    .A(_02611_),
    .B(_02673_));
 sg13g2_nor4_1 _10641_ (.A(_02503_),
    .B(_02524_),
    .C(_02534_),
    .D(_02536_),
    .Y(_02675_));
 sg13g2_nor4_1 _10642_ (.A(_02539_),
    .B(_02542_),
    .C(_02543_),
    .D(_02544_),
    .Y(_02676_));
 sg13g2_xnor2_1 _10643_ (.Y(_02677_),
    .A(_02359_),
    .B(_02547_));
 sg13g2_xnor2_1 _10644_ (.Y(_02678_),
    .A(_02421_),
    .B(_02677_));
 sg13g2_xnor2_1 _10645_ (.Y(_02679_),
    .A(_02436_),
    .B(_02678_));
 sg13g2_nor3_1 _10646_ (.A(_02675_),
    .B(_02676_),
    .C(_02679_),
    .Y(_02680_));
 sg13g2_xor2_1 _10647_ (.B(_02678_),
    .A(_02436_),
    .X(_02681_));
 sg13g2_a21oi_1 _10648_ (.A1(_02538_),
    .A2(_02546_),
    .Y(_02682_),
    .B1(_02681_));
 sg13g2_nand2_2 _10649_ (.Y(_02683_),
    .A(net276),
    .B(net279));
 sg13g2_nand2_1 _10650_ (.Y(_02684_),
    .A(net326),
    .B(net278));
 sg13g2_nand2_1 _10651_ (.Y(_02685_),
    .A(net282),
    .B(net277));
 sg13g2_xor2_1 _10652_ (.B(_02685_),
    .A(_02684_),
    .X(_02686_));
 sg13g2_buf_1 _10653_ (.A(_02686_),
    .X(_02687_));
 sg13g2_nand2b_1 _10654_ (.Y(_02688_),
    .B(_02687_),
    .A_N(_02683_));
 sg13g2_o21ai_1 _10655_ (.B1(_02688_),
    .Y(_02689_),
    .A1(net147),
    .A2(_02645_));
 sg13g2_buf_1 _10656_ (.A(_02689_),
    .X(_02690_));
 sg13g2_nand2_2 _10657_ (.Y(_02691_),
    .A(net234),
    .B(net237));
 sg13g2_a22oi_1 _10658_ (.Y(_02692_),
    .B1(_02539_),
    .B2(_02503_),
    .A2(net236),
    .A1(net276));
 sg13g2_a21oi_1 _10659_ (.A1(_02691_),
    .A2(_02541_),
    .Y(_02693_),
    .B1(_02692_));
 sg13g2_xnor2_1 _10660_ (.Y(_02694_),
    .A(_01725_),
    .B(_02693_));
 sg13g2_nand2_1 _10661_ (.Y(_02695_),
    .A(_02690_),
    .B(_02694_));
 sg13g2_or2_1 _10662_ (.X(_02696_),
    .B(_02694_),
    .A(_02690_));
 sg13g2_nand2_1 _10663_ (.Y(_02697_),
    .A(_02695_),
    .B(_02696_));
 sg13g2_nand2_1 _10664_ (.Y(_02698_),
    .A(net287),
    .B(_01992_));
 sg13g2_buf_2 _10665_ (.A(_02698_),
    .X(_02699_));
 sg13g2_nand2_2 _10666_ (.Y(_02700_),
    .A(net325),
    .B(net280));
 sg13g2_or2_1 _10667_ (.X(_02701_),
    .B(_02700_),
    .A(_02699_));
 sg13g2_buf_1 _10668_ (.A(_02701_),
    .X(_02702_));
 sg13g2_xnor2_1 _10669_ (.Y(_02703_),
    .A(_02445_),
    .B(_02450_));
 sg13g2_nand2_1 _10670_ (.Y(_02704_),
    .A(_02702_),
    .B(_02703_));
 sg13g2_buf_8 _10671_ (.A(_01741_),
    .X(_02705_));
 sg13g2_xnor2_1 _10672_ (.Y(_02706_),
    .A(net39),
    .B(_02450_));
 sg13g2_nand2_1 _10673_ (.Y(_02707_),
    .A(_02702_),
    .B(_02706_));
 sg13g2_o21ai_1 _10674_ (.B1(_02424_),
    .Y(_02708_),
    .A1(_02430_),
    .A2(_02434_));
 sg13g2_buf_1 _10675_ (.A(_02708_),
    .X(_02709_));
 sg13g2_mux2_1 _10676_ (.A0(_02704_),
    .A1(_02707_),
    .S(_02709_),
    .X(_02710_));
 sg13g2_nand2_1 _10677_ (.Y(_02711_),
    .A(_02699_),
    .B(_02700_));
 sg13g2_xnor2_1 _10678_ (.Y(_02712_),
    .A(_02683_),
    .B(_02687_));
 sg13g2_a21oi_1 _10679_ (.A1(_02710_),
    .A2(_02711_),
    .Y(_02713_),
    .B1(_02712_));
 sg13g2_a21oi_1 _10680_ (.A1(net39),
    .A2(_02709_),
    .Y(_02714_),
    .B1(_02450_));
 sg13g2_nor3_2 _10681_ (.A(_01742_),
    .B(_01655_),
    .C(_01657_),
    .Y(_02715_));
 sg13g2_a22oi_1 _10682_ (.Y(_02716_),
    .B1(_02463_),
    .B2(_02530_),
    .A2(_01695_),
    .A1(net62));
 sg13g2_xnor2_1 _10683_ (.Y(_02717_),
    .A(_02691_),
    .B(_02503_));
 sg13g2_nor3_1 _10684_ (.A(_02715_),
    .B(_02716_),
    .C(_02717_),
    .Y(_02718_));
 sg13g2_o21ai_1 _10685_ (.B1(_02717_),
    .Y(_02719_),
    .A1(_02715_),
    .A2(_02716_));
 sg13g2_nand2b_1 _10686_ (.Y(_02720_),
    .B(_02719_),
    .A_N(_02718_));
 sg13g2_xnor2_1 _10687_ (.Y(_02721_),
    .A(_02714_),
    .B(_02720_));
 sg13g2_nand3_1 _10688_ (.B(_02710_),
    .C(_02711_),
    .A(_02712_),
    .Y(_02722_));
 sg13g2_o21ai_1 _10689_ (.B1(_02722_),
    .Y(_02723_),
    .A1(_02713_),
    .A2(_02721_));
 sg13g2_nor4_1 _10690_ (.A(_02680_),
    .B(_02682_),
    .C(_02697_),
    .D(_02723_),
    .Y(_02724_));
 sg13g2_nand3_1 _10691_ (.B(_02546_),
    .C(_02681_),
    .A(_02538_),
    .Y(_02725_));
 sg13g2_buf_1 _10692_ (.A(_02725_),
    .X(_02726_));
 sg13g2_o21ai_1 _10693_ (.B1(_02679_),
    .Y(_02727_),
    .A1(_02675_),
    .A2(_02676_));
 sg13g2_buf_1 _10694_ (.A(_02727_),
    .X(_02728_));
 sg13g2_a221oi_1 _10695_ (.B2(_02696_),
    .C1(_02723_),
    .B1(_02695_),
    .A1(_02726_),
    .Y(_02729_),
    .A2(_02728_));
 sg13g2_inv_1 _10696_ (.Y(_02730_),
    .A(_02697_));
 sg13g2_xor2_1 _10697_ (.B(_02383_),
    .A(_02381_),
    .X(_02731_));
 sg13g2_nor4_1 _10698_ (.A(_02680_),
    .B(_02682_),
    .C(_02730_),
    .D(_02731_),
    .Y(_02732_));
 sg13g2_nand2_1 _10699_ (.Y(_02733_),
    .A(_02730_),
    .B(_02731_));
 sg13g2_a21oi_1 _10700_ (.A1(_02726_),
    .A2(_02728_),
    .Y(_02734_),
    .B1(_02733_));
 sg13g2_nor4_2 _10701_ (.A(_02724_),
    .B(_02729_),
    .C(_02732_),
    .Y(_02735_),
    .D(_02734_));
 sg13g2_a21oi_1 _10702_ (.A1(net174),
    .A2(_02361_),
    .Y(_02736_),
    .B1(net229));
 sg13g2_a21oi_1 _10703_ (.A1(net229),
    .A2(_02363_),
    .Y(_02737_),
    .B1(_02736_));
 sg13g2_nor3_1 _10704_ (.A(net246),
    .B(_01501_),
    .C(net171),
    .Y(_02738_));
 sg13g2_buf_1 _10705_ (.A(net229),
    .X(_02739_));
 sg13g2_a22oi_1 _10706_ (.Y(_02740_),
    .B1(_02738_),
    .B2(net170),
    .A2(_02737_),
    .A1(net246));
 sg13g2_xor2_1 _10707_ (.B(_02740_),
    .A(_02371_),
    .X(_02741_));
 sg13g2_inv_1 _10708_ (.Y(_02742_),
    .A(_01984_));
 sg13g2_nor2_2 _10709_ (.A(_02742_),
    .B(_02358_),
    .Y(_02743_));
 sg13g2_and2_1 _10710_ (.A(net326),
    .B(net282),
    .X(_02744_));
 sg13g2_buf_1 _10711_ (.A(_02744_),
    .X(_02745_));
 sg13g2_xnor2_1 _10712_ (.Y(_02746_),
    .A(_01487_),
    .B(net172));
 sg13g2_nand3_1 _10713_ (.B(_02745_),
    .C(_02746_),
    .A(_02743_),
    .Y(_02747_));
 sg13g2_xnor2_1 _10714_ (.Y(_02748_),
    .A(_01725_),
    .B(_02731_));
 sg13g2_a21o_1 _10715_ (.A2(_02693_),
    .A1(_02690_),
    .B1(_02748_),
    .X(_02749_));
 sg13g2_o21ai_1 _10716_ (.B1(_02749_),
    .Y(_02750_),
    .A1(_02690_),
    .A2(_02693_));
 sg13g2_nor2_1 _10717_ (.A(_02747_),
    .B(_02750_),
    .Y(_02751_));
 sg13g2_nand2_1 _10718_ (.Y(_02752_),
    .A(_02747_),
    .B(_02750_));
 sg13g2_nor2b_1 _10719_ (.A(_02751_),
    .B_N(_02752_),
    .Y(_02753_));
 sg13g2_xnor2_1 _10720_ (.Y(_02754_),
    .A(_02741_),
    .B(_02753_));
 sg13g2_nor2_1 _10721_ (.A(_02560_),
    .B(_02561_),
    .Y(_02755_));
 sg13g2_xnor2_1 _10722_ (.Y(_02756_),
    .A(_02755_),
    .B(_02565_));
 sg13g2_xnor2_1 _10723_ (.Y(_02757_),
    .A(_02501_),
    .B(_02756_));
 sg13g2_nor2_1 _10724_ (.A(_02754_),
    .B(_02757_),
    .Y(_02758_));
 sg13g2_nand2_1 _10725_ (.Y(_02759_),
    .A(_02754_),
    .B(_02757_));
 sg13g2_o21ai_1 _10726_ (.B1(_02759_),
    .Y(_02760_),
    .A1(_02735_),
    .A2(_02758_));
 sg13g2_a21o_1 _10727_ (.A2(_02752_),
    .A1(_02741_),
    .B1(_02751_),
    .X(_02761_));
 sg13g2_xnor2_1 _10728_ (.Y(_02762_),
    .A(_02571_),
    .B(_02605_));
 sg13g2_xnor2_1 _10729_ (.Y(_02763_),
    .A(_02569_),
    .B(_02762_));
 sg13g2_nor2_1 _10730_ (.A(_02761_),
    .B(_02763_),
    .Y(_02764_));
 sg13g2_nand2_1 _10731_ (.Y(_02765_),
    .A(_02761_),
    .B(_02763_));
 sg13g2_o21ai_1 _10732_ (.B1(_02765_),
    .Y(_02766_),
    .A1(_02760_),
    .A2(_02764_));
 sg13g2_nand2_1 _10733_ (.Y(_02767_),
    .A(_02674_),
    .B(_02766_));
 sg13g2_buf_2 _10734_ (.A(_02767_),
    .X(_02768_));
 sg13g2_nand2_1 _10735_ (.Y(_02769_),
    .A(_02672_),
    .B(_02768_));
 sg13g2_buf_1 _10736_ (.A(net172),
    .X(_02770_));
 sg13g2_and2_1 _10737_ (.A(net246),
    .B(net146),
    .X(_02771_));
 sg13g2_buf_1 _10738_ (.A(_02771_),
    .X(_02772_));
 sg13g2_nand3_1 _10739_ (.B(net32),
    .C(_02772_),
    .A(net145),
    .Y(_02773_));
 sg13g2_nand2_1 _10740_ (.Y(_02774_),
    .A(net293),
    .B(net173));
 sg13g2_buf_2 _10741_ (.A(_02774_),
    .X(_02775_));
 sg13g2_nand3_1 _10742_ (.B(net31),
    .C(_02775_),
    .A(net230),
    .Y(_02776_));
 sg13g2_xnor2_1 _10743_ (.Y(_02777_),
    .A(net146),
    .B(net227));
 sg13g2_xnor2_1 _10744_ (.Y(_02778_),
    .A(_01988_),
    .B(_02777_));
 sg13g2_nand4_1 _10745_ (.B(_02773_),
    .C(_02776_),
    .A(net182),
    .Y(_02779_),
    .D(_02778_));
 sg13g2_o21ai_1 _10746_ (.B1(net182),
    .Y(_02780_),
    .A1(net145),
    .A2(_02778_));
 sg13g2_nand3_1 _10747_ (.B(_02775_),
    .C(_02780_),
    .A(net31),
    .Y(_02781_));
 sg13g2_or4_1 _10748_ (.A(net31),
    .B(_02775_),
    .C(_02662_),
    .D(_02778_),
    .X(_02782_));
 sg13g2_and3_1 _10749_ (.X(_02783_),
    .A(_02779_),
    .B(_02781_),
    .C(_02782_));
 sg13g2_buf_1 _10750_ (.A(_02783_),
    .X(_02784_));
 sg13g2_xnor2_1 _10751_ (.Y(_02785_),
    .A(_02775_),
    .B(_02662_));
 sg13g2_buf_2 _10752_ (.A(_02785_),
    .X(_02786_));
 sg13g2_nor2_1 _10753_ (.A(_02663_),
    .B(_02403_),
    .Y(_02787_));
 sg13g2_a21oi_1 _10754_ (.A1(net31),
    .A2(_02786_),
    .Y(_02788_),
    .B1(_02787_));
 sg13g2_nand3b_1 _10755_ (.B(_02327_),
    .C(_02786_),
    .Y(_02789_),
    .A_N(_01946_));
 sg13g2_nor2_1 _10756_ (.A(_02786_),
    .B(_02652_),
    .Y(_02790_));
 sg13g2_o21ai_1 _10757_ (.B1(_02790_),
    .Y(_02791_),
    .A1(_01946_),
    .A2(_01978_));
 sg13g2_xor2_1 _10758_ (.B(_02641_),
    .A(_02309_),
    .X(_02792_));
 sg13g2_nor2_1 _10759_ (.A(_02786_),
    .B(_02792_),
    .Y(_02793_));
 sg13g2_o21ai_1 _10760_ (.B1(_02793_),
    .Y(_02794_),
    .A1(_01946_),
    .A2(_01978_));
 sg13g2_nor2_1 _10761_ (.A(_02786_),
    .B(_02398_),
    .Y(_02795_));
 sg13g2_o21ai_1 _10762_ (.B1(_02663_),
    .Y(_02796_),
    .A1(_02403_),
    .A2(_02795_));
 sg13g2_nand4_1 _10763_ (.B(_02791_),
    .C(_02794_),
    .A(_02789_),
    .Y(_02797_),
    .D(_02796_));
 sg13g2_o21ai_1 _10764_ (.B1(_02797_),
    .Y(_02798_),
    .A1(_02414_),
    .A2(_02788_));
 sg13g2_o21ai_1 _10765_ (.B1(net147),
    .Y(_02799_),
    .A1(_02291_),
    .A2(_02641_));
 sg13g2_nand2_2 _10766_ (.Y(_02800_),
    .A(net238),
    .B(_02799_));
 sg13g2_nor2_2 _10767_ (.A(_02069_),
    .B(_02009_),
    .Y(_02801_));
 sg13g2_xor2_1 _10768_ (.B(_02801_),
    .A(_02800_),
    .X(_02802_));
 sg13g2_inv_1 _10769_ (.Y(_02803_),
    .A(_02802_));
 sg13g2_nor2_1 _10770_ (.A(_02403_),
    .B(_02414_),
    .Y(_02804_));
 sg13g2_o21ai_1 _10771_ (.B1(_02792_),
    .Y(_02805_),
    .A1(net31),
    .A2(_02804_));
 sg13g2_nor2_1 _10772_ (.A(_02792_),
    .B(_02804_),
    .Y(_02806_));
 sg13g2_o21ai_1 _10773_ (.B1(_02802_),
    .Y(_02807_),
    .A1(_02786_),
    .A2(_02806_));
 sg13g2_a21oi_1 _10774_ (.A1(_02329_),
    .A2(_02652_),
    .Y(_02808_),
    .B1(_02807_));
 sg13g2_and2_1 _10775_ (.A(_02792_),
    .B(_02652_),
    .X(_02809_));
 sg13g2_nor4_1 _10776_ (.A(net32),
    .B(_02786_),
    .C(_02803_),
    .D(_02809_),
    .Y(_02810_));
 sg13g2_a221oi_1 _10777_ (.B2(_02808_),
    .C1(_02810_),
    .B1(_02805_),
    .A1(_02798_),
    .Y(_02811_),
    .A2(_02803_));
 sg13g2_xnor2_1 _10778_ (.Y(_02812_),
    .A(_02784_),
    .B(_02811_));
 sg13g2_a22oi_1 _10779_ (.Y(_02813_),
    .B1(_02659_),
    .B2(net235),
    .A2(_02004_),
    .A1(net177));
 sg13g2_nor2b_1 _10780_ (.A(_02813_),
    .B_N(net178),
    .Y(_02814_));
 sg13g2_a21o_1 _10781_ (.A2(_02775_),
    .A1(_02641_),
    .B1(_02642_),
    .X(_02815_));
 sg13g2_o21ai_1 _10782_ (.B1(_02815_),
    .Y(_02816_),
    .A1(_02641_),
    .A2(_02775_));
 sg13g2_buf_1 _10783_ (.A(_02816_),
    .X(_02817_));
 sg13g2_xor2_1 _10784_ (.B(_02817_),
    .A(_02335_),
    .X(_02818_));
 sg13g2_xnor2_1 _10785_ (.Y(_02819_),
    .A(_02775_),
    .B(_02643_));
 sg13g2_nor2_1 _10786_ (.A(_02648_),
    .B(_02819_),
    .Y(_02820_));
 sg13g2_nand2_1 _10787_ (.Y(_02821_),
    .A(_02648_),
    .B(_02819_));
 sg13g2_o21ai_1 _10788_ (.B1(_02821_),
    .Y(_02822_),
    .A1(_02644_),
    .A2(_02820_));
 sg13g2_buf_1 _10789_ (.A(_02822_),
    .X(_02823_));
 sg13g2_xor2_1 _10790_ (.B(_02823_),
    .A(_02818_),
    .X(_02824_));
 sg13g2_xnor2_1 _10791_ (.Y(_02825_),
    .A(_02814_),
    .B(_02824_));
 sg13g2_inv_1 _10792_ (.Y(_02826_),
    .A(_02825_));
 sg13g2_xnor2_1 _10793_ (.Y(_02827_),
    .A(_02786_),
    .B(_02792_));
 sg13g2_xnor2_1 _10794_ (.Y(_02828_),
    .A(_02654_),
    .B(_02827_));
 sg13g2_nor2_1 _10795_ (.A(_02828_),
    .B(_02661_),
    .Y(_02829_));
 sg13g2_nand2_1 _10796_ (.Y(_02830_),
    .A(_02828_),
    .B(_02661_));
 sg13g2_o21ai_1 _10797_ (.B1(_02830_),
    .Y(_02831_),
    .A1(_02829_),
    .A2(_02631_));
 sg13g2_buf_1 _10798_ (.A(_02831_),
    .X(_02832_));
 sg13g2_xnor2_1 _10799_ (.Y(_02833_),
    .A(_02826_),
    .B(_02832_));
 sg13g2_xnor2_1 _10800_ (.Y(_02834_),
    .A(_02812_),
    .B(_02833_));
 sg13g2_buf_1 _10801_ (.A(_02834_),
    .X(_02835_));
 sg13g2_nor2b_1 _10802_ (.A(_02634_),
    .B_N(_02638_),
    .Y(_02836_));
 sg13g2_xor2_1 _10803_ (.B(_02649_),
    .A(_02819_),
    .X(_02837_));
 sg13g2_nand2b_1 _10804_ (.Y(_02838_),
    .B(_02634_),
    .A_N(_02638_));
 sg13g2_o21ai_1 _10805_ (.B1(_02838_),
    .Y(_02839_),
    .A1(_02836_),
    .A2(_02837_));
 sg13g2_buf_2 _10806_ (.A(_02839_),
    .X(_02840_));
 sg13g2_nor2b_1 _10807_ (.A(_02624_),
    .B_N(_02668_),
    .Y(_02841_));
 sg13g2_and2_1 _10808_ (.A(_02772_),
    .B(_02651_),
    .X(_02842_));
 sg13g2_nor2_1 _10809_ (.A(_02772_),
    .B(_02651_),
    .Y(_02843_));
 sg13g2_xnor2_1 _10810_ (.Y(_02844_),
    .A(_02631_),
    .B(_02666_));
 sg13g2_mux2_1 _10811_ (.A0(_02842_),
    .A1(_02843_),
    .S(_02844_),
    .X(_02845_));
 sg13g2_nor2_1 _10812_ (.A(_02841_),
    .B(_02845_),
    .Y(_02846_));
 sg13g2_buf_1 _10813_ (.A(_02846_),
    .X(_02847_));
 sg13g2_or2_1 _10814_ (.X(_02848_),
    .B(_02847_),
    .A(_02840_));
 sg13g2_buf_1 _10815_ (.A(_02848_),
    .X(_02849_));
 sg13g2_xor2_1 _10816_ (.B(_02271_),
    .A(_02269_),
    .X(_02850_));
 sg13g2_xnor2_1 _10817_ (.Y(_02851_),
    .A(_02274_),
    .B(_02850_));
 sg13g2_xnor2_1 _10818_ (.Y(_02852_),
    .A(_02851_),
    .B(_02818_));
 sg13g2_a21o_1 _10819_ (.A2(_02823_),
    .A1(_02814_),
    .B1(_02852_),
    .X(_02853_));
 sg13g2_o21ai_1 _10820_ (.B1(_02853_),
    .Y(_02854_),
    .A1(_02814_),
    .A2(_02823_));
 sg13g2_buf_1 _10821_ (.A(_02854_),
    .X(_02855_));
 sg13g2_xnor2_1 _10822_ (.Y(_02856_),
    .A(_02271_),
    .B(_02784_));
 sg13g2_a21oi_1 _10823_ (.A1(net232),
    .A2(net179),
    .Y(_02857_),
    .B1(_02801_));
 sg13g2_xor2_1 _10824_ (.B(_02857_),
    .A(_02274_),
    .X(_02858_));
 sg13g2_xnor2_1 _10825_ (.Y(_02859_),
    .A(_02800_),
    .B(_02858_));
 sg13g2_nand2_1 _10826_ (.Y(_02860_),
    .A(_02859_),
    .B(_02798_));
 sg13g2_nor2_1 _10827_ (.A(_02859_),
    .B(_02798_),
    .Y(_02861_));
 sg13g2_a21oi_1 _10828_ (.A1(_02856_),
    .A2(_02860_),
    .Y(_02862_),
    .B1(_02861_));
 sg13g2_xnor2_1 _10829_ (.Y(_02863_),
    .A(_02321_),
    .B(_02322_));
 sg13g2_xor2_1 _10830_ (.B(_02863_),
    .A(_02339_),
    .X(_02864_));
 sg13g2_nor3_1 _10831_ (.A(net235),
    .B(net179),
    .C(_02274_),
    .Y(_02865_));
 sg13g2_a21oi_1 _10832_ (.A1(net235),
    .A2(_02274_),
    .Y(_02866_),
    .B1(_02865_));
 sg13g2_xnor2_1 _10833_ (.Y(_02867_),
    .A(net245),
    .B(_02274_));
 sg13g2_nand2_1 _10834_ (.Y(_02868_),
    .A(net235),
    .B(_02867_));
 sg13g2_o21ai_1 _10835_ (.B1(_02868_),
    .Y(_02869_),
    .A1(_02800_),
    .A2(_02867_));
 sg13g2_nand2_1 _10836_ (.Y(_02870_),
    .A(net179),
    .B(_02869_));
 sg13g2_o21ai_1 _10837_ (.B1(_02870_),
    .Y(_02871_),
    .A1(_02800_),
    .A2(_02866_));
 sg13g2_buf_1 _10838_ (.A(_02871_),
    .X(_02872_));
 sg13g2_nor2_1 _10839_ (.A(_02817_),
    .B(_02851_),
    .Y(_02873_));
 sg13g2_nand2_1 _10840_ (.Y(_02874_),
    .A(_02817_),
    .B(_02851_));
 sg13g2_o21ai_1 _10841_ (.B1(_02874_),
    .Y(_02875_),
    .A1(_02335_),
    .A2(_02873_));
 sg13g2_buf_1 _10842_ (.A(_02875_),
    .X(_02876_));
 sg13g2_xnor2_1 _10843_ (.Y(_02877_),
    .A(_02277_),
    .B(_02283_));
 sg13g2_xnor2_1 _10844_ (.Y(_02878_),
    .A(_02876_),
    .B(_02877_));
 sg13g2_xnor2_1 _10845_ (.Y(_02879_),
    .A(_02872_),
    .B(_02878_));
 sg13g2_xor2_1 _10846_ (.B(_02879_),
    .A(_02864_),
    .X(_02880_));
 sg13g2_xor2_1 _10847_ (.B(_02880_),
    .A(_02862_),
    .X(_02881_));
 sg13g2_xor2_1 _10848_ (.B(_02881_),
    .A(_02855_),
    .X(_02882_));
 sg13g2_nand2_1 _10849_ (.Y(_02883_),
    .A(_02825_),
    .B(_02832_));
 sg13g2_o21ai_1 _10850_ (.B1(_02812_),
    .Y(_02884_),
    .A1(_02825_),
    .A2(_02832_));
 sg13g2_nand2_1 _10851_ (.Y(_02885_),
    .A(_02883_),
    .B(_02884_));
 sg13g2_nor2_1 _10852_ (.A(_02826_),
    .B(_02832_),
    .Y(_02886_));
 sg13g2_nand2_1 _10853_ (.Y(_02887_),
    .A(_02826_),
    .B(_02832_));
 sg13g2_o21ai_1 _10854_ (.B1(_02887_),
    .Y(_02888_),
    .A1(_02812_),
    .A2(_02886_));
 sg13g2_mux2_1 _10855_ (.A0(_02885_),
    .A1(_02888_),
    .S(_02851_),
    .X(_02889_));
 sg13g2_xnor2_1 _10856_ (.Y(_02890_),
    .A(_02882_),
    .B(_02889_));
 sg13g2_buf_1 _10857_ (.A(_02890_),
    .X(_02891_));
 sg13g2_o21ai_1 _10858_ (.B1(net24),
    .Y(_02892_),
    .A1(net26),
    .A2(_02849_));
 sg13g2_inv_1 _10859_ (.Y(_02893_),
    .A(net26));
 sg13g2_xor2_1 _10860_ (.B(_02847_),
    .A(_02840_),
    .X(_02894_));
 sg13g2_a21o_1 _10861_ (.A2(_02847_),
    .A1(_02840_),
    .B1(net26),
    .X(_02895_));
 sg13g2_o21ai_1 _10862_ (.B1(_02895_),
    .Y(_02896_),
    .A1(_02893_),
    .A2(_02894_));
 sg13g2_nand2b_1 _10863_ (.Y(_02897_),
    .B(_02896_),
    .A_N(net24));
 sg13g2_nand3_1 _10864_ (.B(_02892_),
    .C(_02897_),
    .A(_02769_),
    .Y(_02898_));
 sg13g2_inv_1 _10865_ (.Y(_02899_),
    .A(net24));
 sg13g2_nor2_1 _10866_ (.A(_02672_),
    .B(_02768_),
    .Y(_02900_));
 sg13g2_and2_1 _10867_ (.A(_02849_),
    .B(_02895_),
    .X(_02901_));
 sg13g2_buf_1 _10868_ (.A(_02901_),
    .X(_02902_));
 sg13g2_inv_1 _10869_ (.Y(_02903_),
    .A(_02902_));
 sg13g2_o21ai_1 _10870_ (.B1(_02903_),
    .Y(_02904_),
    .A1(_02899_),
    .A2(_02900_));
 sg13g2_nand2_1 _10871_ (.Y(_02905_),
    .A(_02835_),
    .B(_02840_));
 sg13g2_nor2_1 _10872_ (.A(net24),
    .B(_02905_),
    .Y(_02906_));
 sg13g2_nand2_1 _10873_ (.Y(_02907_),
    .A(_02900_),
    .B(_02906_));
 sg13g2_nand3_1 _10874_ (.B(_02904_),
    .C(_02907_),
    .A(_02898_),
    .Y(_02908_));
 sg13g2_nor2b_1 _10875_ (.A(_02880_),
    .B_N(_02862_),
    .Y(_02909_));
 sg13g2_nand2_1 _10876_ (.Y(_02910_),
    .A(_02281_),
    .B(_02879_));
 sg13g2_nand3b_1 _10877_ (.B(_02280_),
    .C(_02864_),
    .Y(_02911_),
    .A_N(_02879_));
 sg13g2_o21ai_1 _10878_ (.B1(_02911_),
    .Y(_02912_),
    .A1(_02864_),
    .A2(_02910_));
 sg13g2_nor2_1 _10879_ (.A(_02909_),
    .B(_02912_),
    .Y(_02913_));
 sg13g2_xor2_1 _10880_ (.B(_02302_),
    .A(_02268_),
    .X(_02914_));
 sg13g2_xnor2_1 _10881_ (.Y(_02915_),
    .A(_02342_),
    .B(_02914_));
 sg13g2_nand2_1 _10882_ (.Y(_02916_),
    .A(_02872_),
    .B(_02876_));
 sg13g2_xnor2_1 _10883_ (.Y(_02917_),
    .A(_02281_),
    .B(_02877_));
 sg13g2_o21ai_1 _10884_ (.B1(_02917_),
    .Y(_02918_),
    .A1(_02872_),
    .A2(_02876_));
 sg13g2_nand2_1 _10885_ (.Y(_02919_),
    .A(_02916_),
    .B(_02918_));
 sg13g2_xor2_1 _10886_ (.B(_02919_),
    .A(_02915_),
    .X(_02920_));
 sg13g2_xnor2_1 _10887_ (.Y(_02921_),
    .A(_02913_),
    .B(_02920_));
 sg13g2_buf_1 _10888_ (.A(_02921_),
    .X(_02922_));
 sg13g2_xnor2_1 _10889_ (.Y(_02923_),
    .A(_02699_),
    .B(_02700_));
 sg13g2_nand2_1 _10890_ (.Y(_02924_),
    .A(_02703_),
    .B(_02923_));
 sg13g2_nand2_1 _10891_ (.Y(_02925_),
    .A(_02706_),
    .B(_02923_));
 sg13g2_mux2_1 _10892_ (.A0(_02924_),
    .A1(_02925_),
    .S(_01885_),
    .X(_02926_));
 sg13g2_xor2_1 _10893_ (.B(_02700_),
    .A(_02699_),
    .X(_02927_));
 sg13g2_nand2_1 _10894_ (.Y(_02928_),
    .A(_02703_),
    .B(_02927_));
 sg13g2_nand2_1 _10895_ (.Y(_02929_),
    .A(_02706_),
    .B(_02927_));
 sg13g2_mux2_1 _10896_ (.A0(_02928_),
    .A1(_02929_),
    .S(_02709_),
    .X(_02930_));
 sg13g2_nand2_1 _10897_ (.Y(_02931_),
    .A(_02926_),
    .B(_02930_));
 sg13g2_nand2_1 _10898_ (.Y(_02932_),
    .A(net288),
    .B(_01984_));
 sg13g2_buf_1 _10899_ (.A(_02932_),
    .X(_02933_));
 sg13g2_nand2_2 _10900_ (.Y(_02934_),
    .A(net282),
    .B(_01986_));
 sg13g2_xor2_1 _10901_ (.B(_02934_),
    .A(_02933_),
    .X(_02935_));
 sg13g2_xnor2_1 _10902_ (.Y(_02936_),
    .A(_02002_),
    .B(_02935_));
 sg13g2_o21ai_1 _10903_ (.B1(_02443_),
    .Y(_02937_),
    .A1(_01707_),
    .A2(_01717_));
 sg13g2_buf_2 _10904_ (.A(_02937_),
    .X(_02938_));
 sg13g2_nand3_1 _10905_ (.B(_01880_),
    .C(_01739_),
    .A(_01878_),
    .Y(_02939_));
 sg13g2_buf_2 _10906_ (.A(_02939_),
    .X(_02940_));
 sg13g2_and2_1 _10907_ (.A(net325),
    .B(_01992_),
    .X(_02941_));
 sg13g2_buf_2 _10908_ (.A(_02941_),
    .X(_02942_));
 sg13g2_nand4_1 _10909_ (.B(_02940_),
    .C(_02506_),
    .A(_02938_),
    .Y(_02943_),
    .D(_02942_));
 sg13g2_nor2_1 _10910_ (.A(_01823_),
    .B(_01991_),
    .Y(_02944_));
 sg13g2_nand4_1 _10911_ (.B(_02938_),
    .C(_02940_),
    .A(_02944_),
    .Y(_02945_),
    .D(_02506_));
 sg13g2_a22oi_1 _10912_ (.Y(_02946_),
    .B1(_02943_),
    .B2(_02945_),
    .A2(_02433_),
    .A1(_01852_));
 sg13g2_nand3_1 _10913_ (.B(_01880_),
    .C(_02443_),
    .A(_01878_),
    .Y(_02947_));
 sg13g2_buf_1 _10914_ (.A(_02947_),
    .X(_02948_));
 sg13g2_nand4_1 _10915_ (.B(_02431_),
    .C(net38),
    .A(_01741_),
    .Y(_02949_),
    .D(_02942_));
 sg13g2_nand4_1 _10916_ (.B(_01741_),
    .C(_02431_),
    .A(_02944_),
    .Y(_02950_),
    .D(net38));
 sg13g2_a22oi_1 _10917_ (.Y(_02951_),
    .B1(_02949_),
    .B2(_02950_),
    .A2(_02441_),
    .A1(_01806_));
 sg13g2_nand2_1 _10918_ (.Y(_02952_),
    .A(net325),
    .B(_01992_));
 sg13g2_buf_2 _10919_ (.A(_02952_),
    .X(_02953_));
 sg13g2_nor2_1 _10920_ (.A(_01729_),
    .B(_02953_),
    .Y(_02954_));
 sg13g2_nor3_1 _10921_ (.A(net51),
    .B(net61),
    .C(_02953_),
    .Y(_02955_));
 sg13g2_nand3_1 _10922_ (.B(net38),
    .C(_02955_),
    .A(net39),
    .Y(_02956_));
 sg13g2_nand4_1 _10923_ (.B(_02938_),
    .C(_02940_),
    .A(_01864_),
    .Y(_02957_),
    .D(_02942_));
 sg13g2_nor3_1 _10924_ (.A(_01729_),
    .B(net51),
    .C(net61),
    .Y(_02958_));
 sg13g2_nand3_1 _10925_ (.B(net38),
    .C(_02958_),
    .A(net39),
    .Y(_02959_));
 sg13g2_nand4_1 _10926_ (.B(_01864_),
    .C(_02938_),
    .A(_02944_),
    .Y(_02960_),
    .D(_02940_));
 sg13g2_nand4_1 _10927_ (.B(_02957_),
    .C(_02959_),
    .A(_02956_),
    .Y(_02961_),
    .D(_02960_));
 sg13g2_nor4_1 _10928_ (.A(_02946_),
    .B(_02951_),
    .C(_02954_),
    .D(_02961_),
    .Y(_02962_));
 sg13g2_buf_2 _10929_ (.A(_02962_),
    .X(_02963_));
 sg13g2_nor2_1 _10930_ (.A(_02936_),
    .B(_02963_),
    .Y(_02964_));
 sg13g2_nand2_1 _10931_ (.Y(_02965_),
    .A(_02936_),
    .B(_02963_));
 sg13g2_o21ai_1 _10932_ (.B1(_02965_),
    .Y(_02966_),
    .A1(_02931_),
    .A2(_02964_));
 sg13g2_buf_2 _10933_ (.A(_02966_),
    .X(_02967_));
 sg13g2_nand2_1 _10934_ (.Y(_02968_),
    .A(_02933_),
    .B(_02934_));
 sg13g2_xor2_1 _10935_ (.B(_02968_),
    .A(net276),
    .X(_02969_));
 sg13g2_nor2_1 _10936_ (.A(_02933_),
    .B(_02934_),
    .Y(_02970_));
 sg13g2_mux2_1 _10937_ (.A0(_02969_),
    .A1(_02970_),
    .S(_01823_),
    .X(_02971_));
 sg13g2_inv_1 _10938_ (.Y(_02972_),
    .A(_02711_));
 sg13g2_a21oi_1 _10939_ (.A1(_02702_),
    .A2(_02933_),
    .Y(_02973_),
    .B1(_02972_));
 sg13g2_xnor2_1 _10940_ (.Y(_02974_),
    .A(_02691_),
    .B(_02973_));
 sg13g2_xnor2_1 _10941_ (.Y(_02975_),
    .A(_02971_),
    .B(_02974_));
 sg13g2_mux2_1 _10942_ (.A0(_02503_),
    .A1(_02967_),
    .S(_02975_),
    .X(_02976_));
 sg13g2_xor2_1 _10943_ (.B(_02974_),
    .A(_02971_),
    .X(_02977_));
 sg13g2_buf_1 _10944_ (.A(_02977_),
    .X(_02978_));
 sg13g2_mux2_1 _10945_ (.A0(_02541_),
    .A1(_02967_),
    .S(_02978_),
    .X(_02979_));
 sg13g2_xor2_1 _10946_ (.B(_01695_),
    .A(net62),
    .X(_02980_));
 sg13g2_o21ai_1 _10947_ (.B1(_02010_),
    .Y(_02981_),
    .A1(net279),
    .A2(net237));
 sg13g2_a21oi_1 _10948_ (.A1(net148),
    .A2(_02699_),
    .Y(_02982_),
    .B1(_02683_));
 sg13g2_a21oi_1 _10949_ (.A1(_02699_),
    .A2(_02981_),
    .Y(_02983_),
    .B1(_02982_));
 sg13g2_nand2_1 _10950_ (.Y(_02984_),
    .A(_02980_),
    .B(_02983_));
 sg13g2_nand3_1 _10951_ (.B(net237),
    .C(_01992_),
    .A(net287),
    .Y(_02985_));
 sg13g2_xnor2_1 _10952_ (.Y(_02986_),
    .A(net279),
    .B(_02985_));
 sg13g2_and2_1 _10953_ (.A(_02010_),
    .B(_02986_),
    .X(_02987_));
 sg13g2_nand2_1 _10954_ (.Y(_02988_),
    .A(_02450_),
    .B(_02987_));
 sg13g2_nand4_1 _10955_ (.B(_02709_),
    .C(_02984_),
    .A(net39),
    .Y(_02989_),
    .D(_02988_));
 sg13g2_buf_1 _10956_ (.A(_02989_),
    .X(_02990_));
 sg13g2_nand2_1 _10957_ (.Y(_02991_),
    .A(_02980_),
    .B(_02987_));
 sg13g2_o21ai_1 _10958_ (.B1(_02991_),
    .Y(_02992_),
    .A1(_02980_),
    .A2(_02983_));
 sg13g2_o21ai_1 _10959_ (.B1(_02992_),
    .Y(_02993_),
    .A1(_02445_),
    .A2(_01885_));
 sg13g2_buf_1 _10960_ (.A(_02993_),
    .X(_02994_));
 sg13g2_nand2_1 _10961_ (.Y(_02995_),
    .A(_02990_),
    .B(_02994_));
 sg13g2_o21ai_1 _10962_ (.B1(_02539_),
    .Y(_02996_),
    .A1(_02715_),
    .A2(_02716_));
 sg13g2_buf_1 _10963_ (.A(_02996_),
    .X(_02997_));
 sg13g2_nand3b_1 _10964_ (.B(_02426_),
    .C(_02691_),
    .Y(_02998_),
    .A_N(_02715_));
 sg13g2_buf_1 _10965_ (.A(_02998_),
    .X(_02999_));
 sg13g2_nand2_1 _10966_ (.Y(_03000_),
    .A(_02997_),
    .B(_02999_));
 sg13g2_xnor2_1 _10967_ (.Y(_03001_),
    .A(_02995_),
    .B(_03000_));
 sg13g2_xnor2_1 _10968_ (.Y(_03002_),
    .A(_02687_),
    .B(_03001_));
 sg13g2_mux2_1 _10969_ (.A0(_02976_),
    .A1(_02979_),
    .S(_03002_),
    .X(_03003_));
 sg13g2_buf_1 _10970_ (.A(_03003_),
    .X(_03004_));
 sg13g2_xnor2_1 _10971_ (.Y(_03005_),
    .A(_02683_),
    .B(_02717_));
 sg13g2_a21oi_1 _10972_ (.A1(net175),
    .A2(_02968_),
    .Y(_03006_),
    .B1(_02970_));
 sg13g2_nor2_1 _10973_ (.A(_02973_),
    .B(_03005_),
    .Y(_03007_));
 sg13g2_nor2_1 _10974_ (.A(_03006_),
    .B(_03007_),
    .Y(_03008_));
 sg13g2_a21oi_1 _10975_ (.A1(_02973_),
    .A2(_03005_),
    .Y(_03009_),
    .B1(_03008_));
 sg13g2_buf_1 _10976_ (.A(_03009_),
    .X(_03010_));
 sg13g2_nor2_1 _10977_ (.A(_03004_),
    .B(_03010_),
    .Y(_03011_));
 sg13g2_nand2_1 _10978_ (.Y(_03012_),
    .A(_02726_),
    .B(_02728_));
 sg13g2_xnor2_1 _10979_ (.Y(_03013_),
    .A(_02697_),
    .B(_02723_));
 sg13g2_xnor2_1 _10980_ (.Y(_03014_),
    .A(_03012_),
    .B(_03013_));
 sg13g2_buf_2 _10981_ (.A(_03014_),
    .X(_03015_));
 sg13g2_a21oi_1 _10982_ (.A1(_03004_),
    .A2(_03010_),
    .Y(_03016_),
    .B1(_03015_));
 sg13g2_or2_1 _10983_ (.X(_03017_),
    .B(_03016_),
    .A(_03011_));
 sg13g2_buf_1 _10984_ (.A(_02358_),
    .X(_03018_));
 sg13g2_o21ai_1 _10985_ (.B1(_02360_),
    .Y(_03019_),
    .A1(net232),
    .A2(_02377_));
 sg13g2_nor3_1 _10986_ (.A(net246),
    .B(net245),
    .C(net172),
    .Y(_03020_));
 sg13g2_a21oi_1 _10987_ (.A1(net246),
    .A2(_03019_),
    .Y(_03021_),
    .B1(_03020_));
 sg13g2_nor2_1 _10988_ (.A(net172),
    .B(net174),
    .Y(_03022_));
 sg13g2_a21o_1 _10989_ (.A2(_02389_),
    .A1(net245),
    .B1(_03022_),
    .X(_03023_));
 sg13g2_nor2_1 _10990_ (.A(_02360_),
    .B(_02377_),
    .Y(_03024_));
 sg13g2_a22oi_1 _10991_ (.Y(_03025_),
    .B1(_03024_),
    .B2(net169),
    .A2(_03023_),
    .A1(_02377_));
 sg13g2_o21ai_1 _10992_ (.B1(_03025_),
    .Y(_03026_),
    .A1(net169),
    .A2(_03021_));
 sg13g2_buf_1 _10993_ (.A(_03026_),
    .X(_03027_));
 sg13g2_a21oi_1 _10994_ (.A1(_03004_),
    .A2(_03010_),
    .Y(_03028_),
    .B1(_03027_));
 sg13g2_xor2_1 _10995_ (.B(_02754_),
    .A(_02735_),
    .X(_03029_));
 sg13g2_xor2_1 _10996_ (.B(_03029_),
    .A(_02757_),
    .X(_03030_));
 sg13g2_o21ai_1 _10997_ (.B1(_03030_),
    .Y(_03031_),
    .A1(_03017_),
    .A2(_03028_));
 sg13g2_nor2_1 _10998_ (.A(_03015_),
    .B(_03027_),
    .Y(_03032_));
 sg13g2_o21ai_1 _10999_ (.B1(_03032_),
    .Y(_03033_),
    .A1(_03030_),
    .A2(_03011_));
 sg13g2_and2_1 _11000_ (.A(_03031_),
    .B(_03033_),
    .X(_03034_));
 sg13g2_nand2b_1 _11001_ (.Y(_03035_),
    .B(_02765_),
    .A_N(_02764_));
 sg13g2_xnor2_1 _11002_ (.Y(_03036_),
    .A(_02760_),
    .B(_03035_));
 sg13g2_or2_1 _11003_ (.X(_03037_),
    .B(_03036_),
    .A(_03034_));
 sg13g2_buf_1 _11004_ (.A(_03037_),
    .X(_03038_));
 sg13g2_nand4_1 _11005_ (.B(_02940_),
    .C(net36),
    .A(_02938_),
    .Y(_03039_),
    .D(_02953_));
 sg13g2_nand4_1 _11006_ (.B(net38),
    .C(net36),
    .A(net39),
    .Y(_03040_),
    .D(_02942_));
 sg13g2_a22oi_1 _11007_ (.Y(_03041_),
    .B1(_03039_),
    .B2(_03040_),
    .A2(_02433_),
    .A1(_01852_));
 sg13g2_nand4_1 _11008_ (.B(_02431_),
    .C(net38),
    .A(net39),
    .Y(_03042_),
    .D(_02953_));
 sg13g2_nand4_1 _11009_ (.B(_02938_),
    .C(_02940_),
    .A(_02431_),
    .Y(_03043_),
    .D(_02942_));
 sg13g2_a22oi_1 _11010_ (.Y(_03044_),
    .B1(_03042_),
    .B2(_03043_),
    .A2(_02441_),
    .A1(_01806_));
 sg13g2_nor3_1 _11011_ (.A(net51),
    .B(net61),
    .C(_02942_),
    .Y(_03045_));
 sg13g2_nand3_1 _11012_ (.B(net38),
    .C(_03045_),
    .A(_02705_),
    .Y(_03046_));
 sg13g2_nand4_1 _11013_ (.B(_02938_),
    .C(_02940_),
    .A(_01864_),
    .Y(_03047_),
    .D(_02953_));
 sg13g2_nand4_1 _11014_ (.B(_01864_),
    .C(_02948_),
    .A(_02705_),
    .Y(_03048_),
    .D(_02942_));
 sg13g2_o21ai_1 _11015_ (.B1(_02955_),
    .Y(_03049_),
    .A1(_02445_),
    .A2(_02446_));
 sg13g2_nand4_1 _11016_ (.B(_03047_),
    .C(_03048_),
    .A(_03046_),
    .Y(_03050_),
    .D(_03049_));
 sg13g2_nor3_1 _11017_ (.A(_03041_),
    .B(_03044_),
    .C(_03050_),
    .Y(_03051_));
 sg13g2_o21ai_1 _11018_ (.B1(net36),
    .Y(_03052_),
    .A1(_02430_),
    .A2(_01866_));
 sg13g2_nand3_1 _11019_ (.B(_02433_),
    .C(_02448_),
    .A(_01852_),
    .Y(_03053_));
 sg13g2_buf_1 _11020_ (.A(_03053_),
    .X(_03054_));
 sg13g2_and2_1 _11021_ (.A(_03052_),
    .B(_03054_),
    .X(_03055_));
 sg13g2_nand2_1 _11022_ (.Y(_03056_),
    .A(net288),
    .B(_01985_));
 sg13g2_nand2_2 _11023_ (.Y(_03057_),
    .A(net287),
    .B(_01984_));
 sg13g2_xnor2_1 _11024_ (.Y(_03058_),
    .A(_03056_),
    .B(_03057_));
 sg13g2_a21oi_1 _11025_ (.A1(_02002_),
    .A2(net227),
    .Y(_03059_),
    .B1(net173));
 sg13g2_nor2_1 _11026_ (.A(_03058_),
    .B(_03059_),
    .Y(_03060_));
 sg13g2_nand3_1 _11027_ (.B(_01990_),
    .C(net275),
    .A(net279),
    .Y(_03061_));
 sg13g2_inv_1 _11028_ (.Y(_03062_),
    .A(_03061_));
 sg13g2_xor2_1 _11029_ (.B(_03057_),
    .A(_03056_),
    .X(_03063_));
 sg13g2_a22oi_1 _11030_ (.Y(_03064_),
    .B1(_03062_),
    .B2(_03063_),
    .A2(_03060_),
    .A1(_03055_));
 sg13g2_inv_1 _11031_ (.Y(_03065_),
    .A(_03059_));
 sg13g2_a21oi_1 _11032_ (.A1(_03055_),
    .A2(_03065_),
    .Y(_03066_),
    .B1(_03063_));
 sg13g2_a21oi_1 _11033_ (.A1(_03051_),
    .A2(_03064_),
    .Y(_03067_),
    .B1(_03066_));
 sg13g2_nand2_1 _11034_ (.Y(_03068_),
    .A(_03058_),
    .B(_03051_));
 sg13g2_nand2_1 _11035_ (.Y(_03069_),
    .A(net236),
    .B(net227));
 sg13g2_nor2_1 _11036_ (.A(_02448_),
    .B(_03062_),
    .Y(_03070_));
 sg13g2_nor4_1 _11037_ (.A(_02430_),
    .B(_01866_),
    .C(_02506_),
    .D(_03062_),
    .Y(_03071_));
 sg13g2_a221oi_1 _11038_ (.B2(_02504_),
    .C1(_03071_),
    .B1(_03070_),
    .A1(net148),
    .Y(_03072_),
    .A2(_03069_));
 sg13g2_buf_1 _11039_ (.A(_03072_),
    .X(_03073_));
 sg13g2_o21ai_1 _11040_ (.B1(_03073_),
    .Y(_03074_),
    .A1(_03058_),
    .A2(_03051_));
 sg13g2_a21oi_1 _11041_ (.A1(_03068_),
    .A2(_03074_),
    .Y(_03075_),
    .B1(_01729_));
 sg13g2_a21oi_1 _11042_ (.A1(_01729_),
    .A2(_03067_),
    .Y(_03076_),
    .B1(_03075_));
 sg13g2_or4_1 _11043_ (.A(_02946_),
    .B(_02951_),
    .C(_02954_),
    .D(_02961_),
    .X(_03077_));
 sg13g2_buf_1 _11044_ (.A(_03077_),
    .X(_03078_));
 sg13g2_xnor2_1 _11045_ (.Y(_03079_),
    .A(_01823_),
    .B(_02935_));
 sg13g2_nand2_1 _11046_ (.Y(_03080_),
    .A(_02944_),
    .B(_03063_));
 sg13g2_o21ai_1 _11047_ (.B1(_03080_),
    .Y(_03081_),
    .A1(_02000_),
    .A2(_01506_));
 sg13g2_buf_1 _11048_ (.A(_03081_),
    .X(_03082_));
 sg13g2_xnor2_1 _11049_ (.Y(_03083_),
    .A(_02923_),
    .B(_02933_));
 sg13g2_a21o_1 _11050_ (.A2(_03057_),
    .A1(_02953_),
    .B1(_03056_),
    .X(_03084_));
 sg13g2_o21ai_1 _11051_ (.B1(_03084_),
    .Y(_03085_),
    .A1(_02953_),
    .A2(_03057_));
 sg13g2_buf_1 _11052_ (.A(_03085_),
    .X(_03086_));
 sg13g2_xnor2_1 _11053_ (.Y(_03087_),
    .A(_03083_),
    .B(_03086_));
 sg13g2_xnor2_1 _11054_ (.Y(_03088_),
    .A(_03082_),
    .B(_03087_));
 sg13g2_nor2_1 _11055_ (.A(_03079_),
    .B(_03088_),
    .Y(_03089_));
 sg13g2_nand2_1 _11056_ (.Y(_03090_),
    .A(_03078_),
    .B(_03089_));
 sg13g2_nor2_1 _11057_ (.A(_02936_),
    .B(_03088_),
    .Y(_03091_));
 sg13g2_nand2_1 _11058_ (.Y(_03092_),
    .A(_02963_),
    .B(_03091_));
 sg13g2_a21oi_1 _11059_ (.A1(_03090_),
    .A2(_03092_),
    .Y(_03093_),
    .B1(_02931_));
 sg13g2_nand2_1 _11060_ (.Y(_03094_),
    .A(_02963_),
    .B(_03089_));
 sg13g2_nand2_1 _11061_ (.Y(_03095_),
    .A(_03078_),
    .B(_03091_));
 sg13g2_and2_1 _11062_ (.A(_02926_),
    .B(_02930_),
    .X(_03096_));
 sg13g2_a21oi_1 _11063_ (.A1(_03094_),
    .A2(_03095_),
    .Y(_03097_),
    .B1(_03096_));
 sg13g2_xor2_1 _11064_ (.B(_03087_),
    .A(_03082_),
    .X(_03098_));
 sg13g2_nor2_1 _11065_ (.A(_03079_),
    .B(_03098_),
    .Y(_03099_));
 sg13g2_nand2_1 _11066_ (.Y(_03100_),
    .A(_02963_),
    .B(_03099_));
 sg13g2_nor2_1 _11067_ (.A(_02936_),
    .B(_03098_),
    .Y(_03101_));
 sg13g2_nand2_1 _11068_ (.Y(_03102_),
    .A(_03078_),
    .B(_03101_));
 sg13g2_a21oi_1 _11069_ (.A1(_03100_),
    .A2(_03102_),
    .Y(_03103_),
    .B1(_02931_));
 sg13g2_nand2_1 _11070_ (.Y(_03104_),
    .A(_03078_),
    .B(_03099_));
 sg13g2_nand2_1 _11071_ (.Y(_03105_),
    .A(_02963_),
    .B(_03101_));
 sg13g2_a21oi_1 _11072_ (.A1(_03104_),
    .A2(_03105_),
    .Y(_03106_),
    .B1(_03096_));
 sg13g2_or4_1 _11073_ (.A(_03093_),
    .B(_03097_),
    .C(_03103_),
    .D(_03106_),
    .X(_03107_));
 sg13g2_xnor2_1 _11074_ (.Y(_03108_),
    .A(_03076_),
    .B(_03107_));
 sg13g2_buf_2 _11075_ (.A(_03108_),
    .X(_03109_));
 sg13g2_nor2_1 _11076_ (.A(net245),
    .B(net169),
    .Y(_03110_));
 sg13g2_xnor2_1 _11077_ (.Y(_03111_),
    .A(_02942_),
    .B(_03058_));
 sg13g2_nand2_1 _11078_ (.Y(_03112_),
    .A(net287),
    .B(_01986_));
 sg13g2_nand2_1 _11079_ (.Y(_03113_),
    .A(net276),
    .B(net277));
 sg13g2_xnor2_1 _11080_ (.Y(_03114_),
    .A(_03112_),
    .B(_03113_));
 sg13g2_buf_2 _11081_ (.A(_03114_),
    .X(_03115_));
 sg13g2_nor3_1 _11082_ (.A(_01823_),
    .B(net230),
    .C(_03115_),
    .Y(_03116_));
 sg13g2_nand2_1 _11083_ (.Y(_03117_),
    .A(_03111_),
    .B(_03116_));
 sg13g2_o21ai_1 _11084_ (.B1(_03117_),
    .Y(_03118_),
    .A1(net147),
    .A2(_02024_));
 sg13g2_buf_1 _11085_ (.A(_03118_),
    .X(_03119_));
 sg13g2_a221oi_1 _11086_ (.B2(_02504_),
    .C1(_01864_),
    .B1(net36),
    .A1(net39),
    .Y(_03120_),
    .A2(net38));
 sg13g2_or2_1 _11087_ (.X(_03121_),
    .B(_03120_),
    .A(_01885_));
 sg13g2_buf_1 _11088_ (.A(_03121_),
    .X(_03122_));
 sg13g2_xnor2_1 _11089_ (.Y(_03123_),
    .A(_03073_),
    .B(_03111_));
 sg13g2_xnor2_1 _11090_ (.Y(_03124_),
    .A(_03122_),
    .B(_03123_));
 sg13g2_xor2_1 _11091_ (.B(_03113_),
    .A(_03112_),
    .X(_03125_));
 sg13g2_nor2_1 _11092_ (.A(_02430_),
    .B(_01866_),
    .Y(_03126_));
 sg13g2_xnor2_1 _11093_ (.Y(_03127_),
    .A(net148),
    .B(net36));
 sg13g2_xnor2_1 _11094_ (.Y(_03128_),
    .A(_03126_),
    .B(_03127_));
 sg13g2_a21o_1 _11095_ (.A2(_03128_),
    .A1(_03125_),
    .B1(net172),
    .X(_03129_));
 sg13g2_nand4_1 _11096_ (.B(_01852_),
    .C(_02433_),
    .A(net148),
    .Y(_03130_),
    .D(_02448_));
 sg13g2_nand4_1 _11097_ (.B(_01806_),
    .C(_02441_),
    .A(net148),
    .Y(_03131_),
    .D(net36));
 sg13g2_nand3_1 _11098_ (.B(_02448_),
    .C(_03115_),
    .A(_01866_),
    .Y(_03132_));
 sg13g2_nand3_1 _11099_ (.B(_03131_),
    .C(_03132_),
    .A(_03130_),
    .Y(_03133_));
 sg13g2_nor3_1 _11100_ (.A(net175),
    .B(_01866_),
    .C(_03125_),
    .Y(_03134_));
 sg13g2_xnor2_1 _11101_ (.Y(_03135_),
    .A(_01852_),
    .B(net36));
 sg13g2_nand2_1 _11102_ (.Y(_03136_),
    .A(_02448_),
    .B(_03115_));
 sg13g2_nand2_1 _11103_ (.Y(_03137_),
    .A(net173),
    .B(_02507_));
 sg13g2_a22oi_1 _11104_ (.Y(_03138_),
    .B1(_03136_),
    .B2(_03137_),
    .A2(_02441_),
    .A1(_01806_));
 sg13g2_nand2_1 _11105_ (.Y(_03139_),
    .A(_02507_),
    .B(_03115_));
 sg13g2_nand2_1 _11106_ (.Y(_03140_),
    .A(net173),
    .B(_02448_));
 sg13g2_a22oi_1 _11107_ (.Y(_03141_),
    .B1(_03139_),
    .B2(_03140_),
    .A2(_02433_),
    .A1(_01852_));
 sg13g2_nor4_1 _11108_ (.A(_01823_),
    .B(net230),
    .C(_03138_),
    .D(_03141_),
    .Y(_03142_));
 sg13g2_a221oi_1 _11109_ (.B2(_03135_),
    .C1(_03142_),
    .B1(_03134_),
    .A1(net181),
    .Y(_03143_),
    .A2(_03133_));
 sg13g2_xor2_1 _11110_ (.B(_03116_),
    .A(_03111_),
    .X(_03144_));
 sg13g2_a21oi_1 _11111_ (.A1(_03129_),
    .A2(_03143_),
    .Y(_03145_),
    .B1(_03144_));
 sg13g2_nand3_1 _11112_ (.B(_03129_),
    .C(_03143_),
    .A(_03144_),
    .Y(_03146_));
 sg13g2_o21ai_1 _11113_ (.B1(_03146_),
    .Y(_03147_),
    .A1(_03124_),
    .A2(_03145_));
 sg13g2_buf_1 _11114_ (.A(_03147_),
    .X(_03148_));
 sg13g2_nand3_1 _11115_ (.B(_03119_),
    .C(_03148_),
    .A(_03110_),
    .Y(_03149_));
 sg13g2_nand2_1 _11116_ (.Y(_03150_),
    .A(_03119_),
    .B(_03148_));
 sg13g2_nor2_1 _11117_ (.A(_03119_),
    .B(_03148_),
    .Y(_03151_));
 sg13g2_a21oi_1 _11118_ (.A1(_03150_),
    .A2(_03109_),
    .Y(_03152_),
    .B1(_03151_));
 sg13g2_a21oi_1 _11119_ (.A1(_03151_),
    .A2(_03109_),
    .Y(_03153_),
    .B1(_02934_));
 sg13g2_nor2_1 _11120_ (.A(_03093_),
    .B(_03097_),
    .Y(_03154_));
 sg13g2_or2_1 _11121_ (.X(_03155_),
    .B(_03106_),
    .A(_03103_));
 sg13g2_a21oi_1 _11122_ (.A1(_03076_),
    .A2(_03154_),
    .Y(_03156_),
    .B1(_03155_));
 sg13g2_nor2_1 _11123_ (.A(_03082_),
    .B(_03086_),
    .Y(_03157_));
 sg13g2_nor2_1 _11124_ (.A(_03083_),
    .B(_03157_),
    .Y(_03158_));
 sg13g2_a21oi_1 _11125_ (.A1(_03082_),
    .A2(_03086_),
    .Y(_03159_),
    .B1(_03158_));
 sg13g2_and4_1 _11126_ (.A(_02978_),
    .B(_02990_),
    .C(_02994_),
    .D(_03000_),
    .X(_03160_));
 sg13g2_a221oi_1 _11127_ (.B2(_02999_),
    .C1(_02978_),
    .B1(_02997_),
    .A1(_02990_),
    .Y(_03161_),
    .A2(_02994_));
 sg13g2_and2_1 _11128_ (.A(_02997_),
    .B(_02999_),
    .X(_03162_));
 sg13g2_and4_1 _11129_ (.A(_02975_),
    .B(_02990_),
    .C(_02994_),
    .D(_03162_),
    .X(_03163_));
 sg13g2_nand3_1 _11130_ (.B(_02997_),
    .C(_02999_),
    .A(_02978_),
    .Y(_03164_));
 sg13g2_a21oi_1 _11131_ (.A1(_02990_),
    .A2(_02994_),
    .Y(_03165_),
    .B1(_03164_));
 sg13g2_nor4_1 _11132_ (.A(_03160_),
    .B(_03161_),
    .C(_03163_),
    .D(_03165_),
    .Y(_03166_));
 sg13g2_xnor2_1 _11133_ (.Y(_03167_),
    .A(_02967_),
    .B(_03166_));
 sg13g2_xnor2_1 _11134_ (.Y(_03168_),
    .A(_03159_),
    .B(_03167_));
 sg13g2_xnor2_1 _11135_ (.Y(_03169_),
    .A(_03156_),
    .B(_03168_));
 sg13g2_o21ai_1 _11136_ (.B1(_03169_),
    .Y(_03170_),
    .A1(_03152_),
    .A2(_03153_));
 sg13g2_o21ai_1 _11137_ (.B1(_03170_),
    .Y(_03171_),
    .A1(_03109_),
    .A2(_03149_));
 sg13g2_buf_1 _11138_ (.A(_03171_),
    .X(_03172_));
 sg13g2_xnor2_1 _11139_ (.Y(_03173_),
    .A(_03122_),
    .B(_03073_));
 sg13g2_nand2_1 _11140_ (.Y(_03174_),
    .A(net173),
    .B(_03115_));
 sg13g2_nand3_1 _11141_ (.B(_03054_),
    .C(_03174_),
    .A(_03052_),
    .Y(_03175_));
 sg13g2_nand2_1 _11142_ (.Y(_03176_),
    .A(net181),
    .B(_03125_));
 sg13g2_nand3_1 _11143_ (.B(_03054_),
    .C(_03176_),
    .A(_03052_),
    .Y(_03177_));
 sg13g2_a22oi_1 _11144_ (.Y(_03178_),
    .B1(_03177_),
    .B2(net146),
    .A2(_03175_),
    .A1(net175));
 sg13g2_nand2_1 _11145_ (.Y(_03179_),
    .A(_03125_),
    .B(_03128_));
 sg13g2_o21ai_1 _11146_ (.B1(_03179_),
    .Y(_03180_),
    .A1(net230),
    .A2(_03178_));
 sg13g2_xnor2_1 _11147_ (.Y(_03181_),
    .A(_03173_),
    .B(_03180_));
 sg13g2_nand2_1 _11148_ (.Y(_03182_),
    .A(_02303_),
    .B(_02001_));
 sg13g2_nor3_1 _11149_ (.A(net240),
    .B(_01675_),
    .C(_01676_),
    .Y(_03183_));
 sg13g2_o21ai_1 _11150_ (.B1(_03183_),
    .Y(_03184_),
    .A1(_01775_),
    .A2(_01776_));
 sg13g2_or3_1 _11151_ (.A(_01775_),
    .B(_01776_),
    .C(_03183_),
    .X(_03185_));
 sg13g2_and2_1 _11152_ (.A(_01784_),
    .B(_01798_),
    .X(_03186_));
 sg13g2_a21oi_1 _11153_ (.A1(_03184_),
    .A2(_03185_),
    .Y(_03187_),
    .B1(_03186_));
 sg13g2_and3_1 _11154_ (.X(_03188_),
    .A(_03186_),
    .B(_03184_),
    .C(_03185_));
 sg13g2_and4_1 _11155_ (.A(_01819_),
    .B(_01835_),
    .C(_01838_),
    .D(_01840_),
    .X(_03189_));
 sg13g2_a22oi_1 _11156_ (.Y(_03190_),
    .B1(_01838_),
    .B2(_01840_),
    .A2(_01835_),
    .A1(_01819_));
 sg13g2_nor4_2 _11157_ (.A(_03187_),
    .B(_03188_),
    .C(_03189_),
    .Y(_03191_),
    .D(_03190_));
 sg13g2_a22oi_1 _11158_ (.Y(_03192_),
    .B1(_01843_),
    .B2(_01844_),
    .A2(_01835_),
    .A1(_01819_));
 sg13g2_nor4_2 _11159_ (.A(_01845_),
    .B(_01847_),
    .C(_01848_),
    .Y(_03193_),
    .D(_03192_));
 sg13g2_o21ai_1 _11160_ (.B1(net275),
    .Y(_03194_),
    .A1(_03191_),
    .A2(_03193_));
 sg13g2_nor3_1 _11161_ (.A(net275),
    .B(_03191_),
    .C(_03193_),
    .Y(_03195_));
 sg13g2_a21oi_2 _11162_ (.B1(_03195_),
    .Y(_03196_),
    .A2(_03194_),
    .A1(_03182_));
 sg13g2_xor2_1 _11163_ (.B(_01804_),
    .A(_01768_),
    .X(_03197_));
 sg13g2_a21oi_1 _11164_ (.A1(_01842_),
    .A2(_01850_),
    .Y(_03198_),
    .B1(_03197_));
 sg13g2_and3_1 _11165_ (.X(_03199_),
    .A(_01842_),
    .B(_01850_),
    .C(_03197_));
 sg13g2_buf_1 _11166_ (.A(_03199_),
    .X(_03200_));
 sg13g2_nand2_1 _11167_ (.Y(_03201_),
    .A(net276),
    .B(net228));
 sg13g2_o21ai_1 _11168_ (.B1(_03201_),
    .Y(_03202_),
    .A1(_03198_),
    .A2(_03200_));
 sg13g2_nor3_1 _11169_ (.A(_03201_),
    .B(_03198_),
    .C(_03200_),
    .Y(_03203_));
 sg13g2_a21oi_2 _11170_ (.B1(_03203_),
    .Y(_03204_),
    .A2(_03202_),
    .A1(_03196_));
 sg13g2_nor2_1 _11171_ (.A(net181),
    .B(_02742_),
    .Y(_03205_));
 sg13g2_nand2b_1 _11172_ (.Y(_03206_),
    .B(_03205_),
    .A_N(_03204_));
 sg13g2_nor2_2 _11173_ (.A(net148),
    .B(net275),
    .Y(_03207_));
 sg13g2_xnor2_1 _11174_ (.Y(_03208_),
    .A(_02506_),
    .B(_03207_));
 sg13g2_xnor2_1 _11175_ (.Y(_03209_),
    .A(_03126_),
    .B(_03208_));
 sg13g2_buf_2 _11176_ (.A(_03209_),
    .X(_03210_));
 sg13g2_nand2_1 _11177_ (.Y(_03211_),
    .A(_03125_),
    .B(_03210_));
 sg13g2_a21oi_1 _11178_ (.A1(_03181_),
    .A2(_03206_),
    .Y(_03212_),
    .B1(_03211_));
 sg13g2_buf_1 _11179_ (.A(net175),
    .X(_03213_));
 sg13g2_nand2_1 _11180_ (.Y(_03214_),
    .A(net144),
    .B(net170));
 sg13g2_a21oi_1 _11181_ (.A1(_03204_),
    .A2(_03210_),
    .Y(_03215_),
    .B1(_03214_));
 sg13g2_nor2_1 _11182_ (.A(_03204_),
    .B(_03210_),
    .Y(_03216_));
 sg13g2_nor2_1 _11183_ (.A(_03215_),
    .B(_03216_),
    .Y(_03217_));
 sg13g2_nor2_1 _11184_ (.A(_03181_),
    .B(_03217_),
    .Y(_03218_));
 sg13g2_or2_1 _11185_ (.X(_03219_),
    .B(_03218_),
    .A(_03212_));
 sg13g2_buf_1 _11186_ (.A(_03219_),
    .X(_03220_));
 sg13g2_xnor2_1 _11187_ (.Y(_03221_),
    .A(_03110_),
    .B(_03119_));
 sg13g2_xnor2_1 _11188_ (.Y(_03222_),
    .A(_03148_),
    .B(_03221_));
 sg13g2_xnor2_1 _11189_ (.Y(_03223_),
    .A(_03109_),
    .B(_03222_));
 sg13g2_nor2_1 _11190_ (.A(_03220_),
    .B(_03223_),
    .Y(_03224_));
 sg13g2_and2_1 _11191_ (.A(_03196_),
    .B(_03202_),
    .X(_03225_));
 sg13g2_nor3_1 _11192_ (.A(_03225_),
    .B(_03203_),
    .C(_03210_),
    .Y(_03226_));
 sg13g2_xnor2_1 _11193_ (.Y(_03227_),
    .A(_03115_),
    .B(_03206_));
 sg13g2_a22oi_1 _11194_ (.Y(_03228_),
    .B1(_03227_),
    .B2(_03210_),
    .A2(_03226_),
    .A1(_03214_));
 sg13g2_xor2_1 _11195_ (.B(_03228_),
    .A(_03181_),
    .X(_03229_));
 sg13g2_or2_1 _11196_ (.X(_03230_),
    .B(_03193_),
    .A(_03191_));
 sg13g2_buf_2 _11197_ (.A(_03230_),
    .X(_03231_));
 sg13g2_nor2_1 _11198_ (.A(_02742_),
    .B(_02314_),
    .Y(_03232_));
 sg13g2_o21ai_1 _11199_ (.B1(_03232_),
    .Y(_03233_),
    .A1(net228),
    .A2(_03231_));
 sg13g2_xnor2_1 _11200_ (.Y(_03234_),
    .A(_01819_),
    .B(_01835_));
 sg13g2_inv_1 _11201_ (.Y(_03235_),
    .A(_03234_));
 sg13g2_nand3_1 _11202_ (.B(_01994_),
    .C(_03235_),
    .A(net228),
    .Y(_03236_));
 sg13g2_nand3_1 _11203_ (.B(_03207_),
    .C(_03235_),
    .A(net228),
    .Y(_03237_));
 sg13g2_mux2_1 _11204_ (.A0(_03236_),
    .A1(_03237_),
    .S(_03231_),
    .X(_03238_));
 sg13g2_nand3b_1 _11205_ (.B(_03207_),
    .C(net277),
    .Y(_03239_),
    .A_N(_03231_));
 sg13g2_buf_1 _11206_ (.A(_03234_),
    .X(_03240_));
 sg13g2_nand2_2 _11207_ (.Y(_03241_),
    .A(_02313_),
    .B(_02001_));
 sg13g2_or3_1 _11208_ (.A(_03231_),
    .B(net50),
    .C(_03241_),
    .X(_03242_));
 sg13g2_nand4_1 _11209_ (.B(_03238_),
    .C(_03239_),
    .A(_03233_),
    .Y(_03243_),
    .D(_03242_));
 sg13g2_buf_1 _11210_ (.A(_03243_),
    .X(_03244_));
 sg13g2_nor3_1 _11211_ (.A(net169),
    .B(_02683_),
    .C(_03244_),
    .Y(_03245_));
 sg13g2_and4_1 _11212_ (.A(_03233_),
    .B(_03238_),
    .C(_03239_),
    .D(_03242_),
    .X(_03246_));
 sg13g2_buf_1 _11213_ (.A(_03246_),
    .X(_03247_));
 sg13g2_nor4_1 _11214_ (.A(net178),
    .B(net181),
    .C(net169),
    .D(_03247_),
    .Y(_03248_));
 sg13g2_nor2_1 _11215_ (.A(_03198_),
    .B(_03200_),
    .Y(_03249_));
 sg13g2_xnor2_1 _11216_ (.Y(_03250_),
    .A(_03196_),
    .B(_03249_));
 sg13g2_buf_1 _11217_ (.A(_03250_),
    .X(_03251_));
 sg13g2_nor2_1 _11218_ (.A(_03247_),
    .B(_03251_),
    .Y(_03252_));
 sg13g2_nor2_1 _11219_ (.A(net181),
    .B(_02358_),
    .Y(_03253_));
 sg13g2_nor2b_1 _11220_ (.A(net175),
    .B_N(net233),
    .Y(_03254_));
 sg13g2_and2_1 _11221_ (.A(net174),
    .B(_03254_),
    .X(_03255_));
 sg13g2_mux2_1 _11222_ (.A0(_03253_),
    .A1(_03255_),
    .S(_03251_),
    .X(_03256_));
 sg13g2_nor4_1 _11223_ (.A(_03245_),
    .B(_03248_),
    .C(_03252_),
    .D(_03256_),
    .Y(_03257_));
 sg13g2_xnor2_1 _11224_ (.Y(_03258_),
    .A(_03204_),
    .B(_03210_));
 sg13g2_xnor2_1 _11225_ (.Y(_03259_),
    .A(_03205_),
    .B(_03258_));
 sg13g2_xnor2_1 _11226_ (.Y(_03260_),
    .A(_03257_),
    .B(_03259_));
 sg13g2_xnor2_1 _11227_ (.Y(_03261_),
    .A(_03251_),
    .B(_03253_));
 sg13g2_xnor2_1 _11228_ (.Y(_03262_),
    .A(_03244_),
    .B(_03261_));
 sg13g2_nand2_1 _11229_ (.Y(_03263_),
    .A(_01990_),
    .B(net228));
 sg13g2_nor2_1 _11230_ (.A(_01993_),
    .B(net277),
    .Y(_03264_));
 sg13g2_xor2_1 _11231_ (.B(_03264_),
    .A(_03263_),
    .X(_03265_));
 sg13g2_xnor2_1 _11232_ (.Y(_03266_),
    .A(_03231_),
    .B(_03265_));
 sg13g2_buf_1 _11233_ (.A(_00013_),
    .X(_03267_));
 sg13g2_and2_1 _11234_ (.A(_03267_),
    .B(_02743_),
    .X(_03268_));
 sg13g2_nor2_1 _11235_ (.A(_03267_),
    .B(_02000_),
    .Y(_03269_));
 sg13g2_buf_1 _11236_ (.A(net125),
    .X(_03270_));
 sg13g2_inv_1 _11237_ (.Y(_03271_),
    .A(net105));
 sg13g2_xnor2_1 _11238_ (.Y(_03272_),
    .A(_03271_),
    .B(_01830_));
 sg13g2_nand2_1 _11239_ (.Y(_03273_),
    .A(net183),
    .B(_03272_));
 sg13g2_xor2_1 _11240_ (.B(_03273_),
    .A(_01829_),
    .X(_03274_));
 sg13g2_buf_1 _11241_ (.A(_03274_),
    .X(_03275_));
 sg13g2_mux2_1 _11242_ (.A0(_03268_),
    .A1(_03269_),
    .S(net60),
    .X(_03276_));
 sg13g2_nand2_1 _11243_ (.Y(_03277_),
    .A(_02313_),
    .B(net228));
 sg13g2_buf_1 _11244_ (.A(_03277_),
    .X(_03278_));
 sg13g2_xor2_1 _11245_ (.B(net143),
    .A(net50),
    .X(_03279_));
 sg13g2_and2_1 _11246_ (.A(_03276_),
    .B(_03279_),
    .X(_03280_));
 sg13g2_nand2_1 _11247_ (.Y(_03281_),
    .A(_02335_),
    .B(_01780_));
 sg13g2_buf_2 _11248_ (.A(_03281_),
    .X(_03282_));
 sg13g2_xnor2_1 _11249_ (.Y(_03283_),
    .A(net188),
    .B(net185));
 sg13g2_nand4_1 _11250_ (.B(_02289_),
    .C(_03282_),
    .A(net183),
    .Y(_03284_),
    .D(_03283_));
 sg13g2_buf_1 _11251_ (.A(_03284_),
    .X(_03285_));
 sg13g2_nor4_1 _11252_ (.A(_02743_),
    .B(net50),
    .C(net143),
    .D(_03275_),
    .Y(_03286_));
 sg13g2_and3_1 _11253_ (.X(_03287_),
    .A(net50),
    .B(net143),
    .C(_03275_));
 sg13g2_nand3_1 _11254_ (.B(net50),
    .C(net143),
    .A(net147),
    .Y(_03288_));
 sg13g2_nand3_1 _11255_ (.B(net147),
    .C(net60),
    .A(_03267_),
    .Y(_03289_));
 sg13g2_nand3b_1 _11256_ (.B(_03288_),
    .C(_03289_),
    .Y(_03290_),
    .A_N(_03276_));
 sg13g2_or4_1 _11257_ (.A(_03285_),
    .B(_03286_),
    .C(_03287_),
    .D(_03290_),
    .X(_03291_));
 sg13g2_nor2_1 _11258_ (.A(net50),
    .B(net143),
    .Y(_03292_));
 sg13g2_nor2_1 _11259_ (.A(_03267_),
    .B(net60),
    .Y(_03293_));
 sg13g2_a22oi_1 _11260_ (.Y(_03294_),
    .B1(_03293_),
    .B2(_03279_),
    .A2(_03292_),
    .A1(net60));
 sg13g2_nand2_1 _11261_ (.Y(_03295_),
    .A(_03291_),
    .B(_03294_));
 sg13g2_nor3_2 _11262_ (.A(_03240_),
    .B(net143),
    .C(net60),
    .Y(_03296_));
 sg13g2_xor2_1 _11263_ (.B(_03296_),
    .A(_03266_),
    .X(_03297_));
 sg13g2_a22oi_1 _11264_ (.Y(_03298_),
    .B1(_03295_),
    .B2(_03297_),
    .A2(_03280_),
    .A1(_03266_));
 sg13g2_nand2_1 _11265_ (.Y(_03299_),
    .A(_02304_),
    .B(_02743_));
 sg13g2_nand2_1 _11266_ (.Y(_03300_),
    .A(net50),
    .B(_03241_));
 sg13g2_o21ai_1 _11267_ (.B1(_03263_),
    .Y(_03301_),
    .A1(_03234_),
    .A2(_03241_));
 sg13g2_nand2_1 _11268_ (.Y(_03302_),
    .A(_03300_),
    .B(_03301_));
 sg13g2_xnor2_1 _11269_ (.Y(_03303_),
    .A(_03231_),
    .B(_03302_));
 sg13g2_xor2_1 _11270_ (.B(_03263_),
    .A(_03241_),
    .X(_03304_));
 sg13g2_a21oi_1 _11271_ (.A1(net50),
    .A2(_03304_),
    .Y(_03305_),
    .B1(_03296_));
 sg13g2_a21o_1 _11272_ (.A2(_03303_),
    .A1(net172),
    .B1(_03305_),
    .X(_03306_));
 sg13g2_mux2_1 _11273_ (.A0(net230),
    .A1(_03305_),
    .S(_03303_),
    .X(_03307_));
 sg13g2_a21o_1 _11274_ (.A2(_03306_),
    .A1(_03299_),
    .B1(_03307_),
    .X(_03308_));
 sg13g2_and2_1 _11275_ (.A(_03298_),
    .B(_03308_),
    .X(_03309_));
 sg13g2_or2_1 _11276_ (.X(_03310_),
    .B(_03308_),
    .A(_03298_));
 sg13g2_o21ai_1 _11277_ (.B1(_03310_),
    .Y(_03311_),
    .A1(_03262_),
    .A2(_03309_));
 sg13g2_buf_1 _11278_ (.A(_03311_),
    .X(_03312_));
 sg13g2_nand2b_1 _11279_ (.Y(_03313_),
    .B(_03251_),
    .A_N(_03201_));
 sg13g2_nand2_1 _11280_ (.Y(_03314_),
    .A(_03247_),
    .B(_03251_));
 sg13g2_a21oi_1 _11281_ (.A1(_03253_),
    .A2(_03314_),
    .Y(_03315_),
    .B1(_03252_));
 sg13g2_nand2b_1 _11282_ (.Y(_03316_),
    .B(_03244_),
    .A_N(_03313_));
 sg13g2_mux2_1 _11283_ (.A0(_03205_),
    .A1(_02742_),
    .S(_03258_),
    .X(_03317_));
 sg13g2_and2_1 _11284_ (.A(net181),
    .B(_03258_),
    .X(_03318_));
 sg13g2_a221oi_1 _11285_ (.B2(_03317_),
    .C1(_03318_),
    .B1(_03316_),
    .A1(_03313_),
    .Y(_03319_),
    .A2(_03315_));
 sg13g2_buf_1 _11286_ (.A(_03319_),
    .X(_03320_));
 sg13g2_a21oi_1 _11287_ (.A1(_03260_),
    .A2(_03312_),
    .Y(_03321_),
    .B1(_03320_));
 sg13g2_nand3_1 _11288_ (.B(_03312_),
    .C(_03320_),
    .A(_03260_),
    .Y(_03322_));
 sg13g2_o21ai_1 _11289_ (.B1(_03322_),
    .Y(_03323_),
    .A1(_03229_),
    .A2(_03321_));
 sg13g2_a21oi_1 _11290_ (.A1(_03220_),
    .A2(_03223_),
    .Y(_03324_),
    .B1(_03323_));
 sg13g2_o21ai_1 _11291_ (.B1(_03151_),
    .Y(_03325_),
    .A1(_02934_),
    .A2(_03109_));
 sg13g2_a21o_1 _11292_ (.A2(_03148_),
    .A1(_03119_),
    .B1(_03110_),
    .X(_03326_));
 sg13g2_mux2_1 _11293_ (.A0(_03149_),
    .A1(_03326_),
    .S(_03109_),
    .X(_03327_));
 sg13g2_a21oi_1 _11294_ (.A1(_03325_),
    .A2(_03327_),
    .Y(_03328_),
    .B1(_03169_));
 sg13g2_and3_1 _11295_ (.X(_03329_),
    .A(_03169_),
    .B(_03325_),
    .C(_03327_));
 sg13g2_nor4_2 _11296_ (.A(_03224_),
    .B(_03324_),
    .C(_03328_),
    .Y(_03330_),
    .D(_03329_));
 sg13g2_inv_1 _11297_ (.Y(_03331_),
    .A(_03027_));
 sg13g2_xnor2_1 _11298_ (.Y(_03332_),
    .A(_03331_),
    .B(_03010_));
 sg13g2_xnor2_1 _11299_ (.Y(_03333_),
    .A(_03015_),
    .B(_03332_));
 sg13g2_xnor2_1 _11300_ (.Y(_03334_),
    .A(_03004_),
    .B(_03333_));
 sg13g2_a21o_1 _11301_ (.A2(_03086_),
    .A1(_03082_),
    .B1(_03158_),
    .X(_03335_));
 sg13g2_and4_1 _11302_ (.A(_02687_),
    .B(_03156_),
    .C(_03335_),
    .D(_03167_),
    .X(_03336_));
 sg13g2_nand2_1 _11303_ (.Y(_03337_),
    .A(_03159_),
    .B(_03167_));
 sg13g2_mux2_1 _11304_ (.A0(_03335_),
    .A1(_02687_),
    .S(_03167_),
    .X(_03338_));
 sg13g2_a21o_1 _11305_ (.A2(_03337_),
    .A1(_03156_),
    .B1(_03338_),
    .X(_03339_));
 sg13g2_nand2b_1 _11306_ (.Y(_03340_),
    .B(_03339_),
    .A_N(_03336_));
 sg13g2_xnor2_1 _11307_ (.Y(_03341_),
    .A(_03334_),
    .B(_03340_));
 sg13g2_a21oi_1 _11308_ (.A1(_03172_),
    .A2(_03330_),
    .Y(_03342_),
    .B1(_03341_));
 sg13g2_nor2_1 _11309_ (.A(_03172_),
    .B(_03330_),
    .Y(_03343_));
 sg13g2_nor2_1 _11310_ (.A(_03342_),
    .B(_03343_),
    .Y(_03344_));
 sg13g2_a21oi_2 _11311_ (.B1(_03336_),
    .Y(_03345_),
    .A2(_03339_),
    .A1(_03334_));
 sg13g2_and3_1 _11312_ (.X(_03346_),
    .A(_03015_),
    .B(_03027_),
    .C(_03004_));
 sg13g2_nand2_1 _11313_ (.Y(_03347_),
    .A(_02541_),
    .B(_02978_));
 sg13g2_o21ai_1 _11314_ (.B1(_03347_),
    .Y(_03348_),
    .A1(_02967_),
    .A2(_02978_));
 sg13g2_nand2_1 _11315_ (.Y(_03349_),
    .A(_02503_),
    .B(_02975_));
 sg13g2_o21ai_1 _11316_ (.B1(_03349_),
    .Y(_03350_),
    .A1(_02967_),
    .A2(_02975_));
 sg13g2_mux2_1 _11317_ (.A0(_03348_),
    .A1(_03350_),
    .S(_03002_),
    .X(_03351_));
 sg13g2_inv_1 _11318_ (.Y(_03352_),
    .A(_03010_));
 sg13g2_nor3_1 _11319_ (.A(_03331_),
    .B(_03351_),
    .C(_03352_),
    .Y(_03353_));
 sg13g2_nor4_1 _11320_ (.A(_03015_),
    .B(_03027_),
    .C(_03004_),
    .D(_03010_),
    .Y(_03354_));
 sg13g2_nand2_1 _11321_ (.Y(_03355_),
    .A(_03012_),
    .B(_03013_));
 sg13g2_or2_1 _11322_ (.X(_03356_),
    .B(_03013_),
    .A(_03012_));
 sg13g2_a221oi_1 _11323_ (.B2(_03351_),
    .C1(_03352_),
    .B1(_03331_),
    .A1(_03355_),
    .Y(_03357_),
    .A2(_03356_));
 sg13g2_nor4_1 _11324_ (.A(_03346_),
    .B(_03353_),
    .C(_03354_),
    .D(_03357_),
    .Y(_03358_));
 sg13g2_xnor2_1 _11325_ (.Y(_03359_),
    .A(_03030_),
    .B(_03358_));
 sg13g2_nand2_1 _11326_ (.Y(_03360_),
    .A(net150),
    .B(net169));
 sg13g2_o21ai_1 _11327_ (.B1(_03360_),
    .Y(_03361_),
    .A1(_03345_),
    .A2(_03359_));
 sg13g2_nand2_1 _11328_ (.Y(_03362_),
    .A(_03345_),
    .B(_03359_));
 sg13g2_and2_1 _11329_ (.A(_03361_),
    .B(_03362_),
    .X(_03363_));
 sg13g2_nand3_1 _11330_ (.B(_03345_),
    .C(_03359_),
    .A(_03360_),
    .Y(_03364_));
 sg13g2_o21ai_1 _11331_ (.B1(_03364_),
    .Y(_03365_),
    .A1(_03344_),
    .A2(_03363_));
 sg13g2_buf_1 _11332_ (.A(_03365_),
    .X(_03366_));
 sg13g2_and2_1 _11333_ (.A(_03038_),
    .B(_03366_),
    .X(_03367_));
 sg13g2_xnor2_1 _11334_ (.Y(_03368_),
    .A(_02893_),
    .B(_02672_));
 sg13g2_nand2b_1 _11335_ (.Y(_03369_),
    .B(_02768_),
    .A_N(_03368_));
 sg13g2_and2_1 _11336_ (.A(_02840_),
    .B(_02847_),
    .X(_03370_));
 sg13g2_inv_1 _11337_ (.Y(_03371_),
    .A(_02849_));
 sg13g2_mux2_1 _11338_ (.A0(_03370_),
    .A1(_03371_),
    .S(_02890_),
    .X(_03372_));
 sg13g2_inv_1 _11339_ (.Y(_03373_),
    .A(_02894_));
 sg13g2_nor3_1 _11340_ (.A(net26),
    .B(_02672_),
    .C(_03373_),
    .Y(_03374_));
 sg13g2_nand3_1 _11341_ (.B(_02672_),
    .C(_02894_),
    .A(net26),
    .Y(_03375_));
 sg13g2_nor2_1 _11342_ (.A(net24),
    .B(_03375_),
    .Y(_03376_));
 sg13g2_a221oi_1 _11343_ (.B2(net24),
    .C1(_03376_),
    .B1(_03374_),
    .A1(_03369_),
    .Y(_03377_),
    .A2(_03372_));
 sg13g2_nand2_1 _11344_ (.Y(_03378_),
    .A(_03034_),
    .B(_03036_));
 sg13g2_or2_1 _11345_ (.X(_03379_),
    .B(_02766_),
    .A(_02674_));
 sg13g2_buf_1 _11346_ (.A(_03379_),
    .X(_03380_));
 sg13g2_nand3_1 _11347_ (.B(_03378_),
    .C(_03380_),
    .A(_02768_),
    .Y(_03381_));
 sg13g2_or3_1 _11348_ (.A(_03367_),
    .B(_03377_),
    .C(_03381_),
    .X(_03382_));
 sg13g2_buf_1 _11349_ (.A(_03382_),
    .X(_03383_));
 sg13g2_nand3b_1 _11350_ (.B(_02922_),
    .C(_03383_),
    .Y(_03384_),
    .A_N(_02908_));
 sg13g2_nand2_1 _11351_ (.Y(_03385_),
    .A(_02855_),
    .B(_02881_));
 sg13g2_nor2_1 _11352_ (.A(_02855_),
    .B(_02881_),
    .Y(_03386_));
 sg13g2_a21oi_1 _11353_ (.A1(_03385_),
    .A2(_02889_),
    .Y(_03387_),
    .B1(_03386_));
 sg13g2_buf_2 _11354_ (.A(_03387_),
    .X(_03388_));
 sg13g2_nand2_1 _11355_ (.Y(_03389_),
    .A(_02922_),
    .B(_03388_));
 sg13g2_nand3b_1 _11356_ (.B(_03388_),
    .C(_03383_),
    .Y(_03390_),
    .A_N(_02908_));
 sg13g2_and3_1 _11357_ (.X(_03391_),
    .A(_03384_),
    .B(_03389_),
    .C(_03390_));
 sg13g2_inv_1 _11358_ (.Y(_03392_),
    .A(_02915_));
 sg13g2_nor2_1 _11359_ (.A(_03392_),
    .B(_02919_),
    .Y(_03393_));
 sg13g2_nand2_1 _11360_ (.Y(_03394_),
    .A(_03392_),
    .B(_02919_));
 sg13g2_o21ai_1 _11361_ (.B1(_03394_),
    .Y(_03395_),
    .A1(_02913_),
    .A2(_03393_));
 sg13g2_buf_2 _11362_ (.A(_03395_),
    .X(_03396_));
 sg13g2_o21ai_1 _11363_ (.B1(_03396_),
    .Y(_03397_),
    .A1(_02357_),
    .A2(_03391_));
 sg13g2_nand2_1 _11364_ (.Y(_03398_),
    .A(_02357_),
    .B(_03391_));
 sg13g2_nand2_1 _11365_ (.Y(_03399_),
    .A(_03397_),
    .B(_03398_));
 sg13g2_nor2_2 _11366_ (.A(_02262_),
    .B(_02353_),
    .Y(_03400_));
 sg13g2_a21oi_1 _11367_ (.A1(_02354_),
    .A2(_03399_),
    .Y(_03401_),
    .B1(_03400_));
 sg13g2_xnor2_1 _11368_ (.Y(_03402_),
    .A(_02237_),
    .B(_02250_));
 sg13g2_nor2b_1 _11369_ (.A(_03401_),
    .B_N(_03402_),
    .Y(_03403_));
 sg13g2_a21oi_1 _11370_ (.A1(_02255_),
    .A2(_02260_),
    .Y(_03404_),
    .B1(_03403_));
 sg13g2_nand2b_1 _11371_ (.Y(_03405_),
    .B(_02259_),
    .A_N(_02251_));
 sg13g2_a21oi_1 _11372_ (.A1(_03403_),
    .A2(_02253_),
    .Y(_03406_),
    .B1(_03405_));
 sg13g2_nor3_1 _11373_ (.A(_02163_),
    .B(_03404_),
    .C(_03406_),
    .Y(_03407_));
 sg13g2_xnor2_1 _11374_ (.Y(_03408_),
    .A(_02161_),
    .B(_03407_));
 sg13g2_nor2b_1 _11375_ (.A(_01439_),
    .B_N(_00390_),
    .Y(_03409_));
 sg13g2_xor2_1 _11376_ (.B(_01441_),
    .A(_01457_),
    .X(_03410_));
 sg13g2_or2_1 _11377_ (.X(_03411_),
    .B(_00890_),
    .A(_00893_));
 sg13g2_buf_1 _11378_ (.A(_03411_),
    .X(_03412_));
 sg13g2_o21ai_1 _11379_ (.B1(_03412_),
    .Y(_03413_),
    .A1(_00802_),
    .A2(_00808_));
 sg13g2_or3_1 _11380_ (.A(_00802_),
    .B(_00808_),
    .C(_03412_),
    .X(_03414_));
 sg13g2_a21oi_1 _11381_ (.A1(_03413_),
    .A2(_03414_),
    .Y(_03415_),
    .B1(_00921_));
 sg13g2_nor2_1 _11382_ (.A(_00895_),
    .B(_00916_),
    .Y(_03416_));
 sg13g2_mux2_1 _11383_ (.A0(_03415_),
    .A1(_03416_),
    .S(_00717_),
    .X(_03417_));
 sg13g2_nand3_1 _11384_ (.B(_01416_),
    .C(_03417_),
    .A(_01421_),
    .Y(_03418_));
 sg13g2_nor3_1 _11385_ (.A(_00931_),
    .B(_00941_),
    .C(_01013_),
    .Y(_03419_));
 sg13g2_a21oi_1 _11386_ (.A1(_01017_),
    .A2(_01019_),
    .Y(_03420_),
    .B1(_01020_));
 sg13g2_o21ai_1 _11387_ (.B1(_01104_),
    .Y(_03421_),
    .A1(_03419_),
    .A2(_03420_));
 sg13g2_buf_1 _11388_ (.A(_03421_),
    .X(_03422_));
 sg13g2_nand3_1 _11389_ (.B(_03422_),
    .C(_03417_),
    .A(_00883_),
    .Y(_03423_));
 sg13g2_nand3_1 _11390_ (.B(_00810_),
    .C(_03412_),
    .A(_00895_),
    .Y(_03424_));
 sg13g2_or4_1 _11391_ (.A(net23),
    .B(_01421_),
    .C(_03422_),
    .D(_03424_),
    .X(_03425_));
 sg13g2_or4_1 _11392_ (.A(_01426_),
    .B(_00883_),
    .C(_01416_),
    .D(_03424_),
    .X(_03426_));
 sg13g2_nand4_1 _11393_ (.B(_03423_),
    .C(_03425_),
    .A(_03418_),
    .Y(_03427_),
    .D(_03426_));
 sg13g2_nor2_1 _11394_ (.A(_00883_),
    .B(_03412_),
    .Y(_03428_));
 sg13g2_nor4_1 _11395_ (.A(_01421_),
    .B(_00895_),
    .C(_00892_),
    .D(_01414_),
    .Y(_03429_));
 sg13g2_a221oi_1 _11396_ (.B2(_01023_),
    .C1(net23),
    .B1(_03429_),
    .A1(_03422_),
    .Y(_03430_),
    .A2(_03428_));
 sg13g2_nor3_1 _11397_ (.A(_01421_),
    .B(_03412_),
    .C(_01414_),
    .Y(_03431_));
 sg13g2_a221oi_1 _11398_ (.B2(_01023_),
    .C1(_01426_),
    .B1(_03431_),
    .A1(_00897_),
    .Y(_03432_),
    .A2(_03422_));
 sg13g2_nor3_1 _11399_ (.A(net22),
    .B(_03430_),
    .C(_03432_),
    .Y(_03433_));
 sg13g2_nor2b_1 _11400_ (.A(_01127_),
    .B_N(_01412_),
    .Y(_03434_));
 sg13g2_a21oi_1 _11401_ (.A1(_01015_),
    .A2(_01022_),
    .Y(_03435_),
    .B1(_01104_));
 sg13g2_nor3_1 _11402_ (.A(_01414_),
    .B(_03419_),
    .C(_03420_),
    .Y(_03436_));
 sg13g2_nor3_1 _11403_ (.A(_03434_),
    .B(_03435_),
    .C(_03436_),
    .Y(_03437_));
 sg13g2_o21ai_1 _11404_ (.B1(_03434_),
    .Y(_03438_),
    .A1(_03435_),
    .A2(_03436_));
 sg13g2_o21ai_1 _11405_ (.B1(_03438_),
    .Y(_03439_),
    .A1(_01098_),
    .A2(_03437_));
 sg13g2_o21ai_1 _11406_ (.B1(_03439_),
    .Y(_03440_),
    .A1(_03427_),
    .A2(_03433_));
 sg13g2_o21ai_1 _11407_ (.B1(_00895_),
    .Y(_03441_),
    .A1(_00916_),
    .A2(_00892_));
 sg13g2_buf_1 _11408_ (.A(_03441_),
    .X(_03442_));
 sg13g2_nand2_1 _11409_ (.Y(_03443_),
    .A(_00690_),
    .B(_03442_));
 sg13g2_o21ai_1 _11410_ (.B1(_00636_),
    .Y(_03444_),
    .A1(_00690_),
    .A2(_03442_));
 sg13g2_nand2_1 _11411_ (.Y(_03445_),
    .A(_03443_),
    .B(_03444_));
 sg13g2_nand2_1 _11412_ (.Y(_03446_),
    .A(_00636_),
    .B(_03443_));
 sg13g2_nor3_1 _11413_ (.A(_00690_),
    .B(_00575_),
    .C(_03442_),
    .Y(_03447_));
 sg13g2_or2_1 _11414_ (.X(_03448_),
    .B(_03447_),
    .A(_00636_));
 sg13g2_a22oi_1 _11415_ (.Y(_03449_),
    .B1(_03446_),
    .B2(_03448_),
    .A2(_03445_),
    .A1(_00575_));
 sg13g2_xnor2_1 _11416_ (.Y(_03450_),
    .A(_00706_),
    .B(_03449_));
 sg13g2_or2_1 _11417_ (.X(_03451_),
    .B(_03450_),
    .A(_03440_));
 sg13g2_buf_1 _11418_ (.A(_03451_),
    .X(_03452_));
 sg13g2_nor2b_1 _11419_ (.A(_01464_),
    .B_N(_01461_),
    .Y(_03453_));
 sg13g2_o21ai_1 _11420_ (.B1(_03453_),
    .Y(_03454_),
    .A1(_01472_),
    .A2(_03452_));
 sg13g2_nor2_1 _11421_ (.A(_00883_),
    .B(_01416_),
    .Y(_03455_));
 sg13g2_a21oi_1 _11422_ (.A1(net52),
    .A2(net22),
    .Y(_03456_),
    .B1(_00890_));
 sg13g2_nor2_1 _11423_ (.A(net52),
    .B(net22),
    .Y(_03457_));
 sg13g2_o21ai_1 _11424_ (.B1(net23),
    .Y(_03458_),
    .A1(_03456_),
    .A2(_03457_));
 sg13g2_inv_1 _11425_ (.Y(_03459_),
    .A(_03416_));
 sg13g2_o21ai_1 _11426_ (.B1(_03459_),
    .Y(_03460_),
    .A1(net23),
    .A2(_03457_));
 sg13g2_nand2_1 _11427_ (.Y(_03461_),
    .A(_00883_),
    .B(_01416_));
 sg13g2_nor2_1 _11428_ (.A(net23),
    .B(_03456_),
    .Y(_03462_));
 sg13g2_a221oi_1 _11429_ (.B2(_03461_),
    .C1(_03462_),
    .B1(_03460_),
    .A1(_03455_),
    .Y(_03463_),
    .A2(_03458_));
 sg13g2_o21ai_1 _11430_ (.B1(_00693_),
    .Y(_03464_),
    .A1(_00706_),
    .A2(_03463_));
 sg13g2_nand2_1 _11431_ (.Y(_03465_),
    .A(_00706_),
    .B(_03463_));
 sg13g2_a21o_1 _11432_ (.A2(_03465_),
    .A1(_03464_),
    .B1(_00714_),
    .X(_03466_));
 sg13g2_buf_1 _11433_ (.A(_03466_),
    .X(_03467_));
 sg13g2_nor2b_1 _11434_ (.A(_00708_),
    .B_N(_00714_),
    .Y(_03468_));
 sg13g2_a21oi_1 _11435_ (.A1(_03452_),
    .A2(_03467_),
    .Y(_03469_),
    .B1(_03468_));
 sg13g2_or3_1 _11436_ (.A(_01471_),
    .B(_01469_),
    .C(_03469_),
    .X(_03470_));
 sg13g2_nand3b_1 _11437_ (.B(_03454_),
    .C(_03470_),
    .Y(_03471_),
    .A_N(_03410_));
 sg13g2_nand3_1 _11438_ (.B(_01474_),
    .C(_03471_),
    .A(_00347_),
    .Y(_03472_));
 sg13g2_a21oi_1 _11439_ (.A1(_03409_),
    .A2(_03472_),
    .Y(_03473_),
    .B1(_00412_));
 sg13g2_xnor2_1 _11440_ (.Y(_03474_),
    .A(_00411_),
    .B(_03473_));
 sg13g2_nor2_1 _11441_ (.A(_02922_),
    .B(_03388_),
    .Y(_03475_));
 sg13g2_nor2b_1 _11442_ (.A(_03400_),
    .B_N(_02354_),
    .Y(_03476_));
 sg13g2_buf_1 _11443_ (.A(_03476_),
    .X(_03477_));
 sg13g2_and2_1 _11444_ (.A(_02672_),
    .B(_02847_),
    .X(_03478_));
 sg13g2_buf_1 _11445_ (.A(_03478_),
    .X(_03479_));
 sg13g2_or2_1 _11446_ (.X(_03480_),
    .B(_02847_),
    .A(_02672_));
 sg13g2_buf_1 _11447_ (.A(_03480_),
    .X(_03481_));
 sg13g2_o21ai_1 _11448_ (.B1(_03481_),
    .Y(_03482_),
    .A1(_02840_),
    .A2(_03479_));
 sg13g2_nand2_1 _11449_ (.Y(_03483_),
    .A(_02899_),
    .B(_03482_));
 sg13g2_or2_1 _11450_ (.X(_03484_),
    .B(_02840_),
    .A(net26));
 sg13g2_a21oi_1 _11451_ (.A1(_02891_),
    .A2(_03481_),
    .Y(_03485_),
    .B1(_03484_));
 sg13g2_nor3_1 _11452_ (.A(net26),
    .B(_02891_),
    .C(_03479_),
    .Y(_03486_));
 sg13g2_nor2_1 _11453_ (.A(_03485_),
    .B(_03486_),
    .Y(_03487_));
 sg13g2_xnor2_1 _11454_ (.Y(_03488_),
    .A(_02922_),
    .B(_03388_));
 sg13g2_a21oi_1 _11455_ (.A1(_03483_),
    .A2(_03487_),
    .Y(_03489_),
    .B1(_03488_));
 sg13g2_or2_1 _11456_ (.X(_03490_),
    .B(_03489_),
    .A(_03396_));
 sg13g2_a22oi_1 _11457_ (.Y(_03491_),
    .B1(_03477_),
    .B2(_03490_),
    .A2(_03475_),
    .A1(_02357_));
 sg13g2_o21ai_1 _11458_ (.B1(_03479_),
    .Y(_03492_),
    .A1(net26),
    .A2(_02840_));
 sg13g2_mux2_1 _11459_ (.A0(_03484_),
    .A1(_02905_),
    .S(_03481_),
    .X(_03493_));
 sg13g2_nand2_1 _11460_ (.Y(_03494_),
    .A(_03492_),
    .B(_03493_));
 sg13g2_nor3_1 _11461_ (.A(_02899_),
    .B(_03488_),
    .C(_03494_),
    .Y(_03495_));
 sg13g2_xnor2_1 _11462_ (.Y(_03496_),
    .A(_02903_),
    .B(_03488_));
 sg13g2_nand3_1 _11463_ (.B(_03494_),
    .C(_03496_),
    .A(_02899_),
    .Y(_03497_));
 sg13g2_nand2b_1 _11464_ (.Y(_03498_),
    .B(_03497_),
    .A_N(_03495_));
 sg13g2_nand2_1 _11465_ (.Y(_03499_),
    .A(_03477_),
    .B(_03498_));
 sg13g2_xnor2_1 _11466_ (.Y(_03500_),
    .A(_03368_),
    .B(_02894_));
 sg13g2_nand2b_1 _11467_ (.Y(_03501_),
    .B(_03378_),
    .A_N(_03366_));
 sg13g2_nand3_1 _11468_ (.B(_02768_),
    .C(_03501_),
    .A(_03038_),
    .Y(_03502_));
 sg13g2_nand2_1 _11469_ (.Y(_03503_),
    .A(_03380_),
    .B(_03502_));
 sg13g2_or2_1 _11470_ (.X(_03504_),
    .B(_03503_),
    .A(_03500_));
 sg13g2_buf_1 _11471_ (.A(_03504_),
    .X(_03505_));
 sg13g2_or2_1 _11472_ (.X(_03506_),
    .B(_03475_),
    .A(_02357_));
 sg13g2_a21oi_1 _11473_ (.A1(_03396_),
    .A2(_03489_),
    .Y(_03507_),
    .B1(_03506_));
 sg13g2_nor2b_1 _11474_ (.A(_03507_),
    .B_N(_03477_),
    .Y(_03508_));
 sg13g2_nand2b_1 _11475_ (.Y(_03509_),
    .B(_03508_),
    .A_N(_03491_));
 sg13g2_and2_1 _11476_ (.A(_03477_),
    .B(_03506_),
    .X(_03510_));
 sg13g2_o21ai_1 _11477_ (.B1(_03498_),
    .Y(_03511_),
    .A1(_03396_),
    .A2(_03510_));
 sg13g2_nor2b_1 _11478_ (.A(_03508_),
    .B_N(_03511_),
    .Y(_03512_));
 sg13g2_a221oi_1 _11479_ (.B2(_03509_),
    .C1(_03512_),
    .B1(_03505_),
    .A1(_03491_),
    .Y(_03513_),
    .A2(_03499_));
 sg13g2_and2_1 _11480_ (.A(_03400_),
    .B(_03513_),
    .X(_03514_));
 sg13g2_nor2_1 _11481_ (.A(_03511_),
    .B(_03505_),
    .Y(_03515_));
 sg13g2_o21ai_1 _11482_ (.B1(_03491_),
    .Y(_03516_),
    .A1(_03499_),
    .A2(_03505_));
 sg13g2_o21ai_1 _11483_ (.B1(_03516_),
    .Y(_03517_),
    .A1(_03508_),
    .A2(_03515_));
 sg13g2_nand2b_1 _11484_ (.Y(_03518_),
    .B(_03517_),
    .A_N(_03400_));
 sg13g2_o21ai_1 _11485_ (.B1(_03518_),
    .Y(_03519_),
    .A1(_03402_),
    .A2(_03514_));
 sg13g2_nand2_1 _11486_ (.Y(_03520_),
    .A(_02251_),
    .B(_02253_));
 sg13g2_nand2_1 _11487_ (.Y(_03521_),
    .A(_02259_),
    .B(_03520_));
 sg13g2_nand2_1 _11488_ (.Y(_03522_),
    .A(_02255_),
    .B(_03521_));
 sg13g2_nand2_1 _11489_ (.Y(_03523_),
    .A(_02259_),
    .B(_02255_));
 sg13g2_nand2b_1 _11490_ (.Y(_03524_),
    .B(_03514_),
    .A_N(_03520_));
 sg13g2_nand2b_1 _11491_ (.Y(_03525_),
    .B(_03524_),
    .A_N(_02259_));
 sg13g2_a22oi_1 _11492_ (.Y(_03526_),
    .B1(_03523_),
    .B2(_03525_),
    .A2(_03522_),
    .A1(_03519_));
 sg13g2_xnor2_1 _11493_ (.Y(_03527_),
    .A(_02163_),
    .B(_03526_));
 sg13g2_nand3_1 _11494_ (.B(_03474_),
    .C(_03527_),
    .A(_03408_),
    .Y(_03528_));
 sg13g2_or3_1 _11495_ (.A(_03408_),
    .B(_03474_),
    .C(_03527_),
    .X(_03529_));
 sg13g2_xnor2_1 _11496_ (.Y(_03530_),
    .A(_00351_),
    .B(_00389_));
 sg13g2_xnor2_1 _11497_ (.Y(_03531_),
    .A(_00347_),
    .B(_03530_));
 sg13g2_xnor2_1 _11498_ (.Y(_03532_),
    .A(_01481_),
    .B(_03531_));
 sg13g2_nand3_1 _11499_ (.B(_03520_),
    .C(_02255_),
    .A(_02259_),
    .Y(_03533_));
 sg13g2_o21ai_1 _11500_ (.B1(_03533_),
    .Y(_03534_),
    .A1(_02259_),
    .A2(_02253_));
 sg13g2_xor2_1 _11501_ (.B(_03534_),
    .A(_03403_),
    .X(_03535_));
 sg13g2_nand2_1 _11502_ (.Y(_03536_),
    .A(_03532_),
    .B(_03535_));
 sg13g2_nand2_1 _11503_ (.Y(_03537_),
    .A(_00715_),
    .B(_01466_));
 sg13g2_a21o_1 _11504_ (.A2(_03537_),
    .A1(_01472_),
    .B1(_03452_),
    .X(_03538_));
 sg13g2_nand2b_1 _11505_ (.Y(_03539_),
    .B(_03467_),
    .A_N(_01471_));
 sg13g2_nand2_1 _11506_ (.Y(_03540_),
    .A(_01466_),
    .B(_03539_));
 sg13g2_a21o_1 _11507_ (.A2(_03540_),
    .A1(_03538_),
    .B1(_03410_),
    .X(_03541_));
 sg13g2_inv_1 _11508_ (.Y(_03542_),
    .A(_01469_));
 sg13g2_a22oi_1 _11509_ (.Y(_03543_),
    .B1(_03541_),
    .B2(_03542_),
    .A2(_03538_),
    .A1(_03410_));
 sg13g2_nor2_1 _11510_ (.A(_01438_),
    .B(_01439_),
    .Y(_03544_));
 sg13g2_xnor2_1 _11511_ (.Y(_03545_),
    .A(_03544_),
    .B(_01474_));
 sg13g2_xnor2_1 _11512_ (.Y(_03546_),
    .A(_03543_),
    .B(_03545_));
 sg13g2_buf_1 _11513_ (.A(_03546_),
    .X(_03547_));
 sg13g2_nand2_1 _11514_ (.Y(_03548_),
    .A(_03536_),
    .B(_03547_));
 sg13g2_xor2_1 _11515_ (.B(_03400_),
    .A(_03402_),
    .X(_03549_));
 sg13g2_xnor2_1 _11516_ (.Y(_03550_),
    .A(_03513_),
    .B(_03549_));
 sg13g2_buf_2 _11517_ (.A(_03550_),
    .X(_03551_));
 sg13g2_nand2_1 _11518_ (.Y(_03552_),
    .A(_03536_),
    .B(_03551_));
 sg13g2_nor2b_1 _11519_ (.A(_02908_),
    .B_N(_03383_),
    .Y(_03553_));
 sg13g2_o21ai_1 _11520_ (.B1(_02922_),
    .Y(_03554_),
    .A1(_03388_),
    .A2(_03553_));
 sg13g2_nand2_1 _11521_ (.Y(_03555_),
    .A(_03388_),
    .B(_03553_));
 sg13g2_a22oi_1 _11522_ (.Y(_03556_),
    .B1(_03554_),
    .B2(_03555_),
    .A2(_02357_),
    .A1(_03396_));
 sg13g2_nor2_1 _11523_ (.A(_03396_),
    .B(_02357_),
    .Y(_03557_));
 sg13g2_nor2_1 _11524_ (.A(_03556_),
    .B(_03557_),
    .Y(_03558_));
 sg13g2_xnor2_1 _11525_ (.Y(_03559_),
    .A(_03477_),
    .B(_03558_));
 sg13g2_xor2_1 _11526_ (.B(_03410_),
    .A(_01469_),
    .X(_03560_));
 sg13g2_nand2_1 _11527_ (.Y(_03561_),
    .A(_01471_),
    .B(_01466_));
 sg13g2_nor3_1 _11528_ (.A(_00912_),
    .B(_01432_),
    .C(_00714_),
    .Y(_03562_));
 sg13g2_o21ai_1 _11529_ (.B1(_00714_),
    .Y(_03563_),
    .A1(_00912_),
    .A2(_01432_));
 sg13g2_o21ai_1 _11530_ (.B1(_03563_),
    .Y(_03564_),
    .A1(_00708_),
    .A2(_03562_));
 sg13g2_nor2_1 _11531_ (.A(_01471_),
    .B(_01466_),
    .Y(_03565_));
 sg13g2_a21oi_1 _11532_ (.A1(_03561_),
    .A2(_03564_),
    .Y(_03566_),
    .B1(_03565_));
 sg13g2_a21o_1 _11533_ (.A2(_03563_),
    .A1(_00708_),
    .B1(_03562_),
    .X(_03567_));
 sg13g2_a21o_1 _11534_ (.A2(_01433_),
    .A1(_00708_),
    .B1(_01466_),
    .X(_03568_));
 sg13g2_a221oi_1 _11535_ (.B2(_01471_),
    .C1(_03560_),
    .B1(_03568_),
    .A1(_01466_),
    .Y(_03569_),
    .A2(_03567_));
 sg13g2_a21oi_1 _11536_ (.A1(_03560_),
    .A2(_03566_),
    .Y(_03570_),
    .B1(_03569_));
 sg13g2_buf_1 _11537_ (.A(_03570_),
    .X(_03571_));
 sg13g2_nand2_1 _11538_ (.Y(_03572_),
    .A(_03559_),
    .B(_03571_));
 sg13g2_nor2_1 _11539_ (.A(_02899_),
    .B(_02902_),
    .Y(_03573_));
 sg13g2_o21ai_1 _11540_ (.B1(_02900_),
    .Y(_03574_),
    .A1(_02906_),
    .A2(_03573_));
 sg13g2_nand3_1 _11541_ (.B(_02898_),
    .C(_03574_),
    .A(_03383_),
    .Y(_03575_));
 sg13g2_nor2_1 _11542_ (.A(net24),
    .B(_02902_),
    .Y(_03576_));
 sg13g2_xnor2_1 _11543_ (.Y(_03577_),
    .A(_03576_),
    .B(_03488_));
 sg13g2_xnor2_1 _11544_ (.Y(_03578_),
    .A(_03575_),
    .B(_03577_));
 sg13g2_xor2_1 _11545_ (.B(_00714_),
    .A(_00708_),
    .X(_03579_));
 sg13g2_xnor2_1 _11546_ (.Y(_03580_),
    .A(_01433_),
    .B(_03579_));
 sg13g2_buf_1 _11547_ (.A(_03580_),
    .X(_03581_));
 sg13g2_nor2b_1 _11548_ (.A(_03578_),
    .B_N(_03581_),
    .Y(_03582_));
 sg13g2_buf_2 _11549_ (.A(_03582_),
    .X(_03583_));
 sg13g2_inv_4 _11550_ (.A(_03583_),
    .Y(_03584_));
 sg13g2_nand2b_1 _11551_ (.Y(_03585_),
    .B(_03578_),
    .A_N(_03581_));
 sg13g2_buf_8 _11552_ (.A(_03585_),
    .X(_03586_));
 sg13g2_xnor2_1 _11553_ (.Y(_03587_),
    .A(net24),
    .B(_03494_));
 sg13g2_xnor2_1 _11554_ (.Y(_03588_),
    .A(_03505_),
    .B(_03587_));
 sg13g2_buf_2 _11555_ (.A(_03588_),
    .X(_03589_));
 sg13g2_inv_4 _11556_ (.A(_03589_),
    .Y(_03590_));
 sg13g2_nand3_1 _11557_ (.B(net52),
    .C(net22),
    .A(net23),
    .Y(_03591_));
 sg13g2_nor2_1 _11558_ (.A(_00890_),
    .B(net22),
    .Y(_03592_));
 sg13g2_and2_1 _11559_ (.A(_00890_),
    .B(net22),
    .X(_03593_));
 sg13g2_buf_1 _11560_ (.A(_03593_),
    .X(_03594_));
 sg13g2_nor2_1 _11561_ (.A(net52),
    .B(_03594_),
    .Y(_03595_));
 sg13g2_o21ai_1 _11562_ (.B1(_01426_),
    .Y(_03596_),
    .A1(_03592_),
    .A2(_03595_));
 sg13g2_a21o_1 _11563_ (.A2(_03596_),
    .A1(_03591_),
    .B1(_03461_),
    .X(_03597_));
 sg13g2_mux2_1 _11564_ (.A0(_03592_),
    .A1(_03594_),
    .S(net23),
    .X(_03598_));
 sg13g2_nor3_1 _11565_ (.A(_01426_),
    .B(_03592_),
    .C(_03594_),
    .Y(_03599_));
 sg13g2_mux2_1 _11566_ (.A0(_03598_),
    .A1(_03599_),
    .S(net52),
    .X(_03600_));
 sg13g2_nand2b_1 _11567_ (.Y(_03601_),
    .B(_03600_),
    .A_N(_03455_));
 sg13g2_nand3_1 _11568_ (.B(_03597_),
    .C(_03601_),
    .A(_03440_),
    .Y(_03602_));
 sg13g2_xnor2_1 _11569_ (.Y(_03603_),
    .A(_03450_),
    .B(_03602_));
 sg13g2_or2_1 _11570_ (.X(_03604_),
    .B(_03603_),
    .A(_03590_));
 sg13g2_buf_1 _11571_ (.A(_03604_),
    .X(_03605_));
 sg13g2_nand2_1 _11572_ (.Y(_03606_),
    .A(_03586_),
    .B(_03605_));
 sg13g2_buf_8 _11573_ (.A(_03603_),
    .X(_03607_));
 sg13g2_a22oi_1 _11574_ (.Y(_03608_),
    .B1(_01125_),
    .B2(_01419_),
    .A2(_01106_),
    .A1(_00927_));
 sg13g2_a221oi_1 _11575_ (.B2(_01421_),
    .C1(_03416_),
    .B1(_03442_),
    .A1(_00892_),
    .Y(_03609_),
    .A2(_01422_));
 sg13g2_xnor2_1 _11576_ (.Y(_03610_),
    .A(_01426_),
    .B(_03609_));
 sg13g2_xnor2_1 _11577_ (.Y(_03611_),
    .A(_03608_),
    .B(_03610_));
 sg13g2_buf_1 _11578_ (.A(_03611_),
    .X(_03612_));
 sg13g2_xor2_1 _11579_ (.B(_03503_),
    .A(_03500_),
    .X(_03613_));
 sg13g2_inv_2 _11580_ (.Y(_03614_),
    .A(_03613_));
 sg13g2_nand2b_1 _11581_ (.Y(_03615_),
    .B(_03614_),
    .A_N(_03612_));
 sg13g2_buf_1 _11582_ (.A(_03615_),
    .X(_03616_));
 sg13g2_nand2_1 _11583_ (.Y(_03617_),
    .A(_03038_),
    .B(_03378_));
 sg13g2_nor2_1 _11584_ (.A(_03366_),
    .B(_03617_),
    .Y(_03618_));
 sg13g2_nand2_1 _11585_ (.Y(_03619_),
    .A(_02768_),
    .B(_03380_));
 sg13g2_xnor2_1 _11586_ (.Y(_03620_),
    .A(_03038_),
    .B(_03619_));
 sg13g2_xnor2_1 _11587_ (.Y(_03621_),
    .A(_03618_),
    .B(_03620_));
 sg13g2_buf_1 _11588_ (.A(_03621_),
    .X(_03622_));
 sg13g2_nor2_1 _11589_ (.A(_01417_),
    .B(_01418_),
    .Y(_03623_));
 sg13g2_a21oi_1 _11590_ (.A1(_01098_),
    .A2(_03438_),
    .Y(_03624_),
    .B1(_03437_));
 sg13g2_xnor2_1 _11591_ (.Y(_03625_),
    .A(_03623_),
    .B(_03624_));
 sg13g2_buf_1 _11592_ (.A(_03625_),
    .X(_03626_));
 sg13g2_nor2b_1 _11593_ (.A(net21),
    .B_N(net19),
    .Y(_03627_));
 sg13g2_xnor2_1 _11594_ (.Y(_03628_),
    .A(_01125_),
    .B(_03434_));
 sg13g2_xor2_1 _11595_ (.B(_03617_),
    .A(_03366_),
    .X(_03629_));
 sg13g2_inv_1 _11596_ (.Y(_03630_),
    .A(_03629_));
 sg13g2_xnor2_1 _11597_ (.Y(_03631_),
    .A(_01127_),
    .B(_01412_));
 sg13g2_buf_1 _11598_ (.A(_03631_),
    .X(_03632_));
 sg13g2_xnor2_1 _11599_ (.Y(_03633_),
    .A(_03360_),
    .B(_03345_));
 sg13g2_xnor2_1 _11600_ (.Y(_03634_),
    .A(_03359_),
    .B(_03633_));
 sg13g2_xnor2_1 _11601_ (.Y(_03635_),
    .A(_03344_),
    .B(_03634_));
 sg13g2_buf_2 _11602_ (.A(_03635_),
    .X(_03636_));
 sg13g2_xor2_1 _11603_ (.B(_01409_),
    .A(_01404_),
    .X(_03637_));
 sg13g2_xnor2_1 _11604_ (.Y(_03638_),
    .A(_01398_),
    .B(_03637_));
 sg13g2_buf_1 _11605_ (.A(_03638_),
    .X(_03639_));
 sg13g2_xor2_1 _11606_ (.B(_03330_),
    .A(_03341_),
    .X(_03640_));
 sg13g2_xnor2_1 _11607_ (.Y(_03641_),
    .A(_03172_),
    .B(_03640_));
 sg13g2_buf_2 _11608_ (.A(_03641_),
    .X(_03642_));
 sg13g2_nor2b_1 _11609_ (.A(_03639_),
    .B_N(_03642_),
    .Y(_03643_));
 sg13g2_nor2_1 _11610_ (.A(_03224_),
    .B(_03324_),
    .Y(_03644_));
 sg13g2_nor2_1 _11611_ (.A(_03328_),
    .B(_03329_),
    .Y(_03645_));
 sg13g2_xnor2_1 _11612_ (.Y(_03646_),
    .A(_03644_),
    .B(_03645_));
 sg13g2_buf_1 _11613_ (.A(_03646_),
    .X(_03647_));
 sg13g2_xor2_1 _11614_ (.B(_01393_),
    .A(_01386_),
    .X(_03648_));
 sg13g2_xnor2_1 _11615_ (.Y(_03649_),
    .A(_01199_),
    .B(_03648_));
 sg13g2_xor2_1 _11616_ (.B(_03323_),
    .A(_03220_),
    .X(_03650_));
 sg13g2_xor2_1 _11617_ (.B(_03650_),
    .A(_03223_),
    .X(_03651_));
 sg13g2_nand2_1 _11618_ (.Y(_03652_),
    .A(_03649_),
    .B(_03651_));
 sg13g2_nand2_1 _11619_ (.Y(_03653_),
    .A(net25),
    .B(_03652_));
 sg13g2_xnor2_1 _11620_ (.Y(_03654_),
    .A(_01197_),
    .B(_01396_));
 sg13g2_buf_1 _11621_ (.A(_03654_),
    .X(_03655_));
 sg13g2_o21ai_1 _11622_ (.B1(_03655_),
    .Y(_03656_),
    .A1(net25),
    .A2(_03652_));
 sg13g2_nand2_1 _11623_ (.Y(_03657_),
    .A(_03653_),
    .B(_03656_));
 sg13g2_nand2b_1 _11624_ (.Y(_03658_),
    .B(_03639_),
    .A_N(_03642_));
 sg13g2_o21ai_1 _11625_ (.B1(_03658_),
    .Y(_03659_),
    .A1(_03643_),
    .A2(_03657_));
 sg13g2_and2_1 _11626_ (.A(_03636_),
    .B(_03659_),
    .X(_03660_));
 sg13g2_or2_1 _11627_ (.X(_03661_),
    .B(_03659_),
    .A(_03636_));
 sg13g2_buf_1 _11628_ (.A(_03661_),
    .X(_03662_));
 sg13g2_o21ai_1 _11629_ (.B1(_03662_),
    .Y(_03663_),
    .A1(_03632_),
    .A2(_03660_));
 sg13g2_o21ai_1 _11630_ (.B1(_03663_),
    .Y(_03664_),
    .A1(_03628_),
    .A2(_03630_));
 sg13g2_buf_1 _11631_ (.A(_03664_),
    .X(_03665_));
 sg13g2_nand2_1 _11632_ (.Y(_03666_),
    .A(_03628_),
    .B(_03630_));
 sg13g2_nor2b_1 _11633_ (.A(net19),
    .B_N(net21),
    .Y(_03667_));
 sg13g2_a21oi_1 _11634_ (.A1(_03665_),
    .A2(_03666_),
    .Y(_03668_),
    .B1(_03667_));
 sg13g2_nand2_1 _11635_ (.Y(_03669_),
    .A(_03612_),
    .B(_03613_));
 sg13g2_o21ai_1 _11636_ (.B1(_03669_),
    .Y(_03670_),
    .A1(_03627_),
    .A2(_03668_));
 sg13g2_a22oi_1 _11637_ (.Y(_03671_),
    .B1(_03616_),
    .B2(_03670_),
    .A2(_03607_),
    .A1(_03590_));
 sg13g2_or2_1 _11638_ (.X(_03672_),
    .B(_03671_),
    .A(_03606_));
 sg13g2_nand2b_1 _11639_ (.Y(_03673_),
    .B(_03498_),
    .A_N(_03505_));
 sg13g2_nand2b_1 _11640_ (.Y(_03674_),
    .B(_03673_),
    .A_N(_03489_));
 sg13g2_xor2_1 _11641_ (.B(_03475_),
    .A(_02357_),
    .X(_03675_));
 sg13g2_xnor2_1 _11642_ (.Y(_03676_),
    .A(_03396_),
    .B(_03675_));
 sg13g2_xor2_1 _11643_ (.B(_03676_),
    .A(_03674_),
    .X(_03677_));
 sg13g2_buf_1 _11644_ (.A(_03677_),
    .X(_03678_));
 sg13g2_o21ai_1 _11645_ (.B1(_03467_),
    .Y(_03679_),
    .A1(_03468_),
    .A2(_03452_));
 sg13g2_nor2b_1 _11646_ (.A(_03565_),
    .B_N(_03561_),
    .Y(_03680_));
 sg13g2_xnor2_1 _11647_ (.Y(_03681_),
    .A(_03679_),
    .B(_03680_));
 sg13g2_buf_2 _11648_ (.A(_03681_),
    .X(_03682_));
 sg13g2_a22oi_1 _11649_ (.Y(_03683_),
    .B1(_03678_),
    .B2(_03682_),
    .A2(_03672_),
    .A1(_03584_));
 sg13g2_nor2_1 _11650_ (.A(_03682_),
    .B(_03678_),
    .Y(_03684_));
 sg13g2_or2_1 _11651_ (.X(_03685_),
    .B(_03684_),
    .A(_03683_));
 sg13g2_nor2_1 _11652_ (.A(_03559_),
    .B(_03571_),
    .Y(_03686_));
 sg13g2_a221oi_1 _11653_ (.B2(_03685_),
    .C1(_03686_),
    .B1(_03572_),
    .A1(_03548_),
    .Y(_03687_),
    .A2(_03552_));
 sg13g2_inv_1 _11654_ (.Y(_03688_),
    .A(_03551_));
 sg13g2_nor2_1 _11655_ (.A(_03532_),
    .B(_03535_),
    .Y(_03689_));
 sg13g2_inv_1 _11656_ (.Y(_03690_),
    .A(_03689_));
 sg13g2_o21ai_1 _11657_ (.B1(_03690_),
    .Y(_03691_),
    .A1(_03548_),
    .A2(_03688_));
 sg13g2_nor2_1 _11658_ (.A(_03687_),
    .B(_03691_),
    .Y(_03692_));
 sg13g2_a21o_1 _11659_ (.A2(_03529_),
    .A1(_03528_),
    .B1(_03692_),
    .X(_03693_));
 sg13g2_buf_1 _11660_ (.A(_03693_),
    .X(_03694_));
 sg13g2_nand2_1 _11661_ (.Y(_03695_),
    .A(_03590_),
    .B(net20));
 sg13g2_and2_1 _11662_ (.A(_03612_),
    .B(_03613_),
    .X(_03696_));
 sg13g2_buf_1 _11663_ (.A(_03696_),
    .X(_03697_));
 sg13g2_nand2b_1 _11664_ (.Y(_03698_),
    .B(net21),
    .A_N(net19));
 sg13g2_nand2b_1 _11665_ (.Y(_03699_),
    .B(net19),
    .A_N(net21));
 sg13g2_nand3_1 _11666_ (.B(_03665_),
    .C(_03666_),
    .A(_03699_),
    .Y(_03700_));
 sg13g2_nor2_1 _11667_ (.A(_03612_),
    .B(_03613_),
    .Y(_03701_));
 sg13g2_a21oi_1 _11668_ (.A1(_03698_),
    .A2(_03700_),
    .Y(_03702_),
    .B1(_03701_));
 sg13g2_o21ai_1 _11669_ (.B1(_03605_),
    .Y(_03703_),
    .A1(net18),
    .A2(_03702_));
 sg13g2_nor2b_1 _11670_ (.A(_03581_),
    .B_N(_03578_),
    .Y(_03704_));
 sg13g2_a21o_1 _11671_ (.A2(_03703_),
    .A1(_03695_),
    .B1(_03704_),
    .X(_03705_));
 sg13g2_xor2_1 _11672_ (.B(_03680_),
    .A(_03679_),
    .X(_03706_));
 sg13g2_buf_8 _11673_ (.A(_03706_),
    .X(_03707_));
 sg13g2_xnor2_1 _11674_ (.Y(_03708_),
    .A(_03674_),
    .B(_03676_));
 sg13g2_nor2_1 _11675_ (.A(_03707_),
    .B(_03708_),
    .Y(_03709_));
 sg13g2_a21oi_1 _11676_ (.A1(_03584_),
    .A2(_03705_),
    .Y(_03710_),
    .B1(_03709_));
 sg13g2_or2_1 _11677_ (.X(_03711_),
    .B(_03686_),
    .A(_03684_));
 sg13g2_or2_1 _11678_ (.X(_03712_),
    .B(_03711_),
    .A(_03710_));
 sg13g2_a221oi_1 _11679_ (.B2(_03712_),
    .C1(_03688_),
    .B1(_03572_),
    .A1(_03532_),
    .Y(_03713_),
    .A2(_03535_));
 sg13g2_inv_1 _11680_ (.Y(_03714_),
    .A(_03571_));
 sg13g2_a21oi_1 _11681_ (.A1(_03707_),
    .A2(_03708_),
    .Y(_03715_),
    .B1(_03583_));
 sg13g2_and3_1 _11682_ (.X(_03716_),
    .A(_03699_),
    .B(_03665_),
    .C(_03666_));
 sg13g2_nor4_1 _11683_ (.A(_03607_),
    .B(net18),
    .C(_03667_),
    .D(_03716_),
    .Y(_03717_));
 sg13g2_a21oi_1 _11684_ (.A1(_03590_),
    .A2(_03616_),
    .Y(_03718_),
    .B1(net20));
 sg13g2_nor3_1 _11685_ (.A(_03590_),
    .B(_03616_),
    .C(_03697_),
    .Y(_03719_));
 sg13g2_nor4_1 _11686_ (.A(_03590_),
    .B(_03697_),
    .C(_03667_),
    .D(_03716_),
    .Y(_03720_));
 sg13g2_or4_1 _11687_ (.A(_03717_),
    .B(_03718_),
    .C(_03719_),
    .D(_03720_),
    .X(_03721_));
 sg13g2_o21ai_1 _11688_ (.B1(_03708_),
    .Y(_03722_),
    .A1(_03707_),
    .A2(_03586_));
 sg13g2_nand2_1 _11689_ (.Y(_03723_),
    .A(_03707_),
    .B(_03586_));
 sg13g2_a22oi_1 _11690_ (.Y(_03724_),
    .B1(_03722_),
    .B2(_03723_),
    .A2(_03721_),
    .A1(_03715_));
 sg13g2_inv_2 _11691_ (.Y(_03725_),
    .A(_03559_));
 sg13g2_o21ai_1 _11692_ (.B1(_03725_),
    .Y(_03726_),
    .A1(_03714_),
    .A2(_03724_));
 sg13g2_nand2_1 _11693_ (.Y(_03727_),
    .A(_03714_),
    .B(_03724_));
 sg13g2_a21oi_1 _11694_ (.A1(_03726_),
    .A2(_03727_),
    .Y(_03728_),
    .B1(_03551_));
 sg13g2_o21ai_1 _11695_ (.B1(_03690_),
    .Y(_03729_),
    .A1(_03548_),
    .A2(_03728_));
 sg13g2_o21ai_1 _11696_ (.B1(_03408_),
    .Y(_03730_),
    .A1(_03713_),
    .A2(_03729_));
 sg13g2_or3_1 _11697_ (.A(_03408_),
    .B(_03713_),
    .C(_03729_),
    .X(_03731_));
 sg13g2_xor2_1 _11698_ (.B(_03527_),
    .A(_03474_),
    .X(_03732_));
 sg13g2_nand4_1 _11699_ (.B(_03730_),
    .C(_03731_),
    .A(_03692_),
    .Y(_03733_),
    .D(_03732_));
 sg13g2_buf_1 _11700_ (.A(_03733_),
    .X(_03734_));
 sg13g2_and2_1 _11701_ (.A(_03694_),
    .B(_03734_),
    .X(_03735_));
 sg13g2_buf_8 _11702_ (.A(_03735_),
    .X(_03736_));
 sg13g2_buf_2 _11703_ (.A(\iter[0] ),
    .X(_03737_));
 sg13g2_buf_1 _11704_ (.A(\iter[1] ),
    .X(_03738_));
 sg13g2_nor2_1 _11705_ (.A(_03701_),
    .B(net18),
    .Y(_03739_));
 sg13g2_nand2_1 _11706_ (.Y(_03740_),
    .A(_03665_),
    .B(_03666_));
 sg13g2_nand3b_1 _11707_ (.B(_03627_),
    .C(_03740_),
    .Y(_03741_),
    .A_N(_03739_));
 sg13g2_nor3_1 _11708_ (.A(net21),
    .B(net19),
    .C(_03740_),
    .Y(_03742_));
 sg13g2_xor2_1 _11709_ (.B(_03740_),
    .A(net19),
    .X(_03743_));
 sg13g2_and2_1 _11710_ (.A(net21),
    .B(_03743_),
    .X(_03744_));
 sg13g2_o21ai_1 _11711_ (.B1(_03739_),
    .Y(_03745_),
    .A1(_03742_),
    .A2(_03744_));
 sg13g2_nand2_1 _11712_ (.Y(_03746_),
    .A(_03636_),
    .B(_03659_));
 sg13g2_and3_1 _11713_ (.X(_03747_),
    .A(_03662_),
    .B(_03632_),
    .C(_03746_));
 sg13g2_nor2_1 _11714_ (.A(_03632_),
    .B(_03746_),
    .Y(_03748_));
 sg13g2_xnor2_1 _11715_ (.Y(_03749_),
    .A(_01125_),
    .B(_01413_));
 sg13g2_xnor2_1 _11716_ (.Y(_03750_),
    .A(_03749_),
    .B(_03630_));
 sg13g2_o21ai_1 _11717_ (.B1(_03750_),
    .Y(_03751_),
    .A1(_03747_),
    .A2(_03748_));
 sg13g2_or3_1 _11718_ (.A(_03662_),
    .B(_03632_),
    .C(_03750_),
    .X(_03752_));
 sg13g2_and2_1 _11719_ (.A(_03649_),
    .B(_03651_),
    .X(_03753_));
 sg13g2_inv_1 _11720_ (.Y(_03754_),
    .A(_03655_));
 sg13g2_nor2_1 _11721_ (.A(net25),
    .B(_03754_),
    .Y(_03755_));
 sg13g2_nand2_1 _11722_ (.Y(_03756_),
    .A(net25),
    .B(_03754_));
 sg13g2_nand2b_1 _11723_ (.Y(_03757_),
    .B(_03756_),
    .A_N(_03755_));
 sg13g2_nor2_1 _11724_ (.A(_03649_),
    .B(_03651_),
    .Y(_03758_));
 sg13g2_nor2_1 _11725_ (.A(_03647_),
    .B(_03655_),
    .Y(_03759_));
 sg13g2_a22oi_1 _11726_ (.Y(_03760_),
    .B1(_03758_),
    .B2(_03759_),
    .A2(_03757_),
    .A1(_03753_));
 sg13g2_nand3_1 _11727_ (.B(_03655_),
    .C(_03758_),
    .A(net25),
    .Y(_03761_));
 sg13g2_xor2_1 _11728_ (.B(_03639_),
    .A(_03642_),
    .X(_03762_));
 sg13g2_mux2_1 _11729_ (.A0(_03760_),
    .A1(_03761_),
    .S(_03762_),
    .X(_03763_));
 sg13g2_a221oi_1 _11730_ (.B2(_03752_),
    .C1(_03763_),
    .B1(_03751_),
    .A1(_03741_),
    .Y(_03764_),
    .A2(_03745_));
 sg13g2_nand2_1 _11731_ (.Y(_03765_),
    .A(_03584_),
    .B(_03586_));
 sg13g2_nand3_1 _11732_ (.B(_03698_),
    .C(_03700_),
    .A(_03669_),
    .Y(_03766_));
 sg13g2_nand2_1 _11733_ (.Y(_03767_),
    .A(_03616_),
    .B(_03766_));
 sg13g2_or2_1 _11734_ (.X(_03768_),
    .B(_03709_),
    .A(_03684_));
 sg13g2_or3_1 _11735_ (.A(_03765_),
    .B(_03767_),
    .C(_03768_),
    .X(_03769_));
 sg13g2_nand2_1 _11736_ (.Y(_03770_),
    .A(_03765_),
    .B(_03767_));
 sg13g2_nand2_1 _11737_ (.Y(_03771_),
    .A(_03589_),
    .B(net20));
 sg13g2_nor2_1 _11738_ (.A(_03589_),
    .B(net20),
    .Y(_03772_));
 sg13g2_inv_1 _11739_ (.Y(_03773_),
    .A(_03772_));
 sg13g2_nor3_1 _11740_ (.A(_03701_),
    .B(_03627_),
    .C(_03668_),
    .Y(_03774_));
 sg13g2_nor2_1 _11741_ (.A(net18),
    .B(_03774_),
    .Y(_03775_));
 sg13g2_a221oi_1 _11742_ (.B2(_03773_),
    .C1(_03775_),
    .B1(_03771_),
    .A1(_03769_),
    .Y(_03776_),
    .A2(_03770_));
 sg13g2_a21oi_1 _11743_ (.A1(_03584_),
    .A2(_03586_),
    .Y(_03777_),
    .B1(_03605_));
 sg13g2_nor2_1 _11744_ (.A(_03695_),
    .B(_03765_),
    .Y(_03778_));
 sg13g2_o21ai_1 _11745_ (.B1(_03775_),
    .Y(_03779_),
    .A1(_03777_),
    .A2(_03778_));
 sg13g2_nand2b_1 _11746_ (.Y(_03780_),
    .B(_03779_),
    .A_N(_03776_));
 sg13g2_and2_1 _11747_ (.A(_03725_),
    .B(_03571_),
    .X(_03781_));
 sg13g2_buf_1 _11748_ (.A(_03781_),
    .X(_03782_));
 sg13g2_nor2_1 _11749_ (.A(_03725_),
    .B(_03571_),
    .Y(_03783_));
 sg13g2_or2_1 _11750_ (.X(_03784_),
    .B(_03783_),
    .A(_03782_));
 sg13g2_buf_1 _11751_ (.A(_03784_),
    .X(_03785_));
 sg13g2_or2_1 _11752_ (.X(_03786_),
    .B(_03684_),
    .A(_03583_));
 sg13g2_nor3_1 _11753_ (.A(net20),
    .B(net18),
    .C(_03702_),
    .Y(_03787_));
 sg13g2_o21ai_1 _11754_ (.B1(net20),
    .Y(_03788_),
    .A1(net18),
    .A2(_03702_));
 sg13g2_o21ai_1 _11755_ (.B1(_03788_),
    .Y(_03789_),
    .A1(_03589_),
    .A2(_03787_));
 sg13g2_and2_1 _11756_ (.A(_03586_),
    .B(_03789_),
    .X(_03790_));
 sg13g2_o21ai_1 _11757_ (.B1(_03785_),
    .Y(_03791_),
    .A1(_03786_),
    .A2(_03790_));
 sg13g2_o21ai_1 _11758_ (.B1(_03791_),
    .Y(_03792_),
    .A1(_03710_),
    .A2(_03785_));
 sg13g2_nand2_1 _11759_ (.Y(_03793_),
    .A(_03707_),
    .B(_03678_));
 sg13g2_nand2_1 _11760_ (.Y(_03794_),
    .A(_03682_),
    .B(_03708_));
 sg13g2_o21ai_1 _11761_ (.B1(net20),
    .Y(_03795_),
    .A1(net18),
    .A2(_03774_));
 sg13g2_nor3_1 _11762_ (.A(net20),
    .B(net18),
    .C(_03774_),
    .Y(_03796_));
 sg13g2_a21oi_1 _11763_ (.A1(_03589_),
    .A2(_03795_),
    .Y(_03797_),
    .B1(_03796_));
 sg13g2_o21ai_1 _11764_ (.B1(_03586_),
    .Y(_03798_),
    .A1(_03583_),
    .A2(_03797_));
 sg13g2_a21o_1 _11765_ (.A2(_03794_),
    .A1(_03793_),
    .B1(_03798_),
    .X(_03799_));
 sg13g2_a21o_1 _11766_ (.A2(_03695_),
    .A1(_03584_),
    .B1(_03704_),
    .X(_03800_));
 sg13g2_nand2_1 _11767_ (.Y(_03801_),
    .A(_03709_),
    .B(_03800_));
 sg13g2_or2_1 _11768_ (.X(_03802_),
    .B(_03801_),
    .A(_03785_));
 sg13g2_nand3_1 _11769_ (.B(_03785_),
    .C(_03800_),
    .A(_03684_),
    .Y(_03803_));
 sg13g2_nand3_1 _11770_ (.B(_03802_),
    .C(_03803_),
    .A(_03799_),
    .Y(_03804_));
 sg13g2_and4_1 _11771_ (.A(_03764_),
    .B(_03780_),
    .C(_03792_),
    .D(_03804_),
    .X(_03805_));
 sg13g2_buf_1 _11772_ (.A(_03805_),
    .X(_03806_));
 sg13g2_xnor2_1 _11773_ (.Y(_03807_),
    .A(_03547_),
    .B(_03551_));
 sg13g2_nor2_1 _11774_ (.A(_03682_),
    .B(_03704_),
    .Y(_03808_));
 sg13g2_o21ai_1 _11775_ (.B1(_03808_),
    .Y(_03809_),
    .A1(_03583_),
    .A2(_03797_));
 sg13g2_a22oi_1 _11776_ (.Y(_03810_),
    .B1(_03809_),
    .B2(_03678_),
    .A2(_03798_),
    .A1(_03682_));
 sg13g2_o21ai_1 _11777_ (.B1(_03572_),
    .Y(_03811_),
    .A1(_03686_),
    .A2(_03810_));
 sg13g2_xnor2_1 _11778_ (.Y(_03812_),
    .A(_03807_),
    .B(_03811_));
 sg13g2_and2_1 _11779_ (.A(_03536_),
    .B(_03690_),
    .X(_03813_));
 sg13g2_buf_1 _11780_ (.A(_03813_),
    .X(_03814_));
 sg13g2_o21ai_1 _11781_ (.B1(_03572_),
    .Y(_03815_),
    .A1(_03710_),
    .A2(_03711_));
 sg13g2_a21o_1 _11782_ (.A2(_03727_),
    .A1(_03726_),
    .B1(_03551_),
    .X(_03816_));
 sg13g2_a22oi_1 _11783_ (.Y(_03817_),
    .B1(_03816_),
    .B2(_03547_),
    .A2(_03815_),
    .A1(_03551_));
 sg13g2_xnor2_1 _11784_ (.Y(_03818_),
    .A(_03814_),
    .B(_03817_));
 sg13g2_a21o_1 _11785_ (.A2(_03812_),
    .A1(_03806_),
    .B1(_03818_),
    .X(_03819_));
 sg13g2_nand4_1 _11786_ (.B(_03737_),
    .C(_03738_),
    .A(\iter[2] ),
    .Y(_03820_),
    .D(_03819_));
 sg13g2_or2_1 _11787_ (.X(_03821_),
    .B(_03820_),
    .A(_03736_));
 sg13g2_buf_1 _11788_ (.A(_03821_),
    .X(_03822_));
 sg13g2_nor3_1 _11789_ (.A(_04458_),
    .B(_04439_),
    .C(_03822_),
    .Y(_03823_));
 sg13g2_a21o_1 _11790_ (.A2(_04439_),
    .A1(\last_iter[4] ),
    .B1(_03823_),
    .X(_03824_));
 sg13g2_buf_1 _11791_ (.A(_03824_),
    .X(_00000_));
 sg13g2_and2_1 _11792_ (.A(\last_iter[3] ),
    .B(_04439_),
    .X(_03825_));
 sg13g2_o21ai_1 _11793_ (.B1(_04449_),
    .Y(_03826_),
    .A1(_03736_),
    .A2(_03820_));
 sg13g2_or3_1 _11794_ (.A(_04449_),
    .B(_03736_),
    .C(_03820_),
    .X(_03827_));
 sg13g2_a21oi_1 _11795_ (.A1(_03826_),
    .A2(_03827_),
    .Y(_03828_),
    .B1(_04439_));
 sg13g2_nor2_2 _11796_ (.A(_03825_),
    .B(_03828_),
    .Y(_03829_));
 sg13g2_inv_4 _11797_ (.A(_03829_),
    .Y(_00015_));
 sg13g2_inv_1 _11798_ (.Y(_03830_),
    .A(\last_iter[1] ));
 sg13g2_xor2_1 _11799_ (.B(_03817_),
    .A(_03814_),
    .X(_03831_));
 sg13g2_nand2_1 _11800_ (.Y(_03832_),
    .A(_03806_),
    .B(_03812_));
 sg13g2_inv_1 _11801_ (.Y(_03833_),
    .A(_03737_));
 sg13g2_a221oi_1 _11802_ (.B2(_03832_),
    .C1(_03833_),
    .B1(_03831_),
    .A1(_03694_),
    .Y(_03834_),
    .A2(_03734_));
 sg13g2_xnor2_1 _11803_ (.Y(_03835_),
    .A(_03738_),
    .B(_03834_));
 sg13g2_nand3_1 _11804_ (.B(\step[3] ),
    .C(_03924_),
    .A(_03903_),
    .Y(_03836_));
 sg13g2_buf_1 _11805_ (.A(_03836_),
    .X(_03837_));
 sg13g2_or2_1 _11806_ (.X(_03838_),
    .B(_04391_),
    .A(_04280_));
 sg13g2_buf_1 _11807_ (.A(_03838_),
    .X(_03839_));
 sg13g2_nor2_1 _11808_ (.A(_03837_),
    .B(_03839_),
    .Y(_03840_));
 sg13g2_buf_2 _11809_ (.A(_03840_),
    .X(_03841_));
 sg13g2_mux2_1 _11810_ (.A0(_03830_),
    .A1(_03835_),
    .S(_03841_),
    .X(_03842_));
 sg13g2_buf_8 _11811_ (.A(_03842_),
    .X(_03843_));
 sg13g2_inv_4 _11812_ (.A(_03843_),
    .Y(_00029_));
 sg13g2_inv_1 _11813_ (.Y(_03844_),
    .A(\last_iter[0] ));
 sg13g2_a21oi_1 _11814_ (.A1(_03806_),
    .A2(_03812_),
    .Y(_03845_),
    .B1(_03818_));
 sg13g2_or3_1 _11815_ (.A(_03833_),
    .B(_03694_),
    .C(_03845_),
    .X(_03846_));
 sg13g2_nand2_1 _11816_ (.Y(_03847_),
    .A(_03833_),
    .B(_03845_));
 sg13g2_nand3_1 _11817_ (.B(_03694_),
    .C(_03734_),
    .A(_03833_),
    .Y(_03848_));
 sg13g2_or3_1 _11818_ (.A(_03833_),
    .B(_03734_),
    .C(_03845_),
    .X(_03849_));
 sg13g2_nand4_1 _11819_ (.B(_03847_),
    .C(_03848_),
    .A(_03846_),
    .Y(_03850_),
    .D(_03849_));
 sg13g2_mux2_1 _11820_ (.A0(_03844_),
    .A1(_03850_),
    .S(_03841_),
    .X(_03851_));
 sg13g2_buf_2 _11821_ (.A(_03851_),
    .X(_03852_));
 sg13g2_inv_1 _11822_ (.Y(_00030_),
    .A(_03852_));
 sg13g2_nand3_1 _11823_ (.B(_03738_),
    .C(_03819_),
    .A(_03737_),
    .Y(_03853_));
 sg13g2_inv_1 _11824_ (.Y(_03854_),
    .A(\iter[2] ));
 sg13g2_o21ai_1 _11825_ (.B1(_03854_),
    .Y(_03855_),
    .A1(_03736_),
    .A2(_03853_));
 sg13g2_or3_1 _11826_ (.A(_03854_),
    .B(_03736_),
    .C(_03853_),
    .X(_03856_));
 sg13g2_a21oi_1 _11827_ (.A1(_03855_),
    .A2(_03856_),
    .Y(_03857_),
    .B1(_04439_));
 sg13g2_nor2_1 _11828_ (.A(\last_iter[2] ),
    .B(_03841_),
    .Y(_03858_));
 sg13g2_or2_1 _11829_ (.X(_03859_),
    .B(_03858_),
    .A(_03857_));
 sg13g2_buf_2 _11830_ (.A(_03859_),
    .X(_03860_));
 sg13g2_inv_8 _11831_ (.Y(_00031_),
    .A(_03860_));
 sg13g2_buf_1 _11832_ (.A(_00026_),
    .X(_03861_));
 sg13g2_nand3_1 _11833_ (.B(_03861_),
    .C(_04327_),
    .A(_03964_),
    .Y(_03862_));
 sg13g2_a21o_1 _11834_ (.A2(_03862_),
    .A1(_03998_),
    .B1(_04041_),
    .X(_03863_));
 sg13g2_inv_1 _11835_ (.Y(_03864_),
    .A(_04071_));
 sg13g2_nand2_1 _11836_ (.Y(_03865_),
    .A(_04060_),
    .B(_03864_));
 sg13g2_a21oi_1 _11837_ (.A1(net336),
    .A2(_03863_),
    .Y(_03866_),
    .B1(_03865_));
 sg13g2_nand4_1 _11838_ (.B(_04317_),
    .C(_04071_),
    .A(net336),
    .Y(_03867_),
    .D(_03863_));
 sg13g2_nor2b_1 _11839_ (.A(_03866_),
    .B_N(_03867_),
    .Y(_03868_));
 sg13g2_or3_1 _11840_ (.A(_00033_),
    .B(_04298_),
    .C(_03868_),
    .X(_00002_));
 sg13g2_buf_1 _11841_ (.A(ui_in[3]),
    .X(_03869_));
 sg13g2_buf_1 _11842_ (.A(ui_in[2]),
    .X(_03870_));
 sg13g2_buf_1 _11843_ (.A(ui_in[1]),
    .X(_03871_));
 sg13g2_buf_1 _11844_ (.A(ui_in[0]),
    .X(_03872_));
 sg13g2_nor2_1 _11845_ (.A(_03871_),
    .B(_03872_),
    .Y(_03873_));
 sg13g2_and2_1 _11846_ (.A(_03870_),
    .B(_03873_),
    .X(_03874_));
 sg13g2_buf_2 _11847_ (.A(_03874_),
    .X(_03875_));
 sg13g2_nand2_1 _11848_ (.Y(_03876_),
    .A(_03869_),
    .B(_03875_));
 sg13g2_buf_1 _11849_ (.A(\i_coord.l_xip.data_out[0] ),
    .X(_03877_));
 sg13g2_nand2_1 _11850_ (.Y(_03878_),
    .A(_03870_),
    .B(_03873_));
 sg13g2_buf_2 _11851_ (.A(_03878_),
    .X(_03879_));
 sg13g2_nand2_1 _11852_ (.Y(_03880_),
    .A(_03877_),
    .B(_03879_));
 sg13g2_buf_1 _11853_ (.A(\i_coord.demo_update ),
    .X(_03881_));
 sg13g2_inv_1 _11854_ (.Y(_03882_),
    .A(_03881_));
 sg13g2_buf_1 _11855_ (.A(rst_n),
    .X(_03883_));
 sg13g2_nand2_1 _11856_ (.Y(_03884_),
    .A(_03882_),
    .B(_03883_));
 sg13g2_a21oi_1 _11857_ (.A1(_03876_),
    .A2(_03880_),
    .Y(_00047_),
    .B1(_03884_));
 sg13g2_buf_1 _11858_ (.A(_03881_),
    .X(_03885_));
 sg13g2_buf_1 _11859_ (.A(\i_coord.y_inc_row[-13] ),
    .X(_03886_));
 sg13g2_buf_2 _11860_ (.A(\i_coord.y_inc_row[-11] ),
    .X(_03887_));
 sg13g2_buf_1 _11861_ (.A(\i_coord.y_inc_row[-10] ),
    .X(_03888_));
 sg13g2_buf_2 _11862_ (.A(\i_coord.y_inc_row[-8] ),
    .X(_03889_));
 sg13g2_buf_2 _11863_ (.A(\i_coord.y_inc_row[-9] ),
    .X(_03890_));
 sg13g2_buf_1 _11864_ (.A(\i_coord.y_inc_row[-7] ),
    .X(_03891_));
 sg13g2_inv_1 _11865_ (.Y(_03892_),
    .A(_03891_));
 sg13g2_nor4_1 _11866_ (.A(_03888_),
    .B(_03889_),
    .C(_03890_),
    .D(_03892_),
    .Y(_03893_));
 sg13g2_buf_2 _11867_ (.A(\i_coord.y_inc_row[-12] ),
    .X(_03894_));
 sg13g2_buf_1 _11868_ (.A(\i_coord.y_inc_row[-6] ),
    .X(_03895_));
 sg13g2_nor2_1 _11869_ (.A(_03894_),
    .B(net321),
    .Y(_03896_));
 sg13g2_nand4_1 _11870_ (.B(_03887_),
    .C(_03893_),
    .A(net322),
    .Y(_03897_),
    .D(_03896_));
 sg13g2_buf_2 _11871_ (.A(_03897_),
    .X(_03898_));
 sg13g2_and2_1 _11872_ (.A(net274),
    .B(_03898_),
    .X(_03899_));
 sg13g2_buf_2 _11873_ (.A(_03899_),
    .X(_03900_));
 sg13g2_buf_1 _11874_ (.A(_03900_),
    .X(_03901_));
 sg13g2_inv_1 _11875_ (.Y(_03902_),
    .A(net321));
 sg13g2_buf_1 _11876_ (.A(_03902_),
    .X(_03904_));
 sg13g2_inv_1 _11877_ (.Y(_03905_),
    .A(_03888_));
 sg13g2_nand3_1 _11878_ (.B(net322),
    .C(_03887_),
    .A(_03894_),
    .Y(_03906_));
 sg13g2_nor2_1 _11879_ (.A(_03905_),
    .B(_03906_),
    .Y(_03907_));
 sg13g2_nand3_1 _11880_ (.B(_03890_),
    .C(_03907_),
    .A(_03889_),
    .Y(_03908_));
 sg13g2_buf_1 _11881_ (.A(_03908_),
    .X(_03909_));
 sg13g2_or2_1 _11882_ (.X(_03910_),
    .B(_03909_),
    .A(_03892_));
 sg13g2_xnor2_1 _11883_ (.Y(_03911_),
    .A(net226),
    .B(_03910_));
 sg13g2_buf_2 _11884_ (.A(_03911_),
    .X(_03912_));
 sg13g2_xor2_1 _11885_ (.B(_03912_),
    .A(net322),
    .X(_03913_));
 sg13g2_inv_1 _11886_ (.Y(_03915_),
    .A(net1));
 sg13g2_a21oi_1 _11887_ (.A1(_03915_),
    .A2(_03875_),
    .Y(_03916_),
    .B1(net274));
 sg13g2_a21oi_1 _11888_ (.A1(_03901_),
    .A2(_03913_),
    .Y(_03917_),
    .B1(_03916_));
 sg13g2_buf_1 _11889_ (.A(net274),
    .X(_03918_));
 sg13g2_buf_1 _11890_ (.A(\i_coord.l_xip.data_out[1] ),
    .X(_03919_));
 sg13g2_nor3_1 _11891_ (.A(net225),
    .B(_03919_),
    .C(_03875_),
    .Y(_03920_));
 sg13g2_buf_1 _11892_ (.A(_03883_),
    .X(_03921_));
 sg13g2_buf_1 _11893_ (.A(net320),
    .X(_03922_));
 sg13g2_buf_1 _11894_ (.A(net273),
    .X(_03923_));
 sg13g2_o21ai_1 _11895_ (.B1(net224),
    .Y(_00048_),
    .A1(_03917_),
    .A2(_03920_));
 sg13g2_inv_1 _11896_ (.Y(_03925_),
    .A(_03883_));
 sg13g2_buf_1 _11897_ (.A(_03925_),
    .X(_03926_));
 sg13g2_buf_1 _11898_ (.A(ui_in[5]),
    .X(_03927_));
 sg13g2_mux2_1 _11899_ (.A0(_03927_),
    .A1(\i_coord.l_xip.data_out[2] ),
    .S(_03879_),
    .X(_03928_));
 sg13g2_nor2_1 _11900_ (.A(net225),
    .B(_03928_),
    .Y(_03929_));
 sg13g2_buf_1 _11901_ (.A(_03882_),
    .X(_03930_));
 sg13g2_nand2_2 _11902_ (.Y(_03931_),
    .A(_03898_),
    .B(_03912_));
 sg13g2_xnor2_1 _11903_ (.Y(_03932_),
    .A(_03894_),
    .B(net322));
 sg13g2_xnor2_1 _11904_ (.Y(_03933_),
    .A(_03931_),
    .B(_03932_));
 sg13g2_nor2_1 _11905_ (.A(_03930_),
    .B(_03933_),
    .Y(_03934_));
 sg13g2_nor3_1 _11906_ (.A(net272),
    .B(_03929_),
    .C(_03934_),
    .Y(_00049_));
 sg13g2_buf_1 _11907_ (.A(_03882_),
    .X(_03936_));
 sg13g2_nand2_1 _11908_ (.Y(_03937_),
    .A(_03894_),
    .B(net322));
 sg13g2_xor2_1 _11909_ (.B(_03937_),
    .A(_03887_),
    .X(_03938_));
 sg13g2_inv_1 _11910_ (.Y(_03939_),
    .A(_03938_));
 sg13g2_xnor2_1 _11911_ (.Y(_03940_),
    .A(_03912_),
    .B(_03939_));
 sg13g2_nor2_1 _11912_ (.A(net222),
    .B(_03940_),
    .Y(_03941_));
 sg13g2_buf_1 _11913_ (.A(ui_in[6]),
    .X(_03942_));
 sg13g2_mux2_1 _11914_ (.A0(_03942_),
    .A1(\i_coord.l_xip.data_out[3] ),
    .S(_03879_),
    .X(_03943_));
 sg13g2_nor2_1 _11915_ (.A(net225),
    .B(_03943_),
    .Y(_03944_));
 sg13g2_o21ai_1 _11916_ (.B1(net224),
    .Y(_00050_),
    .A1(_03941_),
    .A2(_03944_));
 sg13g2_xnor2_1 _11917_ (.Y(_03946_),
    .A(_03905_),
    .B(_03906_));
 sg13g2_a21oi_1 _11918_ (.A1(_03898_),
    .A2(_03946_),
    .Y(_03947_),
    .B1(_03882_));
 sg13g2_and2_1 _11919_ (.A(_03875_),
    .B(_03947_),
    .X(_03948_));
 sg13g2_xnor2_1 _11920_ (.Y(_03949_),
    .A(_03931_),
    .B(_03947_));
 sg13g2_buf_1 _11921_ (.A(net274),
    .X(_03950_));
 sg13g2_buf_1 _11922_ (.A(ui_in[7]),
    .X(_03951_));
 sg13g2_mux2_1 _11923_ (.A0(_03951_),
    .A1(\i_coord.l_xip.data_out[4] ),
    .S(_03879_),
    .X(_03952_));
 sg13g2_o21ai_1 _11924_ (.B1(net273),
    .Y(_03953_),
    .A1(_03918_),
    .A2(_03952_));
 sg13g2_a221oi_1 _11925_ (.B2(net221),
    .C1(_03953_),
    .B1(_03949_),
    .A1(_03931_),
    .Y(_00051_),
    .A2(_03948_));
 sg13g2_xnor2_1 _11926_ (.Y(_03955_),
    .A(_03890_),
    .B(_03907_));
 sg13g2_xor2_1 _11927_ (.B(_03955_),
    .A(_03912_),
    .X(_03956_));
 sg13g2_nand2_1 _11928_ (.Y(_03957_),
    .A(net221),
    .B(_03956_));
 sg13g2_buf_1 _11929_ (.A(uio_in[0]),
    .X(_03958_));
 sg13g2_mux2_1 _11930_ (.A0(_03958_),
    .A1(\i_coord.l_xip.data_out[5] ),
    .S(_03879_),
    .X(_03959_));
 sg13g2_nand2_1 _11931_ (.Y(_03960_),
    .A(net223),
    .B(_03959_));
 sg13g2_buf_1 _11932_ (.A(net272),
    .X(_03961_));
 sg13g2_a21oi_1 _11933_ (.A1(_03957_),
    .A2(_03960_),
    .Y(_00052_),
    .B1(net220));
 sg13g2_nand2_1 _11934_ (.Y(_03962_),
    .A(_03890_),
    .B(_03907_));
 sg13g2_xor2_1 _11935_ (.B(_03962_),
    .A(_03889_),
    .X(_03963_));
 sg13g2_xor2_1 _11936_ (.B(_03963_),
    .A(_03912_),
    .X(_03965_));
 sg13g2_inv_1 _11937_ (.Y(_03966_),
    .A(net2));
 sg13g2_a21oi_1 _11938_ (.A1(_03966_),
    .A2(_03875_),
    .Y(_03967_),
    .B1(net274));
 sg13g2_a21oi_1 _11939_ (.A1(net89),
    .A2(_03965_),
    .Y(_03968_),
    .B1(_03967_));
 sg13g2_nor3_1 _11940_ (.A(_03918_),
    .B(\i_coord.l_xip.data_out[6] ),
    .C(_03875_),
    .Y(_03969_));
 sg13g2_nor3_1 _11941_ (.A(net272),
    .B(_03968_),
    .C(_03969_),
    .Y(_00053_));
 sg13g2_buf_1 _11942_ (.A(uio_in[2]),
    .X(_03970_));
 sg13g2_mux2_1 _11943_ (.A0(_03970_),
    .A1(\i_coord.l_xip.data_out[7] ),
    .S(_03879_),
    .X(_03971_));
 sg13g2_nand2_1 _11944_ (.Y(_03972_),
    .A(net223),
    .B(_03971_));
 sg13g2_a21o_1 _11945_ (.A2(_03909_),
    .A1(_03892_),
    .B1(_03904_),
    .X(_03973_));
 sg13g2_nand3_1 _11946_ (.B(_03904_),
    .C(_03909_),
    .A(_03892_),
    .Y(_03975_));
 sg13g2_nand3_1 _11947_ (.B(_03973_),
    .C(_03975_),
    .A(net221),
    .Y(_03976_));
 sg13g2_nand3_1 _11948_ (.B(_03972_),
    .C(_03976_),
    .A(net273),
    .Y(_00054_));
 sg13g2_buf_1 _11949_ (.A(uio_in[3]),
    .X(_03977_));
 sg13g2_nand2_1 _11950_ (.Y(_03978_),
    .A(_03977_),
    .B(_03875_));
 sg13g2_nand2_1 _11951_ (.Y(_03979_),
    .A(\i_coord.l_xip.data_out[8] ),
    .B(_03879_));
 sg13g2_a21oi_1 _11952_ (.A1(_03978_),
    .A2(_03979_),
    .Y(_00055_),
    .B1(_03884_));
 sg13g2_buf_1 _11953_ (.A(uio_in[4]),
    .X(_03980_));
 sg13g2_nand2_1 _11954_ (.Y(_03981_),
    .A(_03980_),
    .B(_03875_));
 sg13g2_buf_1 _11955_ (.A(\i_coord.l_xip.data_out[9] ),
    .X(_03982_));
 sg13g2_nand2_1 _11956_ (.Y(_03984_),
    .A(_03982_),
    .B(_03879_));
 sg13g2_a21oi_1 _11957_ (.A1(_03981_),
    .A2(_03984_),
    .Y(_00056_),
    .B1(_03884_));
 sg13g2_buf_1 _11958_ (.A(\i_coord.l_xir.data_out[0] ),
    .X(_03985_));
 sg13g2_and2_1 _11959_ (.A(net273),
    .B(_03869_),
    .X(_03986_));
 sg13g2_inv_1 _11960_ (.Y(_03987_),
    .A(_03870_));
 sg13g2_nand2b_1 _11961_ (.Y(_03988_),
    .B(_03871_),
    .A_N(_03872_));
 sg13g2_o21ai_1 _11962_ (.B1(net320),
    .Y(_03989_),
    .A1(_03987_),
    .A2(_03988_));
 sg13g2_buf_4 _11963_ (.X(_03990_),
    .A(_03989_));
 sg13g2_mux2_1 _11964_ (.A0(_03985_),
    .A1(_03986_),
    .S(_03990_),
    .X(_00057_));
 sg13g2_nor2_1 _11965_ (.A(net272),
    .B(_03915_),
    .Y(_03991_));
 sg13g2_mux2_1 _11966_ (.A0(\i_coord.l_xir.data_out[1] ),
    .A1(_03991_),
    .S(_03990_),
    .X(_00058_));
 sg13g2_and2_1 _11967_ (.A(net273),
    .B(_03927_),
    .X(_03993_));
 sg13g2_mux2_1 _11968_ (.A0(\i_coord.l_xir.data_out[2] ),
    .A1(_03993_),
    .S(_03990_),
    .X(_00059_));
 sg13g2_and2_1 _11969_ (.A(_03922_),
    .B(_03942_),
    .X(_03994_));
 sg13g2_mux2_1 _11970_ (.A0(\i_coord.l_xir.data_out[3] ),
    .A1(_03994_),
    .S(_03990_),
    .X(_00060_));
 sg13g2_and2_1 _11971_ (.A(_03922_),
    .B(_03951_),
    .X(_03995_));
 sg13g2_mux2_1 _11972_ (.A0(\i_coord.l_xir.data_out[4] ),
    .A1(_03995_),
    .S(_03990_),
    .X(_00061_));
 sg13g2_and2_1 _11973_ (.A(net320),
    .B(_03958_),
    .X(_03996_));
 sg13g2_mux2_1 _11974_ (.A0(\i_coord.l_xir.data_out[5] ),
    .A1(_03996_),
    .S(_03990_),
    .X(_00062_));
 sg13g2_nor2_1 _11975_ (.A(net272),
    .B(_03966_),
    .Y(_03997_));
 sg13g2_mux2_1 _11976_ (.A0(\i_coord.l_xir.data_out[6] ),
    .A1(_03997_),
    .S(_03990_),
    .X(_00063_));
 sg13g2_buf_1 _11977_ (.A(\i_coord.l_xir.data_out[7] ),
    .X(_03999_));
 sg13g2_and2_1 _11978_ (.A(net320),
    .B(_03970_),
    .X(_04000_));
 sg13g2_mux2_1 _11979_ (.A0(_03999_),
    .A1(_04000_),
    .S(_03990_),
    .X(_00064_));
 sg13g2_nand2b_1 _11980_ (.Y(_04001_),
    .B(_03872_),
    .A_N(_03871_));
 sg13g2_nor2_1 _11981_ (.A(_03870_),
    .B(_04001_),
    .Y(_04002_));
 sg13g2_nor2_1 _11982_ (.A(_03926_),
    .B(_04002_),
    .Y(_04003_));
 sg13g2_buf_1 _11983_ (.A(_04003_),
    .X(_04004_));
 sg13g2_nand2_1 _11984_ (.Y(_04005_),
    .A(_03987_),
    .B(net320));
 sg13g2_nor2_1 _11985_ (.A(_04001_),
    .B(_04005_),
    .Y(_04006_));
 sg13g2_buf_1 _11986_ (.A(_04006_),
    .X(_04008_));
 sg13g2_buf_1 _11987_ (.A(_04008_),
    .X(_04009_));
 sg13g2_a22oi_1 _11988_ (.Y(_04010_),
    .B1(_04009_),
    .B2(_03970_),
    .A2(_04004_),
    .A1(\i_coord.l_xl.data_out[10] ));
 sg13g2_inv_1 _11989_ (.Y(_00065_),
    .A(_04010_));
 sg13g2_a22oi_1 _11990_ (.Y(_04011_),
    .B1(net142),
    .B2(_03977_),
    .A2(net168),
    .A1(\i_coord.l_xl.data_out[11] ));
 sg13g2_inv_1 _11991_ (.Y(_00066_),
    .A(_04011_));
 sg13g2_a22oi_1 _11992_ (.Y(_04012_),
    .B1(_04009_),
    .B2(_03980_),
    .A2(_04004_),
    .A1(\i_coord.l_xl.data_out[12] ));
 sg13g2_inv_1 _11993_ (.Y(_00067_),
    .A(_04012_));
 sg13g2_a22oi_1 _11994_ (.Y(_04013_),
    .B1(net142),
    .B2(net3),
    .A2(net168),
    .A1(\i_coord.l_xl.data_out[13] ));
 sg13g2_inv_1 _11995_ (.Y(_00068_),
    .A(_04013_));
 sg13g2_inv_1 _11996_ (.Y(_04015_),
    .A(\i_coord.l_xl.data_out[14] ));
 sg13g2_inv_1 _11997_ (.Y(_04016_),
    .A(net4));
 sg13g2_a22oi_1 _11998_ (.Y(_00069_),
    .B1(net142),
    .B2(_04016_),
    .A2(net168),
    .A1(_04015_));
 sg13g2_inv_1 _11999_ (.Y(_04017_),
    .A(\i_coord.l_xl.data_out[15] ));
 sg13g2_inv_1 _12000_ (.Y(_04018_),
    .A(net5));
 sg13g2_a22oi_1 _12001_ (.Y(_00070_),
    .B1(net142),
    .B2(_04018_),
    .A2(net168),
    .A1(_04017_));
 sg13g2_a22oi_1 _12002_ (.Y(_04019_),
    .B1(net142),
    .B2(_03869_),
    .A2(net168),
    .A1(\i_coord.l_xl.data_out[3] ));
 sg13g2_inv_1 _12003_ (.Y(_00071_),
    .A(_04019_));
 sg13g2_a22oi_1 _12004_ (.Y(_04020_),
    .B1(net142),
    .B2(net1),
    .A2(net168),
    .A1(\i_coord.l_xl.data_out[4] ));
 sg13g2_inv_1 _12005_ (.Y(_00072_),
    .A(_04020_));
 sg13g2_a22oi_1 _12006_ (.Y(_04022_),
    .B1(net142),
    .B2(_03927_),
    .A2(net168),
    .A1(\i_coord.l_xl.data_out[5] ));
 sg13g2_inv_1 _12007_ (.Y(_00073_),
    .A(_04022_));
 sg13g2_a22oi_1 _12008_ (.Y(_04023_),
    .B1(net142),
    .B2(_03942_),
    .A2(net168),
    .A1(\i_coord.l_xl.data_out[6] ));
 sg13g2_inv_1 _12009_ (.Y(_00074_),
    .A(_04023_));
 sg13g2_a22oi_1 _12010_ (.Y(_04024_),
    .B1(_04008_),
    .B2(_03951_),
    .A2(_04003_),
    .A1(\i_coord.l_xl.data_out[7] ));
 sg13g2_inv_1 _12011_ (.Y(_00075_),
    .A(_04024_));
 sg13g2_a22oi_1 _12012_ (.Y(_04025_),
    .B1(_04008_),
    .B2(_03958_),
    .A2(_04003_),
    .A1(\i_coord.l_xl.data_out[8] ));
 sg13g2_inv_1 _12013_ (.Y(_00076_),
    .A(_04025_));
 sg13g2_a22oi_1 _12014_ (.Y(_04026_),
    .B1(_04008_),
    .B2(net2),
    .A2(_04003_),
    .A1(\i_coord.l_xl.data_out[9] ));
 sg13g2_inv_1 _12015_ (.Y(_00077_),
    .A(_04026_));
 sg13g2_buf_1 _12016_ (.A(\i_coord.l_yip.data_out[0] ),
    .X(_04028_));
 sg13g2_o21ai_1 _12017_ (.B1(_03921_),
    .Y(_04029_),
    .A1(_03987_),
    .A2(_04001_));
 sg13g2_buf_1 _12018_ (.A(_04029_),
    .X(_04030_));
 sg13g2_buf_1 _12019_ (.A(_04030_),
    .X(_04031_));
 sg13g2_mux2_1 _12020_ (.A0(_04028_),
    .A1(_03986_),
    .S(net167),
    .X(_00078_));
 sg13g2_buf_1 _12021_ (.A(\i_coord.l_yip.data_out[1] ),
    .X(_04032_));
 sg13g2_mux2_1 _12022_ (.A0(_04032_),
    .A1(_03991_),
    .S(_04031_),
    .X(_00079_));
 sg13g2_buf_1 _12023_ (.A(\i_coord.l_yip.data_out[2] ),
    .X(_04033_));
 sg13g2_mux2_1 _12024_ (.A0(_04033_),
    .A1(_03993_),
    .S(net167),
    .X(_00080_));
 sg13g2_mux2_1 _12025_ (.A0(\i_coord.l_yip.data_out[3] ),
    .A1(_03994_),
    .S(net167),
    .X(_00081_));
 sg13g2_buf_1 _12026_ (.A(\i_coord.l_yip.data_out[4] ),
    .X(_04035_));
 sg13g2_mux2_1 _12027_ (.A0(_04035_),
    .A1(_03995_),
    .S(net167),
    .X(_00082_));
 sg13g2_buf_1 _12028_ (.A(\i_coord.l_yip.data_out[5] ),
    .X(_04036_));
 sg13g2_mux2_1 _12029_ (.A0(_04036_),
    .A1(_03996_),
    .S(_04031_),
    .X(_00083_));
 sg13g2_mux2_1 _12030_ (.A0(\i_coord.l_yip.data_out[6] ),
    .A1(_03997_),
    .S(net167),
    .X(_00084_));
 sg13g2_buf_1 _12031_ (.A(\i_coord.l_yip.data_out[7] ),
    .X(_04037_));
 sg13g2_mux2_1 _12032_ (.A0(_04037_),
    .A1(_04000_),
    .S(net167),
    .X(_00085_));
 sg13g2_buf_1 _12033_ (.A(\i_coord.l_yip.data_out[8] ),
    .X(_04038_));
 sg13g2_inv_1 _12034_ (.Y(_04039_),
    .A(_04038_));
 sg13g2_nand3_1 _12035_ (.B(_03977_),
    .C(_04030_),
    .A(net273),
    .Y(_04040_));
 sg13g2_o21ai_1 _12036_ (.B1(_04040_),
    .Y(_00086_),
    .A1(_04039_),
    .A2(net167));
 sg13g2_buf_1 _12037_ (.A(\i_coord.l_yip.data_out[9] ),
    .X(_04042_));
 sg13g2_inv_1 _12038_ (.Y(_04043_),
    .A(_04042_));
 sg13g2_nand3_1 _12039_ (.B(_03980_),
    .C(_04030_),
    .A(net273),
    .Y(_04044_));
 sg13g2_o21ai_1 _12040_ (.B1(_04044_),
    .Y(_00087_),
    .A1(_04043_),
    .A2(net167));
 sg13g2_nand3b_1 _12041_ (.B(_03898_),
    .C(net320),
    .Y(_04045_),
    .A_N(_00014_));
 sg13g2_buf_2 _12042_ (.A(\i_coord.y0[-13] ),
    .X(_04046_));
 sg13g2_nor2_1 _12043_ (.A(_03870_),
    .B(_03988_),
    .Y(_04047_));
 sg13g2_nor2_1 _12044_ (.A(_03881_),
    .B(_03925_),
    .Y(_04048_));
 sg13g2_nand2b_1 _12045_ (.Y(_04049_),
    .B(_04048_),
    .A_N(_04047_));
 sg13g2_buf_1 _12046_ (.A(_04049_),
    .X(_04051_));
 sg13g2_nand2_1 _12047_ (.Y(_04052_),
    .A(_04046_),
    .B(_04051_));
 sg13g2_nor2_1 _12048_ (.A(_03884_),
    .B(_04047_),
    .Y(_04053_));
 sg13g2_buf_2 _12049_ (.A(_04053_),
    .X(_04054_));
 sg13g2_buf_1 _12050_ (.A(_04054_),
    .X(_04055_));
 sg13g2_nand2_1 _12051_ (.Y(_04056_),
    .A(\i_coord.l_yt.data_out[0] ),
    .B(_04055_));
 sg13g2_o21ai_1 _12052_ (.B1(_04056_),
    .Y(_00088_),
    .A1(_04045_),
    .A2(_04052_));
 sg13g2_buf_1 _12053_ (.A(\i_coord.y0[-5] ),
    .X(_04057_));
 sg13g2_buf_2 _12054_ (.A(\i_coord.y0[-4] ),
    .X(_04058_));
 sg13g2_buf_1 _12055_ (.A(\i_coord.y0[-6] ),
    .X(_04059_));
 sg13g2_inv_1 _12056_ (.Y(_04061_),
    .A(_04059_));
 sg13g2_buf_1 _12057_ (.A(\i_coord.y0[-8] ),
    .X(_04062_));
 sg13g2_buf_2 _12058_ (.A(\i_coord.y0[-9] ),
    .X(_04063_));
 sg13g2_buf_1 _12059_ (.A(\i_coord.y0[-7] ),
    .X(_04064_));
 sg13g2_nand3_1 _12060_ (.B(_04063_),
    .C(_04064_),
    .A(net317),
    .Y(_04065_));
 sg13g2_nor2_2 _12061_ (.A(_04061_),
    .B(_04065_),
    .Y(_04066_));
 sg13g2_or3_1 _12062_ (.A(_04057_),
    .B(_04058_),
    .C(_04066_),
    .X(_04067_));
 sg13g2_buf_1 _12063_ (.A(_04067_),
    .X(_04068_));
 sg13g2_xor2_1 _12064_ (.B(_04068_),
    .A(_00022_),
    .X(_04069_));
 sg13g2_a22oi_1 _12065_ (.Y(_04070_),
    .B1(net89),
    .B2(_04069_),
    .A2(_03977_),
    .A1(net222));
 sg13g2_nand2_1 _12066_ (.Y(_04072_),
    .A(_03921_),
    .B(_04051_));
 sg13g2_buf_2 _12067_ (.A(_04072_),
    .X(_04073_));
 sg13g2_nand2_1 _12068_ (.Y(_04074_),
    .A(\i_coord.l_yt.data_out[10] ),
    .B(net119));
 sg13g2_o21ai_1 _12069_ (.B1(_04074_),
    .Y(_00089_),
    .A1(_04070_),
    .A2(_04073_));
 sg13g2_inv_1 _12070_ (.Y(_04075_),
    .A(\i_coord.l_yt.data_out[11] ));
 sg13g2_buf_2 _12071_ (.A(\i_coord.y0[-3] ),
    .X(_04076_));
 sg13g2_nor2_1 _12072_ (.A(_04076_),
    .B(_04068_),
    .Y(_04077_));
 sg13g2_xnor2_1 _12073_ (.Y(_04078_),
    .A(_00023_),
    .B(_04077_));
 sg13g2_and2_1 _12074_ (.A(net320),
    .B(_03900_),
    .X(_04079_));
 sg13g2_a221oi_1 _12075_ (.B2(_04079_),
    .C1(_04054_),
    .B1(_04078_),
    .A1(_03980_),
    .Y(_04080_),
    .A2(_04048_));
 sg13g2_a21oi_1 _12076_ (.A1(_04075_),
    .A2(net119),
    .Y(_00090_),
    .B1(_04080_));
 sg13g2_inv_1 _12077_ (.Y(_04082_),
    .A(_00024_));
 sg13g2_buf_2 _12078_ (.A(\i_coord.y0[-2] ),
    .X(_04083_));
 sg13g2_nor2_1 _12079_ (.A(_04076_),
    .B(_04083_),
    .Y(_04084_));
 sg13g2_nand2b_1 _12080_ (.Y(_04085_),
    .B(_04084_),
    .A_N(_04068_));
 sg13g2_xnor2_1 _12081_ (.Y(_04086_),
    .A(_04082_),
    .B(_04085_));
 sg13g2_a22oi_1 _12082_ (.Y(_04087_),
    .B1(net89),
    .B2(_04086_),
    .A2(net3),
    .A1(net222));
 sg13g2_nand2_1 _12083_ (.Y(_04088_),
    .A(\i_coord.l_yt.data_out[12] ),
    .B(net119));
 sg13g2_o21ai_1 _12084_ (.B1(_04088_),
    .Y(_00091_),
    .A1(_04073_),
    .A2(_04087_));
 sg13g2_inv_1 _12085_ (.Y(_04089_),
    .A(\i_coord.l_yt.data_out[13] ));
 sg13g2_buf_2 _12086_ (.A(\i_coord.y0[-1] ),
    .X(_04091_));
 sg13g2_nor2_1 _12087_ (.A(_04091_),
    .B(_04085_),
    .Y(_04092_));
 sg13g2_xnor2_1 _12088_ (.Y(_04093_),
    .A(_00025_),
    .B(_04092_));
 sg13g2_a221oi_1 _12089_ (.B2(_04093_),
    .C1(_04054_),
    .B1(_04079_),
    .A1(net4),
    .Y(_04094_),
    .A2(_04048_));
 sg13g2_a21oi_1 _12090_ (.A1(_04089_),
    .A2(net119),
    .Y(_00092_),
    .B1(_04094_));
 sg13g2_inv_1 _12091_ (.Y(_04095_),
    .A(\i_coord.l_yt.data_out[14] ));
 sg13g2_nor2_2 _12092_ (.A(net272),
    .B(_04054_),
    .Y(_04096_));
 sg13g2_buf_2 _12093_ (.A(\i_coord.y0[1] ),
    .X(_04097_));
 sg13g2_buf_1 _12094_ (.A(\i_coord.y0[0] ),
    .X(_04098_));
 sg13g2_nor2_1 _12095_ (.A(_04091_),
    .B(_04098_),
    .Y(_04099_));
 sg13g2_nor2b_1 _12096_ (.A(_04085_),
    .B_N(_04099_),
    .Y(_04101_));
 sg13g2_xnor2_1 _12097_ (.Y(_04102_),
    .A(_04097_),
    .B(_04101_));
 sg13g2_nand2_1 _12098_ (.Y(_04103_),
    .A(_03900_),
    .B(_04102_));
 sg13g2_o21ai_1 _12099_ (.B1(_04103_),
    .Y(_04104_),
    .A1(net225),
    .A2(net5));
 sg13g2_a22oi_1 _12100_ (.Y(_00093_),
    .B1(_04096_),
    .B2(_04104_),
    .A2(net119),
    .A1(_04095_));
 sg13g2_buf_2 _12101_ (.A(\i_coord.y0[-12] ),
    .X(_04105_));
 sg13g2_nand2_1 _12102_ (.Y(_04106_),
    .A(_04105_),
    .B(_04051_));
 sg13g2_nand2_1 _12103_ (.Y(_04107_),
    .A(\i_coord.l_yt.data_out[1] ),
    .B(_04055_));
 sg13g2_o21ai_1 _12104_ (.B1(_04107_),
    .Y(_00094_),
    .A1(_04045_),
    .A2(_04106_));
 sg13g2_buf_2 _12105_ (.A(\i_coord.y0[-11] ),
    .X(_04108_));
 sg13g2_a22oi_1 _12106_ (.Y(_04110_),
    .B1(_04108_),
    .B2(net89),
    .A2(_03869_),
    .A1(net222));
 sg13g2_nand2_1 _12107_ (.Y(_04111_),
    .A(\i_coord.l_yt.data_out[2] ),
    .B(_04054_));
 sg13g2_o21ai_1 _12108_ (.B1(_04111_),
    .Y(_00095_),
    .A1(_04073_),
    .A2(_04110_));
 sg13g2_buf_2 _12109_ (.A(\i_coord.y0[-10] ),
    .X(_04112_));
 sg13g2_a22oi_1 _12110_ (.Y(_04113_),
    .B1(_04112_),
    .B2(net89),
    .A2(net1),
    .A1(net222));
 sg13g2_nand2_1 _12111_ (.Y(_04114_),
    .A(\i_coord.l_yt.data_out[3] ),
    .B(_04054_));
 sg13g2_o21ai_1 _12112_ (.B1(_04114_),
    .Y(_00096_),
    .A1(_04073_),
    .A2(_04113_));
 sg13g2_inv_1 _12113_ (.Y(_04115_),
    .A(\i_coord.l_yt.data_out[4] ));
 sg13g2_nand2b_1 _12114_ (.Y(_04116_),
    .B(_03900_),
    .A_N(_00018_));
 sg13g2_o21ai_1 _12115_ (.B1(_04116_),
    .Y(_04117_),
    .A1(net225),
    .A2(_03927_));
 sg13g2_a22oi_1 _12116_ (.Y(_00097_),
    .B1(_04096_),
    .B2(_04117_),
    .A2(net119),
    .A1(_04115_));
 sg13g2_inv_1 _12117_ (.Y(_04119_),
    .A(\i_coord.l_yt.data_out[5] ));
 sg13g2_xnor2_1 _12118_ (.Y(_04120_),
    .A(net317),
    .B(_04063_));
 sg13g2_nand3_1 _12119_ (.B(_03898_),
    .C(_04120_),
    .A(net274),
    .Y(_04121_));
 sg13g2_o21ai_1 _12120_ (.B1(_04121_),
    .Y(_04122_),
    .A1(net225),
    .A2(_03942_));
 sg13g2_a22oi_1 _12121_ (.Y(_00098_),
    .B1(_04096_),
    .B2(_04122_),
    .A2(net119),
    .A1(_04119_));
 sg13g2_inv_1 _12122_ (.Y(_04123_),
    .A(\i_coord.l_yt.data_out[6] ));
 sg13g2_nand2_1 _12123_ (.Y(_04124_),
    .A(_03936_),
    .B(_03951_));
 sg13g2_nand2_1 _12124_ (.Y(_04125_),
    .A(net317),
    .B(_04063_));
 sg13g2_xor2_1 _12125_ (.B(_04125_),
    .A(_00019_),
    .X(_04126_));
 sg13g2_nand3_1 _12126_ (.B(_03898_),
    .C(_04126_),
    .A(net274),
    .Y(_04128_));
 sg13g2_a21o_1 _12127_ (.A2(_04128_),
    .A1(_04124_),
    .B1(_04073_),
    .X(_04129_));
 sg13g2_o21ai_1 _12128_ (.B1(_04129_),
    .Y(_00099_),
    .A1(_04123_),
    .A2(_04051_));
 sg13g2_inv_1 _12129_ (.Y(_04130_),
    .A(\i_coord.l_yt.data_out[7] ));
 sg13g2_and2_1 _12130_ (.A(_04061_),
    .B(_04065_),
    .X(_04131_));
 sg13g2_o21ai_1 _12131_ (.B1(_03900_),
    .Y(_04132_),
    .A1(_04066_),
    .A2(_04131_));
 sg13g2_o21ai_1 _12132_ (.B1(_04132_),
    .Y(_04133_),
    .A1(net225),
    .A2(_03958_));
 sg13g2_a22oi_1 _12133_ (.Y(_00100_),
    .B1(_04096_),
    .B2(_04133_),
    .A2(net119),
    .A1(_04130_));
 sg13g2_xnor2_1 _12134_ (.Y(_04134_),
    .A(_04057_),
    .B(_04066_));
 sg13g2_a22oi_1 _12135_ (.Y(_04135_),
    .B1(net89),
    .B2(_04134_),
    .A2(net2),
    .A1(net222));
 sg13g2_nand2_1 _12136_ (.Y(_04137_),
    .A(\i_coord.l_yt.data_out[8] ),
    .B(_04054_));
 sg13g2_o21ai_1 _12137_ (.B1(_04137_),
    .Y(_00101_),
    .A1(_04073_),
    .A2(_04135_));
 sg13g2_inv_1 _12138_ (.Y(_04138_),
    .A(_04057_));
 sg13g2_inv_1 _12139_ (.Y(_04139_),
    .A(_00021_));
 sg13g2_a21oi_1 _12140_ (.A1(_04138_),
    .A2(_04066_),
    .Y(_04140_),
    .B1(_04139_));
 sg13g2_xnor2_1 _12141_ (.Y(_04141_),
    .A(_00020_),
    .B(_04140_));
 sg13g2_a22oi_1 _12142_ (.Y(_04142_),
    .B1(net89),
    .B2(_04141_),
    .A2(_03970_),
    .A1(net222));
 sg13g2_nand2_1 _12143_ (.Y(_04143_),
    .A(\i_coord.l_yt.data_out[9] ),
    .B(_04054_));
 sg13g2_o21ai_1 _12144_ (.B1(_04143_),
    .Y(_00102_),
    .A1(_04073_),
    .A2(_04142_));
 sg13g2_buf_1 _12145_ (.A(_04280_),
    .X(_04144_));
 sg13g2_buf_1 _12146_ (.A(net77),
    .X(_04146_));
 sg13g2_buf_1 _12147_ (.A(\i_coord.x_row_start[-13] ),
    .X(_04147_));
 sg13g2_nand4_1 _12148_ (.B(_03964_),
    .C(_04021_),
    .A(_04359_),
    .Y(_04148_),
    .D(_04071_));
 sg13g2_nor4_1 _12149_ (.A(_04007_),
    .B(_04298_),
    .C(_04348_),
    .D(_04148_),
    .Y(_04149_));
 sg13g2_buf_1 _12150_ (.A(_04149_),
    .X(_04150_));
 sg13g2_buf_1 _12151_ (.A(_04150_),
    .X(_04151_));
 sg13g2_nand2_1 _12152_ (.Y(_04152_),
    .A(_03985_),
    .B(net104));
 sg13g2_xor2_1 _12153_ (.B(_04152_),
    .A(_04147_),
    .X(_04153_));
 sg13g2_nor2_1 _12154_ (.A(net66),
    .B(_04153_),
    .Y(_00103_));
 sg13g2_nor4_1 _12155_ (.A(_04298_),
    .B(_04308_),
    .C(_04348_),
    .D(_04381_),
    .Y(_04154_));
 sg13g2_buf_2 _12156_ (.A(_04154_),
    .X(_04156_));
 sg13g2_nor2_1 _12157_ (.A(_04280_),
    .B(_04156_),
    .Y(_04157_));
 sg13g2_buf_2 _12158_ (.A(_04157_),
    .X(_04158_));
 sg13g2_buf_1 _12159_ (.A(_04158_),
    .X(_04159_));
 sg13g2_buf_1 _12160_ (.A(net59),
    .X(_04160_));
 sg13g2_buf_1 _12161_ (.A(net49),
    .X(_04161_));
 sg13g2_or4_1 _12162_ (.A(_04298_),
    .B(_04308_),
    .C(_04348_),
    .D(_04381_),
    .X(_04162_));
 sg13g2_buf_1 _12163_ (.A(_04162_),
    .X(_04163_));
 sg13g2_buf_1 _12164_ (.A(_04163_),
    .X(_04164_));
 sg13g2_inv_2 _12165_ (.Y(_04165_),
    .A(net318));
 sg13g2_buf_2 _12166_ (.A(\i_coord.x_row_start[-4] ),
    .X(_04167_));
 sg13g2_buf_1 _12167_ (.A(\i_coord.x_row_start[-6] ),
    .X(_04168_));
 sg13g2_buf_1 _12168_ (.A(\i_coord.x_row_start[-7] ),
    .X(_04169_));
 sg13g2_inv_1 _12169_ (.Y(_04170_),
    .A(_04169_));
 sg13g2_buf_1 _12170_ (.A(\i_coord.x_row_start[-8] ),
    .X(_04171_));
 sg13g2_buf_1 _12171_ (.A(\i_coord.x_row_start[-9] ),
    .X(_04172_));
 sg13g2_inv_1 _12172_ (.Y(_04173_),
    .A(_04172_));
 sg13g2_buf_1 _12173_ (.A(\i_coord.x_row_start[-10] ),
    .X(_04174_));
 sg13g2_buf_1 _12174_ (.A(\i_coord.x_row_start[-11] ),
    .X(_04175_));
 sg13g2_inv_1 _12175_ (.Y(_04176_),
    .A(\i_coord.l_xir.data_out[1] ));
 sg13g2_buf_1 _12176_ (.A(\i_coord.x_row_start[-12] ),
    .X(_04178_));
 sg13g2_a21oi_1 _12177_ (.A1(_03985_),
    .A2(_04147_),
    .Y(_04179_),
    .B1(_04178_));
 sg13g2_nand3_1 _12178_ (.B(_03985_),
    .C(_04147_),
    .A(_04178_),
    .Y(_04180_));
 sg13g2_o21ai_1 _12179_ (.B1(_04180_),
    .Y(_04181_),
    .A1(_04176_),
    .A2(_04179_));
 sg13g2_buf_1 _12180_ (.A(_04181_),
    .X(_04182_));
 sg13g2_nor2_1 _12181_ (.A(_04175_),
    .B(_04182_),
    .Y(_04183_));
 sg13g2_a21oi_1 _12182_ (.A1(_04175_),
    .A2(_04182_),
    .Y(_04184_),
    .B1(\i_coord.l_xir.data_out[2] ));
 sg13g2_nor2_1 _12183_ (.A(_04183_),
    .B(_04184_),
    .Y(_04185_));
 sg13g2_a21o_1 _12184_ (.A2(_04185_),
    .A1(_04174_),
    .B1(\i_coord.l_xir.data_out[3] ),
    .X(_04186_));
 sg13g2_o21ai_1 _12185_ (.B1(_04186_),
    .Y(_04187_),
    .A1(_04174_),
    .A2(_04185_));
 sg13g2_buf_1 _12186_ (.A(_04187_),
    .X(_04189_));
 sg13g2_inv_1 _12187_ (.Y(_04190_),
    .A(_04189_));
 sg13g2_a21oi_1 _12188_ (.A1(_04172_),
    .A2(_04190_),
    .Y(_04191_),
    .B1(\i_coord.l_xir.data_out[4] ));
 sg13g2_a21oi_1 _12189_ (.A1(_04173_),
    .A2(_04189_),
    .Y(_04192_),
    .B1(_04191_));
 sg13g2_a21o_1 _12190_ (.A2(_04192_),
    .A1(_04171_),
    .B1(\i_coord.l_xir.data_out[5] ),
    .X(_04193_));
 sg13g2_o21ai_1 _12191_ (.B1(_04193_),
    .Y(_04194_),
    .A1(_04171_),
    .A2(_04192_));
 sg13g2_buf_1 _12192_ (.A(_04194_),
    .X(_04195_));
 sg13g2_inv_1 _12193_ (.Y(_04196_),
    .A(_04195_));
 sg13g2_a21oi_1 _12194_ (.A1(_04169_),
    .A2(_04196_),
    .Y(_04197_),
    .B1(\i_coord.l_xir.data_out[6] ));
 sg13g2_a21oi_2 _12195_ (.B1(_04197_),
    .Y(_04198_),
    .A2(_04195_),
    .A1(_04170_));
 sg13g2_and2_1 _12196_ (.A(_04168_),
    .B(_04198_),
    .X(_04200_));
 sg13g2_buf_1 _12197_ (.A(_04200_),
    .X(_04201_));
 sg13g2_a21oi_1 _12198_ (.A1(_04167_),
    .A2(_04201_),
    .Y(_04202_),
    .B1(net318));
 sg13g2_inv_1 _12199_ (.Y(_04203_),
    .A(_04167_));
 sg13g2_nor2_1 _12200_ (.A(_04168_),
    .B(_04198_),
    .Y(_04204_));
 sg13g2_inv_1 _12201_ (.Y(_04205_),
    .A(_04204_));
 sg13g2_a21oi_2 _12202_ (.B1(_04201_),
    .Y(_04206_),
    .A2(_04205_),
    .A1(_03999_));
 sg13g2_nand2_1 _12203_ (.Y(_04207_),
    .A(_04203_),
    .B(_04206_));
 sg13g2_buf_1 _12204_ (.A(\i_coord.x_row_start[-5] ),
    .X(_04208_));
 sg13g2_a21oi_1 _12205_ (.A1(net318),
    .A2(_04207_),
    .Y(_04209_),
    .B1(net316));
 sg13g2_nor2_1 _12206_ (.A(_04202_),
    .B(_04209_),
    .Y(_04211_));
 sg13g2_xnor2_1 _12207_ (.Y(_04212_),
    .A(_04165_),
    .B(_04211_));
 sg13g2_nor2_1 _12208_ (.A(net103),
    .B(_04212_),
    .Y(_04213_));
 sg13g2_buf_1 _12209_ (.A(\i_coord.x_row_start[-3] ),
    .X(_04214_));
 sg13g2_o21ai_1 _12210_ (.B1(net315),
    .Y(_04215_),
    .A1(net43),
    .A2(_04213_));
 sg13g2_buf_1 _12211_ (.A(_04163_),
    .X(_04216_));
 sg13g2_buf_1 _12212_ (.A(net102),
    .X(_04217_));
 sg13g2_nor2_1 _12213_ (.A(net315),
    .B(net88),
    .Y(_04218_));
 sg13g2_a22oi_1 _12214_ (.Y(_04219_),
    .B1(_04212_),
    .B2(_04218_),
    .A2(net66),
    .A1(\i_coord.l_xl.data_out[10] ));
 sg13g2_nand2_1 _12215_ (.Y(_00104_),
    .A(_04215_),
    .B(_04219_));
 sg13g2_nand4_1 _12216_ (.B(_04167_),
    .C(net315),
    .A(net316),
    .Y(_04221_),
    .D(_04198_));
 sg13g2_or4_1 _12217_ (.A(net316),
    .B(_04167_),
    .C(net315),
    .D(_04198_),
    .X(_04222_));
 sg13g2_a21oi_1 _12218_ (.A1(net318),
    .A2(_04222_),
    .Y(_04223_),
    .B1(_04168_));
 sg13g2_a21oi_2 _12219_ (.B1(_04223_),
    .Y(_04224_),
    .A2(_04221_),
    .A1(_04165_));
 sg13g2_xnor2_1 _12220_ (.Y(_04225_),
    .A(_04165_),
    .B(_04224_));
 sg13g2_nor2_1 _12221_ (.A(net103),
    .B(_04225_),
    .Y(_04226_));
 sg13g2_buf_1 _12222_ (.A(\i_coord.x_row_start[-2] ),
    .X(_04227_));
 sg13g2_o21ai_1 _12223_ (.B1(_04227_),
    .Y(_04228_),
    .A1(net43),
    .A2(_04226_));
 sg13g2_nor2_1 _12224_ (.A(_04227_),
    .B(net88),
    .Y(_04229_));
 sg13g2_a22oi_1 _12225_ (.Y(_04230_),
    .B1(_04225_),
    .B2(_04229_),
    .A2(net66),
    .A1(\i_coord.l_xl.data_out[11] ));
 sg13g2_nand2_1 _12226_ (.Y(_00105_),
    .A(_04228_),
    .B(_04230_));
 sg13g2_nor2b_1 _12227_ (.A(net318),
    .B_N(_04227_),
    .Y(_04232_));
 sg13g2_nand4_1 _12228_ (.B(_04167_),
    .C(net315),
    .A(net316),
    .Y(_04233_),
    .D(_04232_));
 sg13g2_nand2b_1 _12229_ (.Y(_04234_),
    .B(net318),
    .A_N(_04227_));
 sg13g2_or4_1 _12230_ (.A(net316),
    .B(_04214_),
    .C(_04207_),
    .D(_04234_),
    .X(_04235_));
 sg13g2_o21ai_1 _12231_ (.B1(_04235_),
    .Y(_04236_),
    .A1(_04206_),
    .A2(_04233_));
 sg13g2_nor2_1 _12232_ (.A(net103),
    .B(_04236_),
    .Y(_04237_));
 sg13g2_buf_1 _12233_ (.A(\i_coord.x_row_start[-1] ),
    .X(_04238_));
 sg13g2_o21ai_1 _12234_ (.B1(_04238_),
    .Y(_04239_),
    .A1(net43),
    .A2(_04237_));
 sg13g2_nor2_1 _12235_ (.A(_04238_),
    .B(net88),
    .Y(_04240_));
 sg13g2_a22oi_1 _12236_ (.Y(_04242_),
    .B1(_04236_),
    .B2(_04240_),
    .A2(net66),
    .A1(\i_coord.l_xl.data_out[12] ));
 sg13g2_nand2_1 _12237_ (.Y(_00106_),
    .A(_04239_),
    .B(_04242_));
 sg13g2_and2_1 _12238_ (.A(_04238_),
    .B(_04232_),
    .X(_04243_));
 sg13g2_buf_1 _12239_ (.A(_04243_),
    .X(_04244_));
 sg13g2_nor3_1 _12240_ (.A(_04238_),
    .B(_04224_),
    .C(_04234_),
    .Y(_04245_));
 sg13g2_a21o_1 _12241_ (.A2(_04244_),
    .A1(_04224_),
    .B1(_04245_),
    .X(_04246_));
 sg13g2_nor2_1 _12242_ (.A(net103),
    .B(_04246_),
    .Y(_04247_));
 sg13g2_buf_1 _12243_ (.A(\i_coord.x_row_start[0] ),
    .X(_04248_));
 sg13g2_o21ai_1 _12244_ (.B1(_04248_),
    .Y(_04249_),
    .A1(net43),
    .A2(_04247_));
 sg13g2_nor2_1 _12245_ (.A(_04248_),
    .B(net88),
    .Y(_04250_));
 sg13g2_a22oi_1 _12246_ (.Y(_04252_),
    .B1(_04246_),
    .B2(_04250_),
    .A2(net66),
    .A1(\i_coord.l_xl.data_out[13] ));
 sg13g2_nand2_1 _12247_ (.Y(_00107_),
    .A(_04249_),
    .B(_04252_));
 sg13g2_buf_1 _12248_ (.A(\i_coord.x_row_start[1] ),
    .X(_04253_));
 sg13g2_inv_1 _12249_ (.Y(_04254_),
    .A(_04253_));
 sg13g2_nor3_1 _12250_ (.A(_04238_),
    .B(_04248_),
    .C(_04234_),
    .Y(_04255_));
 sg13g2_nand2b_1 _12251_ (.Y(_04256_),
    .B(_04255_),
    .A_N(net315));
 sg13g2_nand3_1 _12252_ (.B(_04248_),
    .C(_04244_),
    .A(net315),
    .Y(_04257_));
 sg13g2_mux2_1 _12253_ (.A0(_04256_),
    .A1(_04257_),
    .S(_04211_),
    .X(_04258_));
 sg13g2_a21oi_1 _12254_ (.A1(_04156_),
    .A2(_04258_),
    .Y(_04259_),
    .B1(net49));
 sg13g2_nor3_1 _12255_ (.A(_04253_),
    .B(net102),
    .C(_04258_),
    .Y(_04260_));
 sg13g2_a21oi_1 _12256_ (.A1(\i_coord.l_xl.data_out[14] ),
    .A2(net77),
    .Y(_04262_),
    .B1(_04260_));
 sg13g2_o21ai_1 _12257_ (.B1(_04262_),
    .Y(_00108_),
    .A1(_04254_),
    .A2(_04259_));
 sg13g2_inv_1 _12258_ (.Y(_04263_),
    .A(\i_coord.x_row_start[2] ));
 sg13g2_nand2_1 _12259_ (.Y(_04264_),
    .A(_04254_),
    .B(_04255_));
 sg13g2_nand3_1 _12260_ (.B(_04253_),
    .C(_04244_),
    .A(_04248_),
    .Y(_04265_));
 sg13g2_mux2_1 _12261_ (.A0(_04264_),
    .A1(_04265_),
    .S(_04224_),
    .X(_04266_));
 sg13g2_a21oi_1 _12262_ (.A1(_04156_),
    .A2(_04266_),
    .Y(_04267_),
    .B1(net49));
 sg13g2_nor3_1 _12263_ (.A(\i_coord.x_row_start[2] ),
    .B(net102),
    .C(_04266_),
    .Y(_04268_));
 sg13g2_a21oi_1 _12264_ (.A1(\i_coord.l_xl.data_out[15] ),
    .A2(net77),
    .Y(_04269_),
    .B1(_04268_));
 sg13g2_o21ai_1 _12265_ (.B1(_04269_),
    .Y(_00109_),
    .A1(_04263_),
    .A2(_04267_));
 sg13g2_nand2_1 _12266_ (.Y(_04271_),
    .A(_03985_),
    .B(_04147_));
 sg13g2_xnor2_1 _12267_ (.Y(_04272_),
    .A(\i_coord.l_xir.data_out[1] ),
    .B(_04271_));
 sg13g2_nand2_1 _12268_ (.Y(_04273_),
    .A(net131),
    .B(_04272_));
 sg13g2_nor2_1 _12269_ (.A(net102),
    .B(_04272_),
    .Y(_04274_));
 sg13g2_o21ai_1 _12270_ (.B1(_04178_),
    .Y(_04275_),
    .A1(net49),
    .A2(_04274_));
 sg13g2_o21ai_1 _12271_ (.B1(_04275_),
    .Y(_00110_),
    .A1(_04178_),
    .A2(_04273_));
 sg13g2_xor2_1 _12272_ (.B(_04182_),
    .A(\i_coord.l_xir.data_out[2] ),
    .X(_04276_));
 sg13g2_nand2_1 _12273_ (.Y(_04277_),
    .A(net131),
    .B(_04276_));
 sg13g2_nor2_1 _12274_ (.A(_04216_),
    .B(_04276_),
    .Y(_04278_));
 sg13g2_o21ai_1 _12275_ (.B1(_04175_),
    .Y(_04279_),
    .A1(net49),
    .A2(_04278_));
 sg13g2_o21ai_1 _12276_ (.B1(_04279_),
    .Y(_00111_),
    .A1(_04175_),
    .A2(_04277_));
 sg13g2_xor2_1 _12277_ (.B(_04185_),
    .A(\i_coord.l_xir.data_out[3] ),
    .X(_04281_));
 sg13g2_nor2_1 _12278_ (.A(net103),
    .B(_04281_),
    .Y(_04282_));
 sg13g2_o21ai_1 _12279_ (.B1(_04174_),
    .Y(_04283_),
    .A1(net43),
    .A2(_04282_));
 sg13g2_nor2_1 _12280_ (.A(_04174_),
    .B(net88),
    .Y(_04284_));
 sg13g2_a22oi_1 _12281_ (.Y(_04285_),
    .B1(_04281_),
    .B2(_04284_),
    .A2(_04146_),
    .A1(\i_coord.l_xl.data_out[3] ));
 sg13g2_nand2_1 _12282_ (.Y(_00112_),
    .A(_04283_),
    .B(_04285_));
 sg13g2_xnor2_1 _12283_ (.Y(_04286_),
    .A(\i_coord.l_xir.data_out[4] ),
    .B(_04189_));
 sg13g2_nor2_1 _12284_ (.A(net103),
    .B(_04286_),
    .Y(_04287_));
 sg13g2_o21ai_1 _12285_ (.B1(_04172_),
    .Y(_04288_),
    .A1(net43),
    .A2(_04287_));
 sg13g2_nor2_1 _12286_ (.A(_04172_),
    .B(net88),
    .Y(_04290_));
 sg13g2_a22oi_1 _12287_ (.Y(_04291_),
    .B1(_04286_),
    .B2(_04290_),
    .A2(net66),
    .A1(\i_coord.l_xl.data_out[4] ));
 sg13g2_nand2_1 _12288_ (.Y(_00113_),
    .A(_04288_),
    .B(_04291_));
 sg13g2_xor2_1 _12289_ (.B(_04192_),
    .A(\i_coord.l_xir.data_out[5] ),
    .X(_04292_));
 sg13g2_nor2_1 _12290_ (.A(net103),
    .B(_04292_),
    .Y(_04293_));
 sg13g2_o21ai_1 _12291_ (.B1(_04171_),
    .Y(_04294_),
    .A1(net43),
    .A2(_04293_));
 sg13g2_nor2_1 _12292_ (.A(_04171_),
    .B(net88),
    .Y(_04295_));
 sg13g2_a22oi_1 _12293_ (.Y(_04296_),
    .B1(_04292_),
    .B2(_04295_),
    .A2(_04146_),
    .A1(\i_coord.l_xl.data_out[5] ));
 sg13g2_nand2_1 _12294_ (.Y(_00114_),
    .A(_04294_),
    .B(_04296_));
 sg13g2_xnor2_1 _12295_ (.Y(_04297_),
    .A(\i_coord.l_xir.data_out[6] ),
    .B(_04195_));
 sg13g2_nor2_1 _12296_ (.A(net103),
    .B(_04297_),
    .Y(_04299_));
 sg13g2_o21ai_1 _12297_ (.B1(_04169_),
    .Y(_04300_),
    .A1(net43),
    .A2(_04299_));
 sg13g2_nor2_1 _12298_ (.A(_04169_),
    .B(net88),
    .Y(_04301_));
 sg13g2_a22oi_1 _12299_ (.Y(_04302_),
    .B1(_04297_),
    .B2(_04301_),
    .A2(net77),
    .A1(\i_coord.l_xl.data_out[6] ));
 sg13g2_nand2_1 _12300_ (.Y(_00115_),
    .A(_04300_),
    .B(_04302_));
 sg13g2_xnor2_1 _12301_ (.Y(_04303_),
    .A(_04165_),
    .B(_04198_));
 sg13g2_nor2_1 _12302_ (.A(_04164_),
    .B(_04303_),
    .Y(_04304_));
 sg13g2_o21ai_1 _12303_ (.B1(_04168_),
    .Y(_04305_),
    .A1(_04161_),
    .A2(_04304_));
 sg13g2_nor2_1 _12304_ (.A(_04168_),
    .B(_04217_),
    .Y(_04306_));
 sg13g2_a22oi_1 _12305_ (.Y(_04307_),
    .B1(_04303_),
    .B2(_04306_),
    .A2(net77),
    .A1(\i_coord.l_xl.data_out[7] ));
 sg13g2_nand2_1 _12306_ (.Y(_00116_),
    .A(_04305_),
    .B(_04307_));
 sg13g2_xnor2_1 _12307_ (.Y(_04309_),
    .A(net318),
    .B(_04206_));
 sg13g2_nor2_1 _12308_ (.A(_04164_),
    .B(_04309_),
    .Y(_04310_));
 sg13g2_o21ai_1 _12309_ (.B1(net316),
    .Y(_04311_),
    .A1(_04160_),
    .A2(_04310_));
 sg13g2_nor2_1 _12310_ (.A(net316),
    .B(_04217_),
    .Y(_04312_));
 sg13g2_a22oi_1 _12311_ (.Y(_04313_),
    .B1(_04309_),
    .B2(_04312_),
    .A2(net77),
    .A1(\i_coord.l_xl.data_out[8] ));
 sg13g2_nand2_1 _12312_ (.Y(_00117_),
    .A(_04311_),
    .B(_04313_));
 sg13g2_nor2b_1 _12313_ (.A(net318),
    .B_N(net316),
    .Y(_04314_));
 sg13g2_nor2_1 _12314_ (.A(_04165_),
    .B(_04208_),
    .Y(_04315_));
 sg13g2_a22oi_1 _12315_ (.Y(_04316_),
    .B1(_04315_),
    .B2(_04204_),
    .A2(_04314_),
    .A1(_04201_));
 sg13g2_a21oi_1 _12316_ (.A1(_04156_),
    .A2(_04316_),
    .Y(_04318_),
    .B1(_04160_));
 sg13g2_nor3_1 _12317_ (.A(_04167_),
    .B(_04216_),
    .C(_04316_),
    .Y(_04319_));
 sg13g2_a21oi_1 _12318_ (.A1(\i_coord.l_xl.data_out[9] ),
    .A2(_04144_),
    .Y(_04320_),
    .B1(_04319_));
 sg13g2_o21ai_1 _12319_ (.B1(_04320_),
    .Y(_00118_),
    .A1(_04203_),
    .A2(_04318_));
 sg13g2_buf_1 _12320_ (.A(_04420_),
    .X(_04321_));
 sg13g2_nand2_1 _12321_ (.Y(_04322_),
    .A(_03882_),
    .B(net58));
 sg13g2_buf_1 _12322_ (.A(_04322_),
    .X(_04323_));
 sg13g2_buf_1 _12323_ (.A(_04323_),
    .X(_04324_));
 sg13g2_nor2_1 _12324_ (.A(_03881_),
    .B(_04280_),
    .Y(_04325_));
 sg13g2_buf_1 _12325_ (.A(_04325_),
    .X(_04326_));
 sg13g2_buf_1 _12326_ (.A(_04326_),
    .X(_04328_));
 sg13g2_or2_1 _12327_ (.X(_04329_),
    .B(_04280_),
    .A(net274));
 sg13g2_buf_1 _12328_ (.A(_04329_),
    .X(_04330_));
 sg13g2_buf_1 _12329_ (.A(\i_coord.y_row_start[-13] ),
    .X(_04331_));
 sg13g2_nand2_1 _12330_ (.Y(_04332_),
    .A(net322),
    .B(_04331_));
 sg13g2_or2_1 _12331_ (.X(_04333_),
    .B(_04332_),
    .A(_04330_));
 sg13g2_o21ai_1 _12332_ (.B1(_04333_),
    .Y(_04334_),
    .A1(\i_coord.l_yt.data_out[0] ),
    .A2(_04328_));
 sg13g2_buf_1 _12333_ (.A(_04330_),
    .X(_04335_));
 sg13g2_o21ai_1 _12334_ (.B1(_04324_),
    .Y(_04336_),
    .A1(net322),
    .A2(_04335_));
 sg13g2_inv_1 _12335_ (.Y(_04337_),
    .A(_04331_));
 sg13g2_a22oi_1 _12336_ (.Y(_00127_),
    .B1(_04336_),
    .B2(_04337_),
    .A2(_04334_),
    .A1(_04324_));
 sg13g2_inv_1 _12337_ (.Y(_04339_),
    .A(\i_coord.l_yt.data_out[10] ));
 sg13g2_buf_2 _12338_ (.A(\i_coord.y_row_start[-3] ),
    .X(_04340_));
 sg13g2_buf_1 _12339_ (.A(_03839_),
    .X(_04341_));
 sg13g2_buf_1 _12340_ (.A(net55),
    .X(_04342_));
 sg13g2_buf_2 _12341_ (.A(\i_coord.y_row_start[-5] ),
    .X(_04343_));
 sg13g2_buf_1 _12342_ (.A(\i_coord.y_row_start[-4] ),
    .X(_04344_));
 sg13g2_inv_1 _12343_ (.Y(_04345_),
    .A(\i_coord.y_row_start[-7] ));
 sg13g2_buf_1 _12344_ (.A(\i_coord.y_row_start[-8] ),
    .X(_04346_));
 sg13g2_buf_1 _12345_ (.A(\i_coord.y_row_start[-9] ),
    .X(_04347_));
 sg13g2_buf_1 _12346_ (.A(\i_coord.y_row_start[-10] ),
    .X(_04349_));
 sg13g2_buf_1 _12347_ (.A(\i_coord.y_row_start[-12] ),
    .X(_04350_));
 sg13g2_nand2b_1 _12348_ (.Y(_04351_),
    .B(_04332_),
    .A_N(_04350_));
 sg13g2_and3_1 _12349_ (.X(_04352_),
    .A(net322),
    .B(_04331_),
    .C(_04350_));
 sg13g2_a21oi_1 _12350_ (.A1(_03894_),
    .A2(_04351_),
    .Y(_04353_),
    .B1(_04352_));
 sg13g2_buf_1 _12351_ (.A(\i_coord.y_row_start[-11] ),
    .X(_04354_));
 sg13g2_nand2_1 _12352_ (.Y(_04355_),
    .A(_03887_),
    .B(_04354_));
 sg13g2_nor2_1 _12353_ (.A(_03887_),
    .B(_04354_),
    .Y(_04356_));
 sg13g2_a21oi_2 _12354_ (.B1(_04356_),
    .Y(_04357_),
    .A2(_04355_),
    .A1(_04353_));
 sg13g2_nor2_1 _12355_ (.A(_04349_),
    .B(_04357_),
    .Y(_04358_));
 sg13g2_a21oi_1 _12356_ (.A1(_04349_),
    .A2(_04357_),
    .Y(_04360_),
    .B1(_03888_));
 sg13g2_nor2_1 _12357_ (.A(_04358_),
    .B(_04360_),
    .Y(_04361_));
 sg13g2_nor2_1 _12358_ (.A(_04347_),
    .B(_04361_),
    .Y(_04362_));
 sg13g2_a21oi_1 _12359_ (.A1(_04347_),
    .A2(_04361_),
    .Y(_04363_),
    .B1(_03890_));
 sg13g2_nor2_1 _12360_ (.A(_04362_),
    .B(_04363_),
    .Y(_04364_));
 sg13g2_a21o_1 _12361_ (.A2(_04364_),
    .A1(_04346_),
    .B1(_03889_),
    .X(_04365_));
 sg13g2_o21ai_1 _12362_ (.B1(_04365_),
    .Y(_04366_),
    .A1(_04346_),
    .A2(_04364_));
 sg13g2_buf_1 _12363_ (.A(_04366_),
    .X(_04367_));
 sg13g2_a21o_1 _12364_ (.A2(_04367_),
    .A1(_04345_),
    .B1(_03892_),
    .X(_04368_));
 sg13g2_o21ai_1 _12365_ (.B1(_04368_),
    .Y(_04369_),
    .A1(_04345_),
    .A2(_04367_));
 sg13g2_buf_2 _12366_ (.A(_04369_),
    .X(_04371_));
 sg13g2_nand3_1 _12367_ (.B(_04344_),
    .C(_04371_),
    .A(_04343_),
    .Y(_04372_));
 sg13g2_or3_1 _12368_ (.A(_04343_),
    .B(_04344_),
    .C(_04371_),
    .X(_04373_));
 sg13g2_buf_1 _12369_ (.A(\i_coord.y_row_start[-6] ),
    .X(_04374_));
 sg13g2_a21oi_1 _12370_ (.A1(net321),
    .A2(_04373_),
    .Y(_04375_),
    .B1(_04374_));
 sg13g2_a21oi_2 _12371_ (.B1(_04375_),
    .Y(_04376_),
    .A2(_04372_),
    .A1(net226));
 sg13g2_xor2_1 _12372_ (.B(_04340_),
    .A(net321),
    .X(_04377_));
 sg13g2_xnor2_1 _12373_ (.Y(_04378_),
    .A(_04376_),
    .B(_04377_));
 sg13g2_nand2_1 _12374_ (.Y(_04379_),
    .A(net131),
    .B(_04378_));
 sg13g2_o21ai_1 _12375_ (.B1(_04379_),
    .Y(_04380_),
    .A1(_04340_),
    .A2(net48));
 sg13g2_a22oi_1 _12376_ (.Y(_00128_),
    .B1(_04380_),
    .B2(net223),
    .A2(net56),
    .A1(_04339_));
 sg13g2_buf_2 _12377_ (.A(\i_coord.y_row_start[-2] ),
    .X(_04382_));
 sg13g2_nand4_1 _12378_ (.B(_04344_),
    .C(_04340_),
    .A(_04343_),
    .Y(_04383_),
    .D(_04371_));
 sg13g2_or2_1 _12379_ (.X(_04384_),
    .B(_04373_),
    .A(_04340_));
 sg13g2_a21oi_1 _12380_ (.A1(net321),
    .A2(_04384_),
    .Y(_04385_),
    .B1(_04374_));
 sg13g2_a21oi_1 _12381_ (.A1(net226),
    .A2(_04383_),
    .Y(_04386_),
    .B1(_04385_));
 sg13g2_xor2_1 _12382_ (.B(_04382_),
    .A(net321),
    .X(_04387_));
 sg13g2_xnor2_1 _12383_ (.Y(_04388_),
    .A(_04386_),
    .B(_04387_));
 sg13g2_nand2_1 _12384_ (.Y(_04389_),
    .A(net131),
    .B(_04388_));
 sg13g2_o21ai_1 _12385_ (.B1(_04389_),
    .Y(_04390_),
    .A1(_04382_),
    .A2(net48));
 sg13g2_a22oi_1 _12386_ (.Y(_00129_),
    .B1(_04390_),
    .B2(net223),
    .A2(net56),
    .A1(_04075_));
 sg13g2_buf_1 _12387_ (.A(\i_coord.y_row_start[-1] ),
    .X(_04392_));
 sg13g2_nand2_1 _12388_ (.Y(_04393_),
    .A(net226),
    .B(_04382_));
 sg13g2_nand2_1 _12389_ (.Y(_04394_),
    .A(_04340_),
    .B(_04376_));
 sg13g2_nor2_1 _12390_ (.A(_04340_),
    .B(_04376_),
    .Y(_04395_));
 sg13g2_nand3b_1 _12391_ (.B(_04395_),
    .C(net321),
    .Y(_04396_),
    .A_N(_04382_));
 sg13g2_o21ai_1 _12392_ (.B1(_04396_),
    .Y(_04397_),
    .A1(_04393_),
    .A2(_04394_));
 sg13g2_nand3_1 _12393_ (.B(net57),
    .C(_04397_),
    .A(_04392_),
    .Y(_04398_));
 sg13g2_o21ai_1 _12394_ (.B1(_04398_),
    .Y(_04399_),
    .A1(\i_coord.l_yt.data_out[12] ),
    .A2(net57));
 sg13g2_o21ai_1 _12395_ (.B1(net37),
    .Y(_04400_),
    .A1(net56),
    .A2(_04397_));
 sg13g2_inv_1 _12396_ (.Y(_04402_),
    .A(_04392_));
 sg13g2_a22oi_1 _12397_ (.Y(_00130_),
    .B1(_04400_),
    .B2(_04402_),
    .A2(_04399_),
    .A1(net37));
 sg13g2_nor3_1 _12398_ (.A(net226),
    .B(_04382_),
    .C(_04392_),
    .Y(_04403_));
 sg13g2_and3_1 _12399_ (.X(_04404_),
    .A(net226),
    .B(_04382_),
    .C(_04392_));
 sg13g2_mux2_1 _12400_ (.A0(_04403_),
    .A1(_04404_),
    .S(_04386_),
    .X(_04405_));
 sg13g2_nor2_1 _12401_ (.A(net102),
    .B(_04405_),
    .Y(_04406_));
 sg13g2_buf_1 _12402_ (.A(\i_coord.y_row_start[0] ),
    .X(_04407_));
 sg13g2_inv_1 _12403_ (.Y(_04408_),
    .A(_04407_));
 sg13g2_o21ai_1 _12404_ (.B1(_04408_),
    .Y(_04409_),
    .A1(net49),
    .A2(_04406_));
 sg13g2_nand3_1 _12405_ (.B(net104),
    .C(_04405_),
    .A(_04407_),
    .Y(_04410_));
 sg13g2_nand2_1 _12406_ (.Y(_04412_),
    .A(_04409_),
    .B(_04410_));
 sg13g2_a22oi_1 _12407_ (.Y(_00131_),
    .B1(_04412_),
    .B2(net223),
    .A2(net56),
    .A1(_04089_));
 sg13g2_nand2_1 _12408_ (.Y(_04413_),
    .A(_04407_),
    .B(_04404_));
 sg13g2_nand3_1 _12409_ (.B(_04395_),
    .C(_04403_),
    .A(_04408_),
    .Y(_04414_));
 sg13g2_o21ai_1 _12410_ (.B1(_04414_),
    .Y(_04415_),
    .A1(_04394_),
    .A2(_04413_));
 sg13g2_nand3_1 _12411_ (.B(net57),
    .C(_04415_),
    .A(\i_coord.y_row_start[1] ),
    .Y(_04416_));
 sg13g2_o21ai_1 _12412_ (.B1(_04416_),
    .Y(_04417_),
    .A1(\i_coord.l_yt.data_out[14] ),
    .A2(net57));
 sg13g2_o21ai_1 _12413_ (.B1(net37),
    .Y(_04418_),
    .A1(net56),
    .A2(_04415_));
 sg13g2_inv_1 _12414_ (.Y(_04419_),
    .A(\i_coord.y_row_start[1] ));
 sg13g2_a22oi_1 _12415_ (.Y(_00132_),
    .B1(_04418_),
    .B2(_04419_),
    .A2(_04417_),
    .A1(net37));
 sg13g2_inv_1 _12416_ (.Y(_04421_),
    .A(\i_coord.l_yt.data_out[1] ));
 sg13g2_xnor2_1 _12417_ (.Y(_04422_),
    .A(_03894_),
    .B(_04350_));
 sg13g2_xnor2_1 _12418_ (.Y(_04423_),
    .A(_04332_),
    .B(_04422_));
 sg13g2_nand2_1 _12419_ (.Y(_04424_),
    .A(net131),
    .B(_04423_));
 sg13g2_o21ai_1 _12420_ (.B1(_04424_),
    .Y(_04425_),
    .A1(_04350_),
    .A2(net48));
 sg13g2_a22oi_1 _12421_ (.Y(_00133_),
    .B1(_04425_),
    .B2(net223),
    .A2(net56),
    .A1(_04421_));
 sg13g2_xnor2_1 _12422_ (.Y(_04426_),
    .A(_03887_),
    .B(_04353_));
 sg13g2_nand3_1 _12423_ (.B(_04326_),
    .C(_04426_),
    .A(_04354_),
    .Y(_04427_));
 sg13g2_o21ai_1 _12424_ (.B1(_04427_),
    .Y(_04428_),
    .A1(\i_coord.l_yt.data_out[2] ),
    .A2(_04328_));
 sg13g2_o21ai_1 _12425_ (.B1(_04323_),
    .Y(_04429_),
    .A1(_04330_),
    .A2(_04426_));
 sg13g2_inv_1 _12426_ (.Y(_04431_),
    .A(_04354_));
 sg13g2_a22oi_1 _12427_ (.Y(_00134_),
    .B1(_04429_),
    .B2(_04431_),
    .A2(_04428_),
    .A1(net37));
 sg13g2_buf_1 _12428_ (.A(net58),
    .X(_04432_));
 sg13g2_xor2_1 _12429_ (.B(_04349_),
    .A(_03888_),
    .X(_04433_));
 sg13g2_xnor2_1 _12430_ (.Y(_04434_),
    .A(_04357_),
    .B(_04433_));
 sg13g2_nor2_1 _12431_ (.A(net102),
    .B(_04434_),
    .Y(_04435_));
 sg13g2_a21oi_1 _12432_ (.A1(_04349_),
    .A2(net47),
    .Y(_04436_),
    .B1(_04435_));
 sg13g2_nand2_1 _12433_ (.Y(_04437_),
    .A(\i_coord.l_yt.data_out[3] ),
    .B(_04335_));
 sg13g2_o21ai_1 _12434_ (.B1(_04437_),
    .Y(_00135_),
    .A1(net221),
    .A2(_04436_));
 sg13g2_xor2_1 _12435_ (.B(_04361_),
    .A(_03890_),
    .X(_04438_));
 sg13g2_nand3_1 _12436_ (.B(_04326_),
    .C(_04438_),
    .A(_04347_),
    .Y(_04440_));
 sg13g2_o21ai_1 _12437_ (.B1(_04440_),
    .Y(_04441_),
    .A1(\i_coord.l_yt.data_out[4] ),
    .A2(net57));
 sg13g2_o21ai_1 _12438_ (.B1(_04323_),
    .Y(_04442_),
    .A1(_04330_),
    .A2(_04438_));
 sg13g2_inv_1 _12439_ (.Y(_04443_),
    .A(_04347_));
 sg13g2_a22oi_1 _12440_ (.Y(_00136_),
    .B1(_04442_),
    .B2(_04443_),
    .A2(_04441_),
    .A1(net37));
 sg13g2_xor2_1 _12441_ (.B(_04364_),
    .A(_03889_),
    .X(_04444_));
 sg13g2_nand3_1 _12442_ (.B(_04326_),
    .C(_04444_),
    .A(_04346_),
    .Y(_04445_));
 sg13g2_o21ai_1 _12443_ (.B1(_04445_),
    .Y(_04446_),
    .A1(\i_coord.l_yt.data_out[5] ),
    .A2(net57));
 sg13g2_o21ai_1 _12444_ (.B1(_04323_),
    .Y(_04447_),
    .A1(_04330_),
    .A2(_04444_));
 sg13g2_inv_1 _12445_ (.Y(_04448_),
    .A(_04346_));
 sg13g2_a22oi_1 _12446_ (.Y(_00137_),
    .B1(_04447_),
    .B2(_04448_),
    .A2(_04446_),
    .A1(net37));
 sg13g2_xnor2_1 _12447_ (.Y(_04450_),
    .A(_03892_),
    .B(_04367_));
 sg13g2_a21oi_1 _12448_ (.A1(net131),
    .A2(_04450_),
    .Y(_04451_),
    .B1(net47));
 sg13g2_nor2_1 _12449_ (.A(_04345_),
    .B(_04451_),
    .Y(_04452_));
 sg13g2_nor3_1 _12450_ (.A(\i_coord.y_row_start[-7] ),
    .B(net102),
    .C(_04450_),
    .Y(_04453_));
 sg13g2_o21ai_1 _12451_ (.B1(net223),
    .Y(_04454_),
    .A1(_04452_),
    .A2(_04453_));
 sg13g2_o21ai_1 _12452_ (.B1(_04454_),
    .Y(_00138_),
    .A1(_04123_),
    .A2(net57));
 sg13g2_inv_1 _12453_ (.Y(_04455_),
    .A(_04374_));
 sg13g2_nand2_1 _12454_ (.Y(_04456_),
    .A(net226),
    .B(_04374_));
 sg13g2_nand2_1 _12455_ (.Y(_04457_),
    .A(net321),
    .B(_04455_));
 sg13g2_nand2_1 _12456_ (.Y(_04459_),
    .A(_04456_),
    .B(_04457_));
 sg13g2_xnor2_1 _12457_ (.Y(_04460_),
    .A(_04371_),
    .B(_04459_));
 sg13g2_a22oi_1 _12458_ (.Y(_04461_),
    .B1(_04156_),
    .B2(_04460_),
    .A2(net47),
    .A1(_04455_));
 sg13g2_nor2_1 _12459_ (.A(net221),
    .B(_04461_),
    .Y(_04462_));
 sg13g2_a21oi_1 _12460_ (.A1(_04130_),
    .A2(net56),
    .Y(_00139_),
    .B1(_04462_));
 sg13g2_mux2_1 _12461_ (.A0(_04457_),
    .A1(_04456_),
    .S(_04371_),
    .X(_04463_));
 sg13g2_a21oi_1 _12462_ (.A1(net131),
    .A2(_04463_),
    .Y(_04464_),
    .B1(net47));
 sg13g2_nand2b_1 _12463_ (.Y(_04465_),
    .B(_04343_),
    .A_N(_04464_));
 sg13g2_or3_1 _12464_ (.A(_04343_),
    .B(net102),
    .C(_04463_),
    .X(_04466_));
 sg13g2_a21oi_1 _12465_ (.A1(_04465_),
    .A2(_04466_),
    .Y(_04467_),
    .B1(net221));
 sg13g2_a21o_1 _12466_ (.A2(net56),
    .A1(\i_coord.l_yt.data_out[8] ),
    .B1(_04467_),
    .X(_00140_));
 sg13g2_nor3_1 _12467_ (.A(_04343_),
    .B(_04371_),
    .C(_04457_),
    .Y(_04469_));
 sg13g2_nand4_1 _12468_ (.B(_04374_),
    .C(_04343_),
    .A(net226),
    .Y(_04470_),
    .D(_04371_));
 sg13g2_nand2b_1 _12469_ (.Y(_04471_),
    .B(_04470_),
    .A_N(_04469_));
 sg13g2_nand3_1 _12470_ (.B(_04326_),
    .C(_04471_),
    .A(_04344_),
    .Y(_04472_));
 sg13g2_o21ai_1 _12471_ (.B1(_04472_),
    .Y(_04473_),
    .A1(\i_coord.l_yt.data_out[9] ),
    .A2(net57));
 sg13g2_o21ai_1 _12472_ (.B1(_04323_),
    .Y(_04474_),
    .A1(_04330_),
    .A2(_04471_));
 sg13g2_inv_1 _12473_ (.Y(_04475_),
    .A(_04344_));
 sg13g2_a22oi_1 _12474_ (.Y(_00141_),
    .B1(_04474_),
    .B2(_04475_),
    .A2(_04473_),
    .A1(net37));
 sg13g2_nand2_1 _12475_ (.Y(_04476_),
    .A(_04136_),
    .B(_04118_));
 sg13g2_nor4_1 _12476_ (.A(_04127_),
    .B(_04231_),
    .C(_04251_),
    .D(_04476_),
    .Y(_04478_));
 sg13g2_buf_1 _12477_ (.A(_04478_),
    .X(_04479_));
 sg13g2_buf_1 _12478_ (.A(_04479_),
    .X(_04480_));
 sg13g2_buf_2 _12479_ (.A(\i_coord.x0[-13] ),
    .X(_04481_));
 sg13g2_buf_1 _12480_ (.A(_03945_),
    .X(_04482_));
 sg13g2_buf_1 _12481_ (.A(_03945_),
    .X(_04483_));
 sg13g2_buf_1 _12482_ (.A(_03839_),
    .X(_04484_));
 sg13g2_or4_1 _12483_ (.A(_03998_),
    .B(net336),
    .C(_04071_),
    .D(_04027_),
    .X(_04485_));
 sg13g2_nor3_1 _12484_ (.A(_04081_),
    .B(_04348_),
    .C(_04485_),
    .Y(_04486_));
 sg13g2_nor2b_1 _12485_ (.A(_03964_),
    .B_N(_00033_),
    .Y(_04487_));
 sg13g2_a21oi_1 _12486_ (.A1(_03861_),
    .A2(_04486_),
    .Y(_04489_),
    .B1(_04034_));
 sg13g2_a21oi_1 _12487_ (.A1(_04486_),
    .A2(_04487_),
    .Y(_04490_),
    .B1(_04489_));
 sg13g2_nor2_1 _12488_ (.A(\i_vga.vblank ),
    .B(_04490_),
    .Y(_04491_));
 sg13g2_buf_2 _12489_ (.A(_04491_),
    .X(_04492_));
 sg13g2_o21ai_1 _12490_ (.B1(_04492_),
    .Y(_04493_),
    .A1(_03877_),
    .A2(net54));
 sg13g2_or2_1 _12491_ (.X(_04494_),
    .B(_04490_),
    .A(\i_vga.vblank ));
 sg13g2_buf_1 _12492_ (.A(_04494_),
    .X(_04495_));
 sg13g2_nor2_1 _12493_ (.A(net54),
    .B(net82),
    .Y(_04496_));
 sg13g2_nor2b_1 _12494_ (.A(_04481_),
    .B_N(_03877_),
    .Y(_04497_));
 sg13g2_a22oi_1 _12495_ (.Y(_04498_),
    .B1(_04496_),
    .B2(_04497_),
    .A2(_04493_),
    .A1(_04481_));
 sg13g2_nand2_1 _12496_ (.Y(_04500_),
    .A(net140),
    .B(_04498_));
 sg13g2_o21ai_1 _12497_ (.B1(_04500_),
    .Y(_04501_),
    .A1(_04481_),
    .A2(net141));
 sg13g2_nor3_1 _12498_ (.A(net76),
    .B(net104),
    .C(_04501_),
    .Y(_04502_));
 sg13g2_a21o_1 _12499_ (.A2(_04156_),
    .A1(_04147_),
    .B1(_04502_),
    .X(_00177_));
 sg13g2_buf_1 _12500_ (.A(\i_coord.x0[-3] ),
    .X(_04503_));
 sg13g2_buf_1 _12501_ (.A(\i_coord.x0[-4] ),
    .X(_04504_));
 sg13g2_inv_1 _12502_ (.Y(_04505_),
    .A(_04504_));
 sg13g2_buf_2 _12503_ (.A(\i_coord.x0[-5] ),
    .X(_04506_));
 sg13g2_buf_1 _12504_ (.A(\i_coord.x0[-6] ),
    .X(_04507_));
 sg13g2_inv_1 _12505_ (.Y(_04508_),
    .A(_04507_));
 sg13g2_buf_2 _12506_ (.A(\i_coord.x0[-7] ),
    .X(_04510_));
 sg13g2_buf_1 _12507_ (.A(\i_coord.x0[-8] ),
    .X(_04511_));
 sg13g2_inv_1 _12508_ (.Y(_04512_),
    .A(_04511_));
 sg13g2_buf_1 _12509_ (.A(\i_coord.x0[-9] ),
    .X(_04513_));
 sg13g2_buf_2 _12510_ (.A(\i_coord.x0[-10] ),
    .X(_04514_));
 sg13g2_buf_2 _12511_ (.A(\i_coord.x0[-11] ),
    .X(_04515_));
 sg13g2_buf_2 _12512_ (.A(\i_coord.x0[-12] ),
    .X(_04516_));
 sg13g2_nor2_1 _12513_ (.A(_03919_),
    .B(_04516_),
    .Y(_04517_));
 sg13g2_nand2_1 _12514_ (.Y(_04518_),
    .A(_03877_),
    .B(_04481_));
 sg13g2_nand2_1 _12515_ (.Y(_04519_),
    .A(_03919_),
    .B(_04516_));
 sg13g2_o21ai_1 _12516_ (.B1(_04519_),
    .Y(_04521_),
    .A1(_04517_),
    .A2(_04518_));
 sg13g2_buf_1 _12517_ (.A(_04521_),
    .X(_04522_));
 sg13g2_nor2_1 _12518_ (.A(_04515_),
    .B(_04522_),
    .Y(_04523_));
 sg13g2_a21oi_1 _12519_ (.A1(_04515_),
    .A2(_04522_),
    .Y(_04524_),
    .B1(\i_coord.l_xip.data_out[2] ));
 sg13g2_nor2_1 _12520_ (.A(_04523_),
    .B(_04524_),
    .Y(_04525_));
 sg13g2_nor2_1 _12521_ (.A(_04514_),
    .B(_04525_),
    .Y(_04526_));
 sg13g2_a21oi_1 _12522_ (.A1(_04514_),
    .A2(_04525_),
    .Y(_04527_),
    .B1(\i_coord.l_xip.data_out[3] ));
 sg13g2_nor2_1 _12523_ (.A(_04526_),
    .B(_04527_),
    .Y(_04528_));
 sg13g2_a21o_1 _12524_ (.A2(_04528_),
    .A1(net313),
    .B1(\i_coord.l_xip.data_out[4] ),
    .X(_04529_));
 sg13g2_o21ai_1 _12525_ (.B1(_04529_),
    .Y(_04530_),
    .A1(net313),
    .A2(_04528_));
 sg13g2_buf_1 _12526_ (.A(_04530_),
    .X(_04532_));
 sg13g2_inv_1 _12527_ (.Y(_04533_),
    .A(_04532_));
 sg13g2_a21oi_1 _12528_ (.A1(_04511_),
    .A2(_04533_),
    .Y(_04534_),
    .B1(\i_coord.l_xip.data_out[5] ));
 sg13g2_a21oi_1 _12529_ (.A1(_04512_),
    .A2(_04532_),
    .Y(_04535_),
    .B1(_04534_));
 sg13g2_a21o_1 _12530_ (.A2(_04535_),
    .A1(_04510_),
    .B1(\i_coord.l_xip.data_out[6] ),
    .X(_04536_));
 sg13g2_o21ai_1 _12531_ (.B1(_04536_),
    .Y(_04537_),
    .A1(_04510_),
    .A2(_04535_));
 sg13g2_buf_1 _12532_ (.A(_04537_),
    .X(_04538_));
 sg13g2_inv_1 _12533_ (.Y(_04539_),
    .A(_04538_));
 sg13g2_a21oi_1 _12534_ (.A1(_04507_),
    .A2(_04539_),
    .Y(_04540_),
    .B1(\i_coord.l_xip.data_out[7] ));
 sg13g2_a21oi_1 _12535_ (.A1(_04508_),
    .A2(_04538_),
    .Y(_04541_),
    .B1(_04540_));
 sg13g2_nor2_1 _12536_ (.A(_04506_),
    .B(_04541_),
    .Y(_04543_));
 sg13g2_a21oi_1 _12537_ (.A1(_04506_),
    .A2(_04541_),
    .Y(_04544_),
    .B1(\i_coord.l_xip.data_out[8] ));
 sg13g2_nor3_1 _12538_ (.A(_04505_),
    .B(_04543_),
    .C(_04544_),
    .Y(_04545_));
 sg13g2_nor2_1 _12539_ (.A(net319),
    .B(_04545_),
    .Y(_04546_));
 sg13g2_nor2_2 _12540_ (.A(_04543_),
    .B(_04544_),
    .Y(_04547_));
 sg13g2_nor2_2 _12541_ (.A(_04504_),
    .B(_04547_),
    .Y(_04548_));
 sg13g2_nor2b_1 _12542_ (.A(_04548_),
    .B_N(net319),
    .Y(_04549_));
 sg13g2_o21ai_1 _12543_ (.B1(net58),
    .Y(_04550_),
    .A1(_04546_),
    .A2(_04549_));
 sg13g2_nand2_1 _12544_ (.Y(_04551_),
    .A(_04492_),
    .B(_04550_));
 sg13g2_nor4_1 _12545_ (.A(net314),
    .B(net55),
    .C(_04546_),
    .D(_04549_),
    .Y(_04552_));
 sg13g2_a22oi_1 _12546_ (.Y(_04554_),
    .B1(net104),
    .B2(net315),
    .A2(net76),
    .A1(\i_coord.l_xl.data_out[10] ));
 sg13g2_nand2b_1 _12547_ (.Y(_04555_),
    .B(_04554_),
    .A_N(_04552_));
 sg13g2_buf_1 _12548_ (.A(_04492_),
    .X(_04556_));
 sg13g2_buf_1 _12549_ (.A(_03837_),
    .X(_04557_));
 sg13g2_buf_1 _12550_ (.A(net139),
    .X(_04558_));
 sg13g2_a221oi_1 _12551_ (.B2(net75),
    .C1(net118),
    .B1(_04555_),
    .A1(net314),
    .Y(_04559_),
    .A2(_04551_));
 sg13g2_buf_1 _12552_ (.A(net141),
    .X(_04560_));
 sg13g2_buf_1 _12553_ (.A(_04432_),
    .X(_04561_));
 sg13g2_o21ai_1 _12554_ (.B1(net42),
    .Y(_04562_),
    .A1(net314),
    .A2(net117));
 sg13g2_o21ai_1 _12555_ (.B1(_04554_),
    .Y(_00178_),
    .A1(_04559_),
    .A2(_04562_));
 sg13g2_a21oi_1 _12556_ (.A1(_04503_),
    .A2(_04547_),
    .Y(_04564_),
    .B1(net319));
 sg13g2_o21ai_1 _12557_ (.B1(net319),
    .Y(_04565_),
    .A1(_04503_),
    .A2(_04547_));
 sg13g2_o21ai_1 _12558_ (.B1(_04565_),
    .Y(_04566_),
    .A1(_04505_),
    .A2(_04564_));
 sg13g2_buf_1 _12559_ (.A(_04566_),
    .X(_04567_));
 sg13g2_xnor2_1 _12560_ (.Y(_04568_),
    .A(net319),
    .B(_04567_));
 sg13g2_buf_1 _12561_ (.A(net82),
    .X(_04569_));
 sg13g2_a21oi_1 _12562_ (.A1(net59),
    .A2(_04568_),
    .Y(_04570_),
    .B1(net74));
 sg13g2_buf_2 _12563_ (.A(\i_coord.x0[-2] ),
    .X(_04571_));
 sg13g2_nor2b_1 _12564_ (.A(_04570_),
    .B_N(_04571_),
    .Y(_04572_));
 sg13g2_buf_1 _12565_ (.A(net82),
    .X(_04573_));
 sg13g2_nor3_1 _12566_ (.A(_04571_),
    .B(net55),
    .C(_04568_),
    .Y(_04575_));
 sg13g2_buf_1 _12567_ (.A(_04478_),
    .X(_04576_));
 sg13g2_buf_1 _12568_ (.A(_04150_),
    .X(_04577_));
 sg13g2_a22oi_1 _12569_ (.Y(_04578_),
    .B1(net101),
    .B2(_04227_),
    .A2(net81),
    .A1(\i_coord.l_xl.data_out[11] ));
 sg13g2_nor2b_1 _12570_ (.A(_04575_),
    .B_N(_04578_),
    .Y(_04579_));
 sg13g2_o21ai_1 _12571_ (.B1(net140),
    .Y(_04580_),
    .A1(net73),
    .A2(_04579_));
 sg13g2_nor2_1 _12572_ (.A(_04572_),
    .B(_04580_),
    .Y(_04581_));
 sg13g2_o21ai_1 _12573_ (.B1(net42),
    .Y(_04582_),
    .A1(_04571_),
    .A2(net117));
 sg13g2_o21ai_1 _12574_ (.B1(_04578_),
    .Y(_00179_),
    .A1(_04581_),
    .A2(_04582_));
 sg13g2_buf_1 _12575_ (.A(\i_coord.x0[-1] ),
    .X(_04583_));
 sg13g2_nor2b_1 _12576_ (.A(net319),
    .B_N(_04571_),
    .Y(_04585_));
 sg13g2_and2_1 _12577_ (.A(net314),
    .B(_04585_),
    .X(_04586_));
 sg13g2_nand2b_1 _12578_ (.Y(_04587_),
    .B(net319),
    .A_N(_04571_));
 sg13g2_buf_1 _12579_ (.A(_04587_),
    .X(_04588_));
 sg13g2_nor2_1 _12580_ (.A(net314),
    .B(_04588_),
    .Y(_04589_));
 sg13g2_a22oi_1 _12581_ (.Y(_04590_),
    .B1(_04589_),
    .B2(_04548_),
    .A2(_04586_),
    .A1(_04545_));
 sg13g2_nor3_1 _12582_ (.A(net312),
    .B(net55),
    .C(_04590_),
    .Y(_04591_));
 sg13g2_a22oi_1 _12583_ (.Y(_04592_),
    .B1(net101),
    .B2(_04238_),
    .A2(net81),
    .A1(\i_coord.l_xl.data_out[12] ));
 sg13g2_nor2b_1 _12584_ (.A(_04591_),
    .B_N(_04592_),
    .Y(_04593_));
 sg13g2_a21oi_1 _12585_ (.A1(_04158_),
    .A2(_04590_),
    .Y(_04594_),
    .B1(net82));
 sg13g2_nand2b_1 _12586_ (.Y(_04596_),
    .B(net312),
    .A_N(_04594_));
 sg13g2_o21ai_1 _12587_ (.B1(_04596_),
    .Y(_04597_),
    .A1(net73),
    .A2(_04593_));
 sg13g2_nor2_1 _12588_ (.A(net118),
    .B(_04597_),
    .Y(_04598_));
 sg13g2_o21ai_1 _12589_ (.B1(net42),
    .Y(_04599_),
    .A1(net312),
    .A2(net117));
 sg13g2_o21ai_1 _12590_ (.B1(_04592_),
    .Y(_00180_),
    .A1(_04598_),
    .A2(_04599_));
 sg13g2_buf_1 _12591_ (.A(_04150_),
    .X(_04600_));
 sg13g2_a22oi_1 _12592_ (.Y(_04601_),
    .B1(net100),
    .B2(_04248_),
    .A2(net83),
    .A1(\i_coord.l_xl.data_out[13] ));
 sg13g2_buf_1 _12593_ (.A(\i_coord.x0[0] ),
    .X(_04602_));
 sg13g2_buf_1 _12594_ (.A(_04492_),
    .X(_04603_));
 sg13g2_and2_1 _12595_ (.A(net312),
    .B(_04585_),
    .X(_04604_));
 sg13g2_buf_1 _12596_ (.A(_04604_),
    .X(_04606_));
 sg13g2_nor3_1 _12597_ (.A(net312),
    .B(_04567_),
    .C(_04588_),
    .Y(_04607_));
 sg13g2_a21o_1 _12598_ (.A2(_04606_),
    .A1(_04567_),
    .B1(_04607_),
    .X(_04608_));
 sg13g2_nand4_1 _12599_ (.B(net72),
    .C(_04608_),
    .A(net311),
    .Y(_04609_),
    .D(_04601_));
 sg13g2_nand2b_1 _12600_ (.Y(_04610_),
    .B(_04601_),
    .A_N(_04608_));
 sg13g2_a21o_1 _12601_ (.A2(_04610_),
    .A1(net72),
    .B1(net311),
    .X(_04611_));
 sg13g2_nand3_1 _12602_ (.B(_04609_),
    .C(_04611_),
    .A(_03841_),
    .Y(_04612_));
 sg13g2_buf_1 _12603_ (.A(net118),
    .X(_04613_));
 sg13g2_nand3_1 _12604_ (.B(net99),
    .C(net49),
    .A(net311),
    .Y(_04614_));
 sg13g2_nand3_1 _12605_ (.B(_04612_),
    .C(_04614_),
    .A(_04601_),
    .Y(_00181_));
 sg13g2_buf_2 _12606_ (.A(\i_coord.x0[1] ),
    .X(_04616_));
 sg13g2_buf_1 _12607_ (.A(net72),
    .X(_04617_));
 sg13g2_nand3_1 _12608_ (.B(_04602_),
    .C(_04606_),
    .A(net314),
    .Y(_04618_));
 sg13g2_nor3_1 _12609_ (.A(_04546_),
    .B(_04548_),
    .C(_04618_),
    .Y(_04619_));
 sg13g2_nor4_1 _12610_ (.A(net314),
    .B(net312),
    .C(_04602_),
    .D(_04588_),
    .Y(_04620_));
 sg13g2_o21ai_1 _12611_ (.B1(_04620_),
    .Y(_04621_),
    .A1(_04546_),
    .A2(_04548_));
 sg13g2_nand2b_1 _12612_ (.Y(_04622_),
    .B(_04621_),
    .A_N(_04619_));
 sg13g2_nand3_1 _12613_ (.B(net65),
    .C(_04622_),
    .A(net141),
    .Y(_04623_));
 sg13g2_xor2_1 _12614_ (.B(_04623_),
    .A(_04616_),
    .X(_04624_));
 sg13g2_a22oi_1 _12615_ (.Y(_04625_),
    .B1(net104),
    .B2(_04253_),
    .A2(net76),
    .A1(\i_coord.l_xl.data_out[14] ));
 sg13g2_o21ai_1 _12616_ (.B1(_04625_),
    .Y(_00182_),
    .A1(_04342_),
    .A2(_04624_));
 sg13g2_buf_1 _12617_ (.A(\i_coord.x0[2] ),
    .X(_04627_));
 sg13g2_or4_1 _12618_ (.A(_04583_),
    .B(\i_coord.x0[0] ),
    .C(_04616_),
    .D(_04588_),
    .X(_04628_));
 sg13g2_nand4_1 _12619_ (.B(_04616_),
    .C(_04567_),
    .A(net311),
    .Y(_04629_),
    .D(_04606_));
 sg13g2_o21ai_1 _12620_ (.B1(_04629_),
    .Y(_04630_),
    .A1(_04567_),
    .A2(_04628_));
 sg13g2_nand3_1 _12621_ (.B(net65),
    .C(_04630_),
    .A(net141),
    .Y(_04631_));
 sg13g2_xor2_1 _12622_ (.B(_04631_),
    .A(_04627_),
    .X(_04632_));
 sg13g2_a22oi_1 _12623_ (.Y(_04633_),
    .B1(_04577_),
    .B2(\i_coord.x_row_start[2] ),
    .A2(net81),
    .A1(\i_coord.l_xl.data_out[15] ));
 sg13g2_o21ai_1 _12624_ (.B1(_04633_),
    .Y(_00183_),
    .A1(_04342_),
    .A2(_04632_));
 sg13g2_xor2_1 _12625_ (.B(_04518_),
    .A(_03919_),
    .X(_04634_));
 sg13g2_nor3_1 _12626_ (.A(_04516_),
    .B(_04495_),
    .C(_04634_),
    .Y(_04636_));
 sg13g2_a21o_1 _12627_ (.A2(_04634_),
    .A1(_04516_),
    .B1(_04636_),
    .X(_04637_));
 sg13g2_a221oi_1 _12628_ (.B2(net59),
    .C1(_04557_),
    .B1(_04637_),
    .A1(_04516_),
    .Y(_04638_),
    .A2(net73));
 sg13g2_nor2_1 _12629_ (.A(_04516_),
    .B(_04482_),
    .Y(_04639_));
 sg13g2_nor4_1 _12630_ (.A(net77),
    .B(_04401_),
    .C(_04638_),
    .D(_04639_),
    .Y(_04640_));
 sg13g2_a21o_1 _12631_ (.A2(_04156_),
    .A1(_04178_),
    .B1(_04640_),
    .X(_00184_));
 sg13g2_xor2_1 _12632_ (.B(_04522_),
    .A(\i_coord.l_xip.data_out[2] ),
    .X(_04641_));
 sg13g2_o21ai_1 _12633_ (.B1(_04492_),
    .Y(_04642_),
    .A1(net55),
    .A2(_04641_));
 sg13g2_nor2b_1 _12634_ (.A(_04515_),
    .B_N(_04641_),
    .Y(_04643_));
 sg13g2_a221oi_1 _12635_ (.B2(_04496_),
    .C1(_04557_),
    .B1(_04643_),
    .A1(_04515_),
    .Y(_04644_),
    .A2(_04642_));
 sg13g2_nor2_1 _12636_ (.A(_04515_),
    .B(_04482_),
    .Y(_04646_));
 sg13g2_nor4_1 _12637_ (.A(net77),
    .B(_04401_),
    .C(_04644_),
    .D(_04646_),
    .Y(_04647_));
 sg13g2_a21o_1 _12638_ (.A2(_04156_),
    .A1(_04175_),
    .B1(_04647_),
    .X(_00185_));
 sg13g2_buf_1 _12639_ (.A(_04158_),
    .X(_04648_));
 sg13g2_xnor2_1 _12640_ (.Y(_04649_),
    .A(\i_coord.l_xip.data_out[3] ),
    .B(_04525_));
 sg13g2_buf_1 _12641_ (.A(net82),
    .X(_04650_));
 sg13g2_a21o_1 _12642_ (.A2(_04649_),
    .A1(net53),
    .B1(net71),
    .X(_04651_));
 sg13g2_nor3_1 _12643_ (.A(_04514_),
    .B(net55),
    .C(_04649_),
    .Y(_04652_));
 sg13g2_a22oi_1 _12644_ (.Y(_04653_),
    .B1(net104),
    .B2(_04174_),
    .A2(net76),
    .A1(\i_coord.l_xl.data_out[3] ));
 sg13g2_nand2b_1 _12645_ (.Y(_04654_),
    .B(_04653_),
    .A_N(_04652_));
 sg13g2_a221oi_1 _12646_ (.B2(net75),
    .C1(net118),
    .B1(_04654_),
    .A1(_04514_),
    .Y(_04656_),
    .A2(_04651_));
 sg13g2_o21ai_1 _12647_ (.B1(net42),
    .Y(_04657_),
    .A1(_04514_),
    .A2(net117));
 sg13g2_o21ai_1 _12648_ (.B1(_04653_),
    .Y(_00186_),
    .A1(_04656_),
    .A2(_04657_));
 sg13g2_xnor2_1 _12649_ (.Y(_04658_),
    .A(\i_coord.l_xip.data_out[4] ),
    .B(_04528_));
 sg13g2_a21oi_1 _12650_ (.A1(net59),
    .A2(_04658_),
    .Y(_04659_),
    .B1(net74));
 sg13g2_nor2b_1 _12651_ (.A(_04659_),
    .B_N(net313),
    .Y(_04660_));
 sg13g2_nor3_1 _12652_ (.A(_04513_),
    .B(net54),
    .C(_04658_),
    .Y(_04661_));
 sg13g2_a22oi_1 _12653_ (.Y(_04662_),
    .B1(net100),
    .B2(_04172_),
    .A2(_04576_),
    .A1(\i_coord.l_xl.data_out[4] ));
 sg13g2_nor2b_1 _12654_ (.A(_04661_),
    .B_N(_04662_),
    .Y(_04663_));
 sg13g2_o21ai_1 _12655_ (.B1(net140),
    .Y(_04664_),
    .A1(net73),
    .A2(_04663_));
 sg13g2_nor2_1 _12656_ (.A(_04660_),
    .B(_04664_),
    .Y(_04666_));
 sg13g2_o21ai_1 _12657_ (.B1(net42),
    .Y(_04667_),
    .A1(_04513_),
    .A2(net117));
 sg13g2_o21ai_1 _12658_ (.B1(_04662_),
    .Y(_00187_),
    .A1(_04666_),
    .A2(_04667_));
 sg13g2_xor2_1 _12659_ (.B(_04532_),
    .A(\i_coord.l_xip.data_out[5] ),
    .X(_04668_));
 sg13g2_a21o_1 _12660_ (.A2(_04668_),
    .A1(net53),
    .B1(net71),
    .X(_04669_));
 sg13g2_nand2_1 _12661_ (.Y(_04670_),
    .A(_04512_),
    .B(net58));
 sg13g2_a22oi_1 _12662_ (.Y(_04671_),
    .B1(_04151_),
    .B2(_04171_),
    .A2(net76),
    .A1(\i_coord.l_xl.data_out[5] ));
 sg13g2_o21ai_1 _12663_ (.B1(_04671_),
    .Y(_04672_),
    .A1(_04668_),
    .A2(_04670_));
 sg13g2_a221oi_1 _12664_ (.B2(net75),
    .C1(net118),
    .B1(_04672_),
    .A1(_04511_),
    .Y(_04673_),
    .A2(_04669_));
 sg13g2_o21ai_1 _12665_ (.B1(net42),
    .Y(_04674_),
    .A1(_04511_),
    .A2(net117));
 sg13g2_o21ai_1 _12666_ (.B1(_04671_),
    .Y(_00188_),
    .A1(_04673_),
    .A2(_04674_));
 sg13g2_inv_1 _12667_ (.Y(_04676_),
    .A(_04510_));
 sg13g2_xnor2_1 _12668_ (.Y(_04677_),
    .A(\i_coord.l_xip.data_out[6] ),
    .B(_04535_));
 sg13g2_a21oi_1 _12669_ (.A1(_04159_),
    .A2(_04677_),
    .Y(_04678_),
    .B1(_04569_));
 sg13g2_nor2_1 _12670_ (.A(_04676_),
    .B(_04678_),
    .Y(_04679_));
 sg13g2_nor3_1 _12671_ (.A(_04510_),
    .B(_04484_),
    .C(_04677_),
    .Y(_04680_));
 sg13g2_a22oi_1 _12672_ (.Y(_04681_),
    .B1(_04600_),
    .B2(_04169_),
    .A2(_04576_),
    .A1(\i_coord.l_xl.data_out[6] ));
 sg13g2_nor2b_1 _12673_ (.A(_04680_),
    .B_N(_04681_),
    .Y(_04682_));
 sg13g2_o21ai_1 _12674_ (.B1(_04483_),
    .Y(_04683_),
    .A1(_04573_),
    .A2(_04682_));
 sg13g2_nor2_1 _12675_ (.A(_04679_),
    .B(_04683_),
    .Y(_04684_));
 sg13g2_o21ai_1 _12676_ (.B1(_04561_),
    .Y(_04686_),
    .A1(_04510_),
    .A2(_04560_));
 sg13g2_o21ai_1 _12677_ (.B1(_04681_),
    .Y(_00189_),
    .A1(_04684_),
    .A2(_04686_));
 sg13g2_xor2_1 _12678_ (.B(_04538_),
    .A(\i_coord.l_xip.data_out[7] ),
    .X(_04687_));
 sg13g2_a21o_1 _12679_ (.A2(_04687_),
    .A1(net53),
    .B1(_04650_),
    .X(_04688_));
 sg13g2_nand2_1 _12680_ (.Y(_04689_),
    .A(_04508_),
    .B(_04321_));
 sg13g2_a22oi_1 _12681_ (.Y(_04690_),
    .B1(_04151_),
    .B2(_04168_),
    .A2(_04480_),
    .A1(\i_coord.l_xl.data_out[7] ));
 sg13g2_o21ai_1 _12682_ (.B1(_04690_),
    .Y(_04691_),
    .A1(_04687_),
    .A2(_04689_));
 sg13g2_a221oi_1 _12683_ (.B2(net75),
    .C1(_04558_),
    .B1(_04691_),
    .A1(_04507_),
    .Y(_04692_),
    .A2(_04688_));
 sg13g2_o21ai_1 _12684_ (.B1(_04561_),
    .Y(_04693_),
    .A1(_04507_),
    .A2(_04560_));
 sg13g2_o21ai_1 _12685_ (.B1(_04690_),
    .Y(_00190_),
    .A1(_04692_),
    .A2(_04693_));
 sg13g2_xnor2_1 _12686_ (.Y(_04695_),
    .A(\i_coord.l_xip.data_out[8] ),
    .B(_04541_));
 sg13g2_a21oi_1 _12687_ (.A1(_04159_),
    .A2(_04695_),
    .Y(_04696_),
    .B1(_04569_));
 sg13g2_nor2b_1 _12688_ (.A(_04696_),
    .B_N(_04506_),
    .Y(_04697_));
 sg13g2_nor3_1 _12689_ (.A(_04506_),
    .B(_04484_),
    .C(_04695_),
    .Y(_04698_));
 sg13g2_a22oi_1 _12690_ (.Y(_04699_),
    .B1(_04600_),
    .B2(_04208_),
    .A2(_04479_),
    .A1(\i_coord.l_xl.data_out[8] ));
 sg13g2_nor2b_1 _12691_ (.A(_04698_),
    .B_N(_04699_),
    .Y(_04700_));
 sg13g2_o21ai_1 _12692_ (.B1(_04483_),
    .Y(_04701_),
    .A1(_04573_),
    .A2(_04700_));
 sg13g2_nor2_1 _12693_ (.A(_04697_),
    .B(_04701_),
    .Y(_04702_));
 sg13g2_buf_1 _12694_ (.A(net141),
    .X(_04703_));
 sg13g2_o21ai_1 _12695_ (.B1(net42),
    .Y(_04704_),
    .A1(_04506_),
    .A2(net116));
 sg13g2_o21ai_1 _12696_ (.B1(_04699_),
    .Y(_00191_),
    .A1(_04702_),
    .A2(_04704_));
 sg13g2_xnor2_1 _12697_ (.Y(_04706_),
    .A(net319),
    .B(_04547_));
 sg13g2_a21o_1 _12698_ (.A2(_04706_),
    .A1(_04648_),
    .B1(net71),
    .X(_04707_));
 sg13g2_nand2_1 _12699_ (.Y(_04708_),
    .A(_04505_),
    .B(_04321_));
 sg13g2_a22oi_1 _12700_ (.Y(_04709_),
    .B1(_04577_),
    .B2(_04167_),
    .A2(_04480_),
    .A1(\i_coord.l_xl.data_out[9] ));
 sg13g2_o21ai_1 _12701_ (.B1(_04709_),
    .Y(_04710_),
    .A1(_04706_),
    .A2(_04708_));
 sg13g2_a221oi_1 _12702_ (.B2(_04556_),
    .C1(_04558_),
    .B1(_04710_),
    .A1(_04504_),
    .Y(_04711_),
    .A2(_04707_));
 sg13g2_o21ai_1 _12703_ (.B1(net42),
    .Y(_04712_),
    .A1(_04504_),
    .A2(_04703_));
 sg13g2_o21ai_1 _12704_ (.B1(_04709_),
    .Y(_00192_),
    .A1(_04711_),
    .A2(_04712_));
 sg13g2_nor2_1 _12705_ (.A(_03736_),
    .B(_03845_),
    .Y(_04713_));
 sg13g2_o21ai_1 _12706_ (.B1(_04420_),
    .Y(_04715_),
    .A1(_03945_),
    .A2(_04713_));
 sg13g2_buf_1 _12707_ (.A(_04715_),
    .X(_04716_));
 sg13g2_buf_8 _12708_ (.A(_04716_),
    .X(_04717_));
 sg13g2_buf_1 _12709_ (.A(net17),
    .X(_04718_));
 sg13g2_buf_1 _12710_ (.A(net140),
    .X(_04719_));
 sg13g2_nor3_1 _12711_ (.A(_03267_),
    .B(_02292_),
    .C(_03285_),
    .Y(_04720_));
 sg13g2_or2_1 _12712_ (.X(_04721_),
    .B(_03285_),
    .A(net60));
 sg13g2_nand2_1 _12713_ (.Y(_04722_),
    .A(_03267_),
    .B(_02292_));
 sg13g2_nand2_1 _12714_ (.Y(_04723_),
    .A(_03240_),
    .B(net143));
 sg13g2_o21ai_1 _12715_ (.B1(_04723_),
    .Y(_04724_),
    .A1(_04722_),
    .A2(_03292_));
 sg13g2_a21oi_1 _12716_ (.A1(net60),
    .A2(_03285_),
    .Y(_04726_),
    .B1(_03278_));
 sg13g2_nand3_1 _12717_ (.B(net60),
    .C(_03285_),
    .A(net143),
    .Y(_04727_));
 sg13g2_o21ai_1 _12718_ (.B1(_04727_),
    .Y(_04728_),
    .A1(_03235_),
    .A2(_04726_));
 sg13g2_nor2b_1 _12719_ (.A(_03269_),
    .B_N(_04728_),
    .Y(_04729_));
 sg13g2_a221oi_1 _12720_ (.B2(_04724_),
    .C1(_04729_),
    .B1(_04721_),
    .A1(_03296_),
    .Y(_04730_),
    .A2(_04720_));
 sg13g2_xor2_1 _12721_ (.B(_04730_),
    .A(_03266_),
    .X(_04731_));
 sg13g2_and2_1 _12722_ (.A(_01369_),
    .B(_01372_),
    .X(_04732_));
 sg13g2_nor3_1 _12723_ (.A(_01373_),
    .B(_04731_),
    .C(_04732_),
    .Y(_04733_));
 sg13g2_or3_1 _12724_ (.A(_01373_),
    .B(_01353_),
    .C(_01354_),
    .X(_04734_));
 sg13g2_and2_1 _12725_ (.A(_01374_),
    .B(_04734_),
    .X(_04735_));
 sg13g2_buf_1 _12726_ (.A(_04735_),
    .X(_04737_));
 sg13g2_nand2b_1 _12727_ (.Y(_04738_),
    .B(_03310_),
    .A_N(_03309_));
 sg13g2_xor2_1 _12728_ (.B(_04738_),
    .A(_03262_),
    .X(_04739_));
 sg13g2_xor2_1 _12729_ (.B(_04739_),
    .A(_04481_),
    .X(_04740_));
 sg13g2_xnor2_1 _12730_ (.Y(_04741_),
    .A(_04737_),
    .B(_04740_));
 sg13g2_xnor2_1 _12731_ (.Y(_04742_),
    .A(_04733_),
    .B(_04741_));
 sg13g2_o21ai_1 _12732_ (.B1(_04500_),
    .Y(_04743_),
    .A1(net115),
    .A2(_04742_));
 sg13g2_nand2_1 _12733_ (.Y(_04744_),
    .A(_01926_),
    .B(net17));
 sg13g2_o21ai_1 _12734_ (.B1(_04744_),
    .Y(_00193_),
    .A1(_04718_),
    .A2(_04743_));
 sg13g2_o21ai_1 _12735_ (.B1(_04506_),
    .Y(_04745_),
    .A1(net21),
    .A2(net19));
 sg13g2_nand2_1 _12736_ (.Y(_04747_),
    .A(net21),
    .B(net19));
 sg13g2_nand2_2 _12737_ (.Y(_04748_),
    .A(_04745_),
    .B(_04747_));
 sg13g2_xnor2_1 _12738_ (.Y(_04749_),
    .A(_04504_),
    .B(_03739_));
 sg13g2_xnor2_1 _12739_ (.Y(_04750_),
    .A(_04508_),
    .B(_03750_));
 sg13g2_buf_1 _12740_ (.A(_04750_),
    .X(_04751_));
 sg13g2_inv_1 _12741_ (.Y(_04752_),
    .A(_03632_));
 sg13g2_nand2_1 _12742_ (.Y(_04753_),
    .A(_03636_),
    .B(_04752_));
 sg13g2_a21oi_1 _12743_ (.A1(_04751_),
    .A2(_04753_),
    .Y(_04754_),
    .B1(_04676_));
 sg13g2_nand2b_1 _12744_ (.Y(_04755_),
    .B(_03632_),
    .A_N(_03636_));
 sg13g2_buf_1 _12745_ (.A(_04755_),
    .X(_04756_));
 sg13g2_nor2b_1 _12746_ (.A(_04751_),
    .B_N(_04756_),
    .Y(_04758_));
 sg13g2_xnor2_1 _12747_ (.Y(_04759_),
    .A(_04512_),
    .B(_03762_));
 sg13g2_buf_1 _12748_ (.A(_04759_),
    .X(_04760_));
 sg13g2_nand2b_1 _12749_ (.Y(_04761_),
    .B(_04737_),
    .A_N(_04739_));
 sg13g2_nor2b_1 _12750_ (.A(_04737_),
    .B_N(_04739_),
    .Y(_04762_));
 sg13g2_a21o_1 _12751_ (.A2(_04761_),
    .A1(_04481_),
    .B1(_04762_),
    .X(_04763_));
 sg13g2_buf_1 _12752_ (.A(_04763_),
    .X(_04764_));
 sg13g2_a21o_1 _12753_ (.A2(_01382_),
    .A1(_01321_),
    .B1(_01320_),
    .X(_04765_));
 sg13g2_mux2_1 _12754_ (.A0(_01318_),
    .A1(_01296_),
    .S(_01378_),
    .X(_04766_));
 sg13g2_a21oi_1 _12755_ (.A1(_01312_),
    .A2(_01314_),
    .Y(_04767_),
    .B1(_04766_));
 sg13g2_nor2_1 _12756_ (.A(_01382_),
    .B(_01379_),
    .Y(_04769_));
 sg13g2_o21ai_1 _12757_ (.B1(_04769_),
    .Y(_04770_),
    .A1(_01320_),
    .A2(_04767_));
 sg13g2_nor2_1 _12758_ (.A(_01320_),
    .B(_01321_),
    .Y(_04771_));
 sg13g2_o21ai_1 _12759_ (.B1(_04771_),
    .Y(_04772_),
    .A1(_01379_),
    .A2(_01383_));
 sg13g2_nand2_1 _12760_ (.Y(_04773_),
    .A(_04770_),
    .B(_04772_));
 sg13g2_a21o_1 _12761_ (.A2(_04765_),
    .A1(_01380_),
    .B1(_04773_),
    .X(_04774_));
 sg13g2_buf_1 _12762_ (.A(_04774_),
    .X(_04775_));
 sg13g2_inv_1 _12763_ (.Y(_04776_),
    .A(_04516_));
 sg13g2_xor2_1 _12764_ (.B(_03312_),
    .A(_03260_),
    .X(_04777_));
 sg13g2_xnor2_1 _12765_ (.Y(_04778_),
    .A(_04776_),
    .B(_04777_));
 sg13g2_xnor2_1 _12766_ (.Y(_04780_),
    .A(_04775_),
    .B(_04778_));
 sg13g2_nor2b_1 _12767_ (.A(_04733_),
    .B_N(_04741_),
    .Y(_04781_));
 sg13g2_a21o_1 _12768_ (.A2(_04780_),
    .A1(_04764_),
    .B1(_04781_),
    .X(_04782_));
 sg13g2_o21ai_1 _12769_ (.B1(_04782_),
    .Y(_04783_),
    .A1(_04764_),
    .A2(_04780_));
 sg13g2_xor2_1 _12770_ (.B(_01384_),
    .A(_01250_),
    .X(_04784_));
 sg13g2_xnor2_1 _12771_ (.Y(_04785_),
    .A(_01310_),
    .B(_04784_));
 sg13g2_nand2_1 _12772_ (.Y(_04786_),
    .A(_03260_),
    .B(_03312_));
 sg13g2_xor2_1 _12773_ (.B(_03320_),
    .A(_03229_),
    .X(_04787_));
 sg13g2_xnor2_1 _12774_ (.Y(_04788_),
    .A(_04786_),
    .B(_04787_));
 sg13g2_xnor2_1 _12775_ (.Y(_04789_),
    .A(_04515_),
    .B(_04788_));
 sg13g2_xnor2_1 _12776_ (.Y(_04791_),
    .A(_04785_),
    .B(_04789_));
 sg13g2_inv_1 _12777_ (.Y(_04792_),
    .A(_04777_));
 sg13g2_and2_1 _12778_ (.A(_04775_),
    .B(_04792_),
    .X(_04793_));
 sg13g2_nand2b_1 _12779_ (.Y(_04794_),
    .B(_04777_),
    .A_N(_04775_));
 sg13g2_o21ai_1 _12780_ (.B1(_04794_),
    .Y(_04795_),
    .A1(_04776_),
    .A2(_04793_));
 sg13g2_buf_1 _12781_ (.A(_04795_),
    .X(_04796_));
 sg13g2_nand2_1 _12782_ (.Y(_04797_),
    .A(_04791_),
    .B(_04796_));
 sg13g2_nor2_1 _12783_ (.A(_04791_),
    .B(_04796_),
    .Y(_04798_));
 sg13g2_a21oi_1 _12784_ (.A1(_04783_),
    .A2(_04797_),
    .Y(_04799_),
    .B1(_04798_));
 sg13g2_nand2_1 _12785_ (.Y(_04800_),
    .A(_04785_),
    .B(_04788_));
 sg13g2_nor2_1 _12786_ (.A(_04785_),
    .B(_04788_),
    .Y(_04802_));
 sg13g2_a21oi_2 _12787_ (.B1(_04802_),
    .Y(_04803_),
    .A2(_04800_),
    .A1(_04515_));
 sg13g2_xnor2_1 _12788_ (.Y(_04804_),
    .A(_03223_),
    .B(_03650_));
 sg13g2_nor2_1 _12789_ (.A(_03649_),
    .B(_04804_),
    .Y(_04805_));
 sg13g2_nand2_1 _12790_ (.Y(_04806_),
    .A(_03649_),
    .B(_04804_));
 sg13g2_nand2b_1 _12791_ (.Y(_04807_),
    .B(_04806_),
    .A_N(_04805_));
 sg13g2_xor2_1 _12792_ (.B(_04807_),
    .A(_04514_),
    .X(_04808_));
 sg13g2_nand2_1 _12793_ (.Y(_04809_),
    .A(_04803_),
    .B(_04808_));
 sg13g2_nor2_1 _12794_ (.A(_04803_),
    .B(_04808_),
    .Y(_04810_));
 sg13g2_a21oi_1 _12795_ (.A1(_04799_),
    .A2(_04809_),
    .Y(_04811_),
    .B1(_04810_));
 sg13g2_a21o_1 _12796_ (.A2(_04806_),
    .A1(_04514_),
    .B1(_04805_),
    .X(_04813_));
 sg13g2_buf_1 _12797_ (.A(_04813_),
    .X(_04814_));
 sg13g2_nor2b_1 _12798_ (.A(_04811_),
    .B_N(_04814_),
    .Y(_04815_));
 sg13g2_nor2b_1 _12799_ (.A(_04814_),
    .B_N(_04811_),
    .Y(_04816_));
 sg13g2_or2_1 _12800_ (.X(_04817_),
    .B(_04760_),
    .A(_03755_));
 sg13g2_a22oi_1 _12801_ (.Y(_04818_),
    .B1(_04817_),
    .B2(net313),
    .A2(_04760_),
    .A1(_03756_));
 sg13g2_a21o_1 _12802_ (.A2(_03756_),
    .A1(net313),
    .B1(_03755_),
    .X(_04819_));
 sg13g2_o21ai_1 _12803_ (.B1(_04819_),
    .Y(_04820_),
    .A1(_04760_),
    .A2(_04815_));
 sg13g2_o21ai_1 _12804_ (.B1(_04820_),
    .Y(_04821_),
    .A1(_04816_),
    .A2(_04818_));
 sg13g2_a21o_1 _12805_ (.A2(_04815_),
    .A1(_04760_),
    .B1(_04821_),
    .X(_04822_));
 sg13g2_buf_1 _12806_ (.A(_04822_),
    .X(_04824_));
 sg13g2_nand2_1 _12807_ (.Y(_04825_),
    .A(_03642_),
    .B(_03639_));
 sg13g2_o21ai_1 _12808_ (.B1(_04512_),
    .Y(_04826_),
    .A1(_03642_),
    .A2(_03639_));
 sg13g2_nand2_1 _12809_ (.Y(_04827_),
    .A(_04825_),
    .B(_04826_));
 sg13g2_nand2b_1 _12810_ (.Y(_04828_),
    .B(_04827_),
    .A_N(_04824_));
 sg13g2_buf_1 _12811_ (.A(_04828_),
    .X(_04829_));
 sg13g2_o21ai_1 _12812_ (.B1(_04829_),
    .Y(_04830_),
    .A1(_04754_),
    .A2(_04758_));
 sg13g2_nand2b_1 _12813_ (.Y(_04831_),
    .B(_04824_),
    .A_N(_04827_));
 sg13g2_buf_1 _12814_ (.A(_04831_),
    .X(_04832_));
 sg13g2_inv_1 _12815_ (.Y(_04833_),
    .A(_04753_));
 sg13g2_a21oi_1 _12816_ (.A1(_04510_),
    .A2(_04756_),
    .Y(_04835_),
    .B1(_04833_));
 sg13g2_a21o_1 _12817_ (.A2(_04832_),
    .A1(_04751_),
    .B1(_04835_),
    .X(_04836_));
 sg13g2_or2_1 _12818_ (.X(_04837_),
    .B(_04832_),
    .A(_04751_));
 sg13g2_nand3_1 _12819_ (.B(_04836_),
    .C(_04837_),
    .A(_04830_),
    .Y(_04838_));
 sg13g2_buf_1 _12820_ (.A(_04838_),
    .X(_04839_));
 sg13g2_xnor2_1 _12821_ (.Y(_04840_),
    .A(_04506_),
    .B(_03622_));
 sg13g2_xnor2_1 _12822_ (.Y(_04841_),
    .A(_03626_),
    .B(_04840_));
 sg13g2_a21oi_1 _12823_ (.A1(_03628_),
    .A2(_03629_),
    .Y(_04842_),
    .B1(_04507_));
 sg13g2_a21oi_2 _12824_ (.B1(_04842_),
    .Y(_04843_),
    .A2(_03630_),
    .A1(_03749_));
 sg13g2_o21ai_1 _12825_ (.B1(_04843_),
    .Y(_04844_),
    .A1(_04839_),
    .A2(_04841_));
 sg13g2_nand2_1 _12826_ (.Y(_04846_),
    .A(_04839_),
    .B(_04841_));
 sg13g2_nand2_1 _12827_ (.Y(_04847_),
    .A(_04844_),
    .B(_04846_));
 sg13g2_a21o_1 _12828_ (.A2(_04749_),
    .A1(_04748_),
    .B1(_04847_),
    .X(_04848_));
 sg13g2_o21ai_1 _12829_ (.B1(_04848_),
    .Y(_04849_),
    .A1(_04748_),
    .A2(_04749_));
 sg13g2_o21ai_1 _12830_ (.B1(_04505_),
    .Y(_04850_),
    .A1(_03612_),
    .A2(_03614_));
 sg13g2_nand2_1 _12831_ (.Y(_04851_),
    .A(_03612_),
    .B(_03614_));
 sg13g2_nand2_1 _12832_ (.Y(_04852_),
    .A(_04850_),
    .B(_04851_));
 sg13g2_inv_1 _12833_ (.Y(_04853_),
    .A(\i_coord.x0[-3] ));
 sg13g2_nand2_1 _12834_ (.Y(_04854_),
    .A(_03605_),
    .B(_03695_));
 sg13g2_xnor2_1 _12835_ (.Y(_04855_),
    .A(_04853_),
    .B(_04854_));
 sg13g2_xor2_1 _12836_ (.B(_04855_),
    .A(_04852_),
    .X(_04857_));
 sg13g2_xnor2_1 _12837_ (.Y(_04858_),
    .A(_04849_),
    .B(_04857_));
 sg13g2_a21oi_1 _12838_ (.A1(net99),
    .A2(_04858_),
    .Y(_04859_),
    .B1(_04559_));
 sg13g2_mux2_1 _12839_ (.A0(_04859_),
    .A1(net152),
    .S(net14),
    .X(_00194_));
 sg13g2_inv_1 _12840_ (.Y(_04860_),
    .A(_04855_));
 sg13g2_o21ai_1 _12841_ (.B1(_04841_),
    .Y(_04861_),
    .A1(_04843_),
    .A2(_04839_));
 sg13g2_nand2_1 _12842_ (.Y(_04862_),
    .A(_04843_),
    .B(_04839_));
 sg13g2_inv_1 _12843_ (.Y(_04863_),
    .A(_04749_));
 sg13g2_a21oi_1 _12844_ (.A1(_04861_),
    .A2(_04862_),
    .Y(_04864_),
    .B1(_04863_));
 sg13g2_nand3_1 _12845_ (.B(_04846_),
    .C(_04863_),
    .A(_04844_),
    .Y(_04865_));
 sg13g2_o21ai_1 _12846_ (.B1(_04865_),
    .Y(_04867_),
    .A1(_04748_),
    .A2(_04864_));
 sg13g2_a21o_1 _12847_ (.A2(_04867_),
    .A1(_04860_),
    .B1(_04852_),
    .X(_04868_));
 sg13g2_nand2b_1 _12848_ (.Y(_04869_),
    .B(_04855_),
    .A_N(_04867_));
 sg13g2_nand2_1 _12849_ (.Y(_04870_),
    .A(_04868_),
    .B(_04869_));
 sg13g2_a21oi_1 _12850_ (.A1(net314),
    .A2(_03771_),
    .Y(_04871_),
    .B1(_03772_));
 sg13g2_xor2_1 _12851_ (.B(_03765_),
    .A(_04571_),
    .X(_04872_));
 sg13g2_xnor2_1 _12852_ (.Y(_04873_),
    .A(_04871_),
    .B(_04872_));
 sg13g2_xnor2_1 _12853_ (.Y(_04874_),
    .A(_04870_),
    .B(_04873_));
 sg13g2_a21oi_1 _12854_ (.A1(net99),
    .A2(_04874_),
    .Y(_04875_),
    .B1(_04581_));
 sg13g2_buf_2 _12855_ (.A(_04716_),
    .X(_04876_));
 sg13g2_mux2_1 _12856_ (.A0(_04875_),
    .A1(_02008_),
    .S(_04876_),
    .X(_00195_));
 sg13g2_nand2b_1 _12857_ (.Y(_04878_),
    .B(_04872_),
    .A_N(_04871_));
 sg13g2_nand3_1 _12858_ (.B(_04869_),
    .C(_04878_),
    .A(_04868_),
    .Y(_04879_));
 sg13g2_nand2b_1 _12859_ (.Y(_04880_),
    .B(_04871_),
    .A_N(_04872_));
 sg13g2_nand2_1 _12860_ (.Y(_04881_),
    .A(_04879_),
    .B(_04880_));
 sg13g2_xor2_1 _12861_ (.B(_03768_),
    .A(net312),
    .X(_04882_));
 sg13g2_nand2_1 _12862_ (.Y(_04883_),
    .A(_03578_),
    .B(_03581_));
 sg13g2_nand2_1 _12863_ (.Y(_04884_),
    .A(_04571_),
    .B(_04883_));
 sg13g2_o21ai_1 _12864_ (.B1(_04884_),
    .Y(_04885_),
    .A1(_03578_),
    .A2(_03581_));
 sg13g2_buf_1 _12865_ (.A(_04885_),
    .X(_04886_));
 sg13g2_nor2_1 _12866_ (.A(_04882_),
    .B(_04886_),
    .Y(_04888_));
 sg13g2_nand2_1 _12867_ (.Y(_04889_),
    .A(_04882_),
    .B(_04886_));
 sg13g2_nand2b_1 _12868_ (.Y(_04890_),
    .B(_04889_),
    .A_N(_04888_));
 sg13g2_xnor2_1 _12869_ (.Y(_04891_),
    .A(_04881_),
    .B(_04890_));
 sg13g2_a21oi_1 _12870_ (.A1(_04613_),
    .A2(_04891_),
    .Y(_04892_),
    .B1(_04598_));
 sg13g2_mux2_1 _12871_ (.A0(_04892_),
    .A1(_02032_),
    .S(net16),
    .X(_00196_));
 sg13g2_a22oi_1 _12872_ (.Y(_04893_),
    .B1(_04882_),
    .B2(_04886_),
    .A2(_04880_),
    .A1(_04879_));
 sg13g2_nor2_1 _12873_ (.A(_04888_),
    .B(_04893_),
    .Y(_04894_));
 sg13g2_xor2_1 _12874_ (.B(_03785_),
    .A(net311),
    .X(_04895_));
 sg13g2_nor2_1 _12875_ (.A(_03707_),
    .B(_03678_),
    .Y(_04896_));
 sg13g2_a21oi_1 _12876_ (.A1(net312),
    .A2(_03793_),
    .Y(_04898_),
    .B1(_04896_));
 sg13g2_buf_1 _12877_ (.A(_04898_),
    .X(_04899_));
 sg13g2_xor2_1 _12878_ (.B(_04899_),
    .A(_04895_),
    .X(_04900_));
 sg13g2_xnor2_1 _12879_ (.Y(_04901_),
    .A(_04894_),
    .B(_04900_));
 sg13g2_nand3_1 _12880_ (.B(net53),
    .C(_04713_),
    .A(_03837_),
    .Y(_04902_));
 sg13g2_buf_1 _12881_ (.A(_04902_),
    .X(_04903_));
 sg13g2_nand4_1 _12882_ (.B(net49),
    .C(_04609_),
    .A(net141),
    .Y(_04904_),
    .D(_04611_));
 sg13g2_o21ai_1 _12883_ (.B1(_04904_),
    .Y(_04905_),
    .A1(_04901_),
    .A2(_04903_));
 sg13g2_a21o_1 _12884_ (.A2(net14),
    .A1(_02054_),
    .B1(_04905_),
    .X(_00197_));
 sg13g2_nand4_1 _12885_ (.B(_04617_),
    .C(_04622_),
    .A(_04616_),
    .Y(_04906_),
    .D(_04625_));
 sg13g2_nand2b_1 _12886_ (.Y(_04908_),
    .B(_04625_),
    .A_N(_04622_));
 sg13g2_a21o_1 _12887_ (.A2(_04908_),
    .A1(_04617_),
    .B1(_04616_),
    .X(_04909_));
 sg13g2_nand4_1 _12888_ (.B(_04161_),
    .C(_04906_),
    .A(net117),
    .Y(_04910_),
    .D(_04909_));
 sg13g2_inv_1 _12889_ (.Y(_04911_),
    .A(_04903_));
 sg13g2_xnor2_1 _12890_ (.Y(_04912_),
    .A(_04616_),
    .B(_03807_));
 sg13g2_nor2_1 _12891_ (.A(net311),
    .B(_03782_),
    .Y(_04913_));
 sg13g2_nor2_1 _12892_ (.A(_03783_),
    .B(_04913_),
    .Y(_04914_));
 sg13g2_xnor2_1 _12893_ (.Y(_04915_),
    .A(_04912_),
    .B(_04914_));
 sg13g2_nand2_1 _12894_ (.Y(_04916_),
    .A(_04895_),
    .B(_04899_));
 sg13g2_o21ai_1 _12895_ (.B1(_04889_),
    .Y(_04917_),
    .A1(_04881_),
    .A2(_04888_));
 sg13g2_nor2_1 _12896_ (.A(_04895_),
    .B(_04899_),
    .Y(_04919_));
 sg13g2_a21oi_1 _12897_ (.A1(_04916_),
    .A2(_04917_),
    .Y(_04920_),
    .B1(_04919_));
 sg13g2_xnor2_1 _12898_ (.Y(_04921_),
    .A(_04915_),
    .B(_04920_));
 sg13g2_a22oi_1 _12899_ (.Y(_04922_),
    .B1(_04911_),
    .B2(_04921_),
    .A2(net17),
    .A1(net121));
 sg13g2_nand2_1 _12900_ (.Y(_00198_),
    .A(_04910_),
    .B(_04922_));
 sg13g2_and4_1 _12901_ (.A(_04627_),
    .B(_04603_),
    .C(_04630_),
    .D(_04633_),
    .X(_04923_));
 sg13g2_nand2b_1 _12902_ (.Y(_04924_),
    .B(_04633_),
    .A_N(_04630_));
 sg13g2_a21oi_1 _12903_ (.A1(net72),
    .A2(_04924_),
    .Y(_04925_),
    .B1(_04627_));
 sg13g2_nor3_1 _12904_ (.A(_04439_),
    .B(_04923_),
    .C(_04925_),
    .Y(_04926_));
 sg13g2_nor2_1 _12905_ (.A(_04911_),
    .B(_04926_),
    .Y(_04927_));
 sg13g2_nand2_1 _12906_ (.Y(_04929_),
    .A(net311),
    .B(_03782_));
 sg13g2_nand2_1 _12907_ (.Y(_04930_),
    .A(_04899_),
    .B(_04929_));
 sg13g2_xor2_1 _12908_ (.B(_03807_),
    .A(_04616_),
    .X(_04931_));
 sg13g2_nor2b_1 _12909_ (.A(_04899_),
    .B_N(_03782_),
    .Y(_04932_));
 sg13g2_o21ai_1 _12910_ (.B1(net311),
    .Y(_04933_),
    .A1(_04931_),
    .A2(_04932_));
 sg13g2_o21ai_1 _12911_ (.B1(_04933_),
    .Y(_04934_),
    .A1(_03783_),
    .A2(_04912_));
 sg13g2_a21o_1 _12912_ (.A2(_04930_),
    .A1(_04894_),
    .B1(_04934_),
    .X(_04935_));
 sg13g2_o21ai_1 _12913_ (.B1(_04899_),
    .Y(_04936_),
    .A1(_04888_),
    .A2(_04893_));
 sg13g2_a21o_1 _12914_ (.A2(_04936_),
    .A1(_04931_),
    .B1(_04914_),
    .X(_04937_));
 sg13g2_inv_1 _12915_ (.Y(_04938_),
    .A(_03547_));
 sg13g2_o21ai_1 _12916_ (.B1(_04616_),
    .Y(_04940_),
    .A1(_03547_),
    .A2(_03688_));
 sg13g2_o21ai_1 _12917_ (.B1(_04940_),
    .Y(_04941_),
    .A1(_04938_),
    .A2(_03551_));
 sg13g2_xor2_1 _12918_ (.B(_04941_),
    .A(_03814_),
    .X(_04942_));
 sg13g2_xnor2_1 _12919_ (.Y(_04943_),
    .A(_04627_),
    .B(_04942_));
 sg13g2_a21o_1 _12920_ (.A2(_04937_),
    .A1(_04935_),
    .B1(_04943_),
    .X(_04944_));
 sg13g2_nand3_1 _12921_ (.B(_04937_),
    .C(_04943_),
    .A(_04935_),
    .Y(_04945_));
 sg13g2_a21oi_1 _12922_ (.A1(_04944_),
    .A2(_04945_),
    .Y(_04946_),
    .B1(net117));
 sg13g2_nand2_1 _12923_ (.Y(_04947_),
    .A(_02059_),
    .B(net17));
 sg13g2_o21ai_1 _12924_ (.B1(_04947_),
    .Y(_00199_),
    .A1(_04927_),
    .A2(_04946_));
 sg13g2_or2_1 _12925_ (.X(_04948_),
    .B(_04764_),
    .A(_04781_));
 sg13g2_inv_1 _12926_ (.Y(_04950_),
    .A(_04948_));
 sg13g2_and2_1 _12927_ (.A(_04781_),
    .B(_04764_),
    .X(_04951_));
 sg13g2_nor2_1 _12928_ (.A(_04950_),
    .B(_04951_),
    .Y(_04952_));
 sg13g2_xnor2_1 _12929_ (.Y(_04953_),
    .A(_04780_),
    .B(_04952_));
 sg13g2_a21oi_1 _12930_ (.A1(_04613_),
    .A2(_04953_),
    .Y(_04954_),
    .B1(_04638_));
 sg13g2_buf_1 _12931_ (.A(_01764_),
    .X(_04955_));
 sg13g2_mux2_1 _12932_ (.A0(_04954_),
    .A1(_04955_),
    .S(net16),
    .X(_00200_));
 sg13g2_buf_1 _12933_ (.A(net118),
    .X(_04956_));
 sg13g2_xnor2_1 _12934_ (.Y(_04957_),
    .A(_04791_),
    .B(_04796_));
 sg13g2_xnor2_1 _12935_ (.Y(_04958_),
    .A(_04783_),
    .B(_04957_));
 sg13g2_a21oi_1 _12936_ (.A1(net98),
    .A2(_04958_),
    .Y(_04960_),
    .B1(_04644_));
 sg13g2_buf_1 _12937_ (.A(net187),
    .X(_04961_));
 sg13g2_mux2_1 _12938_ (.A0(_04960_),
    .A1(net137),
    .S(net16),
    .X(_00201_));
 sg13g2_xor2_1 _12939_ (.B(_04808_),
    .A(_04803_),
    .X(_04962_));
 sg13g2_xnor2_1 _12940_ (.Y(_04963_),
    .A(_04799_),
    .B(_04962_));
 sg13g2_a21oi_1 _12941_ (.A1(_04956_),
    .A2(_04963_),
    .Y(_04964_),
    .B1(_04656_));
 sg13g2_buf_1 _12942_ (.A(net323),
    .X(_04965_));
 sg13g2_mux2_1 _12943_ (.A0(_04964_),
    .A1(net271),
    .S(net16),
    .X(_00202_));
 sg13g2_xnor2_1 _12944_ (.Y(_04966_),
    .A(_03757_),
    .B(_04814_));
 sg13g2_xnor2_1 _12945_ (.Y(_04967_),
    .A(net313),
    .B(_04966_));
 sg13g2_xnor2_1 _12946_ (.Y(_04969_),
    .A(_04811_),
    .B(_04967_));
 sg13g2_a21oi_1 _12947_ (.A1(net98),
    .A2(_04969_),
    .Y(_04970_),
    .B1(_04666_));
 sg13g2_buf_1 _12948_ (.A(net174),
    .X(_04971_));
 sg13g2_mux2_1 _12949_ (.A0(_04970_),
    .A1(net136),
    .S(net16),
    .X(_00203_));
 sg13g2_inv_1 _12950_ (.Y(_04972_),
    .A(_03756_));
 sg13g2_inv_1 _12951_ (.Y(_04973_),
    .A(_04815_));
 sg13g2_o21ai_1 _12952_ (.B1(_04973_),
    .Y(_04974_),
    .A1(net25),
    .A2(_04816_));
 sg13g2_nor2_1 _12953_ (.A(net25),
    .B(_04973_),
    .Y(_04975_));
 sg13g2_a21oi_1 _12954_ (.A1(_03655_),
    .A2(_04974_),
    .Y(_04976_),
    .B1(_04975_));
 sg13g2_nand2_1 _12955_ (.Y(_04977_),
    .A(net25),
    .B(_04816_));
 sg13g2_o21ai_1 _12956_ (.B1(_04977_),
    .Y(_04979_),
    .A1(_03655_),
    .A2(_04974_));
 sg13g2_nor2_1 _12957_ (.A(net313),
    .B(_04979_),
    .Y(_04980_));
 sg13g2_a21oi_1 _12958_ (.A1(net313),
    .A2(_04976_),
    .Y(_04981_),
    .B1(_04980_));
 sg13g2_a221oi_1 _12959_ (.B2(_03755_),
    .C1(_04981_),
    .B1(_04815_),
    .A1(_04972_),
    .Y(_04982_),
    .A2(_04816_));
 sg13g2_xnor2_1 _12960_ (.Y(_04983_),
    .A(_04760_),
    .B(_04982_));
 sg13g2_a21oi_1 _12961_ (.A1(net98),
    .A2(_04983_),
    .Y(_04984_),
    .B1(_04673_));
 sg13g2_mux2_1 _12962_ (.A0(_04984_),
    .A1(net170),
    .S(net16),
    .X(_00204_));
 sg13g2_nand2_1 _12963_ (.Y(_04985_),
    .A(_04753_),
    .B(_04756_));
 sg13g2_xor2_1 _12964_ (.B(_04985_),
    .A(_04827_),
    .X(_04986_));
 sg13g2_xnor2_1 _12965_ (.Y(_04987_),
    .A(_04676_),
    .B(_04986_));
 sg13g2_xnor2_1 _12966_ (.Y(_04989_),
    .A(_04824_),
    .B(_04987_));
 sg13g2_a21oi_1 _12967_ (.A1(net98),
    .A2(_04989_),
    .Y(_04990_),
    .B1(_04684_));
 sg13g2_mux2_1 _12968_ (.A0(_04990_),
    .A1(net145),
    .S(net16),
    .X(_00205_));
 sg13g2_inv_1 _12969_ (.Y(_04991_),
    .A(_04832_));
 sg13g2_nand2_1 _12970_ (.Y(_04992_),
    .A(_03636_),
    .B(_04829_));
 sg13g2_nand3_1 _12971_ (.B(_04832_),
    .C(_04992_),
    .A(_03632_),
    .Y(_04993_));
 sg13g2_o21ai_1 _12972_ (.B1(_04993_),
    .Y(_04994_),
    .A1(_03636_),
    .A2(_04829_));
 sg13g2_nand2b_1 _12973_ (.Y(_04995_),
    .B(_04676_),
    .A_N(_04994_));
 sg13g2_nand2_1 _12974_ (.Y(_04996_),
    .A(_04832_),
    .B(_04992_));
 sg13g2_a22oi_1 _12975_ (.Y(_04997_),
    .B1(_04996_),
    .B2(_04752_),
    .A2(_04991_),
    .A1(_03636_));
 sg13g2_nand2_1 _12976_ (.Y(_04999_),
    .A(_04510_),
    .B(_04997_));
 sg13g2_nor2_1 _12977_ (.A(_04829_),
    .B(_04756_),
    .Y(_05000_));
 sg13g2_a221oi_1 _12978_ (.B2(_04999_),
    .C1(_05000_),
    .B1(_04995_),
    .A1(_04833_),
    .Y(_05001_),
    .A2(_04991_));
 sg13g2_xor2_1 _12979_ (.B(_05001_),
    .A(_04751_),
    .X(_05002_));
 sg13g2_a21oi_1 _12980_ (.A1(net98),
    .A2(_05002_),
    .Y(_05003_),
    .B1(_04692_));
 sg13g2_buf_1 _12981_ (.A(net146),
    .X(_05004_));
 sg13g2_mux2_1 _12982_ (.A0(_05003_),
    .A1(_05004_),
    .S(_04876_),
    .X(_00206_));
 sg13g2_xor2_1 _12983_ (.B(_04841_),
    .A(_04843_),
    .X(_05005_));
 sg13g2_xnor2_1 _12984_ (.Y(_05006_),
    .A(_04839_),
    .B(_05005_));
 sg13g2_a21oi_1 _12985_ (.A1(net98),
    .A2(_05006_),
    .Y(_05007_),
    .B1(_04702_));
 sg13g2_mux2_1 _12986_ (.A0(_05007_),
    .A1(net144),
    .S(net16),
    .X(_00207_));
 sg13g2_xor2_1 _12987_ (.B(_04749_),
    .A(_04748_),
    .X(_05009_));
 sg13g2_xnor2_1 _12988_ (.Y(_05010_),
    .A(_04847_),
    .B(_05009_));
 sg13g2_a21oi_1 _12989_ (.A1(net98),
    .A2(_05010_),
    .Y(_05011_),
    .B1(_04711_));
 sg13g2_buf_2 _12990_ (.A(_04716_),
    .X(_05012_));
 sg13g2_mux2_1 _12991_ (.A0(_05011_),
    .A1(net151),
    .S(net15),
    .X(_00208_));
 sg13g2_o21ai_1 _12992_ (.B1(_04492_),
    .Y(_05013_),
    .A1(_04028_),
    .A2(net55));
 sg13g2_nand2b_1 _12993_ (.Y(_05014_),
    .B(_04028_),
    .A_N(_04046_));
 sg13g2_a22oi_1 _12994_ (.Y(_05015_),
    .B1(net101),
    .B2(_04331_),
    .A2(net76),
    .A1(\i_coord.l_yt.data_out[0] ));
 sg13g2_o21ai_1 _12995_ (.B1(_05015_),
    .Y(_05016_),
    .A1(_04341_),
    .A2(_05014_));
 sg13g2_a221oi_1 _12996_ (.B2(_04556_),
    .C1(net118),
    .B1(_05016_),
    .A1(_04046_),
    .Y(_05018_),
    .A2(_05013_));
 sg13g2_buf_1 _12997_ (.A(_04432_),
    .X(_05019_));
 sg13g2_o21ai_1 _12998_ (.B1(net41),
    .Y(_05020_),
    .A1(_04046_),
    .A2(_04703_));
 sg13g2_o21ai_1 _12999_ (.B1(_05015_),
    .Y(_00209_),
    .A1(_05018_),
    .A2(_05020_));
 sg13g2_inv_1 _13000_ (.Y(_05021_),
    .A(_04076_));
 sg13g2_inv_1 _13001_ (.Y(_05022_),
    .A(\i_coord.l_yip.data_out[6] ));
 sg13g2_inv_1 _13002_ (.Y(_05023_),
    .A(\i_coord.l_yip.data_out[3] ));
 sg13g2_nor2_1 _13003_ (.A(_04032_),
    .B(_04105_),
    .Y(_05024_));
 sg13g2_nand2_1 _13004_ (.Y(_05025_),
    .A(_04028_),
    .B(_04046_));
 sg13g2_nand2_1 _13005_ (.Y(_05026_),
    .A(_04032_),
    .B(_04105_));
 sg13g2_o21ai_1 _13006_ (.B1(_05026_),
    .Y(_05028_),
    .A1(_05024_),
    .A2(_05025_));
 sg13g2_a21o_1 _13007_ (.A2(_04033_),
    .A1(_04108_),
    .B1(_05028_),
    .X(_05029_));
 sg13g2_o21ai_1 _13008_ (.B1(_05029_),
    .Y(_05030_),
    .A1(_04108_),
    .A2(_04033_));
 sg13g2_buf_1 _13009_ (.A(_05030_),
    .X(_05031_));
 sg13g2_nand2_1 _13010_ (.Y(_05032_),
    .A(_05023_),
    .B(_05031_));
 sg13g2_nand2_1 _13011_ (.Y(_05033_),
    .A(_04112_),
    .B(_05032_));
 sg13g2_o21ai_1 _13012_ (.B1(_05033_),
    .Y(_05034_),
    .A1(_05023_),
    .A2(_05031_));
 sg13g2_buf_1 _13013_ (.A(_05034_),
    .X(_05035_));
 sg13g2_nor2_1 _13014_ (.A(_04035_),
    .B(_05035_),
    .Y(_05036_));
 sg13g2_a21oi_1 _13015_ (.A1(_04035_),
    .A2(_05035_),
    .Y(_05037_),
    .B1(_04063_));
 sg13g2_nor2_1 _13016_ (.A(_05036_),
    .B(_05037_),
    .Y(_05039_));
 sg13g2_a21o_1 _13017_ (.A2(_05039_),
    .A1(_04036_),
    .B1(net317),
    .X(_05040_));
 sg13g2_o21ai_1 _13018_ (.B1(_05040_),
    .Y(_05041_),
    .A1(_04036_),
    .A2(_05039_));
 sg13g2_buf_1 _13019_ (.A(_05041_),
    .X(_05042_));
 sg13g2_inv_1 _13020_ (.Y(_05043_),
    .A(_05042_));
 sg13g2_a21oi_1 _13021_ (.A1(\i_coord.l_yip.data_out[6] ),
    .A2(_05043_),
    .Y(_05044_),
    .B1(_04064_));
 sg13g2_a21oi_1 _13022_ (.A1(_05022_),
    .A2(_05042_),
    .Y(_05045_),
    .B1(_05044_));
 sg13g2_nor2_1 _13023_ (.A(_04037_),
    .B(_05045_),
    .Y(_05046_));
 sg13g2_a21oi_1 _13024_ (.A1(_04037_),
    .A2(_05045_),
    .Y(_05047_),
    .B1(_04059_));
 sg13g2_nor2_1 _13025_ (.A(_05046_),
    .B(_05047_),
    .Y(_05048_));
 sg13g2_nor2_1 _13026_ (.A(_04038_),
    .B(_05048_),
    .Y(_05050_));
 sg13g2_a21oi_1 _13027_ (.A1(_04038_),
    .A2(_05048_),
    .Y(_05051_),
    .B1(_04057_));
 sg13g2_nor2_2 _13028_ (.A(_05050_),
    .B(_05051_),
    .Y(_05052_));
 sg13g2_a21o_1 _13029_ (.A2(_05052_),
    .A1(_04042_),
    .B1(_04058_),
    .X(_05053_));
 sg13g2_o21ai_1 _13030_ (.B1(_05053_),
    .Y(_05054_),
    .A1(_04042_),
    .A2(_05052_));
 sg13g2_buf_1 _13031_ (.A(_05054_),
    .X(_05055_));
 sg13g2_xnor2_1 _13032_ (.Y(_05056_),
    .A(_04043_),
    .B(_05055_));
 sg13g2_a21oi_1 _13033_ (.A1(net59),
    .A2(_05056_),
    .Y(_05057_),
    .B1(net74));
 sg13g2_nor2_1 _13034_ (.A(_05021_),
    .B(_05057_),
    .Y(_05058_));
 sg13g2_nor3_1 _13035_ (.A(_04076_),
    .B(net54),
    .C(_05056_),
    .Y(_05059_));
 sg13g2_a22oi_1 _13036_ (.Y(_05061_),
    .B1(net100),
    .B2(_04340_),
    .A2(net83),
    .A1(\i_coord.l_yt.data_out[10] ));
 sg13g2_nor2b_1 _13037_ (.A(_05059_),
    .B_N(_05061_),
    .Y(_05062_));
 sg13g2_o21ai_1 _13038_ (.B1(net140),
    .Y(_05063_),
    .A1(net73),
    .A2(_05062_));
 sg13g2_nor2_1 _13039_ (.A(_05058_),
    .B(_05063_),
    .Y(_05064_));
 sg13g2_o21ai_1 _13040_ (.B1(net41),
    .Y(_05065_),
    .A1(_04076_),
    .A2(net116));
 sg13g2_o21ai_1 _13041_ (.B1(_05061_),
    .Y(_00210_),
    .A1(_05064_),
    .A2(_05065_));
 sg13g2_nor2_2 _13042_ (.A(_04043_),
    .B(_05053_),
    .Y(_05066_));
 sg13g2_nor2_1 _13043_ (.A(_05021_),
    .B(_04042_),
    .Y(_05067_));
 sg13g2_and2_1 _13044_ (.A(_04058_),
    .B(_05052_),
    .X(_05068_));
 sg13g2_a22oi_1 _13045_ (.Y(_05069_),
    .B1(_05067_),
    .B2(_05068_),
    .A2(_05066_),
    .A1(_05021_));
 sg13g2_a21o_1 _13046_ (.A2(_05069_),
    .A1(net53),
    .B1(net71),
    .X(_05071_));
 sg13g2_nand2b_1 _13047_ (.Y(_05072_),
    .B(net58),
    .A_N(_04083_));
 sg13g2_a22oi_1 _13048_ (.Y(_05073_),
    .B1(net104),
    .B2(_04382_),
    .A2(net76),
    .A1(\i_coord.l_yt.data_out[11] ));
 sg13g2_o21ai_1 _13049_ (.B1(_05073_),
    .Y(_05074_),
    .A1(_05069_),
    .A2(_05072_));
 sg13g2_a221oi_1 _13050_ (.B2(net75),
    .C1(net118),
    .B1(_05074_),
    .A1(_04083_),
    .Y(_05075_),
    .A2(_05071_));
 sg13g2_o21ai_1 _13051_ (.B1(net41),
    .Y(_05076_),
    .A1(_04083_),
    .A2(net116));
 sg13g2_o21ai_1 _13052_ (.B1(_05073_),
    .Y(_00211_),
    .A1(_05075_),
    .A2(_05076_));
 sg13g2_nand2_1 _13053_ (.Y(_05077_),
    .A(_04083_),
    .B(_05067_));
 sg13g2_nor2_1 _13054_ (.A(_05055_),
    .B(_05077_),
    .Y(_05078_));
 sg13g2_a21oi_1 _13055_ (.A1(_04084_),
    .A2(_05066_),
    .Y(_05079_),
    .B1(_05078_));
 sg13g2_a21o_1 _13056_ (.A2(_05079_),
    .A1(net53),
    .B1(net71),
    .X(_05081_));
 sg13g2_nand2b_1 _13057_ (.Y(_05082_),
    .B(net58),
    .A_N(_04091_));
 sg13g2_a22oi_1 _13058_ (.Y(_05083_),
    .B1(net101),
    .B2(_04392_),
    .A2(net81),
    .A1(\i_coord.l_yt.data_out[12] ));
 sg13g2_o21ai_1 _13059_ (.B1(_05083_),
    .Y(_05084_),
    .A1(_05079_),
    .A2(_05082_));
 sg13g2_a221oi_1 _13060_ (.B2(net75),
    .C1(net139),
    .B1(_05084_),
    .A1(_04091_),
    .Y(_05085_),
    .A2(_05081_));
 sg13g2_o21ai_1 _13061_ (.B1(net41),
    .Y(_05086_),
    .A1(_04091_),
    .A2(net116));
 sg13g2_o21ai_1 _13062_ (.B1(_05083_),
    .Y(_00212_),
    .A1(_05085_),
    .A2(_05086_));
 sg13g2_and3_1 _13063_ (.X(_05087_),
    .A(_04083_),
    .B(_04091_),
    .C(_05067_));
 sg13g2_nor3_1 _13064_ (.A(_04076_),
    .B(_04083_),
    .C(_04091_),
    .Y(_05088_));
 sg13g2_a22oi_1 _13065_ (.Y(_05089_),
    .B1(_05088_),
    .B2(_05066_),
    .A2(_05087_),
    .A1(_05068_));
 sg13g2_a21oi_1 _13066_ (.A1(_04158_),
    .A2(_05089_),
    .Y(_05091_),
    .B1(net82));
 sg13g2_inv_1 _13067_ (.Y(_05092_),
    .A(_05091_));
 sg13g2_nand2b_1 _13068_ (.Y(_05093_),
    .B(net58),
    .A_N(_04098_));
 sg13g2_a22oi_1 _13069_ (.Y(_05094_),
    .B1(net101),
    .B2(_04407_),
    .A2(net81),
    .A1(\i_coord.l_yt.data_out[13] ));
 sg13g2_o21ai_1 _13070_ (.B1(_05094_),
    .Y(_05095_),
    .A1(_05089_),
    .A2(_05093_));
 sg13g2_a221oi_1 _13071_ (.B2(net75),
    .C1(net139),
    .B1(_05095_),
    .A1(_04098_),
    .Y(_05096_),
    .A2(_05092_));
 sg13g2_o21ai_1 _13072_ (.B1(net41),
    .Y(_05097_),
    .A1(_04098_),
    .A2(net116));
 sg13g2_o21ai_1 _13073_ (.B1(_05094_),
    .Y(_00213_),
    .A1(_05096_),
    .A2(_05097_));
 sg13g2_nand2_1 _13074_ (.Y(_05098_),
    .A(_04098_),
    .B(_05087_));
 sg13g2_nand3_1 _13075_ (.B(_04099_),
    .C(_05066_),
    .A(_04084_),
    .Y(_05099_));
 sg13g2_o21ai_1 _13076_ (.B1(_05099_),
    .Y(_05101_),
    .A1(_05055_),
    .A2(_05098_));
 sg13g2_nand3_1 _13077_ (.B(net75),
    .C(_05101_),
    .A(net140),
    .Y(_05102_));
 sg13g2_xor2_1 _13078_ (.B(_05102_),
    .A(_04097_),
    .X(_05103_));
 sg13g2_a22oi_1 _13079_ (.Y(_05104_),
    .B1(net100),
    .B2(\i_coord.y_row_start[1] ),
    .A2(net83),
    .A1(\i_coord.l_yt.data_out[14] ));
 sg13g2_o21ai_1 _13080_ (.B1(_05104_),
    .Y(_00214_),
    .A1(net48),
    .A2(_05103_));
 sg13g2_xor2_1 _13081_ (.B(_05025_),
    .A(_04032_),
    .X(_05105_));
 sg13g2_a21oi_1 _13082_ (.A1(net59),
    .A2(_05105_),
    .Y(_05106_),
    .B1(net74));
 sg13g2_nor2b_1 _13083_ (.A(_05106_),
    .B_N(_04105_),
    .Y(_05107_));
 sg13g2_nor3_1 _13084_ (.A(_04105_),
    .B(net54),
    .C(_05105_),
    .Y(_05108_));
 sg13g2_a22oi_1 _13085_ (.Y(_05109_),
    .B1(net100),
    .B2(_04350_),
    .A2(net83),
    .A1(\i_coord.l_yt.data_out[1] ));
 sg13g2_nor2b_1 _13086_ (.A(_05108_),
    .B_N(_05109_),
    .Y(_05111_));
 sg13g2_o21ai_1 _13087_ (.B1(net140),
    .Y(_05112_),
    .A1(net73),
    .A2(_05111_));
 sg13g2_nor2_1 _13088_ (.A(_05107_),
    .B(_05112_),
    .Y(_05113_));
 sg13g2_o21ai_1 _13089_ (.B1(net41),
    .Y(_05114_),
    .A1(_04105_),
    .A2(net116));
 sg13g2_o21ai_1 _13090_ (.B1(_05109_),
    .Y(_00215_),
    .A1(_05113_),
    .A2(_05114_));
 sg13g2_xnor2_1 _13091_ (.Y(_05115_),
    .A(_04033_),
    .B(_05028_));
 sg13g2_a21oi_1 _13092_ (.A1(net59),
    .A2(_05115_),
    .Y(_05116_),
    .B1(net74));
 sg13g2_nor2b_1 _13093_ (.A(_05116_),
    .B_N(_04108_),
    .Y(_05117_));
 sg13g2_nor3_1 _13094_ (.A(_04108_),
    .B(net54),
    .C(_05115_),
    .Y(_05118_));
 sg13g2_a22oi_1 _13095_ (.Y(_05119_),
    .B1(net100),
    .B2(_04354_),
    .A2(net83),
    .A1(\i_coord.l_yt.data_out[2] ));
 sg13g2_nor2b_1 _13096_ (.A(_05118_),
    .B_N(_05119_),
    .Y(_05121_));
 sg13g2_o21ai_1 _13097_ (.B1(net140),
    .Y(_05122_),
    .A1(net73),
    .A2(_05121_));
 sg13g2_nor2_1 _13098_ (.A(_05117_),
    .B(_05122_),
    .Y(_05123_));
 sg13g2_o21ai_1 _13099_ (.B1(net41),
    .Y(_05124_),
    .A1(_04108_),
    .A2(net116));
 sg13g2_o21ai_1 _13100_ (.B1(_05119_),
    .Y(_00216_),
    .A1(_05123_),
    .A2(_05124_));
 sg13g2_xnor2_1 _13101_ (.Y(_05125_),
    .A(_05023_),
    .B(_05031_));
 sg13g2_a21o_1 _13102_ (.A2(_05125_),
    .A1(_04648_),
    .B1(_04650_),
    .X(_05126_));
 sg13g2_nor3_1 _13103_ (.A(_04112_),
    .B(_04341_),
    .C(_05125_),
    .Y(_05127_));
 sg13g2_a22oi_1 _13104_ (.Y(_05128_),
    .B1(net104),
    .B2(_04349_),
    .A2(net76),
    .A1(\i_coord.l_yt.data_out[3] ));
 sg13g2_nand2b_1 _13105_ (.Y(_05129_),
    .B(_05128_),
    .A_N(_05127_));
 sg13g2_a221oi_1 _13106_ (.B2(net72),
    .C1(net139),
    .B1(_05129_),
    .A1(_04112_),
    .Y(_05131_),
    .A2(_05126_));
 sg13g2_o21ai_1 _13107_ (.B1(net41),
    .Y(_05132_),
    .A1(_04112_),
    .A2(net116));
 sg13g2_o21ai_1 _13108_ (.B1(_05128_),
    .Y(_00217_),
    .A1(_05131_),
    .A2(_05132_));
 sg13g2_xnor2_1 _13109_ (.Y(_05133_),
    .A(_04035_),
    .B(_05035_));
 sg13g2_a21o_1 _13110_ (.A2(_05133_),
    .A1(_04158_),
    .B1(net82),
    .X(_05134_));
 sg13g2_nand2b_1 _13111_ (.Y(_05135_),
    .B(_04420_),
    .A_N(_04063_));
 sg13g2_a22oi_1 _13112_ (.Y(_05136_),
    .B1(net101),
    .B2(_04347_),
    .A2(net81),
    .A1(\i_coord.l_yt.data_out[4] ));
 sg13g2_o21ai_1 _13113_ (.B1(_05136_),
    .Y(_05137_),
    .A1(_05133_),
    .A2(_05135_));
 sg13g2_a221oi_1 _13114_ (.B2(_04603_),
    .C1(net139),
    .B1(_05137_),
    .A1(_04063_),
    .Y(_05138_),
    .A2(_05134_));
 sg13g2_o21ai_1 _13115_ (.B1(_05019_),
    .Y(_05139_),
    .A1(_04063_),
    .A2(net115));
 sg13g2_o21ai_1 _13116_ (.B1(_05136_),
    .Y(_00218_),
    .A1(_05138_),
    .A2(_05139_));
 sg13g2_xnor2_1 _13117_ (.Y(_05141_),
    .A(_04036_),
    .B(_05039_));
 sg13g2_a21oi_1 _13118_ (.A1(net59),
    .A2(_05141_),
    .Y(_05142_),
    .B1(net74));
 sg13g2_nor2b_1 _13119_ (.A(_05142_),
    .B_N(net317),
    .Y(_05143_));
 sg13g2_nor3_1 _13120_ (.A(net317),
    .B(net54),
    .C(_05141_),
    .Y(_05144_));
 sg13g2_a22oi_1 _13121_ (.Y(_05145_),
    .B1(net100),
    .B2(_04346_),
    .A2(net83),
    .A1(\i_coord.l_yt.data_out[5] ));
 sg13g2_nor2b_1 _13122_ (.A(_05144_),
    .B_N(_05145_),
    .Y(_05146_));
 sg13g2_o21ai_1 _13123_ (.B1(_03945_),
    .Y(_05147_),
    .A1(net73),
    .A2(_05146_));
 sg13g2_nor2_1 _13124_ (.A(_05143_),
    .B(_05147_),
    .Y(_05148_));
 sg13g2_o21ai_1 _13125_ (.B1(_05019_),
    .Y(_05149_),
    .A1(_04062_),
    .A2(_04719_));
 sg13g2_o21ai_1 _13126_ (.B1(_05145_),
    .Y(_00219_),
    .A1(_05148_),
    .A2(_05149_));
 sg13g2_xnor2_1 _13127_ (.Y(_05151_),
    .A(_05022_),
    .B(_05042_));
 sg13g2_a21o_1 _13128_ (.A2(_05151_),
    .A1(net53),
    .B1(net71),
    .X(_05152_));
 sg13g2_nand2b_1 _13129_ (.Y(_05153_),
    .B(_04420_),
    .A_N(_04064_));
 sg13g2_a22oi_1 _13130_ (.Y(_05154_),
    .B1(net101),
    .B2(\i_coord.y_row_start[-7] ),
    .A2(net81),
    .A1(\i_coord.l_yt.data_out[6] ));
 sg13g2_o21ai_1 _13131_ (.B1(_05154_),
    .Y(_05155_),
    .A1(_05151_),
    .A2(_05153_));
 sg13g2_a221oi_1 _13132_ (.B2(net72),
    .C1(net139),
    .B1(_05155_),
    .A1(_04064_),
    .Y(_05156_),
    .A2(_05152_));
 sg13g2_o21ai_1 _13133_ (.B1(net47),
    .Y(_05157_),
    .A1(_04064_),
    .A2(net115));
 sg13g2_o21ai_1 _13134_ (.B1(_05154_),
    .Y(_00220_),
    .A1(_05156_),
    .A2(_05157_));
 sg13g2_xnor2_1 _13135_ (.Y(_05158_),
    .A(_04037_),
    .B(_05045_));
 sg13g2_a21oi_1 _13136_ (.A1(net53),
    .A2(_05158_),
    .Y(_05160_),
    .B1(net71));
 sg13g2_nor2_1 _13137_ (.A(_04061_),
    .B(_05160_),
    .Y(_05161_));
 sg13g2_nor3_1 _13138_ (.A(_04059_),
    .B(net54),
    .C(_05158_),
    .Y(_05162_));
 sg13g2_a22oi_1 _13139_ (.Y(_05163_),
    .B1(net100),
    .B2(_04374_),
    .A2(net83),
    .A1(\i_coord.l_yt.data_out[7] ));
 sg13g2_nor2b_1 _13140_ (.A(_05162_),
    .B_N(_05163_),
    .Y(_05164_));
 sg13g2_o21ai_1 _13141_ (.B1(_03945_),
    .Y(_05165_),
    .A1(net74),
    .A2(_05164_));
 sg13g2_nor2_1 _13142_ (.A(_05161_),
    .B(_05165_),
    .Y(_05166_));
 sg13g2_o21ai_1 _13143_ (.B1(net47),
    .Y(_05167_),
    .A1(_04059_),
    .A2(_04719_));
 sg13g2_o21ai_1 _13144_ (.B1(_05163_),
    .Y(_00221_),
    .A1(_05166_),
    .A2(_05167_));
 sg13g2_xnor2_1 _13145_ (.Y(_05168_),
    .A(_04038_),
    .B(_05048_));
 sg13g2_a21o_1 _13146_ (.A2(_05168_),
    .A1(_04158_),
    .B1(net71),
    .X(_05170_));
 sg13g2_nand2_1 _13147_ (.Y(_05171_),
    .A(_04138_),
    .B(net58));
 sg13g2_a22oi_1 _13148_ (.Y(_05172_),
    .B1(net101),
    .B2(_04343_),
    .A2(net81),
    .A1(\i_coord.l_yt.data_out[8] ));
 sg13g2_o21ai_1 _13149_ (.B1(_05172_),
    .Y(_05173_),
    .A1(_05168_),
    .A2(_05171_));
 sg13g2_a221oi_1 _13150_ (.B2(net72),
    .C1(net139),
    .B1(_05173_),
    .A1(_04057_),
    .Y(_05174_),
    .A2(_05170_));
 sg13g2_o21ai_1 _13151_ (.B1(net47),
    .Y(_05175_),
    .A1(_04057_),
    .A2(net115));
 sg13g2_o21ai_1 _13152_ (.B1(_05172_),
    .Y(_00222_),
    .A1(_05174_),
    .A2(_05175_));
 sg13g2_xnor2_1 _13153_ (.Y(_05176_),
    .A(_04042_),
    .B(_05052_));
 sg13g2_a21oi_1 _13154_ (.A1(_04158_),
    .A2(_05176_),
    .Y(_05177_),
    .B1(net82));
 sg13g2_nor2b_1 _13155_ (.A(_05177_),
    .B_N(_04058_),
    .Y(_05178_));
 sg13g2_nor3_1 _13156_ (.A(_04058_),
    .B(_03839_),
    .C(_05176_),
    .Y(_05180_));
 sg13g2_a22oi_1 _13157_ (.Y(_05181_),
    .B1(_04150_),
    .B2(_04344_),
    .A2(net83),
    .A1(\i_coord.l_yt.data_out[9] ));
 sg13g2_nor2b_1 _13158_ (.A(_05180_),
    .B_N(_05181_),
    .Y(_05182_));
 sg13g2_o21ai_1 _13159_ (.B1(_03945_),
    .Y(_05183_),
    .A1(net74),
    .A2(_05182_));
 sg13g2_nor2_1 _13160_ (.A(_05178_),
    .B(_05183_),
    .Y(_05184_));
 sg13g2_o21ai_1 _13161_ (.B1(net47),
    .Y(_05185_),
    .A1(_04058_),
    .A2(net115));
 sg13g2_o21ai_1 _13162_ (.B1(_05181_),
    .Y(_00223_),
    .A1(_05184_),
    .A2(_05185_));
 sg13g2_or2_1 _13163_ (.X(_05186_),
    .B(net147),
    .A(_01267_));
 sg13g2_buf_1 _13164_ (.A(_05186_),
    .X(_05187_));
 sg13g2_buf_1 _13165_ (.A(_00034_),
    .X(_05188_));
 sg13g2_nor3_2 _13166_ (.A(_05188_),
    .B(_05376_),
    .C(_05420_),
    .Y(_05190_));
 sg13g2_nor2_2 _13167_ (.A(net188),
    .B(_07296_),
    .Y(_05191_));
 sg13g2_buf_1 _13168_ (.A(_01538_),
    .X(_05192_));
 sg13g2_nor2_1 _13169_ (.A(net166),
    .B(net160),
    .Y(_05193_));
 sg13g2_xnor2_1 _13170_ (.Y(_05194_),
    .A(_05191_),
    .B(_05193_));
 sg13g2_xnor2_1 _13171_ (.Y(_05195_),
    .A(_05190_),
    .B(_05194_));
 sg13g2_inv_1 _13172_ (.Y(_05196_),
    .A(_05188_));
 sg13g2_nand4_1 _13173_ (.B(_05196_),
    .C(net161),
    .A(net184),
    .Y(_05197_),
    .D(net209));
 sg13g2_buf_1 _13174_ (.A(_05197_),
    .X(_05198_));
 sg13g2_a22oi_1 _13175_ (.Y(_05199_),
    .B1(net209),
    .B2(net184),
    .A2(net161),
    .A1(_05196_));
 sg13g2_a21oi_1 _13176_ (.A1(net166),
    .A2(_05198_),
    .Y(_05201_),
    .B1(_05199_));
 sg13g2_or3_1 _13177_ (.A(net323),
    .B(net166),
    .C(_05199_),
    .X(_05202_));
 sg13g2_o21ai_1 _13178_ (.B1(_05202_),
    .Y(_05203_),
    .A1(_01922_),
    .A2(_05201_));
 sg13g2_nand2_1 _13179_ (.Y(_05204_),
    .A(net323),
    .B(net210));
 sg13g2_nor2b_1 _13180_ (.A(_05198_),
    .B_N(_05204_),
    .Y(_05205_));
 sg13g2_a21o_1 _13181_ (.A2(_05203_),
    .A1(net210),
    .B1(_05205_),
    .X(_05206_));
 sg13g2_xnor2_1 _13182_ (.Y(_05207_),
    .A(_05195_),
    .B(_05206_));
 sg13g2_nand2_1 _13183_ (.Y(_05208_),
    .A(net138),
    .B(net209));
 sg13g2_nand2_1 _13184_ (.Y(_05209_),
    .A(_05196_),
    .B(net161));
 sg13g2_nand2_1 _13185_ (.Y(_05210_),
    .A(net187),
    .B(net210));
 sg13g2_xnor2_1 _13186_ (.Y(_05212_),
    .A(_05209_),
    .B(_05210_));
 sg13g2_xor2_1 _13187_ (.B(_05212_),
    .A(_05208_),
    .X(_05213_));
 sg13g2_nand2_1 _13188_ (.Y(_05214_),
    .A(_01560_),
    .B(_06420_));
 sg13g2_nand4_1 _13189_ (.B(_05196_),
    .C(net209),
    .A(net184),
    .Y(_05215_),
    .D(net210));
 sg13g2_a22oi_1 _13190_ (.Y(_05216_),
    .B1(net210),
    .B2(net184),
    .A2(net209),
    .A1(_05196_));
 sg13g2_a21o_1 _13191_ (.A2(_05215_),
    .A1(_05214_),
    .B1(_05216_),
    .X(_05217_));
 sg13g2_buf_1 _13192_ (.A(_05217_),
    .X(_05218_));
 sg13g2_inv_1 _13193_ (.Y(_05219_),
    .A(_05218_));
 sg13g2_nor2_1 _13194_ (.A(_05213_),
    .B(_05219_),
    .Y(_05220_));
 sg13g2_o21ai_1 _13195_ (.B1(net166),
    .Y(_05221_),
    .A1(_05188_),
    .A2(net160));
 sg13g2_buf_1 _13196_ (.A(_05221_),
    .X(_05223_));
 sg13g2_nor2_1 _13197_ (.A(_05188_),
    .B(net160),
    .Y(_05224_));
 sg13g2_nand2_1 _13198_ (.Y(_05225_),
    .A(net137),
    .B(_05224_));
 sg13g2_nor2_1 _13199_ (.A(net301),
    .B(_00043_),
    .Y(_05226_));
 sg13g2_a22oi_1 _13200_ (.Y(_05227_),
    .B1(_05226_),
    .B2(net304),
    .A2(_00502_),
    .A1(net302));
 sg13g2_nand2_1 _13201_ (.Y(_05228_),
    .A(_01764_),
    .B(_01611_));
 sg13g2_nor2_1 _13202_ (.A(_05227_),
    .B(_05228_),
    .Y(_05229_));
 sg13g2_inv_1 _13203_ (.Y(_05230_),
    .A(_05229_));
 sg13g2_a21oi_1 _13204_ (.A1(_05223_),
    .A2(_05225_),
    .Y(_05231_),
    .B1(_05230_));
 sg13g2_a21oi_1 _13205_ (.A1(_05213_),
    .A2(_05219_),
    .Y(_05232_),
    .B1(_05231_));
 sg13g2_nand2_2 _13206_ (.Y(_05234_),
    .A(_01908_),
    .B(_06420_));
 sg13g2_o21ai_1 _13207_ (.B1(_05234_),
    .Y(_05235_),
    .A1(_05220_),
    .A2(_05232_));
 sg13g2_a21o_1 _13208_ (.A2(_05225_),
    .A1(_05223_),
    .B1(_05230_),
    .X(_05236_));
 sg13g2_xnor2_1 _13209_ (.Y(_05237_),
    .A(_05208_),
    .B(_05212_));
 sg13g2_nor2_1 _13210_ (.A(_05237_),
    .B(_05236_),
    .Y(_05238_));
 sg13g2_nor2_1 _13211_ (.A(_05234_),
    .B(_05218_),
    .Y(_05239_));
 sg13g2_a22oi_1 _13212_ (.Y(_05240_),
    .B1(_05238_),
    .B2(_05239_),
    .A2(_05236_),
    .A1(_05220_));
 sg13g2_and3_1 _13213_ (.X(_05241_),
    .A(_05207_),
    .B(_05235_),
    .C(_05240_));
 sg13g2_buf_1 _13214_ (.A(_05241_),
    .X(_05242_));
 sg13g2_a21oi_2 _13215_ (.B1(_05207_),
    .Y(_05243_),
    .A2(_05240_),
    .A1(_05235_));
 sg13g2_nor2_1 _13216_ (.A(net252),
    .B(_02040_),
    .Y(_05245_));
 sg13g2_o21ai_1 _13217_ (.B1(_05245_),
    .Y(_05246_),
    .A1(_05242_),
    .A2(_05243_));
 sg13g2_or3_1 _13218_ (.A(_05245_),
    .B(_05242_),
    .C(_05243_),
    .X(_05247_));
 sg13g2_nand2_1 _13219_ (.Y(_05248_),
    .A(net253),
    .B(net126));
 sg13g2_nand2_1 _13220_ (.Y(_05249_),
    .A(net207),
    .B(net105));
 sg13g2_nor3_1 _13221_ (.A(net259),
    .B(_01675_),
    .C(_01676_),
    .Y(_05250_));
 sg13g2_xnor2_1 _13222_ (.Y(_05251_),
    .A(_05249_),
    .B(_05250_));
 sg13g2_xnor2_1 _13223_ (.Y(_05252_),
    .A(_05248_),
    .B(_05251_));
 sg13g2_a21o_1 _13224_ (.A2(_01757_),
    .A1(_01594_),
    .B1(_01759_),
    .X(_05253_));
 sg13g2_buf_1 _13225_ (.A(_05253_),
    .X(_05254_));
 sg13g2_nand4_1 _13226_ (.B(net253),
    .C(net126),
    .A(net205),
    .Y(_05256_),
    .D(_03270_));
 sg13g2_a22oi_1 _13227_ (.Y(_05257_),
    .B1(_03270_),
    .B2(net253),
    .A2(net126),
    .A1(net205));
 sg13g2_a21o_1 _13228_ (.A2(_05256_),
    .A1(net206),
    .B1(_05257_),
    .X(_05258_));
 sg13g2_nor2_1 _13229_ (.A(_06233_),
    .B(_05257_),
    .Y(_05259_));
 sg13g2_a21oi_1 _13230_ (.A1(net297),
    .A2(_05258_),
    .Y(_05260_),
    .B1(_05259_));
 sg13g2_nand2_1 _13231_ (.Y(_05261_),
    .A(net299),
    .B(net125));
 sg13g2_and2_1 _13232_ (.A(_07466_),
    .B(net126),
    .X(_05262_));
 sg13g2_buf_1 _13233_ (.A(_05262_),
    .X(_05263_));
 sg13g2_nor2b_1 _13234_ (.A(_05261_),
    .B_N(_05263_),
    .Y(_05264_));
 sg13g2_o21ai_1 _13235_ (.B1(_05264_),
    .Y(_05265_),
    .A1(net257),
    .A2(_05254_));
 sg13g2_o21ai_1 _13236_ (.B1(_05265_),
    .Y(_05267_),
    .A1(_05254_),
    .A2(_05260_));
 sg13g2_xor2_1 _13237_ (.B(_05267_),
    .A(_05252_),
    .X(_05268_));
 sg13g2_nand2_2 _13238_ (.Y(_05269_),
    .A(net254),
    .B(_03282_));
 sg13g2_nand3_1 _13239_ (.B(net207),
    .C(net105),
    .A(net205),
    .Y(_05270_));
 sg13g2_a21o_1 _13240_ (.A2(net105),
    .A1(net205),
    .B1(net207),
    .X(_05271_));
 sg13g2_nand3_1 _13241_ (.B(net294),
    .C(_01783_),
    .A(net253),
    .Y(_05272_));
 sg13g2_a21oi_1 _13242_ (.A1(_05270_),
    .A2(_05271_),
    .Y(_05273_),
    .B1(_05272_));
 sg13g2_nand2_1 _13243_ (.Y(_05274_),
    .A(net207),
    .B(_03282_));
 sg13g2_a22oi_1 _13244_ (.Y(_05275_),
    .B1(net185),
    .B2(_07480_),
    .A2(net105),
    .A1(net205));
 sg13g2_nand4_1 _13245_ (.B(_07480_),
    .C(net105),
    .A(net205),
    .Y(_05276_),
    .D(net185));
 sg13g2_o21ai_1 _13246_ (.B1(_05276_),
    .Y(_05278_),
    .A1(_05274_),
    .A2(_05275_));
 sg13g2_or2_1 _13247_ (.X(_05279_),
    .B(_05278_),
    .A(_05273_));
 sg13g2_xnor2_1 _13248_ (.Y(_05280_),
    .A(_05261_),
    .B(_05263_));
 sg13g2_nand2_1 _13249_ (.Y(_05281_),
    .A(_01330_),
    .B(net185));
 sg13g2_xnor2_1 _13250_ (.Y(_05282_),
    .A(_05280_),
    .B(_05281_));
 sg13g2_and2_1 _13251_ (.A(_05273_),
    .B(_05278_),
    .X(_05283_));
 sg13g2_a21oi_1 _13252_ (.A1(_05279_),
    .A2(_05282_),
    .Y(_05284_),
    .B1(_05283_));
 sg13g2_nor2b_1 _13253_ (.A(_05269_),
    .B_N(_05282_),
    .Y(_05285_));
 sg13g2_nor2_1 _13254_ (.A(_05279_),
    .B(_05282_),
    .Y(_05286_));
 sg13g2_a221oi_1 _13255_ (.B2(_05283_),
    .C1(_05286_),
    .B1(_05285_),
    .A1(_05269_),
    .Y(_05287_),
    .A2(_05284_));
 sg13g2_xor2_1 _13256_ (.B(_05287_),
    .A(_05268_),
    .X(_05289_));
 sg13g2_a21o_1 _13257_ (.A2(_05247_),
    .A1(_05246_),
    .B1(_05289_),
    .X(_05290_));
 sg13g2_buf_1 _13258_ (.A(_05290_),
    .X(_05291_));
 sg13g2_nand3_1 _13259_ (.B(_05246_),
    .C(_05247_),
    .A(_05289_),
    .Y(_05292_));
 sg13g2_buf_1 _13260_ (.A(_05292_),
    .X(_05293_));
 sg13g2_nand2_1 _13261_ (.Y(_05294_),
    .A(net250),
    .B(net227));
 sg13g2_nand2_1 _13262_ (.Y(_05295_),
    .A(net266),
    .B(net228));
 sg13g2_nand2_1 _13263_ (.Y(_05296_),
    .A(net265),
    .B(net277));
 sg13g2_xnor2_1 _13264_ (.Y(_05297_),
    .A(_05295_),
    .B(_05296_));
 sg13g2_xnor2_1 _13265_ (.Y(_05298_),
    .A(_05294_),
    .B(_05297_));
 sg13g2_xor2_1 _13266_ (.B(_05218_),
    .A(_05234_),
    .X(_05300_));
 sg13g2_xnor2_1 _13267_ (.Y(_05301_),
    .A(_05213_),
    .B(_05231_));
 sg13g2_xnor2_1 _13268_ (.Y(_05302_),
    .A(_05300_),
    .B(_05301_));
 sg13g2_a21o_1 _13269_ (.A2(_02332_),
    .A1(net251),
    .B1(_05302_),
    .X(_05303_));
 sg13g2_nand2_1 _13270_ (.Y(_05304_),
    .A(net205),
    .B(net105));
 sg13g2_buf_1 _13271_ (.A(net253),
    .X(_05305_));
 sg13g2_nand2_1 _13272_ (.Y(_05306_),
    .A(_05305_),
    .B(net185));
 sg13g2_nor2_1 _13273_ (.A(_05304_),
    .B(_05306_),
    .Y(_05307_));
 sg13g2_nand2_1 _13274_ (.Y(_05308_),
    .A(_05270_),
    .B(_05306_));
 sg13g2_a21oi_1 _13275_ (.A1(_05271_),
    .A2(_05308_),
    .Y(_05309_),
    .B1(net257));
 sg13g2_nor2_1 _13276_ (.A(_06233_),
    .B(_05275_),
    .Y(_05311_));
 sg13g2_or2_1 _13277_ (.X(_05312_),
    .B(_05311_),
    .A(_05309_));
 sg13g2_a22oi_1 _13278_ (.Y(_05313_),
    .B1(_05312_),
    .B2(_03282_),
    .A2(_05307_),
    .A1(_05269_));
 sg13g2_buf_1 _13279_ (.A(net294),
    .X(_05314_));
 sg13g2_and3_1 _13280_ (.X(_05315_),
    .A(net165),
    .B(net219),
    .C(_01783_));
 sg13g2_nor2_1 _13281_ (.A(net259),
    .B(_03271_),
    .Y(_05316_));
 sg13g2_buf_1 _13282_ (.A(net155),
    .X(_05317_));
 sg13g2_nand2_1 _13283_ (.Y(_05318_),
    .A(net113),
    .B(_05254_));
 sg13g2_o21ai_1 _13284_ (.B1(_05318_),
    .Y(_05319_),
    .A1(net113),
    .A2(_05315_));
 sg13g2_a21oi_1 _13285_ (.A1(_05315_),
    .A2(_05316_),
    .Y(_05320_),
    .B1(_05319_));
 sg13g2_xor2_1 _13286_ (.B(_05320_),
    .A(_05280_),
    .X(_05322_));
 sg13g2_xnor2_1 _13287_ (.Y(_05323_),
    .A(_05313_),
    .B(_05322_));
 sg13g2_nand2_1 _13288_ (.Y(_05324_),
    .A(net251),
    .B(net227));
 sg13g2_nor2b_1 _13289_ (.A(_05324_),
    .B_N(_05302_),
    .Y(_05325_));
 sg13g2_a21oi_2 _13290_ (.B1(_05325_),
    .Y(_05326_),
    .A2(_05323_),
    .A1(_05303_));
 sg13g2_xor2_1 _13291_ (.B(_05326_),
    .A(_05298_),
    .X(_05327_));
 sg13g2_a21oi_1 _13292_ (.A1(_05291_),
    .A2(_05293_),
    .Y(_05328_),
    .B1(_05327_));
 sg13g2_and3_1 _13293_ (.X(_05329_),
    .A(_05291_),
    .B(_05293_),
    .C(_05327_));
 sg13g2_buf_1 _13294_ (.A(_05329_),
    .X(_05330_));
 sg13g2_or3_1 _13295_ (.A(_05187_),
    .B(_05328_),
    .C(_05330_),
    .X(_05331_));
 sg13g2_o21ai_1 _13296_ (.B1(_05187_),
    .Y(_05333_),
    .A1(_05328_),
    .A2(_05330_));
 sg13g2_xnor2_1 _13297_ (.Y(_05334_),
    .A(_05324_),
    .B(_05302_));
 sg13g2_xnor2_1 _13298_ (.Y(_05335_),
    .A(_05323_),
    .B(_05334_));
 sg13g2_nand2_1 _13299_ (.Y(_05336_),
    .A(net215),
    .B(net174));
 sg13g2_nand2_1 _13300_ (.Y(_05337_),
    .A(net250),
    .B(net229));
 sg13g2_xor2_1 _13301_ (.B(_05337_),
    .A(_05336_),
    .X(_05338_));
 sg13g2_buf_1 _13302_ (.A(_05305_),
    .X(_05339_));
 sg13g2_nand3_1 _13303_ (.B(_01329_),
    .C(net185),
    .A(net135),
    .Y(_05340_));
 sg13g2_nand2b_1 _13304_ (.Y(_05341_),
    .B(_05340_),
    .A_N(_01332_));
 sg13g2_a22oi_1 _13305_ (.Y(_05342_),
    .B1(_05341_),
    .B2(_03282_),
    .A2(_05274_),
    .A1(_05306_));
 sg13g2_xnor2_1 _13306_ (.Y(_05344_),
    .A(_05316_),
    .B(_05342_));
 sg13g2_nand2_1 _13307_ (.Y(_05345_),
    .A(net138),
    .B(net210));
 sg13g2_a21oi_1 _13308_ (.A1(net183),
    .A2(_06420_),
    .Y(_05346_),
    .B1(_05345_));
 sg13g2_nor2_1 _13309_ (.A(_05345_),
    .B(_05214_),
    .Y(_05347_));
 sg13g2_a22oi_1 _13310_ (.Y(_05348_),
    .B1(_05347_),
    .B2(net240),
    .A2(_05345_),
    .A1(_06771_));
 sg13g2_o21ai_1 _13311_ (.B1(_05348_),
    .Y(_05349_),
    .A1(net137),
    .A2(_05346_));
 sg13g2_xor2_1 _13312_ (.B(_05349_),
    .A(_05224_),
    .X(_05350_));
 sg13g2_nand2_1 _13313_ (.Y(_05351_),
    .A(_05344_),
    .B(_05350_));
 sg13g2_nand2_1 _13314_ (.Y(_05352_),
    .A(net251),
    .B(net229));
 sg13g2_o21ai_1 _13315_ (.B1(_05352_),
    .Y(_05353_),
    .A1(_05344_),
    .A2(_05350_));
 sg13g2_nand3_1 _13316_ (.B(_05351_),
    .C(_05353_),
    .A(_05338_),
    .Y(_05355_));
 sg13g2_or2_1 _13317_ (.X(_05356_),
    .B(_05355_),
    .A(_05335_));
 sg13g2_a21oi_1 _13318_ (.A1(_05331_),
    .A2(_05333_),
    .Y(_05357_),
    .B1(_05356_));
 sg13g2_nand2_1 _13319_ (.Y(_05358_),
    .A(_05351_),
    .B(_05353_));
 sg13g2_nand2b_1 _13320_ (.Y(_05359_),
    .B(_05335_),
    .A_N(_05338_));
 sg13g2_xnor2_1 _13321_ (.Y(_05360_),
    .A(_05335_),
    .B(_05338_));
 sg13g2_nand2_1 _13322_ (.Y(_05361_),
    .A(_05358_),
    .B(_05360_));
 sg13g2_o21ai_1 _13323_ (.B1(_05361_),
    .Y(_05362_),
    .A1(_05358_),
    .A2(_05359_));
 sg13g2_and3_1 _13324_ (.X(_05363_),
    .A(_05331_),
    .B(_05333_),
    .C(_05362_));
 sg13g2_xnor2_1 _13325_ (.Y(_05364_),
    .A(_05344_),
    .B(_05352_));
 sg13g2_xnor2_1 _13326_ (.Y(_05366_),
    .A(_05350_),
    .B(_05364_));
 sg13g2_a22oi_1 _13327_ (.Y(_05367_),
    .B1(_03282_),
    .B2(_01331_),
    .A2(_02307_),
    .A1(_01758_));
 sg13g2_nor2_1 _13328_ (.A(net255),
    .B(_05367_),
    .Y(_05368_));
 sg13g2_or2_1 _13329_ (.X(_05369_),
    .B(_01758_),
    .A(_01981_));
 sg13g2_o21ai_1 _13330_ (.B1(_02283_),
    .Y(_05370_),
    .A1(net135),
    .A2(net146));
 sg13g2_o21ai_1 _13331_ (.B1(_05370_),
    .Y(_05371_),
    .A1(net146),
    .A2(_05369_));
 sg13g2_a21oi_1 _13332_ (.A1(_01781_),
    .A2(_05369_),
    .Y(_05372_),
    .B1(net135));
 sg13g2_o21ai_1 _13333_ (.B1(_05314_),
    .Y(_05373_),
    .A1(_05371_),
    .A2(_05372_));
 sg13g2_nor2b_1 _13334_ (.A(_05368_),
    .B_N(_05373_),
    .Y(_05374_));
 sg13g2_nor2_1 _13335_ (.A(_00043_),
    .B(net240),
    .Y(_05375_));
 sg13g2_nand2_1 _13336_ (.Y(_05377_),
    .A(_04959_),
    .B(_04955_));
 sg13g2_xnor2_1 _13337_ (.Y(_05378_),
    .A(_05375_),
    .B(_05377_));
 sg13g2_nand2_1 _13338_ (.Y(_05379_),
    .A(net266),
    .B(net183));
 sg13g2_o21ai_1 _13339_ (.B1(_05379_),
    .Y(_05380_),
    .A1(net216),
    .A2(net188));
 sg13g2_nand3_1 _13340_ (.B(net188),
    .C(net183),
    .A(net264),
    .Y(_05381_));
 sg13g2_o21ai_1 _13341_ (.B1(_05381_),
    .Y(_05382_),
    .A1(net188),
    .A2(_01926_));
 sg13g2_a22oi_1 _13342_ (.Y(_05383_),
    .B1(_05382_),
    .B2(_00932_),
    .A2(_05380_),
    .A1(_00449_));
 sg13g2_nand2_1 _13343_ (.Y(_05384_),
    .A(net263),
    .B(_05383_));
 sg13g2_o21ai_1 _13344_ (.B1(_05384_),
    .Y(_05385_),
    .A1(_00245_),
    .A2(_05378_));
 sg13g2_or2_1 _13345_ (.X(_05386_),
    .B(_05385_),
    .A(_05374_));
 sg13g2_a21oi_1 _13346_ (.A1(_05366_),
    .A2(_05386_),
    .Y(_05388_),
    .B1(net204));
 sg13g2_a221oi_1 _13347_ (.B2(_05385_),
    .C1(net252),
    .B1(_05374_),
    .A1(net204),
    .Y(_05389_),
    .A2(_05366_));
 sg13g2_o21ai_1 _13348_ (.B1(_04971_),
    .Y(_05390_),
    .A1(_05388_),
    .A2(_05389_));
 sg13g2_o21ai_1 _13349_ (.B1(_05390_),
    .Y(_05391_),
    .A1(_05366_),
    .A2(_05386_));
 sg13g2_o21ai_1 _13350_ (.B1(_05391_),
    .Y(_05392_),
    .A1(_05357_),
    .A2(_05363_));
 sg13g2_a21oi_1 _13351_ (.A1(_05351_),
    .A2(_05353_),
    .Y(_05393_),
    .B1(_05338_));
 sg13g2_o21ai_1 _13352_ (.B1(_05355_),
    .Y(_05394_),
    .A1(_05335_),
    .A2(_05393_));
 sg13g2_nor3_1 _13353_ (.A(_05187_),
    .B(_05328_),
    .C(_05330_),
    .Y(_05395_));
 sg13g2_a21oi_1 _13354_ (.A1(_05333_),
    .A2(_05394_),
    .Y(_05396_),
    .B1(_05395_));
 sg13g2_o21ai_1 _13355_ (.B1(_05284_),
    .Y(_05397_),
    .A1(_05269_),
    .A2(_05286_));
 sg13g2_nand2_1 _13356_ (.Y(_05399_),
    .A(_05314_),
    .B(_07467_));
 sg13g2_nor4_1 _13357_ (.A(_05254_),
    .B(_05269_),
    .C(_05304_),
    .D(_05399_),
    .Y(_05400_));
 sg13g2_a22oi_1 _13358_ (.Y(_05401_),
    .B1(_05400_),
    .B2(_05282_),
    .A2(_05397_),
    .A1(_05268_));
 sg13g2_buf_1 _13359_ (.A(_05401_),
    .X(_05402_));
 sg13g2_nor2_1 _13360_ (.A(net206),
    .B(_05257_),
    .Y(_05403_));
 sg13g2_o21ai_1 _13361_ (.B1(_05403_),
    .Y(_05404_),
    .A1(net254),
    .A2(_05252_));
 sg13g2_o21ai_1 _13362_ (.B1(net254),
    .Y(_05405_),
    .A1(_05252_),
    .A2(_05264_));
 sg13g2_nand2_1 _13363_ (.Y(_05406_),
    .A(_05404_),
    .B(_05405_));
 sg13g2_a22oi_1 _13364_ (.Y(_05407_),
    .B1(_05406_),
    .B2(net185),
    .A2(_05264_),
    .A1(_05252_));
 sg13g2_buf_2 _13365_ (.A(_05407_),
    .X(_05408_));
 sg13g2_nand2_1 _13366_ (.Y(_05410_),
    .A(net165),
    .B(net108));
 sg13g2_nand2_1 _13367_ (.Y(_05411_),
    .A(net207),
    .B(_01679_));
 sg13g2_nand3_1 _13368_ (.B(_01602_),
    .C(_01604_),
    .A(_06684_),
    .Y(_05412_));
 sg13g2_buf_1 _13369_ (.A(_05412_),
    .X(_05413_));
 sg13g2_xor2_1 _13370_ (.B(_05413_),
    .A(_05411_),
    .X(_05414_));
 sg13g2_xnor2_1 _13371_ (.Y(_05415_),
    .A(_05410_),
    .B(_05414_));
 sg13g2_nand2_1 _13372_ (.Y(_05416_),
    .A(net205),
    .B(net108));
 sg13g2_nand3_1 _13373_ (.B(_01678_),
    .C(_05263_),
    .A(net253),
    .Y(_05417_));
 sg13g2_buf_1 _13374_ (.A(_05417_),
    .X(_05418_));
 sg13g2_a22oi_1 _13375_ (.Y(_05419_),
    .B1(_05418_),
    .B2(_07453_),
    .A2(_05416_),
    .A1(_05248_));
 sg13g2_a21o_1 _13376_ (.A2(_01679_),
    .A1(net165),
    .B1(_05250_),
    .X(_05421_));
 sg13g2_nand2_1 _13377_ (.Y(_05422_),
    .A(_07416_),
    .B(_05421_));
 sg13g2_o21ai_1 _13378_ (.B1(_05422_),
    .Y(_05423_),
    .A1(net257),
    .A2(_05419_));
 sg13g2_nor2_1 _13379_ (.A(net257),
    .B(_03271_),
    .Y(_05424_));
 sg13g2_nor2_1 _13380_ (.A(_05418_),
    .B(_05424_),
    .Y(_05425_));
 sg13g2_a21oi_1 _13381_ (.A1(net105),
    .A2(_05423_),
    .Y(_05426_),
    .B1(_05425_));
 sg13g2_xor2_1 _13382_ (.B(_05426_),
    .A(_05415_),
    .X(_05427_));
 sg13g2_buf_2 _13383_ (.A(_05427_),
    .X(_05428_));
 sg13g2_xnor2_1 _13384_ (.Y(_05429_),
    .A(_05408_),
    .B(_05428_));
 sg13g2_xnor2_1 _13385_ (.Y(_05430_),
    .A(_05402_),
    .B(_05429_));
 sg13g2_nand2_1 _13386_ (.Y(_05432_),
    .A(net251),
    .B(net175));
 sg13g2_o21ai_1 _13387_ (.B1(_01922_),
    .Y(_05433_),
    .A1(net166),
    .A2(_05216_));
 sg13g2_nand2_1 _13388_ (.Y(_05434_),
    .A(_06420_),
    .B(_05433_));
 sg13g2_or2_1 _13389_ (.X(_05435_),
    .B(_05223_),
    .A(_05230_));
 sg13g2_and3_1 _13390_ (.X(_05436_),
    .A(_05215_),
    .B(_05434_),
    .C(_05435_));
 sg13g2_o21ai_1 _13391_ (.B1(_05225_),
    .Y(_05437_),
    .A1(_05234_),
    .A2(_05223_));
 sg13g2_a21oi_1 _13392_ (.A1(_05229_),
    .A2(_05437_),
    .Y(_05438_),
    .B1(_05239_));
 sg13g2_o21ai_1 _13393_ (.B1(_05438_),
    .Y(_05439_),
    .A1(_05237_),
    .A2(_05436_));
 sg13g2_xor2_1 _13394_ (.B(_05206_),
    .A(_05195_),
    .X(_05440_));
 sg13g2_a22oi_1 _13395_ (.Y(_05441_),
    .B1(_05439_),
    .B2(_05440_),
    .A2(_05239_),
    .A1(_05238_));
 sg13g2_a21o_1 _13396_ (.A2(_05210_),
    .A1(_05198_),
    .B1(_05199_),
    .X(_05443_));
 sg13g2_nand2_1 _13397_ (.Y(_05444_),
    .A(_05204_),
    .B(_05443_));
 sg13g2_nor2_1 _13398_ (.A(_05204_),
    .B(_05443_),
    .Y(_05445_));
 sg13g2_a21oi_1 _13399_ (.A1(_05195_),
    .A2(_05444_),
    .Y(_05446_),
    .B1(_05445_));
 sg13g2_nand2_1 _13400_ (.Y(_05447_),
    .A(_01560_),
    .B(net161));
 sg13g2_or3_1 _13401_ (.A(_01542_),
    .B(_05376_),
    .C(_05420_),
    .X(_05448_));
 sg13g2_buf_1 _13402_ (.A(_05448_),
    .X(_05449_));
 sg13g2_or2_1 _13403_ (.X(_05450_),
    .B(_06024_),
    .A(net208));
 sg13g2_nand3_1 _13404_ (.B(_07021_),
    .C(_05450_),
    .A(net239),
    .Y(_05451_));
 sg13g2_xor2_1 _13405_ (.B(_05451_),
    .A(_05449_),
    .X(_05452_));
 sg13g2_xnor2_1 _13406_ (.Y(_05454_),
    .A(_05447_),
    .B(_05452_));
 sg13g2_nand2_1 _13407_ (.Y(_05455_),
    .A(_05190_),
    .B(_05191_));
 sg13g2_o21ai_1 _13408_ (.B1(net137),
    .Y(_05456_),
    .A1(_05190_),
    .A2(_05191_));
 sg13g2_buf_1 _13409_ (.A(_05456_),
    .X(_05457_));
 sg13g2_nand2_1 _13410_ (.Y(_05458_),
    .A(net271),
    .B(net209));
 sg13g2_a21o_1 _13411_ (.A2(_05457_),
    .A1(_05455_),
    .B1(_05458_),
    .X(_05459_));
 sg13g2_a21oi_1 _13412_ (.A1(_05190_),
    .A2(_05191_),
    .Y(_05460_),
    .B1(_01908_));
 sg13g2_a22oi_1 _13413_ (.Y(_05461_),
    .B1(_05457_),
    .B2(_05460_),
    .A2(_05455_),
    .A1(net160));
 sg13g2_and3_1 _13414_ (.X(_05462_),
    .A(_05454_),
    .B(_05459_),
    .C(_05461_));
 sg13g2_a21oi_1 _13415_ (.A1(_05459_),
    .A2(_05461_),
    .Y(_05463_),
    .B1(_05454_));
 sg13g2_nor2_1 _13416_ (.A(_05462_),
    .B(_05463_),
    .Y(_05465_));
 sg13g2_xor2_1 _13417_ (.B(_05465_),
    .A(_05446_),
    .X(_05466_));
 sg13g2_xnor2_1 _13418_ (.Y(_05467_),
    .A(_05441_),
    .B(_05466_));
 sg13g2_xor2_1 _13419_ (.B(_05467_),
    .A(_05432_),
    .X(_05468_));
 sg13g2_xnor2_1 _13420_ (.Y(_05469_),
    .A(_05430_),
    .B(_05468_));
 sg13g2_nand2_1 _13421_ (.Y(_05470_),
    .A(net216),
    .B(_02288_));
 sg13g2_nand2_1 _13422_ (.Y(_05471_),
    .A(net250),
    .B(_02304_));
 sg13g2_nand2_1 _13423_ (.Y(_05472_),
    .A(net215),
    .B(_02333_));
 sg13g2_xnor2_1 _13424_ (.Y(_05473_),
    .A(_05471_),
    .B(_05472_));
 sg13g2_xnor2_1 _13425_ (.Y(_05474_),
    .A(_05470_),
    .B(_05473_));
 sg13g2_nand2_1 _13426_ (.Y(_05476_),
    .A(net196),
    .B(net146));
 sg13g2_nor3_1 _13427_ (.A(_05289_),
    .B(_05242_),
    .C(_05243_),
    .Y(_05477_));
 sg13g2_o21ai_1 _13428_ (.B1(_05289_),
    .Y(_05478_),
    .A1(_05242_),
    .A2(_05243_));
 sg13g2_o21ai_1 _13429_ (.B1(_05478_),
    .Y(_05479_),
    .A1(_05476_),
    .A2(_05477_));
 sg13g2_xor2_1 _13430_ (.B(_05479_),
    .A(_05474_),
    .X(_05480_));
 sg13g2_xnor2_1 _13431_ (.Y(_05481_),
    .A(_05469_),
    .B(_05480_));
 sg13g2_nor2_1 _13432_ (.A(_05294_),
    .B(_05296_),
    .Y(_05482_));
 sg13g2_nand2_1 _13433_ (.Y(_05483_),
    .A(net214),
    .B(_04971_));
 sg13g2_nor2_1 _13434_ (.A(net216),
    .B(_05482_),
    .Y(_05484_));
 sg13g2_a21oi_1 _13435_ (.A1(_05294_),
    .A2(_05296_),
    .Y(_05485_),
    .B1(_05484_));
 sg13g2_nand2_1 _13436_ (.Y(_05487_),
    .A(_05294_),
    .B(_05296_));
 sg13g2_a21oi_1 _13437_ (.A1(net216),
    .A2(_05487_),
    .Y(_05488_),
    .B1(_05027_));
 sg13g2_a21oi_1 _13438_ (.A1(_05027_),
    .A2(_05485_),
    .Y(_05489_),
    .B1(_05488_));
 sg13g2_a22oi_1 _13439_ (.Y(_05490_),
    .B1(_05489_),
    .B2(net136),
    .A2(_05483_),
    .A1(_05482_));
 sg13g2_buf_1 _13440_ (.A(_05490_),
    .X(_05491_));
 sg13g2_nor2_1 _13441_ (.A(_05298_),
    .B(_05326_),
    .Y(_05492_));
 sg13g2_a21oi_1 _13442_ (.A1(_05291_),
    .A2(_05293_),
    .Y(_05493_),
    .B1(_05492_));
 sg13g2_a21oi_2 _13443_ (.B1(_05493_),
    .Y(_05494_),
    .A2(_05326_),
    .A1(_05298_));
 sg13g2_xnor2_1 _13444_ (.Y(_05495_),
    .A(_05491_),
    .B(_05494_));
 sg13g2_xnor2_1 _13445_ (.Y(_05496_),
    .A(_05481_),
    .B(_05495_));
 sg13g2_xnor2_1 _13446_ (.Y(_05498_),
    .A(_05396_),
    .B(_05496_));
 sg13g2_xor2_1 _13447_ (.B(_05498_),
    .A(_05392_),
    .X(_05499_));
 sg13g2_xnor2_1 _13448_ (.Y(_05500_),
    .A(_04046_),
    .B(_05499_));
 sg13g2_a21oi_1 _13449_ (.A1(_04956_),
    .A2(_05500_),
    .Y(_05501_),
    .B1(_05018_));
 sg13g2_mux2_1 _13450_ (.A0(_05501_),
    .A1(net219),
    .S(net15),
    .X(_00224_));
 sg13g2_nand2_2 _13451_ (.Y(_05502_),
    .A(net219),
    .B(net124));
 sg13g2_nand2_1 _13452_ (.Y(_05503_),
    .A(net155),
    .B(net107));
 sg13g2_nand2_1 _13453_ (.Y(_05504_),
    .A(net165),
    .B(net110));
 sg13g2_xnor2_1 _13454_ (.Y(_05505_),
    .A(_05503_),
    .B(_05504_));
 sg13g2_xnor2_1 _13455_ (.Y(_05506_),
    .A(_05502_),
    .B(_05505_));
 sg13g2_and4_1 _13456_ (.A(net165),
    .B(net294),
    .C(net107),
    .D(net110),
    .X(_05508_));
 sg13g2_buf_1 _13457_ (.A(_05508_),
    .X(_05509_));
 sg13g2_buf_1 _13458_ (.A(net254),
    .X(_05510_));
 sg13g2_nand2_1 _13459_ (.Y(_05511_),
    .A(net164),
    .B(_01854_));
 sg13g2_a22oi_1 _13460_ (.Y(_05512_),
    .B1(net110),
    .B2(net294),
    .A2(net107),
    .A1(net165));
 sg13g2_nor2_1 _13461_ (.A(net155),
    .B(_05509_),
    .Y(_05513_));
 sg13g2_o21ai_1 _13462_ (.B1(net164),
    .Y(_05514_),
    .A1(_05512_),
    .A2(_05513_));
 sg13g2_o21ai_1 _13463_ (.B1(_05514_),
    .Y(_05515_),
    .A1(_06233_),
    .A2(_05512_));
 sg13g2_a22oi_1 _13464_ (.Y(_05516_),
    .B1(_05515_),
    .B2(_01854_),
    .A2(_05511_),
    .A1(_05509_));
 sg13g2_xnor2_1 _13465_ (.Y(_05517_),
    .A(_05506_),
    .B(_05516_));
 sg13g2_a22oi_1 _13466_ (.Y(_05519_),
    .B1(_05421_),
    .B2(net155),
    .A2(_05415_),
    .A1(net254));
 sg13g2_o21ai_1 _13467_ (.B1(_05418_),
    .Y(_05520_),
    .A1(_03271_),
    .A2(_05519_));
 sg13g2_o21ai_1 _13468_ (.B1(_05520_),
    .Y(_05521_),
    .A1(_05415_),
    .A2(_05424_));
 sg13g2_buf_1 _13469_ (.A(_05521_),
    .X(_05522_));
 sg13g2_nand2_1 _13470_ (.Y(_05523_),
    .A(net155),
    .B(net108));
 sg13g2_o21ai_1 _13471_ (.B1(_01604_),
    .Y(_05524_),
    .A1(net253),
    .A2(_01533_));
 sg13g2_nor2_1 _13472_ (.A(_01628_),
    .B(_01527_),
    .Y(_05525_));
 sg13g2_a22oi_1 _13473_ (.Y(_05526_),
    .B1(_01629_),
    .B2(net255),
    .A2(_05525_),
    .A1(_01600_));
 sg13g2_nor2_1 _13474_ (.A(_01506_),
    .B(net190),
    .Y(_05527_));
 sg13g2_nor2b_1 _13475_ (.A(_05526_),
    .B_N(_05527_),
    .Y(_05528_));
 sg13g2_a21o_1 _13476_ (.A2(_05524_),
    .A1(_01626_),
    .B1(_05528_),
    .X(_05530_));
 sg13g2_nand3_1 _13477_ (.B(_01628_),
    .C(_01569_),
    .A(net294),
    .Y(_05531_));
 sg13g2_nand3_1 _13478_ (.B(_01602_),
    .C(_01604_),
    .A(_01331_),
    .Y(_05532_));
 sg13g2_nand3_1 _13479_ (.B(_05531_),
    .C(_05532_),
    .A(_01568_),
    .Y(_05533_));
 sg13g2_a22oi_1 _13480_ (.Y(_05534_),
    .B1(_05533_),
    .B2(net165),
    .A2(_05530_),
    .A1(_01328_));
 sg13g2_xnor2_1 _13481_ (.Y(_05535_),
    .A(_05523_),
    .B(_05534_));
 sg13g2_and2_1 _13482_ (.A(_05411_),
    .B(_05413_),
    .X(_05536_));
 sg13g2_or2_1 _13483_ (.X(_05537_),
    .B(_05413_),
    .A(_05411_));
 sg13g2_o21ai_1 _13484_ (.B1(_05537_),
    .Y(_05538_),
    .A1(_05410_),
    .A2(_05536_));
 sg13g2_buf_1 _13485_ (.A(_05538_),
    .X(_05539_));
 sg13g2_nand2_1 _13486_ (.Y(_05541_),
    .A(net254),
    .B(net126));
 sg13g2_xor2_1 _13487_ (.B(_05541_),
    .A(_05539_),
    .X(_05542_));
 sg13g2_xnor2_1 _13488_ (.Y(_05543_),
    .A(_05535_),
    .B(_05542_));
 sg13g2_nand2_1 _13489_ (.Y(_05544_),
    .A(_05522_),
    .B(_05543_));
 sg13g2_nor2_1 _13490_ (.A(_05408_),
    .B(_05428_),
    .Y(_05545_));
 sg13g2_a21oi_1 _13491_ (.A1(_05408_),
    .A2(_05428_),
    .Y(_05546_),
    .B1(_05402_));
 sg13g2_nor2_1 _13492_ (.A(_05522_),
    .B(_05543_),
    .Y(_05547_));
 sg13g2_or3_1 _13493_ (.A(_05545_),
    .B(_05546_),
    .C(_05547_),
    .X(_05548_));
 sg13g2_buf_1 _13494_ (.A(_05548_),
    .X(_05549_));
 sg13g2_nand4_1 _13495_ (.B(net219),
    .C(net107),
    .A(net155),
    .Y(_05550_),
    .D(net108));
 sg13g2_nand2_1 _13496_ (.Y(_05552_),
    .A(net135),
    .B(_01854_));
 sg13g2_a22oi_1 _13497_ (.Y(_05553_),
    .B1(net108),
    .B2(net113),
    .A2(net107),
    .A1(net219));
 sg13g2_a21o_1 _13498_ (.A2(_05552_),
    .A1(_05550_),
    .B1(_05553_),
    .X(_05554_));
 sg13g2_buf_1 _13499_ (.A(_05554_),
    .X(_05555_));
 sg13g2_nor2b_1 _13500_ (.A(_05539_),
    .B_N(_05541_),
    .Y(_05556_));
 sg13g2_nand3_1 _13501_ (.B(net126),
    .C(_05539_),
    .A(net164),
    .Y(_05557_));
 sg13g2_o21ai_1 _13502_ (.B1(_05557_),
    .Y(_05558_),
    .A1(_05535_),
    .A2(_05556_));
 sg13g2_buf_2 _13503_ (.A(_05558_),
    .X(_05559_));
 sg13g2_nand2_1 _13504_ (.Y(_05560_),
    .A(net165),
    .B(net107));
 sg13g2_and3_1 _13505_ (.X(_05561_),
    .A(net206),
    .B(net281),
    .C(_02745_));
 sg13g2_nor3_1 _13506_ (.A(net281),
    .B(_01516_),
    .C(_02745_),
    .Y(_05563_));
 sg13g2_o21ai_1 _13507_ (.B1(_05527_),
    .Y(_05564_),
    .A1(_05561_),
    .A2(_05563_));
 sg13g2_o21ai_1 _13508_ (.B1(net206),
    .Y(_05565_),
    .A1(_01544_),
    .A2(_01512_));
 sg13g2_a21o_1 _13509_ (.A2(_05565_),
    .A1(_01604_),
    .B1(_01640_),
    .X(_05566_));
 sg13g2_nand2_1 _13510_ (.Y(_05567_),
    .A(_05564_),
    .B(_05566_));
 sg13g2_nor3_1 _13511_ (.A(_02745_),
    .B(_01512_),
    .C(_01566_),
    .Y(_05568_));
 sg13g2_o21ai_1 _13512_ (.B1(net281),
    .Y(_05569_),
    .A1(_01564_),
    .A2(_05568_));
 sg13g2_xor2_1 _13513_ (.B(_01516_),
    .A(_01640_),
    .X(_05570_));
 sg13g2_nand3_1 _13514_ (.B(_02745_),
    .C(_05570_),
    .A(net294),
    .Y(_05571_));
 sg13g2_nand3_1 _13515_ (.B(_05569_),
    .C(_05571_),
    .A(_05532_),
    .Y(_05572_));
 sg13g2_a22oi_1 _13516_ (.Y(_05574_),
    .B1(_05572_),
    .B2(net155),
    .A2(_05567_),
    .A1(net294));
 sg13g2_xnor2_1 _13517_ (.Y(_05575_),
    .A(_05560_),
    .B(_05574_));
 sg13g2_buf_2 _13518_ (.A(_05575_),
    .X(_05576_));
 sg13g2_nand2_1 _13519_ (.Y(_05577_),
    .A(net254),
    .B(net108));
 sg13g2_buf_2 _13520_ (.A(_05577_),
    .X(_05578_));
 sg13g2_nor2_1 _13521_ (.A(_05576_),
    .B(_05578_),
    .Y(_05579_));
 sg13g2_nand2_1 _13522_ (.Y(_05580_),
    .A(_05576_),
    .B(_05578_));
 sg13g2_o21ai_1 _13523_ (.B1(_05580_),
    .Y(_05581_),
    .A1(_05559_),
    .A2(_05579_));
 sg13g2_nor2_1 _13524_ (.A(_05559_),
    .B(_05580_),
    .Y(_05582_));
 sg13g2_a21oi_1 _13525_ (.A1(net70),
    .A2(_05581_),
    .Y(_05583_),
    .B1(_05582_));
 sg13g2_a21oi_1 _13526_ (.A1(_05544_),
    .A2(_05549_),
    .Y(_05585_),
    .B1(_05583_));
 sg13g2_nor3_1 _13527_ (.A(_05576_),
    .B(_05578_),
    .C(net70),
    .Y(_05586_));
 sg13g2_a22oi_1 _13528_ (.Y(_05587_),
    .B1(_05582_),
    .B2(net70),
    .A2(_05586_),
    .A1(_05559_));
 sg13g2_inv_1 _13529_ (.Y(_05588_),
    .A(_05587_));
 sg13g2_inv_1 _13530_ (.Y(_05589_),
    .A(_05544_));
 sg13g2_nor3_1 _13531_ (.A(_05545_),
    .B(_05546_),
    .C(_05547_),
    .Y(_05590_));
 sg13g2_nor2_1 _13532_ (.A(net70),
    .B(_05581_),
    .Y(_05591_));
 sg13g2_a21oi_1 _13533_ (.A1(_05559_),
    .A2(_05579_),
    .Y(_05592_),
    .B1(_05591_));
 sg13g2_nor3_1 _13534_ (.A(_05589_),
    .B(_05590_),
    .C(_05592_),
    .Y(_05593_));
 sg13g2_nor3_1 _13535_ (.A(_05585_),
    .B(_05588_),
    .C(_05593_),
    .Y(_05594_));
 sg13g2_xor2_1 _13536_ (.B(_05594_),
    .A(_05517_),
    .X(_05596_));
 sg13g2_nand2_1 _13537_ (.Y(_05597_),
    .A(net138),
    .B(net130));
 sg13g2_nor3_1 _13538_ (.A(net240),
    .B(_07313_),
    .C(_07321_),
    .Y(_05598_));
 sg13g2_nor3_1 _13539_ (.A(net239),
    .B(_05980_),
    .C(_06035_),
    .Y(_05599_));
 sg13g2_nor3_1 _13540_ (.A(_07317_),
    .B(_05598_),
    .C(_05599_),
    .Y(_05600_));
 sg13g2_nand3_1 _13541_ (.B(_04705_),
    .C(_07313_),
    .A(_07316_),
    .Y(_05601_));
 sg13g2_nand3_1 _13542_ (.B(_01538_),
    .C(_00737_),
    .A(_07315_),
    .Y(_05602_));
 sg13g2_nand2_1 _13543_ (.Y(_05603_),
    .A(net211),
    .B(_05958_));
 sg13g2_a21oi_1 _13544_ (.A1(_05601_),
    .A2(_05602_),
    .Y(_05604_),
    .B1(_05603_));
 sg13g2_o21ai_1 _13545_ (.B1(net166),
    .Y(_05605_),
    .A1(net208),
    .A2(_07325_));
 sg13g2_a21oi_1 _13546_ (.A1(_07021_),
    .A2(_05605_),
    .Y(_05607_),
    .B1(net330));
 sg13g2_o21ai_1 _13547_ (.B1(net239),
    .Y(_05608_),
    .A1(_05604_),
    .A2(_05607_));
 sg13g2_o21ai_1 _13548_ (.B1(_05608_),
    .Y(_05609_),
    .A1(_05192_),
    .A2(_05600_));
 sg13g2_xor2_1 _13549_ (.B(_05609_),
    .A(_05597_),
    .X(_05610_));
 sg13g2_nand3_1 _13550_ (.B(_07021_),
    .C(_05450_),
    .A(net138),
    .Y(_05611_));
 sg13g2_nor3_1 _13551_ (.A(_05192_),
    .B(_05376_),
    .C(_05420_),
    .Y(_05612_));
 sg13g2_a21oi_1 _13552_ (.A1(net239),
    .A2(net130),
    .Y(_05613_),
    .B1(_05612_));
 sg13g2_nand4_1 _13553_ (.B(_05343_),
    .C(net261),
    .A(net301),
    .Y(_05614_),
    .D(_04563_));
 sg13g2_o21ai_1 _13554_ (.B1(_05354_),
    .Y(_05615_),
    .A1(_04823_),
    .A2(_05398_));
 sg13g2_nand3_1 _13555_ (.B(_05614_),
    .C(_05615_),
    .A(_06912_),
    .Y(_05616_));
 sg13g2_nand3_1 _13556_ (.B(_05343_),
    .C(net261),
    .A(net301),
    .Y(_05618_));
 sg13g2_o21ai_1 _13557_ (.B1(_06902_),
    .Y(_05619_),
    .A1(_04563_),
    .A2(_05618_));
 sg13g2_nand4_1 _13558_ (.B(net239),
    .C(_05616_),
    .A(net137),
    .Y(_05620_),
    .D(_05619_));
 sg13g2_o21ai_1 _13559_ (.B1(_05620_),
    .Y(_05621_),
    .A1(_05611_),
    .A2(_05613_));
 sg13g2_buf_1 _13560_ (.A(_05621_),
    .X(_05622_));
 sg13g2_or2_1 _13561_ (.X(_05623_),
    .B(_07336_),
    .A(_01922_));
 sg13g2_buf_1 _13562_ (.A(_05623_),
    .X(_05624_));
 sg13g2_xnor2_1 _13563_ (.Y(_05625_),
    .A(_05622_),
    .B(_05624_));
 sg13g2_xnor2_1 _13564_ (.Y(_05626_),
    .A(_05610_),
    .B(_05625_));
 sg13g2_nand2_1 _13565_ (.Y(_05627_),
    .A(_05447_),
    .B(_05449_));
 sg13g2_o21ai_1 _13566_ (.B1(_05451_),
    .Y(_05629_),
    .A1(_05447_),
    .A2(_05449_));
 sg13g2_nand2_1 _13567_ (.Y(_05630_),
    .A(_05627_),
    .B(_05629_));
 sg13g2_nand2_1 _13568_ (.Y(_05631_),
    .A(net239),
    .B(net130));
 sg13g2_xnor2_1 _13569_ (.Y(_05632_),
    .A(_05611_),
    .B(_05612_));
 sg13g2_xor2_1 _13570_ (.B(_05632_),
    .A(_05631_),
    .X(_05633_));
 sg13g2_nand2_1 _13571_ (.Y(_05634_),
    .A(net271),
    .B(_05925_));
 sg13g2_a21o_1 _13572_ (.A2(_05633_),
    .A1(_05630_),
    .B1(_05634_),
    .X(_05635_));
 sg13g2_o21ai_1 _13573_ (.B1(_05635_),
    .Y(_05636_),
    .A1(_05630_),
    .A2(_05633_));
 sg13g2_buf_1 _13574_ (.A(_05636_),
    .X(_05637_));
 sg13g2_nand2_2 _13575_ (.Y(_05638_),
    .A(_05626_),
    .B(_05637_));
 sg13g2_xor2_1 _13576_ (.B(_05634_),
    .A(_05630_),
    .X(_05640_));
 sg13g2_xnor2_1 _13577_ (.Y(_05641_),
    .A(_05633_),
    .B(_05640_));
 sg13g2_nand2_1 _13578_ (.Y(_05642_),
    .A(_05455_),
    .B(_05457_));
 sg13g2_o21ai_1 _13579_ (.B1(net271),
    .Y(_05643_),
    .A1(_05454_),
    .A2(_05642_));
 sg13g2_nand2b_1 _13580_ (.Y(_05644_),
    .B(_05454_),
    .A_N(_05457_));
 sg13g2_a21oi_1 _13581_ (.A1(_05643_),
    .A2(_05644_),
    .Y(_05645_),
    .B1(_06189_));
 sg13g2_nor2b_1 _13582_ (.A(_05455_),
    .B_N(_05454_),
    .Y(_05646_));
 sg13g2_nor3_1 _13583_ (.A(_05641_),
    .B(_05645_),
    .C(_05646_),
    .Y(_05647_));
 sg13g2_nor2b_1 _13584_ (.A(_05465_),
    .B_N(_05446_),
    .Y(_05648_));
 sg13g2_nor3_1 _13585_ (.A(_05446_),
    .B(_05462_),
    .C(_05463_),
    .Y(_05649_));
 sg13g2_a221oi_1 _13586_ (.B2(_05440_),
    .C1(_05649_),
    .B1(_05439_),
    .A1(_05238_),
    .Y(_05651_),
    .A2(_05239_));
 sg13g2_buf_1 _13587_ (.A(_05651_),
    .X(_05652_));
 sg13g2_nor3_1 _13588_ (.A(_05647_),
    .B(_05648_),
    .C(_05652_),
    .Y(_05653_));
 sg13g2_or2_1 _13589_ (.X(_05654_),
    .B(_05646_),
    .A(_05645_));
 sg13g2_and2_1 _13590_ (.A(_05641_),
    .B(_05654_),
    .X(_05655_));
 sg13g2_or2_1 _13591_ (.X(_05656_),
    .B(_05637_),
    .A(_05626_));
 sg13g2_o21ai_1 _13592_ (.B1(_05656_),
    .Y(_05657_),
    .A1(_05653_),
    .A2(_05655_));
 sg13g2_nand2b_1 _13593_ (.Y(_05658_),
    .B(_05622_),
    .A_N(_05624_));
 sg13g2_nor2b_1 _13594_ (.A(_05622_),
    .B_N(_05624_),
    .Y(_05659_));
 sg13g2_a21o_1 _13595_ (.A2(_05658_),
    .A1(_05610_),
    .B1(_05659_),
    .X(_05660_));
 sg13g2_buf_1 _13596_ (.A(_05660_),
    .X(_05662_));
 sg13g2_nand2_2 _13597_ (.Y(_05663_),
    .A(net138),
    .B(net94));
 sg13g2_or3_1 _13598_ (.A(_01538_),
    .B(_06923_),
    .C(_06956_),
    .X(_05664_));
 sg13g2_buf_1 _13599_ (.A(_05664_),
    .X(_05665_));
 sg13g2_and2_1 _13600_ (.A(net239),
    .B(net129),
    .X(_05666_));
 sg13g2_xnor2_1 _13601_ (.Y(_05667_),
    .A(_05665_),
    .B(_05666_));
 sg13g2_xor2_1 _13602_ (.B(_05667_),
    .A(_05663_),
    .X(_05668_));
 sg13g2_buf_2 _13603_ (.A(_05668_),
    .X(_05669_));
 sg13g2_a22oi_1 _13604_ (.Y(_05670_),
    .B1(_07483_),
    .B2(_01925_),
    .A2(net130),
    .A1(net138));
 sg13g2_nand2_1 _13605_ (.Y(_05671_),
    .A(net137),
    .B(_07411_));
 sg13g2_nand4_1 _13606_ (.B(_01925_),
    .C(net130),
    .A(net138),
    .Y(_05673_),
    .D(net94));
 sg13g2_o21ai_1 _13607_ (.B1(_05673_),
    .Y(_05674_),
    .A1(_05670_),
    .A2(_05671_));
 sg13g2_buf_1 _13608_ (.A(_05674_),
    .X(_05675_));
 sg13g2_nand2_2 _13609_ (.Y(_05676_),
    .A(net271),
    .B(_07411_));
 sg13g2_xnor2_1 _13610_ (.Y(_05677_),
    .A(net64),
    .B(_05676_));
 sg13g2_xor2_1 _13611_ (.B(_05677_),
    .A(_05669_),
    .X(_05678_));
 sg13g2_xnor2_1 _13612_ (.Y(_05679_),
    .A(_05662_),
    .B(_05678_));
 sg13g2_a21o_1 _13613_ (.A2(_05657_),
    .A1(_05638_),
    .B1(_05679_),
    .X(_05680_));
 sg13g2_nand3_1 _13614_ (.B(_05638_),
    .C(_05657_),
    .A(_05679_),
    .Y(_05681_));
 sg13g2_and2_1 _13615_ (.A(_05680_),
    .B(_05681_),
    .X(_05682_));
 sg13g2_buf_1 _13616_ (.A(_05682_),
    .X(_05684_));
 sg13g2_nand2_1 _13617_ (.Y(_05685_),
    .A(net196),
    .B(_02007_));
 sg13g2_nor2b_1 _13618_ (.A(_05684_),
    .B_N(_05685_),
    .Y(_05686_));
 sg13g2_nand2b_1 _13619_ (.Y(_05687_),
    .B(_05684_),
    .A_N(_05685_));
 sg13g2_o21ai_1 _13620_ (.B1(_05687_),
    .Y(_05688_),
    .A1(_05596_),
    .A2(_05686_));
 sg13g2_a21oi_1 _13621_ (.A1(_05576_),
    .A2(_05578_),
    .Y(_05689_),
    .B1(net70));
 sg13g2_xor2_1 _13622_ (.B(_05578_),
    .A(_05576_),
    .X(_05690_));
 sg13g2_nor2b_1 _13623_ (.A(_05690_),
    .B_N(net70),
    .Y(_05691_));
 sg13g2_nor2_1 _13624_ (.A(_05689_),
    .B(_05691_),
    .Y(_05692_));
 sg13g2_mux2_1 _13625_ (.A0(_05692_),
    .A1(_05586_),
    .S(_05517_),
    .X(_05693_));
 sg13g2_a22oi_1 _13626_ (.Y(_05695_),
    .B1(_05559_),
    .B2(_05693_),
    .A2(_05549_),
    .A1(_05544_));
 sg13g2_buf_2 _13627_ (.A(_05695_),
    .X(_05696_));
 sg13g2_nor2b_1 _13628_ (.A(_05559_),
    .B_N(net70),
    .Y(_05697_));
 sg13g2_nor2_1 _13629_ (.A(_05580_),
    .B(_05697_),
    .Y(_05698_));
 sg13g2_a21oi_1 _13630_ (.A1(net70),
    .A2(_05690_),
    .Y(_05699_),
    .B1(_05698_));
 sg13g2_mux2_1 _13631_ (.A0(_05699_),
    .A1(_05592_),
    .S(_05517_),
    .X(_05700_));
 sg13g2_buf_1 _13632_ (.A(_05700_),
    .X(_05701_));
 sg13g2_nor2_1 _13633_ (.A(_05696_),
    .B(_05701_),
    .Y(_05702_));
 sg13g2_nand2_1 _13634_ (.Y(_05703_),
    .A(_05502_),
    .B(_05504_));
 sg13g2_o21ai_1 _13635_ (.B1(net107),
    .Y(_05704_),
    .A1(net164),
    .A2(_05703_));
 sg13g2_nand3_1 _13636_ (.B(net164),
    .C(_05703_),
    .A(net113),
    .Y(_05706_));
 sg13g2_nor2b_1 _13637_ (.A(_05704_),
    .B_N(_05706_),
    .Y(_05707_));
 sg13g2_nor2_1 _13638_ (.A(_05502_),
    .B(_05504_),
    .Y(_05708_));
 sg13g2_o21ai_1 _13639_ (.B1(net206),
    .Y(_05709_),
    .A1(net257),
    .A2(_05708_));
 sg13g2_nand2_1 _13640_ (.Y(_05710_),
    .A(net164),
    .B(net107));
 sg13g2_a22oi_1 _13641_ (.Y(_05711_),
    .B1(_05710_),
    .B2(_05708_),
    .A2(_05709_),
    .A1(_05707_));
 sg13g2_nand2_1 _13642_ (.Y(_05712_),
    .A(net113),
    .B(net110));
 sg13g2_xor2_1 _13643_ (.B(net219),
    .A(net135),
    .X(_05713_));
 sg13g2_nand2_1 _13644_ (.Y(_05714_),
    .A(net124),
    .B(_05713_));
 sg13g2_xnor2_1 _13645_ (.Y(_05715_),
    .A(_05712_),
    .B(_05714_));
 sg13g2_xnor2_1 _13646_ (.Y(_05717_),
    .A(_05711_),
    .B(_05715_));
 sg13g2_inv_1 _13647_ (.Y(_05718_),
    .A(_05717_));
 sg13g2_a21oi_1 _13648_ (.A1(net113),
    .A2(_01854_),
    .Y(_05719_),
    .B1(_05509_));
 sg13g2_or2_1 _13649_ (.X(_05720_),
    .B(_05719_),
    .A(_05512_));
 sg13g2_buf_1 _13650_ (.A(_05720_),
    .X(_05721_));
 sg13g2_nor2_1 _13651_ (.A(_05579_),
    .B(_05689_),
    .Y(_05722_));
 sg13g2_nor2_1 _13652_ (.A(_05721_),
    .B(_05722_),
    .Y(_05723_));
 sg13g2_nor2_2 _13653_ (.A(_05506_),
    .B(_05511_),
    .Y(_05724_));
 sg13g2_nand2_1 _13654_ (.Y(_05725_),
    .A(_05721_),
    .B(_05722_));
 sg13g2_and2_1 _13655_ (.A(_05506_),
    .B(_05511_),
    .X(_05726_));
 sg13g2_o21ai_1 _13656_ (.B1(_05726_),
    .Y(_05728_),
    .A1(_05721_),
    .A2(_05722_));
 sg13g2_o21ai_1 _13657_ (.B1(_05728_),
    .Y(_05729_),
    .A1(_05724_),
    .A2(_05725_));
 sg13g2_a21oi_1 _13658_ (.A1(_05723_),
    .A2(_05724_),
    .Y(_05730_),
    .B1(_05729_));
 sg13g2_xnor2_1 _13659_ (.Y(_05731_),
    .A(_05718_),
    .B(_05730_));
 sg13g2_xnor2_1 _13660_ (.Y(_05732_),
    .A(_05702_),
    .B(_05731_));
 sg13g2_nand2_1 _13661_ (.Y(_05733_),
    .A(net196),
    .B(_02031_));
 sg13g2_nor2_1 _13662_ (.A(_05663_),
    .B(_05665_),
    .Y(_05734_));
 sg13g2_nand2_1 _13663_ (.Y(_05735_),
    .A(_05663_),
    .B(_05665_));
 sg13g2_o21ai_1 _13664_ (.B1(_05735_),
    .Y(_05736_),
    .A1(_05666_),
    .A2(_05734_));
 sg13g2_nand2_1 _13665_ (.Y(_05737_),
    .A(net271),
    .B(net130));
 sg13g2_nand2_1 _13666_ (.Y(_05739_),
    .A(net137),
    .B(_07483_));
 sg13g2_nand2_1 _13667_ (.Y(_05740_),
    .A(net129),
    .B(_01651_));
 sg13g2_xor2_1 _13668_ (.B(_05740_),
    .A(_05739_),
    .X(_05741_));
 sg13g2_xnor2_1 _13669_ (.Y(_05742_),
    .A(_05737_),
    .B(_05741_));
 sg13g2_xnor2_1 _13670_ (.Y(_05743_),
    .A(_05736_),
    .B(_05742_));
 sg13g2_buf_1 _13671_ (.A(_05743_),
    .X(_05744_));
 sg13g2_nor2_1 _13672_ (.A(_05669_),
    .B(_05676_),
    .Y(_05745_));
 sg13g2_nand2_1 _13673_ (.Y(_05746_),
    .A(_05669_),
    .B(_05676_));
 sg13g2_o21ai_1 _13674_ (.B1(_05746_),
    .Y(_05747_),
    .A1(net64),
    .A2(_05745_));
 sg13g2_nand2_1 _13675_ (.Y(_05748_),
    .A(_05663_),
    .B(_05667_));
 sg13g2_or2_1 _13676_ (.X(_05750_),
    .B(_05667_),
    .A(_05663_));
 sg13g2_a221oi_1 _13677_ (.B2(_05750_),
    .C1(_05659_),
    .B1(_05748_),
    .A1(_05610_),
    .Y(_05751_),
    .A2(_05658_));
 sg13g2_nand3_1 _13678_ (.B(_07411_),
    .C(net64),
    .A(net271),
    .Y(_05752_));
 sg13g2_buf_1 _13679_ (.A(_05752_),
    .X(_05753_));
 sg13g2_inv_1 _13680_ (.Y(_05754_),
    .A(_05753_));
 sg13g2_nor2_1 _13681_ (.A(net64),
    .B(_05746_),
    .Y(_05755_));
 sg13g2_a221oi_1 _13682_ (.B2(_05754_),
    .C1(_05755_),
    .B1(_05751_),
    .A1(_05662_),
    .Y(_05756_),
    .A2(_05747_));
 sg13g2_xnor2_1 _13683_ (.Y(_05757_),
    .A(net46),
    .B(_05756_));
 sg13g2_xnor2_1 _13684_ (.Y(_05758_),
    .A(_05680_),
    .B(_05757_));
 sg13g2_xnor2_1 _13685_ (.Y(_05759_),
    .A(_05733_),
    .B(_05758_));
 sg13g2_xnor2_1 _13686_ (.Y(_05761_),
    .A(_05732_),
    .B(_05759_));
 sg13g2_nand2_1 _13687_ (.Y(_05762_),
    .A(net162),
    .B(net151));
 sg13g2_buf_1 _13688_ (.A(net250),
    .X(_05763_));
 sg13g2_nand2_1 _13689_ (.Y(_05764_),
    .A(_05763_),
    .B(net180));
 sg13g2_buf_1 _13690_ (.A(net215),
    .X(_05765_));
 sg13g2_nand2_1 _13691_ (.Y(_05766_),
    .A(net134),
    .B(_02014_));
 sg13g2_xnor2_1 _13692_ (.Y(_05767_),
    .A(_05764_),
    .B(_05766_));
 sg13g2_xnor2_1 _13693_ (.Y(_05768_),
    .A(_05762_),
    .B(_05767_));
 sg13g2_xnor2_1 _13694_ (.Y(_05769_),
    .A(_05761_),
    .B(_05768_));
 sg13g2_xnor2_1 _13695_ (.Y(_05770_),
    .A(_05688_),
    .B(_05769_));
 sg13g2_buf_2 _13696_ (.A(_05770_),
    .X(_05772_));
 sg13g2_xnor2_1 _13697_ (.Y(_05773_),
    .A(_05685_),
    .B(_05684_));
 sg13g2_xnor2_1 _13698_ (.Y(_05774_),
    .A(_05596_),
    .B(_05773_));
 sg13g2_xor2_1 _13699_ (.B(_05555_),
    .A(_05578_),
    .X(_05775_));
 sg13g2_xnor2_1 _13700_ (.Y(_05776_),
    .A(_05576_),
    .B(_05775_));
 sg13g2_xnor2_1 _13701_ (.Y(_05777_),
    .A(_05559_),
    .B(_05776_));
 sg13g2_inv_1 _13702_ (.Y(_05778_),
    .A(_05777_));
 sg13g2_a21oi_1 _13703_ (.A1(_05544_),
    .A2(_05549_),
    .Y(_05779_),
    .B1(_05778_));
 sg13g2_nor3_1 _13704_ (.A(_05589_),
    .B(_05590_),
    .C(_05777_),
    .Y(_05780_));
 sg13g2_nor2_1 _13705_ (.A(_05653_),
    .B(_05655_),
    .Y(_05781_));
 sg13g2_nand2_1 _13706_ (.Y(_05783_),
    .A(_05638_),
    .B(_05656_));
 sg13g2_xnor2_1 _13707_ (.Y(_05784_),
    .A(_05781_),
    .B(_05783_));
 sg13g2_o21ai_1 _13708_ (.B1(_05784_),
    .Y(_05785_),
    .A1(_05779_),
    .A2(_05780_));
 sg13g2_nor2_1 _13709_ (.A(net252),
    .B(_02188_),
    .Y(_05786_));
 sg13g2_nor3_1 _13710_ (.A(_05784_),
    .B(_05779_),
    .C(_05780_),
    .Y(_05787_));
 sg13g2_a21oi_2 _13711_ (.B1(_05787_),
    .Y(_05788_),
    .A2(_05786_),
    .A1(_05785_));
 sg13g2_nand2_1 _13712_ (.Y(_05789_),
    .A(_04968_),
    .B(net144));
 sg13g2_nand2_1 _13713_ (.Y(_05790_),
    .A(_05763_),
    .B(net179));
 sg13g2_nand2_1 _13714_ (.Y(_05791_),
    .A(_05765_),
    .B(_02016_));
 sg13g2_xnor2_1 _13715_ (.Y(_05792_),
    .A(_05790_),
    .B(_05791_));
 sg13g2_xnor2_1 _13716_ (.Y(_05794_),
    .A(_05789_),
    .B(_05792_));
 sg13g2_nand2_1 _13717_ (.Y(_05795_),
    .A(_05788_),
    .B(_05794_));
 sg13g2_nor2_1 _13718_ (.A(_05788_),
    .B(_05794_),
    .Y(_05796_));
 sg13g2_a21oi_2 _13719_ (.B1(_05796_),
    .Y(_05797_),
    .A2(_05795_),
    .A1(_05774_));
 sg13g2_nor2_1 _13720_ (.A(_05772_),
    .B(_05797_),
    .Y(_05798_));
 sg13g2_nand2_1 _13721_ (.Y(_05799_),
    .A(net212),
    .B(net145));
 sg13g2_nand2_1 _13722_ (.Y(_05800_),
    .A(net268),
    .B(net114));
 sg13g2_buf_1 _13723_ (.A(net214),
    .X(_05801_));
 sg13g2_nand2_1 _13724_ (.Y(_05802_),
    .A(net133),
    .B(_03213_));
 sg13g2_xnor2_1 _13725_ (.Y(_05803_),
    .A(_05800_),
    .B(_05802_));
 sg13g2_xnor2_1 _13726_ (.Y(_05805_),
    .A(_05799_),
    .B(_05803_));
 sg13g2_and2_1 _13727_ (.A(_05790_),
    .B(_05791_),
    .X(_05806_));
 sg13g2_or2_1 _13728_ (.X(_05807_),
    .B(_05791_),
    .A(_05790_));
 sg13g2_o21ai_1 _13729_ (.B1(_05807_),
    .Y(_05808_),
    .A1(_05789_),
    .A2(_05806_));
 sg13g2_buf_1 _13730_ (.A(_05808_),
    .X(_05809_));
 sg13g2_nand2_1 _13731_ (.Y(_05810_),
    .A(_05233_),
    .B(net170));
 sg13g2_nand2_1 _13732_ (.Y(_05811_),
    .A(net268),
    .B(net145));
 sg13g2_nand2_1 _13733_ (.Y(_05812_),
    .A(net214),
    .B(net114));
 sg13g2_and2_1 _13734_ (.A(_05811_),
    .B(_05812_),
    .X(_05813_));
 sg13g2_or2_1 _13735_ (.X(_05814_),
    .B(_05812_),
    .A(_05811_));
 sg13g2_o21ai_1 _13736_ (.B1(_05814_),
    .Y(_05816_),
    .A1(_05810_),
    .A2(_05813_));
 sg13g2_buf_1 _13737_ (.A(_05816_),
    .X(_05817_));
 sg13g2_xor2_1 _13738_ (.B(_05817_),
    .A(_05809_),
    .X(_05818_));
 sg13g2_xnor2_1 _13739_ (.Y(_05819_),
    .A(_05805_),
    .B(_05818_));
 sg13g2_inv_1 _13740_ (.Y(_05820_),
    .A(_05819_));
 sg13g2_a21oi_1 _13741_ (.A1(_05772_),
    .A2(_05797_),
    .Y(_05821_),
    .B1(_05820_));
 sg13g2_nand2_1 _13742_ (.Y(_05822_),
    .A(_05809_),
    .B(_05817_));
 sg13g2_nor2_1 _13743_ (.A(_05809_),
    .B(_05817_),
    .Y(_05823_));
 sg13g2_a21oi_1 _13744_ (.A1(_05805_),
    .A2(_05822_),
    .Y(_05824_),
    .B1(_05823_));
 sg13g2_nand2_1 _13745_ (.Y(_05825_),
    .A(net213),
    .B(net170));
 sg13g2_nand2_1 _13746_ (.Y(_05827_),
    .A(net201),
    .B(net145));
 sg13g2_o21ai_1 _13747_ (.B1(_05827_),
    .Y(_05828_),
    .A1(net201),
    .A2(_05825_));
 sg13g2_nor2_1 _13748_ (.A(net249),
    .B(net202),
    .Y(_05829_));
 sg13g2_a221oi_1 _13749_ (.B2(_02041_),
    .C1(net169),
    .B1(_05829_),
    .A1(net199),
    .Y(_05830_),
    .A2(_05828_));
 sg13g2_or2_1 _13750_ (.X(_05831_),
    .B(_05827_),
    .A(_05825_));
 sg13g2_and2_1 _13751_ (.A(_03018_),
    .B(_05831_),
    .X(_05832_));
 sg13g2_a21oi_1 _13752_ (.A1(net249),
    .A2(net136),
    .Y(_05833_),
    .B1(net201));
 sg13g2_o21ai_1 _13753_ (.B1(_05825_),
    .Y(_05834_),
    .A1(_03022_),
    .A2(_05833_));
 sg13g2_o21ai_1 _13754_ (.B1(_05834_),
    .Y(_05835_),
    .A1(_05830_),
    .A2(_05832_));
 sg13g2_nand2b_1 _13755_ (.Y(_05836_),
    .B(_05835_),
    .A_N(_05824_));
 sg13g2_buf_1 _13756_ (.A(_05836_),
    .X(_05838_));
 sg13g2_nand2b_1 _13757_ (.Y(_05839_),
    .B(_05824_),
    .A_N(_05835_));
 sg13g2_nand2_1 _13758_ (.Y(_05840_),
    .A(_05838_),
    .B(_05839_));
 sg13g2_nor3_1 _13759_ (.A(_05798_),
    .B(_05821_),
    .C(_05840_),
    .Y(_05841_));
 sg13g2_nand2_1 _13760_ (.Y(_05842_),
    .A(_05772_),
    .B(_05797_));
 sg13g2_o21ai_1 _13761_ (.B1(_05820_),
    .Y(_05843_),
    .A1(_05772_),
    .A2(_05797_));
 sg13g2_and3_1 _13762_ (.X(_05844_),
    .A(_05842_),
    .B(_05843_),
    .C(_05840_));
 sg13g2_o21ai_1 _13763_ (.B1(_05729_),
    .Y(_05845_),
    .A1(_05696_),
    .A2(_05701_));
 sg13g2_inv_1 _13764_ (.Y(_05846_),
    .A(_05726_));
 sg13g2_a21o_1 _13765_ (.A2(_05846_),
    .A1(_05725_),
    .B1(_05724_),
    .X(_05847_));
 sg13g2_a22oi_1 _13766_ (.Y(_05849_),
    .B1(_05847_),
    .B2(_05702_),
    .A2(_05845_),
    .A1(_05718_));
 sg13g2_inv_1 _13767_ (.Y(_05850_),
    .A(_05725_));
 sg13g2_nor3_1 _13768_ (.A(_05696_),
    .B(_05701_),
    .C(_05850_),
    .Y(_05851_));
 sg13g2_o21ai_1 _13769_ (.B1(_05723_),
    .Y(_05852_),
    .A1(_05724_),
    .A2(_05851_));
 sg13g2_nor2_1 _13770_ (.A(net257),
    .B(_01553_),
    .Y(_05853_));
 sg13g2_nor2_1 _13771_ (.A(_05317_),
    .B(net219),
    .Y(_05854_));
 sg13g2_nand2_1 _13772_ (.Y(_05855_),
    .A(_07456_),
    .B(_05854_));
 sg13g2_nand3_1 _13773_ (.B(_05399_),
    .C(_05855_),
    .A(net124),
    .Y(_05856_));
 sg13g2_nand2_1 _13774_ (.Y(_05857_),
    .A(net219),
    .B(_01553_));
 sg13g2_a21oi_1 _13775_ (.A1(_07454_),
    .A2(_05857_),
    .Y(_05858_),
    .B1(_01332_));
 sg13g2_nand2_1 _13776_ (.Y(_05860_),
    .A(net257),
    .B(_01331_));
 sg13g2_nor2_1 _13777_ (.A(_01553_),
    .B(_05860_),
    .Y(_05861_));
 sg13g2_nor2_1 _13778_ (.A(net113),
    .B(net110),
    .Y(_05862_));
 sg13g2_o21ai_1 _13779_ (.B1(net135),
    .Y(_05863_),
    .A1(_05861_),
    .A2(_05862_));
 sg13g2_o21ai_1 _13780_ (.B1(_05863_),
    .Y(_05864_),
    .A1(_05853_),
    .A2(_05858_));
 sg13g2_a22oi_1 _13781_ (.Y(_05865_),
    .B1(_05864_),
    .B2(net124),
    .A2(_05856_),
    .A1(_05853_));
 sg13g2_a21oi_1 _13782_ (.A1(_01331_),
    .A2(net124),
    .Y(_05866_),
    .B1(net255));
 sg13g2_nor2_1 _13783_ (.A(net164),
    .B(_05866_),
    .Y(_05867_));
 sg13g2_a21oi_1 _13784_ (.A1(_01332_),
    .A2(_01553_),
    .Y(_05868_),
    .B1(net257));
 sg13g2_a21oi_1 _13785_ (.A1(net113),
    .A2(_01553_),
    .Y(_05869_),
    .B1(net164));
 sg13g2_nor3_1 _13786_ (.A(net135),
    .B(_01331_),
    .C(_05869_),
    .Y(_05871_));
 sg13g2_a21oi_1 _13787_ (.A1(net135),
    .A2(_05868_),
    .Y(_05872_),
    .B1(_05871_));
 sg13g2_nand2b_1 _13788_ (.Y(_05873_),
    .B(_01921_),
    .A_N(_05872_));
 sg13g2_o21ai_1 _13789_ (.B1(_05873_),
    .Y(_05874_),
    .A1(_05712_),
    .A2(_05867_));
 sg13g2_nor2_1 _13790_ (.A(_07481_),
    .B(_05502_),
    .Y(_05875_));
 sg13g2_a22oi_1 _13791_ (.Y(_05876_),
    .B1(_05875_),
    .B2(net110),
    .A2(_05874_),
    .A1(_01737_));
 sg13g2_xnor2_1 _13792_ (.Y(_05877_),
    .A(_05865_),
    .B(_05876_));
 sg13g2_inv_1 _13793_ (.Y(_05878_),
    .A(_05877_));
 sg13g2_a21o_1 _13794_ (.A2(_05852_),
    .A1(_05849_),
    .B1(_05878_),
    .X(_05879_));
 sg13g2_buf_1 _13795_ (.A(_05879_),
    .X(_05880_));
 sg13g2_nand3_1 _13796_ (.B(_05849_),
    .C(_05852_),
    .A(_05878_),
    .Y(_05882_));
 sg13g2_buf_1 _13797_ (.A(_05882_),
    .X(_05883_));
 sg13g2_nand2_1 _13798_ (.Y(_05884_),
    .A(net196),
    .B(_01500_));
 sg13g2_or3_1 _13799_ (.A(_05647_),
    .B(_05648_),
    .C(_05652_),
    .X(_05885_));
 sg13g2_o21ai_1 _13800_ (.B1(_05641_),
    .Y(_05886_),
    .A1(_05645_),
    .A2(_05646_));
 sg13g2_nand2b_1 _13801_ (.Y(_05887_),
    .B(_05637_),
    .A_N(_05626_));
 sg13g2_nand2b_1 _13802_ (.Y(_05888_),
    .B(_05626_),
    .A_N(_05637_));
 sg13g2_a221oi_1 _13803_ (.B2(_05888_),
    .C1(_05757_),
    .B1(_05887_),
    .A1(_05885_),
    .Y(_05889_),
    .A2(_05886_));
 sg13g2_o21ai_1 _13804_ (.B1(_05638_),
    .Y(_05890_),
    .A1(_05662_),
    .A2(_05669_));
 sg13g2_nor2b_1 _13805_ (.A(net64),
    .B_N(_05676_),
    .Y(_05891_));
 sg13g2_nand2_1 _13806_ (.Y(_05893_),
    .A(_05891_),
    .B(net46));
 sg13g2_o21ai_1 _13807_ (.B1(_05893_),
    .Y(_05894_),
    .A1(_05753_),
    .A2(net46));
 sg13g2_or2_1 _13808_ (.X(_05895_),
    .B(_05891_),
    .A(_05669_));
 sg13g2_nand2_1 _13809_ (.Y(_05896_),
    .A(_05669_),
    .B(_05753_));
 sg13g2_mux2_1 _13810_ (.A0(_05895_),
    .A1(_05896_),
    .S(net46),
    .X(_05897_));
 sg13g2_a21oi_1 _13811_ (.A1(_05610_),
    .A2(_05658_),
    .Y(_05898_),
    .B1(_05659_));
 sg13g2_nand4_1 _13812_ (.B(_05669_),
    .C(_05677_),
    .A(_05898_),
    .Y(_05899_),
    .D(net46));
 sg13g2_o21ai_1 _13813_ (.B1(_05899_),
    .Y(_05900_),
    .A1(_05638_),
    .A2(_05897_));
 sg13g2_a21o_1 _13814_ (.A2(_05894_),
    .A1(_05890_),
    .B1(_05900_),
    .X(_05901_));
 sg13g2_xor2_1 _13815_ (.B(_05676_),
    .A(_05669_),
    .X(_05902_));
 sg13g2_nor3_1 _13816_ (.A(_05662_),
    .B(net64),
    .C(net46),
    .Y(_05904_));
 sg13g2_a21o_1 _13817_ (.A2(net64),
    .A1(_05662_),
    .B1(_05904_),
    .X(_05905_));
 sg13g2_or2_1 _13818_ (.X(_05906_),
    .B(_05746_),
    .A(net46));
 sg13g2_nand2_1 _13819_ (.Y(_05907_),
    .A(_05744_),
    .B(_05745_));
 sg13g2_a21oi_1 _13820_ (.A1(_05906_),
    .A2(_05907_),
    .Y(_05908_),
    .B1(_05662_));
 sg13g2_nor3_1 _13821_ (.A(_05898_),
    .B(net64),
    .C(_05902_),
    .Y(_05909_));
 sg13g2_a221oi_1 _13822_ (.B2(_05675_),
    .C1(_05909_),
    .B1(_05908_),
    .A1(_05902_),
    .Y(_05910_),
    .A2(_05905_));
 sg13g2_o21ai_1 _13823_ (.B1(_05910_),
    .Y(_05911_),
    .A1(_05889_),
    .A2(_05901_));
 sg13g2_nor2_1 _13824_ (.A(net138),
    .B(net183),
    .Y(_05912_));
 sg13g2_inv_1 _13825_ (.Y(_05913_),
    .A(_05912_));
 sg13g2_o21ai_1 _13826_ (.B1(net129),
    .Y(_05915_),
    .A1(net137),
    .A2(_05913_));
 sg13g2_nand3_1 _13827_ (.B(net129),
    .C(_05228_),
    .A(_01922_),
    .Y(_05916_));
 sg13g2_o21ai_1 _13828_ (.B1(_05916_),
    .Y(_05917_),
    .A1(_01922_),
    .A2(_05228_));
 sg13g2_a22oi_1 _13829_ (.Y(_05918_),
    .B1(_05917_),
    .B2(_04961_),
    .A2(_05915_),
    .A1(_04965_));
 sg13g2_inv_1 _13830_ (.Y(_05919_),
    .A(_05918_));
 sg13g2_nand2_1 _13831_ (.Y(_05920_),
    .A(_04961_),
    .B(_05912_));
 sg13g2_nand2_1 _13832_ (.Y(_05921_),
    .A(_04965_),
    .B(net94));
 sg13g2_nand3_1 _13833_ (.B(_05913_),
    .C(_05921_),
    .A(net166),
    .Y(_05922_));
 sg13g2_o21ai_1 _13834_ (.B1(_05922_),
    .Y(_05923_),
    .A1(net94),
    .A2(_05920_));
 sg13g2_a22oi_1 _13835_ (.Y(_05924_),
    .B1(_05923_),
    .B2(net129),
    .A2(_05919_),
    .A1(net94));
 sg13g2_nor2b_1 _13836_ (.A(_05741_),
    .B_N(_05737_),
    .Y(_05926_));
 sg13g2_nand2b_1 _13837_ (.Y(_05927_),
    .B(_05741_),
    .A_N(_05737_));
 sg13g2_o21ai_1 _13838_ (.B1(_05927_),
    .Y(_05928_),
    .A1(_05736_),
    .A2(_05926_));
 sg13g2_xor2_1 _13839_ (.B(_05928_),
    .A(_05924_),
    .X(_05929_));
 sg13g2_nand3b_1 _13840_ (.B(net46),
    .C(_05896_),
    .Y(_05930_),
    .A_N(_05891_));
 sg13g2_xnor2_1 _13841_ (.Y(_05931_),
    .A(_05929_),
    .B(_05930_));
 sg13g2_xnor2_1 _13842_ (.Y(_05932_),
    .A(_05911_),
    .B(_05931_));
 sg13g2_xnor2_1 _13843_ (.Y(_05933_),
    .A(_05884_),
    .B(_05932_));
 sg13g2_inv_1 _13844_ (.Y(_05934_),
    .A(_05933_));
 sg13g2_a21oi_1 _13845_ (.A1(_05880_),
    .A2(_05883_),
    .Y(_05935_),
    .B1(_05934_));
 sg13g2_and3_1 _13846_ (.X(_05937_),
    .A(_05880_),
    .B(_05883_),
    .C(_05934_));
 sg13g2_buf_1 _13847_ (.A(_05937_),
    .X(_05938_));
 sg13g2_nand2_1 _13848_ (.Y(_05939_),
    .A(net162),
    .B(net179));
 sg13g2_nand2_1 _13849_ (.Y(_05940_),
    .A(net163),
    .B(_02031_));
 sg13g2_nand2_1 _13850_ (.Y(_05941_),
    .A(net134),
    .B(net235));
 sg13g2_xnor2_1 _13851_ (.Y(_05942_),
    .A(_05940_),
    .B(_05941_));
 sg13g2_xnor2_1 _13852_ (.Y(_05943_),
    .A(_05939_),
    .B(_05942_));
 sg13g2_nand2_1 _13853_ (.Y(_05944_),
    .A(_05733_),
    .B(_05758_));
 sg13g2_nor2_1 _13854_ (.A(_05733_),
    .B(_05758_),
    .Y(_05945_));
 sg13g2_a21oi_1 _13855_ (.A1(_05732_),
    .A2(_05944_),
    .Y(_05946_),
    .B1(_05945_));
 sg13g2_xnor2_1 _13856_ (.Y(_05948_),
    .A(_05943_),
    .B(_05946_));
 sg13g2_o21ai_1 _13857_ (.B1(_05948_),
    .Y(_05949_),
    .A1(_05935_),
    .A2(_05938_));
 sg13g2_or3_1 _13858_ (.A(_05935_),
    .B(_05938_),
    .C(_05948_),
    .X(_05950_));
 sg13g2_buf_1 _13859_ (.A(_05950_),
    .X(_05951_));
 sg13g2_and2_1 _13860_ (.A(_05949_),
    .B(_05951_),
    .X(_05952_));
 sg13g2_buf_1 _13861_ (.A(_05952_),
    .X(_05953_));
 sg13g2_inv_1 _13862_ (.Y(_05954_),
    .A(_05761_));
 sg13g2_inv_1 _13863_ (.Y(_05955_),
    .A(_05768_));
 sg13g2_o21ai_1 _13864_ (.B1(_05688_),
    .Y(_05956_),
    .A1(_05761_),
    .A2(_05955_));
 sg13g2_o21ai_1 _13865_ (.B1(_05956_),
    .Y(_05957_),
    .A1(_05954_),
    .A2(_05768_));
 sg13g2_nand2_1 _13866_ (.Y(_05959_),
    .A(net212),
    .B(net114));
 sg13g2_nand2_1 _13867_ (.Y(_05960_),
    .A(_04801_),
    .B(net144));
 sg13g2_nand2_1 _13868_ (.Y(_05961_),
    .A(_05801_),
    .B(net151));
 sg13g2_xnor2_1 _13869_ (.Y(_05962_),
    .A(_05960_),
    .B(_05961_));
 sg13g2_xnor2_1 _13870_ (.Y(_05963_),
    .A(_05959_),
    .B(_05962_));
 sg13g2_and2_1 _13871_ (.A(_05764_),
    .B(_05766_),
    .X(_05964_));
 sg13g2_or2_1 _13872_ (.X(_05965_),
    .B(_05766_),
    .A(_05764_));
 sg13g2_o21ai_1 _13873_ (.B1(_05965_),
    .Y(_05966_),
    .A1(_05762_),
    .A2(_05964_));
 sg13g2_buf_1 _13874_ (.A(_05966_),
    .X(_05967_));
 sg13g2_and2_1 _13875_ (.A(_05800_),
    .B(_05802_),
    .X(_05968_));
 sg13g2_or2_1 _13876_ (.X(_05970_),
    .B(_05802_),
    .A(_05800_));
 sg13g2_o21ai_1 _13877_ (.B1(_05970_),
    .Y(_05971_),
    .A1(_05799_),
    .A2(_05968_));
 sg13g2_buf_1 _13878_ (.A(_05971_),
    .X(_05972_));
 sg13g2_xnor2_1 _13879_ (.Y(_05973_),
    .A(_05967_),
    .B(_05972_));
 sg13g2_xnor2_1 _13880_ (.Y(_05974_),
    .A(_05963_),
    .B(_05973_));
 sg13g2_xnor2_1 _13881_ (.Y(_05975_),
    .A(_05957_),
    .B(_05974_));
 sg13g2_xor2_1 _13882_ (.B(_05975_),
    .A(_05953_),
    .X(_05976_));
 sg13g2_o21ai_1 _13883_ (.B1(_05976_),
    .Y(_05977_),
    .A1(_05841_),
    .A2(_05844_));
 sg13g2_buf_1 _13884_ (.A(_05977_),
    .X(_05978_));
 sg13g2_or3_1 _13885_ (.A(_05976_),
    .B(_05841_),
    .C(_05844_),
    .X(_05979_));
 sg13g2_buf_1 _13886_ (.A(_05979_),
    .X(_05981_));
 sg13g2_xnor2_1 _13887_ (.Y(_05982_),
    .A(_05788_),
    .B(_05794_));
 sg13g2_xnor2_1 _13888_ (.Y(_05983_),
    .A(_05774_),
    .B(_05982_));
 sg13g2_xor2_1 _13889_ (.B(_05812_),
    .A(_05811_),
    .X(_05984_));
 sg13g2_xnor2_1 _13890_ (.Y(_05985_),
    .A(_05810_),
    .B(_05984_));
 sg13g2_nand2_1 _13891_ (.Y(_05986_),
    .A(net305),
    .B(_02288_));
 sg13g2_nand2_1 _13892_ (.Y(_05987_),
    .A(net264),
    .B(_02333_));
 sg13g2_and2_1 _13893_ (.A(_05986_),
    .B(_05987_),
    .X(_05988_));
 sg13g2_nand2_1 _13894_ (.Y(_05989_),
    .A(net270),
    .B(_02290_));
 sg13g2_or2_1 _13895_ (.X(_05990_),
    .B(_05987_),
    .A(_05986_));
 sg13g2_o21ai_1 _13896_ (.B1(_05990_),
    .Y(_05992_),
    .A1(_05988_),
    .A2(_05989_));
 sg13g2_nand2_1 _13897_ (.Y(_05993_),
    .A(net250),
    .B(net178));
 sg13g2_nand2_1 _13898_ (.Y(_05994_),
    .A(net215),
    .B(_02282_));
 sg13g2_and2_1 _13899_ (.A(_05993_),
    .B(_05994_),
    .X(_05995_));
 sg13g2_nand2_1 _13900_ (.Y(_05996_),
    .A(net216),
    .B(_05004_));
 sg13g2_or2_1 _13901_ (.X(_05997_),
    .B(_05994_),
    .A(_05993_));
 sg13g2_o21ai_1 _13902_ (.B1(_05997_),
    .Y(_05998_),
    .A1(_05995_),
    .A2(_05996_));
 sg13g2_buf_1 _13903_ (.A(_05998_),
    .X(_05999_));
 sg13g2_xor2_1 _13904_ (.B(_05999_),
    .A(_05992_),
    .X(_06000_));
 sg13g2_xnor2_1 _13905_ (.Y(_06001_),
    .A(_05985_),
    .B(_06000_));
 sg13g2_nor2_1 _13906_ (.A(_05779_),
    .B(_05780_),
    .Y(_06003_));
 sg13g2_xnor2_1 _13907_ (.Y(_06004_),
    .A(_05784_),
    .B(_05786_));
 sg13g2_xor2_1 _13908_ (.B(_06004_),
    .A(_06003_),
    .X(_06005_));
 sg13g2_xor2_1 _13909_ (.B(_05994_),
    .A(_05993_),
    .X(_06006_));
 sg13g2_xnor2_1 _13910_ (.Y(_06007_),
    .A(_05996_),
    .B(_06006_));
 sg13g2_xor2_1 _13911_ (.B(_05543_),
    .A(_05522_),
    .X(_06008_));
 sg13g2_nor3_1 _13912_ (.A(_05545_),
    .B(_05546_),
    .C(_06008_),
    .Y(_06009_));
 sg13g2_nand2_1 _13913_ (.Y(_06010_),
    .A(_05408_),
    .B(_05428_));
 sg13g2_o21ai_1 _13914_ (.B1(_05402_),
    .Y(_06011_),
    .A1(_05408_),
    .A2(_05428_));
 sg13g2_and3_1 _13915_ (.X(_06012_),
    .A(_06010_),
    .B(_06011_),
    .C(_06008_));
 sg13g2_buf_1 _13916_ (.A(_06012_),
    .X(_06014_));
 sg13g2_nor2_1 _13917_ (.A(_05648_),
    .B(_05652_),
    .Y(_06015_));
 sg13g2_nor2b_1 _13918_ (.A(_05647_),
    .B_N(_05886_),
    .Y(_06016_));
 sg13g2_xnor2_1 _13919_ (.Y(_06017_),
    .A(_06015_),
    .B(_06016_));
 sg13g2_o21ai_1 _13920_ (.B1(_06017_),
    .Y(_06018_),
    .A1(_06009_),
    .A2(_06014_));
 sg13g2_nand2_1 _13921_ (.Y(_06019_),
    .A(net251),
    .B(_02015_));
 sg13g2_inv_1 _13922_ (.Y(_06020_),
    .A(_06019_));
 sg13g2_nor3_1 _13923_ (.A(_06017_),
    .B(_06009_),
    .C(_06014_),
    .Y(_06021_));
 sg13g2_a21oi_2 _13924_ (.B1(_06021_),
    .Y(_06022_),
    .A2(_06020_),
    .A1(_06018_));
 sg13g2_nand2b_1 _13925_ (.Y(_06023_),
    .B(_06022_),
    .A_N(_06007_));
 sg13g2_nor2b_1 _13926_ (.A(_06022_),
    .B_N(_06007_),
    .Y(_06025_));
 sg13g2_a21oi_2 _13927_ (.B1(_06025_),
    .Y(_06026_),
    .A2(_06023_),
    .A1(_06005_));
 sg13g2_nand2_1 _13928_ (.Y(_06027_),
    .A(_06001_),
    .B(_06026_));
 sg13g2_nor2_1 _13929_ (.A(_06001_),
    .B(_06026_),
    .Y(_06028_));
 sg13g2_a21o_1 _13930_ (.A2(_06027_),
    .A1(_05983_),
    .B1(_06028_),
    .X(_06029_));
 sg13g2_buf_1 _13931_ (.A(_06029_),
    .X(_06030_));
 sg13g2_nand2_1 _13932_ (.Y(_06031_),
    .A(_05985_),
    .B(_05999_));
 sg13g2_o21ai_1 _13933_ (.B1(_05992_),
    .Y(_06032_),
    .A1(_05985_),
    .A2(_05999_));
 sg13g2_nand2_1 _13934_ (.Y(_06033_),
    .A(_06031_),
    .B(_06032_));
 sg13g2_nand2_1 _13935_ (.Y(_06034_),
    .A(_06030_),
    .B(_06033_));
 sg13g2_nand3_1 _13936_ (.B(_05981_),
    .C(_06034_),
    .A(_05978_),
    .Y(_06036_));
 sg13g2_xnor2_1 _13937_ (.Y(_06037_),
    .A(_05797_),
    .B(_05820_));
 sg13g2_xnor2_1 _13938_ (.Y(_06038_),
    .A(_05772_),
    .B(_06037_));
 sg13g2_buf_1 _13939_ (.A(_06038_),
    .X(_06039_));
 sg13g2_nand2_1 _13940_ (.Y(_06040_),
    .A(_00331_),
    .B(net136));
 sg13g2_nand2_1 _13941_ (.Y(_06041_),
    .A(net201),
    .B(_02739_));
 sg13g2_xnor2_1 _13942_ (.Y(_06042_),
    .A(_06040_),
    .B(_06041_));
 sg13g2_buf_1 _13943_ (.A(_06042_),
    .X(_06043_));
 sg13g2_nor2_1 _13944_ (.A(_06039_),
    .B(_06043_),
    .Y(_06044_));
 sg13g2_nor2_1 _13945_ (.A(_06030_),
    .B(_06033_),
    .Y(_06045_));
 sg13g2_inv_1 _13946_ (.Y(_06047_),
    .A(_06043_));
 sg13g2_a21oi_1 _13947_ (.A1(_06030_),
    .A2(_06033_),
    .Y(_06048_),
    .B1(_06047_));
 sg13g2_or2_1 _13948_ (.X(_06049_),
    .B(_06048_),
    .A(_06045_));
 sg13g2_or2_1 _13949_ (.X(_06050_),
    .B(_06045_),
    .A(_06039_));
 sg13g2_a22oi_1 _13950_ (.Y(_06051_),
    .B1(_06049_),
    .B2(_06050_),
    .A2(_05981_),
    .A1(_05978_));
 sg13g2_a21oi_2 _13951_ (.B1(_06051_),
    .Y(_06052_),
    .A2(_06044_),
    .A1(_06036_));
 sg13g2_a22oi_1 _13952_ (.Y(_06053_),
    .B1(_05884_),
    .B2(_05932_),
    .A2(_05883_),
    .A1(_05880_));
 sg13g2_nor2_1 _13953_ (.A(_05884_),
    .B(_05932_),
    .Y(_06054_));
 sg13g2_nor2_1 _13954_ (.A(_06053_),
    .B(_06054_),
    .Y(_06055_));
 sg13g2_nand2_1 _13955_ (.Y(_06056_),
    .A(_05718_),
    .B(_05725_));
 sg13g2_o21ai_1 _13956_ (.B1(_06056_),
    .Y(_06058_),
    .A1(_05696_),
    .A2(_05701_));
 sg13g2_nand2_1 _13957_ (.Y(_06059_),
    .A(_05717_),
    .B(_05850_));
 sg13g2_a21oi_1 _13958_ (.A1(_06058_),
    .A2(_06059_),
    .Y(_06060_),
    .B1(_05724_));
 sg13g2_a21oi_1 _13959_ (.A1(_05718_),
    .A2(_05846_),
    .Y(_06061_),
    .B1(_05723_));
 sg13g2_o21ai_1 _13960_ (.B1(_06061_),
    .Y(_06062_),
    .A1(_05696_),
    .A2(_05701_));
 sg13g2_nand2b_1 _13961_ (.Y(_06063_),
    .B(_05717_),
    .A_N(_05728_));
 sg13g2_nand3_1 _13962_ (.B(_06062_),
    .C(_06063_),
    .A(_05878_),
    .Y(_06064_));
 sg13g2_nor2_1 _13963_ (.A(_07453_),
    .B(_01331_),
    .Y(_06065_));
 sg13g2_o21ai_1 _13964_ (.B1(_05339_),
    .Y(_06066_),
    .A1(_01553_),
    .A2(_06065_));
 sg13g2_o21ai_1 _13965_ (.B1(_06066_),
    .Y(_06067_),
    .A1(_01557_),
    .A2(_05854_));
 sg13g2_o21ai_1 _13966_ (.B1(_01921_),
    .Y(_06069_),
    .A1(_07468_),
    .A2(_05860_));
 sg13g2_a21oi_1 _13967_ (.A1(_05510_),
    .A2(_06067_),
    .Y(_06070_),
    .B1(_06069_));
 sg13g2_nor2_1 _13968_ (.A(_05865_),
    .B(_05876_),
    .Y(_06071_));
 sg13g2_nor2_1 _13969_ (.A(_06070_),
    .B(_06071_),
    .Y(_06072_));
 sg13g2_o21ai_1 _13970_ (.B1(_06072_),
    .Y(_06073_),
    .A1(_06060_),
    .A2(_06064_));
 sg13g2_or3_1 _13971_ (.A(_06072_),
    .B(_06060_),
    .C(_06064_),
    .X(_06074_));
 sg13g2_buf_1 _13972_ (.A(_06074_),
    .X(_06075_));
 sg13g2_nand2_1 _13973_ (.Y(_06076_),
    .A(_06073_),
    .B(_06075_));
 sg13g2_inv_1 _13974_ (.Y(_06077_),
    .A(_05924_));
 sg13g2_a21o_1 _13975_ (.A2(_05228_),
    .A1(net94),
    .B1(net166),
    .X(_06078_));
 sg13g2_o21ai_1 _13976_ (.B1(_06078_),
    .Y(_06080_),
    .A1(net94),
    .A2(_05912_));
 sg13g2_nand2_1 _13977_ (.Y(_06081_),
    .A(net129),
    .B(_01924_));
 sg13g2_a21oi_1 _13978_ (.A1(net271),
    .A2(_06080_),
    .Y(_06082_),
    .B1(_06081_));
 sg13g2_a21oi_1 _13979_ (.A1(_06077_),
    .A2(_05928_),
    .Y(_06083_),
    .B1(_06082_));
 sg13g2_a21oi_1 _13980_ (.A1(_05911_),
    .A2(_05930_),
    .Y(_06084_),
    .B1(_05929_));
 sg13g2_xnor2_1 _13981_ (.Y(_06085_),
    .A(_06083_),
    .B(_06084_));
 sg13g2_and2_1 _13982_ (.A(net196),
    .B(_01489_),
    .X(_06086_));
 sg13g2_xnor2_1 _13983_ (.Y(_06087_),
    .A(_06085_),
    .B(_06086_));
 sg13g2_xnor2_1 _13984_ (.Y(_06088_),
    .A(_06076_),
    .B(_06087_));
 sg13g2_nand2_1 _13985_ (.Y(_06089_),
    .A(net162),
    .B(net180));
 sg13g2_nand2_1 _13986_ (.Y(_06091_),
    .A(net163),
    .B(net231));
 sg13g2_nand2_1 _13987_ (.Y(_06092_),
    .A(net134),
    .B(net177));
 sg13g2_xor2_1 _13988_ (.B(_06092_),
    .A(_06091_),
    .X(_06093_));
 sg13g2_xnor2_1 _13989_ (.Y(_06094_),
    .A(_06089_),
    .B(_06093_));
 sg13g2_xor2_1 _13990_ (.B(_06094_),
    .A(_06088_),
    .X(_06095_));
 sg13g2_xnor2_1 _13991_ (.Y(_06096_),
    .A(_06055_),
    .B(_06095_));
 sg13g2_or2_1 _13992_ (.X(_06097_),
    .B(_05938_),
    .A(_05935_));
 sg13g2_nand2_1 _13993_ (.Y(_06098_),
    .A(_05943_),
    .B(_05946_));
 sg13g2_nor2_1 _13994_ (.A(_05943_),
    .B(_05946_),
    .Y(_06099_));
 sg13g2_a21oi_1 _13995_ (.A1(_06097_),
    .A2(_06098_),
    .Y(_06100_),
    .B1(_06099_));
 sg13g2_nand2_1 _13996_ (.Y(_06102_),
    .A(net212),
    .B(net144));
 sg13g2_nand2_1 _13997_ (.Y(_06103_),
    .A(net268),
    .B(_02016_));
 sg13g2_nand2_1 _13998_ (.Y(_06104_),
    .A(net214),
    .B(_02013_));
 sg13g2_xnor2_1 _13999_ (.Y(_06105_),
    .A(_06103_),
    .B(_06104_));
 sg13g2_xnor2_1 _14000_ (.Y(_06106_),
    .A(_06102_),
    .B(_06105_));
 sg13g2_and2_1 _14001_ (.A(_05940_),
    .B(_05941_),
    .X(_06107_));
 sg13g2_or2_1 _14002_ (.X(_06108_),
    .B(_05941_),
    .A(_05940_));
 sg13g2_o21ai_1 _14003_ (.B1(_06108_),
    .Y(_06109_),
    .A1(_05939_),
    .A2(_06107_));
 sg13g2_buf_1 _14004_ (.A(_06109_),
    .X(_06110_));
 sg13g2_and2_1 _14005_ (.A(_05960_),
    .B(_05961_),
    .X(_06111_));
 sg13g2_or2_1 _14006_ (.X(_06113_),
    .B(_05961_),
    .A(_05960_));
 sg13g2_o21ai_1 _14007_ (.B1(_06113_),
    .Y(_06114_),
    .A1(_05959_),
    .A2(_06111_));
 sg13g2_buf_1 _14008_ (.A(_06114_),
    .X(_06115_));
 sg13g2_xnor2_1 _14009_ (.Y(_06116_),
    .A(_06110_),
    .B(_06115_));
 sg13g2_xnor2_1 _14010_ (.Y(_06117_),
    .A(_06106_),
    .B(_06116_));
 sg13g2_xor2_1 _14011_ (.B(_06117_),
    .A(_06100_),
    .X(_06118_));
 sg13g2_xnor2_1 _14012_ (.Y(_06119_),
    .A(_06096_),
    .B(_06118_));
 sg13g2_nand3_1 _14013_ (.B(_05951_),
    .C(_05974_),
    .A(_05949_),
    .Y(_06120_));
 sg13g2_a21oi_1 _14014_ (.A1(_05949_),
    .A2(_05951_),
    .Y(_06121_),
    .B1(_05974_));
 sg13g2_a21oi_2 _14015_ (.B1(_06121_),
    .Y(_06122_),
    .A2(_06120_),
    .A1(_05957_));
 sg13g2_nand2_1 _14016_ (.Y(_06124_),
    .A(net199),
    .B(net136));
 sg13g2_and2_1 _14017_ (.A(_06124_),
    .B(_05831_),
    .X(_06125_));
 sg13g2_a21oi_1 _14018_ (.A1(_05825_),
    .A2(_05827_),
    .Y(_06126_),
    .B1(_06125_));
 sg13g2_nand2_1 _14019_ (.Y(_06127_),
    .A(net249),
    .B(net170));
 sg13g2_nand2_1 _14020_ (.Y(_06128_),
    .A(net213),
    .B(_02770_));
 sg13g2_nand2_1 _14021_ (.Y(_06129_),
    .A(net201),
    .B(net114));
 sg13g2_xnor2_1 _14022_ (.Y(_06130_),
    .A(_06128_),
    .B(_06129_));
 sg13g2_xnor2_1 _14023_ (.Y(_06131_),
    .A(_06127_),
    .B(_06130_));
 sg13g2_nand2_1 _14024_ (.Y(_06132_),
    .A(_00333_),
    .B(net136));
 sg13g2_xor2_1 _14025_ (.B(_06132_),
    .A(_06131_),
    .X(_06133_));
 sg13g2_xnor2_1 _14026_ (.Y(_06135_),
    .A(_06126_),
    .B(_06133_));
 sg13g2_inv_1 _14027_ (.Y(_06136_),
    .A(_06135_));
 sg13g2_nor2_1 _14028_ (.A(_05967_),
    .B(_05972_),
    .Y(_06137_));
 sg13g2_nor2_1 _14029_ (.A(_05963_),
    .B(_06137_),
    .Y(_06138_));
 sg13g2_a21oi_1 _14030_ (.A1(_05967_),
    .A2(_05972_),
    .Y(_06139_),
    .B1(_06138_));
 sg13g2_xor2_1 _14031_ (.B(net145),
    .A(net199),
    .X(_06140_));
 sg13g2_nor3_2 _14032_ (.A(_04563_),
    .B(net147),
    .C(_06140_),
    .Y(_06141_));
 sg13g2_xnor2_1 _14033_ (.Y(_06142_),
    .A(_06139_),
    .B(_06141_));
 sg13g2_xnor2_1 _14034_ (.Y(_06143_),
    .A(_06136_),
    .B(_06142_));
 sg13g2_xnor2_1 _14035_ (.Y(_06144_),
    .A(_06122_),
    .B(_06143_));
 sg13g2_xor2_1 _14036_ (.B(_06144_),
    .A(_06119_),
    .X(_06146_));
 sg13g2_inv_1 _14037_ (.Y(_06147_),
    .A(_05839_));
 sg13g2_nand2_1 _14038_ (.Y(_06148_),
    .A(_05842_),
    .B(_05843_));
 sg13g2_nor2_1 _14039_ (.A(_06148_),
    .B(_05976_),
    .Y(_06149_));
 sg13g2_xnor2_1 _14040_ (.Y(_06150_),
    .A(_05953_),
    .B(_05975_));
 sg13g2_o21ai_1 _14041_ (.B1(_05838_),
    .Y(_06151_),
    .A1(_06150_),
    .A2(_06147_));
 sg13g2_nor2_1 _14042_ (.A(_06150_),
    .B(_05838_),
    .Y(_06152_));
 sg13g2_a221oi_1 _14043_ (.B2(_06148_),
    .C1(_06152_),
    .B1(_06151_),
    .A1(_06147_),
    .Y(_06153_),
    .A2(_06149_));
 sg13g2_xor2_1 _14044_ (.B(_06153_),
    .A(_06146_),
    .X(_06154_));
 sg13g2_xor2_1 _14045_ (.B(_06026_),
    .A(_06001_),
    .X(_06155_));
 sg13g2_xnor2_1 _14046_ (.Y(_06157_),
    .A(_05983_),
    .B(_06155_));
 sg13g2_xor2_1 _14047_ (.B(_05987_),
    .A(_05986_),
    .X(_06158_));
 sg13g2_xnor2_1 _14048_ (.Y(_06159_),
    .A(_05989_),
    .B(_06158_));
 sg13g2_nand2_1 _14049_ (.Y(_06160_),
    .A(net250),
    .B(_02282_));
 sg13g2_nand2_1 _14050_ (.Y(_06161_),
    .A(net215),
    .B(_02303_));
 sg13g2_nand2_1 _14051_ (.Y(_06162_),
    .A(net216),
    .B(net172));
 sg13g2_a21o_1 _14052_ (.A2(_06161_),
    .A1(_06160_),
    .B1(_06162_),
    .X(_06163_));
 sg13g2_o21ai_1 _14053_ (.B1(_06163_),
    .Y(_06164_),
    .A1(_06160_),
    .A2(_06161_));
 sg13g2_buf_1 _14054_ (.A(_06164_),
    .X(_06165_));
 sg13g2_nand2_1 _14055_ (.Y(_06166_),
    .A(_00814_),
    .B(_02743_));
 sg13g2_xnor2_1 _14056_ (.Y(_06168_),
    .A(_06165_),
    .B(_06166_));
 sg13g2_xnor2_1 _14057_ (.Y(_06169_),
    .A(_06159_),
    .B(_06168_));
 sg13g2_or2_1 _14058_ (.X(_06170_),
    .B(_06014_),
    .A(_06009_));
 sg13g2_xnor2_1 _14059_ (.Y(_06171_),
    .A(_06017_),
    .B(_06020_));
 sg13g2_xnor2_1 _14060_ (.Y(_06172_),
    .A(_06170_),
    .B(_06171_));
 sg13g2_or2_1 _14061_ (.X(_06173_),
    .B(_05467_),
    .A(_05430_));
 sg13g2_buf_1 _14062_ (.A(_06173_),
    .X(_06174_));
 sg13g2_a21o_1 _14063_ (.A2(_05467_),
    .A1(_05430_),
    .B1(_05432_),
    .X(_06175_));
 sg13g2_buf_1 _14064_ (.A(_06175_),
    .X(_06176_));
 sg13g2_xor2_1 _14065_ (.B(_06161_),
    .A(_06160_),
    .X(_06177_));
 sg13g2_xnor2_1 _14066_ (.Y(_06179_),
    .A(_06162_),
    .B(_06177_));
 sg13g2_inv_1 _14067_ (.Y(_06180_),
    .A(_06179_));
 sg13g2_nand3_1 _14068_ (.B(_06176_),
    .C(_06180_),
    .A(_06174_),
    .Y(_06181_));
 sg13g2_a21oi_1 _14069_ (.A1(_06174_),
    .A2(_06176_),
    .Y(_06182_),
    .B1(_06180_));
 sg13g2_a21oi_1 _14070_ (.A1(_06172_),
    .A2(_06181_),
    .Y(_06183_),
    .B1(_06182_));
 sg13g2_or2_1 _14071_ (.X(_06184_),
    .B(_06183_),
    .A(_06169_));
 sg13g2_xnor2_1 _14072_ (.Y(_06185_),
    .A(_06022_),
    .B(_06007_));
 sg13g2_xnor2_1 _14073_ (.Y(_06186_),
    .A(_06005_),
    .B(_06185_));
 sg13g2_and2_1 _14074_ (.A(_06169_),
    .B(_06183_),
    .X(_06187_));
 sg13g2_a21o_1 _14075_ (.A2(_06186_),
    .A1(_06184_),
    .B1(_06187_),
    .X(_06188_));
 sg13g2_buf_1 _14076_ (.A(_06188_),
    .X(_06190_));
 sg13g2_nand2_1 _14077_ (.Y(_06191_),
    .A(_00289_),
    .B(net136));
 sg13g2_nor2_1 _14078_ (.A(_06165_),
    .B(_06159_),
    .Y(_06192_));
 sg13g2_nand2_1 _14079_ (.Y(_06193_),
    .A(_06165_),
    .B(_06159_));
 sg13g2_o21ai_1 _14080_ (.B1(_06193_),
    .Y(_06194_),
    .A1(_06166_),
    .A2(_06192_));
 sg13g2_buf_1 _14081_ (.A(_06194_),
    .X(_06195_));
 sg13g2_nand2b_1 _14082_ (.Y(_06196_),
    .B(_06195_),
    .A_N(_06191_));
 sg13g2_nor3_1 _14083_ (.A(_06157_),
    .B(_06190_),
    .C(_06196_),
    .Y(_06197_));
 sg13g2_xnor2_1 _14084_ (.Y(_06198_),
    .A(_06191_),
    .B(_06195_));
 sg13g2_xnor2_1 _14085_ (.Y(_06199_),
    .A(_06190_),
    .B(_06198_));
 sg13g2_xnor2_1 _14086_ (.Y(_06201_),
    .A(_06157_),
    .B(_06199_));
 sg13g2_inv_1 _14087_ (.Y(_06202_),
    .A(_06201_));
 sg13g2_xor2_1 _14088_ (.B(_06183_),
    .A(_06169_),
    .X(_06203_));
 sg13g2_xnor2_1 _14089_ (.Y(_06204_),
    .A(_06186_),
    .B(_06203_));
 sg13g2_nand2_1 _14090_ (.Y(_06205_),
    .A(net268),
    .B(_02290_));
 sg13g2_nand2_1 _14091_ (.Y(_06206_),
    .A(net214),
    .B(_02739_));
 sg13g2_xor2_1 _14092_ (.B(_06206_),
    .A(_06205_),
    .X(_06207_));
 sg13g2_buf_1 _14093_ (.A(_06207_),
    .X(_06208_));
 sg13g2_nor2b_1 _14094_ (.A(_05474_),
    .B_N(_05479_),
    .Y(_06209_));
 sg13g2_nand2b_1 _14095_ (.Y(_06210_),
    .B(_05474_),
    .A_N(_05479_));
 sg13g2_o21ai_1 _14096_ (.B1(_06210_),
    .Y(_06212_),
    .A1(_05469_),
    .A2(_06209_));
 sg13g2_buf_1 _14097_ (.A(_06212_),
    .X(_06213_));
 sg13g2_nand2_1 _14098_ (.Y(_06214_),
    .A(_05471_),
    .B(_05472_));
 sg13g2_o21ai_1 _14099_ (.B1(_05470_),
    .Y(_06215_),
    .A1(_05471_),
    .A2(_05472_));
 sg13g2_nand2_1 _14100_ (.Y(_06216_),
    .A(_06214_),
    .B(_06215_));
 sg13g2_nand2_1 _14101_ (.Y(_06217_),
    .A(_06213_),
    .B(_06216_));
 sg13g2_nor2_1 _14102_ (.A(_06213_),
    .B(_06216_),
    .Y(_06218_));
 sg13g2_a21o_1 _14103_ (.A2(_06217_),
    .A1(_06208_),
    .B1(_06218_),
    .X(_06219_));
 sg13g2_and2_1 _14104_ (.A(_06204_),
    .B(_06219_),
    .X(_06220_));
 sg13g2_buf_1 _14105_ (.A(_06220_),
    .X(_06221_));
 sg13g2_o21ai_1 _14106_ (.B1(_06208_),
    .Y(_06223_),
    .A1(_06204_),
    .A2(_06218_));
 sg13g2_nand2_1 _14107_ (.Y(_06224_),
    .A(_06204_),
    .B(_06217_));
 sg13g2_and3_1 _14108_ (.X(_06225_),
    .A(_06174_),
    .B(_06176_),
    .C(_06180_));
 sg13g2_o21ai_1 _14109_ (.B1(_06172_),
    .Y(_06226_),
    .A1(_06182_),
    .A2(_06225_));
 sg13g2_or3_1 _14110_ (.A(_06172_),
    .B(_06182_),
    .C(_06225_),
    .X(_06227_));
 sg13g2_and2_1 _14111_ (.A(_06226_),
    .B(_06227_),
    .X(_06228_));
 sg13g2_buf_1 _14112_ (.A(_06228_),
    .X(_06229_));
 sg13g2_a21oi_1 _14113_ (.A1(_06223_),
    .A2(_06224_),
    .Y(_06230_),
    .B1(_06229_));
 sg13g2_nor2_1 _14114_ (.A(net195),
    .B(_03018_),
    .Y(_06231_));
 sg13g2_nand2_1 _14115_ (.Y(_06232_),
    .A(_05481_),
    .B(_05494_));
 sg13g2_nor2_1 _14116_ (.A(_05481_),
    .B(_05494_),
    .Y(_06234_));
 sg13g2_a21oi_1 _14117_ (.A1(_05491_),
    .A2(_06232_),
    .Y(_06235_),
    .B1(_06234_));
 sg13g2_and2_1 _14118_ (.A(_06214_),
    .B(_06215_),
    .X(_06236_));
 sg13g2_xnor2_1 _14119_ (.Y(_06237_),
    .A(_06208_),
    .B(_06236_));
 sg13g2_xor2_1 _14120_ (.B(_06237_),
    .A(_06213_),
    .X(_06238_));
 sg13g2_xnor2_1 _14121_ (.Y(_06239_),
    .A(_06229_),
    .B(_06238_));
 sg13g2_a21oi_1 _14122_ (.A1(_05392_),
    .A2(_05396_),
    .Y(_06240_),
    .B1(_05496_));
 sg13g2_a221oi_1 _14123_ (.B2(_06239_),
    .C1(_06240_),
    .B1(_06235_),
    .A1(_06231_),
    .Y(_06241_),
    .A2(_05485_));
 sg13g2_nand2_1 _14124_ (.Y(_06242_),
    .A(_05491_),
    .B(_06232_));
 sg13g2_or2_1 _14125_ (.X(_06243_),
    .B(_05494_),
    .A(_05481_));
 sg13g2_and2_1 _14126_ (.A(_06231_),
    .B(_05485_),
    .X(_06245_));
 sg13g2_a221oi_1 _14127_ (.B2(_06240_),
    .C1(_06239_),
    .B1(_06245_),
    .A1(_06242_),
    .Y(_06246_),
    .A2(_06243_));
 sg13g2_nor2b_1 _14128_ (.A(_06208_),
    .B_N(_06213_),
    .Y(_06247_));
 sg13g2_a21oi_1 _14129_ (.A1(_06208_),
    .A2(_06217_),
    .Y(_06248_),
    .B1(_06218_));
 sg13g2_nand2_1 _14130_ (.Y(_06249_),
    .A(_06208_),
    .B(_06236_));
 sg13g2_or2_1 _14131_ (.X(_06250_),
    .B(_06249_),
    .A(_06213_));
 sg13g2_a21oi_1 _14132_ (.A1(_06226_),
    .A2(_06227_),
    .Y(_06251_),
    .B1(_06250_));
 sg13g2_a221oi_1 _14133_ (.B2(_06229_),
    .C1(_06251_),
    .B1(_06248_),
    .A1(_06216_),
    .Y(_06252_),
    .A2(_06247_));
 sg13g2_xnor2_1 _14134_ (.Y(_06253_),
    .A(_06204_),
    .B(_06252_));
 sg13g2_nor3_1 _14135_ (.A(_06241_),
    .B(_06246_),
    .C(_06253_),
    .Y(_06254_));
 sg13g2_o21ai_1 _14136_ (.B1(_06254_),
    .Y(_06256_),
    .A1(_06221_),
    .A2(_06230_));
 sg13g2_buf_1 _14137_ (.A(_06256_),
    .X(_06257_));
 sg13g2_nor3_1 _14138_ (.A(_06221_),
    .B(_06230_),
    .C(_06254_),
    .Y(_06258_));
 sg13g2_a21o_1 _14139_ (.A2(_06257_),
    .A1(_06202_),
    .B1(_06258_),
    .X(_06259_));
 sg13g2_buf_1 _14140_ (.A(_06259_),
    .X(_06260_));
 sg13g2_xnor2_1 _14141_ (.Y(_06261_),
    .A(_06043_),
    .B(_06033_));
 sg13g2_xnor2_1 _14142_ (.Y(_06262_),
    .A(_06030_),
    .B(_06261_));
 sg13g2_xnor2_1 _14143_ (.Y(_06263_),
    .A(_06039_),
    .B(_06262_));
 sg13g2_nand3b_1 _14144_ (.B(_06260_),
    .C(_06263_),
    .Y(_06264_),
    .A_N(_06197_));
 sg13g2_a21oi_1 _14145_ (.A1(net157),
    .A2(net136),
    .Y(_06265_),
    .B1(_06195_));
 sg13g2_a21o_1 _14146_ (.A2(_06196_),
    .A1(_06190_),
    .B1(_06265_),
    .X(_06267_));
 sg13g2_and2_1 _14147_ (.A(_06190_),
    .B(_06265_),
    .X(_06268_));
 sg13g2_a21o_1 _14148_ (.A2(_06267_),
    .A1(_06157_),
    .B1(_06268_),
    .X(_06269_));
 sg13g2_o21ai_1 _14149_ (.B1(_06269_),
    .Y(_06270_),
    .A1(_06260_),
    .A2(_06263_));
 sg13g2_o21ai_1 _14150_ (.B1(_06039_),
    .Y(_06271_),
    .A1(_06045_),
    .A2(_06048_));
 sg13g2_or3_1 _14151_ (.A(_06039_),
    .B(_06043_),
    .C(_06034_),
    .X(_06272_));
 sg13g2_nand2_1 _14152_ (.Y(_06273_),
    .A(_06043_),
    .B(_06045_));
 sg13g2_nand3_1 _14153_ (.B(_06272_),
    .C(_06273_),
    .A(_06271_),
    .Y(_06274_));
 sg13g2_nand3_1 _14154_ (.B(_05981_),
    .C(_06274_),
    .A(_05978_),
    .Y(_06275_));
 sg13g2_a21o_1 _14155_ (.A2(_05981_),
    .A1(_05978_),
    .B1(_06274_),
    .X(_06276_));
 sg13g2_nand4_1 _14156_ (.B(_06270_),
    .C(_06275_),
    .A(_06264_),
    .Y(_06278_),
    .D(_06276_));
 sg13g2_o21ai_1 _14157_ (.B1(_06278_),
    .Y(_06279_),
    .A1(_06052_),
    .A2(_06154_));
 sg13g2_nand2_1 _14158_ (.Y(_06280_),
    .A(_06052_),
    .B(_06154_));
 sg13g2_nand2_1 _14159_ (.Y(_06281_),
    .A(_06279_),
    .B(_06280_));
 sg13g2_nand2_1 _14160_ (.Y(_06282_),
    .A(_05839_),
    .B(_06146_));
 sg13g2_o21ai_1 _14161_ (.B1(_05838_),
    .Y(_06283_),
    .A1(_05798_),
    .A2(_05821_));
 sg13g2_a21oi_1 _14162_ (.A1(_06151_),
    .A2(_06283_),
    .Y(_06284_),
    .B1(_06146_));
 sg13g2_a21oi_1 _14163_ (.A1(_06149_),
    .A2(_06282_),
    .Y(_06285_),
    .B1(_06284_));
 sg13g2_a21o_1 _14164_ (.A2(_06075_),
    .A1(_06073_),
    .B1(_06085_),
    .X(_06286_));
 sg13g2_and3_1 _14165_ (.X(_06287_),
    .A(_06073_),
    .B(_06075_),
    .C(_06085_));
 sg13g2_a21oi_1 _14166_ (.A1(_06086_),
    .A2(_06286_),
    .Y(_06289_),
    .B1(_06287_));
 sg13g2_nor2_1 _14167_ (.A(net252),
    .B(net191),
    .Y(_06290_));
 sg13g2_buf_1 _14168_ (.A(_06290_),
    .X(_06291_));
 sg13g2_buf_1 _14169_ (.A(_06291_),
    .X(_06292_));
 sg13g2_nand2_1 _14170_ (.Y(_06293_),
    .A(net134),
    .B(net292));
 sg13g2_nand2_1 _14171_ (.Y(_06294_),
    .A(net163),
    .B(_01489_));
 sg13g2_xor2_1 _14172_ (.B(_06294_),
    .A(_06293_),
    .X(_06295_));
 sg13g2_xnor2_1 _14173_ (.Y(_06296_),
    .A(net97),
    .B(_06295_));
 sg13g2_inv_1 _14174_ (.Y(_06297_),
    .A(_06069_));
 sg13g2_and2_1 _14175_ (.A(_06297_),
    .B(_06075_),
    .X(_06298_));
 sg13g2_buf_1 _14176_ (.A(_06298_),
    .X(_06300_));
 sg13g2_nor2b_1 _14177_ (.A(_06083_),
    .B_N(_06084_),
    .Y(_06301_));
 sg13g2_nor2_1 _14178_ (.A(_06081_),
    .B(_06301_),
    .Y(_06302_));
 sg13g2_buf_2 _14179_ (.A(_06302_),
    .X(_06303_));
 sg13g2_xnor2_1 _14180_ (.Y(_06304_),
    .A(net267),
    .B(_06303_));
 sg13g2_xnor2_1 _14181_ (.Y(_06305_),
    .A(_06300_),
    .B(_06304_));
 sg13g2_xnor2_1 _14182_ (.Y(_06306_),
    .A(_06296_),
    .B(_06305_));
 sg13g2_xnor2_1 _14183_ (.Y(_06307_),
    .A(_06289_),
    .B(_06306_));
 sg13g2_o21ai_1 _14184_ (.B1(_06094_),
    .Y(_06308_),
    .A1(_06053_),
    .A2(_06054_));
 sg13g2_nor3_1 _14185_ (.A(_06053_),
    .B(_06054_),
    .C(_06094_),
    .Y(_06309_));
 sg13g2_a21oi_2 _14186_ (.B1(_06309_),
    .Y(_06311_),
    .A2(_06308_),
    .A1(_06088_));
 sg13g2_nand2_1 _14187_ (.Y(_06312_),
    .A(net268),
    .B(_02013_));
 sg13g2_nand2_1 _14188_ (.Y(_06313_),
    .A(net162),
    .B(net177));
 sg13g2_nand2_1 _14189_ (.Y(_06314_),
    .A(net214),
    .B(_02007_));
 sg13g2_xnor2_1 _14190_ (.Y(_06315_),
    .A(_06313_),
    .B(_06314_));
 sg13g2_xnor2_1 _14191_ (.Y(_06316_),
    .A(_06312_),
    .B(_06315_));
 sg13g2_and2_1 _14192_ (.A(_06091_),
    .B(_06092_),
    .X(_06317_));
 sg13g2_or2_1 _14193_ (.X(_06318_),
    .B(_06092_),
    .A(_06091_));
 sg13g2_o21ai_1 _14194_ (.B1(_06318_),
    .Y(_06319_),
    .A1(_06089_),
    .A2(_06317_));
 sg13g2_buf_1 _14195_ (.A(_06319_),
    .X(_06320_));
 sg13g2_and2_1 _14196_ (.A(_06103_),
    .B(_06104_),
    .X(_06322_));
 sg13g2_or2_1 _14197_ (.X(_06323_),
    .B(_06104_),
    .A(_06103_));
 sg13g2_o21ai_1 _14198_ (.B1(_06323_),
    .Y(_06324_),
    .A1(_06102_),
    .A2(_06322_));
 sg13g2_buf_1 _14199_ (.A(_06324_),
    .X(_06325_));
 sg13g2_xor2_1 _14200_ (.B(_06325_),
    .A(_06320_),
    .X(_06326_));
 sg13g2_xnor2_1 _14201_ (.Y(_06327_),
    .A(_06316_),
    .B(_06326_));
 sg13g2_xor2_1 _14202_ (.B(_06327_),
    .A(_06311_),
    .X(_06328_));
 sg13g2_xnor2_1 _14203_ (.Y(_06329_),
    .A(_06307_),
    .B(_06328_));
 sg13g2_nand2_1 _14204_ (.Y(_06330_),
    .A(net213),
    .B(net114));
 sg13g2_nand2_1 _14205_ (.Y(_06331_),
    .A(net212),
    .B(net178));
 sg13g2_nand2_1 _14206_ (.Y(_06333_),
    .A(net269),
    .B(net144));
 sg13g2_xnor2_1 _14207_ (.Y(_06334_),
    .A(_06331_),
    .B(_06333_));
 sg13g2_xnor2_1 _14208_ (.Y(_06335_),
    .A(_06330_),
    .B(_06334_));
 sg13g2_and2_1 _14209_ (.A(_06128_),
    .B(_06129_),
    .X(_06336_));
 sg13g2_or2_1 _14210_ (.X(_06337_),
    .B(_06129_),
    .A(_06128_));
 sg13g2_o21ai_1 _14211_ (.B1(_06337_),
    .Y(_06338_),
    .A1(_06127_),
    .A2(_06336_));
 sg13g2_nand2_1 _14212_ (.Y(_06339_),
    .A(net203),
    .B(net169));
 sg13g2_nand2_1 _14213_ (.Y(_06340_),
    .A(net249),
    .B(_02770_));
 sg13g2_nand2_1 _14214_ (.Y(_06341_),
    .A(net306),
    .B(net170));
 sg13g2_xnor2_1 _14215_ (.Y(_06342_),
    .A(_06340_),
    .B(_06341_));
 sg13g2_xnor2_1 _14216_ (.Y(_06344_),
    .A(_06339_),
    .B(_06342_));
 sg13g2_xor2_1 _14217_ (.B(_06344_),
    .A(_06338_),
    .X(_06345_));
 sg13g2_xnor2_1 _14218_ (.Y(_06346_),
    .A(_06335_),
    .B(_06345_));
 sg13g2_nand2_1 _14219_ (.Y(_06347_),
    .A(_06110_),
    .B(_06115_));
 sg13g2_nor2_1 _14220_ (.A(_06110_),
    .B(_06115_),
    .Y(_06348_));
 sg13g2_or2_1 _14221_ (.X(_06349_),
    .B(_06348_),
    .A(_06106_));
 sg13g2_nand2b_1 _14222_ (.Y(_06350_),
    .B(_06126_),
    .A_N(_06131_));
 sg13g2_nand2b_1 _14223_ (.Y(_06351_),
    .B(_06131_),
    .A_N(_06126_));
 sg13g2_nand2b_1 _14224_ (.Y(_06352_),
    .B(_06351_),
    .A_N(_06132_));
 sg13g2_and4_1 _14225_ (.A(_06347_),
    .B(_06349_),
    .C(_06350_),
    .D(_06352_),
    .X(_06353_));
 sg13g2_a22oi_1 _14226_ (.Y(_06355_),
    .B1(_06350_),
    .B2(_06352_),
    .A2(_06349_),
    .A1(_06347_));
 sg13g2_nor2_1 _14227_ (.A(_06353_),
    .B(_06355_),
    .Y(_06356_));
 sg13g2_xnor2_1 _14228_ (.Y(_06357_),
    .A(_06346_),
    .B(_06356_));
 sg13g2_or2_1 _14229_ (.X(_06358_),
    .B(_06117_),
    .A(_06100_));
 sg13g2_and2_1 _14230_ (.A(_06100_),
    .B(_06117_),
    .X(_06359_));
 sg13g2_a21o_1 _14231_ (.A2(_06358_),
    .A1(_06096_),
    .B1(_06359_),
    .X(_06360_));
 sg13g2_xnor2_1 _14232_ (.Y(_06361_),
    .A(_06357_),
    .B(_06360_));
 sg13g2_xnor2_1 _14233_ (.Y(_06362_),
    .A(_06329_),
    .B(_06361_));
 sg13g2_nand2_1 _14234_ (.Y(_06363_),
    .A(_06122_),
    .B(_06143_));
 sg13g2_nor2_1 _14235_ (.A(_06122_),
    .B(_06143_),
    .Y(_06364_));
 sg13g2_a21oi_1 _14236_ (.A1(_06119_),
    .A2(_06363_),
    .Y(_06366_),
    .B1(_06364_));
 sg13g2_inv_1 _14237_ (.Y(_06367_),
    .A(_06141_));
 sg13g2_a21oi_1 _14238_ (.A1(_06135_),
    .A2(_06367_),
    .Y(_06368_),
    .B1(_06139_));
 sg13g2_a21oi_1 _14239_ (.A1(_06136_),
    .A2(_06141_),
    .Y(_06369_),
    .B1(_06368_));
 sg13g2_xor2_1 _14240_ (.B(_06369_),
    .A(_06366_),
    .X(_06370_));
 sg13g2_xnor2_1 _14241_ (.Y(_06371_),
    .A(_06362_),
    .B(_06370_));
 sg13g2_xnor2_1 _14242_ (.Y(_06372_),
    .A(_06285_),
    .B(_06371_));
 sg13g2_xnor2_1 _14243_ (.Y(_06373_),
    .A(_06281_),
    .B(_06372_));
 sg13g2_nand2_1 _14244_ (.Y(_06374_),
    .A(_06264_),
    .B(_06270_));
 sg13g2_nand2_1 _14245_ (.Y(_06375_),
    .A(_06275_),
    .B(_06276_));
 sg13g2_xnor2_1 _14246_ (.Y(_06377_),
    .A(_06374_),
    .B(_06375_));
 sg13g2_or3_1 _14247_ (.A(_06221_),
    .B(_06230_),
    .C(_06254_),
    .X(_06378_));
 sg13g2_and3_1 _14248_ (.X(_06379_),
    .A(_06202_),
    .B(_06257_),
    .C(_06378_));
 sg13g2_buf_1 _14249_ (.A(_06379_),
    .X(_06380_));
 sg13g2_a21oi_1 _14250_ (.A1(_06257_),
    .A2(_06378_),
    .Y(_06381_),
    .B1(_06202_));
 sg13g2_nor3_1 _14251_ (.A(_04112_),
    .B(_06380_),
    .C(_06381_),
    .Y(_06382_));
 sg13g2_nor2_1 _14252_ (.A(_06241_),
    .B(_06246_),
    .Y(_06383_));
 sg13g2_xnor2_1 _14253_ (.Y(_06384_),
    .A(_06383_),
    .B(_06253_));
 sg13g2_and2_1 _14254_ (.A(_04046_),
    .B(_05499_),
    .X(_06385_));
 sg13g2_buf_1 _14255_ (.A(_06385_),
    .X(_06386_));
 sg13g2_xor2_1 _14256_ (.B(_06245_),
    .A(_06235_),
    .X(_06388_));
 sg13g2_xnor2_1 _14257_ (.Y(_06389_),
    .A(_06240_),
    .B(_06388_));
 sg13g2_xnor2_1 _14258_ (.Y(_06390_),
    .A(_06239_),
    .B(_06389_));
 sg13g2_or2_1 _14259_ (.X(_06391_),
    .B(_06390_),
    .A(_06386_));
 sg13g2_a21o_1 _14260_ (.A2(_06390_),
    .A1(_06386_),
    .B1(_04105_),
    .X(_06392_));
 sg13g2_and3_1 _14261_ (.X(_06393_),
    .A(_06384_),
    .B(_06391_),
    .C(_06392_));
 sg13g2_a21o_1 _14262_ (.A2(_06392_),
    .A1(_06391_),
    .B1(_06384_),
    .X(_06394_));
 sg13g2_o21ai_1 _14263_ (.B1(_06394_),
    .Y(_06395_),
    .A1(_04108_),
    .A2(_06393_));
 sg13g2_o21ai_1 _14264_ (.B1(_04112_),
    .Y(_06396_),
    .A1(_06380_),
    .A2(_06381_));
 sg13g2_o21ai_1 _14265_ (.B1(_06396_),
    .Y(_06397_),
    .A1(_06382_),
    .A2(_06395_));
 sg13g2_nor2_1 _14266_ (.A(_06197_),
    .B(_06269_),
    .Y(_06399_));
 sg13g2_xor2_1 _14267_ (.B(_06399_),
    .A(_06263_),
    .X(_06400_));
 sg13g2_xnor2_1 _14268_ (.Y(_06401_),
    .A(_06260_),
    .B(_06400_));
 sg13g2_xnor2_1 _14269_ (.Y(_06402_),
    .A(_04063_),
    .B(_06401_));
 sg13g2_nor2_1 _14270_ (.A(_00018_),
    .B(_06401_),
    .Y(_06403_));
 sg13g2_a21oi_2 _14271_ (.B1(_06403_),
    .Y(_06404_),
    .A2(_06402_),
    .A1(_06397_));
 sg13g2_nor2_1 _14272_ (.A(_06377_),
    .B(_06404_),
    .Y(_06405_));
 sg13g2_nand2_1 _14273_ (.Y(_06406_),
    .A(_06377_),
    .B(_06404_));
 sg13g2_o21ai_1 _14274_ (.B1(_06406_),
    .Y(_06407_),
    .A1(net317),
    .A2(_06405_));
 sg13g2_xnor2_1 _14275_ (.Y(_06408_),
    .A(_06278_),
    .B(_06154_));
 sg13g2_xor2_1 _14276_ (.B(_06408_),
    .A(_06052_),
    .X(_06410_));
 sg13g2_xnor2_1 _14277_ (.Y(_06411_),
    .A(_04064_),
    .B(_06410_));
 sg13g2_nand2b_1 _14278_ (.Y(_06412_),
    .B(_06410_),
    .A_N(_00019_));
 sg13g2_o21ai_1 _14279_ (.B1(_06412_),
    .Y(_06413_),
    .A1(_06407_),
    .A2(_06411_));
 sg13g2_buf_1 _14280_ (.A(_06413_),
    .X(_06414_));
 sg13g2_o21ai_1 _14281_ (.B1(_04059_),
    .Y(_06415_),
    .A1(_06373_),
    .A2(_06414_));
 sg13g2_nand2_1 _14282_ (.Y(_06416_),
    .A(_06373_),
    .B(_06414_));
 sg13g2_nand2_1 _14283_ (.Y(_06417_),
    .A(_06329_),
    .B(_06357_));
 sg13g2_nor2_1 _14284_ (.A(_06329_),
    .B(_06357_),
    .Y(_06418_));
 sg13g2_a21o_1 _14285_ (.A2(_06417_),
    .A1(_06360_),
    .B1(_06418_),
    .X(_06419_));
 sg13g2_buf_1 _14286_ (.A(_06419_),
    .X(_06421_));
 sg13g2_nor2_1 _14287_ (.A(_06346_),
    .B(_06353_),
    .Y(_06422_));
 sg13g2_nor2_1 _14288_ (.A(_06355_),
    .B(_06422_),
    .Y(_06423_));
 sg13g2_nand2_1 _14289_ (.Y(_06424_),
    .A(_06311_),
    .B(_06327_));
 sg13g2_nor2_1 _14290_ (.A(_06311_),
    .B(_06327_),
    .Y(_06425_));
 sg13g2_a21oi_1 _14291_ (.A1(_06307_),
    .A2(_06424_),
    .Y(_06426_),
    .B1(_06425_));
 sg13g2_or2_1 _14292_ (.X(_06427_),
    .B(_06296_),
    .A(_06289_));
 sg13g2_buf_2 _14293_ (.A(_06427_),
    .X(_06428_));
 sg13g2_nand2_1 _14294_ (.Y(_06429_),
    .A(net249),
    .B(net114));
 sg13g2_nand2_1 _14295_ (.Y(_06430_),
    .A(net269),
    .B(net178));
 sg13g2_nand2_1 _14296_ (.Y(_06432_),
    .A(net213),
    .B(_03213_));
 sg13g2_xnor2_1 _14297_ (.Y(_06433_),
    .A(_06430_),
    .B(_06432_));
 sg13g2_xnor2_1 _14298_ (.Y(_06434_),
    .A(_06429_),
    .B(_06433_));
 sg13g2_and2_1 _14299_ (.A(_06331_),
    .B(_06333_),
    .X(_06435_));
 sg13g2_or2_1 _14300_ (.X(_06436_),
    .B(_06333_),
    .A(_06331_));
 sg13g2_o21ai_1 _14301_ (.B1(_06436_),
    .Y(_06437_),
    .A1(_06330_),
    .A2(_06435_));
 sg13g2_nand2_1 _14302_ (.Y(_06438_),
    .A(net203),
    .B(_02742_));
 sg13g2_nand2_1 _14303_ (.Y(_06439_),
    .A(net306),
    .B(net145));
 sg13g2_xnor2_1 _14304_ (.Y(_06440_),
    .A(_06438_),
    .B(_06439_));
 sg13g2_xnor2_1 _14305_ (.Y(_06441_),
    .A(_06437_),
    .B(_06440_));
 sg13g2_xnor2_1 _14306_ (.Y(_06443_),
    .A(_06434_),
    .B(_06441_));
 sg13g2_nand2_1 _14307_ (.Y(_06444_),
    .A(_06320_),
    .B(_06325_));
 sg13g2_nor2_1 _14308_ (.A(_06320_),
    .B(_06325_),
    .Y(_06445_));
 sg13g2_a21oi_1 _14309_ (.A1(_06316_),
    .A2(_06444_),
    .Y(_06446_),
    .B1(_06445_));
 sg13g2_nor2_1 _14310_ (.A(_06335_),
    .B(_06344_),
    .Y(_06447_));
 sg13g2_nor2_1 _14311_ (.A(_06338_),
    .B(_06447_),
    .Y(_06448_));
 sg13g2_a21oi_2 _14312_ (.B1(_06448_),
    .Y(_06449_),
    .A2(_06344_),
    .A1(_06335_));
 sg13g2_xnor2_1 _14313_ (.Y(_06450_),
    .A(_06446_),
    .B(_06449_));
 sg13g2_xor2_1 _14314_ (.B(_06450_),
    .A(_06443_),
    .X(_06451_));
 sg13g2_inv_1 _14315_ (.Y(_06452_),
    .A(_06451_));
 sg13g2_a21o_1 _14316_ (.A2(_06296_),
    .A1(_06289_),
    .B1(_06305_),
    .X(_06454_));
 sg13g2_buf_2 _14317_ (.A(_06454_),
    .X(_06455_));
 sg13g2_nand2_1 _14318_ (.Y(_06456_),
    .A(net212),
    .B(net152));
 sg13g2_nand2_1 _14319_ (.Y(_06457_),
    .A(net133),
    .B(net177));
 sg13g2_nand2_1 _14320_ (.Y(_06458_),
    .A(net217),
    .B(net180));
 sg13g2_xnor2_1 _14321_ (.Y(_06459_),
    .A(_06457_),
    .B(_06458_));
 sg13g2_xnor2_1 _14322_ (.Y(_06460_),
    .A(_06456_),
    .B(_06459_));
 sg13g2_nor2b_1 _14323_ (.A(_06291_),
    .B_N(_06293_),
    .Y(_06461_));
 sg13g2_nand3_1 _14324_ (.B(net231),
    .C(_06291_),
    .A(net134),
    .Y(_06462_));
 sg13g2_o21ai_1 _14325_ (.B1(_06462_),
    .Y(_06463_),
    .A1(_06294_),
    .A2(_06461_));
 sg13g2_buf_1 _14326_ (.A(_06463_),
    .X(_06465_));
 sg13g2_and2_1 _14327_ (.A(_06313_),
    .B(_06314_),
    .X(_06466_));
 sg13g2_or2_1 _14328_ (.X(_06467_),
    .B(_06314_),
    .A(_06313_));
 sg13g2_o21ai_1 _14329_ (.B1(_06467_),
    .Y(_06468_),
    .A1(_06312_),
    .A2(_06466_));
 sg13g2_xnor2_1 _14330_ (.Y(_06469_),
    .A(_06465_),
    .B(_06468_));
 sg13g2_xnor2_1 _14331_ (.Y(_06470_),
    .A(_06460_),
    .B(_06469_));
 sg13g2_buf_1 _14332_ (.A(_06470_),
    .X(_06471_));
 sg13g2_nand2_1 _14333_ (.Y(_06472_),
    .A(net163),
    .B(net150));
 sg13g2_nand2_1 _14334_ (.Y(_06473_),
    .A(net134),
    .B(net192));
 sg13g2_nand2_1 _14335_ (.Y(_06474_),
    .A(net162),
    .B(net231));
 sg13g2_xnor2_1 _14336_ (.Y(_06476_),
    .A(_06473_),
    .B(_06474_));
 sg13g2_xnor2_1 _14337_ (.Y(_06477_),
    .A(_06472_),
    .B(_06476_));
 sg13g2_xor2_1 _14338_ (.B(_06477_),
    .A(_06291_),
    .X(_06478_));
 sg13g2_or2_1 _14339_ (.X(_06479_),
    .B(_06478_),
    .A(_06471_));
 sg13g2_nand2_1 _14340_ (.Y(_06480_),
    .A(_06471_),
    .B(_06478_));
 sg13g2_o21ai_1 _14341_ (.B1(_00281_),
    .Y(_06481_),
    .A1(_06081_),
    .A2(_06301_));
 sg13g2_and3_1 _14342_ (.X(_06482_),
    .A(_06297_),
    .B(_06075_),
    .C(_06481_));
 sg13g2_buf_1 _14343_ (.A(_06482_),
    .X(_06483_));
 sg13g2_a21o_1 _14344_ (.A2(_06480_),
    .A1(_06479_),
    .B1(_06483_),
    .X(_06484_));
 sg13g2_buf_1 _14345_ (.A(_06484_),
    .X(_06485_));
 sg13g2_nor2b_1 _14346_ (.A(_06478_),
    .B_N(_06471_),
    .Y(_06487_));
 sg13g2_nor2b_1 _14347_ (.A(_06471_),
    .B_N(_06478_),
    .Y(_06488_));
 sg13g2_o21ai_1 _14348_ (.B1(_06483_),
    .Y(_06489_),
    .A1(_06487_),
    .A2(_06488_));
 sg13g2_buf_1 _14349_ (.A(_06489_),
    .X(_06490_));
 sg13g2_and2_1 _14350_ (.A(_06485_),
    .B(_06490_),
    .X(_06491_));
 sg13g2_and4_1 _14351_ (.A(_06428_),
    .B(_06452_),
    .C(_06455_),
    .D(_06491_),
    .X(_06492_));
 sg13g2_a221oi_1 _14352_ (.B2(_06490_),
    .C1(_06451_),
    .B1(_06485_),
    .A1(_06428_),
    .Y(_06493_),
    .A2(_06455_));
 sg13g2_nand3_1 _14353_ (.B(_06485_),
    .C(_06490_),
    .A(_06451_),
    .Y(_06494_));
 sg13g2_a21oi_1 _14354_ (.A1(_06428_),
    .A2(_06455_),
    .Y(_06495_),
    .B1(_06494_));
 sg13g2_a21oi_1 _14355_ (.A1(_06485_),
    .A2(_06490_),
    .Y(_06496_),
    .B1(_06452_));
 sg13g2_and3_1 _14356_ (.X(_06498_),
    .A(_06428_),
    .B(_06455_),
    .C(_06496_));
 sg13g2_nor4_1 _14357_ (.A(_06492_),
    .B(_06493_),
    .C(_06495_),
    .D(_06498_),
    .Y(_06499_));
 sg13g2_xnor2_1 _14358_ (.Y(_06500_),
    .A(_06426_),
    .B(_06499_));
 sg13g2_xor2_1 _14359_ (.B(_06500_),
    .A(_06423_),
    .X(_06501_));
 sg13g2_xnor2_1 _14360_ (.Y(_06502_),
    .A(_06421_),
    .B(_06501_));
 sg13g2_nand2_1 _14361_ (.Y(_06503_),
    .A(_06340_),
    .B(_06339_));
 sg13g2_o21ai_1 _14362_ (.B1(_06341_),
    .Y(_06504_),
    .A1(_06340_),
    .A2(_06339_));
 sg13g2_nand2_1 _14363_ (.Y(_06505_),
    .A(_06503_),
    .B(_06504_));
 sg13g2_and2_1 _14364_ (.A(_06366_),
    .B(_06369_),
    .X(_06506_));
 sg13g2_or2_1 _14365_ (.X(_06507_),
    .B(_06369_),
    .A(_06366_));
 sg13g2_o21ai_1 _14366_ (.B1(_06507_),
    .Y(_06509_),
    .A1(_06362_),
    .A2(_06506_));
 sg13g2_buf_1 _14367_ (.A(_06509_),
    .X(_06510_));
 sg13g2_xor2_1 _14368_ (.B(_06510_),
    .A(_06505_),
    .X(_06511_));
 sg13g2_xnor2_1 _14369_ (.Y(_06512_),
    .A(_06502_),
    .B(_06511_));
 sg13g2_a21oi_1 _14370_ (.A1(_06279_),
    .A2(_06280_),
    .Y(_06513_),
    .B1(_06371_));
 sg13g2_nand3_1 _14371_ (.B(_06280_),
    .C(_06371_),
    .A(_06279_),
    .Y(_06514_));
 sg13g2_o21ai_1 _14372_ (.B1(_06514_),
    .Y(_06515_),
    .A1(_06285_),
    .A2(_06513_));
 sg13g2_buf_2 _14373_ (.A(_06515_),
    .X(_06516_));
 sg13g2_xnor2_1 _14374_ (.Y(_06517_),
    .A(_06512_),
    .B(_06516_));
 sg13g2_xnor2_1 _14375_ (.Y(_06518_),
    .A(_04138_),
    .B(_06517_));
 sg13g2_a21o_1 _14376_ (.A2(_06416_),
    .A1(_06415_),
    .B1(_06518_),
    .X(_06520_));
 sg13g2_buf_1 _14377_ (.A(_06520_),
    .X(_06521_));
 sg13g2_nand2b_1 _14378_ (.Y(_06522_),
    .B(_04139_),
    .A_N(_06517_));
 sg13g2_nand2_1 _14379_ (.Y(_06523_),
    .A(_06512_),
    .B(_06516_));
 sg13g2_nand2_1 _14380_ (.Y(_06524_),
    .A(_06421_),
    .B(_06500_));
 sg13g2_o21ai_1 _14381_ (.B1(_06423_),
    .Y(_06525_),
    .A1(_06421_),
    .A2(_06500_));
 sg13g2_nand2_1 _14382_ (.Y(_06526_),
    .A(_06524_),
    .B(_06525_));
 sg13g2_nor3_2 _14383_ (.A(_02041_),
    .B(net170),
    .C(_02131_),
    .Y(_06527_));
 sg13g2_a21o_1 _14384_ (.A2(_06449_),
    .A1(_06443_),
    .B1(_06446_),
    .X(_06528_));
 sg13g2_o21ai_1 _14385_ (.B1(_06528_),
    .Y(_06529_),
    .A1(_06443_),
    .A2(_06449_));
 sg13g2_xor2_1 _14386_ (.B(_06478_),
    .A(_06483_),
    .X(_06531_));
 sg13g2_inv_1 _14387_ (.Y(_06532_),
    .A(_06531_));
 sg13g2_nand3_1 _14388_ (.B(_06455_),
    .C(_06471_),
    .A(_06428_),
    .Y(_06533_));
 sg13g2_a21oi_1 _14389_ (.A1(_06428_),
    .A2(_06455_),
    .Y(_06534_),
    .B1(_06471_));
 sg13g2_a21oi_1 _14390_ (.A1(_06532_),
    .A2(_06533_),
    .Y(_06535_),
    .B1(_06534_));
 sg13g2_nand2_1 _14391_ (.Y(_06536_),
    .A(net249),
    .B(net144));
 sg13g2_nand2_1 _14392_ (.Y(_06537_),
    .A(net201),
    .B(net152));
 sg13g2_nand2_1 _14393_ (.Y(_06538_),
    .A(net158),
    .B(net151));
 sg13g2_xnor2_1 _14394_ (.Y(_06539_),
    .A(_06537_),
    .B(_06538_));
 sg13g2_xnor2_1 _14395_ (.Y(_06540_),
    .A(_06536_),
    .B(_06539_));
 sg13g2_and2_1 _14396_ (.A(_06430_),
    .B(_06432_),
    .X(_06542_));
 sg13g2_or2_1 _14397_ (.X(_06543_),
    .B(_06432_),
    .A(_06430_));
 sg13g2_o21ai_1 _14398_ (.B1(_06543_),
    .Y(_06544_),
    .A1(_06429_),
    .A2(_06542_));
 sg13g2_nand2_1 _14399_ (.Y(_06545_),
    .A(net159),
    .B(net230));
 sg13g2_nand2_1 _14400_ (.Y(_06546_),
    .A(net248),
    .B(net114));
 sg13g2_xnor2_1 _14401_ (.Y(_06547_),
    .A(_06545_),
    .B(_06546_));
 sg13g2_xnor2_1 _14402_ (.Y(_06548_),
    .A(_06544_),
    .B(_06547_));
 sg13g2_xnor2_1 _14403_ (.Y(_06549_),
    .A(_06540_),
    .B(_06548_));
 sg13g2_or2_1 _14404_ (.X(_06550_),
    .B(_06468_),
    .A(_06465_));
 sg13g2_nand2_1 _14405_ (.Y(_06551_),
    .A(_06465_),
    .B(_06468_));
 sg13g2_nand2_1 _14406_ (.Y(_06553_),
    .A(_06460_),
    .B(_06551_));
 sg13g2_nand2_1 _14407_ (.Y(_06554_),
    .A(_06434_),
    .B(_06440_));
 sg13g2_nand2_1 _14408_ (.Y(_06555_),
    .A(_06437_),
    .B(_06554_));
 sg13g2_o21ai_1 _14409_ (.B1(_06555_),
    .Y(_06556_),
    .A1(_06434_),
    .A2(_06440_));
 sg13g2_a21oi_1 _14410_ (.A1(_06550_),
    .A2(_06553_),
    .Y(_06557_),
    .B1(_06556_));
 sg13g2_and3_1 _14411_ (.X(_06558_),
    .A(_06550_),
    .B(_06553_),
    .C(_06556_));
 sg13g2_nor2_1 _14412_ (.A(_06557_),
    .B(_06558_),
    .Y(_06559_));
 sg13g2_xnor2_1 _14413_ (.Y(_06560_),
    .A(_06549_),
    .B(_06559_));
 sg13g2_buf_1 _14414_ (.A(_06560_),
    .X(_06561_));
 sg13g2_nand2_1 _14415_ (.Y(_06562_),
    .A(net212),
    .B(net180));
 sg13g2_nand2_1 _14416_ (.Y(_06564_),
    .A(net133),
    .B(net231));
 sg13g2_nand2_1 _14417_ (.Y(_06565_),
    .A(net217),
    .B(net177));
 sg13g2_xnor2_1 _14418_ (.Y(_06566_),
    .A(_06564_),
    .B(_06565_));
 sg13g2_xnor2_1 _14419_ (.Y(_06567_),
    .A(_06562_),
    .B(_06566_));
 sg13g2_and2_1 _14420_ (.A(_06472_),
    .B(_06473_),
    .X(_06568_));
 sg13g2_or2_1 _14421_ (.X(_06569_),
    .B(_06473_),
    .A(_06472_));
 sg13g2_o21ai_1 _14422_ (.B1(_06569_),
    .Y(_06570_),
    .A1(_06474_),
    .A2(_06568_));
 sg13g2_buf_1 _14423_ (.A(_06570_),
    .X(_06571_));
 sg13g2_and2_1 _14424_ (.A(_06457_),
    .B(_06458_),
    .X(_06572_));
 sg13g2_or2_1 _14425_ (.X(_06573_),
    .B(_06458_),
    .A(_06457_));
 sg13g2_o21ai_1 _14426_ (.B1(_06573_),
    .Y(_06575_),
    .A1(_06456_),
    .A2(_06572_));
 sg13g2_buf_1 _14427_ (.A(_06575_),
    .X(_06576_));
 sg13g2_xnor2_1 _14428_ (.Y(_06577_),
    .A(_06571_),
    .B(_06576_));
 sg13g2_xnor2_1 _14429_ (.Y(_06578_),
    .A(_06567_),
    .B(_06577_));
 sg13g2_nand2_1 _14430_ (.Y(_06579_),
    .A(net162),
    .B(net192));
 sg13g2_nand2_1 _14431_ (.Y(_06580_),
    .A(net150),
    .B(_01362_));
 sg13g2_xor2_1 _14432_ (.B(_06580_),
    .A(_06579_),
    .X(_06581_));
 sg13g2_and2_1 _14433_ (.A(_06578_),
    .B(_06581_),
    .X(_06582_));
 sg13g2_nand2_1 _14434_ (.Y(_06583_),
    .A(_06561_),
    .B(_06582_));
 sg13g2_xor2_1 _14435_ (.B(_06559_),
    .A(_06549_),
    .X(_06584_));
 sg13g2_nor2b_1 _14436_ (.A(_06578_),
    .B_N(_06581_),
    .Y(_06586_));
 sg13g2_nand2_1 _14437_ (.Y(_06587_),
    .A(_06584_),
    .B(_06586_));
 sg13g2_nand2_1 _14438_ (.Y(_06588_),
    .A(_06483_),
    .B(_06477_));
 sg13g2_o21ai_1 _14439_ (.B1(net97),
    .Y(_06589_),
    .A1(_06483_),
    .A2(_06477_));
 sg13g2_and2_1 _14440_ (.A(_06588_),
    .B(_06589_),
    .X(_06590_));
 sg13g2_buf_1 _14441_ (.A(_06590_),
    .X(_06591_));
 sg13g2_a21o_1 _14442_ (.A2(_06587_),
    .A1(_06583_),
    .B1(_06591_),
    .X(_06592_));
 sg13g2_inv_1 _14443_ (.Y(_06593_),
    .A(_06578_));
 sg13g2_buf_1 _14444_ (.A(_06581_),
    .X(_06594_));
 sg13g2_nor2_1 _14445_ (.A(_06593_),
    .B(net87),
    .Y(_06595_));
 sg13g2_nand2_1 _14446_ (.Y(_06597_),
    .A(_06584_),
    .B(_06595_));
 sg13g2_nor2_1 _14447_ (.A(_06578_),
    .B(net87),
    .Y(_06598_));
 sg13g2_nand2_1 _14448_ (.Y(_06599_),
    .A(_06561_),
    .B(_06598_));
 sg13g2_a21o_1 _14449_ (.A2(_06599_),
    .A1(_06597_),
    .B1(_06591_),
    .X(_06600_));
 sg13g2_and2_1 _14450_ (.A(_06584_),
    .B(_06582_),
    .X(_06601_));
 sg13g2_and2_1 _14451_ (.A(_06561_),
    .B(_06586_),
    .X(_06602_));
 sg13g2_o21ai_1 _14452_ (.B1(_06591_),
    .Y(_06603_),
    .A1(_06601_),
    .A2(_06602_));
 sg13g2_and2_1 _14453_ (.A(_06561_),
    .B(_06595_),
    .X(_06604_));
 sg13g2_and2_1 _14454_ (.A(_06584_),
    .B(_06598_),
    .X(_06605_));
 sg13g2_o21ai_1 _14455_ (.B1(_06591_),
    .Y(_06606_),
    .A1(_06604_),
    .A2(_06605_));
 sg13g2_nand4_1 _14456_ (.B(_06600_),
    .C(_06603_),
    .A(_06592_),
    .Y(_06608_),
    .D(_06606_));
 sg13g2_xor2_1 _14457_ (.B(_06608_),
    .A(_06535_),
    .X(_06609_));
 sg13g2_nand2_1 _14458_ (.Y(_06610_),
    .A(_06428_),
    .B(_06455_));
 sg13g2_nor2_1 _14459_ (.A(_06451_),
    .B(_06491_),
    .Y(_06611_));
 sg13g2_nor2_1 _14460_ (.A(_06495_),
    .B(_06498_),
    .Y(_06612_));
 sg13g2_a221oi_1 _14461_ (.B2(_06426_),
    .C1(_06492_),
    .B1(_06612_),
    .A1(_06610_),
    .Y(_06613_),
    .A2(_06611_));
 sg13g2_xnor2_1 _14462_ (.Y(_06614_),
    .A(_06609_),
    .B(_06613_));
 sg13g2_xnor2_1 _14463_ (.Y(_06615_),
    .A(_06529_),
    .B(_06614_));
 sg13g2_xor2_1 _14464_ (.B(_06615_),
    .A(_06527_),
    .X(_06616_));
 sg13g2_xnor2_1 _14465_ (.Y(_06617_),
    .A(_06526_),
    .B(_06616_));
 sg13g2_buf_1 _14466_ (.A(_06617_),
    .X(_06619_));
 sg13g2_nand2_1 _14467_ (.Y(_06620_),
    .A(_06510_),
    .B(_06502_));
 sg13g2_nor2_1 _14468_ (.A(_06510_),
    .B(_06502_),
    .Y(_06621_));
 sg13g2_a21oi_2 _14469_ (.B1(_06621_),
    .Y(_06622_),
    .A2(_06620_),
    .A1(_06505_));
 sg13g2_xnor2_1 _14470_ (.Y(_06623_),
    .A(_06619_),
    .B(_06622_));
 sg13g2_xnor2_1 _14471_ (.Y(_06624_),
    .A(_06523_),
    .B(_06623_));
 sg13g2_or2_1 _14472_ (.X(_06625_),
    .B(_06624_),
    .A(_04058_));
 sg13g2_nand2_1 _14473_ (.Y(_06626_),
    .A(_04058_),
    .B(_06624_));
 sg13g2_a22oi_1 _14474_ (.Y(_06627_),
    .B1(_06625_),
    .B2(_06626_),
    .A2(_06522_),
    .A1(_06521_));
 sg13g2_nor2_1 _14475_ (.A(_00020_),
    .B(_06624_),
    .Y(_06628_));
 sg13g2_inv_1 _14476_ (.Y(_06630_),
    .A(_06622_));
 sg13g2_a21oi_1 _14477_ (.A1(_06512_),
    .A2(_06516_),
    .Y(_06631_),
    .B1(_06619_));
 sg13g2_nand3_1 _14478_ (.B(_06516_),
    .C(_06619_),
    .A(_06512_),
    .Y(_06632_));
 sg13g2_o21ai_1 _14479_ (.B1(_06632_),
    .Y(_06633_),
    .A1(_06630_),
    .A2(_06631_));
 sg13g2_nor2_1 _14480_ (.A(_06527_),
    .B(_06615_),
    .Y(_06634_));
 sg13g2_nand2_1 _14481_ (.Y(_06635_),
    .A(_06527_),
    .B(_06615_));
 sg13g2_o21ai_1 _14482_ (.B1(_06635_),
    .Y(_06636_),
    .A1(_06526_),
    .A2(_06634_));
 sg13g2_nand2b_1 _14483_ (.Y(_06637_),
    .B(_06609_),
    .A_N(_06529_));
 sg13g2_nor2b_1 _14484_ (.A(_06609_),
    .B_N(_06529_),
    .Y(_06638_));
 sg13g2_a21oi_1 _14485_ (.A1(_06613_),
    .A2(_06637_),
    .Y(_06639_),
    .B1(_06638_));
 sg13g2_inv_1 _14486_ (.Y(_06641_),
    .A(_02131_));
 sg13g2_nand2_1 _14487_ (.Y(_06642_),
    .A(_03207_),
    .B(_06641_));
 sg13g2_xnor2_1 _14488_ (.Y(_06643_),
    .A(_06591_),
    .B(net87));
 sg13g2_xnor2_1 _14489_ (.Y(_06644_),
    .A(_06593_),
    .B(_06643_));
 sg13g2_a21o_1 _14490_ (.A2(_06644_),
    .A1(_06561_),
    .B1(_06535_),
    .X(_06645_));
 sg13g2_o21ai_1 _14491_ (.B1(_06645_),
    .Y(_06646_),
    .A1(_06561_),
    .A2(_06644_));
 sg13g2_buf_1 _14492_ (.A(_06300_),
    .X(_06647_));
 sg13g2_nand3_1 _14493_ (.B(_06647_),
    .C(_06481_),
    .A(net97),
    .Y(_06648_));
 sg13g2_nor3_1 _14494_ (.A(net97),
    .B(_06300_),
    .C(_06303_),
    .Y(_06649_));
 sg13g2_a21oi_1 _14495_ (.A1(net97),
    .A2(_06477_),
    .Y(_06650_),
    .B1(_06649_));
 sg13g2_nand3_1 _14496_ (.B(_06648_),
    .C(_06650_),
    .A(_06588_),
    .Y(_06652_));
 sg13g2_nand2_1 _14497_ (.Y(_06653_),
    .A(net97),
    .B(_06303_));
 sg13g2_inv_1 _14498_ (.Y(_06654_),
    .A(_06653_));
 sg13g2_nand3_1 _14499_ (.B(_06594_),
    .C(_06654_),
    .A(_06647_),
    .Y(_06655_));
 sg13g2_o21ai_1 _14500_ (.B1(_06655_),
    .Y(_06656_),
    .A1(net87),
    .A2(_06652_));
 sg13g2_a21oi_2 _14501_ (.B1(_06656_),
    .Y(_06657_),
    .A2(_06643_),
    .A1(_06593_));
 sg13g2_nand2_1 _14502_ (.Y(_06658_),
    .A(_06594_),
    .B(_06653_));
 sg13g2_nor2_1 _14503_ (.A(net97),
    .B(_06303_),
    .Y(_06659_));
 sg13g2_nor2_1 _14504_ (.A(net87),
    .B(_06659_),
    .Y(_06660_));
 sg13g2_a21oi_1 _14505_ (.A1(net28),
    .A2(_06658_),
    .Y(_06661_),
    .B1(_06660_));
 sg13g2_xnor2_1 _14506_ (.Y(_06663_),
    .A(net163),
    .B(_00246_));
 sg13g2_nand2_2 _14507_ (.Y(_06664_),
    .A(net122),
    .B(_06663_));
 sg13g2_buf_1 _14508_ (.A(net212),
    .X(_06665_));
 sg13g2_nand2_1 _14509_ (.Y(_06666_),
    .A(net132),
    .B(net149));
 sg13g2_nand2_1 _14510_ (.Y(_06667_),
    .A(net133),
    .B(net192));
 sg13g2_nand2_1 _14511_ (.Y(_06668_),
    .A(net217),
    .B(net231));
 sg13g2_xnor2_1 _14512_ (.Y(_06669_),
    .A(_06667_),
    .B(_06668_));
 sg13g2_xnor2_1 _14513_ (.Y(_06670_),
    .A(_06666_),
    .B(_06669_));
 sg13g2_nor2_1 _14514_ (.A(net163),
    .B(net134),
    .Y(_06671_));
 sg13g2_o21ai_1 _14515_ (.B1(_01267_),
    .Y(_06672_),
    .A1(_06579_),
    .A2(_06671_));
 sg13g2_nand2_1 _14516_ (.Y(_06674_),
    .A(net150),
    .B(_06672_));
 sg13g2_and2_1 _14517_ (.A(_06564_),
    .B(_06565_),
    .X(_06675_));
 sg13g2_or2_1 _14518_ (.X(_06676_),
    .B(_06565_),
    .A(_06564_));
 sg13g2_o21ai_1 _14519_ (.B1(_06676_),
    .Y(_06677_),
    .A1(_06562_),
    .A2(_06675_));
 sg13g2_xnor2_1 _14520_ (.Y(_06678_),
    .A(_06674_),
    .B(_06677_));
 sg13g2_xor2_1 _14521_ (.B(_06678_),
    .A(_06670_),
    .X(_06679_));
 sg13g2_xnor2_1 _14522_ (.Y(_06680_),
    .A(_06664_),
    .B(_06679_));
 sg13g2_xnor2_1 _14523_ (.Y(_06681_),
    .A(_06661_),
    .B(_06680_));
 sg13g2_buf_1 _14524_ (.A(_06681_),
    .X(_06682_));
 sg13g2_nand2_1 _14525_ (.Y(_06683_),
    .A(net199),
    .B(net151));
 sg13g2_nand2_1 _14526_ (.Y(_06685_),
    .A(net157),
    .B(net153));
 sg13g2_nand2_1 _14527_ (.Y(_06686_),
    .A(net158),
    .B(net152));
 sg13g2_xnor2_1 _14528_ (.Y(_06687_),
    .A(_06685_),
    .B(_06686_));
 sg13g2_xnor2_1 _14529_ (.Y(_06688_),
    .A(_06683_),
    .B(_06687_));
 sg13g2_and2_1 _14530_ (.A(_06537_),
    .B(_06538_),
    .X(_06689_));
 sg13g2_or2_1 _14531_ (.X(_06690_),
    .B(_06538_),
    .A(_06537_));
 sg13g2_o21ai_1 _14532_ (.B1(_06690_),
    .Y(_06691_),
    .A1(_06536_),
    .A2(_06689_));
 sg13g2_nand2_1 _14533_ (.Y(_06692_),
    .A(net159),
    .B(_02040_));
 sg13g2_nand2_1 _14534_ (.Y(_06693_),
    .A(net248),
    .B(net144));
 sg13g2_xnor2_1 _14535_ (.Y(_06694_),
    .A(_06692_),
    .B(_06693_));
 sg13g2_xor2_1 _14536_ (.B(_06694_),
    .A(_06691_),
    .X(_06696_));
 sg13g2_xnor2_1 _14537_ (.Y(_06697_),
    .A(_06688_),
    .B(_06696_));
 sg13g2_inv_1 _14538_ (.Y(_06698_),
    .A(_06697_));
 sg13g2_nand2_1 _14539_ (.Y(_06699_),
    .A(_06540_),
    .B(_06547_));
 sg13g2_nand2_1 _14540_ (.Y(_06700_),
    .A(_06544_),
    .B(_06699_));
 sg13g2_o21ai_1 _14541_ (.B1(_06700_),
    .Y(_06701_),
    .A1(_06540_),
    .A2(_06547_));
 sg13g2_nand2_1 _14542_ (.Y(_06702_),
    .A(_06571_),
    .B(_06576_));
 sg13g2_nor2_1 _14543_ (.A(_06571_),
    .B(_06576_),
    .Y(_06703_));
 sg13g2_a21oi_1 _14544_ (.A1(_06567_),
    .A2(_06702_),
    .Y(_06704_),
    .B1(_06703_));
 sg13g2_nor2_1 _14545_ (.A(_06701_),
    .B(_06704_),
    .Y(_06705_));
 sg13g2_buf_1 _14546_ (.A(_06705_),
    .X(_06707_));
 sg13g2_and2_1 _14547_ (.A(_06701_),
    .B(_06704_),
    .X(_06708_));
 sg13g2_buf_1 _14548_ (.A(_06708_),
    .X(_06709_));
 sg13g2_nor2_1 _14549_ (.A(_06707_),
    .B(_06709_),
    .Y(_06710_));
 sg13g2_xnor2_1 _14550_ (.Y(_06711_),
    .A(_06698_),
    .B(_06710_));
 sg13g2_xnor2_1 _14551_ (.Y(_06712_),
    .A(_06682_),
    .B(_06711_));
 sg13g2_xnor2_1 _14552_ (.Y(_06713_),
    .A(_06657_),
    .B(_06712_));
 sg13g2_nor2_1 _14553_ (.A(_06549_),
    .B(_06558_),
    .Y(_06714_));
 sg13g2_nor2_1 _14554_ (.A(_06557_),
    .B(_06714_),
    .Y(_06715_));
 sg13g2_xnor2_1 _14555_ (.Y(_06716_),
    .A(_06713_),
    .B(_06715_));
 sg13g2_xnor2_1 _14556_ (.Y(_06718_),
    .A(_06646_),
    .B(_06716_));
 sg13g2_xor2_1 _14557_ (.B(_06718_),
    .A(_06642_),
    .X(_06719_));
 sg13g2_xnor2_1 _14558_ (.Y(_06720_),
    .A(_06639_),
    .B(_06719_));
 sg13g2_xnor2_1 _14559_ (.Y(_06721_),
    .A(_06636_),
    .B(_06720_));
 sg13g2_xnor2_1 _14560_ (.Y(_06722_),
    .A(_06633_),
    .B(_06721_));
 sg13g2_xnor2_1 _14561_ (.Y(_06723_),
    .A(_04076_),
    .B(_06722_));
 sg13g2_o21ai_1 _14562_ (.B1(_06723_),
    .Y(_06724_),
    .A1(_06627_),
    .A2(_06628_));
 sg13g2_or3_1 _14563_ (.A(_06627_),
    .B(_06628_),
    .C(_06723_),
    .X(_06725_));
 sg13g2_nand2_1 _14564_ (.Y(_06726_),
    .A(_06724_),
    .B(_06725_));
 sg13g2_a21oi_1 _14565_ (.A1(net98),
    .A2(_06726_),
    .Y(_06727_),
    .B1(_05064_));
 sg13g2_mux2_1 _14566_ (.A0(_06727_),
    .A1(_06665_),
    .S(net15),
    .X(_00225_));
 sg13g2_or2_1 _14567_ (.X(_06729_),
    .B(_06722_),
    .A(_00022_));
 sg13g2_inv_1 _14568_ (.Y(_06730_),
    .A(_06636_));
 sg13g2_nor2_1 _14569_ (.A(_06730_),
    .B(_06720_),
    .Y(_06731_));
 sg13g2_nand2_1 _14570_ (.Y(_06732_),
    .A(_06619_),
    .B(_06622_));
 sg13g2_nor2_1 _14571_ (.A(_06619_),
    .B(_06622_),
    .Y(_06733_));
 sg13g2_a21oi_1 _14572_ (.A1(_06523_),
    .A2(_06732_),
    .Y(_06734_),
    .B1(_06733_));
 sg13g2_nand2_1 _14573_ (.Y(_06735_),
    .A(_06730_),
    .B(_06720_));
 sg13g2_o21ai_1 _14574_ (.B1(_06735_),
    .Y(_06736_),
    .A1(_06731_),
    .A2(_06734_));
 sg13g2_nand2_1 _14575_ (.Y(_06737_),
    .A(_06642_),
    .B(_06718_));
 sg13g2_nor2_1 _14576_ (.A(_06642_),
    .B(_06718_),
    .Y(_06739_));
 sg13g2_a21oi_1 _14577_ (.A1(_06639_),
    .A2(_06737_),
    .Y(_06740_),
    .B1(_06739_));
 sg13g2_nand2b_1 _14578_ (.Y(_06741_),
    .B(_06713_),
    .A_N(_06715_));
 sg13g2_nor2b_1 _14579_ (.A(_06713_),
    .B_N(_06715_),
    .Y(_06742_));
 sg13g2_a21o_1 _14580_ (.A2(_06741_),
    .A1(_06646_),
    .B1(_06742_),
    .X(_06743_));
 sg13g2_buf_1 _14581_ (.A(_06743_),
    .X(_06744_));
 sg13g2_and2_1 _14582_ (.A(net122),
    .B(_06663_),
    .X(_06745_));
 sg13g2_buf_1 _14583_ (.A(_06745_),
    .X(_06746_));
 sg13g2_a21oi_1 _14584_ (.A1(net28),
    .A2(_06746_),
    .Y(_06747_),
    .B1(_06679_));
 sg13g2_nand2_1 _14585_ (.Y(_06748_),
    .A(_06746_),
    .B(_06679_));
 sg13g2_o21ai_1 _14586_ (.B1(_06748_),
    .Y(_06750_),
    .A1(net87),
    .A2(_06747_));
 sg13g2_a21oi_1 _14587_ (.A1(net97),
    .A2(_06746_),
    .Y(_06751_),
    .B1(_06679_));
 sg13g2_o21ai_1 _14588_ (.B1(_06748_),
    .Y(_06752_),
    .A1(net87),
    .A2(_06751_));
 sg13g2_a21oi_1 _14589_ (.A1(_06659_),
    .A2(_06664_),
    .Y(_06753_),
    .B1(_06752_));
 sg13g2_and4_1 _14590_ (.A(_06292_),
    .B(net28),
    .C(_06664_),
    .D(_06679_),
    .X(_06754_));
 sg13g2_nor3_1 _14591_ (.A(net28),
    .B(net87),
    .C(_06664_),
    .Y(_06755_));
 sg13g2_o21ai_1 _14592_ (.B1(_06303_),
    .Y(_06756_),
    .A1(_06754_),
    .A2(_06755_));
 sg13g2_o21ai_1 _14593_ (.B1(_06756_),
    .Y(_06757_),
    .A1(net28),
    .A2(_06753_));
 sg13g2_a21o_1 _14594_ (.A2(_06750_),
    .A1(_06653_),
    .B1(_06757_),
    .X(_06758_));
 sg13g2_buf_1 _14595_ (.A(_06758_),
    .X(_06759_));
 sg13g2_nand2_1 _14596_ (.Y(_06761_),
    .A(net199),
    .B(net152));
 sg13g2_nand2_1 _14597_ (.Y(_06762_),
    .A(net157),
    .B(net149));
 sg13g2_nand2_1 _14598_ (.Y(_06763_),
    .A(net158),
    .B(net153));
 sg13g2_xnor2_1 _14599_ (.Y(_06764_),
    .A(_06762_),
    .B(_06763_));
 sg13g2_xnor2_1 _14600_ (.Y(_06765_),
    .A(_06761_),
    .B(_06764_));
 sg13g2_and2_1 _14601_ (.A(_06685_),
    .B(_06686_),
    .X(_06766_));
 sg13g2_or2_1 _14602_ (.X(_06767_),
    .B(_06686_),
    .A(_06685_));
 sg13g2_o21ai_1 _14603_ (.B1(_06767_),
    .Y(_06768_),
    .A1(_06683_),
    .A2(_06766_));
 sg13g2_nand2_1 _14604_ (.Y(_06769_),
    .A(net159),
    .B(_01983_));
 sg13g2_nand2_1 _14605_ (.Y(_06770_),
    .A(net248),
    .B(_02017_));
 sg13g2_xnor2_1 _14606_ (.Y(_06772_),
    .A(_06769_),
    .B(_06770_));
 sg13g2_xnor2_1 _14607_ (.Y(_06773_),
    .A(_06768_),
    .B(_06772_));
 sg13g2_xnor2_1 _14608_ (.Y(_06774_),
    .A(_06765_),
    .B(_06773_));
 sg13g2_inv_1 _14609_ (.Y(_06775_),
    .A(_06677_));
 sg13g2_nand2_1 _14610_ (.Y(_06776_),
    .A(_06674_),
    .B(_06775_));
 sg13g2_o21ai_1 _14611_ (.B1(_06670_),
    .Y(_06777_),
    .A1(_06674_),
    .A2(_06775_));
 sg13g2_nand2_1 _14612_ (.Y(_06778_),
    .A(_06776_),
    .B(_06777_));
 sg13g2_nand2_1 _14613_ (.Y(_06779_),
    .A(_06688_),
    .B(_06694_));
 sg13g2_nor2_1 _14614_ (.A(_06688_),
    .B(_06694_),
    .Y(_06780_));
 sg13g2_a21oi_1 _14615_ (.A1(_06691_),
    .A2(_06779_),
    .Y(_06781_),
    .B1(_06780_));
 sg13g2_xnor2_1 _14616_ (.Y(_06783_),
    .A(_06778_),
    .B(_06781_));
 sg13g2_xnor2_1 _14617_ (.Y(_06784_),
    .A(_06774_),
    .B(_06783_));
 sg13g2_nand3_1 _14618_ (.B(_06654_),
    .C(_06746_),
    .A(net28),
    .Y(_06785_));
 sg13g2_buf_1 _14619_ (.A(_06785_),
    .X(_06786_));
 sg13g2_nand3b_1 _14620_ (.B(_06659_),
    .C(_06664_),
    .Y(_06787_),
    .A_N(net28));
 sg13g2_nand2_1 _14621_ (.Y(_06788_),
    .A(_06786_),
    .B(_06787_));
 sg13g2_nand2_1 _14622_ (.Y(_06789_),
    .A(net133),
    .B(net122));
 sg13g2_nand2_1 _14623_ (.Y(_06790_),
    .A(net217),
    .B(net192));
 sg13g2_nand2_1 _14624_ (.Y(_06791_),
    .A(net132),
    .B(net231));
 sg13g2_xnor2_1 _14625_ (.Y(_06792_),
    .A(_06790_),
    .B(_06791_));
 sg13g2_xnor2_1 _14626_ (.Y(_06794_),
    .A(_06789_),
    .B(_06792_));
 sg13g2_and2_1 _14627_ (.A(_06667_),
    .B(_06668_),
    .X(_06795_));
 sg13g2_or2_1 _14628_ (.X(_06796_),
    .B(_06668_),
    .A(_06667_));
 sg13g2_o21ai_1 _14629_ (.B1(_06796_),
    .Y(_06797_),
    .A1(_06666_),
    .A2(_06795_));
 sg13g2_buf_1 _14630_ (.A(_06797_),
    .X(_06798_));
 sg13g2_xnor2_1 _14631_ (.Y(_06799_),
    .A(_06794_),
    .B(_06798_));
 sg13g2_o21ai_1 _14632_ (.B1(net162),
    .Y(_06800_),
    .A1(net163),
    .A2(net134));
 sg13g2_a21oi_1 _14633_ (.A1(_01267_),
    .A2(_06800_),
    .Y(_06801_),
    .B1(net191));
 sg13g2_buf_1 _14634_ (.A(_06801_),
    .X(_06802_));
 sg13g2_xnor2_1 _14635_ (.Y(_06803_),
    .A(_06799_),
    .B(net86));
 sg13g2_xnor2_1 _14636_ (.Y(_06805_),
    .A(_06788_),
    .B(_06803_));
 sg13g2_xor2_1 _14637_ (.B(_06805_),
    .A(_06784_),
    .X(_06806_));
 sg13g2_xnor2_1 _14638_ (.Y(_06807_),
    .A(_06759_),
    .B(_06806_));
 sg13g2_buf_1 _14639_ (.A(_06807_),
    .X(_06808_));
 sg13g2_nor2_1 _14640_ (.A(_06682_),
    .B(_06697_),
    .Y(_06809_));
 sg13g2_and2_1 _14641_ (.A(_06682_),
    .B(_06697_),
    .X(_06810_));
 sg13g2_buf_1 _14642_ (.A(_06810_),
    .X(_06811_));
 sg13g2_a22oi_1 _14643_ (.Y(_06812_),
    .B1(_06811_),
    .B2(_06707_),
    .A2(_06809_),
    .A1(_06709_));
 sg13g2_nor2_1 _14644_ (.A(_06697_),
    .B(_06707_),
    .Y(_06813_));
 sg13g2_nor2_1 _14645_ (.A(_06709_),
    .B(_06813_),
    .Y(_06814_));
 sg13g2_nor2_1 _14646_ (.A(_06682_),
    .B(_06814_),
    .Y(_06816_));
 sg13g2_a21oi_1 _14647_ (.A1(_06698_),
    .A2(_06709_),
    .Y(_06817_),
    .B1(_06816_));
 sg13g2_a22oi_1 _14648_ (.Y(_06818_),
    .B1(_06814_),
    .B2(_06682_),
    .A2(_06707_),
    .A1(_06697_));
 sg13g2_mux2_1 _14649_ (.A0(_06817_),
    .A1(_06818_),
    .S(_06657_),
    .X(_06819_));
 sg13g2_nand2_1 _14650_ (.Y(_06820_),
    .A(_06812_),
    .B(_06819_));
 sg13g2_xor2_1 _14651_ (.B(_06820_),
    .A(_06808_),
    .X(_06821_));
 sg13g2_nor3_1 _14652_ (.A(_01983_),
    .B(net114),
    .C(_02131_),
    .Y(_06822_));
 sg13g2_xor2_1 _14653_ (.B(_06822_),
    .A(_06821_),
    .X(_06823_));
 sg13g2_xnor2_1 _14654_ (.Y(_06824_),
    .A(_06744_),
    .B(_06823_));
 sg13g2_and2_1 _14655_ (.A(_06740_),
    .B(_06824_),
    .X(_06825_));
 sg13g2_or2_1 _14656_ (.X(_06827_),
    .B(_06824_),
    .A(_06740_));
 sg13g2_nor2b_1 _14657_ (.A(_06825_),
    .B_N(_06827_),
    .Y(_06828_));
 sg13g2_xnor2_1 _14658_ (.Y(_06829_),
    .A(_06736_),
    .B(_06828_));
 sg13g2_xnor2_1 _14659_ (.Y(_06830_),
    .A(_04083_),
    .B(_06829_));
 sg13g2_a21oi_1 _14660_ (.A1(_06724_),
    .A2(_06729_),
    .Y(_06831_),
    .B1(_06830_));
 sg13g2_and3_1 _14661_ (.X(_06832_),
    .A(_06724_),
    .B(_06729_),
    .C(_06830_));
 sg13g2_buf_1 _14662_ (.A(net139),
    .X(_06833_));
 sg13g2_o21ai_1 _14663_ (.B1(net112),
    .Y(_06834_),
    .A1(_06831_),
    .A2(_06832_));
 sg13g2_nor2b_1 _14664_ (.A(_05075_),
    .B_N(_06834_),
    .Y(_06835_));
 sg13g2_mux2_1 _14665_ (.A0(_06835_),
    .A1(net157),
    .S(_05012_),
    .X(_00226_));
 sg13g2_inv_1 _14666_ (.Y(_06837_),
    .A(_00023_));
 sg13g2_a21oi_1 _14667_ (.A1(_06837_),
    .A2(_06829_),
    .Y(_06838_),
    .B1(_06831_));
 sg13g2_a21o_1 _14668_ (.A2(_06827_),
    .A1(_06736_),
    .B1(_06825_),
    .X(_06839_));
 sg13g2_buf_1 _14669_ (.A(_06839_),
    .X(_06840_));
 sg13g2_inv_1 _14670_ (.Y(_06841_),
    .A(_06809_));
 sg13g2_or2_1 _14671_ (.X(_06842_),
    .B(_06811_),
    .A(_06808_));
 sg13g2_a22oi_1 _14672_ (.Y(_06843_),
    .B1(_06842_),
    .B2(_06657_),
    .A2(_06841_),
    .A1(_06808_));
 sg13g2_a21oi_1 _14673_ (.A1(_06657_),
    .A2(_06841_),
    .Y(_06844_),
    .B1(_06811_));
 sg13g2_nor2_1 _14674_ (.A(_06707_),
    .B(_06808_),
    .Y(_06845_));
 sg13g2_nor2_1 _14675_ (.A(_06844_),
    .B(_06845_),
    .Y(_06846_));
 sg13g2_a21oi_1 _14676_ (.A1(_06707_),
    .A2(_06808_),
    .Y(_06848_),
    .B1(_06846_));
 sg13g2_o21ai_1 _14677_ (.B1(_06848_),
    .Y(_06849_),
    .A1(_06709_),
    .A2(_06843_));
 sg13g2_nor2_1 _14678_ (.A(_06759_),
    .B(_06805_),
    .Y(_06850_));
 sg13g2_nand2_1 _14679_ (.Y(_06851_),
    .A(_06759_),
    .B(_06805_));
 sg13g2_o21ai_1 _14680_ (.B1(_06851_),
    .Y(_06852_),
    .A1(_06784_),
    .A2(_06850_));
 sg13g2_nor2_1 _14681_ (.A(_06778_),
    .B(_06781_),
    .Y(_06853_));
 sg13g2_nand2_1 _14682_ (.Y(_06854_),
    .A(_06778_),
    .B(_06781_));
 sg13g2_o21ai_1 _14683_ (.B1(_06854_),
    .Y(_06855_),
    .A1(_06774_),
    .A2(_06853_));
 sg13g2_nor4_2 _14684_ (.A(_06292_),
    .B(net28),
    .C(_06303_),
    .Y(_06856_),
    .D(_06746_));
 sg13g2_nor2_1 _14685_ (.A(_06786_),
    .B(net86),
    .Y(_06857_));
 sg13g2_a21oi_1 _14686_ (.A1(_06856_),
    .A2(net86),
    .Y(_06859_),
    .B1(_06857_));
 sg13g2_o21ai_1 _14687_ (.B1(_06859_),
    .Y(_06860_),
    .A1(_06788_),
    .A2(_06799_));
 sg13g2_nand2_1 _14688_ (.Y(_06861_),
    .A(net132),
    .B(net154));
 sg13g2_xnor2_1 _14689_ (.Y(_06862_),
    .A(net217),
    .B(net133));
 sg13g2_nor2_1 _14690_ (.A(_01497_),
    .B(_06862_),
    .Y(_06863_));
 sg13g2_xnor2_1 _14691_ (.Y(_06864_),
    .A(_06861_),
    .B(_06863_));
 sg13g2_and2_1 _14692_ (.A(_06789_),
    .B(_06790_),
    .X(_06865_));
 sg13g2_or2_1 _14693_ (.X(_06866_),
    .B(_06790_),
    .A(_06789_));
 sg13g2_o21ai_1 _14694_ (.B1(_06866_),
    .Y(_06867_),
    .A1(_06791_),
    .A2(_06865_));
 sg13g2_buf_1 _14695_ (.A(_06867_),
    .X(_06868_));
 sg13g2_xnor2_1 _14696_ (.Y(_06870_),
    .A(_06864_),
    .B(_06868_));
 sg13g2_a21o_1 _14697_ (.A2(_06763_),
    .A1(_06762_),
    .B1(_06761_),
    .X(_06871_));
 sg13g2_o21ai_1 _14698_ (.B1(_06871_),
    .Y(_06872_),
    .A1(_06762_),
    .A2(_06763_));
 sg13g2_nand2_1 _14699_ (.Y(_06873_),
    .A(net199),
    .B(net153));
 sg13g2_nand2_1 _14700_ (.Y(_06874_),
    .A(net157),
    .B(net231));
 sg13g2_nand2_1 _14701_ (.Y(_06875_),
    .A(net158),
    .B(net149));
 sg13g2_xor2_1 _14702_ (.B(_06875_),
    .A(_06874_),
    .X(_06876_));
 sg13g2_xnor2_1 _14703_ (.Y(_06877_),
    .A(_06873_),
    .B(_06876_));
 sg13g2_nor2_1 _14704_ (.A(net200),
    .B(_02017_),
    .Y(_06878_));
 sg13g2_nand2_1 _14705_ (.Y(_06879_),
    .A(net248),
    .B(_02014_));
 sg13g2_xnor2_1 _14706_ (.Y(_06881_),
    .A(_06878_),
    .B(_06879_));
 sg13g2_xnor2_1 _14707_ (.Y(_06882_),
    .A(_06877_),
    .B(_06881_));
 sg13g2_xnor2_1 _14708_ (.Y(_06883_),
    .A(_06872_),
    .B(_06882_));
 sg13g2_nand2_1 _14709_ (.Y(_06884_),
    .A(_06798_),
    .B(net86));
 sg13g2_nand2_1 _14710_ (.Y(_06885_),
    .A(_06794_),
    .B(_06884_));
 sg13g2_o21ai_1 _14711_ (.B1(_06885_),
    .Y(_06886_),
    .A1(_06798_),
    .A2(net86));
 sg13g2_buf_1 _14712_ (.A(_06886_),
    .X(_06887_));
 sg13g2_nand2_1 _14713_ (.Y(_06888_),
    .A(_06765_),
    .B(_06772_));
 sg13g2_nor2_1 _14714_ (.A(_06765_),
    .B(_06772_),
    .Y(_06889_));
 sg13g2_a21oi_2 _14715_ (.B1(_06889_),
    .Y(_06890_),
    .A2(_06888_),
    .A1(_06768_));
 sg13g2_xnor2_1 _14716_ (.Y(_06892_),
    .A(_06887_),
    .B(_06890_));
 sg13g2_xnor2_1 _14717_ (.Y(_06893_),
    .A(_06883_),
    .B(_06892_));
 sg13g2_xor2_1 _14718_ (.B(_06893_),
    .A(_06870_),
    .X(_06894_));
 sg13g2_xnor2_1 _14719_ (.Y(_06895_),
    .A(_06860_),
    .B(_06894_));
 sg13g2_xnor2_1 _14720_ (.Y(_06896_),
    .A(_06855_),
    .B(_06895_));
 sg13g2_xnor2_1 _14721_ (.Y(_06897_),
    .A(_06852_),
    .B(_06896_));
 sg13g2_nand2_1 _14722_ (.Y(_06898_),
    .A(_03254_),
    .B(_06641_));
 sg13g2_xor2_1 _14723_ (.B(_06898_),
    .A(_06897_),
    .X(_06899_));
 sg13g2_xnor2_1 _14724_ (.Y(_06900_),
    .A(_06849_),
    .B(_06899_));
 sg13g2_buf_1 _14725_ (.A(_06900_),
    .X(_06901_));
 sg13g2_a21o_1 _14726_ (.A2(_06821_),
    .A1(_06744_),
    .B1(_06822_),
    .X(_06903_));
 sg13g2_o21ai_1 _14727_ (.B1(_06903_),
    .Y(_06904_),
    .A1(_06744_),
    .A2(_06821_));
 sg13g2_buf_1 _14728_ (.A(_06904_),
    .X(_06905_));
 sg13g2_xor2_1 _14729_ (.B(_06905_),
    .A(_06901_),
    .X(_06906_));
 sg13g2_xnor2_1 _14730_ (.Y(_06907_),
    .A(_06840_),
    .B(_06906_));
 sg13g2_xnor2_1 _14731_ (.Y(_06908_),
    .A(_04091_),
    .B(_06907_));
 sg13g2_xnor2_1 _14732_ (.Y(_06909_),
    .A(_06838_),
    .B(_06908_));
 sg13g2_a21oi_1 _14733_ (.A1(net112),
    .A2(_06909_),
    .Y(_06910_),
    .B1(_05085_));
 sg13g2_mux2_1 _14734_ (.A0(_06910_),
    .A1(_00361_),
    .S(net15),
    .X(_00227_));
 sg13g2_a21o_1 _14735_ (.A2(_06905_),
    .A1(_06901_),
    .B1(_06840_),
    .X(_06911_));
 sg13g2_o21ai_1 _14736_ (.B1(_06911_),
    .Y(_06913_),
    .A1(_06901_),
    .A2(_06905_));
 sg13g2_inv_1 _14737_ (.Y(_06914_),
    .A(_06852_));
 sg13g2_nor2_1 _14738_ (.A(_06914_),
    .B(_06895_),
    .Y(_06915_));
 sg13g2_nand2_1 _14739_ (.Y(_06916_),
    .A(_06914_),
    .B(_06895_));
 sg13g2_o21ai_1 _14740_ (.B1(_06916_),
    .Y(_06917_),
    .A1(_06855_),
    .A2(_06915_));
 sg13g2_buf_1 _14741_ (.A(_06917_),
    .X(_06918_));
 sg13g2_xor2_1 _14742_ (.B(_06870_),
    .A(_06799_),
    .X(_06919_));
 sg13g2_a21o_1 _14743_ (.A2(_06800_),
    .A1(_01267_),
    .B1(_01497_),
    .X(_06920_));
 sg13g2_buf_1 _14744_ (.A(_06920_),
    .X(_06921_));
 sg13g2_nor2_1 _14745_ (.A(_06921_),
    .B(_06870_),
    .Y(_06922_));
 sg13g2_and2_1 _14746_ (.A(_06921_),
    .B(_06870_),
    .X(_06924_));
 sg13g2_mux2_1 _14747_ (.A0(_06922_),
    .A1(_06924_),
    .S(_06799_),
    .X(_06925_));
 sg13g2_a22oi_1 _14748_ (.Y(_06926_),
    .B1(_06925_),
    .B2(_06786_),
    .A2(_06919_),
    .A1(_06893_));
 sg13g2_inv_1 _14749_ (.Y(_06927_),
    .A(_06786_));
 sg13g2_nor2_1 _14750_ (.A(_06922_),
    .B(_06924_),
    .Y(_06928_));
 sg13g2_a21o_1 _14751_ (.A2(_06893_),
    .A1(_06856_),
    .B1(_06927_),
    .X(_06929_));
 sg13g2_a22oi_1 _14752_ (.Y(_06930_),
    .B1(_06928_),
    .B2(_06929_),
    .A2(_06893_),
    .A1(_06927_));
 sg13g2_o21ai_1 _14753_ (.B1(_06930_),
    .Y(_06931_),
    .A1(_06856_),
    .A2(_06926_));
 sg13g2_o21ai_1 _14754_ (.B1(_06786_),
    .Y(_06932_),
    .A1(_06856_),
    .A2(_06928_));
 sg13g2_nand2_1 _14755_ (.Y(_06933_),
    .A(net199),
    .B(net149));
 sg13g2_nand2_1 _14756_ (.Y(_06935_),
    .A(net157),
    .B(_01490_));
 sg13g2_nand2_1 _14757_ (.Y(_06936_),
    .A(net158),
    .B(net176));
 sg13g2_xnor2_1 _14758_ (.Y(_06937_),
    .A(_06935_),
    .B(_06936_));
 sg13g2_xnor2_1 _14759_ (.Y(_06938_),
    .A(_06933_),
    .B(_06937_));
 sg13g2_and2_1 _14760_ (.A(_06874_),
    .B(_06875_),
    .X(_06939_));
 sg13g2_or2_1 _14761_ (.X(_06940_),
    .B(_06875_),
    .A(_06874_));
 sg13g2_o21ai_1 _14762_ (.B1(_06940_),
    .Y(_06941_),
    .A1(_06873_),
    .A2(_06939_));
 sg13g2_nand2_1 _14763_ (.Y(_06942_),
    .A(net127),
    .B(_02188_));
 sg13g2_nand2_1 _14764_ (.Y(_06943_),
    .A(net248),
    .B(net153));
 sg13g2_xnor2_1 _14765_ (.Y(_06944_),
    .A(_06942_),
    .B(_06943_));
 sg13g2_xnor2_1 _14766_ (.Y(_06946_),
    .A(_06941_),
    .B(_06944_));
 sg13g2_xnor2_1 _14767_ (.Y(_06947_),
    .A(_06938_),
    .B(_06946_));
 sg13g2_nor2_1 _14768_ (.A(_06864_),
    .B(_06868_),
    .Y(_06948_));
 sg13g2_a21oi_1 _14769_ (.A1(_06864_),
    .A2(_06868_),
    .Y(_06949_),
    .B1(net86));
 sg13g2_nor2_1 _14770_ (.A(_06948_),
    .B(_06949_),
    .Y(_06950_));
 sg13g2_nand2_1 _14771_ (.Y(_06951_),
    .A(_06877_),
    .B(_06881_));
 sg13g2_o21ai_1 _14772_ (.B1(_06872_),
    .Y(_06952_),
    .A1(_06877_),
    .A2(_06881_));
 sg13g2_nand2_1 _14773_ (.Y(_06953_),
    .A(_06951_),
    .B(_06952_));
 sg13g2_xnor2_1 _14774_ (.Y(_06954_),
    .A(_06950_),
    .B(_06953_));
 sg13g2_xnor2_1 _14775_ (.Y(_06955_),
    .A(_06947_),
    .B(_06954_));
 sg13g2_a21o_1 _14776_ (.A2(net121),
    .A1(net195),
    .B1(_00532_),
    .X(_06957_));
 sg13g2_o21ai_1 _14777_ (.B1(_06957_),
    .Y(_06958_),
    .A1(net195),
    .A2(net121));
 sg13g2_nor3_1 _14778_ (.A(net132),
    .B(net217),
    .C(net133),
    .Y(_06959_));
 sg13g2_nand2b_1 _14779_ (.Y(_06960_),
    .B(net106),
    .A_N(_06959_));
 sg13g2_a21oi_1 _14780_ (.A1(_06665_),
    .A2(_06958_),
    .Y(_06961_),
    .B1(_06960_));
 sg13g2_xnor2_1 _14781_ (.Y(_06962_),
    .A(net86),
    .B(_06961_));
 sg13g2_nand2b_1 _14782_ (.Y(_06963_),
    .B(_06962_),
    .A_N(_06955_));
 sg13g2_nand2b_1 _14783_ (.Y(_06964_),
    .B(_06955_),
    .A_N(_06962_));
 sg13g2_and2_1 _14784_ (.A(_06963_),
    .B(_06964_),
    .X(_06965_));
 sg13g2_xnor2_1 _14785_ (.Y(_06966_),
    .A(_06932_),
    .B(_06965_));
 sg13g2_nor2_1 _14786_ (.A(_06887_),
    .B(_06890_),
    .Y(_06968_));
 sg13g2_nand2_1 _14787_ (.Y(_06969_),
    .A(_06887_),
    .B(_06890_));
 sg13g2_o21ai_1 _14788_ (.B1(_06969_),
    .Y(_06970_),
    .A1(_06883_),
    .A2(_06968_));
 sg13g2_buf_1 _14789_ (.A(_06970_),
    .X(_06971_));
 sg13g2_xnor2_1 _14790_ (.Y(_06972_),
    .A(_06966_),
    .B(_06971_));
 sg13g2_xnor2_1 _14791_ (.Y(_06973_),
    .A(_06931_),
    .B(_06972_));
 sg13g2_nor3_1 _14792_ (.A(_02188_),
    .B(net151),
    .C(_02131_),
    .Y(_06974_));
 sg13g2_xor2_1 _14793_ (.B(_06974_),
    .A(_06973_),
    .X(_06975_));
 sg13g2_xnor2_1 _14794_ (.Y(_06976_),
    .A(_06918_),
    .B(_06975_));
 sg13g2_inv_1 _14795_ (.Y(_06977_),
    .A(_06849_));
 sg13g2_nor2_1 _14796_ (.A(_06977_),
    .B(_06897_),
    .Y(_06979_));
 sg13g2_nand2_1 _14797_ (.Y(_06980_),
    .A(_06977_),
    .B(_06897_));
 sg13g2_o21ai_1 _14798_ (.B1(_06980_),
    .Y(_06981_),
    .A1(_06898_),
    .A2(_06979_));
 sg13g2_xnor2_1 _14799_ (.Y(_06982_),
    .A(_06976_),
    .B(_06981_));
 sg13g2_xnor2_1 _14800_ (.Y(_06983_),
    .A(_04098_),
    .B(_06982_));
 sg13g2_xnor2_1 _14801_ (.Y(_06984_),
    .A(_06913_),
    .B(_06983_));
 sg13g2_nor2_1 _14802_ (.A(_06838_),
    .B(_06908_),
    .Y(_06985_));
 sg13g2_a21oi_1 _14803_ (.A1(_04082_),
    .A2(_06907_),
    .Y(_06986_),
    .B1(_06985_));
 sg13g2_xor2_1 _14804_ (.B(_06986_),
    .A(_06984_),
    .X(_06987_));
 sg13g2_a21oi_1 _14805_ (.A1(net112),
    .A2(_06987_),
    .Y(_06988_),
    .B1(_05096_));
 sg13g2_mux2_1 _14806_ (.A0(_06988_),
    .A1(_02109_),
    .S(net15),
    .X(_00228_));
 sg13g2_nand2b_1 _14807_ (.Y(_06990_),
    .B(_05104_),
    .A_N(_05101_));
 sg13g2_a21oi_1 _14808_ (.A1(net72),
    .A2(_06990_),
    .Y(_06991_),
    .B1(_04097_));
 sg13g2_nand4_1 _14809_ (.B(_04492_),
    .C(_05101_),
    .A(_04097_),
    .Y(_06992_),
    .D(_05104_));
 sg13g2_nor2b_1 _14810_ (.A(_06991_),
    .B_N(_06992_),
    .Y(_06993_));
 sg13g2_o21ai_1 _14811_ (.B1(_04903_),
    .Y(_06994_),
    .A1(_04439_),
    .A2(_06993_));
 sg13g2_xnor2_1 _14812_ (.Y(_06995_),
    .A(_06913_),
    .B(_06982_));
 sg13g2_nand2b_1 _14813_ (.Y(_06996_),
    .B(_06984_),
    .A_N(_06986_));
 sg13g2_o21ai_1 _14814_ (.B1(_06996_),
    .Y(_06997_),
    .A1(_00025_),
    .A2(_06995_));
 sg13g2_inv_1 _14815_ (.Y(_06998_),
    .A(_06981_));
 sg13g2_nand2_1 _14816_ (.Y(_07000_),
    .A(_06976_),
    .B(_06998_));
 sg13g2_a21o_1 _14817_ (.A2(_06901_),
    .A1(_06840_),
    .B1(_06905_),
    .X(_07001_));
 sg13g2_o21ai_1 _14818_ (.B1(_07001_),
    .Y(_07002_),
    .A1(_06840_),
    .A2(_06901_));
 sg13g2_nor2_1 _14819_ (.A(_06976_),
    .B(_06998_),
    .Y(_07003_));
 sg13g2_a21oi_2 _14820_ (.B1(_07003_),
    .Y(_07004_),
    .A2(_07002_),
    .A1(_07000_));
 sg13g2_a21o_1 _14821_ (.A2(_06973_),
    .A1(_06918_),
    .B1(_06974_),
    .X(_07005_));
 sg13g2_o21ai_1 _14822_ (.B1(_07005_),
    .Y(_07006_),
    .A1(_06918_),
    .A2(_06973_));
 sg13g2_nor2_1 _14823_ (.A(_06966_),
    .B(_06971_),
    .Y(_07007_));
 sg13g2_nor2_1 _14824_ (.A(_06931_),
    .B(_07007_),
    .Y(_07008_));
 sg13g2_a21oi_1 _14825_ (.A1(_06966_),
    .A2(_06971_),
    .Y(_07009_),
    .B1(_07008_));
 sg13g2_inv_1 _14826_ (.Y(_07011_),
    .A(_06928_));
 sg13g2_o21ai_1 _14827_ (.B1(_06955_),
    .Y(_07012_),
    .A1(_06856_),
    .A2(_06962_));
 sg13g2_nand2_1 _14828_ (.Y(_07013_),
    .A(_06787_),
    .B(_06962_));
 sg13g2_a221oi_1 _14829_ (.B2(_06964_),
    .C1(_06927_),
    .B1(_07013_),
    .A1(_07011_),
    .Y(_07014_),
    .A2(_07012_));
 sg13g2_a21o_1 _14830_ (.A2(_06963_),
    .A1(_06927_),
    .B1(_07014_),
    .X(_07015_));
 sg13g2_buf_1 _14831_ (.A(_07015_),
    .X(_07016_));
 sg13g2_nand2_1 _14832_ (.Y(_07017_),
    .A(_06786_),
    .B(_07013_));
 sg13g2_a21oi_1 _14833_ (.A1(net132),
    .A2(_00814_),
    .Y(_07018_),
    .B1(_06960_));
 sg13g2_xnor2_1 _14834_ (.Y(_07019_),
    .A(_06921_),
    .B(_07018_));
 sg13g2_nand2_1 _14835_ (.Y(_07020_),
    .A(net128),
    .B(net121));
 sg13g2_nand2_1 _14836_ (.Y(_07022_),
    .A(net157),
    .B(net106));
 sg13g2_nand2_1 _14837_ (.Y(_07023_),
    .A(net120),
    .B(_02054_));
 sg13g2_xnor2_1 _14838_ (.Y(_07024_),
    .A(_07022_),
    .B(_07023_));
 sg13g2_xnor2_1 _14839_ (.Y(_07025_),
    .A(_07020_),
    .B(_07024_));
 sg13g2_buf_1 _14840_ (.A(_07025_),
    .X(_07026_));
 sg13g2_and2_1 _14841_ (.A(_06935_),
    .B(_06936_),
    .X(_07027_));
 sg13g2_or2_1 _14842_ (.X(_07028_),
    .B(_06936_),
    .A(_06935_));
 sg13g2_o21ai_1 _14843_ (.B1(_07028_),
    .Y(_07029_),
    .A1(_06933_),
    .A2(_07027_));
 sg13g2_buf_1 _14844_ (.A(_07029_),
    .X(_07030_));
 sg13g2_nor2_1 _14845_ (.A(net200),
    .B(_02008_),
    .Y(_07031_));
 sg13g2_nand2_1 _14846_ (.Y(_07033_),
    .A(net198),
    .B(_02032_));
 sg13g2_xnor2_1 _14847_ (.Y(_07034_),
    .A(_07031_),
    .B(_07033_));
 sg13g2_xnor2_1 _14848_ (.Y(_07035_),
    .A(_07030_),
    .B(_07034_));
 sg13g2_xnor2_1 _14849_ (.Y(_07036_),
    .A(_07026_),
    .B(_07035_));
 sg13g2_nand2_1 _14850_ (.Y(_07037_),
    .A(_06938_),
    .B(_06944_));
 sg13g2_nor2_1 _14851_ (.A(_06938_),
    .B(_06944_),
    .Y(_07038_));
 sg13g2_a21oi_2 _14852_ (.B1(_07038_),
    .Y(_07039_),
    .A2(_07037_),
    .A1(_06941_));
 sg13g2_nor2_1 _14853_ (.A(net217),
    .B(net133),
    .Y(_07040_));
 sg13g2_nor2_1 _14854_ (.A(net121),
    .B(_07040_),
    .Y(_07041_));
 sg13g2_a21oi_1 _14855_ (.A1(net132),
    .A2(_07041_),
    .Y(_07042_),
    .B1(_06959_));
 sg13g2_a22oi_1 _14856_ (.Y(_07044_),
    .B1(net86),
    .B2(_07042_),
    .A2(_00814_),
    .A1(net132));
 sg13g2_nand2b_1 _14857_ (.Y(_07045_),
    .B(net106),
    .A_N(_07044_));
 sg13g2_xnor2_1 _14858_ (.Y(_07046_),
    .A(_07039_),
    .B(_07045_));
 sg13g2_xnor2_1 _14859_ (.Y(_07047_),
    .A(_07036_),
    .B(_07046_));
 sg13g2_xnor2_1 _14860_ (.Y(_07048_),
    .A(_07019_),
    .B(_07047_));
 sg13g2_xnor2_1 _14861_ (.Y(_07049_),
    .A(_07017_),
    .B(_07048_));
 sg13g2_nand2_1 _14862_ (.Y(_07050_),
    .A(_06950_),
    .B(_06953_));
 sg13g2_o21ai_1 _14863_ (.B1(_06947_),
    .Y(_07051_),
    .A1(_06950_),
    .A2(_06953_));
 sg13g2_nand2_1 _14864_ (.Y(_07052_),
    .A(_07050_),
    .B(_07051_));
 sg13g2_nand3_1 _14865_ (.B(_06641_),
    .C(_07052_),
    .A(_02801_),
    .Y(_07053_));
 sg13g2_buf_1 _14866_ (.A(_07053_),
    .X(_07055_));
 sg13g2_a21oi_1 _14867_ (.A1(_02801_),
    .A2(_06641_),
    .Y(_07056_),
    .B1(_07052_));
 sg13g2_inv_1 _14868_ (.Y(_07057_),
    .A(_07056_));
 sg13g2_nand2_1 _14869_ (.Y(_07058_),
    .A(_07055_),
    .B(_07057_));
 sg13g2_xnor2_1 _14870_ (.Y(_07059_),
    .A(_07049_),
    .B(_07058_));
 sg13g2_xnor2_1 _14871_ (.Y(_07060_),
    .A(_07016_),
    .B(_07059_));
 sg13g2_xnor2_1 _14872_ (.Y(_07061_),
    .A(_07009_),
    .B(_07060_));
 sg13g2_xnor2_1 _14873_ (.Y(_07062_),
    .A(_07006_),
    .B(_07061_));
 sg13g2_xnor2_1 _14874_ (.Y(_07063_),
    .A(_07004_),
    .B(_07062_));
 sg13g2_xor2_1 _14875_ (.B(_07063_),
    .A(_04097_),
    .X(_07064_));
 sg13g2_xnor2_1 _14876_ (.Y(_07066_),
    .A(_06997_),
    .B(_07064_));
 sg13g2_nand2_1 _14877_ (.Y(_07067_),
    .A(net99),
    .B(_07066_));
 sg13g2_a22oi_1 _14878_ (.Y(_00229_),
    .B1(_06994_),
    .B2(_07067_),
    .A2(net14),
    .A1(_00406_));
 sg13g2_a21oi_1 _14879_ (.A1(_07049_),
    .A2(_07055_),
    .Y(_07068_),
    .B1(_07056_));
 sg13g2_nand2_1 _14880_ (.Y(_07069_),
    .A(_07049_),
    .B(_07056_));
 sg13g2_o21ai_1 _14881_ (.B1(_07069_),
    .Y(_07070_),
    .A1(_07016_),
    .A2(_07068_));
 sg13g2_nor2b_1 _14882_ (.A(_07009_),
    .B_N(_07070_),
    .Y(_07071_));
 sg13g2_nor2_1 _14883_ (.A(_07049_),
    .B(_07055_),
    .Y(_07072_));
 sg13g2_nand2_1 _14884_ (.Y(_07073_),
    .A(_07016_),
    .B(_07072_));
 sg13g2_o21ai_1 _14885_ (.B1(_07073_),
    .Y(_07074_),
    .A1(_07016_),
    .A2(_07069_));
 sg13g2_a21oi_1 _14886_ (.A1(_07016_),
    .A2(_07068_),
    .Y(_07076_),
    .B1(_07072_));
 sg13g2_nor2b_1 _14887_ (.A(_07076_),
    .B_N(_07009_),
    .Y(_07077_));
 sg13g2_nor3_1 _14888_ (.A(_07071_),
    .B(_07074_),
    .C(_07077_),
    .Y(_07078_));
 sg13g2_nor2_1 _14889_ (.A(_07039_),
    .B(_07045_),
    .Y(_07079_));
 sg13g2_nand2_1 _14890_ (.Y(_07080_),
    .A(_07039_),
    .B(_07045_));
 sg13g2_o21ai_1 _14891_ (.B1(_07080_),
    .Y(_07081_),
    .A1(_07034_),
    .A2(_07079_));
 sg13g2_nor2_1 _14892_ (.A(_07034_),
    .B(_07080_),
    .Y(_07082_));
 sg13g2_a21oi_1 _14893_ (.A1(_07026_),
    .A2(_07081_),
    .Y(_07083_),
    .B1(_07082_));
 sg13g2_nand2_1 _14894_ (.Y(_07084_),
    .A(_07034_),
    .B(_07079_));
 sg13g2_o21ai_1 _14895_ (.B1(_07084_),
    .Y(_07085_),
    .A1(_07026_),
    .A2(_07081_));
 sg13g2_nor2_1 _14896_ (.A(_07026_),
    .B(_07084_),
    .Y(_07087_));
 sg13g2_a221oi_1 _14897_ (.B2(_07030_),
    .C1(_07087_),
    .B1(_07085_),
    .A1(_07026_),
    .Y(_07088_),
    .A2(_07082_));
 sg13g2_o21ai_1 _14898_ (.B1(_07088_),
    .Y(_07089_),
    .A1(_07030_),
    .A2(_07083_));
 sg13g2_a21oi_1 _14899_ (.A1(net127),
    .A2(_01493_),
    .Y(_07090_),
    .B1(net198));
 sg13g2_a21oi_1 _14900_ (.A1(net127),
    .A2(_02164_),
    .Y(_07091_),
    .B1(net176));
 sg13g2_and3_1 _14901_ (.X(_07092_),
    .A(net176),
    .B(_02164_),
    .C(_06641_));
 sg13g2_nor3_1 _14902_ (.A(_07090_),
    .B(_07091_),
    .C(_07092_),
    .Y(_07093_));
 sg13g2_nand3_1 _14903_ (.B(_02057_),
    .C(net106),
    .A(net202),
    .Y(_07094_));
 sg13g2_a21oi_1 _14904_ (.A1(net128),
    .A2(_07094_),
    .Y(_07095_),
    .B1(_07023_));
 sg13g2_o21ai_1 _14905_ (.B1(_02059_),
    .Y(_07096_),
    .A1(net121),
    .A2(_04563_));
 sg13g2_o21ai_1 _14906_ (.B1(_02077_),
    .Y(_07098_),
    .A1(net128),
    .A2(net157));
 sg13g2_a21oi_1 _14907_ (.A1(_07023_),
    .A2(_07096_),
    .Y(_07099_),
    .B1(_07098_));
 sg13g2_nand2b_1 _14908_ (.Y(_07100_),
    .B(_07099_),
    .A_N(_07095_));
 sg13g2_nand2_1 _14909_ (.Y(_07101_),
    .A(net120),
    .B(_02057_));
 sg13g2_xnor2_1 _14910_ (.Y(_07102_),
    .A(_04097_),
    .B(_07101_));
 sg13g2_xnor2_1 _14911_ (.Y(_07103_),
    .A(_07100_),
    .B(_07102_));
 sg13g2_xnor2_1 _14912_ (.Y(_07104_),
    .A(_07093_),
    .B(_07103_));
 sg13g2_o21ai_1 _14913_ (.B1(net132),
    .Y(_07105_),
    .A1(_00814_),
    .A2(_06802_));
 sg13g2_o21ai_1 _14914_ (.B1(_07105_),
    .Y(_07106_),
    .A1(_06921_),
    .A2(_07040_));
 sg13g2_nand2_1 _14915_ (.Y(_07107_),
    .A(net106),
    .B(_07106_));
 sg13g2_xnor2_1 _14916_ (.Y(_07109_),
    .A(_07104_),
    .B(_07107_));
 sg13g2_xnor2_1 _14917_ (.Y(_07110_),
    .A(_07089_),
    .B(_07109_));
 sg13g2_nand2_1 _14918_ (.Y(_07111_),
    .A(_07019_),
    .B(_07047_));
 sg13g2_o21ai_1 _14919_ (.B1(_07017_),
    .Y(_07112_),
    .A1(_07019_),
    .A2(_07047_));
 sg13g2_nand2_1 _14920_ (.Y(_07113_),
    .A(_07111_),
    .B(_07112_));
 sg13g2_xnor2_1 _14921_ (.Y(_07114_),
    .A(_07110_),
    .B(_07113_));
 sg13g2_xnor2_1 _14922_ (.Y(_07115_),
    .A(_07078_),
    .B(_07114_));
 sg13g2_a21o_1 _14923_ (.A2(_07061_),
    .A1(_07004_),
    .B1(_07006_),
    .X(_07116_));
 sg13g2_o21ai_1 _14924_ (.B1(_07116_),
    .Y(_07117_),
    .A1(_07004_),
    .A2(_07061_));
 sg13g2_xnor2_1 _14925_ (.Y(_07118_),
    .A(_07115_),
    .B(_07117_));
 sg13g2_nand2b_1 _14926_ (.Y(_07120_),
    .B(_07063_),
    .A_N(_06997_));
 sg13g2_nor2b_1 _14927_ (.A(_07063_),
    .B_N(_06997_),
    .Y(_07121_));
 sg13g2_a21oi_1 _14928_ (.A1(_04097_),
    .A2(_07120_),
    .Y(_07122_),
    .B1(_07121_));
 sg13g2_xnor2_1 _14929_ (.Y(_07123_),
    .A(_07118_),
    .B(_07122_));
 sg13g2_nand2_1 _14930_ (.Y(_07124_),
    .A(net99),
    .B(_07123_));
 sg13g2_a22oi_1 _14931_ (.Y(_00230_),
    .B1(_06994_),
    .B2(_07124_),
    .A2(net14),
    .A1(_00363_));
 sg13g2_xor2_1 _14932_ (.B(_06386_),
    .A(_04105_),
    .X(_07125_));
 sg13g2_xnor2_1 _14933_ (.Y(_07126_),
    .A(_06390_),
    .B(_07125_));
 sg13g2_a21oi_1 _14934_ (.A1(net112),
    .A2(_07126_),
    .Y(_07127_),
    .B1(_05113_));
 sg13g2_mux2_1 _14935_ (.A0(_07127_),
    .A1(_05339_),
    .S(net15),
    .X(_00231_));
 sg13g2_nor2b_1 _14936_ (.A(_06393_),
    .B_N(_06394_),
    .Y(_07129_));
 sg13g2_xnor2_1 _14937_ (.Y(_07130_),
    .A(_04108_),
    .B(_07129_));
 sg13g2_a21oi_1 _14938_ (.A1(net112),
    .A2(_07130_),
    .Y(_07131_),
    .B1(_05123_));
 sg13g2_mux2_1 _14939_ (.A0(_07131_),
    .A1(_05317_),
    .S(net15),
    .X(_00232_));
 sg13g2_or2_1 _14940_ (.X(_07132_),
    .B(_06381_),
    .A(_06380_));
 sg13g2_xnor2_1 _14941_ (.Y(_07133_),
    .A(_04112_),
    .B(_06395_));
 sg13g2_xnor2_1 _14942_ (.Y(_07134_),
    .A(_07132_),
    .B(_07133_));
 sg13g2_a21oi_1 _14943_ (.A1(net112),
    .A2(_07134_),
    .Y(_07135_),
    .B1(_05131_));
 sg13g2_mux2_1 _14944_ (.A0(_07135_),
    .A1(_05510_),
    .S(_05012_),
    .X(_00233_));
 sg13g2_xnor2_1 _14945_ (.Y(_07136_),
    .A(_06397_),
    .B(_06402_));
 sg13g2_a21o_1 _14946_ (.A2(_07136_),
    .A1(_06833_),
    .B1(_05138_),
    .X(_07138_));
 sg13g2_nand2_1 _14947_ (.Y(_07139_),
    .A(net196),
    .B(net17));
 sg13g2_o21ai_1 _14948_ (.B1(_07139_),
    .Y(_00234_),
    .A1(net14),
    .A2(_07138_));
 sg13g2_xor2_1 _14949_ (.B(_06377_),
    .A(net317),
    .X(_07140_));
 sg13g2_xnor2_1 _14950_ (.Y(_07141_),
    .A(_06404_),
    .B(_07140_));
 sg13g2_a21oi_1 _14951_ (.A1(_06833_),
    .A2(_07141_),
    .Y(_07142_),
    .B1(_05148_));
 sg13g2_mux2_1 _14952_ (.A0(_07142_),
    .A1(net163),
    .S(net15),
    .X(_00235_));
 sg13g2_xor2_1 _14953_ (.B(_06411_),
    .A(_06407_),
    .X(_07143_));
 sg13g2_nor2_1 _14954_ (.A(net115),
    .B(_07143_),
    .Y(_07144_));
 sg13g2_nor3_1 _14955_ (.A(net17),
    .B(_05156_),
    .C(_07144_),
    .Y(_07145_));
 sg13g2_a21o_1 _14956_ (.A2(net14),
    .A1(_05765_),
    .B1(_07145_),
    .X(_00236_));
 sg13g2_xnor2_1 _14957_ (.Y(_07147_),
    .A(_06373_),
    .B(_06414_));
 sg13g2_xnor2_1 _14958_ (.Y(_07148_),
    .A(_04061_),
    .B(_07147_));
 sg13g2_a21o_1 _14959_ (.A2(_07148_),
    .A1(net112),
    .B1(_05166_),
    .X(_07149_));
 sg13g2_nand2_1 _14960_ (.Y(_07150_),
    .A(net162),
    .B(_04717_));
 sg13g2_o21ai_1 _14961_ (.B1(_07150_),
    .Y(_00237_),
    .A1(net14),
    .A2(_07149_));
 sg13g2_nand3_1 _14962_ (.B(_06416_),
    .C(_06518_),
    .A(_06415_),
    .Y(_07151_));
 sg13g2_a21oi_1 _14963_ (.A1(_06521_),
    .A2(_07151_),
    .Y(_07152_),
    .B1(net141));
 sg13g2_nor3_1 _14964_ (.A(net17),
    .B(_05174_),
    .C(_07152_),
    .Y(_07153_));
 sg13g2_a21o_1 _14965_ (.A2(net14),
    .A1(_05801_),
    .B1(_07153_),
    .X(_00238_));
 sg13g2_nand2_1 _14966_ (.Y(_07155_),
    .A(_06521_),
    .B(_06522_));
 sg13g2_and2_1 _14967_ (.A(_06625_),
    .B(_06626_),
    .X(_07156_));
 sg13g2_xnor2_1 _14968_ (.Y(_07157_),
    .A(_07155_),
    .B(_07156_));
 sg13g2_nor2_1 _14969_ (.A(net141),
    .B(_07157_),
    .Y(_07158_));
 sg13g2_or2_1 _14970_ (.X(_07159_),
    .B(_07158_),
    .A(_05184_));
 sg13g2_nand2_1 _14971_ (.Y(_07160_),
    .A(_04801_),
    .B(_04717_));
 sg13g2_o21ai_1 _14972_ (.B1(_07160_),
    .Y(_00239_),
    .A1(_04718_),
    .A2(_07159_));
 sg13g2_nand2_1 _14973_ (.Y(_07161_),
    .A(_03737_),
    .B(net17));
 sg13g2_o21ai_1 _14974_ (.B1(_07161_),
    .Y(_00163_),
    .A1(_03737_),
    .A2(_04903_));
 sg13g2_nand2_1 _14975_ (.Y(_07162_),
    .A(_03737_),
    .B(_04713_));
 sg13g2_a21o_1 _14976_ (.A2(_07162_),
    .A1(net112),
    .B1(net48),
    .X(_07164_));
 sg13g2_nor3_1 _14977_ (.A(_03833_),
    .B(_03738_),
    .C(_04903_),
    .Y(_07165_));
 sg13g2_a21o_1 _14978_ (.A2(_07164_),
    .A1(_03738_),
    .B1(_07165_),
    .X(_00164_));
 sg13g2_or2_1 _14979_ (.X(_07166_),
    .B(_03853_),
    .A(_03736_));
 sg13g2_a21oi_1 _14980_ (.A1(net99),
    .A2(_07166_),
    .Y(_07167_),
    .B1(net48));
 sg13g2_or4_1 _14981_ (.A(\iter[2] ),
    .B(net115),
    .C(net48),
    .D(_07166_),
    .X(_07168_));
 sg13g2_o21ai_1 _14982_ (.B1(_07168_),
    .Y(_00165_),
    .A1(_03854_),
    .A2(_07167_));
 sg13g2_a21oi_1 _14983_ (.A1(net99),
    .A2(_03822_),
    .Y(_07169_),
    .B1(net48));
 sg13g2_or4_1 _14984_ (.A(_04449_),
    .B(net115),
    .C(net55),
    .D(_03822_),
    .X(_07170_));
 sg13g2_o21ai_1 _14985_ (.B1(_07170_),
    .Y(_00166_),
    .A1(_04458_),
    .A2(_07169_));
 sg13g2_and3_1 _14986_ (.X(_00167_),
    .A(net273),
    .B(_00044_),
    .C(net99));
 sg13g2_xnor2_1 _14987_ (.Y(_07172_),
    .A(\step[1] ),
    .B(\step[0] ));
 sg13g2_nor2_1 _14988_ (.A(net220),
    .B(_07172_),
    .Y(_00168_));
 sg13g2_xnor2_1 _14989_ (.Y(_07173_),
    .A(_03903_),
    .B(_03924_));
 sg13g2_nor2_1 _14990_ (.A(net220),
    .B(_07173_),
    .Y(_00169_));
 sg13g2_nand2_1 _14991_ (.Y(_07174_),
    .A(_03903_),
    .B(_03924_));
 sg13g2_xor2_1 _14992_ (.B(_07174_),
    .A(\step[3] ),
    .X(_07175_));
 sg13g2_nor2_1 _14993_ (.A(net220),
    .B(_07175_),
    .Y(_00170_));
 sg13g2_nand3_1 _14994_ (.B(_03852_),
    .C(_03860_),
    .A(_03829_),
    .Y(_07176_));
 sg13g2_nor3_1 _14995_ (.A(_00029_),
    .B(_03857_),
    .C(_03858_),
    .Y(_07177_));
 sg13g2_o21ai_1 _14996_ (.B1(_00015_),
    .Y(_07179_),
    .A1(_00030_),
    .A2(_07177_));
 sg13g2_a21oi_1 _14997_ (.A1(_07176_),
    .A2(_07179_),
    .Y(_00171_),
    .B1(_00000_));
 sg13g2_nor3_1 _14998_ (.A(_03829_),
    .B(_00029_),
    .C(_00031_),
    .Y(_07180_));
 sg13g2_a21oi_1 _14999_ (.A1(_03843_),
    .A2(_03860_),
    .Y(_07181_),
    .B1(_00015_));
 sg13g2_nor3_1 _15000_ (.A(_03843_),
    .B(_03852_),
    .C(_03860_),
    .Y(_07182_));
 sg13g2_nor4_1 _15001_ (.A(_00000_),
    .B(_07180_),
    .C(_07181_),
    .D(_07182_),
    .Y(_00172_));
 sg13g2_inv_1 _15002_ (.Y(_07183_),
    .A(_00000_));
 sg13g2_nand2_1 _15003_ (.Y(_07184_),
    .A(_00030_),
    .B(_07177_));
 sg13g2_o21ai_1 _15004_ (.B1(_00029_),
    .Y(_07185_),
    .A1(_03825_),
    .A2(_03828_));
 sg13g2_nand2b_1 _15005_ (.Y(_07186_),
    .B(_00030_),
    .A_N(_07185_));
 sg13g2_mux2_1 _15006_ (.A0(_00015_),
    .A1(_07185_),
    .S(_00031_),
    .X(_07188_));
 sg13g2_and4_1 _15007_ (.A(_07183_),
    .B(_07184_),
    .C(_07186_),
    .D(_07188_),
    .X(_00173_));
 sg13g2_nand2_1 _15008_ (.Y(_07189_),
    .A(_03843_),
    .B(_03852_));
 sg13g2_nand3_1 _15009_ (.B(_00031_),
    .C(_07189_),
    .A(_03829_),
    .Y(_07190_));
 sg13g2_a21o_1 _15010_ (.A2(_04439_),
    .A1(_00032_),
    .B1(_03857_),
    .X(_07191_));
 sg13g2_nand2_1 _15011_ (.Y(_07192_),
    .A(_00015_),
    .B(_07191_));
 sg13g2_a21oi_1 _15012_ (.A1(_07190_),
    .A2(_07192_),
    .Y(_00174_),
    .B1(_00000_));
 sg13g2_xnor2_1 _15013_ (.Y(_07193_),
    .A(_00029_),
    .B(_00031_));
 sg13g2_and2_1 _15014_ (.A(_04458_),
    .B(_03822_),
    .X(_07194_));
 sg13g2_nor3_1 _15015_ (.A(\last_iter[4] ),
    .B(\last_iter[3] ),
    .C(_03841_),
    .Y(_07195_));
 sg13g2_a21oi_1 _15016_ (.A1(_03841_),
    .A2(_07194_),
    .Y(_07197_),
    .B1(_07195_));
 sg13g2_a21oi_1 _15017_ (.A1(_03852_),
    .A2(_07193_),
    .Y(_00175_),
    .B1(_07197_));
 sg13g2_nor3_1 _15018_ (.A(_03843_),
    .B(_03852_),
    .C(_07191_),
    .Y(_07198_));
 sg13g2_nor2_1 _15019_ (.A(_07197_),
    .B(_07198_),
    .Y(_00176_));
 sg13g2_nor4_1 _15020_ (.A(_03871_),
    .B(_03872_),
    .C(\i_coord.demo_update_delay ),
    .D(_04005_),
    .Y(_07199_));
 sg13g2_and2_1 _15021_ (.A(net66),
    .B(_07199_),
    .X(_00045_));
 sg13g2_nand2b_1 _15022_ (.Y(_07200_),
    .B(\i_coord.demo_update_delay ),
    .A_N(_04144_));
 sg13g2_nand2_1 _15023_ (.Y(_07201_),
    .A(_00001_),
    .B(net66));
 sg13g2_a21oi_1 _15024_ (.A1(_07200_),
    .A2(_07201_),
    .Y(_00046_),
    .B1(_03926_));
 sg13g2_nand3_1 _15025_ (.B(_03872_),
    .C(_03870_),
    .A(_03871_),
    .Y(_07202_));
 sg13g2_buf_1 _15026_ (.A(_07202_),
    .X(_07204_));
 sg13g2_buf_1 _15027_ (.A(_07204_),
    .X(_07205_));
 sg13g2_mux2_1 _15028_ (.A0(_03869_),
    .A1(_03886_),
    .S(_07205_),
    .X(_07206_));
 sg13g2_nand3_1 _15029_ (.B(_03886_),
    .C(_03898_),
    .A(_03885_),
    .Y(_07207_));
 sg13g2_o21ai_1 _15030_ (.B1(_07207_),
    .Y(_07208_),
    .A1(net221),
    .A2(_07206_));
 sg13g2_nand2_1 _15031_ (.Y(_00119_),
    .A(net224),
    .B(_07208_));
 sg13g2_nand2_1 _15032_ (.Y(_07209_),
    .A(_03894_),
    .B(net218));
 sg13g2_o21ai_1 _15033_ (.B1(_07209_),
    .Y(_07210_),
    .A1(_03915_),
    .A2(_07205_));
 sg13g2_nand2_1 _15034_ (.Y(_07211_),
    .A(_03885_),
    .B(_03932_));
 sg13g2_o21ai_1 _15035_ (.B1(_07211_),
    .Y(_07212_),
    .A1(_03950_),
    .A2(_07210_));
 sg13g2_nand2_1 _15036_ (.Y(_00120_),
    .A(net224),
    .B(_07212_));
 sg13g2_mux2_1 _15037_ (.A0(_03927_),
    .A1(_03887_),
    .S(net218),
    .X(_07214_));
 sg13g2_a22oi_1 _15038_ (.Y(_07215_),
    .B1(_07214_),
    .B2(_03930_),
    .A2(_03939_),
    .A1(_03901_));
 sg13g2_nor2_1 _15039_ (.A(_03961_),
    .B(_07215_),
    .Y(_00121_));
 sg13g2_o21ai_1 _15040_ (.B1(_03882_),
    .Y(_07216_),
    .A1(_03942_),
    .A2(net218));
 sg13g2_nor2b_1 _15041_ (.A(_03947_),
    .B_N(_07216_),
    .Y(_07217_));
 sg13g2_inv_1 _15042_ (.Y(_07218_),
    .A(_07204_));
 sg13g2_nor3_1 _15043_ (.A(net225),
    .B(_03888_),
    .C(_07218_),
    .Y(_07219_));
 sg13g2_o21ai_1 _15044_ (.B1(_03923_),
    .Y(_00122_),
    .A1(_07217_),
    .A2(_07219_));
 sg13g2_mux2_1 _15045_ (.A0(_03951_),
    .A1(_03890_),
    .S(net218),
    .X(_07220_));
 sg13g2_nand2_1 _15046_ (.Y(_07222_),
    .A(_03900_),
    .B(_03955_));
 sg13g2_o21ai_1 _15047_ (.B1(_07222_),
    .Y(_07223_),
    .A1(_03950_),
    .A2(_07220_));
 sg13g2_nand2_1 _15048_ (.Y(_00123_),
    .A(_03923_),
    .B(_07223_));
 sg13g2_mux2_1 _15049_ (.A0(_03958_),
    .A1(_03889_),
    .S(net218),
    .X(_07224_));
 sg13g2_nand2_1 _15050_ (.Y(_07225_),
    .A(_03900_),
    .B(_03963_));
 sg13g2_o21ai_1 _15051_ (.B1(_07225_),
    .Y(_07226_),
    .A1(net221),
    .A2(_07224_));
 sg13g2_nand2_1 _15052_ (.Y(_00124_),
    .A(net224),
    .B(_07226_));
 sg13g2_nand2_1 _15053_ (.Y(_07227_),
    .A(_03891_),
    .B(net218));
 sg13g2_o21ai_1 _15054_ (.B1(_07227_),
    .Y(_07228_),
    .A1(_03966_),
    .A2(net218));
 sg13g2_xnor2_1 _15055_ (.Y(_07229_),
    .A(_03891_),
    .B(_03909_));
 sg13g2_a22oi_1 _15056_ (.Y(_07231_),
    .B1(_07229_),
    .B2(net89),
    .A2(_07228_),
    .A1(net223));
 sg13g2_nor2_1 _15057_ (.A(_03961_),
    .B(_07231_),
    .Y(_00125_));
 sg13g2_nor2_1 _15058_ (.A(_03970_),
    .B(net218),
    .Y(_07232_));
 sg13g2_nor2_1 _15059_ (.A(_03895_),
    .B(_07218_),
    .Y(_07233_));
 sg13g2_o21ai_1 _15060_ (.B1(net222),
    .Y(_07234_),
    .A1(_07232_),
    .A2(_07233_));
 sg13g2_o21ai_1 _15061_ (.B1(_07234_),
    .Y(_07235_),
    .A1(_03936_),
    .A2(_03931_));
 sg13g2_nand2_1 _15062_ (.Y(_00126_),
    .A(net224),
    .B(_07235_));
 sg13g2_nand2_1 _15063_ (.Y(_07236_),
    .A(_03861_),
    .B(_03924_));
 sg13g2_nand2_2 _15064_ (.Y(_07237_),
    .A(\step[1] ),
    .B(\step[0] ));
 sg13g2_nand2_1 _15065_ (.Y(_07238_),
    .A(_03964_),
    .B(_07237_));
 sg13g2_buf_1 _15066_ (.A(_04118_),
    .X(_07240_));
 sg13g2_nand2b_1 _15067_ (.Y(_07241_),
    .B(net320),
    .A_N(net96));
 sg13g2_buf_1 _15068_ (.A(_07241_),
    .X(_07242_));
 sg13g2_a21oi_1 _15069_ (.A1(_07236_),
    .A2(_07238_),
    .Y(_00142_),
    .B1(_07242_));
 sg13g2_nor2_1 _15070_ (.A(net272),
    .B(net96),
    .Y(_07243_));
 sg13g2_nand3_1 _15071_ (.B(net336),
    .C(_04014_),
    .A(_04041_),
    .Y(_07244_));
 sg13g2_nor3_1 _15072_ (.A(_04317_),
    .B(_03864_),
    .C(_07244_),
    .Y(_07245_));
 sg13g2_nand3_1 _15073_ (.B(_04027_),
    .C(_07245_),
    .A(_04081_),
    .Y(_07246_));
 sg13g2_xor2_1 _15074_ (.B(_07246_),
    .A(_04034_),
    .X(_07247_));
 sg13g2_nand2_1 _15075_ (.Y(_00143_),
    .A(_07243_),
    .B(_07247_));
 sg13g2_xor2_1 _15076_ (.B(_04308_),
    .A(_03954_),
    .X(_07249_));
 sg13g2_nor2_1 _15077_ (.A(_07242_),
    .B(_07249_),
    .Y(_00144_));
 sg13g2_nand3_1 _15078_ (.B(_03964_),
    .C(_03924_),
    .A(_03954_),
    .Y(_07250_));
 sg13g2_xor2_1 _15079_ (.B(_07250_),
    .A(_03974_),
    .X(_07251_));
 sg13g2_nor2_1 _15080_ (.A(net220),
    .B(_07251_),
    .Y(_00145_));
 sg13g2_xnor2_1 _15081_ (.Y(_07252_),
    .A(_00027_),
    .B(_03992_));
 sg13g2_nor3_1 _15082_ (.A(_07237_),
    .B(net96),
    .C(_07252_),
    .Y(_07253_));
 sg13g2_a21oi_1 _15083_ (.A1(_03998_),
    .A2(_07237_),
    .Y(_07254_),
    .B1(_07253_));
 sg13g2_nor2_1 _15084_ (.A(net220),
    .B(_07254_),
    .Y(_00146_));
 sg13g2_xnor2_1 _15085_ (.Y(_07255_),
    .A(_04041_),
    .B(_04014_));
 sg13g2_nand2_1 _15086_ (.Y(_00147_),
    .A(net224),
    .B(_07255_));
 sg13g2_nand2_1 _15087_ (.Y(_07257_),
    .A(_03954_),
    .B(_03974_));
 sg13g2_nor4_1 _15088_ (.A(_04050_),
    .B(_03861_),
    .C(_07257_),
    .D(_04007_),
    .Y(_07258_));
 sg13g2_xnor2_1 _15089_ (.Y(_07259_),
    .A(net336),
    .B(_07258_));
 sg13g2_nor2_1 _15090_ (.A(_07242_),
    .B(_07259_),
    .Y(_00148_));
 sg13g2_xor2_1 _15091_ (.B(_07244_),
    .A(_04071_),
    .X(_07260_));
 sg13g2_nand2_1 _15092_ (.Y(_00149_),
    .A(_07243_),
    .B(_07260_));
 sg13g2_nand4_1 _15093_ (.B(_04041_),
    .C(net336),
    .A(_03998_),
    .Y(_07261_),
    .D(_04071_));
 sg13g2_nor2_1 _15094_ (.A(_03992_),
    .B(_07261_),
    .Y(_07262_));
 sg13g2_xnor2_1 _15095_ (.Y(_07263_),
    .A(_00028_),
    .B(_07262_));
 sg13g2_nor2_1 _15096_ (.A(_07237_),
    .B(net96),
    .Y(_07265_));
 sg13g2_a22oi_1 _15097_ (.Y(_07266_),
    .B1(_07263_),
    .B2(_07265_),
    .A2(_07237_),
    .A1(_04060_));
 sg13g2_nor2_1 _15098_ (.A(net220),
    .B(_07266_),
    .Y(_00150_));
 sg13g2_or2_1 _15099_ (.X(_07267_),
    .B(_07245_),
    .A(_04027_));
 sg13g2_nand2_1 _15100_ (.Y(_07268_),
    .A(_04027_),
    .B(_07245_));
 sg13g2_a21o_1 _15101_ (.A2(_07268_),
    .A1(_07267_),
    .B1(_07242_),
    .X(_00151_));
 sg13g2_xor2_1 _15102_ (.B(_07268_),
    .A(_04081_),
    .X(_07269_));
 sg13g2_nand2_1 _15103_ (.Y(_00152_),
    .A(_07243_),
    .B(_07269_));
 sg13g2_nor3_1 _15104_ (.A(_04155_),
    .B(_04166_),
    .C(_04199_),
    .Y(_07270_));
 sg13g2_nand3_1 _15105_ (.B(_04136_),
    .C(net96),
    .A(_04127_),
    .Y(_07271_));
 sg13g2_nor2_1 _15106_ (.A(_04251_),
    .B(_07271_),
    .Y(_07273_));
 sg13g2_and2_1 _15107_ (.A(\i_vga.timing_ver.counter[4] ),
    .B(_07273_),
    .X(_07274_));
 sg13g2_buf_1 _15108_ (.A(_07274_),
    .X(_07275_));
 sg13g2_a21oi_1 _15109_ (.A1(_07270_),
    .A2(_07275_),
    .Y(_07276_),
    .B1(net272));
 sg13g2_buf_1 _15110_ (.A(_07276_),
    .X(_07277_));
 sg13g2_nand2b_1 _15111_ (.Y(_07278_),
    .B(net96),
    .A_N(_00017_));
 sg13g2_o21ai_1 _15112_ (.B1(_07278_),
    .Y(_07279_),
    .A1(_04127_),
    .A2(_07240_));
 sg13g2_nand2_1 _15113_ (.Y(_00153_),
    .A(net45),
    .B(_07279_));
 sg13g2_nand3b_1 _15114_ (.B(net96),
    .C(net45),
    .Y(_07280_),
    .A_N(_04127_));
 sg13g2_and2_1 _15115_ (.A(_07242_),
    .B(_07280_),
    .X(_07281_));
 sg13g2_nand4_1 _15116_ (.B(_04145_),
    .C(net96),
    .A(_04127_),
    .Y(_07283_),
    .D(_07277_));
 sg13g2_o21ai_1 _15117_ (.B1(_07283_),
    .Y(_00154_),
    .A1(_04145_),
    .A2(_07281_));
 sg13g2_xor2_1 _15118_ (.B(_07271_),
    .A(_04241_),
    .X(_07284_));
 sg13g2_nand2_1 _15119_ (.Y(_00155_),
    .A(net45),
    .B(_07284_));
 sg13g2_nand4_1 _15120_ (.B(_04136_),
    .C(_04241_),
    .A(_04127_),
    .Y(_07285_),
    .D(_07240_));
 sg13g2_xor2_1 _15121_ (.B(_07285_),
    .A(\i_vga.timing_ver.counter[3] ),
    .X(_07286_));
 sg13g2_nand2_1 _15122_ (.Y(_00156_),
    .A(net45),
    .B(_07286_));
 sg13g2_xnor2_1 _15123_ (.Y(_07287_),
    .A(\i_vga.timing_ver.counter[4] ),
    .B(_07273_));
 sg13g2_nor2_1 _15124_ (.A(net220),
    .B(_07287_),
    .Y(_00157_));
 sg13g2_xnor2_1 _15125_ (.Y(_07288_),
    .A(_04155_),
    .B(_07275_));
 sg13g2_nand2_1 _15126_ (.Y(_00158_),
    .A(net224),
    .B(_07288_));
 sg13g2_nand2_1 _15127_ (.Y(_07290_),
    .A(_04155_),
    .B(_07275_));
 sg13g2_xor2_1 _15128_ (.B(_07290_),
    .A(_04177_),
    .X(_07291_));
 sg13g2_nand2_1 _15129_ (.Y(_00159_),
    .A(net45),
    .B(_07291_));
 sg13g2_nand3_1 _15130_ (.B(_04177_),
    .C(_07275_),
    .A(_04155_),
    .Y(_07292_));
 sg13g2_xor2_1 _15131_ (.B(_07292_),
    .A(\i_vga.timing_ver.counter[7] ),
    .X(_07293_));
 sg13g2_nand2_1 _15132_ (.Y(_00160_),
    .A(net45),
    .B(_07293_));
 sg13g2_nand4_1 _15133_ (.B(\i_vga.timing_ver.counter[7] ),
    .C(_04177_),
    .A(_04155_),
    .Y(_07294_),
    .D(_07275_));
 sg13g2_xor2_1 _15134_ (.B(_07294_),
    .A(\i_vga.timing_ver.counter[8] ),
    .X(_07295_));
 sg13g2_nand2_1 _15135_ (.Y(_00161_),
    .A(net45),
    .B(_07295_));
 sg13g2_nor2_1 _15136_ (.A(_04199_),
    .B(_07290_),
    .Y(_07297_));
 sg13g2_xnor2_1 _15137_ (.Y(_07298_),
    .A(_04166_),
    .B(_07297_));
 sg13g2_nand2_1 _15138_ (.Y(_00162_),
    .A(net45),
    .B(_07298_));
 sg13g2_o21ai_1 _15139_ (.B1(\i_vga.timing_ver.counter[3] ),
    .Y(_07299_),
    .A1(_04136_),
    .A2(_04241_));
 sg13g2_inv_1 _15140_ (.Y(_07300_),
    .A(_07299_));
 sg13g2_nor3_1 _15141_ (.A(_00016_),
    .B(_04231_),
    .C(_07300_),
    .Y(\i_vga.timing_ver.sync_tmp ));
 sg13g2_buf_1 _15142_ (.A(_04166_),
    .X(\i_vga.timing_ver.blank ));
 sg13g2_and2_1 _15143_ (.A(\video_colour[5] ),
    .B(net65),
    .X(net6));
 sg13g2_and2_1 _15144_ (.A(\video_colour[3] ),
    .B(net65),
    .X(net7));
 sg13g2_and2_1 _15145_ (.A(\video_colour[1] ),
    .B(net65),
    .X(net8));
 sg13g2_and2_1 _15146_ (.A(\video_colour[4] ),
    .B(net65),
    .X(net10));
 sg13g2_and2_1 _15147_ (.A(\video_colour[2] ),
    .B(net65),
    .X(net11));
 sg13g2_and2_1 _15148_ (.A(\video_colour[0] ),
    .B(net65),
    .X(net12));
 sg13g2_buf_4 clkbuf_leaf_0_clk (.X(clknet_leaf_0_clk),
    .A(clknet_2_1__leaf_clk));
 sg13g2_tiehi \i_coord.demo_update$_SDFF_PN0__353  (.L_HI(net353));
 sg13g2_buf_1 _15151_ (.A(net337),
    .X(uio_oe[0]));
 sg13g2_buf_1 _15152_ (.A(net338),
    .X(uio_oe[1]));
 sg13g2_buf_1 _15153_ (.A(net339),
    .X(uio_oe[2]));
 sg13g2_buf_1 _15154_ (.A(net340),
    .X(uio_oe[3]));
 sg13g2_buf_1 _15155_ (.A(net341),
    .X(uio_oe[4]));
 sg13g2_buf_1 _15156_ (.A(net342),
    .X(uio_oe[5]));
 sg13g2_buf_1 _15157_ (.A(net343),
    .X(uio_oe[6]));
 sg13g2_buf_1 _15158_ (.A(net344),
    .X(uio_oe[7]));
 sg13g2_buf_1 _15159_ (.A(net345),
    .X(uio_out[0]));
 sg13g2_buf_1 _15160_ (.A(net346),
    .X(uio_out[1]));
 sg13g2_buf_1 _15161_ (.A(net347),
    .X(uio_out[2]));
 sg13g2_buf_1 _15162_ (.A(net348),
    .X(uio_out[3]));
 sg13g2_buf_1 _15163_ (.A(net349),
    .X(uio_out[4]));
 sg13g2_buf_1 _15164_ (.A(net350),
    .X(uio_out[5]));
 sg13g2_buf_1 _15165_ (.A(net351),
    .X(uio_out[6]));
 sg13g2_buf_1 _15166_ (.A(net352),
    .X(uio_out[7]));
 sg13g2_buf_1 _15167_ (.A(\i_vga.timing_ver.sync ),
    .X(net9));
 sg13g2_buf_1 _15168_ (.A(\i_vga.hsync ),
    .X(net13));
 sg13g2_dfrbp_1 \i_coord.demo_update$_SDFF_PN0_  (.CLK(clknet_leaf_12_clk),
    .RESET_B(net353),
    .D(_00045_),
    .Q_N(_00014_),
    .Q(\i_coord.demo_update ));
 sg13g2_dfrbp_1 \i_coord.demo_update_delay$_SDFFE_PN0P_  (.CLK(clknet_leaf_13_clk),
    .RESET_B(net354),
    .D(_00046_),
    .Q_N(_00001_),
    .Q(\i_coord.demo_update_delay ));
 sg13g2_dfrbp_1 \i_coord.l_xip.state[0]$_SDFFCE_PP0P_  (.CLK(clknet_leaf_14_clk),
    .RESET_B(net355),
    .D(_00047_),
    .Q_N(_07668_),
    .Q(\i_coord.l_xip.data_out[0] ));
 sg13g2_dfrbp_1 \i_coord.l_xip.state[1]$_SDFFCE_PN1P_  (.CLK(clknet_leaf_12_clk),
    .RESET_B(net356),
    .D(_00048_),
    .Q_N(_07667_),
    .Q(\i_coord.l_xip.data_out[1] ));
 sg13g2_dfrbp_1 \i_coord.l_xip.state[2]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_13_clk),
    .RESET_B(net357),
    .D(_00049_),
    .Q_N(_07666_),
    .Q(\i_coord.l_xip.data_out[2] ));
 sg13g2_dfrbp_1 \i_coord.l_xip.state[3]$_SDFFCE_PN1P_  (.CLK(clknet_leaf_13_clk),
    .RESET_B(net358),
    .D(_00050_),
    .Q_N(_07665_),
    .Q(\i_coord.l_xip.data_out[3] ));
 sg13g2_dfrbp_1 \i_coord.l_xip.state[4]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_13_clk),
    .RESET_B(net359),
    .D(_00051_),
    .Q_N(_07664_),
    .Q(\i_coord.l_xip.data_out[4] ));
 sg13g2_dfrbp_1 \i_coord.l_xip.state[5]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_13_clk),
    .RESET_B(net360),
    .D(_00052_),
    .Q_N(_07663_),
    .Q(\i_coord.l_xip.data_out[5] ));
 sg13g2_dfrbp_1 \i_coord.l_xip.state[6]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_14_clk),
    .RESET_B(net361),
    .D(_00053_),
    .Q_N(_07662_),
    .Q(\i_coord.l_xip.data_out[6] ));
 sg13g2_dfrbp_1 \i_coord.l_xip.state[7]$_SDFFCE_PN1P_  (.CLK(clknet_leaf_14_clk),
    .RESET_B(net362),
    .D(_00054_),
    .Q_N(_07661_),
    .Q(\i_coord.l_xip.data_out[7] ));
 sg13g2_dfrbp_1 \i_coord.l_xip.state[8]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_14_clk),
    .RESET_B(net363),
    .D(_00055_),
    .Q_N(_07660_),
    .Q(\i_coord.l_xip.data_out[8] ));
 sg13g2_dfrbp_1 \i_coord.l_xip.state[9]$_SDFFCE_PP0P_  (.CLK(clknet_leaf_13_clk),
    .RESET_B(net364),
    .D(_00056_),
    .Q_N(_07659_),
    .Q(\i_coord.l_xip.data_out[9] ));
 sg13g2_dfrbp_1 \i_coord.l_xir.state[0]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_19_clk),
    .RESET_B(net365),
    .D(_00057_),
    .Q_N(_07658_),
    .Q(\i_coord.l_xir.data_out[0] ));
 sg13g2_dfrbp_1 \i_coord.l_xir.state[1]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_19_clk),
    .RESET_B(net366),
    .D(_00058_),
    .Q_N(_07657_),
    .Q(\i_coord.l_xir.data_out[1] ));
 sg13g2_dfrbp_1 \i_coord.l_xir.state[2]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_19_clk),
    .RESET_B(net367),
    .D(_00059_),
    .Q_N(_07656_),
    .Q(\i_coord.l_xir.data_out[2] ));
 sg13g2_dfrbp_1 \i_coord.l_xir.state[3]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_18_clk),
    .RESET_B(net368),
    .D(_00060_),
    .Q_N(_07655_),
    .Q(\i_coord.l_xir.data_out[3] ));
 sg13g2_dfrbp_1 \i_coord.l_xir.state[4]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_14_clk),
    .RESET_B(net369),
    .D(_00061_),
    .Q_N(_07654_),
    .Q(\i_coord.l_xir.data_out[4] ));
 sg13g2_dfrbp_1 \i_coord.l_xir.state[5]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_16_clk),
    .RESET_B(net370),
    .D(_00062_),
    .Q_N(_07653_),
    .Q(\i_coord.l_xir.data_out[5] ));
 sg13g2_dfrbp_1 \i_coord.l_xir.state[6]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_17_clk),
    .RESET_B(net371),
    .D(_00063_),
    .Q_N(_07652_),
    .Q(\i_coord.l_xir.data_out[6] ));
 sg13g2_dfrbp_1 \i_coord.l_xir.state[7]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_18_clk),
    .RESET_B(net372),
    .D(_00064_),
    .Q_N(_07651_),
    .Q(\i_coord.l_xir.data_out[7] ));
 sg13g2_dfrbp_1 \i_coord.l_xl.state[10]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_16_clk),
    .RESET_B(net373),
    .D(_00065_),
    .Q_N(_07650_),
    .Q(\i_coord.l_xl.data_out[10] ));
 sg13g2_dfrbp_1 \i_coord.l_xl.state[11]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_16_clk),
    .RESET_B(net374),
    .D(_00066_),
    .Q_N(_07649_),
    .Q(\i_coord.l_xl.data_out[11] ));
 sg13g2_dfrbp_1 \i_coord.l_xl.state[12]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_16_clk),
    .RESET_B(net375),
    .D(_00067_),
    .Q_N(_07648_),
    .Q(\i_coord.l_xl.data_out[12] ));
 sg13g2_dfrbp_1 \i_coord.l_xl.state[13]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_15_clk),
    .RESET_B(net376),
    .D(_00068_),
    .Q_N(_07647_),
    .Q(\i_coord.l_xl.data_out[13] ));
 sg13g2_dfrbp_1 \i_coord.l_xl.state[14]$_SDFFCE_PN1P_  (.CLK(clknet_leaf_20_clk),
    .RESET_B(net377),
    .D(_00069_),
    .Q_N(_07646_),
    .Q(\i_coord.l_xl.data_out[14] ));
 sg13g2_dfrbp_1 \i_coord.l_xl.state[15]$_SDFFCE_PN1P_  (.CLK(clknet_leaf_16_clk),
    .RESET_B(net378),
    .D(_00070_),
    .Q_N(_07645_),
    .Q(\i_coord.l_xl.data_out[15] ));
 sg13g2_dfrbp_1 \i_coord.l_xl.state[3]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_17_clk),
    .RESET_B(net379),
    .D(_00071_),
    .Q_N(_07644_),
    .Q(\i_coord.l_xl.data_out[3] ));
 sg13g2_dfrbp_1 \i_coord.l_xl.state[4]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_16_clk),
    .RESET_B(net380),
    .D(_00072_),
    .Q_N(_07643_),
    .Q(\i_coord.l_xl.data_out[4] ));
 sg13g2_dfrbp_1 \i_coord.l_xl.state[5]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_17_clk),
    .RESET_B(net381),
    .D(_00073_),
    .Q_N(_07642_),
    .Q(\i_coord.l_xl.data_out[5] ));
 sg13g2_dfrbp_1 \i_coord.l_xl.state[6]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_16_clk),
    .RESET_B(net382),
    .D(_00074_),
    .Q_N(_07641_),
    .Q(\i_coord.l_xl.data_out[6] ));
 sg13g2_dfrbp_1 \i_coord.l_xl.state[7]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_14_clk),
    .RESET_B(net383),
    .D(_00075_),
    .Q_N(_07640_),
    .Q(\i_coord.l_xl.data_out[7] ));
 sg13g2_dfrbp_1 \i_coord.l_xl.state[8]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_17_clk),
    .RESET_B(net384),
    .D(_00076_),
    .Q_N(_07639_),
    .Q(\i_coord.l_xl.data_out[8] ));
 sg13g2_dfrbp_1 \i_coord.l_xl.state[9]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_14_clk),
    .RESET_B(net385),
    .D(_00077_),
    .Q_N(_07638_),
    .Q(\i_coord.l_xl.data_out[9] ));
 sg13g2_dfrbp_1 \i_coord.l_yip.state[0]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_15_clk),
    .RESET_B(net386),
    .D(_00078_),
    .Q_N(_07637_),
    .Q(\i_coord.l_yip.data_out[0] ));
 sg13g2_dfrbp_1 \i_coord.l_yip.state[1]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_11_clk),
    .RESET_B(net387),
    .D(_00079_),
    .Q_N(_07636_),
    .Q(\i_coord.l_yip.data_out[1] ));
 sg13g2_dfrbp_1 \i_coord.l_yip.state[2]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_15_clk),
    .RESET_B(net388),
    .D(_00080_),
    .Q_N(_07635_),
    .Q(\i_coord.l_yip.data_out[2] ));
 sg13g2_dfrbp_1 \i_coord.l_yip.state[3]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_15_clk),
    .RESET_B(net389),
    .D(_00081_),
    .Q_N(_07634_),
    .Q(\i_coord.l_yip.data_out[3] ));
 sg13g2_dfrbp_1 \i_coord.l_yip.state[4]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_14_clk),
    .RESET_B(net390),
    .D(_00082_),
    .Q_N(_07633_),
    .Q(\i_coord.l_yip.data_out[4] ));
 sg13g2_dfrbp_1 \i_coord.l_yip.state[5]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_15_clk),
    .RESET_B(net391),
    .D(_00083_),
    .Q_N(_07632_),
    .Q(\i_coord.l_yip.data_out[5] ));
 sg13g2_dfrbp_1 \i_coord.l_yip.state[6]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_9_clk),
    .RESET_B(net392),
    .D(_00084_),
    .Q_N(_07631_),
    .Q(\i_coord.l_yip.data_out[6] ));
 sg13g2_dfrbp_1 \i_coord.l_yip.state[7]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_9_clk),
    .RESET_B(net393),
    .D(_00085_),
    .Q_N(_07630_),
    .Q(\i_coord.l_yip.data_out[7] ));
 sg13g2_dfrbp_1 \i_coord.l_yip.state[8]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_9_clk),
    .RESET_B(net394),
    .D(_00086_),
    .Q_N(_07629_),
    .Q(\i_coord.l_yip.data_out[8] ));
 sg13g2_dfrbp_1 \i_coord.l_yip.state[9]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_9_clk),
    .RESET_B(net395),
    .D(_00087_),
    .Q_N(_07628_),
    .Q(\i_coord.l_yip.data_out[9] ));
 sg13g2_dfrbp_1 \i_coord.l_yt.state[0]$_SDFFCE_PP0P_  (.CLK(clknet_leaf_12_clk),
    .RESET_B(net396),
    .D(_00088_),
    .Q_N(_07627_),
    .Q(\i_coord.l_yt.data_out[0] ));
 sg13g2_dfrbp_1 \i_coord.l_yt.state[10]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_6_clk),
    .RESET_B(net397),
    .D(_00089_),
    .Q_N(_07626_),
    .Q(\i_coord.l_yt.data_out[10] ));
 sg13g2_dfrbp_1 \i_coord.l_yt.state[11]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_6_clk),
    .RESET_B(net398),
    .D(_00090_),
    .Q_N(_07625_),
    .Q(\i_coord.l_yt.data_out[11] ));
 sg13g2_dfrbp_1 \i_coord.l_yt.state[12]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_6_clk),
    .RESET_B(net399),
    .D(_00091_),
    .Q_N(_07624_),
    .Q(\i_coord.l_yt.data_out[12] ));
 sg13g2_dfrbp_1 \i_coord.l_yt.state[13]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_6_clk),
    .RESET_B(net400),
    .D(_00092_),
    .Q_N(_07623_),
    .Q(\i_coord.l_yt.data_out[13] ));
 sg13g2_dfrbp_1 \i_coord.l_yt.state[14]$_SDFFCE_PN1P_  (.CLK(clknet_leaf_7_clk),
    .RESET_B(net401),
    .D(_00093_),
    .Q_N(_07622_),
    .Q(\i_coord.l_yt.data_out[14] ));
 sg13g2_dfrbp_1 \i_coord.l_yt.state[1]$_SDFFCE_PP0P_  (.CLK(clknet_leaf_12_clk),
    .RESET_B(net402),
    .D(_00094_),
    .Q_N(_07621_),
    .Q(\i_coord.l_yt.data_out[1] ));
 sg13g2_dfrbp_1 \i_coord.l_yt.state[2]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_9_clk),
    .RESET_B(net403),
    .D(_00095_),
    .Q_N(_07620_),
    .Q(\i_coord.l_yt.data_out[2] ));
 sg13g2_dfrbp_1 \i_coord.l_yt.state[3]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_8_clk),
    .RESET_B(net404),
    .D(_00096_),
    .Q_N(_07619_),
    .Q(\i_coord.l_yt.data_out[3] ));
 sg13g2_dfrbp_1 \i_coord.l_yt.state[4]$_SDFFCE_PN1P_  (.CLK(clknet_leaf_7_clk),
    .RESET_B(net405),
    .D(_00097_),
    .Q_N(_07618_),
    .Q(\i_coord.l_yt.data_out[4] ));
 sg13g2_dfrbp_1 \i_coord.l_yt.state[5]$_SDFFCE_PN1P_  (.CLK(clknet_leaf_7_clk),
    .RESET_B(net406),
    .D(_00098_),
    .Q_N(_07617_),
    .Q(\i_coord.l_yt.data_out[5] ));
 sg13g2_dfrbp_1 \i_coord.l_yt.state[6]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_9_clk),
    .RESET_B(net407),
    .D(_00099_),
    .Q_N(_07616_),
    .Q(\i_coord.l_yt.data_out[6] ));
 sg13g2_dfrbp_1 \i_coord.l_yt.state[7]$_SDFFCE_PN1P_  (.CLK(clknet_leaf_7_clk),
    .RESET_B(net408),
    .D(_00100_),
    .Q_N(_07615_),
    .Q(\i_coord.l_yt.data_out[7] ));
 sg13g2_dfrbp_1 \i_coord.l_yt.state[8]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_6_clk),
    .RESET_B(net409),
    .D(_00101_),
    .Q_N(_07614_),
    .Q(\i_coord.l_yt.data_out[8] ));
 sg13g2_dfrbp_1 \i_coord.l_yt.state[9]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_5_clk),
    .RESET_B(net410),
    .D(_00102_),
    .Q_N(_07613_),
    .Q(\i_coord.l_yt.data_out[9] ));
 sg13g2_dfrbp_1 \i_coord.x_row_start[0]$_SDFFCE_PP0P_  (.CLK(clknet_leaf_19_clk),
    .RESET_B(net411),
    .D(_00103_),
    .Q_N(_07612_),
    .Q(\i_coord.x_row_start[-13] ));
 sg13g2_dfrbp_1 \i_coord.x_row_start[10]$_DFFE_PP_  (.CLK(clknet_leaf_18_clk),
    .RESET_B(net412),
    .D(_00104_),
    .Q_N(_07611_),
    .Q(\i_coord.x_row_start[-3] ));
 sg13g2_dfrbp_1 \i_coord.x_row_start[11]$_DFFE_PP_  (.CLK(clknet_leaf_18_clk),
    .RESET_B(net413),
    .D(_00105_),
    .Q_N(_07610_),
    .Q(\i_coord.x_row_start[-2] ));
 sg13g2_dfrbp_1 \i_coord.x_row_start[12]$_DFFE_PP_  (.CLK(clknet_leaf_18_clk),
    .RESET_B(net414),
    .D(_00106_),
    .Q_N(_07609_),
    .Q(\i_coord.x_row_start[-1] ));
 sg13g2_dfrbp_1 \i_coord.x_row_start[13]$_DFFE_PP_  (.CLK(clknet_leaf_20_clk),
    .RESET_B(net415),
    .D(_00107_),
    .Q_N(_07608_),
    .Q(\i_coord.x_row_start[0] ));
 sg13g2_dfrbp_1 \i_coord.x_row_start[14]$_DFFE_PP_  (.CLK(clknet_leaf_20_clk),
    .RESET_B(net416),
    .D(_00108_),
    .Q_N(_07607_),
    .Q(\i_coord.x_row_start[1] ));
 sg13g2_dfrbp_1 \i_coord.x_row_start[15]$_DFFE_PP_  (.CLK(clknet_leaf_16_clk),
    .RESET_B(net417),
    .D(_00109_),
    .Q_N(_07606_),
    .Q(\i_coord.x_row_start[2] ));
 sg13g2_dfrbp_1 \i_coord.x_row_start[1]$_SDFFCE_PP0P_  (.CLK(clknet_leaf_19_clk),
    .RESET_B(net418),
    .D(_00110_),
    .Q_N(_07605_),
    .Q(\i_coord.x_row_start[-12] ));
 sg13g2_dfrbp_1 \i_coord.x_row_start[2]$_SDFFCE_PP0P_  (.CLK(clknet_leaf_19_clk),
    .RESET_B(net419),
    .D(_00111_),
    .Q_N(_07604_),
    .Q(\i_coord.x_row_start[-11] ));
 sg13g2_dfrbp_1 \i_coord.x_row_start[3]$_DFFE_PP_  (.CLK(clknet_leaf_18_clk),
    .RESET_B(net420),
    .D(_00112_),
    .Q_N(_07603_),
    .Q(\i_coord.x_row_start[-10] ));
 sg13g2_dfrbp_1 \i_coord.x_row_start[4]$_DFFE_PP_  (.CLK(clknet_leaf_17_clk),
    .RESET_B(net421),
    .D(_00113_),
    .Q_N(_07602_),
    .Q(\i_coord.x_row_start[-9] ));
 sg13g2_dfrbp_1 \i_coord.x_row_start[5]$_DFFE_PP_  (.CLK(clknet_leaf_17_clk),
    .RESET_B(net422),
    .D(_00114_),
    .Q_N(_07601_),
    .Q(\i_coord.x_row_start[-8] ));
 sg13g2_dfrbp_1 \i_coord.x_row_start[6]$_DFFE_PP_  (.CLK(clknet_leaf_17_clk),
    .RESET_B(net423),
    .D(_00115_),
    .Q_N(_07600_),
    .Q(\i_coord.x_row_start[-7] ));
 sg13g2_dfrbp_1 \i_coord.x_row_start[7]$_DFFE_PP_  (.CLK(clknet_leaf_17_clk),
    .RESET_B(net424),
    .D(_00116_),
    .Q_N(_07599_),
    .Q(\i_coord.x_row_start[-6] ));
 sg13g2_dfrbp_1 \i_coord.x_row_start[8]$_DFFE_PP_  (.CLK(clknet_leaf_18_clk),
    .RESET_B(net425),
    .D(_00117_),
    .Q_N(_07598_),
    .Q(\i_coord.x_row_start[-5] ));
 sg13g2_dfrbp_1 \i_coord.x_row_start[9]$_DFFE_PP_  (.CLK(clknet_leaf_18_clk),
    .RESET_B(net426),
    .D(_00118_),
    .Q_N(_07597_),
    .Q(\i_coord.x_row_start[-4] ));
 sg13g2_dfrbp_1 \i_coord.y_inc_row[0]$_SDFFE_PN1P_  (.CLK(clknet_leaf_13_clk),
    .RESET_B(net427),
    .D(_00119_),
    .Q_N(_07596_),
    .Q(\i_coord.y_inc_row[-13] ));
 sg13g2_dfrbp_1 \i_coord.y_inc_row[1]$_SDFFE_PN1P_  (.CLK(clknet_leaf_13_clk),
    .RESET_B(net428),
    .D(_00120_),
    .Q_N(_07595_),
    .Q(\i_coord.y_inc_row[-12] ));
 sg13g2_dfrbp_1 \i_coord.y_inc_row[2]$_SDFFE_PN0P_  (.CLK(clknet_leaf_12_clk),
    .RESET_B(net429),
    .D(_00121_),
    .Q_N(_07594_),
    .Q(\i_coord.y_inc_row[-11] ));
 sg13g2_dfrbp_1 \i_coord.y_inc_row[3]$_SDFFE_PN1P_  (.CLK(clknet_leaf_8_clk),
    .RESET_B(net430),
    .D(_00122_),
    .Q_N(_07593_),
    .Q(\i_coord.y_inc_row[-10] ));
 sg13g2_dfrbp_1 \i_coord.y_inc_row[4]$_SDFFE_PN1P_  (.CLK(clknet_leaf_8_clk),
    .RESET_B(net431),
    .D(_00123_),
    .Q_N(_07592_),
    .Q(\i_coord.y_inc_row[-9] ));
 sg13g2_dfrbp_1 \i_coord.y_inc_row[5]$_SDFFE_PN1P_  (.CLK(clknet_leaf_7_clk),
    .RESET_B(net432),
    .D(_00124_),
    .Q_N(_07591_),
    .Q(\i_coord.y_inc_row[-8] ));
 sg13g2_dfrbp_1 \i_coord.y_inc_row[6]$_SDFFE_PN0P_  (.CLK(clknet_leaf_8_clk),
    .RESET_B(net433),
    .D(_00125_),
    .Q_N(_07590_),
    .Q(\i_coord.y_inc_row[-7] ));
 sg13g2_dfrbp_1 \i_coord.y_inc_row[7]$_SDFFE_PN1P_  (.CLK(clknet_leaf_5_clk),
    .RESET_B(net434),
    .D(_00126_),
    .Q_N(_07589_),
    .Q(\i_coord.y_inc_row[-6] ));
 sg13g2_dfrbp_1 \i_coord.y_row_start[0]$_DFFE_PP_  (.CLK(clknet_leaf_9_clk),
    .RESET_B(net435),
    .D(_00127_),
    .Q_N(_07588_),
    .Q(\i_coord.y_row_start[-13] ));
 sg13g2_dfrbp_1 \i_coord.y_row_start[10]$_DFFE_PP_  (.CLK(clknet_leaf_2_clk),
    .RESET_B(net436),
    .D(_00128_),
    .Q_N(_07587_),
    .Q(\i_coord.y_row_start[-3] ));
 sg13g2_dfrbp_1 \i_coord.y_row_start[11]$_DFFE_PP_  (.CLK(clknet_leaf_2_clk),
    .RESET_B(net437),
    .D(_00129_),
    .Q_N(_07586_),
    .Q(\i_coord.y_row_start[-2] ));
 sg13g2_dfrbp_1 \i_coord.y_row_start[12]$_DFFE_PP_  (.CLK(clknet_leaf_6_clk),
    .RESET_B(net438),
    .D(_00130_),
    .Q_N(_07585_),
    .Q(\i_coord.y_row_start[-1] ));
 sg13g2_dfrbp_1 \i_coord.y_row_start[13]$_DFFE_PP_  (.CLK(clknet_leaf_6_clk),
    .RESET_B(net439),
    .D(_00131_),
    .Q_N(_07584_),
    .Q(\i_coord.y_row_start[0] ));
 sg13g2_dfrbp_1 \i_coord.y_row_start[14]$_DFFE_PP_  (.CLK(clknet_leaf_7_clk),
    .RESET_B(net440),
    .D(_00132_),
    .Q_N(_07583_),
    .Q(\i_coord.y_row_start[1] ));
 sg13g2_dfrbp_1 \i_coord.y_row_start[1]$_DFFE_PP_  (.CLK(clknet_leaf_12_clk),
    .RESET_B(net441),
    .D(_00133_),
    .Q_N(_07582_),
    .Q(\i_coord.y_row_start[-12] ));
 sg13g2_dfrbp_1 \i_coord.y_row_start[2]$_DFFE_PP_  (.CLK(clknet_leaf_8_clk),
    .RESET_B(net442),
    .D(_00134_),
    .Q_N(_07581_),
    .Q(\i_coord.y_row_start[-11] ));
 sg13g2_dfrbp_1 \i_coord.y_row_start[3]$_DFFE_PP_  (.CLK(clknet_leaf_8_clk),
    .RESET_B(net443),
    .D(_00135_),
    .Q_N(_07580_),
    .Q(\i_coord.y_row_start[-10] ));
 sg13g2_dfrbp_1 \i_coord.y_row_start[4]$_DFFE_PP_  (.CLK(clknet_leaf_8_clk),
    .RESET_B(net444),
    .D(_00136_),
    .Q_N(_07579_),
    .Q(\i_coord.y_row_start[-9] ));
 sg13g2_dfrbp_1 \i_coord.y_row_start[5]$_DFFE_PP_  (.CLK(clknet_leaf_7_clk),
    .RESET_B(net445),
    .D(_00137_),
    .Q_N(_07578_),
    .Q(\i_coord.y_row_start[-8] ));
 sg13g2_dfrbp_1 \i_coord.y_row_start[6]$_DFFE_PP_  (.CLK(clknet_leaf_8_clk),
    .RESET_B(net446),
    .D(_00138_),
    .Q_N(_07577_),
    .Q(\i_coord.y_row_start[-7] ));
 sg13g2_dfrbp_1 \i_coord.y_row_start[7]$_DFFE_PP_  (.CLK(clknet_leaf_5_clk),
    .RESET_B(net447),
    .D(_00139_),
    .Q_N(_07576_),
    .Q(\i_coord.y_row_start[-6] ));
 sg13g2_dfrbp_1 \i_coord.y_row_start[8]$_DFFE_PP_  (.CLK(clknet_leaf_5_clk),
    .RESET_B(net448),
    .D(_00140_),
    .Q_N(_07575_),
    .Q(\i_coord.y_row_start[-5] ));
 sg13g2_dfrbp_1 \i_coord.y_row_start[9]$_DFFE_PP_  (.CLK(clknet_leaf_5_clk),
    .RESET_B(net449),
    .D(_00141_),
    .Q_N(_07574_),
    .Q(\i_coord.y_row_start[-4] ));
 sg13g2_dfrbp_1 \i_vga.timing_hor.counter[0]$_SDFFE_PN0P_  (.CLK(clknet_leaf_0_clk),
    .RESET_B(net450),
    .D(_00142_),
    .Q_N(_00026_),
    .Q(\i_vga.timing_hor.counter[0] ));
 sg13g2_dfrbp_1 \i_vga.timing_hor.counter[10]$_SDFFE_PN1P_  (.CLK(clknet_leaf_3_clk),
    .RESET_B(net451),
    .D(_00143_),
    .Q_N(_00033_),
    .Q(\i_vga.timing_hor.counter[10] ));
 sg13g2_dfrbp_1 \i_vga.timing_hor.counter[1]$_SDFFE_PN0P_  (.CLK(clknet_leaf_2_clk),
    .RESET_B(net452),
    .D(_00144_),
    .Q_N(_07573_),
    .Q(\i_vga.timing_hor.counter[1] ));
 sg13g2_dfrbp_1 \i_vga.timing_hor.counter[2]$_SDFFE_PN0P_  (.CLK(clknet_leaf_0_clk),
    .RESET_B(net453),
    .D(_00145_),
    .Q_N(_07572_),
    .Q(\i_vga.timing_hor.counter[2] ));
 sg13g2_dfrbp_1 \i_vga.timing_hor.counter[3]$_SDFFE_PN0P_  (.CLK(clknet_leaf_2_clk),
    .RESET_B(net454),
    .D(_00146_),
    .Q_N(_00027_),
    .Q(\i_vga.timing_hor.counter[3] ));
 sg13g2_dfrbp_1 \i_vga.timing_hor.counter[4]$_SDFFE_PN1P_  (.CLK(clknet_leaf_3_clk),
    .RESET_B(net455),
    .D(_00147_),
    .Q_N(_07571_),
    .Q(\i_vga.timing_hor.counter[4] ));
 sg13g2_dfrbp_1 \i_vga.timing_hor.counter[5]$_SDFFE_PN0P_  (.CLK(clknet_leaf_2_clk),
    .RESET_B(net456),
    .D(_00148_),
    .Q_N(_07570_),
    .Q(\i_vga.timing_hor.counter[5] ));
 sg13g2_dfrbp_1 \i_vga.timing_hor.counter[6]$_SDFFE_PN1P_  (.CLK(clknet_leaf_3_clk),
    .RESET_B(net457),
    .D(_00149_),
    .Q_N(_07569_),
    .Q(\i_vga.timing_hor.counter[6] ));
 sg13g2_dfrbp_1 \i_vga.timing_hor.counter[7]$_SDFFE_PN0P_  (.CLK(clknet_leaf_3_clk),
    .RESET_B(net458),
    .D(_00150_),
    .Q_N(_00028_),
    .Q(\i_vga.timing_hor.counter[7] ));
 sg13g2_dfrbp_1 \i_vga.timing_hor.counter[8]$_SDFFE_PN1P_  (.CLK(clknet_leaf_3_clk),
    .RESET_B(net459),
    .D(_00151_),
    .Q_N(_07568_),
    .Q(\i_vga.timing_hor.counter[8] ));
 sg13g2_dfrbp_1 \i_vga.timing_hor.counter[9]$_SDFFE_PN1P_  (.CLK(clknet_leaf_3_clk),
    .RESET_B(net460),
    .D(_00152_),
    .Q_N(_07669_),
    .Q(\i_vga.timing_hor.counter[9] ));
 sg13g2_dfrbp_1 \i_vga.timing_hor.sync$_DFF_P_  (.CLK(clknet_leaf_5_clk),
    .RESET_B(net461),
    .D(_00002_),
    .Q_N(_07567_),
    .Q(\i_vga.hsync ));
 sg13g2_dfrbp_1 \i_vga.timing_ver.counter[0]$_SDFFE_PN1P_  (.CLK(clknet_leaf_3_clk),
    .RESET_B(net462),
    .D(_00153_),
    .Q_N(_00017_),
    .Q(\i_vga.timing_ver.counter[0] ));
 sg13g2_dfrbp_1 \i_vga.timing_ver.counter[1]$_SDFFE_PN0P_  (.CLK(clknet_leaf_4_clk),
    .RESET_B(net463),
    .D(_00154_),
    .Q_N(_07566_),
    .Q(\i_vga.timing_ver.counter[1] ));
 sg13g2_dfrbp_1 \i_vga.timing_ver.counter[2]$_SDFFE_PN1P_  (.CLK(clknet_leaf_4_clk),
    .RESET_B(net464),
    .D(_00155_),
    .Q_N(_07565_),
    .Q(\i_vga.timing_ver.counter[2] ));
 sg13g2_dfrbp_1 \i_vga.timing_ver.counter[3]$_SDFFE_PN1P_  (.CLK(clknet_leaf_3_clk),
    .RESET_B(net465),
    .D(_00156_),
    .Q_N(_07564_),
    .Q(\i_vga.timing_ver.counter[3] ));
 sg13g2_dfrbp_1 \i_vga.timing_ver.counter[4]$_SDFFE_PN0P_  (.CLK(clknet_leaf_4_clk),
    .RESET_B(net466),
    .D(_00157_),
    .Q_N(_07563_),
    .Q(\i_vga.timing_ver.counter[4] ));
 sg13g2_dfrbp_1 \i_vga.timing_ver.counter[5]$_SDFFE_PN1P_  (.CLK(clknet_leaf_4_clk),
    .RESET_B(net467),
    .D(_00158_),
    .Q_N(_07562_),
    .Q(\i_vga.timing_ver.counter[5] ));
 sg13g2_dfrbp_1 \i_vga.timing_ver.counter[6]$_SDFFE_PN1P_  (.CLK(clknet_leaf_4_clk),
    .RESET_B(net468),
    .D(_00159_),
    .Q_N(_07561_),
    .Q(\i_vga.timing_ver.counter[6] ));
 sg13g2_dfrbp_1 \i_vga.timing_ver.counter[7]$_SDFFE_PN1P_  (.CLK(clknet_leaf_4_clk),
    .RESET_B(net469),
    .D(_00160_),
    .Q_N(_07560_),
    .Q(\i_vga.timing_ver.counter[7] ));
 sg13g2_dfrbp_1 \i_vga.timing_ver.counter[8]$_SDFFE_PN1P_  (.CLK(clknet_leaf_4_clk),
    .RESET_B(net470),
    .D(_00161_),
    .Q_N(_07559_),
    .Q(\i_vga.timing_ver.counter[8] ));
 sg13g2_dfrbp_1 \i_vga.timing_ver.counter[9]$_SDFFE_PN1P_  (.CLK(clknet_leaf_4_clk),
    .RESET_B(net471),
    .D(_00162_),
    .Q_N(_00016_),
    .Q(\i_vga.timing_ver.counter[9] ));
 sg13g2_dfrbp_1 \i_vga.timing_ver.sync$_DFF_P_  (.CLK(clknet_leaf_5_clk),
    .RESET_B(net472),
    .D(\i_vga.timing_ver.sync_tmp ),
    .Q_N(_07670_),
    .Q(\i_vga.timing_ver.sync ));
 sg13g2_dfrbp_1 \i_vga.vblank$_DFF_P_  (.CLK(clknet_leaf_5_clk),
    .RESET_B(net473),
    .D(\i_vga.timing_ver.blank ),
    .Q_N(_07558_),
    .Q(\i_vga.vblank ));
 sg13g2_dfrbp_1 \iter[0]$_SDFFCE_PP0N_  (.CLK(clknet_leaf_25_clk),
    .RESET_B(net474),
    .D(_00163_),
    .Q_N(_07557_),
    .Q(\iter[0] ));
 sg13g2_dfrbp_1 \iter[1]$_SDFFCE_PP0N_  (.CLK(clknet_leaf_10_clk),
    .RESET_B(net475),
    .D(_00164_),
    .Q_N(_07556_),
    .Q(\iter[1] ));
 sg13g2_dfrbp_1 \iter[2]$_SDFFCE_PP0N_  (.CLK(clknet_leaf_0_clk),
    .RESET_B(net476),
    .D(_00165_),
    .Q_N(_07555_),
    .Q(\iter[2] ));
 sg13g2_dfrbp_1 \iter[3]$_SDFFCE_PP0N_  (.CLK(clknet_leaf_1_clk),
    .RESET_B(net477),
    .D(_00166_),
    .Q_N(_07554_),
    .Q(\iter[3] ));
 sg13g2_dfrbp_1 \last_iter[0]$_DFFE_PP_  (.CLK(clknet_leaf_0_clk),
    .RESET_B(net478),
    .D(_00030_),
    .Q_N(_07553_),
    .Q(\last_iter[0] ));
 sg13g2_dfrbp_1 \last_iter[1]$_DFFE_PP_  (.CLK(clknet_leaf_1_clk),
    .RESET_B(net479),
    .D(_00029_),
    .Q_N(_07552_),
    .Q(\last_iter[1] ));
 sg13g2_dfrbp_1 \last_iter[2]$_DFFE_PP_  (.CLK(clknet_leaf_1_clk),
    .RESET_B(net480),
    .D(_00031_),
    .Q_N(_00032_),
    .Q(\last_iter[2] ));
 sg13g2_dfrbp_1 \last_iter[3]$_DFFE_PP_  (.CLK(clknet_leaf_0_clk),
    .RESET_B(net481),
    .D(_00015_),
    .Q_N(_07551_),
    .Q(\last_iter[3] ));
 sg13g2_dfrbp_1 \last_iter[4]$_DFFE_PP_  (.CLK(clknet_leaf_1_clk),
    .RESET_B(net482),
    .D(_00000_),
    .Q_N(_07550_),
    .Q(\last_iter[4] ));
 sg13g2_dfrbp_1 \step[0]$_SDFF_PP0_  (.CLK(clknet_leaf_1_clk),
    .RESET_B(net483),
    .D(_00167_),
    .Q_N(_00044_),
    .Q(\step[0] ));
 sg13g2_dfrbp_1 \step[1]$_SDFF_PP0_  (.CLK(clknet_leaf_0_clk),
    .RESET_B(net484),
    .D(_00168_),
    .Q_N(_07549_),
    .Q(\step[1] ));
 sg13g2_dfrbp_1 \step[2]$_SDFF_PP0_  (.CLK(clknet_leaf_0_clk),
    .RESET_B(net485),
    .D(_00169_),
    .Q_N(_07548_),
    .Q(\step[2] ));
 sg13g2_dfrbp_1 \step[3]$_SDFF_PP0_  (.CLK(clknet_leaf_0_clk),
    .RESET_B(net486),
    .D(_00170_),
    .Q_N(_07547_),
    .Q(\step[3] ));
 sg13g2_dfrbp_1 \video_colour[0]$_SDFF_PP0_  (.CLK(clknet_leaf_2_clk),
    .RESET_B(net487),
    .D(_00171_),
    .Q_N(_07546_),
    .Q(\video_colour[0] ));
 sg13g2_dfrbp_1 \video_colour[1]$_SDFF_PP0_  (.CLK(clknet_leaf_2_clk),
    .RESET_B(net488),
    .D(_00172_),
    .Q_N(_07545_),
    .Q(\video_colour[1] ));
 sg13g2_dfrbp_1 \video_colour[2]$_SDFF_PP0_  (.CLK(clknet_leaf_2_clk),
    .RESET_B(net489),
    .D(_00173_),
    .Q_N(_07544_),
    .Q(\video_colour[2] ));
 sg13g2_dfrbp_1 \video_colour[3]$_SDFF_PP0_  (.CLK(clknet_leaf_1_clk),
    .RESET_B(net490),
    .D(_00174_),
    .Q_N(_07543_),
    .Q(\video_colour[3] ));
 sg13g2_dfrbp_1 \video_colour[4]$_SDFF_PP0_  (.CLK(clknet_leaf_1_clk),
    .RESET_B(net491),
    .D(_00175_),
    .Q_N(_07542_),
    .Q(\video_colour[4] ));
 sg13g2_dfrbp_1 \video_colour[5]$_SDFF_PP0_  (.CLK(clknet_leaf_1_clk),
    .RESET_B(net492),
    .D(_00176_),
    .Q_N(_07541_),
    .Q(\video_colour[5] ));
 sg13g2_dfrbp_1 \x0[0]$_DFFE_PP_  (.CLK(clknet_leaf_19_clk),
    .RESET_B(net493),
    .D(_00177_),
    .Q_N(_07540_),
    .Q(\i_coord.x0[-13] ));
 sg13g2_dfrbp_1 \x0[10]$_DFFE_PP_  (.CLK(clknet_leaf_11_clk),
    .RESET_B(net494),
    .D(_00178_),
    .Q_N(_07539_),
    .Q(\i_coord.x0[-3] ));
 sg13g2_dfrbp_1 \x0[11]$_DFFE_PP_  (.CLK(clknet_leaf_11_clk),
    .RESET_B(net495),
    .D(_00179_),
    .Q_N(_07538_),
    .Q(\i_coord.x0[-2] ));
 sg13g2_dfrbp_1 \x0[12]$_DFFE_PP_  (.CLK(clknet_leaf_11_clk),
    .RESET_B(net496),
    .D(_00180_),
    .Q_N(_07537_),
    .Q(\i_coord.x0[-1] ));
 sg13g2_dfrbp_1 \x0[13]$_DFFE_PP_  (.CLK(clknet_leaf_11_clk),
    .RESET_B(net497),
    .D(_00181_),
    .Q_N(_07536_),
    .Q(\i_coord.x0[0] ));
 sg13g2_dfrbp_1 \x0[14]$_DFFE_PP_  (.CLK(clknet_leaf_11_clk),
    .RESET_B(net498),
    .D(_00182_),
    .Q_N(_07535_),
    .Q(\i_coord.x0[1] ));
 sg13g2_dfrbp_1 \x0[15]$_DFFE_PP_  (.CLK(clknet_leaf_10_clk),
    .RESET_B(net499),
    .D(_00183_),
    .Q_N(_07534_),
    .Q(\i_coord.x0[2] ));
 sg13g2_dfrbp_1 \x0[1]$_DFFE_PP_  (.CLK(clknet_leaf_20_clk),
    .RESET_B(net500),
    .D(_00184_),
    .Q_N(_07533_),
    .Q(\i_coord.x0[-12] ));
 sg13g2_dfrbp_1 \x0[2]$_DFFE_PP_  (.CLK(clknet_leaf_19_clk),
    .RESET_B(net501),
    .D(_00185_),
    .Q_N(_07532_),
    .Q(\i_coord.x0[-11] ));
 sg13g2_dfrbp_1 \x0[3]$_DFFE_PP_  (.CLK(clknet_leaf_15_clk),
    .RESET_B(net502),
    .D(_00186_),
    .Q_N(_07531_),
    .Q(\i_coord.x0[-10] ));
 sg13g2_dfrbp_1 \x0[4]$_DFFE_PP_  (.CLK(clknet_leaf_15_clk),
    .RESET_B(net503),
    .D(_00187_),
    .Q_N(_07530_),
    .Q(\i_coord.x0[-9] ));
 sg13g2_dfrbp_1 \x0[5]$_DFFE_PP_  (.CLK(clknet_leaf_15_clk),
    .RESET_B(net504),
    .D(_00188_),
    .Q_N(_07529_),
    .Q(\i_coord.x0[-8] ));
 sg13g2_dfrbp_1 \x0[6]$_DFFE_PP_  (.CLK(clknet_leaf_20_clk),
    .RESET_B(net505),
    .D(_00189_),
    .Q_N(_07528_),
    .Q(\i_coord.x0[-7] ));
 sg13g2_dfrbp_1 \x0[7]$_DFFE_PP_  (.CLK(clknet_leaf_20_clk),
    .RESET_B(net506),
    .D(_00190_),
    .Q_N(_07527_),
    .Q(\i_coord.x0[-6] ));
 sg13g2_dfrbp_1 \x0[8]$_DFFE_PP_  (.CLK(clknet_leaf_20_clk),
    .RESET_B(net507),
    .D(_00191_),
    .Q_N(_07526_),
    .Q(\i_coord.x0[-5] ));
 sg13g2_dfrbp_1 \x0[9]$_DFFE_PP_  (.CLK(clknet_leaf_20_clk),
    .RESET_B(net508),
    .D(_00192_),
    .Q_N(_07525_),
    .Q(\i_coord.x0[-4] ));
 sg13g2_dfrbp_1 \x[0]$_DFFE_PP_  (.CLK(clknet_leaf_22_clk),
    .RESET_B(net509),
    .D(_00193_),
    .Q_N(_00034_),
    .Q(\i_mandel.i_sq_x.x[-13] ));
 sg13g2_dfrbp_1 \x[10]$_DFFE_PP_  (.CLK(clknet_leaf_24_clk),
    .RESET_B(net510),
    .D(_00194_),
    .Q_N(_00010_),
    .Q(\i_mandel.i_sq_x.x[-3] ));
 sg13g2_dfrbp_1 \x[11]$_DFFE_PP_  (.CLK(clknet_leaf_24_clk),
    .RESET_B(net511),
    .D(_00195_),
    .Q_N(_00009_),
    .Q(\i_mandel.i_sq_x.x[-2] ));
 sg13g2_dfrbp_1 \x[12]$_DFFE_PP_  (.CLK(clknet_leaf_22_clk),
    .RESET_B(net512),
    .D(_00196_),
    .Q_N(_00008_),
    .Q(\i_mandel.i_sq_x.x[-1] ));
 sg13g2_dfrbp_1 \x[13]$_DFFE_PP_  (.CLK(clknet_leaf_24_clk),
    .RESET_B(net513),
    .D(_00197_),
    .Q_N(_00007_),
    .Q(\i_mandel.i_sq_x.x[0] ));
 sg13g2_dfrbp_1 \x[14]$_DFFE_PP_  (.CLK(clknet_leaf_22_clk),
    .RESET_B(net514),
    .D(_00198_),
    .Q_N(_00005_),
    .Q(\i_mandel.i_sq_x.x[1] ));
 sg13g2_dfrbp_1 \x[15]$_DFFE_PP_  (.CLK(clknet_leaf_24_clk),
    .RESET_B(net515),
    .D(_00199_),
    .Q_N(_00004_),
    .Q(\i_mandel.i_sq_x.x[2] ));
 sg13g2_dfrbp_1 \x[1]$_DFFE_PP_  (.CLK(clknet_leaf_22_clk),
    .RESET_B(net516),
    .D(_00200_),
    .Q_N(_07524_),
    .Q(\i_mandel.i_sq_x.x[-12] ));
 sg13g2_dfrbp_1 \x[2]$_DFFE_PP_  (.CLK(clknet_leaf_22_clk),
    .RESET_B(net517),
    .D(_00201_),
    .Q_N(_07523_),
    .Q(\i_mandel.i_sq_x.x[-11] ));
 sg13g2_dfrbp_1 \x[3]$_DFFE_PP_  (.CLK(clknet_leaf_22_clk),
    .RESET_B(net518),
    .D(_00202_),
    .Q_N(_00006_),
    .Q(\i_mandel.i_sq_x.x[-10] ));
 sg13g2_dfrbp_1 \x[4]$_DFFE_PP_  (.CLK(clknet_leaf_23_clk),
    .RESET_B(net519),
    .D(_00203_),
    .Q_N(_07522_),
    .Q(\i_mandel.i_sq_x.x[-9] ));
 sg13g2_dfrbp_1 \x[5]$_DFFE_PP_  (.CLK(clknet_leaf_24_clk),
    .RESET_B(net520),
    .D(_00204_),
    .Q_N(_00013_),
    .Q(\i_mandel.i_sq_x.x[-8] ));
 sg13g2_dfrbp_1 \x[6]$_DFFE_PP_  (.CLK(clknet_leaf_24_clk),
    .RESET_B(net521),
    .D(_00205_),
    .Q_N(_07521_),
    .Q(\i_mandel.i_sq_x.x[-7] ));
 sg13g2_dfrbp_1 \x[7]$_DFFE_PP_  (.CLK(clknet_leaf_23_clk),
    .RESET_B(net522),
    .D(_00206_),
    .Q_N(_07520_),
    .Q(\i_mandel.i_sq_x.x[-6] ));
 sg13g2_dfrbp_1 \x[8]$_DFFE_PP_  (.CLK(clknet_leaf_24_clk),
    .RESET_B(net523),
    .D(_00207_),
    .Q_N(_00012_),
    .Q(\i_mandel.i_sq_x.x[-5] ));
 sg13g2_dfrbp_1 \x[9]$_DFFE_PP_  (.CLK(clknet_leaf_24_clk),
    .RESET_B(net524),
    .D(_00208_),
    .Q_N(_00011_),
    .Q(\i_mandel.i_sq_x.x[-4] ));
 sg13g2_dfrbp_1 \y0[0]$_DFFE_PP_  (.CLK(clknet_leaf_11_clk),
    .RESET_B(net525),
    .D(_00209_),
    .Q_N(_07519_),
    .Q(\i_coord.y0[-13] ));
 sg13g2_dfrbp_1 \y0[10]$_DFFE_PP_  (.CLK(clknet_leaf_10_clk),
    .RESET_B(net526),
    .D(_00210_),
    .Q_N(_00022_),
    .Q(\i_coord.y0[-3] ));
 sg13g2_dfrbp_1 \y0[11]$_DFFE_PP_  (.CLK(clknet_leaf_25_clk),
    .RESET_B(net527),
    .D(_00211_),
    .Q_N(_00023_),
    .Q(\i_coord.y0[-2] ));
 sg13g2_dfrbp_1 \y0[12]$_DFFE_PP_  (.CLK(clknet_leaf_25_clk),
    .RESET_B(net528),
    .D(_00212_),
    .Q_N(_00024_),
    .Q(\i_coord.y0[-1] ));
 sg13g2_dfrbp_1 \y0[13]$_DFFE_PP_  (.CLK(clknet_leaf_6_clk),
    .RESET_B(net529),
    .D(_00213_),
    .Q_N(_00025_),
    .Q(\i_coord.y0[0] ));
 sg13g2_dfrbp_1 \y0[14]$_DFFE_PP_  (.CLK(clknet_leaf_7_clk),
    .RESET_B(net530),
    .D(_00214_),
    .Q_N(_07518_),
    .Q(\i_coord.y0[1] ));
 sg13g2_dfrbp_1 \y0[1]$_DFFE_PP_  (.CLK(clknet_leaf_12_clk),
    .RESET_B(net531),
    .D(_00215_),
    .Q_N(_07517_),
    .Q(\i_coord.y0[-12] ));
 sg13g2_dfrbp_1 \y0[2]$_DFFE_PP_  (.CLK(clknet_leaf_12_clk),
    .RESET_B(net532),
    .D(_00216_),
    .Q_N(_07516_),
    .Q(\i_coord.y0[-11] ));
 sg13g2_dfrbp_1 \y0[3]$_DFFE_PP_  (.CLK(clknet_leaf_11_clk),
    .RESET_B(net533),
    .D(_00217_),
    .Q_N(_07515_),
    .Q(\i_coord.y0[-10] ));
 sg13g2_dfrbp_1 \y0[4]$_DFFE_PP_  (.CLK(clknet_leaf_9_clk),
    .RESET_B(net534),
    .D(_00218_),
    .Q_N(_00018_),
    .Q(\i_coord.y0[-9] ));
 sg13g2_dfrbp_1 \y0[5]$_DFFE_PP_  (.CLK(clknet_leaf_10_clk),
    .RESET_B(net535),
    .D(_00219_),
    .Q_N(_07514_),
    .Q(\i_coord.y0[-8] ));
 sg13g2_dfrbp_1 \y0[6]$_DFFE_PP_  (.CLK(clknet_leaf_10_clk),
    .RESET_B(net536),
    .D(_00220_),
    .Q_N(_00019_),
    .Q(\i_coord.y0[-7] ));
 sg13g2_dfrbp_1 \y0[7]$_DFFE_PP_  (.CLK(clknet_leaf_10_clk),
    .RESET_B(net537),
    .D(_00221_),
    .Q_N(_07513_),
    .Q(\i_coord.y0[-6] ));
 sg13g2_dfrbp_1 \y0[8]$_DFFE_PP_  (.CLK(clknet_leaf_10_clk),
    .RESET_B(net538),
    .D(_00222_),
    .Q_N(_00021_),
    .Q(\i_coord.y0[-5] ));
 sg13g2_dfrbp_1 \y0[9]$_DFFE_PP_  (.CLK(clknet_leaf_10_clk),
    .RESET_B(net539),
    .D(_00223_),
    .Q_N(_00020_),
    .Q(\i_coord.y0[-4] ));
 sg13g2_dfrbp_1 \y[0]$_DFFE_PP_  (.CLK(clknet_leaf_22_clk),
    .RESET_B(net540),
    .D(_00224_),
    .Q_N(_00035_),
    .Q(\i_mandel.i_sq_y.x[-13] ));
 sg13g2_dfrbp_1 \y[10]$_DFFE_PP_  (.CLK(clknet_leaf_21_clk),
    .RESET_B(net541),
    .D(_00225_),
    .Q_N(_00041_),
    .Q(\i_mandel.i_sq_y.x[-3] ));
 sg13g2_dfrbp_1 \y[11]$_DFFE_PP_  (.CLK(clknet_leaf_21_clk),
    .RESET_B(net542),
    .D(_00226_),
    .Q_N(_00040_),
    .Q(\i_mandel.i_sq_y.x[-2] ));
 sg13g2_dfrbp_1 \y[12]$_DFFE_PP_  (.CLK(clknet_leaf_23_clk),
    .RESET_B(net543),
    .D(_00227_),
    .Q_N(_00039_),
    .Q(\i_mandel.i_sq_y.x[-1] ));
 sg13g2_dfrbp_1 \y[13]$_DFFE_PP_  (.CLK(clknet_leaf_21_clk),
    .RESET_B(net544),
    .D(_00228_),
    .Q_N(_00038_),
    .Q(\i_mandel.i_sq_y.x[0] ));
 sg13g2_dfrbp_1 \y[14]$_DFFE_PP_  (.CLK(clknet_leaf_21_clk),
    .RESET_B(net545),
    .D(_00229_),
    .Q_N(_00037_),
    .Q(\i_mandel.i_sq_y.x[1] ));
 sg13g2_dfrbp_1 \y[15]$_DFFE_PP_  (.CLK(clknet_leaf_21_clk),
    .RESET_B(net546),
    .D(_00230_),
    .Q_N(_00036_),
    .Q(\i_mandel.i_sq_y.x[2] ));
 sg13g2_dfrbp_1 \y[1]$_DFFE_PP_  (.CLK(clknet_leaf_21_clk),
    .RESET_B(net547),
    .D(_00231_),
    .Q_N(_07512_),
    .Q(\i_mandel.i_sq_y.x[-12] ));
 sg13g2_dfrbp_1 \y[2]$_DFFE_PP_  (.CLK(clknet_leaf_22_clk),
    .RESET_B(net548),
    .D(_00232_),
    .Q_N(_07511_),
    .Q(\i_mandel.i_sq_y.x[-11] ));
 sg13g2_dfrbp_1 \y[3]$_DFFE_PP_  (.CLK(clknet_leaf_21_clk),
    .RESET_B(net549),
    .D(_00233_),
    .Q_N(_07510_),
    .Q(\i_mandel.i_sq_y.x[-10] ));
 sg13g2_dfrbp_1 \y[4]$_DFFE_PP_  (.CLK(clknet_leaf_23_clk),
    .RESET_B(net550),
    .D(_00234_),
    .Q_N(_07509_),
    .Q(\i_mandel.i_sq_y.x[-9] ));
 sg13g2_dfrbp_1 \y[5]$_DFFE_PP_  (.CLK(clknet_leaf_23_clk),
    .RESET_B(net551),
    .D(_00235_),
    .Q_N(_07508_),
    .Q(\i_mandel.i_sq_y.x[-8] ));
 sg13g2_dfrbp_1 \y[6]$_DFFE_PP_  (.CLK(clknet_leaf_23_clk),
    .RESET_B(net552),
    .D(_00236_),
    .Q_N(_07507_),
    .Q(\i_mandel.i_sq_y.x[-7] ));
 sg13g2_dfrbp_1 \y[7]$_DFFE_PP_  (.CLK(clknet_leaf_23_clk),
    .RESET_B(net553),
    .D(_00237_),
    .Q_N(_00003_),
    .Q(\i_mandel.i_sq_y.x[-6] ));
 sg13g2_dfrbp_1 \y[8]$_DFFE_PP_  (.CLK(clknet_leaf_23_clk),
    .RESET_B(net554),
    .D(_00238_),
    .Q_N(_00043_),
    .Q(\i_mandel.i_sq_y.x[-5] ));
 sg13g2_dfrbp_1 \y[9]$_DFFE_PP_  (.CLK(clknet_leaf_21_clk),
    .RESET_B(net555),
    .D(_00239_),
    .Q_N(_00042_),
    .Q(\i_mandel.i_sq_y.x[-4] ));
 sg13g2_buf_1 input1 (.A(ui_in[4]),
    .X(net1));
 sg13g2_buf_1 input2 (.A(uio_in[1]),
    .X(net2));
 sg13g2_buf_1 input3 (.A(uio_in[5]),
    .X(net3));
 sg13g2_buf_1 input4 (.A(uio_in[6]),
    .X(net4));
 sg13g2_buf_1 input5 (.A(uio_in[7]),
    .X(net5));
 sg13g2_buf_1 output6 (.A(net6),
    .X(uo_out[0]));
 sg13g2_buf_1 output7 (.A(net7),
    .X(uo_out[1]));
 sg13g2_buf_1 output8 (.A(net8),
    .X(uo_out[2]));
 sg13g2_buf_1 output9 (.A(net9),
    .X(uo_out[3]));
 sg13g2_buf_1 output10 (.A(net10),
    .X(uo_out[4]));
 sg13g2_buf_1 output11 (.A(net11),
    .X(uo_out[5]));
 sg13g2_buf_1 output12 (.A(net12),
    .X(uo_out[6]));
 sg13g2_buf_1 output13 (.A(net13),
    .X(uo_out[7]));
 sg13g2_buf_2 fanout14 (.A(_04718_),
    .X(net14));
 sg13g2_buf_4 fanout15 (.X(net15),
    .A(_05012_));
 sg13g2_buf_4 fanout16 (.X(net16),
    .A(_04876_));
 sg13g2_buf_2 fanout17 (.A(_04717_),
    .X(net17));
 sg13g2_buf_2 fanout18 (.A(_03697_),
    .X(net18));
 sg13g2_buf_2 fanout19 (.A(_03626_),
    .X(net19));
 sg13g2_buf_2 fanout20 (.A(_03607_),
    .X(net20));
 sg13g2_buf_2 fanout21 (.A(_03622_),
    .X(net21));
 sg13g2_buf_2 fanout22 (.A(_00810_),
    .X(net22));
 sg13g2_buf_2 fanout23 (.A(_00718_),
    .X(net23));
 sg13g2_buf_2 fanout24 (.A(_02891_),
    .X(net24));
 sg13g2_buf_2 fanout25 (.A(_03647_),
    .X(net25));
 sg13g2_buf_2 fanout26 (.A(_02835_),
    .X(net26));
 sg13g2_buf_2 fanout27 (.A(_00377_),
    .X(net27));
 sg13g2_buf_2 fanout28 (.A(_06647_),
    .X(net28));
 sg13g2_buf_2 fanout29 (.A(_01998_),
    .X(net29));
 sg13g2_buf_2 fanout30 (.A(_07503_),
    .X(net30));
 sg13g2_buf_2 fanout31 (.A(_02329_),
    .X(net31));
 sg13g2_buf_2 fanout32 (.A(_01980_),
    .X(net32));
 sg13g2_buf_2 fanout33 (.A(_00974_),
    .X(net33));
 sg13g2_buf_2 fanout34 (.A(_07282_),
    .X(net34));
 sg13g2_buf_2 fanout35 (.A(_01659_),
    .X(net35));
 sg13g2_buf_2 fanout36 (.A(_02507_),
    .X(net36));
 sg13g2_buf_2 fanout37 (.A(_04324_),
    .X(net37));
 sg13g2_buf_2 fanout38 (.A(_02948_),
    .X(net38));
 sg13g2_buf_2 fanout39 (.A(_02705_),
    .X(net39));
 sg13g2_buf_2 fanout40 (.A(_02468_),
    .X(net40));
 sg13g2_buf_2 fanout41 (.A(_05019_),
    .X(net41));
 sg13g2_buf_2 fanout42 (.A(_04561_),
    .X(net42));
 sg13g2_buf_2 fanout43 (.A(_04161_),
    .X(net43));
 sg13g2_buf_2 fanout44 (.A(_01151_),
    .X(net44));
 sg13g2_buf_2 fanout45 (.A(_07277_),
    .X(net45));
 sg13g2_buf_2 fanout46 (.A(_05744_),
    .X(net46));
 sg13g2_buf_2 fanout47 (.A(_04432_),
    .X(net47));
 sg13g2_buf_2 fanout48 (.A(_04342_),
    .X(net48));
 sg13g2_buf_2 fanout49 (.A(_04160_),
    .X(net49));
 sg13g2_buf_2 fanout50 (.A(_03240_),
    .X(net50));
 sg13g2_buf_2 fanout51 (.A(_01871_),
    .X(net51));
 sg13g2_buf_2 fanout52 (.A(_00893_),
    .X(net52));
 sg13g2_buf_2 fanout53 (.A(_04648_),
    .X(net53));
 sg13g2_buf_2 fanout54 (.A(_04484_),
    .X(net54));
 sg13g2_buf_2 fanout55 (.A(_04341_),
    .X(net55));
 sg13g2_buf_2 fanout56 (.A(_04335_),
    .X(net56));
 sg13g2_buf_2 fanout57 (.A(_04328_),
    .X(net57));
 sg13g2_buf_2 fanout58 (.A(_04321_),
    .X(net58));
 sg13g2_buf_2 fanout59 (.A(_04159_),
    .X(net59));
 sg13g2_buf_2 fanout60 (.A(_03275_),
    .X(net60));
 sg13g2_buf_2 fanout61 (.A(_01862_),
    .X(net61));
 sg13g2_buf_2 fanout62 (.A(_01691_),
    .X(net62));
 sg13g2_buf_2 fanout63 (.A(_01620_),
    .X(net63));
 sg13g2_buf_2 fanout64 (.A(_05675_),
    .X(net64));
 sg13g2_buf_2 fanout65 (.A(_04617_),
    .X(net65));
 sg13g2_buf_2 fanout66 (.A(_04146_),
    .X(net66));
 sg13g2_buf_2 fanout67 (.A(_00381_),
    .X(net67));
 sg13g2_buf_2 fanout68 (.A(_00260_),
    .X(net68));
 sg13g2_buf_2 fanout69 (.A(_06826_),
    .X(net69));
 sg13g2_buf_2 fanout70 (.A(_05555_),
    .X(net70));
 sg13g2_buf_2 fanout71 (.A(_04650_),
    .X(net71));
 sg13g2_buf_2 fanout72 (.A(_04603_),
    .X(net72));
 sg13g2_buf_2 fanout73 (.A(_04573_),
    .X(net73));
 sg13g2_buf_2 fanout74 (.A(_04569_),
    .X(net74));
 sg13g2_buf_2 fanout75 (.A(_04556_),
    .X(net75));
 sg13g2_buf_2 fanout76 (.A(_04480_),
    .X(net76));
 sg13g2_buf_2 fanout77 (.A(_04144_),
    .X(net77));
 sg13g2_buf_2 fanout78 (.A(_02028_),
    .X(net78));
 sg13g2_buf_2 fanout79 (.A(_02023_),
    .X(net79));
 sg13g2_buf_2 fanout80 (.A(_07075_),
    .X(net80));
 sg13g2_buf_2 fanout81 (.A(_04576_),
    .X(net81));
 sg13g2_buf_2 fanout82 (.A(_04495_),
    .X(net82));
 sg13g2_buf_2 fanout83 (.A(_04479_),
    .X(net83));
 sg13g2_buf_2 fanout84 (.A(_01609_),
    .X(net84));
 sg13g2_buf_2 fanout85 (.A(_00267_),
    .X(net85));
 sg13g2_buf_2 fanout86 (.A(_06802_),
    .X(net86));
 sg13g2_buf_2 fanout87 (.A(_06594_),
    .X(net87));
 sg13g2_buf_2 fanout88 (.A(_04217_),
    .X(net88));
 sg13g2_buf_2 fanout89 (.A(_03901_),
    .X(net89));
 sg13g2_buf_2 fanout90 (.A(_01927_),
    .X(net90));
 sg13g2_buf_2 fanout91 (.A(_01684_),
    .X(net91));
 sg13g2_buf_2 fanout92 (.A(_01202_),
    .X(net92));
 sg13g2_buf_2 fanout93 (.A(_00551_),
    .X(net93));
 sg13g2_buf_2 fanout94 (.A(_07483_),
    .X(net94));
 sg13g2_buf_2 fanout95 (.A(_05060_),
    .X(net95));
 sg13g2_buf_2 fanout96 (.A(_07240_),
    .X(net96));
 sg13g2_buf_2 fanout97 (.A(_06292_),
    .X(net97));
 sg13g2_buf_2 fanout98 (.A(_04956_),
    .X(net98));
 sg13g2_buf_2 fanout99 (.A(_04613_),
    .X(net99));
 sg13g2_buf_2 fanout100 (.A(_04600_),
    .X(net100));
 sg13g2_buf_2 fanout101 (.A(_04577_),
    .X(net101));
 sg13g2_buf_2 fanout102 (.A(_04216_),
    .X(net102));
 sg13g2_buf_2 fanout103 (.A(_04164_),
    .X(net103));
 sg13g2_buf_2 fanout104 (.A(_04151_),
    .X(net104));
 sg13g2_buf_2 fanout105 (.A(_03270_),
    .X(net105));
 sg13g2_buf_2 fanout106 (.A(_02059_),
    .X(net106));
 sg13g2_buf_2 fanout107 (.A(_01737_),
    .X(net107));
 sg13g2_buf_2 fanout108 (.A(_01678_),
    .X(net108));
 sg13g2_buf_2 fanout109 (.A(_01661_),
    .X(net109));
 sg13g2_buf_2 fanout110 (.A(_01557_),
    .X(net110));
 sg13g2_buf_2 fanout111 (.A(_00819_),
    .X(net111));
 sg13g2_buf_2 fanout112 (.A(_06833_),
    .X(net112));
 sg13g2_buf_2 fanout113 (.A(_05317_),
    .X(net113));
 sg13g2_buf_2 fanout114 (.A(_05004_),
    .X(net114));
 sg13g2_buf_2 fanout115 (.A(_04719_),
    .X(net115));
 sg13g2_buf_2 fanout116 (.A(_04703_),
    .X(net116));
 sg13g2_buf_2 fanout117 (.A(_04560_),
    .X(net117));
 sg13g2_buf_2 fanout118 (.A(_04558_),
    .X(net118));
 sg13g2_buf_2 fanout119 (.A(_04055_),
    .X(net119));
 sg13g2_buf_2 fanout120 (.A(_02109_),
    .X(net120));
 sg13g2_buf_2 fanout121 (.A(_02057_),
    .X(net121));
 sg13g2_buf_2 fanout122 (.A(_02029_),
    .X(net122));
 sg13g2_buf_2 fanout123 (.A(_02005_),
    .X(net123));
 sg13g2_buf_2 fanout124 (.A(_01921_),
    .X(net124));
 sg13g2_buf_2 fanout125 (.A(_01732_),
    .X(net125));
 sg13g2_buf_2 fanout126 (.A(_01679_),
    .X(net126));
 sg13g2_buf_2 fanout127 (.A(_00382_),
    .X(net127));
 sg13g2_buf_2 fanout128 (.A(_00361_),
    .X(net128));
 sg13g2_buf_2 fanout129 (.A(_07452_),
    .X(net129));
 sg13g2_buf_2 fanout130 (.A(_07309_),
    .X(net130));
 sg13g2_buf_2 fanout131 (.A(_04401_),
    .X(net131));
 sg13g2_buf_2 fanout132 (.A(_06665_),
    .X(net132));
 sg13g2_buf_2 fanout133 (.A(_05801_),
    .X(net133));
 sg13g2_buf_2 fanout134 (.A(_05765_),
    .X(net134));
 sg13g2_buf_2 fanout135 (.A(_05339_),
    .X(net135));
 sg13g2_buf_2 fanout136 (.A(_04971_),
    .X(net136));
 sg13g2_buf_2 fanout137 (.A(_04961_),
    .X(net137));
 sg13g2_buf_2 fanout138 (.A(_04955_),
    .X(net138));
 sg13g2_buf_2 fanout139 (.A(_04557_),
    .X(net139));
 sg13g2_buf_2 fanout140 (.A(_04483_),
    .X(net140));
 sg13g2_buf_2 fanout141 (.A(_04482_),
    .X(net141));
 sg13g2_buf_2 fanout142 (.A(_04009_),
    .X(net142));
 sg13g2_buf_2 fanout143 (.A(_03278_),
    .X(net143));
 sg13g2_buf_2 fanout144 (.A(_03213_),
    .X(net144));
 sg13g2_buf_2 fanout145 (.A(_02770_),
    .X(net145));
 sg13g2_buf_2 fanout146 (.A(_02304_),
    .X(net146));
 sg13g2_buf_2 fanout147 (.A(_02292_),
    .X(net147));
 sg13g2_buf_2 fanout148 (.A(_02040_),
    .X(net148));
 sg13g2_buf_2 fanout149 (.A(_02032_),
    .X(net149));
 sg13g2_buf_2 fanout150 (.A(_02019_),
    .X(net150));
 sg13g2_buf_2 fanout151 (.A(_02017_),
    .X(net151));
 sg13g2_buf_2 fanout152 (.A(_02014_),
    .X(net152));
 sg13g2_buf_2 fanout153 (.A(_02008_),
    .X(net153));
 sg13g2_buf_2 fanout154 (.A(_01490_),
    .X(net154));
 sg13g2_buf_2 fanout155 (.A(_01330_),
    .X(net155));
 sg13g2_buf_2 fanout156 (.A(_00371_),
    .X(net156));
 sg13g2_buf_2 fanout157 (.A(_00362_),
    .X(net157));
 sg13g2_buf_2 fanout158 (.A(_00331_),
    .X(net158));
 sg13g2_buf_2 fanout159 (.A(_00281_),
    .X(net159));
 sg13g2_buf_2 fanout160 (.A(_06189_),
    .X(net160));
 sg13g2_buf_2 fanout161 (.A(_05925_),
    .X(net161));
 sg13g2_buf_2 fanout162 (.A(_04968_),
    .X(net162));
 sg13g2_buf_2 fanout163 (.A(_05763_),
    .X(net163));
 sg13g2_buf_2 fanout164 (.A(_05510_),
    .X(net164));
 sg13g2_buf_2 fanout165 (.A(_05305_),
    .X(net165));
 sg13g2_buf_2 fanout166 (.A(_05192_),
    .X(net166));
 sg13g2_buf_2 fanout167 (.A(_04031_),
    .X(net167));
 sg13g2_buf_2 fanout168 (.A(_04004_),
    .X(net168));
 sg13g2_buf_2 fanout169 (.A(_03018_),
    .X(net169));
 sg13g2_buf_2 fanout170 (.A(_02739_),
    .X(net170));
 sg13g2_buf_2 fanout171 (.A(_02360_),
    .X(net171));
 sg13g2_buf_2 fanout172 (.A(_02333_),
    .X(net172));
 sg13g2_buf_2 fanout173 (.A(_02303_),
    .X(net173));
 sg13g2_buf_2 fanout174 (.A(_02290_),
    .X(net174));
 sg13g2_buf_2 fanout175 (.A(_02282_),
    .X(net175));
 sg13g2_buf_2 fanout176 (.A(_02054_),
    .X(net176));
 sg13g2_buf_2 fanout177 (.A(_02031_),
    .X(net177));
 sg13g2_buf_2 fanout178 (.A(_02016_),
    .X(net178));
 sg13g2_buf_2 fanout179 (.A(_02013_),
    .X(net179));
 sg13g2_buf_2 fanout180 (.A(_02007_),
    .X(net180));
 sg13g2_buf_2 fanout181 (.A(_01983_),
    .X(net181));
 sg13g2_buf_2 fanout182 (.A(_01982_),
    .X(net182));
 sg13g2_buf_2 fanout183 (.A(_01926_),
    .X(net183));
 sg13g2_buf_2 fanout184 (.A(_01764_),
    .X(net184));
 sg13g2_buf_2 fanout185 (.A(_01761_),
    .X(net185));
 sg13g2_buf_2 fanout186 (.A(_01624_),
    .X(net186));
 sg13g2_buf_2 fanout187 (.A(_01560_),
    .X(net187));
 sg13g2_buf_2 fanout188 (.A(_01542_),
    .X(net188));
 sg13g2_buf_2 fanout189 (.A(_01523_),
    .X(net189));
 sg13g2_buf_2 fanout190 (.A(_01512_),
    .X(net190));
 sg13g2_buf_2 fanout191 (.A(_01497_),
    .X(net191));
 sg13g2_buf_2 fanout192 (.A(_01489_),
    .X(net192));
 sg13g2_buf_2 fanout193 (.A(_00830_),
    .X(net193));
 sg13g2_buf_2 fanout194 (.A(_00753_),
    .X(net194));
 sg13g2_buf_2 fanout195 (.A(_00450_),
    .X(net195));
 sg13g2_buf_2 fanout196 (.A(_00429_),
    .X(net196));
 sg13g2_buf_2 fanout197 (.A(_00415_),
    .X(net197));
 sg13g2_buf_2 fanout198 (.A(_00368_),
    .X(net198));
 sg13g2_buf_2 fanout199 (.A(_00366_),
    .X(net199));
 sg13g2_buf_2 fanout200 (.A(_00363_),
    .X(net200));
 sg13g2_buf_2 fanout201 (.A(_00289_),
    .X(net201));
 sg13g2_buf_2 fanout202 (.A(_00283_),
    .X(net202));
 sg13g2_buf_2 fanout203 (.A(_00245_),
    .X(net203));
 sg13g2_buf_2 fanout204 (.A(_07500_),
    .X(net204));
 sg13g2_buf_2 fanout205 (.A(_07466_),
    .X(net205));
 sg13g2_buf_2 fanout206 (.A(_07453_),
    .X(net206));
 sg13g2_buf_2 fanout207 (.A(_07357_),
    .X(net207));
 sg13g2_buf_2 fanout208 (.A(_06255_),
    .X(net208));
 sg13g2_buf_2 fanout209 (.A(_05793_),
    .X(net209));
 sg13g2_buf_2 fanout210 (.A(_05694_),
    .X(net210));
 sg13g2_buf_2 fanout211 (.A(_05507_),
    .X(net211));
 sg13g2_buf_2 fanout212 (.A(_05233_),
    .X(net212));
 sg13g2_buf_2 fanout213 (.A(_05179_),
    .X(net213));
 sg13g2_buf_2 fanout214 (.A(_05027_),
    .X(net214));
 sg13g2_buf_2 fanout215 (.A(_04988_),
    .X(net215));
 sg13g2_buf_2 fanout216 (.A(_04959_),
    .X(net216));
 sg13g2_buf_2 fanout217 (.A(_04801_),
    .X(net217));
 sg13g2_buf_2 fanout218 (.A(_07205_),
    .X(net218));
 sg13g2_buf_2 fanout219 (.A(_05314_),
    .X(net219));
 sg13g2_buf_2 fanout220 (.A(_03961_),
    .X(net220));
 sg13g2_buf_2 fanout221 (.A(_03950_),
    .X(net221));
 sg13g2_buf_2 fanout222 (.A(_03936_),
    .X(net222));
 sg13g2_buf_2 fanout223 (.A(_03930_),
    .X(net223));
 sg13g2_buf_2 fanout224 (.A(_03923_),
    .X(net224));
 sg13g2_buf_2 fanout225 (.A(_03918_),
    .X(net225));
 sg13g2_buf_2 fanout226 (.A(_03904_),
    .X(net226));
 sg13g2_buf_2 fanout227 (.A(_02332_),
    .X(net227));
 sg13g2_buf_2 fanout228 (.A(_02289_),
    .X(net228));
 sg13g2_buf_2 fanout229 (.A(_02288_),
    .X(net229));
 sg13g2_buf_2 fanout230 (.A(_02041_),
    .X(net230));
 sg13g2_buf_2 fanout231 (.A(_02034_),
    .X(net231));
 sg13g2_buf_2 fanout232 (.A(_02030_),
    .X(net232));
 sg13g2_buf_2 fanout233 (.A(_02015_),
    .X(net233));
 sg13g2_buf_2 fanout234 (.A(_02009_),
    .X(net234));
 sg13g2_buf_2 fanout235 (.A(_02006_),
    .X(net235));
 sg13g2_buf_2 fanout236 (.A(_02002_),
    .X(net236));
 sg13g2_buf_2 fanout237 (.A(_01990_),
    .X(net237));
 sg13g2_buf_2 fanout238 (.A(_01981_),
    .X(net238));
 sg13g2_buf_2 fanout239 (.A(_01925_),
    .X(net239));
 sg13g2_buf_2 fanout240 (.A(_01833_),
    .X(net240));
 sg13g2_buf_2 fanout241 (.A(_01559_),
    .X(net241));
 sg13g2_buf_2 fanout242 (.A(_01555_),
    .X(net242));
 sg13g2_buf_2 fanout243 (.A(_01522_),
    .X(net243));
 sg13g2_buf_2 fanout244 (.A(_01496_),
    .X(net244));
 sg13g2_buf_2 fanout245 (.A(_01493_),
    .X(net245));
 sg13g2_buf_2 fanout246 (.A(_01488_),
    .X(net246));
 sg13g2_buf_2 fanout247 (.A(_00537_),
    .X(net247));
 sg13g2_buf_2 fanout248 (.A(_00333_),
    .X(net248));
 sg13g2_buf_2 fanout249 (.A(_00298_),
    .X(net249));
 sg13g2_buf_2 fanout250 (.A(_07506_),
    .X(net250));
 sg13g2_buf_2 fanout251 (.A(_07505_),
    .X(net251));
 sg13g2_buf_2 fanout252 (.A(_07496_),
    .X(net252));
 sg13g2_buf_2 fanout253 (.A(_07480_),
    .X(net253));
 sg13g2_buf_2 fanout254 (.A(_07479_),
    .X(net254));
 sg13g2_buf_2 fanout255 (.A(_07456_),
    .X(net255));
 sg13g2_buf_2 fanout256 (.A(_07319_),
    .X(net256));
 sg13g2_buf_2 fanout257 (.A(_07213_),
    .X(net257));
 sg13g2_buf_2 fanout258 (.A(_06651_),
    .X(net258));
 sg13g2_buf_2 fanout259 (.A(_06552_),
    .X(net259));
 sg13g2_buf_2 fanout260 (.A(_05562_),
    .X(net260));
 sg13g2_buf_2 fanout261 (.A(_05332_),
    .X(net261));
 sg13g2_buf_2 fanout262 (.A(_05169_),
    .X(net262));
 sg13g2_buf_2 fanout263 (.A(_05080_),
    .X(net263));
 sg13g2_buf_2 fanout264 (.A(_05017_),
    .X(net264));
 sg13g2_buf_2 fanout265 (.A(_04978_),
    .X(net265));
 sg13g2_buf_2 fanout266 (.A(_04907_),
    .X(net266));
 sg13g2_buf_2 fanout267 (.A(_04834_),
    .X(net267));
 sg13g2_buf_2 fanout268 (.A(_04790_),
    .X(net268));
 sg13g2_buf_2 fanout269 (.A(_04746_),
    .X(net269));
 sg13g2_buf_2 fanout270 (.A(_04595_),
    .X(net270));
 sg13g2_buf_2 fanout271 (.A(_04965_),
    .X(net271));
 sg13g2_buf_2 fanout272 (.A(_03926_),
    .X(net272));
 sg13g2_buf_2 fanout273 (.A(_03922_),
    .X(net273));
 sg13g2_buf_2 fanout274 (.A(_03885_),
    .X(net274));
 sg13g2_buf_2 fanout275 (.A(_02313_),
    .X(net275));
 sg13g2_buf_2 fanout276 (.A(_02010_),
    .X(net276));
 sg13g2_buf_2 fanout277 (.A(_02001_),
    .X(net277));
 sg13g2_buf_2 fanout278 (.A(_01986_),
    .X(net278));
 sg13g2_buf_2 fanout279 (.A(_01790_),
    .X(net279));
 sg13g2_buf_2 fanout280 (.A(_01779_),
    .X(net280));
 sg13g2_buf_2 fanout281 (.A(_01640_),
    .X(net281));
 sg13g2_buf_2 fanout282 (.A(_01628_),
    .X(net282));
 sg13g2_buf_2 fanout283 (.A(_01611_),
    .X(net283));
 sg13g2_buf_2 fanout284 (.A(_01594_),
    .X(net284));
 sg13g2_buf_2 fanout285 (.A(_01540_),
    .X(net285));
 sg13g2_buf_2 fanout286 (.A(_01537_),
    .X(net286));
 sg13g2_buf_2 fanout287 (.A(_01530_),
    .X(net287));
 sg13g2_buf_2 fanout288 (.A(_01529_),
    .X(net288));
 sg13g2_buf_2 fanout289 (.A(_01527_),
    .X(net289));
 sg13g2_buf_2 fanout290 (.A(_01516_),
    .X(net290));
 sg13g2_buf_2 fanout291 (.A(_01514_),
    .X(net291));
 sg13g2_buf_2 fanout292 (.A(_01500_),
    .X(net292));
 sg13g2_buf_2 fanout293 (.A(_01487_),
    .X(net293));
 sg13g2_buf_2 fanout294 (.A(_01328_),
    .X(net294));
 sg13g2_buf_2 fanout295 (.A(_07504_),
    .X(net295));
 sg13g2_buf_2 fanout296 (.A(_07498_),
    .X(net296));
 sg13g2_buf_2 fanout297 (.A(_07355_),
    .X(net297));
 sg13g2_buf_2 fanout298 (.A(_05782_),
    .X(net298));
 sg13g2_buf_2 fanout299 (.A(_05771_),
    .X(net299));
 sg13g2_buf_2 fanout300 (.A(_05310_),
    .X(net300));
 sg13g2_buf_2 fanout301 (.A(_05070_),
    .X(net301));
 sg13g2_buf_2 fanout302 (.A(_05008_),
    .X(net302));
 sg13g2_buf_2 fanout303 (.A(_04928_),
    .X(net303));
 sg13g2_buf_2 fanout304 (.A(_04897_),
    .X(net304));
 sg13g2_buf_2 fanout305 (.A(_04645_),
    .X(net305));
 sg13g2_buf_2 fanout306 (.A(_04626_),
    .X(net306));
 sg13g2_buf_2 fanout307 (.A(_04584_),
    .X(net307));
 sg13g2_buf_2 fanout308 (.A(_04574_),
    .X(net308));
 sg13g2_buf_2 fanout309 (.A(_04542_),
    .X(net309));
 sg13g2_buf_2 fanout310 (.A(_04488_),
    .X(net310));
 sg13g2_buf_2 fanout311 (.A(_04602_),
    .X(net311));
 sg13g2_buf_2 fanout312 (.A(_04583_),
    .X(net312));
 sg13g2_buf_2 fanout313 (.A(_04513_),
    .X(net313));
 sg13g2_buf_2 fanout314 (.A(_04503_),
    .X(net314));
 sg13g2_buf_2 fanout315 (.A(_04214_),
    .X(net315));
 sg13g2_buf_2 fanout316 (.A(_04208_),
    .X(net316));
 sg13g2_buf_2 fanout317 (.A(_04062_),
    .X(net317));
 sg13g2_buf_2 fanout318 (.A(_03999_),
    .X(net318));
 sg13g2_buf_2 fanout319 (.A(_03982_),
    .X(net319));
 sg13g2_buf_2 fanout320 (.A(_03921_),
    .X(net320));
 sg13g2_buf_2 fanout321 (.A(_03895_),
    .X(net321));
 sg13g2_buf_2 fanout322 (.A(_03886_),
    .X(net322));
 sg13g2_buf_2 fanout323 (.A(_01908_),
    .X(net323));
 sg13g2_buf_2 fanout324 (.A(_01508_),
    .X(net324));
 sg13g2_buf_2 fanout325 (.A(_01507_),
    .X(net325));
 sg13g2_buf_2 fanout326 (.A(_01499_),
    .X(net326));
 sg13g2_buf_2 fanout327 (.A(_01494_),
    .X(net327));
 sg13g2_buf_2 fanout328 (.A(_01491_),
    .X(net328));
 sg13g2_buf_2 fanout329 (.A(_07497_),
    .X(net329));
 sg13g2_buf_2 fanout330 (.A(_07315_),
    .X(net330));
 sg13g2_buf_2 fanout331 (.A(_05650_),
    .X(net331));
 sg13g2_buf_2 fanout332 (.A(_05453_),
    .X(net332));
 sg13g2_buf_2 fanout333 (.A(_04887_),
    .X(net333));
 sg13g2_buf_2 fanout334 (.A(_04812_),
    .X(net334));
 sg13g2_buf_2 fanout335 (.A(_04635_),
    .X(net335));
 sg13g2_buf_2 fanout336 (.A(_04021_),
    .X(net336));
 sg13g2_tielo _15151__337 (.L_LO(net337));
 sg13g2_tielo _15152__338 (.L_LO(net338));
 sg13g2_tielo _15153__339 (.L_LO(net339));
 sg13g2_tielo _15154__340 (.L_LO(net340));
 sg13g2_tielo _15155__341 (.L_LO(net341));
 sg13g2_tielo _15156__342 (.L_LO(net342));
 sg13g2_tielo _15157__343 (.L_LO(net343));
 sg13g2_tielo _15158__344 (.L_LO(net344));
 sg13g2_tielo _15159__345 (.L_LO(net345));
 sg13g2_tielo _15160__346 (.L_LO(net346));
 sg13g2_tielo _15161__347 (.L_LO(net347));
 sg13g2_tielo _15162__348 (.L_LO(net348));
 sg13g2_tielo _15163__349 (.L_LO(net349));
 sg13g2_tielo _15164__350 (.L_LO(net350));
 sg13g2_tielo _15165__351 (.L_LO(net351));
 sg13g2_tielo _15166__352 (.L_LO(net352));
 sg13g2_tiehi \i_coord.demo_update_delay$_SDFFE_PN0P__354  (.L_HI(net354));
 sg13g2_tiehi \i_coord.l_xip.state[0]$_SDFFCE_PP0P__355  (.L_HI(net355));
 sg13g2_tiehi \i_coord.l_xip.state[1]$_SDFFCE_PN1P__356  (.L_HI(net356));
 sg13g2_tiehi \i_coord.l_xip.state[2]$_SDFFCE_PN0P__357  (.L_HI(net357));
 sg13g2_tiehi \i_coord.l_xip.state[3]$_SDFFCE_PN1P__358  (.L_HI(net358));
 sg13g2_tiehi \i_coord.l_xip.state[4]$_SDFFCE_PN0P__359  (.L_HI(net359));
 sg13g2_tiehi \i_coord.l_xip.state[5]$_SDFFCE_PN0P__360  (.L_HI(net360));
 sg13g2_tiehi \i_coord.l_xip.state[6]$_SDFFCE_PN0P__361  (.L_HI(net361));
 sg13g2_tiehi \i_coord.l_xip.state[7]$_SDFFCE_PN1P__362  (.L_HI(net362));
 sg13g2_tiehi \i_coord.l_xip.state[8]$_SDFFCE_PN0P__363  (.L_HI(net363));
 sg13g2_tiehi \i_coord.l_xip.state[9]$_SDFFCE_PP0P__364  (.L_HI(net364));
 sg13g2_tiehi \i_coord.l_xir.state[0]$_SDFFCE_PN0P__365  (.L_HI(net365));
 sg13g2_tiehi \i_coord.l_xir.state[1]$_SDFFCE_PN0P__366  (.L_HI(net366));
 sg13g2_tiehi \i_coord.l_xir.state[2]$_SDFFCE_PN0P__367  (.L_HI(net367));
 sg13g2_tiehi \i_coord.l_xir.state[3]$_SDFFCE_PN0P__368  (.L_HI(net368));
 sg13g2_tiehi \i_coord.l_xir.state[4]$_SDFFCE_PN0P__369  (.L_HI(net369));
 sg13g2_tiehi \i_coord.l_xir.state[5]$_SDFFCE_PN0P__370  (.L_HI(net370));
 sg13g2_tiehi \i_coord.l_xir.state[6]$_SDFFCE_PN0P__371  (.L_HI(net371));
 sg13g2_tiehi \i_coord.l_xir.state[7]$_SDFFCE_PN0P__372  (.L_HI(net372));
 sg13g2_tiehi \i_coord.l_xl.state[10]$_SDFFCE_PN0P__373  (.L_HI(net373));
 sg13g2_tiehi \i_coord.l_xl.state[11]$_SDFFCE_PN0P__374  (.L_HI(net374));
 sg13g2_tiehi \i_coord.l_xl.state[12]$_SDFFCE_PN0P__375  (.L_HI(net375));
 sg13g2_tiehi \i_coord.l_xl.state[13]$_SDFFCE_PN0P__376  (.L_HI(net376));
 sg13g2_tiehi \i_coord.l_xl.state[14]$_SDFFCE_PN1P__377  (.L_HI(net377));
 sg13g2_tiehi \i_coord.l_xl.state[15]$_SDFFCE_PN1P__378  (.L_HI(net378));
 sg13g2_tiehi \i_coord.l_xl.state[3]$_SDFFCE_PN0P__379  (.L_HI(net379));
 sg13g2_tiehi \i_coord.l_xl.state[4]$_SDFFCE_PN0P__380  (.L_HI(net380));
 sg13g2_tiehi \i_coord.l_xl.state[5]$_SDFFCE_PN0P__381  (.L_HI(net381));
 sg13g2_tiehi \i_coord.l_xl.state[6]$_SDFFCE_PN0P__382  (.L_HI(net382));
 sg13g2_tiehi \i_coord.l_xl.state[7]$_SDFFCE_PN0P__383  (.L_HI(net383));
 sg13g2_tiehi \i_coord.l_xl.state[8]$_SDFFCE_PN0P__384  (.L_HI(net384));
 sg13g2_tiehi \i_coord.l_xl.state[9]$_SDFFCE_PN0P__385  (.L_HI(net385));
 sg13g2_tiehi \i_coord.l_yip.state[0]$_SDFFCE_PN0P__386  (.L_HI(net386));
 sg13g2_tiehi \i_coord.l_yip.state[1]$_SDFFCE_PN0P__387  (.L_HI(net387));
 sg13g2_tiehi \i_coord.l_yip.state[2]$_SDFFCE_PN0P__388  (.L_HI(net388));
 sg13g2_tiehi \i_coord.l_yip.state[3]$_SDFFCE_PN0P__389  (.L_HI(net389));
 sg13g2_tiehi \i_coord.l_yip.state[4]$_SDFFCE_PN0P__390  (.L_HI(net390));
 sg13g2_tiehi \i_coord.l_yip.state[5]$_SDFFCE_PN0P__391  (.L_HI(net391));
 sg13g2_tiehi \i_coord.l_yip.state[6]$_SDFFCE_PN0P__392  (.L_HI(net392));
 sg13g2_tiehi \i_coord.l_yip.state[7]$_SDFFCE_PN0P__393  (.L_HI(net393));
 sg13g2_tiehi \i_coord.l_yip.state[8]$_SDFFCE_PN0P__394  (.L_HI(net394));
 sg13g2_tiehi \i_coord.l_yip.state[9]$_SDFFCE_PN0P__395  (.L_HI(net395));
 sg13g2_tiehi \i_coord.l_yt.state[0]$_SDFFCE_PP0P__396  (.L_HI(net396));
 sg13g2_tiehi \i_coord.l_yt.state[10]$_SDFFCE_PN0P__397  (.L_HI(net397));
 sg13g2_tiehi \i_coord.l_yt.state[11]$_SDFFCE_PN0P__398  (.L_HI(net398));
 sg13g2_tiehi \i_coord.l_yt.state[12]$_SDFFCE_PN0P__399  (.L_HI(net399));
 sg13g2_tiehi \i_coord.l_yt.state[13]$_SDFFCE_PN0P__400  (.L_HI(net400));
 sg13g2_tiehi \i_coord.l_yt.state[14]$_SDFFCE_PN1P__401  (.L_HI(net401));
 sg13g2_tiehi \i_coord.l_yt.state[1]$_SDFFCE_PP0P__402  (.L_HI(net402));
 sg13g2_tiehi \i_coord.l_yt.state[2]$_SDFFCE_PN0P__403  (.L_HI(net403));
 sg13g2_tiehi \i_coord.l_yt.state[3]$_SDFFCE_PN0P__404  (.L_HI(net404));
 sg13g2_tiehi \i_coord.l_yt.state[4]$_SDFFCE_PN1P__405  (.L_HI(net405));
 sg13g2_tiehi \i_coord.l_yt.state[5]$_SDFFCE_PN1P__406  (.L_HI(net406));
 sg13g2_tiehi \i_coord.l_yt.state[6]$_SDFFCE_PN0P__407  (.L_HI(net407));
 sg13g2_tiehi \i_coord.l_yt.state[7]$_SDFFCE_PN1P__408  (.L_HI(net408));
 sg13g2_tiehi \i_coord.l_yt.state[8]$_SDFFCE_PN0P__409  (.L_HI(net409));
 sg13g2_tiehi \i_coord.l_yt.state[9]$_SDFFCE_PN0P__410  (.L_HI(net410));
 sg13g2_tiehi \i_coord.x_row_start[0]$_SDFFCE_PP0P__411  (.L_HI(net411));
 sg13g2_tiehi \i_coord.x_row_start[10]$_DFFE_PP__412  (.L_HI(net412));
 sg13g2_tiehi \i_coord.x_row_start[11]$_DFFE_PP__413  (.L_HI(net413));
 sg13g2_tiehi \i_coord.x_row_start[12]$_DFFE_PP__414  (.L_HI(net414));
 sg13g2_tiehi \i_coord.x_row_start[13]$_DFFE_PP__415  (.L_HI(net415));
 sg13g2_tiehi \i_coord.x_row_start[14]$_DFFE_PP__416  (.L_HI(net416));
 sg13g2_tiehi \i_coord.x_row_start[15]$_DFFE_PP__417  (.L_HI(net417));
 sg13g2_tiehi \i_coord.x_row_start[1]$_SDFFCE_PP0P__418  (.L_HI(net418));
 sg13g2_tiehi \i_coord.x_row_start[2]$_SDFFCE_PP0P__419  (.L_HI(net419));
 sg13g2_tiehi \i_coord.x_row_start[3]$_DFFE_PP__420  (.L_HI(net420));
 sg13g2_tiehi \i_coord.x_row_start[4]$_DFFE_PP__421  (.L_HI(net421));
 sg13g2_tiehi \i_coord.x_row_start[5]$_DFFE_PP__422  (.L_HI(net422));
 sg13g2_tiehi \i_coord.x_row_start[6]$_DFFE_PP__423  (.L_HI(net423));
 sg13g2_tiehi \i_coord.x_row_start[7]$_DFFE_PP__424  (.L_HI(net424));
 sg13g2_tiehi \i_coord.x_row_start[8]$_DFFE_PP__425  (.L_HI(net425));
 sg13g2_tiehi \i_coord.x_row_start[9]$_DFFE_PP__426  (.L_HI(net426));
 sg13g2_tiehi \i_coord.y_inc_row[0]$_SDFFE_PN1P__427  (.L_HI(net427));
 sg13g2_tiehi \i_coord.y_inc_row[1]$_SDFFE_PN1P__428  (.L_HI(net428));
 sg13g2_tiehi \i_coord.y_inc_row[2]$_SDFFE_PN0P__429  (.L_HI(net429));
 sg13g2_tiehi \i_coord.y_inc_row[3]$_SDFFE_PN1P__430  (.L_HI(net430));
 sg13g2_tiehi \i_coord.y_inc_row[4]$_SDFFE_PN1P__431  (.L_HI(net431));
 sg13g2_tiehi \i_coord.y_inc_row[5]$_SDFFE_PN1P__432  (.L_HI(net432));
 sg13g2_tiehi \i_coord.y_inc_row[6]$_SDFFE_PN0P__433  (.L_HI(net433));
 sg13g2_tiehi \i_coord.y_inc_row[7]$_SDFFE_PN1P__434  (.L_HI(net434));
 sg13g2_tiehi \i_coord.y_row_start[0]$_DFFE_PP__435  (.L_HI(net435));
 sg13g2_tiehi \i_coord.y_row_start[10]$_DFFE_PP__436  (.L_HI(net436));
 sg13g2_tiehi \i_coord.y_row_start[11]$_DFFE_PP__437  (.L_HI(net437));
 sg13g2_tiehi \i_coord.y_row_start[12]$_DFFE_PP__438  (.L_HI(net438));
 sg13g2_tiehi \i_coord.y_row_start[13]$_DFFE_PP__439  (.L_HI(net439));
 sg13g2_tiehi \i_coord.y_row_start[14]$_DFFE_PP__440  (.L_HI(net440));
 sg13g2_tiehi \i_coord.y_row_start[1]$_DFFE_PP__441  (.L_HI(net441));
 sg13g2_tiehi \i_coord.y_row_start[2]$_DFFE_PP__442  (.L_HI(net442));
 sg13g2_tiehi \i_coord.y_row_start[3]$_DFFE_PP__443  (.L_HI(net443));
 sg13g2_tiehi \i_coord.y_row_start[4]$_DFFE_PP__444  (.L_HI(net444));
 sg13g2_tiehi \i_coord.y_row_start[5]$_DFFE_PP__445  (.L_HI(net445));
 sg13g2_tiehi \i_coord.y_row_start[6]$_DFFE_PP__446  (.L_HI(net446));
 sg13g2_tiehi \i_coord.y_row_start[7]$_DFFE_PP__447  (.L_HI(net447));
 sg13g2_tiehi \i_coord.y_row_start[8]$_DFFE_PP__448  (.L_HI(net448));
 sg13g2_tiehi \i_coord.y_row_start[9]$_DFFE_PP__449  (.L_HI(net449));
 sg13g2_tiehi \i_vga.timing_hor.counter[0]$_SDFFE_PN0P__450  (.L_HI(net450));
 sg13g2_tiehi \i_vga.timing_hor.counter[10]$_SDFFE_PN1P__451  (.L_HI(net451));
 sg13g2_tiehi \i_vga.timing_hor.counter[1]$_SDFFE_PN0P__452  (.L_HI(net452));
 sg13g2_tiehi \i_vga.timing_hor.counter[2]$_SDFFE_PN0P__453  (.L_HI(net453));
 sg13g2_tiehi \i_vga.timing_hor.counter[3]$_SDFFE_PN0P__454  (.L_HI(net454));
 sg13g2_tiehi \i_vga.timing_hor.counter[4]$_SDFFE_PN1P__455  (.L_HI(net455));
 sg13g2_tiehi \i_vga.timing_hor.counter[5]$_SDFFE_PN0P__456  (.L_HI(net456));
 sg13g2_tiehi \i_vga.timing_hor.counter[6]$_SDFFE_PN1P__457  (.L_HI(net457));
 sg13g2_tiehi \i_vga.timing_hor.counter[7]$_SDFFE_PN0P__458  (.L_HI(net458));
 sg13g2_tiehi \i_vga.timing_hor.counter[8]$_SDFFE_PN1P__459  (.L_HI(net459));
 sg13g2_tiehi \i_vga.timing_hor.counter[9]$_SDFFE_PN1P__460  (.L_HI(net460));
 sg13g2_tiehi \i_vga.timing_hor.sync$_DFF_P__461  (.L_HI(net461));
 sg13g2_tiehi \i_vga.timing_ver.counter[0]$_SDFFE_PN1P__462  (.L_HI(net462));
 sg13g2_tiehi \i_vga.timing_ver.counter[1]$_SDFFE_PN0P__463  (.L_HI(net463));
 sg13g2_tiehi \i_vga.timing_ver.counter[2]$_SDFFE_PN1P__464  (.L_HI(net464));
 sg13g2_tiehi \i_vga.timing_ver.counter[3]$_SDFFE_PN1P__465  (.L_HI(net465));
 sg13g2_tiehi \i_vga.timing_ver.counter[4]$_SDFFE_PN0P__466  (.L_HI(net466));
 sg13g2_tiehi \i_vga.timing_ver.counter[5]$_SDFFE_PN1P__467  (.L_HI(net467));
 sg13g2_tiehi \i_vga.timing_ver.counter[6]$_SDFFE_PN1P__468  (.L_HI(net468));
 sg13g2_tiehi \i_vga.timing_ver.counter[7]$_SDFFE_PN1P__469  (.L_HI(net469));
 sg13g2_tiehi \i_vga.timing_ver.counter[8]$_SDFFE_PN1P__470  (.L_HI(net470));
 sg13g2_tiehi \i_vga.timing_ver.counter[9]$_SDFFE_PN1P__471  (.L_HI(net471));
 sg13g2_tiehi \i_vga.timing_ver.sync$_DFF_P__472  (.L_HI(net472));
 sg13g2_tiehi \i_vga.vblank$_DFF_P__473  (.L_HI(net473));
 sg13g2_tiehi \iter[0]$_SDFFCE_PP0N__474  (.L_HI(net474));
 sg13g2_tiehi \iter[1]$_SDFFCE_PP0N__475  (.L_HI(net475));
 sg13g2_tiehi \iter[2]$_SDFFCE_PP0N__476  (.L_HI(net476));
 sg13g2_tiehi \iter[3]$_SDFFCE_PP0N__477  (.L_HI(net477));
 sg13g2_tiehi \last_iter[0]$_DFFE_PP__478  (.L_HI(net478));
 sg13g2_tiehi \last_iter[1]$_DFFE_PP__479  (.L_HI(net479));
 sg13g2_tiehi \last_iter[2]$_DFFE_PP__480  (.L_HI(net480));
 sg13g2_tiehi \last_iter[3]$_DFFE_PP__481  (.L_HI(net481));
 sg13g2_tiehi \last_iter[4]$_DFFE_PP__482  (.L_HI(net482));
 sg13g2_tiehi \step[0]$_SDFF_PP0__483  (.L_HI(net483));
 sg13g2_tiehi \step[1]$_SDFF_PP0__484  (.L_HI(net484));
 sg13g2_tiehi \step[2]$_SDFF_PP0__485  (.L_HI(net485));
 sg13g2_tiehi \step[3]$_SDFF_PP0__486  (.L_HI(net486));
 sg13g2_tiehi \video_colour[0]$_SDFF_PP0__487  (.L_HI(net487));
 sg13g2_tiehi \video_colour[1]$_SDFF_PP0__488  (.L_HI(net488));
 sg13g2_tiehi \video_colour[2]$_SDFF_PP0__489  (.L_HI(net489));
 sg13g2_tiehi \video_colour[3]$_SDFF_PP0__490  (.L_HI(net490));
 sg13g2_tiehi \video_colour[4]$_SDFF_PP0__491  (.L_HI(net491));
 sg13g2_tiehi \video_colour[5]$_SDFF_PP0__492  (.L_HI(net492));
 sg13g2_tiehi \x0[0]$_DFFE_PP__493  (.L_HI(net493));
 sg13g2_tiehi \x0[10]$_DFFE_PP__494  (.L_HI(net494));
 sg13g2_tiehi \x0[11]$_DFFE_PP__495  (.L_HI(net495));
 sg13g2_tiehi \x0[12]$_DFFE_PP__496  (.L_HI(net496));
 sg13g2_tiehi \x0[13]$_DFFE_PP__497  (.L_HI(net497));
 sg13g2_tiehi \x0[14]$_DFFE_PP__498  (.L_HI(net498));
 sg13g2_tiehi \x0[15]$_DFFE_PP__499  (.L_HI(net499));
 sg13g2_tiehi \x0[1]$_DFFE_PP__500  (.L_HI(net500));
 sg13g2_tiehi \x0[2]$_DFFE_PP__501  (.L_HI(net501));
 sg13g2_tiehi \x0[3]$_DFFE_PP__502  (.L_HI(net502));
 sg13g2_tiehi \x0[4]$_DFFE_PP__503  (.L_HI(net503));
 sg13g2_tiehi \x0[5]$_DFFE_PP__504  (.L_HI(net504));
 sg13g2_tiehi \x0[6]$_DFFE_PP__505  (.L_HI(net505));
 sg13g2_tiehi \x0[7]$_DFFE_PP__506  (.L_HI(net506));
 sg13g2_tiehi \x0[8]$_DFFE_PP__507  (.L_HI(net507));
 sg13g2_tiehi \x0[9]$_DFFE_PP__508  (.L_HI(net508));
 sg13g2_tiehi \x[0]$_DFFE_PP__509  (.L_HI(net509));
 sg13g2_tiehi \x[10]$_DFFE_PP__510  (.L_HI(net510));
 sg13g2_tiehi \x[11]$_DFFE_PP__511  (.L_HI(net511));
 sg13g2_tiehi \x[12]$_DFFE_PP__512  (.L_HI(net512));
 sg13g2_tiehi \x[13]$_DFFE_PP__513  (.L_HI(net513));
 sg13g2_tiehi \x[14]$_DFFE_PP__514  (.L_HI(net514));
 sg13g2_tiehi \x[15]$_DFFE_PP__515  (.L_HI(net515));
 sg13g2_tiehi \x[1]$_DFFE_PP__516  (.L_HI(net516));
 sg13g2_tiehi \x[2]$_DFFE_PP__517  (.L_HI(net517));
 sg13g2_tiehi \x[3]$_DFFE_PP__518  (.L_HI(net518));
 sg13g2_tiehi \x[4]$_DFFE_PP__519  (.L_HI(net519));
 sg13g2_tiehi \x[5]$_DFFE_PP__520  (.L_HI(net520));
 sg13g2_tiehi \x[6]$_DFFE_PP__521  (.L_HI(net521));
 sg13g2_tiehi \x[7]$_DFFE_PP__522  (.L_HI(net522));
 sg13g2_tiehi \x[8]$_DFFE_PP__523  (.L_HI(net523));
 sg13g2_tiehi \x[9]$_DFFE_PP__524  (.L_HI(net524));
 sg13g2_tiehi \y0[0]$_DFFE_PP__525  (.L_HI(net525));
 sg13g2_tiehi \y0[10]$_DFFE_PP__526  (.L_HI(net526));
 sg13g2_tiehi \y0[11]$_DFFE_PP__527  (.L_HI(net527));
 sg13g2_tiehi \y0[12]$_DFFE_PP__528  (.L_HI(net528));
 sg13g2_tiehi \y0[13]$_DFFE_PP__529  (.L_HI(net529));
 sg13g2_tiehi \y0[14]$_DFFE_PP__530  (.L_HI(net530));
 sg13g2_tiehi \y0[1]$_DFFE_PP__531  (.L_HI(net531));
 sg13g2_tiehi \y0[2]$_DFFE_PP__532  (.L_HI(net532));
 sg13g2_tiehi \y0[3]$_DFFE_PP__533  (.L_HI(net533));
 sg13g2_tiehi \y0[4]$_DFFE_PP__534  (.L_HI(net534));
 sg13g2_tiehi \y0[5]$_DFFE_PP__535  (.L_HI(net535));
 sg13g2_tiehi \y0[6]$_DFFE_PP__536  (.L_HI(net536));
 sg13g2_tiehi \y0[7]$_DFFE_PP__537  (.L_HI(net537));
 sg13g2_tiehi \y0[8]$_DFFE_PP__538  (.L_HI(net538));
 sg13g2_tiehi \y0[9]$_DFFE_PP__539  (.L_HI(net539));
 sg13g2_tiehi \y[0]$_DFFE_PP__540  (.L_HI(net540));
 sg13g2_tiehi \y[10]$_DFFE_PP__541  (.L_HI(net541));
 sg13g2_tiehi \y[11]$_DFFE_PP__542  (.L_HI(net542));
 sg13g2_tiehi \y[12]$_DFFE_PP__543  (.L_HI(net543));
 sg13g2_tiehi \y[13]$_DFFE_PP__544  (.L_HI(net544));
 sg13g2_tiehi \y[14]$_DFFE_PP__545  (.L_HI(net545));
 sg13g2_tiehi \y[15]$_DFFE_PP__546  (.L_HI(net546));
 sg13g2_tiehi \y[1]$_DFFE_PP__547  (.L_HI(net547));
 sg13g2_tiehi \y[2]$_DFFE_PP__548  (.L_HI(net548));
 sg13g2_tiehi \y[3]$_DFFE_PP__549  (.L_HI(net549));
 sg13g2_tiehi \y[4]$_DFFE_PP__550  (.L_HI(net550));
 sg13g2_tiehi \y[5]$_DFFE_PP__551  (.L_HI(net551));
 sg13g2_tiehi \y[6]$_DFFE_PP__552  (.L_HI(net552));
 sg13g2_tiehi \y[7]$_DFFE_PP__553  (.L_HI(net553));
 sg13g2_tiehi \y[8]$_DFFE_PP__554  (.L_HI(net554));
 sg13g2_tiehi \y[9]$_DFFE_PP__555  (.L_HI(net555));
 sg13g2_buf_4 clkbuf_leaf_1_clk (.X(clknet_leaf_1_clk),
    .A(clknet_2_0__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_2_clk (.X(clknet_leaf_2_clk),
    .A(clknet_2_1__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_3_clk (.X(clknet_leaf_3_clk),
    .A(clknet_2_1__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_4_clk (.X(clknet_leaf_4_clk),
    .A(clknet_2_1__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_5_clk (.X(clknet_leaf_5_clk),
    .A(clknet_2_1__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_6_clk (.X(clknet_leaf_6_clk),
    .A(clknet_2_0__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_7_clk (.X(clknet_leaf_7_clk),
    .A(clknet_2_0__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_8_clk (.X(clknet_leaf_8_clk),
    .A(clknet_2_0__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_9_clk (.X(clknet_leaf_9_clk),
    .A(clknet_2_0__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_10_clk (.X(clknet_leaf_10_clk),
    .A(clknet_2_0__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_11_clk (.X(clknet_leaf_11_clk),
    .A(clknet_2_2__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_12_clk (.X(clknet_leaf_12_clk),
    .A(clknet_2_2__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_13_clk (.X(clknet_leaf_13_clk),
    .A(clknet_2_2__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_14_clk (.X(clknet_leaf_14_clk),
    .A(clknet_2_3__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_15_clk (.X(clknet_leaf_15_clk),
    .A(clknet_2_2__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_16_clk (.X(clknet_leaf_16_clk),
    .A(clknet_2_3__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_17_clk (.X(clknet_leaf_17_clk),
    .A(clknet_2_3__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_18_clk (.X(clknet_leaf_18_clk),
    .A(clknet_2_3__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_19_clk (.X(clknet_leaf_19_clk),
    .A(clknet_2_3__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_20_clk (.X(clknet_leaf_20_clk),
    .A(clknet_2_3__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_21_clk (.X(clknet_leaf_21_clk),
    .A(clknet_2_2__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_22_clk (.X(clknet_leaf_22_clk),
    .A(clknet_2_2__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_23_clk (.X(clknet_leaf_23_clk),
    .A(clknet_2_2__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_24_clk (.X(clknet_leaf_24_clk),
    .A(clknet_2_0__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_25_clk (.X(clknet_leaf_25_clk),
    .A(clknet_2_1__leaf_clk));
 sg13g2_buf_2 clkbuf_0_clk (.A(clk),
    .X(clknet_0_clk));
 sg13g2_buf_2 clkbuf_2_0__f_clk (.A(clknet_0_clk),
    .X(clknet_2_0__leaf_clk));
 sg13g2_buf_2 clkbuf_2_1__f_clk (.A(clknet_0_clk),
    .X(clknet_2_1__leaf_clk));
 sg13g2_buf_2 clkbuf_2_2__f_clk (.A(clknet_0_clk),
    .X(clknet_2_2__leaf_clk));
 sg13g2_buf_2 clkbuf_2_3__f_clk (.A(clknet_0_clk),
    .X(clknet_2_3__leaf_clk));
 sg13g2_buf_4 clkload0 (.A(clknet_2_1__leaf_clk));
 sg13g2_buf_4 clkload1 (.A(clknet_2_3__leaf_clk));
 sg13g2_buf_16 clkload2 (.A(clknet_leaf_25_clk));
 sg13g2_antennanp ANTENNA_1 (.A(_00198_));
 sg13g2_antennanp ANTENNA_2 (.A(_00199_));
 sg13g2_antennanp ANTENNA_3 (.A(_00225_));
 sg13g2_antennanp ANTENNA_4 (.A(_00225_));
 sg13g2_antennanp ANTENNA_5 (.A(_00227_));
 sg13g2_antennanp ANTENNA_6 (.A(_00228_));
 sg13g2_antennanp ANTENNA_7 (.A(_00228_));
 sg13g2_antennanp ANTENNA_8 (.A(_00229_));
 sg13g2_antennanp ANTENNA_9 (.A(_00229_));
 sg13g2_antennanp ANTENNA_10 (.A(_00230_));
 sg13g2_antennanp ANTENNA_11 (.A(_00238_));
 sg13g2_antennanp ANTENNA_12 (.A(_00239_));
 sg13g2_antennanp ANTENNA_13 (.A(_03588_));
 sg13g2_antennanp ANTENNA_14 (.A(_03588_));
 sg13g2_antennanp ANTENNA_15 (.A(_03621_));
 sg13g2_antennanp ANTENNA_16 (.A(_03621_));
 sg13g2_antennanp ANTENNA_17 (.A(_03635_));
 sg13g2_antennanp ANTENNA_18 (.A(_03635_));
 sg13g2_antennanp ANTENNA_19 (.A(_03677_));
 sg13g2_antennanp ANTENNA_20 (.A(_03677_));
 sg13g2_antennanp ANTENNA_21 (.A(_04990_));
 sg13g2_antennanp ANTENNA_22 (.A(_05003_));
 sg13g2_antennanp ANTENNA_23 (.A(_05007_));
 sg13g2_antennanp ANTENNA_24 (.A(net102));
 sg13g2_antennanp ANTENNA_25 (.A(net102));
 sg13g2_antennanp ANTENNA_26 (.A(net102));
 sg13g2_antennanp ANTENNA_27 (.A(net102));
 sg13g2_antennanp ANTENNA_28 (.A(net102));
 sg13g2_antennanp ANTENNA_29 (.A(net102));
 sg13g2_antennanp ANTENNA_30 (.A(net102));
 sg13g2_antennanp ANTENNA_31 (.A(net102));
 sg13g2_antennanp ANTENNA_32 (.A(net102));
 sg13g2_antennanp ANTENNA_33 (.A(net102));
 sg13g2_antennanp ANTENNA_34 (.A(net102));
 sg13g2_antennanp ANTENNA_35 (.A(net102));
 sg13g2_antennanp ANTENNA_36 (.A(net102));
 sg13g2_antennanp ANTENNA_37 (.A(net102));
 sg13g2_antennanp ANTENNA_38 (.A(net102));
 sg13g2_antennanp ANTENNA_39 (.A(_00198_));
 sg13g2_antennanp ANTENNA_40 (.A(_00199_));
 sg13g2_antennanp ANTENNA_41 (.A(_00225_));
 sg13g2_antennanp ANTENNA_42 (.A(_00225_));
 sg13g2_antennanp ANTENNA_43 (.A(_00227_));
 sg13g2_antennanp ANTENNA_44 (.A(_00228_));
 sg13g2_antennanp ANTENNA_45 (.A(_00228_));
 sg13g2_antennanp ANTENNA_46 (.A(_00229_));
 sg13g2_antennanp ANTENNA_47 (.A(_00230_));
 sg13g2_antennanp ANTENNA_48 (.A(_00238_));
 sg13g2_antennanp ANTENNA_49 (.A(_03635_));
 sg13g2_antennanp ANTENNA_50 (.A(_03635_));
 sg13g2_antennanp ANTENNA_51 (.A(_03677_));
 sg13g2_antennanp ANTENNA_52 (.A(_03677_));
 sg13g2_antennanp ANTENNA_53 (.A(_04990_));
 sg13g2_antennanp ANTENNA_54 (.A(_05003_));
 sg13g2_antennanp ANTENNA_55 (.A(_05007_));
 sg13g2_antennanp ANTENNA_56 (.A(_00198_));
 sg13g2_antennanp ANTENNA_57 (.A(_00199_));
 sg13g2_antennanp ANTENNA_58 (.A(_00225_));
 sg13g2_antennanp ANTENNA_59 (.A(_00227_));
 sg13g2_antennanp ANTENNA_60 (.A(_00228_));
 sg13g2_antennanp ANTENNA_61 (.A(_00229_));
 sg13g2_antennanp ANTENNA_62 (.A(_00230_));
 sg13g2_antennanp ANTENNA_63 (.A(_03677_));
 sg13g2_antennanp ANTENNA_64 (.A(_03677_));
 sg13g2_antennanp ANTENNA_65 (.A(_04990_));
 sg13g2_antennanp ANTENNA_66 (.A(_05007_));
 sg13g2_antennanp ANTENNA_67 (.A(_00198_));
 sg13g2_antennanp ANTENNA_68 (.A(_00199_));
 sg13g2_antennanp ANTENNA_69 (.A(_00225_));
 sg13g2_antennanp ANTENNA_70 (.A(_00227_));
 sg13g2_antennanp ANTENNA_71 (.A(_00228_));
 sg13g2_antennanp ANTENNA_72 (.A(_00229_));
 sg13g2_antennanp ANTENNA_73 (.A(_03677_));
 sg13g2_antennanp ANTENNA_74 (.A(_03677_));
 sg13g2_antennanp ANTENNA_75 (.A(_04990_));
 sg13g2_antennanp ANTENNA_76 (.A(_05007_));
 sg13g2_antennanp ANTENNA_77 (.A(_00198_));
 sg13g2_antennanp ANTENNA_78 (.A(_00199_));
 sg13g2_antennanp ANTENNA_79 (.A(_00225_));
 sg13g2_antennanp ANTENNA_80 (.A(_00227_));
 sg13g2_antennanp ANTENNA_81 (.A(_00228_));
 sg13g2_antennanp ANTENNA_82 (.A(_00229_));
 sg13g2_antennanp ANTENNA_83 (.A(_03677_));
 sg13g2_antennanp ANTENNA_84 (.A(_03677_));
 sg13g2_antennanp ANTENNA_85 (.A(_04990_));
 sg13g2_antennanp ANTENNA_86 (.A(_05007_));
 sg13g2_decap_8 FILLER_0_0 ();
 sg13g2_decap_8 FILLER_0_7 ();
 sg13g2_decap_8 FILLER_0_14 ();
 sg13g2_decap_8 FILLER_0_21 ();
 sg13g2_decap_8 FILLER_0_28 ();
 sg13g2_decap_8 FILLER_0_35 ();
 sg13g2_decap_8 FILLER_0_42 ();
 sg13g2_decap_8 FILLER_0_49 ();
 sg13g2_decap_8 FILLER_0_56 ();
 sg13g2_decap_8 FILLER_0_63 ();
 sg13g2_decap_8 FILLER_0_70 ();
 sg13g2_decap_8 FILLER_0_77 ();
 sg13g2_decap_8 FILLER_0_84 ();
 sg13g2_decap_8 FILLER_0_91 ();
 sg13g2_decap_8 FILLER_0_98 ();
 sg13g2_decap_8 FILLER_0_105 ();
 sg13g2_decap_8 FILLER_0_112 ();
 sg13g2_decap_8 FILLER_0_119 ();
 sg13g2_decap_8 FILLER_0_126 ();
 sg13g2_decap_8 FILLER_0_133 ();
 sg13g2_decap_8 FILLER_0_140 ();
 sg13g2_decap_8 FILLER_0_147 ();
 sg13g2_decap_8 FILLER_0_154 ();
 sg13g2_decap_8 FILLER_0_161 ();
 sg13g2_decap_8 FILLER_0_168 ();
 sg13g2_decap_8 FILLER_0_175 ();
 sg13g2_decap_8 FILLER_0_182 ();
 sg13g2_decap_8 FILLER_0_189 ();
 sg13g2_decap_8 FILLER_0_196 ();
 sg13g2_decap_8 FILLER_0_203 ();
 sg13g2_decap_8 FILLER_0_210 ();
 sg13g2_decap_8 FILLER_0_217 ();
 sg13g2_decap_8 FILLER_0_224 ();
 sg13g2_decap_8 FILLER_0_231 ();
 sg13g2_decap_8 FILLER_0_238 ();
 sg13g2_decap_8 FILLER_0_245 ();
 sg13g2_decap_8 FILLER_0_252 ();
 sg13g2_decap_8 FILLER_0_259 ();
 sg13g2_decap_8 FILLER_0_266 ();
 sg13g2_decap_8 FILLER_0_273 ();
 sg13g2_decap_8 FILLER_0_280 ();
 sg13g2_decap_8 FILLER_0_287 ();
 sg13g2_decap_8 FILLER_0_294 ();
 sg13g2_decap_8 FILLER_0_301 ();
 sg13g2_decap_8 FILLER_0_308 ();
 sg13g2_decap_8 FILLER_0_315 ();
 sg13g2_decap_8 FILLER_0_322 ();
 sg13g2_decap_8 FILLER_0_329 ();
 sg13g2_decap_8 FILLER_0_336 ();
 sg13g2_decap_8 FILLER_0_343 ();
 sg13g2_decap_8 FILLER_0_350 ();
 sg13g2_fill_1 FILLER_0_357 ();
 sg13g2_fill_2 FILLER_0_363 ();
 sg13g2_decap_4 FILLER_0_370 ();
 sg13g2_fill_2 FILLER_0_374 ();
 sg13g2_decap_8 FILLER_0_381 ();
 sg13g2_fill_2 FILLER_0_388 ();
 sg13g2_decap_8 FILLER_0_396 ();
 sg13g2_decap_8 FILLER_0_403 ();
 sg13g2_decap_8 FILLER_0_410 ();
 sg13g2_decap_8 FILLER_0_417 ();
 sg13g2_decap_8 FILLER_0_424 ();
 sg13g2_decap_4 FILLER_0_431 ();
 sg13g2_fill_2 FILLER_0_435 ();
 sg13g2_fill_2 FILLER_0_451 ();
 sg13g2_fill_1 FILLER_0_453 ();
 sg13g2_decap_4 FILLER_0_467 ();
 sg13g2_fill_2 FILLER_0_471 ();
 sg13g2_decap_8 FILLER_0_478 ();
 sg13g2_decap_4 FILLER_0_485 ();
 sg13g2_fill_1 FILLER_0_499 ();
 sg13g2_decap_8 FILLER_0_507 ();
 sg13g2_decap_8 FILLER_0_514 ();
 sg13g2_decap_8 FILLER_0_521 ();
 sg13g2_decap_8 FILLER_0_528 ();
 sg13g2_decap_8 FILLER_0_535 ();
 sg13g2_decap_8 FILLER_0_542 ();
 sg13g2_decap_8 FILLER_0_549 ();
 sg13g2_decap_8 FILLER_0_556 ();
 sg13g2_decap_8 FILLER_0_563 ();
 sg13g2_decap_8 FILLER_0_570 ();
 sg13g2_decap_8 FILLER_0_577 ();
 sg13g2_decap_8 FILLER_0_584 ();
 sg13g2_decap_8 FILLER_0_591 ();
 sg13g2_decap_8 FILLER_0_598 ();
 sg13g2_decap_8 FILLER_0_605 ();
 sg13g2_decap_8 FILLER_0_612 ();
 sg13g2_decap_8 FILLER_0_619 ();
 sg13g2_decap_8 FILLER_0_626 ();
 sg13g2_decap_8 FILLER_0_633 ();
 sg13g2_decap_8 FILLER_0_640 ();
 sg13g2_decap_8 FILLER_0_647 ();
 sg13g2_decap_8 FILLER_0_654 ();
 sg13g2_decap_8 FILLER_0_661 ();
 sg13g2_decap_8 FILLER_0_668 ();
 sg13g2_decap_8 FILLER_0_675 ();
 sg13g2_decap_8 FILLER_0_682 ();
 sg13g2_decap_8 FILLER_0_689 ();
 sg13g2_decap_8 FILLER_0_696 ();
 sg13g2_decap_8 FILLER_0_703 ();
 sg13g2_decap_8 FILLER_0_710 ();
 sg13g2_decap_8 FILLER_0_717 ();
 sg13g2_decap_8 FILLER_0_724 ();
 sg13g2_decap_8 FILLER_0_731 ();
 sg13g2_decap_8 FILLER_0_738 ();
 sg13g2_decap_8 FILLER_0_745 ();
 sg13g2_decap_8 FILLER_0_752 ();
 sg13g2_decap_8 FILLER_0_759 ();
 sg13g2_decap_8 FILLER_0_766 ();
 sg13g2_decap_8 FILLER_0_773 ();
 sg13g2_decap_8 FILLER_0_780 ();
 sg13g2_decap_8 FILLER_0_787 ();
 sg13g2_decap_8 FILLER_0_794 ();
 sg13g2_decap_8 FILLER_0_801 ();
 sg13g2_decap_8 FILLER_0_808 ();
 sg13g2_decap_8 FILLER_0_815 ();
 sg13g2_decap_8 FILLER_0_822 ();
 sg13g2_decap_8 FILLER_0_829 ();
 sg13g2_decap_8 FILLER_0_836 ();
 sg13g2_decap_8 FILLER_0_843 ();
 sg13g2_decap_8 FILLER_0_850 ();
 sg13g2_decap_8 FILLER_0_857 ();
 sg13g2_decap_8 FILLER_0_864 ();
 sg13g2_decap_8 FILLER_0_871 ();
 sg13g2_decap_8 FILLER_1_0 ();
 sg13g2_decap_8 FILLER_1_7 ();
 sg13g2_decap_8 FILLER_1_14 ();
 sg13g2_decap_8 FILLER_1_21 ();
 sg13g2_decap_8 FILLER_1_28 ();
 sg13g2_decap_8 FILLER_1_35 ();
 sg13g2_decap_8 FILLER_1_42 ();
 sg13g2_decap_8 FILLER_1_49 ();
 sg13g2_decap_8 FILLER_1_56 ();
 sg13g2_decap_8 FILLER_1_63 ();
 sg13g2_decap_8 FILLER_1_70 ();
 sg13g2_decap_8 FILLER_1_77 ();
 sg13g2_decap_8 FILLER_1_84 ();
 sg13g2_decap_8 FILLER_1_91 ();
 sg13g2_decap_8 FILLER_1_98 ();
 sg13g2_decap_8 FILLER_1_105 ();
 sg13g2_decap_8 FILLER_1_112 ();
 sg13g2_decap_8 FILLER_1_119 ();
 sg13g2_decap_8 FILLER_1_126 ();
 sg13g2_decap_8 FILLER_1_133 ();
 sg13g2_decap_8 FILLER_1_140 ();
 sg13g2_decap_8 FILLER_1_147 ();
 sg13g2_decap_8 FILLER_1_154 ();
 sg13g2_decap_8 FILLER_1_161 ();
 sg13g2_decap_8 FILLER_1_168 ();
 sg13g2_decap_8 FILLER_1_175 ();
 sg13g2_decap_8 FILLER_1_182 ();
 sg13g2_decap_8 FILLER_1_189 ();
 sg13g2_decap_8 FILLER_1_196 ();
 sg13g2_decap_4 FILLER_1_203 ();
 sg13g2_fill_1 FILLER_1_211 ();
 sg13g2_decap_8 FILLER_1_221 ();
 sg13g2_decap_8 FILLER_1_228 ();
 sg13g2_decap_4 FILLER_1_235 ();
 sg13g2_decap_4 FILLER_1_245 ();
 sg13g2_decap_8 FILLER_1_254 ();
 sg13g2_fill_2 FILLER_1_261 ();
 sg13g2_fill_2 FILLER_1_276 ();
 sg13g2_decap_8 FILLER_1_285 ();
 sg13g2_decap_8 FILLER_1_292 ();
 sg13g2_decap_8 FILLER_1_299 ();
 sg13g2_decap_8 FILLER_1_306 ();
 sg13g2_decap_4 FILLER_1_313 ();
 sg13g2_fill_2 FILLER_1_317 ();
 sg13g2_decap_8 FILLER_1_323 ();
 sg13g2_fill_2 FILLER_1_330 ();
 sg13g2_decap_4 FILLER_1_337 ();
 sg13g2_fill_1 FILLER_1_341 ();
 sg13g2_fill_2 FILLER_1_375 ();
 sg13g2_fill_1 FILLER_1_377 ();
 sg13g2_decap_4 FILLER_1_388 ();
 sg13g2_decap_8 FILLER_1_412 ();
 sg13g2_decap_8 FILLER_1_419 ();
 sg13g2_decap_8 FILLER_1_426 ();
 sg13g2_fill_1 FILLER_1_453 ();
 sg13g2_fill_1 FILLER_1_473 ();
 sg13g2_decap_4 FILLER_1_493 ();
 sg13g2_decap_8 FILLER_1_504 ();
 sg13g2_decap_8 FILLER_1_511 ();
 sg13g2_decap_4 FILLER_1_518 ();
 sg13g2_fill_1 FILLER_1_522 ();
 sg13g2_decap_8 FILLER_1_531 ();
 sg13g2_decap_8 FILLER_1_538 ();
 sg13g2_decap_8 FILLER_1_545 ();
 sg13g2_decap_8 FILLER_1_552 ();
 sg13g2_decap_8 FILLER_1_559 ();
 sg13g2_decap_8 FILLER_1_566 ();
 sg13g2_decap_8 FILLER_1_573 ();
 sg13g2_decap_8 FILLER_1_580 ();
 sg13g2_decap_8 FILLER_1_587 ();
 sg13g2_decap_8 FILLER_1_594 ();
 sg13g2_decap_8 FILLER_1_601 ();
 sg13g2_decap_8 FILLER_1_608 ();
 sg13g2_decap_8 FILLER_1_615 ();
 sg13g2_decap_8 FILLER_1_622 ();
 sg13g2_decap_8 FILLER_1_629 ();
 sg13g2_decap_8 FILLER_1_636 ();
 sg13g2_decap_8 FILLER_1_643 ();
 sg13g2_decap_8 FILLER_1_650 ();
 sg13g2_decap_8 FILLER_1_657 ();
 sg13g2_decap_8 FILLER_1_664 ();
 sg13g2_decap_8 FILLER_1_671 ();
 sg13g2_decap_8 FILLER_1_678 ();
 sg13g2_decap_8 FILLER_1_685 ();
 sg13g2_decap_8 FILLER_1_692 ();
 sg13g2_decap_8 FILLER_1_699 ();
 sg13g2_decap_8 FILLER_1_706 ();
 sg13g2_decap_8 FILLER_1_713 ();
 sg13g2_decap_8 FILLER_1_720 ();
 sg13g2_decap_8 FILLER_1_727 ();
 sg13g2_decap_8 FILLER_1_734 ();
 sg13g2_decap_8 FILLER_1_741 ();
 sg13g2_decap_8 FILLER_1_748 ();
 sg13g2_decap_8 FILLER_1_755 ();
 sg13g2_decap_8 FILLER_1_762 ();
 sg13g2_decap_8 FILLER_1_769 ();
 sg13g2_decap_8 FILLER_1_776 ();
 sg13g2_decap_8 FILLER_1_783 ();
 sg13g2_decap_8 FILLER_1_790 ();
 sg13g2_decap_8 FILLER_1_797 ();
 sg13g2_decap_8 FILLER_1_804 ();
 sg13g2_decap_8 FILLER_1_811 ();
 sg13g2_decap_8 FILLER_1_818 ();
 sg13g2_decap_8 FILLER_1_825 ();
 sg13g2_decap_8 FILLER_1_832 ();
 sg13g2_decap_8 FILLER_1_839 ();
 sg13g2_decap_8 FILLER_1_846 ();
 sg13g2_decap_8 FILLER_1_853 ();
 sg13g2_decap_8 FILLER_1_860 ();
 sg13g2_decap_8 FILLER_1_867 ();
 sg13g2_decap_4 FILLER_1_874 ();
 sg13g2_decap_8 FILLER_2_0 ();
 sg13g2_decap_8 FILLER_2_7 ();
 sg13g2_decap_8 FILLER_2_14 ();
 sg13g2_decap_8 FILLER_2_21 ();
 sg13g2_decap_8 FILLER_2_28 ();
 sg13g2_decap_8 FILLER_2_35 ();
 sg13g2_decap_8 FILLER_2_42 ();
 sg13g2_decap_8 FILLER_2_49 ();
 sg13g2_decap_8 FILLER_2_56 ();
 sg13g2_decap_8 FILLER_2_63 ();
 sg13g2_decap_8 FILLER_2_70 ();
 sg13g2_decap_8 FILLER_2_77 ();
 sg13g2_decap_8 FILLER_2_84 ();
 sg13g2_decap_8 FILLER_2_91 ();
 sg13g2_decap_8 FILLER_2_98 ();
 sg13g2_decap_8 FILLER_2_105 ();
 sg13g2_decap_8 FILLER_2_112 ();
 sg13g2_decap_8 FILLER_2_119 ();
 sg13g2_decap_8 FILLER_2_126 ();
 sg13g2_decap_8 FILLER_2_133 ();
 sg13g2_fill_2 FILLER_2_140 ();
 sg13g2_fill_1 FILLER_2_142 ();
 sg13g2_decap_4 FILLER_2_151 ();
 sg13g2_fill_2 FILLER_2_160 ();
 sg13g2_fill_1 FILLER_2_162 ();
 sg13g2_decap_8 FILLER_2_179 ();
 sg13g2_decap_8 FILLER_2_186 ();
 sg13g2_fill_1 FILLER_2_193 ();
 sg13g2_decap_4 FILLER_2_198 ();
 sg13g2_fill_1 FILLER_2_207 ();
 sg13g2_fill_2 FILLER_2_227 ();
 sg13g2_fill_1 FILLER_2_229 ();
 sg13g2_fill_2 FILLER_2_260 ();
 sg13g2_fill_1 FILLER_2_262 ();
 sg13g2_decap_8 FILLER_2_282 ();
 sg13g2_decap_8 FILLER_2_289 ();
 sg13g2_decap_8 FILLER_2_296 ();
 sg13g2_decap_4 FILLER_2_303 ();
 sg13g2_fill_1 FILLER_2_307 ();
 sg13g2_decap_4 FILLER_2_313 ();
 sg13g2_fill_1 FILLER_2_317 ();
 sg13g2_decap_8 FILLER_2_323 ();
 sg13g2_decap_8 FILLER_2_330 ();
 sg13g2_fill_2 FILLER_2_337 ();
 sg13g2_fill_1 FILLER_2_339 ();
 sg13g2_fill_2 FILLER_2_371 ();
 sg13g2_fill_2 FILLER_2_377 ();
 sg13g2_fill_2 FILLER_2_384 ();
 sg13g2_fill_2 FILLER_2_390 ();
 sg13g2_fill_1 FILLER_2_392 ();
 sg13g2_fill_1 FILLER_2_402 ();
 sg13g2_decap_8 FILLER_2_408 ();
 sg13g2_decap_4 FILLER_2_415 ();
 sg13g2_fill_2 FILLER_2_419 ();
 sg13g2_fill_1 FILLER_2_445 ();
 sg13g2_fill_2 FILLER_2_466 ();
 sg13g2_fill_1 FILLER_2_486 ();
 sg13g2_fill_1 FILLER_2_501 ();
 sg13g2_decap_8 FILLER_2_506 ();
 sg13g2_decap_4 FILLER_2_513 ();
 sg13g2_decap_8 FILLER_2_537 ();
 sg13g2_decap_8 FILLER_2_544 ();
 sg13g2_decap_8 FILLER_2_551 ();
 sg13g2_decap_8 FILLER_2_558 ();
 sg13g2_decap_8 FILLER_2_565 ();
 sg13g2_decap_8 FILLER_2_572 ();
 sg13g2_decap_8 FILLER_2_579 ();
 sg13g2_decap_8 FILLER_2_586 ();
 sg13g2_decap_8 FILLER_2_593 ();
 sg13g2_decap_8 FILLER_2_600 ();
 sg13g2_decap_8 FILLER_2_607 ();
 sg13g2_decap_8 FILLER_2_614 ();
 sg13g2_decap_8 FILLER_2_621 ();
 sg13g2_decap_8 FILLER_2_628 ();
 sg13g2_decap_8 FILLER_2_635 ();
 sg13g2_decap_8 FILLER_2_642 ();
 sg13g2_decap_8 FILLER_2_649 ();
 sg13g2_decap_8 FILLER_2_656 ();
 sg13g2_decap_8 FILLER_2_663 ();
 sg13g2_decap_8 FILLER_2_670 ();
 sg13g2_decap_8 FILLER_2_677 ();
 sg13g2_decap_8 FILLER_2_684 ();
 sg13g2_decap_8 FILLER_2_691 ();
 sg13g2_decap_8 FILLER_2_698 ();
 sg13g2_decap_8 FILLER_2_705 ();
 sg13g2_decap_8 FILLER_2_712 ();
 sg13g2_decap_8 FILLER_2_719 ();
 sg13g2_decap_8 FILLER_2_726 ();
 sg13g2_decap_8 FILLER_2_733 ();
 sg13g2_decap_8 FILLER_2_740 ();
 sg13g2_decap_8 FILLER_2_747 ();
 sg13g2_decap_8 FILLER_2_754 ();
 sg13g2_decap_8 FILLER_2_761 ();
 sg13g2_decap_8 FILLER_2_768 ();
 sg13g2_decap_8 FILLER_2_775 ();
 sg13g2_decap_8 FILLER_2_782 ();
 sg13g2_decap_8 FILLER_2_789 ();
 sg13g2_decap_8 FILLER_2_796 ();
 sg13g2_decap_8 FILLER_2_803 ();
 sg13g2_decap_8 FILLER_2_810 ();
 sg13g2_decap_8 FILLER_2_817 ();
 sg13g2_decap_8 FILLER_2_824 ();
 sg13g2_decap_8 FILLER_2_831 ();
 sg13g2_decap_8 FILLER_2_838 ();
 sg13g2_decap_8 FILLER_2_845 ();
 sg13g2_decap_8 FILLER_2_852 ();
 sg13g2_decap_8 FILLER_2_859 ();
 sg13g2_decap_8 FILLER_2_866 ();
 sg13g2_decap_4 FILLER_2_873 ();
 sg13g2_fill_1 FILLER_2_877 ();
 sg13g2_decap_8 FILLER_3_0 ();
 sg13g2_decap_8 FILLER_3_7 ();
 sg13g2_decap_8 FILLER_3_14 ();
 sg13g2_decap_8 FILLER_3_21 ();
 sg13g2_decap_8 FILLER_3_28 ();
 sg13g2_decap_8 FILLER_3_35 ();
 sg13g2_decap_8 FILLER_3_42 ();
 sg13g2_decap_8 FILLER_3_49 ();
 sg13g2_decap_8 FILLER_3_56 ();
 sg13g2_decap_8 FILLER_3_63 ();
 sg13g2_decap_8 FILLER_3_70 ();
 sg13g2_decap_8 FILLER_3_77 ();
 sg13g2_decap_8 FILLER_3_84 ();
 sg13g2_decap_8 FILLER_3_91 ();
 sg13g2_decap_8 FILLER_3_98 ();
 sg13g2_decap_8 FILLER_3_105 ();
 sg13g2_decap_8 FILLER_3_112 ();
 sg13g2_decap_8 FILLER_3_119 ();
 sg13g2_decap_8 FILLER_3_126 ();
 sg13g2_fill_2 FILLER_3_133 ();
 sg13g2_decap_4 FILLER_3_139 ();
 sg13g2_fill_1 FILLER_3_143 ();
 sg13g2_fill_2 FILLER_3_152 ();
 sg13g2_fill_1 FILLER_3_154 ();
 sg13g2_fill_1 FILLER_3_159 ();
 sg13g2_fill_2 FILLER_3_169 ();
 sg13g2_decap_4 FILLER_3_193 ();
 sg13g2_decap_8 FILLER_3_205 ();
 sg13g2_decap_8 FILLER_3_212 ();
 sg13g2_fill_2 FILLER_3_219 ();
 sg13g2_fill_1 FILLER_3_221 ();
 sg13g2_fill_1 FILLER_3_238 ();
 sg13g2_fill_2 FILLER_3_253 ();
 sg13g2_fill_1 FILLER_3_255 ();
 sg13g2_decap_8 FILLER_3_277 ();
 sg13g2_fill_1 FILLER_3_284 ();
 sg13g2_decap_8 FILLER_3_291 ();
 sg13g2_decap_8 FILLER_3_298 ();
 sg13g2_decap_8 FILLER_3_305 ();
 sg13g2_fill_2 FILLER_3_312 ();
 sg13g2_fill_1 FILLER_3_314 ();
 sg13g2_decap_8 FILLER_3_329 ();
 sg13g2_decap_4 FILLER_3_336 ();
 sg13g2_fill_2 FILLER_3_350 ();
 sg13g2_fill_1 FILLER_3_356 ();
 sg13g2_fill_2 FILLER_3_367 ();
 sg13g2_fill_2 FILLER_3_383 ();
 sg13g2_fill_1 FILLER_3_385 ();
 sg13g2_fill_1 FILLER_3_433 ();
 sg13g2_fill_1 FILLER_3_438 ();
 sg13g2_fill_2 FILLER_3_443 ();
 sg13g2_fill_1 FILLER_3_445 ();
 sg13g2_decap_4 FILLER_3_469 ();
 sg13g2_fill_2 FILLER_3_487 ();
 sg13g2_fill_1 FILLER_3_489 ();
 sg13g2_fill_2 FILLER_3_496 ();
 sg13g2_fill_1 FILLER_3_502 ();
 sg13g2_fill_2 FILLER_3_507 ();
 sg13g2_decap_4 FILLER_3_518 ();
 sg13g2_fill_1 FILLER_3_531 ();
 sg13g2_decap_8 FILLER_3_542 ();
 sg13g2_decap_8 FILLER_3_549 ();
 sg13g2_decap_8 FILLER_3_556 ();
 sg13g2_decap_8 FILLER_3_563 ();
 sg13g2_decap_8 FILLER_3_570 ();
 sg13g2_decap_8 FILLER_3_577 ();
 sg13g2_decap_8 FILLER_3_584 ();
 sg13g2_decap_8 FILLER_3_591 ();
 sg13g2_decap_8 FILLER_3_598 ();
 sg13g2_decap_8 FILLER_3_605 ();
 sg13g2_decap_8 FILLER_3_612 ();
 sg13g2_decap_8 FILLER_3_619 ();
 sg13g2_decap_8 FILLER_3_626 ();
 sg13g2_decap_8 FILLER_3_633 ();
 sg13g2_decap_8 FILLER_3_640 ();
 sg13g2_decap_8 FILLER_3_647 ();
 sg13g2_decap_8 FILLER_3_654 ();
 sg13g2_decap_8 FILLER_3_661 ();
 sg13g2_decap_8 FILLER_3_668 ();
 sg13g2_decap_8 FILLER_3_675 ();
 sg13g2_decap_8 FILLER_3_682 ();
 sg13g2_decap_8 FILLER_3_689 ();
 sg13g2_decap_8 FILLER_3_696 ();
 sg13g2_decap_8 FILLER_3_703 ();
 sg13g2_decap_8 FILLER_3_710 ();
 sg13g2_decap_8 FILLER_3_717 ();
 sg13g2_decap_8 FILLER_3_724 ();
 sg13g2_decap_8 FILLER_3_731 ();
 sg13g2_decap_8 FILLER_3_738 ();
 sg13g2_decap_8 FILLER_3_745 ();
 sg13g2_decap_8 FILLER_3_752 ();
 sg13g2_decap_8 FILLER_3_759 ();
 sg13g2_decap_8 FILLER_3_766 ();
 sg13g2_decap_8 FILLER_3_773 ();
 sg13g2_decap_8 FILLER_3_780 ();
 sg13g2_decap_8 FILLER_3_787 ();
 sg13g2_decap_8 FILLER_3_794 ();
 sg13g2_decap_8 FILLER_3_801 ();
 sg13g2_decap_8 FILLER_3_808 ();
 sg13g2_decap_8 FILLER_3_815 ();
 sg13g2_decap_8 FILLER_3_822 ();
 sg13g2_decap_8 FILLER_3_829 ();
 sg13g2_decap_8 FILLER_3_836 ();
 sg13g2_decap_8 FILLER_3_843 ();
 sg13g2_decap_8 FILLER_3_850 ();
 sg13g2_decap_8 FILLER_3_857 ();
 sg13g2_decap_8 FILLER_3_864 ();
 sg13g2_decap_8 FILLER_3_871 ();
 sg13g2_decap_8 FILLER_4_0 ();
 sg13g2_decap_8 FILLER_4_7 ();
 sg13g2_decap_8 FILLER_4_14 ();
 sg13g2_decap_8 FILLER_4_21 ();
 sg13g2_decap_8 FILLER_4_28 ();
 sg13g2_decap_8 FILLER_4_35 ();
 sg13g2_decap_8 FILLER_4_42 ();
 sg13g2_decap_8 FILLER_4_49 ();
 sg13g2_decap_8 FILLER_4_56 ();
 sg13g2_decap_8 FILLER_4_63 ();
 sg13g2_decap_8 FILLER_4_70 ();
 sg13g2_decap_8 FILLER_4_77 ();
 sg13g2_decap_8 FILLER_4_84 ();
 sg13g2_decap_8 FILLER_4_91 ();
 sg13g2_fill_1 FILLER_4_98 ();
 sg13g2_fill_1 FILLER_4_107 ();
 sg13g2_fill_2 FILLER_4_124 ();
 sg13g2_decap_4 FILLER_4_143 ();
 sg13g2_fill_2 FILLER_4_159 ();
 sg13g2_decap_4 FILLER_4_174 ();
 sg13g2_fill_1 FILLER_4_178 ();
 sg13g2_fill_1 FILLER_4_196 ();
 sg13g2_decap_4 FILLER_4_201 ();
 sg13g2_fill_1 FILLER_4_205 ();
 sg13g2_decap_8 FILLER_4_211 ();
 sg13g2_fill_1 FILLER_4_218 ();
 sg13g2_fill_1 FILLER_4_233 ();
 sg13g2_decap_8 FILLER_4_250 ();
 sg13g2_fill_1 FILLER_4_257 ();
 sg13g2_fill_1 FILLER_4_264 ();
 sg13g2_decap_4 FILLER_4_280 ();
 sg13g2_fill_2 FILLER_4_284 ();
 sg13g2_fill_1 FILLER_4_316 ();
 sg13g2_decap_4 FILLER_4_354 ();
 sg13g2_fill_1 FILLER_4_358 ();
 sg13g2_decap_8 FILLER_4_363 ();
 sg13g2_fill_1 FILLER_4_375 ();
 sg13g2_fill_1 FILLER_4_381 ();
 sg13g2_fill_2 FILLER_4_396 ();
 sg13g2_fill_1 FILLER_4_405 ();
 sg13g2_decap_8 FILLER_4_410 ();
 sg13g2_decap_4 FILLER_4_417 ();
 sg13g2_fill_1 FILLER_4_421 ();
 sg13g2_decap_8 FILLER_4_426 ();
 sg13g2_decap_8 FILLER_4_433 ();
 sg13g2_fill_1 FILLER_4_445 ();
 sg13g2_decap_4 FILLER_4_453 ();
 sg13g2_decap_4 FILLER_4_462 ();
 sg13g2_fill_1 FILLER_4_515 ();
 sg13g2_fill_1 FILLER_4_521 ();
 sg13g2_fill_1 FILLER_4_527 ();
 sg13g2_fill_2 FILLER_4_533 ();
 sg13g2_fill_2 FILLER_4_544 ();
 sg13g2_fill_1 FILLER_4_546 ();
 sg13g2_decap_4 FILLER_4_551 ();
 sg13g2_fill_1 FILLER_4_555 ();
 sg13g2_fill_1 FILLER_4_564 ();
 sg13g2_decap_8 FILLER_4_570 ();
 sg13g2_decap_8 FILLER_4_577 ();
 sg13g2_decap_8 FILLER_4_584 ();
 sg13g2_decap_8 FILLER_4_591 ();
 sg13g2_decap_8 FILLER_4_598 ();
 sg13g2_decap_8 FILLER_4_605 ();
 sg13g2_decap_8 FILLER_4_612 ();
 sg13g2_decap_8 FILLER_4_619 ();
 sg13g2_decap_8 FILLER_4_626 ();
 sg13g2_decap_8 FILLER_4_633 ();
 sg13g2_decap_8 FILLER_4_640 ();
 sg13g2_decap_8 FILLER_4_647 ();
 sg13g2_decap_8 FILLER_4_654 ();
 sg13g2_decap_8 FILLER_4_661 ();
 sg13g2_decap_8 FILLER_4_668 ();
 sg13g2_decap_8 FILLER_4_675 ();
 sg13g2_decap_8 FILLER_4_682 ();
 sg13g2_decap_8 FILLER_4_689 ();
 sg13g2_decap_8 FILLER_4_696 ();
 sg13g2_decap_8 FILLER_4_703 ();
 sg13g2_decap_8 FILLER_4_710 ();
 sg13g2_decap_8 FILLER_4_717 ();
 sg13g2_decap_8 FILLER_4_724 ();
 sg13g2_decap_8 FILLER_4_731 ();
 sg13g2_decap_8 FILLER_4_738 ();
 sg13g2_decap_8 FILLER_4_745 ();
 sg13g2_decap_8 FILLER_4_752 ();
 sg13g2_decap_8 FILLER_4_759 ();
 sg13g2_decap_8 FILLER_4_766 ();
 sg13g2_decap_8 FILLER_4_773 ();
 sg13g2_decap_8 FILLER_4_780 ();
 sg13g2_decap_8 FILLER_4_787 ();
 sg13g2_decap_8 FILLER_4_794 ();
 sg13g2_decap_8 FILLER_4_801 ();
 sg13g2_decap_8 FILLER_4_808 ();
 sg13g2_decap_8 FILLER_4_815 ();
 sg13g2_decap_8 FILLER_4_822 ();
 sg13g2_decap_8 FILLER_4_829 ();
 sg13g2_decap_8 FILLER_4_836 ();
 sg13g2_decap_8 FILLER_4_843 ();
 sg13g2_decap_8 FILLER_4_850 ();
 sg13g2_decap_8 FILLER_4_857 ();
 sg13g2_decap_8 FILLER_4_864 ();
 sg13g2_decap_8 FILLER_4_871 ();
 sg13g2_decap_8 FILLER_5_0 ();
 sg13g2_decap_8 FILLER_5_7 ();
 sg13g2_decap_8 FILLER_5_14 ();
 sg13g2_decap_8 FILLER_5_21 ();
 sg13g2_decap_8 FILLER_5_28 ();
 sg13g2_decap_8 FILLER_5_35 ();
 sg13g2_decap_8 FILLER_5_42 ();
 sg13g2_decap_8 FILLER_5_49 ();
 sg13g2_decap_8 FILLER_5_56 ();
 sg13g2_decap_8 FILLER_5_63 ();
 sg13g2_decap_8 FILLER_5_70 ();
 sg13g2_decap_8 FILLER_5_77 ();
 sg13g2_decap_8 FILLER_5_84 ();
 sg13g2_fill_1 FILLER_5_113 ();
 sg13g2_decap_8 FILLER_5_122 ();
 sg13g2_fill_1 FILLER_5_129 ();
 sg13g2_decap_4 FILLER_5_139 ();
 sg13g2_fill_2 FILLER_5_143 ();
 sg13g2_fill_2 FILLER_5_149 ();
 sg13g2_fill_2 FILLER_5_156 ();
 sg13g2_fill_1 FILLER_5_158 ();
 sg13g2_fill_1 FILLER_5_181 ();
 sg13g2_fill_1 FILLER_5_188 ();
 sg13g2_fill_1 FILLER_5_198 ();
 sg13g2_fill_1 FILLER_5_206 ();
 sg13g2_fill_2 FILLER_5_230 ();
 sg13g2_fill_2 FILLER_5_258 ();
 sg13g2_fill_2 FILLER_5_265 ();
 sg13g2_fill_1 FILLER_5_267 ();
 sg13g2_fill_1 FILLER_5_273 ();
 sg13g2_fill_1 FILLER_5_306 ();
 sg13g2_decap_4 FILLER_5_327 ();
 sg13g2_fill_1 FILLER_5_351 ();
 sg13g2_fill_2 FILLER_5_367 ();
 sg13g2_decap_8 FILLER_5_377 ();
 sg13g2_fill_2 FILLER_5_384 ();
 sg13g2_fill_1 FILLER_5_386 ();
 sg13g2_fill_1 FILLER_5_408 ();
 sg13g2_fill_2 FILLER_5_457 ();
 sg13g2_decap_8 FILLER_5_467 ();
 sg13g2_fill_2 FILLER_5_474 ();
 sg13g2_fill_1 FILLER_5_476 ();
 sg13g2_decap_4 FILLER_5_486 ();
 sg13g2_decap_4 FILLER_5_494 ();
 sg13g2_fill_1 FILLER_5_498 ();
 sg13g2_fill_1 FILLER_5_507 ();
 sg13g2_fill_2 FILLER_5_516 ();
 sg13g2_decap_4 FILLER_5_542 ();
 sg13g2_decap_8 FILLER_5_578 ();
 sg13g2_decap_8 FILLER_5_585 ();
 sg13g2_decap_8 FILLER_5_592 ();
 sg13g2_decap_8 FILLER_5_599 ();
 sg13g2_decap_8 FILLER_5_606 ();
 sg13g2_decap_8 FILLER_5_613 ();
 sg13g2_decap_8 FILLER_5_620 ();
 sg13g2_decap_8 FILLER_5_627 ();
 sg13g2_decap_8 FILLER_5_634 ();
 sg13g2_decap_8 FILLER_5_641 ();
 sg13g2_decap_8 FILLER_5_648 ();
 sg13g2_decap_8 FILLER_5_655 ();
 sg13g2_decap_8 FILLER_5_662 ();
 sg13g2_decap_8 FILLER_5_669 ();
 sg13g2_decap_8 FILLER_5_676 ();
 sg13g2_decap_8 FILLER_5_683 ();
 sg13g2_decap_8 FILLER_5_690 ();
 sg13g2_decap_8 FILLER_5_697 ();
 sg13g2_decap_8 FILLER_5_704 ();
 sg13g2_decap_8 FILLER_5_711 ();
 sg13g2_decap_8 FILLER_5_718 ();
 sg13g2_decap_8 FILLER_5_725 ();
 sg13g2_decap_8 FILLER_5_732 ();
 sg13g2_decap_8 FILLER_5_739 ();
 sg13g2_decap_8 FILLER_5_746 ();
 sg13g2_decap_8 FILLER_5_753 ();
 sg13g2_decap_8 FILLER_5_760 ();
 sg13g2_decap_8 FILLER_5_767 ();
 sg13g2_decap_8 FILLER_5_774 ();
 sg13g2_decap_8 FILLER_5_781 ();
 sg13g2_decap_8 FILLER_5_788 ();
 sg13g2_decap_8 FILLER_5_795 ();
 sg13g2_decap_8 FILLER_5_802 ();
 sg13g2_decap_8 FILLER_5_809 ();
 sg13g2_decap_8 FILLER_5_816 ();
 sg13g2_decap_8 FILLER_5_823 ();
 sg13g2_decap_8 FILLER_5_830 ();
 sg13g2_decap_8 FILLER_5_837 ();
 sg13g2_decap_8 FILLER_5_844 ();
 sg13g2_decap_8 FILLER_5_851 ();
 sg13g2_decap_8 FILLER_5_858 ();
 sg13g2_decap_8 FILLER_5_865 ();
 sg13g2_decap_4 FILLER_5_872 ();
 sg13g2_fill_2 FILLER_5_876 ();
 sg13g2_decap_8 FILLER_6_0 ();
 sg13g2_decap_8 FILLER_6_7 ();
 sg13g2_decap_8 FILLER_6_14 ();
 sg13g2_decap_8 FILLER_6_21 ();
 sg13g2_decap_8 FILLER_6_28 ();
 sg13g2_decap_8 FILLER_6_35 ();
 sg13g2_decap_8 FILLER_6_42 ();
 sg13g2_decap_8 FILLER_6_49 ();
 sg13g2_decap_8 FILLER_6_56 ();
 sg13g2_decap_8 FILLER_6_63 ();
 sg13g2_decap_4 FILLER_6_70 ();
 sg13g2_fill_1 FILLER_6_74 ();
 sg13g2_decap_4 FILLER_6_84 ();
 sg13g2_fill_1 FILLER_6_101 ();
 sg13g2_fill_1 FILLER_6_118 ();
 sg13g2_decap_8 FILLER_6_131 ();
 sg13g2_fill_2 FILLER_6_138 ();
 sg13g2_fill_1 FILLER_6_140 ();
 sg13g2_fill_2 FILLER_6_155 ();
 sg13g2_fill_1 FILLER_6_157 ();
 sg13g2_fill_2 FILLER_6_192 ();
 sg13g2_decap_4 FILLER_6_221 ();
 sg13g2_fill_2 FILLER_6_234 ();
 sg13g2_decap_4 FILLER_6_240 ();
 sg13g2_decap_8 FILLER_6_262 ();
 sg13g2_fill_1 FILLER_6_269 ();
 sg13g2_fill_2 FILLER_6_286 ();
 sg13g2_fill_1 FILLER_6_321 ();
 sg13g2_fill_2 FILLER_6_328 ();
 sg13g2_decap_4 FILLER_6_334 ();
 sg13g2_fill_1 FILLER_6_343 ();
 sg13g2_fill_1 FILLER_6_352 ();
 sg13g2_fill_2 FILLER_6_374 ();
 sg13g2_fill_1 FILLER_6_376 ();
 sg13g2_fill_1 FILLER_6_390 ();
 sg13g2_fill_2 FILLER_6_396 ();
 sg13g2_decap_4 FILLER_6_407 ();
 sg13g2_fill_2 FILLER_6_411 ();
 sg13g2_fill_1 FILLER_6_417 ();
 sg13g2_decap_4 FILLER_6_434 ();
 sg13g2_decap_8 FILLER_6_442 ();
 sg13g2_fill_2 FILLER_6_449 ();
 sg13g2_fill_2 FILLER_6_495 ();
 sg13g2_decap_8 FILLER_6_522 ();
 sg13g2_decap_8 FILLER_6_529 ();
 sg13g2_decap_4 FILLER_6_536 ();
 sg13g2_fill_2 FILLER_6_540 ();
 sg13g2_fill_2 FILLER_6_546 ();
 sg13g2_fill_1 FILLER_6_548 ();
 sg13g2_fill_2 FILLER_6_557 ();
 sg13g2_fill_1 FILLER_6_563 ();
 sg13g2_fill_1 FILLER_6_570 ();
 sg13g2_decap_8 FILLER_6_576 ();
 sg13g2_decap_8 FILLER_6_583 ();
 sg13g2_decap_8 FILLER_6_590 ();
 sg13g2_decap_8 FILLER_6_597 ();
 sg13g2_decap_8 FILLER_6_604 ();
 sg13g2_decap_8 FILLER_6_611 ();
 sg13g2_decap_8 FILLER_6_618 ();
 sg13g2_decap_4 FILLER_6_625 ();
 sg13g2_fill_1 FILLER_6_629 ();
 sg13g2_decap_8 FILLER_6_634 ();
 sg13g2_decap_8 FILLER_6_641 ();
 sg13g2_decap_8 FILLER_6_648 ();
 sg13g2_decap_8 FILLER_6_655 ();
 sg13g2_decap_8 FILLER_6_662 ();
 sg13g2_decap_8 FILLER_6_669 ();
 sg13g2_decap_8 FILLER_6_676 ();
 sg13g2_decap_4 FILLER_6_683 ();
 sg13g2_decap_8 FILLER_6_695 ();
 sg13g2_decap_4 FILLER_6_710 ();
 sg13g2_fill_2 FILLER_6_714 ();
 sg13g2_decap_8 FILLER_6_721 ();
 sg13g2_decap_8 FILLER_6_728 ();
 sg13g2_fill_2 FILLER_6_743 ();
 sg13g2_decap_8 FILLER_6_775 ();
 sg13g2_decap_8 FILLER_6_782 ();
 sg13g2_decap_8 FILLER_6_789 ();
 sg13g2_decap_8 FILLER_6_796 ();
 sg13g2_decap_8 FILLER_6_803 ();
 sg13g2_decap_8 FILLER_6_810 ();
 sg13g2_decap_8 FILLER_6_817 ();
 sg13g2_decap_8 FILLER_6_824 ();
 sg13g2_decap_8 FILLER_6_831 ();
 sg13g2_decap_8 FILLER_6_838 ();
 sg13g2_decap_8 FILLER_6_845 ();
 sg13g2_decap_8 FILLER_6_852 ();
 sg13g2_decap_8 FILLER_6_859 ();
 sg13g2_decap_8 FILLER_6_866 ();
 sg13g2_decap_4 FILLER_6_873 ();
 sg13g2_fill_1 FILLER_6_877 ();
 sg13g2_decap_8 FILLER_7_0 ();
 sg13g2_decap_8 FILLER_7_7 ();
 sg13g2_decap_8 FILLER_7_14 ();
 sg13g2_decap_8 FILLER_7_21 ();
 sg13g2_decap_8 FILLER_7_28 ();
 sg13g2_decap_8 FILLER_7_35 ();
 sg13g2_decap_8 FILLER_7_42 ();
 sg13g2_decap_8 FILLER_7_49 ();
 sg13g2_decap_8 FILLER_7_56 ();
 sg13g2_decap_8 FILLER_7_63 ();
 sg13g2_decap_4 FILLER_7_70 ();
 sg13g2_decap_4 FILLER_7_105 ();
 sg13g2_fill_1 FILLER_7_109 ();
 sg13g2_fill_1 FILLER_7_114 ();
 sg13g2_fill_2 FILLER_7_132 ();
 sg13g2_decap_4 FILLER_7_138 ();
 sg13g2_fill_2 FILLER_7_142 ();
 sg13g2_decap_8 FILLER_7_172 ();
 sg13g2_fill_2 FILLER_7_179 ();
 sg13g2_fill_1 FILLER_7_197 ();
 sg13g2_fill_1 FILLER_7_206 ();
 sg13g2_fill_1 FILLER_7_212 ();
 sg13g2_fill_1 FILLER_7_217 ();
 sg13g2_decap_4 FILLER_7_240 ();
 sg13g2_decap_8 FILLER_7_252 ();
 sg13g2_decap_4 FILLER_7_259 ();
 sg13g2_decap_4 FILLER_7_271 ();
 sg13g2_decap_4 FILLER_7_281 ();
 sg13g2_fill_1 FILLER_7_291 ();
 sg13g2_decap_4 FILLER_7_298 ();
 sg13g2_fill_2 FILLER_7_322 ();
 sg13g2_fill_2 FILLER_7_355 ();
 sg13g2_fill_1 FILLER_7_357 ();
 sg13g2_decap_8 FILLER_7_370 ();
 sg13g2_decap_4 FILLER_7_377 ();
 sg13g2_decap_8 FILLER_7_385 ();
 sg13g2_decap_8 FILLER_7_392 ();
 sg13g2_fill_1 FILLER_7_403 ();
 sg13g2_fill_1 FILLER_7_416 ();
 sg13g2_fill_2 FILLER_7_421 ();
 sg13g2_decap_8 FILLER_7_432 ();
 sg13g2_fill_2 FILLER_7_453 ();
 sg13g2_fill_2 FILLER_7_462 ();
 sg13g2_fill_1 FILLER_7_464 ();
 sg13g2_fill_2 FILLER_7_470 ();
 sg13g2_fill_1 FILLER_7_472 ();
 sg13g2_fill_2 FILLER_7_479 ();
 sg13g2_decap_8 FILLER_7_497 ();
 sg13g2_decap_4 FILLER_7_522 ();
 sg13g2_fill_1 FILLER_7_526 ();
 sg13g2_decap_4 FILLER_7_532 ();
 sg13g2_fill_2 FILLER_7_536 ();
 sg13g2_fill_1 FILLER_7_547 ();
 sg13g2_fill_1 FILLER_7_552 ();
 sg13g2_fill_1 FILLER_7_558 ();
 sg13g2_fill_1 FILLER_7_563 ();
 sg13g2_fill_1 FILLER_7_569 ();
 sg13g2_fill_1 FILLER_7_574 ();
 sg13g2_fill_1 FILLER_7_579 ();
 sg13g2_fill_1 FILLER_7_585 ();
 sg13g2_fill_1 FILLER_7_590 ();
 sg13g2_fill_2 FILLER_7_596 ();
 sg13g2_decap_8 FILLER_7_602 ();
 sg13g2_decap_8 FILLER_7_609 ();
 sg13g2_fill_2 FILLER_7_635 ();
 sg13g2_fill_1 FILLER_7_637 ();
 sg13g2_decap_8 FILLER_7_651 ();
 sg13g2_fill_1 FILLER_7_658 ();
 sg13g2_fill_1 FILLER_7_669 ();
 sg13g2_decap_4 FILLER_7_678 ();
 sg13g2_fill_1 FILLER_7_682 ();
 sg13g2_fill_1 FILLER_7_696 ();
 sg13g2_fill_2 FILLER_7_721 ();
 sg13g2_decap_4 FILLER_7_727 ();
 sg13g2_fill_2 FILLER_7_753 ();
 sg13g2_fill_1 FILLER_7_755 ();
 sg13g2_decap_8 FILLER_7_769 ();
 sg13g2_decap_8 FILLER_7_776 ();
 sg13g2_decap_8 FILLER_7_783 ();
 sg13g2_decap_8 FILLER_7_790 ();
 sg13g2_decap_8 FILLER_7_797 ();
 sg13g2_decap_8 FILLER_7_804 ();
 sg13g2_decap_8 FILLER_7_811 ();
 sg13g2_decap_8 FILLER_7_818 ();
 sg13g2_decap_8 FILLER_7_825 ();
 sg13g2_decap_8 FILLER_7_832 ();
 sg13g2_decap_8 FILLER_7_839 ();
 sg13g2_decap_8 FILLER_7_846 ();
 sg13g2_decap_8 FILLER_7_853 ();
 sg13g2_decap_8 FILLER_7_860 ();
 sg13g2_decap_8 FILLER_7_867 ();
 sg13g2_decap_4 FILLER_7_874 ();
 sg13g2_decap_8 FILLER_8_0 ();
 sg13g2_decap_8 FILLER_8_7 ();
 sg13g2_decap_8 FILLER_8_14 ();
 sg13g2_decap_8 FILLER_8_21 ();
 sg13g2_decap_8 FILLER_8_28 ();
 sg13g2_decap_8 FILLER_8_35 ();
 sg13g2_decap_8 FILLER_8_42 ();
 sg13g2_decap_8 FILLER_8_49 ();
 sg13g2_decap_8 FILLER_8_56 ();
 sg13g2_decap_8 FILLER_8_63 ();
 sg13g2_decap_4 FILLER_8_70 ();
 sg13g2_fill_1 FILLER_8_74 ();
 sg13g2_decap_4 FILLER_8_79 ();
 sg13g2_decap_4 FILLER_8_104 ();
 sg13g2_decap_4 FILLER_8_132 ();
 sg13g2_fill_2 FILLER_8_136 ();
 sg13g2_decap_8 FILLER_8_164 ();
 sg13g2_fill_1 FILLER_8_171 ();
 sg13g2_decap_8 FILLER_8_176 ();
 sg13g2_decap_4 FILLER_8_183 ();
 sg13g2_fill_1 FILLER_8_187 ();
 sg13g2_decap_8 FILLER_8_210 ();
 sg13g2_fill_1 FILLER_8_217 ();
 sg13g2_fill_2 FILLER_8_231 ();
 sg13g2_fill_1 FILLER_8_233 ();
 sg13g2_decap_4 FILLER_8_266 ();
 sg13g2_fill_1 FILLER_8_274 ();
 sg13g2_fill_2 FILLER_8_285 ();
 sg13g2_decap_4 FILLER_8_299 ();
 sg13g2_fill_1 FILLER_8_303 ();
 sg13g2_decap_8 FILLER_8_322 ();
 sg13g2_decap_8 FILLER_8_329 ();
 sg13g2_decap_8 FILLER_8_336 ();
 sg13g2_fill_1 FILLER_8_343 ();
 sg13g2_fill_1 FILLER_8_363 ();
 sg13g2_fill_1 FILLER_8_371 ();
 sg13g2_fill_1 FILLER_8_376 ();
 sg13g2_fill_2 FILLER_8_382 ();
 sg13g2_decap_8 FILLER_8_395 ();
 sg13g2_fill_2 FILLER_8_402 ();
 sg13g2_fill_1 FILLER_8_404 ();
 sg13g2_fill_2 FILLER_8_429 ();
 sg13g2_decap_4 FILLER_8_442 ();
 sg13g2_fill_1 FILLER_8_450 ();
 sg13g2_fill_1 FILLER_8_457 ();
 sg13g2_decap_8 FILLER_8_463 ();
 sg13g2_decap_4 FILLER_8_470 ();
 sg13g2_decap_8 FILLER_8_482 ();
 sg13g2_decap_8 FILLER_8_489 ();
 sg13g2_decap_4 FILLER_8_496 ();
 sg13g2_fill_1 FILLER_8_505 ();
 sg13g2_fill_2 FILLER_8_516 ();
 sg13g2_fill_1 FILLER_8_558 ();
 sg13g2_decap_8 FILLER_8_563 ();
 sg13g2_decap_4 FILLER_8_570 ();
 sg13g2_fill_2 FILLER_8_574 ();
 sg13g2_fill_1 FILLER_8_596 ();
 sg13g2_decap_8 FILLER_8_601 ();
 sg13g2_fill_1 FILLER_8_608 ();
 sg13g2_fill_1 FILLER_8_629 ();
 sg13g2_decap_4 FILLER_8_634 ();
 sg13g2_fill_2 FILLER_8_652 ();
 sg13g2_decap_8 FILLER_8_666 ();
 sg13g2_fill_2 FILLER_8_673 ();
 sg13g2_fill_1 FILLER_8_675 ();
 sg13g2_decap_8 FILLER_8_690 ();
 sg13g2_decap_4 FILLER_8_697 ();
 sg13g2_fill_2 FILLER_8_701 ();
 sg13g2_fill_1 FILLER_8_707 ();
 sg13g2_fill_1 FILLER_8_713 ();
 sg13g2_fill_2 FILLER_8_719 ();
 sg13g2_decap_4 FILLER_8_739 ();
 sg13g2_fill_1 FILLER_8_755 ();
 sg13g2_decap_8 FILLER_8_769 ();
 sg13g2_decap_8 FILLER_8_776 ();
 sg13g2_decap_8 FILLER_8_783 ();
 sg13g2_decap_8 FILLER_8_790 ();
 sg13g2_decap_8 FILLER_8_797 ();
 sg13g2_decap_8 FILLER_8_804 ();
 sg13g2_decap_8 FILLER_8_811 ();
 sg13g2_decap_8 FILLER_8_818 ();
 sg13g2_decap_8 FILLER_8_825 ();
 sg13g2_decap_8 FILLER_8_832 ();
 sg13g2_decap_8 FILLER_8_839 ();
 sg13g2_decap_8 FILLER_8_846 ();
 sg13g2_decap_8 FILLER_8_853 ();
 sg13g2_decap_8 FILLER_8_860 ();
 sg13g2_decap_8 FILLER_8_867 ();
 sg13g2_decap_4 FILLER_8_874 ();
 sg13g2_decap_8 FILLER_9_0 ();
 sg13g2_decap_8 FILLER_9_7 ();
 sg13g2_decap_8 FILLER_9_14 ();
 sg13g2_decap_8 FILLER_9_21 ();
 sg13g2_decap_8 FILLER_9_28 ();
 sg13g2_decap_8 FILLER_9_35 ();
 sg13g2_decap_8 FILLER_9_42 ();
 sg13g2_decap_8 FILLER_9_49 ();
 sg13g2_decap_8 FILLER_9_56 ();
 sg13g2_decap_4 FILLER_9_63 ();
 sg13g2_fill_2 FILLER_9_67 ();
 sg13g2_decap_4 FILLER_9_82 ();
 sg13g2_fill_1 FILLER_9_86 ();
 sg13g2_fill_1 FILLER_9_92 ();
 sg13g2_decap_8 FILLER_9_101 ();
 sg13g2_decap_4 FILLER_9_108 ();
 sg13g2_fill_2 FILLER_9_112 ();
 sg13g2_decap_8 FILLER_9_121 ();
 sg13g2_decap_8 FILLER_9_128 ();
 sg13g2_decap_4 FILLER_9_135 ();
 sg13g2_decap_8 FILLER_9_160 ();
 sg13g2_decap_4 FILLER_9_167 ();
 sg13g2_fill_1 FILLER_9_171 ();
 sg13g2_decap_4 FILLER_9_196 ();
 sg13g2_decap_8 FILLER_9_204 ();
 sg13g2_fill_2 FILLER_9_211 ();
 sg13g2_fill_1 FILLER_9_213 ();
 sg13g2_fill_1 FILLER_9_219 ();
 sg13g2_fill_1 FILLER_9_234 ();
 sg13g2_decap_8 FILLER_9_243 ();
 sg13g2_decap_8 FILLER_9_250 ();
 sg13g2_decap_4 FILLER_9_257 ();
 sg13g2_fill_2 FILLER_9_261 ();
 sg13g2_decap_4 FILLER_9_267 ();
 sg13g2_fill_2 FILLER_9_271 ();
 sg13g2_decap_8 FILLER_9_293 ();
 sg13g2_decap_4 FILLER_9_300 ();
 sg13g2_fill_2 FILLER_9_308 ();
 sg13g2_fill_1 FILLER_9_310 ();
 sg13g2_fill_1 FILLER_9_330 ();
 sg13g2_decap_8 FILLER_9_365 ();
 sg13g2_fill_2 FILLER_9_372 ();
 sg13g2_fill_1 FILLER_9_374 ();
 sg13g2_fill_2 FILLER_9_380 ();
 sg13g2_fill_2 FILLER_9_386 ();
 sg13g2_fill_1 FILLER_9_393 ();
 sg13g2_fill_1 FILLER_9_422 ();
 sg13g2_decap_4 FILLER_9_430 ();
 sg13g2_fill_1 FILLER_9_434 ();
 sg13g2_decap_4 FILLER_9_442 ();
 sg13g2_fill_1 FILLER_9_450 ();
 sg13g2_fill_2 FILLER_9_466 ();
 sg13g2_fill_2 FILLER_9_502 ();
 sg13g2_fill_2 FILLER_9_529 ();
 sg13g2_fill_2 FILLER_9_543 ();
 sg13g2_fill_1 FILLER_9_545 ();
 sg13g2_decap_8 FILLER_9_554 ();
 sg13g2_decap_8 FILLER_9_561 ();
 sg13g2_decap_4 FILLER_9_568 ();
 sg13g2_fill_2 FILLER_9_580 ();
 sg13g2_fill_2 FILLER_9_592 ();
 sg13g2_fill_2 FILLER_9_610 ();
 sg13g2_fill_2 FILLER_9_628 ();
 sg13g2_fill_1 FILLER_9_630 ();
 sg13g2_fill_1 FILLER_9_639 ();
 sg13g2_decap_4 FILLER_9_653 ();
 sg13g2_decap_4 FILLER_9_667 ();
 sg13g2_fill_1 FILLER_9_680 ();
 sg13g2_fill_2 FILLER_9_723 ();
 sg13g2_fill_1 FILLER_9_725 ();
 sg13g2_fill_2 FILLER_9_747 ();
 sg13g2_fill_1 FILLER_9_749 ();
 sg13g2_fill_2 FILLER_9_755 ();
 sg13g2_decap_8 FILLER_9_771 ();
 sg13g2_decap_8 FILLER_9_778 ();
 sg13g2_decap_8 FILLER_9_785 ();
 sg13g2_decap_8 FILLER_9_792 ();
 sg13g2_decap_8 FILLER_9_799 ();
 sg13g2_decap_8 FILLER_9_806 ();
 sg13g2_decap_8 FILLER_9_813 ();
 sg13g2_decap_8 FILLER_9_820 ();
 sg13g2_decap_8 FILLER_9_827 ();
 sg13g2_decap_8 FILLER_9_834 ();
 sg13g2_decap_8 FILLER_9_841 ();
 sg13g2_decap_8 FILLER_9_848 ();
 sg13g2_decap_8 FILLER_9_855 ();
 sg13g2_decap_8 FILLER_9_862 ();
 sg13g2_decap_8 FILLER_9_869 ();
 sg13g2_fill_2 FILLER_9_876 ();
 sg13g2_decap_8 FILLER_10_0 ();
 sg13g2_decap_8 FILLER_10_7 ();
 sg13g2_decap_8 FILLER_10_14 ();
 sg13g2_decap_8 FILLER_10_21 ();
 sg13g2_decap_8 FILLER_10_28 ();
 sg13g2_decap_8 FILLER_10_35 ();
 sg13g2_decap_8 FILLER_10_42 ();
 sg13g2_decap_8 FILLER_10_49 ();
 sg13g2_decap_8 FILLER_10_56 ();
 sg13g2_decap_4 FILLER_10_63 ();
 sg13g2_fill_2 FILLER_10_67 ();
 sg13g2_decap_8 FILLER_10_73 ();
 sg13g2_fill_1 FILLER_10_104 ();
 sg13g2_fill_2 FILLER_10_134 ();
 sg13g2_fill_1 FILLER_10_136 ();
 sg13g2_fill_2 FILLER_10_146 ();
 sg13g2_fill_2 FILLER_10_152 ();
 sg13g2_decap_4 FILLER_10_162 ();
 sg13g2_fill_1 FILLER_10_166 ();
 sg13g2_decap_4 FILLER_10_195 ();
 sg13g2_fill_1 FILLER_10_212 ();
 sg13g2_decap_8 FILLER_10_223 ();
 sg13g2_fill_2 FILLER_10_230 ();
 sg13g2_fill_1 FILLER_10_232 ();
 sg13g2_decap_8 FILLER_10_243 ();
 sg13g2_fill_2 FILLER_10_259 ();
 sg13g2_fill_2 FILLER_10_269 ();
 sg13g2_fill_1 FILLER_10_271 ();
 sg13g2_decap_4 FILLER_10_277 ();
 sg13g2_fill_1 FILLER_10_299 ();
 sg13g2_fill_1 FILLER_10_305 ();
 sg13g2_fill_1 FILLER_10_310 ();
 sg13g2_fill_1 FILLER_10_319 ();
 sg13g2_fill_1 FILLER_10_326 ();
 sg13g2_decap_8 FILLER_10_343 ();
 sg13g2_decap_4 FILLER_10_350 ();
 sg13g2_fill_1 FILLER_10_359 ();
 sg13g2_fill_1 FILLER_10_365 ();
 sg13g2_fill_2 FILLER_10_370 ();
 sg13g2_fill_1 FILLER_10_377 ();
 sg13g2_fill_2 FILLER_10_390 ();
 sg13g2_decap_4 FILLER_10_412 ();
 sg13g2_fill_1 FILLER_10_416 ();
 sg13g2_fill_1 FILLER_10_426 ();
 sg13g2_decap_4 FILLER_10_448 ();
 sg13g2_fill_2 FILLER_10_452 ();
 sg13g2_fill_1 FILLER_10_461 ();
 sg13g2_fill_2 FILLER_10_466 ();
 sg13g2_fill_1 FILLER_10_501 ();
 sg13g2_fill_1 FILLER_10_509 ();
 sg13g2_decap_4 FILLER_10_519 ();
 sg13g2_fill_2 FILLER_10_535 ();
 sg13g2_decap_4 FILLER_10_551 ();
 sg13g2_fill_2 FILLER_10_568 ();
 sg13g2_decap_4 FILLER_10_583 ();
 sg13g2_fill_2 FILLER_10_587 ();
 sg13g2_decap_4 FILLER_10_602 ();
 sg13g2_decap_4 FILLER_10_623 ();
 sg13g2_fill_2 FILLER_10_627 ();
 sg13g2_fill_1 FILLER_10_647 ();
 sg13g2_fill_1 FILLER_10_652 ();
 sg13g2_fill_2 FILLER_10_658 ();
 sg13g2_fill_2 FILLER_10_664 ();
 sg13g2_fill_2 FILLER_10_670 ();
 sg13g2_fill_1 FILLER_10_693 ();
 sg13g2_fill_1 FILLER_10_698 ();
 sg13g2_decap_4 FILLER_10_704 ();
 sg13g2_fill_1 FILLER_10_708 ();
 sg13g2_decap_8 FILLER_10_721 ();
 sg13g2_decap_8 FILLER_10_728 ();
 sg13g2_decap_8 FILLER_10_775 ();
 sg13g2_decap_8 FILLER_10_782 ();
 sg13g2_decap_8 FILLER_10_789 ();
 sg13g2_decap_8 FILLER_10_796 ();
 sg13g2_decap_8 FILLER_10_803 ();
 sg13g2_decap_8 FILLER_10_810 ();
 sg13g2_decap_8 FILLER_10_817 ();
 sg13g2_decap_8 FILLER_10_824 ();
 sg13g2_decap_8 FILLER_10_831 ();
 sg13g2_decap_8 FILLER_10_838 ();
 sg13g2_decap_8 FILLER_10_845 ();
 sg13g2_decap_8 FILLER_10_852 ();
 sg13g2_decap_8 FILLER_10_859 ();
 sg13g2_decap_8 FILLER_10_866 ();
 sg13g2_decap_4 FILLER_10_873 ();
 sg13g2_fill_1 FILLER_10_877 ();
 sg13g2_decap_8 FILLER_11_0 ();
 sg13g2_decap_8 FILLER_11_7 ();
 sg13g2_decap_8 FILLER_11_14 ();
 sg13g2_decap_8 FILLER_11_21 ();
 sg13g2_decap_8 FILLER_11_28 ();
 sg13g2_decap_8 FILLER_11_35 ();
 sg13g2_decap_8 FILLER_11_42 ();
 sg13g2_decap_8 FILLER_11_49 ();
 sg13g2_fill_2 FILLER_11_56 ();
 sg13g2_fill_1 FILLER_11_58 ();
 sg13g2_fill_1 FILLER_11_79 ();
 sg13g2_decap_8 FILLER_11_84 ();
 sg13g2_decap_4 FILLER_11_101 ();
 sg13g2_fill_2 FILLER_11_113 ();
 sg13g2_fill_1 FILLER_11_115 ();
 sg13g2_fill_1 FILLER_11_122 ();
 sg13g2_fill_1 FILLER_11_130 ();
 sg13g2_fill_2 FILLER_11_153 ();
 sg13g2_fill_1 FILLER_11_160 ();
 sg13g2_fill_1 FILLER_11_165 ();
 sg13g2_fill_2 FILLER_11_170 ();
 sg13g2_fill_1 FILLER_11_182 ();
 sg13g2_fill_2 FILLER_11_191 ();
 sg13g2_fill_1 FILLER_11_201 ();
 sg13g2_decap_4 FILLER_11_210 ();
 sg13g2_fill_2 FILLER_11_217 ();
 sg13g2_fill_2 FILLER_11_223 ();
 sg13g2_decap_8 FILLER_11_233 ();
 sg13g2_decap_4 FILLER_11_282 ();
 sg13g2_fill_2 FILLER_11_286 ();
 sg13g2_fill_2 FILLER_11_293 ();
 sg13g2_fill_1 FILLER_11_303 ();
 sg13g2_decap_8 FILLER_11_309 ();
 sg13g2_fill_2 FILLER_11_316 ();
 sg13g2_fill_2 FILLER_11_337 ();
 sg13g2_fill_2 FILLER_11_358 ();
 sg13g2_fill_1 FILLER_11_360 ();
 sg13g2_fill_2 FILLER_11_366 ();
 sg13g2_fill_2 FILLER_11_410 ();
 sg13g2_fill_1 FILLER_11_412 ();
 sg13g2_decap_4 FILLER_11_423 ();
 sg13g2_decap_8 FILLER_11_432 ();
 sg13g2_decap_8 FILLER_11_444 ();
 sg13g2_fill_1 FILLER_11_456 ();
 sg13g2_fill_2 FILLER_11_466 ();
 sg13g2_fill_1 FILLER_11_473 ();
 sg13g2_fill_2 FILLER_11_479 ();
 sg13g2_fill_2 FILLER_11_494 ();
 sg13g2_fill_2 FILLER_11_518 ();
 sg13g2_decap_4 FILLER_11_525 ();
 sg13g2_fill_1 FILLER_11_529 ();
 sg13g2_fill_1 FILLER_11_534 ();
 sg13g2_decap_8 FILLER_11_548 ();
 sg13g2_decap_4 FILLER_11_555 ();
 sg13g2_fill_1 FILLER_11_559 ();
 sg13g2_decap_4 FILLER_11_573 ();
 sg13g2_fill_1 FILLER_11_577 ();
 sg13g2_fill_1 FILLER_11_589 ();
 sg13g2_fill_1 FILLER_11_598 ();
 sg13g2_fill_2 FILLER_11_640 ();
 sg13g2_fill_1 FILLER_11_642 ();
 sg13g2_fill_2 FILLER_11_658 ();
 sg13g2_fill_2 FILLER_11_669 ();
 sg13g2_fill_1 FILLER_11_671 ();
 sg13g2_fill_2 FILLER_11_677 ();
 sg13g2_fill_2 FILLER_11_700 ();
 sg13g2_decap_4 FILLER_11_706 ();
 sg13g2_fill_2 FILLER_11_715 ();
 sg13g2_fill_1 FILLER_11_717 ();
 sg13g2_fill_1 FILLER_11_735 ();
 sg13g2_fill_1 FILLER_11_741 ();
 sg13g2_fill_1 FILLER_11_747 ();
 sg13g2_fill_1 FILLER_11_758 ();
 sg13g2_fill_1 FILLER_11_765 ();
 sg13g2_decap_8 FILLER_11_774 ();
 sg13g2_decap_8 FILLER_11_781 ();
 sg13g2_decap_8 FILLER_11_788 ();
 sg13g2_decap_8 FILLER_11_795 ();
 sg13g2_decap_8 FILLER_11_802 ();
 sg13g2_decap_8 FILLER_11_809 ();
 sg13g2_decap_8 FILLER_11_816 ();
 sg13g2_decap_8 FILLER_11_823 ();
 sg13g2_decap_8 FILLER_11_830 ();
 sg13g2_decap_8 FILLER_11_837 ();
 sg13g2_decap_8 FILLER_11_844 ();
 sg13g2_decap_8 FILLER_11_851 ();
 sg13g2_decap_8 FILLER_11_858 ();
 sg13g2_decap_8 FILLER_11_865 ();
 sg13g2_decap_4 FILLER_11_872 ();
 sg13g2_fill_2 FILLER_11_876 ();
 sg13g2_decap_8 FILLER_12_0 ();
 sg13g2_decap_8 FILLER_12_7 ();
 sg13g2_decap_8 FILLER_12_14 ();
 sg13g2_decap_8 FILLER_12_21 ();
 sg13g2_decap_8 FILLER_12_28 ();
 sg13g2_decap_8 FILLER_12_35 ();
 sg13g2_decap_8 FILLER_12_42 ();
 sg13g2_decap_8 FILLER_12_49 ();
 sg13g2_decap_4 FILLER_12_56 ();
 sg13g2_fill_1 FILLER_12_80 ();
 sg13g2_fill_1 FILLER_12_86 ();
 sg13g2_fill_1 FILLER_12_97 ();
 sg13g2_decap_8 FILLER_12_102 ();
 sg13g2_fill_2 FILLER_12_109 ();
 sg13g2_fill_1 FILLER_12_111 ();
 sg13g2_fill_1 FILLER_12_117 ();
 sg13g2_fill_2 FILLER_12_132 ();
 sg13g2_fill_2 FILLER_12_142 ();
 sg13g2_fill_1 FILLER_12_155 ();
 sg13g2_fill_2 FILLER_12_164 ();
 sg13g2_fill_2 FILLER_12_174 ();
 sg13g2_fill_2 FILLER_12_181 ();
 sg13g2_decap_8 FILLER_12_203 ();
 sg13g2_decap_4 FILLER_12_210 ();
 sg13g2_fill_1 FILLER_12_214 ();
 sg13g2_decap_4 FILLER_12_237 ();
 sg13g2_fill_2 FILLER_12_241 ();
 sg13g2_decap_4 FILLER_12_274 ();
 sg13g2_fill_2 FILLER_12_278 ();
 sg13g2_decap_4 FILLER_12_299 ();
 sg13g2_fill_1 FILLER_12_303 ();
 sg13g2_fill_2 FILLER_12_308 ();
 sg13g2_fill_1 FILLER_12_310 ();
 sg13g2_decap_8 FILLER_12_336 ();
 sg13g2_decap_4 FILLER_12_343 ();
 sg13g2_fill_1 FILLER_12_347 ();
 sg13g2_fill_2 FILLER_12_391 ();
 sg13g2_fill_2 FILLER_12_421 ();
 sg13g2_decap_4 FILLER_12_429 ();
 sg13g2_fill_1 FILLER_12_433 ();
 sg13g2_fill_1 FILLER_12_450 ();
 sg13g2_fill_1 FILLER_12_463 ();
 sg13g2_decap_8 FILLER_12_470 ();
 sg13g2_fill_2 FILLER_12_477 ();
 sg13g2_fill_1 FILLER_12_479 ();
 sg13g2_fill_1 FILLER_12_485 ();
 sg13g2_fill_1 FILLER_12_491 ();
 sg13g2_fill_1 FILLER_12_509 ();
 sg13g2_decap_4 FILLER_12_515 ();
 sg13g2_fill_2 FILLER_12_519 ();
 sg13g2_fill_1 FILLER_12_530 ();
 sg13g2_fill_1 FILLER_12_536 ();
 sg13g2_fill_1 FILLER_12_544 ();
 sg13g2_decap_8 FILLER_12_549 ();
 sg13g2_decap_8 FILLER_12_556 ();
 sg13g2_decap_8 FILLER_12_563 ();
 sg13g2_fill_2 FILLER_12_570 ();
 sg13g2_fill_2 FILLER_12_629 ();
 sg13g2_decap_4 FILLER_12_645 ();
 sg13g2_fill_1 FILLER_12_649 ();
 sg13g2_fill_1 FILLER_12_686 ();
 sg13g2_fill_2 FILLER_12_705 ();
 sg13g2_fill_1 FILLER_12_707 ();
 sg13g2_fill_2 FILLER_12_736 ();
 sg13g2_fill_2 FILLER_12_745 ();
 sg13g2_fill_1 FILLER_12_747 ();
 sg13g2_decap_8 FILLER_12_756 ();
 sg13g2_decap_8 FILLER_12_763 ();
 sg13g2_decap_8 FILLER_12_770 ();
 sg13g2_decap_8 FILLER_12_777 ();
 sg13g2_decap_8 FILLER_12_784 ();
 sg13g2_decap_8 FILLER_12_791 ();
 sg13g2_decap_8 FILLER_12_798 ();
 sg13g2_decap_8 FILLER_12_805 ();
 sg13g2_decap_8 FILLER_12_812 ();
 sg13g2_decap_8 FILLER_12_819 ();
 sg13g2_decap_8 FILLER_12_826 ();
 sg13g2_decap_8 FILLER_12_833 ();
 sg13g2_decap_8 FILLER_12_840 ();
 sg13g2_decap_8 FILLER_12_847 ();
 sg13g2_decap_8 FILLER_12_854 ();
 sg13g2_decap_8 FILLER_12_861 ();
 sg13g2_decap_8 FILLER_12_868 ();
 sg13g2_fill_2 FILLER_12_875 ();
 sg13g2_fill_1 FILLER_12_877 ();
 sg13g2_decap_8 FILLER_13_0 ();
 sg13g2_decap_8 FILLER_13_7 ();
 sg13g2_decap_8 FILLER_13_14 ();
 sg13g2_decap_8 FILLER_13_21 ();
 sg13g2_decap_8 FILLER_13_28 ();
 sg13g2_decap_8 FILLER_13_35 ();
 sg13g2_decap_8 FILLER_13_42 ();
 sg13g2_decap_8 FILLER_13_49 ();
 sg13g2_decap_4 FILLER_13_56 ();
 sg13g2_decap_8 FILLER_13_64 ();
 sg13g2_fill_2 FILLER_13_71 ();
 sg13g2_fill_1 FILLER_13_79 ();
 sg13g2_decap_8 FILLER_13_98 ();
 sg13g2_decap_8 FILLER_13_105 ();
 sg13g2_fill_2 FILLER_13_112 ();
 sg13g2_fill_1 FILLER_13_119 ();
 sg13g2_fill_1 FILLER_13_124 ();
 sg13g2_decap_8 FILLER_13_151 ();
 sg13g2_fill_1 FILLER_13_158 ();
 sg13g2_decap_8 FILLER_13_171 ();
 sg13g2_decap_4 FILLER_13_178 ();
 sg13g2_decap_4 FILLER_13_209 ();
 sg13g2_fill_2 FILLER_13_229 ();
 sg13g2_decap_8 FILLER_13_247 ();
 sg13g2_decap_4 FILLER_13_254 ();
 sg13g2_fill_2 FILLER_13_275 ();
 sg13g2_fill_1 FILLER_13_289 ();
 sg13g2_fill_1 FILLER_13_295 ();
 sg13g2_decap_8 FILLER_13_301 ();
 sg13g2_fill_2 FILLER_13_308 ();
 sg13g2_fill_1 FILLER_13_310 ();
 sg13g2_decap_8 FILLER_13_323 ();
 sg13g2_decap_8 FILLER_13_330 ();
 sg13g2_decap_8 FILLER_13_337 ();
 sg13g2_fill_2 FILLER_13_344 ();
 sg13g2_fill_1 FILLER_13_346 ();
 sg13g2_decap_4 FILLER_13_362 ();
 sg13g2_decap_4 FILLER_13_378 ();
 sg13g2_fill_1 FILLER_13_382 ();
 sg13g2_fill_2 FILLER_13_388 ();
 sg13g2_fill_1 FILLER_13_390 ();
 sg13g2_fill_1 FILLER_13_394 ();
 sg13g2_fill_2 FILLER_13_421 ();
 sg13g2_fill_1 FILLER_13_426 ();
 sg13g2_decap_4 FILLER_13_459 ();
 sg13g2_fill_1 FILLER_13_463 ();
 sg13g2_fill_2 FILLER_13_474 ();
 sg13g2_fill_1 FILLER_13_476 ();
 sg13g2_fill_1 FILLER_13_481 ();
 sg13g2_fill_2 FILLER_13_491 ();
 sg13g2_fill_1 FILLER_13_493 ();
 sg13g2_fill_1 FILLER_13_503 ();
 sg13g2_decap_8 FILLER_13_508 ();
 sg13g2_decap_4 FILLER_13_515 ();
 sg13g2_fill_2 FILLER_13_519 ();
 sg13g2_fill_2 FILLER_13_552 ();
 sg13g2_decap_8 FILLER_13_559 ();
 sg13g2_decap_8 FILLER_13_566 ();
 sg13g2_decap_8 FILLER_13_573 ();
 sg13g2_fill_2 FILLER_13_580 ();
 sg13g2_fill_2 FILLER_13_599 ();
 sg13g2_fill_2 FILLER_13_619 ();
 sg13g2_fill_1 FILLER_13_621 ();
 sg13g2_decap_4 FILLER_13_627 ();
 sg13g2_fill_1 FILLER_13_631 ();
 sg13g2_fill_2 FILLER_13_640 ();
 sg13g2_fill_1 FILLER_13_642 ();
 sg13g2_decap_4 FILLER_13_651 ();
 sg13g2_fill_1 FILLER_13_655 ();
 sg13g2_decap_4 FILLER_13_660 ();
 sg13g2_fill_1 FILLER_13_664 ();
 sg13g2_fill_1 FILLER_13_670 ();
 sg13g2_fill_1 FILLER_13_677 ();
 sg13g2_fill_1 FILLER_13_682 ();
 sg13g2_fill_2 FILLER_13_692 ();
 sg13g2_fill_2 FILLER_13_699 ();
 sg13g2_fill_1 FILLER_13_701 ();
 sg13g2_decap_4 FILLER_13_707 ();
 sg13g2_fill_1 FILLER_13_711 ();
 sg13g2_decap_8 FILLER_13_716 ();
 sg13g2_decap_4 FILLER_13_723 ();
 sg13g2_fill_1 FILLER_13_727 ();
 sg13g2_fill_1 FILLER_13_767 ();
 sg13g2_decap_8 FILLER_13_773 ();
 sg13g2_decap_8 FILLER_13_780 ();
 sg13g2_decap_8 FILLER_13_787 ();
 sg13g2_decap_8 FILLER_13_794 ();
 sg13g2_decap_8 FILLER_13_801 ();
 sg13g2_decap_8 FILLER_13_808 ();
 sg13g2_decap_8 FILLER_13_815 ();
 sg13g2_decap_8 FILLER_13_822 ();
 sg13g2_decap_8 FILLER_13_829 ();
 sg13g2_decap_8 FILLER_13_836 ();
 sg13g2_decap_8 FILLER_13_843 ();
 sg13g2_decap_8 FILLER_13_850 ();
 sg13g2_decap_8 FILLER_13_857 ();
 sg13g2_decap_8 FILLER_13_864 ();
 sg13g2_decap_8 FILLER_13_871 ();
 sg13g2_decap_8 FILLER_14_0 ();
 sg13g2_decap_8 FILLER_14_7 ();
 sg13g2_decap_8 FILLER_14_14 ();
 sg13g2_decap_8 FILLER_14_21 ();
 sg13g2_decap_8 FILLER_14_28 ();
 sg13g2_decap_4 FILLER_14_35 ();
 sg13g2_fill_1 FILLER_14_39 ();
 sg13g2_fill_2 FILLER_14_45 ();
 sg13g2_fill_1 FILLER_14_47 ();
 sg13g2_fill_2 FILLER_14_68 ();
 sg13g2_decap_4 FILLER_14_106 ();
 sg13g2_fill_1 FILLER_14_110 ();
 sg13g2_decap_4 FILLER_14_123 ();
 sg13g2_fill_1 FILLER_14_127 ();
 sg13g2_decap_4 FILLER_14_138 ();
 sg13g2_fill_2 FILLER_14_142 ();
 sg13g2_fill_1 FILLER_14_151 ();
 sg13g2_fill_1 FILLER_14_160 ();
 sg13g2_fill_1 FILLER_14_169 ();
 sg13g2_fill_2 FILLER_14_181 ();
 sg13g2_fill_2 FILLER_14_187 ();
 sg13g2_decap_8 FILLER_14_202 ();
 sg13g2_fill_1 FILLER_14_209 ();
 sg13g2_fill_1 FILLER_14_224 ();
 sg13g2_fill_2 FILLER_14_230 ();
 sg13g2_decap_8 FILLER_14_248 ();
 sg13g2_fill_2 FILLER_14_255 ();
 sg13g2_fill_1 FILLER_14_257 ();
 sg13g2_fill_2 FILLER_14_271 ();
 sg13g2_fill_1 FILLER_14_273 ();
 sg13g2_fill_2 FILLER_14_294 ();
 sg13g2_fill_1 FILLER_14_296 ();
 sg13g2_decap_4 FILLER_14_307 ();
 sg13g2_fill_1 FILLER_14_311 ();
 sg13g2_decap_4 FILLER_14_316 ();
 sg13g2_fill_1 FILLER_14_320 ();
 sg13g2_fill_2 FILLER_14_360 ();
 sg13g2_decap_8 FILLER_14_367 ();
 sg13g2_fill_1 FILLER_14_374 ();
 sg13g2_decap_8 FILLER_14_380 ();
 sg13g2_fill_2 FILLER_14_387 ();
 sg13g2_fill_2 FILLER_14_393 ();
 sg13g2_decap_8 FILLER_14_409 ();
 sg13g2_decap_4 FILLER_14_416 ();
 sg13g2_fill_2 FILLER_14_420 ();
 sg13g2_fill_1 FILLER_14_444 ();
 sg13g2_fill_2 FILLER_14_449 ();
 sg13g2_fill_1 FILLER_14_455 ();
 sg13g2_fill_2 FILLER_14_461 ();
 sg13g2_fill_2 FILLER_14_495 ();
 sg13g2_fill_1 FILLER_14_500 ();
 sg13g2_fill_1 FILLER_14_506 ();
 sg13g2_decap_4 FILLER_14_512 ();
 sg13g2_fill_1 FILLER_14_516 ();
 sg13g2_fill_2 FILLER_14_521 ();
 sg13g2_fill_1 FILLER_14_523 ();
 sg13g2_fill_1 FILLER_14_547 ();
 sg13g2_decap_4 FILLER_14_560 ();
 sg13g2_fill_2 FILLER_14_569 ();
 sg13g2_decap_8 FILLER_14_575 ();
 sg13g2_fill_2 FILLER_14_582 ();
 sg13g2_fill_1 FILLER_14_619 ();
 sg13g2_fill_1 FILLER_14_624 ();
 sg13g2_decap_8 FILLER_14_630 ();
 sg13g2_fill_2 FILLER_14_637 ();
 sg13g2_decap_8 FILLER_14_647 ();
 sg13g2_decap_8 FILLER_14_692 ();
 sg13g2_fill_1 FILLER_14_699 ();
 sg13g2_fill_1 FILLER_14_705 ();
 sg13g2_decap_4 FILLER_14_722 ();
 sg13g2_fill_2 FILLER_14_726 ();
 sg13g2_fill_2 FILLER_14_736 ();
 sg13g2_fill_2 FILLER_14_754 ();
 sg13g2_fill_1 FILLER_14_756 ();
 sg13g2_decap_8 FILLER_14_762 ();
 sg13g2_decap_8 FILLER_14_769 ();
 sg13g2_decap_8 FILLER_14_776 ();
 sg13g2_decap_8 FILLER_14_783 ();
 sg13g2_decap_8 FILLER_14_790 ();
 sg13g2_decap_8 FILLER_14_797 ();
 sg13g2_decap_8 FILLER_14_804 ();
 sg13g2_decap_8 FILLER_14_811 ();
 sg13g2_decap_8 FILLER_14_818 ();
 sg13g2_decap_8 FILLER_14_825 ();
 sg13g2_decap_8 FILLER_14_832 ();
 sg13g2_decap_8 FILLER_14_839 ();
 sg13g2_decap_8 FILLER_14_846 ();
 sg13g2_decap_8 FILLER_14_853 ();
 sg13g2_decap_8 FILLER_14_860 ();
 sg13g2_decap_8 FILLER_14_867 ();
 sg13g2_decap_4 FILLER_14_874 ();
 sg13g2_decap_8 FILLER_15_0 ();
 sg13g2_decap_8 FILLER_15_7 ();
 sg13g2_decap_8 FILLER_15_14 ();
 sg13g2_decap_8 FILLER_15_21 ();
 sg13g2_decap_8 FILLER_15_28 ();
 sg13g2_fill_2 FILLER_15_35 ();
 sg13g2_fill_1 FILLER_15_37 ();
 sg13g2_fill_1 FILLER_15_46 ();
 sg13g2_fill_2 FILLER_15_55 ();
 sg13g2_decap_8 FILLER_15_65 ();
 sg13g2_decap_8 FILLER_15_72 ();
 sg13g2_decap_8 FILLER_15_79 ();
 sg13g2_decap_8 FILLER_15_86 ();
 sg13g2_decap_4 FILLER_15_93 ();
 sg13g2_fill_2 FILLER_15_97 ();
 sg13g2_fill_1 FILLER_15_103 ();
 sg13g2_fill_1 FILLER_15_109 ();
 sg13g2_decap_8 FILLER_15_118 ();
 sg13g2_fill_2 FILLER_15_129 ();
 sg13g2_fill_2 FILLER_15_162 ();
 sg13g2_fill_1 FILLER_15_173 ();
 sg13g2_fill_2 FILLER_15_188 ();
 sg13g2_fill_2 FILLER_15_208 ();
 sg13g2_fill_2 FILLER_15_223 ();
 sg13g2_decap_8 FILLER_15_238 ();
 sg13g2_fill_1 FILLER_15_245 ();
 sg13g2_fill_2 FILLER_15_256 ();
 sg13g2_decap_4 FILLER_15_264 ();
 sg13g2_fill_1 FILLER_15_268 ();
 sg13g2_fill_2 FILLER_15_298 ();
 sg13g2_decap_8 FILLER_15_315 ();
 sg13g2_decap_4 FILLER_15_322 ();
 sg13g2_fill_2 FILLER_15_326 ();
 sg13g2_fill_1 FILLER_15_347 ();
 sg13g2_fill_2 FILLER_15_358 ();
 sg13g2_decap_8 FILLER_15_391 ();
 sg13g2_fill_1 FILLER_15_398 ();
 sg13g2_decap_4 FILLER_15_405 ();
 sg13g2_fill_1 FILLER_15_409 ();
 sg13g2_fill_2 FILLER_15_414 ();
 sg13g2_fill_1 FILLER_15_416 ();
 sg13g2_decap_8 FILLER_15_422 ();
 sg13g2_fill_1 FILLER_15_429 ();
 sg13g2_fill_1 FILLER_15_441 ();
 sg13g2_fill_2 FILLER_15_455 ();
 sg13g2_fill_1 FILLER_15_461 ();
 sg13g2_fill_1 FILLER_15_467 ();
 sg13g2_fill_1 FILLER_15_473 ();
 sg13g2_fill_1 FILLER_15_479 ();
 sg13g2_fill_1 FILLER_15_496 ();
 sg13g2_fill_1 FILLER_15_502 ();
 sg13g2_fill_2 FILLER_15_510 ();
 sg13g2_decap_8 FILLER_15_526 ();
 sg13g2_decap_8 FILLER_15_533 ();
 sg13g2_fill_2 FILLER_15_540 ();
 sg13g2_fill_2 FILLER_15_547 ();
 sg13g2_fill_1 FILLER_15_554 ();
 sg13g2_fill_2 FILLER_15_584 ();
 sg13g2_fill_2 FILLER_15_590 ();
 sg13g2_fill_1 FILLER_15_592 ();
 sg13g2_decap_8 FILLER_15_605 ();
 sg13g2_decap_8 FILLER_15_612 ();
 sg13g2_decap_8 FILLER_15_619 ();
 sg13g2_decap_8 FILLER_15_626 ();
 sg13g2_decap_4 FILLER_15_633 ();
 sg13g2_fill_1 FILLER_15_645 ();
 sg13g2_fill_2 FILLER_15_650 ();
 sg13g2_decap_8 FILLER_15_660 ();
 sg13g2_decap_8 FILLER_15_667 ();
 sg13g2_fill_1 FILLER_15_674 ();
 sg13g2_fill_2 FILLER_15_680 ();
 sg13g2_fill_1 FILLER_15_682 ();
 sg13g2_fill_2 FILLER_15_688 ();
 sg13g2_fill_1 FILLER_15_690 ();
 sg13g2_decap_8 FILLER_15_725 ();
 sg13g2_decap_8 FILLER_15_732 ();
 sg13g2_fill_2 FILLER_15_739 ();
 sg13g2_decap_4 FILLER_15_753 ();
 sg13g2_fill_1 FILLER_15_757 ();
 sg13g2_decap_4 FILLER_15_762 ();
 sg13g2_fill_1 FILLER_15_766 ();
 sg13g2_fill_2 FILLER_15_772 ();
 sg13g2_fill_2 FILLER_15_778 ();
 sg13g2_fill_1 FILLER_15_780 ();
 sg13g2_decap_8 FILLER_15_785 ();
 sg13g2_decap_8 FILLER_15_792 ();
 sg13g2_decap_8 FILLER_15_799 ();
 sg13g2_decap_8 FILLER_15_806 ();
 sg13g2_decap_8 FILLER_15_813 ();
 sg13g2_decap_8 FILLER_15_820 ();
 sg13g2_decap_8 FILLER_15_827 ();
 sg13g2_decap_8 FILLER_15_834 ();
 sg13g2_decap_8 FILLER_15_841 ();
 sg13g2_decap_8 FILLER_15_848 ();
 sg13g2_decap_8 FILLER_15_855 ();
 sg13g2_decap_8 FILLER_15_862 ();
 sg13g2_decap_8 FILLER_15_869 ();
 sg13g2_fill_2 FILLER_15_876 ();
 sg13g2_decap_4 FILLER_16_0 ();
 sg13g2_fill_2 FILLER_16_7 ();
 sg13g2_fill_1 FILLER_16_9 ();
 sg13g2_decap_4 FILLER_16_25 ();
 sg13g2_fill_1 FILLER_16_41 ();
 sg13g2_fill_2 FILLER_16_55 ();
 sg13g2_fill_1 FILLER_16_57 ();
 sg13g2_decap_4 FILLER_16_74 ();
 sg13g2_fill_2 FILLER_16_110 ();
 sg13g2_fill_1 FILLER_16_112 ();
 sg13g2_fill_2 FILLER_16_126 ();
 sg13g2_fill_1 FILLER_16_141 ();
 sg13g2_decap_4 FILLER_16_146 ();
 sg13g2_fill_1 FILLER_16_150 ();
 sg13g2_fill_1 FILLER_16_155 ();
 sg13g2_fill_2 FILLER_16_165 ();
 sg13g2_fill_2 FILLER_16_172 ();
 sg13g2_fill_1 FILLER_16_174 ();
 sg13g2_fill_1 FILLER_16_183 ();
 sg13g2_fill_2 FILLER_16_193 ();
 sg13g2_fill_1 FILLER_16_195 ();
 sg13g2_fill_1 FILLER_16_214 ();
 sg13g2_fill_2 FILLER_16_223 ();
 sg13g2_fill_2 FILLER_16_236 ();
 sg13g2_decap_4 FILLER_16_242 ();
 sg13g2_fill_2 FILLER_16_274 ();
 sg13g2_fill_2 FILLER_16_280 ();
 sg13g2_fill_2 FILLER_16_287 ();
 sg13g2_fill_2 FILLER_16_314 ();
 sg13g2_fill_1 FILLER_16_316 ();
 sg13g2_decap_8 FILLER_16_322 ();
 sg13g2_fill_2 FILLER_16_329 ();
 sg13g2_fill_1 FILLER_16_331 ();
 sg13g2_decap_4 FILLER_16_342 ();
 sg13g2_fill_1 FILLER_16_358 ();
 sg13g2_fill_2 FILLER_16_364 ();
 sg13g2_fill_1 FILLER_16_366 ();
 sg13g2_decap_8 FILLER_16_384 ();
 sg13g2_decap_8 FILLER_16_409 ();
 sg13g2_fill_2 FILLER_16_429 ();
 sg13g2_fill_2 FILLER_16_434 ();
 sg13g2_fill_1 FILLER_16_436 ();
 sg13g2_fill_2 FILLER_16_455 ();
 sg13g2_fill_1 FILLER_16_475 ();
 sg13g2_fill_2 FILLER_16_500 ();
 sg13g2_decap_8 FILLER_16_508 ();
 sg13g2_fill_1 FILLER_16_515 ();
 sg13g2_fill_2 FILLER_16_525 ();
 sg13g2_fill_1 FILLER_16_527 ();
 sg13g2_fill_1 FILLER_16_537 ();
 sg13g2_fill_2 FILLER_16_548 ();
 sg13g2_fill_1 FILLER_16_554 ();
 sg13g2_decap_4 FILLER_16_559 ();
 sg13g2_fill_1 FILLER_16_563 ();
 sg13g2_fill_1 FILLER_16_569 ();
 sg13g2_fill_2 FILLER_16_607 ();
 sg13g2_decap_8 FILLER_16_632 ();
 sg13g2_fill_1 FILLER_16_639 ();
 sg13g2_fill_1 FILLER_16_648 ();
 sg13g2_fill_2 FILLER_16_659 ();
 sg13g2_fill_1 FILLER_16_666 ();
 sg13g2_fill_1 FILLER_16_674 ();
 sg13g2_fill_2 FILLER_16_704 ();
 sg13g2_decap_4 FILLER_16_713 ();
 sg13g2_fill_2 FILLER_16_721 ();
 sg13g2_fill_1 FILLER_16_723 ();
 sg13g2_fill_2 FILLER_16_728 ();
 sg13g2_fill_1 FILLER_16_730 ();
 sg13g2_fill_1 FILLER_16_747 ();
 sg13g2_fill_2 FILLER_16_769 ();
 sg13g2_fill_1 FILLER_16_775 ();
 sg13g2_decap_4 FILLER_16_801 ();
 sg13g2_fill_1 FILLER_16_805 ();
 sg13g2_decap_8 FILLER_16_810 ();
 sg13g2_decap_8 FILLER_16_835 ();
 sg13g2_decap_8 FILLER_16_842 ();
 sg13g2_decap_8 FILLER_16_849 ();
 sg13g2_decap_8 FILLER_16_856 ();
 sg13g2_decap_8 FILLER_16_863 ();
 sg13g2_decap_8 FILLER_16_870 ();
 sg13g2_fill_1 FILLER_16_877 ();
 sg13g2_decap_4 FILLER_17_0 ();
 sg13g2_fill_2 FILLER_17_30 ();
 sg13g2_fill_1 FILLER_17_32 ();
 sg13g2_fill_1 FILLER_17_45 ();
 sg13g2_decap_4 FILLER_17_62 ();
 sg13g2_fill_1 FILLER_17_66 ();
 sg13g2_fill_2 FILLER_17_76 ();
 sg13g2_decap_4 FILLER_17_103 ();
 sg13g2_fill_1 FILLER_17_107 ();
 sg13g2_fill_1 FILLER_17_121 ();
 sg13g2_decap_4 FILLER_17_134 ();
 sg13g2_fill_2 FILLER_17_138 ();
 sg13g2_fill_2 FILLER_17_144 ();
 sg13g2_fill_1 FILLER_17_146 ();
 sg13g2_fill_1 FILLER_17_169 ();
 sg13g2_fill_2 FILLER_17_174 ();
 sg13g2_decap_4 FILLER_17_181 ();
 sg13g2_fill_1 FILLER_17_195 ();
 sg13g2_fill_2 FILLER_17_215 ();
 sg13g2_decap_4 FILLER_17_234 ();
 sg13g2_fill_2 FILLER_17_238 ();
 sg13g2_fill_1 FILLER_17_254 ();
 sg13g2_fill_1 FILLER_17_273 ();
 sg13g2_fill_1 FILLER_17_283 ();
 sg13g2_fill_1 FILLER_17_289 ();
 sg13g2_fill_1 FILLER_17_312 ();
 sg13g2_decap_4 FILLER_17_325 ();
 sg13g2_fill_2 FILLER_17_334 ();
 sg13g2_fill_2 FILLER_17_340 ();
 sg13g2_fill_1 FILLER_17_342 ();
 sg13g2_fill_1 FILLER_17_347 ();
 sg13g2_fill_2 FILLER_17_378 ();
 sg13g2_decap_4 FILLER_17_384 ();
 sg13g2_fill_2 FILLER_17_393 ();
 sg13g2_decap_4 FILLER_17_402 ();
 sg13g2_fill_2 FILLER_17_429 ();
 sg13g2_decap_4 FILLER_17_435 ();
 sg13g2_fill_1 FILLER_17_439 ();
 sg13g2_fill_2 FILLER_17_445 ();
 sg13g2_fill_1 FILLER_17_451 ();
 sg13g2_fill_2 FILLER_17_456 ();
 sg13g2_decap_8 FILLER_17_462 ();
 sg13g2_decap_4 FILLER_17_474 ();
 sg13g2_fill_1 FILLER_17_478 ();
 sg13g2_decap_4 FILLER_17_484 ();
 sg13g2_fill_1 FILLER_17_488 ();
 sg13g2_fill_1 FILLER_17_518 ();
 sg13g2_fill_1 FILLER_17_531 ();
 sg13g2_fill_1 FILLER_17_545 ();
 sg13g2_fill_2 FILLER_17_561 ();
 sg13g2_fill_1 FILLER_17_563 ();
 sg13g2_fill_1 FILLER_17_569 ();
 sg13g2_fill_2 FILLER_17_579 ();
 sg13g2_fill_1 FILLER_17_581 ();
 sg13g2_fill_2 FILLER_17_603 ();
 sg13g2_fill_1 FILLER_17_609 ();
 sg13g2_decap_8 FILLER_17_631 ();
 sg13g2_decap_4 FILLER_17_648 ();
 sg13g2_fill_2 FILLER_17_665 ();
 sg13g2_fill_1 FILLER_17_692 ();
 sg13g2_fill_1 FILLER_17_698 ();
 sg13g2_fill_1 FILLER_17_706 ();
 sg13g2_fill_1 FILLER_17_721 ();
 sg13g2_decap_8 FILLER_17_727 ();
 sg13g2_decap_4 FILLER_17_734 ();
 sg13g2_fill_2 FILLER_17_738 ();
 sg13g2_fill_1 FILLER_17_753 ();
 sg13g2_decap_4 FILLER_17_759 ();
 sg13g2_fill_1 FILLER_17_763 ();
 sg13g2_fill_2 FILLER_17_772 ();
 sg13g2_fill_1 FILLER_17_774 ();
 sg13g2_fill_2 FILLER_17_793 ();
 sg13g2_fill_1 FILLER_17_795 ();
 sg13g2_fill_1 FILLER_17_804 ();
 sg13g2_decap_8 FILLER_17_810 ();
 sg13g2_decap_4 FILLER_17_817 ();
 sg13g2_fill_1 FILLER_17_821 ();
 sg13g2_decap_8 FILLER_17_835 ();
 sg13g2_decap_8 FILLER_17_842 ();
 sg13g2_decap_8 FILLER_17_849 ();
 sg13g2_decap_8 FILLER_17_856 ();
 sg13g2_decap_8 FILLER_17_863 ();
 sg13g2_decap_8 FILLER_17_870 ();
 sg13g2_fill_1 FILLER_17_877 ();
 sg13g2_decap_8 FILLER_18_0 ();
 sg13g2_fill_1 FILLER_18_7 ();
 sg13g2_decap_8 FILLER_18_24 ();
 sg13g2_fill_2 FILLER_18_38 ();
 sg13g2_fill_1 FILLER_18_40 ();
 sg13g2_decap_4 FILLER_18_49 ();
 sg13g2_fill_1 FILLER_18_53 ();
 sg13g2_decap_8 FILLER_18_58 ();
 sg13g2_fill_2 FILLER_18_82 ();
 sg13g2_fill_1 FILLER_18_84 ();
 sg13g2_fill_2 FILLER_18_114 ();
 sg13g2_fill_2 FILLER_18_132 ();
 sg13g2_fill_1 FILLER_18_134 ();
 sg13g2_decap_8 FILLER_18_143 ();
 sg13g2_decap_4 FILLER_18_150 ();
 sg13g2_fill_2 FILLER_18_154 ();
 sg13g2_decap_8 FILLER_18_164 ();
 sg13g2_fill_2 FILLER_18_171 ();
 sg13g2_fill_2 FILLER_18_182 ();
 sg13g2_fill_1 FILLER_18_189 ();
 sg13g2_decap_8 FILLER_18_209 ();
 sg13g2_decap_4 FILLER_18_216 ();
 sg13g2_fill_2 FILLER_18_220 ();
 sg13g2_fill_2 FILLER_18_249 ();
 sg13g2_decap_4 FILLER_18_264 ();
 sg13g2_fill_1 FILLER_18_276 ();
 sg13g2_fill_2 FILLER_18_285 ();
 sg13g2_fill_2 FILLER_18_292 ();
 sg13g2_fill_1 FILLER_18_298 ();
 sg13g2_decap_8 FILLER_18_311 ();
 sg13g2_fill_2 FILLER_18_318 ();
 sg13g2_fill_1 FILLER_18_324 ();
 sg13g2_fill_2 FILLER_18_339 ();
 sg13g2_decap_8 FILLER_18_351 ();
 sg13g2_fill_2 FILLER_18_358 ();
 sg13g2_fill_2 FILLER_18_378 ();
 sg13g2_fill_1 FILLER_18_406 ();
 sg13g2_decap_8 FILLER_18_454 ();
 sg13g2_fill_2 FILLER_18_461 ();
 sg13g2_fill_1 FILLER_18_463 ();
 sg13g2_fill_1 FILLER_18_494 ();
 sg13g2_fill_1 FILLER_18_501 ();
 sg13g2_fill_1 FILLER_18_519 ();
 sg13g2_decap_4 FILLER_18_525 ();
 sg13g2_fill_1 FILLER_18_549 ();
 sg13g2_fill_2 FILLER_18_566 ();
 sg13g2_fill_2 FILLER_18_574 ();
 sg13g2_fill_2 FILLER_18_581 ();
 sg13g2_fill_2 FILLER_18_595 ();
 sg13g2_fill_1 FILLER_18_597 ();
 sg13g2_fill_1 FILLER_18_612 ();
 sg13g2_decap_4 FILLER_18_644 ();
 sg13g2_fill_2 FILLER_18_661 ();
 sg13g2_fill_2 FILLER_18_666 ();
 sg13g2_fill_1 FILLER_18_683 ();
 sg13g2_fill_1 FILLER_18_694 ();
 sg13g2_fill_2 FILLER_18_704 ();
 sg13g2_fill_1 FILLER_18_706 ();
 sg13g2_decap_4 FILLER_18_712 ();
 sg13g2_decap_4 FILLER_18_721 ();
 sg13g2_fill_1 FILLER_18_725 ();
 sg13g2_fill_2 FILLER_18_731 ();
 sg13g2_fill_1 FILLER_18_733 ();
 sg13g2_decap_4 FILLER_18_739 ();
 sg13g2_fill_1 FILLER_18_743 ();
 sg13g2_decap_4 FILLER_18_774 ();
 sg13g2_fill_2 FILLER_18_803 ();
 sg13g2_fill_1 FILLER_18_805 ();
 sg13g2_fill_1 FILLER_18_810 ();
 sg13g2_fill_2 FILLER_18_816 ();
 sg13g2_decap_8 FILLER_18_823 ();
 sg13g2_fill_2 FILLER_18_830 ();
 sg13g2_fill_1 FILLER_18_832 ();
 sg13g2_decap_8 FILLER_18_841 ();
 sg13g2_decap_8 FILLER_18_848 ();
 sg13g2_decap_8 FILLER_18_855 ();
 sg13g2_decap_8 FILLER_18_862 ();
 sg13g2_decap_8 FILLER_18_869 ();
 sg13g2_fill_2 FILLER_18_876 ();
 sg13g2_fill_2 FILLER_19_20 ();
 sg13g2_decap_8 FILLER_19_30 ();
 sg13g2_fill_2 FILLER_19_37 ();
 sg13g2_fill_1 FILLER_19_39 ();
 sg13g2_decap_4 FILLER_19_45 ();
 sg13g2_fill_1 FILLER_19_54 ();
 sg13g2_fill_1 FILLER_19_68 ();
 sg13g2_fill_1 FILLER_19_75 ();
 sg13g2_fill_1 FILLER_19_81 ();
 sg13g2_fill_1 FILLER_19_99 ();
 sg13g2_fill_2 FILLER_19_105 ();
 sg13g2_fill_2 FILLER_19_111 ();
 sg13g2_fill_2 FILLER_19_117 ();
 sg13g2_fill_1 FILLER_19_131 ();
 sg13g2_decap_4 FILLER_19_144 ();
 sg13g2_fill_2 FILLER_19_214 ();
 sg13g2_fill_1 FILLER_19_221 ();
 sg13g2_fill_1 FILLER_19_226 ();
 sg13g2_fill_1 FILLER_19_235 ();
 sg13g2_fill_1 FILLER_19_257 ();
 sg13g2_fill_1 FILLER_19_262 ();
 sg13g2_decap_4 FILLER_19_275 ();
 sg13g2_fill_1 FILLER_19_284 ();
 sg13g2_decap_4 FILLER_19_290 ();
 sg13g2_decap_4 FILLER_19_298 ();
 sg13g2_decap_8 FILLER_19_306 ();
 sg13g2_fill_2 FILLER_19_313 ();
 sg13g2_fill_1 FILLER_19_315 ();
 sg13g2_fill_2 FILLER_19_362 ();
 sg13g2_fill_1 FILLER_19_372 ();
 sg13g2_fill_2 FILLER_19_428 ();
 sg13g2_decap_8 FILLER_19_438 ();
 sg13g2_fill_2 FILLER_19_445 ();
 sg13g2_fill_1 FILLER_19_447 ();
 sg13g2_decap_8 FILLER_19_452 ();
 sg13g2_decap_8 FILLER_19_459 ();
 sg13g2_decap_8 FILLER_19_466 ();
 sg13g2_fill_2 FILLER_19_473 ();
 sg13g2_decap_8 FILLER_19_479 ();
 sg13g2_fill_2 FILLER_19_486 ();
 sg13g2_fill_1 FILLER_19_488 ();
 sg13g2_fill_2 FILLER_19_503 ();
 sg13g2_fill_1 FILLER_19_523 ();
 sg13g2_fill_2 FILLER_19_529 ();
 sg13g2_fill_1 FILLER_19_531 ();
 sg13g2_fill_2 FILLER_19_554 ();
 sg13g2_fill_2 FILLER_19_561 ();
 sg13g2_fill_1 FILLER_19_563 ();
 sg13g2_fill_1 FILLER_19_574 ();
 sg13g2_fill_2 FILLER_19_589 ();
 sg13g2_fill_1 FILLER_19_591 ();
 sg13g2_fill_2 FILLER_19_596 ();
 sg13g2_fill_1 FILLER_19_598 ();
 sg13g2_decap_4 FILLER_19_603 ();
 sg13g2_fill_1 FILLER_19_607 ();
 sg13g2_fill_1 FILLER_19_627 ();
 sg13g2_fill_1 FILLER_19_633 ();
 sg13g2_decap_4 FILLER_19_639 ();
 sg13g2_fill_1 FILLER_19_643 ();
 sg13g2_fill_2 FILLER_19_654 ();
 sg13g2_fill_2 FILLER_19_667 ();
 sg13g2_decap_8 FILLER_19_705 ();
 sg13g2_fill_2 FILLER_19_738 ();
 sg13g2_fill_1 FILLER_19_740 ();
 sg13g2_fill_2 FILLER_19_745 ();
 sg13g2_fill_2 FILLER_19_752 ();
 sg13g2_fill_1 FILLER_19_754 ();
 sg13g2_fill_1 FILLER_19_760 ();
 sg13g2_decap_8 FILLER_19_782 ();
 sg13g2_fill_2 FILLER_19_789 ();
 sg13g2_fill_1 FILLER_19_795 ();
 sg13g2_fill_1 FILLER_19_803 ();
 sg13g2_fill_1 FILLER_19_824 ();
 sg13g2_fill_2 FILLER_19_829 ();
 sg13g2_fill_1 FILLER_19_836 ();
 sg13g2_decap_8 FILLER_19_845 ();
 sg13g2_decap_8 FILLER_19_852 ();
 sg13g2_decap_8 FILLER_19_859 ();
 sg13g2_decap_8 FILLER_19_866 ();
 sg13g2_decap_4 FILLER_19_873 ();
 sg13g2_fill_1 FILLER_19_877 ();
 sg13g2_decap_8 FILLER_20_16 ();
 sg13g2_fill_2 FILLER_20_23 ();
 sg13g2_fill_1 FILLER_20_25 ();
 sg13g2_decap_4 FILLER_20_30 ();
 sg13g2_fill_1 FILLER_20_42 ();
 sg13g2_fill_2 FILLER_20_79 ();
 sg13g2_fill_2 FILLER_20_86 ();
 sg13g2_fill_2 FILLER_20_93 ();
 sg13g2_fill_1 FILLER_20_99 ();
 sg13g2_fill_1 FILLER_20_105 ();
 sg13g2_fill_1 FILLER_20_110 ();
 sg13g2_fill_1 FILLER_20_116 ();
 sg13g2_fill_1 FILLER_20_121 ();
 sg13g2_fill_1 FILLER_20_131 ();
 sg13g2_decap_8 FILLER_20_137 ();
 sg13g2_decap_8 FILLER_20_144 ();
 sg13g2_fill_2 FILLER_20_151 ();
 sg13g2_fill_1 FILLER_20_153 ();
 sg13g2_decap_8 FILLER_20_187 ();
 sg13g2_decap_4 FILLER_20_194 ();
 sg13g2_fill_2 FILLER_20_198 ();
 sg13g2_fill_2 FILLER_20_204 ();
 sg13g2_fill_1 FILLER_20_206 ();
 sg13g2_fill_2 FILLER_20_214 ();
 sg13g2_decap_8 FILLER_20_248 ();
 sg13g2_decap_8 FILLER_20_272 ();
 sg13g2_fill_2 FILLER_20_279 ();
 sg13g2_fill_1 FILLER_20_281 ();
 sg13g2_decap_4 FILLER_20_304 ();
 sg13g2_fill_1 FILLER_20_308 ();
 sg13g2_fill_2 FILLER_20_327 ();
 sg13g2_fill_1 FILLER_20_329 ();
 sg13g2_decap_8 FILLER_20_334 ();
 sg13g2_decap_8 FILLER_20_341 ();
 sg13g2_fill_2 FILLER_20_348 ();
 sg13g2_fill_1 FILLER_20_350 ();
 sg13g2_fill_2 FILLER_20_384 ();
 sg13g2_decap_4 FILLER_20_454 ();
 sg13g2_fill_2 FILLER_20_551 ();
 sg13g2_decap_8 FILLER_20_594 ();
 sg13g2_decap_4 FILLER_20_601 ();
 sg13g2_fill_1 FILLER_20_605 ();
 sg13g2_fill_1 FILLER_20_611 ();
 sg13g2_fill_2 FILLER_20_616 ();
 sg13g2_fill_2 FILLER_20_621 ();
 sg13g2_fill_2 FILLER_20_628 ();
 sg13g2_decap_8 FILLER_20_634 ();
 sg13g2_fill_2 FILLER_20_641 ();
 sg13g2_fill_2 FILLER_20_647 ();
 sg13g2_fill_1 FILLER_20_649 ();
 sg13g2_fill_1 FILLER_20_661 ();
 sg13g2_fill_1 FILLER_20_672 ();
 sg13g2_fill_1 FILLER_20_683 ();
 sg13g2_fill_2 FILLER_20_694 ();
 sg13g2_fill_1 FILLER_20_696 ();
 sg13g2_decap_4 FILLER_20_706 ();
 sg13g2_fill_1 FILLER_20_716 ();
 sg13g2_fill_2 FILLER_20_733 ();
 sg13g2_fill_2 FILLER_20_739 ();
 sg13g2_fill_2 FILLER_20_746 ();
 sg13g2_decap_8 FILLER_20_755 ();
 sg13g2_fill_2 FILLER_20_762 ();
 sg13g2_fill_1 FILLER_20_764 ();
 sg13g2_decap_8 FILLER_20_773 ();
 sg13g2_decap_8 FILLER_20_790 ();
 sg13g2_fill_1 FILLER_20_797 ();
 sg13g2_fill_2 FILLER_20_803 ();
 sg13g2_fill_1 FILLER_20_809 ();
 sg13g2_fill_1 FILLER_20_816 ();
 sg13g2_fill_1 FILLER_20_822 ();
 sg13g2_fill_1 FILLER_20_831 ();
 sg13g2_decap_8 FILLER_20_836 ();
 sg13g2_fill_2 FILLER_20_843 ();
 sg13g2_fill_1 FILLER_20_845 ();
 sg13g2_fill_1 FILLER_20_858 ();
 sg13g2_decap_8 FILLER_20_863 ();
 sg13g2_decap_8 FILLER_20_870 ();
 sg13g2_fill_1 FILLER_20_877 ();
 sg13g2_decap_4 FILLER_21_14 ();
 sg13g2_fill_1 FILLER_21_18 ();
 sg13g2_decap_8 FILLER_21_28 ();
 sg13g2_decap_4 FILLER_21_35 ();
 sg13g2_fill_2 FILLER_21_47 ();
 sg13g2_fill_2 FILLER_21_57 ();
 sg13g2_fill_1 FILLER_21_59 ();
 sg13g2_decap_8 FILLER_21_79 ();
 sg13g2_decap_4 FILLER_21_90 ();
 sg13g2_decap_8 FILLER_21_98 ();
 sg13g2_decap_4 FILLER_21_105 ();
 sg13g2_fill_2 FILLER_21_117 ();
 sg13g2_fill_1 FILLER_21_132 ();
 sg13g2_fill_1 FILLER_21_142 ();
 sg13g2_fill_1 FILLER_21_148 ();
 sg13g2_decap_4 FILLER_21_190 ();
 sg13g2_decap_4 FILLER_21_198 ();
 sg13g2_fill_1 FILLER_21_202 ();
 sg13g2_fill_2 FILLER_21_216 ();
 sg13g2_fill_1 FILLER_21_218 ();
 sg13g2_fill_2 FILLER_21_233 ();
 sg13g2_decap_4 FILLER_21_264 ();
 sg13g2_fill_2 FILLER_21_276 ();
 sg13g2_decap_4 FILLER_21_310 ();
 sg13g2_fill_1 FILLER_21_314 ();
 sg13g2_decap_8 FILLER_21_324 ();
 sg13g2_fill_1 FILLER_21_331 ();
 sg13g2_fill_2 FILLER_21_337 ();
 sg13g2_fill_2 FILLER_21_367 ();
 sg13g2_fill_2 FILLER_21_374 ();
 sg13g2_decap_4 FILLER_21_391 ();
 sg13g2_fill_1 FILLER_21_407 ();
 sg13g2_decap_8 FILLER_21_447 ();
 sg13g2_fill_2 FILLER_21_454 ();
 sg13g2_decap_8 FILLER_21_461 ();
 sg13g2_fill_1 FILLER_21_481 ();
 sg13g2_fill_2 FILLER_21_486 ();
 sg13g2_fill_1 FILLER_21_488 ();
 sg13g2_fill_2 FILLER_21_494 ();
 sg13g2_decap_4 FILLER_21_513 ();
 sg13g2_fill_2 FILLER_21_525 ();
 sg13g2_fill_1 FILLER_21_532 ();
 sg13g2_fill_1 FILLER_21_556 ();
 sg13g2_fill_2 FILLER_21_562 ();
 sg13g2_decap_4 FILLER_21_568 ();
 sg13g2_fill_1 FILLER_21_572 ();
 sg13g2_decap_4 FILLER_21_585 ();
 sg13g2_decap_8 FILLER_21_594 ();
 sg13g2_decap_8 FILLER_21_601 ();
 sg13g2_decap_4 FILLER_21_608 ();
 sg13g2_fill_1 FILLER_21_621 ();
 sg13g2_fill_2 FILLER_21_627 ();
 sg13g2_decap_8 FILLER_21_634 ();
 sg13g2_fill_2 FILLER_21_653 ();
 sg13g2_fill_2 FILLER_21_660 ();
 sg13g2_fill_2 FILLER_21_671 ();
 sg13g2_decap_8 FILLER_21_698 ();
 sg13g2_fill_2 FILLER_21_713 ();
 sg13g2_fill_1 FILLER_21_715 ();
 sg13g2_decap_8 FILLER_21_721 ();
 sg13g2_fill_2 FILLER_21_728 ();
 sg13g2_fill_1 FILLER_21_734 ();
 sg13g2_decap_4 FILLER_21_740 ();
 sg13g2_fill_1 FILLER_21_744 ();
 sg13g2_fill_1 FILLER_21_770 ();
 sg13g2_fill_2 FILLER_21_776 ();
 sg13g2_fill_2 FILLER_21_782 ();
 sg13g2_fill_1 FILLER_21_788 ();
 sg13g2_fill_2 FILLER_21_795 ();
 sg13g2_decap_4 FILLER_21_801 ();
 sg13g2_fill_2 FILLER_21_805 ();
 sg13g2_decap_4 FILLER_21_818 ();
 sg13g2_fill_1 FILLER_21_822 ();
 sg13g2_fill_1 FILLER_21_841 ();
 sg13g2_fill_2 FILLER_21_847 ();
 sg13g2_fill_1 FILLER_21_849 ();
 sg13g2_fill_2 FILLER_21_855 ();
 sg13g2_fill_1 FILLER_21_857 ();
 sg13g2_decap_8 FILLER_21_871 ();
 sg13g2_fill_1 FILLER_22_0 ();
 sg13g2_decap_4 FILLER_22_10 ();
 sg13g2_fill_1 FILLER_22_14 ();
 sg13g2_decap_8 FILLER_22_23 ();
 sg13g2_fill_2 FILLER_22_30 ();
 sg13g2_fill_2 FILLER_22_48 ();
 sg13g2_fill_1 FILLER_22_50 ();
 sg13g2_fill_1 FILLER_22_81 ();
 sg13g2_decap_8 FILLER_22_86 ();
 sg13g2_decap_8 FILLER_22_93 ();
 sg13g2_fill_2 FILLER_22_100 ();
 sg13g2_fill_2 FILLER_22_122 ();
 sg13g2_fill_2 FILLER_22_132 ();
 sg13g2_fill_1 FILLER_22_156 ();
 sg13g2_decap_4 FILLER_22_180 ();
 sg13g2_fill_2 FILLER_22_188 ();
 sg13g2_fill_1 FILLER_22_190 ();
 sg13g2_fill_2 FILLER_22_195 ();
 sg13g2_fill_1 FILLER_22_197 ();
 sg13g2_fill_2 FILLER_22_201 ();
 sg13g2_fill_1 FILLER_22_203 ();
 sg13g2_fill_1 FILLER_22_226 ();
 sg13g2_decap_8 FILLER_22_243 ();
 sg13g2_fill_1 FILLER_22_255 ();
 sg13g2_fill_2 FILLER_22_274 ();
 sg13g2_fill_2 FILLER_22_292 ();
 sg13g2_fill_2 FILLER_22_304 ();
 sg13g2_fill_1 FILLER_22_319 ();
 sg13g2_decap_8 FILLER_22_371 ();
 sg13g2_fill_2 FILLER_22_378 ();
 sg13g2_fill_1 FILLER_22_380 ();
 sg13g2_fill_2 FILLER_22_399 ();
 sg13g2_fill_1 FILLER_22_401 ();
 sg13g2_decap_4 FILLER_22_412 ();
 sg13g2_fill_2 FILLER_22_416 ();
 sg13g2_fill_1 FILLER_22_443 ();
 sg13g2_decap_4 FILLER_22_460 ();
 sg13g2_fill_2 FILLER_22_464 ();
 sg13g2_fill_2 FILLER_22_475 ();
 sg13g2_fill_1 FILLER_22_477 ();
 sg13g2_fill_1 FILLER_22_495 ();
 sg13g2_fill_2 FILLER_22_504 ();
 sg13g2_fill_2 FILLER_22_511 ();
 sg13g2_decap_4 FILLER_22_527 ();
 sg13g2_fill_1 FILLER_22_531 ();
 sg13g2_decap_4 FILLER_22_540 ();
 sg13g2_fill_1 FILLER_22_567 ();
 sg13g2_fill_1 FILLER_22_577 ();
 sg13g2_fill_1 FILLER_22_582 ();
 sg13g2_decap_8 FILLER_22_588 ();
 sg13g2_decap_4 FILLER_22_595 ();
 sg13g2_fill_2 FILLER_22_604 ();
 sg13g2_fill_1 FILLER_22_613 ();
 sg13g2_fill_1 FILLER_22_631 ();
 sg13g2_decap_4 FILLER_22_637 ();
 sg13g2_fill_1 FILLER_22_678 ();
 sg13g2_decap_8 FILLER_22_688 ();
 sg13g2_fill_1 FILLER_22_695 ();
 sg13g2_fill_2 FILLER_22_727 ();
 sg13g2_fill_1 FILLER_22_734 ();
 sg13g2_fill_1 FILLER_22_739 ();
 sg13g2_fill_1 FILLER_22_744 ();
 sg13g2_fill_1 FILLER_22_750 ();
 sg13g2_fill_1 FILLER_22_755 ();
 sg13g2_fill_2 FILLER_22_765 ();
 sg13g2_fill_2 FILLER_22_776 ();
 sg13g2_fill_1 FILLER_22_808 ();
 sg13g2_fill_1 FILLER_22_813 ();
 sg13g2_fill_2 FILLER_22_819 ();
 sg13g2_decap_8 FILLER_22_834 ();
 sg13g2_decap_8 FILLER_22_845 ();
 sg13g2_fill_2 FILLER_22_857 ();
 sg13g2_decap_8 FILLER_22_870 ();
 sg13g2_fill_1 FILLER_22_877 ();
 sg13g2_fill_2 FILLER_23_0 ();
 sg13g2_fill_2 FILLER_23_15 ();
 sg13g2_fill_2 FILLER_23_26 ();
 sg13g2_fill_1 FILLER_23_28 ();
 sg13g2_fill_2 FILLER_23_41 ();
 sg13g2_fill_1 FILLER_23_43 ();
 sg13g2_fill_1 FILLER_23_52 ();
 sg13g2_fill_2 FILLER_23_58 ();
 sg13g2_fill_1 FILLER_23_68 ();
 sg13g2_fill_1 FILLER_23_77 ();
 sg13g2_fill_2 FILLER_23_102 ();
 sg13g2_fill_1 FILLER_23_109 ();
 sg13g2_fill_2 FILLER_23_114 ();
 sg13g2_fill_1 FILLER_23_116 ();
 sg13g2_fill_2 FILLER_23_130 ();
 sg13g2_decap_4 FILLER_23_146 ();
 sg13g2_fill_1 FILLER_23_150 ();
 sg13g2_fill_2 FILLER_23_182 ();
 sg13g2_decap_8 FILLER_23_188 ();
 sg13g2_decap_4 FILLER_23_195 ();
 sg13g2_fill_1 FILLER_23_199 ();
 sg13g2_fill_1 FILLER_23_222 ();
 sg13g2_decap_4 FILLER_23_227 ();
 sg13g2_fill_1 FILLER_23_231 ();
 sg13g2_decap_4 FILLER_23_242 ();
 sg13g2_fill_1 FILLER_23_246 ();
 sg13g2_fill_1 FILLER_23_265 ();
 sg13g2_fill_2 FILLER_23_271 ();
 sg13g2_fill_1 FILLER_23_308 ();
 sg13g2_fill_1 FILLER_23_328 ();
 sg13g2_fill_1 FILLER_23_337 ();
 sg13g2_fill_2 FILLER_23_347 ();
 sg13g2_fill_1 FILLER_23_358 ();
 sg13g2_fill_1 FILLER_23_364 ();
 sg13g2_fill_1 FILLER_23_383 ();
 sg13g2_fill_2 FILLER_23_389 ();
 sg13g2_fill_1 FILLER_23_391 ();
 sg13g2_fill_1 FILLER_23_405 ();
 sg13g2_decap_8 FILLER_23_411 ();
 sg13g2_fill_1 FILLER_23_427 ();
 sg13g2_fill_2 FILLER_23_454 ();
 sg13g2_decap_4 FILLER_23_461 ();
 sg13g2_fill_1 FILLER_23_465 ();
 sg13g2_decap_4 FILLER_23_490 ();
 sg13g2_fill_1 FILLER_23_508 ();
 sg13g2_fill_1 FILLER_23_519 ();
 sg13g2_decap_4 FILLER_23_535 ();
 sg13g2_fill_1 FILLER_23_544 ();
 sg13g2_fill_2 FILLER_23_550 ();
 sg13g2_fill_1 FILLER_23_565 ();
 sg13g2_fill_1 FILLER_23_570 ();
 sg13g2_fill_2 FILLER_23_576 ();
 sg13g2_fill_2 FILLER_23_595 ();
 sg13g2_fill_1 FILLER_23_602 ();
 sg13g2_fill_1 FILLER_23_620 ();
 sg13g2_decap_4 FILLER_23_643 ();
 sg13g2_fill_1 FILLER_23_647 ();
 sg13g2_fill_2 FILLER_23_664 ();
 sg13g2_fill_1 FILLER_23_666 ();
 sg13g2_decap_8 FILLER_23_672 ();
 sg13g2_decap_8 FILLER_23_679 ();
 sg13g2_decap_4 FILLER_23_686 ();
 sg13g2_decap_8 FILLER_23_718 ();
 sg13g2_fill_1 FILLER_23_725 ();
 sg13g2_decap_4 FILLER_23_730 ();
 sg13g2_fill_2 FILLER_23_739 ();
 sg13g2_fill_1 FILLER_23_746 ();
 sg13g2_fill_1 FILLER_23_771 ();
 sg13g2_decap_8 FILLER_23_782 ();
 sg13g2_fill_1 FILLER_23_789 ();
 sg13g2_fill_2 FILLER_23_806 ();
 sg13g2_fill_1 FILLER_23_813 ();
 sg13g2_decap_8 FILLER_23_818 ();
 sg13g2_fill_1 FILLER_23_825 ();
 sg13g2_fill_1 FILLER_23_831 ();
 sg13g2_fill_2 FILLER_23_837 ();
 sg13g2_fill_1 FILLER_23_839 ();
 sg13g2_fill_2 FILLER_23_876 ();
 sg13g2_decap_8 FILLER_24_0 ();
 sg13g2_decap_4 FILLER_24_7 ();
 sg13g2_decap_4 FILLER_24_16 ();
 sg13g2_fill_2 FILLER_24_53 ();
 sg13g2_fill_1 FILLER_24_60 ();
 sg13g2_fill_2 FILLER_24_76 ();
 sg13g2_decap_4 FILLER_24_82 ();
 sg13g2_fill_2 FILLER_24_93 ();
 sg13g2_fill_1 FILLER_24_129 ();
 sg13g2_fill_1 FILLER_24_138 ();
 sg13g2_fill_2 FILLER_24_148 ();
 sg13g2_fill_2 FILLER_24_167 ();
 sg13g2_fill_1 FILLER_24_180 ();
 sg13g2_fill_2 FILLER_24_186 ();
 sg13g2_fill_1 FILLER_24_188 ();
 sg13g2_fill_2 FILLER_24_198 ();
 sg13g2_fill_1 FILLER_24_208 ();
 sg13g2_fill_2 FILLER_24_252 ();
 sg13g2_fill_1 FILLER_24_254 ();
 sg13g2_fill_2 FILLER_24_259 ();
 sg13g2_fill_1 FILLER_24_261 ();
 sg13g2_decap_8 FILLER_24_267 ();
 sg13g2_decap_4 FILLER_24_274 ();
 sg13g2_decap_8 FILLER_24_283 ();
 sg13g2_decap_8 FILLER_24_290 ();
 sg13g2_decap_4 FILLER_24_297 ();
 sg13g2_fill_2 FILLER_24_340 ();
 sg13g2_fill_2 FILLER_24_347 ();
 sg13g2_fill_2 FILLER_24_353 ();
 sg13g2_decap_8 FILLER_24_389 ();
 sg13g2_decap_8 FILLER_24_396 ();
 sg13g2_decap_4 FILLER_24_403 ();
 sg13g2_decap_4 FILLER_24_429 ();
 sg13g2_fill_1 FILLER_24_438 ();
 sg13g2_fill_2 FILLER_24_452 ();
 sg13g2_fill_1 FILLER_24_454 ();
 sg13g2_decap_4 FILLER_24_460 ();
 sg13g2_fill_2 FILLER_24_464 ();
 sg13g2_decap_4 FILLER_24_488 ();
 sg13g2_fill_1 FILLER_24_492 ();
 sg13g2_fill_1 FILLER_24_515 ();
 sg13g2_decap_4 FILLER_24_532 ();
 sg13g2_fill_1 FILLER_24_536 ();
 sg13g2_fill_2 FILLER_24_541 ();
 sg13g2_fill_1 FILLER_24_543 ();
 sg13g2_fill_2 FILLER_24_559 ();
 sg13g2_fill_1 FILLER_24_561 ();
 sg13g2_fill_1 FILLER_24_567 ();
 sg13g2_decap_4 FILLER_24_574 ();
 sg13g2_fill_1 FILLER_24_578 ();
 sg13g2_fill_1 FILLER_24_583 ();
 sg13g2_decap_8 FILLER_24_592 ();
 sg13g2_fill_1 FILLER_24_599 ();
 sg13g2_fill_2 FILLER_24_621 ();
 sg13g2_decap_4 FILLER_24_628 ();
 sg13g2_fill_2 FILLER_24_632 ();
 sg13g2_fill_2 FILLER_24_646 ();
 sg13g2_fill_1 FILLER_24_648 ();
 sg13g2_fill_1 FILLER_24_672 ();
 sg13g2_fill_1 FILLER_24_686 ();
 sg13g2_fill_1 FILLER_24_711 ();
 sg13g2_fill_2 FILLER_24_725 ();
 sg13g2_fill_1 FILLER_24_732 ();
 sg13g2_decap_8 FILLER_24_750 ();
 sg13g2_fill_2 FILLER_24_757 ();
 sg13g2_fill_2 FILLER_24_772 ();
 sg13g2_fill_1 FILLER_24_779 ();
 sg13g2_decap_4 FILLER_24_786 ();
 sg13g2_fill_2 FILLER_24_790 ();
 sg13g2_fill_1 FILLER_24_798 ();
 sg13g2_fill_1 FILLER_24_803 ();
 sg13g2_decap_8 FILLER_24_818 ();
 sg13g2_decap_4 FILLER_24_825 ();
 sg13g2_fill_1 FILLER_24_829 ();
 sg13g2_decap_4 FILLER_24_846 ();
 sg13g2_fill_1 FILLER_24_850 ();
 sg13g2_decap_8 FILLER_24_870 ();
 sg13g2_fill_1 FILLER_24_877 ();
 sg13g2_decap_4 FILLER_25_0 ();
 sg13g2_fill_2 FILLER_25_4 ();
 sg13g2_fill_2 FILLER_25_18 ();
 sg13g2_decap_4 FILLER_25_24 ();
 sg13g2_fill_1 FILLER_25_28 ();
 sg13g2_fill_2 FILLER_25_49 ();
 sg13g2_decap_4 FILLER_25_63 ();
 sg13g2_fill_1 FILLER_25_67 ();
 sg13g2_fill_2 FILLER_25_98 ();
 sg13g2_decap_4 FILLER_25_114 ();
 sg13g2_fill_1 FILLER_25_118 ();
 sg13g2_fill_1 FILLER_25_145 ();
 sg13g2_fill_2 FILLER_25_169 ();
 sg13g2_fill_1 FILLER_25_171 ();
 sg13g2_fill_2 FILLER_25_183 ();
 sg13g2_fill_2 FILLER_25_200 ();
 sg13g2_fill_2 FILLER_25_207 ();
 sg13g2_fill_2 FILLER_25_233 ();
 sg13g2_fill_2 FILLER_25_240 ();
 sg13g2_decap_8 FILLER_25_285 ();
 sg13g2_decap_8 FILLER_25_292 ();
 sg13g2_decap_8 FILLER_25_299 ();
 sg13g2_fill_2 FILLER_25_323 ();
 sg13g2_fill_1 FILLER_25_325 ();
 sg13g2_fill_2 FILLER_25_340 ();
 sg13g2_decap_4 FILLER_25_395 ();
 sg13g2_fill_2 FILLER_25_399 ();
 sg13g2_fill_1 FILLER_25_414 ();
 sg13g2_fill_2 FILLER_25_420 ();
 sg13g2_decap_8 FILLER_25_432 ();
 sg13g2_fill_1 FILLER_25_439 ();
 sg13g2_fill_1 FILLER_25_460 ();
 sg13g2_fill_1 FILLER_25_473 ();
 sg13g2_fill_2 FILLER_25_493 ();
 sg13g2_fill_1 FILLER_25_495 ();
 sg13g2_fill_2 FILLER_25_512 ();
 sg13g2_fill_1 FILLER_25_514 ();
 sg13g2_fill_1 FILLER_25_523 ();
 sg13g2_fill_2 FILLER_25_559 ();
 sg13g2_fill_2 FILLER_25_565 ();
 sg13g2_decap_8 FILLER_25_571 ();
 sg13g2_fill_2 FILLER_25_582 ();
 sg13g2_fill_2 FILLER_25_592 ();
 sg13g2_fill_1 FILLER_25_594 ();
 sg13g2_fill_2 FILLER_25_600 ();
 sg13g2_fill_1 FILLER_25_602 ();
 sg13g2_fill_2 FILLER_25_607 ();
 sg13g2_fill_1 FILLER_25_635 ();
 sg13g2_fill_1 FILLER_25_641 ();
 sg13g2_fill_1 FILLER_25_653 ();
 sg13g2_decap_4 FILLER_25_659 ();
 sg13g2_fill_2 FILLER_25_663 ();
 sg13g2_decap_8 FILLER_25_675 ();
 sg13g2_decap_8 FILLER_25_682 ();
 sg13g2_fill_1 FILLER_25_689 ();
 sg13g2_fill_2 FILLER_25_694 ();
 sg13g2_fill_1 FILLER_25_696 ();
 sg13g2_fill_2 FILLER_25_702 ();
 sg13g2_decap_4 FILLER_25_708 ();
 sg13g2_fill_1 FILLER_25_722 ();
 sg13g2_fill_1 FILLER_25_737 ();
 sg13g2_fill_2 FILLER_25_750 ();
 sg13g2_fill_2 FILLER_25_757 ();
 sg13g2_fill_1 FILLER_25_779 ();
 sg13g2_fill_1 FILLER_25_805 ();
 sg13g2_fill_2 FILLER_25_825 ();
 sg13g2_decap_4 FILLER_25_847 ();
 sg13g2_decap_4 FILLER_25_872 ();
 sg13g2_fill_2 FILLER_25_876 ();
 sg13g2_fill_1 FILLER_26_0 ();
 sg13g2_fill_1 FILLER_26_9 ();
 sg13g2_fill_1 FILLER_26_19 ();
 sg13g2_decap_8 FILLER_26_24 ();
 sg13g2_decap_4 FILLER_26_31 ();
 sg13g2_fill_1 FILLER_26_35 ();
 sg13g2_decap_4 FILLER_26_51 ();
 sg13g2_fill_1 FILLER_26_59 ();
 sg13g2_fill_1 FILLER_26_64 ();
 sg13g2_fill_1 FILLER_26_69 ();
 sg13g2_fill_1 FILLER_26_74 ();
 sg13g2_fill_2 FILLER_26_91 ();
 sg13g2_fill_1 FILLER_26_93 ();
 sg13g2_fill_2 FILLER_26_98 ();
 sg13g2_fill_1 FILLER_26_100 ();
 sg13g2_fill_2 FILLER_26_109 ();
 sg13g2_decap_8 FILLER_26_119 ();
 sg13g2_decap_4 FILLER_26_126 ();
 sg13g2_fill_1 FILLER_26_135 ();
 sg13g2_fill_1 FILLER_26_147 ();
 sg13g2_decap_4 FILLER_26_160 ();
 sg13g2_fill_2 FILLER_26_171 ();
 sg13g2_fill_1 FILLER_26_173 ();
 sg13g2_decap_4 FILLER_26_189 ();
 sg13g2_decap_4 FILLER_26_228 ();
 sg13g2_fill_1 FILLER_26_232 ();
 sg13g2_fill_1 FILLER_26_241 ();
 sg13g2_fill_2 FILLER_26_267 ();
 sg13g2_fill_2 FILLER_26_277 ();
 sg13g2_decap_8 FILLER_26_291 ();
 sg13g2_fill_1 FILLER_26_303 ();
 sg13g2_fill_2 FILLER_26_309 ();
 sg13g2_fill_2 FILLER_26_318 ();
 sg13g2_fill_1 FILLER_26_320 ();
 sg13g2_fill_1 FILLER_26_359 ();
 sg13g2_fill_2 FILLER_26_378 ();
 sg13g2_decap_8 FILLER_26_393 ();
 sg13g2_fill_1 FILLER_26_400 ();
 sg13g2_decap_4 FILLER_26_422 ();
 sg13g2_fill_2 FILLER_26_426 ();
 sg13g2_fill_1 FILLER_26_447 ();
 sg13g2_fill_1 FILLER_26_459 ();
 sg13g2_fill_2 FILLER_26_468 ();
 sg13g2_decap_8 FILLER_26_474 ();
 sg13g2_fill_1 FILLER_26_481 ();
 sg13g2_decap_8 FILLER_26_509 ();
 sg13g2_fill_2 FILLER_26_540 ();
 sg13g2_fill_1 FILLER_26_542 ();
 sg13g2_fill_2 FILLER_26_547 ();
 sg13g2_fill_2 FILLER_26_554 ();
 sg13g2_decap_4 FILLER_26_592 ();
 sg13g2_fill_1 FILLER_26_596 ();
 sg13g2_fill_1 FILLER_26_623 ();
 sg13g2_decap_8 FILLER_26_631 ();
 sg13g2_fill_1 FILLER_26_643 ();
 sg13g2_decap_8 FILLER_26_662 ();
 sg13g2_fill_1 FILLER_26_669 ();
 sg13g2_decap_8 FILLER_26_675 ();
 sg13g2_decap_4 FILLER_26_682 ();
 sg13g2_fill_2 FILLER_26_693 ();
 sg13g2_decap_8 FILLER_26_725 ();
 sg13g2_decap_8 FILLER_26_737 ();
 sg13g2_decap_8 FILLER_26_744 ();
 sg13g2_decap_8 FILLER_26_751 ();
 sg13g2_decap_8 FILLER_26_758 ();
 sg13g2_fill_1 FILLER_26_773 ();
 sg13g2_fill_1 FILLER_26_778 ();
 sg13g2_fill_1 FILLER_26_783 ();
 sg13g2_fill_2 FILLER_26_788 ();
 sg13g2_decap_8 FILLER_26_802 ();
 sg13g2_decap_8 FILLER_26_809 ();
 sg13g2_decap_8 FILLER_26_816 ();
 sg13g2_decap_4 FILLER_26_823 ();
 sg13g2_fill_1 FILLER_26_827 ();
 sg13g2_decap_4 FILLER_26_833 ();
 sg13g2_decap_4 FILLER_26_841 ();
 sg13g2_fill_1 FILLER_26_866 ();
 sg13g2_decap_8 FILLER_26_871 ();
 sg13g2_decap_4 FILLER_27_0 ();
 sg13g2_fill_2 FILLER_27_12 ();
 sg13g2_fill_2 FILLER_27_24 ();
 sg13g2_fill_1 FILLER_27_26 ();
 sg13g2_fill_1 FILLER_27_31 ();
 sg13g2_fill_2 FILLER_27_40 ();
 sg13g2_fill_1 FILLER_27_42 ();
 sg13g2_decap_4 FILLER_27_48 ();
 sg13g2_fill_2 FILLER_27_52 ();
 sg13g2_fill_2 FILLER_27_63 ();
 sg13g2_fill_1 FILLER_27_65 ();
 sg13g2_fill_2 FILLER_27_71 ();
 sg13g2_fill_2 FILLER_27_77 ();
 sg13g2_fill_2 FILLER_27_84 ();
 sg13g2_fill_2 FILLER_27_95 ();
 sg13g2_fill_1 FILLER_27_97 ();
 sg13g2_fill_2 FILLER_27_106 ();
 sg13g2_fill_1 FILLER_27_108 ();
 sg13g2_fill_2 FILLER_27_122 ();
 sg13g2_fill_1 FILLER_27_130 ();
 sg13g2_fill_2 FILLER_27_135 ();
 sg13g2_fill_2 FILLER_27_167 ();
 sg13g2_fill_2 FILLER_27_179 ();
 sg13g2_fill_1 FILLER_27_181 ();
 sg13g2_decap_4 FILLER_27_186 ();
 sg13g2_fill_1 FILLER_27_190 ();
 sg13g2_fill_2 FILLER_27_196 ();
 sg13g2_fill_1 FILLER_27_198 ();
 sg13g2_fill_2 FILLER_27_209 ();
 sg13g2_fill_1 FILLER_27_211 ();
 sg13g2_decap_8 FILLER_27_234 ();
 sg13g2_fill_2 FILLER_27_241 ();
 sg13g2_fill_1 FILLER_27_248 ();
 sg13g2_decap_8 FILLER_27_267 ();
 sg13g2_fill_2 FILLER_27_274 ();
 sg13g2_fill_2 FILLER_27_294 ();
 sg13g2_fill_2 FILLER_27_300 ();
 sg13g2_fill_1 FILLER_27_302 ();
 sg13g2_fill_1 FILLER_27_308 ();
 sg13g2_fill_2 FILLER_27_314 ();
 sg13g2_fill_1 FILLER_27_316 ();
 sg13g2_fill_1 FILLER_27_325 ();
 sg13g2_fill_1 FILLER_27_355 ();
 sg13g2_decap_8 FILLER_27_382 ();
 sg13g2_fill_2 FILLER_27_389 ();
 sg13g2_fill_1 FILLER_27_391 ();
 sg13g2_decap_8 FILLER_27_410 ();
 sg13g2_decap_8 FILLER_27_417 ();
 sg13g2_fill_2 FILLER_27_424 ();
 sg13g2_fill_1 FILLER_27_432 ();
 sg13g2_fill_2 FILLER_27_469 ();
 sg13g2_decap_8 FILLER_27_474 ();
 sg13g2_fill_2 FILLER_27_481 ();
 sg13g2_fill_2 FILLER_27_488 ();
 sg13g2_fill_1 FILLER_27_490 ();
 sg13g2_fill_2 FILLER_27_501 ();
 sg13g2_decap_8 FILLER_27_513 ();
 sg13g2_decap_8 FILLER_27_520 ();
 sg13g2_decap_8 FILLER_27_527 ();
 sg13g2_fill_1 FILLER_27_534 ();
 sg13g2_fill_2 FILLER_27_543 ();
 sg13g2_fill_1 FILLER_27_545 ();
 sg13g2_decap_4 FILLER_27_550 ();
 sg13g2_fill_1 FILLER_27_554 ();
 sg13g2_decap_8 FILLER_27_581 ();
 sg13g2_fill_1 FILLER_27_592 ();
 sg13g2_decap_8 FILLER_27_609 ();
 sg13g2_decap_8 FILLER_27_625 ();
 sg13g2_fill_2 FILLER_27_659 ();
 sg13g2_fill_2 FILLER_27_681 ();
 sg13g2_fill_1 FILLER_27_687 ();
 sg13g2_decap_4 FILLER_27_691 ();
 sg13g2_fill_2 FILLER_27_705 ();
 sg13g2_decap_8 FILLER_27_712 ();
 sg13g2_decap_8 FILLER_27_719 ();
 sg13g2_fill_2 FILLER_27_726 ();
 sg13g2_fill_1 FILLER_27_733 ();
 sg13g2_fill_1 FILLER_27_742 ();
 sg13g2_fill_2 FILLER_27_748 ();
 sg13g2_decap_8 FILLER_27_753 ();
 sg13g2_decap_8 FILLER_27_760 ();
 sg13g2_decap_8 FILLER_27_774 ();
 sg13g2_fill_2 FILLER_27_781 ();
 sg13g2_fill_1 FILLER_27_783 ();
 sg13g2_fill_1 FILLER_27_834 ();
 sg13g2_decap_4 FILLER_27_839 ();
 sg13g2_decap_8 FILLER_27_847 ();
 sg13g2_fill_2 FILLER_27_854 ();
 sg13g2_fill_1 FILLER_27_856 ();
 sg13g2_fill_1 FILLER_27_862 ();
 sg13g2_decap_8 FILLER_27_871 ();
 sg13g2_decap_4 FILLER_28_0 ();
 sg13g2_fill_2 FILLER_28_4 ();
 sg13g2_fill_1 FILLER_28_15 ();
 sg13g2_fill_2 FILLER_28_32 ();
 sg13g2_fill_2 FILLER_28_39 ();
 sg13g2_fill_1 FILLER_28_41 ();
 sg13g2_fill_2 FILLER_28_50 ();
 sg13g2_fill_1 FILLER_28_75 ();
 sg13g2_fill_2 FILLER_28_80 ();
 sg13g2_fill_1 FILLER_28_90 ();
 sg13g2_fill_1 FILLER_28_95 ();
 sg13g2_fill_1 FILLER_28_106 ();
 sg13g2_fill_1 FILLER_28_115 ();
 sg13g2_decap_8 FILLER_28_121 ();
 sg13g2_decap_8 FILLER_28_128 ();
 sg13g2_fill_1 FILLER_28_135 ();
 sg13g2_fill_1 FILLER_28_149 ();
 sg13g2_fill_1 FILLER_28_155 ();
 sg13g2_fill_1 FILLER_28_161 ();
 sg13g2_fill_2 FILLER_28_171 ();
 sg13g2_decap_4 FILLER_28_187 ();
 sg13g2_fill_1 FILLER_28_191 ();
 sg13g2_fill_1 FILLER_28_232 ();
 sg13g2_fill_1 FILLER_28_245 ();
 sg13g2_fill_1 FILLER_28_250 ();
 sg13g2_decap_4 FILLER_28_255 ();
 sg13g2_fill_2 FILLER_28_263 ();
 sg13g2_fill_1 FILLER_28_270 ();
 sg13g2_fill_2 FILLER_28_295 ();
 sg13g2_fill_2 FILLER_28_301 ();
 sg13g2_fill_1 FILLER_28_303 ();
 sg13g2_decap_4 FILLER_28_318 ();
 sg13g2_fill_1 FILLER_28_322 ();
 sg13g2_decap_4 FILLER_28_327 ();
 sg13g2_fill_2 FILLER_28_362 ();
 sg13g2_fill_1 FILLER_28_368 ();
 sg13g2_fill_1 FILLER_28_404 ();
 sg13g2_decap_4 FILLER_28_409 ();
 sg13g2_fill_1 FILLER_28_413 ();
 sg13g2_decap_4 FILLER_28_426 ();
 sg13g2_fill_2 FILLER_28_442 ();
 sg13g2_fill_1 FILLER_28_444 ();
 sg13g2_decap_8 FILLER_28_487 ();
 sg13g2_decap_4 FILLER_28_494 ();
 sg13g2_decap_4 FILLER_28_508 ();
 sg13g2_fill_1 FILLER_28_512 ();
 sg13g2_decap_8 FILLER_28_577 ();
 sg13g2_fill_2 FILLER_28_584 ();
 sg13g2_fill_1 FILLER_28_586 ();
 sg13g2_fill_2 FILLER_28_590 ();
 sg13g2_fill_1 FILLER_28_592 ();
 sg13g2_fill_2 FILLER_28_597 ();
 sg13g2_decap_8 FILLER_28_609 ();
 sg13g2_fill_2 FILLER_28_616 ();
 sg13g2_fill_1 FILLER_28_640 ();
 sg13g2_decap_8 FILLER_28_648 ();
 sg13g2_fill_1 FILLER_28_655 ();
 sg13g2_fill_1 FILLER_28_669 ();
 sg13g2_fill_2 FILLER_28_676 ();
 sg13g2_fill_1 FILLER_28_684 ();
 sg13g2_decap_4 FILLER_28_694 ();
 sg13g2_fill_1 FILLER_28_698 ();
 sg13g2_decap_4 FILLER_28_717 ();
 sg13g2_decap_4 FILLER_28_728 ();
 sg13g2_fill_1 FILLER_28_732 ();
 sg13g2_decap_4 FILLER_28_742 ();
 sg13g2_fill_1 FILLER_28_762 ();
 sg13g2_fill_1 FILLER_28_768 ();
 sg13g2_decap_4 FILLER_28_774 ();
 sg13g2_fill_1 FILLER_28_778 ();
 sg13g2_decap_4 FILLER_28_783 ();
 sg13g2_fill_2 FILLER_28_787 ();
 sg13g2_decap_4 FILLER_28_794 ();
 sg13g2_decap_4 FILLER_28_802 ();
 sg13g2_fill_2 FILLER_28_811 ();
 sg13g2_fill_1 FILLER_28_813 ();
 sg13g2_decap_4 FILLER_28_819 ();
 sg13g2_decap_8 FILLER_28_827 ();
 sg13g2_decap_4 FILLER_28_834 ();
 sg13g2_fill_2 FILLER_28_868 ();
 sg13g2_decap_4 FILLER_28_873 ();
 sg13g2_fill_1 FILLER_28_877 ();
 sg13g2_decap_8 FILLER_29_0 ();
 sg13g2_fill_2 FILLER_29_7 ();
 sg13g2_fill_1 FILLER_29_9 ();
 sg13g2_fill_1 FILLER_29_14 ();
 sg13g2_decap_8 FILLER_29_28 ();
 sg13g2_fill_2 FILLER_29_35 ();
 sg13g2_fill_1 FILLER_29_37 ();
 sg13g2_decap_4 FILLER_29_42 ();
 sg13g2_fill_1 FILLER_29_63 ();
 sg13g2_fill_2 FILLER_29_80 ();
 sg13g2_decap_4 FILLER_29_95 ();
 sg13g2_fill_2 FILLER_29_103 ();
 sg13g2_fill_2 FILLER_29_110 ();
 sg13g2_fill_1 FILLER_29_112 ();
 sg13g2_decap_8 FILLER_29_153 ();
 sg13g2_decap_4 FILLER_29_160 ();
 sg13g2_fill_2 FILLER_29_172 ();
 sg13g2_fill_2 FILLER_29_179 ();
 sg13g2_decap_4 FILLER_29_198 ();
 sg13g2_fill_1 FILLER_29_202 ();
 sg13g2_fill_1 FILLER_29_207 ();
 sg13g2_decap_8 FILLER_29_228 ();
 sg13g2_fill_2 FILLER_29_235 ();
 sg13g2_fill_1 FILLER_29_237 ();
 sg13g2_decap_4 FILLER_29_250 ();
 sg13g2_fill_2 FILLER_29_265 ();
 sg13g2_decap_8 FILLER_29_298 ();
 sg13g2_decap_4 FILLER_29_305 ();
 sg13g2_fill_1 FILLER_29_309 ();
 sg13g2_decap_4 FILLER_29_325 ();
 sg13g2_fill_2 FILLER_29_329 ();
 sg13g2_decap_4 FILLER_29_335 ();
 sg13g2_decap_4 FILLER_29_380 ();
 sg13g2_fill_1 FILLER_29_384 ();
 sg13g2_decap_4 FILLER_29_393 ();
 sg13g2_decap_8 FILLER_29_413 ();
 sg13g2_decap_8 FILLER_29_428 ();
 sg13g2_decap_8 FILLER_29_435 ();
 sg13g2_decap_8 FILLER_29_442 ();
 sg13g2_fill_2 FILLER_29_461 ();
 sg13g2_fill_1 FILLER_29_463 ();
 sg13g2_decap_8 FILLER_29_491 ();
 sg13g2_fill_2 FILLER_29_498 ();
 sg13g2_fill_1 FILLER_29_500 ();
 sg13g2_fill_1 FILLER_29_511 ();
 sg13g2_fill_2 FILLER_29_517 ();
 sg13g2_fill_1 FILLER_29_519 ();
 sg13g2_fill_1 FILLER_29_528 ();
 sg13g2_fill_2 FILLER_29_533 ();
 sg13g2_fill_2 FILLER_29_540 ();
 sg13g2_fill_1 FILLER_29_542 ();
 sg13g2_decap_8 FILLER_29_546 ();
 sg13g2_fill_2 FILLER_29_553 ();
 sg13g2_fill_1 FILLER_29_555 ();
 sg13g2_fill_2 FILLER_29_560 ();
 sg13g2_fill_1 FILLER_29_562 ();
 sg13g2_decap_8 FILLER_29_567 ();
 sg13g2_decap_4 FILLER_29_574 ();
 sg13g2_fill_2 FILLER_29_578 ();
 sg13g2_fill_1 FILLER_29_616 ();
 sg13g2_fill_2 FILLER_29_647 ();
 sg13g2_decap_8 FILLER_29_661 ();
 sg13g2_decap_4 FILLER_29_668 ();
 sg13g2_decap_4 FILLER_29_676 ();
 sg13g2_fill_2 FILLER_29_689 ();
 sg13g2_fill_1 FILLER_29_691 ();
 sg13g2_fill_2 FILLER_29_697 ();
 sg13g2_fill_1 FILLER_29_699 ();
 sg13g2_fill_2 FILLER_29_706 ();
 sg13g2_fill_2 FILLER_29_717 ();
 sg13g2_fill_1 FILLER_29_719 ();
 sg13g2_decap_8 FILLER_29_728 ();
 sg13g2_fill_1 FILLER_29_739 ();
 sg13g2_fill_2 FILLER_29_752 ();
 sg13g2_fill_1 FILLER_29_754 ();
 sg13g2_decap_8 FILLER_29_760 ();
 sg13g2_decap_8 FILLER_29_767 ();
 sg13g2_fill_2 FILLER_29_774 ();
 sg13g2_fill_1 FILLER_29_776 ();
 sg13g2_fill_2 FILLER_29_810 ();
 sg13g2_fill_2 FILLER_29_825 ();
 sg13g2_fill_2 FILLER_29_832 ();
 sg13g2_fill_1 FILLER_29_834 ();
 sg13g2_decap_8 FILLER_29_839 ();
 sg13g2_decap_4 FILLER_29_846 ();
 sg13g2_fill_2 FILLER_29_850 ();
 sg13g2_fill_1 FILLER_29_869 ();
 sg13g2_fill_2 FILLER_29_875 ();
 sg13g2_fill_1 FILLER_29_877 ();
 sg13g2_fill_2 FILLER_30_0 ();
 sg13g2_fill_1 FILLER_30_2 ();
 sg13g2_decap_4 FILLER_30_22 ();
 sg13g2_fill_1 FILLER_30_26 ();
 sg13g2_decap_8 FILLER_30_32 ();
 sg13g2_decap_4 FILLER_30_39 ();
 sg13g2_fill_1 FILLER_30_43 ();
 sg13g2_fill_2 FILLER_30_57 ();
 sg13g2_fill_1 FILLER_30_59 ();
 sg13g2_decap_8 FILLER_30_68 ();
 sg13g2_decap_8 FILLER_30_75 ();
 sg13g2_fill_1 FILLER_30_82 ();
 sg13g2_fill_1 FILLER_30_87 ();
 sg13g2_fill_1 FILLER_30_96 ();
 sg13g2_fill_1 FILLER_30_100 ();
 sg13g2_fill_1 FILLER_30_111 ();
 sg13g2_decap_4 FILLER_30_117 ();
 sg13g2_decap_8 FILLER_30_129 ();
 sg13g2_decap_8 FILLER_30_136 ();
 sg13g2_decap_4 FILLER_30_143 ();
 sg13g2_fill_2 FILLER_30_147 ();
 sg13g2_fill_2 FILLER_30_153 ();
 sg13g2_fill_2 FILLER_30_175 ();
 sg13g2_fill_1 FILLER_30_177 ();
 sg13g2_fill_1 FILLER_30_183 ();
 sg13g2_fill_2 FILLER_30_189 ();
 sg13g2_decap_8 FILLER_30_199 ();
 sg13g2_decap_8 FILLER_30_206 ();
 sg13g2_decap_4 FILLER_30_213 ();
 sg13g2_decap_8 FILLER_30_221 ();
 sg13g2_decap_8 FILLER_30_228 ();
 sg13g2_decap_4 FILLER_30_247 ();
 sg13g2_fill_2 FILLER_30_251 ();
 sg13g2_decap_4 FILLER_30_268 ();
 sg13g2_decap_8 FILLER_30_280 ();
 sg13g2_fill_1 FILLER_30_287 ();
 sg13g2_decap_4 FILLER_30_292 ();
 sg13g2_fill_2 FILLER_30_304 ();
 sg13g2_fill_2 FILLER_30_314 ();
 sg13g2_fill_2 FILLER_30_332 ();
 sg13g2_decap_4 FILLER_30_338 ();
 sg13g2_decap_4 FILLER_30_350 ();
 sg13g2_fill_1 FILLER_30_354 ();
 sg13g2_decap_4 FILLER_30_370 ();
 sg13g2_decap_8 FILLER_30_382 ();
 sg13g2_decap_8 FILLER_30_389 ();
 sg13g2_fill_2 FILLER_30_396 ();
 sg13g2_fill_2 FILLER_30_424 ();
 sg13g2_fill_1 FILLER_30_444 ();
 sg13g2_fill_2 FILLER_30_455 ();
 sg13g2_fill_2 FILLER_30_461 ();
 sg13g2_fill_2 FILLER_30_467 ();
 sg13g2_fill_2 FILLER_30_478 ();
 sg13g2_decap_4 FILLER_30_488 ();
 sg13g2_fill_1 FILLER_30_492 ();
 sg13g2_decap_4 FILLER_30_497 ();
 sg13g2_fill_2 FILLER_30_501 ();
 sg13g2_decap_8 FILLER_30_548 ();
 sg13g2_fill_1 FILLER_30_555 ();
 sg13g2_fill_2 FILLER_30_560 ();
 sg13g2_fill_2 FILLER_30_571 ();
 sg13g2_fill_1 FILLER_30_573 ();
 sg13g2_decap_8 FILLER_30_586 ();
 sg13g2_decap_8 FILLER_30_593 ();
 sg13g2_fill_2 FILLER_30_600 ();
 sg13g2_fill_1 FILLER_30_602 ();
 sg13g2_decap_8 FILLER_30_608 ();
 sg13g2_fill_2 FILLER_30_615 ();
 sg13g2_fill_1 FILLER_30_628 ();
 sg13g2_fill_1 FILLER_30_636 ();
 sg13g2_fill_1 FILLER_30_643 ();
 sg13g2_fill_1 FILLER_30_649 ();
 sg13g2_fill_1 FILLER_30_655 ();
 sg13g2_decap_8 FILLER_30_668 ();
 sg13g2_fill_2 FILLER_30_675 ();
 sg13g2_decap_4 FILLER_30_704 ();
 sg13g2_fill_1 FILLER_30_708 ();
 sg13g2_fill_2 FILLER_30_714 ();
 sg13g2_fill_1 FILLER_30_716 ();
 sg13g2_fill_2 FILLER_30_722 ();
 sg13g2_fill_1 FILLER_30_724 ();
 sg13g2_fill_2 FILLER_30_750 ();
 sg13g2_decap_8 FILLER_30_762 ();
 sg13g2_decap_4 FILLER_30_769 ();
 sg13g2_fill_2 FILLER_30_773 ();
 sg13g2_fill_1 FILLER_30_780 ();
 sg13g2_fill_2 FILLER_30_785 ();
 sg13g2_decap_8 FILLER_30_791 ();
 sg13g2_decap_8 FILLER_30_798 ();
 sg13g2_decap_8 FILLER_30_805 ();
 sg13g2_decap_4 FILLER_30_812 ();
 sg13g2_fill_2 FILLER_30_816 ();
 sg13g2_fill_1 FILLER_30_847 ();
 sg13g2_fill_2 FILLER_30_876 ();
 sg13g2_decap_4 FILLER_31_0 ();
 sg13g2_fill_2 FILLER_31_4 ();
 sg13g2_fill_1 FILLER_31_10 ();
 sg13g2_fill_1 FILLER_31_16 ();
 sg13g2_fill_1 FILLER_31_39 ();
 sg13g2_fill_1 FILLER_31_45 ();
 sg13g2_fill_1 FILLER_31_50 ();
 sg13g2_fill_1 FILLER_31_55 ();
 sg13g2_decap_8 FILLER_31_60 ();
 sg13g2_decap_4 FILLER_31_78 ();
 sg13g2_decap_4 FILLER_31_90 ();
 sg13g2_fill_2 FILLER_31_119 ();
 sg13g2_decap_8 FILLER_31_126 ();
 sg13g2_fill_1 FILLER_31_141 ();
 sg13g2_fill_1 FILLER_31_147 ();
 sg13g2_fill_1 FILLER_31_168 ();
 sg13g2_fill_1 FILLER_31_177 ();
 sg13g2_fill_1 FILLER_31_187 ();
 sg13g2_decap_4 FILLER_31_192 ();
 sg13g2_fill_2 FILLER_31_204 ();
 sg13g2_decap_8 FILLER_31_210 ();
 sg13g2_decap_8 FILLER_31_217 ();
 sg13g2_fill_1 FILLER_31_224 ();
 sg13g2_fill_2 FILLER_31_241 ();
 sg13g2_fill_1 FILLER_31_243 ();
 sg13g2_decap_8 FILLER_31_262 ();
 sg13g2_fill_2 FILLER_31_281 ();
 sg13g2_fill_1 FILLER_31_283 ();
 sg13g2_decap_4 FILLER_31_292 ();
 sg13g2_fill_2 FILLER_31_296 ();
 sg13g2_decap_8 FILLER_31_303 ();
 sg13g2_decap_4 FILLER_31_310 ();
 sg13g2_fill_2 FILLER_31_314 ();
 sg13g2_fill_2 FILLER_31_331 ();
 sg13g2_fill_1 FILLER_31_340 ();
 sg13g2_fill_1 FILLER_31_344 ();
 sg13g2_fill_2 FILLER_31_350 ();
 sg13g2_fill_1 FILLER_31_352 ();
 sg13g2_decap_8 FILLER_31_361 ();
 sg13g2_decap_4 FILLER_31_368 ();
 sg13g2_decap_8 FILLER_31_376 ();
 sg13g2_fill_2 FILLER_31_383 ();
 sg13g2_fill_1 FILLER_31_385 ();
 sg13g2_fill_1 FILLER_31_403 ();
 sg13g2_fill_2 FILLER_31_408 ();
 sg13g2_fill_1 FILLER_31_410 ();
 sg13g2_decap_8 FILLER_31_415 ();
 sg13g2_fill_2 FILLER_31_422 ();
 sg13g2_fill_1 FILLER_31_424 ();
 sg13g2_fill_1 FILLER_31_433 ();
 sg13g2_fill_2 FILLER_31_454 ();
 sg13g2_fill_2 FILLER_31_461 ();
 sg13g2_fill_1 FILLER_31_463 ();
 sg13g2_fill_2 FILLER_31_468 ();
 sg13g2_fill_1 FILLER_31_470 ();
 sg13g2_fill_2 FILLER_31_478 ();
 sg13g2_fill_1 FILLER_31_480 ();
 sg13g2_decap_8 FILLER_31_489 ();
 sg13g2_decap_8 FILLER_31_496 ();
 sg13g2_fill_1 FILLER_31_503 ();
 sg13g2_fill_2 FILLER_31_508 ();
 sg13g2_fill_1 FILLER_31_510 ();
 sg13g2_fill_2 FILLER_31_531 ();
 sg13g2_fill_1 FILLER_31_533 ();
 sg13g2_fill_2 FILLER_31_555 ();
 sg13g2_decap_8 FILLER_31_575 ();
 sg13g2_decap_8 FILLER_31_582 ();
 sg13g2_decap_8 FILLER_31_589 ();
 sg13g2_decap_4 FILLER_31_596 ();
 sg13g2_fill_1 FILLER_31_600 ();
 sg13g2_decap_4 FILLER_31_605 ();
 sg13g2_fill_2 FILLER_31_638 ();
 sg13g2_fill_1 FILLER_31_640 ();
 sg13g2_decap_8 FILLER_31_659 ();
 sg13g2_decap_4 FILLER_31_671 ();
 sg13g2_fill_1 FILLER_31_675 ();
 sg13g2_decap_4 FILLER_31_719 ();
 sg13g2_fill_2 FILLER_31_723 ();
 sg13g2_fill_2 FILLER_31_747 ();
 sg13g2_fill_1 FILLER_31_749 ();
 sg13g2_fill_1 FILLER_31_755 ();
 sg13g2_fill_2 FILLER_31_768 ();
 sg13g2_decap_4 FILLER_31_774 ();
 sg13g2_fill_1 FILLER_31_778 ();
 sg13g2_decap_4 FILLER_31_799 ();
 sg13g2_decap_8 FILLER_31_816 ();
 sg13g2_fill_2 FILLER_31_823 ();
 sg13g2_fill_1 FILLER_31_825 ();
 sg13g2_fill_1 FILLER_31_839 ();
 sg13g2_decap_8 FILLER_31_869 ();
 sg13g2_fill_2 FILLER_31_876 ();
 sg13g2_decap_4 FILLER_32_0 ();
 sg13g2_fill_2 FILLER_32_4 ();
 sg13g2_fill_1 FILLER_32_35 ();
 sg13g2_fill_1 FILLER_32_59 ();
 sg13g2_fill_2 FILLER_32_68 ();
 sg13g2_fill_1 FILLER_32_70 ();
 sg13g2_fill_2 FILLER_32_79 ();
 sg13g2_fill_1 FILLER_32_81 ();
 sg13g2_fill_1 FILLER_32_91 ();
 sg13g2_decap_8 FILLER_32_100 ();
 sg13g2_fill_2 FILLER_32_107 ();
 sg13g2_fill_1 FILLER_32_109 ();
 sg13g2_fill_1 FILLER_32_118 ();
 sg13g2_fill_2 FILLER_32_127 ();
 sg13g2_fill_2 FILLER_32_134 ();
 sg13g2_fill_2 FILLER_32_140 ();
 sg13g2_fill_1 FILLER_32_142 ();
 sg13g2_fill_2 FILLER_32_151 ();
 sg13g2_decap_8 FILLER_32_157 ();
 sg13g2_decap_4 FILLER_32_164 ();
 sg13g2_fill_2 FILLER_32_168 ();
 sg13g2_fill_2 FILLER_32_195 ();
 sg13g2_decap_4 FILLER_32_222 ();
 sg13g2_fill_1 FILLER_32_226 ();
 sg13g2_decap_4 FILLER_32_243 ();
 sg13g2_fill_1 FILLER_32_247 ();
 sg13g2_fill_2 FILLER_32_264 ();
 sg13g2_fill_2 FILLER_32_270 ();
 sg13g2_fill_1 FILLER_32_276 ();
 sg13g2_decap_8 FILLER_32_293 ();
 sg13g2_fill_1 FILLER_32_308 ();
 sg13g2_decap_8 FILLER_32_317 ();
 sg13g2_decap_8 FILLER_32_347 ();
 sg13g2_fill_1 FILLER_32_354 ();
 sg13g2_fill_1 FILLER_32_359 ();
 sg13g2_fill_1 FILLER_32_391 ();
 sg13g2_fill_2 FILLER_32_409 ();
 sg13g2_fill_1 FILLER_32_432 ();
 sg13g2_fill_1 FILLER_32_438 ();
 sg13g2_decap_4 FILLER_32_443 ();
 sg13g2_fill_1 FILLER_32_455 ();
 sg13g2_fill_1 FILLER_32_461 ();
 sg13g2_decap_4 FILLER_32_474 ();
 sg13g2_decap_4 FILLER_32_496 ();
 sg13g2_decap_4 FILLER_32_504 ();
 sg13g2_fill_1 FILLER_32_508 ();
 sg13g2_fill_2 FILLER_32_522 ();
 sg13g2_decap_8 FILLER_32_536 ();
 sg13g2_fill_2 FILLER_32_543 ();
 sg13g2_fill_1 FILLER_32_545 ();
 sg13g2_fill_2 FILLER_32_555 ();
 sg13g2_decap_4 FILLER_32_583 ();
 sg13g2_fill_2 FILLER_32_587 ();
 sg13g2_fill_1 FILLER_32_605 ();
 sg13g2_fill_1 FILLER_32_610 ();
 sg13g2_fill_1 FILLER_32_614 ();
 sg13g2_fill_1 FILLER_32_619 ();
 sg13g2_fill_2 FILLER_32_624 ();
 sg13g2_fill_1 FILLER_32_641 ();
 sg13g2_decap_8 FILLER_32_646 ();
 sg13g2_decap_4 FILLER_32_653 ();
 sg13g2_fill_1 FILLER_32_657 ();
 sg13g2_fill_2 FILLER_32_666 ();
 sg13g2_fill_1 FILLER_32_668 ();
 sg13g2_fill_1 FILLER_32_688 ();
 sg13g2_fill_2 FILLER_32_705 ();
 sg13g2_decap_4 FILLER_32_715 ();
 sg13g2_decap_8 FILLER_32_740 ();
 sg13g2_fill_1 FILLER_32_747 ();
 sg13g2_decap_8 FILLER_32_784 ();
 sg13g2_decap_8 FILLER_32_799 ();
 sg13g2_decap_4 FILLER_32_806 ();
 sg13g2_fill_2 FILLER_32_810 ();
 sg13g2_fill_2 FILLER_32_836 ();
 sg13g2_fill_1 FILLER_32_838 ();
 sg13g2_decap_4 FILLER_32_844 ();
 sg13g2_decap_8 FILLER_32_869 ();
 sg13g2_fill_2 FILLER_32_876 ();
 sg13g2_decap_8 FILLER_33_0 ();
 sg13g2_decap_4 FILLER_33_7 ();
 sg13g2_fill_2 FILLER_33_11 ();
 sg13g2_decap_8 FILLER_33_37 ();
 sg13g2_decap_8 FILLER_33_44 ();
 sg13g2_fill_2 FILLER_33_51 ();
 sg13g2_decap_4 FILLER_33_80 ();
 sg13g2_fill_1 FILLER_33_88 ();
 sg13g2_fill_2 FILLER_33_105 ();
 sg13g2_fill_1 FILLER_33_107 ();
 sg13g2_fill_1 FILLER_33_137 ();
 sg13g2_decap_4 FILLER_33_148 ();
 sg13g2_decap_8 FILLER_33_170 ();
 sg13g2_decap_4 FILLER_33_204 ();
 sg13g2_fill_1 FILLER_33_218 ();
 sg13g2_fill_1 FILLER_33_234 ();
 sg13g2_fill_1 FILLER_33_248 ();
 sg13g2_fill_2 FILLER_33_275 ();
 sg13g2_fill_1 FILLER_33_282 ();
 sg13g2_fill_2 FILLER_33_288 ();
 sg13g2_fill_1 FILLER_33_290 ();
 sg13g2_decap_4 FILLER_33_295 ();
 sg13g2_fill_1 FILLER_33_299 ();
 sg13g2_fill_2 FILLER_33_315 ();
 sg13g2_fill_1 FILLER_33_330 ();
 sg13g2_fill_1 FILLER_33_335 ();
 sg13g2_fill_1 FILLER_33_344 ();
 sg13g2_fill_1 FILLER_33_349 ();
 sg13g2_fill_1 FILLER_33_354 ();
 sg13g2_fill_1 FILLER_33_360 ();
 sg13g2_fill_2 FILLER_33_370 ();
 sg13g2_fill_2 FILLER_33_393 ();
 sg13g2_fill_2 FILLER_33_424 ();
 sg13g2_fill_1 FILLER_33_431 ();
 sg13g2_fill_1 FILLER_33_447 ();
 sg13g2_fill_1 FILLER_33_460 ();
 sg13g2_decap_4 FILLER_33_486 ();
 sg13g2_fill_1 FILLER_33_494 ();
 sg13g2_fill_2 FILLER_33_520 ();
 sg13g2_fill_1 FILLER_33_527 ();
 sg13g2_decap_8 FILLER_33_557 ();
 sg13g2_decap_8 FILLER_33_564 ();
 sg13g2_decap_8 FILLER_33_586 ();
 sg13g2_fill_1 FILLER_33_593 ();
 sg13g2_fill_1 FILLER_33_602 ();
 sg13g2_fill_2 FILLER_33_607 ();
 sg13g2_fill_1 FILLER_33_609 ();
 sg13g2_fill_1 FILLER_33_619 ();
 sg13g2_fill_1 FILLER_33_624 ();
 sg13g2_decap_8 FILLER_33_642 ();
 sg13g2_decap_4 FILLER_33_649 ();
 sg13g2_fill_2 FILLER_33_658 ();
 sg13g2_fill_2 FILLER_33_665 ();
 sg13g2_decap_8 FILLER_33_700 ();
 sg13g2_fill_1 FILLER_33_707 ();
 sg13g2_fill_1 FILLER_33_729 ();
 sg13g2_decap_8 FILLER_33_744 ();
 sg13g2_fill_2 FILLER_33_751 ();
 sg13g2_fill_1 FILLER_33_753 ();
 sg13g2_fill_2 FILLER_33_790 ();
 sg13g2_fill_1 FILLER_33_792 ();
 sg13g2_fill_1 FILLER_33_842 ();
 sg13g2_fill_2 FILLER_33_876 ();
 sg13g2_fill_2 FILLER_34_0 ();
 sg13g2_fill_1 FILLER_34_2 ();
 sg13g2_decap_4 FILLER_34_33 ();
 sg13g2_fill_2 FILLER_34_37 ();
 sg13g2_decap_8 FILLER_34_44 ();
 sg13g2_fill_1 FILLER_34_51 ();
 sg13g2_decap_4 FILLER_34_72 ();
 sg13g2_fill_1 FILLER_34_76 ();
 sg13g2_decap_8 FILLER_34_81 ();
 sg13g2_fill_1 FILLER_34_88 ();
 sg13g2_fill_2 FILLER_34_123 ();
 sg13g2_fill_1 FILLER_34_125 ();
 sg13g2_fill_2 FILLER_34_131 ();
 sg13g2_decap_8 FILLER_34_138 ();
 sg13g2_fill_1 FILLER_34_153 ();
 sg13g2_fill_1 FILLER_34_164 ();
 sg13g2_fill_1 FILLER_34_170 ();
 sg13g2_fill_1 FILLER_34_176 ();
 sg13g2_decap_8 FILLER_34_185 ();
 sg13g2_fill_2 FILLER_34_192 ();
 sg13g2_fill_1 FILLER_34_194 ();
 sg13g2_decap_4 FILLER_34_212 ();
 sg13g2_fill_1 FILLER_34_216 ();
 sg13g2_fill_1 FILLER_34_221 ();
 sg13g2_decap_8 FILLER_34_227 ();
 sg13g2_fill_2 FILLER_34_239 ();
 sg13g2_fill_1 FILLER_34_245 ();
 sg13g2_fill_2 FILLER_34_250 ();
 sg13g2_decap_4 FILLER_34_260 ();
 sg13g2_fill_2 FILLER_34_264 ();
 sg13g2_fill_2 FILLER_34_270 ();
 sg13g2_decap_8 FILLER_34_277 ();
 sg13g2_fill_2 FILLER_34_288 ();
 sg13g2_decap_8 FILLER_34_294 ();
 sg13g2_decap_8 FILLER_34_301 ();
 sg13g2_fill_2 FILLER_34_308 ();
 sg13g2_fill_1 FILLER_34_310 ();
 sg13g2_decap_4 FILLER_34_315 ();
 sg13g2_fill_1 FILLER_34_319 ();
 sg13g2_decap_4 FILLER_34_328 ();
 sg13g2_fill_1 FILLER_34_373 ();
 sg13g2_fill_1 FILLER_34_382 ();
 sg13g2_fill_1 FILLER_34_387 ();
 sg13g2_fill_2 FILLER_34_404 ();
 sg13g2_fill_1 FILLER_34_406 ();
 sg13g2_fill_2 FILLER_34_411 ();
 sg13g2_fill_1 FILLER_34_413 ();
 sg13g2_decap_4 FILLER_34_434 ();
 sg13g2_decap_8 FILLER_34_454 ();
 sg13g2_fill_2 FILLER_34_461 ();
 sg13g2_decap_4 FILLER_34_467 ();
 sg13g2_decap_4 FILLER_34_484 ();
 sg13g2_fill_1 FILLER_34_488 ();
 sg13g2_fill_1 FILLER_34_498 ();
 sg13g2_fill_1 FILLER_34_507 ();
 sg13g2_fill_1 FILLER_34_516 ();
 sg13g2_fill_2 FILLER_34_543 ();
 sg13g2_decap_8 FILLER_34_559 ();
 sg13g2_fill_1 FILLER_34_571 ();
 sg13g2_fill_2 FILLER_34_576 ();
 sg13g2_decap_8 FILLER_34_584 ();
 sg13g2_fill_2 FILLER_34_591 ();
 sg13g2_decap_4 FILLER_34_657 ();
 sg13g2_fill_2 FILLER_34_669 ();
 sg13g2_decap_8 FILLER_34_677 ();
 sg13g2_decap_8 FILLER_34_684 ();
 sg13g2_fill_2 FILLER_34_691 ();
 sg13g2_fill_1 FILLER_34_693 ();
 sg13g2_fill_1 FILLER_34_730 ();
 sg13g2_fill_1 FILLER_34_751 ();
 sg13g2_fill_2 FILLER_34_761 ();
 sg13g2_fill_2 FILLER_34_784 ();
 sg13g2_decap_4 FILLER_34_791 ();
 sg13g2_fill_1 FILLER_34_795 ();
 sg13g2_fill_2 FILLER_34_804 ();
 sg13g2_fill_1 FILLER_34_806 ();
 sg13g2_fill_1 FILLER_34_811 ();
 sg13g2_decap_4 FILLER_34_838 ();
 sg13g2_decap_4 FILLER_34_849 ();
 sg13g2_decap_4 FILLER_34_859 ();
 sg13g2_decap_4 FILLER_34_873 ();
 sg13g2_fill_1 FILLER_34_877 ();
 sg13g2_fill_1 FILLER_35_13 ();
 sg13g2_decap_8 FILLER_35_47 ();
 sg13g2_fill_1 FILLER_35_54 ();
 sg13g2_fill_2 FILLER_35_63 ();
 sg13g2_fill_1 FILLER_35_65 ();
 sg13g2_decap_4 FILLER_35_78 ();
 sg13g2_fill_2 FILLER_35_82 ();
 sg13g2_fill_1 FILLER_35_100 ();
 sg13g2_fill_2 FILLER_35_106 ();
 sg13g2_fill_1 FILLER_35_169 ();
 sg13g2_fill_2 FILLER_35_174 ();
 sg13g2_decap_4 FILLER_35_181 ();
 sg13g2_fill_1 FILLER_35_185 ();
 sg13g2_fill_2 FILLER_35_197 ();
 sg13g2_decap_4 FILLER_35_209 ();
 sg13g2_fill_2 FILLER_35_213 ();
 sg13g2_fill_1 FILLER_35_232 ();
 sg13g2_decap_8 FILLER_35_238 ();
 sg13g2_fill_1 FILLER_35_245 ();
 sg13g2_fill_2 FILLER_35_251 ();
 sg13g2_fill_1 FILLER_35_253 ();
 sg13g2_fill_1 FILLER_35_285 ();
 sg13g2_fill_1 FILLER_35_303 ();
 sg13g2_decap_4 FILLER_35_309 ();
 sg13g2_fill_2 FILLER_35_330 ();
 sg13g2_fill_1 FILLER_35_332 ();
 sg13g2_decap_8 FILLER_35_351 ();
 sg13g2_fill_1 FILLER_35_358 ();
 sg13g2_decap_4 FILLER_35_363 ();
 sg13g2_fill_1 FILLER_35_371 ();
 sg13g2_decap_8 FILLER_35_375 ();
 sg13g2_decap_8 FILLER_35_382 ();
 sg13g2_decap_4 FILLER_35_389 ();
 sg13g2_fill_2 FILLER_35_393 ();
 sg13g2_decap_4 FILLER_35_400 ();
 sg13g2_fill_2 FILLER_35_417 ();
 sg13g2_decap_8 FILLER_35_432 ();
 sg13g2_fill_1 FILLER_35_439 ();
 sg13g2_fill_2 FILLER_35_450 ();
 sg13g2_decap_8 FILLER_35_457 ();
 sg13g2_fill_2 FILLER_35_464 ();
 sg13g2_fill_2 FILLER_35_475 ();
 sg13g2_fill_1 FILLER_35_477 ();
 sg13g2_decap_4 FILLER_35_487 ();
 sg13g2_fill_1 FILLER_35_491 ();
 sg13g2_fill_1 FILLER_35_517 ();
 sg13g2_fill_2 FILLER_35_535 ();
 sg13g2_fill_1 FILLER_35_542 ();
 sg13g2_fill_2 FILLER_35_550 ();
 sg13g2_fill_1 FILLER_35_552 ();
 sg13g2_fill_2 FILLER_35_571 ();
 sg13g2_fill_1 FILLER_35_578 ();
 sg13g2_fill_2 FILLER_35_583 ();
 sg13g2_fill_1 FILLER_35_585 ();
 sg13g2_fill_2 FILLER_35_590 ();
 sg13g2_fill_1 FILLER_35_596 ();
 sg13g2_fill_1 FILLER_35_607 ();
 sg13g2_fill_1 FILLER_35_615 ();
 sg13g2_fill_1 FILLER_35_621 ();
 sg13g2_fill_2 FILLER_35_627 ();
 sg13g2_fill_2 FILLER_35_639 ();
 sg13g2_fill_1 FILLER_35_641 ();
 sg13g2_fill_2 FILLER_35_649 ();
 sg13g2_fill_1 FILLER_35_651 ();
 sg13g2_fill_1 FILLER_35_659 ();
 sg13g2_fill_1 FILLER_35_665 ();
 sg13g2_fill_1 FILLER_35_679 ();
 sg13g2_decap_8 FILLER_35_708 ();
 sg13g2_fill_2 FILLER_35_715 ();
 sg13g2_fill_1 FILLER_35_717 ();
 sg13g2_decap_4 FILLER_35_723 ();
 sg13g2_fill_2 FILLER_35_759 ();
 sg13g2_fill_1 FILLER_35_761 ();
 sg13g2_fill_1 FILLER_35_770 ();
 sg13g2_fill_1 FILLER_35_784 ();
 sg13g2_fill_2 FILLER_35_789 ();
 sg13g2_fill_1 FILLER_35_791 ();
 sg13g2_fill_1 FILLER_35_796 ();
 sg13g2_fill_1 FILLER_35_810 ();
 sg13g2_fill_2 FILLER_35_827 ();
 sg13g2_decap_4 FILLER_35_839 ();
 sg13g2_fill_1 FILLER_35_843 ();
 sg13g2_fill_2 FILLER_35_854 ();
 sg13g2_fill_2 FILLER_35_875 ();
 sg13g2_fill_1 FILLER_35_877 ();
 sg13g2_decap_4 FILLER_36_0 ();
 sg13g2_fill_1 FILLER_36_4 ();
 sg13g2_decap_8 FILLER_36_25 ();
 sg13g2_fill_1 FILLER_36_32 ();
 sg13g2_decap_8 FILLER_36_46 ();
 sg13g2_decap_8 FILLER_36_72 ();
 sg13g2_decap_4 FILLER_36_79 ();
 sg13g2_fill_2 FILLER_36_83 ();
 sg13g2_decap_8 FILLER_36_118 ();
 sg13g2_decap_4 FILLER_36_125 ();
 sg13g2_decap_8 FILLER_36_138 ();
 sg13g2_decap_8 FILLER_36_145 ();
 sg13g2_decap_8 FILLER_36_152 ();
 sg13g2_fill_2 FILLER_36_159 ();
 sg13g2_fill_1 FILLER_36_186 ();
 sg13g2_decap_4 FILLER_36_205 ();
 sg13g2_fill_2 FILLER_36_233 ();
 sg13g2_fill_2 FILLER_36_245 ();
 sg13g2_fill_1 FILLER_36_247 ();
 sg13g2_fill_2 FILLER_36_256 ();
 sg13g2_decap_4 FILLER_36_262 ();
 sg13g2_decap_8 FILLER_36_278 ();
 sg13g2_fill_1 FILLER_36_301 ();
 sg13g2_fill_1 FILLER_36_314 ();
 sg13g2_fill_1 FILLER_36_327 ();
 sg13g2_fill_1 FILLER_36_345 ();
 sg13g2_fill_1 FILLER_36_354 ();
 sg13g2_fill_1 FILLER_36_375 ();
 sg13g2_fill_1 FILLER_36_380 ();
 sg13g2_fill_2 FILLER_36_402 ();
 sg13g2_fill_1 FILLER_36_404 ();
 sg13g2_fill_2 FILLER_36_421 ();
 sg13g2_fill_1 FILLER_36_423 ();
 sg13g2_decap_8 FILLER_36_428 ();
 sg13g2_decap_4 FILLER_36_435 ();
 sg13g2_fill_1 FILLER_36_443 ();
 sg13g2_decap_8 FILLER_36_448 ();
 sg13g2_decap_4 FILLER_36_455 ();
 sg13g2_fill_2 FILLER_36_459 ();
 sg13g2_fill_1 FILLER_36_465 ();
 sg13g2_fill_1 FILLER_36_480 ();
 sg13g2_decap_4 FILLER_36_486 ();
 sg13g2_fill_1 FILLER_36_490 ();
 sg13g2_fill_1 FILLER_36_501 ();
 sg13g2_decap_8 FILLER_36_506 ();
 sg13g2_decap_8 FILLER_36_513 ();
 sg13g2_decap_8 FILLER_36_520 ();
 sg13g2_decap_4 FILLER_36_527 ();
 sg13g2_decap_4 FILLER_36_536 ();
 sg13g2_fill_2 FILLER_36_545 ();
 sg13g2_fill_2 FILLER_36_552 ();
 sg13g2_fill_1 FILLER_36_554 ();
 sg13g2_decap_4 FILLER_36_565 ();
 sg13g2_fill_1 FILLER_36_569 ();
 sg13g2_fill_2 FILLER_36_574 ();
 sg13g2_fill_1 FILLER_36_589 ();
 sg13g2_fill_1 FILLER_36_603 ();
 sg13g2_fill_1 FILLER_36_609 ();
 sg13g2_fill_1 FILLER_36_614 ();
 sg13g2_fill_2 FILLER_36_619 ();
 sg13g2_fill_2 FILLER_36_645 ();
 sg13g2_fill_1 FILLER_36_647 ();
 sg13g2_fill_2 FILLER_36_652 ();
 sg13g2_fill_1 FILLER_36_666 ();
 sg13g2_decap_8 FILLER_36_679 ();
 sg13g2_decap_4 FILLER_36_686 ();
 sg13g2_fill_1 FILLER_36_690 ();
 sg13g2_fill_1 FILLER_36_698 ();
 sg13g2_decap_4 FILLER_36_707 ();
 sg13g2_fill_2 FILLER_36_711 ();
 sg13g2_decap_8 FILLER_36_721 ();
 sg13g2_decap_4 FILLER_36_728 ();
 sg13g2_fill_1 FILLER_36_755 ();
 sg13g2_fill_1 FILLER_36_768 ();
 sg13g2_decap_4 FILLER_36_787 ();
 sg13g2_fill_2 FILLER_36_791 ();
 sg13g2_fill_2 FILLER_36_797 ();
 sg13g2_decap_4 FILLER_36_804 ();
 sg13g2_fill_1 FILLER_36_808 ();
 sg13g2_decap_4 FILLER_36_814 ();
 sg13g2_fill_1 FILLER_36_818 ();
 sg13g2_fill_1 FILLER_36_829 ();
 sg13g2_fill_1 FILLER_36_835 ();
 sg13g2_fill_2 FILLER_36_848 ();
 sg13g2_fill_1 FILLER_36_861 ();
 sg13g2_fill_2 FILLER_36_867 ();
 sg13g2_decap_8 FILLER_37_0 ();
 sg13g2_fill_2 FILLER_37_34 ();
 sg13g2_fill_1 FILLER_37_36 ();
 sg13g2_decap_8 FILLER_37_41 ();
 sg13g2_decap_8 FILLER_37_48 ();
 sg13g2_fill_1 FILLER_37_55 ();
 sg13g2_fill_1 FILLER_37_64 ();
 sg13g2_fill_2 FILLER_37_86 ();
 sg13g2_fill_2 FILLER_37_105 ();
 sg13g2_decap_8 FILLER_37_119 ();
 sg13g2_fill_2 FILLER_37_126 ();
 sg13g2_fill_1 FILLER_37_141 ();
 sg13g2_fill_2 FILLER_37_154 ();
 sg13g2_fill_1 FILLER_37_156 ();
 sg13g2_fill_1 FILLER_37_189 ();
 sg13g2_fill_2 FILLER_37_198 ();
 sg13g2_fill_1 FILLER_37_200 ();
 sg13g2_decap_8 FILLER_37_209 ();
 sg13g2_decap_8 FILLER_37_216 ();
 sg13g2_decap_4 FILLER_37_235 ();
 sg13g2_decap_4 FILLER_37_251 ();
 sg13g2_fill_2 FILLER_37_268 ();
 sg13g2_fill_1 FILLER_37_270 ();
 sg13g2_fill_2 FILLER_37_275 ();
 sg13g2_fill_1 FILLER_37_277 ();
 sg13g2_decap_4 FILLER_37_298 ();
 sg13g2_fill_2 FILLER_37_302 ();
 sg13g2_fill_1 FILLER_37_318 ();
 sg13g2_fill_2 FILLER_37_328 ();
 sg13g2_decap_8 FILLER_37_335 ();
 sg13g2_decap_8 FILLER_37_342 ();
 sg13g2_decap_8 FILLER_37_349 ();
 sg13g2_fill_1 FILLER_37_356 ();
 sg13g2_fill_2 FILLER_37_373 ();
 sg13g2_fill_1 FILLER_37_383 ();
 sg13g2_decap_8 FILLER_37_398 ();
 sg13g2_fill_2 FILLER_37_405 ();
 sg13g2_fill_1 FILLER_37_411 ();
 sg13g2_fill_1 FILLER_37_419 ();
 sg13g2_fill_1 FILLER_37_424 ();
 sg13g2_fill_1 FILLER_37_433 ();
 sg13g2_fill_2 FILLER_37_438 ();
 sg13g2_fill_1 FILLER_37_448 ();
 sg13g2_fill_2 FILLER_37_453 ();
 sg13g2_fill_1 FILLER_37_474 ();
 sg13g2_fill_1 FILLER_37_522 ();
 sg13g2_fill_2 FILLER_37_528 ();
 sg13g2_decap_8 FILLER_37_538 ();
 sg13g2_decap_8 FILLER_37_545 ();
 sg13g2_decap_8 FILLER_37_552 ();
 sg13g2_decap_4 FILLER_37_572 ();
 sg13g2_fill_1 FILLER_37_580 ();
 sg13g2_fill_1 FILLER_37_611 ();
 sg13g2_fill_2 FILLER_37_624 ();
 sg13g2_fill_1 FILLER_37_631 ();
 sg13g2_fill_2 FILLER_37_643 ();
 sg13g2_fill_1 FILLER_37_645 ();
 sg13g2_fill_2 FILLER_37_652 ();
 sg13g2_fill_2 FILLER_37_663 ();
 sg13g2_fill_1 FILLER_37_665 ();
 sg13g2_decap_8 FILLER_37_702 ();
 sg13g2_fill_2 FILLER_37_713 ();
 sg13g2_fill_1 FILLER_37_715 ();
 sg13g2_fill_1 FILLER_37_728 ();
 sg13g2_fill_1 FILLER_37_741 ();
 sg13g2_fill_1 FILLER_37_775 ();
 sg13g2_decap_8 FILLER_37_786 ();
 sg13g2_decap_8 FILLER_37_793 ();
 sg13g2_fill_1 FILLER_37_800 ();
 sg13g2_decap_4 FILLER_37_805 ();
 sg13g2_fill_1 FILLER_37_809 ();
 sg13g2_decap_4 FILLER_37_826 ();
 sg13g2_fill_2 FILLER_37_838 ();
 sg13g2_fill_1 FILLER_37_840 ();
 sg13g2_fill_2 FILLER_37_846 ();
 sg13g2_fill_2 FILLER_37_852 ();
 sg13g2_fill_1 FILLER_37_854 ();
 sg13g2_decap_8 FILLER_37_860 ();
 sg13g2_fill_2 FILLER_37_867 ();
 sg13g2_fill_1 FILLER_37_869 ();
 sg13g2_decap_4 FILLER_38_0 ();
 sg13g2_fill_2 FILLER_38_15 ();
 sg13g2_fill_1 FILLER_38_31 ();
 sg13g2_decap_8 FILLER_38_37 ();
 sg13g2_decap_8 FILLER_38_44 ();
 sg13g2_fill_1 FILLER_38_74 ();
 sg13g2_decap_8 FILLER_38_78 ();
 sg13g2_fill_2 FILLER_38_85 ();
 sg13g2_fill_1 FILLER_38_87 ();
 sg13g2_decap_8 FILLER_38_114 ();
 sg13g2_fill_2 FILLER_38_125 ();
 sg13g2_fill_2 FILLER_38_131 ();
 sg13g2_fill_1 FILLER_38_133 ();
 sg13g2_fill_1 FILLER_38_139 ();
 sg13g2_fill_2 FILLER_38_144 ();
 sg13g2_fill_1 FILLER_38_146 ();
 sg13g2_fill_2 FILLER_38_155 ();
 sg13g2_fill_1 FILLER_38_165 ();
 sg13g2_fill_2 FILLER_38_170 ();
 sg13g2_fill_1 FILLER_38_172 ();
 sg13g2_fill_1 FILLER_38_178 ();
 sg13g2_decap_4 FILLER_38_184 ();
 sg13g2_fill_2 FILLER_38_192 ();
 sg13g2_fill_2 FILLER_38_207 ();
 sg13g2_fill_1 FILLER_38_209 ();
 sg13g2_fill_1 FILLER_38_238 ();
 sg13g2_fill_1 FILLER_38_247 ();
 sg13g2_fill_2 FILLER_38_261 ();
 sg13g2_decap_8 FILLER_38_268 ();
 sg13g2_decap_4 FILLER_38_275 ();
 sg13g2_fill_1 FILLER_38_279 ();
 sg13g2_fill_1 FILLER_38_288 ();
 sg13g2_decap_8 FILLER_38_294 ();
 sg13g2_fill_1 FILLER_38_312 ();
 sg13g2_fill_2 FILLER_38_317 ();
 sg13g2_fill_1 FILLER_38_335 ();
 sg13g2_fill_2 FILLER_38_341 ();
 sg13g2_fill_1 FILLER_38_343 ();
 sg13g2_fill_1 FILLER_38_353 ();
 sg13g2_fill_2 FILLER_38_357 ();
 sg13g2_fill_2 FILLER_38_363 ();
 sg13g2_fill_2 FILLER_38_375 ();
 sg13g2_fill_1 FILLER_38_377 ();
 sg13g2_decap_8 FILLER_38_386 ();
 sg13g2_decap_4 FILLER_38_393 ();
 sg13g2_fill_1 FILLER_38_397 ();
 sg13g2_fill_2 FILLER_38_401 ();
 sg13g2_decap_8 FILLER_38_407 ();
 sg13g2_decap_8 FILLER_38_434 ();
 sg13g2_decap_8 FILLER_38_441 ();
 sg13g2_decap_4 FILLER_38_448 ();
 sg13g2_fill_1 FILLER_38_459 ();
 sg13g2_fill_1 FILLER_38_464 ();
 sg13g2_fill_1 FILLER_38_481 ();
 sg13g2_fill_1 FILLER_38_490 ();
 sg13g2_fill_1 FILLER_38_499 ();
 sg13g2_fill_2 FILLER_38_504 ();
 sg13g2_decap_4 FILLER_38_562 ();
 sg13g2_fill_2 FILLER_38_570 ();
 sg13g2_fill_1 FILLER_38_591 ();
 sg13g2_fill_2 FILLER_38_617 ();
 sg13g2_fill_1 FILLER_38_619 ();
 sg13g2_fill_1 FILLER_38_623 ();
 sg13g2_fill_2 FILLER_38_630 ();
 sg13g2_fill_1 FILLER_38_646 ();
 sg13g2_fill_2 FILLER_38_672 ();
 sg13g2_fill_1 FILLER_38_674 ();
 sg13g2_decap_8 FILLER_38_700 ();
 sg13g2_decap_8 FILLER_38_707 ();
 sg13g2_fill_1 FILLER_38_714 ();
 sg13g2_fill_2 FILLER_38_719 ();
 sg13g2_fill_1 FILLER_38_742 ();
 sg13g2_fill_2 FILLER_38_748 ();
 sg13g2_fill_1 FILLER_38_759 ();
 sg13g2_fill_1 FILLER_38_779 ();
 sg13g2_decap_4 FILLER_38_792 ();
 sg13g2_fill_1 FILLER_38_796 ();
 sg13g2_fill_1 FILLER_38_807 ();
 sg13g2_decap_4 FILLER_38_821 ();
 sg13g2_fill_2 FILLER_38_825 ();
 sg13g2_fill_2 FILLER_38_835 ();
 sg13g2_fill_1 FILLER_38_837 ();
 sg13g2_decap_8 FILLER_38_859 ();
 sg13g2_fill_1 FILLER_38_866 ();
 sg13g2_fill_1 FILLER_38_877 ();
 sg13g2_decap_4 FILLER_39_0 ();
 sg13g2_fill_1 FILLER_39_4 ();
 sg13g2_fill_1 FILLER_39_30 ();
 sg13g2_decap_8 FILLER_39_47 ();
 sg13g2_fill_2 FILLER_39_54 ();
 sg13g2_fill_1 FILLER_39_72 ();
 sg13g2_decap_4 FILLER_39_82 ();
 sg13g2_fill_1 FILLER_39_86 ();
 sg13g2_fill_2 FILLER_39_117 ();
 sg13g2_fill_1 FILLER_39_124 ();
 sg13g2_fill_1 FILLER_39_134 ();
 sg13g2_fill_1 FILLER_39_139 ();
 sg13g2_decap_4 FILLER_39_161 ();
 sg13g2_fill_2 FILLER_39_197 ();
 sg13g2_decap_8 FILLER_39_207 ();
 sg13g2_decap_8 FILLER_39_214 ();
 sg13g2_decap_4 FILLER_39_221 ();
 sg13g2_fill_1 FILLER_39_225 ();
 sg13g2_fill_2 FILLER_39_236 ();
 sg13g2_fill_1 FILLER_39_238 ();
 sg13g2_fill_1 FILLER_39_244 ();
 sg13g2_fill_2 FILLER_39_253 ();
 sg13g2_fill_2 FILLER_39_263 ();
 sg13g2_decap_8 FILLER_39_269 ();
 sg13g2_fill_2 FILLER_39_292 ();
 sg13g2_fill_1 FILLER_39_311 ();
 sg13g2_fill_1 FILLER_39_320 ();
 sg13g2_fill_1 FILLER_39_326 ();
 sg13g2_fill_1 FILLER_39_335 ();
 sg13g2_fill_2 FILLER_39_358 ();
 sg13g2_fill_1 FILLER_39_360 ();
 sg13g2_fill_1 FILLER_39_366 ();
 sg13g2_fill_2 FILLER_39_386 ();
 sg13g2_fill_1 FILLER_39_392 ();
 sg13g2_fill_1 FILLER_39_423 ();
 sg13g2_decap_8 FILLER_39_440 ();
 sg13g2_decap_4 FILLER_39_447 ();
 sg13g2_fill_2 FILLER_39_456 ();
 sg13g2_fill_1 FILLER_39_463 ();
 sg13g2_decap_8 FILLER_39_472 ();
 sg13g2_decap_4 FILLER_39_479 ();
 sg13g2_fill_1 FILLER_39_513 ();
 sg13g2_fill_1 FILLER_39_542 ();
 sg13g2_decap_4 FILLER_39_547 ();
 sg13g2_decap_4 FILLER_39_558 ();
 sg13g2_fill_2 FILLER_39_562 ();
 sg13g2_decap_4 FILLER_39_568 ();
 sg13g2_fill_1 FILLER_39_572 ();
 sg13g2_fill_1 FILLER_39_581 ();
 sg13g2_fill_1 FILLER_39_590 ();
 sg13g2_decap_4 FILLER_39_595 ();
 sg13g2_decap_4 FILLER_39_608 ();
 sg13g2_decap_4 FILLER_39_615 ();
 sg13g2_fill_1 FILLER_39_623 ();
 sg13g2_fill_2 FILLER_39_634 ();
 sg13g2_decap_8 FILLER_39_640 ();
 sg13g2_fill_2 FILLER_39_647 ();
 sg13g2_fill_1 FILLER_39_649 ();
 sg13g2_fill_1 FILLER_39_662 ();
 sg13g2_fill_1 FILLER_39_696 ();
 sg13g2_fill_2 FILLER_39_715 ();
 sg13g2_decap_4 FILLER_39_721 ();
 sg13g2_fill_1 FILLER_39_730 ();
 sg13g2_fill_2 FILLER_39_739 ();
 sg13g2_fill_1 FILLER_39_741 ();
 sg13g2_fill_2 FILLER_39_760 ();
 sg13g2_fill_1 FILLER_39_762 ();
 sg13g2_fill_2 FILLER_39_771 ();
 sg13g2_fill_1 FILLER_39_773 ();
 sg13g2_fill_2 FILLER_39_787 ();
 sg13g2_fill_1 FILLER_39_797 ();
 sg13g2_fill_2 FILLER_39_807 ();
 sg13g2_decap_4 FILLER_39_824 ();
 sg13g2_decap_4 FILLER_39_837 ();
 sg13g2_fill_2 FILLER_39_849 ();
 sg13g2_fill_1 FILLER_39_851 ();
 sg13g2_fill_2 FILLER_39_865 ();
 sg13g2_decap_4 FILLER_39_872 ();
 sg13g2_fill_2 FILLER_39_876 ();
 sg13g2_decap_8 FILLER_40_0 ();
 sg13g2_fill_1 FILLER_40_22 ();
 sg13g2_fill_1 FILLER_40_53 ();
 sg13g2_fill_1 FILLER_40_63 ();
 sg13g2_decap_8 FILLER_40_73 ();
 sg13g2_decap_8 FILLER_40_80 ();
 sg13g2_fill_2 FILLER_40_87 ();
 sg13g2_fill_2 FILLER_40_97 ();
 sg13g2_fill_2 FILLER_40_128 ();
 sg13g2_fill_1 FILLER_40_130 ();
 sg13g2_fill_2 FILLER_40_144 ();
 sg13g2_decap_4 FILLER_40_150 ();
 sg13g2_fill_2 FILLER_40_154 ();
 sg13g2_fill_1 FILLER_40_163 ();
 sg13g2_fill_1 FILLER_40_187 ();
 sg13g2_fill_2 FILLER_40_199 ();
 sg13g2_decap_4 FILLER_40_213 ();
 sg13g2_fill_1 FILLER_40_217 ();
 sg13g2_fill_1 FILLER_40_226 ();
 sg13g2_decap_4 FILLER_40_244 ();
 sg13g2_fill_2 FILLER_40_265 ();
 sg13g2_decap_4 FILLER_40_271 ();
 sg13g2_fill_1 FILLER_40_275 ();
 sg13g2_fill_1 FILLER_40_283 ();
 sg13g2_decap_8 FILLER_40_292 ();
 sg13g2_decap_8 FILLER_40_299 ();
 sg13g2_fill_1 FILLER_40_306 ();
 sg13g2_decap_8 FILLER_40_325 ();
 sg13g2_decap_4 FILLER_40_332 ();
 sg13g2_fill_1 FILLER_40_336 ();
 sg13g2_decap_8 FILLER_40_358 ();
 sg13g2_fill_1 FILLER_40_365 ();
 sg13g2_decap_4 FILLER_40_383 ();
 sg13g2_fill_1 FILLER_40_387 ();
 sg13g2_fill_2 FILLER_40_402 ();
 sg13g2_decap_4 FILLER_40_419 ();
 sg13g2_decap_8 FILLER_40_433 ();
 sg13g2_fill_1 FILLER_40_440 ();
 sg13g2_fill_2 FILLER_40_449 ();
 sg13g2_fill_2 FILLER_40_460 ();
 sg13g2_fill_1 FILLER_40_495 ();
 sg13g2_fill_2 FILLER_40_500 ();
 sg13g2_fill_1 FILLER_40_502 ();
 sg13g2_fill_2 FILLER_40_511 ();
 sg13g2_fill_1 FILLER_40_513 ();
 sg13g2_decap_8 FILLER_40_557 ();
 sg13g2_decap_4 FILLER_40_564 ();
 sg13g2_fill_1 FILLER_40_568 ();
 sg13g2_fill_2 FILLER_40_574 ();
 sg13g2_fill_1 FILLER_40_576 ();
 sg13g2_fill_1 FILLER_40_585 ();
 sg13g2_decap_4 FILLER_40_604 ();
 sg13g2_fill_1 FILLER_40_638 ();
 sg13g2_fill_2 FILLER_40_652 ();
 sg13g2_fill_2 FILLER_40_669 ();
 sg13g2_fill_1 FILLER_40_671 ();
 sg13g2_decap_4 FILLER_40_680 ();
 sg13g2_fill_1 FILLER_40_697 ();
 sg13g2_fill_1 FILLER_40_704 ();
 sg13g2_decap_8 FILLER_40_730 ();
 sg13g2_fill_2 FILLER_40_737 ();
 sg13g2_fill_1 FILLER_40_751 ();
 sg13g2_fill_2 FILLER_40_757 ();
 sg13g2_fill_1 FILLER_40_759 ();
 sg13g2_fill_2 FILLER_40_764 ();
 sg13g2_fill_2 FILLER_40_770 ();
 sg13g2_fill_2 FILLER_40_776 ();
 sg13g2_fill_1 FILLER_40_778 ();
 sg13g2_decap_8 FILLER_40_783 ();
 sg13g2_fill_2 FILLER_40_790 ();
 sg13g2_fill_1 FILLER_40_792 ();
 sg13g2_decap_8 FILLER_40_801 ();
 sg13g2_fill_1 FILLER_40_808 ();
 sg13g2_fill_1 FILLER_40_823 ();
 sg13g2_decap_4 FILLER_40_842 ();
 sg13g2_fill_2 FILLER_40_846 ();
 sg13g2_decap_4 FILLER_40_874 ();
 sg13g2_decap_8 FILLER_41_0 ();
 sg13g2_decap_8 FILLER_41_7 ();
 sg13g2_fill_2 FILLER_41_14 ();
 sg13g2_decap_8 FILLER_41_31 ();
 sg13g2_fill_1 FILLER_41_38 ();
 sg13g2_fill_2 FILLER_41_43 ();
 sg13g2_fill_1 FILLER_41_45 ();
 sg13g2_decap_4 FILLER_41_50 ();
 sg13g2_decap_4 FILLER_41_80 ();
 sg13g2_fill_1 FILLER_41_84 ();
 sg13g2_fill_1 FILLER_41_97 ();
 sg13g2_fill_1 FILLER_41_111 ();
 sg13g2_decap_4 FILLER_41_118 ();
 sg13g2_decap_8 FILLER_41_127 ();
 sg13g2_decap_8 FILLER_41_134 ();
 sg13g2_decap_8 FILLER_41_146 ();
 sg13g2_decap_4 FILLER_41_153 ();
 sg13g2_fill_2 FILLER_41_183 ();
 sg13g2_fill_1 FILLER_41_185 ();
 sg13g2_fill_1 FILLER_41_194 ();
 sg13g2_fill_1 FILLER_41_203 ();
 sg13g2_decap_4 FILLER_41_220 ();
 sg13g2_fill_1 FILLER_41_224 ();
 sg13g2_fill_1 FILLER_41_246 ();
 sg13g2_fill_2 FILLER_41_273 ();
 sg13g2_fill_1 FILLER_41_275 ();
 sg13g2_fill_1 FILLER_41_284 ();
 sg13g2_fill_2 FILLER_41_301 ();
 sg13g2_fill_1 FILLER_41_321 ();
 sg13g2_fill_1 FILLER_41_326 ();
 sg13g2_fill_2 FILLER_41_339 ();
 sg13g2_fill_1 FILLER_41_349 ();
 sg13g2_decap_8 FILLER_41_354 ();
 sg13g2_decap_8 FILLER_41_361 ();
 sg13g2_decap_8 FILLER_41_368 ();
 sg13g2_fill_1 FILLER_41_387 ();
 sg13g2_fill_2 FILLER_41_416 ();
 sg13g2_decap_4 FILLER_41_442 ();
 sg13g2_fill_2 FILLER_41_446 ();
 sg13g2_fill_1 FILLER_41_451 ();
 sg13g2_fill_2 FILLER_41_472 ();
 sg13g2_fill_1 FILLER_41_474 ();
 sg13g2_decap_4 FILLER_41_479 ();
 sg13g2_decap_4 FILLER_41_492 ();
 sg13g2_fill_1 FILLER_41_496 ();
 sg13g2_fill_2 FILLER_41_502 ();
 sg13g2_fill_2 FILLER_41_508 ();
 sg13g2_fill_1 FILLER_41_510 ();
 sg13g2_fill_2 FILLER_41_519 ();
 sg13g2_fill_2 FILLER_41_530 ();
 sg13g2_fill_1 FILLER_41_549 ();
 sg13g2_fill_2 FILLER_41_554 ();
 sg13g2_fill_2 FILLER_41_565 ();
 sg13g2_fill_1 FILLER_41_571 ();
 sg13g2_decap_4 FILLER_41_589 ();
 sg13g2_decap_4 FILLER_41_625 ();
 sg13g2_fill_2 FILLER_41_653 ();
 sg13g2_fill_2 FILLER_41_668 ();
 sg13g2_fill_2 FILLER_41_674 ();
 sg13g2_fill_2 FILLER_41_680 ();
 sg13g2_decap_4 FILLER_41_690 ();
 sg13g2_fill_2 FILLER_41_694 ();
 sg13g2_decap_4 FILLER_41_700 ();
 sg13g2_fill_1 FILLER_41_704 ();
 sg13g2_decap_4 FILLER_41_714 ();
 sg13g2_fill_2 FILLER_41_740 ();
 sg13g2_fill_1 FILLER_41_773 ();
 sg13g2_fill_2 FILLER_41_778 ();
 sg13g2_fill_2 FILLER_41_785 ();
 sg13g2_fill_1 FILLER_41_787 ();
 sg13g2_fill_2 FILLER_41_795 ();
 sg13g2_fill_1 FILLER_41_797 ();
 sg13g2_decap_8 FILLER_41_803 ();
 sg13g2_fill_1 FILLER_41_810 ();
 sg13g2_fill_1 FILLER_41_833 ();
 sg13g2_fill_2 FILLER_41_842 ();
 sg13g2_fill_1 FILLER_41_852 ();
 sg13g2_fill_2 FILLER_41_858 ();
 sg13g2_decap_4 FILLER_41_873 ();
 sg13g2_fill_1 FILLER_41_877 ();
 sg13g2_decap_8 FILLER_42_0 ();
 sg13g2_fill_2 FILLER_42_30 ();
 sg13g2_fill_1 FILLER_42_32 ();
 sg13g2_fill_1 FILLER_42_43 ();
 sg13g2_decap_4 FILLER_42_52 ();
 sg13g2_decap_8 FILLER_42_68 ();
 sg13g2_decap_8 FILLER_42_75 ();
 sg13g2_decap_4 FILLER_42_82 ();
 sg13g2_fill_2 FILLER_42_86 ();
 sg13g2_decap_4 FILLER_42_104 ();
 sg13g2_fill_1 FILLER_42_108 ();
 sg13g2_fill_2 FILLER_42_121 ();
 sg13g2_fill_1 FILLER_42_123 ();
 sg13g2_fill_1 FILLER_42_132 ();
 sg13g2_fill_2 FILLER_42_148 ();
 sg13g2_fill_2 FILLER_42_155 ();
 sg13g2_fill_2 FILLER_42_162 ();
 sg13g2_fill_2 FILLER_42_168 ();
 sg13g2_fill_1 FILLER_42_170 ();
 sg13g2_fill_1 FILLER_42_179 ();
 sg13g2_fill_2 FILLER_42_188 ();
 sg13g2_fill_2 FILLER_42_197 ();
 sg13g2_fill_2 FILLER_42_204 ();
 sg13g2_fill_1 FILLER_42_206 ();
 sg13g2_decap_4 FILLER_42_223 ();
 sg13g2_fill_1 FILLER_42_227 ();
 sg13g2_decap_8 FILLER_42_246 ();
 sg13g2_fill_1 FILLER_42_253 ();
 sg13g2_fill_1 FILLER_42_267 ();
 sg13g2_fill_1 FILLER_42_272 ();
 sg13g2_fill_2 FILLER_42_291 ();
 sg13g2_fill_1 FILLER_42_293 ();
 sg13g2_fill_1 FILLER_42_299 ();
 sg13g2_decap_8 FILLER_42_317 ();
 sg13g2_decap_8 FILLER_42_324 ();
 sg13g2_decap_4 FILLER_42_331 ();
 sg13g2_fill_1 FILLER_42_335 ();
 sg13g2_fill_1 FILLER_42_341 ();
 sg13g2_fill_2 FILLER_42_347 ();
 sg13g2_fill_1 FILLER_42_349 ();
 sg13g2_fill_2 FILLER_42_367 ();
 sg13g2_fill_1 FILLER_42_369 ();
 sg13g2_decap_4 FILLER_42_380 ();
 sg13g2_decap_8 FILLER_42_402 ();
 sg13g2_fill_2 FILLER_42_421 ();
 sg13g2_fill_1 FILLER_42_423 ();
 sg13g2_decap_4 FILLER_42_428 ();
 sg13g2_decap_4 FILLER_42_442 ();
 sg13g2_fill_2 FILLER_42_446 ();
 sg13g2_decap_8 FILLER_42_459 ();
 sg13g2_decap_8 FILLER_42_466 ();
 sg13g2_decap_8 FILLER_42_473 ();
 sg13g2_decap_8 FILLER_42_480 ();
 sg13g2_decap_4 FILLER_42_487 ();
 sg13g2_fill_1 FILLER_42_491 ();
 sg13g2_fill_1 FILLER_42_497 ();
 sg13g2_fill_2 FILLER_42_507 ();
 sg13g2_fill_1 FILLER_42_509 ();
 sg13g2_fill_1 FILLER_42_534 ();
 sg13g2_fill_1 FILLER_42_543 ();
 sg13g2_decap_8 FILLER_42_553 ();
 sg13g2_decap_8 FILLER_42_560 ();
 sg13g2_decap_4 FILLER_42_567 ();
 sg13g2_fill_1 FILLER_42_571 ();
 sg13g2_decap_8 FILLER_42_595 ();
 sg13g2_fill_2 FILLER_42_602 ();
 sg13g2_fill_1 FILLER_42_620 ();
 sg13g2_fill_1 FILLER_42_663 ();
 sg13g2_fill_1 FILLER_42_675 ();
 sg13g2_fill_1 FILLER_42_681 ();
 sg13g2_fill_2 FILLER_42_702 ();
 sg13g2_fill_1 FILLER_42_704 ();
 sg13g2_fill_1 FILLER_42_710 ();
 sg13g2_fill_2 FILLER_42_742 ();
 sg13g2_fill_1 FILLER_42_744 ();
 sg13g2_fill_2 FILLER_42_767 ();
 sg13g2_fill_1 FILLER_42_769 ();
 sg13g2_decap_8 FILLER_42_774 ();
 sg13g2_fill_1 FILLER_42_781 ();
 sg13g2_fill_2 FILLER_42_791 ();
 sg13g2_fill_1 FILLER_42_793 ();
 sg13g2_decap_4 FILLER_42_798 ();
 sg13g2_fill_1 FILLER_42_802 ();
 sg13g2_fill_2 FILLER_42_807 ();
 sg13g2_fill_1 FILLER_42_809 ();
 sg13g2_decap_8 FILLER_42_814 ();
 sg13g2_decap_8 FILLER_42_821 ();
 sg13g2_fill_1 FILLER_42_828 ();
 sg13g2_decap_8 FILLER_42_834 ();
 sg13g2_decap_4 FILLER_42_841 ();
 sg13g2_fill_2 FILLER_42_845 ();
 sg13g2_decap_4 FILLER_42_852 ();
 sg13g2_fill_1 FILLER_42_856 ();
 sg13g2_decap_4 FILLER_42_873 ();
 sg13g2_fill_1 FILLER_42_877 ();
 sg13g2_fill_1 FILLER_43_0 ();
 sg13g2_fill_1 FILLER_43_7 ();
 sg13g2_fill_2 FILLER_43_26 ();
 sg13g2_decap_4 FILLER_43_38 ();
 sg13g2_decap_8 FILLER_43_46 ();
 sg13g2_decap_8 FILLER_43_79 ();
 sg13g2_fill_1 FILLER_43_86 ();
 sg13g2_fill_2 FILLER_43_99 ();
 sg13g2_fill_1 FILLER_43_101 ();
 sg13g2_fill_2 FILLER_43_117 ();
 sg13g2_fill_1 FILLER_43_162 ();
 sg13g2_fill_1 FILLER_43_167 ();
 sg13g2_fill_1 FILLER_43_173 ();
 sg13g2_fill_1 FILLER_43_178 ();
 sg13g2_decap_8 FILLER_43_192 ();
 sg13g2_decap_8 FILLER_43_199 ();
 sg13g2_fill_2 FILLER_43_206 ();
 sg13g2_decap_8 FILLER_43_237 ();
 sg13g2_fill_2 FILLER_43_244 ();
 sg13g2_fill_1 FILLER_43_246 ();
 sg13g2_fill_2 FILLER_43_255 ();
 sg13g2_fill_1 FILLER_43_265 ();
 sg13g2_fill_1 FILLER_43_270 ();
 sg13g2_fill_1 FILLER_43_279 ();
 sg13g2_fill_1 FILLER_43_284 ();
 sg13g2_decap_8 FILLER_43_303 ();
 sg13g2_fill_1 FILLER_43_310 ();
 sg13g2_fill_2 FILLER_43_324 ();
 sg13g2_decap_4 FILLER_43_331 ();
 sg13g2_fill_1 FILLER_43_335 ();
 sg13g2_fill_1 FILLER_43_341 ();
 sg13g2_decap_8 FILLER_43_350 ();
 sg13g2_decap_4 FILLER_43_357 ();
 sg13g2_fill_1 FILLER_43_361 ();
 sg13g2_decap_8 FILLER_43_374 ();
 sg13g2_decap_4 FILLER_43_381 ();
 sg13g2_decap_4 FILLER_43_401 ();
 sg13g2_fill_2 FILLER_43_405 ();
 sg13g2_fill_2 FILLER_43_419 ();
 sg13g2_decap_8 FILLER_43_433 ();
 sg13g2_decap_8 FILLER_43_440 ();
 sg13g2_fill_1 FILLER_43_447 ();
 sg13g2_fill_1 FILLER_43_506 ();
 sg13g2_decap_4 FILLER_43_520 ();
 sg13g2_fill_1 FILLER_43_524 ();
 sg13g2_fill_1 FILLER_43_545 ();
 sg13g2_fill_2 FILLER_43_556 ();
 sg13g2_decap_8 FILLER_43_563 ();
 sg13g2_decap_8 FILLER_43_579 ();
 sg13g2_fill_1 FILLER_43_591 ();
 sg13g2_decap_4 FILLER_43_601 ();
 sg13g2_fill_1 FILLER_43_605 ();
 sg13g2_fill_2 FILLER_43_618 ();
 sg13g2_fill_1 FILLER_43_620 ();
 sg13g2_fill_2 FILLER_43_626 ();
 sg13g2_fill_1 FILLER_43_628 ();
 sg13g2_decap_8 FILLER_43_643 ();
 sg13g2_fill_2 FILLER_43_650 ();
 sg13g2_decap_4 FILLER_43_661 ();
 sg13g2_fill_2 FILLER_43_679 ();
 sg13g2_fill_2 FILLER_43_699 ();
 sg13g2_fill_2 FILLER_43_747 ();
 sg13g2_fill_1 FILLER_43_755 ();
 sg13g2_decap_8 FILLER_43_761 ();
 sg13g2_fill_2 FILLER_43_768 ();
 sg13g2_fill_1 FILLER_43_770 ();
 sg13g2_fill_1 FILLER_43_775 ();
 sg13g2_fill_1 FILLER_43_781 ();
 sg13g2_decap_8 FILLER_43_796 ();
 sg13g2_fill_1 FILLER_43_803 ();
 sg13g2_decap_4 FILLER_43_825 ();
 sg13g2_fill_1 FILLER_43_829 ();
 sg13g2_fill_2 FILLER_43_834 ();
 sg13g2_decap_8 FILLER_43_840 ();
 sg13g2_decap_4 FILLER_43_847 ();
 sg13g2_fill_2 FILLER_43_851 ();
 sg13g2_fill_1 FILLER_43_877 ();
 sg13g2_decap_4 FILLER_44_0 ();
 sg13g2_fill_2 FILLER_44_16 ();
 sg13g2_fill_1 FILLER_44_18 ();
 sg13g2_fill_2 FILLER_44_46 ();
 sg13g2_decap_4 FILLER_44_52 ();
 sg13g2_fill_1 FILLER_44_66 ();
 sg13g2_decap_8 FILLER_44_78 ();
 sg13g2_decap_8 FILLER_44_85 ();
 sg13g2_decap_4 FILLER_44_92 ();
 sg13g2_fill_2 FILLER_44_96 ();
 sg13g2_fill_1 FILLER_44_111 ();
 sg13g2_decap_4 FILLER_44_134 ();
 sg13g2_fill_2 FILLER_44_138 ();
 sg13g2_fill_1 FILLER_44_145 ();
 sg13g2_fill_2 FILLER_44_151 ();
 sg13g2_fill_1 FILLER_44_157 ();
 sg13g2_fill_2 FILLER_44_163 ();
 sg13g2_fill_2 FILLER_44_168 ();
 sg13g2_fill_2 FILLER_44_174 ();
 sg13g2_fill_1 FILLER_44_184 ();
 sg13g2_decap_8 FILLER_44_190 ();
 sg13g2_decap_8 FILLER_44_197 ();
 sg13g2_decap_4 FILLER_44_204 ();
 sg13g2_decap_8 FILLER_44_213 ();
 sg13g2_fill_2 FILLER_44_220 ();
 sg13g2_fill_1 FILLER_44_222 ();
 sg13g2_decap_4 FILLER_44_227 ();
 sg13g2_decap_4 FILLER_44_235 ();
 sg13g2_decap_8 FILLER_44_247 ();
 sg13g2_decap_8 FILLER_44_254 ();
 sg13g2_fill_2 FILLER_44_261 ();
 sg13g2_fill_1 FILLER_44_267 ();
 sg13g2_fill_2 FILLER_44_280 ();
 sg13g2_decap_4 FILLER_44_296 ();
 sg13g2_fill_2 FILLER_44_300 ();
 sg13g2_fill_1 FILLER_44_306 ();
 sg13g2_fill_1 FILLER_44_315 ();
 sg13g2_fill_1 FILLER_44_340 ();
 sg13g2_fill_2 FILLER_44_348 ();
 sg13g2_decap_4 FILLER_44_381 ();
 sg13g2_fill_1 FILLER_44_385 ();
 sg13g2_fill_2 FILLER_44_390 ();
 sg13g2_fill_1 FILLER_44_392 ();
 sg13g2_fill_1 FILLER_44_398 ();
 sg13g2_fill_1 FILLER_44_407 ();
 sg13g2_fill_1 FILLER_44_413 ();
 sg13g2_fill_1 FILLER_44_419 ();
 sg13g2_fill_1 FILLER_44_428 ();
 sg13g2_fill_2 FILLER_44_434 ();
 sg13g2_decap_8 FILLER_44_484 ();
 sg13g2_fill_2 FILLER_44_491 ();
 sg13g2_decap_4 FILLER_44_498 ();
 sg13g2_fill_2 FILLER_44_502 ();
 sg13g2_fill_2 FILLER_44_517 ();
 sg13g2_fill_1 FILLER_44_519 ();
 sg13g2_fill_2 FILLER_44_562 ();
 sg13g2_decap_8 FILLER_44_600 ();
 sg13g2_fill_1 FILLER_44_622 ();
 sg13g2_fill_2 FILLER_44_634 ();
 sg13g2_decap_8 FILLER_44_653 ();
 sg13g2_fill_2 FILLER_44_730 ();
 sg13g2_fill_1 FILLER_44_739 ();
 sg13g2_fill_1 FILLER_44_744 ();
 sg13g2_fill_1 FILLER_44_761 ();
 sg13g2_fill_1 FILLER_44_767 ();
 sg13g2_fill_1 FILLER_44_774 ();
 sg13g2_decap_4 FILLER_44_786 ();
 sg13g2_fill_1 FILLER_44_795 ();
 sg13g2_fill_2 FILLER_44_801 ();
 sg13g2_decap_4 FILLER_44_819 ();
 sg13g2_fill_1 FILLER_44_823 ();
 sg13g2_decap_8 FILLER_44_844 ();
 sg13g2_decap_8 FILLER_44_851 ();
 sg13g2_fill_2 FILLER_44_858 ();
 sg13g2_fill_1 FILLER_44_860 ();
 sg13g2_fill_1 FILLER_44_877 ();
 sg13g2_decap_4 FILLER_45_0 ();
 sg13g2_fill_1 FILLER_45_4 ();
 sg13g2_decap_8 FILLER_45_10 ();
 sg13g2_decap_8 FILLER_45_17 ();
 sg13g2_decap_4 FILLER_45_28 ();
 sg13g2_fill_1 FILLER_45_32 ();
 sg13g2_decap_8 FILLER_45_41 ();
 sg13g2_fill_1 FILLER_45_48 ();
 sg13g2_fill_1 FILLER_45_66 ();
 sg13g2_decap_4 FILLER_45_77 ();
 sg13g2_fill_1 FILLER_45_81 ();
 sg13g2_fill_1 FILLER_45_92 ();
 sg13g2_fill_1 FILLER_45_101 ();
 sg13g2_fill_2 FILLER_45_111 ();
 sg13g2_fill_1 FILLER_45_113 ();
 sg13g2_fill_2 FILLER_45_144 ();
 sg13g2_fill_2 FILLER_45_154 ();
 sg13g2_fill_1 FILLER_45_173 ();
 sg13g2_fill_2 FILLER_45_198 ();
 sg13g2_fill_2 FILLER_45_213 ();
 sg13g2_fill_1 FILLER_45_215 ();
 sg13g2_fill_2 FILLER_45_247 ();
 sg13g2_fill_1 FILLER_45_249 ();
 sg13g2_fill_2 FILLER_45_280 ();
 sg13g2_fill_2 FILLER_45_286 ();
 sg13g2_fill_2 FILLER_45_296 ();
 sg13g2_fill_1 FILLER_45_298 ();
 sg13g2_fill_1 FILLER_45_303 ();
 sg13g2_fill_2 FILLER_45_308 ();
 sg13g2_fill_2 FILLER_45_319 ();
 sg13g2_fill_1 FILLER_45_326 ();
 sg13g2_decap_4 FILLER_45_332 ();
 sg13g2_fill_1 FILLER_45_336 ();
 sg13g2_fill_2 FILLER_45_341 ();
 sg13g2_decap_4 FILLER_45_352 ();
 sg13g2_fill_2 FILLER_45_377 ();
 sg13g2_fill_2 FILLER_45_437 ();
 sg13g2_fill_2 FILLER_45_447 ();
 sg13g2_fill_2 FILLER_45_453 ();
 sg13g2_fill_1 FILLER_45_455 ();
 sg13g2_fill_2 FILLER_45_464 ();
 sg13g2_fill_1 FILLER_45_466 ();
 sg13g2_fill_2 FILLER_45_472 ();
 sg13g2_decap_4 FILLER_45_514 ();
 sg13g2_fill_1 FILLER_45_518 ();
 sg13g2_fill_1 FILLER_45_528 ();
 sg13g2_fill_2 FILLER_45_533 ();
 sg13g2_fill_2 FILLER_45_548 ();
 sg13g2_decap_4 FILLER_45_558 ();
 sg13g2_fill_2 FILLER_45_562 ();
 sg13g2_fill_1 FILLER_45_572 ();
 sg13g2_fill_1 FILLER_45_577 ();
 sg13g2_fill_2 FILLER_45_586 ();
 sg13g2_fill_1 FILLER_45_596 ();
 sg13g2_fill_2 FILLER_45_601 ();
 sg13g2_fill_1 FILLER_45_607 ();
 sg13g2_fill_2 FILLER_45_618 ();
 sg13g2_fill_1 FILLER_45_632 ();
 sg13g2_fill_1 FILLER_45_667 ();
 sg13g2_fill_1 FILLER_45_689 ();
 sg13g2_fill_2 FILLER_45_724 ();
 sg13g2_fill_1 FILLER_45_726 ();
 sg13g2_fill_2 FILLER_45_738 ();
 sg13g2_fill_1 FILLER_45_781 ();
 sg13g2_fill_1 FILLER_45_791 ();
 sg13g2_decap_4 FILLER_45_797 ();
 sg13g2_fill_1 FILLER_45_821 ();
 sg13g2_fill_2 FILLER_45_832 ();
 sg13g2_fill_1 FILLER_45_834 ();
 sg13g2_fill_2 FILLER_45_859 ();
 sg13g2_decap_8 FILLER_45_869 ();
 sg13g2_fill_2 FILLER_45_876 ();
 sg13g2_fill_2 FILLER_46_0 ();
 sg13g2_fill_1 FILLER_46_12 ();
 sg13g2_fill_1 FILLER_46_27 ();
 sg13g2_fill_1 FILLER_46_36 ();
 sg13g2_fill_2 FILLER_46_51 ();
 sg13g2_fill_1 FILLER_46_53 ();
 sg13g2_fill_1 FILLER_46_81 ();
 sg13g2_fill_1 FILLER_46_123 ();
 sg13g2_fill_1 FILLER_46_129 ();
 sg13g2_decap_8 FILLER_46_134 ();
 sg13g2_decap_8 FILLER_46_141 ();
 sg13g2_fill_2 FILLER_46_148 ();
 sg13g2_fill_1 FILLER_46_158 ();
 sg13g2_fill_1 FILLER_46_169 ();
 sg13g2_fill_1 FILLER_46_176 ();
 sg13g2_decap_8 FILLER_46_194 ();
 sg13g2_decap_4 FILLER_46_201 ();
 sg13g2_fill_1 FILLER_46_205 ();
 sg13g2_fill_1 FILLER_46_214 ();
 sg13g2_decap_4 FILLER_46_223 ();
 sg13g2_fill_1 FILLER_46_227 ();
 sg13g2_fill_1 FILLER_46_232 ();
 sg13g2_decap_4 FILLER_46_259 ();
 sg13g2_fill_1 FILLER_46_271 ();
 sg13g2_fill_1 FILLER_46_292 ();
 sg13g2_decap_8 FILLER_46_297 ();
 sg13g2_fill_1 FILLER_46_304 ();
 sg13g2_fill_1 FILLER_46_310 ();
 sg13g2_fill_2 FILLER_46_325 ();
 sg13g2_fill_2 FILLER_46_335 ();
 sg13g2_fill_1 FILLER_46_337 ();
 sg13g2_fill_2 FILLER_46_342 ();
 sg13g2_fill_2 FILLER_46_349 ();
 sg13g2_fill_1 FILLER_46_361 ();
 sg13g2_decap_4 FILLER_46_385 ();
 sg13g2_fill_2 FILLER_46_389 ();
 sg13g2_fill_2 FILLER_46_422 ();
 sg13g2_fill_2 FILLER_46_428 ();
 sg13g2_fill_1 FILLER_46_430 ();
 sg13g2_fill_2 FILLER_46_445 ();
 sg13g2_decap_4 FILLER_46_454 ();
 sg13g2_decap_4 FILLER_46_463 ();
 sg13g2_fill_2 FILLER_46_475 ();
 sg13g2_fill_1 FILLER_46_477 ();
 sg13g2_fill_1 FILLER_46_482 ();
 sg13g2_fill_2 FILLER_46_491 ();
 sg13g2_fill_2 FILLER_46_501 ();
 sg13g2_fill_1 FILLER_46_503 ();
 sg13g2_fill_1 FILLER_46_508 ();
 sg13g2_fill_2 FILLER_46_513 ();
 sg13g2_fill_1 FILLER_46_515 ();
 sg13g2_fill_2 FILLER_46_540 ();
 sg13g2_fill_1 FILLER_46_542 ();
 sg13g2_decap_8 FILLER_46_555 ();
 sg13g2_fill_2 FILLER_46_575 ();
 sg13g2_fill_1 FILLER_46_590 ();
 sg13g2_fill_2 FILLER_46_596 ();
 sg13g2_fill_1 FILLER_46_598 ();
 sg13g2_fill_1 FILLER_46_614 ();
 sg13g2_decap_4 FILLER_46_619 ();
 sg13g2_fill_1 FILLER_46_634 ();
 sg13g2_decap_4 FILLER_46_651 ();
 sg13g2_fill_1 FILLER_46_655 ();
 sg13g2_decap_4 FILLER_46_664 ();
 sg13g2_fill_1 FILLER_46_668 ();
 sg13g2_fill_1 FILLER_46_723 ();
 sg13g2_fill_2 FILLER_46_744 ();
 sg13g2_decap_8 FILLER_46_754 ();
 sg13g2_fill_1 FILLER_46_771 ();
 sg13g2_fill_1 FILLER_46_794 ();
 sg13g2_fill_2 FILLER_46_809 ();
 sg13g2_decap_8 FILLER_46_815 ();
 sg13g2_decap_4 FILLER_46_832 ();
 sg13g2_fill_2 FILLER_46_836 ();
 sg13g2_decap_4 FILLER_46_874 ();
 sg13g2_fill_2 FILLER_47_0 ();
 sg13g2_fill_1 FILLER_47_2 ();
 sg13g2_fill_2 FILLER_47_22 ();
 sg13g2_fill_1 FILLER_47_24 ();
 sg13g2_fill_1 FILLER_47_30 ();
 sg13g2_fill_1 FILLER_47_75 ();
 sg13g2_fill_1 FILLER_47_81 ();
 sg13g2_fill_2 FILLER_47_87 ();
 sg13g2_fill_1 FILLER_47_89 ();
 sg13g2_fill_1 FILLER_47_105 ();
 sg13g2_fill_2 FILLER_47_125 ();
 sg13g2_fill_1 FILLER_47_147 ();
 sg13g2_decap_4 FILLER_47_156 ();
 sg13g2_fill_2 FILLER_47_160 ();
 sg13g2_fill_1 FILLER_47_167 ();
 sg13g2_fill_2 FILLER_47_197 ();
 sg13g2_fill_1 FILLER_47_199 ();
 sg13g2_fill_1 FILLER_47_216 ();
 sg13g2_fill_2 FILLER_47_245 ();
 sg13g2_fill_1 FILLER_47_255 ();
 sg13g2_decap_4 FILLER_47_268 ();
 sg13g2_fill_2 FILLER_47_272 ();
 sg13g2_fill_1 FILLER_47_278 ();
 sg13g2_fill_1 FILLER_47_283 ();
 sg13g2_fill_2 FILLER_47_304 ();
 sg13g2_fill_1 FILLER_47_306 ();
 sg13g2_decap_8 FILLER_47_334 ();
 sg13g2_fill_2 FILLER_47_341 ();
 sg13g2_fill_1 FILLER_47_343 ();
 sg13g2_fill_2 FILLER_47_348 ();
 sg13g2_fill_2 FILLER_47_372 ();
 sg13g2_fill_1 FILLER_47_387 ();
 sg13g2_fill_2 FILLER_47_393 ();
 sg13g2_fill_1 FILLER_47_395 ();
 sg13g2_fill_2 FILLER_47_400 ();
 sg13g2_decap_4 FILLER_47_414 ();
 sg13g2_decap_8 FILLER_47_440 ();
 sg13g2_decap_8 FILLER_47_447 ();
 sg13g2_decap_4 FILLER_47_454 ();
 sg13g2_decap_4 FILLER_47_468 ();
 sg13g2_fill_1 FILLER_47_472 ();
 sg13g2_fill_1 FILLER_47_494 ();
 sg13g2_fill_1 FILLER_47_503 ();
 sg13g2_fill_1 FILLER_47_510 ();
 sg13g2_decap_4 FILLER_47_516 ();
 sg13g2_fill_2 FILLER_47_525 ();
 sg13g2_fill_1 FILLER_47_527 ();
 sg13g2_decap_8 FILLER_47_542 ();
 sg13g2_fill_1 FILLER_47_549 ();
 sg13g2_fill_2 FILLER_47_563 ();
 sg13g2_decap_4 FILLER_47_572 ();
 sg13g2_fill_2 FILLER_47_576 ();
 sg13g2_decap_4 FILLER_47_583 ();
 sg13g2_fill_1 FILLER_47_587 ();
 sg13g2_fill_2 FILLER_47_593 ();
 sg13g2_decap_4 FILLER_47_603 ();
 sg13g2_fill_2 FILLER_47_607 ();
 sg13g2_fill_2 FILLER_47_621 ();
 sg13g2_decap_4 FILLER_47_674 ();
 sg13g2_decap_4 FILLER_47_715 ();
 sg13g2_fill_1 FILLER_47_719 ();
 sg13g2_fill_1 FILLER_47_729 ();
 sg13g2_fill_2 FILLER_47_743 ();
 sg13g2_decap_8 FILLER_47_753 ();
 sg13g2_decap_8 FILLER_47_760 ();
 sg13g2_fill_1 FILLER_47_767 ();
 sg13g2_fill_1 FILLER_47_776 ();
 sg13g2_fill_2 FILLER_47_781 ();
 sg13g2_fill_1 FILLER_47_783 ();
 sg13g2_decap_4 FILLER_47_792 ();
 sg13g2_decap_8 FILLER_47_812 ();
 sg13g2_decap_4 FILLER_47_819 ();
 sg13g2_decap_8 FILLER_47_832 ();
 sg13g2_decap_4 FILLER_47_839 ();
 sg13g2_decap_4 FILLER_47_860 ();
 sg13g2_fill_1 FILLER_47_864 ();
 sg13g2_decap_8 FILLER_47_869 ();
 sg13g2_fill_2 FILLER_47_876 ();
 sg13g2_fill_2 FILLER_48_0 ();
 sg13g2_fill_1 FILLER_48_29 ();
 sg13g2_fill_2 FILLER_48_38 ();
 sg13g2_fill_1 FILLER_48_40 ();
 sg13g2_fill_1 FILLER_48_49 ();
 sg13g2_fill_2 FILLER_48_60 ();
 sg13g2_decap_8 FILLER_48_70 ();
 sg13g2_decap_8 FILLER_48_77 ();
 sg13g2_decap_4 FILLER_48_84 ();
 sg13g2_fill_1 FILLER_48_96 ();
 sg13g2_fill_1 FILLER_48_102 ();
 sg13g2_fill_1 FILLER_48_107 ();
 sg13g2_fill_2 FILLER_48_113 ();
 sg13g2_fill_1 FILLER_48_126 ();
 sg13g2_fill_1 FILLER_48_136 ();
 sg13g2_decap_4 FILLER_48_145 ();
 sg13g2_decap_4 FILLER_48_162 ();
 sg13g2_fill_1 FILLER_48_166 ();
 sg13g2_fill_2 FILLER_48_171 ();
 sg13g2_fill_1 FILLER_48_181 ();
 sg13g2_fill_2 FILLER_48_187 ();
 sg13g2_decap_8 FILLER_48_197 ();
 sg13g2_fill_1 FILLER_48_204 ();
 sg13g2_decap_8 FILLER_48_242 ();
 sg13g2_fill_2 FILLER_48_249 ();
 sg13g2_decap_8 FILLER_48_256 ();
 sg13g2_fill_1 FILLER_48_263 ();
 sg13g2_fill_1 FILLER_48_277 ();
 sg13g2_fill_2 FILLER_48_283 ();
 sg13g2_fill_2 FILLER_48_290 ();
 sg13g2_fill_1 FILLER_48_292 ();
 sg13g2_decap_8 FILLER_48_301 ();
 sg13g2_fill_1 FILLER_48_308 ();
 sg13g2_fill_1 FILLER_48_355 ();
 sg13g2_fill_1 FILLER_48_360 ();
 sg13g2_decap_4 FILLER_48_374 ();
 sg13g2_fill_2 FILLER_48_378 ();
 sg13g2_decap_8 FILLER_48_396 ();
 sg13g2_decap_8 FILLER_48_403 ();
 sg13g2_decap_8 FILLER_48_410 ();
 sg13g2_fill_2 FILLER_48_417 ();
 sg13g2_fill_1 FILLER_48_419 ();
 sg13g2_fill_2 FILLER_48_433 ();
 sg13g2_fill_1 FILLER_48_457 ();
 sg13g2_fill_1 FILLER_48_462 ();
 sg13g2_fill_2 FILLER_48_476 ();
 sg13g2_fill_1 FILLER_48_496 ();
 sg13g2_fill_1 FILLER_48_505 ();
 sg13g2_fill_1 FILLER_48_523 ();
 sg13g2_fill_1 FILLER_48_539 ();
 sg13g2_fill_2 FILLER_48_545 ();
 sg13g2_decap_8 FILLER_48_555 ();
 sg13g2_fill_2 FILLER_48_562 ();
 sg13g2_fill_1 FILLER_48_564 ();
 sg13g2_fill_2 FILLER_48_576 ();
 sg13g2_fill_1 FILLER_48_578 ();
 sg13g2_fill_2 FILLER_48_584 ();
 sg13g2_fill_1 FILLER_48_586 ();
 sg13g2_fill_1 FILLER_48_592 ();
 sg13g2_fill_1 FILLER_48_607 ();
 sg13g2_fill_2 FILLER_48_613 ();
 sg13g2_decap_4 FILLER_48_620 ();
 sg13g2_fill_2 FILLER_48_628 ();
 sg13g2_fill_1 FILLER_48_630 ();
 sg13g2_decap_4 FILLER_48_670 ();
 sg13g2_fill_2 FILLER_48_674 ();
 sg13g2_decap_8 FILLER_48_722 ();
 sg13g2_fill_2 FILLER_48_745 ();
 sg13g2_fill_1 FILLER_48_800 ();
 sg13g2_decap_4 FILLER_48_814 ();
 sg13g2_fill_1 FILLER_48_818 ();
 sg13g2_decap_8 FILLER_48_832 ();
 sg13g2_decap_8 FILLER_48_839 ();
 sg13g2_fill_2 FILLER_48_851 ();
 sg13g2_decap_8 FILLER_48_868 ();
 sg13g2_fill_2 FILLER_48_875 ();
 sg13g2_fill_1 FILLER_48_877 ();
 sg13g2_decap_4 FILLER_49_0 ();
 sg13g2_fill_1 FILLER_49_4 ();
 sg13g2_decap_8 FILLER_49_15 ();
 sg13g2_decap_8 FILLER_49_22 ();
 sg13g2_fill_2 FILLER_49_29 ();
 sg13g2_fill_1 FILLER_49_31 ();
 sg13g2_decap_4 FILLER_49_40 ();
 sg13g2_decap_8 FILLER_49_52 ();
 sg13g2_decap_8 FILLER_49_59 ();
 sg13g2_decap_8 FILLER_49_66 ();
 sg13g2_decap_8 FILLER_49_77 ();
 sg13g2_decap_8 FILLER_49_84 ();
 sg13g2_fill_2 FILLER_49_91 ();
 sg13g2_fill_2 FILLER_49_99 ();
 sg13g2_fill_1 FILLER_49_101 ();
 sg13g2_fill_1 FILLER_49_106 ();
 sg13g2_fill_1 FILLER_49_117 ();
 sg13g2_fill_2 FILLER_49_123 ();
 sg13g2_fill_2 FILLER_49_135 ();
 sg13g2_fill_1 FILLER_49_141 ();
 sg13g2_fill_2 FILLER_49_147 ();
 sg13g2_fill_2 FILLER_49_157 ();
 sg13g2_fill_1 FILLER_49_159 ();
 sg13g2_fill_1 FILLER_49_168 ();
 sg13g2_fill_1 FILLER_49_174 ();
 sg13g2_fill_1 FILLER_49_183 ();
 sg13g2_decap_8 FILLER_49_189 ();
 sg13g2_decap_8 FILLER_49_196 ();
 sg13g2_decap_4 FILLER_49_203 ();
 sg13g2_decap_8 FILLER_49_219 ();
 sg13g2_fill_1 FILLER_49_226 ();
 sg13g2_fill_2 FILLER_49_235 ();
 sg13g2_decap_8 FILLER_49_249 ();
 sg13g2_decap_8 FILLER_49_256 ();
 sg13g2_fill_2 FILLER_49_263 ();
 sg13g2_decap_8 FILLER_49_288 ();
 sg13g2_fill_2 FILLER_49_308 ();
 sg13g2_fill_1 FILLER_49_310 ();
 sg13g2_fill_1 FILLER_49_337 ();
 sg13g2_fill_2 FILLER_49_351 ();
 sg13g2_fill_2 FILLER_49_357 ();
 sg13g2_fill_1 FILLER_49_368 ();
 sg13g2_fill_2 FILLER_49_374 ();
 sg13g2_fill_1 FILLER_49_384 ();
 sg13g2_decap_4 FILLER_49_393 ();
 sg13g2_fill_1 FILLER_49_397 ();
 sg13g2_fill_2 FILLER_49_424 ();
 sg13g2_fill_2 FILLER_49_431 ();
 sg13g2_decap_8 FILLER_49_441 ();
 sg13g2_fill_1 FILLER_49_452 ();
 sg13g2_decap_4 FILLER_49_466 ();
 sg13g2_fill_1 FILLER_49_470 ();
 sg13g2_decap_4 FILLER_49_479 ();
 sg13g2_fill_1 FILLER_49_483 ();
 sg13g2_fill_2 FILLER_49_488 ();
 sg13g2_fill_1 FILLER_49_490 ();
 sg13g2_fill_2 FILLER_49_499 ();
 sg13g2_fill_2 FILLER_49_506 ();
 sg13g2_fill_1 FILLER_49_508 ();
 sg13g2_fill_1 FILLER_49_517 ();
 sg13g2_fill_2 FILLER_49_522 ();
 sg13g2_fill_1 FILLER_49_524 ();
 sg13g2_fill_2 FILLER_49_547 ();
 sg13g2_decap_4 FILLER_49_557 ();
 sg13g2_decap_4 FILLER_49_569 ();
 sg13g2_fill_1 FILLER_49_595 ();
 sg13g2_fill_2 FILLER_49_604 ();
 sg13g2_fill_2 FILLER_49_614 ();
 sg13g2_fill_1 FILLER_49_616 ();
 sg13g2_decap_8 FILLER_49_662 ();
 sg13g2_decap_8 FILLER_49_669 ();
 sg13g2_decap_8 FILLER_49_676 ();
 sg13g2_fill_2 FILLER_49_683 ();
 sg13g2_fill_1 FILLER_49_685 ();
 sg13g2_decap_4 FILLER_49_706 ();
 sg13g2_fill_2 FILLER_49_710 ();
 sg13g2_decap_4 FILLER_49_749 ();
 sg13g2_fill_2 FILLER_49_757 ();
 sg13g2_fill_1 FILLER_49_759 ();
 sg13g2_fill_2 FILLER_49_764 ();
 sg13g2_fill_1 FILLER_49_766 ();
 sg13g2_decap_8 FILLER_49_779 ();
 sg13g2_fill_2 FILLER_49_803 ();
 sg13g2_fill_1 FILLER_49_805 ();
 sg13g2_fill_2 FILLER_49_810 ();
 sg13g2_decap_4 FILLER_49_835 ();
 sg13g2_fill_1 FILLER_49_839 ();
 sg13g2_fill_1 FILLER_49_844 ();
 sg13g2_decap_4 FILLER_49_872 ();
 sg13g2_fill_2 FILLER_49_876 ();
 sg13g2_decap_8 FILLER_50_0 ();
 sg13g2_fill_1 FILLER_50_7 ();
 sg13g2_decap_4 FILLER_50_13 ();
 sg13g2_fill_2 FILLER_50_30 ();
 sg13g2_fill_1 FILLER_50_74 ();
 sg13g2_decap_8 FILLER_50_80 ();
 sg13g2_decap_4 FILLER_50_87 ();
 sg13g2_decap_8 FILLER_50_95 ();
 sg13g2_fill_1 FILLER_50_106 ();
 sg13g2_fill_1 FILLER_50_117 ();
 sg13g2_fill_1 FILLER_50_130 ();
 sg13g2_fill_1 FILLER_50_135 ();
 sg13g2_fill_1 FILLER_50_160 ();
 sg13g2_fill_1 FILLER_50_179 ();
 sg13g2_fill_2 FILLER_50_187 ();
 sg13g2_fill_2 FILLER_50_193 ();
 sg13g2_fill_2 FILLER_50_199 ();
 sg13g2_fill_2 FILLER_50_205 ();
 sg13g2_fill_1 FILLER_50_207 ();
 sg13g2_fill_2 FILLER_50_213 ();
 sg13g2_fill_1 FILLER_50_215 ();
 sg13g2_fill_2 FILLER_50_220 ();
 sg13g2_fill_1 FILLER_50_230 ();
 sg13g2_fill_1 FILLER_50_236 ();
 sg13g2_fill_2 FILLER_50_253 ();
 sg13g2_fill_1 FILLER_50_255 ();
 sg13g2_decap_8 FILLER_50_260 ();
 sg13g2_fill_1 FILLER_50_267 ();
 sg13g2_fill_1 FILLER_50_273 ();
 sg13g2_fill_1 FILLER_50_278 ();
 sg13g2_fill_1 FILLER_50_306 ();
 sg13g2_fill_1 FILLER_50_311 ();
 sg13g2_fill_2 FILLER_50_330 ();
 sg13g2_fill_1 FILLER_50_332 ();
 sg13g2_fill_1 FILLER_50_338 ();
 sg13g2_fill_1 FILLER_50_349 ();
 sg13g2_fill_2 FILLER_50_386 ();
 sg13g2_fill_2 FILLER_50_421 ();
 sg13g2_fill_1 FILLER_50_430 ();
 sg13g2_decap_8 FILLER_50_436 ();
 sg13g2_decap_8 FILLER_50_443 ();
 sg13g2_fill_2 FILLER_50_450 ();
 sg13g2_fill_1 FILLER_50_452 ();
 sg13g2_fill_2 FILLER_50_474 ();
 sg13g2_fill_1 FILLER_50_476 ();
 sg13g2_decap_8 FILLER_50_485 ();
 sg13g2_fill_2 FILLER_50_492 ();
 sg13g2_fill_2 FILLER_50_502 ();
 sg13g2_fill_1 FILLER_50_504 ();
 sg13g2_fill_1 FILLER_50_509 ();
 sg13g2_fill_1 FILLER_50_530 ();
 sg13g2_decap_8 FILLER_50_549 ();
 sg13g2_decap_4 FILLER_50_556 ();
 sg13g2_fill_1 FILLER_50_572 ();
 sg13g2_fill_1 FILLER_50_581 ();
 sg13g2_fill_2 FILLER_50_586 ();
 sg13g2_fill_1 FILLER_50_592 ();
 sg13g2_fill_1 FILLER_50_598 ();
 sg13g2_decap_8 FILLER_50_604 ();
 sg13g2_decap_8 FILLER_50_611 ();
 sg13g2_decap_4 FILLER_50_618 ();
 sg13g2_fill_2 FILLER_50_622 ();
 sg13g2_fill_1 FILLER_50_659 ();
 sg13g2_fill_2 FILLER_50_664 ();
 sg13g2_fill_2 FILLER_50_670 ();
 sg13g2_decap_8 FILLER_50_680 ();
 sg13g2_decap_8 FILLER_50_687 ();
 sg13g2_decap_8 FILLER_50_694 ();
 sg13g2_decap_4 FILLER_50_701 ();
 sg13g2_fill_2 FILLER_50_713 ();
 sg13g2_decap_4 FILLER_50_719 ();
 sg13g2_decap_8 FILLER_50_736 ();
 sg13g2_fill_1 FILLER_50_743 ();
 sg13g2_fill_1 FILLER_50_747 ();
 sg13g2_decap_8 FILLER_50_752 ();
 sg13g2_decap_8 FILLER_50_759 ();
 sg13g2_fill_1 FILLER_50_773 ();
 sg13g2_decap_8 FILLER_50_782 ();
 sg13g2_fill_2 FILLER_50_789 ();
 sg13g2_fill_1 FILLER_50_791 ();
 sg13g2_decap_8 FILLER_50_810 ();
 sg13g2_fill_1 FILLER_50_817 ();
 sg13g2_decap_8 FILLER_50_826 ();
 sg13g2_decap_4 FILLER_50_833 ();
 sg13g2_fill_2 FILLER_50_837 ();
 sg13g2_fill_2 FILLER_50_859 ();
 sg13g2_decap_8 FILLER_50_866 ();
 sg13g2_decap_4 FILLER_50_873 ();
 sg13g2_fill_1 FILLER_50_877 ();
 sg13g2_decap_4 FILLER_51_0 ();
 sg13g2_fill_2 FILLER_51_4 ();
 sg13g2_fill_2 FILLER_51_16 ();
 sg13g2_fill_1 FILLER_51_18 ();
 sg13g2_decap_8 FILLER_51_27 ();
 sg13g2_fill_1 FILLER_51_34 ();
 sg13g2_decap_4 FILLER_51_60 ();
 sg13g2_fill_2 FILLER_51_64 ();
 sg13g2_fill_2 FILLER_51_78 ();
 sg13g2_fill_1 FILLER_51_80 ();
 sg13g2_fill_1 FILLER_51_95 ();
 sg13g2_decap_4 FILLER_51_113 ();
 sg13g2_fill_2 FILLER_51_117 ();
 sg13g2_fill_1 FILLER_51_123 ();
 sg13g2_fill_1 FILLER_51_131 ();
 sg13g2_fill_1 FILLER_51_140 ();
 sg13g2_fill_1 FILLER_51_149 ();
 sg13g2_decap_8 FILLER_51_154 ();
 sg13g2_decap_8 FILLER_51_170 ();
 sg13g2_fill_2 FILLER_51_177 ();
 sg13g2_fill_1 FILLER_51_179 ();
 sg13g2_fill_1 FILLER_51_189 ();
 sg13g2_fill_2 FILLER_51_205 ();
 sg13g2_fill_1 FILLER_51_223 ();
 sg13g2_fill_1 FILLER_51_245 ();
 sg13g2_decap_4 FILLER_51_266 ();
 sg13g2_fill_2 FILLER_51_270 ();
 sg13g2_fill_1 FILLER_51_280 ();
 sg13g2_fill_1 FILLER_51_313 ();
 sg13g2_fill_2 FILLER_51_329 ();
 sg13g2_fill_1 FILLER_51_345 ();
 sg13g2_fill_2 FILLER_51_350 ();
 sg13g2_fill_2 FILLER_51_374 ();
 sg13g2_fill_2 FILLER_51_384 ();
 sg13g2_decap_4 FILLER_51_398 ();
 sg13g2_fill_1 FILLER_51_402 ();
 sg13g2_fill_1 FILLER_51_431 ();
 sg13g2_fill_2 FILLER_51_437 ();
 sg13g2_decap_4 FILLER_51_451 ();
 sg13g2_fill_2 FILLER_51_463 ();
 sg13g2_fill_1 FILLER_51_470 ();
 sg13g2_decap_4 FILLER_51_504 ();
 sg13g2_decap_4 FILLER_51_516 ();
 sg13g2_fill_2 FILLER_51_520 ();
 sg13g2_fill_2 FILLER_51_550 ();
 sg13g2_fill_1 FILLER_51_560 ();
 sg13g2_decap_8 FILLER_51_570 ();
 sg13g2_decap_8 FILLER_51_577 ();
 sg13g2_fill_1 FILLER_51_605 ();
 sg13g2_fill_2 FILLER_51_611 ();
 sg13g2_fill_1 FILLER_51_622 ();
 sg13g2_decap_8 FILLER_51_632 ();
 sg13g2_fill_2 FILLER_51_639 ();
 sg13g2_fill_1 FILLER_51_641 ();
 sg13g2_decap_8 FILLER_51_655 ();
 sg13g2_fill_2 FILLER_51_662 ();
 sg13g2_fill_1 FILLER_51_664 ();
 sg13g2_decap_8 FILLER_51_682 ();
 sg13g2_decap_8 FILLER_51_689 ();
 sg13g2_decap_4 FILLER_51_696 ();
 sg13g2_fill_2 FILLER_51_711 ();
 sg13g2_fill_1 FILLER_51_713 ();
 sg13g2_decap_8 FILLER_51_730 ();
 sg13g2_fill_1 FILLER_51_737 ();
 sg13g2_decap_4 FILLER_51_760 ();
 sg13g2_fill_2 FILLER_51_764 ();
 sg13g2_fill_1 FILLER_51_792 ();
 sg13g2_fill_1 FILLER_51_800 ();
 sg13g2_fill_2 FILLER_51_814 ();
 sg13g2_decap_4 FILLER_51_820 ();
 sg13g2_fill_1 FILLER_51_828 ();
 sg13g2_fill_2 FILLER_51_858 ();
 sg13g2_decap_8 FILLER_51_870 ();
 sg13g2_fill_1 FILLER_51_877 ();
 sg13g2_fill_2 FILLER_52_0 ();
 sg13g2_fill_1 FILLER_52_2 ();
 sg13g2_fill_1 FILLER_52_13 ();
 sg13g2_decap_8 FILLER_52_42 ();
 sg13g2_decap_8 FILLER_52_49 ();
 sg13g2_fill_2 FILLER_52_56 ();
 sg13g2_fill_1 FILLER_52_66 ();
 sg13g2_fill_2 FILLER_52_75 ();
 sg13g2_fill_1 FILLER_52_77 ();
 sg13g2_fill_1 FILLER_52_99 ();
 sg13g2_fill_2 FILLER_52_112 ();
 sg13g2_fill_1 FILLER_52_114 ();
 sg13g2_fill_1 FILLER_52_119 ();
 sg13g2_fill_1 FILLER_52_130 ();
 sg13g2_fill_2 FILLER_52_135 ();
 sg13g2_fill_2 FILLER_52_154 ();
 sg13g2_fill_1 FILLER_52_156 ();
 sg13g2_fill_2 FILLER_52_175 ();
 sg13g2_fill_1 FILLER_52_177 ();
 sg13g2_fill_1 FILLER_52_183 ();
 sg13g2_decap_8 FILLER_52_217 ();
 sg13g2_decap_4 FILLER_52_224 ();
 sg13g2_fill_1 FILLER_52_228 ();
 sg13g2_fill_1 FILLER_52_245 ();
 sg13g2_fill_2 FILLER_52_254 ();
 sg13g2_fill_2 FILLER_52_264 ();
 sg13g2_fill_2 FILLER_52_270 ();
 sg13g2_fill_1 FILLER_52_272 ();
 sg13g2_decap_4 FILLER_52_285 ();
 sg13g2_fill_1 FILLER_52_289 ();
 sg13g2_fill_1 FILLER_52_295 ();
 sg13g2_fill_2 FILLER_52_311 ();
 sg13g2_fill_1 FILLER_52_313 ();
 sg13g2_fill_2 FILLER_52_328 ();
 sg13g2_fill_1 FILLER_52_336 ();
 sg13g2_fill_2 FILLER_52_358 ();
 sg13g2_fill_1 FILLER_52_360 ();
 sg13g2_decap_8 FILLER_52_369 ();
 sg13g2_decap_8 FILLER_52_376 ();
 sg13g2_decap_8 FILLER_52_392 ();
 sg13g2_decap_8 FILLER_52_399 ();
 sg13g2_decap_4 FILLER_52_406 ();
 sg13g2_fill_1 FILLER_52_415 ();
 sg13g2_fill_2 FILLER_52_429 ();
 sg13g2_fill_1 FILLER_52_431 ();
 sg13g2_decap_8 FILLER_52_454 ();
 sg13g2_fill_2 FILLER_52_461 ();
 sg13g2_fill_1 FILLER_52_463 ();
 sg13g2_fill_2 FILLER_52_471 ();
 sg13g2_fill_1 FILLER_52_478 ();
 sg13g2_fill_2 FILLER_52_501 ();
 sg13g2_fill_2 FILLER_52_519 ();
 sg13g2_fill_1 FILLER_52_521 ();
 sg13g2_fill_2 FILLER_52_527 ();
 sg13g2_fill_1 FILLER_52_529 ();
 sg13g2_decap_4 FILLER_52_538 ();
 sg13g2_fill_2 FILLER_52_542 ();
 sg13g2_fill_2 FILLER_52_552 ();
 sg13g2_fill_1 FILLER_52_554 ();
 sg13g2_decap_8 FILLER_52_567 ();
 sg13g2_decap_4 FILLER_52_574 ();
 sg13g2_fill_1 FILLER_52_578 ();
 sg13g2_fill_1 FILLER_52_595 ();
 sg13g2_decap_4 FILLER_52_601 ();
 sg13g2_fill_1 FILLER_52_632 ();
 sg13g2_fill_1 FILLER_52_645 ();
 sg13g2_decap_8 FILLER_52_656 ();
 sg13g2_fill_1 FILLER_52_675 ();
 sg13g2_decap_4 FILLER_52_686 ();
 sg13g2_fill_2 FILLER_52_715 ();
 sg13g2_fill_1 FILLER_52_717 ();
 sg13g2_decap_4 FILLER_52_722 ();
 sg13g2_fill_2 FILLER_52_731 ();
 sg13g2_fill_1 FILLER_52_733 ();
 sg13g2_decap_4 FILLER_52_759 ();
 sg13g2_fill_1 FILLER_52_772 ();
 sg13g2_fill_2 FILLER_52_809 ();
 sg13g2_decap_8 FILLER_52_819 ();
 sg13g2_decap_8 FILLER_52_826 ();
 sg13g2_fill_2 FILLER_52_845 ();
 sg13g2_fill_1 FILLER_52_851 ();
 sg13g2_decap_4 FILLER_52_872 ();
 sg13g2_fill_2 FILLER_52_876 ();
 sg13g2_fill_1 FILLER_53_0 ();
 sg13g2_fill_1 FILLER_53_15 ();
 sg13g2_fill_1 FILLER_53_20 ();
 sg13g2_fill_2 FILLER_53_57 ();
 sg13g2_fill_2 FILLER_53_76 ();
 sg13g2_fill_1 FILLER_53_78 ();
 sg13g2_fill_1 FILLER_53_87 ();
 sg13g2_fill_2 FILLER_53_92 ();
 sg13g2_decap_4 FILLER_53_111 ();
 sg13g2_fill_1 FILLER_53_115 ();
 sg13g2_decap_4 FILLER_53_128 ();
 sg13g2_fill_1 FILLER_53_140 ();
 sg13g2_fill_2 FILLER_53_146 ();
 sg13g2_decap_8 FILLER_53_153 ();
 sg13g2_fill_1 FILLER_53_172 ();
 sg13g2_fill_2 FILLER_53_177 ();
 sg13g2_fill_1 FILLER_53_179 ();
 sg13g2_decap_4 FILLER_53_185 ();
 sg13g2_fill_2 FILLER_53_189 ();
 sg13g2_decap_8 FILLER_53_200 ();
 sg13g2_decap_8 FILLER_53_207 ();
 sg13g2_fill_2 FILLER_53_214 ();
 sg13g2_decap_4 FILLER_53_233 ();
 sg13g2_fill_1 FILLER_53_237 ();
 sg13g2_fill_2 FILLER_53_247 ();
 sg13g2_fill_2 FILLER_53_261 ();
 sg13g2_decap_4 FILLER_53_271 ();
 sg13g2_fill_2 FILLER_53_279 ();
 sg13g2_fill_1 FILLER_53_281 ();
 sg13g2_fill_2 FILLER_53_290 ();
 sg13g2_fill_1 FILLER_53_292 ();
 sg13g2_decap_8 FILLER_53_298 ();
 sg13g2_decap_8 FILLER_53_305 ();
 sg13g2_decap_8 FILLER_53_312 ();
 sg13g2_fill_2 FILLER_53_319 ();
 sg13g2_fill_1 FILLER_53_321 ();
 sg13g2_fill_1 FILLER_53_332 ();
 sg13g2_fill_2 FILLER_53_338 ();
 sg13g2_fill_2 FILLER_53_353 ();
 sg13g2_fill_2 FILLER_53_360 ();
 sg13g2_fill_1 FILLER_53_362 ();
 sg13g2_decap_4 FILLER_53_380 ();
 sg13g2_fill_2 FILLER_53_384 ();
 sg13g2_fill_2 FILLER_53_398 ();
 sg13g2_fill_1 FILLER_53_400 ();
 sg13g2_decap_8 FILLER_53_405 ();
 sg13g2_fill_2 FILLER_53_418 ();
 sg13g2_fill_2 FILLER_53_424 ();
 sg13g2_fill_1 FILLER_53_426 ();
 sg13g2_decap_4 FILLER_53_438 ();
 sg13g2_fill_2 FILLER_53_442 ();
 sg13g2_fill_1 FILLER_53_449 ();
 sg13g2_fill_2 FILLER_53_459 ();
 sg13g2_fill_1 FILLER_53_461 ();
 sg13g2_decap_8 FILLER_53_484 ();
 sg13g2_decap_4 FILLER_53_491 ();
 sg13g2_fill_1 FILLER_53_505 ();
 sg13g2_fill_2 FILLER_53_511 ();
 sg13g2_decap_4 FILLER_53_521 ();
 sg13g2_fill_1 FILLER_53_525 ();
 sg13g2_fill_2 FILLER_53_581 ();
 sg13g2_fill_2 FILLER_53_610 ();
 sg13g2_decap_8 FILLER_53_627 ();
 sg13g2_decap_4 FILLER_53_634 ();
 sg13g2_fill_1 FILLER_53_652 ();
 sg13g2_fill_2 FILLER_53_668 ();
 sg13g2_fill_1 FILLER_53_670 ();
 sg13g2_fill_2 FILLER_53_676 ();
 sg13g2_decap_4 FILLER_53_683 ();
 sg13g2_fill_1 FILLER_53_691 ();
 sg13g2_fill_1 FILLER_53_700 ();
 sg13g2_fill_1 FILLER_53_709 ();
 sg13g2_decap_4 FILLER_53_722 ();
 sg13g2_fill_2 FILLER_53_726 ();
 sg13g2_decap_8 FILLER_53_744 ();
 sg13g2_fill_2 FILLER_53_751 ();
 sg13g2_decap_8 FILLER_53_758 ();
 sg13g2_fill_1 FILLER_53_769 ();
 sg13g2_fill_2 FILLER_53_800 ();
 sg13g2_decap_8 FILLER_53_807 ();
 sg13g2_fill_2 FILLER_53_814 ();
 sg13g2_decap_4 FILLER_53_824 ();
 sg13g2_fill_1 FILLER_53_828 ();
 sg13g2_decap_8 FILLER_53_834 ();
 sg13g2_decap_8 FILLER_53_841 ();
 sg13g2_fill_2 FILLER_53_848 ();
 sg13g2_fill_1 FILLER_53_850 ();
 sg13g2_decap_8 FILLER_54_0 ();
 sg13g2_decap_8 FILLER_54_7 ();
 sg13g2_decap_8 FILLER_54_14 ();
 sg13g2_decap_4 FILLER_54_21 ();
 sg13g2_fill_1 FILLER_54_41 ();
 sg13g2_fill_2 FILLER_54_47 ();
 sg13g2_fill_1 FILLER_54_53 ();
 sg13g2_fill_1 FILLER_54_62 ();
 sg13g2_fill_2 FILLER_54_71 ();
 sg13g2_fill_1 FILLER_54_78 ();
 sg13g2_fill_2 FILLER_54_84 ();
 sg13g2_decap_8 FILLER_54_94 ();
 sg13g2_fill_2 FILLER_54_105 ();
 sg13g2_fill_1 FILLER_54_107 ();
 sg13g2_fill_2 FILLER_54_112 ();
 sg13g2_fill_1 FILLER_54_114 ();
 sg13g2_decap_8 FILLER_54_127 ();
 sg13g2_fill_2 FILLER_54_134 ();
 sg13g2_fill_2 FILLER_54_152 ();
 sg13g2_decap_8 FILLER_54_179 ();
 sg13g2_fill_2 FILLER_54_186 ();
 sg13g2_fill_1 FILLER_54_188 ();
 sg13g2_fill_2 FILLER_54_201 ();
 sg13g2_fill_2 FILLER_54_237 ();
 sg13g2_fill_1 FILLER_54_239 ();
 sg13g2_decap_8 FILLER_54_261 ();
 sg13g2_fill_2 FILLER_54_268 ();
 sg13g2_fill_1 FILLER_54_270 ();
 sg13g2_fill_2 FILLER_54_279 ();
 sg13g2_fill_2 FILLER_54_285 ();
 sg13g2_fill_1 FILLER_54_292 ();
 sg13g2_fill_2 FILLER_54_310 ();
 sg13g2_fill_1 FILLER_54_312 ();
 sg13g2_decap_8 FILLER_54_343 ();
 sg13g2_decap_8 FILLER_54_350 ();
 sg13g2_decap_8 FILLER_54_377 ();
 sg13g2_decap_8 FILLER_54_384 ();
 sg13g2_fill_2 FILLER_54_391 ();
 sg13g2_fill_1 FILLER_54_404 ();
 sg13g2_decap_8 FILLER_54_413 ();
 sg13g2_decap_8 FILLER_54_420 ();
 sg13g2_decap_4 FILLER_54_427 ();
 sg13g2_fill_2 FILLER_54_444 ();
 sg13g2_fill_1 FILLER_54_446 ();
 sg13g2_fill_2 FILLER_54_462 ();
 sg13g2_fill_1 FILLER_54_492 ();
 sg13g2_decap_8 FILLER_54_496 ();
 sg13g2_decap_8 FILLER_54_503 ();
 sg13g2_fill_2 FILLER_54_510 ();
 sg13g2_decap_4 FILLER_54_517 ();
 sg13g2_fill_2 FILLER_54_521 ();
 sg13g2_decap_8 FILLER_54_539 ();
 sg13g2_decap_4 FILLER_54_546 ();
 sg13g2_fill_1 FILLER_54_550 ();
 sg13g2_fill_2 FILLER_54_575 ();
 sg13g2_fill_1 FILLER_54_577 ();
 sg13g2_decap_8 FILLER_54_599 ();
 sg13g2_fill_2 FILLER_54_606 ();
 sg13g2_fill_1 FILLER_54_608 ();
 sg13g2_decap_8 FILLER_54_631 ();
 sg13g2_fill_1 FILLER_54_638 ();
 sg13g2_decap_8 FILLER_54_647 ();
 sg13g2_decap_4 FILLER_54_654 ();
 sg13g2_decap_8 FILLER_54_693 ();
 sg13g2_fill_2 FILLER_54_700 ();
 sg13g2_fill_1 FILLER_54_702 ();
 sg13g2_fill_2 FILLER_54_711 ();
 sg13g2_fill_1 FILLER_54_718 ();
 sg13g2_decap_4 FILLER_54_723 ();
 sg13g2_fill_2 FILLER_54_731 ();
 sg13g2_fill_1 FILLER_54_733 ();
 sg13g2_fill_2 FILLER_54_744 ();
 sg13g2_decap_8 FILLER_54_751 ();
 sg13g2_fill_2 FILLER_54_758 ();
 sg13g2_fill_1 FILLER_54_760 ();
 sg13g2_decap_4 FILLER_54_765 ();
 sg13g2_fill_1 FILLER_54_769 ();
 sg13g2_fill_1 FILLER_54_783 ();
 sg13g2_decap_4 FILLER_54_807 ();
 sg13g2_fill_1 FILLER_54_811 ();
 sg13g2_fill_2 FILLER_54_820 ();
 sg13g2_fill_1 FILLER_54_822 ();
 sg13g2_decap_4 FILLER_54_826 ();
 sg13g2_fill_1 FILLER_54_830 ();
 sg13g2_fill_2 FILLER_54_846 ();
 sg13g2_fill_1 FILLER_54_848 ();
 sg13g2_decap_8 FILLER_54_867 ();
 sg13g2_decap_4 FILLER_54_874 ();
 sg13g2_decap_8 FILLER_55_0 ();
 sg13g2_decap_8 FILLER_55_7 ();
 sg13g2_decap_8 FILLER_55_14 ();
 sg13g2_decap_8 FILLER_55_21 ();
 sg13g2_decap_8 FILLER_55_28 ();
 sg13g2_fill_2 FILLER_55_35 ();
 sg13g2_fill_2 FILLER_55_59 ();
 sg13g2_fill_1 FILLER_55_69 ();
 sg13g2_fill_1 FILLER_55_86 ();
 sg13g2_fill_2 FILLER_55_91 ();
 sg13g2_fill_1 FILLER_55_93 ();
 sg13g2_decap_8 FILLER_55_119 ();
 sg13g2_decap_4 FILLER_55_126 ();
 sg13g2_fill_1 FILLER_55_130 ();
 sg13g2_decap_4 FILLER_55_139 ();
 sg13g2_fill_2 FILLER_55_143 ();
 sg13g2_fill_1 FILLER_55_160 ();
 sg13g2_decap_4 FILLER_55_208 ();
 sg13g2_fill_1 FILLER_55_212 ();
 sg13g2_decap_8 FILLER_55_235 ();
 sg13g2_fill_1 FILLER_55_242 ();
 sg13g2_decap_4 FILLER_55_247 ();
 sg13g2_fill_1 FILLER_55_251 ();
 sg13g2_decap_8 FILLER_55_260 ();
 sg13g2_decap_8 FILLER_55_267 ();
 sg13g2_decap_4 FILLER_55_274 ();
 sg13g2_fill_2 FILLER_55_278 ();
 sg13g2_fill_2 FILLER_55_313 ();
 sg13g2_decap_4 FILLER_55_328 ();
 sg13g2_decap_4 FILLER_55_341 ();
 sg13g2_fill_1 FILLER_55_345 ();
 sg13g2_fill_1 FILLER_55_354 ();
 sg13g2_decap_8 FILLER_55_362 ();
 sg13g2_fill_1 FILLER_55_402 ();
 sg13g2_fill_2 FILLER_55_419 ();
 sg13g2_fill_1 FILLER_55_421 ();
 sg13g2_fill_1 FILLER_55_435 ();
 sg13g2_decap_4 FILLER_55_462 ();
 sg13g2_fill_1 FILLER_55_496 ();
 sg13g2_fill_1 FILLER_55_507 ();
 sg13g2_fill_2 FILLER_55_526 ();
 sg13g2_decap_8 FILLER_55_546 ();
 sg13g2_decap_4 FILLER_55_553 ();
 sg13g2_fill_2 FILLER_55_557 ();
 sg13g2_decap_8 FILLER_55_564 ();
 sg13g2_decap_8 FILLER_55_571 ();
 sg13g2_fill_2 FILLER_55_590 ();
 sg13g2_fill_1 FILLER_55_598 ();
 sg13g2_fill_2 FILLER_55_604 ();
 sg13g2_decap_8 FILLER_55_630 ();
 sg13g2_decap_4 FILLER_55_637 ();
 sg13g2_fill_1 FILLER_55_641 ();
 sg13g2_fill_2 FILLER_55_650 ();
 sg13g2_fill_1 FILLER_55_652 ();
 sg13g2_fill_2 FILLER_55_684 ();
 sg13g2_decap_4 FILLER_55_695 ();
 sg13g2_decap_4 FILLER_55_704 ();
 sg13g2_fill_2 FILLER_55_712 ();
 sg13g2_fill_1 FILLER_55_714 ();
 sg13g2_fill_1 FILLER_55_720 ();
 sg13g2_fill_1 FILLER_55_726 ();
 sg13g2_fill_1 FILLER_55_740 ();
 sg13g2_decap_8 FILLER_55_749 ();
 sg13g2_decap_8 FILLER_55_756 ();
 sg13g2_decap_8 FILLER_55_763 ();
 sg13g2_decap_4 FILLER_55_770 ();
 sg13g2_fill_1 FILLER_55_774 ();
 sg13g2_decap_8 FILLER_55_785 ();
 sg13g2_fill_2 FILLER_55_792 ();
 sg13g2_fill_1 FILLER_55_794 ();
 sg13g2_decap_8 FILLER_55_808 ();
 sg13g2_fill_2 FILLER_55_815 ();
 sg13g2_fill_2 FILLER_55_828 ();
 sg13g2_fill_2 FILLER_55_838 ();
 sg13g2_fill_2 FILLER_55_849 ();
 sg13g2_fill_1 FILLER_55_851 ();
 sg13g2_fill_2 FILLER_55_856 ();
 sg13g2_fill_2 FILLER_55_875 ();
 sg13g2_fill_1 FILLER_55_877 ();
 sg13g2_decap_8 FILLER_56_0 ();
 sg13g2_decap_8 FILLER_56_7 ();
 sg13g2_decap_8 FILLER_56_14 ();
 sg13g2_decap_8 FILLER_56_21 ();
 sg13g2_decap_8 FILLER_56_28 ();
 sg13g2_decap_8 FILLER_56_35 ();
 sg13g2_fill_1 FILLER_56_42 ();
 sg13g2_decap_4 FILLER_56_51 ();
 sg13g2_fill_2 FILLER_56_55 ();
 sg13g2_decap_4 FILLER_56_94 ();
 sg13g2_fill_2 FILLER_56_98 ();
 sg13g2_decap_4 FILLER_56_139 ();
 sg13g2_fill_2 FILLER_56_147 ();
 sg13g2_fill_1 FILLER_56_149 ();
 sg13g2_fill_2 FILLER_56_163 ();
 sg13g2_fill_1 FILLER_56_165 ();
 sg13g2_decap_4 FILLER_56_174 ();
 sg13g2_decap_4 FILLER_56_203 ();
 sg13g2_decap_8 FILLER_56_242 ();
 sg13g2_fill_2 FILLER_56_249 ();
 sg13g2_fill_1 FILLER_56_251 ();
 sg13g2_decap_4 FILLER_56_272 ();
 sg13g2_decap_4 FILLER_56_280 ();
 sg13g2_decap_8 FILLER_56_320 ();
 sg13g2_fill_1 FILLER_56_327 ();
 sg13g2_fill_1 FILLER_56_353 ();
 sg13g2_decap_4 FILLER_56_358 ();
 sg13g2_decap_8 FILLER_56_366 ();
 sg13g2_decap_8 FILLER_56_373 ();
 sg13g2_decap_8 FILLER_56_380 ();
 sg13g2_fill_2 FILLER_56_387 ();
 sg13g2_fill_1 FILLER_56_389 ();
 sg13g2_fill_2 FILLER_56_406 ();
 sg13g2_fill_2 FILLER_56_431 ();
 sg13g2_fill_1 FILLER_56_433 ();
 sg13g2_fill_2 FILLER_56_446 ();
 sg13g2_fill_2 FILLER_56_453 ();
 sg13g2_decap_8 FILLER_56_460 ();
 sg13g2_decap_4 FILLER_56_467 ();
 sg13g2_fill_1 FILLER_56_471 ();
 sg13g2_fill_1 FILLER_56_480 ();
 sg13g2_fill_1 FILLER_56_493 ();
 sg13g2_fill_1 FILLER_56_516 ();
 sg13g2_fill_2 FILLER_56_526 ();
 sg13g2_decap_8 FILLER_56_532 ();
 sg13g2_fill_2 FILLER_56_539 ();
 sg13g2_fill_1 FILLER_56_541 ();
 sg13g2_fill_2 FILLER_56_553 ();
 sg13g2_fill_1 FILLER_56_555 ();
 sg13g2_decap_8 FILLER_56_561 ();
 sg13g2_decap_4 FILLER_56_568 ();
 sg13g2_fill_1 FILLER_56_572 ();
 sg13g2_decap_4 FILLER_56_578 ();
 sg13g2_fill_2 FILLER_56_582 ();
 sg13g2_fill_2 FILLER_56_599 ();
 sg13g2_fill_1 FILLER_56_601 ();
 sg13g2_decap_4 FILLER_56_614 ();
 sg13g2_fill_1 FILLER_56_618 ();
 sg13g2_fill_2 FILLER_56_648 ();
 sg13g2_fill_1 FILLER_56_650 ();
 sg13g2_fill_2 FILLER_56_658 ();
 sg13g2_fill_2 FILLER_56_676 ();
 sg13g2_fill_1 FILLER_56_678 ();
 sg13g2_fill_1 FILLER_56_708 ();
 sg13g2_decap_4 FILLER_56_714 ();
 sg13g2_fill_2 FILLER_56_718 ();
 sg13g2_fill_2 FILLER_56_725 ();
 sg13g2_fill_1 FILLER_56_735 ();
 sg13g2_decap_4 FILLER_56_746 ();
 sg13g2_fill_2 FILLER_56_759 ();
 sg13g2_fill_2 FILLER_56_782 ();
 sg13g2_fill_1 FILLER_56_784 ();
 sg13g2_decap_4 FILLER_56_798 ();
 sg13g2_fill_2 FILLER_56_802 ();
 sg13g2_decap_8 FILLER_56_825 ();
 sg13g2_decap_8 FILLER_56_832 ();
 sg13g2_decap_8 FILLER_56_839 ();
 sg13g2_decap_4 FILLER_56_846 ();
 sg13g2_fill_1 FILLER_56_854 ();
 sg13g2_fill_2 FILLER_56_867 ();
 sg13g2_decap_4 FILLER_56_874 ();
 sg13g2_decap_8 FILLER_57_0 ();
 sg13g2_decap_8 FILLER_57_7 ();
 sg13g2_decap_8 FILLER_57_14 ();
 sg13g2_decap_8 FILLER_57_21 ();
 sg13g2_decap_8 FILLER_57_28 ();
 sg13g2_decap_8 FILLER_57_35 ();
 sg13g2_decap_8 FILLER_57_42 ();
 sg13g2_fill_2 FILLER_57_57 ();
 sg13g2_fill_2 FILLER_57_92 ();
 sg13g2_fill_1 FILLER_57_99 ();
 sg13g2_fill_2 FILLER_57_104 ();
 sg13g2_fill_1 FILLER_57_110 ();
 sg13g2_fill_2 FILLER_57_114 ();
 sg13g2_decap_8 FILLER_57_128 ();
 sg13g2_fill_1 FILLER_57_135 ();
 sg13g2_fill_1 FILLER_57_144 ();
 sg13g2_fill_1 FILLER_57_172 ();
 sg13g2_fill_1 FILLER_57_181 ();
 sg13g2_decap_4 FILLER_57_190 ();
 sg13g2_fill_1 FILLER_57_194 ();
 sg13g2_fill_1 FILLER_57_198 ();
 sg13g2_fill_2 FILLER_57_203 ();
 sg13g2_decap_8 FILLER_57_209 ();
 sg13g2_decap_4 FILLER_57_216 ();
 sg13g2_fill_2 FILLER_57_220 ();
 sg13g2_fill_2 FILLER_57_230 ();
 sg13g2_fill_1 FILLER_57_232 ();
 sg13g2_decap_8 FILLER_57_238 ();
 sg13g2_decap_4 FILLER_57_245 ();
 sg13g2_fill_2 FILLER_57_267 ();
 sg13g2_fill_1 FILLER_57_269 ();
 sg13g2_fill_1 FILLER_57_275 ();
 sg13g2_fill_1 FILLER_57_300 ();
 sg13g2_decap_8 FILLER_57_305 ();
 sg13g2_fill_1 FILLER_57_312 ();
 sg13g2_decap_8 FILLER_57_318 ();
 sg13g2_decap_8 FILLER_57_325 ();
 sg13g2_fill_2 FILLER_57_335 ();
 sg13g2_fill_1 FILLER_57_337 ();
 sg13g2_fill_1 FILLER_57_343 ();
 sg13g2_fill_1 FILLER_57_362 ();
 sg13g2_fill_2 FILLER_57_368 ();
 sg13g2_decap_8 FILLER_57_374 ();
 sg13g2_fill_2 FILLER_57_381 ();
 sg13g2_decap_4 FILLER_57_400 ();
 sg13g2_fill_2 FILLER_57_404 ();
 sg13g2_fill_2 FILLER_57_411 ();
 sg13g2_fill_1 FILLER_57_421 ();
 sg13g2_decap_8 FILLER_57_430 ();
 sg13g2_fill_1 FILLER_57_437 ();
 sg13g2_fill_2 FILLER_57_442 ();
 sg13g2_fill_1 FILLER_57_444 ();
 sg13g2_decap_4 FILLER_57_455 ();
 sg13g2_fill_1 FILLER_57_459 ();
 sg13g2_decap_8 FILLER_57_464 ();
 sg13g2_fill_1 FILLER_57_471 ();
 sg13g2_decap_4 FILLER_57_477 ();
 sg13g2_fill_2 FILLER_57_505 ();
 sg13g2_fill_1 FILLER_57_514 ();
 sg13g2_fill_2 FILLER_57_526 ();
 sg13g2_fill_1 FILLER_57_528 ();
 sg13g2_fill_2 FILLER_57_538 ();
 sg13g2_decap_4 FILLER_57_584 ();
 sg13g2_decap_4 FILLER_57_593 ();
 sg13g2_fill_1 FILLER_57_597 ();
 sg13g2_fill_1 FILLER_57_608 ();
 sg13g2_fill_1 FILLER_57_633 ();
 sg13g2_decap_8 FILLER_57_638 ();
 sg13g2_decap_8 FILLER_57_645 ();
 sg13g2_decap_4 FILLER_57_652 ();
 sg13g2_fill_1 FILLER_57_656 ();
 sg13g2_fill_1 FILLER_57_668 ();
 sg13g2_fill_2 FILLER_57_674 ();
 sg13g2_decap_8 FILLER_57_693 ();
 sg13g2_decap_4 FILLER_57_706 ();
 sg13g2_fill_1 FILLER_57_749 ();
 sg13g2_fill_1 FILLER_57_754 ();
 sg13g2_fill_2 FILLER_57_760 ();
 sg13g2_fill_1 FILLER_57_766 ();
 sg13g2_fill_2 FILLER_57_777 ();
 sg13g2_fill_1 FILLER_57_787 ();
 sg13g2_fill_1 FILLER_57_799 ();
 sg13g2_fill_2 FILLER_57_805 ();
 sg13g2_fill_2 FILLER_57_812 ();
 sg13g2_fill_2 FILLER_57_818 ();
 sg13g2_fill_1 FILLER_57_820 ();
 sg13g2_fill_2 FILLER_57_837 ();
 sg13g2_fill_1 FILLER_57_847 ();
 sg13g2_decap_4 FILLER_57_874 ();
 sg13g2_decap_8 FILLER_58_0 ();
 sg13g2_decap_8 FILLER_58_7 ();
 sg13g2_decap_8 FILLER_58_14 ();
 sg13g2_decap_8 FILLER_58_21 ();
 sg13g2_decap_8 FILLER_58_28 ();
 sg13g2_decap_8 FILLER_58_35 ();
 sg13g2_decap_4 FILLER_58_42 ();
 sg13g2_fill_2 FILLER_58_46 ();
 sg13g2_fill_2 FILLER_58_52 ();
 sg13g2_fill_1 FILLER_58_54 ();
 sg13g2_fill_2 FILLER_58_81 ();
 sg13g2_fill_2 FILLER_58_87 ();
 sg13g2_fill_2 FILLER_58_104 ();
 sg13g2_fill_2 FILLER_58_111 ();
 sg13g2_fill_2 FILLER_58_117 ();
 sg13g2_fill_1 FILLER_58_119 ();
 sg13g2_decap_8 FILLER_58_128 ();
 sg13g2_decap_8 FILLER_58_135 ();
 sg13g2_decap_8 FILLER_58_142 ();
 sg13g2_decap_8 FILLER_58_149 ();
 sg13g2_decap_4 FILLER_58_156 ();
 sg13g2_fill_1 FILLER_58_160 ();
 sg13g2_decap_8 FILLER_58_169 ();
 sg13g2_decap_8 FILLER_58_176 ();
 sg13g2_decap_8 FILLER_58_183 ();
 sg13g2_fill_1 FILLER_58_190 ();
 sg13g2_fill_1 FILLER_58_215 ();
 sg13g2_fill_1 FILLER_58_232 ();
 sg13g2_fill_2 FILLER_58_251 ();
 sg13g2_fill_2 FILLER_58_258 ();
 sg13g2_fill_1 FILLER_58_326 ();
 sg13g2_decap_4 FILLER_58_363 ();
 sg13g2_decap_4 FILLER_58_391 ();
 sg13g2_fill_1 FILLER_58_395 ();
 sg13g2_fill_2 FILLER_58_399 ();
 sg13g2_decap_4 FILLER_58_414 ();
 sg13g2_fill_1 FILLER_58_434 ();
 sg13g2_fill_1 FILLER_58_448 ();
 sg13g2_fill_2 FILLER_58_458 ();
 sg13g2_fill_1 FILLER_58_468 ();
 sg13g2_decap_8 FILLER_58_473 ();
 sg13g2_fill_2 FILLER_58_480 ();
 sg13g2_fill_1 FILLER_58_496 ();
 sg13g2_decap_4 FILLER_58_502 ();
 sg13g2_fill_1 FILLER_58_513 ();
 sg13g2_fill_1 FILLER_58_518 ();
 sg13g2_fill_1 FILLER_58_526 ();
 sg13g2_fill_1 FILLER_58_563 ();
 sg13g2_fill_1 FILLER_58_569 ();
 sg13g2_fill_2 FILLER_58_598 ();
 sg13g2_fill_1 FILLER_58_600 ();
 sg13g2_fill_1 FILLER_58_623 ();
 sg13g2_decap_8 FILLER_58_641 ();
 sg13g2_decap_4 FILLER_58_648 ();
 sg13g2_fill_1 FILLER_58_652 ();
 sg13g2_decap_8 FILLER_58_657 ();
 sg13g2_decap_4 FILLER_58_664 ();
 sg13g2_fill_1 FILLER_58_668 ();
 sg13g2_decap_8 FILLER_58_678 ();
 sg13g2_fill_1 FILLER_58_685 ();
 sg13g2_fill_1 FILLER_58_693 ();
 sg13g2_fill_2 FILLER_58_704 ();
 sg13g2_fill_1 FILLER_58_706 ();
 sg13g2_decap_8 FILLER_58_712 ();
 sg13g2_decap_8 FILLER_58_719 ();
 sg13g2_decap_8 FILLER_58_726 ();
 sg13g2_decap_4 FILLER_58_733 ();
 sg13g2_fill_2 FILLER_58_737 ();
 sg13g2_fill_2 FILLER_58_743 ();
 sg13g2_fill_1 FILLER_58_763 ();
 sg13g2_decap_4 FILLER_58_776 ();
 sg13g2_fill_1 FILLER_58_780 ();
 sg13g2_fill_1 FILLER_58_786 ();
 sg13g2_fill_1 FILLER_58_791 ();
 sg13g2_fill_2 FILLER_58_801 ();
 sg13g2_fill_1 FILLER_58_803 ();
 sg13g2_decap_8 FILLER_58_813 ();
 sg13g2_decap_8 FILLER_58_820 ();
 sg13g2_fill_2 FILLER_58_827 ();
 sg13g2_fill_1 FILLER_58_829 ();
 sg13g2_decap_4 FILLER_58_840 ();
 sg13g2_fill_2 FILLER_58_862 ();
 sg13g2_fill_2 FILLER_58_870 ();
 sg13g2_fill_2 FILLER_58_876 ();
 sg13g2_decap_8 FILLER_59_0 ();
 sg13g2_decap_8 FILLER_59_7 ();
 sg13g2_decap_8 FILLER_59_14 ();
 sg13g2_decap_8 FILLER_59_21 ();
 sg13g2_decap_8 FILLER_59_28 ();
 sg13g2_decap_8 FILLER_59_35 ();
 sg13g2_decap_8 FILLER_59_42 ();
 sg13g2_decap_8 FILLER_59_49 ();
 sg13g2_fill_2 FILLER_59_56 ();
 sg13g2_fill_1 FILLER_59_58 ();
 sg13g2_decap_8 FILLER_59_63 ();
 sg13g2_decap_8 FILLER_59_70 ();
 sg13g2_decap_8 FILLER_59_77 ();
 sg13g2_decap_8 FILLER_59_84 ();
 sg13g2_fill_2 FILLER_59_91 ();
 sg13g2_fill_1 FILLER_59_98 ();
 sg13g2_fill_2 FILLER_59_104 ();
 sg13g2_fill_1 FILLER_59_110 ();
 sg13g2_fill_2 FILLER_59_119 ();
 sg13g2_fill_1 FILLER_59_203 ();
 sg13g2_fill_1 FILLER_59_212 ();
 sg13g2_fill_2 FILLER_59_218 ();
 sg13g2_decap_4 FILLER_59_228 ();
 sg13g2_fill_1 FILLER_59_232 ();
 sg13g2_fill_1 FILLER_59_251 ();
 sg13g2_decap_8 FILLER_59_304 ();
 sg13g2_fill_1 FILLER_59_311 ();
 sg13g2_fill_2 FILLER_59_316 ();
 sg13g2_fill_1 FILLER_59_318 ();
 sg13g2_fill_1 FILLER_59_326 ();
 sg13g2_fill_1 FILLER_59_331 ();
 sg13g2_fill_1 FILLER_59_336 ();
 sg13g2_decap_8 FILLER_59_355 ();
 sg13g2_fill_2 FILLER_59_367 ();
 sg13g2_fill_2 FILLER_59_377 ();
 sg13g2_fill_1 FILLER_59_379 ();
 sg13g2_fill_1 FILLER_59_409 ();
 sg13g2_decap_4 FILLER_59_418 ();
 sg13g2_fill_1 FILLER_59_422 ();
 sg13g2_fill_2 FILLER_59_431 ();
 sg13g2_decap_4 FILLER_59_440 ();
 sg13g2_fill_1 FILLER_59_444 ();
 sg13g2_fill_2 FILLER_59_462 ();
 sg13g2_decap_8 FILLER_59_474 ();
 sg13g2_decap_8 FILLER_59_506 ();
 sg13g2_decap_8 FILLER_59_513 ();
 sg13g2_fill_2 FILLER_59_520 ();
 sg13g2_fill_1 FILLER_59_545 ();
 sg13g2_fill_2 FILLER_59_559 ();
 sg13g2_fill_2 FILLER_59_574 ();
 sg13g2_fill_1 FILLER_59_576 ();
 sg13g2_decap_4 FILLER_59_586 ();
 sg13g2_decap_4 FILLER_59_607 ();
 sg13g2_fill_2 FILLER_59_611 ();
 sg13g2_fill_1 FILLER_59_622 ();
 sg13g2_fill_1 FILLER_59_645 ();
 sg13g2_fill_1 FILLER_59_658 ();
 sg13g2_fill_1 FILLER_59_688 ();
 sg13g2_decap_8 FILLER_59_693 ();
 sg13g2_decap_8 FILLER_59_700 ();
 sg13g2_decap_4 FILLER_59_707 ();
 sg13g2_fill_2 FILLER_59_727 ();
 sg13g2_fill_2 FILLER_59_734 ();
 sg13g2_fill_2 FILLER_59_744 ();
 sg13g2_fill_1 FILLER_59_750 ();
 sg13g2_fill_2 FILLER_59_791 ();
 sg13g2_fill_1 FILLER_59_793 ();
 sg13g2_fill_2 FILLER_59_812 ();
 sg13g2_fill_1 FILLER_59_814 ();
 sg13g2_decap_4 FILLER_59_820 ();
 sg13g2_fill_1 FILLER_59_824 ();
 sg13g2_decap_4 FILLER_59_841 ();
 sg13g2_decap_4 FILLER_59_873 ();
 sg13g2_fill_1 FILLER_59_877 ();
 sg13g2_decap_8 FILLER_60_0 ();
 sg13g2_decap_8 FILLER_60_7 ();
 sg13g2_decap_8 FILLER_60_14 ();
 sg13g2_decap_8 FILLER_60_21 ();
 sg13g2_decap_8 FILLER_60_28 ();
 sg13g2_decap_8 FILLER_60_35 ();
 sg13g2_decap_4 FILLER_60_42 ();
 sg13g2_fill_2 FILLER_60_50 ();
 sg13g2_decap_4 FILLER_60_78 ();
 sg13g2_decap_8 FILLER_60_111 ();
 sg13g2_fill_2 FILLER_60_118 ();
 sg13g2_decap_8 FILLER_60_126 ();
 sg13g2_fill_2 FILLER_60_133 ();
 sg13g2_decap_8 FILLER_60_139 ();
 sg13g2_decap_4 FILLER_60_146 ();
 sg13g2_decap_4 FILLER_60_154 ();
 sg13g2_decap_4 FILLER_60_176 ();
 sg13g2_decap_8 FILLER_60_184 ();
 sg13g2_fill_2 FILLER_60_191 ();
 sg13g2_fill_1 FILLER_60_193 ();
 sg13g2_decap_8 FILLER_60_216 ();
 sg13g2_decap_4 FILLER_60_223 ();
 sg13g2_fill_1 FILLER_60_227 ();
 sg13g2_fill_2 FILLER_60_244 ();
 sg13g2_decap_8 FILLER_60_327 ();
 sg13g2_fill_1 FILLER_60_339 ();
 sg13g2_decap_8 FILLER_60_352 ();
 sg13g2_fill_2 FILLER_60_359 ();
 sg13g2_fill_1 FILLER_60_361 ();
 sg13g2_fill_1 FILLER_60_384 ();
 sg13g2_fill_2 FILLER_60_393 ();
 sg13g2_fill_2 FILLER_60_416 ();
 sg13g2_fill_1 FILLER_60_418 ();
 sg13g2_fill_2 FILLER_60_427 ();
 sg13g2_decap_4 FILLER_60_441 ();
 sg13g2_fill_1 FILLER_60_452 ();
 sg13g2_decap_4 FILLER_60_461 ();
 sg13g2_fill_2 FILLER_60_478 ();
 sg13g2_fill_2 FILLER_60_493 ();
 sg13g2_fill_1 FILLER_60_495 ();
 sg13g2_decap_4 FILLER_60_500 ();
 sg13g2_fill_1 FILLER_60_504 ();
 sg13g2_fill_1 FILLER_60_511 ();
 sg13g2_decap_4 FILLER_60_516 ();
 sg13g2_fill_2 FILLER_60_520 ();
 sg13g2_fill_1 FILLER_60_527 ();
 sg13g2_decap_8 FILLER_60_538 ();
 sg13g2_decap_8 FILLER_60_545 ();
 sg13g2_fill_1 FILLER_60_552 ();
 sg13g2_fill_1 FILLER_60_565 ();
 sg13g2_fill_2 FILLER_60_573 ();
 sg13g2_decap_8 FILLER_60_588 ();
 sg13g2_fill_2 FILLER_60_595 ();
 sg13g2_fill_1 FILLER_60_597 ();
 sg13g2_decap_4 FILLER_60_611 ();
 sg13g2_fill_2 FILLER_60_615 ();
 sg13g2_fill_1 FILLER_60_628 ();
 sg13g2_decap_4 FILLER_60_633 ();
 sg13g2_fill_1 FILLER_60_637 ();
 sg13g2_fill_1 FILLER_60_648 ();
 sg13g2_fill_1 FILLER_60_657 ();
 sg13g2_fill_2 FILLER_60_678 ();
 sg13g2_fill_1 FILLER_60_680 ();
 sg13g2_decap_8 FILLER_60_697 ();
 sg13g2_decap_8 FILLER_60_704 ();
 sg13g2_decap_4 FILLER_60_711 ();
 sg13g2_fill_1 FILLER_60_715 ();
 sg13g2_decap_4 FILLER_60_720 ();
 sg13g2_fill_1 FILLER_60_732 ();
 sg13g2_fill_2 FILLER_60_741 ();
 sg13g2_fill_2 FILLER_60_746 ();
 sg13g2_fill_2 FILLER_60_753 ();
 sg13g2_fill_1 FILLER_60_776 ();
 sg13g2_fill_2 FILLER_60_786 ();
 sg13g2_decap_4 FILLER_60_795 ();
 sg13g2_fill_2 FILLER_60_804 ();
 sg13g2_fill_1 FILLER_60_806 ();
 sg13g2_decap_8 FILLER_60_812 ();
 sg13g2_decap_8 FILLER_60_819 ();
 sg13g2_decap_4 FILLER_60_826 ();
 sg13g2_decap_8 FILLER_60_842 ();
 sg13g2_fill_1 FILLER_60_849 ();
 sg13g2_decap_8 FILLER_60_868 ();
 sg13g2_fill_2 FILLER_60_875 ();
 sg13g2_fill_1 FILLER_60_877 ();
 sg13g2_decap_8 FILLER_61_0 ();
 sg13g2_decap_8 FILLER_61_7 ();
 sg13g2_decap_8 FILLER_61_14 ();
 sg13g2_decap_8 FILLER_61_21 ();
 sg13g2_fill_2 FILLER_61_28 ();
 sg13g2_decap_4 FILLER_61_60 ();
 sg13g2_fill_2 FILLER_61_69 ();
 sg13g2_fill_1 FILLER_61_71 ();
 sg13g2_fill_1 FILLER_61_76 ();
 sg13g2_decap_8 FILLER_61_81 ();
 sg13g2_fill_1 FILLER_61_88 ();
 sg13g2_fill_1 FILLER_61_93 ();
 sg13g2_fill_1 FILLER_61_99 ();
 sg13g2_fill_2 FILLER_61_110 ();
 sg13g2_fill_1 FILLER_61_112 ();
 sg13g2_fill_1 FILLER_61_126 ();
 sg13g2_decap_4 FILLER_61_160 ();
 sg13g2_fill_1 FILLER_61_164 ();
 sg13g2_decap_4 FILLER_61_169 ();
 sg13g2_decap_8 FILLER_61_178 ();
 sg13g2_decap_8 FILLER_61_185 ();
 sg13g2_fill_2 FILLER_61_192 ();
 sg13g2_fill_2 FILLER_61_208 ();
 sg13g2_fill_2 FILLER_61_217 ();
 sg13g2_fill_1 FILLER_61_219 ();
 sg13g2_fill_2 FILLER_61_263 ();
 sg13g2_fill_2 FILLER_61_291 ();
 sg13g2_decap_8 FILLER_61_327 ();
 sg13g2_decap_4 FILLER_61_334 ();
 sg13g2_fill_2 FILLER_61_341 ();
 sg13g2_fill_2 FILLER_61_352 ();
 sg13g2_fill_1 FILLER_61_354 ();
 sg13g2_fill_2 FILLER_61_359 ();
 sg13g2_fill_1 FILLER_61_361 ();
 sg13g2_decap_4 FILLER_61_366 ();
 sg13g2_fill_2 FILLER_61_370 ();
 sg13g2_decap_8 FILLER_61_376 ();
 sg13g2_decap_8 FILLER_61_383 ();
 sg13g2_fill_2 FILLER_61_390 ();
 sg13g2_fill_2 FILLER_61_405 ();
 sg13g2_fill_1 FILLER_61_407 ();
 sg13g2_decap_8 FILLER_61_415 ();
 sg13g2_fill_1 FILLER_61_422 ();
 sg13g2_fill_1 FILLER_61_427 ();
 sg13g2_decap_8 FILLER_61_433 ();
 sg13g2_fill_2 FILLER_61_440 ();
 sg13g2_fill_1 FILLER_61_442 ();
 sg13g2_decap_4 FILLER_61_448 ();
 sg13g2_fill_1 FILLER_61_452 ();
 sg13g2_fill_1 FILLER_61_457 ();
 sg13g2_fill_2 FILLER_61_471 ();
 sg13g2_fill_1 FILLER_61_473 ();
 sg13g2_fill_2 FILLER_61_478 ();
 sg13g2_fill_1 FILLER_61_480 ();
 sg13g2_decap_8 FILLER_61_511 ();
 sg13g2_decap_4 FILLER_61_518 ();
 sg13g2_fill_2 FILLER_61_522 ();
 sg13g2_fill_2 FILLER_61_549 ();
 sg13g2_fill_1 FILLER_61_574 ();
 sg13g2_decap_4 FILLER_61_583 ();
 sg13g2_decap_8 FILLER_61_590 ();
 sg13g2_fill_1 FILLER_61_605 ();
 sg13g2_fill_2 FILLER_61_626 ();
 sg13g2_fill_1 FILLER_61_642 ();
 sg13g2_decap_8 FILLER_61_661 ();
 sg13g2_decap_8 FILLER_61_668 ();
 sg13g2_fill_2 FILLER_61_675 ();
 sg13g2_decap_8 FILLER_61_695 ();
 sg13g2_decap_4 FILLER_61_711 ();
 sg13g2_fill_2 FILLER_61_715 ();
 sg13g2_decap_8 FILLER_61_721 ();
 sg13g2_decap_8 FILLER_61_728 ();
 sg13g2_fill_1 FILLER_61_735 ();
 sg13g2_fill_2 FILLER_61_758 ();
 sg13g2_fill_1 FILLER_61_760 ();
 sg13g2_decap_4 FILLER_61_790 ();
 sg13g2_fill_1 FILLER_61_808 ();
 sg13g2_fill_1 FILLER_61_819 ();
 sg13g2_fill_1 FILLER_61_823 ();
 sg13g2_fill_1 FILLER_61_829 ();
 sg13g2_decap_8 FILLER_61_839 ();
 sg13g2_fill_1 FILLER_61_846 ();
 sg13g2_decap_8 FILLER_61_868 ();
 sg13g2_fill_2 FILLER_61_875 ();
 sg13g2_fill_1 FILLER_61_877 ();
 sg13g2_decap_8 FILLER_62_0 ();
 sg13g2_decap_8 FILLER_62_7 ();
 sg13g2_decap_8 FILLER_62_14 ();
 sg13g2_decap_8 FILLER_62_21 ();
 sg13g2_decap_8 FILLER_62_28 ();
 sg13g2_fill_1 FILLER_62_35 ();
 sg13g2_fill_2 FILLER_62_40 ();
 sg13g2_fill_1 FILLER_62_42 ();
 sg13g2_fill_1 FILLER_62_63 ();
 sg13g2_fill_2 FILLER_62_105 ();
 sg13g2_fill_1 FILLER_62_117 ();
 sg13g2_fill_2 FILLER_62_138 ();
 sg13g2_fill_1 FILLER_62_140 ();
 sg13g2_decap_4 FILLER_62_195 ();
 sg13g2_decap_8 FILLER_62_211 ();
 sg13g2_fill_2 FILLER_62_218 ();
 sg13g2_fill_1 FILLER_62_225 ();
 sg13g2_fill_1 FILLER_62_265 ();
 sg13g2_decap_4 FILLER_62_279 ();
 sg13g2_fill_2 FILLER_62_283 ();
 sg13g2_decap_8 FILLER_62_290 ();
 sg13g2_decap_8 FILLER_62_297 ();
 sg13g2_fill_1 FILLER_62_311 ();
 sg13g2_fill_1 FILLER_62_325 ();
 sg13g2_decap_4 FILLER_62_334 ();
 sg13g2_decap_8 FILLER_62_343 ();
 sg13g2_fill_2 FILLER_62_376 ();
 sg13g2_fill_2 FILLER_62_382 ();
 sg13g2_decap_4 FILLER_62_399 ();
 sg13g2_fill_1 FILLER_62_429 ();
 sg13g2_fill_2 FILLER_62_436 ();
 sg13g2_fill_2 FILLER_62_443 ();
 sg13g2_fill_2 FILLER_62_471 ();
 sg13g2_decap_4 FILLER_62_485 ();
 sg13g2_fill_2 FILLER_62_489 ();
 sg13g2_decap_8 FILLER_62_495 ();
 sg13g2_fill_2 FILLER_62_502 ();
 sg13g2_fill_2 FILLER_62_510 ();
 sg13g2_fill_2 FILLER_62_520 ();
 sg13g2_fill_2 FILLER_62_527 ();
 sg13g2_decap_4 FILLER_62_539 ();
 sg13g2_fill_2 FILLER_62_577 ();
 sg13g2_fill_1 FILLER_62_596 ();
 sg13g2_decap_4 FILLER_62_602 ();
 sg13g2_decap_8 FILLER_62_614 ();
 sg13g2_decap_8 FILLER_62_621 ();
 sg13g2_decap_8 FILLER_62_628 ();
 sg13g2_decap_4 FILLER_62_635 ();
 sg13g2_fill_2 FILLER_62_643 ();
 sg13g2_fill_1 FILLER_62_645 ();
 sg13g2_fill_2 FILLER_62_659 ();
 sg13g2_fill_1 FILLER_62_661 ();
 sg13g2_fill_1 FILLER_62_670 ();
 sg13g2_fill_2 FILLER_62_692 ();
 sg13g2_fill_1 FILLER_62_703 ();
 sg13g2_fill_2 FILLER_62_728 ();
 sg13g2_decap_4 FILLER_62_760 ();
 sg13g2_fill_2 FILLER_62_764 ();
 sg13g2_decap_4 FILLER_62_774 ();
 sg13g2_fill_1 FILLER_62_788 ();
 sg13g2_fill_1 FILLER_62_794 ();
 sg13g2_fill_1 FILLER_62_801 ();
 sg13g2_fill_1 FILLER_62_819 ();
 sg13g2_fill_2 FILLER_62_840 ();
 sg13g2_fill_2 FILLER_62_863 ();
 sg13g2_fill_1 FILLER_62_865 ();
 sg13g2_decap_4 FILLER_62_873 ();
 sg13g2_fill_1 FILLER_62_877 ();
 sg13g2_decap_8 FILLER_63_0 ();
 sg13g2_decap_8 FILLER_63_7 ();
 sg13g2_decap_8 FILLER_63_14 ();
 sg13g2_fill_1 FILLER_63_21 ();
 sg13g2_fill_2 FILLER_63_26 ();
 sg13g2_fill_1 FILLER_63_28 ();
 sg13g2_fill_2 FILLER_63_33 ();
 sg13g2_fill_1 FILLER_63_43 ();
 sg13g2_fill_2 FILLER_63_48 ();
 sg13g2_fill_1 FILLER_63_55 ();
 sg13g2_fill_2 FILLER_63_60 ();
 sg13g2_decap_8 FILLER_63_70 ();
 sg13g2_decap_8 FILLER_63_77 ();
 sg13g2_decap_4 FILLER_63_84 ();
 sg13g2_decap_4 FILLER_63_92 ();
 sg13g2_fill_1 FILLER_63_96 ();
 sg13g2_fill_1 FILLER_63_114 ();
 sg13g2_fill_1 FILLER_63_129 ();
 sg13g2_fill_2 FILLER_63_142 ();
 sg13g2_fill_1 FILLER_63_156 ();
 sg13g2_fill_1 FILLER_63_162 ();
 sg13g2_fill_1 FILLER_63_168 ();
 sg13g2_fill_2 FILLER_63_173 ();
 sg13g2_fill_2 FILLER_63_180 ();
 sg13g2_fill_1 FILLER_63_197 ();
 sg13g2_fill_1 FILLER_63_215 ();
 sg13g2_fill_2 FILLER_63_221 ();
 sg13g2_fill_1 FILLER_63_240 ();
 sg13g2_fill_1 FILLER_63_246 ();
 sg13g2_decap_4 FILLER_63_279 ();
 sg13g2_fill_1 FILLER_63_283 ();
 sg13g2_fill_1 FILLER_63_314 ();
 sg13g2_fill_2 FILLER_63_372 ();
 sg13g2_fill_2 FILLER_63_382 ();
 sg13g2_decap_8 FILLER_63_402 ();
 sg13g2_fill_1 FILLER_63_409 ();
 sg13g2_decap_8 FILLER_63_414 ();
 sg13g2_decap_4 FILLER_63_421 ();
 sg13g2_fill_1 FILLER_63_454 ();
 sg13g2_fill_2 FILLER_63_460 ();
 sg13g2_fill_1 FILLER_63_462 ();
 sg13g2_fill_2 FILLER_63_475 ();
 sg13g2_fill_1 FILLER_63_477 ();
 sg13g2_fill_1 FILLER_63_483 ();
 sg13g2_fill_1 FILLER_63_504 ();
 sg13g2_decap_4 FILLER_63_520 ();
 sg13g2_fill_2 FILLER_63_524 ();
 sg13g2_fill_2 FILLER_63_537 ();
 sg13g2_fill_1 FILLER_63_539 ();
 sg13g2_fill_2 FILLER_63_554 ();
 sg13g2_fill_1 FILLER_63_556 ();
 sg13g2_fill_1 FILLER_63_576 ();
 sg13g2_fill_2 FILLER_63_583 ();
 sg13g2_fill_2 FILLER_63_592 ();
 sg13g2_fill_2 FILLER_63_606 ();
 sg13g2_fill_2 FILLER_63_639 ();
 sg13g2_fill_1 FILLER_63_641 ();
 sg13g2_decap_8 FILLER_63_652 ();
 sg13g2_fill_2 FILLER_63_659 ();
 sg13g2_fill_1 FILLER_63_661 ();
 sg13g2_decap_4 FILLER_63_674 ();
 sg13g2_fill_2 FILLER_63_678 ();
 sg13g2_decap_8 FILLER_63_729 ();
 sg13g2_fill_1 FILLER_63_736 ();
 sg13g2_decap_4 FILLER_63_750 ();
 sg13g2_fill_2 FILLER_63_754 ();
 sg13g2_decap_4 FILLER_63_769 ();
 sg13g2_fill_1 FILLER_63_773 ();
 sg13g2_fill_1 FILLER_63_803 ();
 sg13g2_decap_8 FILLER_63_809 ();
 sg13g2_fill_1 FILLER_63_816 ();
 sg13g2_decap_4 FILLER_63_839 ();
 sg13g2_decap_8 FILLER_63_847 ();
 sg13g2_decap_8 FILLER_63_854 ();
 sg13g2_decap_8 FILLER_63_861 ();
 sg13g2_decap_8 FILLER_63_868 ();
 sg13g2_fill_2 FILLER_63_875 ();
 sg13g2_fill_1 FILLER_63_877 ();
 sg13g2_decap_8 FILLER_64_0 ();
 sg13g2_decap_4 FILLER_64_7 ();
 sg13g2_fill_2 FILLER_64_11 ();
 sg13g2_fill_1 FILLER_64_69 ();
 sg13g2_decap_8 FILLER_64_101 ();
 sg13g2_decap_8 FILLER_64_108 ();
 sg13g2_decap_4 FILLER_64_115 ();
 sg13g2_decap_4 FILLER_64_124 ();
 sg13g2_fill_1 FILLER_64_128 ();
 sg13g2_decap_4 FILLER_64_132 ();
 sg13g2_fill_2 FILLER_64_150 ();
 sg13g2_fill_1 FILLER_64_152 ();
 sg13g2_fill_1 FILLER_64_222 ();
 sg13g2_fill_1 FILLER_64_231 ();
 sg13g2_fill_1 FILLER_64_237 ();
 sg13g2_fill_1 FILLER_64_245 ();
 sg13g2_fill_1 FILLER_64_251 ();
 sg13g2_fill_1 FILLER_64_257 ();
 sg13g2_decap_4 FILLER_64_272 ();
 sg13g2_fill_1 FILLER_64_276 ();
 sg13g2_decap_4 FILLER_64_290 ();
 sg13g2_fill_1 FILLER_64_299 ();
 sg13g2_fill_1 FILLER_64_318 ();
 sg13g2_fill_1 FILLER_64_344 ();
 sg13g2_fill_1 FILLER_64_349 ();
 sg13g2_fill_2 FILLER_64_368 ();
 sg13g2_fill_2 FILLER_64_400 ();
 sg13g2_fill_1 FILLER_64_420 ();
 sg13g2_decap_4 FILLER_64_439 ();
 sg13g2_fill_2 FILLER_64_443 ();
 sg13g2_decap_4 FILLER_64_455 ();
 sg13g2_fill_1 FILLER_64_459 ();
 sg13g2_decap_8 FILLER_64_469 ();
 sg13g2_fill_2 FILLER_64_520 ();
 sg13g2_decap_4 FILLER_64_544 ();
 sg13g2_fill_2 FILLER_64_553 ();
 sg13g2_decap_4 FILLER_64_563 ();
 sg13g2_fill_2 FILLER_64_577 ();
 sg13g2_fill_1 FILLER_64_579 ();
 sg13g2_fill_1 FILLER_64_591 ();
 sg13g2_fill_2 FILLER_64_604 ();
 sg13g2_decap_4 FILLER_64_611 ();
 sg13g2_fill_2 FILLER_64_615 ();
 sg13g2_decap_8 FILLER_64_625 ();
 sg13g2_decap_4 FILLER_64_632 ();
 sg13g2_fill_1 FILLER_64_636 ();
 sg13g2_decap_4 FILLER_64_677 ();
 sg13g2_fill_1 FILLER_64_681 ();
 sg13g2_fill_2 FILLER_64_686 ();
 sg13g2_decap_4 FILLER_64_695 ();
 sg13g2_fill_2 FILLER_64_704 ();
 sg13g2_fill_1 FILLER_64_706 ();
 sg13g2_decap_8 FILLER_64_716 ();
 sg13g2_decap_8 FILLER_64_723 ();
 sg13g2_decap_4 FILLER_64_730 ();
 sg13g2_decap_4 FILLER_64_764 ();
 sg13g2_fill_2 FILLER_64_768 ();
 sg13g2_decap_4 FILLER_64_774 ();
 sg13g2_fill_1 FILLER_64_778 ();
 sg13g2_decap_8 FILLER_64_785 ();
 sg13g2_decap_4 FILLER_64_792 ();
 sg13g2_decap_8 FILLER_64_805 ();
 sg13g2_decap_8 FILLER_64_812 ();
 sg13g2_decap_8 FILLER_64_819 ();
 sg13g2_decap_8 FILLER_64_826 ();
 sg13g2_decap_8 FILLER_64_833 ();
 sg13g2_decap_8 FILLER_64_840 ();
 sg13g2_decap_8 FILLER_64_847 ();
 sg13g2_decap_8 FILLER_64_854 ();
 sg13g2_decap_8 FILLER_64_861 ();
 sg13g2_decap_8 FILLER_64_868 ();
 sg13g2_fill_2 FILLER_64_875 ();
 sg13g2_fill_1 FILLER_64_877 ();
 sg13g2_decap_8 FILLER_65_0 ();
 sg13g2_decap_8 FILLER_65_11 ();
 sg13g2_fill_1 FILLER_65_18 ();
 sg13g2_decap_8 FILLER_65_32 ();
 sg13g2_fill_1 FILLER_65_39 ();
 sg13g2_fill_1 FILLER_65_50 ();
 sg13g2_decap_4 FILLER_65_56 ();
 sg13g2_fill_2 FILLER_65_60 ();
 sg13g2_fill_1 FILLER_65_76 ();
 sg13g2_fill_1 FILLER_65_81 ();
 sg13g2_fill_1 FILLER_65_90 ();
 sg13g2_fill_2 FILLER_65_95 ();
 sg13g2_fill_2 FILLER_65_101 ();
 sg13g2_fill_2 FILLER_65_107 ();
 sg13g2_fill_1 FILLER_65_109 ();
 sg13g2_decap_4 FILLER_65_136 ();
 sg13g2_fill_2 FILLER_65_140 ();
 sg13g2_decap_4 FILLER_65_168 ();
 sg13g2_fill_2 FILLER_65_172 ();
 sg13g2_decap_8 FILLER_65_178 ();
 sg13g2_decap_8 FILLER_65_185 ();
 sg13g2_fill_1 FILLER_65_197 ();
 sg13g2_decap_4 FILLER_65_202 ();
 sg13g2_decap_4 FILLER_65_210 ();
 sg13g2_fill_2 FILLER_65_251 ();
 sg13g2_fill_2 FILLER_65_276 ();
 sg13g2_fill_1 FILLER_65_278 ();
 sg13g2_fill_2 FILLER_65_283 ();
 sg13g2_fill_1 FILLER_65_285 ();
 sg13g2_fill_2 FILLER_65_294 ();
 sg13g2_fill_1 FILLER_65_306 ();
 sg13g2_decap_8 FILLER_65_325 ();
 sg13g2_fill_1 FILLER_65_340 ();
 sg13g2_fill_1 FILLER_65_345 ();
 sg13g2_fill_1 FILLER_65_350 ();
 sg13g2_fill_2 FILLER_65_356 ();
 sg13g2_fill_2 FILLER_65_376 ();
 sg13g2_fill_2 FILLER_65_382 ();
 sg13g2_fill_1 FILLER_65_384 ();
 sg13g2_decap_8 FILLER_65_411 ();
 sg13g2_fill_2 FILLER_65_448 ();
 sg13g2_fill_1 FILLER_65_485 ();
 sg13g2_fill_1 FILLER_65_505 ();
 sg13g2_fill_2 FILLER_65_521 ();
 sg13g2_fill_1 FILLER_65_528 ();
 sg13g2_fill_2 FILLER_65_538 ();
 sg13g2_decap_8 FILLER_65_594 ();
 sg13g2_decap_8 FILLER_65_662 ();
 sg13g2_fill_1 FILLER_65_669 ();
 sg13g2_fill_1 FILLER_65_673 ();
 sg13g2_decap_4 FILLER_65_704 ();
 sg13g2_decap_8 FILLER_65_734 ();
 sg13g2_fill_2 FILLER_65_741 ();
 sg13g2_fill_1 FILLER_65_743 ();
 sg13g2_decap_4 FILLER_65_748 ();
 sg13g2_decap_8 FILLER_65_760 ();
 sg13g2_decap_8 FILLER_65_767 ();
 sg13g2_decap_4 FILLER_65_774 ();
 sg13g2_fill_1 FILLER_65_778 ();
 sg13g2_decap_8 FILLER_65_783 ();
 sg13g2_decap_4 FILLER_65_790 ();
 sg13g2_fill_2 FILLER_65_794 ();
 sg13g2_decap_8 FILLER_65_800 ();
 sg13g2_decap_8 FILLER_65_807 ();
 sg13g2_decap_8 FILLER_65_814 ();
 sg13g2_decap_8 FILLER_65_821 ();
 sg13g2_decap_8 FILLER_65_828 ();
 sg13g2_decap_8 FILLER_65_835 ();
 sg13g2_decap_8 FILLER_65_842 ();
 sg13g2_decap_8 FILLER_65_849 ();
 sg13g2_decap_8 FILLER_65_856 ();
 sg13g2_decap_8 FILLER_65_863 ();
 sg13g2_decap_8 FILLER_65_870 ();
 sg13g2_fill_1 FILLER_65_877 ();
 sg13g2_fill_2 FILLER_66_26 ();
 sg13g2_fill_1 FILLER_66_28 ();
 sg13g2_fill_2 FILLER_66_34 ();
 sg13g2_fill_1 FILLER_66_87 ();
 sg13g2_fill_1 FILLER_66_114 ();
 sg13g2_fill_2 FILLER_66_119 ();
 sg13g2_fill_2 FILLER_66_147 ();
 sg13g2_fill_1 FILLER_66_175 ();
 sg13g2_decap_4 FILLER_66_180 ();
 sg13g2_fill_2 FILLER_66_184 ();
 sg13g2_decap_8 FILLER_66_191 ();
 sg13g2_fill_2 FILLER_66_228 ();
 sg13g2_fill_1 FILLER_66_242 ();
 sg13g2_decap_8 FILLER_66_277 ();
 sg13g2_fill_1 FILLER_66_289 ();
 sg13g2_fill_1 FILLER_66_296 ();
 sg13g2_fill_1 FILLER_66_304 ();
 sg13g2_fill_2 FILLER_66_313 ();
 sg13g2_fill_1 FILLER_66_330 ();
 sg13g2_fill_2 FILLER_66_351 ();
 sg13g2_fill_1 FILLER_66_367 ();
 sg13g2_fill_1 FILLER_66_376 ();
 sg13g2_fill_1 FILLER_66_401 ();
 sg13g2_decap_8 FILLER_66_407 ();
 sg13g2_fill_2 FILLER_66_414 ();
 sg13g2_fill_1 FILLER_66_416 ();
 sg13g2_fill_1 FILLER_66_425 ();
 sg13g2_decap_8 FILLER_66_431 ();
 sg13g2_fill_2 FILLER_66_438 ();
 sg13g2_fill_1 FILLER_66_458 ();
 sg13g2_decap_8 FILLER_66_471 ();
 sg13g2_fill_1 FILLER_66_504 ();
 sg13g2_decap_8 FILLER_66_536 ();
 sg13g2_decap_4 FILLER_66_563 ();
 sg13g2_fill_1 FILLER_66_567 ();
 sg13g2_fill_2 FILLER_66_573 ();
 sg13g2_decap_8 FILLER_66_584 ();
 sg13g2_decap_4 FILLER_66_591 ();
 sg13g2_fill_1 FILLER_66_600 ();
 sg13g2_fill_1 FILLER_66_630 ();
 sg13g2_fill_1 FILLER_66_636 ();
 sg13g2_fill_1 FILLER_66_665 ();
 sg13g2_fill_1 FILLER_66_670 ();
 sg13g2_decap_4 FILLER_66_691 ();
 sg13g2_fill_1 FILLER_66_705 ();
 sg13g2_fill_2 FILLER_66_713 ();
 sg13g2_decap_4 FILLER_66_719 ();
 sg13g2_decap_4 FILLER_66_728 ();
 sg13g2_fill_2 FILLER_66_732 ();
 sg13g2_decap_8 FILLER_66_739 ();
 sg13g2_fill_2 FILLER_66_798 ();
 sg13g2_fill_1 FILLER_66_800 ();
 sg13g2_decap_8 FILLER_66_827 ();
 sg13g2_decap_8 FILLER_66_834 ();
 sg13g2_decap_8 FILLER_66_841 ();
 sg13g2_decap_8 FILLER_66_848 ();
 sg13g2_decap_8 FILLER_66_855 ();
 sg13g2_decap_8 FILLER_66_862 ();
 sg13g2_decap_8 FILLER_66_869 ();
 sg13g2_fill_2 FILLER_66_876 ();
 sg13g2_decap_8 FILLER_67_0 ();
 sg13g2_decap_8 FILLER_67_7 ();
 sg13g2_decap_8 FILLER_67_14 ();
 sg13g2_decap_4 FILLER_67_21 ();
 sg13g2_fill_2 FILLER_67_41 ();
 sg13g2_fill_2 FILLER_67_47 ();
 sg13g2_fill_1 FILLER_67_49 ();
 sg13g2_fill_2 FILLER_67_58 ();
 sg13g2_fill_1 FILLER_67_60 ();
 sg13g2_fill_2 FILLER_67_80 ();
 sg13g2_fill_2 FILLER_67_104 ();
 sg13g2_decap_8 FILLER_67_110 ();
 sg13g2_fill_1 FILLER_67_117 ();
 sg13g2_decap_4 FILLER_67_123 ();
 sg13g2_fill_1 FILLER_67_127 ();
 sg13g2_decap_8 FILLER_67_132 ();
 sg13g2_fill_2 FILLER_67_139 ();
 sg13g2_fill_1 FILLER_67_141 ();
 sg13g2_fill_1 FILLER_67_146 ();
 sg13g2_fill_1 FILLER_67_151 ();
 sg13g2_fill_1 FILLER_67_157 ();
 sg13g2_fill_2 FILLER_67_193 ();
 sg13g2_decap_8 FILLER_67_199 ();
 sg13g2_decap_4 FILLER_67_206 ();
 sg13g2_fill_1 FILLER_67_214 ();
 sg13g2_decap_4 FILLER_67_247 ();
 sg13g2_fill_1 FILLER_67_259 ();
 sg13g2_fill_2 FILLER_67_265 ();
 sg13g2_fill_2 FILLER_67_283 ();
 sg13g2_fill_1 FILLER_67_295 ();
 sg13g2_fill_2 FILLER_67_305 ();
 sg13g2_fill_1 FILLER_67_307 ();
 sg13g2_decap_8 FILLER_67_312 ();
 sg13g2_fill_1 FILLER_67_319 ();
 sg13g2_fill_1 FILLER_67_326 ();
 sg13g2_fill_1 FILLER_67_335 ();
 sg13g2_fill_2 FILLER_67_346 ();
 sg13g2_fill_2 FILLER_67_352 ();
 sg13g2_fill_2 FILLER_67_358 ();
 sg13g2_fill_2 FILLER_67_393 ();
 sg13g2_decap_4 FILLER_67_402 ();
 sg13g2_fill_1 FILLER_67_406 ();
 sg13g2_fill_2 FILLER_67_443 ();
 sg13g2_decap_8 FILLER_67_450 ();
 sg13g2_fill_1 FILLER_67_457 ();
 sg13g2_fill_1 FILLER_67_468 ();
 sg13g2_decap_8 FILLER_67_474 ();
 sg13g2_decap_4 FILLER_67_481 ();
 sg13g2_fill_1 FILLER_67_485 ();
 sg13g2_decap_8 FILLER_67_491 ();
 sg13g2_fill_2 FILLER_67_498 ();
 sg13g2_fill_1 FILLER_67_500 ();
 sg13g2_fill_1 FILLER_67_506 ();
 sg13g2_fill_2 FILLER_67_514 ();
 sg13g2_fill_1 FILLER_67_516 ();
 sg13g2_fill_2 FILLER_67_521 ();
 sg13g2_fill_1 FILLER_67_523 ();
 sg13g2_decap_8 FILLER_67_529 ();
 sg13g2_fill_2 FILLER_67_536 ();
 sg13g2_fill_1 FILLER_67_538 ();
 sg13g2_decap_8 FILLER_67_544 ();
 sg13g2_fill_2 FILLER_67_551 ();
 sg13g2_fill_2 FILLER_67_558 ();
 sg13g2_fill_2 FILLER_67_565 ();
 sg13g2_fill_1 FILLER_67_567 ();
 sg13g2_decap_8 FILLER_67_592 ();
 sg13g2_decap_8 FILLER_67_599 ();
 sg13g2_fill_2 FILLER_67_606 ();
 sg13g2_fill_1 FILLER_67_608 ();
 sg13g2_fill_1 FILLER_67_618 ();
 sg13g2_fill_1 FILLER_67_626 ();
 sg13g2_decap_4 FILLER_67_632 ();
 sg13g2_fill_1 FILLER_67_636 ();
 sg13g2_fill_2 FILLER_67_642 ();
 sg13g2_fill_1 FILLER_67_644 ();
 sg13g2_fill_2 FILLER_67_681 ();
 sg13g2_fill_1 FILLER_67_683 ();
 sg13g2_fill_2 FILLER_67_697 ();
 sg13g2_fill_2 FILLER_67_735 ();
 sg13g2_fill_2 FILLER_67_740 ();
 sg13g2_fill_1 FILLER_67_742 ();
 sg13g2_decap_8 FILLER_67_754 ();
 sg13g2_fill_1 FILLER_67_761 ();
 sg13g2_fill_1 FILLER_67_766 ();
 sg13g2_decap_8 FILLER_67_783 ();
 sg13g2_fill_2 FILLER_67_812 ();
 sg13g2_decap_8 FILLER_67_825 ();
 sg13g2_decap_8 FILLER_67_832 ();
 sg13g2_decap_8 FILLER_67_839 ();
 sg13g2_decap_8 FILLER_67_846 ();
 sg13g2_decap_8 FILLER_67_853 ();
 sg13g2_decap_8 FILLER_67_860 ();
 sg13g2_decap_8 FILLER_67_867 ();
 sg13g2_decap_4 FILLER_67_874 ();
 sg13g2_decap_4 FILLER_68_0 ();
 sg13g2_fill_2 FILLER_68_4 ();
 sg13g2_decap_8 FILLER_68_10 ();
 sg13g2_decap_4 FILLER_68_17 ();
 sg13g2_fill_1 FILLER_68_33 ();
 sg13g2_decap_4 FILLER_68_40 ();
 sg13g2_fill_2 FILLER_68_44 ();
 sg13g2_fill_1 FILLER_68_63 ();
 sg13g2_fill_1 FILLER_68_101 ();
 sg13g2_fill_1 FILLER_68_108 ();
 sg13g2_fill_1 FILLER_68_115 ();
 sg13g2_fill_1 FILLER_68_122 ();
 sg13g2_fill_2 FILLER_68_135 ();
 sg13g2_fill_1 FILLER_68_137 ();
 sg13g2_fill_2 FILLER_68_171 ();
 sg13g2_fill_2 FILLER_68_177 ();
 sg13g2_decap_4 FILLER_68_183 ();
 sg13g2_decap_4 FILLER_68_192 ();
 sg13g2_fill_1 FILLER_68_196 ();
 sg13g2_decap_4 FILLER_68_202 ();
 sg13g2_decap_4 FILLER_68_211 ();
 sg13g2_fill_1 FILLER_68_215 ();
 sg13g2_decap_4 FILLER_68_222 ();
 sg13g2_fill_1 FILLER_68_226 ();
 sg13g2_decap_8 FILLER_68_232 ();
 sg13g2_fill_2 FILLER_68_239 ();
 sg13g2_fill_1 FILLER_68_249 ();
 sg13g2_decap_8 FILLER_68_276 ();
 sg13g2_decap_4 FILLER_68_288 ();
 sg13g2_fill_1 FILLER_68_292 ();
 sg13g2_decap_8 FILLER_68_296 ();
 sg13g2_fill_1 FILLER_68_307 ();
 sg13g2_fill_2 FILLER_68_316 ();
 sg13g2_fill_1 FILLER_68_322 ();
 sg13g2_fill_2 FILLER_68_328 ();
 sg13g2_fill_1 FILLER_68_334 ();
 sg13g2_fill_1 FILLER_68_341 ();
 sg13g2_fill_2 FILLER_68_347 ();
 sg13g2_fill_2 FILLER_68_353 ();
 sg13g2_fill_1 FILLER_68_355 ();
 sg13g2_fill_1 FILLER_68_364 ();
 sg13g2_fill_1 FILLER_68_368 ();
 sg13g2_decap_4 FILLER_68_374 ();
 sg13g2_fill_1 FILLER_68_378 ();
 sg13g2_decap_8 FILLER_68_387 ();
 sg13g2_decap_4 FILLER_68_394 ();
 sg13g2_fill_2 FILLER_68_398 ();
 sg13g2_fill_2 FILLER_68_413 ();
 sg13g2_fill_1 FILLER_68_420 ();
 sg13g2_fill_1 FILLER_68_426 ();
 sg13g2_decap_8 FILLER_68_432 ();
 sg13g2_decap_4 FILLER_68_439 ();
 sg13g2_fill_1 FILLER_68_443 ();
 sg13g2_fill_2 FILLER_68_463 ();
 sg13g2_fill_2 FILLER_68_504 ();
 sg13g2_fill_1 FILLER_68_506 ();
 sg13g2_decap_4 FILLER_68_528 ();
 sg13g2_fill_1 FILLER_68_536 ();
 sg13g2_decap_8 FILLER_68_562 ();
 sg13g2_decap_4 FILLER_68_569 ();
 sg13g2_fill_1 FILLER_68_623 ();
 sg13g2_fill_2 FILLER_68_634 ();
 sg13g2_fill_1 FILLER_68_636 ();
 sg13g2_decap_8 FILLER_68_647 ();
 sg13g2_decap_8 FILLER_68_654 ();
 sg13g2_decap_4 FILLER_68_661 ();
 sg13g2_fill_2 FILLER_68_665 ();
 sg13g2_fill_1 FILLER_68_677 ();
 sg13g2_decap_8 FILLER_68_682 ();
 sg13g2_fill_1 FILLER_68_689 ();
 sg13g2_fill_2 FILLER_68_722 ();
 sg13g2_fill_1 FILLER_68_768 ();
 sg13g2_fill_1 FILLER_68_803 ();
 sg13g2_fill_2 FILLER_68_809 ();
 sg13g2_decap_8 FILLER_68_827 ();
 sg13g2_decap_8 FILLER_68_834 ();
 sg13g2_decap_8 FILLER_68_841 ();
 sg13g2_decap_8 FILLER_68_848 ();
 sg13g2_decap_8 FILLER_68_855 ();
 sg13g2_decap_8 FILLER_68_862 ();
 sg13g2_decap_8 FILLER_68_869 ();
 sg13g2_fill_2 FILLER_68_876 ();
 sg13g2_fill_1 FILLER_69_0 ();
 sg13g2_fill_1 FILLER_69_51 ();
 sg13g2_fill_1 FILLER_69_62 ();
 sg13g2_decap_4 FILLER_69_79 ();
 sg13g2_fill_2 FILLER_69_83 ();
 sg13g2_decap_4 FILLER_69_103 ();
 sg13g2_fill_2 FILLER_69_107 ();
 sg13g2_decap_8 FILLER_69_117 ();
 sg13g2_decap_8 FILLER_69_124 ();
 sg13g2_fill_1 FILLER_69_131 ();
 sg13g2_decap_8 FILLER_69_136 ();
 sg13g2_fill_2 FILLER_69_143 ();
 sg13g2_fill_2 FILLER_69_179 ();
 sg13g2_fill_1 FILLER_69_181 ();
 sg13g2_fill_2 FILLER_69_219 ();
 sg13g2_fill_1 FILLER_69_221 ();
 sg13g2_fill_2 FILLER_69_251 ();
 sg13g2_fill_1 FILLER_69_259 ();
 sg13g2_fill_1 FILLER_69_286 ();
 sg13g2_fill_1 FILLER_69_313 ();
 sg13g2_fill_1 FILLER_69_317 ();
 sg13g2_decap_8 FILLER_69_326 ();
 sg13g2_decap_4 FILLER_69_350 ();
 sg13g2_fill_1 FILLER_69_367 ();
 sg13g2_fill_1 FILLER_69_376 ();
 sg13g2_fill_1 FILLER_69_381 ();
 sg13g2_fill_1 FILLER_69_387 ();
 sg13g2_fill_1 FILLER_69_395 ();
 sg13g2_decap_8 FILLER_69_409 ();
 sg13g2_fill_2 FILLER_69_416 ();
 sg13g2_fill_1 FILLER_69_418 ();
 sg13g2_fill_1 FILLER_69_475 ();
 sg13g2_decap_8 FILLER_69_484 ();
 sg13g2_decap_4 FILLER_69_491 ();
 sg13g2_fill_1 FILLER_69_495 ();
 sg13g2_fill_1 FILLER_69_501 ();
 sg13g2_fill_2 FILLER_69_520 ();
 sg13g2_decap_8 FILLER_69_539 ();
 sg13g2_fill_1 FILLER_69_546 ();
 sg13g2_fill_2 FILLER_69_568 ();
 sg13g2_decap_4 FILLER_69_578 ();
 sg13g2_fill_2 FILLER_69_629 ();
 sg13g2_fill_2 FILLER_69_660 ();
 sg13g2_fill_2 FILLER_69_667 ();
 sg13g2_fill_1 FILLER_69_698 ();
 sg13g2_fill_1 FILLER_69_742 ();
 sg13g2_decap_8 FILLER_69_752 ();
 sg13g2_decap_4 FILLER_69_759 ();
 sg13g2_fill_2 FILLER_69_773 ();
 sg13g2_decap_4 FILLER_69_779 ();
 sg13g2_fill_1 FILLER_69_783 ();
 sg13g2_decap_8 FILLER_69_840 ();
 sg13g2_decap_8 FILLER_69_847 ();
 sg13g2_decap_8 FILLER_69_854 ();
 sg13g2_decap_8 FILLER_69_861 ();
 sg13g2_decap_8 FILLER_69_868 ();
 sg13g2_fill_2 FILLER_69_875 ();
 sg13g2_fill_1 FILLER_69_877 ();
 sg13g2_fill_2 FILLER_70_26 ();
 sg13g2_decap_8 FILLER_70_46 ();
 sg13g2_decap_8 FILLER_70_76 ();
 sg13g2_fill_2 FILLER_70_83 ();
 sg13g2_fill_1 FILLER_70_85 ();
 sg13g2_fill_2 FILLER_70_99 ();
 sg13g2_decap_8 FILLER_70_112 ();
 sg13g2_decap_4 FILLER_70_150 ();
 sg13g2_fill_2 FILLER_70_154 ();
 sg13g2_fill_2 FILLER_70_167 ();
 sg13g2_fill_1 FILLER_70_169 ();
 sg13g2_fill_2 FILLER_70_178 ();
 sg13g2_fill_1 FILLER_70_190 ();
 sg13g2_fill_1 FILLER_70_196 ();
 sg13g2_fill_1 FILLER_70_205 ();
 sg13g2_fill_1 FILLER_70_211 ();
 sg13g2_fill_1 FILLER_70_231 ();
 sg13g2_fill_1 FILLER_70_237 ();
 sg13g2_fill_1 FILLER_70_270 ();
 sg13g2_decap_8 FILLER_70_275 ();
 sg13g2_fill_1 FILLER_70_282 ();
 sg13g2_decap_8 FILLER_70_286 ();
 sg13g2_fill_2 FILLER_70_293 ();
 sg13g2_fill_2 FILLER_70_299 ();
 sg13g2_fill_2 FILLER_70_337 ();
 sg13g2_fill_1 FILLER_70_339 ();
 sg13g2_fill_1 FILLER_70_378 ();
 sg13g2_fill_1 FILLER_70_389 ();
 sg13g2_fill_1 FILLER_70_416 ();
 sg13g2_fill_1 FILLER_70_443 ();
 sg13g2_fill_2 FILLER_70_448 ();
 sg13g2_decap_8 FILLER_70_454 ();
 sg13g2_decap_4 FILLER_70_486 ();
 sg13g2_fill_2 FILLER_70_516 ();
 sg13g2_fill_1 FILLER_70_518 ();
 sg13g2_decap_8 FILLER_70_522 ();
 sg13g2_decap_8 FILLER_70_529 ();
 sg13g2_fill_1 FILLER_70_536 ();
 sg13g2_decap_4 FILLER_70_568 ();
 sg13g2_fill_2 FILLER_70_572 ();
 sg13g2_decap_4 FILLER_70_581 ();
 sg13g2_fill_2 FILLER_70_585 ();
 sg13g2_fill_2 FILLER_70_626 ();
 sg13g2_decap_8 FILLER_70_634 ();
 sg13g2_fill_1 FILLER_70_641 ();
 sg13g2_fill_2 FILLER_70_646 ();
 sg13g2_fill_2 FILLER_70_654 ();
 sg13g2_fill_1 FILLER_70_656 ();
 sg13g2_fill_1 FILLER_70_661 ();
 sg13g2_decap_8 FILLER_70_674 ();
 sg13g2_decap_8 FILLER_70_681 ();
 sg13g2_decap_8 FILLER_70_697 ();
 sg13g2_fill_2 FILLER_70_704 ();
 sg13g2_fill_1 FILLER_70_706 ();
 sg13g2_fill_2 FILLER_70_711 ();
 sg13g2_decap_4 FILLER_70_717 ();
 sg13g2_fill_2 FILLER_70_726 ();
 sg13g2_fill_1 FILLER_70_728 ();
 sg13g2_fill_2 FILLER_70_753 ();
 sg13g2_fill_1 FILLER_70_804 ();
 sg13g2_fill_1 FILLER_70_809 ();
 sg13g2_decap_8 FILLER_70_840 ();
 sg13g2_decap_8 FILLER_70_847 ();
 sg13g2_decap_8 FILLER_70_854 ();
 sg13g2_decap_8 FILLER_70_861 ();
 sg13g2_decap_8 FILLER_70_868 ();
 sg13g2_fill_2 FILLER_70_875 ();
 sg13g2_fill_1 FILLER_70_877 ();
 sg13g2_fill_2 FILLER_71_0 ();
 sg13g2_fill_1 FILLER_71_2 ();
 sg13g2_fill_1 FILLER_71_29 ();
 sg13g2_fill_2 FILLER_71_45 ();
 sg13g2_decap_8 FILLER_71_51 ();
 sg13g2_fill_1 FILLER_71_58 ();
 sg13g2_fill_1 FILLER_71_63 ();
 sg13g2_fill_1 FILLER_71_69 ();
 sg13g2_fill_1 FILLER_71_104 ();
 sg13g2_fill_2 FILLER_71_109 ();
 sg13g2_fill_1 FILLER_71_111 ();
 sg13g2_fill_2 FILLER_71_142 ();
 sg13g2_fill_1 FILLER_71_149 ();
 sg13g2_fill_2 FILLER_71_154 ();
 sg13g2_fill_1 FILLER_71_161 ();
 sg13g2_fill_1 FILLER_71_168 ();
 sg13g2_fill_2 FILLER_71_183 ();
 sg13g2_fill_1 FILLER_71_185 ();
 sg13g2_fill_2 FILLER_71_194 ();
 sg13g2_fill_2 FILLER_71_231 ();
 sg13g2_fill_1 FILLER_71_233 ();
 sg13g2_fill_1 FILLER_71_256 ();
 sg13g2_fill_2 FILLER_71_262 ();
 sg13g2_fill_1 FILLER_71_264 ();
 sg13g2_fill_1 FILLER_71_285 ();
 sg13g2_decap_4 FILLER_71_298 ();
 sg13g2_fill_2 FILLER_71_307 ();
 sg13g2_decap_4 FILLER_71_314 ();
 sg13g2_fill_1 FILLER_71_318 ();
 sg13g2_decap_8 FILLER_71_323 ();
 sg13g2_decap_4 FILLER_71_330 ();
 sg13g2_fill_2 FILLER_71_344 ();
 sg13g2_fill_1 FILLER_71_346 ();
 sg13g2_decap_4 FILLER_71_351 ();
 sg13g2_fill_1 FILLER_71_365 ();
 sg13g2_fill_1 FILLER_71_396 ();
 sg13g2_decap_4 FILLER_71_401 ();
 sg13g2_decap_4 FILLER_71_411 ();
 sg13g2_fill_1 FILLER_71_433 ();
 sg13g2_fill_1 FILLER_71_440 ();
 sg13g2_fill_2 FILLER_71_450 ();
 sg13g2_fill_2 FILLER_71_457 ();
 sg13g2_fill_2 FILLER_71_485 ();
 sg13g2_decap_4 FILLER_71_491 ();
 sg13g2_fill_2 FILLER_71_495 ();
 sg13g2_decap_4 FILLER_71_501 ();
 sg13g2_fill_1 FILLER_71_505 ();
 sg13g2_decap_4 FILLER_71_540 ();
 sg13g2_fill_1 FILLER_71_548 ();
 sg13g2_decap_8 FILLER_71_553 ();
 sg13g2_decap_4 FILLER_71_560 ();
 sg13g2_fill_1 FILLER_71_564 ();
 sg13g2_fill_2 FILLER_71_575 ();
 sg13g2_fill_1 FILLER_71_581 ();
 sg13g2_fill_1 FILLER_71_600 ();
 sg13g2_fill_1 FILLER_71_605 ();
 sg13g2_fill_1 FILLER_71_610 ();
 sg13g2_decap_8 FILLER_71_615 ();
 sg13g2_decap_4 FILLER_71_622 ();
 sg13g2_fill_1 FILLER_71_667 ();
 sg13g2_fill_2 FILLER_71_704 ();
 sg13g2_fill_1 FILLER_71_706 ();
 sg13g2_fill_2 FILLER_71_717 ();
 sg13g2_fill_1 FILLER_71_719 ();
 sg13g2_fill_2 FILLER_71_724 ();
 sg13g2_fill_2 FILLER_71_738 ();
 sg13g2_fill_2 FILLER_71_772 ();
 sg13g2_fill_1 FILLER_71_774 ();
 sg13g2_decap_8 FILLER_71_779 ();
 sg13g2_decap_4 FILLER_71_790 ();
 sg13g2_fill_2 FILLER_71_798 ();
 sg13g2_fill_1 FILLER_71_812 ();
 sg13g2_fill_2 FILLER_71_818 ();
 sg13g2_fill_1 FILLER_71_820 ();
 sg13g2_decap_8 FILLER_71_825 ();
 sg13g2_decap_8 FILLER_71_832 ();
 sg13g2_decap_8 FILLER_71_839 ();
 sg13g2_decap_8 FILLER_71_846 ();
 sg13g2_decap_8 FILLER_71_853 ();
 sg13g2_decap_8 FILLER_71_860 ();
 sg13g2_decap_8 FILLER_71_867 ();
 sg13g2_decap_4 FILLER_71_874 ();
 sg13g2_decap_8 FILLER_72_0 ();
 sg13g2_decap_8 FILLER_72_15 ();
 sg13g2_fill_2 FILLER_72_22 ();
 sg13g2_fill_2 FILLER_72_66 ();
 sg13g2_fill_2 FILLER_72_72 ();
 sg13g2_fill_1 FILLER_72_74 ();
 sg13g2_decap_4 FILLER_72_118 ();
 sg13g2_decap_8 FILLER_72_130 ();
 sg13g2_decap_4 FILLER_72_137 ();
 sg13g2_fill_2 FILLER_72_141 ();
 sg13g2_fill_1 FILLER_72_159 ();
 sg13g2_fill_2 FILLER_72_164 ();
 sg13g2_fill_2 FILLER_72_173 ();
 sg13g2_fill_1 FILLER_72_180 ();
 sg13g2_fill_2 FILLER_72_188 ();
 sg13g2_fill_1 FILLER_72_211 ();
 sg13g2_decap_4 FILLER_72_228 ();
 sg13g2_fill_1 FILLER_72_232 ();
 sg13g2_decap_4 FILLER_72_236 ();
 sg13g2_fill_1 FILLER_72_240 ();
 sg13g2_fill_2 FILLER_72_262 ();
 sg13g2_decap_4 FILLER_72_270 ();
 sg13g2_fill_1 FILLER_72_274 ();
 sg13g2_fill_2 FILLER_72_280 ();
 sg13g2_decap_8 FILLER_72_287 ();
 sg13g2_decap_4 FILLER_72_294 ();
 sg13g2_fill_2 FILLER_72_298 ();
 sg13g2_decap_4 FILLER_72_304 ();
 sg13g2_fill_1 FILLER_72_314 ();
 sg13g2_decap_4 FILLER_72_345 ();
 sg13g2_fill_1 FILLER_72_375 ();
 sg13g2_fill_2 FILLER_72_381 ();
 sg13g2_fill_1 FILLER_72_387 ();
 sg13g2_fill_1 FILLER_72_392 ();
 sg13g2_fill_1 FILLER_72_419 ();
 sg13g2_fill_2 FILLER_72_424 ();
 sg13g2_decap_4 FILLER_72_430 ();
 sg13g2_decap_4 FILLER_72_482 ();
 sg13g2_fill_1 FILLER_72_486 ();
 sg13g2_fill_1 FILLER_72_517 ();
 sg13g2_fill_1 FILLER_72_522 ();
 sg13g2_fill_1 FILLER_72_528 ();
 sg13g2_fill_1 FILLER_72_539 ();
 sg13g2_fill_2 FILLER_72_566 ();
 sg13g2_fill_1 FILLER_72_594 ();
 sg13g2_decap_8 FILLER_72_625 ();
 sg13g2_fill_2 FILLER_72_632 ();
 sg13g2_fill_1 FILLER_72_634 ();
 sg13g2_fill_1 FILLER_72_664 ();
 sg13g2_decap_8 FILLER_72_681 ();
 sg13g2_fill_1 FILLER_72_725 ();
 sg13g2_fill_1 FILLER_72_736 ();
 sg13g2_fill_2 FILLER_72_747 ();
 sg13g2_fill_2 FILLER_72_769 ();
 sg13g2_fill_1 FILLER_72_771 ();
 sg13g2_fill_1 FILLER_72_798 ();
 sg13g2_fill_1 FILLER_72_809 ();
 sg13g2_decap_8 FILLER_72_836 ();
 sg13g2_decap_8 FILLER_72_843 ();
 sg13g2_decap_8 FILLER_72_850 ();
 sg13g2_decap_8 FILLER_72_857 ();
 sg13g2_decap_8 FILLER_72_864 ();
 sg13g2_decap_8 FILLER_72_871 ();
 sg13g2_fill_1 FILLER_73_31 ();
 sg13g2_fill_1 FILLER_73_37 ();
 sg13g2_decap_4 FILLER_73_42 ();
 sg13g2_fill_1 FILLER_73_46 ();
 sg13g2_fill_1 FILLER_73_57 ();
 sg13g2_decap_4 FILLER_73_68 ();
 sg13g2_decap_4 FILLER_73_82 ();
 sg13g2_decap_8 FILLER_73_90 ();
 sg13g2_fill_2 FILLER_73_97 ();
 sg13g2_decap_8 FILLER_73_103 ();
 sg13g2_decap_4 FILLER_73_110 ();
 sg13g2_fill_1 FILLER_73_114 ();
 sg13g2_fill_2 FILLER_73_174 ();
 sg13g2_fill_1 FILLER_73_176 ();
 sg13g2_fill_2 FILLER_73_181 ();
 sg13g2_fill_1 FILLER_73_183 ();
 sg13g2_fill_2 FILLER_73_202 ();
 sg13g2_fill_1 FILLER_73_213 ();
 sg13g2_fill_1 FILLER_73_254 ();
 sg13g2_fill_2 FILLER_73_287 ();
 sg13g2_decap_4 FILLER_73_294 ();
 sg13g2_fill_1 FILLER_73_298 ();
 sg13g2_decap_4 FILLER_73_349 ();
 sg13g2_fill_1 FILLER_73_353 ();
 sg13g2_fill_1 FILLER_73_366 ();
 sg13g2_fill_1 FILLER_73_372 ();
 sg13g2_fill_2 FILLER_73_378 ();
 sg13g2_fill_2 FILLER_73_385 ();
 sg13g2_fill_1 FILLER_73_414 ();
 sg13g2_decap_8 FILLER_73_436 ();
 sg13g2_fill_1 FILLER_73_443 ();
 sg13g2_fill_1 FILLER_73_449 ();
 sg13g2_decap_8 FILLER_73_461 ();
 sg13g2_decap_4 FILLER_73_472 ();
 sg13g2_fill_1 FILLER_73_476 ();
 sg13g2_decap_8 FILLER_73_482 ();
 sg13g2_fill_1 FILLER_73_489 ();
 sg13g2_fill_1 FILLER_73_495 ();
 sg13g2_fill_2 FILLER_73_500 ();
 sg13g2_fill_1 FILLER_73_507 ();
 sg13g2_fill_1 FILLER_73_512 ();
 sg13g2_fill_1 FILLER_73_539 ();
 sg13g2_fill_2 FILLER_73_545 ();
 sg13g2_fill_2 FILLER_73_551 ();
 sg13g2_fill_1 FILLER_73_553 ();
 sg13g2_decap_4 FILLER_73_625 ();
 sg13g2_fill_1 FILLER_73_629 ();
 sg13g2_fill_2 FILLER_73_658 ();
 sg13g2_decap_4 FILLER_73_694 ();
 sg13g2_fill_2 FILLER_73_698 ();
 sg13g2_decap_8 FILLER_73_704 ();
 sg13g2_decap_8 FILLER_73_711 ();
 sg13g2_fill_2 FILLER_73_729 ();
 sg13g2_fill_2 FILLER_73_735 ();
 sg13g2_fill_1 FILLER_73_745 ();
 sg13g2_fill_1 FILLER_73_759 ();
 sg13g2_fill_2 FILLER_73_782 ();
 sg13g2_decap_8 FILLER_73_798 ();
 sg13g2_decap_8 FILLER_73_805 ();
 sg13g2_decap_4 FILLER_73_812 ();
 sg13g2_fill_1 FILLER_73_816 ();
 sg13g2_decap_8 FILLER_73_821 ();
 sg13g2_decap_8 FILLER_73_828 ();
 sg13g2_decap_8 FILLER_73_835 ();
 sg13g2_decap_8 FILLER_73_842 ();
 sg13g2_decap_8 FILLER_73_849 ();
 sg13g2_decap_8 FILLER_73_856 ();
 sg13g2_decap_8 FILLER_73_863 ();
 sg13g2_decap_8 FILLER_73_870 ();
 sg13g2_fill_1 FILLER_73_877 ();
 sg13g2_decap_8 FILLER_74_0 ();
 sg13g2_fill_2 FILLER_74_7 ();
 sg13g2_decap_8 FILLER_74_13 ();
 sg13g2_fill_2 FILLER_74_20 ();
 sg13g2_fill_1 FILLER_74_22 ();
 sg13g2_fill_2 FILLER_74_82 ();
 sg13g2_fill_2 FILLER_74_89 ();
 sg13g2_decap_4 FILLER_74_121 ();
 sg13g2_fill_2 FILLER_74_125 ();
 sg13g2_fill_1 FILLER_74_157 ();
 sg13g2_fill_1 FILLER_74_163 ();
 sg13g2_fill_1 FILLER_74_174 ();
 sg13g2_decap_4 FILLER_74_207 ();
 sg13g2_fill_1 FILLER_74_211 ();
 sg13g2_fill_1 FILLER_74_223 ();
 sg13g2_fill_1 FILLER_74_228 ();
 sg13g2_fill_1 FILLER_74_234 ();
 sg13g2_fill_2 FILLER_74_245 ();
 sg13g2_fill_2 FILLER_74_260 ();
 sg13g2_decap_8 FILLER_74_272 ();
 sg13g2_fill_1 FILLER_74_317 ();
 sg13g2_decap_8 FILLER_74_352 ();
 sg13g2_decap_4 FILLER_74_359 ();
 sg13g2_fill_2 FILLER_74_372 ();
 sg13g2_fill_1 FILLER_74_374 ();
 sg13g2_decap_4 FILLER_74_382 ();
 sg13g2_fill_1 FILLER_74_386 ();
 sg13g2_decap_8 FILLER_74_392 ();
 sg13g2_fill_2 FILLER_74_410 ();
 sg13g2_fill_1 FILLER_74_412 ();
 sg13g2_fill_1 FILLER_74_435 ();
 sg13g2_fill_1 FILLER_74_440 ();
 sg13g2_fill_2 FILLER_74_467 ();
 sg13g2_decap_4 FILLER_74_482 ();
 sg13g2_fill_1 FILLER_74_486 ();
 sg13g2_fill_1 FILLER_74_494 ();
 sg13g2_decap_8 FILLER_74_499 ();
 sg13g2_fill_2 FILLER_74_534 ();
 sg13g2_decap_8 FILLER_74_577 ();
 sg13g2_decap_8 FILLER_74_584 ();
 sg13g2_fill_2 FILLER_74_591 ();
 sg13g2_decap_4 FILLER_74_598 ();
 sg13g2_decap_8 FILLER_74_606 ();
 sg13g2_decap_4 FILLER_74_613 ();
 sg13g2_fill_2 FILLER_74_617 ();
 sg13g2_fill_2 FILLER_74_657 ();
 sg13g2_decap_8 FILLER_74_668 ();
 sg13g2_fill_1 FILLER_74_675 ();
 sg13g2_fill_2 FILLER_74_680 ();
 sg13g2_fill_1 FILLER_74_734 ();
 sg13g2_fill_1 FILLER_74_740 ();
 sg13g2_fill_1 FILLER_74_746 ();
 sg13g2_fill_1 FILLER_74_752 ();
 sg13g2_fill_2 FILLER_74_762 ();
 sg13g2_fill_1 FILLER_74_764 ();
 sg13g2_fill_1 FILLER_74_778 ();
 sg13g2_fill_2 FILLER_74_805 ();
 sg13g2_fill_1 FILLER_74_807 ();
 sg13g2_decap_8 FILLER_74_838 ();
 sg13g2_decap_8 FILLER_74_845 ();
 sg13g2_decap_8 FILLER_74_852 ();
 sg13g2_decap_8 FILLER_74_859 ();
 sg13g2_decap_8 FILLER_74_866 ();
 sg13g2_decap_4 FILLER_74_873 ();
 sg13g2_fill_1 FILLER_74_877 ();
 sg13g2_decap_8 FILLER_75_0 ();
 sg13g2_fill_2 FILLER_75_37 ();
 sg13g2_fill_1 FILLER_75_43 ();
 sg13g2_decap_8 FILLER_75_68 ();
 sg13g2_fill_2 FILLER_75_75 ();
 sg13g2_fill_1 FILLER_75_80 ();
 sg13g2_fill_1 FILLER_75_93 ();
 sg13g2_fill_2 FILLER_75_99 ();
 sg13g2_fill_2 FILLER_75_105 ();
 sg13g2_fill_1 FILLER_75_107 ();
 sg13g2_fill_1 FILLER_75_134 ();
 sg13g2_fill_2 FILLER_75_139 ();
 sg13g2_fill_1 FILLER_75_141 ();
 sg13g2_decap_8 FILLER_75_146 ();
 sg13g2_decap_4 FILLER_75_153 ();
 sg13g2_fill_2 FILLER_75_157 ();
 sg13g2_fill_2 FILLER_75_178 ();
 sg13g2_decap_4 FILLER_75_205 ();
 sg13g2_fill_1 FILLER_75_226 ();
 sg13g2_fill_1 FILLER_75_232 ();
 sg13g2_fill_1 FILLER_75_253 ();
 sg13g2_decap_8 FILLER_75_303 ();
 sg13g2_fill_1 FILLER_75_310 ();
 sg13g2_fill_2 FILLER_75_337 ();
 sg13g2_fill_2 FILLER_75_344 ();
 sg13g2_fill_1 FILLER_75_351 ();
 sg13g2_fill_2 FILLER_75_357 ();
 sg13g2_fill_1 FILLER_75_359 ();
 sg13g2_fill_2 FILLER_75_365 ();
 sg13g2_fill_1 FILLER_75_367 ();
 sg13g2_fill_2 FILLER_75_373 ();
 sg13g2_fill_2 FILLER_75_379 ();
 sg13g2_fill_1 FILLER_75_381 ();
 sg13g2_fill_1 FILLER_75_393 ();
 sg13g2_fill_1 FILLER_75_411 ();
 sg13g2_fill_2 FILLER_75_416 ();
 sg13g2_fill_2 FILLER_75_426 ();
 sg13g2_fill_1 FILLER_75_432 ();
 sg13g2_decap_8 FILLER_75_438 ();
 sg13g2_fill_2 FILLER_75_445 ();
 sg13g2_fill_1 FILLER_75_447 ();
 sg13g2_decap_4 FILLER_75_457 ();
 sg13g2_fill_1 FILLER_75_465 ();
 sg13g2_fill_1 FILLER_75_481 ();
 sg13g2_fill_1 FILLER_75_487 ();
 sg13g2_fill_1 FILLER_75_514 ();
 sg13g2_fill_2 FILLER_75_519 ();
 sg13g2_fill_2 FILLER_75_531 ();
 sg13g2_fill_1 FILLER_75_533 ();
 sg13g2_fill_2 FILLER_75_539 ();
 sg13g2_fill_1 FILLER_75_541 ();
 sg13g2_fill_1 FILLER_75_556 ();
 sg13g2_decap_4 FILLER_75_561 ();
 sg13g2_fill_2 FILLER_75_565 ();
 sg13g2_fill_2 FILLER_75_571 ();
 sg13g2_fill_1 FILLER_75_573 ();
 sg13g2_fill_1 FILLER_75_578 ();
 sg13g2_fill_2 FILLER_75_584 ();
 sg13g2_decap_4 FILLER_75_591 ();
 sg13g2_decap_4 FILLER_75_605 ();
 sg13g2_decap_4 FILLER_75_619 ();
 sg13g2_fill_2 FILLER_75_623 ();
 sg13g2_decap_8 FILLER_75_638 ();
 sg13g2_fill_1 FILLER_75_645 ();
 sg13g2_decap_4 FILLER_75_650 ();
 sg13g2_fill_1 FILLER_75_689 ();
 sg13g2_fill_1 FILLER_75_702 ();
 sg13g2_decap_4 FILLER_75_707 ();
 sg13g2_fill_2 FILLER_75_711 ();
 sg13g2_decap_4 FILLER_75_721 ();
 sg13g2_fill_1 FILLER_75_745 ();
 sg13g2_fill_1 FILLER_75_749 ();
 sg13g2_fill_1 FILLER_75_758 ();
 sg13g2_fill_1 FILLER_75_769 ();
 sg13g2_fill_2 FILLER_75_775 ();
 sg13g2_fill_2 FILLER_75_781 ();
 sg13g2_fill_2 FILLER_75_791 ();
 sg13g2_fill_2 FILLER_75_812 ();
 sg13g2_fill_1 FILLER_75_814 ();
 sg13g2_decap_8 FILLER_75_819 ();
 sg13g2_decap_8 FILLER_75_826 ();
 sg13g2_decap_8 FILLER_75_833 ();
 sg13g2_decap_8 FILLER_75_840 ();
 sg13g2_decap_8 FILLER_75_847 ();
 sg13g2_decap_8 FILLER_75_854 ();
 sg13g2_decap_8 FILLER_75_861 ();
 sg13g2_decap_8 FILLER_75_868 ();
 sg13g2_fill_2 FILLER_75_875 ();
 sg13g2_fill_1 FILLER_75_877 ();
 sg13g2_decap_8 FILLER_76_0 ();
 sg13g2_decap_8 FILLER_76_7 ();
 sg13g2_fill_2 FILLER_76_14 ();
 sg13g2_fill_1 FILLER_76_20 ();
 sg13g2_fill_1 FILLER_76_63 ();
 sg13g2_fill_1 FILLER_76_69 ();
 sg13g2_fill_2 FILLER_76_112 ();
 sg13g2_fill_1 FILLER_76_114 ();
 sg13g2_decap_8 FILLER_76_119 ();
 sg13g2_decap_4 FILLER_76_126 ();
 sg13g2_fill_1 FILLER_76_130 ();
 sg13g2_fill_2 FILLER_76_157 ();
 sg13g2_decap_4 FILLER_76_171 ();
 sg13g2_fill_2 FILLER_76_193 ();
 sg13g2_fill_2 FILLER_76_199 ();
 sg13g2_fill_1 FILLER_76_201 ();
 sg13g2_decap_8 FILLER_76_208 ();
 sg13g2_fill_2 FILLER_76_253 ();
 sg13g2_fill_2 FILLER_76_260 ();
 sg13g2_fill_1 FILLER_76_262 ();
 sg13g2_fill_2 FILLER_76_269 ();
 sg13g2_decap_8 FILLER_76_275 ();
 sg13g2_decap_8 FILLER_76_294 ();
 sg13g2_fill_1 FILLER_76_301 ();
 sg13g2_fill_1 FILLER_76_330 ();
 sg13g2_fill_1 FILLER_76_343 ();
 sg13g2_decap_8 FILLER_76_352 ();
 sg13g2_fill_1 FILLER_76_359 ();
 sg13g2_fill_1 FILLER_76_395 ();
 sg13g2_fill_2 FILLER_76_403 ();
 sg13g2_fill_1 FILLER_76_417 ();
 sg13g2_decap_4 FILLER_76_426 ();
 sg13g2_fill_2 FILLER_76_444 ();
 sg13g2_fill_1 FILLER_76_446 ();
 sg13g2_fill_1 FILLER_76_450 ();
 sg13g2_fill_1 FILLER_76_480 ();
 sg13g2_fill_1 FILLER_76_485 ();
 sg13g2_fill_2 FILLER_76_503 ();
 sg13g2_decap_4 FILLER_76_510 ();
 sg13g2_fill_2 FILLER_76_514 ();
 sg13g2_decap_4 FILLER_76_556 ();
 sg13g2_decap_4 FILLER_76_595 ();
 sg13g2_fill_1 FILLER_76_651 ();
 sg13g2_fill_2 FILLER_76_687 ();
 sg13g2_decap_4 FILLER_76_723 ();
 sg13g2_fill_1 FILLER_76_765 ();
 sg13g2_fill_1 FILLER_76_770 ();
 sg13g2_decap_8 FILLER_76_831 ();
 sg13g2_decap_8 FILLER_76_838 ();
 sg13g2_decap_8 FILLER_76_845 ();
 sg13g2_decap_8 FILLER_76_852 ();
 sg13g2_decap_8 FILLER_76_859 ();
 sg13g2_decap_8 FILLER_76_866 ();
 sg13g2_decap_4 FILLER_76_873 ();
 sg13g2_fill_1 FILLER_76_877 ();
 sg13g2_decap_8 FILLER_77_0 ();
 sg13g2_decap_8 FILLER_77_7 ();
 sg13g2_decap_8 FILLER_77_14 ();
 sg13g2_decap_8 FILLER_77_21 ();
 sg13g2_fill_2 FILLER_77_28 ();
 sg13g2_fill_1 FILLER_77_30 ();
 sg13g2_decap_4 FILLER_77_35 ();
 sg13g2_decap_8 FILLER_77_43 ();
 sg13g2_fill_1 FILLER_77_50 ();
 sg13g2_fill_2 FILLER_77_87 ();
 sg13g2_decap_8 FILLER_77_93 ();
 sg13g2_decap_8 FILLER_77_100 ();
 sg13g2_fill_2 FILLER_77_107 ();
 sg13g2_fill_1 FILLER_77_139 ();
 sg13g2_fill_1 FILLER_77_197 ();
 sg13g2_fill_1 FILLER_77_203 ();
 sg13g2_fill_1 FILLER_77_209 ();
 sg13g2_fill_1 FILLER_77_215 ();
 sg13g2_fill_1 FILLER_77_221 ();
 sg13g2_fill_1 FILLER_77_227 ();
 sg13g2_fill_1 FILLER_77_254 ();
 sg13g2_fill_1 FILLER_77_260 ();
 sg13g2_fill_2 FILLER_77_266 ();
 sg13g2_fill_1 FILLER_77_276 ();
 sg13g2_fill_2 FILLER_77_291 ();
 sg13g2_fill_2 FILLER_77_298 ();
 sg13g2_fill_2 FILLER_77_304 ();
 sg13g2_fill_1 FILLER_77_306 ();
 sg13g2_fill_2 FILLER_77_326 ();
 sg13g2_fill_2 FILLER_77_341 ();
 sg13g2_decap_4 FILLER_77_357 ();
 sg13g2_decap_4 FILLER_77_371 ();
 sg13g2_fill_2 FILLER_77_378 ();
 sg13g2_fill_2 FILLER_77_384 ();
 sg13g2_fill_1 FILLER_77_386 ();
 sg13g2_fill_1 FILLER_77_392 ();
 sg13g2_fill_2 FILLER_77_398 ();
 sg13g2_fill_1 FILLER_77_400 ();
 sg13g2_decap_4 FILLER_77_435 ();
 sg13g2_fill_1 FILLER_77_439 ();
 sg13g2_decap_4 FILLER_77_471 ();
 sg13g2_fill_1 FILLER_77_475 ();
 sg13g2_fill_2 FILLER_77_501 ();
 sg13g2_fill_1 FILLER_77_503 ();
 sg13g2_fill_2 FILLER_77_539 ();
 sg13g2_decap_8 FILLER_77_545 ();
 sg13g2_decap_4 FILLER_77_552 ();
 sg13g2_fill_2 FILLER_77_573 ();
 sg13g2_fill_1 FILLER_77_575 ();
 sg13g2_fill_2 FILLER_77_580 ();
 sg13g2_fill_1 FILLER_77_582 ();
 sg13g2_fill_2 FILLER_77_603 ();
 sg13g2_decap_8 FILLER_77_609 ();
 sg13g2_decap_8 FILLER_77_616 ();
 sg13g2_fill_1 FILLER_77_623 ();
 sg13g2_fill_1 FILLER_77_628 ();
 sg13g2_fill_1 FILLER_77_644 ();
 sg13g2_fill_2 FILLER_77_660 ();
 sg13g2_fill_2 FILLER_77_666 ();
 sg13g2_fill_2 FILLER_77_673 ();
 sg13g2_fill_1 FILLER_77_675 ();
 sg13g2_decap_4 FILLER_77_694 ();
 sg13g2_fill_2 FILLER_77_738 ();
 sg13g2_decap_4 FILLER_77_744 ();
 sg13g2_fill_1 FILLER_77_748 ();
 sg13g2_fill_2 FILLER_77_759 ();
 sg13g2_fill_1 FILLER_77_761 ();
 sg13g2_decap_8 FILLER_77_770 ();
 sg13g2_decap_8 FILLER_77_777 ();
 sg13g2_decap_8 FILLER_77_784 ();
 sg13g2_fill_2 FILLER_77_791 ();
 sg13g2_fill_1 FILLER_77_793 ();
 sg13g2_decap_8 FILLER_77_814 ();
 sg13g2_decap_8 FILLER_77_821 ();
 sg13g2_decap_8 FILLER_77_828 ();
 sg13g2_decap_8 FILLER_77_835 ();
 sg13g2_decap_8 FILLER_77_842 ();
 sg13g2_decap_8 FILLER_77_849 ();
 sg13g2_decap_8 FILLER_77_856 ();
 sg13g2_decap_8 FILLER_77_863 ();
 sg13g2_decap_8 FILLER_77_870 ();
 sg13g2_fill_1 FILLER_77_877 ();
 sg13g2_decap_8 FILLER_78_0 ();
 sg13g2_fill_1 FILLER_78_7 ();
 sg13g2_fill_1 FILLER_78_12 ();
 sg13g2_fill_2 FILLER_78_39 ();
 sg13g2_fill_1 FILLER_78_66 ();
 sg13g2_fill_1 FILLER_78_71 ();
 sg13g2_fill_1 FILLER_78_77 ();
 sg13g2_fill_2 FILLER_78_82 ();
 sg13g2_fill_1 FILLER_78_84 ();
 sg13g2_decap_8 FILLER_78_123 ();
 sg13g2_decap_4 FILLER_78_130 ();
 sg13g2_decap_8 FILLER_78_138 ();
 sg13g2_decap_4 FILLER_78_145 ();
 sg13g2_fill_1 FILLER_78_153 ();
 sg13g2_fill_1 FILLER_78_184 ();
 sg13g2_fill_2 FILLER_78_189 ();
 sg13g2_fill_1 FILLER_78_195 ();
 sg13g2_fill_2 FILLER_78_200 ();
 sg13g2_fill_2 FILLER_78_209 ();
 sg13g2_decap_4 FILLER_78_217 ();
 sg13g2_fill_1 FILLER_78_221 ();
 sg13g2_fill_1 FILLER_78_226 ();
 sg13g2_decap_4 FILLER_78_245 ();
 sg13g2_fill_2 FILLER_78_255 ();
 sg13g2_fill_1 FILLER_78_264 ();
 sg13g2_fill_2 FILLER_78_277 ();
 sg13g2_fill_1 FILLER_78_283 ();
 sg13g2_fill_1 FILLER_78_295 ();
 sg13g2_fill_1 FILLER_78_304 ();
 sg13g2_fill_1 FILLER_78_309 ();
 sg13g2_decap_4 FILLER_78_314 ();
 sg13g2_fill_2 FILLER_78_318 ();
 sg13g2_fill_2 FILLER_78_324 ();
 sg13g2_decap_4 FILLER_78_329 ();
 sg13g2_fill_1 FILLER_78_333 ();
 sg13g2_fill_1 FILLER_78_355 ();
 sg13g2_fill_1 FILLER_78_361 ();
 sg13g2_fill_1 FILLER_78_366 ();
 sg13g2_fill_1 FILLER_78_375 ();
 sg13g2_decap_8 FILLER_78_393 ();
 sg13g2_fill_2 FILLER_78_400 ();
 sg13g2_fill_2 FILLER_78_426 ();
 sg13g2_fill_1 FILLER_78_432 ();
 sg13g2_fill_1 FILLER_78_443 ();
 sg13g2_fill_1 FILLER_78_448 ();
 sg13g2_fill_1 FILLER_78_464 ();
 sg13g2_fill_1 FILLER_78_474 ();
 sg13g2_fill_1 FILLER_78_480 ();
 sg13g2_fill_1 FILLER_78_490 ();
 sg13g2_fill_2 FILLER_78_499 ();
 sg13g2_fill_1 FILLER_78_509 ();
 sg13g2_fill_1 FILLER_78_532 ();
 sg13g2_fill_2 FILLER_78_538 ();
 sg13g2_decap_4 FILLER_78_544 ();
 sg13g2_fill_1 FILLER_78_548 ();
 sg13g2_fill_2 FILLER_78_558 ();
 sg13g2_fill_1 FILLER_78_596 ();
 sg13g2_decap_8 FILLER_78_635 ();
 sg13g2_fill_2 FILLER_78_642 ();
 sg13g2_fill_1 FILLER_78_657 ();
 sg13g2_decap_4 FILLER_78_667 ();
 sg13g2_fill_1 FILLER_78_694 ();
 sg13g2_fill_2 FILLER_78_698 ();
 sg13g2_decap_8 FILLER_78_710 ();
 sg13g2_fill_2 FILLER_78_717 ();
 sg13g2_decap_4 FILLER_78_725 ();
 sg13g2_fill_1 FILLER_78_737 ();
 sg13g2_fill_2 FILLER_78_751 ();
 sg13g2_fill_1 FILLER_78_758 ();
 sg13g2_fill_1 FILLER_78_774 ();
 sg13g2_decap_8 FILLER_78_805 ();
 sg13g2_decap_8 FILLER_78_812 ();
 sg13g2_decap_8 FILLER_78_819 ();
 sg13g2_decap_8 FILLER_78_826 ();
 sg13g2_decap_8 FILLER_78_833 ();
 sg13g2_decap_8 FILLER_78_840 ();
 sg13g2_decap_8 FILLER_78_847 ();
 sg13g2_decap_8 FILLER_78_854 ();
 sg13g2_decap_8 FILLER_78_861 ();
 sg13g2_decap_8 FILLER_78_868 ();
 sg13g2_fill_2 FILLER_78_875 ();
 sg13g2_fill_1 FILLER_78_877 ();
 sg13g2_decap_8 FILLER_79_0 ();
 sg13g2_decap_8 FILLER_79_7 ();
 sg13g2_decap_8 FILLER_79_14 ();
 sg13g2_decap_8 FILLER_79_21 ();
 sg13g2_fill_2 FILLER_79_28 ();
 sg13g2_fill_1 FILLER_79_30 ();
 sg13g2_decap_8 FILLER_79_35 ();
 sg13g2_fill_2 FILLER_79_42 ();
 sg13g2_fill_1 FILLER_79_44 ();
 sg13g2_fill_2 FILLER_79_50 ();
 sg13g2_fill_2 FILLER_79_58 ();
 sg13g2_fill_2 FILLER_79_68 ();
 sg13g2_fill_1 FILLER_79_70 ();
 sg13g2_fill_1 FILLER_79_103 ();
 sg13g2_decap_8 FILLER_79_108 ();
 sg13g2_fill_2 FILLER_79_115 ();
 sg13g2_fill_1 FILLER_79_121 ();
 sg13g2_decap_4 FILLER_79_152 ();
 sg13g2_fill_1 FILLER_79_156 ();
 sg13g2_fill_2 FILLER_79_161 ();
 sg13g2_fill_1 FILLER_79_163 ();
 sg13g2_fill_1 FILLER_79_168 ();
 sg13g2_fill_1 FILLER_79_177 ();
 sg13g2_fill_1 FILLER_79_213 ();
 sg13g2_fill_1 FILLER_79_222 ();
 sg13g2_fill_2 FILLER_79_262 ();
 sg13g2_decap_4 FILLER_79_268 ();
 sg13g2_fill_2 FILLER_79_284 ();
 sg13g2_fill_1 FILLER_79_301 ();
 sg13g2_decap_8 FILLER_79_310 ();
 sg13g2_fill_1 FILLER_79_317 ();
 sg13g2_decap_8 FILLER_79_337 ();
 sg13g2_fill_1 FILLER_79_344 ();
 sg13g2_decap_4 FILLER_79_363 ();
 sg13g2_fill_1 FILLER_79_367 ();
 sg13g2_decap_4 FILLER_79_373 ();
 sg13g2_fill_1 FILLER_79_377 ();
 sg13g2_fill_2 FILLER_79_396 ();
 sg13g2_fill_1 FILLER_79_402 ();
 sg13g2_fill_2 FILLER_79_407 ();
 sg13g2_fill_2 FILLER_79_414 ();
 sg13g2_fill_1 FILLER_79_416 ();
 sg13g2_fill_1 FILLER_79_428 ();
 sg13g2_fill_1 FILLER_79_469 ();
 sg13g2_fill_2 FILLER_79_474 ();
 sg13g2_fill_2 FILLER_79_480 ();
 sg13g2_fill_1 FILLER_79_482 ();
 sg13g2_fill_1 FILLER_79_513 ();
 sg13g2_fill_1 FILLER_79_519 ();
 sg13g2_fill_1 FILLER_79_524 ();
 sg13g2_fill_1 FILLER_79_531 ();
 sg13g2_fill_2 FILLER_79_562 ();
 sg13g2_decap_4 FILLER_79_581 ();
 sg13g2_fill_1 FILLER_79_585 ();
 sg13g2_decap_8 FILLER_79_596 ();
 sg13g2_decap_8 FILLER_79_611 ();
 sg13g2_fill_1 FILLER_79_618 ();
 sg13g2_decap_4 FILLER_79_625 ();
 sg13g2_decap_4 FILLER_79_668 ();
 sg13g2_fill_1 FILLER_79_676 ();
 sg13g2_fill_1 FILLER_79_734 ();
 sg13g2_fill_2 FILLER_79_739 ();
 sg13g2_fill_1 FILLER_79_741 ();
 sg13g2_fill_2 FILLER_79_746 ();
 sg13g2_fill_2 FILLER_79_778 ();
 sg13g2_fill_1 FILLER_79_780 ();
 sg13g2_decap_8 FILLER_79_785 ();
 sg13g2_decap_8 FILLER_79_792 ();
 sg13g2_decap_8 FILLER_79_799 ();
 sg13g2_decap_8 FILLER_79_806 ();
 sg13g2_decap_8 FILLER_79_813 ();
 sg13g2_decap_8 FILLER_79_820 ();
 sg13g2_decap_8 FILLER_79_827 ();
 sg13g2_decap_8 FILLER_79_834 ();
 sg13g2_decap_8 FILLER_79_841 ();
 sg13g2_decap_8 FILLER_79_848 ();
 sg13g2_decap_8 FILLER_79_855 ();
 sg13g2_decap_8 FILLER_79_862 ();
 sg13g2_decap_8 FILLER_79_869 ();
 sg13g2_fill_2 FILLER_79_876 ();
 sg13g2_decap_8 FILLER_80_0 ();
 sg13g2_decap_8 FILLER_80_7 ();
 sg13g2_decap_8 FILLER_80_14 ();
 sg13g2_fill_2 FILLER_80_59 ();
 sg13g2_fill_2 FILLER_80_199 ();
 sg13g2_fill_1 FILLER_80_235 ();
 sg13g2_fill_1 FILLER_80_296 ();
 sg13g2_decap_4 FILLER_80_331 ();
 sg13g2_fill_1 FILLER_80_335 ();
 sg13g2_fill_1 FILLER_80_340 ();
 sg13g2_fill_1 FILLER_80_375 ();
 sg13g2_fill_2 FILLER_80_422 ();
 sg13g2_fill_1 FILLER_80_424 ();
 sg13g2_decap_8 FILLER_80_430 ();
 sg13g2_fill_1 FILLER_80_437 ();
 sg13g2_decap_8 FILLER_80_442 ();
 sg13g2_decap_8 FILLER_80_449 ();
 sg13g2_decap_4 FILLER_80_456 ();
 sg13g2_decap_8 FILLER_80_486 ();
 sg13g2_fill_1 FILLER_80_493 ();
 sg13g2_decap_8 FILLER_80_498 ();
 sg13g2_fill_2 FILLER_80_505 ();
 sg13g2_fill_1 FILLER_80_507 ();
 sg13g2_fill_2 FILLER_80_521 ();
 sg13g2_fill_1 FILLER_80_523 ();
 sg13g2_decap_4 FILLER_80_529 ();
 sg13g2_decap_8 FILLER_80_538 ();
 sg13g2_fill_2 FILLER_80_549 ();
 sg13g2_decap_8 FILLER_80_556 ();
 sg13g2_fill_2 FILLER_80_563 ();
 sg13g2_fill_1 FILLER_80_649 ();
 sg13g2_fill_2 FILLER_80_676 ();
 sg13g2_fill_1 FILLER_80_678 ();
 sg13g2_fill_1 FILLER_80_705 ();
 sg13g2_decap_8 FILLER_80_710 ();
 sg13g2_decap_8 FILLER_80_717 ();
 sg13g2_decap_8 FILLER_80_758 ();
 sg13g2_fill_2 FILLER_80_765 ();
 sg13g2_fill_1 FILLER_80_767 ();
 sg13g2_decap_8 FILLER_80_772 ();
 sg13g2_decap_8 FILLER_80_779 ();
 sg13g2_decap_8 FILLER_80_786 ();
 sg13g2_decap_8 FILLER_80_793 ();
 sg13g2_decap_8 FILLER_80_800 ();
 sg13g2_decap_8 FILLER_80_807 ();
 sg13g2_decap_8 FILLER_80_814 ();
 sg13g2_decap_8 FILLER_80_821 ();
 sg13g2_decap_8 FILLER_80_828 ();
 sg13g2_decap_8 FILLER_80_835 ();
 sg13g2_decap_8 FILLER_80_842 ();
 sg13g2_decap_8 FILLER_80_849 ();
 sg13g2_decap_8 FILLER_80_856 ();
 sg13g2_decap_8 FILLER_80_863 ();
 sg13g2_decap_8 FILLER_80_870 ();
 sg13g2_fill_1 FILLER_80_877 ();
endmodule
