module tt_um_vc32_cpu (clk,
    ena,
    rst_n,
    ui_in,
    uio_in,
    uio_oe,
    uio_out,
    uo_out);
 input clk;
 input ena;
 input rst_n;
 input [7:0] ui_in;
 input [7:0] uio_in;
 output [7:0] uio_oe;
 output [7:0] uio_out;
 output [7:0] uo_out;

 wire _00000_;
 wire _00001_;
 wire _00002_;
 wire _00003_;
 wire _00004_;
 wire _00005_;
 wire _00006_;
 wire _00007_;
 wire _00008_;
 wire _00009_;
 wire _00010_;
 wire _00011_;
 wire _00012_;
 wire _00013_;
 wire _00014_;
 wire _00015_;
 wire _00016_;
 wire _00017_;
 wire _00018_;
 wire _00019_;
 wire _00020_;
 wire _00021_;
 wire _00022_;
 wire _00023_;
 wire _00024_;
 wire _00025_;
 wire _00026_;
 wire _00027_;
 wire _00028_;
 wire _00029_;
 wire _00030_;
 wire _00031_;
 wire _00032_;
 wire _00033_;
 wire _00034_;
 wire _00035_;
 wire _00036_;
 wire _00037_;
 wire _00038_;
 wire _00039_;
 wire _00040_;
 wire _00041_;
 wire _00042_;
 wire _00043_;
 wire _00044_;
 wire _00045_;
 wire _00046_;
 wire _00047_;
 wire _00048_;
 wire _00049_;
 wire _00050_;
 wire _00051_;
 wire _00052_;
 wire _00053_;
 wire _00054_;
 wire _00055_;
 wire _00056_;
 wire _00057_;
 wire _00058_;
 wire _00059_;
 wire _00060_;
 wire _00061_;
 wire _00062_;
 wire _00063_;
 wire _00064_;
 wire _00065_;
 wire _00066_;
 wire _00067_;
 wire _00068_;
 wire _00069_;
 wire _00070_;
 wire _00071_;
 wire _00072_;
 wire _00073_;
 wire _00074_;
 wire _00075_;
 wire _00076_;
 wire _00077_;
 wire _00078_;
 wire _00079_;
 wire _00080_;
 wire _00081_;
 wire _00082_;
 wire _00083_;
 wire _00084_;
 wire _00085_;
 wire _00086_;
 wire _00087_;
 wire _00088_;
 wire _00089_;
 wire _00090_;
 wire _00091_;
 wire _00092_;
 wire _00093_;
 wire _00094_;
 wire _00095_;
 wire _00096_;
 wire _00097_;
 wire _00098_;
 wire _00099_;
 wire _00100_;
 wire _00101_;
 wire _00102_;
 wire _00103_;
 wire _00104_;
 wire _00105_;
 wire _00106_;
 wire _00107_;
 wire _00108_;
 wire _00109_;
 wire _00110_;
 wire _00111_;
 wire _00112_;
 wire _00113_;
 wire _00114_;
 wire _00115_;
 wire _00116_;
 wire _00117_;
 wire _00118_;
 wire _00119_;
 wire _00120_;
 wire _00121_;
 wire _00122_;
 wire _00123_;
 wire _00124_;
 wire _00125_;
 wire _00126_;
 wire _00127_;
 wire _00128_;
 wire _00129_;
 wire _00130_;
 wire _00131_;
 wire _00132_;
 wire _00133_;
 wire _00134_;
 wire _00135_;
 wire _00136_;
 wire _00137_;
 wire _00138_;
 wire _00139_;
 wire _00140_;
 wire _00141_;
 wire _00142_;
 wire _00143_;
 wire _00144_;
 wire _00145_;
 wire _00146_;
 wire _00147_;
 wire _00148_;
 wire _00149_;
 wire _00150_;
 wire _00151_;
 wire _00152_;
 wire _00153_;
 wire _00154_;
 wire _00155_;
 wire _00156_;
 wire _00157_;
 wire _00158_;
 wire _00159_;
 wire _00160_;
 wire _00161_;
 wire _00162_;
 wire _00163_;
 wire _00164_;
 wire _00165_;
 wire _00166_;
 wire _00167_;
 wire _00168_;
 wire _00169_;
 wire _00170_;
 wire _00171_;
 wire _00172_;
 wire _00173_;
 wire _00174_;
 wire _00175_;
 wire _00176_;
 wire _00177_;
 wire _00178_;
 wire _00179_;
 wire _00180_;
 wire _00181_;
 wire _00182_;
 wire _00183_;
 wire _00184_;
 wire _00185_;
 wire _00186_;
 wire _00187_;
 wire _00188_;
 wire _00189_;
 wire _00190_;
 wire _00191_;
 wire _00192_;
 wire _00193_;
 wire _00194_;
 wire _00195_;
 wire _00196_;
 wire _00197_;
 wire _00198_;
 wire _00199_;
 wire _00200_;
 wire _00201_;
 wire _00202_;
 wire _00203_;
 wire _00204_;
 wire _00205_;
 wire _00206_;
 wire _00207_;
 wire _00208_;
 wire _00209_;
 wire _00210_;
 wire _00211_;
 wire _00212_;
 wire _00213_;
 wire _00214_;
 wire _00215_;
 wire _00216_;
 wire _00217_;
 wire _00218_;
 wire _00219_;
 wire _00220_;
 wire _00221_;
 wire _00222_;
 wire _00223_;
 wire _00224_;
 wire _00225_;
 wire _00226_;
 wire _00227_;
 wire _00228_;
 wire _00229_;
 wire _00230_;
 wire _00231_;
 wire _00232_;
 wire _00233_;
 wire _00234_;
 wire _00235_;
 wire _00236_;
 wire _00237_;
 wire _00238_;
 wire _00239_;
 wire _00240_;
 wire _00241_;
 wire _00242_;
 wire _00243_;
 wire _00244_;
 wire _00245_;
 wire _00246_;
 wire _00247_;
 wire _00248_;
 wire _00249_;
 wire _00250_;
 wire _00251_;
 wire _00252_;
 wire _00253_;
 wire _00254_;
 wire _00255_;
 wire _00256_;
 wire _00257_;
 wire _00258_;
 wire _00259_;
 wire _00260_;
 wire _00261_;
 wire _00262_;
 wire _00263_;
 wire _00264_;
 wire _00265_;
 wire _00266_;
 wire _00267_;
 wire _00268_;
 wire _00269_;
 wire _00270_;
 wire _00271_;
 wire _00272_;
 wire _00273_;
 wire _00274_;
 wire _00275_;
 wire _00276_;
 wire _00277_;
 wire _00278_;
 wire _00279_;
 wire _00280_;
 wire _00281_;
 wire _00282_;
 wire _00283_;
 wire _00284_;
 wire _00285_;
 wire _00286_;
 wire _00287_;
 wire _00288_;
 wire _00289_;
 wire _00290_;
 wire _00291_;
 wire _00292_;
 wire _00293_;
 wire _00294_;
 wire _00295_;
 wire _00296_;
 wire _00297_;
 wire _00298_;
 wire _00299_;
 wire _00300_;
 wire _00301_;
 wire _00302_;
 wire _00303_;
 wire _00304_;
 wire _00305_;
 wire _00306_;
 wire _00307_;
 wire _00308_;
 wire _00309_;
 wire _00310_;
 wire _00311_;
 wire _00312_;
 wire _00313_;
 wire _00314_;
 wire _00315_;
 wire _00316_;
 wire _00317_;
 wire _00318_;
 wire _00319_;
 wire _00320_;
 wire _00321_;
 wire _00322_;
 wire _00323_;
 wire _00324_;
 wire _00325_;
 wire _00326_;
 wire _00327_;
 wire _00328_;
 wire _00329_;
 wire _00330_;
 wire _00331_;
 wire _00332_;
 wire _00333_;
 wire _00334_;
 wire _00335_;
 wire _00336_;
 wire _00337_;
 wire _00338_;
 wire _00339_;
 wire _00340_;
 wire _00341_;
 wire _00342_;
 wire _00343_;
 wire _00344_;
 wire _00345_;
 wire _00346_;
 wire _00347_;
 wire _00348_;
 wire _00349_;
 wire _00350_;
 wire _00351_;
 wire _00352_;
 wire _00353_;
 wire _00354_;
 wire _00355_;
 wire _00356_;
 wire _00357_;
 wire _00358_;
 wire _00359_;
 wire _00360_;
 wire _00361_;
 wire _00362_;
 wire _00363_;
 wire _00364_;
 wire _00365_;
 wire _00366_;
 wire _00367_;
 wire _00368_;
 wire _00369_;
 wire _00370_;
 wire _00371_;
 wire _00372_;
 wire _00373_;
 wire _00374_;
 wire _00375_;
 wire _00376_;
 wire _00377_;
 wire _00378_;
 wire _00379_;
 wire _00380_;
 wire _00381_;
 wire _00382_;
 wire _00383_;
 wire _00384_;
 wire _00385_;
 wire _00386_;
 wire _00387_;
 wire _00388_;
 wire _00389_;
 wire _00390_;
 wire _00391_;
 wire _00392_;
 wire _00393_;
 wire _00394_;
 wire _00395_;
 wire _00396_;
 wire _00397_;
 wire _00398_;
 wire _00399_;
 wire _00400_;
 wire _00401_;
 wire _00402_;
 wire _00403_;
 wire _00404_;
 wire _00405_;
 wire _00406_;
 wire _00407_;
 wire _00408_;
 wire _00409_;
 wire _00410_;
 wire _00411_;
 wire _00412_;
 wire _00413_;
 wire _00414_;
 wire _00415_;
 wire _00416_;
 wire _00417_;
 wire _00418_;
 wire _00419_;
 wire _00420_;
 wire _00421_;
 wire _00422_;
 wire _00423_;
 wire _00424_;
 wire _00425_;
 wire _00426_;
 wire _00427_;
 wire _00428_;
 wire _00429_;
 wire _00430_;
 wire _00431_;
 wire _00432_;
 wire _00433_;
 wire _00434_;
 wire _00435_;
 wire _00436_;
 wire _00437_;
 wire _00438_;
 wire _00439_;
 wire _00440_;
 wire _00441_;
 wire _00442_;
 wire _00443_;
 wire _00444_;
 wire _00445_;
 wire _00446_;
 wire _00447_;
 wire _00448_;
 wire _00449_;
 wire _00450_;
 wire _00451_;
 wire _00452_;
 wire _00453_;
 wire _00454_;
 wire _00455_;
 wire _00456_;
 wire _00457_;
 wire _00458_;
 wire _00459_;
 wire _00460_;
 wire _00461_;
 wire _00462_;
 wire _00463_;
 wire _00464_;
 wire _00465_;
 wire _00466_;
 wire _00467_;
 wire _00468_;
 wire _00469_;
 wire _00470_;
 wire _00471_;
 wire _00472_;
 wire _00473_;
 wire _00474_;
 wire _00475_;
 wire _00476_;
 wire _00477_;
 wire _00478_;
 wire _00479_;
 wire _00480_;
 wire _00481_;
 wire _00482_;
 wire _00483_;
 wire _00484_;
 wire _00485_;
 wire _00486_;
 wire _00487_;
 wire _00488_;
 wire _00489_;
 wire _00490_;
 wire _00491_;
 wire _00492_;
 wire _00493_;
 wire _00494_;
 wire _00495_;
 wire _00496_;
 wire _00497_;
 wire _00498_;
 wire _00499_;
 wire _00500_;
 wire _00501_;
 wire _00502_;
 wire _00503_;
 wire _00504_;
 wire _00505_;
 wire _00506_;
 wire _00507_;
 wire _00508_;
 wire _00509_;
 wire _00510_;
 wire _00511_;
 wire _00512_;
 wire _00513_;
 wire _00514_;
 wire _00515_;
 wire _00516_;
 wire _00517_;
 wire _00518_;
 wire _00519_;
 wire _00520_;
 wire _00521_;
 wire _00522_;
 wire _00523_;
 wire _00524_;
 wire _00525_;
 wire _00526_;
 wire _00527_;
 wire _00528_;
 wire _00529_;
 wire _00530_;
 wire _00531_;
 wire _00532_;
 wire _00533_;
 wire _00534_;
 wire _00535_;
 wire _00536_;
 wire _00537_;
 wire _00538_;
 wire _00539_;
 wire _00540_;
 wire _00541_;
 wire _00542_;
 wire _00543_;
 wire _00544_;
 wire _00545_;
 wire _00546_;
 wire _00547_;
 wire _00548_;
 wire _00549_;
 wire _00550_;
 wire _00551_;
 wire _00552_;
 wire _00553_;
 wire _00554_;
 wire _00555_;
 wire _00556_;
 wire _00557_;
 wire _00558_;
 wire _00559_;
 wire _00560_;
 wire _00561_;
 wire _00562_;
 wire _00563_;
 wire _00564_;
 wire _00565_;
 wire _00566_;
 wire _00567_;
 wire _00568_;
 wire _00569_;
 wire _00570_;
 wire _00571_;
 wire _00572_;
 wire _00573_;
 wire _00574_;
 wire _00575_;
 wire _00576_;
 wire _00577_;
 wire _00578_;
 wire _00579_;
 wire _00580_;
 wire _00581_;
 wire _00582_;
 wire _00583_;
 wire _00584_;
 wire _00585_;
 wire _00586_;
 wire _00587_;
 wire _00588_;
 wire _00589_;
 wire _00590_;
 wire _00591_;
 wire _00592_;
 wire _00593_;
 wire _00594_;
 wire _00595_;
 wire _00596_;
 wire _00597_;
 wire _00598_;
 wire _00599_;
 wire _00600_;
 wire _00601_;
 wire _00602_;
 wire _00603_;
 wire _00604_;
 wire _00605_;
 wire _00606_;
 wire _00607_;
 wire _00608_;
 wire _00609_;
 wire _00610_;
 wire _00611_;
 wire _00612_;
 wire _00613_;
 wire _00614_;
 wire _00615_;
 wire _00616_;
 wire _00617_;
 wire _00618_;
 wire _00619_;
 wire _00620_;
 wire _00621_;
 wire _00622_;
 wire _00623_;
 wire _00624_;
 wire _00625_;
 wire _00626_;
 wire _00627_;
 wire _00628_;
 wire _00629_;
 wire _00630_;
 wire _00631_;
 wire _00632_;
 wire _00633_;
 wire _00634_;
 wire _00635_;
 wire _00636_;
 wire _00637_;
 wire _00638_;
 wire _00639_;
 wire _00640_;
 wire _00641_;
 wire _00642_;
 wire _00643_;
 wire _00644_;
 wire _00645_;
 wire _00646_;
 wire _00647_;
 wire _00648_;
 wire _00649_;
 wire _00650_;
 wire _00651_;
 wire _00652_;
 wire _00653_;
 wire _00654_;
 wire _00655_;
 wire _00656_;
 wire _00657_;
 wire _00658_;
 wire _00659_;
 wire _00660_;
 wire _00661_;
 wire _00662_;
 wire _00663_;
 wire _00664_;
 wire _00665_;
 wire _00666_;
 wire _00667_;
 wire _00668_;
 wire _00669_;
 wire _00670_;
 wire _00671_;
 wire _00672_;
 wire _00673_;
 wire _00674_;
 wire _00675_;
 wire _00676_;
 wire _00677_;
 wire _00678_;
 wire _00679_;
 wire _00680_;
 wire _00681_;
 wire _00682_;
 wire _00683_;
 wire _00684_;
 wire _00685_;
 wire _00686_;
 wire _00687_;
 wire _00688_;
 wire _00689_;
 wire _00690_;
 wire _00691_;
 wire _00692_;
 wire _00693_;
 wire _00694_;
 wire _00695_;
 wire _00696_;
 wire _00697_;
 wire _00698_;
 wire _00699_;
 wire _00700_;
 wire _00701_;
 wire _00702_;
 wire _00703_;
 wire _00704_;
 wire _00705_;
 wire _00706_;
 wire _00707_;
 wire _00708_;
 wire _00709_;
 wire _00710_;
 wire _00711_;
 wire _00712_;
 wire _00713_;
 wire _00714_;
 wire _00715_;
 wire _00716_;
 wire _00717_;
 wire _00718_;
 wire _00719_;
 wire _00720_;
 wire _00721_;
 wire _00722_;
 wire _00723_;
 wire _00724_;
 wire _00725_;
 wire _00726_;
 wire _00727_;
 wire _00728_;
 wire _00729_;
 wire _00730_;
 wire _00731_;
 wire _00732_;
 wire _00733_;
 wire _00734_;
 wire _00735_;
 wire _00736_;
 wire _00737_;
 wire _00738_;
 wire _00739_;
 wire _00740_;
 wire _00741_;
 wire _00742_;
 wire _00743_;
 wire _00744_;
 wire _00745_;
 wire _00746_;
 wire _00747_;
 wire _00748_;
 wire _00749_;
 wire _00750_;
 wire _00751_;
 wire _00752_;
 wire _00753_;
 wire _00754_;
 wire _00755_;
 wire _00756_;
 wire _00757_;
 wire _00758_;
 wire _00759_;
 wire _00760_;
 wire _00761_;
 wire _00762_;
 wire _00763_;
 wire _00764_;
 wire _00765_;
 wire _00766_;
 wire _00767_;
 wire _00768_;
 wire _00769_;
 wire _00770_;
 wire _00771_;
 wire _00772_;
 wire _00773_;
 wire _00774_;
 wire _00775_;
 wire _00776_;
 wire _00777_;
 wire _00778_;
 wire _00779_;
 wire _00780_;
 wire _00781_;
 wire _00782_;
 wire _00783_;
 wire _00784_;
 wire _00785_;
 wire _00786_;
 wire _00787_;
 wire _00788_;
 wire _00789_;
 wire _00790_;
 wire _00791_;
 wire _00792_;
 wire _00793_;
 wire _00794_;
 wire _00795_;
 wire _00796_;
 wire _00797_;
 wire _00798_;
 wire _00799_;
 wire _00800_;
 wire _00801_;
 wire _00802_;
 wire _00803_;
 wire _00804_;
 wire _00805_;
 wire _00806_;
 wire _00807_;
 wire _00808_;
 wire _00809_;
 wire _00810_;
 wire _00811_;
 wire _00812_;
 wire _00813_;
 wire _00814_;
 wire _00815_;
 wire _00816_;
 wire _00817_;
 wire _00818_;
 wire _00819_;
 wire _00820_;
 wire _00821_;
 wire _00822_;
 wire _00823_;
 wire _00824_;
 wire _00825_;
 wire _00826_;
 wire _00827_;
 wire _00828_;
 wire _00829_;
 wire _00830_;
 wire _00831_;
 wire _00832_;
 wire _00833_;
 wire _00834_;
 wire _00835_;
 wire _00836_;
 wire _00837_;
 wire _00838_;
 wire _00839_;
 wire _00840_;
 wire _00841_;
 wire _00842_;
 wire _00843_;
 wire _00844_;
 wire _00845_;
 wire _00846_;
 wire _00847_;
 wire _00848_;
 wire _00849_;
 wire _00850_;
 wire _00851_;
 wire _00852_;
 wire _00853_;
 wire _00854_;
 wire _00855_;
 wire _00856_;
 wire _00857_;
 wire _00858_;
 wire _00859_;
 wire _00860_;
 wire _00861_;
 wire _00862_;
 wire _00863_;
 wire _00864_;
 wire _00865_;
 wire _00866_;
 wire _00867_;
 wire _00868_;
 wire _00869_;
 wire _00870_;
 wire _00871_;
 wire _00872_;
 wire _00873_;
 wire _00874_;
 wire _00875_;
 wire _00876_;
 wire _00877_;
 wire _00878_;
 wire _00879_;
 wire _00880_;
 wire _00881_;
 wire _00882_;
 wire _00883_;
 wire _00884_;
 wire _00885_;
 wire _00886_;
 wire _00887_;
 wire _00888_;
 wire _00889_;
 wire _00890_;
 wire _00891_;
 wire _00892_;
 wire _00893_;
 wire _00894_;
 wire _00895_;
 wire _00896_;
 wire _00897_;
 wire _00898_;
 wire _00899_;
 wire _00900_;
 wire _00901_;
 wire _00902_;
 wire _00903_;
 wire _00904_;
 wire _00905_;
 wire _00906_;
 wire _00907_;
 wire _00908_;
 wire _00909_;
 wire _00910_;
 wire _00911_;
 wire _00912_;
 wire _00913_;
 wire _00914_;
 wire _00915_;
 wire _00916_;
 wire _00917_;
 wire _00918_;
 wire _00919_;
 wire _00920_;
 wire _00921_;
 wire _00922_;
 wire _00923_;
 wire _00924_;
 wire _00925_;
 wire _00926_;
 wire _00927_;
 wire _00928_;
 wire _00929_;
 wire _00930_;
 wire _00931_;
 wire _00932_;
 wire _00933_;
 wire _00934_;
 wire _00935_;
 wire _00936_;
 wire _00937_;
 wire _00938_;
 wire _00939_;
 wire _00940_;
 wire _00941_;
 wire _00942_;
 wire _00943_;
 wire _00944_;
 wire _00945_;
 wire _00946_;
 wire _00947_;
 wire _00948_;
 wire _00949_;
 wire _00950_;
 wire _00951_;
 wire _00952_;
 wire _00953_;
 wire _00954_;
 wire _00955_;
 wire _00956_;
 wire _00957_;
 wire _00958_;
 wire _00959_;
 wire _00960_;
 wire _00961_;
 wire _00962_;
 wire _00963_;
 wire _00964_;
 wire _00965_;
 wire _00966_;
 wire _00967_;
 wire _00968_;
 wire _00969_;
 wire _00970_;
 wire _00971_;
 wire _00972_;
 wire _00973_;
 wire _00974_;
 wire _00975_;
 wire _00976_;
 wire _00977_;
 wire _00978_;
 wire _00979_;
 wire _00980_;
 wire _00981_;
 wire _00982_;
 wire _00983_;
 wire _00984_;
 wire _00985_;
 wire _00986_;
 wire _00987_;
 wire _00988_;
 wire _00989_;
 wire _00990_;
 wire _00991_;
 wire _00992_;
 wire _00993_;
 wire _00994_;
 wire _00995_;
 wire _00996_;
 wire _00997_;
 wire _00998_;
 wire _00999_;
 wire _01000_;
 wire _01001_;
 wire _01002_;
 wire _01003_;
 wire _01004_;
 wire _01005_;
 wire _01006_;
 wire _01007_;
 wire _01008_;
 wire _01009_;
 wire _01010_;
 wire _01011_;
 wire _01012_;
 wire _01013_;
 wire _01014_;
 wire _01015_;
 wire _01016_;
 wire _01017_;
 wire _01018_;
 wire _01019_;
 wire _01020_;
 wire _01021_;
 wire _01022_;
 wire _01023_;
 wire _01024_;
 wire _01025_;
 wire _01026_;
 wire _01027_;
 wire _01028_;
 wire _01029_;
 wire _01030_;
 wire _01031_;
 wire _01032_;
 wire _01033_;
 wire _01034_;
 wire _01035_;
 wire _01036_;
 wire _01037_;
 wire _01038_;
 wire _01039_;
 wire _01040_;
 wire _01041_;
 wire _01042_;
 wire _01043_;
 wire _01044_;
 wire _01045_;
 wire _01046_;
 wire _01047_;
 wire _01048_;
 wire _01049_;
 wire _01050_;
 wire _01051_;
 wire _01052_;
 wire _01053_;
 wire _01054_;
 wire _01055_;
 wire _01056_;
 wire _01057_;
 wire _01058_;
 wire _01059_;
 wire _01060_;
 wire _01061_;
 wire _01062_;
 wire _01063_;
 wire _01064_;
 wire _01065_;
 wire _01066_;
 wire _01067_;
 wire _01068_;
 wire _01069_;
 wire _01070_;
 wire _01071_;
 wire _01072_;
 wire _01073_;
 wire _01074_;
 wire _01075_;
 wire _01076_;
 wire _01077_;
 wire _01078_;
 wire _01079_;
 wire _01080_;
 wire _01081_;
 wire _01082_;
 wire _01083_;
 wire _01084_;
 wire _01085_;
 wire _01086_;
 wire _01087_;
 wire _01088_;
 wire _01089_;
 wire _01090_;
 wire _01091_;
 wire _01092_;
 wire _01093_;
 wire _01094_;
 wire _01095_;
 wire _01096_;
 wire _01097_;
 wire _01098_;
 wire _01099_;
 wire _01100_;
 wire _01101_;
 wire _01102_;
 wire _01103_;
 wire _01104_;
 wire _01105_;
 wire _01106_;
 wire _01107_;
 wire _01108_;
 wire _01109_;
 wire _01110_;
 wire _01111_;
 wire _01112_;
 wire _01113_;
 wire _01114_;
 wire _01115_;
 wire _01116_;
 wire _01117_;
 wire _01118_;
 wire _01119_;
 wire _01120_;
 wire _01121_;
 wire _01122_;
 wire _01123_;
 wire _01124_;
 wire _01125_;
 wire _01126_;
 wire _01127_;
 wire _01128_;
 wire _01129_;
 wire _01130_;
 wire _01131_;
 wire _01132_;
 wire _01133_;
 wire _01134_;
 wire _01135_;
 wire _01136_;
 wire _01137_;
 wire _01138_;
 wire _01139_;
 wire _01140_;
 wire _01141_;
 wire _01142_;
 wire _01143_;
 wire _01144_;
 wire _01145_;
 wire _01146_;
 wire _01147_;
 wire _01148_;
 wire _01149_;
 wire _01150_;
 wire _01151_;
 wire _01152_;
 wire _01153_;
 wire _01154_;
 wire _01155_;
 wire _01156_;
 wire _01157_;
 wire _01158_;
 wire _01159_;
 wire _01160_;
 wire _01161_;
 wire _01162_;
 wire _01163_;
 wire _01164_;
 wire _01165_;
 wire _01166_;
 wire _01167_;
 wire _01168_;
 wire _01169_;
 wire _01170_;
 wire _01171_;
 wire _01172_;
 wire _01173_;
 wire _01174_;
 wire _01175_;
 wire _01176_;
 wire _01177_;
 wire _01178_;
 wire _01179_;
 wire _01180_;
 wire _01181_;
 wire _01182_;
 wire _01183_;
 wire _01184_;
 wire _01185_;
 wire _01186_;
 wire _01187_;
 wire _01188_;
 wire _01189_;
 wire _01190_;
 wire _01191_;
 wire _01192_;
 wire _01193_;
 wire _01194_;
 wire _01195_;
 wire _01196_;
 wire _01197_;
 wire _01198_;
 wire _01199_;
 wire _01200_;
 wire _01201_;
 wire _01202_;
 wire _01203_;
 wire _01204_;
 wire _01205_;
 wire _01206_;
 wire _01207_;
 wire _01208_;
 wire _01209_;
 wire _01210_;
 wire _01211_;
 wire _01212_;
 wire _01213_;
 wire _01214_;
 wire _01215_;
 wire _01216_;
 wire _01217_;
 wire _01218_;
 wire _01219_;
 wire _01220_;
 wire _01221_;
 wire _01222_;
 wire _01223_;
 wire _01224_;
 wire _01225_;
 wire _01226_;
 wire _01227_;
 wire _01228_;
 wire _01229_;
 wire _01230_;
 wire _01231_;
 wire _01232_;
 wire _01233_;
 wire _01234_;
 wire _01235_;
 wire _01236_;
 wire _01237_;
 wire _01238_;
 wire _01239_;
 wire _01240_;
 wire _01241_;
 wire _01242_;
 wire _01243_;
 wire _01244_;
 wire _01245_;
 wire _01246_;
 wire _01247_;
 wire _01248_;
 wire _01249_;
 wire _01250_;
 wire _01251_;
 wire _01252_;
 wire _01253_;
 wire _01254_;
 wire _01255_;
 wire _01256_;
 wire _01257_;
 wire _01258_;
 wire _01259_;
 wire _01260_;
 wire _01261_;
 wire _01262_;
 wire _01263_;
 wire _01264_;
 wire _01265_;
 wire _01266_;
 wire _01267_;
 wire _01268_;
 wire _01269_;
 wire _01270_;
 wire _01271_;
 wire _01272_;
 wire _01273_;
 wire _01274_;
 wire _01275_;
 wire _01276_;
 wire _01277_;
 wire _01278_;
 wire _01279_;
 wire _01280_;
 wire _01281_;
 wire _01282_;
 wire _01283_;
 wire _01284_;
 wire _01285_;
 wire _01286_;
 wire _01287_;
 wire _01288_;
 wire _01289_;
 wire _01290_;
 wire _01291_;
 wire _01292_;
 wire _01293_;
 wire _01294_;
 wire _01295_;
 wire _01296_;
 wire _01297_;
 wire _01298_;
 wire _01299_;
 wire _01300_;
 wire _01301_;
 wire _01302_;
 wire _01303_;
 wire _01304_;
 wire _01305_;
 wire _01306_;
 wire _01307_;
 wire _01308_;
 wire _01309_;
 wire _01310_;
 wire _01311_;
 wire _01312_;
 wire _01313_;
 wire _01314_;
 wire _01315_;
 wire _01316_;
 wire _01317_;
 wire _01318_;
 wire _01319_;
 wire _01320_;
 wire _01321_;
 wire _01322_;
 wire _01323_;
 wire _01324_;
 wire _01325_;
 wire _01326_;
 wire _01327_;
 wire _01328_;
 wire _01329_;
 wire _01330_;
 wire _01331_;
 wire _01332_;
 wire _01333_;
 wire _01334_;
 wire _01335_;
 wire _01336_;
 wire _01337_;
 wire _01338_;
 wire _01339_;
 wire _01340_;
 wire _01341_;
 wire _01342_;
 wire _01343_;
 wire _01344_;
 wire _01345_;
 wire _01346_;
 wire _01347_;
 wire _01348_;
 wire _01349_;
 wire _01350_;
 wire _01351_;
 wire _01352_;
 wire _01353_;
 wire _01354_;
 wire _01355_;
 wire _01356_;
 wire _01357_;
 wire _01358_;
 wire _01359_;
 wire _01360_;
 wire _01361_;
 wire _01362_;
 wire _01363_;
 wire _01364_;
 wire _01365_;
 wire _01366_;
 wire _01367_;
 wire _01368_;
 wire _01369_;
 wire _01370_;
 wire _01371_;
 wire _01372_;
 wire _01373_;
 wire _01374_;
 wire _01375_;
 wire _01376_;
 wire _01377_;
 wire _01378_;
 wire _01379_;
 wire _01380_;
 wire _01381_;
 wire _01382_;
 wire _01383_;
 wire _01384_;
 wire _01385_;
 wire _01386_;
 wire _01387_;
 wire _01388_;
 wire _01389_;
 wire _01390_;
 wire _01391_;
 wire _01392_;
 wire _01393_;
 wire _01394_;
 wire _01395_;
 wire _01396_;
 wire _01397_;
 wire _01398_;
 wire _01399_;
 wire _01400_;
 wire _01401_;
 wire _01402_;
 wire _01403_;
 wire _01404_;
 wire _01405_;
 wire _01406_;
 wire _01407_;
 wire _01408_;
 wire _01409_;
 wire _01410_;
 wire _01411_;
 wire _01412_;
 wire _01413_;
 wire _01414_;
 wire _01415_;
 wire _01416_;
 wire _01417_;
 wire _01418_;
 wire _01419_;
 wire _01420_;
 wire _01421_;
 wire _01422_;
 wire _01423_;
 wire _01424_;
 wire _01425_;
 wire _01426_;
 wire _01427_;
 wire _01428_;
 wire _01429_;
 wire _01430_;
 wire _01431_;
 wire _01432_;
 wire _01433_;
 wire _01434_;
 wire _01435_;
 wire _01436_;
 wire _01437_;
 wire _01438_;
 wire _01439_;
 wire _01440_;
 wire _01441_;
 wire _01442_;
 wire _01443_;
 wire _01444_;
 wire _01445_;
 wire _01446_;
 wire _01447_;
 wire _01448_;
 wire _01449_;
 wire _01450_;
 wire _01451_;
 wire _01452_;
 wire _01453_;
 wire _01454_;
 wire _01455_;
 wire _01456_;
 wire _01457_;
 wire _01458_;
 wire _01459_;
 wire _01460_;
 wire _01461_;
 wire _01462_;
 wire _01463_;
 wire _01464_;
 wire _01465_;
 wire _01466_;
 wire _01467_;
 wire _01468_;
 wire _01469_;
 wire _01470_;
 wire _01471_;
 wire _01472_;
 wire _01473_;
 wire _01474_;
 wire _01475_;
 wire _01476_;
 wire _01477_;
 wire _01478_;
 wire _01479_;
 wire _01480_;
 wire _01481_;
 wire _01482_;
 wire _01483_;
 wire _01484_;
 wire _01485_;
 wire _01486_;
 wire _01487_;
 wire _01488_;
 wire _01489_;
 wire _01490_;
 wire _01491_;
 wire _01492_;
 wire _01493_;
 wire _01494_;
 wire _01495_;
 wire _01496_;
 wire _01497_;
 wire _01498_;
 wire _01499_;
 wire _01500_;
 wire _01501_;
 wire _01502_;
 wire _01503_;
 wire _01504_;
 wire _01505_;
 wire _01506_;
 wire _01507_;
 wire _01508_;
 wire _01509_;
 wire _01510_;
 wire _01511_;
 wire _01512_;
 wire _01513_;
 wire _01514_;
 wire _01515_;
 wire _01516_;
 wire _01517_;
 wire _01518_;
 wire _01519_;
 wire _01520_;
 wire _01521_;
 wire _01522_;
 wire _01523_;
 wire _01524_;
 wire _01525_;
 wire _01526_;
 wire _01527_;
 wire _01528_;
 wire _01529_;
 wire _01530_;
 wire _01531_;
 wire _01532_;
 wire _01533_;
 wire _01534_;
 wire _01535_;
 wire _01536_;
 wire _01537_;
 wire _01538_;
 wire _01539_;
 wire _01540_;
 wire _01541_;
 wire _01542_;
 wire _01543_;
 wire _01544_;
 wire _01545_;
 wire _01546_;
 wire _01547_;
 wire _01548_;
 wire _01549_;
 wire _01550_;
 wire _01551_;
 wire _01552_;
 wire _01553_;
 wire _01554_;
 wire _01555_;
 wire _01556_;
 wire _01557_;
 wire _01558_;
 wire _01559_;
 wire _01560_;
 wire _01561_;
 wire _01562_;
 wire _01563_;
 wire _01564_;
 wire _01565_;
 wire _01566_;
 wire _01567_;
 wire _01568_;
 wire _01569_;
 wire _01570_;
 wire _01571_;
 wire _01572_;
 wire _01573_;
 wire _01574_;
 wire _01575_;
 wire _01576_;
 wire _01577_;
 wire _01578_;
 wire _01579_;
 wire _01580_;
 wire _01581_;
 wire _01582_;
 wire _01583_;
 wire _01584_;
 wire _01585_;
 wire _01586_;
 wire _01587_;
 wire _01588_;
 wire _01589_;
 wire _01590_;
 wire _01591_;
 wire _01592_;
 wire _01593_;
 wire _01594_;
 wire _01595_;
 wire _01596_;
 wire _01597_;
 wire _01598_;
 wire _01599_;
 wire _01600_;
 wire _01601_;
 wire _01602_;
 wire _01603_;
 wire _01604_;
 wire _01605_;
 wire _01606_;
 wire _01607_;
 wire _01608_;
 wire _01609_;
 wire _01610_;
 wire _01611_;
 wire _01612_;
 wire _01613_;
 wire _01614_;
 wire _01615_;
 wire _01616_;
 wire _01617_;
 wire _01618_;
 wire _01619_;
 wire _01620_;
 wire _01621_;
 wire _01622_;
 wire _01623_;
 wire _01624_;
 wire _01625_;
 wire _01626_;
 wire _01627_;
 wire _01628_;
 wire _01629_;
 wire _01630_;
 wire _01631_;
 wire _01632_;
 wire _01633_;
 wire _01634_;
 wire _01635_;
 wire _01636_;
 wire _01637_;
 wire _01638_;
 wire _01639_;
 wire _01640_;
 wire _01641_;
 wire _01642_;
 wire _01643_;
 wire _01644_;
 wire _01645_;
 wire _01646_;
 wire _01647_;
 wire _01648_;
 wire _01649_;
 wire _01650_;
 wire _01651_;
 wire _01652_;
 wire _01653_;
 wire _01654_;
 wire _01655_;
 wire _01656_;
 wire _01657_;
 wire _01658_;
 wire _01659_;
 wire _01660_;
 wire _01661_;
 wire _01662_;
 wire _01663_;
 wire _01664_;
 wire _01665_;
 wire _01666_;
 wire _01667_;
 wire _01668_;
 wire _01669_;
 wire _01670_;
 wire _01671_;
 wire _01672_;
 wire _01673_;
 wire _01674_;
 wire _01675_;
 wire _01676_;
 wire _01677_;
 wire _01678_;
 wire _01679_;
 wire _01680_;
 wire _01681_;
 wire _01682_;
 wire _01683_;
 wire _01684_;
 wire _01685_;
 wire _01686_;
 wire _01687_;
 wire _01688_;
 wire _01689_;
 wire _01690_;
 wire _01691_;
 wire _01692_;
 wire _01693_;
 wire _01694_;
 wire _01695_;
 wire _01696_;
 wire _01697_;
 wire _01698_;
 wire _01699_;
 wire _01700_;
 wire _01701_;
 wire _01702_;
 wire _01703_;
 wire _01704_;
 wire _01705_;
 wire _01706_;
 wire _01707_;
 wire _01708_;
 wire _01709_;
 wire _01710_;
 wire _01711_;
 wire _01712_;
 wire _01713_;
 wire _01714_;
 wire _01715_;
 wire _01716_;
 wire _01717_;
 wire _01718_;
 wire _01719_;
 wire _01720_;
 wire _01721_;
 wire _01722_;
 wire _01723_;
 wire _01724_;
 wire _01725_;
 wire _01726_;
 wire _01727_;
 wire _01728_;
 wire _01729_;
 wire _01730_;
 wire _01731_;
 wire _01732_;
 wire _01733_;
 wire _01734_;
 wire _01735_;
 wire _01736_;
 wire _01737_;
 wire _01738_;
 wire _01739_;
 wire _01740_;
 wire _01741_;
 wire _01742_;
 wire _01743_;
 wire _01744_;
 wire _01745_;
 wire _01746_;
 wire _01747_;
 wire _01748_;
 wire _01749_;
 wire _01750_;
 wire _01751_;
 wire _01752_;
 wire _01753_;
 wire _01754_;
 wire _01755_;
 wire _01756_;
 wire _01757_;
 wire _01758_;
 wire _01759_;
 wire _01760_;
 wire _01761_;
 wire _01762_;
 wire _01763_;
 wire _01764_;
 wire _01765_;
 wire _01766_;
 wire _01767_;
 wire _01768_;
 wire _01769_;
 wire _01770_;
 wire _01771_;
 wire _01772_;
 wire _01773_;
 wire _01774_;
 wire _01775_;
 wire _01776_;
 wire _01777_;
 wire _01778_;
 wire _01779_;
 wire _01780_;
 wire _01781_;
 wire _01782_;
 wire _01783_;
 wire _01784_;
 wire _01785_;
 wire _01786_;
 wire _01787_;
 wire _01788_;
 wire _01789_;
 wire _01790_;
 wire _01791_;
 wire _01792_;
 wire _01793_;
 wire _01794_;
 wire _01795_;
 wire _01796_;
 wire _01797_;
 wire _01798_;
 wire _01799_;
 wire _01800_;
 wire _01801_;
 wire _01802_;
 wire _01803_;
 wire _01804_;
 wire _01805_;
 wire _01806_;
 wire _01807_;
 wire _01808_;
 wire _01809_;
 wire _01810_;
 wire _01811_;
 wire _01812_;
 wire _01813_;
 wire _01814_;
 wire _01815_;
 wire _01816_;
 wire _01817_;
 wire _01818_;
 wire _01819_;
 wire _01820_;
 wire _01821_;
 wire _01822_;
 wire _01823_;
 wire _01824_;
 wire _01825_;
 wire _01826_;
 wire _01827_;
 wire _01828_;
 wire _01829_;
 wire _01830_;
 wire _01831_;
 wire _01832_;
 wire _01833_;
 wire _01834_;
 wire _01835_;
 wire _01836_;
 wire _01837_;
 wire _01838_;
 wire _01839_;
 wire _01840_;
 wire _01841_;
 wire _01842_;
 wire _01843_;
 wire _01844_;
 wire _01845_;
 wire _01846_;
 wire _01847_;
 wire _01848_;
 wire _01849_;
 wire _01850_;
 wire _01851_;
 wire _01852_;
 wire _01853_;
 wire _01854_;
 wire _01855_;
 wire _01856_;
 wire _01857_;
 wire _01858_;
 wire _01859_;
 wire _01860_;
 wire _01861_;
 wire _01862_;
 wire _01863_;
 wire _01864_;
 wire _01865_;
 wire _01866_;
 wire _01867_;
 wire _01868_;
 wire _01869_;
 wire _01870_;
 wire _01871_;
 wire _01872_;
 wire _01873_;
 wire _01874_;
 wire _01875_;
 wire _01876_;
 wire _01877_;
 wire _01878_;
 wire _01879_;
 wire _01880_;
 wire _01881_;
 wire _01882_;
 wire _01883_;
 wire _01884_;
 wire _01885_;
 wire _01886_;
 wire _01887_;
 wire _01888_;
 wire _01889_;
 wire _01890_;
 wire _01891_;
 wire _01892_;
 wire _01893_;
 wire _01894_;
 wire _01895_;
 wire _01896_;
 wire _01897_;
 wire _01898_;
 wire _01899_;
 wire _01900_;
 wire _01901_;
 wire _01902_;
 wire _01903_;
 wire _01904_;
 wire _01905_;
 wire _01906_;
 wire _01907_;
 wire _01908_;
 wire _01909_;
 wire _01910_;
 wire _01911_;
 wire _01912_;
 wire _01913_;
 wire _01914_;
 wire _01915_;
 wire _01916_;
 wire _01917_;
 wire _01918_;
 wire _01919_;
 wire _01920_;
 wire _01921_;
 wire _01922_;
 wire _01923_;
 wire _01924_;
 wire _01925_;
 wire _01926_;
 wire _01927_;
 wire _01928_;
 wire _01929_;
 wire _01930_;
 wire _01931_;
 wire _01932_;
 wire _01933_;
 wire _01934_;
 wire _01935_;
 wire _01936_;
 wire _01937_;
 wire _01938_;
 wire _01939_;
 wire _01940_;
 wire _01941_;
 wire _01942_;
 wire _01943_;
 wire _01944_;
 wire _01945_;
 wire _01946_;
 wire _01947_;
 wire _01948_;
 wire _01949_;
 wire _01950_;
 wire _01951_;
 wire _01952_;
 wire _01953_;
 wire _01954_;
 wire _01955_;
 wire _01956_;
 wire _01957_;
 wire _01958_;
 wire _01959_;
 wire _01960_;
 wire _01961_;
 wire _01962_;
 wire _01963_;
 wire _01964_;
 wire _01965_;
 wire _01966_;
 wire _01967_;
 wire _01968_;
 wire _01969_;
 wire _01970_;
 wire _01971_;
 wire _01972_;
 wire _01973_;
 wire _01974_;
 wire _01975_;
 wire _01976_;
 wire _01977_;
 wire _01978_;
 wire _01979_;
 wire _01980_;
 wire _01981_;
 wire _01982_;
 wire _01983_;
 wire _01984_;
 wire _01985_;
 wire _01986_;
 wire _01987_;
 wire _01988_;
 wire _01989_;
 wire _01990_;
 wire _01991_;
 wire _01992_;
 wire _01993_;
 wire _01994_;
 wire _01995_;
 wire _01996_;
 wire _01997_;
 wire _01998_;
 wire _01999_;
 wire _02000_;
 wire _02001_;
 wire _02002_;
 wire _02003_;
 wire _02004_;
 wire _02005_;
 wire _02006_;
 wire _02007_;
 wire _02008_;
 wire _02009_;
 wire _02010_;
 wire _02011_;
 wire _02012_;
 wire _02013_;
 wire _02014_;
 wire _02015_;
 wire _02016_;
 wire _02017_;
 wire _02018_;
 wire _02019_;
 wire _02020_;
 wire _02021_;
 wire _02022_;
 wire _02023_;
 wire _02024_;
 wire _02025_;
 wire _02026_;
 wire _02027_;
 wire _02028_;
 wire _02029_;
 wire _02030_;
 wire _02031_;
 wire _02032_;
 wire _02033_;
 wire _02034_;
 wire _02035_;
 wire _02036_;
 wire _02037_;
 wire _02038_;
 wire _02039_;
 wire _02040_;
 wire _02041_;
 wire _02042_;
 wire _02043_;
 wire _02044_;
 wire _02045_;
 wire _02046_;
 wire _02047_;
 wire _02048_;
 wire _02049_;
 wire _02050_;
 wire _02051_;
 wire _02052_;
 wire _02053_;
 wire _02054_;
 wire _02055_;
 wire _02056_;
 wire _02057_;
 wire _02058_;
 wire _02059_;
 wire _02060_;
 wire _02061_;
 wire _02062_;
 wire _02063_;
 wire _02064_;
 wire _02065_;
 wire _02066_;
 wire _02067_;
 wire _02068_;
 wire _02069_;
 wire _02070_;
 wire _02071_;
 wire _02072_;
 wire _02073_;
 wire _02074_;
 wire _02075_;
 wire _02076_;
 wire _02077_;
 wire _02078_;
 wire _02079_;
 wire _02080_;
 wire _02081_;
 wire _02082_;
 wire _02083_;
 wire _02084_;
 wire _02085_;
 wire _02086_;
 wire _02087_;
 wire _02088_;
 wire _02089_;
 wire _02090_;
 wire _02091_;
 wire _02092_;
 wire _02093_;
 wire _02094_;
 wire _02095_;
 wire _02096_;
 wire _02097_;
 wire _02098_;
 wire _02099_;
 wire _02100_;
 wire _02101_;
 wire _02102_;
 wire _02103_;
 wire _02104_;
 wire _02105_;
 wire _02106_;
 wire _02107_;
 wire _02108_;
 wire _02109_;
 wire _02110_;
 wire _02111_;
 wire _02112_;
 wire _02113_;
 wire _02114_;
 wire _02115_;
 wire _02116_;
 wire _02117_;
 wire _02118_;
 wire _02119_;
 wire _02120_;
 wire _02121_;
 wire _02122_;
 wire _02123_;
 wire _02124_;
 wire _02125_;
 wire _02126_;
 wire _02127_;
 wire _02128_;
 wire _02129_;
 wire _02130_;
 wire _02131_;
 wire _02132_;
 wire _02133_;
 wire _02134_;
 wire _02135_;
 wire _02136_;
 wire _02137_;
 wire _02138_;
 wire _02139_;
 wire _02140_;
 wire _02141_;
 wire _02142_;
 wire _02143_;
 wire _02144_;
 wire _02145_;
 wire _02146_;
 wire _02147_;
 wire _02148_;
 wire _02149_;
 wire _02150_;
 wire _02151_;
 wire _02152_;
 wire _02153_;
 wire _02154_;
 wire _02155_;
 wire _02156_;
 wire _02157_;
 wire _02158_;
 wire _02159_;
 wire _02160_;
 wire _02161_;
 wire _02162_;
 wire _02163_;
 wire _02164_;
 wire _02165_;
 wire _02166_;
 wire _02167_;
 wire _02168_;
 wire _02169_;
 wire _02170_;
 wire _02171_;
 wire _02172_;
 wire _02173_;
 wire _02174_;
 wire _02175_;
 wire _02176_;
 wire _02177_;
 wire _02178_;
 wire _02179_;
 wire _02180_;
 wire _02181_;
 wire _02182_;
 wire _02183_;
 wire _02184_;
 wire _02185_;
 wire _02186_;
 wire _02187_;
 wire _02188_;
 wire _02189_;
 wire _02190_;
 wire _02191_;
 wire _02192_;
 wire _02193_;
 wire _02194_;
 wire _02195_;
 wire _02196_;
 wire _02197_;
 wire _02198_;
 wire _02199_;
 wire _02200_;
 wire _02201_;
 wire _02202_;
 wire _02203_;
 wire _02204_;
 wire _02205_;
 wire _02206_;
 wire _02207_;
 wire _02208_;
 wire _02209_;
 wire _02210_;
 wire _02211_;
 wire _02212_;
 wire _02213_;
 wire _02214_;
 wire _02215_;
 wire _02216_;
 wire _02217_;
 wire _02218_;
 wire _02219_;
 wire _02220_;
 wire _02221_;
 wire _02222_;
 wire _02223_;
 wire _02224_;
 wire _02225_;
 wire _02226_;
 wire _02227_;
 wire _02228_;
 wire _02229_;
 wire _02230_;
 wire _02231_;
 wire _02232_;
 wire _02233_;
 wire _02234_;
 wire _02235_;
 wire _02236_;
 wire _02237_;
 wire _02238_;
 wire _02239_;
 wire _02240_;
 wire _02241_;
 wire _02242_;
 wire _02243_;
 wire _02244_;
 wire _02245_;
 wire _02246_;
 wire _02247_;
 wire _02248_;
 wire _02249_;
 wire _02250_;
 wire _02251_;
 wire _02252_;
 wire _02253_;
 wire _02254_;
 wire _02255_;
 wire _02256_;
 wire _02257_;
 wire _02258_;
 wire _02259_;
 wire _02260_;
 wire _02261_;
 wire _02262_;
 wire _02263_;
 wire _02264_;
 wire _02265_;
 wire _02266_;
 wire _02267_;
 wire _02268_;
 wire _02269_;
 wire _02270_;
 wire _02271_;
 wire _02272_;
 wire _02273_;
 wire _02274_;
 wire _02275_;
 wire _02276_;
 wire _02277_;
 wire _02278_;
 wire _02279_;
 wire _02280_;
 wire _02281_;
 wire _02282_;
 wire _02283_;
 wire _02284_;
 wire _02285_;
 wire _02286_;
 wire _02287_;
 wire _02288_;
 wire _02289_;
 wire _02290_;
 wire _02291_;
 wire _02292_;
 wire _02293_;
 wire _02294_;
 wire _02295_;
 wire _02296_;
 wire _02297_;
 wire _02298_;
 wire _02299_;
 wire _02300_;
 wire _02301_;
 wire _02302_;
 wire _02303_;
 wire _02304_;
 wire _02305_;
 wire _02306_;
 wire _02307_;
 wire _02308_;
 wire _02309_;
 wire _02310_;
 wire _02311_;
 wire _02312_;
 wire _02313_;
 wire _02314_;
 wire _02315_;
 wire _02316_;
 wire _02317_;
 wire _02318_;
 wire _02319_;
 wire _02320_;
 wire _02321_;
 wire _02322_;
 wire _02323_;
 wire _02324_;
 wire _02325_;
 wire _02326_;
 wire _02327_;
 wire _02328_;
 wire _02329_;
 wire _02330_;
 wire _02331_;
 wire _02332_;
 wire _02333_;
 wire _02334_;
 wire _02335_;
 wire _02336_;
 wire _02337_;
 wire _02338_;
 wire _02339_;
 wire _02340_;
 wire _02341_;
 wire _02342_;
 wire _02343_;
 wire _02344_;
 wire _02345_;
 wire _02346_;
 wire _02347_;
 wire _02348_;
 wire _02349_;
 wire _02350_;
 wire _02351_;
 wire _02352_;
 wire _02353_;
 wire _02354_;
 wire _02355_;
 wire _02356_;
 wire _02357_;
 wire _02358_;
 wire _02359_;
 wire _02360_;
 wire _02361_;
 wire _02362_;
 wire _02363_;
 wire _02364_;
 wire _02365_;
 wire _02366_;
 wire _02367_;
 wire _02368_;
 wire _02369_;
 wire _02370_;
 wire _02371_;
 wire _02372_;
 wire _02373_;
 wire _02374_;
 wire _02375_;
 wire _02376_;
 wire _02377_;
 wire _02378_;
 wire _02379_;
 wire _02380_;
 wire _02381_;
 wire _02382_;
 wire _02383_;
 wire _02384_;
 wire _02385_;
 wire _02386_;
 wire _02387_;
 wire _02388_;
 wire _02389_;
 wire _02390_;
 wire _02391_;
 wire _02392_;
 wire _02393_;
 wire _02394_;
 wire _02395_;
 wire _02396_;
 wire _02397_;
 wire _02398_;
 wire _02399_;
 wire _02400_;
 wire _02401_;
 wire _02402_;
 wire _02403_;
 wire _02404_;
 wire _02405_;
 wire _02406_;
 wire _02407_;
 wire _02408_;
 wire _02409_;
 wire _02410_;
 wire _02411_;
 wire _02412_;
 wire _02413_;
 wire _02414_;
 wire _02415_;
 wire _02416_;
 wire _02417_;
 wire _02418_;
 wire _02419_;
 wire _02420_;
 wire _02421_;
 wire _02422_;
 wire _02423_;
 wire _02424_;
 wire _02425_;
 wire _02426_;
 wire _02427_;
 wire _02428_;
 wire _02429_;
 wire _02430_;
 wire _02431_;
 wire _02432_;
 wire _02433_;
 wire _02434_;
 wire _02435_;
 wire _02436_;
 wire _02437_;
 wire _02438_;
 wire _02439_;
 wire _02440_;
 wire _02441_;
 wire _02442_;
 wire _02443_;
 wire _02444_;
 wire _02445_;
 wire _02446_;
 wire _02447_;
 wire _02448_;
 wire _02449_;
 wire _02450_;
 wire _02451_;
 wire _02452_;
 wire _02453_;
 wire _02454_;
 wire _02455_;
 wire _02456_;
 wire _02457_;
 wire _02458_;
 wire _02459_;
 wire _02460_;
 wire _02461_;
 wire _02462_;
 wire _02463_;
 wire _02464_;
 wire _02465_;
 wire _02466_;
 wire _02467_;
 wire _02468_;
 wire _02469_;
 wire _02470_;
 wire _02471_;
 wire _02472_;
 wire _02473_;
 wire _02474_;
 wire _02475_;
 wire _02476_;
 wire _02477_;
 wire _02478_;
 wire _02479_;
 wire _02480_;
 wire _02481_;
 wire _02482_;
 wire _02483_;
 wire _02484_;
 wire _02485_;
 wire _02486_;
 wire _02487_;
 wire _02488_;
 wire _02489_;
 wire _02490_;
 wire _02491_;
 wire _02492_;
 wire _02493_;
 wire _02494_;
 wire _02495_;
 wire _02496_;
 wire _02497_;
 wire _02498_;
 wire _02499_;
 wire _02500_;
 wire _02501_;
 wire _02502_;
 wire _02503_;
 wire _02504_;
 wire _02505_;
 wire _02506_;
 wire _02507_;
 wire _02508_;
 wire _02509_;
 wire _02510_;
 wire _02511_;
 wire _02512_;
 wire _02513_;
 wire _02514_;
 wire _02515_;
 wire _02516_;
 wire _02517_;
 wire _02518_;
 wire _02519_;
 wire _02520_;
 wire _02521_;
 wire _02522_;
 wire _02523_;
 wire _02524_;
 wire _02525_;
 wire _02526_;
 wire _02527_;
 wire _02528_;
 wire _02529_;
 wire _02530_;
 wire _02531_;
 wire _02532_;
 wire _02533_;
 wire _02534_;
 wire _02535_;
 wire _02536_;
 wire _02537_;
 wire _02538_;
 wire _02539_;
 wire _02540_;
 wire _02541_;
 wire _02542_;
 wire _02543_;
 wire _02544_;
 wire _02545_;
 wire _02546_;
 wire _02547_;
 wire _02548_;
 wire _02549_;
 wire _02550_;
 wire _02551_;
 wire _02552_;
 wire _02553_;
 wire _02554_;
 wire _02555_;
 wire _02556_;
 wire _02557_;
 wire _02558_;
 wire _02559_;
 wire _02560_;
 wire _02561_;
 wire _02562_;
 wire _02563_;
 wire _02564_;
 wire _02565_;
 wire _02566_;
 wire _02567_;
 wire _02568_;
 wire _02569_;
 wire _02570_;
 wire _02571_;
 wire _02572_;
 wire _02573_;
 wire _02574_;
 wire _02575_;
 wire _02576_;
 wire _02577_;
 wire _02578_;
 wire _02579_;
 wire _02580_;
 wire _02581_;
 wire _02582_;
 wire _02583_;
 wire _02584_;
 wire _02585_;
 wire _02586_;
 wire _02587_;
 wire _02588_;
 wire _02589_;
 wire _02590_;
 wire _02591_;
 wire _02592_;
 wire _02593_;
 wire _02594_;
 wire _02595_;
 wire _02596_;
 wire _02597_;
 wire _02598_;
 wire _02599_;
 wire _02600_;
 wire _02601_;
 wire _02602_;
 wire _02603_;
 wire _02604_;
 wire _02605_;
 wire _02606_;
 wire _02607_;
 wire _02608_;
 wire _02609_;
 wire _02610_;
 wire _02611_;
 wire _02612_;
 wire _02613_;
 wire _02614_;
 wire _02615_;
 wire _02616_;
 wire _02617_;
 wire _02618_;
 wire _02619_;
 wire _02620_;
 wire _02621_;
 wire _02622_;
 wire _02623_;
 wire _02624_;
 wire _02625_;
 wire _02626_;
 wire _02627_;
 wire _02628_;
 wire _02629_;
 wire _02630_;
 wire _02631_;
 wire _02632_;
 wire _02633_;
 wire _02634_;
 wire _02635_;
 wire _02636_;
 wire _02637_;
 wire _02638_;
 wire _02639_;
 wire _02640_;
 wire _02641_;
 wire _02642_;
 wire _02643_;
 wire _02644_;
 wire _02645_;
 wire _02646_;
 wire _02647_;
 wire _02648_;
 wire _02649_;
 wire _02650_;
 wire _02651_;
 wire _02652_;
 wire _02653_;
 wire _02654_;
 wire _02655_;
 wire _02656_;
 wire _02657_;
 wire _02658_;
 wire _02659_;
 wire _02660_;
 wire _02661_;
 wire _02662_;
 wire _02663_;
 wire _02664_;
 wire _02665_;
 wire _02666_;
 wire _02667_;
 wire _02668_;
 wire _02669_;
 wire _02670_;
 wire _02671_;
 wire _02672_;
 wire _02673_;
 wire _02674_;
 wire _02675_;
 wire _02676_;
 wire _02677_;
 wire _02678_;
 wire _02679_;
 wire _02680_;
 wire _02681_;
 wire _02682_;
 wire _02683_;
 wire _02684_;
 wire _02685_;
 wire _02686_;
 wire _02687_;
 wire _02688_;
 wire _02689_;
 wire _02690_;
 wire _02691_;
 wire _02692_;
 wire _02693_;
 wire _02694_;
 wire _02695_;
 wire _02696_;
 wire _02697_;
 wire _02698_;
 wire _02699_;
 wire _02700_;
 wire _02701_;
 wire _02702_;
 wire _02703_;
 wire _02704_;
 wire _02705_;
 wire _02706_;
 wire _02707_;
 wire _02708_;
 wire _02709_;
 wire _02710_;
 wire _02711_;
 wire _02712_;
 wire _02713_;
 wire _02714_;
 wire _02715_;
 wire _02716_;
 wire _02717_;
 wire _02718_;
 wire _02719_;
 wire _02720_;
 wire _02721_;
 wire _02722_;
 wire _02723_;
 wire _02724_;
 wire _02725_;
 wire _02726_;
 wire _02727_;
 wire _02728_;
 wire _02729_;
 wire _02730_;
 wire _02731_;
 wire _02732_;
 wire _02733_;
 wire _02734_;
 wire _02735_;
 wire _02736_;
 wire _02737_;
 wire _02738_;
 wire _02739_;
 wire _02740_;
 wire _02741_;
 wire _02742_;
 wire _02743_;
 wire _02744_;
 wire _02745_;
 wire _02746_;
 wire _02747_;
 wire _02748_;
 wire _02749_;
 wire _02750_;
 wire _02751_;
 wire _02752_;
 wire _02753_;
 wire _02754_;
 wire _02755_;
 wire _02756_;
 wire _02757_;
 wire _02758_;
 wire _02759_;
 wire _02760_;
 wire _02761_;
 wire _02762_;
 wire _02763_;
 wire _02764_;
 wire _02765_;
 wire _02766_;
 wire _02767_;
 wire _02768_;
 wire _02769_;
 wire _02770_;
 wire _02771_;
 wire _02772_;
 wire _02773_;
 wire _02774_;
 wire _02775_;
 wire _02776_;
 wire _02777_;
 wire _02778_;
 wire _02779_;
 wire _02780_;
 wire _02781_;
 wire _02782_;
 wire _02783_;
 wire _02784_;
 wire _02785_;
 wire _02786_;
 wire _02787_;
 wire _02788_;
 wire _02789_;
 wire _02790_;
 wire _02791_;
 wire _02792_;
 wire _02793_;
 wire _02794_;
 wire _02795_;
 wire _02796_;
 wire _02797_;
 wire _02798_;
 wire _02799_;
 wire _02800_;
 wire _02801_;
 wire _02802_;
 wire _02803_;
 wire _02804_;
 wire _02805_;
 wire _02806_;
 wire _02807_;
 wire _02808_;
 wire _02809_;
 wire _02810_;
 wire _02811_;
 wire _02812_;
 wire _02813_;
 wire _02814_;
 wire _02815_;
 wire _02816_;
 wire _02817_;
 wire _02818_;
 wire _02819_;
 wire _02820_;
 wire _02821_;
 wire _02822_;
 wire _02823_;
 wire _02824_;
 wire _02825_;
 wire _02826_;
 wire _02827_;
 wire _02828_;
 wire _02829_;
 wire _02830_;
 wire _02831_;
 wire _02832_;
 wire _02833_;
 wire _02834_;
 wire _02835_;
 wire _02836_;
 wire _02837_;
 wire _02838_;
 wire _02839_;
 wire _02840_;
 wire _02841_;
 wire _02842_;
 wire _02843_;
 wire _02844_;
 wire _02845_;
 wire _02846_;
 wire _02847_;
 wire _02848_;
 wire _02849_;
 wire _02850_;
 wire _02851_;
 wire _02852_;
 wire _02853_;
 wire _02854_;
 wire _02855_;
 wire _02856_;
 wire _02857_;
 wire _02858_;
 wire _02859_;
 wire _02860_;
 wire _02861_;
 wire _02862_;
 wire _02863_;
 wire _02864_;
 wire _02865_;
 wire _02866_;
 wire _02867_;
 wire _02868_;
 wire _02869_;
 wire _02870_;
 wire _02871_;
 wire _02872_;
 wire _02873_;
 wire _02874_;
 wire _02875_;
 wire _02876_;
 wire _02877_;
 wire _02878_;
 wire _02879_;
 wire _02880_;
 wire _02881_;
 wire _02882_;
 wire _02883_;
 wire _02884_;
 wire _02885_;
 wire _02886_;
 wire _02887_;
 wire _02888_;
 wire _02889_;
 wire _02890_;
 wire _02891_;
 wire _02892_;
 wire _02893_;
 wire _02894_;
 wire _02895_;
 wire _02896_;
 wire _02897_;
 wire _02898_;
 wire _02899_;
 wire _02900_;
 wire _02901_;
 wire _02902_;
 wire _02903_;
 wire _02904_;
 wire _02905_;
 wire _02906_;
 wire _02907_;
 wire _02908_;
 wire _02909_;
 wire _02910_;
 wire _02911_;
 wire _02912_;
 wire _02913_;
 wire _02914_;
 wire _02915_;
 wire _02916_;
 wire _02917_;
 wire _02918_;
 wire _02919_;
 wire _02920_;
 wire _02921_;
 wire _02922_;
 wire _02923_;
 wire _02924_;
 wire _02925_;
 wire _02926_;
 wire _02927_;
 wire _02928_;
 wire _02929_;
 wire _02930_;
 wire _02931_;
 wire _02932_;
 wire _02933_;
 wire _02934_;
 wire _02935_;
 wire _02936_;
 wire _02937_;
 wire _02938_;
 wire _02939_;
 wire _02940_;
 wire _02941_;
 wire _02942_;
 wire _02943_;
 wire _02944_;
 wire _02945_;
 wire _02946_;
 wire _02947_;
 wire _02948_;
 wire _02949_;
 wire _02950_;
 wire _02951_;
 wire _02952_;
 wire _02953_;
 wire _02954_;
 wire _02955_;
 wire _02956_;
 wire _02957_;
 wire _02958_;
 wire _02959_;
 wire _02960_;
 wire _02961_;
 wire _02962_;
 wire _02963_;
 wire _02964_;
 wire _02965_;
 wire _02966_;
 wire _02967_;
 wire _02968_;
 wire _02969_;
 wire _02970_;
 wire _02971_;
 wire _02972_;
 wire _02973_;
 wire _02974_;
 wire _02975_;
 wire _02976_;
 wire _02977_;
 wire _02978_;
 wire _02979_;
 wire _02980_;
 wire _02981_;
 wire _02982_;
 wire _02983_;
 wire _02984_;
 wire _02985_;
 wire _02986_;
 wire _02987_;
 wire _02988_;
 wire _02989_;
 wire _02990_;
 wire _02991_;
 wire _02992_;
 wire _02993_;
 wire _02994_;
 wire _02995_;
 wire _02996_;
 wire _02997_;
 wire _02998_;
 wire _02999_;
 wire _03000_;
 wire _03001_;
 wire _03002_;
 wire _03003_;
 wire _03004_;
 wire _03005_;
 wire _03006_;
 wire _03007_;
 wire _03008_;
 wire _03009_;
 wire _03010_;
 wire _03011_;
 wire _03012_;
 wire _03013_;
 wire _03014_;
 wire _03015_;
 wire _03016_;
 wire _03017_;
 wire _03018_;
 wire _03019_;
 wire _03020_;
 wire _03021_;
 wire _03022_;
 wire _03023_;
 wire _03024_;
 wire _03025_;
 wire _03026_;
 wire _03027_;
 wire _03028_;
 wire _03029_;
 wire _03030_;
 wire _03031_;
 wire _03032_;
 wire _03033_;
 wire _03034_;
 wire _03035_;
 wire _03036_;
 wire _03037_;
 wire _03038_;
 wire _03039_;
 wire _03040_;
 wire _03041_;
 wire _03042_;
 wire _03043_;
 wire _03044_;
 wire _03045_;
 wire _03046_;
 wire _03047_;
 wire _03048_;
 wire _03049_;
 wire _03050_;
 wire _03051_;
 wire _03052_;
 wire _03053_;
 wire _03054_;
 wire _03055_;
 wire _03056_;
 wire _03057_;
 wire _03058_;
 wire _03059_;
 wire _03060_;
 wire _03061_;
 wire _03062_;
 wire _03063_;
 wire _03064_;
 wire _03065_;
 wire _03066_;
 wire _03067_;
 wire _03068_;
 wire _03069_;
 wire _03070_;
 wire _03071_;
 wire _03072_;
 wire _03073_;
 wire _03074_;
 wire _03075_;
 wire _03076_;
 wire _03077_;
 wire _03078_;
 wire _03079_;
 wire _03080_;
 wire _03081_;
 wire _03082_;
 wire _03083_;
 wire _03084_;
 wire _03085_;
 wire _03086_;
 wire _03087_;
 wire _03088_;
 wire _03089_;
 wire _03090_;
 wire _03091_;
 wire _03092_;
 wire _03093_;
 wire _03094_;
 wire _03095_;
 wire _03096_;
 wire _03097_;
 wire _03098_;
 wire _03099_;
 wire _03100_;
 wire _03101_;
 wire _03102_;
 wire _03103_;
 wire _03104_;
 wire _03105_;
 wire _03106_;
 wire _03107_;
 wire _03108_;
 wire _03109_;
 wire _03110_;
 wire _03111_;
 wire _03112_;
 wire _03113_;
 wire _03114_;
 wire _03115_;
 wire _03116_;
 wire _03117_;
 wire _03118_;
 wire _03119_;
 wire _03120_;
 wire _03121_;
 wire _03122_;
 wire _03123_;
 wire _03124_;
 wire _03125_;
 wire _03126_;
 wire _03127_;
 wire _03128_;
 wire _03129_;
 wire _03130_;
 wire _03131_;
 wire _03132_;
 wire _03133_;
 wire _03134_;
 wire _03135_;
 wire _03136_;
 wire _03137_;
 wire _03138_;
 wire _03139_;
 wire _03140_;
 wire _03141_;
 wire _03142_;
 wire _03143_;
 wire _03144_;
 wire _03145_;
 wire _03146_;
 wire _03147_;
 wire _03148_;
 wire _03149_;
 wire _03150_;
 wire _03151_;
 wire _03152_;
 wire _03153_;
 wire _03154_;
 wire _03155_;
 wire _03156_;
 wire _03157_;
 wire _03158_;
 wire _03159_;
 wire _03160_;
 wire _03161_;
 wire _03162_;
 wire _03163_;
 wire _03164_;
 wire _03165_;
 wire _03166_;
 wire _03167_;
 wire _03168_;
 wire _03169_;
 wire _03170_;
 wire _03171_;
 wire _03172_;
 wire _03173_;
 wire _03174_;
 wire _03175_;
 wire _03176_;
 wire _03177_;
 wire _03178_;
 wire _03179_;
 wire _03180_;
 wire _03181_;
 wire _03182_;
 wire _03183_;
 wire _03184_;
 wire _03185_;
 wire _03186_;
 wire _03187_;
 wire _03188_;
 wire _03189_;
 wire _03190_;
 wire _03191_;
 wire _03192_;
 wire _03193_;
 wire _03194_;
 wire _03195_;
 wire _03196_;
 wire _03197_;
 wire _03198_;
 wire _03199_;
 wire _03200_;
 wire _03201_;
 wire _03202_;
 wire _03203_;
 wire _03204_;
 wire _03205_;
 wire _03206_;
 wire _03207_;
 wire _03208_;
 wire _03209_;
 wire _03210_;
 wire _03211_;
 wire _03212_;
 wire _03213_;
 wire _03214_;
 wire _03215_;
 wire _03216_;
 wire _03217_;
 wire _03218_;
 wire _03219_;
 wire _03220_;
 wire _03221_;
 wire _03222_;
 wire _03223_;
 wire _03224_;
 wire _03225_;
 wire _03226_;
 wire _03227_;
 wire _03228_;
 wire _03229_;
 wire _03230_;
 wire _03231_;
 wire _03232_;
 wire _03233_;
 wire _03234_;
 wire _03235_;
 wire _03236_;
 wire _03237_;
 wire _03238_;
 wire _03239_;
 wire _03240_;
 wire _03241_;
 wire _03242_;
 wire _03243_;
 wire _03244_;
 wire _03245_;
 wire _03246_;
 wire _03247_;
 wire _03248_;
 wire _03249_;
 wire _03250_;
 wire _03251_;
 wire _03252_;
 wire _03253_;
 wire _03254_;
 wire _03255_;
 wire _03256_;
 wire _03257_;
 wire _03258_;
 wire _03259_;
 wire _03260_;
 wire _03261_;
 wire _03262_;
 wire _03263_;
 wire _03264_;
 wire _03265_;
 wire _03266_;
 wire _03267_;
 wire _03268_;
 wire _03269_;
 wire _03270_;
 wire _03271_;
 wire _03272_;
 wire _03273_;
 wire _03274_;
 wire _03275_;
 wire _03276_;
 wire _03277_;
 wire _03278_;
 wire _03279_;
 wire _03280_;
 wire _03281_;
 wire _03282_;
 wire _03283_;
 wire _03284_;
 wire _03285_;
 wire _03286_;
 wire _03287_;
 wire _03288_;
 wire _03289_;
 wire _03290_;
 wire _03291_;
 wire _03292_;
 wire _03293_;
 wire _03294_;
 wire _03295_;
 wire _03296_;
 wire _03297_;
 wire _03298_;
 wire _03299_;
 wire _03300_;
 wire _03301_;
 wire _03302_;
 wire _03303_;
 wire _03304_;
 wire _03305_;
 wire _03306_;
 wire _03307_;
 wire _03308_;
 wire _03309_;
 wire _03310_;
 wire _03311_;
 wire _03312_;
 wire _03313_;
 wire _03314_;
 wire _03315_;
 wire _03316_;
 wire _03317_;
 wire _03318_;
 wire _03319_;
 wire _03320_;
 wire _03321_;
 wire _03322_;
 wire _03323_;
 wire _03324_;
 wire _03325_;
 wire _03326_;
 wire _03327_;
 wire _03328_;
 wire _03329_;
 wire _03330_;
 wire _03331_;
 wire _03332_;
 wire _03333_;
 wire _03334_;
 wire _03335_;
 wire _03336_;
 wire _03337_;
 wire _03338_;
 wire _03339_;
 wire _03340_;
 wire _03341_;
 wire _03342_;
 wire _03343_;
 wire _03344_;
 wire _03345_;
 wire _03346_;
 wire _03347_;
 wire _03348_;
 wire _03349_;
 wire _03350_;
 wire _03351_;
 wire _03352_;
 wire _03353_;
 wire _03354_;
 wire _03355_;
 wire _03356_;
 wire _03357_;
 wire _03358_;
 wire _03359_;
 wire _03360_;
 wire _03361_;
 wire _03362_;
 wire _03363_;
 wire _03364_;
 wire _03365_;
 wire _03366_;
 wire _03367_;
 wire _03368_;
 wire _03369_;
 wire _03370_;
 wire _03371_;
 wire _03372_;
 wire _03373_;
 wire _03374_;
 wire _03375_;
 wire _03376_;
 wire _03377_;
 wire _03378_;
 wire _03379_;
 wire _03380_;
 wire _03381_;
 wire _03382_;
 wire _03383_;
 wire _03384_;
 wire _03385_;
 wire _03386_;
 wire _03387_;
 wire _03388_;
 wire _03389_;
 wire _03390_;
 wire _03391_;
 wire _03392_;
 wire _03393_;
 wire _03394_;
 wire _03395_;
 wire _03396_;
 wire _03397_;
 wire _03398_;
 wire _03399_;
 wire _03400_;
 wire _03401_;
 wire _03402_;
 wire _03403_;
 wire _03404_;
 wire _03405_;
 wire _03406_;
 wire _03407_;
 wire _03408_;
 wire _03409_;
 wire _03410_;
 wire _03411_;
 wire _03412_;
 wire _03413_;
 wire _03414_;
 wire _03415_;
 wire _03416_;
 wire _03417_;
 wire _03418_;
 wire _03419_;
 wire _03420_;
 wire _03421_;
 wire _03422_;
 wire _03423_;
 wire _03424_;
 wire _03425_;
 wire _03426_;
 wire _03427_;
 wire _03428_;
 wire _03429_;
 wire _03430_;
 wire _03431_;
 wire _03432_;
 wire _03433_;
 wire _03434_;
 wire _03435_;
 wire _03436_;
 wire _03437_;
 wire _03438_;
 wire _03439_;
 wire _03440_;
 wire _03441_;
 wire _03442_;
 wire _03443_;
 wire _03444_;
 wire _03445_;
 wire _03446_;
 wire _03447_;
 wire _03448_;
 wire _03449_;
 wire _03450_;
 wire _03451_;
 wire _03452_;
 wire _03453_;
 wire _03454_;
 wire _03455_;
 wire _03456_;
 wire _03457_;
 wire _03458_;
 wire _03459_;
 wire _03460_;
 wire _03461_;
 wire _03462_;
 wire _03463_;
 wire _03464_;
 wire _03465_;
 wire _03466_;
 wire _03467_;
 wire _03468_;
 wire _03469_;
 wire _03470_;
 wire _03471_;
 wire _03472_;
 wire _03473_;
 wire _03474_;
 wire _03475_;
 wire _03476_;
 wire _03477_;
 wire _03478_;
 wire _03479_;
 wire _03480_;
 wire _03481_;
 wire _03482_;
 wire _03483_;
 wire _03484_;
 wire _03485_;
 wire _03486_;
 wire _03487_;
 wire _03488_;
 wire _03489_;
 wire _03490_;
 wire _03491_;
 wire _03492_;
 wire _03493_;
 wire _03494_;
 wire _03495_;
 wire _03496_;
 wire _03497_;
 wire _03498_;
 wire _03499_;
 wire _03500_;
 wire _03501_;
 wire _03502_;
 wire _03503_;
 wire _03504_;
 wire _03505_;
 wire _03506_;
 wire _03507_;
 wire _03508_;
 wire _03509_;
 wire _03510_;
 wire _03511_;
 wire _03512_;
 wire _03513_;
 wire _03514_;
 wire _03515_;
 wire _03516_;
 wire _03517_;
 wire _03518_;
 wire _03519_;
 wire _03520_;
 wire _03521_;
 wire _03522_;
 wire _03523_;
 wire _03524_;
 wire _03525_;
 wire _03526_;
 wire _03527_;
 wire _03528_;
 wire _03529_;
 wire _03530_;
 wire _03531_;
 wire _03532_;
 wire _03533_;
 wire _03534_;
 wire _03535_;
 wire _03536_;
 wire _03537_;
 wire _03538_;
 wire _03539_;
 wire _03540_;
 wire _03541_;
 wire _03542_;
 wire _03543_;
 wire _03544_;
 wire _03545_;
 wire _03546_;
 wire _03547_;
 wire _03548_;
 wire _03549_;
 wire _03550_;
 wire _03551_;
 wire _03552_;
 wire _03553_;
 wire _03554_;
 wire _03555_;
 wire _03556_;
 wire _03557_;
 wire _03558_;
 wire _03559_;
 wire _03560_;
 wire _03561_;
 wire _03562_;
 wire _03563_;
 wire _03564_;
 wire _03565_;
 wire _03566_;
 wire _03567_;
 wire _03568_;
 wire _03569_;
 wire _03570_;
 wire _03571_;
 wire _03572_;
 wire _03573_;
 wire _03574_;
 wire _03575_;
 wire _03576_;
 wire _03577_;
 wire _03578_;
 wire _03579_;
 wire _03580_;
 wire _03581_;
 wire _03582_;
 wire _03583_;
 wire _03584_;
 wire _03585_;
 wire _03586_;
 wire _03587_;
 wire _03588_;
 wire _03589_;
 wire _03590_;
 wire _03591_;
 wire _03592_;
 wire _03593_;
 wire _03594_;
 wire _03595_;
 wire _03596_;
 wire _03597_;
 wire _03598_;
 wire _03599_;
 wire _03600_;
 wire _03601_;
 wire _03602_;
 wire _03603_;
 wire _03604_;
 wire _03605_;
 wire _03606_;
 wire _03607_;
 wire _03608_;
 wire _03609_;
 wire _03610_;
 wire _03611_;
 wire _03612_;
 wire _03613_;
 wire _03614_;
 wire _03615_;
 wire _03616_;
 wire _03617_;
 wire _03618_;
 wire _03619_;
 wire _03620_;
 wire _03621_;
 wire _03622_;
 wire _03623_;
 wire _03624_;
 wire _03625_;
 wire _03626_;
 wire _03627_;
 wire _03628_;
 wire _03629_;
 wire _03630_;
 wire _03631_;
 wire _03632_;
 wire _03633_;
 wire _03634_;
 wire _03635_;
 wire _03636_;
 wire _03637_;
 wire _03638_;
 wire _03639_;
 wire _03640_;
 wire _03641_;
 wire _03642_;
 wire _03643_;
 wire _03644_;
 wire _03645_;
 wire _03646_;
 wire _03647_;
 wire _03648_;
 wire _03649_;
 wire _03650_;
 wire _03651_;
 wire _03652_;
 wire _03653_;
 wire _03654_;
 wire _03655_;
 wire _03656_;
 wire _03657_;
 wire _03658_;
 wire _03659_;
 wire _03660_;
 wire _03661_;
 wire _03662_;
 wire _03663_;
 wire _03664_;
 wire _03665_;
 wire _03666_;
 wire _03667_;
 wire _03668_;
 wire _03669_;
 wire _03670_;
 wire _03671_;
 wire _03672_;
 wire _03673_;
 wire _03674_;
 wire _03675_;
 wire _03676_;
 wire _03677_;
 wire _03678_;
 wire _03679_;
 wire _03680_;
 wire _03681_;
 wire _03682_;
 wire _03683_;
 wire _03684_;
 wire _03685_;
 wire _03686_;
 wire _03687_;
 wire _03688_;
 wire _03689_;
 wire _03690_;
 wire _03691_;
 wire _03692_;
 wire _03693_;
 wire _03694_;
 wire _03695_;
 wire _03696_;
 wire _03697_;
 wire _03698_;
 wire _03699_;
 wire _03700_;
 wire _03701_;
 wire _03702_;
 wire _03703_;
 wire _03704_;
 wire _03705_;
 wire _03706_;
 wire _03707_;
 wire _03708_;
 wire _03709_;
 wire _03710_;
 wire _03711_;
 wire _03712_;
 wire _03713_;
 wire _03714_;
 wire _03715_;
 wire _03716_;
 wire _03717_;
 wire _03718_;
 wire _03719_;
 wire _03720_;
 wire _03721_;
 wire _03722_;
 wire _03723_;
 wire _03724_;
 wire _03725_;
 wire _03726_;
 wire _03727_;
 wire _03728_;
 wire _03729_;
 wire _03730_;
 wire _03731_;
 wire _03732_;
 wire _03733_;
 wire _03734_;
 wire _03735_;
 wire _03736_;
 wire _03737_;
 wire _03738_;
 wire _03739_;
 wire _03740_;
 wire _03741_;
 wire _03742_;
 wire _03743_;
 wire _03744_;
 wire _03745_;
 wire _03746_;
 wire _03747_;
 wire _03748_;
 wire _03749_;
 wire _03750_;
 wire _03751_;
 wire _03752_;
 wire _03753_;
 wire _03754_;
 wire _03755_;
 wire _03756_;
 wire _03757_;
 wire _03758_;
 wire _03759_;
 wire _03760_;
 wire _03761_;
 wire _03762_;
 wire _03763_;
 wire _03764_;
 wire _03765_;
 wire _03766_;
 wire _03767_;
 wire _03768_;
 wire _03769_;
 wire _03770_;
 wire _03771_;
 wire _03772_;
 wire _03773_;
 wire _03774_;
 wire _03775_;
 wire _03776_;
 wire _03777_;
 wire _03778_;
 wire _03779_;
 wire _03780_;
 wire _03781_;
 wire _03782_;
 wire _03783_;
 wire _03784_;
 wire _03785_;
 wire _03786_;
 wire _03787_;
 wire _03788_;
 wire _03789_;
 wire _03790_;
 wire _03791_;
 wire _03792_;
 wire _03793_;
 wire _03794_;
 wire _03795_;
 wire _03796_;
 wire _03797_;
 wire _03798_;
 wire _03799_;
 wire _03800_;
 wire _03801_;
 wire _03802_;
 wire _03803_;
 wire _03804_;
 wire _03805_;
 wire _03806_;
 wire _03807_;
 wire _03808_;
 wire _03809_;
 wire _03810_;
 wire _03811_;
 wire _03812_;
 wire _03813_;
 wire _03814_;
 wire _03815_;
 wire _03816_;
 wire _03817_;
 wire _03818_;
 wire _03819_;
 wire _03820_;
 wire _03821_;
 wire _03822_;
 wire _03823_;
 wire _03824_;
 wire _03825_;
 wire _03826_;
 wire _03827_;
 wire _03828_;
 wire _03829_;
 wire _03830_;
 wire _03831_;
 wire _03832_;
 wire _03833_;
 wire _03834_;
 wire _03835_;
 wire _03836_;
 wire _03837_;
 wire _03838_;
 wire _03839_;
 wire _03840_;
 wire _03841_;
 wire _03842_;
 wire _03843_;
 wire _03844_;
 wire _03845_;
 wire _03846_;
 wire _03847_;
 wire _03848_;
 wire _03849_;
 wire _03850_;
 wire _03851_;
 wire _03852_;
 wire _03853_;
 wire _03854_;
 wire _03855_;
 wire _03856_;
 wire _03857_;
 wire _03858_;
 wire _03859_;
 wire _03860_;
 wire _03861_;
 wire _03862_;
 wire _03863_;
 wire _03864_;
 wire _03865_;
 wire _03866_;
 wire _03867_;
 wire _03868_;
 wire _03869_;
 wire _03870_;
 wire _03871_;
 wire _03872_;
 wire _03873_;
 wire _03874_;
 wire _03875_;
 wire _03876_;
 wire _03877_;
 wire _03878_;
 wire _03879_;
 wire _03880_;
 wire _03881_;
 wire _03882_;
 wire _03883_;
 wire _03884_;
 wire _03885_;
 wire _03886_;
 wire _03887_;
 wire _03888_;
 wire _03889_;
 wire _03890_;
 wire _03891_;
 wire _03892_;
 wire _03893_;
 wire _03894_;
 wire _03895_;
 wire _03896_;
 wire _03897_;
 wire _03898_;
 wire _03899_;
 wire _03900_;
 wire _03901_;
 wire _03902_;
 wire _03903_;
 wire _03904_;
 wire _03905_;
 wire _03906_;
 wire _03907_;
 wire _03908_;
 wire _03909_;
 wire _03910_;
 wire _03911_;
 wire _03912_;
 wire _03913_;
 wire _03914_;
 wire _03915_;
 wire _03916_;
 wire _03917_;
 wire _03918_;
 wire _03919_;
 wire _03920_;
 wire _03921_;
 wire _03922_;
 wire _03923_;
 wire _03924_;
 wire _03925_;
 wire _03926_;
 wire _03927_;
 wire _03928_;
 wire _03929_;
 wire _03930_;
 wire _03931_;
 wire _03932_;
 wire _03933_;
 wire _03934_;
 wire _03935_;
 wire _03936_;
 wire _03937_;
 wire _03938_;
 wire _03939_;
 wire _03940_;
 wire _03941_;
 wire _03942_;
 wire _03943_;
 wire _03944_;
 wire _03945_;
 wire _03946_;
 wire _03947_;
 wire _03948_;
 wire _03949_;
 wire _03950_;
 wire _03951_;
 wire _03952_;
 wire _03953_;
 wire _03954_;
 wire _03955_;
 wire _03956_;
 wire _03957_;
 wire _03958_;
 wire _03959_;
 wire _03960_;
 wire _03961_;
 wire _03962_;
 wire _03963_;
 wire _03964_;
 wire _03965_;
 wire _03966_;
 wire _03967_;
 wire _03968_;
 wire _03969_;
 wire _03970_;
 wire _03971_;
 wire _03972_;
 wire _03973_;
 wire _03974_;
 wire _03975_;
 wire _03976_;
 wire _03977_;
 wire _03978_;
 wire _03979_;
 wire _03980_;
 wire _03981_;
 wire _03982_;
 wire _03983_;
 wire _03984_;
 wire _03985_;
 wire _03986_;
 wire _03987_;
 wire _03988_;
 wire _03989_;
 wire _03990_;
 wire _03991_;
 wire _03992_;
 wire _03993_;
 wire _03994_;
 wire _03995_;
 wire _03996_;
 wire _03997_;
 wire _03998_;
 wire _03999_;
 wire _04000_;
 wire _04001_;
 wire _04002_;
 wire _04003_;
 wire _04004_;
 wire _04005_;
 wire _04006_;
 wire _04007_;
 wire _04008_;
 wire _04009_;
 wire _04010_;
 wire _04011_;
 wire _04012_;
 wire _04013_;
 wire _04014_;
 wire _04015_;
 wire _04016_;
 wire _04017_;
 wire _04018_;
 wire _04019_;
 wire _04020_;
 wire _04021_;
 wire _04022_;
 wire _04023_;
 wire _04024_;
 wire _04025_;
 wire _04026_;
 wire _04027_;
 wire _04028_;
 wire _04029_;
 wire _04030_;
 wire _04031_;
 wire _04032_;
 wire _04033_;
 wire _04034_;
 wire _04035_;
 wire _04036_;
 wire _04037_;
 wire _04038_;
 wire _04039_;
 wire _04040_;
 wire _04041_;
 wire _04042_;
 wire _04043_;
 wire _04044_;
 wire _04045_;
 wire _04046_;
 wire _04047_;
 wire _04048_;
 wire _04049_;
 wire _04050_;
 wire _04051_;
 wire _04052_;
 wire _04053_;
 wire _04054_;
 wire _04055_;
 wire _04056_;
 wire _04057_;
 wire _04058_;
 wire _04059_;
 wire _04060_;
 wire _04061_;
 wire _04062_;
 wire _04063_;
 wire _04064_;
 wire _04065_;
 wire _04066_;
 wire _04067_;
 wire _04068_;
 wire _04069_;
 wire _04070_;
 wire _04071_;
 wire _04072_;
 wire _04073_;
 wire _04074_;
 wire _04075_;
 wire _04076_;
 wire _04077_;
 wire _04078_;
 wire _04079_;
 wire _04080_;
 wire _04081_;
 wire _04082_;
 wire _04083_;
 wire _04084_;
 wire _04085_;
 wire _04086_;
 wire _04087_;
 wire _04088_;
 wire _04089_;
 wire _04090_;
 wire _04091_;
 wire _04092_;
 wire _04093_;
 wire _04094_;
 wire _04095_;
 wire _04096_;
 wire _04097_;
 wire _04098_;
 wire _04099_;
 wire _04100_;
 wire _04101_;
 wire _04102_;
 wire _04103_;
 wire _04104_;
 wire _04105_;
 wire _04106_;
 wire _04107_;
 wire _04108_;
 wire _04109_;
 wire _04110_;
 wire _04111_;
 wire _04112_;
 wire _04113_;
 wire _04114_;
 wire _04115_;
 wire _04116_;
 wire _04117_;
 wire _04118_;
 wire _04119_;
 wire _04120_;
 wire _04121_;
 wire _04122_;
 wire _04123_;
 wire _04124_;
 wire _04125_;
 wire _04126_;
 wire _04127_;
 wire _04128_;
 wire _04129_;
 wire _04130_;
 wire _04131_;
 wire _04132_;
 wire _04133_;
 wire _04134_;
 wire _04135_;
 wire _04136_;
 wire _04137_;
 wire _04138_;
 wire _04139_;
 wire _04140_;
 wire _04141_;
 wire _04142_;
 wire _04143_;
 wire _04144_;
 wire _04145_;
 wire _04146_;
 wire _04147_;
 wire _04148_;
 wire _04149_;
 wire _04150_;
 wire _04151_;
 wire _04152_;
 wire _04153_;
 wire _04154_;
 wire _04155_;
 wire _04156_;
 wire _04157_;
 wire _04158_;
 wire _04159_;
 wire _04160_;
 wire _04161_;
 wire _04162_;
 wire _04163_;
 wire _04164_;
 wire _04165_;
 wire _04166_;
 wire _04167_;
 wire _04168_;
 wire _04169_;
 wire _04170_;
 wire _04171_;
 wire _04172_;
 wire _04173_;
 wire _04174_;
 wire _04175_;
 wire _04176_;
 wire _04177_;
 wire _04178_;
 wire _04179_;
 wire _04180_;
 wire _04181_;
 wire _04182_;
 wire _04183_;
 wire _04184_;
 wire _04185_;
 wire _04186_;
 wire _04187_;
 wire _04188_;
 wire _04189_;
 wire _04190_;
 wire _04191_;
 wire _04192_;
 wire _04193_;
 wire _04194_;
 wire _04195_;
 wire _04196_;
 wire _04197_;
 wire _04198_;
 wire _04199_;
 wire _04200_;
 wire _04201_;
 wire _04202_;
 wire _04203_;
 wire _04204_;
 wire _04205_;
 wire _04206_;
 wire _04207_;
 wire _04208_;
 wire _04209_;
 wire _04210_;
 wire _04211_;
 wire _04212_;
 wire _04213_;
 wire _04214_;
 wire _04215_;
 wire _04216_;
 wire _04217_;
 wire _04218_;
 wire _04219_;
 wire _04220_;
 wire _04221_;
 wire _04222_;
 wire _04223_;
 wire _04224_;
 wire _04225_;
 wire _04226_;
 wire _04227_;
 wire _04228_;
 wire _04229_;
 wire _04230_;
 wire _04231_;
 wire _04232_;
 wire _04233_;
 wire _04234_;
 wire _04235_;
 wire _04236_;
 wire _04237_;
 wire _04238_;
 wire _04239_;
 wire _04240_;
 wire _04241_;
 wire _04242_;
 wire _04243_;
 wire _04244_;
 wire _04245_;
 wire _04246_;
 wire _04247_;
 wire _04248_;
 wire _04249_;
 wire _04250_;
 wire _04251_;
 wire _04252_;
 wire _04253_;
 wire _04254_;
 wire _04255_;
 wire _04256_;
 wire _04257_;
 wire _04258_;
 wire _04259_;
 wire _04260_;
 wire _04261_;
 wire _04262_;
 wire _04263_;
 wire _04264_;
 wire _04265_;
 wire _04266_;
 wire _04267_;
 wire _04268_;
 wire _04269_;
 wire _04270_;
 wire _04271_;
 wire _04272_;
 wire _04273_;
 wire _04274_;
 wire _04275_;
 wire _04276_;
 wire _04277_;
 wire _04278_;
 wire _04279_;
 wire _04280_;
 wire _04281_;
 wire _04282_;
 wire _04283_;
 wire _04284_;
 wire _04285_;
 wire _04286_;
 wire _04287_;
 wire _04288_;
 wire _04289_;
 wire _04290_;
 wire _04291_;
 wire _04292_;
 wire _04293_;
 wire _04294_;
 wire _04295_;
 wire _04296_;
 wire _04297_;
 wire _04298_;
 wire _04299_;
 wire _04300_;
 wire _04301_;
 wire _04302_;
 wire _04303_;
 wire _04304_;
 wire _04305_;
 wire _04306_;
 wire _04307_;
 wire _04308_;
 wire _04309_;
 wire _04310_;
 wire _04311_;
 wire _04312_;
 wire _04313_;
 wire _04314_;
 wire _04315_;
 wire _04316_;
 wire _04317_;
 wire _04318_;
 wire _04319_;
 wire _04320_;
 wire _04321_;
 wire _04322_;
 wire _04323_;
 wire _04324_;
 wire _04325_;
 wire _04326_;
 wire _04327_;
 wire _04328_;
 wire _04329_;
 wire _04330_;
 wire _04331_;
 wire _04332_;
 wire _04333_;
 wire _04334_;
 wire _04335_;
 wire _04336_;
 wire _04337_;
 wire _04338_;
 wire _04339_;
 wire _04340_;
 wire _04341_;
 wire _04342_;
 wire _04343_;
 wire _04344_;
 wire _04345_;
 wire _04346_;
 wire _04347_;
 wire _04348_;
 wire _04349_;
 wire _04350_;
 wire _04351_;
 wire _04352_;
 wire _04353_;
 wire _04354_;
 wire _04355_;
 wire _04356_;
 wire _04357_;
 wire _04358_;
 wire _04359_;
 wire _04360_;
 wire _04361_;
 wire _04362_;
 wire _04363_;
 wire _04364_;
 wire _04365_;
 wire _04366_;
 wire _04367_;
 wire _04368_;
 wire _04369_;
 wire _04370_;
 wire _04371_;
 wire _04372_;
 wire _04373_;
 wire _04374_;
 wire _04375_;
 wire _04376_;
 wire _04377_;
 wire _04378_;
 wire _04379_;
 wire _04380_;
 wire _04381_;
 wire _04382_;
 wire _04383_;
 wire _04384_;
 wire _04385_;
 wire _04386_;
 wire _04387_;
 wire _04388_;
 wire _04389_;
 wire _04390_;
 wire _04391_;
 wire _04392_;
 wire _04393_;
 wire _04394_;
 wire _04395_;
 wire _04396_;
 wire _04397_;
 wire _04398_;
 wire _04399_;
 wire _04400_;
 wire _04401_;
 wire _04402_;
 wire _04403_;
 wire _04404_;
 wire _04405_;
 wire _04406_;
 wire _04407_;
 wire _04408_;
 wire _04409_;
 wire _04410_;
 wire _04411_;
 wire _04412_;
 wire _04413_;
 wire _04414_;
 wire _04415_;
 wire _04416_;
 wire _04417_;
 wire _04418_;
 wire _04419_;
 wire _04420_;
 wire _04421_;
 wire _04422_;
 wire _04423_;
 wire _04424_;
 wire _04425_;
 wire _04426_;
 wire _04427_;
 wire _04428_;
 wire _04429_;
 wire _04430_;
 wire _04431_;
 wire _04432_;
 wire _04433_;
 wire _04434_;
 wire _04435_;
 wire _04436_;
 wire _04437_;
 wire _04438_;
 wire _04439_;
 wire _04440_;
 wire _04441_;
 wire _04442_;
 wire _04443_;
 wire _04444_;
 wire _04445_;
 wire _04446_;
 wire _04447_;
 wire _04448_;
 wire _04449_;
 wire _04450_;
 wire _04451_;
 wire _04452_;
 wire _04453_;
 wire _04454_;
 wire _04455_;
 wire _04456_;
 wire _04457_;
 wire _04458_;
 wire _04459_;
 wire _04460_;
 wire _04461_;
 wire _04462_;
 wire _04463_;
 wire _04464_;
 wire _04465_;
 wire _04466_;
 wire _04467_;
 wire _04468_;
 wire _04469_;
 wire _04470_;
 wire _04471_;
 wire _04472_;
 wire _04473_;
 wire _04474_;
 wire _04475_;
 wire _04476_;
 wire _04477_;
 wire _04478_;
 wire _04479_;
 wire _04480_;
 wire _04481_;
 wire _04482_;
 wire _04483_;
 wire _04484_;
 wire _04485_;
 wire _04486_;
 wire _04487_;
 wire _04488_;
 wire _04489_;
 wire _04490_;
 wire _04491_;
 wire _04492_;
 wire _04493_;
 wire _04494_;
 wire _04495_;
 wire _04496_;
 wire _04497_;
 wire _04498_;
 wire _04499_;
 wire _04500_;
 wire _04501_;
 wire _04502_;
 wire _04503_;
 wire _04504_;
 wire _04505_;
 wire _04506_;
 wire _04507_;
 wire _04508_;
 wire _04509_;
 wire _04510_;
 wire _04511_;
 wire _04512_;
 wire _04513_;
 wire _04514_;
 wire _04515_;
 wire _04516_;
 wire _04517_;
 wire _04518_;
 wire _04519_;
 wire _04520_;
 wire _04521_;
 wire _04522_;
 wire _04523_;
 wire _04524_;
 wire _04525_;
 wire _04526_;
 wire _04527_;
 wire _04528_;
 wire _04529_;
 wire _04530_;
 wire _04531_;
 wire _04532_;
 wire _04533_;
 wire _04534_;
 wire _04535_;
 wire _04536_;
 wire _04537_;
 wire _04538_;
 wire _04539_;
 wire _04540_;
 wire _04541_;
 wire _04542_;
 wire _04543_;
 wire _04544_;
 wire _04545_;
 wire _04546_;
 wire _04547_;
 wire _04548_;
 wire _04549_;
 wire _04550_;
 wire _04551_;
 wire _04552_;
 wire _04553_;
 wire _04554_;
 wire _04555_;
 wire _04556_;
 wire _04557_;
 wire _04558_;
 wire _04559_;
 wire _04560_;
 wire _04561_;
 wire _04562_;
 wire _04563_;
 wire _04564_;
 wire _04565_;
 wire _04566_;
 wire _04567_;
 wire _04568_;
 wire _04569_;
 wire _04570_;
 wire _04571_;
 wire _04572_;
 wire _04573_;
 wire _04574_;
 wire _04575_;
 wire _04576_;
 wire _04577_;
 wire _04578_;
 wire _04579_;
 wire _04580_;
 wire _04581_;
 wire _04582_;
 wire _04583_;
 wire _04584_;
 wire _04585_;
 wire _04586_;
 wire _04587_;
 wire _04588_;
 wire _04589_;
 wire _04590_;
 wire _04591_;
 wire _04592_;
 wire _04593_;
 wire _04594_;
 wire _04595_;
 wire _04596_;
 wire _04597_;
 wire _04598_;
 wire _04599_;
 wire _04600_;
 wire _04601_;
 wire _04602_;
 wire _04603_;
 wire _04604_;
 wire _04605_;
 wire _04606_;
 wire _04607_;
 wire _04608_;
 wire _04609_;
 wire _04610_;
 wire _04611_;
 wire _04612_;
 wire _04613_;
 wire _04614_;
 wire _04615_;
 wire _04616_;
 wire _04617_;
 wire _04618_;
 wire _04619_;
 wire _04620_;
 wire _04621_;
 wire _04622_;
 wire _04623_;
 wire _04624_;
 wire _04625_;
 wire _04626_;
 wire _04627_;
 wire _04628_;
 wire _04629_;
 wire _04630_;
 wire _04631_;
 wire _04632_;
 wire _04633_;
 wire _04634_;
 wire _04635_;
 wire _04636_;
 wire _04637_;
 wire _04638_;
 wire _04639_;
 wire _04640_;
 wire _04641_;
 wire _04642_;
 wire _04643_;
 wire _04644_;
 wire _04645_;
 wire _04646_;
 wire _04647_;
 wire _04648_;
 wire _04649_;
 wire _04650_;
 wire _04651_;
 wire _04652_;
 wire _04653_;
 wire _04654_;
 wire _04655_;
 wire _04656_;
 wire _04657_;
 wire _04658_;
 wire _04659_;
 wire _04660_;
 wire _04661_;
 wire _04662_;
 wire _04663_;
 wire _04664_;
 wire _04665_;
 wire _04666_;
 wire _04667_;
 wire _04668_;
 wire _04669_;
 wire _04670_;
 wire _04671_;
 wire _04672_;
 wire _04673_;
 wire _04674_;
 wire _04675_;
 wire _04676_;
 wire _04677_;
 wire _04678_;
 wire _04679_;
 wire _04680_;
 wire _04681_;
 wire _04682_;
 wire _04683_;
 wire _04684_;
 wire _04685_;
 wire _04686_;
 wire _04687_;
 wire _04688_;
 wire _04689_;
 wire _04690_;
 wire _04691_;
 wire _04692_;
 wire _04693_;
 wire _04694_;
 wire _04695_;
 wire _04696_;
 wire _04697_;
 wire _04698_;
 wire _04699_;
 wire _04700_;
 wire _04701_;
 wire _04702_;
 wire _04703_;
 wire _04704_;
 wire _04705_;
 wire _04706_;
 wire _04707_;
 wire _04708_;
 wire _04709_;
 wire _04710_;
 wire _04711_;
 wire _04712_;
 wire _04713_;
 wire _04714_;
 wire _04715_;
 wire _04716_;
 wire _04717_;
 wire _04718_;
 wire _04719_;
 wire _04720_;
 wire _04721_;
 wire _04722_;
 wire _04723_;
 wire _04724_;
 wire _04725_;
 wire _04726_;
 wire _04727_;
 wire _04728_;
 wire _04729_;
 wire _04730_;
 wire _04731_;
 wire _04732_;
 wire _04733_;
 wire _04734_;
 wire _04735_;
 wire _04736_;
 wire _04737_;
 wire _04738_;
 wire _04739_;
 wire _04740_;
 wire _04741_;
 wire _04742_;
 wire _04743_;
 wire _04744_;
 wire _04745_;
 wire _04746_;
 wire _04747_;
 wire _04748_;
 wire _04749_;
 wire _04750_;
 wire _04751_;
 wire _04752_;
 wire _04753_;
 wire _04754_;
 wire _04755_;
 wire _04756_;
 wire _04757_;
 wire _04758_;
 wire _04759_;
 wire _04760_;
 wire _04761_;
 wire _04762_;
 wire _04763_;
 wire _04764_;
 wire _04765_;
 wire _04766_;
 wire _04767_;
 wire _04768_;
 wire _04769_;
 wire _04770_;
 wire _04771_;
 wire _04772_;
 wire _04773_;
 wire _04774_;
 wire _04775_;
 wire _04776_;
 wire _04777_;
 wire _04778_;
 wire _04779_;
 wire _04780_;
 wire _04781_;
 wire _04782_;
 wire _04783_;
 wire _04784_;
 wire _04785_;
 wire _04786_;
 wire _04787_;
 wire _04788_;
 wire _04789_;
 wire _04790_;
 wire _04791_;
 wire _04792_;
 wire _04793_;
 wire _04794_;
 wire _04795_;
 wire _04796_;
 wire _04797_;
 wire _04798_;
 wire _04799_;
 wire _04800_;
 wire _04801_;
 wire _04802_;
 wire _04803_;
 wire _04804_;
 wire _04805_;
 wire _04806_;
 wire _04807_;
 wire _04808_;
 wire _04809_;
 wire _04810_;
 wire _04811_;
 wire _04812_;
 wire _04813_;
 wire _04814_;
 wire _04815_;
 wire _04816_;
 wire _04817_;
 wire _04818_;
 wire _04819_;
 wire _04820_;
 wire _04821_;
 wire _04822_;
 wire _04823_;
 wire _04824_;
 wire _04825_;
 wire _04826_;
 wire _04827_;
 wire _04828_;
 wire _04829_;
 wire _04830_;
 wire _04831_;
 wire _04832_;
 wire _04833_;
 wire _04834_;
 wire _04835_;
 wire _04836_;
 wire _04837_;
 wire _04838_;
 wire _04839_;
 wire _04840_;
 wire _04841_;
 wire _04842_;
 wire _04843_;
 wire _04844_;
 wire _04845_;
 wire _04846_;
 wire _04847_;
 wire _04848_;
 wire _04849_;
 wire _04850_;
 wire _04851_;
 wire _04852_;
 wire _04853_;
 wire _04854_;
 wire _04855_;
 wire _04856_;
 wire _04857_;
 wire _04858_;
 wire _04859_;
 wire _04860_;
 wire _04861_;
 wire _04862_;
 wire _04863_;
 wire _04864_;
 wire _04865_;
 wire _04866_;
 wire _04867_;
 wire _04868_;
 wire _04869_;
 wire _04870_;
 wire _04871_;
 wire _04872_;
 wire _04873_;
 wire _04874_;
 wire _04875_;
 wire _04876_;
 wire _04877_;
 wire _04878_;
 wire _04879_;
 wire _04880_;
 wire _04881_;
 wire _04882_;
 wire _04883_;
 wire _04884_;
 wire _04885_;
 wire _04886_;
 wire _04887_;
 wire _04888_;
 wire _04889_;
 wire _04890_;
 wire _04891_;
 wire _04892_;
 wire _04893_;
 wire _04894_;
 wire _04895_;
 wire _04896_;
 wire _04897_;
 wire _04898_;
 wire _04899_;
 wire _04900_;
 wire _04901_;
 wire _04902_;
 wire _04903_;
 wire _04904_;
 wire _04905_;
 wire _04906_;
 wire _04907_;
 wire _04908_;
 wire _04909_;
 wire _04910_;
 wire _04911_;
 wire _04912_;
 wire _04913_;
 wire _04914_;
 wire _04915_;
 wire _04916_;
 wire _04917_;
 wire _04918_;
 wire _04919_;
 wire _04920_;
 wire _04921_;
 wire _04922_;
 wire _04923_;
 wire _04924_;
 wire _04925_;
 wire _04926_;
 wire _04927_;
 wire _04928_;
 wire _04929_;
 wire _04930_;
 wire _04931_;
 wire _04932_;
 wire _04933_;
 wire _04934_;
 wire _04935_;
 wire _04936_;
 wire _04937_;
 wire _04938_;
 wire _04939_;
 wire _04940_;
 wire _04941_;
 wire _04942_;
 wire _04943_;
 wire _04944_;
 wire _04945_;
 wire _04946_;
 wire _04947_;
 wire _04948_;
 wire _04949_;
 wire _04950_;
 wire _04951_;
 wire _04952_;
 wire _04953_;
 wire _04954_;
 wire _04955_;
 wire _04956_;
 wire _04957_;
 wire _04958_;
 wire _04959_;
 wire _04960_;
 wire _04961_;
 wire _04962_;
 wire _04963_;
 wire _04964_;
 wire _04965_;
 wire _04966_;
 wire _04967_;
 wire _04968_;
 wire _04969_;
 wire _04970_;
 wire _04971_;
 wire _04972_;
 wire _04973_;
 wire _04974_;
 wire _04975_;
 wire _04976_;
 wire _04977_;
 wire _04978_;
 wire _04979_;
 wire _04980_;
 wire _04981_;
 wire _04982_;
 wire _04983_;
 wire _04984_;
 wire _04985_;
 wire _04986_;
 wire _04987_;
 wire _04988_;
 wire _04989_;
 wire _04990_;
 wire _04991_;
 wire _04992_;
 wire _04993_;
 wire _04994_;
 wire _04995_;
 wire _04996_;
 wire _04997_;
 wire _04998_;
 wire _04999_;
 wire _05000_;
 wire _05001_;
 wire _05002_;
 wire _05003_;
 wire _05004_;
 wire _05005_;
 wire _05006_;
 wire _05007_;
 wire _05008_;
 wire _05009_;
 wire _05010_;
 wire _05011_;
 wire _05012_;
 wire _05013_;
 wire _05014_;
 wire _05015_;
 wire _05016_;
 wire _05017_;
 wire _05018_;
 wire _05019_;
 wire _05020_;
 wire _05021_;
 wire _05022_;
 wire _05023_;
 wire _05024_;
 wire _05025_;
 wire _05026_;
 wire _05027_;
 wire _05028_;
 wire _05029_;
 wire _05030_;
 wire _05031_;
 wire _05032_;
 wire _05033_;
 wire _05034_;
 wire _05035_;
 wire _05036_;
 wire _05037_;
 wire _05038_;
 wire _05039_;
 wire _05040_;
 wire _05041_;
 wire _05042_;
 wire _05043_;
 wire _05044_;
 wire _05045_;
 wire _05046_;
 wire _05047_;
 wire _05048_;
 wire _05049_;
 wire _05050_;
 wire _05051_;
 wire _05052_;
 wire _05053_;
 wire _05054_;
 wire _05055_;
 wire _05056_;
 wire _05057_;
 wire _05058_;
 wire _05059_;
 wire _05060_;
 wire _05061_;
 wire _05062_;
 wire _05063_;
 wire _05064_;
 wire _05065_;
 wire _05066_;
 wire _05067_;
 wire _05068_;
 wire _05069_;
 wire _05070_;
 wire _05071_;
 wire _05072_;
 wire _05073_;
 wire _05074_;
 wire _05075_;
 wire _05076_;
 wire _05077_;
 wire _05078_;
 wire _05079_;
 wire _05080_;
 wire _05081_;
 wire _05082_;
 wire _05083_;
 wire _05084_;
 wire _05085_;
 wire _05086_;
 wire _05087_;
 wire _05088_;
 wire _05089_;
 wire _05090_;
 wire _05091_;
 wire _05092_;
 wire _05093_;
 wire _05094_;
 wire _05095_;
 wire _05096_;
 wire _05097_;
 wire _05098_;
 wire _05099_;
 wire _05100_;
 wire _05101_;
 wire _05102_;
 wire _05103_;
 wire _05104_;
 wire _05105_;
 wire _05106_;
 wire _05107_;
 wire _05108_;
 wire _05109_;
 wire _05110_;
 wire _05111_;
 wire _05112_;
 wire _05113_;
 wire _05114_;
 wire _05115_;
 wire _05116_;
 wire _05117_;
 wire _05118_;
 wire _05119_;
 wire _05120_;
 wire _05121_;
 wire _05122_;
 wire _05123_;
 wire _05124_;
 wire _05125_;
 wire _05126_;
 wire _05127_;
 wire _05128_;
 wire _05129_;
 wire _05130_;
 wire _05131_;
 wire _05132_;
 wire _05133_;
 wire _05134_;
 wire _05135_;
 wire _05136_;
 wire _05137_;
 wire _05138_;
 wire _05139_;
 wire _05140_;
 wire _05141_;
 wire _05142_;
 wire _05143_;
 wire _05144_;
 wire _05145_;
 wire _05146_;
 wire _05147_;
 wire _05148_;
 wire _05149_;
 wire _05150_;
 wire _05151_;
 wire _05152_;
 wire _05153_;
 wire _05154_;
 wire _05155_;
 wire _05156_;
 wire _05157_;
 wire _05158_;
 wire _05159_;
 wire _05160_;
 wire _05161_;
 wire _05162_;
 wire _05163_;
 wire _05164_;
 wire _05165_;
 wire _05166_;
 wire _05167_;
 wire _05168_;
 wire _05169_;
 wire _05170_;
 wire _05171_;
 wire _05172_;
 wire _05173_;
 wire _05174_;
 wire _05175_;
 wire _05176_;
 wire _05177_;
 wire _05178_;
 wire _05179_;
 wire _05180_;
 wire _05181_;
 wire _05182_;
 wire _05183_;
 wire _05184_;
 wire _05185_;
 wire _05186_;
 wire _05187_;
 wire _05188_;
 wire _05189_;
 wire _05190_;
 wire _05191_;
 wire _05192_;
 wire _05193_;
 wire _05194_;
 wire _05195_;
 wire _05196_;
 wire _05197_;
 wire _05198_;
 wire _05199_;
 wire _05200_;
 wire _05201_;
 wire _05202_;
 wire _05203_;
 wire _05204_;
 wire _05205_;
 wire _05206_;
 wire _05207_;
 wire _05208_;
 wire _05209_;
 wire _05210_;
 wire _05211_;
 wire _05212_;
 wire _05213_;
 wire _05214_;
 wire _05215_;
 wire _05216_;
 wire _05217_;
 wire _05218_;
 wire _05219_;
 wire _05220_;
 wire _05221_;
 wire _05222_;
 wire _05223_;
 wire _05224_;
 wire _05225_;
 wire _05226_;
 wire _05227_;
 wire _05228_;
 wire _05229_;
 wire _05230_;
 wire _05231_;
 wire _05232_;
 wire _05233_;
 wire _05234_;
 wire _05235_;
 wire _05236_;
 wire _05237_;
 wire _05238_;
 wire _05239_;
 wire _05240_;
 wire _05241_;
 wire _05242_;
 wire _05243_;
 wire _05244_;
 wire _05245_;
 wire _05246_;
 wire _05247_;
 wire _05248_;
 wire _05249_;
 wire _05250_;
 wire _05251_;
 wire _05252_;
 wire _05253_;
 wire _05254_;
 wire _05255_;
 wire _05256_;
 wire _05257_;
 wire _05258_;
 wire _05259_;
 wire _05260_;
 wire _05261_;
 wire _05262_;
 wire _05263_;
 wire _05264_;
 wire _05265_;
 wire _05266_;
 wire _05267_;
 wire _05268_;
 wire _05269_;
 wire _05270_;
 wire _05271_;
 wire _05272_;
 wire _05273_;
 wire _05274_;
 wire _05275_;
 wire _05276_;
 wire _05277_;
 wire _05278_;
 wire _05279_;
 wire _05280_;
 wire _05281_;
 wire _05282_;
 wire _05283_;
 wire _05284_;
 wire _05285_;
 wire _05286_;
 wire _05287_;
 wire _05288_;
 wire _05289_;
 wire _05290_;
 wire _05291_;
 wire _05292_;
 wire _05293_;
 wire _05294_;
 wire _05295_;
 wire _05296_;
 wire _05297_;
 wire _05298_;
 wire _05299_;
 wire _05300_;
 wire _05301_;
 wire _05302_;
 wire _05303_;
 wire _05304_;
 wire _05305_;
 wire _05306_;
 wire _05307_;
 wire _05308_;
 wire _05309_;
 wire _05310_;
 wire _05311_;
 wire _05312_;
 wire _05313_;
 wire _05314_;
 wire _05315_;
 wire _05316_;
 wire _05317_;
 wire _05318_;
 wire _05319_;
 wire _05320_;
 wire _05321_;
 wire _05322_;
 wire _05323_;
 wire _05324_;
 wire _05325_;
 wire _05326_;
 wire _05327_;
 wire _05328_;
 wire _05329_;
 wire _05330_;
 wire _05331_;
 wire _05332_;
 wire _05333_;
 wire _05334_;
 wire _05335_;
 wire _05336_;
 wire _05337_;
 wire _05338_;
 wire _05339_;
 wire _05340_;
 wire _05341_;
 wire _05342_;
 wire _05343_;
 wire _05344_;
 wire _05345_;
 wire _05346_;
 wire _05347_;
 wire _05348_;
 wire _05349_;
 wire _05350_;
 wire _05351_;
 wire _05352_;
 wire _05353_;
 wire _05354_;
 wire _05355_;
 wire _05356_;
 wire _05357_;
 wire _05358_;
 wire _05359_;
 wire _05360_;
 wire _05361_;
 wire _05362_;
 wire _05363_;
 wire _05364_;
 wire _05365_;
 wire _05366_;
 wire _05367_;
 wire _05368_;
 wire _05369_;
 wire _05370_;
 wire _05371_;
 wire _05372_;
 wire _05373_;
 wire _05374_;
 wire _05375_;
 wire _05376_;
 wire _05377_;
 wire _05378_;
 wire _05379_;
 wire _05380_;
 wire _05381_;
 wire _05382_;
 wire _05383_;
 wire _05384_;
 wire _05385_;
 wire _05386_;
 wire _05387_;
 wire _05388_;
 wire _05389_;
 wire _05390_;
 wire _05391_;
 wire _05392_;
 wire _05393_;
 wire _05394_;
 wire _05395_;
 wire _05396_;
 wire _05397_;
 wire _05398_;
 wire _05399_;
 wire _05400_;
 wire _05401_;
 wire _05402_;
 wire _05403_;
 wire _05404_;
 wire _05405_;
 wire _05406_;
 wire _05407_;
 wire _05408_;
 wire _05409_;
 wire _05410_;
 wire _05411_;
 wire _05412_;
 wire _05413_;
 wire _05414_;
 wire _05415_;
 wire _05416_;
 wire _05417_;
 wire _05418_;
 wire _05419_;
 wire _05420_;
 wire _05421_;
 wire _05422_;
 wire _05423_;
 wire _05424_;
 wire _05425_;
 wire _05426_;
 wire _05427_;
 wire _05428_;
 wire _05429_;
 wire _05430_;
 wire _05431_;
 wire _05432_;
 wire _05433_;
 wire _05434_;
 wire _05435_;
 wire _05436_;
 wire _05437_;
 wire _05438_;
 wire _05439_;
 wire _05440_;
 wire _05441_;
 wire _05442_;
 wire _05443_;
 wire _05444_;
 wire _05445_;
 wire _05446_;
 wire _05447_;
 wire _05448_;
 wire _05449_;
 wire _05450_;
 wire _05451_;
 wire _05452_;
 wire _05453_;
 wire _05454_;
 wire _05455_;
 wire _05456_;
 wire _05457_;
 wire _05458_;
 wire _05459_;
 wire _05460_;
 wire _05461_;
 wire _05462_;
 wire _05463_;
 wire _05464_;
 wire _05465_;
 wire _05466_;
 wire _05467_;
 wire _05468_;
 wire _05469_;
 wire _05470_;
 wire _05471_;
 wire _05472_;
 wire _05473_;
 wire _05474_;
 wire _05475_;
 wire _05476_;
 wire _05477_;
 wire _05478_;
 wire _05479_;
 wire _05480_;
 wire _05481_;
 wire _05482_;
 wire _05483_;
 wire _05484_;
 wire _05485_;
 wire _05486_;
 wire _05487_;
 wire _05488_;
 wire _05489_;
 wire _05490_;
 wire _05491_;
 wire _05492_;
 wire _05493_;
 wire _05494_;
 wire _05495_;
 wire _05496_;
 wire _05497_;
 wire _05498_;
 wire _05499_;
 wire _05500_;
 wire _05501_;
 wire _05502_;
 wire _05503_;
 wire _05504_;
 wire _05505_;
 wire _05506_;
 wire _05507_;
 wire _05508_;
 wire _05509_;
 wire _05510_;
 wire _05511_;
 wire _05512_;
 wire _05513_;
 wire _05514_;
 wire _05515_;
 wire _05516_;
 wire _05517_;
 wire _05518_;
 wire _05519_;
 wire _05520_;
 wire _05521_;
 wire _05522_;
 wire _05523_;
 wire _05524_;
 wire _05525_;
 wire _05526_;
 wire _05527_;
 wire _05528_;
 wire _05529_;
 wire _05530_;
 wire _05531_;
 wire _05532_;
 wire _05533_;
 wire _05534_;
 wire _05535_;
 wire _05536_;
 wire _05537_;
 wire _05538_;
 wire _05539_;
 wire _05540_;
 wire _05541_;
 wire _05542_;
 wire _05543_;
 wire _05544_;
 wire _05545_;
 wire _05546_;
 wire _05547_;
 wire _05548_;
 wire _05549_;
 wire _05550_;
 wire _05551_;
 wire _05552_;
 wire _05553_;
 wire _05554_;
 wire _05555_;
 wire _05556_;
 wire _05557_;
 wire _05558_;
 wire _05559_;
 wire _05560_;
 wire _05561_;
 wire _05562_;
 wire _05563_;
 wire _05564_;
 wire _05565_;
 wire _05566_;
 wire _05567_;
 wire _05568_;
 wire _05569_;
 wire _05570_;
 wire _05571_;
 wire _05572_;
 wire _05573_;
 wire _05574_;
 wire _05575_;
 wire _05576_;
 wire _05577_;
 wire _05578_;
 wire _05579_;
 wire _05580_;
 wire _05581_;
 wire _05582_;
 wire _05583_;
 wire _05584_;
 wire _05585_;
 wire _05586_;
 wire _05587_;
 wire _05588_;
 wire _05589_;
 wire _05590_;
 wire _05591_;
 wire _05592_;
 wire _05593_;
 wire _05594_;
 wire _05595_;
 wire _05596_;
 wire _05597_;
 wire _05598_;
 wire _05599_;
 wire _05600_;
 wire _05601_;
 wire _05602_;
 wire _05603_;
 wire _05604_;
 wire _05605_;
 wire _05606_;
 wire _05607_;
 wire _05608_;
 wire _05609_;
 wire _05610_;
 wire _05611_;
 wire _05612_;
 wire _05613_;
 wire _05614_;
 wire _05615_;
 wire _05616_;
 wire _05617_;
 wire _05618_;
 wire _05619_;
 wire _05620_;
 wire _05621_;
 wire _05622_;
 wire _05623_;
 wire _05624_;
 wire _05625_;
 wire _05626_;
 wire _05627_;
 wire _05628_;
 wire _05629_;
 wire _05630_;
 wire _05631_;
 wire _05632_;
 wire _05633_;
 wire _05634_;
 wire _05635_;
 wire _05636_;
 wire _05637_;
 wire _05638_;
 wire _05639_;
 wire _05640_;
 wire _05641_;
 wire _05642_;
 wire _05643_;
 wire _05644_;
 wire _05645_;
 wire _05646_;
 wire _05647_;
 wire _05648_;
 wire _05649_;
 wire _05650_;
 wire _05651_;
 wire _05652_;
 wire _05653_;
 wire _05654_;
 wire _05655_;
 wire _05656_;
 wire _05657_;
 wire _05658_;
 wire _05659_;
 wire _05660_;
 wire _05661_;
 wire _05662_;
 wire _05663_;
 wire _05664_;
 wire _05665_;
 wire _05666_;
 wire _05667_;
 wire _05668_;
 wire _05669_;
 wire _05670_;
 wire _05671_;
 wire _05672_;
 wire _05673_;
 wire _05674_;
 wire _05675_;
 wire _05676_;
 wire _05677_;
 wire _05678_;
 wire _05679_;
 wire _05680_;
 wire _05681_;
 wire _05682_;
 wire _05683_;
 wire _05684_;
 wire _05685_;
 wire _05686_;
 wire _05687_;
 wire _05688_;
 wire _05689_;
 wire _05690_;
 wire _05691_;
 wire _05692_;
 wire _05693_;
 wire _05694_;
 wire _05695_;
 wire _05696_;
 wire _05697_;
 wire _05698_;
 wire _05699_;
 wire _05700_;
 wire _05701_;
 wire _05702_;
 wire _05703_;
 wire _05704_;
 wire _05705_;
 wire _05706_;
 wire _05707_;
 wire _05708_;
 wire _05709_;
 wire _05710_;
 wire _05711_;
 wire _05712_;
 wire _05713_;
 wire _05714_;
 wire _05715_;
 wire _05716_;
 wire _05717_;
 wire _05718_;
 wire _05719_;
 wire _05720_;
 wire _05721_;
 wire _05722_;
 wire _05723_;
 wire _05724_;
 wire _05725_;
 wire _05726_;
 wire _05727_;
 wire _05728_;
 wire _05729_;
 wire _05730_;
 wire _05731_;
 wire _05732_;
 wire _05733_;
 wire _05734_;
 wire _05735_;
 wire _05736_;
 wire _05737_;
 wire _05738_;
 wire _05739_;
 wire _05740_;
 wire _05741_;
 wire _05742_;
 wire _05743_;
 wire _05744_;
 wire _05745_;
 wire _05746_;
 wire _05747_;
 wire _05748_;
 wire _05749_;
 wire _05750_;
 wire _05751_;
 wire _05752_;
 wire _05753_;
 wire _05754_;
 wire _05755_;
 wire _05756_;
 wire _05757_;
 wire _05758_;
 wire _05759_;
 wire _05760_;
 wire _05761_;
 wire _05762_;
 wire _05763_;
 wire _05764_;
 wire _05765_;
 wire _05766_;
 wire _05767_;
 wire _05768_;
 wire _05769_;
 wire _05770_;
 wire _05771_;
 wire _05772_;
 wire _05773_;
 wire _05774_;
 wire _05775_;
 wire _05776_;
 wire _05777_;
 wire _05778_;
 wire _05779_;
 wire _05780_;
 wire _05781_;
 wire _05782_;
 wire _05783_;
 wire _05784_;
 wire _05785_;
 wire _05786_;
 wire _05787_;
 wire _05788_;
 wire _05789_;
 wire _05790_;
 wire _05791_;
 wire _05792_;
 wire _05793_;
 wire _05794_;
 wire _05795_;
 wire _05796_;
 wire _05797_;
 wire _05798_;
 wire _05799_;
 wire _05800_;
 wire _05801_;
 wire _05802_;
 wire _05803_;
 wire _05804_;
 wire _05805_;
 wire _05806_;
 wire _05807_;
 wire _05808_;
 wire _05809_;
 wire _05810_;
 wire _05811_;
 wire _05812_;
 wire _05813_;
 wire _05814_;
 wire _05815_;
 wire _05816_;
 wire _05817_;
 wire _05818_;
 wire _05819_;
 wire _05820_;
 wire _05821_;
 wire _05822_;
 wire _05823_;
 wire _05824_;
 wire _05825_;
 wire _05826_;
 wire _05827_;
 wire _05828_;
 wire _05829_;
 wire _05830_;
 wire _05831_;
 wire _05832_;
 wire _05833_;
 wire _05834_;
 wire _05835_;
 wire _05836_;
 wire _05837_;
 wire _05838_;
 wire _05839_;
 wire _05840_;
 wire _05841_;
 wire _05842_;
 wire _05843_;
 wire _05844_;
 wire _05845_;
 wire _05846_;
 wire _05847_;
 wire _05848_;
 wire _05849_;
 wire _05850_;
 wire _05851_;
 wire _05852_;
 wire _05853_;
 wire _05854_;
 wire _05855_;
 wire _05856_;
 wire _05857_;
 wire _05858_;
 wire _05859_;
 wire _05860_;
 wire _05861_;
 wire _05862_;
 wire _05863_;
 wire _05864_;
 wire _05865_;
 wire _05866_;
 wire _05867_;
 wire _05868_;
 wire _05869_;
 wire _05870_;
 wire _05871_;
 wire _05872_;
 wire _05873_;
 wire _05874_;
 wire _05875_;
 wire _05876_;
 wire _05877_;
 wire _05878_;
 wire _05879_;
 wire _05880_;
 wire _05881_;
 wire _05882_;
 wire _05883_;
 wire _05884_;
 wire _05885_;
 wire _05886_;
 wire _05887_;
 wire _05888_;
 wire _05889_;
 wire _05890_;
 wire _05891_;
 wire _05892_;
 wire _05893_;
 wire _05894_;
 wire _05895_;
 wire _05896_;
 wire _05897_;
 wire _05898_;
 wire _05899_;
 wire _05900_;
 wire _05901_;
 wire _05902_;
 wire _05903_;
 wire _05904_;
 wire _05905_;
 wire _05906_;
 wire _05907_;
 wire _05908_;
 wire _05909_;
 wire _05910_;
 wire _05911_;
 wire _05912_;
 wire _05913_;
 wire _05914_;
 wire _05915_;
 wire _05916_;
 wire _05917_;
 wire _05918_;
 wire _05919_;
 wire _05920_;
 wire _05921_;
 wire _05922_;
 wire _05923_;
 wire _05924_;
 wire _05925_;
 wire _05926_;
 wire _05927_;
 wire _05928_;
 wire _05929_;
 wire _05930_;
 wire _05931_;
 wire _05932_;
 wire _05933_;
 wire _05934_;
 wire _05935_;
 wire _05936_;
 wire _05937_;
 wire _05938_;
 wire _05939_;
 wire _05940_;
 wire _05941_;
 wire _05942_;
 wire _05943_;
 wire _05944_;
 wire _05945_;
 wire _05946_;
 wire _05947_;
 wire _05948_;
 wire _05949_;
 wire _05950_;
 wire _05951_;
 wire _05952_;
 wire _05953_;
 wire _05954_;
 wire _05955_;
 wire _05956_;
 wire _05957_;
 wire _05958_;
 wire _05959_;
 wire _05960_;
 wire _05961_;
 wire _05962_;
 wire _05963_;
 wire _05964_;
 wire _05965_;
 wire _05966_;
 wire _05967_;
 wire _05968_;
 wire _05969_;
 wire _05970_;
 wire _05971_;
 wire _05972_;
 wire _05973_;
 wire _05974_;
 wire _05975_;
 wire _05976_;
 wire _05977_;
 wire _05978_;
 wire _05979_;
 wire _05980_;
 wire _05981_;
 wire _05982_;
 wire _05983_;
 wire _05984_;
 wire _05985_;
 wire _05986_;
 wire _05987_;
 wire _05988_;
 wire _05989_;
 wire _05990_;
 wire _05991_;
 wire _05992_;
 wire _05993_;
 wire _05994_;
 wire _05995_;
 wire _05996_;
 wire _05997_;
 wire _05998_;
 wire _05999_;
 wire _06000_;
 wire _06001_;
 wire _06002_;
 wire _06003_;
 wire _06004_;
 wire _06005_;
 wire _06006_;
 wire _06007_;
 wire _06008_;
 wire _06009_;
 wire _06010_;
 wire _06011_;
 wire _06012_;
 wire _06013_;
 wire _06014_;
 wire _06015_;
 wire _06016_;
 wire _06017_;
 wire _06018_;
 wire _06019_;
 wire _06020_;
 wire _06021_;
 wire _06022_;
 wire _06023_;
 wire _06024_;
 wire _06025_;
 wire _06026_;
 wire _06027_;
 wire _06028_;
 wire _06029_;
 wire _06030_;
 wire _06031_;
 wire _06032_;
 wire _06033_;
 wire _06034_;
 wire _06035_;
 wire _06036_;
 wire _06037_;
 wire _06038_;
 wire _06039_;
 wire _06040_;
 wire _06041_;
 wire _06042_;
 wire _06043_;
 wire _06044_;
 wire _06045_;
 wire _06046_;
 wire _06047_;
 wire _06048_;
 wire _06049_;
 wire _06050_;
 wire _06051_;
 wire _06052_;
 wire _06053_;
 wire _06054_;
 wire _06055_;
 wire _06056_;
 wire _06057_;
 wire _06058_;
 wire _06059_;
 wire _06060_;
 wire _06061_;
 wire _06062_;
 wire _06063_;
 wire _06064_;
 wire _06065_;
 wire _06066_;
 wire _06067_;
 wire _06068_;
 wire _06069_;
 wire _06070_;
 wire _06071_;
 wire _06072_;
 wire _06073_;
 wire _06074_;
 wire _06075_;
 wire _06076_;
 wire _06077_;
 wire _06078_;
 wire _06079_;
 wire _06080_;
 wire _06081_;
 wire _06082_;
 wire _06083_;
 wire _06084_;
 wire _06085_;
 wire _06086_;
 wire _06087_;
 wire _06088_;
 wire _06089_;
 wire _06090_;
 wire _06091_;
 wire _06092_;
 wire _06093_;
 wire _06094_;
 wire _06095_;
 wire _06096_;
 wire _06097_;
 wire _06098_;
 wire _06099_;
 wire _06100_;
 wire _06101_;
 wire _06102_;
 wire _06103_;
 wire _06104_;
 wire _06105_;
 wire _06106_;
 wire _06107_;
 wire _06108_;
 wire _06109_;
 wire _06110_;
 wire _06111_;
 wire _06112_;
 wire _06113_;
 wire _06114_;
 wire _06115_;
 wire _06116_;
 wire _06117_;
 wire _06118_;
 wire _06119_;
 wire _06120_;
 wire _06121_;
 wire _06122_;
 wire _06123_;
 wire _06124_;
 wire _06125_;
 wire _06126_;
 wire _06127_;
 wire _06128_;
 wire _06129_;
 wire _06130_;
 wire _06131_;
 wire _06132_;
 wire _06133_;
 wire _06134_;
 wire _06135_;
 wire _06136_;
 wire _06137_;
 wire _06138_;
 wire _06139_;
 wire _06140_;
 wire _06141_;
 wire _06142_;
 wire _06143_;
 wire _06144_;
 wire _06145_;
 wire _06146_;
 wire _06147_;
 wire _06148_;
 wire _06149_;
 wire _06150_;
 wire _06151_;
 wire _06152_;
 wire _06153_;
 wire _06154_;
 wire _06155_;
 wire _06156_;
 wire _06157_;
 wire _06158_;
 wire _06159_;
 wire _06160_;
 wire _06161_;
 wire _06162_;
 wire _06163_;
 wire _06164_;
 wire _06165_;
 wire _06166_;
 wire _06167_;
 wire _06168_;
 wire _06169_;
 wire _06170_;
 wire _06171_;
 wire _06172_;
 wire _06173_;
 wire _06174_;
 wire _06175_;
 wire _06176_;
 wire _06177_;
 wire _06178_;
 wire _06179_;
 wire _06180_;
 wire _06181_;
 wire _06182_;
 wire _06183_;
 wire _06184_;
 wire _06185_;
 wire _06186_;
 wire _06187_;
 wire _06188_;
 wire _06189_;
 wire _06190_;
 wire _06191_;
 wire _06192_;
 wire _06193_;
 wire _06194_;
 wire _06195_;
 wire _06196_;
 wire _06197_;
 wire _06198_;
 wire _06199_;
 wire _06200_;
 wire _06201_;
 wire _06202_;
 wire _06203_;
 wire _06204_;
 wire _06205_;
 wire _06206_;
 wire _06207_;
 wire _06208_;
 wire _06209_;
 wire _06210_;
 wire _06211_;
 wire _06212_;
 wire _06213_;
 wire _06214_;
 wire _06215_;
 wire _06216_;
 wire _06217_;
 wire _06218_;
 wire _06219_;
 wire _06220_;
 wire _06221_;
 wire _06222_;
 wire _06223_;
 wire _06224_;
 wire _06225_;
 wire _06226_;
 wire _06227_;
 wire _06228_;
 wire _06229_;
 wire _06230_;
 wire _06231_;
 wire _06232_;
 wire _06233_;
 wire _06234_;
 wire _06235_;
 wire _06236_;
 wire _06237_;
 wire _06238_;
 wire _06239_;
 wire _06240_;
 wire _06241_;
 wire _06242_;
 wire _06243_;
 wire _06244_;
 wire _06245_;
 wire _06246_;
 wire _06247_;
 wire _06248_;
 wire _06249_;
 wire _06250_;
 wire _06251_;
 wire _06252_;
 wire _06253_;
 wire _06254_;
 wire _06255_;
 wire _06256_;
 wire _06257_;
 wire _06258_;
 wire _06259_;
 wire _06260_;
 wire _06261_;
 wire _06262_;
 wire _06263_;
 wire _06264_;
 wire _06265_;
 wire _06266_;
 wire _06267_;
 wire _06268_;
 wire _06269_;
 wire _06270_;
 wire _06271_;
 wire _06272_;
 wire _06273_;
 wire _06274_;
 wire _06275_;
 wire _06276_;
 wire _06277_;
 wire _06278_;
 wire _06279_;
 wire _06280_;
 wire _06281_;
 wire _06282_;
 wire _06283_;
 wire _06284_;
 wire _06285_;
 wire _06286_;
 wire _06287_;
 wire _06288_;
 wire _06289_;
 wire _06290_;
 wire _06291_;
 wire _06292_;
 wire _06293_;
 wire _06294_;
 wire _06295_;
 wire _06296_;
 wire _06297_;
 wire _06298_;
 wire _06299_;
 wire _06300_;
 wire _06301_;
 wire _06302_;
 wire _06303_;
 wire _06304_;
 wire _06305_;
 wire _06306_;
 wire _06307_;
 wire _06308_;
 wire _06309_;
 wire _06310_;
 wire _06311_;
 wire _06312_;
 wire _06313_;
 wire _06314_;
 wire _06315_;
 wire _06316_;
 wire _06317_;
 wire _06318_;
 wire _06319_;
 wire _06320_;
 wire _06321_;
 wire _06322_;
 wire _06323_;
 wire _06324_;
 wire _06325_;
 wire _06326_;
 wire _06327_;
 wire _06328_;
 wire _06329_;
 wire _06330_;
 wire _06331_;
 wire _06332_;
 wire _06333_;
 wire _06334_;
 wire _06335_;
 wire _06336_;
 wire _06337_;
 wire _06338_;
 wire _06339_;
 wire _06340_;
 wire _06341_;
 wire _06342_;
 wire _06343_;
 wire _06344_;
 wire _06345_;
 wire _06346_;
 wire _06347_;
 wire _06348_;
 wire _06349_;
 wire _06350_;
 wire _06351_;
 wire _06352_;
 wire _06353_;
 wire _06354_;
 wire _06355_;
 wire _06356_;
 wire _06357_;
 wire _06358_;
 wire _06359_;
 wire _06360_;
 wire _06361_;
 wire _06362_;
 wire _06363_;
 wire _06364_;
 wire _06365_;
 wire _06366_;
 wire _06367_;
 wire _06368_;
 wire _06369_;
 wire _06370_;
 wire _06371_;
 wire _06372_;
 wire _06373_;
 wire _06374_;
 wire _06375_;
 wire _06376_;
 wire _06377_;
 wire _06378_;
 wire _06379_;
 wire _06380_;
 wire _06381_;
 wire _06382_;
 wire _06383_;
 wire _06384_;
 wire _06385_;
 wire _06386_;
 wire _06387_;
 wire _06388_;
 wire _06389_;
 wire _06390_;
 wire _06391_;
 wire _06392_;
 wire _06393_;
 wire _06394_;
 wire _06395_;
 wire _06396_;
 wire _06397_;
 wire _06398_;
 wire _06399_;
 wire _06400_;
 wire _06401_;
 wire _06402_;
 wire _06403_;
 wire _06404_;
 wire _06405_;
 wire _06406_;
 wire _06407_;
 wire _06408_;
 wire _06409_;
 wire _06410_;
 wire _06411_;
 wire _06412_;
 wire _06413_;
 wire _06414_;
 wire _06415_;
 wire _06416_;
 wire _06417_;
 wire _06418_;
 wire _06419_;
 wire _06420_;
 wire _06421_;
 wire _06422_;
 wire _06423_;
 wire _06424_;
 wire _06425_;
 wire _06426_;
 wire _06427_;
 wire _06428_;
 wire _06429_;
 wire _06430_;
 wire _06431_;
 wire _06432_;
 wire _06433_;
 wire _06434_;
 wire _06435_;
 wire _06436_;
 wire _06437_;
 wire _06438_;
 wire _06439_;
 wire _06440_;
 wire _06441_;
 wire _06442_;
 wire _06443_;
 wire _06444_;
 wire _06445_;
 wire _06446_;
 wire _06447_;
 wire _06448_;
 wire _06449_;
 wire _06450_;
 wire _06451_;
 wire _06452_;
 wire _06453_;
 wire _06454_;
 wire _06455_;
 wire _06456_;
 wire _06457_;
 wire _06458_;
 wire _06459_;
 wire _06460_;
 wire _06461_;
 wire _06462_;
 wire _06463_;
 wire _06464_;
 wire _06465_;
 wire _06466_;
 wire _06467_;
 wire _06468_;
 wire _06469_;
 wire _06470_;
 wire _06471_;
 wire _06472_;
 wire _06473_;
 wire _06474_;
 wire _06475_;
 wire _06476_;
 wire _06477_;
 wire _06478_;
 wire _06479_;
 wire _06480_;
 wire _06481_;
 wire _06482_;
 wire _06483_;
 wire _06484_;
 wire _06485_;
 wire _06486_;
 wire _06487_;
 wire _06488_;
 wire _06489_;
 wire _06490_;
 wire _06491_;
 wire _06492_;
 wire _06493_;
 wire _06494_;
 wire _06495_;
 wire _06496_;
 wire _06497_;
 wire _06498_;
 wire _06499_;
 wire _06500_;
 wire _06501_;
 wire _06502_;
 wire _06503_;
 wire _06504_;
 wire _06505_;
 wire _06506_;
 wire _06507_;
 wire _06508_;
 wire _06509_;
 wire _06510_;
 wire _06511_;
 wire _06512_;
 wire _06513_;
 wire _06514_;
 wire _06515_;
 wire _06516_;
 wire _06517_;
 wire _06518_;
 wire _06519_;
 wire _06520_;
 wire _06521_;
 wire _06522_;
 wire _06523_;
 wire _06524_;
 wire _06525_;
 wire _06526_;
 wire _06527_;
 wire _06528_;
 wire _06529_;
 wire _06530_;
 wire _06531_;
 wire _06532_;
 wire _06533_;
 wire _06534_;
 wire _06535_;
 wire _06536_;
 wire _06537_;
 wire _06538_;
 wire _06539_;
 wire _06540_;
 wire _06541_;
 wire _06542_;
 wire _06543_;
 wire _06544_;
 wire _06545_;
 wire _06546_;
 wire _06547_;
 wire _06548_;
 wire _06549_;
 wire _06550_;
 wire _06551_;
 wire _06552_;
 wire _06553_;
 wire _06554_;
 wire _06555_;
 wire _06556_;
 wire _06557_;
 wire _06558_;
 wire _06559_;
 wire _06560_;
 wire _06561_;
 wire _06562_;
 wire _06563_;
 wire _06564_;
 wire _06565_;
 wire _06566_;
 wire _06567_;
 wire _06568_;
 wire _06569_;
 wire _06570_;
 wire _06571_;
 wire _06572_;
 wire _06573_;
 wire _06574_;
 wire _06575_;
 wire _06576_;
 wire _06577_;
 wire _06578_;
 wire _06579_;
 wire _06580_;
 wire _06581_;
 wire _06582_;
 wire _06583_;
 wire _06584_;
 wire _06585_;
 wire _06586_;
 wire _06587_;
 wire _06588_;
 wire _06589_;
 wire _06590_;
 wire _06591_;
 wire _06592_;
 wire _06593_;
 wire _06594_;
 wire _06595_;
 wire _06596_;
 wire _06597_;
 wire _06598_;
 wire _06599_;
 wire _06600_;
 wire _06601_;
 wire _06602_;
 wire _06603_;
 wire _06604_;
 wire _06605_;
 wire _06606_;
 wire _06607_;
 wire _06608_;
 wire _06609_;
 wire _06610_;
 wire _06611_;
 wire _06612_;
 wire _06613_;
 wire _06614_;
 wire _06615_;
 wire _06616_;
 wire _06617_;
 wire _06618_;
 wire _06619_;
 wire _06620_;
 wire _06621_;
 wire _06622_;
 wire _06623_;
 wire _06624_;
 wire _06625_;
 wire _06626_;
 wire _06627_;
 wire _06628_;
 wire _06629_;
 wire _06630_;
 wire _06631_;
 wire _06632_;
 wire _06633_;
 wire _06634_;
 wire _06635_;
 wire _06636_;
 wire _06637_;
 wire _06638_;
 wire _06639_;
 wire _06640_;
 wire _06641_;
 wire _06642_;
 wire _06643_;
 wire _06644_;
 wire _06645_;
 wire _06646_;
 wire _06647_;
 wire _06648_;
 wire _06649_;
 wire _06650_;
 wire _06651_;
 wire _06652_;
 wire _06653_;
 wire _06654_;
 wire _06655_;
 wire _06656_;
 wire _06657_;
 wire _06658_;
 wire _06659_;
 wire _06660_;
 wire _06661_;
 wire _06662_;
 wire _06663_;
 wire _06664_;
 wire _06665_;
 wire _06666_;
 wire _06667_;
 wire _06668_;
 wire _06669_;
 wire _06670_;
 wire _06671_;
 wire _06672_;
 wire _06673_;
 wire _06674_;
 wire _06675_;
 wire _06676_;
 wire _06677_;
 wire _06678_;
 wire _06679_;
 wire _06680_;
 wire _06681_;
 wire _06682_;
 wire _06683_;
 wire _06684_;
 wire _06685_;
 wire _06686_;
 wire _06687_;
 wire _06688_;
 wire _06689_;
 wire _06690_;
 wire _06691_;
 wire _06692_;
 wire _06693_;
 wire _06694_;
 wire _06695_;
 wire _06696_;
 wire _06697_;
 wire _06698_;
 wire _06699_;
 wire _06700_;
 wire _06701_;
 wire _06702_;
 wire _06703_;
 wire _06704_;
 wire _06705_;
 wire _06706_;
 wire _06707_;
 wire _06708_;
 wire _06709_;
 wire _06710_;
 wire _06711_;
 wire _06712_;
 wire _06713_;
 wire _06714_;
 wire _06715_;
 wire _06716_;
 wire _06717_;
 wire _06718_;
 wire _06719_;
 wire _06720_;
 wire _06721_;
 wire _06722_;
 wire _06723_;
 wire _06724_;
 wire _06725_;
 wire _06726_;
 wire _06727_;
 wire _06728_;
 wire _06729_;
 wire _06730_;
 wire _06731_;
 wire _06732_;
 wire _06733_;
 wire _06734_;
 wire _06735_;
 wire _06736_;
 wire _06737_;
 wire _06738_;
 wire _06739_;
 wire _06740_;
 wire _06741_;
 wire _06742_;
 wire _06743_;
 wire _06744_;
 wire _06745_;
 wire _06746_;
 wire _06747_;
 wire _06748_;
 wire _06749_;
 wire _06750_;
 wire _06751_;
 wire _06752_;
 wire _06753_;
 wire _06754_;
 wire _06755_;
 wire _06756_;
 wire _06757_;
 wire _06758_;
 wire _06759_;
 wire _06760_;
 wire _06761_;
 wire _06762_;
 wire _06763_;
 wire _06764_;
 wire _06765_;
 wire _06766_;
 wire _06767_;
 wire _06768_;
 wire _06769_;
 wire _06770_;
 wire _06771_;
 wire _06772_;
 wire _06773_;
 wire _06774_;
 wire _06775_;
 wire _06776_;
 wire _06777_;
 wire _06778_;
 wire _06779_;
 wire _06780_;
 wire _06781_;
 wire _06782_;
 wire _06783_;
 wire _06784_;
 wire _06785_;
 wire _06786_;
 wire _06787_;
 wire _06788_;
 wire _06789_;
 wire _06790_;
 wire _06791_;
 wire _06792_;
 wire _06793_;
 wire _06794_;
 wire _06795_;
 wire _06796_;
 wire _06797_;
 wire _06798_;
 wire _06799_;
 wire _06800_;
 wire _06801_;
 wire _06802_;
 wire _06803_;
 wire _06804_;
 wire _06805_;
 wire _06806_;
 wire _06807_;
 wire _06808_;
 wire _06809_;
 wire _06810_;
 wire _06811_;
 wire _06812_;
 wire _06813_;
 wire _06814_;
 wire _06815_;
 wire _06816_;
 wire _06817_;
 wire _06818_;
 wire _06819_;
 wire _06820_;
 wire _06821_;
 wire _06822_;
 wire _06823_;
 wire _06824_;
 wire _06825_;
 wire _06826_;
 wire _06827_;
 wire _06828_;
 wire _06829_;
 wire _06830_;
 wire _06831_;
 wire _06832_;
 wire _06833_;
 wire _06834_;
 wire _06835_;
 wire _06836_;
 wire _06837_;
 wire _06838_;
 wire _06839_;
 wire _06840_;
 wire _06841_;
 wire _06842_;
 wire _06843_;
 wire _06844_;
 wire _06845_;
 wire _06846_;
 wire _06847_;
 wire _06848_;
 wire _06849_;
 wire _06850_;
 wire _06851_;
 wire _06852_;
 wire _06853_;
 wire _06854_;
 wire _06855_;
 wire _06856_;
 wire _06857_;
 wire _06858_;
 wire _06859_;
 wire _06860_;
 wire _06861_;
 wire _06862_;
 wire _06863_;
 wire _06864_;
 wire _06865_;
 wire _06866_;
 wire _06867_;
 wire _06868_;
 wire _06869_;
 wire _06870_;
 wire _06871_;
 wire _06872_;
 wire _06873_;
 wire _06874_;
 wire _06875_;
 wire _06876_;
 wire _06877_;
 wire _06878_;
 wire _06879_;
 wire _06880_;
 wire _06881_;
 wire _06882_;
 wire _06883_;
 wire _06884_;
 wire _06885_;
 wire _06886_;
 wire _06887_;
 wire _06888_;
 wire _06889_;
 wire _06890_;
 wire _06891_;
 wire _06892_;
 wire _06893_;
 wire _06894_;
 wire _06895_;
 wire _06896_;
 wire _06897_;
 wire _06898_;
 wire _06899_;
 wire _06900_;
 wire _06901_;
 wire _06902_;
 wire _06903_;
 wire _06904_;
 wire _06905_;
 wire _06906_;
 wire _06907_;
 wire _06908_;
 wire _06909_;
 wire _06910_;
 wire _06911_;
 wire _06912_;
 wire _06913_;
 wire _06914_;
 wire _06915_;
 wire _06916_;
 wire _06917_;
 wire _06918_;
 wire _06919_;
 wire _06920_;
 wire _06921_;
 wire _06922_;
 wire _06923_;
 wire _06924_;
 wire _06925_;
 wire _06926_;
 wire _06927_;
 wire _06928_;
 wire _06929_;
 wire _06930_;
 wire _06931_;
 wire _06932_;
 wire _06933_;
 wire _06934_;
 wire _06935_;
 wire _06936_;
 wire _06937_;
 wire _06938_;
 wire _06939_;
 wire _06940_;
 wire _06941_;
 wire _06942_;
 wire _06943_;
 wire _06944_;
 wire _06945_;
 wire _06946_;
 wire _06947_;
 wire _06948_;
 wire _06949_;
 wire _06950_;
 wire _06951_;
 wire _06952_;
 wire _06953_;
 wire _06954_;
 wire _06955_;
 wire _06956_;
 wire _06957_;
 wire _06958_;
 wire _06959_;
 wire _06960_;
 wire _06961_;
 wire _06962_;
 wire _06963_;
 wire _06964_;
 wire _06965_;
 wire _06966_;
 wire _06967_;
 wire _06968_;
 wire _06969_;
 wire _06970_;
 wire _06971_;
 wire _06972_;
 wire _06973_;
 wire _06974_;
 wire _06975_;
 wire _06976_;
 wire _06977_;
 wire _06978_;
 wire _06979_;
 wire _06980_;
 wire _06981_;
 wire _06982_;
 wire _06983_;
 wire _06984_;
 wire _06985_;
 wire _06986_;
 wire _06987_;
 wire _06988_;
 wire _06989_;
 wire _06990_;
 wire _06991_;
 wire _06992_;
 wire _06993_;
 wire _06994_;
 wire _06995_;
 wire _06996_;
 wire _06997_;
 wire _06998_;
 wire _06999_;
 wire _07000_;
 wire _07001_;
 wire _07002_;
 wire _07003_;
 wire _07004_;
 wire _07005_;
 wire _07006_;
 wire _07007_;
 wire _07008_;
 wire _07009_;
 wire _07010_;
 wire _07011_;
 wire _07012_;
 wire _07013_;
 wire _07014_;
 wire _07015_;
 wire _07016_;
 wire _07017_;
 wire _07018_;
 wire _07019_;
 wire _07020_;
 wire _07021_;
 wire _07022_;
 wire _07023_;
 wire _07024_;
 wire _07025_;
 wire _07026_;
 wire _07027_;
 wire _07028_;
 wire _07029_;
 wire _07030_;
 wire _07031_;
 wire _07032_;
 wire _07033_;
 wire _07034_;
 wire _07035_;
 wire _07036_;
 wire _07037_;
 wire _07038_;
 wire _07039_;
 wire _07040_;
 wire _07041_;
 wire _07042_;
 wire _07043_;
 wire _07044_;
 wire _07045_;
 wire _07046_;
 wire _07047_;
 wire _07048_;
 wire _07049_;
 wire _07050_;
 wire _07051_;
 wire _07052_;
 wire _07053_;
 wire _07054_;
 wire _07055_;
 wire _07056_;
 wire _07057_;
 wire _07058_;
 wire _07059_;
 wire _07060_;
 wire _07061_;
 wire _07062_;
 wire _07063_;
 wire _07064_;
 wire _07065_;
 wire _07066_;
 wire _07067_;
 wire _07068_;
 wire _07069_;
 wire _07070_;
 wire _07071_;
 wire _07072_;
 wire _07073_;
 wire _07074_;
 wire _07075_;
 wire _07076_;
 wire _07077_;
 wire _07078_;
 wire _07079_;
 wire _07080_;
 wire _07081_;
 wire _07082_;
 wire _07083_;
 wire _07084_;
 wire _07085_;
 wire _07086_;
 wire _07087_;
 wire _07088_;
 wire _07089_;
 wire _07090_;
 wire _07091_;
 wire _07092_;
 wire _07093_;
 wire _07094_;
 wire _07095_;
 wire _07096_;
 wire _07097_;
 wire _07098_;
 wire _07099_;
 wire _07100_;
 wire _07101_;
 wire _07102_;
 wire _07103_;
 wire _07104_;
 wire _07105_;
 wire _07106_;
 wire _07107_;
 wire _07108_;
 wire _07109_;
 wire _07110_;
 wire _07111_;
 wire _07112_;
 wire _07113_;
 wire _07114_;
 wire _07115_;
 wire _07116_;
 wire _07117_;
 wire _07118_;
 wire _07119_;
 wire _07120_;
 wire _07121_;
 wire _07122_;
 wire _07123_;
 wire _07124_;
 wire _07125_;
 wire _07126_;
 wire _07127_;
 wire _07128_;
 wire _07129_;
 wire _07130_;
 wire _07131_;
 wire _07132_;
 wire _07133_;
 wire _07134_;
 wire _07135_;
 wire _07136_;
 wire _07137_;
 wire _07138_;
 wire _07139_;
 wire _07140_;
 wire _07141_;
 wire _07142_;
 wire _07143_;
 wire _07144_;
 wire _07145_;
 wire _07146_;
 wire _07147_;
 wire _07148_;
 wire _07149_;
 wire _07150_;
 wire _07151_;
 wire _07152_;
 wire _07153_;
 wire _07154_;
 wire _07155_;
 wire _07156_;
 wire _07157_;
 wire _07158_;
 wire _07159_;
 wire _07160_;
 wire _07161_;
 wire _07162_;
 wire _07163_;
 wire _07164_;
 wire _07165_;
 wire _07166_;
 wire _07167_;
 wire _07168_;
 wire _07169_;
 wire _07170_;
 wire _07171_;
 wire _07172_;
 wire _07173_;
 wire _07174_;
 wire _07175_;
 wire _07176_;
 wire _07177_;
 wire _07178_;
 wire _07179_;
 wire _07180_;
 wire _07181_;
 wire _07182_;
 wire _07183_;
 wire _07184_;
 wire _07185_;
 wire _07186_;
 wire _07187_;
 wire _07188_;
 wire _07189_;
 wire _07190_;
 wire _07191_;
 wire _07192_;
 wire _07193_;
 wire _07194_;
 wire _07195_;
 wire _07196_;
 wire _07197_;
 wire _07198_;
 wire _07199_;
 wire _07200_;
 wire _07201_;
 wire _07202_;
 wire _07203_;
 wire _07204_;
 wire _07205_;
 wire _07206_;
 wire _07207_;
 wire _07208_;
 wire _07209_;
 wire _07210_;
 wire _07211_;
 wire _07212_;
 wire _07213_;
 wire _07214_;
 wire _07215_;
 wire _07216_;
 wire _07217_;
 wire _07218_;
 wire _07219_;
 wire _07220_;
 wire _07221_;
 wire _07222_;
 wire _07223_;
 wire _07224_;
 wire _07225_;
 wire _07226_;
 wire _07227_;
 wire _07228_;
 wire _07229_;
 wire _07230_;
 wire _07231_;
 wire _07232_;
 wire _07233_;
 wire _07234_;
 wire _07235_;
 wire _07236_;
 wire _07237_;
 wire _07238_;
 wire _07239_;
 wire _07240_;
 wire _07241_;
 wire _07242_;
 wire _07243_;
 wire _07244_;
 wire _07245_;
 wire _07246_;
 wire _07247_;
 wire _07248_;
 wire _07249_;
 wire _07250_;
 wire _07251_;
 wire _07252_;
 wire _07253_;
 wire _07254_;
 wire _07255_;
 wire _07256_;
 wire _07257_;
 wire _07258_;
 wire _07259_;
 wire _07260_;
 wire _07261_;
 wire _07262_;
 wire _07263_;
 wire _07264_;
 wire _07265_;
 wire _07266_;
 wire _07267_;
 wire _07268_;
 wire _07269_;
 wire _07270_;
 wire _07271_;
 wire _07272_;
 wire _07273_;
 wire _07274_;
 wire _07275_;
 wire _07276_;
 wire _07277_;
 wire _07278_;
 wire _07279_;
 wire _07280_;
 wire _07281_;
 wire _07282_;
 wire _07283_;
 wire _07284_;
 wire _07285_;
 wire _07286_;
 wire _07287_;
 wire _07288_;
 wire _07289_;
 wire _07290_;
 wire _07291_;
 wire _07292_;
 wire _07293_;
 wire _07294_;
 wire _07295_;
 wire _07296_;
 wire _07297_;
 wire _07298_;
 wire _07299_;
 wire _07300_;
 wire _07301_;
 wire _07302_;
 wire _07303_;
 wire _07304_;
 wire _07305_;
 wire _07306_;
 wire _07307_;
 wire _07308_;
 wire _07309_;
 wire _07310_;
 wire _07311_;
 wire _07312_;
 wire _07313_;
 wire _07314_;
 wire _07315_;
 wire _07316_;
 wire _07317_;
 wire _07318_;
 wire _07319_;
 wire _07320_;
 wire _07321_;
 wire _07322_;
 wire _07323_;
 wire _07324_;
 wire _07325_;
 wire _07326_;
 wire _07327_;
 wire _07328_;
 wire _07329_;
 wire _07330_;
 wire _07331_;
 wire _07332_;
 wire _07333_;
 wire _07334_;
 wire _07335_;
 wire _07336_;
 wire _07337_;
 wire _07338_;
 wire _07339_;
 wire _07340_;
 wire _07341_;
 wire _07342_;
 wire _07343_;
 wire _07344_;
 wire _07345_;
 wire _07346_;
 wire _07347_;
 wire _07348_;
 wire _07349_;
 wire _07350_;
 wire _07351_;
 wire _07352_;
 wire _07353_;
 wire _07354_;
 wire _07355_;
 wire _07356_;
 wire _07357_;
 wire _07358_;
 wire _07359_;
 wire _07360_;
 wire _07361_;
 wire _07362_;
 wire _07363_;
 wire _07364_;
 wire _07365_;
 wire _07366_;
 wire _07367_;
 wire _07368_;
 wire _07369_;
 wire _07370_;
 wire _07371_;
 wire _07372_;
 wire _07373_;
 wire _07374_;
 wire _07375_;
 wire _07376_;
 wire _07377_;
 wire _07378_;
 wire _07379_;
 wire _07380_;
 wire _07381_;
 wire _07382_;
 wire _07383_;
 wire _07384_;
 wire _07385_;
 wire _07386_;
 wire _07387_;
 wire _07388_;
 wire _07389_;
 wire _07390_;
 wire _07391_;
 wire _07392_;
 wire _07393_;
 wire _07394_;
 wire _07395_;
 wire _07396_;
 wire _07397_;
 wire _07398_;
 wire _07399_;
 wire _07400_;
 wire _07401_;
 wire _07402_;
 wire _07403_;
 wire _07404_;
 wire _07405_;
 wire _07406_;
 wire _07407_;
 wire _07408_;
 wire _07409_;
 wire _07410_;
 wire _07411_;
 wire _07412_;
 wire _07413_;
 wire _07414_;
 wire _07415_;
 wire _07416_;
 wire _07417_;
 wire _07418_;
 wire _07419_;
 wire _07420_;
 wire _07421_;
 wire _07422_;
 wire _07423_;
 wire _07424_;
 wire _07425_;
 wire _07426_;
 wire _07427_;
 wire _07428_;
 wire _07429_;
 wire _07430_;
 wire _07431_;
 wire _07432_;
 wire _07433_;
 wire _07434_;
 wire _07435_;
 wire _07436_;
 wire _07437_;
 wire _07438_;
 wire _07439_;
 wire _07440_;
 wire _07441_;
 wire _07442_;
 wire _07443_;
 wire _07444_;
 wire _07445_;
 wire _07446_;
 wire _07447_;
 wire _07448_;
 wire _07449_;
 wire _07450_;
 wire _07451_;
 wire _07452_;
 wire _07453_;
 wire _07454_;
 wire _07455_;
 wire _07456_;
 wire _07457_;
 wire _07458_;
 wire _07459_;
 wire _07460_;
 wire _07461_;
 wire _07462_;
 wire _07463_;
 wire _07464_;
 wire _07465_;
 wire _07466_;
 wire _07467_;
 wire _07468_;
 wire _07469_;
 wire _07470_;
 wire _07471_;
 wire _07472_;
 wire _07473_;
 wire _07474_;
 wire _07475_;
 wire _07476_;
 wire _07477_;
 wire _07478_;
 wire _07479_;
 wire _07480_;
 wire _07481_;
 wire _07482_;
 wire _07483_;
 wire _07484_;
 wire _07485_;
 wire _07486_;
 wire _07487_;
 wire _07488_;
 wire _07489_;
 wire _07490_;
 wire _07491_;
 wire _07492_;
 wire _07493_;
 wire _07494_;
 wire _07495_;
 wire _07496_;
 wire _07497_;
 wire _07498_;
 wire _07499_;
 wire _07500_;
 wire _07501_;
 wire _07502_;
 wire _07503_;
 wire _07504_;
 wire _07505_;
 wire _07506_;
 wire _07507_;
 wire _07508_;
 wire _07509_;
 wire _07510_;
 wire _07511_;
 wire _07512_;
 wire _07513_;
 wire _07514_;
 wire _07515_;
 wire _07516_;
 wire _07517_;
 wire _07518_;
 wire _07519_;
 wire _07520_;
 wire _07521_;
 wire _07522_;
 wire _07523_;
 wire _07524_;
 wire _07525_;
 wire _07526_;
 wire _07527_;
 wire _07528_;
 wire _07529_;
 wire _07530_;
 wire _07531_;
 wire _07532_;
 wire _07533_;
 wire _07534_;
 wire _07535_;
 wire _07536_;
 wire _07537_;
 wire _07538_;
 wire _07539_;
 wire _07540_;
 wire _07541_;
 wire _07542_;
 wire _07543_;
 wire _07544_;
 wire _07545_;
 wire _07546_;
 wire _07547_;
 wire _07548_;
 wire _07549_;
 wire _07550_;
 wire _07551_;
 wire _07552_;
 wire _07553_;
 wire _07554_;
 wire _07555_;
 wire _07556_;
 wire _07557_;
 wire _07558_;
 wire _07559_;
 wire _07560_;
 wire _07561_;
 wire _07562_;
 wire _07563_;
 wire _07564_;
 wire _07565_;
 wire _07566_;
 wire _07567_;
 wire _07568_;
 wire _07569_;
 wire _07570_;
 wire _07571_;
 wire _07572_;
 wire _07573_;
 wire _07574_;
 wire _07575_;
 wire _07576_;
 wire _07577_;
 wire _07578_;
 wire _07579_;
 wire _07580_;
 wire _07581_;
 wire _07582_;
 wire _07583_;
 wire _07584_;
 wire _07585_;
 wire _07586_;
 wire _07587_;
 wire _07588_;
 wire _07589_;
 wire _07590_;
 wire _07591_;
 wire _07592_;
 wire _07593_;
 wire _07594_;
 wire _07595_;
 wire _07596_;
 wire _07597_;
 wire _07598_;
 wire _07599_;
 wire _07600_;
 wire _07601_;
 wire _07602_;
 wire _07603_;
 wire _07604_;
 wire _07605_;
 wire _07606_;
 wire _07607_;
 wire _07608_;
 wire _07609_;
 wire _07610_;
 wire _07611_;
 wire _07612_;
 wire _07613_;
 wire _07614_;
 wire _07615_;
 wire _07616_;
 wire _07617_;
 wire _07618_;
 wire _07619_;
 wire _07620_;
 wire _07621_;
 wire _07622_;
 wire _07623_;
 wire _07624_;
 wire _07625_;
 wire _07626_;
 wire _07627_;
 wire _07628_;
 wire _07629_;
 wire _07630_;
 wire _07631_;
 wire _07632_;
 wire _07633_;
 wire _07634_;
 wire _07635_;
 wire _07636_;
 wire _07637_;
 wire _07638_;
 wire _07639_;
 wire _07640_;
 wire _07641_;
 wire _07642_;
 wire _07643_;
 wire _07644_;
 wire _07645_;
 wire _07646_;
 wire _07647_;
 wire _07648_;
 wire _07649_;
 wire _07650_;
 wire _07651_;
 wire _07652_;
 wire _07653_;
 wire _07654_;
 wire _07655_;
 wire _07656_;
 wire _07657_;
 wire _07658_;
 wire _07659_;
 wire _07660_;
 wire _07661_;
 wire _07662_;
 wire _07663_;
 wire _07664_;
 wire _07665_;
 wire _07666_;
 wire _07667_;
 wire _07668_;
 wire _07669_;
 wire _07670_;
 wire _07671_;
 wire _07672_;
 wire _07673_;
 wire _07674_;
 wire _07675_;
 wire _07676_;
 wire _07677_;
 wire _07678_;
 wire _07679_;
 wire _07680_;
 wire _07681_;
 wire _07682_;
 wire _07683_;
 wire _07684_;
 wire _07685_;
 wire _07686_;
 wire _07687_;
 wire _07688_;
 wire _07689_;
 wire _07690_;
 wire _07691_;
 wire _07692_;
 wire _07693_;
 wire _07694_;
 wire _07695_;
 wire _07696_;
 wire _07697_;
 wire _07698_;
 wire _07699_;
 wire _07700_;
 wire _07701_;
 wire _07702_;
 wire _07703_;
 wire _07704_;
 wire _07705_;
 wire _07706_;
 wire _07707_;
 wire _07708_;
 wire _07709_;
 wire _07710_;
 wire _07711_;
 wire _07712_;
 wire _07713_;
 wire _07714_;
 wire _07715_;
 wire _07716_;
 wire _07717_;
 wire _07718_;
 wire _07719_;
 wire _07720_;
 wire _07721_;
 wire _07722_;
 wire _07723_;
 wire _07724_;
 wire _07725_;
 wire _07726_;
 wire _07727_;
 wire _07728_;
 wire _07729_;
 wire _07730_;
 wire _07731_;
 wire _07732_;
 wire _07733_;
 wire _07734_;
 wire _07735_;
 wire _07736_;
 wire _07737_;
 wire _07738_;
 wire _07739_;
 wire _07740_;
 wire _07741_;
 wire _07742_;
 wire _07743_;
 wire _07744_;
 wire _07745_;
 wire _07746_;
 wire _07747_;
 wire _07748_;
 wire _07749_;
 wire _07750_;
 wire _07751_;
 wire _07752_;
 wire _07753_;
 wire _07754_;
 wire _07755_;
 wire _07756_;
 wire _07757_;
 wire _07758_;
 wire _07759_;
 wire _07760_;
 wire _07761_;
 wire _07762_;
 wire _07763_;
 wire _07764_;
 wire _07765_;
 wire _07766_;
 wire _07767_;
 wire _07768_;
 wire _07769_;
 wire _07770_;
 wire _07771_;
 wire _07772_;
 wire _07773_;
 wire _07774_;
 wire _07775_;
 wire _07776_;
 wire _07777_;
 wire _07778_;
 wire _07779_;
 wire _07780_;
 wire _07781_;
 wire _07782_;
 wire _07783_;
 wire _07784_;
 wire _07785_;
 wire _07786_;
 wire _07787_;
 wire _07788_;
 wire _07789_;
 wire _07790_;
 wire _07791_;
 wire _07792_;
 wire _07793_;
 wire _07794_;
 wire _07795_;
 wire _07796_;
 wire _07797_;
 wire _07798_;
 wire _07799_;
 wire _07800_;
 wire _07801_;
 wire _07802_;
 wire _07803_;
 wire _07804_;
 wire _07805_;
 wire _07806_;
 wire _07807_;
 wire _07808_;
 wire _07809_;
 wire _07810_;
 wire _07811_;
 wire _07812_;
 wire _07813_;
 wire _07814_;
 wire _07815_;
 wire _07816_;
 wire _07817_;
 wire _07818_;
 wire _07819_;
 wire _07820_;
 wire _07821_;
 wire _07822_;
 wire _07823_;
 wire _07824_;
 wire _07825_;
 wire _07826_;
 wire _07827_;
 wire _07828_;
 wire _07829_;
 wire _07830_;
 wire _07831_;
 wire _07832_;
 wire _07833_;
 wire _07834_;
 wire _07835_;
 wire _07836_;
 wire _07837_;
 wire _07838_;
 wire _07839_;
 wire _07840_;
 wire _07841_;
 wire _07842_;
 wire _07843_;
 wire _07844_;
 wire _07845_;
 wire _07846_;
 wire _07847_;
 wire _07848_;
 wire _07849_;
 wire _07850_;
 wire _07851_;
 wire _07852_;
 wire _07853_;
 wire _07854_;
 wire _07855_;
 wire _07856_;
 wire _07857_;
 wire _07858_;
 wire _07859_;
 wire _07860_;
 wire _07861_;
 wire _07862_;
 wire _07863_;
 wire _07864_;
 wire _07865_;
 wire _07866_;
 wire _07867_;
 wire _07868_;
 wire _07869_;
 wire _07870_;
 wire _07871_;
 wire _07872_;
 wire _07873_;
 wire _07874_;
 wire _07875_;
 wire _07876_;
 wire _07877_;
 wire _07878_;
 wire _07879_;
 wire _07880_;
 wire _07881_;
 wire _07882_;
 wire _07883_;
 wire _07884_;
 wire _07885_;
 wire _07886_;
 wire _07887_;
 wire _07888_;
 wire _07889_;
 wire _07890_;
 wire _07891_;
 wire _07892_;
 wire _07893_;
 wire _07894_;
 wire _07895_;
 wire _07896_;
 wire _07897_;
 wire _07898_;
 wire _07899_;
 wire _07900_;
 wire _07901_;
 wire _07902_;
 wire _07903_;
 wire _07904_;
 wire _07905_;
 wire _07906_;
 wire _07907_;
 wire _07908_;
 wire _07909_;
 wire _07910_;
 wire _07911_;
 wire _07912_;
 wire _07913_;
 wire _07914_;
 wire _07915_;
 wire _07916_;
 wire _07917_;
 wire _07918_;
 wire _07919_;
 wire _07920_;
 wire _07921_;
 wire _07922_;
 wire _07923_;
 wire _07924_;
 wire _07925_;
 wire _07926_;
 wire _07927_;
 wire _07928_;
 wire _07929_;
 wire _07930_;
 wire _07931_;
 wire _07932_;
 wire _07933_;
 wire _07934_;
 wire _07935_;
 wire _07936_;
 wire _07937_;
 wire _07938_;
 wire _07939_;
 wire _07940_;
 wire _07941_;
 wire _07942_;
 wire _07943_;
 wire _07944_;
 wire _07945_;
 wire _07946_;
 wire _07947_;
 wire _07948_;
 wire _07949_;
 wire _07950_;
 wire _07951_;
 wire _07952_;
 wire _07953_;
 wire _07954_;
 wire _07955_;
 wire _07956_;
 wire _07957_;
 wire _07958_;
 wire _07959_;
 wire _07960_;
 wire _07961_;
 wire _07962_;
 wire _07963_;
 wire _07964_;
 wire _07965_;
 wire _07966_;
 wire _07967_;
 wire _07968_;
 wire _07969_;
 wire _07970_;
 wire _07971_;
 wire _07972_;
 wire _07973_;
 wire _07974_;
 wire _07975_;
 wire _07976_;
 wire _07977_;
 wire _07978_;
 wire _07979_;
 wire _07980_;
 wire _07981_;
 wire _07982_;
 wire _07983_;
 wire _07984_;
 wire _07985_;
 wire _07986_;
 wire _07987_;
 wire _07988_;
 wire _07989_;
 wire _07990_;
 wire _07991_;
 wire _07992_;
 wire _07993_;
 wire _07994_;
 wire _07995_;
 wire _07996_;
 wire _07997_;
 wire _07998_;
 wire _07999_;
 wire _08000_;
 wire _08001_;
 wire _08002_;
 wire _08003_;
 wire _08004_;
 wire _08005_;
 wire _08006_;
 wire _08007_;
 wire _08008_;
 wire _08009_;
 wire _08010_;
 wire _08011_;
 wire _08012_;
 wire _08013_;
 wire _08014_;
 wire _08015_;
 wire _08016_;
 wire _08017_;
 wire _08018_;
 wire _08019_;
 wire _08020_;
 wire _08021_;
 wire _08022_;
 wire _08023_;
 wire _08024_;
 wire _08025_;
 wire _08026_;
 wire _08027_;
 wire _08028_;
 wire _08029_;
 wire _08030_;
 wire _08031_;
 wire _08032_;
 wire _08033_;
 wire _08034_;
 wire _08035_;
 wire _08036_;
 wire _08037_;
 wire _08038_;
 wire _08039_;
 wire _08040_;
 wire _08041_;
 wire _08042_;
 wire _08043_;
 wire _08044_;
 wire _08045_;
 wire _08046_;
 wire _08047_;
 wire _08048_;
 wire _08049_;
 wire _08050_;
 wire _08051_;
 wire _08052_;
 wire _08053_;
 wire _08054_;
 wire _08055_;
 wire _08056_;
 wire _08057_;
 wire _08058_;
 wire _08059_;
 wire _08060_;
 wire _08061_;
 wire _08062_;
 wire _08063_;
 wire _08064_;
 wire _08065_;
 wire _08066_;
 wire _08067_;
 wire _08068_;
 wire _08069_;
 wire _08070_;
 wire _08071_;
 wire _08072_;
 wire _08073_;
 wire _08074_;
 wire _08075_;
 wire _08076_;
 wire _08077_;
 wire _08078_;
 wire _08079_;
 wire _08080_;
 wire _08081_;
 wire _08082_;
 wire _08083_;
 wire _08084_;
 wire _08085_;
 wire _08086_;
 wire _08087_;
 wire _08088_;
 wire _08089_;
 wire _08090_;
 wire _08091_;
 wire _08092_;
 wire _08093_;
 wire _08094_;
 wire _08095_;
 wire _08096_;
 wire _08097_;
 wire _08098_;
 wire _08099_;
 wire _08100_;
 wire _08101_;
 wire _08102_;
 wire _08103_;
 wire _08104_;
 wire _08105_;
 wire _08106_;
 wire _08107_;
 wire _08108_;
 wire _08109_;
 wire _08110_;
 wire _08111_;
 wire _08112_;
 wire _08113_;
 wire _08114_;
 wire _08115_;
 wire _08116_;
 wire _08117_;
 wire _08118_;
 wire _08119_;
 wire _08120_;
 wire _08121_;
 wire _08122_;
 wire _08123_;
 wire _08124_;
 wire _08125_;
 wire _08126_;
 wire _08127_;
 wire _08128_;
 wire _08129_;
 wire _08130_;
 wire _08131_;
 wire _08132_;
 wire _08133_;
 wire _08134_;
 wire _08135_;
 wire _08136_;
 wire _08137_;
 wire _08138_;
 wire _08139_;
 wire _08140_;
 wire _08141_;
 wire _08142_;
 wire _08143_;
 wire _08144_;
 wire _08145_;
 wire _08146_;
 wire _08147_;
 wire _08148_;
 wire _08149_;
 wire _08150_;
 wire _08151_;
 wire _08152_;
 wire _08153_;
 wire _08154_;
 wire _08155_;
 wire _08156_;
 wire _08157_;
 wire _08158_;
 wire _08159_;
 wire _08160_;
 wire _08161_;
 wire _08162_;
 wire _08163_;
 wire _08164_;
 wire _08165_;
 wire _08166_;
 wire _08167_;
 wire _08168_;
 wire _08169_;
 wire _08170_;
 wire _08171_;
 wire _08172_;
 wire _08173_;
 wire _08174_;
 wire _08175_;
 wire _08176_;
 wire _08177_;
 wire _08178_;
 wire _08179_;
 wire _08180_;
 wire _08181_;
 wire _08182_;
 wire _08183_;
 wire _08184_;
 wire _08185_;
 wire _08186_;
 wire _08187_;
 wire _08188_;
 wire _08189_;
 wire _08190_;
 wire _08191_;
 wire _08192_;
 wire _08193_;
 wire _08194_;
 wire _08195_;
 wire _08196_;
 wire _08197_;
 wire _08198_;
 wire _08199_;
 wire _08200_;
 wire _08201_;
 wire _08202_;
 wire _08203_;
 wire _08204_;
 wire _08205_;
 wire _08206_;
 wire _08207_;
 wire _08208_;
 wire _08209_;
 wire _08210_;
 wire _08211_;
 wire _08212_;
 wire _08213_;
 wire _08214_;
 wire _08215_;
 wire _08216_;
 wire _08217_;
 wire _08218_;
 wire _08219_;
 wire _08220_;
 wire _08221_;
 wire _08222_;
 wire _08223_;
 wire _08224_;
 wire _08225_;
 wire _08226_;
 wire _08227_;
 wire _08228_;
 wire _08229_;
 wire _08230_;
 wire _08231_;
 wire _08232_;
 wire _08233_;
 wire _08234_;
 wire _08235_;
 wire _08236_;
 wire _08237_;
 wire _08238_;
 wire _08239_;
 wire _08240_;
 wire _08241_;
 wire _08242_;
 wire _08243_;
 wire _08244_;
 wire _08245_;
 wire _08246_;
 wire _08247_;
 wire _08248_;
 wire _08249_;
 wire _08250_;
 wire _08251_;
 wire _08252_;
 wire _08253_;
 wire _08254_;
 wire _08255_;
 wire _08256_;
 wire _08257_;
 wire _08258_;
 wire _08259_;
 wire _08260_;
 wire _08261_;
 wire _08262_;
 wire _08263_;
 wire _08264_;
 wire _08265_;
 wire _08266_;
 wire _08267_;
 wire _08268_;
 wire _08269_;
 wire _08270_;
 wire _08271_;
 wire _08272_;
 wire _08273_;
 wire _08274_;
 wire _08275_;
 wire _08276_;
 wire _08277_;
 wire _08278_;
 wire _08279_;
 wire _08280_;
 wire _08281_;
 wire _08282_;
 wire _08283_;
 wire _08284_;
 wire _08285_;
 wire _08286_;
 wire _08287_;
 wire _08288_;
 wire _08289_;
 wire _08290_;
 wire _08291_;
 wire _08292_;
 wire _08293_;
 wire _08294_;
 wire _08295_;
 wire _08296_;
 wire _08297_;
 wire _08298_;
 wire _08299_;
 wire _08300_;
 wire _08301_;
 wire _08302_;
 wire _08303_;
 wire _08304_;
 wire _08305_;
 wire _08306_;
 wire _08307_;
 wire _08308_;
 wire _08309_;
 wire _08310_;
 wire _08311_;
 wire _08312_;
 wire _08313_;
 wire _08314_;
 wire _08315_;
 wire _08316_;
 wire _08317_;
 wire _08318_;
 wire _08319_;
 wire _08320_;
 wire _08321_;
 wire _08322_;
 wire _08323_;
 wire _08324_;
 wire _08325_;
 wire _08326_;
 wire _08327_;
 wire _08328_;
 wire _08329_;
 wire _08330_;
 wire _08331_;
 wire _08332_;
 wire _08333_;
 wire _08334_;
 wire _08335_;
 wire _08336_;
 wire _08337_;
 wire _08338_;
 wire _08339_;
 wire _08340_;
 wire _08341_;
 wire _08342_;
 wire _08343_;
 wire _08344_;
 wire _08345_;
 wire _08346_;
 wire _08347_;
 wire _08348_;
 wire _08349_;
 wire _08350_;
 wire _08351_;
 wire _08352_;
 wire _08353_;
 wire _08354_;
 wire _08355_;
 wire _08356_;
 wire _08357_;
 wire _08358_;
 wire _08359_;
 wire _08360_;
 wire _08361_;
 wire _08362_;
 wire _08363_;
 wire _08364_;
 wire _08365_;
 wire _08366_;
 wire _08367_;
 wire _08368_;
 wire _08369_;
 wire _08370_;
 wire _08371_;
 wire _08372_;
 wire _08373_;
 wire _08374_;
 wire _08375_;
 wire _08376_;
 wire _08377_;
 wire _08378_;
 wire _08379_;
 wire _08380_;
 wire _08381_;
 wire _08382_;
 wire _08383_;
 wire _08384_;
 wire _08385_;
 wire _08386_;
 wire _08387_;
 wire _08388_;
 wire _08389_;
 wire _08390_;
 wire _08391_;
 wire _08392_;
 wire _08393_;
 wire _08394_;
 wire _08395_;
 wire _08396_;
 wire _08397_;
 wire _08398_;
 wire _08399_;
 wire _08400_;
 wire _08401_;
 wire _08402_;
 wire _08403_;
 wire _08404_;
 wire _08405_;
 wire _08406_;
 wire _08407_;
 wire _08408_;
 wire _08409_;
 wire _08410_;
 wire _08411_;
 wire _08412_;
 wire _08413_;
 wire _08414_;
 wire _08415_;
 wire _08416_;
 wire _08417_;
 wire _08418_;
 wire _08419_;
 wire _08420_;
 wire _08421_;
 wire _08422_;
 wire _08423_;
 wire _08424_;
 wire _08425_;
 wire _08426_;
 wire _08427_;
 wire _08428_;
 wire _08429_;
 wire _08430_;
 wire _08431_;
 wire _08432_;
 wire _08433_;
 wire _08434_;
 wire _08435_;
 wire _08436_;
 wire _08437_;
 wire _08438_;
 wire _08439_;
 wire _08440_;
 wire _08441_;
 wire _08442_;
 wire _08443_;
 wire _08444_;
 wire _08445_;
 wire _08446_;
 wire _08447_;
 wire _08448_;
 wire _08449_;
 wire _08450_;
 wire _08451_;
 wire _08452_;
 wire _08453_;
 wire _08454_;
 wire _08455_;
 wire _08456_;
 wire _08457_;
 wire _08458_;
 wire _08459_;
 wire _08460_;
 wire _08461_;
 wire _08462_;
 wire _08463_;
 wire _08464_;
 wire _08465_;
 wire _08466_;
 wire _08467_;
 wire _08468_;
 wire _08469_;
 wire _08470_;
 wire _08471_;
 wire _08472_;
 wire _08473_;
 wire _08474_;
 wire _08475_;
 wire _08476_;
 wire _08477_;
 wire _08478_;
 wire _08479_;
 wire _08480_;
 wire _08481_;
 wire _08482_;
 wire _08483_;
 wire _08484_;
 wire _08485_;
 wire _08486_;
 wire _08487_;
 wire _08488_;
 wire _08489_;
 wire _08490_;
 wire _08491_;
 wire _08492_;
 wire _08493_;
 wire _08494_;
 wire _08495_;
 wire _08496_;
 wire _08497_;
 wire _08498_;
 wire _08499_;
 wire _08500_;
 wire _08501_;
 wire _08502_;
 wire _08503_;
 wire _08504_;
 wire _08505_;
 wire _08506_;
 wire _08507_;
 wire _08508_;
 wire _08509_;
 wire _08510_;
 wire _08511_;
 wire _08512_;
 wire _08513_;
 wire _08514_;
 wire _08515_;
 wire _08516_;
 wire _08517_;
 wire _08518_;
 wire _08519_;
 wire _08520_;
 wire _08521_;
 wire _08522_;
 wire _08523_;
 wire _08524_;
 wire _08525_;
 wire _08526_;
 wire _08527_;
 wire _08528_;
 wire _08529_;
 wire _08530_;
 wire _08531_;
 wire _08532_;
 wire _08533_;
 wire _08534_;
 wire _08535_;
 wire _08536_;
 wire _08537_;
 wire _08538_;
 wire _08539_;
 wire _08540_;
 wire _08541_;
 wire _08542_;
 wire _08543_;
 wire _08544_;
 wire _08545_;
 wire _08546_;
 wire _08547_;
 wire _08548_;
 wire _08549_;
 wire _08550_;
 wire _08551_;
 wire _08552_;
 wire _08553_;
 wire _08554_;
 wire _08555_;
 wire _08556_;
 wire _08557_;
 wire _08558_;
 wire _08559_;
 wire _08560_;
 wire _08561_;
 wire _08562_;
 wire _08563_;
 wire _08564_;
 wire _08565_;
 wire _08566_;
 wire _08567_;
 wire _08568_;
 wire _08569_;
 wire _08570_;
 wire _08571_;
 wire _08572_;
 wire _08573_;
 wire _08574_;
 wire _08575_;
 wire _08576_;
 wire _08577_;
 wire _08578_;
 wire _08579_;
 wire _08580_;
 wire _08581_;
 wire _08582_;
 wire _08583_;
 wire _08584_;
 wire _08585_;
 wire _08586_;
 wire _08587_;
 wire _08588_;
 wire _08589_;
 wire _08590_;
 wire _08591_;
 wire _08592_;
 wire _08593_;
 wire _08594_;
 wire _08595_;
 wire _08596_;
 wire _08597_;
 wire _08598_;
 wire _08599_;
 wire _08600_;
 wire _08601_;
 wire _08602_;
 wire _08603_;
 wire _08604_;
 wire _08605_;
 wire _08606_;
 wire _08607_;
 wire _08608_;
 wire _08609_;
 wire _08610_;
 wire _08611_;
 wire _08612_;
 wire _08613_;
 wire _08614_;
 wire _08615_;
 wire _08616_;
 wire _08617_;
 wire _08618_;
 wire _08619_;
 wire _08620_;
 wire _08621_;
 wire _08622_;
 wire _08623_;
 wire _08624_;
 wire _08625_;
 wire _08626_;
 wire _08627_;
 wire _08628_;
 wire _08629_;
 wire _08630_;
 wire _08631_;
 wire _08632_;
 wire _08633_;
 wire _08634_;
 wire _08635_;
 wire _08636_;
 wire _08637_;
 wire _08638_;
 wire _08639_;
 wire _08640_;
 wire _08641_;
 wire _08642_;
 wire _08643_;
 wire _08644_;
 wire _08645_;
 wire _08646_;
 wire _08647_;
 wire _08648_;
 wire _08649_;
 wire _08650_;
 wire _08651_;
 wire _08652_;
 wire _08653_;
 wire _08654_;
 wire _08655_;
 wire _08656_;
 wire _08657_;
 wire _08658_;
 wire _08659_;
 wire _08660_;
 wire _08661_;
 wire _08662_;
 wire _08663_;
 wire _08664_;
 wire _08665_;
 wire _08666_;
 wire _08667_;
 wire _08668_;
 wire _08669_;
 wire _08670_;
 wire _08671_;
 wire _08672_;
 wire _08673_;
 wire _08674_;
 wire _08675_;
 wire _08676_;
 wire _08677_;
 wire _08678_;
 wire _08679_;
 wire _08680_;
 wire _08681_;
 wire _08682_;
 wire _08683_;
 wire _08684_;
 wire _08685_;
 wire _08686_;
 wire _08687_;
 wire _08688_;
 wire _08689_;
 wire _08690_;
 wire _08691_;
 wire _08692_;
 wire _08693_;
 wire _08694_;
 wire _08695_;
 wire _08696_;
 wire _08697_;
 wire _08698_;
 wire _08699_;
 wire _08700_;
 wire _08701_;
 wire _08702_;
 wire _08703_;
 wire _08704_;
 wire _08705_;
 wire _08706_;
 wire _08707_;
 wire _08708_;
 wire _08709_;
 wire _08710_;
 wire _08711_;
 wire _08712_;
 wire _08713_;
 wire _08714_;
 wire _08715_;
 wire _08716_;
 wire _08717_;
 wire _08718_;
 wire _08719_;
 wire _08720_;
 wire _08721_;
 wire _08722_;
 wire _08723_;
 wire _08724_;
 wire _08725_;
 wire _08726_;
 wire _08727_;
 wire _08728_;
 wire _08729_;
 wire _08730_;
 wire _08731_;
 wire _08732_;
 wire _08733_;
 wire _08734_;
 wire _08735_;
 wire _08736_;
 wire _08737_;
 wire _08738_;
 wire _08739_;
 wire _08740_;
 wire _08741_;
 wire _08742_;
 wire _08743_;
 wire _08744_;
 wire _08745_;
 wire _08746_;
 wire _08747_;
 wire _08748_;
 wire _08749_;
 wire _08750_;
 wire _08751_;
 wire _08752_;
 wire _08753_;
 wire _08754_;
 wire _08755_;
 wire _08756_;
 wire _08757_;
 wire _08758_;
 wire _08759_;
 wire _08760_;
 wire _08761_;
 wire _08762_;
 wire _08763_;
 wire _08764_;
 wire _08765_;
 wire _08766_;
 wire _08767_;
 wire _08768_;
 wire _08769_;
 wire _08770_;
 wire _08771_;
 wire _08772_;
 wire _08773_;
 wire _08774_;
 wire _08775_;
 wire _08776_;
 wire _08777_;
 wire _08778_;
 wire _08779_;
 wire _08780_;
 wire _08781_;
 wire _08782_;
 wire _08783_;
 wire _08784_;
 wire _08785_;
 wire _08786_;
 wire _08787_;
 wire _08788_;
 wire _08789_;
 wire _08790_;
 wire _08791_;
 wire _08792_;
 wire _08793_;
 wire _08794_;
 wire _08795_;
 wire _08796_;
 wire _08797_;
 wire _08798_;
 wire _08799_;
 wire _08800_;
 wire _08801_;
 wire _08802_;
 wire _08803_;
 wire _08804_;
 wire _08805_;
 wire _08806_;
 wire _08807_;
 wire _08808_;
 wire _08809_;
 wire _08810_;
 wire _08811_;
 wire _08812_;
 wire _08813_;
 wire _08814_;
 wire _08815_;
 wire _08816_;
 wire _08817_;
 wire _08818_;
 wire _08819_;
 wire _08820_;
 wire _08821_;
 wire _08822_;
 wire _08823_;
 wire _08824_;
 wire _08825_;
 wire _08826_;
 wire _08827_;
 wire _08828_;
 wire _08829_;
 wire _08830_;
 wire _08831_;
 wire _08832_;
 wire _08833_;
 wire _08834_;
 wire _08835_;
 wire _08836_;
 wire _08837_;
 wire _08838_;
 wire _08839_;
 wire _08840_;
 wire _08841_;
 wire _08842_;
 wire _08843_;
 wire _08844_;
 wire _08845_;
 wire _08846_;
 wire _08847_;
 wire _08848_;
 wire _08849_;
 wire _08850_;
 wire _08851_;
 wire _08852_;
 wire _08853_;
 wire _08854_;
 wire _08855_;
 wire _08856_;
 wire _08857_;
 wire _08858_;
 wire _08859_;
 wire _08860_;
 wire _08861_;
 wire _08862_;
 wire _08863_;
 wire _08864_;
 wire _08865_;
 wire _08866_;
 wire _08867_;
 wire _08868_;
 wire _08869_;
 wire _08870_;
 wire _08871_;
 wire _08872_;
 wire _08873_;
 wire _08874_;
 wire _08875_;
 wire _08876_;
 wire _08877_;
 wire _08878_;
 wire _08879_;
 wire _08880_;
 wire _08881_;
 wire _08882_;
 wire _08883_;
 wire _08884_;
 wire _08885_;
 wire _08886_;
 wire _08887_;
 wire _08888_;
 wire _08889_;
 wire _08890_;
 wire _08891_;
 wire _08892_;
 wire _08893_;
 wire _08894_;
 wire _08895_;
 wire _08896_;
 wire _08897_;
 wire _08898_;
 wire _08899_;
 wire _08900_;
 wire _08901_;
 wire _08902_;
 wire _08903_;
 wire _08904_;
 wire _08905_;
 wire _08906_;
 wire _08907_;
 wire _08908_;
 wire _08909_;
 wire _08910_;
 wire _08911_;
 wire _08912_;
 wire _08913_;
 wire _08914_;
 wire _08915_;
 wire _08916_;
 wire _08917_;
 wire _08918_;
 wire _08919_;
 wire _08920_;
 wire _08921_;
 wire _08922_;
 wire _08923_;
 wire _08924_;
 wire _08925_;
 wire _08926_;
 wire _08927_;
 wire _08928_;
 wire _08929_;
 wire _08930_;
 wire _08931_;
 wire _08932_;
 wire _08933_;
 wire _08934_;
 wire _08935_;
 wire _08936_;
 wire _08937_;
 wire _08938_;
 wire _08939_;
 wire _08940_;
 wire _08941_;
 wire _08942_;
 wire _08943_;
 wire _08944_;
 wire _08945_;
 wire _08946_;
 wire _08947_;
 wire _08948_;
 wire _08949_;
 wire _08950_;
 wire _08951_;
 wire _08952_;
 wire _08953_;
 wire _08954_;
 wire _08955_;
 wire _08956_;
 wire _08957_;
 wire _08958_;
 wire _08959_;
 wire _08960_;
 wire _08961_;
 wire _08962_;
 wire _08963_;
 wire _08964_;
 wire _08965_;
 wire _08966_;
 wire _08967_;
 wire _08968_;
 wire _08969_;
 wire _08970_;
 wire _08971_;
 wire _08972_;
 wire _08973_;
 wire _08974_;
 wire _08975_;
 wire _08976_;
 wire _08977_;
 wire _08978_;
 wire _08979_;
 wire _08980_;
 wire _08981_;
 wire _08982_;
 wire _08983_;
 wire _08984_;
 wire _08985_;
 wire _08986_;
 wire _08987_;
 wire _08988_;
 wire _08989_;
 wire _08990_;
 wire _08991_;
 wire _08992_;
 wire _08993_;
 wire _08994_;
 wire _08995_;
 wire _08996_;
 wire _08997_;
 wire _08998_;
 wire _08999_;
 wire _09000_;
 wire _09001_;
 wire _09002_;
 wire _09003_;
 wire _09004_;
 wire _09005_;
 wire _09006_;
 wire _09007_;
 wire _09008_;
 wire _09009_;
 wire _09010_;
 wire _09011_;
 wire _09012_;
 wire _09013_;
 wire _09014_;
 wire _09015_;
 wire _09016_;
 wire _09017_;
 wire _09018_;
 wire _09019_;
 wire _09020_;
 wire _09021_;
 wire _09022_;
 wire _09023_;
 wire _09024_;
 wire _09025_;
 wire _09026_;
 wire _09027_;
 wire _09028_;
 wire _09029_;
 wire _09030_;
 wire _09031_;
 wire _09032_;
 wire _09033_;
 wire _09034_;
 wire _09035_;
 wire _09036_;
 wire _09037_;
 wire _09038_;
 wire _09039_;
 wire _09040_;
 wire _09041_;
 wire _09042_;
 wire _09043_;
 wire _09044_;
 wire _09045_;
 wire _09046_;
 wire _09047_;
 wire _09048_;
 wire _09049_;
 wire _09050_;
 wire _09051_;
 wire _09052_;
 wire _09053_;
 wire _09054_;
 wire _09055_;
 wire _09056_;
 wire _09057_;
 wire _09058_;
 wire _09059_;
 wire _09060_;
 wire _09061_;
 wire _09062_;
 wire _09063_;
 wire _09064_;
 wire _09065_;
 wire _09066_;
 wire _09067_;
 wire _09068_;
 wire _09069_;
 wire _09070_;
 wire _09071_;
 wire _09072_;
 wire _09073_;
 wire _09074_;
 wire _09075_;
 wire _09076_;
 wire _09077_;
 wire _09078_;
 wire _09079_;
 wire _09080_;
 wire _09081_;
 wire _09082_;
 wire _09083_;
 wire _09084_;
 wire _09085_;
 wire _09086_;
 wire _09087_;
 wire _09088_;
 wire _09089_;
 wire _09090_;
 wire _09091_;
 wire _09092_;
 wire _09093_;
 wire _09094_;
 wire _09095_;
 wire _09096_;
 wire _09097_;
 wire _09098_;
 wire _09099_;
 wire _09100_;
 wire _09101_;
 wire _09102_;
 wire _09103_;
 wire _09104_;
 wire _09105_;
 wire _09106_;
 wire _09107_;
 wire _09108_;
 wire _09109_;
 wire _09110_;
 wire _09111_;
 wire _09112_;
 wire _09113_;
 wire _09114_;
 wire _09115_;
 wire _09116_;
 wire _09117_;
 wire _09118_;
 wire _09119_;
 wire _09120_;
 wire _09121_;
 wire _09122_;
 wire _09123_;
 wire _09124_;
 wire _09125_;
 wire _09126_;
 wire _09127_;
 wire _09128_;
 wire _09129_;
 wire _09130_;
 wire _09131_;
 wire _09132_;
 wire _09133_;
 wire _09134_;
 wire _09135_;
 wire _09136_;
 wire _09137_;
 wire _09138_;
 wire _09139_;
 wire _09140_;
 wire _09141_;
 wire _09142_;
 wire _09143_;
 wire _09144_;
 wire _09145_;
 wire _09146_;
 wire _09147_;
 wire _09148_;
 wire _09149_;
 wire _09150_;
 wire _09151_;
 wire _09152_;
 wire _09153_;
 wire _09154_;
 wire _09155_;
 wire _09156_;
 wire _09157_;
 wire _09158_;
 wire _09159_;
 wire _09160_;
 wire _09161_;
 wire _09162_;
 wire _09163_;
 wire _09164_;
 wire _09165_;
 wire _09166_;
 wire _09167_;
 wire _09168_;
 wire _09169_;
 wire _09170_;
 wire _09171_;
 wire _09172_;
 wire _09173_;
 wire _09174_;
 wire _09175_;
 wire _09176_;
 wire _09177_;
 wire _09178_;
 wire _09179_;
 wire _09180_;
 wire _09181_;
 wire _09182_;
 wire _09183_;
 wire _09184_;
 wire _09185_;
 wire _09186_;
 wire _09187_;
 wire _09188_;
 wire _09189_;
 wire _09190_;
 wire _09191_;
 wire _09192_;
 wire _09193_;
 wire _09194_;
 wire _09195_;
 wire _09196_;
 wire _09197_;
 wire _09198_;
 wire _09199_;
 wire _09200_;
 wire _09201_;
 wire _09202_;
 wire _09203_;
 wire _09204_;
 wire _09205_;
 wire _09206_;
 wire _09207_;
 wire _09208_;
 wire _09209_;
 wire _09210_;
 wire _09211_;
 wire _09212_;
 wire _09213_;
 wire _09214_;
 wire _09215_;
 wire _09216_;
 wire _09217_;
 wire _09218_;
 wire _09219_;
 wire _09220_;
 wire _09221_;
 wire _09222_;
 wire _09223_;
 wire _09224_;
 wire _09225_;
 wire _09226_;
 wire _09227_;
 wire _09228_;
 wire _09229_;
 wire _09230_;
 wire _09231_;
 wire _09232_;
 wire _09233_;
 wire _09234_;
 wire _09235_;
 wire _09236_;
 wire _09237_;
 wire _09238_;
 wire _09239_;
 wire _09240_;
 wire _09241_;
 wire _09242_;
 wire _09243_;
 wire _09244_;
 wire _09245_;
 wire _09246_;
 wire _09247_;
 wire _09248_;
 wire _09249_;
 wire _09250_;
 wire _09251_;
 wire _09252_;
 wire _09253_;
 wire _09254_;
 wire _09255_;
 wire _09256_;
 wire _09257_;
 wire _09258_;
 wire _09259_;
 wire _09260_;
 wire _09261_;
 wire _09262_;
 wire _09263_;
 wire _09264_;
 wire _09265_;
 wire _09266_;
 wire _09267_;
 wire _09268_;
 wire _09269_;
 wire _09270_;
 wire _09271_;
 wire _09272_;
 wire _09273_;
 wire _09274_;
 wire _09275_;
 wire _09276_;
 wire _09277_;
 wire _09278_;
 wire _09279_;
 wire _09280_;
 wire _09281_;
 wire _09282_;
 wire _09283_;
 wire _09284_;
 wire _09285_;
 wire _09286_;
 wire _09287_;
 wire _09288_;
 wire _09289_;
 wire _09290_;
 wire _09291_;
 wire _09292_;
 wire _09293_;
 wire _09294_;
 wire _09295_;
 wire _09296_;
 wire _09297_;
 wire _09298_;
 wire _09299_;
 wire _09300_;
 wire _09301_;
 wire _09302_;
 wire _09303_;
 wire _09304_;
 wire _09305_;
 wire _09306_;
 wire _09307_;
 wire _09308_;
 wire _09309_;
 wire _09310_;
 wire _09311_;
 wire _09312_;
 wire _09313_;
 wire _09314_;
 wire _09315_;
 wire _09316_;
 wire _09317_;
 wire _09318_;
 wire _09319_;
 wire _09320_;
 wire _09321_;
 wire _09322_;
 wire _09323_;
 wire _09324_;
 wire _09325_;
 wire _09326_;
 wire _09327_;
 wire _09328_;
 wire _09329_;
 wire _09330_;
 wire _09331_;
 wire _09332_;
 wire _09333_;
 wire _09334_;
 wire _09335_;
 wire _09336_;
 wire _09337_;
 wire _09338_;
 wire _09339_;
 wire _09340_;
 wire _09341_;
 wire _09342_;
 wire _09343_;
 wire _09344_;
 wire _09345_;
 wire _09346_;
 wire _09347_;
 wire _09348_;
 wire _09349_;
 wire _09350_;
 wire _09351_;
 wire _09352_;
 wire _09353_;
 wire _09354_;
 wire _09355_;
 wire _09356_;
 wire _09357_;
 wire _09358_;
 wire _09359_;
 wire _09360_;
 wire _09361_;
 wire _09362_;
 wire _09363_;
 wire _09364_;
 wire _09365_;
 wire _09366_;
 wire _09367_;
 wire _09368_;
 wire _09369_;
 wire _09370_;
 wire _09371_;
 wire _09372_;
 wire _09373_;
 wire _09374_;
 wire _09375_;
 wire _09376_;
 wire _09377_;
 wire _09378_;
 wire _09379_;
 wire _09380_;
 wire _09381_;
 wire _09382_;
 wire _09383_;
 wire _09384_;
 wire _09385_;
 wire _09386_;
 wire _09387_;
 wire _09388_;
 wire _09389_;
 wire _09390_;
 wire _09391_;
 wire _09392_;
 wire _09393_;
 wire _09394_;
 wire _09395_;
 wire _09396_;
 wire _09397_;
 wire _09398_;
 wire _09399_;
 wire _09400_;
 wire _09401_;
 wire _09402_;
 wire _09403_;
 wire _09404_;
 wire _09405_;
 wire _09406_;
 wire _09407_;
 wire _09408_;
 wire _09409_;
 wire _09410_;
 wire _09411_;
 wire _09412_;
 wire _09413_;
 wire _09414_;
 wire _09415_;
 wire _09416_;
 wire _09417_;
 wire _09418_;
 wire _09419_;
 wire _09420_;
 wire _09421_;
 wire _09422_;
 wire _09423_;
 wire _09424_;
 wire _09425_;
 wire _09426_;
 wire _09427_;
 wire _09428_;
 wire _09429_;
 wire _09430_;
 wire _09431_;
 wire _09432_;
 wire _09433_;
 wire _09434_;
 wire _09435_;
 wire _09436_;
 wire _09437_;
 wire _09438_;
 wire _09439_;
 wire _09440_;
 wire _09441_;
 wire _09442_;
 wire _09443_;
 wire _09444_;
 wire _09445_;
 wire _09446_;
 wire _09447_;
 wire _09448_;
 wire _09449_;
 wire _09450_;
 wire _09451_;
 wire _09452_;
 wire _09453_;
 wire _09454_;
 wire _09455_;
 wire _09456_;
 wire _09457_;
 wire _09458_;
 wire _09459_;
 wire _09460_;
 wire _09461_;
 wire _09462_;
 wire _09463_;
 wire _09464_;
 wire _09465_;
 wire _09466_;
 wire _09467_;
 wire _09468_;
 wire _09469_;
 wire _09470_;
 wire _09471_;
 wire _09472_;
 wire _09473_;
 wire _09474_;
 wire _09475_;
 wire _09476_;
 wire _09477_;
 wire _09478_;
 wire _09479_;
 wire _09480_;
 wire _09481_;
 wire _09482_;
 wire _09483_;
 wire _09484_;
 wire _09485_;
 wire _09486_;
 wire _09487_;
 wire _09488_;
 wire _09489_;
 wire _09490_;
 wire _09491_;
 wire _09492_;
 wire _09493_;
 wire _09494_;
 wire _09495_;
 wire _09496_;
 wire _09497_;
 wire _09498_;
 wire _09499_;
 wire _09500_;
 wire _09501_;
 wire _09502_;
 wire _09503_;
 wire _09504_;
 wire _09505_;
 wire _09506_;
 wire _09507_;
 wire _09508_;
 wire _09509_;
 wire _09510_;
 wire _09511_;
 wire _09512_;
 wire _09513_;
 wire _09514_;
 wire _09515_;
 wire _09516_;
 wire _09517_;
 wire _09518_;
 wire _09519_;
 wire _09520_;
 wire _09521_;
 wire _09522_;
 wire _09523_;
 wire _09524_;
 wire _09525_;
 wire _09526_;
 wire _09527_;
 wire _09528_;
 wire _09529_;
 wire _09530_;
 wire _09531_;
 wire _09532_;
 wire _09533_;
 wire _09534_;
 wire _09535_;
 wire _09536_;
 wire _09537_;
 wire _09538_;
 wire _09539_;
 wire _09540_;
 wire _09541_;
 wire _09542_;
 wire _09543_;
 wire _09544_;
 wire _09545_;
 wire _09546_;
 wire _09547_;
 wire _09548_;
 wire _09549_;
 wire _09550_;
 wire _09551_;
 wire _09552_;
 wire _09553_;
 wire _09554_;
 wire _09555_;
 wire _09556_;
 wire _09557_;
 wire _09558_;
 wire _09559_;
 wire _09560_;
 wire _09561_;
 wire _09562_;
 wire _09563_;
 wire _09564_;
 wire _09565_;
 wire _09566_;
 wire _09567_;
 wire _09568_;
 wire _09569_;
 wire _09570_;
 wire _09571_;
 wire _09572_;
 wire _09573_;
 wire _09574_;
 wire _09575_;
 wire _09576_;
 wire _09577_;
 wire _09578_;
 wire _09579_;
 wire _09580_;
 wire _09581_;
 wire _09582_;
 wire _09583_;
 wire _09584_;
 wire _09585_;
 wire _09586_;
 wire _09587_;
 wire _09588_;
 wire _09589_;
 wire _09590_;
 wire _09591_;
 wire _09592_;
 wire _09593_;
 wire _09594_;
 wire _09595_;
 wire _09596_;
 wire _09597_;
 wire _09598_;
 wire _09599_;
 wire _09600_;
 wire _09601_;
 wire _09602_;
 wire _09603_;
 wire _09604_;
 wire _09605_;
 wire _09606_;
 wire _09607_;
 wire _09608_;
 wire _09609_;
 wire _09610_;
 wire _09611_;
 wire _09612_;
 wire _09613_;
 wire _09614_;
 wire _09615_;
 wire _09616_;
 wire _09617_;
 wire _09618_;
 wire _09619_;
 wire _09620_;
 wire _09621_;
 wire _09622_;
 wire _09623_;
 wire _09624_;
 wire _09625_;
 wire _09626_;
 wire _09627_;
 wire _09628_;
 wire _09629_;
 wire _09630_;
 wire _09631_;
 wire _09632_;
 wire _09633_;
 wire _09634_;
 wire _09635_;
 wire _09636_;
 wire _09637_;
 wire _09638_;
 wire _09639_;
 wire _09640_;
 wire _09641_;
 wire _09642_;
 wire _09643_;
 wire _09644_;
 wire _09645_;
 wire _09646_;
 wire _09647_;
 wire _09648_;
 wire _09649_;
 wire _09650_;
 wire _09651_;
 wire _09652_;
 wire _09653_;
 wire _09654_;
 wire _09655_;
 wire _09656_;
 wire _09657_;
 wire _09658_;
 wire _09659_;
 wire _09660_;
 wire _09661_;
 wire _09662_;
 wire _09663_;
 wire _09664_;
 wire _09665_;
 wire _09666_;
 wire _09667_;
 wire _09668_;
 wire _09669_;
 wire _09670_;
 wire _09671_;
 wire _09672_;
 wire _09673_;
 wire _09674_;
 wire _09675_;
 wire _09676_;
 wire _09677_;
 wire _09678_;
 wire _09679_;
 wire _09680_;
 wire _09681_;
 wire _09682_;
 wire _09683_;
 wire _09684_;
 wire _09685_;
 wire _09686_;
 wire _09687_;
 wire _09688_;
 wire _09689_;
 wire _09690_;
 wire _09691_;
 wire _09692_;
 wire _09693_;
 wire _09694_;
 wire _09695_;
 wire _09696_;
 wire _09697_;
 wire _09698_;
 wire _09699_;
 wire _09700_;
 wire _09701_;
 wire _09702_;
 wire _09703_;
 wire _09704_;
 wire _09705_;
 wire _09706_;
 wire _09707_;
 wire _09708_;
 wire _09709_;
 wire _09710_;
 wire _09711_;
 wire _09712_;
 wire _09713_;
 wire _09714_;
 wire _09715_;
 wire _09716_;
 wire _09717_;
 wire _09718_;
 wire _09719_;
 wire _09720_;
 wire _09721_;
 wire _09722_;
 wire _09723_;
 wire _09724_;
 wire _09725_;
 wire _09726_;
 wire _09727_;
 wire _09728_;
 wire _09729_;
 wire _09730_;
 wire _09731_;
 wire _09732_;
 wire _09733_;
 wire _09734_;
 wire _09735_;
 wire _09736_;
 wire _09737_;
 wire _09738_;
 wire _09739_;
 wire _09740_;
 wire _09741_;
 wire _09742_;
 wire _09743_;
 wire _09744_;
 wire _09745_;
 wire _09746_;
 wire _09747_;
 wire _09748_;
 wire _09749_;
 wire _09750_;
 wire _09751_;
 wire _09752_;
 wire _09753_;
 wire _09754_;
 wire _09755_;
 wire _09756_;
 wire _09757_;
 wire _09758_;
 wire _09759_;
 wire _09760_;
 wire _09761_;
 wire _09762_;
 wire _09763_;
 wire _09764_;
 wire _09765_;
 wire _09766_;
 wire _09767_;
 wire _09768_;
 wire _09769_;
 wire _09770_;
 wire _09771_;
 wire _09772_;
 wire _09773_;
 wire _09774_;
 wire _09775_;
 wire _09776_;
 wire _09777_;
 wire _09778_;
 wire _09779_;
 wire _09780_;
 wire _09781_;
 wire _09782_;
 wire _09783_;
 wire _09784_;
 wire _09785_;
 wire _09786_;
 wire _09787_;
 wire _09788_;
 wire _09789_;
 wire _09790_;
 wire _09791_;
 wire _09792_;
 wire _09793_;
 wire _09794_;
 wire _09795_;
 wire _09796_;
 wire _09797_;
 wire _09798_;
 wire _09799_;
 wire _09800_;
 wire _09801_;
 wire _09802_;
 wire _09803_;
 wire _09804_;
 wire _09805_;
 wire _09806_;
 wire _09807_;
 wire _09808_;
 wire _09809_;
 wire _09810_;
 wire _09811_;
 wire _09812_;
 wire _09813_;
 wire _09814_;
 wire _09815_;
 wire _09816_;
 wire _09817_;
 wire _09818_;
 wire _09819_;
 wire _09820_;
 wire _09821_;
 wire _09822_;
 wire _09823_;
 wire _09824_;
 wire _09825_;
 wire _09826_;
 wire _09827_;
 wire _09828_;
 wire _09829_;
 wire _09830_;
 wire _09831_;
 wire _09832_;
 wire _09833_;
 wire _09834_;
 wire _09835_;
 wire _09836_;
 wire _09837_;
 wire _09838_;
 wire _09839_;
 wire _09840_;
 wire _09841_;
 wire _09842_;
 wire _09843_;
 wire _09844_;
 wire _09845_;
 wire _09846_;
 wire _09847_;
 wire _09848_;
 wire _09849_;
 wire _09850_;
 wire _09851_;
 wire _09852_;
 wire _09853_;
 wire _09854_;
 wire _09855_;
 wire _09856_;
 wire _09857_;
 wire _09858_;
 wire _09859_;
 wire _09860_;
 wire _09861_;
 wire _09862_;
 wire _09863_;
 wire _09864_;
 wire _09865_;
 wire _09866_;
 wire _09867_;
 wire _09868_;
 wire _09869_;
 wire _09870_;
 wire _09871_;
 wire _09872_;
 wire _09873_;
 wire _09874_;
 wire _09875_;
 wire _09876_;
 wire _09877_;
 wire _09878_;
 wire _09879_;
 wire _09880_;
 wire _09881_;
 wire _09882_;
 wire _09883_;
 wire _09884_;
 wire _09885_;
 wire _09886_;
 wire _09887_;
 wire _09888_;
 wire _09889_;
 wire _09890_;
 wire _09891_;
 wire _09892_;
 wire _09893_;
 wire _09894_;
 wire _09895_;
 wire _09896_;
 wire _09897_;
 wire _09898_;
 wire _09899_;
 wire _09900_;
 wire _09901_;
 wire _09902_;
 wire _09903_;
 wire _09904_;
 wire _09905_;
 wire _09906_;
 wire _09907_;
 wire _09908_;
 wire _09909_;
 wire _09910_;
 wire _09911_;
 wire _09912_;
 wire _09913_;
 wire _09914_;
 wire _09915_;
 wire _09916_;
 wire _09917_;
 wire _09918_;
 wire _09919_;
 wire _09920_;
 wire _09921_;
 wire _09922_;
 wire _09923_;
 wire _09924_;
 wire _09925_;
 wire _09926_;
 wire _09927_;
 wire _09928_;
 wire _09929_;
 wire _09930_;
 wire _09931_;
 wire _09932_;
 wire _09933_;
 wire _09934_;
 wire _09935_;
 wire _09936_;
 wire _09937_;
 wire _09938_;
 wire _09939_;
 wire _09940_;
 wire _09941_;
 wire _09942_;
 wire _09943_;
 wire _09944_;
 wire _09945_;
 wire _09946_;
 wire _09947_;
 wire _09948_;
 wire _09949_;
 wire _09950_;
 wire _09951_;
 wire _09952_;
 wire _09953_;
 wire _09954_;
 wire _09955_;
 wire _09956_;
 wire _09957_;
 wire _09958_;
 wire _09959_;
 wire _09960_;
 wire _09961_;
 wire _09962_;
 wire _09963_;
 wire _09964_;
 wire _09965_;
 wire _09966_;
 wire _09967_;
 wire _09968_;
 wire _09969_;
 wire _09970_;
 wire _09971_;
 wire _09972_;
 wire _09973_;
 wire _09974_;
 wire _09975_;
 wire _09976_;
 wire _09977_;
 wire _09978_;
 wire _09979_;
 wire _09980_;
 wire _09981_;
 wire _09982_;
 wire _09983_;
 wire _09984_;
 wire _09985_;
 wire _09986_;
 wire _09987_;
 wire _09988_;
 wire _09989_;
 wire _09990_;
 wire _09991_;
 wire _09992_;
 wire _09993_;
 wire _09994_;
 wire _09995_;
 wire _09996_;
 wire _09997_;
 wire _09998_;
 wire _09999_;
 wire _10000_;
 wire _10001_;
 wire _10002_;
 wire _10003_;
 wire _10004_;
 wire _10005_;
 wire _10006_;
 wire _10007_;
 wire _10008_;
 wire _10009_;
 wire _10010_;
 wire _10011_;
 wire _10012_;
 wire _10013_;
 wire _10014_;
 wire _10015_;
 wire _10016_;
 wire _10017_;
 wire _10018_;
 wire _10019_;
 wire _10020_;
 wire _10021_;
 wire _10022_;
 wire _10023_;
 wire _10024_;
 wire _10025_;
 wire _10026_;
 wire _10027_;
 wire _10028_;
 wire _10029_;
 wire _10030_;
 wire _10031_;
 wire _10032_;
 wire _10033_;
 wire _10034_;
 wire _10035_;
 wire _10036_;
 wire _10037_;
 wire _10038_;
 wire _10039_;
 wire _10040_;
 wire _10041_;
 wire _10042_;
 wire _10043_;
 wire _10044_;
 wire _10045_;
 wire _10046_;
 wire _10047_;
 wire _10048_;
 wire _10049_;
 wire _10050_;
 wire _10051_;
 wire _10052_;
 wire _10053_;
 wire _10054_;
 wire _10055_;
 wire _10056_;
 wire _10057_;
 wire _10058_;
 wire _10059_;
 wire _10060_;
 wire _10061_;
 wire _10062_;
 wire _10063_;
 wire _10064_;
 wire _10065_;
 wire _10066_;
 wire _10067_;
 wire _10068_;
 wire _10069_;
 wire _10070_;
 wire _10071_;
 wire _10072_;
 wire _10073_;
 wire _10074_;
 wire _10075_;
 wire _10076_;
 wire _10077_;
 wire _10078_;
 wire _10079_;
 wire _10080_;
 wire _10081_;
 wire _10082_;
 wire _10083_;
 wire _10084_;
 wire _10085_;
 wire _10086_;
 wire _10087_;
 wire _10088_;
 wire _10089_;
 wire _10090_;
 wire _10091_;
 wire _10092_;
 wire _10093_;
 wire _10094_;
 wire _10095_;
 wire _10096_;
 wire _10097_;
 wire _10098_;
 wire _10099_;
 wire _10100_;
 wire _10101_;
 wire _10102_;
 wire _10103_;
 wire _10104_;
 wire _10105_;
 wire _10106_;
 wire _10107_;
 wire _10108_;
 wire _10109_;
 wire _10110_;
 wire _10111_;
 wire _10112_;
 wire _10113_;
 wire _10114_;
 wire _10115_;
 wire _10116_;
 wire _10117_;
 wire _10118_;
 wire _10119_;
 wire _10120_;
 wire _10121_;
 wire _10122_;
 wire _10123_;
 wire _10124_;
 wire _10125_;
 wire _10126_;
 wire _10127_;
 wire _10128_;
 wire _10129_;
 wire _10130_;
 wire _10131_;
 wire _10132_;
 wire _10133_;
 wire _10134_;
 wire _10135_;
 wire _10136_;
 wire _10137_;
 wire _10138_;
 wire _10139_;
 wire _10140_;
 wire _10141_;
 wire _10142_;
 wire _10143_;
 wire _10144_;
 wire _10145_;
 wire _10146_;
 wire _10147_;
 wire _10148_;
 wire _10149_;
 wire _10150_;
 wire _10151_;
 wire _10152_;
 wire _10153_;
 wire _10154_;
 wire _10155_;
 wire _10156_;
 wire _10157_;
 wire _10158_;
 wire _10159_;
 wire _10160_;
 wire _10161_;
 wire _10162_;
 wire _10163_;
 wire _10164_;
 wire _10165_;
 wire _10166_;
 wire _10167_;
 wire _10168_;
 wire _10169_;
 wire _10170_;
 wire _10171_;
 wire _10172_;
 wire _10173_;
 wire _10174_;
 wire _10175_;
 wire _10176_;
 wire _10177_;
 wire _10178_;
 wire _10179_;
 wire _10180_;
 wire _10181_;
 wire _10182_;
 wire _10183_;
 wire _10184_;
 wire _10185_;
 wire _10186_;
 wire _10187_;
 wire _10188_;
 wire _10189_;
 wire _10190_;
 wire _10191_;
 wire _10192_;
 wire _10193_;
 wire _10194_;
 wire _10195_;
 wire _10196_;
 wire _10197_;
 wire _10198_;
 wire _10199_;
 wire _10200_;
 wire _10201_;
 wire _10202_;
 wire _10203_;
 wire _10204_;
 wire _10205_;
 wire _10206_;
 wire _10207_;
 wire _10208_;
 wire _10209_;
 wire _10210_;
 wire _10211_;
 wire _10212_;
 wire _10213_;
 wire _10214_;
 wire _10215_;
 wire _10216_;
 wire _10217_;
 wire _10218_;
 wire _10219_;
 wire _10220_;
 wire _10221_;
 wire _10222_;
 wire _10223_;
 wire _10224_;
 wire _10225_;
 wire _10226_;
 wire _10227_;
 wire _10228_;
 wire _10229_;
 wire _10230_;
 wire _10231_;
 wire _10232_;
 wire _10233_;
 wire _10234_;
 wire _10235_;
 wire _10236_;
 wire _10237_;
 wire _10238_;
 wire _10239_;
 wire _10240_;
 wire _10241_;
 wire _10242_;
 wire _10243_;
 wire _10244_;
 wire _10245_;
 wire _10246_;
 wire _10247_;
 wire _10248_;
 wire _10249_;
 wire _10250_;
 wire _10251_;
 wire _10252_;
 wire _10253_;
 wire _10254_;
 wire _10255_;
 wire _10256_;
 wire _10257_;
 wire _10258_;
 wire _10259_;
 wire _10260_;
 wire _10261_;
 wire _10262_;
 wire _10263_;
 wire _10264_;
 wire _10265_;
 wire _10266_;
 wire _10267_;
 wire _10268_;
 wire _10269_;
 wire _10270_;
 wire _10271_;
 wire _10272_;
 wire _10273_;
 wire _10274_;
 wire _10275_;
 wire _10276_;
 wire _10277_;
 wire _10278_;
 wire _10279_;
 wire _10280_;
 wire _10281_;
 wire _10282_;
 wire _10283_;
 wire _10284_;
 wire _10285_;
 wire _10286_;
 wire _10287_;
 wire _10288_;
 wire _10289_;
 wire _10290_;
 wire _10291_;
 wire _10292_;
 wire _10293_;
 wire _10294_;
 wire _10295_;
 wire _10296_;
 wire _10297_;
 wire _10298_;
 wire _10299_;
 wire _10300_;
 wire _10301_;
 wire _10302_;
 wire _10303_;
 wire _10304_;
 wire _10305_;
 wire _10306_;
 wire _10307_;
 wire _10308_;
 wire _10309_;
 wire _10310_;
 wire _10311_;
 wire _10312_;
 wire _10313_;
 wire _10314_;
 wire _10315_;
 wire _10316_;
 wire _10317_;
 wire _10318_;
 wire _10319_;
 wire _10320_;
 wire _10321_;
 wire _10322_;
 wire _10323_;
 wire _10324_;
 wire _10325_;
 wire _10326_;
 wire _10327_;
 wire _10328_;
 wire _10329_;
 wire _10330_;
 wire _10331_;
 wire _10332_;
 wire _10333_;
 wire _10334_;
 wire _10335_;
 wire _10336_;
 wire _10337_;
 wire _10338_;
 wire _10339_;
 wire _10340_;
 wire _10341_;
 wire _10342_;
 wire _10343_;
 wire _10344_;
 wire _10345_;
 wire _10346_;
 wire _10347_;
 wire _10348_;
 wire _10349_;
 wire _10350_;
 wire _10351_;
 wire _10352_;
 wire _10353_;
 wire _10354_;
 wire _10355_;
 wire _10356_;
 wire _10357_;
 wire _10358_;
 wire _10359_;
 wire _10360_;
 wire _10361_;
 wire _10362_;
 wire _10363_;
 wire _10364_;
 wire _10365_;
 wire _10366_;
 wire _10367_;
 wire _10368_;
 wire _10369_;
 wire _10370_;
 wire _10371_;
 wire _10372_;
 wire _10373_;
 wire _10374_;
 wire _10375_;
 wire _10376_;
 wire _10377_;
 wire _10378_;
 wire _10379_;
 wire _10380_;
 wire _10381_;
 wire _10382_;
 wire _10383_;
 wire _10384_;
 wire _10385_;
 wire _10386_;
 wire _10387_;
 wire _10388_;
 wire _10389_;
 wire _10390_;
 wire _10391_;
 wire _10392_;
 wire _10393_;
 wire _10394_;
 wire _10395_;
 wire _10396_;
 wire _10397_;
 wire _10398_;
 wire _10399_;
 wire _10400_;
 wire _10401_;
 wire _10402_;
 wire _10403_;
 wire _10404_;
 wire _10405_;
 wire _10406_;
 wire _10407_;
 wire _10408_;
 wire _10409_;
 wire _10410_;
 wire _10411_;
 wire _10412_;
 wire _10413_;
 wire _10414_;
 wire _10415_;
 wire _10416_;
 wire _10417_;
 wire _10418_;
 wire _10419_;
 wire _10420_;
 wire _10421_;
 wire _10422_;
 wire _10423_;
 wire _10424_;
 wire _10425_;
 wire _10426_;
 wire _10427_;
 wire _10428_;
 wire _10429_;
 wire _10430_;
 wire _10431_;
 wire _10432_;
 wire _10433_;
 wire _10434_;
 wire _10435_;
 wire _10436_;
 wire _10437_;
 wire _10438_;
 wire _10439_;
 wire _10440_;
 wire _10441_;
 wire _10442_;
 wire _10443_;
 wire _10444_;
 wire _10445_;
 wire _10446_;
 wire _10447_;
 wire _10448_;
 wire _10449_;
 wire _10450_;
 wire _10451_;
 wire _10452_;
 wire _10453_;
 wire _10454_;
 wire _10455_;
 wire _10456_;
 wire _10457_;
 wire _10458_;
 wire _10459_;
 wire _10460_;
 wire _10461_;
 wire _10462_;
 wire _10463_;
 wire _10464_;
 wire _10465_;
 wire _10466_;
 wire _10467_;
 wire _10468_;
 wire _10469_;
 wire _10470_;
 wire _10471_;
 wire _10472_;
 wire _10473_;
 wire _10474_;
 wire _10475_;
 wire _10476_;
 wire _10477_;
 wire _10478_;
 wire _10479_;
 wire _10480_;
 wire _10481_;
 wire _10482_;
 wire _10483_;
 wire _10484_;
 wire _10485_;
 wire _10486_;
 wire _10487_;
 wire _10488_;
 wire _10489_;
 wire _10490_;
 wire _10491_;
 wire _10492_;
 wire _10493_;
 wire _10494_;
 wire _10495_;
 wire _10496_;
 wire _10497_;
 wire _10498_;
 wire _10499_;
 wire _10500_;
 wire _10501_;
 wire _10502_;
 wire _10503_;
 wire _10504_;
 wire _10505_;
 wire _10506_;
 wire _10507_;
 wire _10508_;
 wire _10509_;
 wire _10510_;
 wire _10511_;
 wire _10512_;
 wire _10513_;
 wire _10514_;
 wire _10515_;
 wire _10516_;
 wire _10517_;
 wire _10518_;
 wire _10519_;
 wire _10520_;
 wire _10521_;
 wire _10522_;
 wire _10523_;
 wire _10524_;
 wire _10525_;
 wire _10526_;
 wire _10527_;
 wire _10528_;
 wire _10529_;
 wire _10530_;
 wire _10531_;
 wire _10532_;
 wire _10533_;
 wire _10534_;
 wire _10535_;
 wire _10536_;
 wire _10537_;
 wire _10538_;
 wire _10539_;
 wire _10540_;
 wire _10541_;
 wire _10542_;
 wire _10543_;
 wire _10544_;
 wire _10545_;
 wire _10546_;
 wire _10547_;
 wire _10548_;
 wire _10549_;
 wire _10550_;
 wire _10551_;
 wire _10552_;
 wire _10553_;
 wire _10554_;
 wire _10555_;
 wire _10556_;
 wire _10557_;
 wire _10558_;
 wire _10559_;
 wire _10560_;
 wire _10561_;
 wire _10562_;
 wire _10563_;
 wire _10564_;
 wire _10565_;
 wire _10566_;
 wire _10567_;
 wire _10568_;
 wire _10569_;
 wire _10570_;
 wire _10571_;
 wire _10572_;
 wire _10573_;
 wire _10574_;
 wire _10575_;
 wire _10576_;
 wire _10577_;
 wire _10578_;
 wire _10579_;
 wire _10580_;
 wire _10581_;
 wire _10582_;
 wire _10583_;
 wire _10584_;
 wire _10585_;
 wire _10586_;
 wire _10587_;
 wire _10588_;
 wire _10589_;
 wire _10590_;
 wire _10591_;
 wire _10592_;
 wire _10593_;
 wire _10594_;
 wire _10595_;
 wire _10596_;
 wire _10597_;
 wire _10598_;
 wire _10599_;
 wire _10600_;
 wire _10601_;
 wire _10602_;
 wire _10603_;
 wire _10604_;
 wire _10605_;
 wire _10606_;
 wire _10607_;
 wire _10608_;
 wire _10609_;
 wire _10610_;
 wire _10611_;
 wire _10612_;
 wire _10613_;
 wire _10614_;
 wire _10615_;
 wire _10616_;
 wire _10617_;
 wire _10618_;
 wire _10619_;
 wire _10620_;
 wire _10621_;
 wire _10622_;
 wire _10623_;
 wire _10624_;
 wire _10625_;
 wire _10626_;
 wire _10627_;
 wire _10628_;
 wire _10629_;
 wire _10630_;
 wire _10631_;
 wire _10632_;
 wire _10633_;
 wire _10634_;
 wire _10635_;
 wire _10636_;
 wire _10637_;
 wire _10638_;
 wire _10639_;
 wire _10640_;
 wire _10641_;
 wire _10642_;
 wire _10643_;
 wire _10644_;
 wire _10645_;
 wire _10646_;
 wire _10647_;
 wire _10648_;
 wire _10649_;
 wire _10650_;
 wire _10651_;
 wire _10652_;
 wire _10653_;
 wire _10654_;
 wire _10655_;
 wire _10656_;
 wire _10657_;
 wire _10658_;
 wire _10659_;
 wire _10660_;
 wire _10661_;
 wire _10662_;
 wire _10663_;
 wire _10664_;
 wire _10665_;
 wire _10666_;
 wire _10667_;
 wire _10668_;
 wire _10669_;
 wire _10670_;
 wire _10671_;
 wire _10672_;
 wire _10673_;
 wire _10674_;
 wire _10675_;
 wire _10676_;
 wire _10677_;
 wire _10678_;
 wire _10679_;
 wire _10680_;
 wire _10681_;
 wire _10682_;
 wire _10683_;
 wire _10684_;
 wire _10685_;
 wire _10686_;
 wire _10687_;
 wire _10688_;
 wire _10689_;
 wire _10690_;
 wire _10691_;
 wire _10692_;
 wire _10693_;
 wire _10694_;
 wire _10695_;
 wire _10696_;
 wire _10697_;
 wire _10698_;
 wire _10699_;
 wire _10700_;
 wire _10701_;
 wire _10702_;
 wire _10703_;
 wire _10704_;
 wire _10705_;
 wire _10706_;
 wire _10707_;
 wire _10708_;
 wire _10709_;
 wire _10710_;
 wire _10711_;
 wire _10712_;
 wire _10713_;
 wire _10714_;
 wire _10715_;
 wire _10716_;
 wire _10717_;
 wire _10718_;
 wire _10719_;
 wire _10720_;
 wire _10721_;
 wire _10722_;
 wire _10723_;
 wire _10724_;
 wire _10725_;
 wire _10726_;
 wire _10727_;
 wire _10728_;
 wire _10729_;
 wire _10730_;
 wire _10731_;
 wire _10732_;
 wire _10733_;
 wire _10734_;
 wire _10735_;
 wire _10736_;
 wire _10737_;
 wire _10738_;
 wire _10739_;
 wire _10740_;
 wire _10741_;
 wire _10742_;
 wire _10743_;
 wire _10744_;
 wire _10745_;
 wire _10746_;
 wire _10747_;
 wire _10748_;
 wire _10749_;
 wire _10750_;
 wire _10751_;
 wire _10752_;
 wire _10753_;
 wire _10754_;
 wire _10755_;
 wire _10756_;
 wire _10757_;
 wire _10758_;
 wire _10759_;
 wire _10760_;
 wire _10761_;
 wire _10762_;
 wire _10763_;
 wire _10764_;
 wire _10765_;
 wire _10766_;
 wire _10767_;
 wire _10768_;
 wire _10769_;
 wire _10770_;
 wire _10771_;
 wire _10772_;
 wire _10773_;
 wire _10774_;
 wire _10775_;
 wire _10776_;
 wire _10777_;
 wire _10778_;
 wire _10779_;
 wire _10780_;
 wire _10781_;
 wire _10782_;
 wire _10783_;
 wire _10784_;
 wire _10785_;
 wire _10786_;
 wire _10787_;
 wire _10788_;
 wire _10789_;
 wire _10790_;
 wire _10791_;
 wire _10792_;
 wire _10793_;
 wire _10794_;
 wire _10795_;
 wire _10796_;
 wire _10797_;
 wire _10798_;
 wire _10799_;
 wire _10800_;
 wire _10801_;
 wire _10802_;
 wire _10803_;
 wire _10804_;
 wire _10805_;
 wire _10806_;
 wire _10807_;
 wire _10808_;
 wire _10809_;
 wire _10810_;
 wire _10811_;
 wire _10812_;
 wire _10813_;
 wire _10814_;
 wire _10815_;
 wire _10816_;
 wire _10817_;
 wire _10818_;
 wire _10819_;
 wire _10820_;
 wire _10821_;
 wire _10822_;
 wire _10823_;
 wire _10824_;
 wire _10825_;
 wire _10826_;
 wire _10827_;
 wire _10828_;
 wire _10829_;
 wire _10830_;
 wire _10831_;
 wire _10832_;
 wire _10833_;
 wire _10834_;
 wire _10835_;
 wire _10836_;
 wire _10837_;
 wire _10838_;
 wire _10839_;
 wire _10840_;
 wire _10841_;
 wire _10842_;
 wire _10843_;
 wire _10844_;
 wire _10845_;
 wire _10846_;
 wire _10847_;
 wire _10848_;
 wire _10849_;
 wire _10850_;
 wire _10851_;
 wire _10852_;
 wire _10853_;
 wire _10854_;
 wire _10855_;
 wire _10856_;
 wire _10857_;
 wire _10858_;
 wire _10859_;
 wire _10860_;
 wire _10861_;
 wire _10862_;
 wire _10863_;
 wire _10864_;
 wire _10865_;
 wire _10866_;
 wire _10867_;
 wire _10868_;
 wire _10869_;
 wire _10870_;
 wire _10871_;
 wire _10872_;
 wire _10873_;
 wire _10874_;
 wire _10875_;
 wire _10876_;
 wire _10877_;
 wire _10878_;
 wire _10879_;
 wire _10880_;
 wire _10881_;
 wire _10882_;
 wire _10883_;
 wire _10884_;
 wire _10885_;
 wire _10886_;
 wire _10887_;
 wire _10888_;
 wire _10889_;
 wire _10890_;
 wire _10891_;
 wire _10892_;
 wire _10893_;
 wire _10894_;
 wire _10895_;
 wire _10896_;
 wire _10897_;
 wire _10898_;
 wire _10899_;
 wire _10900_;
 wire _10901_;
 wire _10902_;
 wire _10903_;
 wire _10904_;
 wire _10905_;
 wire _10906_;
 wire _10907_;
 wire _10908_;
 wire _10909_;
 wire _10910_;
 wire _10911_;
 wire _10912_;
 wire _10913_;
 wire _10914_;
 wire _10915_;
 wire _10916_;
 wire _10917_;
 wire _10918_;
 wire _10919_;
 wire _10920_;
 wire _10921_;
 wire _10922_;
 wire _10923_;
 wire _10924_;
 wire _10925_;
 wire _10926_;
 wire _10927_;
 wire _10928_;
 wire _10929_;
 wire _10930_;
 wire _10931_;
 wire _10932_;
 wire _10933_;
 wire _10934_;
 wire _10935_;
 wire _10936_;
 wire _10937_;
 wire _10938_;
 wire _10939_;
 wire _10940_;
 wire _10941_;
 wire _10942_;
 wire _10943_;
 wire _10944_;
 wire _10945_;
 wire _10946_;
 wire _10947_;
 wire _10948_;
 wire _10949_;
 wire _10950_;
 wire _10951_;
 wire _10952_;
 wire _10953_;
 wire _10954_;
 wire _10955_;
 wire _10956_;
 wire _10957_;
 wire _10958_;
 wire _10959_;
 wire _10960_;
 wire _10961_;
 wire _10962_;
 wire _10963_;
 wire _10964_;
 wire _10965_;
 wire _10966_;
 wire _10967_;
 wire _10968_;
 wire _10969_;
 wire _10970_;
 wire _10971_;
 wire _10972_;
 wire _10973_;
 wire _10974_;
 wire _10975_;
 wire _10976_;
 wire _10977_;
 wire _10978_;
 wire _10979_;
 wire _10980_;
 wire _10981_;
 wire _10982_;
 wire _10983_;
 wire _10984_;
 wire _10985_;
 wire _10986_;
 wire _10987_;
 wire _10988_;
 wire _10989_;
 wire _10990_;
 wire _10991_;
 wire _10992_;
 wire _10993_;
 wire _10994_;
 wire _10995_;
 wire _10996_;
 wire _10997_;
 wire _10998_;
 wire _10999_;
 wire _11000_;
 wire _11001_;
 wire _11002_;
 wire _11003_;
 wire _11004_;
 wire _11005_;
 wire _11006_;
 wire _11007_;
 wire _11008_;
 wire _11009_;
 wire _11010_;
 wire _11011_;
 wire _11012_;
 wire _11013_;
 wire _11014_;
 wire _11015_;
 wire _11016_;
 wire _11017_;
 wire _11018_;
 wire _11019_;
 wire _11020_;
 wire _11021_;
 wire _11022_;
 wire _11023_;
 wire _11024_;
 wire _11025_;
 wire _11026_;
 wire _11027_;
 wire _11028_;
 wire _11029_;
 wire _11030_;
 wire _11031_;
 wire _11032_;
 wire _11033_;
 wire _11034_;
 wire _11035_;
 wire _11036_;
 wire _11037_;
 wire _11038_;
 wire _11039_;
 wire _11040_;
 wire _11041_;
 wire _11042_;
 wire _11043_;
 wire _11044_;
 wire _11045_;
 wire _11046_;
 wire _11047_;
 wire _11048_;
 wire _11049_;
 wire _11050_;
 wire _11051_;
 wire _11052_;
 wire _11053_;
 wire _11054_;
 wire _11055_;
 wire _11056_;
 wire _11057_;
 wire _11058_;
 wire _11059_;
 wire _11060_;
 wire _11061_;
 wire _11062_;
 wire _11063_;
 wire _11064_;
 wire _11065_;
 wire _11066_;
 wire _11067_;
 wire _11068_;
 wire _11069_;
 wire _11070_;
 wire _11071_;
 wire _11072_;
 wire _11073_;
 wire _11074_;
 wire _11075_;
 wire _11076_;
 wire _11077_;
 wire _11078_;
 wire _11079_;
 wire _11080_;
 wire _11081_;
 wire _11082_;
 wire _11083_;
 wire _11084_;
 wire _11085_;
 wire _11086_;
 wire _11087_;
 wire _11088_;
 wire _11089_;
 wire _11090_;
 wire _11091_;
 wire _11092_;
 wire _11093_;
 wire _11094_;
 wire _11095_;
 wire _11096_;
 wire _11097_;
 wire _11098_;
 wire _11099_;
 wire _11100_;
 wire _11101_;
 wire _11102_;
 wire _11103_;
 wire _11104_;
 wire _11105_;
 wire _11106_;
 wire _11107_;
 wire _11108_;
 wire _11109_;
 wire _11110_;
 wire _11111_;
 wire _11112_;
 wire _11113_;
 wire _11114_;
 wire _11115_;
 wire _11116_;
 wire _11117_;
 wire _11118_;
 wire _11119_;
 wire _11120_;
 wire _11121_;
 wire _11122_;
 wire _11123_;
 wire _11124_;
 wire _11125_;
 wire _11126_;
 wire _11127_;
 wire _11128_;
 wire _11129_;
 wire _11130_;
 wire _11131_;
 wire _11132_;
 wire _11133_;
 wire _11134_;
 wire _11135_;
 wire _11136_;
 wire _11137_;
 wire _11138_;
 wire _11139_;
 wire _11140_;
 wire _11141_;
 wire _11142_;
 wire _11143_;
 wire _11144_;
 wire _11145_;
 wire _11146_;
 wire _11147_;
 wire _11148_;
 wire _11149_;
 wire _11150_;
 wire _11151_;
 wire _11152_;
 wire _11153_;
 wire _11154_;
 wire _11155_;
 wire _11156_;
 wire _11157_;
 wire _11158_;
 wire _11159_;
 wire _11160_;
 wire _11161_;
 wire _11162_;
 wire _11163_;
 wire _11164_;
 wire _11165_;
 wire _11166_;
 wire _11167_;
 wire _11168_;
 wire _11169_;
 wire _11170_;
 wire _11171_;
 wire _11172_;
 wire _11173_;
 wire _11174_;
 wire _11175_;
 wire _11176_;
 wire _11177_;
 wire _11178_;
 wire _11179_;
 wire _11180_;
 wire _11181_;
 wire _11182_;
 wire _11183_;
 wire _11184_;
 wire _11185_;
 wire _11186_;
 wire _11187_;
 wire _11188_;
 wire _11189_;
 wire _11190_;
 wire _11191_;
 wire _11192_;
 wire _11193_;
 wire _11194_;
 wire _11195_;
 wire _11196_;
 wire _11197_;
 wire _11198_;
 wire _11199_;
 wire _11200_;
 wire _11201_;
 wire _11202_;
 wire _11203_;
 wire _11204_;
 wire _11205_;
 wire _11206_;
 wire _11207_;
 wire _11208_;
 wire _11209_;
 wire _11210_;
 wire _11211_;
 wire _11212_;
 wire _11213_;
 wire _11214_;
 wire _11215_;
 wire _11216_;
 wire _11217_;
 wire _11218_;
 wire _11219_;
 wire _11220_;
 wire _11221_;
 wire _11222_;
 wire _11223_;
 wire _11224_;
 wire _11225_;
 wire _11226_;
 wire _11227_;
 wire _11228_;
 wire _11229_;
 wire _11230_;
 wire _11231_;
 wire _11232_;
 wire _11233_;
 wire _11234_;
 wire _11235_;
 wire _11236_;
 wire _11237_;
 wire _11238_;
 wire _11239_;
 wire _11240_;
 wire _11241_;
 wire _11242_;
 wire _11243_;
 wire _11244_;
 wire _11245_;
 wire _11246_;
 wire _11247_;
 wire _11248_;
 wire _11249_;
 wire _11250_;
 wire _11251_;
 wire _11252_;
 wire _11253_;
 wire _11254_;
 wire _11255_;
 wire _11256_;
 wire _11257_;
 wire _11258_;
 wire _11259_;
 wire _11260_;
 wire _11261_;
 wire _11262_;
 wire _11263_;
 wire _11264_;
 wire _11265_;
 wire _11266_;
 wire _11267_;
 wire _11268_;
 wire _11269_;
 wire _11270_;
 wire _11271_;
 wire _11272_;
 wire _11273_;
 wire _11274_;
 wire _11275_;
 wire _11276_;
 wire _11277_;
 wire _11278_;
 wire _11279_;
 wire _11280_;
 wire _11281_;
 wire _11282_;
 wire _11283_;
 wire _11284_;
 wire _11285_;
 wire _11286_;
 wire _11287_;
 wire _11288_;
 wire _11289_;
 wire _11290_;
 wire _11291_;
 wire _11292_;
 wire _11293_;
 wire _11294_;
 wire _11295_;
 wire _11296_;
 wire _11297_;
 wire _11298_;
 wire _11299_;
 wire _11300_;
 wire _11301_;
 wire _11302_;
 wire _11303_;
 wire _11304_;
 wire _11305_;
 wire _11306_;
 wire _11307_;
 wire _11308_;
 wire _11309_;
 wire _11310_;
 wire _11311_;
 wire _11312_;
 wire _11313_;
 wire _11314_;
 wire _11315_;
 wire _11316_;
 wire _11317_;
 wire _11318_;
 wire _11319_;
 wire _11320_;
 wire _11321_;
 wire _11322_;
 wire _11323_;
 wire _11324_;
 wire _11325_;
 wire _11326_;
 wire _11327_;
 wire _11328_;
 wire _11329_;
 wire _11330_;
 wire _11331_;
 wire _11332_;
 wire _11333_;
 wire _11334_;
 wire _11335_;
 wire _11336_;
 wire _11337_;
 wire _11338_;
 wire _11339_;
 wire _11340_;
 wire _11341_;
 wire _11342_;
 wire _11343_;
 wire _11344_;
 wire _11345_;
 wire _11346_;
 wire _11347_;
 wire _11348_;
 wire _11349_;
 wire _11350_;
 wire _11351_;
 wire _11352_;
 wire _11353_;
 wire _11354_;
 wire _11355_;
 wire _11356_;
 wire _11357_;
 wire _11358_;
 wire _11359_;
 wire _11360_;
 wire _11361_;
 wire _11362_;
 wire _11363_;
 wire _11364_;
 wire _11365_;
 wire _11366_;
 wire _11367_;
 wire _11368_;
 wire _11369_;
 wire _11370_;
 wire _11371_;
 wire _11372_;
 wire _11373_;
 wire _11374_;
 wire _11375_;
 wire _11376_;
 wire _11377_;
 wire _11378_;
 wire _11379_;
 wire _11380_;
 wire _11381_;
 wire _11382_;
 wire _11383_;
 wire _11384_;
 wire _11385_;
 wire _11386_;
 wire _11387_;
 wire _11388_;
 wire _11389_;
 wire _11390_;
 wire _11391_;
 wire _11392_;
 wire _11393_;
 wire _11394_;
 wire _11395_;
 wire _11396_;
 wire _11397_;
 wire _11398_;
 wire _11399_;
 wire _11400_;
 wire _11401_;
 wire _11402_;
 wire _11403_;
 wire _11404_;
 wire _11405_;
 wire _11406_;
 wire _11407_;
 wire _11408_;
 wire _11409_;
 wire _11410_;
 wire _11411_;
 wire _11412_;
 wire _11413_;
 wire _11414_;
 wire _11415_;
 wire _11416_;
 wire _11417_;
 wire _11418_;
 wire _11419_;
 wire _11420_;
 wire _11421_;
 wire _11422_;
 wire _11423_;
 wire _11424_;
 wire _11425_;
 wire _11426_;
 wire _11427_;
 wire _11428_;
 wire _11429_;
 wire _11430_;
 wire _11431_;
 wire _11432_;
 wire _11433_;
 wire _11434_;
 wire _11435_;
 wire _11436_;
 wire _11437_;
 wire _11438_;
 wire _11439_;
 wire _11440_;
 wire _11441_;
 wire _11442_;
 wire _11443_;
 wire _11444_;
 wire _11445_;
 wire _11446_;
 wire _11447_;
 wire _11448_;
 wire _11449_;
 wire _11450_;
 wire _11451_;
 wire _11452_;
 wire _11453_;
 wire _11454_;
 wire _11455_;
 wire _11456_;
 wire _11457_;
 wire _11458_;
 wire _11459_;
 wire _11460_;
 wire _11461_;
 wire _11462_;
 wire _11463_;
 wire _11464_;
 wire _11465_;
 wire _11466_;
 wire _11467_;
 wire _11468_;
 wire _11469_;
 wire _11470_;
 wire _11471_;
 wire _11472_;
 wire _11473_;
 wire _11474_;
 wire _11475_;
 wire _11476_;
 wire _11477_;
 wire _11478_;
 wire _11479_;
 wire _11480_;
 wire _11481_;
 wire _11482_;
 wire _11483_;
 wire _11484_;
 wire _11485_;
 wire _11486_;
 wire _11487_;
 wire _11488_;
 wire _11489_;
 wire _11490_;
 wire _11491_;
 wire _11492_;
 wire _11493_;
 wire _11494_;
 wire _11495_;
 wire _11496_;
 wire _11497_;
 wire _11498_;
 wire _11499_;
 wire _11500_;
 wire _11501_;
 wire _11502_;
 wire _11503_;
 wire _11504_;
 wire _11505_;
 wire _11506_;
 wire _11507_;
 wire _11508_;
 wire _11509_;
 wire _11510_;
 wire _11511_;
 wire _11512_;
 wire _11513_;
 wire _11514_;
 wire _11515_;
 wire _11516_;
 wire _11517_;
 wire _11518_;
 wire _11519_;
 wire _11520_;
 wire _11521_;
 wire _11522_;
 wire _11523_;
 wire _11524_;
 wire _11525_;
 wire _11526_;
 wire _11527_;
 wire _11528_;
 wire _11529_;
 wire _11530_;
 wire _11531_;
 wire _11532_;
 wire _11533_;
 wire _11534_;
 wire _11535_;
 wire _11536_;
 wire _11537_;
 wire _11538_;
 wire _11539_;
 wire _11540_;
 wire _11541_;
 wire _11542_;
 wire _11543_;
 wire _11544_;
 wire _11545_;
 wire _11546_;
 wire _11547_;
 wire _11548_;
 wire _11549_;
 wire _11550_;
 wire _11551_;
 wire _11552_;
 wire _11553_;
 wire _11554_;
 wire _11555_;
 wire _11556_;
 wire _11557_;
 wire _11558_;
 wire _11559_;
 wire _11560_;
 wire _11561_;
 wire _11562_;
 wire _11563_;
 wire _11564_;
 wire _11565_;
 wire _11566_;
 wire _11567_;
 wire _11568_;
 wire _11569_;
 wire _11570_;
 wire _11571_;
 wire _11572_;
 wire _11573_;
 wire _11574_;
 wire _11575_;
 wire _11576_;
 wire _11577_;
 wire _11578_;
 wire _11579_;
 wire _11580_;
 wire _11581_;
 wire _11582_;
 wire _11583_;
 wire _11584_;
 wire _11585_;
 wire _11586_;
 wire _11587_;
 wire _11588_;
 wire _11589_;
 wire _11590_;
 wire _11591_;
 wire _11592_;
 wire _11593_;
 wire _11594_;
 wire _11595_;
 wire _11596_;
 wire _11597_;
 wire _11598_;
 wire _11599_;
 wire _11600_;
 wire _11601_;
 wire _11602_;
 wire _11603_;
 wire _11604_;
 wire _11605_;
 wire _11606_;
 wire _11607_;
 wire _11608_;
 wire _11609_;
 wire _11610_;
 wire _11611_;
 wire _11612_;
 wire _11613_;
 wire _11614_;
 wire _11615_;
 wire _11616_;
 wire _11617_;
 wire _11618_;
 wire _11619_;
 wire _11620_;
 wire _11621_;
 wire _11622_;
 wire _11623_;
 wire _11624_;
 wire _11625_;
 wire _11626_;
 wire _11627_;
 wire _11628_;
 wire _11629_;
 wire _11630_;
 wire _11631_;
 wire _11632_;
 wire _11633_;
 wire _11634_;
 wire _11635_;
 wire _11636_;
 wire _11637_;
 wire _11638_;
 wire _11639_;
 wire _11640_;
 wire _11641_;
 wire _11642_;
 wire _11643_;
 wire _11644_;
 wire _11645_;
 wire _11646_;
 wire _11647_;
 wire _11648_;
 wire _11649_;
 wire _11650_;
 wire _11651_;
 wire _11652_;
 wire _11653_;
 wire _11654_;
 wire _11655_;
 wire _11656_;
 wire _11657_;
 wire _11658_;
 wire _11659_;
 wire _11660_;
 wire _11661_;
 wire _11662_;
 wire _11663_;
 wire _11664_;
 wire _11665_;
 wire _11666_;
 wire _11667_;
 wire _11668_;
 wire _11669_;
 wire _11670_;
 wire _11671_;
 wire _11672_;
 wire _11673_;
 wire _11674_;
 wire _11675_;
 wire _11676_;
 wire _11677_;
 wire _11678_;
 wire _11679_;
 wire _11680_;
 wire _11681_;
 wire _11682_;
 wire _11683_;
 wire _11684_;
 wire _11685_;
 wire _11686_;
 wire _11687_;
 wire _11688_;
 wire _11689_;
 wire _11690_;
 wire _11691_;
 wire _11692_;
 wire _11693_;
 wire _11694_;
 wire _11695_;
 wire _11696_;
 wire _11697_;
 wire _11698_;
 wire _11699_;
 wire _11700_;
 wire _11701_;
 wire _11702_;
 wire _11703_;
 wire _11704_;
 wire _11705_;
 wire _11706_;
 wire _11707_;
 wire _11708_;
 wire _11709_;
 wire _11710_;
 wire _11711_;
 wire _11712_;
 wire _11713_;
 wire _11714_;
 wire _11715_;
 wire _11716_;
 wire _11717_;
 wire _11718_;
 wire _11719_;
 wire _11720_;
 wire _11721_;
 wire _11722_;
 wire _11723_;
 wire _11724_;
 wire _11725_;
 wire _11726_;
 wire _11727_;
 wire _11728_;
 wire _11729_;
 wire _11730_;
 wire _11731_;
 wire _11732_;
 wire _11733_;
 wire _11734_;
 wire _11735_;
 wire _11736_;
 wire _11737_;
 wire _11738_;
 wire _11739_;
 wire _11740_;
 wire _11741_;
 wire _11742_;
 wire _11743_;
 wire _11744_;
 wire _11745_;
 wire _11746_;
 wire _11747_;
 wire _11748_;
 wire _11749_;
 wire _11750_;
 wire _11751_;
 wire _11752_;
 wire _11753_;
 wire _11754_;
 wire _11755_;
 wire _11756_;
 wire _11757_;
 wire _11758_;
 wire _11759_;
 wire _11760_;
 wire _11761_;
 wire _11762_;
 wire _11763_;
 wire _11764_;
 wire _11765_;
 wire _11766_;
 wire _11767_;
 wire _11768_;
 wire _11769_;
 wire _11770_;
 wire _11771_;
 wire _11772_;
 wire _11773_;
 wire _11774_;
 wire _11775_;
 wire _11776_;
 wire _11777_;
 wire _11778_;
 wire _11779_;
 wire _11780_;
 wire _11781_;
 wire _11782_;
 wire _11783_;
 wire _11784_;
 wire _11785_;
 wire _11786_;
 wire _11787_;
 wire _11788_;
 wire _11789_;
 wire _11790_;
 wire _11791_;
 wire _11792_;
 wire _11793_;
 wire _11794_;
 wire _11795_;
 wire _11796_;
 wire _11797_;
 wire _11798_;
 wire _11799_;
 wire _11800_;
 wire _11801_;
 wire _11802_;
 wire _11803_;
 wire _11804_;
 wire _11805_;
 wire _11806_;
 wire _11807_;
 wire _11808_;
 wire _11809_;
 wire _11810_;
 wire _11811_;
 wire _11812_;
 wire _11813_;
 wire _11814_;
 wire _11815_;
 wire _11816_;
 wire _11817_;
 wire _11818_;
 wire _11819_;
 wire _11820_;
 wire _11821_;
 wire _11822_;
 wire _11823_;
 wire _11824_;
 wire _11825_;
 wire _11826_;
 wire _11827_;
 wire _11828_;
 wire _11829_;
 wire _11830_;
 wire _11831_;
 wire _11832_;
 wire _11833_;
 wire _11834_;
 wire _11835_;
 wire _11836_;
 wire _11837_;
 wire _11838_;
 wire _11839_;
 wire _11840_;
 wire _11841_;
 wire _11842_;
 wire _11843_;
 wire _11844_;
 wire _11845_;
 wire _11846_;
 wire _11847_;
 wire _11848_;
 wire _11849_;
 wire _11850_;
 wire _11851_;
 wire _11852_;
 wire _11853_;
 wire _11854_;
 wire _11855_;
 wire _11856_;
 wire _11857_;
 wire _11858_;
 wire _11859_;
 wire _11860_;
 wire _11861_;
 wire _11862_;
 wire _11863_;
 wire _11864_;
 wire _11865_;
 wire _11866_;
 wire _11867_;
 wire _11868_;
 wire _11869_;
 wire _11870_;
 wire _11871_;
 wire _11872_;
 wire _11873_;
 wire _11874_;
 wire _11875_;
 wire _11876_;
 wire _11877_;
 wire _11878_;
 wire _11879_;
 wire _11880_;
 wire _11881_;
 wire _11882_;
 wire _11883_;
 wire _11884_;
 wire _11885_;
 wire _11886_;
 wire _11887_;
 wire _11888_;
 wire _11889_;
 wire _11890_;
 wire _11891_;
 wire _11892_;
 wire _11893_;
 wire _11894_;
 wire _11895_;
 wire _11896_;
 wire _11897_;
 wire _11898_;
 wire _11899_;
 wire _11900_;
 wire _11901_;
 wire _11902_;
 wire _11903_;
 wire _11904_;
 wire _11905_;
 wire _11906_;
 wire _11907_;
 wire _11908_;
 wire _11909_;
 wire _11910_;
 wire _11911_;
 wire _11912_;
 wire _11913_;
 wire _11914_;
 wire _11915_;
 wire _11916_;
 wire _11917_;
 wire _11918_;
 wire _11919_;
 wire _11920_;
 wire _11921_;
 wire _11922_;
 wire _11923_;
 wire _11924_;
 wire _11925_;
 wire _11926_;
 wire _11927_;
 wire _11928_;
 wire _11929_;
 wire _11930_;
 wire _11931_;
 wire _11932_;
 wire _11933_;
 wire _11934_;
 wire _11935_;
 wire _11936_;
 wire _11937_;
 wire _11938_;
 wire _11939_;
 wire _11940_;
 wire _11941_;
 wire _11942_;
 wire _11943_;
 wire _11944_;
 wire _11945_;
 wire _11946_;
 wire _11947_;
 wire _11948_;
 wire _11949_;
 wire _11950_;
 wire _11951_;
 wire _11952_;
 wire _11953_;
 wire _11954_;
 wire _11955_;
 wire _11956_;
 wire _11957_;
 wire _11958_;
 wire _11959_;
 wire _11960_;
 wire _11961_;
 wire _11962_;
 wire _11963_;
 wire _11964_;
 wire _11965_;
 wire _11966_;
 wire _11967_;
 wire _11968_;
 wire _11969_;
 wire _11970_;
 wire _11971_;
 wire _11972_;
 wire _11973_;
 wire _11974_;
 wire _11975_;
 wire _11976_;
 wire _11977_;
 wire _11978_;
 wire _11979_;
 wire _11980_;
 wire _11981_;
 wire _11982_;
 wire _11983_;
 wire _11984_;
 wire _11985_;
 wire _11986_;
 wire _11987_;
 wire _11988_;
 wire _11989_;
 wire _11990_;
 wire _11991_;
 wire _11992_;
 wire _11993_;
 wire _11994_;
 wire _11995_;
 wire _11996_;
 wire _11997_;
 wire _11998_;
 wire _11999_;
 wire _12000_;
 wire _12001_;
 wire _12002_;
 wire _12003_;
 wire _12004_;
 wire _12005_;
 wire _12006_;
 wire _12007_;
 wire _12008_;
 wire _12009_;
 wire _12010_;
 wire _12011_;
 wire _12012_;
 wire _12013_;
 wire _12014_;
 wire _12015_;
 wire _12016_;
 wire _12017_;
 wire _12018_;
 wire _12019_;
 wire _12020_;
 wire _12021_;
 wire _12022_;
 wire _12023_;
 wire _12024_;
 wire _12025_;
 wire _12026_;
 wire _12027_;
 wire _12028_;
 wire _12029_;
 wire _12030_;
 wire _12031_;
 wire _12032_;
 wire _12033_;
 wire _12034_;
 wire _12035_;
 wire _12036_;
 wire _12037_;
 wire _12038_;
 wire _12039_;
 wire _12040_;
 wire _12041_;
 wire _12042_;
 wire _12043_;
 wire _12044_;
 wire _12045_;
 wire _12046_;
 wire _12047_;
 wire _12048_;
 wire _12049_;
 wire _12050_;
 wire _12051_;
 wire _12052_;
 wire _12053_;
 wire _12054_;
 wire _12055_;
 wire _12056_;
 wire _12057_;
 wire _12058_;
 wire _12059_;
 wire _12060_;
 wire _12061_;
 wire _12062_;
 wire _12063_;
 wire _12064_;
 wire _12065_;
 wire _12066_;
 wire _12067_;
 wire _12068_;
 wire _12069_;
 wire _12070_;
 wire _12071_;
 wire _12072_;
 wire _12073_;
 wire _12074_;
 wire _12075_;
 wire _12076_;
 wire _12077_;
 wire _12078_;
 wire _12079_;
 wire _12080_;
 wire _12081_;
 wire _12082_;
 wire _12083_;
 wire _12084_;
 wire _12085_;
 wire _12086_;
 wire _12087_;
 wire _12088_;
 wire _12089_;
 wire _12090_;
 wire _12091_;
 wire _12092_;
 wire _12093_;
 wire _12094_;
 wire _12095_;
 wire _12096_;
 wire _12097_;
 wire _12098_;
 wire _12099_;
 wire _12100_;
 wire _12101_;
 wire _12102_;
 wire _12103_;
 wire _12104_;
 wire _12105_;
 wire _12106_;
 wire _12107_;
 wire _12108_;
 wire _12109_;
 wire _12110_;
 wire _12111_;
 wire _12112_;
 wire _12113_;
 wire _12114_;
 wire _12115_;
 wire _12116_;
 wire _12117_;
 wire _12118_;
 wire _12119_;
 wire _12120_;
 wire _12121_;
 wire _12122_;
 wire _12123_;
 wire _12124_;
 wire _12125_;
 wire _12126_;
 wire _12127_;
 wire _12128_;
 wire _12129_;
 wire _12130_;
 wire _12131_;
 wire _12132_;
 wire _12133_;
 wire _12134_;
 wire _12135_;
 wire _12136_;
 wire _12137_;
 wire _12138_;
 wire _12139_;
 wire _12140_;
 wire _12141_;
 wire _12142_;
 wire _12143_;
 wire _12144_;
 wire _12145_;
 wire _12146_;
 wire _12147_;
 wire _12148_;
 wire _12149_;
 wire _12150_;
 wire _12151_;
 wire _12152_;
 wire _12153_;
 wire _12154_;
 wire _12155_;
 wire _12156_;
 wire _12157_;
 wire _12158_;
 wire _12159_;
 wire _12160_;
 wire _12161_;
 wire _12162_;
 wire _12163_;
 wire _12164_;
 wire _12165_;
 wire _12166_;
 wire _12167_;
 wire _12168_;
 wire _12169_;
 wire _12170_;
 wire _12171_;
 wire _12172_;
 wire _12173_;
 wire _12174_;
 wire _12175_;
 wire _12176_;
 wire _12177_;
 wire _12178_;
 wire _12179_;
 wire _12180_;
 wire _12181_;
 wire _12182_;
 wire _12183_;
 wire _12184_;
 wire _12185_;
 wire _12186_;
 wire _12187_;
 wire _12188_;
 wire _12189_;
 wire _12190_;
 wire _12191_;
 wire _12192_;
 wire _12193_;
 wire _12194_;
 wire _12195_;
 wire _12196_;
 wire _12197_;
 wire _12198_;
 wire _12199_;
 wire _12200_;
 wire _12201_;
 wire _12202_;
 wire _12203_;
 wire _12204_;
 wire _12205_;
 wire _12206_;
 wire _12207_;
 wire _12208_;
 wire _12209_;
 wire _12210_;
 wire _12211_;
 wire _12212_;
 wire _12213_;
 wire _12214_;
 wire _12215_;
 wire _12216_;
 wire _12217_;
 wire _12218_;
 wire _12219_;
 wire _12220_;
 wire _12221_;
 wire _12222_;
 wire _12223_;
 wire _12224_;
 wire _12225_;
 wire _12226_;
 wire _12227_;
 wire _12228_;
 wire _12229_;
 wire _12230_;
 wire _12231_;
 wire _12232_;
 wire _12233_;
 wire _12234_;
 wire _12235_;
 wire _12236_;
 wire _12237_;
 wire _12238_;
 wire _12239_;
 wire _12240_;
 wire _12241_;
 wire _12242_;
 wire _12243_;
 wire _12244_;
 wire _12245_;
 wire _12246_;
 wire _12247_;
 wire _12248_;
 wire _12249_;
 wire _12250_;
 wire _12251_;
 wire _12252_;
 wire _12253_;
 wire _12254_;
 wire _12255_;
 wire _12256_;
 wire _12257_;
 wire _12258_;
 wire _12259_;
 wire _12260_;
 wire _12261_;
 wire _12262_;
 wire _12263_;
 wire _12264_;
 wire _12265_;
 wire _12266_;
 wire _12267_;
 wire _12268_;
 wire _12269_;
 wire _12270_;
 wire _12271_;
 wire _12272_;
 wire _12273_;
 wire _12274_;
 wire _12275_;
 wire _12276_;
 wire _12277_;
 wire _12278_;
 wire _12279_;
 wire _12280_;
 wire _12281_;
 wire _12282_;
 wire _12283_;
 wire _12284_;
 wire _12285_;
 wire _12286_;
 wire _12287_;
 wire _12288_;
 wire _12289_;
 wire _12290_;
 wire _12291_;
 wire _12292_;
 wire _12293_;
 wire _12294_;
 wire _12295_;
 wire _12296_;
 wire _12297_;
 wire _12298_;
 wire _12299_;
 wire _12300_;
 wire _12301_;
 wire _12302_;
 wire _12303_;
 wire _12304_;
 wire _12305_;
 wire _12306_;
 wire _12307_;
 wire _12308_;
 wire _12309_;
 wire _12310_;
 wire _12311_;
 wire _12312_;
 wire _12313_;
 wire _12314_;
 wire _12315_;
 wire _12316_;
 wire _12317_;
 wire _12318_;
 wire _12319_;
 wire _12320_;
 wire _12321_;
 wire _12322_;
 wire _12323_;
 wire _12324_;
 wire _12325_;
 wire _12326_;
 wire _12327_;
 wire _12328_;
 wire _12329_;
 wire _12330_;
 wire _12331_;
 wire _12332_;
 wire _12333_;
 wire _12334_;
 wire _12335_;
 wire _12336_;
 wire _12337_;
 wire _12338_;
 wire _12339_;
 wire _12340_;
 wire _12341_;
 wire _12342_;
 wire _12343_;
 wire _12344_;
 wire _12345_;
 wire _12346_;
 wire _12347_;
 wire _12348_;
 wire _12349_;
 wire _12350_;
 wire _12351_;
 wire _12352_;
 wire _12353_;
 wire _12354_;
 wire _12355_;
 wire _12356_;
 wire _12357_;
 wire _12358_;
 wire _12359_;
 wire _12360_;
 wire _12361_;
 wire _12362_;
 wire _12363_;
 wire _12364_;
 wire _12365_;
 wire _12366_;
 wire _12367_;
 wire _12368_;
 wire _12369_;
 wire _12370_;
 wire _12371_;
 wire _12372_;
 wire _12373_;
 wire _12374_;
 wire _12375_;
 wire _12376_;
 wire _12377_;
 wire _12378_;
 wire _12379_;
 wire _12380_;
 wire _12381_;
 wire _12382_;
 wire _12383_;
 wire _12384_;
 wire _12385_;
 wire _12386_;
 wire _12387_;
 wire _12388_;
 wire _12389_;
 wire _12390_;
 wire _12391_;
 wire _12392_;
 wire _12393_;
 wire _12394_;
 wire _12395_;
 wire _12396_;
 wire _12397_;
 wire _12398_;
 wire _12399_;
 wire _12400_;
 wire _12401_;
 wire _12402_;
 wire _12403_;
 wire _12404_;
 wire _12405_;
 wire _12406_;
 wire _12407_;
 wire _12408_;
 wire _12409_;
 wire _12410_;
 wire _12411_;
 wire _12412_;
 wire _12413_;
 wire _12414_;
 wire _12415_;
 wire _12416_;
 wire _12417_;
 wire _12418_;
 wire _12419_;
 wire _12420_;
 wire _12421_;
 wire _12422_;
 wire _12423_;
 wire _12424_;
 wire _12425_;
 wire _12426_;
 wire _12427_;
 wire _12428_;
 wire _12429_;
 wire _12430_;
 wire _12431_;
 wire _12432_;
 wire _12433_;
 wire _12434_;
 wire _12435_;
 wire _12436_;
 wire _12437_;
 wire _12438_;
 wire _12439_;
 wire _12440_;
 wire _12441_;
 wire _12442_;
 wire _12443_;
 wire _12444_;
 wire _12445_;
 wire _12446_;
 wire _12447_;
 wire _12448_;
 wire _12449_;
 wire _12450_;
 wire _12451_;
 wire _12452_;
 wire _12453_;
 wire _12454_;
 wire _12455_;
 wire _12456_;
 wire _12457_;
 wire _12458_;
 wire _12459_;
 wire _12460_;
 wire _12461_;
 wire _12462_;
 wire _12463_;
 wire _12464_;
 wire _12465_;
 wire _12466_;
 wire _12467_;
 wire _12468_;
 wire _12469_;
 wire _12470_;
 wire _12471_;
 wire _12472_;
 wire _12473_;
 wire _12474_;
 wire _12475_;
 wire _12476_;
 wire _12477_;
 wire _12478_;
 wire _12479_;
 wire _12480_;
 wire _12481_;
 wire _12482_;
 wire _12483_;
 wire _12484_;
 wire _12485_;
 wire _12486_;
 wire _12487_;
 wire _12488_;
 wire _12489_;
 wire _12490_;
 wire _12491_;
 wire _12492_;
 wire _12493_;
 wire _12494_;
 wire _12495_;
 wire _12496_;
 wire _12497_;
 wire _12498_;
 wire _12499_;
 wire _12500_;
 wire _12501_;
 wire _12502_;
 wire _12503_;
 wire _12504_;
 wire _12505_;
 wire _12506_;
 wire _12507_;
 wire _12508_;
 wire _12509_;
 wire _12510_;
 wire _12511_;
 wire _12512_;
 wire _12513_;
 wire _12514_;
 wire _12515_;
 wire _12516_;
 wire _12517_;
 wire _12518_;
 wire _12519_;
 wire _12520_;
 wire _12521_;
 wire _12522_;
 wire _12523_;
 wire _12524_;
 wire _12525_;
 wire _12526_;
 wire _12527_;
 wire _12528_;
 wire _12529_;
 wire _12530_;
 wire _12531_;
 wire _12532_;
 wire _12533_;
 wire _12534_;
 wire _12535_;
 wire _12536_;
 wire _12537_;
 wire _12538_;
 wire _12539_;
 wire _12540_;
 wire _12541_;
 wire _12542_;
 wire _12543_;
 wire _12544_;
 wire _12545_;
 wire _12546_;
 wire _12547_;
 wire _12548_;
 wire _12549_;
 wire _12550_;
 wire _12551_;
 wire _12552_;
 wire _12553_;
 wire _12554_;
 wire _12555_;
 wire _12556_;
 wire _12557_;
 wire _12558_;
 wire _12559_;
 wire _12560_;
 wire _12561_;
 wire _12562_;
 wire _12563_;
 wire _12564_;
 wire _12565_;
 wire _12566_;
 wire _12567_;
 wire _12568_;
 wire _12569_;
 wire _12570_;
 wire _12571_;
 wire _12572_;
 wire _12573_;
 wire _12574_;
 wire _12575_;
 wire _12576_;
 wire _12577_;
 wire _12578_;
 wire _12579_;
 wire _12580_;
 wire _12581_;
 wire _12582_;
 wire _12583_;
 wire _12584_;
 wire _12585_;
 wire _12586_;
 wire _12587_;
 wire _12588_;
 wire _12589_;
 wire _12590_;
 wire _12591_;
 wire _12592_;
 wire _12593_;
 wire _12594_;
 wire _12595_;
 wire _12596_;
 wire _12597_;
 wire _12598_;
 wire _12599_;
 wire _12600_;
 wire _12601_;
 wire _12602_;
 wire _12603_;
 wire _12604_;
 wire _12605_;
 wire _12606_;
 wire _12607_;
 wire _12608_;
 wire _12609_;
 wire _12610_;
 wire _12611_;
 wire _12612_;
 wire _12613_;
 wire _12614_;
 wire _12615_;
 wire _12616_;
 wire _12617_;
 wire _12618_;
 wire _12619_;
 wire _12620_;
 wire _12621_;
 wire _12622_;
 wire _12623_;
 wire _12624_;
 wire _12625_;
 wire _12626_;
 wire _12627_;
 wire _12628_;
 wire _12629_;
 wire _12630_;
 wire _12631_;
 wire _12632_;
 wire _12633_;
 wire _12634_;
 wire _12635_;
 wire _12636_;
 wire _12637_;
 wire _12638_;
 wire _12639_;
 wire _12640_;
 wire _12641_;
 wire _12642_;
 wire _12643_;
 wire _12644_;
 wire _12645_;
 wire _12646_;
 wire _12647_;
 wire _12648_;
 wire _12649_;
 wire _12650_;
 wire _12651_;
 wire _12652_;
 wire _12653_;
 wire _12654_;
 wire _12655_;
 wire _12656_;
 wire _12657_;
 wire _12658_;
 wire _12659_;
 wire _12660_;
 wire _12661_;
 wire _12662_;
 wire _12663_;
 wire _12664_;
 wire _12665_;
 wire _12666_;
 wire _12667_;
 wire _12668_;
 wire _12669_;
 wire _12670_;
 wire _12671_;
 wire _12672_;
 wire _12673_;
 wire _12674_;
 wire _12675_;
 wire _12676_;
 wire _12677_;
 wire _12678_;
 wire _12679_;
 wire _12680_;
 wire _12681_;
 wire _12682_;
 wire _12683_;
 wire _12684_;
 wire _12685_;
 wire _12686_;
 wire _12687_;
 wire _12688_;
 wire _12689_;
 wire _12690_;
 wire _12691_;
 wire _12692_;
 wire _12693_;
 wire _12694_;
 wire _12695_;
 wire _12696_;
 wire _12697_;
 wire _12698_;
 wire _12699_;
 wire _12700_;
 wire _12701_;
 wire _12702_;
 wire _12703_;
 wire _12704_;
 wire _12705_;
 wire _12706_;
 wire _12707_;
 wire _12708_;
 wire _12709_;
 wire _12710_;
 wire _12711_;
 wire _12712_;
 wire _12713_;
 wire _12714_;
 wire _12715_;
 wire _12716_;
 wire _12717_;
 wire _12718_;
 wire _12719_;
 wire _12720_;
 wire _12721_;
 wire _12722_;
 wire _12723_;
 wire _12724_;
 wire _12725_;
 wire _12726_;
 wire _12727_;
 wire _12728_;
 wire _12729_;
 wire _12730_;
 wire _12731_;
 wire _12732_;
 wire _12733_;
 wire _12734_;
 wire _12735_;
 wire _12736_;
 wire _12737_;
 wire _12738_;
 wire _12739_;
 wire _12740_;
 wire _12741_;
 wire _12742_;
 wire _12743_;
 wire _12744_;
 wire _12745_;
 wire _12746_;
 wire _12747_;
 wire _12748_;
 wire _12749_;
 wire _12750_;
 wire _12751_;
 wire _12752_;
 wire _12753_;
 wire _12754_;
 wire _12755_;
 wire _12756_;
 wire _12757_;
 wire _12758_;
 wire _12759_;
 wire _12760_;
 wire _12761_;
 wire _12762_;
 wire _12763_;
 wire _12764_;
 wire _12765_;
 wire _12766_;
 wire _12767_;
 wire _12768_;
 wire _12769_;
 wire _12770_;
 wire _12771_;
 wire _12772_;
 wire _12773_;
 wire _12774_;
 wire _12775_;
 wire _12776_;
 wire _12777_;
 wire _12778_;
 wire _12779_;
 wire _12780_;
 wire _12781_;
 wire _12782_;
 wire _12783_;
 wire _12784_;
 wire _12785_;
 wire _12786_;
 wire _12787_;
 wire _12788_;
 wire _12789_;
 wire _12790_;
 wire _12791_;
 wire _12792_;
 wire _12793_;
 wire _12794_;
 wire _12795_;
 wire _12796_;
 wire _12797_;
 wire _12798_;
 wire _12799_;
 wire _12800_;
 wire _12801_;
 wire _12802_;
 wire _12803_;
 wire _12804_;
 wire _12805_;
 wire _12806_;
 wire _12807_;
 wire _12808_;
 wire _12809_;
 wire _12810_;
 wire _12811_;
 wire _12812_;
 wire _12813_;
 wire _12814_;
 wire _12815_;
 wire _12816_;
 wire _12817_;
 wire _12818_;
 wire _12819_;
 wire _12820_;
 wire _12821_;
 wire _12822_;
 wire _12823_;
 wire _12824_;
 wire _12825_;
 wire _12826_;
 wire _12827_;
 wire _12828_;
 wire _12829_;
 wire _12830_;
 wire _12831_;
 wire _12832_;
 wire _12833_;
 wire _12834_;
 wire _12835_;
 wire _12836_;
 wire _12837_;
 wire _12838_;
 wire _12839_;
 wire _12840_;
 wire _12841_;
 wire _12842_;
 wire _12843_;
 wire _12844_;
 wire _12845_;
 wire _12846_;
 wire _12847_;
 wire _12848_;
 wire _12849_;
 wire _12850_;
 wire _12851_;
 wire _12852_;
 wire _12853_;
 wire _12854_;
 wire _12855_;
 wire _12856_;
 wire _12857_;
 wire _12858_;
 wire _12859_;
 wire _12860_;
 wire _12861_;
 wire _12862_;
 wire _12863_;
 wire _12864_;
 wire _12865_;
 wire _12866_;
 wire _12867_;
 wire _12868_;
 wire _12869_;
 wire _12870_;
 wire _12871_;
 wire _12872_;
 wire _12873_;
 wire _12874_;
 wire _12875_;
 wire _12876_;
 wire _12877_;
 wire _12878_;
 wire _12879_;
 wire _12880_;
 wire _12881_;
 wire _12882_;
 wire _12883_;
 wire _12884_;
 wire _12885_;
 wire _12886_;
 wire _12887_;
 wire _12888_;
 wire _12889_;
 wire _12890_;
 wire _12891_;
 wire _12892_;
 wire _12893_;
 wire _12894_;
 wire _12895_;
 wire _12896_;
 wire _12897_;
 wire _12898_;
 wire _12899_;
 wire _12900_;
 wire _12901_;
 wire _12902_;
 wire _12903_;
 wire _12904_;
 wire _12905_;
 wire _12906_;
 wire _12907_;
 wire _12908_;
 wire _12909_;
 wire _12910_;
 wire _12911_;
 wire _12912_;
 wire _12913_;
 wire _12914_;
 wire _12915_;
 wire _12916_;
 wire _12917_;
 wire _12918_;
 wire _12919_;
 wire _12920_;
 wire _12921_;
 wire _12922_;
 wire _12923_;
 wire _12924_;
 wire _12925_;
 wire _12926_;
 wire _12927_;
 wire _12928_;
 wire _12929_;
 wire _12930_;
 wire _12931_;
 wire _12932_;
 wire _12933_;
 wire _12934_;
 wire _12935_;
 wire _12936_;
 wire _12937_;
 wire _12938_;
 wire _12939_;
 wire _12940_;
 wire _12941_;
 wire _12942_;
 wire _12943_;
 wire _12944_;
 wire _12945_;
 wire _12946_;
 wire _12947_;
 wire _12948_;
 wire _12949_;
 wire _12950_;
 wire _12951_;
 wire _12952_;
 wire _12953_;
 wire _12954_;
 wire _12955_;
 wire _12956_;
 wire _12957_;
 wire _12958_;
 wire _12959_;
 wire _12960_;
 wire _12961_;
 wire _12962_;
 wire _12963_;
 wire _12964_;
 wire _12965_;
 wire _12966_;
 wire _12967_;
 wire _12968_;
 wire _12969_;
 wire _12970_;
 wire _12971_;
 wire _12972_;
 wire _12973_;
 wire _12974_;
 wire _12975_;
 wire _12976_;
 wire _12977_;
 wire _12978_;
 wire _12979_;
 wire _12980_;
 wire _12981_;
 wire _12982_;
 wire _12983_;
 wire _12984_;
 wire _12985_;
 wire _12986_;
 wire _12987_;
 wire _12988_;
 wire _12989_;
 wire _12990_;
 wire _12991_;
 wire _12992_;
 wire _12993_;
 wire _12994_;
 wire _12995_;
 wire _12996_;
 wire _12997_;
 wire _12998_;
 wire _12999_;
 wire _13000_;
 wire _13001_;
 wire _13002_;
 wire _13003_;
 wire _13004_;
 wire _13005_;
 wire _13006_;
 wire _13007_;
 wire _13008_;
 wire _13009_;
 wire _13010_;
 wire _13011_;
 wire _13012_;
 wire _13013_;
 wire _13014_;
 wire _13015_;
 wire _13016_;
 wire _13017_;
 wire _13018_;
 wire _13019_;
 wire _13020_;
 wire _13021_;
 wire _13022_;
 wire _13023_;
 wire _13024_;
 wire _13025_;
 wire _13026_;
 wire _13027_;
 wire _13028_;
 wire _13029_;
 wire _13030_;
 wire _13031_;
 wire _13032_;
 wire _13033_;
 wire _13034_;
 wire _13035_;
 wire _13036_;
 wire _13037_;
 wire _13038_;
 wire _13039_;
 wire _13040_;
 wire _13041_;
 wire _13042_;
 wire _13043_;
 wire _13044_;
 wire _13045_;
 wire _13046_;
 wire _13047_;
 wire _13048_;
 wire _13049_;
 wire _13050_;
 wire _13051_;
 wire _13052_;
 wire _13053_;
 wire _13054_;
 wire _13055_;
 wire _13056_;
 wire _13057_;
 wire _13058_;
 wire _13059_;
 wire _13060_;
 wire _13061_;
 wire _13062_;
 wire _13063_;
 wire _13064_;
 wire _13065_;
 wire _13066_;
 wire _13067_;
 wire _13068_;
 wire _13069_;
 wire _13070_;
 wire _13071_;
 wire _13072_;
 wire _13073_;
 wire _13074_;
 wire _13075_;
 wire _13076_;
 wire _13077_;
 wire _13078_;
 wire _13079_;
 wire _13080_;
 wire _13081_;
 wire _13082_;
 wire _13083_;
 wire _13084_;
 wire _13085_;
 wire _13086_;
 wire _13087_;
 wire _13088_;
 wire _13089_;
 wire _13090_;
 wire _13091_;
 wire _13092_;
 wire _13093_;
 wire _13094_;
 wire _13095_;
 wire _13096_;
 wire _13097_;
 wire _13098_;
 wire _13099_;
 wire _13100_;
 wire _13101_;
 wire _13102_;
 wire _13103_;
 wire _13104_;
 wire _13105_;
 wire _13106_;
 wire _13107_;
 wire _13108_;
 wire _13109_;
 wire _13110_;
 wire _13111_;
 wire _13112_;
 wire _13113_;
 wire _13114_;
 wire _13115_;
 wire _13116_;
 wire _13117_;
 wire _13118_;
 wire _13119_;
 wire _13120_;
 wire _13121_;
 wire _13122_;
 wire _13123_;
 wire _13124_;
 wire _13125_;
 wire _13126_;
 wire _13127_;
 wire _13128_;
 wire _13129_;
 wire _13130_;
 wire _13131_;
 wire _13132_;
 wire _13133_;
 wire _13134_;
 wire _13135_;
 wire _13136_;
 wire _13137_;
 wire _13138_;
 wire _13139_;
 wire _13140_;
 wire _13141_;
 wire _13142_;
 wire _13143_;
 wire _13144_;
 wire _13145_;
 wire _13146_;
 wire _13147_;
 wire _13148_;
 wire _13149_;
 wire _13150_;
 wire _13151_;
 wire _13152_;
 wire _13153_;
 wire _13154_;
 wire _13155_;
 wire _13156_;
 wire _13157_;
 wire _13158_;
 wire _13159_;
 wire _13160_;
 wire _13161_;
 wire _13162_;
 wire _13163_;
 wire _13164_;
 wire _13165_;
 wire _13166_;
 wire _13167_;
 wire _13168_;
 wire _13169_;
 wire _13170_;
 wire _13171_;
 wire _13172_;
 wire _13173_;
 wire _13174_;
 wire _13175_;
 wire _13176_;
 wire _13177_;
 wire _13178_;
 wire _13179_;
 wire _13180_;
 wire _13181_;
 wire _13182_;
 wire _13183_;
 wire _13184_;
 wire _13185_;
 wire _13186_;
 wire _13187_;
 wire _13188_;
 wire _13189_;
 wire _13190_;
 wire _13191_;
 wire _13192_;
 wire _13193_;
 wire _13194_;
 wire _13195_;
 wire _13196_;
 wire _13197_;
 wire _13198_;
 wire _13199_;
 wire _13200_;
 wire _13201_;
 wire _13202_;
 wire _13203_;
 wire _13204_;
 wire _13205_;
 wire _13206_;
 wire _13207_;
 wire _13208_;
 wire _13209_;
 wire _13210_;
 wire _13211_;
 wire _13212_;
 wire _13213_;
 wire _13214_;
 wire _13215_;
 wire _13216_;
 wire _13217_;
 wire _13218_;
 wire _13219_;
 wire _13220_;
 wire _13221_;
 wire _13222_;
 wire _13223_;
 wire _13224_;
 wire _13225_;
 wire _13226_;
 wire _13227_;
 wire _13228_;
 wire _13229_;
 wire _13230_;
 wire _13231_;
 wire _13232_;
 wire _13233_;
 wire _13234_;
 wire _13235_;
 wire _13236_;
 wire _13237_;
 wire _13238_;
 wire _13239_;
 wire _13240_;
 wire _13241_;
 wire _13242_;
 wire _13243_;
 wire _13244_;
 wire _13245_;
 wire _13246_;
 wire _13247_;
 wire _13248_;
 wire _13249_;
 wire _13250_;
 wire _13251_;
 wire _13252_;
 wire _13253_;
 wire _13254_;
 wire _13255_;
 wire _13256_;
 wire _13257_;
 wire _13258_;
 wire _13259_;
 wire _13260_;
 wire _13261_;
 wire _13262_;
 wire _13263_;
 wire _13264_;
 wire _13265_;
 wire _13266_;
 wire _13267_;
 wire _13268_;
 wire _13269_;
 wire _13270_;
 wire _13271_;
 wire _13272_;
 wire _13273_;
 wire _13274_;
 wire _13275_;
 wire _13276_;
 wire _13277_;
 wire _13278_;
 wire _13279_;
 wire _13280_;
 wire _13281_;
 wire _13282_;
 wire _13283_;
 wire _13284_;
 wire _13285_;
 wire _13286_;
 wire _13287_;
 wire _13288_;
 wire _13289_;
 wire _13290_;
 wire _13291_;
 wire _13292_;
 wire _13293_;
 wire _13294_;
 wire _13295_;
 wire _13296_;
 wire _13297_;
 wire _13298_;
 wire _13299_;
 wire _13300_;
 wire _13301_;
 wire _13302_;
 wire _13303_;
 wire _13304_;
 wire _13305_;
 wire _13306_;
 wire _13307_;
 wire _13308_;
 wire _13309_;
 wire _13310_;
 wire _13311_;
 wire _13312_;
 wire _13313_;
 wire _13314_;
 wire _13315_;
 wire _13316_;
 wire _13317_;
 wire _13318_;
 wire _13319_;
 wire _13320_;
 wire _13321_;
 wire _13322_;
 wire _13323_;
 wire _13324_;
 wire _13325_;
 wire _13326_;
 wire _13327_;
 wire _13328_;
 wire _13329_;
 wire _13330_;
 wire _13331_;
 wire _13332_;
 wire _13333_;
 wire _13334_;
 wire _13335_;
 wire _13336_;
 wire _13337_;
 wire _13338_;
 wire _13339_;
 wire _13340_;
 wire _13341_;
 wire _13342_;
 wire _13343_;
 wire _13344_;
 wire _13345_;
 wire _13346_;
 wire _13347_;
 wire _13348_;
 wire _13349_;
 wire _13350_;
 wire _13351_;
 wire _13352_;
 wire _13353_;
 wire _13354_;
 wire _13355_;
 wire _13356_;
 wire _13357_;
 wire _13358_;
 wire _13359_;
 wire _13360_;
 wire _13361_;
 wire _13362_;
 wire _13363_;
 wire _13364_;
 wire _13365_;
 wire _13366_;
 wire _13367_;
 wire _13368_;
 wire _13369_;
 wire _13370_;
 wire _13371_;
 wire _13372_;
 wire _13373_;
 wire _13374_;
 wire _13375_;
 wire _13376_;
 wire _13377_;
 wire _13378_;
 wire _13379_;
 wire _13380_;
 wire _13381_;
 wire _13382_;
 wire _13383_;
 wire _13384_;
 wire _13385_;
 wire _13386_;
 wire _13387_;
 wire _13388_;
 wire _13389_;
 wire _13390_;
 wire _13391_;
 wire _13392_;
 wire _13393_;
 wire _13394_;
 wire _13395_;
 wire _13396_;
 wire _13397_;
 wire _13398_;
 wire _13399_;
 wire _13400_;
 wire _13401_;
 wire _13402_;
 wire _13403_;
 wire _13404_;
 wire _13405_;
 wire _13406_;
 wire _13407_;
 wire _13408_;
 wire _13409_;
 wire _13410_;
 wire _13411_;
 wire _13412_;
 wire _13413_;
 wire _13414_;
 wire _13415_;
 wire _13416_;
 wire _13417_;
 wire _13418_;
 wire _13419_;
 wire _13420_;
 wire _13421_;
 wire _13422_;
 wire _13423_;
 wire _13424_;
 wire _13425_;
 wire _13426_;
 wire _13427_;
 wire _13428_;
 wire _13429_;
 wire _13430_;
 wire _13431_;
 wire _13432_;
 wire _13433_;
 wire _13434_;
 wire _13435_;
 wire _13436_;
 wire _13437_;
 wire _13438_;
 wire _13439_;
 wire _13440_;
 wire _13441_;
 wire _13442_;
 wire _13443_;
 wire _13444_;
 wire _13445_;
 wire _13446_;
 wire _13447_;
 wire _13448_;
 wire _13449_;
 wire _13450_;
 wire _13451_;
 wire _13452_;
 wire _13453_;
 wire _13454_;
 wire _13455_;
 wire _13456_;
 wire _13457_;
 wire _13458_;
 wire _13459_;
 wire _13460_;
 wire _13461_;
 wire _13462_;
 wire _13463_;
 wire _13464_;
 wire _13465_;
 wire _13466_;
 wire _13467_;
 wire _13468_;
 wire _13469_;
 wire _13470_;
 wire _13471_;
 wire _13472_;
 wire _13473_;
 wire _13474_;
 wire _13475_;
 wire _13476_;
 wire _13477_;
 wire _13478_;
 wire _13479_;
 wire _13480_;
 wire _13481_;
 wire _13482_;
 wire _13483_;
 wire _13484_;
 wire _13485_;
 wire _13486_;
 wire _13487_;
 wire _13488_;
 wire _13489_;
 wire _13490_;
 wire _13491_;
 wire _13492_;
 wire _13493_;
 wire _13494_;
 wire _13495_;
 wire _13496_;
 wire _13497_;
 wire _13498_;
 wire _13499_;
 wire _13500_;
 wire _13501_;
 wire _13502_;
 wire _13503_;
 wire _13504_;
 wire _13505_;
 wire _13506_;
 wire _13507_;
 wire _13508_;
 wire _13509_;
 wire _13510_;
 wire _13511_;
 wire _13512_;
 wire _13513_;
 wire _13514_;
 wire _13515_;
 wire _13516_;
 wire _13517_;
 wire _13518_;
 wire _13519_;
 wire _13520_;
 wire _13521_;
 wire _13522_;
 wire _13523_;
 wire _13524_;
 wire _13525_;
 wire _13526_;
 wire _13527_;
 wire _13528_;
 wire _13529_;
 wire _13530_;
 wire _13531_;
 wire _13532_;
 wire _13533_;
 wire _13534_;
 wire _13535_;
 wire _13536_;
 wire _13537_;
 wire _13538_;
 wire _13539_;
 wire _13540_;
 wire _13541_;
 wire _13542_;
 wire _13543_;
 wire _13544_;
 wire _13545_;
 wire _13546_;
 wire _13547_;
 wire _13548_;
 wire _13549_;
 wire _13550_;
 wire _13551_;
 wire _13552_;
 wire _13553_;
 wire _13554_;
 wire _13555_;
 wire _13556_;
 wire _13557_;
 wire _13558_;
 wire _13559_;
 wire _13560_;
 wire _13561_;
 wire _13562_;
 wire _13563_;
 wire _13564_;
 wire _13565_;
 wire _13566_;
 wire _13567_;
 wire _13568_;
 wire _13569_;
 wire _13570_;
 wire _13571_;
 wire _13572_;
 wire _13573_;
 wire _13574_;
 wire _13575_;
 wire _13576_;
 wire _13577_;
 wire _13578_;
 wire _13579_;
 wire _13580_;
 wire _13581_;
 wire _13582_;
 wire _13583_;
 wire _13584_;
 wire _13585_;
 wire _13586_;
 wire _13587_;
 wire _13588_;
 wire _13589_;
 wire _13590_;
 wire _13591_;
 wire _13592_;
 wire _13593_;
 wire _13594_;
 wire _13595_;
 wire _13596_;
 wire _13597_;
 wire _13598_;
 wire _13599_;
 wire _13600_;
 wire _13601_;
 wire _13602_;
 wire _13603_;
 wire _13604_;
 wire _13605_;
 wire _13606_;
 wire _13607_;
 wire _13608_;
 wire _13609_;
 wire _13610_;
 wire _13611_;
 wire _13612_;
 wire _13613_;
 wire _13614_;
 wire _13615_;
 wire _13616_;
 wire _13617_;
 wire _13618_;
 wire _13619_;
 wire _13620_;
 wire _13621_;
 wire _13622_;
 wire _13623_;
 wire _13624_;
 wire _13625_;
 wire _13626_;
 wire _13627_;
 wire _13628_;
 wire _13629_;
 wire _13630_;
 wire _13631_;
 wire _13632_;
 wire _13633_;
 wire _13634_;
 wire _13635_;
 wire _13636_;
 wire _13637_;
 wire _13638_;
 wire _13639_;
 wire _13640_;
 wire _13641_;
 wire _13642_;
 wire _13643_;
 wire _13644_;
 wire _13645_;
 wire _13646_;
 wire _13647_;
 wire _13648_;
 wire _13649_;
 wire _13650_;
 wire _13651_;
 wire _13652_;
 wire _13653_;
 wire _13654_;
 wire _13655_;
 wire _13656_;
 wire _13657_;
 wire _13658_;
 wire _13659_;
 wire _13660_;
 wire _13661_;
 wire _13662_;
 wire _13663_;
 wire _13664_;
 wire _13665_;
 wire _13666_;
 wire _13667_;
 wire _13668_;
 wire _13669_;
 wire _13670_;
 wire _13671_;
 wire _13672_;
 wire _13673_;
 wire _13674_;
 wire _13675_;
 wire _13676_;
 wire _13677_;
 wire _13678_;
 wire _13679_;
 wire _13680_;
 wire _13681_;
 wire _13682_;
 wire _13683_;
 wire _13684_;
 wire _13685_;
 wire _13686_;
 wire _13687_;
 wire _13688_;
 wire _13689_;
 wire _13690_;
 wire _13691_;
 wire _13692_;
 wire _13693_;
 wire _13694_;
 wire _13695_;
 wire _13696_;
 wire _13697_;
 wire _13698_;
 wire _13699_;
 wire _13700_;
 wire _13701_;
 wire _13702_;
 wire _13703_;
 wire _13704_;
 wire _13705_;
 wire _13706_;
 wire _13707_;
 wire _13708_;
 wire _13709_;
 wire _13710_;
 wire _13711_;
 wire _13712_;
 wire _13713_;
 wire _13714_;
 wire _13715_;
 wire _13716_;
 wire _13717_;
 wire _13718_;
 wire _13719_;
 wire _13720_;
 wire _13721_;
 wire _13722_;
 wire _13723_;
 wire _13724_;
 wire _13725_;
 wire _13726_;
 wire _13727_;
 wire _13728_;
 wire _13729_;
 wire _13730_;
 wire _13731_;
 wire _13732_;
 wire _13733_;
 wire _13734_;
 wire _13735_;
 wire _13736_;
 wire _13737_;
 wire _13738_;
 wire _13739_;
 wire _13740_;
 wire _13741_;
 wire _13742_;
 wire _13743_;
 wire _13744_;
 wire _13745_;
 wire _13746_;
 wire _13747_;
 wire _13748_;
 wire _13749_;
 wire _13750_;
 wire _13751_;
 wire _13752_;
 wire _13753_;
 wire _13754_;
 wire _13755_;
 wire _13756_;
 wire _13757_;
 wire _13758_;
 wire _13759_;
 wire _13760_;
 wire _13761_;
 wire _13762_;
 wire _13763_;
 wire _13764_;
 wire _13765_;
 wire _13766_;
 wire _13767_;
 wire _13768_;
 wire _13769_;
 wire _13770_;
 wire _13771_;
 wire _13772_;
 wire _13773_;
 wire _13774_;
 wire _13775_;
 wire _13776_;
 wire _13777_;
 wire _13778_;
 wire _13779_;
 wire _13780_;
 wire _13781_;
 wire _13782_;
 wire _13783_;
 wire _13784_;
 wire _13785_;
 wire _13786_;
 wire _13787_;
 wire _13788_;
 wire _13789_;
 wire _13790_;
 wire _13791_;
 wire _13792_;
 wire _13793_;
 wire _13794_;
 wire _13795_;
 wire _13796_;
 wire _13797_;
 wire _13798_;
 wire _13799_;
 wire _13800_;
 wire _13801_;
 wire _13802_;
 wire _13803_;
 wire _13804_;
 wire _13805_;
 wire _13806_;
 wire _13807_;
 wire _13808_;
 wire _13809_;
 wire _13810_;
 wire _13811_;
 wire _13812_;
 wire _13813_;
 wire _13814_;
 wire _13815_;
 wire _13816_;
 wire _13817_;
 wire _13818_;
 wire _13819_;
 wire _13820_;
 wire _13821_;
 wire _13822_;
 wire _13823_;
 wire _13824_;
 wire _13825_;
 wire _13826_;
 wire _13827_;
 wire _13828_;
 wire _13829_;
 wire _13830_;
 wire _13831_;
 wire _13832_;
 wire _13833_;
 wire _13834_;
 wire _13835_;
 wire _13836_;
 wire _13837_;
 wire _13838_;
 wire _13839_;
 wire _13840_;
 wire _13841_;
 wire _13842_;
 wire _13843_;
 wire _13844_;
 wire _13845_;
 wire _13846_;
 wire _13847_;
 wire _13848_;
 wire _13849_;
 wire _13850_;
 wire _13851_;
 wire _13852_;
 wire _13853_;
 wire _13854_;
 wire _13855_;
 wire _13856_;
 wire _13857_;
 wire _13858_;
 wire _13859_;
 wire _13860_;
 wire _13861_;
 wire _13862_;
 wire _13863_;
 wire _13864_;
 wire _13865_;
 wire _13866_;
 wire _13867_;
 wire _13868_;
 wire _13869_;
 wire _13870_;
 wire _13871_;
 wire _13872_;
 wire _13873_;
 wire _13874_;
 wire _13875_;
 wire _13876_;
 wire _13877_;
 wire _13878_;
 wire _13879_;
 wire _13880_;
 wire _13881_;
 wire _13882_;
 wire _13883_;
 wire _13884_;
 wire _13885_;
 wire _13886_;
 wire _13887_;
 wire _13888_;
 wire _13889_;
 wire _13890_;
 wire _13891_;
 wire _13892_;
 wire _13893_;
 wire _13894_;
 wire _13895_;
 wire _13896_;
 wire _13897_;
 wire _13898_;
 wire _13899_;
 wire _13900_;
 wire _13901_;
 wire _13902_;
 wire _13903_;
 wire _13904_;
 wire _13905_;
 wire _13906_;
 wire _13907_;
 wire _13908_;
 wire _13909_;
 wire _13910_;
 wire _13911_;
 wire _13912_;
 wire _13913_;
 wire _13914_;
 wire _13915_;
 wire _13916_;
 wire _13917_;
 wire _13918_;
 wire _13919_;
 wire _13920_;
 wire _13921_;
 wire _13922_;
 wire _13923_;
 wire _13924_;
 wire _13925_;
 wire _13926_;
 wire _13927_;
 wire _13928_;
 wire _13929_;
 wire _13930_;
 wire _13931_;
 wire _13932_;
 wire _13933_;
 wire _13934_;
 wire _13935_;
 wire _13936_;
 wire _13937_;
 wire _13938_;
 wire _13939_;
 wire _13940_;
 wire _13941_;
 wire _13942_;
 wire _13943_;
 wire _13944_;
 wire _13945_;
 wire _13946_;
 wire _13947_;
 wire _13948_;
 wire _13949_;
 wire _13950_;
 wire _13951_;
 wire _13952_;
 wire _13953_;
 wire _13954_;
 wire _13955_;
 wire _13956_;
 wire _13957_;
 wire _13958_;
 wire _13959_;
 wire _13960_;
 wire _13961_;
 wire _13962_;
 wire _13963_;
 wire _13964_;
 wire _13965_;
 wire _13966_;
 wire _13967_;
 wire _13968_;
 wire _13969_;
 wire _13970_;
 wire _13971_;
 wire _13972_;
 wire _13973_;
 wire _13974_;
 wire _13975_;
 wire _13976_;
 wire _13977_;
 wire _13978_;
 wire _13979_;
 wire _13980_;
 wire _13981_;
 wire _13982_;
 wire _13983_;
 wire _13984_;
 wire _13985_;
 wire _13986_;
 wire _13987_;
 wire _13988_;
 wire _13989_;
 wire _13990_;
 wire _13991_;
 wire _13992_;
 wire _13993_;
 wire _13994_;
 wire _13995_;
 wire _13996_;
 wire _13997_;
 wire _13998_;
 wire _13999_;
 wire _14000_;
 wire _14001_;
 wire _14002_;
 wire _14003_;
 wire _14004_;
 wire _14005_;
 wire _14006_;
 wire _14007_;
 wire _14008_;
 wire _14009_;
 wire _14010_;
 wire _14011_;
 wire _14012_;
 wire _14013_;
 wire _14014_;
 wire _14015_;
 wire _14016_;
 wire _14017_;
 wire _14018_;
 wire _14019_;
 wire _14020_;
 wire _14021_;
 wire _14022_;
 wire _14023_;
 wire _14024_;
 wire _14025_;
 wire _14026_;
 wire _14027_;
 wire _14028_;
 wire _14029_;
 wire _14030_;
 wire _14031_;
 wire _14032_;
 wire _14033_;
 wire _14034_;
 wire _14035_;
 wire _14036_;
 wire _14037_;
 wire _14038_;
 wire _14039_;
 wire _14040_;
 wire _14041_;
 wire _14042_;
 wire _14043_;
 wire _14044_;
 wire _14045_;
 wire _14046_;
 wire _14047_;
 wire _14048_;
 wire _14049_;
 wire _14050_;
 wire _14051_;
 wire _14052_;
 wire _14053_;
 wire _14054_;
 wire _14055_;
 wire _14056_;
 wire _14057_;
 wire _14058_;
 wire _14059_;
 wire _14060_;
 wire _14061_;
 wire _14062_;
 wire _14063_;
 wire _14064_;
 wire _14065_;
 wire _14066_;
 wire _14067_;
 wire _14068_;
 wire _14069_;
 wire _14070_;
 wire _14071_;
 wire _14072_;
 wire _14073_;
 wire _14074_;
 wire _14075_;
 wire _14076_;
 wire _14077_;
 wire _14078_;
 wire _14079_;
 wire _14080_;
 wire _14081_;
 wire _14082_;
 wire _14083_;
 wire _14084_;
 wire _14085_;
 wire _14086_;
 wire _14087_;
 wire _14088_;
 wire _14089_;
 wire _14090_;
 wire _14091_;
 wire _14092_;
 wire _14093_;
 wire _14094_;
 wire _14095_;
 wire _14096_;
 wire _14097_;
 wire _14098_;
 wire _14099_;
 wire _14100_;
 wire _14101_;
 wire _14102_;
 wire _14103_;
 wire _14104_;
 wire _14105_;
 wire _14106_;
 wire _14107_;
 wire _14108_;
 wire _14109_;
 wire _14110_;
 wire _14111_;
 wire _14112_;
 wire _14113_;
 wire _14114_;
 wire _14115_;
 wire _14116_;
 wire _14117_;
 wire _14118_;
 wire _14119_;
 wire _14120_;
 wire _14121_;
 wire _14122_;
 wire _14123_;
 wire _14124_;
 wire _14125_;
 wire _14126_;
 wire _14127_;
 wire _14128_;
 wire _14129_;
 wire _14130_;
 wire _14131_;
 wire _14132_;
 wire _14133_;
 wire _14134_;
 wire _14135_;
 wire _14136_;
 wire _14137_;
 wire _14138_;
 wire _14139_;
 wire _14140_;
 wire _14141_;
 wire _14142_;
 wire _14143_;
 wire _14144_;
 wire _14145_;
 wire _14146_;
 wire _14147_;
 wire _14148_;
 wire _14149_;
 wire _14150_;
 wire _14151_;
 wire _14152_;
 wire _14153_;
 wire _14154_;
 wire _14155_;
 wire _14156_;
 wire _14157_;
 wire _14158_;
 wire _14159_;
 wire _14160_;
 wire _14161_;
 wire _14162_;
 wire _14163_;
 wire _14164_;
 wire _14165_;
 wire _14166_;
 wire _14167_;
 wire _14168_;
 wire _14169_;
 wire _14170_;
 wire _14171_;
 wire _14172_;
 wire _14173_;
 wire _14174_;
 wire _14175_;
 wire _14176_;
 wire _14177_;
 wire _14178_;
 wire _14179_;
 wire _14180_;
 wire _14181_;
 wire _14182_;
 wire _14183_;
 wire _14184_;
 wire _14185_;
 wire _14186_;
 wire _14187_;
 wire _14188_;
 wire _14189_;
 wire _14190_;
 wire _14191_;
 wire _14192_;
 wire _14193_;
 wire _14194_;
 wire _14195_;
 wire _14196_;
 wire _14197_;
 wire _14198_;
 wire _14199_;
 wire _14200_;
 wire _14201_;
 wire _14202_;
 wire _14203_;
 wire _14204_;
 wire _14205_;
 wire _14206_;
 wire _14207_;
 wire _14208_;
 wire _14209_;
 wire _14210_;
 wire _14211_;
 wire _14212_;
 wire _14213_;
 wire _14214_;
 wire _14215_;
 wire _14216_;
 wire _14217_;
 wire _14218_;
 wire _14219_;
 wire _14220_;
 wire _14221_;
 wire _14222_;
 wire _14223_;
 wire _14224_;
 wire _14225_;
 wire _14226_;
 wire _14227_;
 wire _14228_;
 wire _14229_;
 wire _14230_;
 wire _14231_;
 wire _14232_;
 wire _14233_;
 wire _14234_;
 wire _14235_;
 wire _14236_;
 wire _14237_;
 wire _14238_;
 wire _14239_;
 wire _14240_;
 wire _14241_;
 wire _14242_;
 wire _14243_;
 wire _14244_;
 wire _14245_;
 wire _14246_;
 wire _14247_;
 wire _14248_;
 wire _14249_;
 wire _14250_;
 wire _14251_;
 wire _14252_;
 wire _14253_;
 wire _14254_;
 wire _14255_;
 wire _14256_;
 wire _14257_;
 wire _14258_;
 wire _14259_;
 wire _14260_;
 wire _14261_;
 wire _14262_;
 wire _14263_;
 wire _14264_;
 wire _14265_;
 wire _14266_;
 wire _14267_;
 wire _14268_;
 wire _14269_;
 wire _14270_;
 wire _14271_;
 wire _14272_;
 wire _14273_;
 wire _14274_;
 wire _14275_;
 wire _14276_;
 wire _14277_;
 wire _14278_;
 wire _14279_;
 wire _14280_;
 wire _14281_;
 wire _14282_;
 wire _14283_;
 wire _14284_;
 wire _14285_;
 wire _14286_;
 wire _14287_;
 wire _14288_;
 wire _14289_;
 wire _14290_;
 wire _14291_;
 wire _14292_;
 wire _14293_;
 wire _14294_;
 wire _14295_;
 wire _14296_;
 wire _14297_;
 wire _14298_;
 wire _14299_;
 wire _14300_;
 wire _14301_;
 wire _14302_;
 wire _14303_;
 wire _14304_;
 wire _14305_;
 wire _14306_;
 wire _14307_;
 wire _14308_;
 wire _14309_;
 wire _14310_;
 wire _14311_;
 wire _14312_;
 wire _14313_;
 wire _14314_;
 wire _14315_;
 wire _14316_;
 wire _14317_;
 wire _14318_;
 wire _14319_;
 wire _14320_;
 wire _14321_;
 wire _14322_;
 wire _14323_;
 wire _14324_;
 wire _14325_;
 wire _14326_;
 wire _14327_;
 wire _14328_;
 wire _14329_;
 wire _14330_;
 wire _14331_;
 wire _14332_;
 wire _14333_;
 wire _14334_;
 wire _14335_;
 wire _14336_;
 wire _14337_;
 wire _14338_;
 wire _14339_;
 wire _14340_;
 wire _14341_;
 wire _14342_;
 wire _14343_;
 wire _14344_;
 wire _14345_;
 wire _14346_;
 wire _14347_;
 wire _14348_;
 wire _14349_;
 wire _14350_;
 wire _14351_;
 wire _14352_;
 wire _14353_;
 wire _14354_;
 wire _14355_;
 wire _14356_;
 wire _14357_;
 wire _14358_;
 wire _14359_;
 wire _14360_;
 wire _14361_;
 wire _14362_;
 wire _14363_;
 wire _14364_;
 wire _14365_;
 wire _14366_;
 wire _14367_;
 wire _14368_;
 wire _14369_;
 wire _14370_;
 wire _14371_;
 wire _14372_;
 wire _14373_;
 wire _14374_;
 wire _14375_;
 wire _14376_;
 wire _14377_;
 wire _14378_;
 wire _14379_;
 wire _14380_;
 wire _14381_;
 wire _14382_;
 wire _14383_;
 wire _14384_;
 wire _14385_;
 wire _14386_;
 wire _14387_;
 wire _14388_;
 wire _14389_;
 wire _14390_;
 wire _14391_;
 wire _14392_;
 wire _14393_;
 wire _14394_;
 wire _14395_;
 wire _14396_;
 wire _14397_;
 wire _14398_;
 wire _14399_;
 wire _14400_;
 wire _14401_;
 wire _14402_;
 wire _14403_;
 wire _14404_;
 wire _14405_;
 wire _14406_;
 wire _14407_;
 wire _14408_;
 wire _14409_;
 wire _14410_;
 wire _14411_;
 wire _14412_;
 wire _14413_;
 wire _14414_;
 wire _14415_;
 wire _14416_;
 wire _14417_;
 wire _14418_;
 wire _14419_;
 wire _14420_;
 wire _14421_;
 wire _14422_;
 wire _14423_;
 wire _14424_;
 wire _14425_;
 wire _14426_;
 wire _14427_;
 wire _14428_;
 wire _14429_;
 wire _14430_;
 wire _14431_;
 wire _14432_;
 wire _14433_;
 wire _14434_;
 wire _14435_;
 wire _14436_;
 wire _14437_;
 wire _14438_;
 wire _14439_;
 wire _14440_;
 wire _14441_;
 wire _14442_;
 wire _14443_;
 wire _14444_;
 wire _14445_;
 wire _14446_;
 wire _14447_;
 wire _14448_;
 wire _14449_;
 wire _14450_;
 wire _14451_;
 wire _14452_;
 wire _14453_;
 wire _14454_;
 wire _14455_;
 wire _14456_;
 wire _14457_;
 wire _14458_;
 wire _14459_;
 wire _14460_;
 wire _14461_;
 wire _14462_;
 wire _14463_;
 wire _14464_;
 wire _14465_;
 wire _14466_;
 wire _14467_;
 wire _14468_;
 wire _14469_;
 wire _14470_;
 wire _14471_;
 wire _14472_;
 wire _14473_;
 wire _14474_;
 wire _14475_;
 wire _14476_;
 wire _14477_;
 wire _14478_;
 wire _14479_;
 wire _14480_;
 wire _14481_;
 wire _14482_;
 wire _14483_;
 wire _14484_;
 wire _14485_;
 wire _14486_;
 wire _14487_;
 wire _14488_;
 wire _14489_;
 wire _14490_;
 wire _14491_;
 wire _14492_;
 wire _14493_;
 wire _14494_;
 wire _14495_;
 wire _14496_;
 wire _14497_;
 wire _14498_;
 wire _14499_;
 wire _14500_;
 wire _14501_;
 wire _14502_;
 wire _14503_;
 wire _14504_;
 wire _14505_;
 wire _14506_;
 wire _14507_;
 wire _14508_;
 wire _14509_;
 wire _14510_;
 wire _14511_;
 wire _14512_;
 wire _14513_;
 wire _14514_;
 wire _14515_;
 wire _14516_;
 wire _14517_;
 wire _14518_;
 wire _14519_;
 wire _14520_;
 wire _14521_;
 wire _14522_;
 wire _14523_;
 wire _14524_;
 wire _14525_;
 wire _14526_;
 wire _14527_;
 wire _14528_;
 wire _14529_;
 wire _14530_;
 wire _14531_;
 wire _14532_;
 wire _14533_;
 wire _14534_;
 wire _14535_;
 wire _14536_;
 wire _14537_;
 wire _14538_;
 wire _14539_;
 wire _14540_;
 wire _14541_;
 wire _14542_;
 wire _14543_;
 wire _14544_;
 wire _14545_;
 wire _14546_;
 wire _14547_;
 wire _14548_;
 wire _14549_;
 wire _14550_;
 wire _14551_;
 wire _14552_;
 wire _14553_;
 wire _14554_;
 wire _14555_;
 wire _14556_;
 wire _14557_;
 wire _14558_;
 wire _14559_;
 wire _14560_;
 wire _14561_;
 wire _14562_;
 wire _14563_;
 wire _14564_;
 wire _14565_;
 wire _14566_;
 wire _14567_;
 wire _14568_;
 wire _14569_;
 wire _14570_;
 wire _14571_;
 wire _14572_;
 wire _14573_;
 wire _14574_;
 wire _14575_;
 wire _14576_;
 wire _14577_;
 wire _14578_;
 wire _14579_;
 wire _14580_;
 wire _14581_;
 wire _14582_;
 wire _14583_;
 wire _14584_;
 wire _14585_;
 wire _14586_;
 wire _14587_;
 wire _14588_;
 wire _14589_;
 wire _14590_;
 wire _14591_;
 wire _14592_;
 wire _14593_;
 wire _14594_;
 wire _14595_;
 wire _14596_;
 wire _14597_;
 wire _14598_;
 wire _14599_;
 wire _14600_;
 wire _14601_;
 wire _14602_;
 wire _14603_;
 wire _14604_;
 wire _14605_;
 wire _14606_;
 wire _14607_;
 wire _14608_;
 wire _14609_;
 wire _14610_;
 wire _14611_;
 wire _14612_;
 wire _14613_;
 wire _14614_;
 wire _14615_;
 wire _14616_;
 wire _14617_;
 wire _14618_;
 wire _14619_;
 wire _14620_;
 wire _14621_;
 wire _14622_;
 wire _14623_;
 wire _14624_;
 wire _14625_;
 wire _14626_;
 wire _14627_;
 wire _14628_;
 wire _14629_;
 wire _14630_;
 wire _14631_;
 wire _14632_;
 wire _14633_;
 wire _14634_;
 wire _14635_;
 wire _14636_;
 wire _14637_;
 wire _14638_;
 wire _14639_;
 wire _14640_;
 wire _14641_;
 wire _14642_;
 wire _14643_;
 wire _14644_;
 wire _14645_;
 wire _14646_;
 wire _14647_;
 wire _14648_;
 wire _14649_;
 wire _14650_;
 wire _14651_;
 wire _14652_;
 wire _14653_;
 wire _14654_;
 wire _14655_;
 wire _14656_;
 wire _14657_;
 wire _14658_;
 wire _14659_;
 wire _14660_;
 wire _14661_;
 wire _14662_;
 wire _14663_;
 wire _14664_;
 wire _14665_;
 wire _14666_;
 wire _14667_;
 wire _14668_;
 wire _14669_;
 wire _14670_;
 wire _14671_;
 wire _14672_;
 wire _14673_;
 wire _14674_;
 wire _14675_;
 wire _14676_;
 wire _14677_;
 wire _14678_;
 wire _14679_;
 wire _14680_;
 wire _14681_;
 wire _14682_;
 wire _14683_;
 wire _14684_;
 wire _14685_;
 wire _14686_;
 wire _14687_;
 wire _14688_;
 wire _14689_;
 wire _14690_;
 wire _14691_;
 wire _14692_;
 wire _14693_;
 wire _14694_;
 wire _14695_;
 wire _14696_;
 wire _14697_;
 wire _14698_;
 wire _14699_;
 wire _14700_;
 wire _14701_;
 wire _14702_;
 wire _14703_;
 wire _14704_;
 wire _14705_;
 wire _14706_;
 wire _14707_;
 wire _14708_;
 wire _14709_;
 wire _14710_;
 wire _14711_;
 wire _14712_;
 wire _14713_;
 wire _14714_;
 wire _14715_;
 wire _14716_;
 wire _14717_;
 wire _14718_;
 wire _14719_;
 wire _14720_;
 wire _14721_;
 wire _14722_;
 wire _14723_;
 wire _14724_;
 wire _14725_;
 wire _14726_;
 wire _14727_;
 wire _14728_;
 wire _14729_;
 wire _14730_;
 wire _14731_;
 wire _14732_;
 wire _14733_;
 wire _14734_;
 wire _14735_;
 wire _14736_;
 wire _14737_;
 wire _14738_;
 wire _14739_;
 wire _14740_;
 wire _14741_;
 wire _14742_;
 wire _14743_;
 wire _14744_;
 wire _14745_;
 wire _14746_;
 wire _14747_;
 wire _14748_;
 wire _14749_;
 wire _14750_;
 wire _14751_;
 wire _14752_;
 wire _14753_;
 wire _14754_;
 wire _14755_;
 wire _14756_;
 wire _14757_;
 wire _14758_;
 wire _14759_;
 wire _14760_;
 wire _14761_;
 wire _14762_;
 wire _14763_;
 wire _14764_;
 wire _14765_;
 wire _14766_;
 wire _14767_;
 wire _14768_;
 wire _14769_;
 wire _14770_;
 wire _14771_;
 wire _14772_;
 wire _14773_;
 wire _14774_;
 wire _14775_;
 wire _14776_;
 wire _14777_;
 wire _14778_;
 wire _14779_;
 wire _14780_;
 wire _14781_;
 wire _14782_;
 wire _14783_;
 wire _14784_;
 wire _14785_;
 wire _14786_;
 wire _14787_;
 wire _14788_;
 wire _14789_;
 wire _14790_;
 wire _14791_;
 wire _14792_;
 wire _14793_;
 wire _14794_;
 wire _14795_;
 wire _14796_;
 wire _14797_;
 wire _14798_;
 wire _14799_;
 wire _14800_;
 wire _14801_;
 wire _14802_;
 wire _14803_;
 wire _14804_;
 wire _14805_;
 wire _14806_;
 wire _14807_;
 wire _14808_;
 wire _14809_;
 wire _14810_;
 wire _14811_;
 wire _14812_;
 wire _14813_;
 wire _14814_;
 wire _14815_;
 wire _14816_;
 wire _14817_;
 wire _14818_;
 wire _14819_;
 wire _14820_;
 wire _14821_;
 wire _14822_;
 wire _14823_;
 wire _14824_;
 wire _14825_;
 wire _14826_;
 wire _14827_;
 wire _14828_;
 wire _14829_;
 wire _14830_;
 wire _14831_;
 wire _14832_;
 wire _14833_;
 wire _14834_;
 wire _14835_;
 wire _14836_;
 wire _14837_;
 wire _14838_;
 wire _14839_;
 wire _14840_;
 wire _14841_;
 wire _14842_;
 wire _14843_;
 wire _14844_;
 wire _14845_;
 wire _14846_;
 wire _14847_;
 wire _14848_;
 wire _14849_;
 wire _14850_;
 wire _14851_;
 wire _14852_;
 wire _14853_;
 wire _14854_;
 wire _14855_;
 wire _14856_;
 wire _14857_;
 wire _14858_;
 wire _14859_;
 wire _14860_;
 wire _14861_;
 wire _14862_;
 wire _14863_;
 wire _14864_;
 wire _14865_;
 wire _14866_;
 wire _14867_;
 wire _14868_;
 wire _14869_;
 wire _14870_;
 wire _14871_;
 wire _14872_;
 wire _14873_;
 wire _14874_;
 wire _14875_;
 wire _14876_;
 wire _14877_;
 wire _14878_;
 wire _14879_;
 wire _14880_;
 wire _14881_;
 wire _14882_;
 wire _14883_;
 wire _14884_;
 wire _14885_;
 wire _14886_;
 wire _14887_;
 wire _14888_;
 wire _14889_;
 wire _14890_;
 wire _14891_;
 wire _14892_;
 wire _14893_;
 wire _14894_;
 wire _14895_;
 wire _14896_;
 wire _14897_;
 wire _14898_;
 wire _14899_;
 wire _14900_;
 wire _14901_;
 wire _14902_;
 wire _14903_;
 wire _14904_;
 wire _14905_;
 wire _14906_;
 wire _14907_;
 wire _14908_;
 wire _14909_;
 wire _14910_;
 wire _14911_;
 wire _14912_;
 wire _14913_;
 wire _14914_;
 wire _14915_;
 wire _14916_;
 wire _14917_;
 wire _14918_;
 wire _14919_;
 wire _14920_;
 wire _14921_;
 wire _14922_;
 wire _14923_;
 wire _14924_;
 wire _14925_;
 wire _14926_;
 wire _14927_;
 wire _14928_;
 wire _14929_;
 wire _14930_;
 wire _14931_;
 wire _14932_;
 wire _14933_;
 wire _14934_;
 wire _14935_;
 wire _14936_;
 wire _14937_;
 wire _14938_;
 wire _14939_;
 wire _14940_;
 wire _14941_;
 wire _14942_;
 wire _14943_;
 wire _14944_;
 wire _14945_;
 wire _14946_;
 wire _14947_;
 wire _14948_;
 wire _14949_;
 wire _14950_;
 wire _14951_;
 wire _14952_;
 wire _14953_;
 wire _14954_;
 wire _14955_;
 wire _14956_;
 wire _14957_;
 wire _14958_;
 wire _14959_;
 wire _14960_;
 wire _14961_;
 wire _14962_;
 wire _14963_;
 wire _14964_;
 wire _14965_;
 wire _14966_;
 wire _14967_;
 wire _14968_;
 wire _14969_;
 wire _14970_;
 wire _14971_;
 wire _14972_;
 wire _14973_;
 wire _14974_;
 wire _14975_;
 wire _14976_;
 wire _14977_;
 wire _14978_;
 wire _14979_;
 wire _14980_;
 wire _14981_;
 wire _14982_;
 wire _14983_;
 wire _14984_;
 wire _14985_;
 wire _14986_;
 wire _14987_;
 wire _14988_;
 wire _14989_;
 wire _14990_;
 wire _14991_;
 wire _14992_;
 wire _14993_;
 wire _14994_;
 wire _14995_;
 wire _14996_;
 wire _14997_;
 wire _14998_;
 wire _14999_;
 wire _15000_;
 wire _15001_;
 wire _15002_;
 wire _15003_;
 wire _15004_;
 wire _15005_;
 wire _15006_;
 wire _15007_;
 wire _15008_;
 wire _15009_;
 wire _15010_;
 wire _15011_;
 wire _15012_;
 wire _15013_;
 wire _15014_;
 wire _15015_;
 wire _15016_;
 wire _15017_;
 wire _15018_;
 wire _15019_;
 wire _15020_;
 wire _15021_;
 wire _15022_;
 wire _15023_;
 wire _15024_;
 wire _15025_;
 wire _15026_;
 wire _15027_;
 wire _15028_;
 wire _15029_;
 wire _15030_;
 wire _15031_;
 wire _15032_;
 wire _15033_;
 wire _15034_;
 wire _15035_;
 wire _15036_;
 wire _15037_;
 wire _15038_;
 wire _15039_;
 wire _15040_;
 wire _15041_;
 wire _15042_;
 wire _15043_;
 wire _15044_;
 wire _15045_;
 wire _15046_;
 wire _15047_;
 wire _15048_;
 wire _15049_;
 wire _15050_;
 wire _15051_;
 wire _15052_;
 wire _15053_;
 wire _15054_;
 wire _15055_;
 wire _15056_;
 wire _15057_;
 wire _15058_;
 wire _15059_;
 wire _15060_;
 wire _15061_;
 wire _15062_;
 wire _15063_;
 wire _15064_;
 wire _15065_;
 wire _15066_;
 wire _15067_;
 wire _15068_;
 wire _15069_;
 wire _15070_;
 wire _15071_;
 wire _15072_;
 wire _15073_;
 wire _15074_;
 wire _15075_;
 wire _15076_;
 wire _15077_;
 wire _15078_;
 wire _15079_;
 wire _15080_;
 wire _15081_;
 wire _15082_;
 wire clknet_leaf_0_clk;
 wire \cpu.addr[10] ;
 wire \cpu.addr[11] ;
 wire \cpu.addr[12] ;
 wire \cpu.addr[13] ;
 wire \cpu.addr[14] ;
 wire \cpu.addr[15] ;
 wire \cpu.addr[1] ;
 wire \cpu.addr[2] ;
 wire \cpu.addr[3] ;
 wire \cpu.addr[4] ;
 wire \cpu.addr[5] ;
 wire \cpu.addr[6] ;
 wire \cpu.addr[7] ;
 wire \cpu.addr[8] ;
 wire \cpu.addr[9] ;
 wire \cpu.br ;
 wire \cpu.cond[0] ;
 wire \cpu.cond[1] ;
 wire \cpu.cond[2] ;
 wire \cpu.d_flush_all ;
 wire \cpu.d_rstrobe_d ;
 wire \cpu.d_wstrobe_d ;
 wire \cpu.dcache.flush_write ;
 wire \cpu.dcache.r_data[0][0] ;
 wire \cpu.dcache.r_data[0][10] ;
 wire \cpu.dcache.r_data[0][11] ;
 wire \cpu.dcache.r_data[0][12] ;
 wire \cpu.dcache.r_data[0][13] ;
 wire \cpu.dcache.r_data[0][14] ;
 wire \cpu.dcache.r_data[0][15] ;
 wire \cpu.dcache.r_data[0][16] ;
 wire \cpu.dcache.r_data[0][17] ;
 wire \cpu.dcache.r_data[0][18] ;
 wire \cpu.dcache.r_data[0][19] ;
 wire \cpu.dcache.r_data[0][1] ;
 wire \cpu.dcache.r_data[0][20] ;
 wire \cpu.dcache.r_data[0][21] ;
 wire \cpu.dcache.r_data[0][22] ;
 wire \cpu.dcache.r_data[0][23] ;
 wire \cpu.dcache.r_data[0][24] ;
 wire \cpu.dcache.r_data[0][25] ;
 wire \cpu.dcache.r_data[0][26] ;
 wire \cpu.dcache.r_data[0][27] ;
 wire \cpu.dcache.r_data[0][28] ;
 wire \cpu.dcache.r_data[0][29] ;
 wire \cpu.dcache.r_data[0][2] ;
 wire \cpu.dcache.r_data[0][30] ;
 wire \cpu.dcache.r_data[0][31] ;
 wire \cpu.dcache.r_data[0][3] ;
 wire \cpu.dcache.r_data[0][4] ;
 wire \cpu.dcache.r_data[0][5] ;
 wire \cpu.dcache.r_data[0][6] ;
 wire \cpu.dcache.r_data[0][7] ;
 wire \cpu.dcache.r_data[0][8] ;
 wire \cpu.dcache.r_data[0][9] ;
 wire \cpu.dcache.r_data[1][0] ;
 wire \cpu.dcache.r_data[1][10] ;
 wire \cpu.dcache.r_data[1][11] ;
 wire \cpu.dcache.r_data[1][12] ;
 wire \cpu.dcache.r_data[1][13] ;
 wire \cpu.dcache.r_data[1][14] ;
 wire \cpu.dcache.r_data[1][15] ;
 wire \cpu.dcache.r_data[1][16] ;
 wire \cpu.dcache.r_data[1][17] ;
 wire \cpu.dcache.r_data[1][18] ;
 wire \cpu.dcache.r_data[1][19] ;
 wire \cpu.dcache.r_data[1][1] ;
 wire \cpu.dcache.r_data[1][20] ;
 wire \cpu.dcache.r_data[1][21] ;
 wire \cpu.dcache.r_data[1][22] ;
 wire \cpu.dcache.r_data[1][23] ;
 wire \cpu.dcache.r_data[1][24] ;
 wire \cpu.dcache.r_data[1][25] ;
 wire \cpu.dcache.r_data[1][26] ;
 wire \cpu.dcache.r_data[1][27] ;
 wire \cpu.dcache.r_data[1][28] ;
 wire \cpu.dcache.r_data[1][29] ;
 wire \cpu.dcache.r_data[1][2] ;
 wire \cpu.dcache.r_data[1][30] ;
 wire \cpu.dcache.r_data[1][31] ;
 wire \cpu.dcache.r_data[1][3] ;
 wire \cpu.dcache.r_data[1][4] ;
 wire \cpu.dcache.r_data[1][5] ;
 wire \cpu.dcache.r_data[1][6] ;
 wire \cpu.dcache.r_data[1][7] ;
 wire \cpu.dcache.r_data[1][8] ;
 wire \cpu.dcache.r_data[1][9] ;
 wire \cpu.dcache.r_data[2][0] ;
 wire \cpu.dcache.r_data[2][10] ;
 wire \cpu.dcache.r_data[2][11] ;
 wire \cpu.dcache.r_data[2][12] ;
 wire \cpu.dcache.r_data[2][13] ;
 wire \cpu.dcache.r_data[2][14] ;
 wire \cpu.dcache.r_data[2][15] ;
 wire \cpu.dcache.r_data[2][16] ;
 wire \cpu.dcache.r_data[2][17] ;
 wire \cpu.dcache.r_data[2][18] ;
 wire \cpu.dcache.r_data[2][19] ;
 wire \cpu.dcache.r_data[2][1] ;
 wire \cpu.dcache.r_data[2][20] ;
 wire \cpu.dcache.r_data[2][21] ;
 wire \cpu.dcache.r_data[2][22] ;
 wire \cpu.dcache.r_data[2][23] ;
 wire \cpu.dcache.r_data[2][24] ;
 wire \cpu.dcache.r_data[2][25] ;
 wire \cpu.dcache.r_data[2][26] ;
 wire \cpu.dcache.r_data[2][27] ;
 wire \cpu.dcache.r_data[2][28] ;
 wire \cpu.dcache.r_data[2][29] ;
 wire \cpu.dcache.r_data[2][2] ;
 wire \cpu.dcache.r_data[2][30] ;
 wire \cpu.dcache.r_data[2][31] ;
 wire \cpu.dcache.r_data[2][3] ;
 wire \cpu.dcache.r_data[2][4] ;
 wire \cpu.dcache.r_data[2][5] ;
 wire \cpu.dcache.r_data[2][6] ;
 wire \cpu.dcache.r_data[2][7] ;
 wire \cpu.dcache.r_data[2][8] ;
 wire \cpu.dcache.r_data[2][9] ;
 wire \cpu.dcache.r_data[3][0] ;
 wire \cpu.dcache.r_data[3][10] ;
 wire \cpu.dcache.r_data[3][11] ;
 wire \cpu.dcache.r_data[3][12] ;
 wire \cpu.dcache.r_data[3][13] ;
 wire \cpu.dcache.r_data[3][14] ;
 wire \cpu.dcache.r_data[3][15] ;
 wire \cpu.dcache.r_data[3][16] ;
 wire \cpu.dcache.r_data[3][17] ;
 wire \cpu.dcache.r_data[3][18] ;
 wire \cpu.dcache.r_data[3][19] ;
 wire \cpu.dcache.r_data[3][1] ;
 wire \cpu.dcache.r_data[3][20] ;
 wire \cpu.dcache.r_data[3][21] ;
 wire \cpu.dcache.r_data[3][22] ;
 wire \cpu.dcache.r_data[3][23] ;
 wire \cpu.dcache.r_data[3][24] ;
 wire \cpu.dcache.r_data[3][25] ;
 wire \cpu.dcache.r_data[3][26] ;
 wire \cpu.dcache.r_data[3][27] ;
 wire \cpu.dcache.r_data[3][28] ;
 wire \cpu.dcache.r_data[3][29] ;
 wire \cpu.dcache.r_data[3][2] ;
 wire \cpu.dcache.r_data[3][30] ;
 wire \cpu.dcache.r_data[3][31] ;
 wire \cpu.dcache.r_data[3][3] ;
 wire \cpu.dcache.r_data[3][4] ;
 wire \cpu.dcache.r_data[3][5] ;
 wire \cpu.dcache.r_data[3][6] ;
 wire \cpu.dcache.r_data[3][7] ;
 wire \cpu.dcache.r_data[3][8] ;
 wire \cpu.dcache.r_data[3][9] ;
 wire \cpu.dcache.r_data[4][0] ;
 wire \cpu.dcache.r_data[4][10] ;
 wire \cpu.dcache.r_data[4][11] ;
 wire \cpu.dcache.r_data[4][12] ;
 wire \cpu.dcache.r_data[4][13] ;
 wire \cpu.dcache.r_data[4][14] ;
 wire \cpu.dcache.r_data[4][15] ;
 wire \cpu.dcache.r_data[4][16] ;
 wire \cpu.dcache.r_data[4][17] ;
 wire \cpu.dcache.r_data[4][18] ;
 wire \cpu.dcache.r_data[4][19] ;
 wire \cpu.dcache.r_data[4][1] ;
 wire \cpu.dcache.r_data[4][20] ;
 wire \cpu.dcache.r_data[4][21] ;
 wire \cpu.dcache.r_data[4][22] ;
 wire \cpu.dcache.r_data[4][23] ;
 wire \cpu.dcache.r_data[4][24] ;
 wire \cpu.dcache.r_data[4][25] ;
 wire \cpu.dcache.r_data[4][26] ;
 wire \cpu.dcache.r_data[4][27] ;
 wire \cpu.dcache.r_data[4][28] ;
 wire \cpu.dcache.r_data[4][29] ;
 wire \cpu.dcache.r_data[4][2] ;
 wire \cpu.dcache.r_data[4][30] ;
 wire \cpu.dcache.r_data[4][31] ;
 wire \cpu.dcache.r_data[4][3] ;
 wire \cpu.dcache.r_data[4][4] ;
 wire \cpu.dcache.r_data[4][5] ;
 wire \cpu.dcache.r_data[4][6] ;
 wire \cpu.dcache.r_data[4][7] ;
 wire \cpu.dcache.r_data[4][8] ;
 wire \cpu.dcache.r_data[4][9] ;
 wire \cpu.dcache.r_data[5][0] ;
 wire \cpu.dcache.r_data[5][10] ;
 wire \cpu.dcache.r_data[5][11] ;
 wire \cpu.dcache.r_data[5][12] ;
 wire \cpu.dcache.r_data[5][13] ;
 wire \cpu.dcache.r_data[5][14] ;
 wire \cpu.dcache.r_data[5][15] ;
 wire \cpu.dcache.r_data[5][16] ;
 wire \cpu.dcache.r_data[5][17] ;
 wire \cpu.dcache.r_data[5][18] ;
 wire \cpu.dcache.r_data[5][19] ;
 wire \cpu.dcache.r_data[5][1] ;
 wire \cpu.dcache.r_data[5][20] ;
 wire \cpu.dcache.r_data[5][21] ;
 wire \cpu.dcache.r_data[5][22] ;
 wire \cpu.dcache.r_data[5][23] ;
 wire \cpu.dcache.r_data[5][24] ;
 wire \cpu.dcache.r_data[5][25] ;
 wire \cpu.dcache.r_data[5][26] ;
 wire \cpu.dcache.r_data[5][27] ;
 wire \cpu.dcache.r_data[5][28] ;
 wire \cpu.dcache.r_data[5][29] ;
 wire \cpu.dcache.r_data[5][2] ;
 wire \cpu.dcache.r_data[5][30] ;
 wire \cpu.dcache.r_data[5][31] ;
 wire \cpu.dcache.r_data[5][3] ;
 wire \cpu.dcache.r_data[5][4] ;
 wire \cpu.dcache.r_data[5][5] ;
 wire \cpu.dcache.r_data[5][6] ;
 wire \cpu.dcache.r_data[5][7] ;
 wire \cpu.dcache.r_data[5][8] ;
 wire \cpu.dcache.r_data[5][9] ;
 wire \cpu.dcache.r_data[6][0] ;
 wire \cpu.dcache.r_data[6][10] ;
 wire \cpu.dcache.r_data[6][11] ;
 wire \cpu.dcache.r_data[6][12] ;
 wire \cpu.dcache.r_data[6][13] ;
 wire \cpu.dcache.r_data[6][14] ;
 wire \cpu.dcache.r_data[6][15] ;
 wire \cpu.dcache.r_data[6][16] ;
 wire \cpu.dcache.r_data[6][17] ;
 wire \cpu.dcache.r_data[6][18] ;
 wire \cpu.dcache.r_data[6][19] ;
 wire \cpu.dcache.r_data[6][1] ;
 wire \cpu.dcache.r_data[6][20] ;
 wire \cpu.dcache.r_data[6][21] ;
 wire \cpu.dcache.r_data[6][22] ;
 wire \cpu.dcache.r_data[6][23] ;
 wire \cpu.dcache.r_data[6][24] ;
 wire \cpu.dcache.r_data[6][25] ;
 wire \cpu.dcache.r_data[6][26] ;
 wire \cpu.dcache.r_data[6][27] ;
 wire \cpu.dcache.r_data[6][28] ;
 wire \cpu.dcache.r_data[6][29] ;
 wire \cpu.dcache.r_data[6][2] ;
 wire \cpu.dcache.r_data[6][30] ;
 wire \cpu.dcache.r_data[6][31] ;
 wire \cpu.dcache.r_data[6][3] ;
 wire \cpu.dcache.r_data[6][4] ;
 wire \cpu.dcache.r_data[6][5] ;
 wire \cpu.dcache.r_data[6][6] ;
 wire \cpu.dcache.r_data[6][7] ;
 wire \cpu.dcache.r_data[6][8] ;
 wire \cpu.dcache.r_data[6][9] ;
 wire \cpu.dcache.r_data[7][0] ;
 wire \cpu.dcache.r_data[7][10] ;
 wire \cpu.dcache.r_data[7][11] ;
 wire \cpu.dcache.r_data[7][12] ;
 wire \cpu.dcache.r_data[7][13] ;
 wire \cpu.dcache.r_data[7][14] ;
 wire \cpu.dcache.r_data[7][15] ;
 wire \cpu.dcache.r_data[7][16] ;
 wire \cpu.dcache.r_data[7][17] ;
 wire \cpu.dcache.r_data[7][18] ;
 wire \cpu.dcache.r_data[7][19] ;
 wire \cpu.dcache.r_data[7][1] ;
 wire \cpu.dcache.r_data[7][20] ;
 wire \cpu.dcache.r_data[7][21] ;
 wire \cpu.dcache.r_data[7][22] ;
 wire \cpu.dcache.r_data[7][23] ;
 wire \cpu.dcache.r_data[7][24] ;
 wire \cpu.dcache.r_data[7][25] ;
 wire \cpu.dcache.r_data[7][26] ;
 wire \cpu.dcache.r_data[7][27] ;
 wire \cpu.dcache.r_data[7][28] ;
 wire \cpu.dcache.r_data[7][29] ;
 wire \cpu.dcache.r_data[7][2] ;
 wire \cpu.dcache.r_data[7][30] ;
 wire \cpu.dcache.r_data[7][31] ;
 wire \cpu.dcache.r_data[7][3] ;
 wire \cpu.dcache.r_data[7][4] ;
 wire \cpu.dcache.r_data[7][5] ;
 wire \cpu.dcache.r_data[7][6] ;
 wire \cpu.dcache.r_data[7][7] ;
 wire \cpu.dcache.r_data[7][8] ;
 wire \cpu.dcache.r_data[7][9] ;
 wire \cpu.dcache.r_dirty[0] ;
 wire \cpu.dcache.r_dirty[1] ;
 wire \cpu.dcache.r_dirty[2] ;
 wire \cpu.dcache.r_dirty[3] ;
 wire \cpu.dcache.r_dirty[4] ;
 wire \cpu.dcache.r_dirty[5] ;
 wire \cpu.dcache.r_dirty[6] ;
 wire \cpu.dcache.r_dirty[7] ;
 wire \cpu.dcache.r_offset[0] ;
 wire \cpu.dcache.r_offset[1] ;
 wire \cpu.dcache.r_offset[2] ;
 wire \cpu.dcache.r_tag[0][10] ;
 wire \cpu.dcache.r_tag[0][11] ;
 wire \cpu.dcache.r_tag[0][12] ;
 wire \cpu.dcache.r_tag[0][13] ;
 wire \cpu.dcache.r_tag[0][14] ;
 wire \cpu.dcache.r_tag[0][15] ;
 wire \cpu.dcache.r_tag[0][16] ;
 wire \cpu.dcache.r_tag[0][17] ;
 wire \cpu.dcache.r_tag[0][18] ;
 wire \cpu.dcache.r_tag[0][19] ;
 wire \cpu.dcache.r_tag[0][20] ;
 wire \cpu.dcache.r_tag[0][21] ;
 wire \cpu.dcache.r_tag[0][22] ;
 wire \cpu.dcache.r_tag[0][23] ;
 wire \cpu.dcache.r_tag[0][5] ;
 wire \cpu.dcache.r_tag[0][6] ;
 wire \cpu.dcache.r_tag[0][7] ;
 wire \cpu.dcache.r_tag[0][8] ;
 wire \cpu.dcache.r_tag[0][9] ;
 wire \cpu.dcache.r_tag[1][10] ;
 wire \cpu.dcache.r_tag[1][11] ;
 wire \cpu.dcache.r_tag[1][12] ;
 wire \cpu.dcache.r_tag[1][13] ;
 wire \cpu.dcache.r_tag[1][14] ;
 wire \cpu.dcache.r_tag[1][15] ;
 wire \cpu.dcache.r_tag[1][16] ;
 wire \cpu.dcache.r_tag[1][17] ;
 wire \cpu.dcache.r_tag[1][18] ;
 wire \cpu.dcache.r_tag[1][19] ;
 wire \cpu.dcache.r_tag[1][20] ;
 wire \cpu.dcache.r_tag[1][21] ;
 wire \cpu.dcache.r_tag[1][22] ;
 wire \cpu.dcache.r_tag[1][23] ;
 wire \cpu.dcache.r_tag[1][5] ;
 wire \cpu.dcache.r_tag[1][6] ;
 wire \cpu.dcache.r_tag[1][7] ;
 wire \cpu.dcache.r_tag[1][8] ;
 wire \cpu.dcache.r_tag[1][9] ;
 wire \cpu.dcache.r_tag[2][10] ;
 wire \cpu.dcache.r_tag[2][11] ;
 wire \cpu.dcache.r_tag[2][12] ;
 wire \cpu.dcache.r_tag[2][13] ;
 wire \cpu.dcache.r_tag[2][14] ;
 wire \cpu.dcache.r_tag[2][15] ;
 wire \cpu.dcache.r_tag[2][16] ;
 wire \cpu.dcache.r_tag[2][17] ;
 wire \cpu.dcache.r_tag[2][18] ;
 wire \cpu.dcache.r_tag[2][19] ;
 wire \cpu.dcache.r_tag[2][20] ;
 wire \cpu.dcache.r_tag[2][21] ;
 wire \cpu.dcache.r_tag[2][22] ;
 wire \cpu.dcache.r_tag[2][23] ;
 wire \cpu.dcache.r_tag[2][5] ;
 wire \cpu.dcache.r_tag[2][6] ;
 wire \cpu.dcache.r_tag[2][7] ;
 wire \cpu.dcache.r_tag[2][8] ;
 wire \cpu.dcache.r_tag[2][9] ;
 wire \cpu.dcache.r_tag[3][10] ;
 wire \cpu.dcache.r_tag[3][11] ;
 wire \cpu.dcache.r_tag[3][12] ;
 wire \cpu.dcache.r_tag[3][13] ;
 wire \cpu.dcache.r_tag[3][14] ;
 wire \cpu.dcache.r_tag[3][15] ;
 wire \cpu.dcache.r_tag[3][16] ;
 wire \cpu.dcache.r_tag[3][17] ;
 wire \cpu.dcache.r_tag[3][18] ;
 wire \cpu.dcache.r_tag[3][19] ;
 wire \cpu.dcache.r_tag[3][20] ;
 wire \cpu.dcache.r_tag[3][21] ;
 wire \cpu.dcache.r_tag[3][22] ;
 wire \cpu.dcache.r_tag[3][23] ;
 wire \cpu.dcache.r_tag[3][5] ;
 wire \cpu.dcache.r_tag[3][6] ;
 wire \cpu.dcache.r_tag[3][7] ;
 wire \cpu.dcache.r_tag[3][8] ;
 wire \cpu.dcache.r_tag[3][9] ;
 wire \cpu.dcache.r_tag[4][10] ;
 wire \cpu.dcache.r_tag[4][11] ;
 wire \cpu.dcache.r_tag[4][12] ;
 wire \cpu.dcache.r_tag[4][13] ;
 wire \cpu.dcache.r_tag[4][14] ;
 wire \cpu.dcache.r_tag[4][15] ;
 wire \cpu.dcache.r_tag[4][16] ;
 wire \cpu.dcache.r_tag[4][17] ;
 wire \cpu.dcache.r_tag[4][18] ;
 wire \cpu.dcache.r_tag[4][19] ;
 wire \cpu.dcache.r_tag[4][20] ;
 wire \cpu.dcache.r_tag[4][21] ;
 wire \cpu.dcache.r_tag[4][22] ;
 wire \cpu.dcache.r_tag[4][23] ;
 wire \cpu.dcache.r_tag[4][5] ;
 wire \cpu.dcache.r_tag[4][6] ;
 wire \cpu.dcache.r_tag[4][7] ;
 wire \cpu.dcache.r_tag[4][8] ;
 wire \cpu.dcache.r_tag[4][9] ;
 wire \cpu.dcache.r_tag[5][10] ;
 wire \cpu.dcache.r_tag[5][11] ;
 wire \cpu.dcache.r_tag[5][12] ;
 wire \cpu.dcache.r_tag[5][13] ;
 wire \cpu.dcache.r_tag[5][14] ;
 wire \cpu.dcache.r_tag[5][15] ;
 wire \cpu.dcache.r_tag[5][16] ;
 wire \cpu.dcache.r_tag[5][17] ;
 wire \cpu.dcache.r_tag[5][18] ;
 wire \cpu.dcache.r_tag[5][19] ;
 wire \cpu.dcache.r_tag[5][20] ;
 wire \cpu.dcache.r_tag[5][21] ;
 wire \cpu.dcache.r_tag[5][22] ;
 wire \cpu.dcache.r_tag[5][23] ;
 wire \cpu.dcache.r_tag[5][5] ;
 wire \cpu.dcache.r_tag[5][6] ;
 wire \cpu.dcache.r_tag[5][7] ;
 wire \cpu.dcache.r_tag[5][8] ;
 wire \cpu.dcache.r_tag[5][9] ;
 wire \cpu.dcache.r_tag[6][10] ;
 wire \cpu.dcache.r_tag[6][11] ;
 wire \cpu.dcache.r_tag[6][12] ;
 wire \cpu.dcache.r_tag[6][13] ;
 wire \cpu.dcache.r_tag[6][14] ;
 wire \cpu.dcache.r_tag[6][15] ;
 wire \cpu.dcache.r_tag[6][16] ;
 wire \cpu.dcache.r_tag[6][17] ;
 wire \cpu.dcache.r_tag[6][18] ;
 wire \cpu.dcache.r_tag[6][19] ;
 wire \cpu.dcache.r_tag[6][20] ;
 wire \cpu.dcache.r_tag[6][21] ;
 wire \cpu.dcache.r_tag[6][22] ;
 wire \cpu.dcache.r_tag[6][23] ;
 wire \cpu.dcache.r_tag[6][5] ;
 wire \cpu.dcache.r_tag[6][6] ;
 wire \cpu.dcache.r_tag[6][7] ;
 wire \cpu.dcache.r_tag[6][8] ;
 wire \cpu.dcache.r_tag[6][9] ;
 wire \cpu.dcache.r_tag[7][10] ;
 wire \cpu.dcache.r_tag[7][11] ;
 wire \cpu.dcache.r_tag[7][12] ;
 wire \cpu.dcache.r_tag[7][13] ;
 wire \cpu.dcache.r_tag[7][14] ;
 wire \cpu.dcache.r_tag[7][15] ;
 wire \cpu.dcache.r_tag[7][16] ;
 wire \cpu.dcache.r_tag[7][17] ;
 wire \cpu.dcache.r_tag[7][18] ;
 wire \cpu.dcache.r_tag[7][19] ;
 wire \cpu.dcache.r_tag[7][20] ;
 wire \cpu.dcache.r_tag[7][21] ;
 wire \cpu.dcache.r_tag[7][22] ;
 wire \cpu.dcache.r_tag[7][23] ;
 wire \cpu.dcache.r_tag[7][5] ;
 wire \cpu.dcache.r_tag[7][6] ;
 wire \cpu.dcache.r_tag[7][7] ;
 wire \cpu.dcache.r_tag[7][8] ;
 wire \cpu.dcache.r_tag[7][9] ;
 wire \cpu.dcache.r_valid[0] ;
 wire \cpu.dcache.r_valid[1] ;
 wire \cpu.dcache.r_valid[2] ;
 wire \cpu.dcache.r_valid[3] ;
 wire \cpu.dcache.r_valid[4] ;
 wire \cpu.dcache.r_valid[5] ;
 wire \cpu.dcache.r_valid[6] ;
 wire \cpu.dcache.r_valid[7] ;
 wire \cpu.dcache.wdata[0] ;
 wire \cpu.dcache.wdata[10] ;
 wire \cpu.dcache.wdata[11] ;
 wire \cpu.dcache.wdata[12] ;
 wire \cpu.dcache.wdata[13] ;
 wire \cpu.dcache.wdata[14] ;
 wire \cpu.dcache.wdata[15] ;
 wire \cpu.dcache.wdata[1] ;
 wire \cpu.dcache.wdata[2] ;
 wire \cpu.dcache.wdata[3] ;
 wire \cpu.dcache.wdata[4] ;
 wire \cpu.dcache.wdata[5] ;
 wire \cpu.dcache.wdata[6] ;
 wire \cpu.dcache.wdata[7] ;
 wire \cpu.dcache.wdata[8] ;
 wire \cpu.dcache.wdata[9] ;
 wire \cpu.dec.div ;
 wire \cpu.dec.do_flush_all ;
 wire \cpu.dec.do_flush_write ;
 wire \cpu.dec.do_inv_mmu ;
 wire \cpu.dec.imm[0] ;
 wire \cpu.dec.imm[10] ;
 wire \cpu.dec.imm[11] ;
 wire \cpu.dec.imm[12] ;
 wire \cpu.dec.imm[13] ;
 wire \cpu.dec.imm[14] ;
 wire \cpu.dec.imm[15] ;
 wire \cpu.dec.imm[1] ;
 wire \cpu.dec.imm[2] ;
 wire \cpu.dec.imm[3] ;
 wire \cpu.dec.imm[4] ;
 wire \cpu.dec.imm[5] ;
 wire \cpu.dec.imm[6] ;
 wire \cpu.dec.imm[7] ;
 wire \cpu.dec.imm[8] ;
 wire \cpu.dec.imm[9] ;
 wire \cpu.dec.io ;
 wire \cpu.dec.iready ;
 wire \cpu.dec.jmp ;
 wire \cpu.dec.load ;
 wire \cpu.dec.mult ;
 wire \cpu.dec.needs_rs2 ;
 wire \cpu.dec.r_op[10] ;
 wire \cpu.dec.r_op[1] ;
 wire \cpu.dec.r_op[2] ;
 wire \cpu.dec.r_op[3] ;
 wire \cpu.dec.r_op[4] ;
 wire \cpu.dec.r_op[5] ;
 wire \cpu.dec.r_op[6] ;
 wire \cpu.dec.r_op[7] ;
 wire \cpu.dec.r_op[8] ;
 wire \cpu.dec.r_op[9] ;
 wire \cpu.dec.r_rd[0] ;
 wire \cpu.dec.r_rd[1] ;
 wire \cpu.dec.r_rd[2] ;
 wire \cpu.dec.r_rd[3] ;
 wire \cpu.dec.r_rs1[0] ;
 wire \cpu.dec.r_rs1[1] ;
 wire \cpu.dec.r_rs1[2] ;
 wire \cpu.dec.r_rs1[3] ;
 wire \cpu.dec.r_rs2[0] ;
 wire \cpu.dec.r_rs2[1] ;
 wire \cpu.dec.r_rs2[2] ;
 wire \cpu.dec.r_rs2[3] ;
 wire \cpu.dec.r_rs2_pc ;
 wire \cpu.dec.r_set_cc ;
 wire \cpu.dec.r_store ;
 wire \cpu.dec.r_swapsp ;
 wire \cpu.dec.r_sys_call ;
 wire \cpu.dec.r_trap ;
 wire \cpu.dec.supmode ;
 wire \cpu.dec.user_io ;
 wire \cpu.ex.c_div_running ;
 wire \cpu.ex.c_mult[0] ;
 wire \cpu.ex.c_mult[10] ;
 wire \cpu.ex.c_mult[11] ;
 wire \cpu.ex.c_mult[12] ;
 wire \cpu.ex.c_mult[13] ;
 wire \cpu.ex.c_mult[14] ;
 wire \cpu.ex.c_mult[15] ;
 wire \cpu.ex.c_mult[1] ;
 wire \cpu.ex.c_mult[2] ;
 wire \cpu.ex.c_mult[3] ;
 wire \cpu.ex.c_mult[4] ;
 wire \cpu.ex.c_mult[5] ;
 wire \cpu.ex.c_mult[6] ;
 wire \cpu.ex.c_mult[7] ;
 wire \cpu.ex.c_mult[8] ;
 wire \cpu.ex.c_mult[9] ;
 wire \cpu.ex.c_mult_off[0] ;
 wire \cpu.ex.c_mult_off[1] ;
 wire \cpu.ex.c_mult_off[2] ;
 wire \cpu.ex.c_mult_off[3] ;
 wire \cpu.ex.c_mult_running ;
 wire \cpu.ex.genblk3.c_supmode ;
 wire \cpu.ex.genblk3.r_mmu_d_proxy ;
 wire \cpu.ex.genblk3.r_mmu_enable ;
 wire \cpu.ex.genblk3.r_prev_supmode ;
 wire \cpu.ex.i_flush_all ;
 wire \cpu.ex.ifetch ;
 wire \cpu.ex.io_access ;
 wire \cpu.ex.mmu_read[12] ;
 wire \cpu.ex.mmu_read[13] ;
 wire \cpu.ex.mmu_read[14] ;
 wire \cpu.ex.mmu_read[15] ;
 wire \cpu.ex.mmu_read[1] ;
 wire \cpu.ex.mmu_read[2] ;
 wire \cpu.ex.mmu_read[3] ;
 wire \cpu.ex.mmu_reg_data[0] ;
 wire \cpu.ex.pc[10] ;
 wire \cpu.ex.pc[11] ;
 wire \cpu.ex.pc[12] ;
 wire \cpu.ex.pc[13] ;
 wire \cpu.ex.pc[14] ;
 wire \cpu.ex.pc[15] ;
 wire \cpu.ex.pc[1] ;
 wire \cpu.ex.pc[2] ;
 wire \cpu.ex.pc[3] ;
 wire \cpu.ex.pc[4] ;
 wire \cpu.ex.pc[5] ;
 wire \cpu.ex.pc[6] ;
 wire \cpu.ex.pc[7] ;
 wire \cpu.ex.pc[8] ;
 wire \cpu.ex.pc[9] ;
 wire \cpu.ex.r_10[0] ;
 wire \cpu.ex.r_10[10] ;
 wire \cpu.ex.r_10[11] ;
 wire \cpu.ex.r_10[12] ;
 wire \cpu.ex.r_10[13] ;
 wire \cpu.ex.r_10[14] ;
 wire \cpu.ex.r_10[15] ;
 wire \cpu.ex.r_10[1] ;
 wire \cpu.ex.r_10[2] ;
 wire \cpu.ex.r_10[3] ;
 wire \cpu.ex.r_10[4] ;
 wire \cpu.ex.r_10[5] ;
 wire \cpu.ex.r_10[6] ;
 wire \cpu.ex.r_10[7] ;
 wire \cpu.ex.r_10[8] ;
 wire \cpu.ex.r_10[9] ;
 wire \cpu.ex.r_11[0] ;
 wire \cpu.ex.r_11[10] ;
 wire \cpu.ex.r_11[11] ;
 wire \cpu.ex.r_11[12] ;
 wire \cpu.ex.r_11[13] ;
 wire \cpu.ex.r_11[14] ;
 wire \cpu.ex.r_11[15] ;
 wire \cpu.ex.r_11[1] ;
 wire \cpu.ex.r_11[2] ;
 wire \cpu.ex.r_11[3] ;
 wire \cpu.ex.r_11[4] ;
 wire \cpu.ex.r_11[5] ;
 wire \cpu.ex.r_11[6] ;
 wire \cpu.ex.r_11[7] ;
 wire \cpu.ex.r_11[8] ;
 wire \cpu.ex.r_11[9] ;
 wire \cpu.ex.r_12[0] ;
 wire \cpu.ex.r_12[10] ;
 wire \cpu.ex.r_12[11] ;
 wire \cpu.ex.r_12[12] ;
 wire \cpu.ex.r_12[13] ;
 wire \cpu.ex.r_12[14] ;
 wire \cpu.ex.r_12[15] ;
 wire \cpu.ex.r_12[1] ;
 wire \cpu.ex.r_12[2] ;
 wire \cpu.ex.r_12[3] ;
 wire \cpu.ex.r_12[4] ;
 wire \cpu.ex.r_12[5] ;
 wire \cpu.ex.r_12[6] ;
 wire \cpu.ex.r_12[7] ;
 wire \cpu.ex.r_12[8] ;
 wire \cpu.ex.r_12[9] ;
 wire \cpu.ex.r_13[0] ;
 wire \cpu.ex.r_13[10] ;
 wire \cpu.ex.r_13[11] ;
 wire \cpu.ex.r_13[12] ;
 wire \cpu.ex.r_13[13] ;
 wire \cpu.ex.r_13[14] ;
 wire \cpu.ex.r_13[15] ;
 wire \cpu.ex.r_13[1] ;
 wire \cpu.ex.r_13[2] ;
 wire \cpu.ex.r_13[3] ;
 wire \cpu.ex.r_13[4] ;
 wire \cpu.ex.r_13[5] ;
 wire \cpu.ex.r_13[6] ;
 wire \cpu.ex.r_13[7] ;
 wire \cpu.ex.r_13[8] ;
 wire \cpu.ex.r_13[9] ;
 wire \cpu.ex.r_14[0] ;
 wire \cpu.ex.r_14[10] ;
 wire \cpu.ex.r_14[11] ;
 wire \cpu.ex.r_14[12] ;
 wire \cpu.ex.r_14[13] ;
 wire \cpu.ex.r_14[14] ;
 wire \cpu.ex.r_14[15] ;
 wire \cpu.ex.r_14[1] ;
 wire \cpu.ex.r_14[2] ;
 wire \cpu.ex.r_14[3] ;
 wire \cpu.ex.r_14[4] ;
 wire \cpu.ex.r_14[5] ;
 wire \cpu.ex.r_14[6] ;
 wire \cpu.ex.r_14[7] ;
 wire \cpu.ex.r_14[8] ;
 wire \cpu.ex.r_14[9] ;
 wire \cpu.ex.r_15[0] ;
 wire \cpu.ex.r_15[10] ;
 wire \cpu.ex.r_15[11] ;
 wire \cpu.ex.r_15[12] ;
 wire \cpu.ex.r_15[13] ;
 wire \cpu.ex.r_15[14] ;
 wire \cpu.ex.r_15[15] ;
 wire \cpu.ex.r_15[1] ;
 wire \cpu.ex.r_15[2] ;
 wire \cpu.ex.r_15[3] ;
 wire \cpu.ex.r_15[4] ;
 wire \cpu.ex.r_15[5] ;
 wire \cpu.ex.r_15[6] ;
 wire \cpu.ex.r_15[7] ;
 wire \cpu.ex.r_15[8] ;
 wire \cpu.ex.r_15[9] ;
 wire \cpu.ex.r_8[0] ;
 wire \cpu.ex.r_8[10] ;
 wire \cpu.ex.r_8[11] ;
 wire \cpu.ex.r_8[12] ;
 wire \cpu.ex.r_8[13] ;
 wire \cpu.ex.r_8[14] ;
 wire \cpu.ex.r_8[15] ;
 wire \cpu.ex.r_8[1] ;
 wire \cpu.ex.r_8[2] ;
 wire \cpu.ex.r_8[3] ;
 wire \cpu.ex.r_8[4] ;
 wire \cpu.ex.r_8[5] ;
 wire \cpu.ex.r_8[6] ;
 wire \cpu.ex.r_8[7] ;
 wire \cpu.ex.r_8[8] ;
 wire \cpu.ex.r_8[9] ;
 wire \cpu.ex.r_9[0] ;
 wire \cpu.ex.r_9[10] ;
 wire \cpu.ex.r_9[11] ;
 wire \cpu.ex.r_9[12] ;
 wire \cpu.ex.r_9[13] ;
 wire \cpu.ex.r_9[14] ;
 wire \cpu.ex.r_9[15] ;
 wire \cpu.ex.r_9[1] ;
 wire \cpu.ex.r_9[2] ;
 wire \cpu.ex.r_9[3] ;
 wire \cpu.ex.r_9[4] ;
 wire \cpu.ex.r_9[5] ;
 wire \cpu.ex.r_9[6] ;
 wire \cpu.ex.r_9[7] ;
 wire \cpu.ex.r_9[8] ;
 wire \cpu.ex.r_9[9] ;
 wire \cpu.ex.r_branch_stall ;
 wire \cpu.ex.r_cc ;
 wire \cpu.ex.r_div_running ;
 wire \cpu.ex.r_epc[10] ;
 wire \cpu.ex.r_epc[11] ;
 wire \cpu.ex.r_epc[12] ;
 wire \cpu.ex.r_epc[13] ;
 wire \cpu.ex.r_epc[14] ;
 wire \cpu.ex.r_epc[15] ;
 wire \cpu.ex.r_epc[1] ;
 wire \cpu.ex.r_epc[2] ;
 wire \cpu.ex.r_epc[3] ;
 wire \cpu.ex.r_epc[4] ;
 wire \cpu.ex.r_epc[5] ;
 wire \cpu.ex.r_epc[6] ;
 wire \cpu.ex.r_epc[7] ;
 wire \cpu.ex.r_epc[8] ;
 wire \cpu.ex.r_epc[9] ;
 wire \cpu.ex.r_ie ;
 wire \cpu.ex.r_lr[10] ;
 wire \cpu.ex.r_lr[11] ;
 wire \cpu.ex.r_lr[12] ;
 wire \cpu.ex.r_lr[13] ;
 wire \cpu.ex.r_lr[14] ;
 wire \cpu.ex.r_lr[15] ;
 wire \cpu.ex.r_lr[1] ;
 wire \cpu.ex.r_lr[2] ;
 wire \cpu.ex.r_lr[3] ;
 wire \cpu.ex.r_lr[4] ;
 wire \cpu.ex.r_lr[5] ;
 wire \cpu.ex.r_lr[6] ;
 wire \cpu.ex.r_lr[7] ;
 wire \cpu.ex.r_lr[8] ;
 wire \cpu.ex.r_lr[9] ;
 wire \cpu.ex.r_mult[0] ;
 wire \cpu.ex.r_mult[10] ;
 wire \cpu.ex.r_mult[11] ;
 wire \cpu.ex.r_mult[12] ;
 wire \cpu.ex.r_mult[13] ;
 wire \cpu.ex.r_mult[14] ;
 wire \cpu.ex.r_mult[15] ;
 wire \cpu.ex.r_mult[16] ;
 wire \cpu.ex.r_mult[17] ;
 wire \cpu.ex.r_mult[18] ;
 wire \cpu.ex.r_mult[19] ;
 wire \cpu.ex.r_mult[1] ;
 wire \cpu.ex.r_mult[20] ;
 wire \cpu.ex.r_mult[21] ;
 wire \cpu.ex.r_mult[22] ;
 wire \cpu.ex.r_mult[23] ;
 wire \cpu.ex.r_mult[24] ;
 wire \cpu.ex.r_mult[25] ;
 wire \cpu.ex.r_mult[26] ;
 wire \cpu.ex.r_mult[27] ;
 wire \cpu.ex.r_mult[28] ;
 wire \cpu.ex.r_mult[29] ;
 wire \cpu.ex.r_mult[2] ;
 wire \cpu.ex.r_mult[30] ;
 wire \cpu.ex.r_mult[31] ;
 wire \cpu.ex.r_mult[3] ;
 wire \cpu.ex.r_mult[4] ;
 wire \cpu.ex.r_mult[5] ;
 wire \cpu.ex.r_mult[6] ;
 wire \cpu.ex.r_mult[7] ;
 wire \cpu.ex.r_mult[8] ;
 wire \cpu.ex.r_mult[9] ;
 wire \cpu.ex.r_mult_off[0] ;
 wire \cpu.ex.r_mult_off[1] ;
 wire \cpu.ex.r_mult_off[2] ;
 wire \cpu.ex.r_mult_off[3] ;
 wire \cpu.ex.r_mult_running ;
 wire \cpu.ex.r_prev_ie ;
 wire \cpu.ex.r_read_stall ;
 wire \cpu.ex.r_set_cc ;
 wire \cpu.ex.r_sp[10] ;
 wire \cpu.ex.r_sp[11] ;
 wire \cpu.ex.r_sp[12] ;
 wire \cpu.ex.r_sp[13] ;
 wire \cpu.ex.r_sp[14] ;
 wire \cpu.ex.r_sp[15] ;
 wire \cpu.ex.r_sp[1] ;
 wire \cpu.ex.r_sp[2] ;
 wire \cpu.ex.r_sp[3] ;
 wire \cpu.ex.r_sp[4] ;
 wire \cpu.ex.r_sp[5] ;
 wire \cpu.ex.r_sp[6] ;
 wire \cpu.ex.r_sp[7] ;
 wire \cpu.ex.r_sp[8] ;
 wire \cpu.ex.r_sp[9] ;
 wire \cpu.ex.r_stmp[0] ;
 wire \cpu.ex.r_stmp[10] ;
 wire \cpu.ex.r_stmp[11] ;
 wire \cpu.ex.r_stmp[12] ;
 wire \cpu.ex.r_stmp[13] ;
 wire \cpu.ex.r_stmp[14] ;
 wire \cpu.ex.r_stmp[15] ;
 wire \cpu.ex.r_stmp[1] ;
 wire \cpu.ex.r_stmp[2] ;
 wire \cpu.ex.r_stmp[3] ;
 wire \cpu.ex.r_stmp[4] ;
 wire \cpu.ex.r_stmp[5] ;
 wire \cpu.ex.r_stmp[6] ;
 wire \cpu.ex.r_stmp[7] ;
 wire \cpu.ex.r_stmp[8] ;
 wire \cpu.ex.r_stmp[9] ;
 wire \cpu.ex.r_wb_addr[0] ;
 wire \cpu.ex.r_wb_addr[1] ;
 wire \cpu.ex.r_wb_addr[2] ;
 wire \cpu.ex.r_wb_addr[3] ;
 wire \cpu.ex.r_wb_swapsp ;
 wire \cpu.ex.r_wb_valid ;
 wire \cpu.ex.r_wmask[0] ;
 wire \cpu.ex.r_wmask[1] ;
 wire \cpu.genblk1.mmu.r_valid_d[0] ;
 wire \cpu.genblk1.mmu.r_valid_d[10] ;
 wire \cpu.genblk1.mmu.r_valid_d[11] ;
 wire \cpu.genblk1.mmu.r_valid_d[12] ;
 wire \cpu.genblk1.mmu.r_valid_d[13] ;
 wire \cpu.genblk1.mmu.r_valid_d[14] ;
 wire \cpu.genblk1.mmu.r_valid_d[15] ;
 wire \cpu.genblk1.mmu.r_valid_d[16] ;
 wire \cpu.genblk1.mmu.r_valid_d[17] ;
 wire \cpu.genblk1.mmu.r_valid_d[18] ;
 wire \cpu.genblk1.mmu.r_valid_d[19] ;
 wire \cpu.genblk1.mmu.r_valid_d[1] ;
 wire \cpu.genblk1.mmu.r_valid_d[20] ;
 wire \cpu.genblk1.mmu.r_valid_d[21] ;
 wire \cpu.genblk1.mmu.r_valid_d[22] ;
 wire \cpu.genblk1.mmu.r_valid_d[23] ;
 wire \cpu.genblk1.mmu.r_valid_d[24] ;
 wire \cpu.genblk1.mmu.r_valid_d[25] ;
 wire \cpu.genblk1.mmu.r_valid_d[26] ;
 wire \cpu.genblk1.mmu.r_valid_d[27] ;
 wire \cpu.genblk1.mmu.r_valid_d[28] ;
 wire \cpu.genblk1.mmu.r_valid_d[29] ;
 wire \cpu.genblk1.mmu.r_valid_d[2] ;
 wire \cpu.genblk1.mmu.r_valid_d[30] ;
 wire \cpu.genblk1.mmu.r_valid_d[31] ;
 wire \cpu.genblk1.mmu.r_valid_d[3] ;
 wire \cpu.genblk1.mmu.r_valid_d[4] ;
 wire \cpu.genblk1.mmu.r_valid_d[5] ;
 wire \cpu.genblk1.mmu.r_valid_d[6] ;
 wire \cpu.genblk1.mmu.r_valid_d[7] ;
 wire \cpu.genblk1.mmu.r_valid_d[8] ;
 wire \cpu.genblk1.mmu.r_valid_d[9] ;
 wire \cpu.genblk1.mmu.r_valid_i[0] ;
 wire \cpu.genblk1.mmu.r_valid_i[10] ;
 wire \cpu.genblk1.mmu.r_valid_i[11] ;
 wire \cpu.genblk1.mmu.r_valid_i[12] ;
 wire \cpu.genblk1.mmu.r_valid_i[13] ;
 wire \cpu.genblk1.mmu.r_valid_i[14] ;
 wire \cpu.genblk1.mmu.r_valid_i[15] ;
 wire \cpu.genblk1.mmu.r_valid_i[16] ;
 wire \cpu.genblk1.mmu.r_valid_i[17] ;
 wire \cpu.genblk1.mmu.r_valid_i[18] ;
 wire \cpu.genblk1.mmu.r_valid_i[19] ;
 wire \cpu.genblk1.mmu.r_valid_i[1] ;
 wire \cpu.genblk1.mmu.r_valid_i[20] ;
 wire \cpu.genblk1.mmu.r_valid_i[21] ;
 wire \cpu.genblk1.mmu.r_valid_i[22] ;
 wire \cpu.genblk1.mmu.r_valid_i[23] ;
 wire \cpu.genblk1.mmu.r_valid_i[24] ;
 wire \cpu.genblk1.mmu.r_valid_i[25] ;
 wire \cpu.genblk1.mmu.r_valid_i[26] ;
 wire \cpu.genblk1.mmu.r_valid_i[27] ;
 wire \cpu.genblk1.mmu.r_valid_i[28] ;
 wire \cpu.genblk1.mmu.r_valid_i[29] ;
 wire \cpu.genblk1.mmu.r_valid_i[2] ;
 wire \cpu.genblk1.mmu.r_valid_i[30] ;
 wire \cpu.genblk1.mmu.r_valid_i[31] ;
 wire \cpu.genblk1.mmu.r_valid_i[3] ;
 wire \cpu.genblk1.mmu.r_valid_i[4] ;
 wire \cpu.genblk1.mmu.r_valid_i[5] ;
 wire \cpu.genblk1.mmu.r_valid_i[6] ;
 wire \cpu.genblk1.mmu.r_valid_i[7] ;
 wire \cpu.genblk1.mmu.r_valid_i[8] ;
 wire \cpu.genblk1.mmu.r_valid_i[9] ;
 wire \cpu.genblk1.mmu.r_vtop_d[0][0] ;
 wire \cpu.genblk1.mmu.r_vtop_d[0][10] ;
 wire \cpu.genblk1.mmu.r_vtop_d[0][11] ;
 wire \cpu.genblk1.mmu.r_vtop_d[0][1] ;
 wire \cpu.genblk1.mmu.r_vtop_d[0][2] ;
 wire \cpu.genblk1.mmu.r_vtop_d[0][3] ;
 wire \cpu.genblk1.mmu.r_vtop_d[0][4] ;
 wire \cpu.genblk1.mmu.r_vtop_d[0][5] ;
 wire \cpu.genblk1.mmu.r_vtop_d[0][6] ;
 wire \cpu.genblk1.mmu.r_vtop_d[0][7] ;
 wire \cpu.genblk1.mmu.r_vtop_d[0][8] ;
 wire \cpu.genblk1.mmu.r_vtop_d[0][9] ;
 wire \cpu.genblk1.mmu.r_vtop_d[10][0] ;
 wire \cpu.genblk1.mmu.r_vtop_d[10][10] ;
 wire \cpu.genblk1.mmu.r_vtop_d[10][11] ;
 wire \cpu.genblk1.mmu.r_vtop_d[10][1] ;
 wire \cpu.genblk1.mmu.r_vtop_d[10][2] ;
 wire \cpu.genblk1.mmu.r_vtop_d[10][3] ;
 wire \cpu.genblk1.mmu.r_vtop_d[10][4] ;
 wire \cpu.genblk1.mmu.r_vtop_d[10][5] ;
 wire \cpu.genblk1.mmu.r_vtop_d[10][6] ;
 wire \cpu.genblk1.mmu.r_vtop_d[10][7] ;
 wire \cpu.genblk1.mmu.r_vtop_d[10][8] ;
 wire \cpu.genblk1.mmu.r_vtop_d[10][9] ;
 wire \cpu.genblk1.mmu.r_vtop_d[11][0] ;
 wire \cpu.genblk1.mmu.r_vtop_d[11][10] ;
 wire \cpu.genblk1.mmu.r_vtop_d[11][11] ;
 wire \cpu.genblk1.mmu.r_vtop_d[11][1] ;
 wire \cpu.genblk1.mmu.r_vtop_d[11][2] ;
 wire \cpu.genblk1.mmu.r_vtop_d[11][3] ;
 wire \cpu.genblk1.mmu.r_vtop_d[11][4] ;
 wire \cpu.genblk1.mmu.r_vtop_d[11][5] ;
 wire \cpu.genblk1.mmu.r_vtop_d[11][6] ;
 wire \cpu.genblk1.mmu.r_vtop_d[11][7] ;
 wire \cpu.genblk1.mmu.r_vtop_d[11][8] ;
 wire \cpu.genblk1.mmu.r_vtop_d[11][9] ;
 wire \cpu.genblk1.mmu.r_vtop_d[12][0] ;
 wire \cpu.genblk1.mmu.r_vtop_d[12][10] ;
 wire \cpu.genblk1.mmu.r_vtop_d[12][11] ;
 wire \cpu.genblk1.mmu.r_vtop_d[12][1] ;
 wire \cpu.genblk1.mmu.r_vtop_d[12][2] ;
 wire \cpu.genblk1.mmu.r_vtop_d[12][3] ;
 wire \cpu.genblk1.mmu.r_vtop_d[12][4] ;
 wire \cpu.genblk1.mmu.r_vtop_d[12][5] ;
 wire \cpu.genblk1.mmu.r_vtop_d[12][6] ;
 wire \cpu.genblk1.mmu.r_vtop_d[12][7] ;
 wire \cpu.genblk1.mmu.r_vtop_d[12][8] ;
 wire \cpu.genblk1.mmu.r_vtop_d[12][9] ;
 wire \cpu.genblk1.mmu.r_vtop_d[13][0] ;
 wire \cpu.genblk1.mmu.r_vtop_d[13][10] ;
 wire \cpu.genblk1.mmu.r_vtop_d[13][11] ;
 wire \cpu.genblk1.mmu.r_vtop_d[13][1] ;
 wire \cpu.genblk1.mmu.r_vtop_d[13][2] ;
 wire \cpu.genblk1.mmu.r_vtop_d[13][3] ;
 wire \cpu.genblk1.mmu.r_vtop_d[13][4] ;
 wire \cpu.genblk1.mmu.r_vtop_d[13][5] ;
 wire \cpu.genblk1.mmu.r_vtop_d[13][6] ;
 wire \cpu.genblk1.mmu.r_vtop_d[13][7] ;
 wire \cpu.genblk1.mmu.r_vtop_d[13][8] ;
 wire \cpu.genblk1.mmu.r_vtop_d[13][9] ;
 wire \cpu.genblk1.mmu.r_vtop_d[14][0] ;
 wire \cpu.genblk1.mmu.r_vtop_d[14][10] ;
 wire \cpu.genblk1.mmu.r_vtop_d[14][11] ;
 wire \cpu.genblk1.mmu.r_vtop_d[14][1] ;
 wire \cpu.genblk1.mmu.r_vtop_d[14][2] ;
 wire \cpu.genblk1.mmu.r_vtop_d[14][3] ;
 wire \cpu.genblk1.mmu.r_vtop_d[14][4] ;
 wire \cpu.genblk1.mmu.r_vtop_d[14][5] ;
 wire \cpu.genblk1.mmu.r_vtop_d[14][6] ;
 wire \cpu.genblk1.mmu.r_vtop_d[14][7] ;
 wire \cpu.genblk1.mmu.r_vtop_d[14][8] ;
 wire \cpu.genblk1.mmu.r_vtop_d[14][9] ;
 wire \cpu.genblk1.mmu.r_vtop_d[15][0] ;
 wire \cpu.genblk1.mmu.r_vtop_d[15][10] ;
 wire \cpu.genblk1.mmu.r_vtop_d[15][11] ;
 wire \cpu.genblk1.mmu.r_vtop_d[15][1] ;
 wire \cpu.genblk1.mmu.r_vtop_d[15][2] ;
 wire \cpu.genblk1.mmu.r_vtop_d[15][3] ;
 wire \cpu.genblk1.mmu.r_vtop_d[15][4] ;
 wire \cpu.genblk1.mmu.r_vtop_d[15][5] ;
 wire \cpu.genblk1.mmu.r_vtop_d[15][6] ;
 wire \cpu.genblk1.mmu.r_vtop_d[15][7] ;
 wire \cpu.genblk1.mmu.r_vtop_d[15][8] ;
 wire \cpu.genblk1.mmu.r_vtop_d[15][9] ;
 wire \cpu.genblk1.mmu.r_vtop_d[16][0] ;
 wire \cpu.genblk1.mmu.r_vtop_d[16][10] ;
 wire \cpu.genblk1.mmu.r_vtop_d[16][11] ;
 wire \cpu.genblk1.mmu.r_vtop_d[16][1] ;
 wire \cpu.genblk1.mmu.r_vtop_d[16][2] ;
 wire \cpu.genblk1.mmu.r_vtop_d[16][3] ;
 wire \cpu.genblk1.mmu.r_vtop_d[16][4] ;
 wire \cpu.genblk1.mmu.r_vtop_d[16][5] ;
 wire \cpu.genblk1.mmu.r_vtop_d[16][6] ;
 wire \cpu.genblk1.mmu.r_vtop_d[16][7] ;
 wire \cpu.genblk1.mmu.r_vtop_d[16][8] ;
 wire \cpu.genblk1.mmu.r_vtop_d[16][9] ;
 wire \cpu.genblk1.mmu.r_vtop_d[17][0] ;
 wire \cpu.genblk1.mmu.r_vtop_d[17][10] ;
 wire \cpu.genblk1.mmu.r_vtop_d[17][11] ;
 wire \cpu.genblk1.mmu.r_vtop_d[17][1] ;
 wire \cpu.genblk1.mmu.r_vtop_d[17][2] ;
 wire \cpu.genblk1.mmu.r_vtop_d[17][3] ;
 wire \cpu.genblk1.mmu.r_vtop_d[17][4] ;
 wire \cpu.genblk1.mmu.r_vtop_d[17][5] ;
 wire \cpu.genblk1.mmu.r_vtop_d[17][6] ;
 wire \cpu.genblk1.mmu.r_vtop_d[17][7] ;
 wire \cpu.genblk1.mmu.r_vtop_d[17][8] ;
 wire \cpu.genblk1.mmu.r_vtop_d[17][9] ;
 wire \cpu.genblk1.mmu.r_vtop_d[18][0] ;
 wire \cpu.genblk1.mmu.r_vtop_d[18][10] ;
 wire \cpu.genblk1.mmu.r_vtop_d[18][11] ;
 wire \cpu.genblk1.mmu.r_vtop_d[18][1] ;
 wire \cpu.genblk1.mmu.r_vtop_d[18][2] ;
 wire \cpu.genblk1.mmu.r_vtop_d[18][3] ;
 wire \cpu.genblk1.mmu.r_vtop_d[18][4] ;
 wire \cpu.genblk1.mmu.r_vtop_d[18][5] ;
 wire \cpu.genblk1.mmu.r_vtop_d[18][6] ;
 wire \cpu.genblk1.mmu.r_vtop_d[18][7] ;
 wire \cpu.genblk1.mmu.r_vtop_d[18][8] ;
 wire \cpu.genblk1.mmu.r_vtop_d[18][9] ;
 wire \cpu.genblk1.mmu.r_vtop_d[19][0] ;
 wire \cpu.genblk1.mmu.r_vtop_d[19][10] ;
 wire \cpu.genblk1.mmu.r_vtop_d[19][11] ;
 wire \cpu.genblk1.mmu.r_vtop_d[19][1] ;
 wire \cpu.genblk1.mmu.r_vtop_d[19][2] ;
 wire \cpu.genblk1.mmu.r_vtop_d[19][3] ;
 wire \cpu.genblk1.mmu.r_vtop_d[19][4] ;
 wire \cpu.genblk1.mmu.r_vtop_d[19][5] ;
 wire \cpu.genblk1.mmu.r_vtop_d[19][6] ;
 wire \cpu.genblk1.mmu.r_vtop_d[19][7] ;
 wire \cpu.genblk1.mmu.r_vtop_d[19][8] ;
 wire \cpu.genblk1.mmu.r_vtop_d[19][9] ;
 wire \cpu.genblk1.mmu.r_vtop_d[1][0] ;
 wire \cpu.genblk1.mmu.r_vtop_d[1][10] ;
 wire \cpu.genblk1.mmu.r_vtop_d[1][11] ;
 wire \cpu.genblk1.mmu.r_vtop_d[1][1] ;
 wire \cpu.genblk1.mmu.r_vtop_d[1][2] ;
 wire \cpu.genblk1.mmu.r_vtop_d[1][3] ;
 wire \cpu.genblk1.mmu.r_vtop_d[1][4] ;
 wire \cpu.genblk1.mmu.r_vtop_d[1][5] ;
 wire \cpu.genblk1.mmu.r_vtop_d[1][6] ;
 wire \cpu.genblk1.mmu.r_vtop_d[1][7] ;
 wire \cpu.genblk1.mmu.r_vtop_d[1][8] ;
 wire \cpu.genblk1.mmu.r_vtop_d[1][9] ;
 wire \cpu.genblk1.mmu.r_vtop_d[20][0] ;
 wire \cpu.genblk1.mmu.r_vtop_d[20][10] ;
 wire \cpu.genblk1.mmu.r_vtop_d[20][11] ;
 wire \cpu.genblk1.mmu.r_vtop_d[20][1] ;
 wire \cpu.genblk1.mmu.r_vtop_d[20][2] ;
 wire \cpu.genblk1.mmu.r_vtop_d[20][3] ;
 wire \cpu.genblk1.mmu.r_vtop_d[20][4] ;
 wire \cpu.genblk1.mmu.r_vtop_d[20][5] ;
 wire \cpu.genblk1.mmu.r_vtop_d[20][6] ;
 wire \cpu.genblk1.mmu.r_vtop_d[20][7] ;
 wire \cpu.genblk1.mmu.r_vtop_d[20][8] ;
 wire \cpu.genblk1.mmu.r_vtop_d[20][9] ;
 wire \cpu.genblk1.mmu.r_vtop_d[21][0] ;
 wire \cpu.genblk1.mmu.r_vtop_d[21][10] ;
 wire \cpu.genblk1.mmu.r_vtop_d[21][11] ;
 wire \cpu.genblk1.mmu.r_vtop_d[21][1] ;
 wire \cpu.genblk1.mmu.r_vtop_d[21][2] ;
 wire \cpu.genblk1.mmu.r_vtop_d[21][3] ;
 wire \cpu.genblk1.mmu.r_vtop_d[21][4] ;
 wire \cpu.genblk1.mmu.r_vtop_d[21][5] ;
 wire \cpu.genblk1.mmu.r_vtop_d[21][6] ;
 wire \cpu.genblk1.mmu.r_vtop_d[21][7] ;
 wire \cpu.genblk1.mmu.r_vtop_d[21][8] ;
 wire \cpu.genblk1.mmu.r_vtop_d[21][9] ;
 wire \cpu.genblk1.mmu.r_vtop_d[22][0] ;
 wire \cpu.genblk1.mmu.r_vtop_d[22][10] ;
 wire \cpu.genblk1.mmu.r_vtop_d[22][11] ;
 wire \cpu.genblk1.mmu.r_vtop_d[22][1] ;
 wire \cpu.genblk1.mmu.r_vtop_d[22][2] ;
 wire \cpu.genblk1.mmu.r_vtop_d[22][3] ;
 wire \cpu.genblk1.mmu.r_vtop_d[22][4] ;
 wire \cpu.genblk1.mmu.r_vtop_d[22][5] ;
 wire \cpu.genblk1.mmu.r_vtop_d[22][6] ;
 wire \cpu.genblk1.mmu.r_vtop_d[22][7] ;
 wire \cpu.genblk1.mmu.r_vtop_d[22][8] ;
 wire \cpu.genblk1.mmu.r_vtop_d[22][9] ;
 wire \cpu.genblk1.mmu.r_vtop_d[23][0] ;
 wire \cpu.genblk1.mmu.r_vtop_d[23][10] ;
 wire \cpu.genblk1.mmu.r_vtop_d[23][11] ;
 wire \cpu.genblk1.mmu.r_vtop_d[23][1] ;
 wire \cpu.genblk1.mmu.r_vtop_d[23][2] ;
 wire \cpu.genblk1.mmu.r_vtop_d[23][3] ;
 wire \cpu.genblk1.mmu.r_vtop_d[23][4] ;
 wire \cpu.genblk1.mmu.r_vtop_d[23][5] ;
 wire \cpu.genblk1.mmu.r_vtop_d[23][6] ;
 wire \cpu.genblk1.mmu.r_vtop_d[23][7] ;
 wire \cpu.genblk1.mmu.r_vtop_d[23][8] ;
 wire \cpu.genblk1.mmu.r_vtop_d[23][9] ;
 wire \cpu.genblk1.mmu.r_vtop_d[24][0] ;
 wire \cpu.genblk1.mmu.r_vtop_d[24][10] ;
 wire \cpu.genblk1.mmu.r_vtop_d[24][11] ;
 wire \cpu.genblk1.mmu.r_vtop_d[24][1] ;
 wire \cpu.genblk1.mmu.r_vtop_d[24][2] ;
 wire \cpu.genblk1.mmu.r_vtop_d[24][3] ;
 wire \cpu.genblk1.mmu.r_vtop_d[24][4] ;
 wire \cpu.genblk1.mmu.r_vtop_d[24][5] ;
 wire \cpu.genblk1.mmu.r_vtop_d[24][6] ;
 wire \cpu.genblk1.mmu.r_vtop_d[24][7] ;
 wire \cpu.genblk1.mmu.r_vtop_d[24][8] ;
 wire \cpu.genblk1.mmu.r_vtop_d[24][9] ;
 wire \cpu.genblk1.mmu.r_vtop_d[25][0] ;
 wire \cpu.genblk1.mmu.r_vtop_d[25][10] ;
 wire \cpu.genblk1.mmu.r_vtop_d[25][11] ;
 wire \cpu.genblk1.mmu.r_vtop_d[25][1] ;
 wire \cpu.genblk1.mmu.r_vtop_d[25][2] ;
 wire \cpu.genblk1.mmu.r_vtop_d[25][3] ;
 wire \cpu.genblk1.mmu.r_vtop_d[25][4] ;
 wire \cpu.genblk1.mmu.r_vtop_d[25][5] ;
 wire \cpu.genblk1.mmu.r_vtop_d[25][6] ;
 wire \cpu.genblk1.mmu.r_vtop_d[25][7] ;
 wire \cpu.genblk1.mmu.r_vtop_d[25][8] ;
 wire \cpu.genblk1.mmu.r_vtop_d[25][9] ;
 wire \cpu.genblk1.mmu.r_vtop_d[26][0] ;
 wire \cpu.genblk1.mmu.r_vtop_d[26][10] ;
 wire \cpu.genblk1.mmu.r_vtop_d[26][11] ;
 wire \cpu.genblk1.mmu.r_vtop_d[26][1] ;
 wire \cpu.genblk1.mmu.r_vtop_d[26][2] ;
 wire \cpu.genblk1.mmu.r_vtop_d[26][3] ;
 wire \cpu.genblk1.mmu.r_vtop_d[26][4] ;
 wire \cpu.genblk1.mmu.r_vtop_d[26][5] ;
 wire \cpu.genblk1.mmu.r_vtop_d[26][6] ;
 wire \cpu.genblk1.mmu.r_vtop_d[26][7] ;
 wire \cpu.genblk1.mmu.r_vtop_d[26][8] ;
 wire \cpu.genblk1.mmu.r_vtop_d[26][9] ;
 wire \cpu.genblk1.mmu.r_vtop_d[27][0] ;
 wire \cpu.genblk1.mmu.r_vtop_d[27][10] ;
 wire \cpu.genblk1.mmu.r_vtop_d[27][11] ;
 wire \cpu.genblk1.mmu.r_vtop_d[27][1] ;
 wire \cpu.genblk1.mmu.r_vtop_d[27][2] ;
 wire \cpu.genblk1.mmu.r_vtop_d[27][3] ;
 wire \cpu.genblk1.mmu.r_vtop_d[27][4] ;
 wire \cpu.genblk1.mmu.r_vtop_d[27][5] ;
 wire \cpu.genblk1.mmu.r_vtop_d[27][6] ;
 wire \cpu.genblk1.mmu.r_vtop_d[27][7] ;
 wire \cpu.genblk1.mmu.r_vtop_d[27][8] ;
 wire \cpu.genblk1.mmu.r_vtop_d[27][9] ;
 wire \cpu.genblk1.mmu.r_vtop_d[28][0] ;
 wire \cpu.genblk1.mmu.r_vtop_d[28][10] ;
 wire \cpu.genblk1.mmu.r_vtop_d[28][11] ;
 wire \cpu.genblk1.mmu.r_vtop_d[28][1] ;
 wire \cpu.genblk1.mmu.r_vtop_d[28][2] ;
 wire \cpu.genblk1.mmu.r_vtop_d[28][3] ;
 wire \cpu.genblk1.mmu.r_vtop_d[28][4] ;
 wire \cpu.genblk1.mmu.r_vtop_d[28][5] ;
 wire \cpu.genblk1.mmu.r_vtop_d[28][6] ;
 wire \cpu.genblk1.mmu.r_vtop_d[28][7] ;
 wire \cpu.genblk1.mmu.r_vtop_d[28][8] ;
 wire \cpu.genblk1.mmu.r_vtop_d[28][9] ;
 wire \cpu.genblk1.mmu.r_vtop_d[29][0] ;
 wire \cpu.genblk1.mmu.r_vtop_d[29][10] ;
 wire \cpu.genblk1.mmu.r_vtop_d[29][11] ;
 wire \cpu.genblk1.mmu.r_vtop_d[29][1] ;
 wire \cpu.genblk1.mmu.r_vtop_d[29][2] ;
 wire \cpu.genblk1.mmu.r_vtop_d[29][3] ;
 wire \cpu.genblk1.mmu.r_vtop_d[29][4] ;
 wire \cpu.genblk1.mmu.r_vtop_d[29][5] ;
 wire \cpu.genblk1.mmu.r_vtop_d[29][6] ;
 wire \cpu.genblk1.mmu.r_vtop_d[29][7] ;
 wire \cpu.genblk1.mmu.r_vtop_d[29][8] ;
 wire \cpu.genblk1.mmu.r_vtop_d[29][9] ;
 wire \cpu.genblk1.mmu.r_vtop_d[2][0] ;
 wire \cpu.genblk1.mmu.r_vtop_d[2][10] ;
 wire \cpu.genblk1.mmu.r_vtop_d[2][11] ;
 wire \cpu.genblk1.mmu.r_vtop_d[2][1] ;
 wire \cpu.genblk1.mmu.r_vtop_d[2][2] ;
 wire \cpu.genblk1.mmu.r_vtop_d[2][3] ;
 wire \cpu.genblk1.mmu.r_vtop_d[2][4] ;
 wire \cpu.genblk1.mmu.r_vtop_d[2][5] ;
 wire \cpu.genblk1.mmu.r_vtop_d[2][6] ;
 wire \cpu.genblk1.mmu.r_vtop_d[2][7] ;
 wire \cpu.genblk1.mmu.r_vtop_d[2][8] ;
 wire \cpu.genblk1.mmu.r_vtop_d[2][9] ;
 wire \cpu.genblk1.mmu.r_vtop_d[30][0] ;
 wire \cpu.genblk1.mmu.r_vtop_d[30][10] ;
 wire \cpu.genblk1.mmu.r_vtop_d[30][11] ;
 wire \cpu.genblk1.mmu.r_vtop_d[30][1] ;
 wire \cpu.genblk1.mmu.r_vtop_d[30][2] ;
 wire \cpu.genblk1.mmu.r_vtop_d[30][3] ;
 wire \cpu.genblk1.mmu.r_vtop_d[30][4] ;
 wire \cpu.genblk1.mmu.r_vtop_d[30][5] ;
 wire \cpu.genblk1.mmu.r_vtop_d[30][6] ;
 wire \cpu.genblk1.mmu.r_vtop_d[30][7] ;
 wire \cpu.genblk1.mmu.r_vtop_d[30][8] ;
 wire \cpu.genblk1.mmu.r_vtop_d[30][9] ;
 wire \cpu.genblk1.mmu.r_vtop_d[31][0] ;
 wire \cpu.genblk1.mmu.r_vtop_d[31][10] ;
 wire \cpu.genblk1.mmu.r_vtop_d[31][11] ;
 wire \cpu.genblk1.mmu.r_vtop_d[31][1] ;
 wire \cpu.genblk1.mmu.r_vtop_d[31][2] ;
 wire \cpu.genblk1.mmu.r_vtop_d[31][3] ;
 wire \cpu.genblk1.mmu.r_vtop_d[31][4] ;
 wire \cpu.genblk1.mmu.r_vtop_d[31][5] ;
 wire \cpu.genblk1.mmu.r_vtop_d[31][6] ;
 wire \cpu.genblk1.mmu.r_vtop_d[31][7] ;
 wire \cpu.genblk1.mmu.r_vtop_d[31][8] ;
 wire \cpu.genblk1.mmu.r_vtop_d[31][9] ;
 wire \cpu.genblk1.mmu.r_vtop_d[3][0] ;
 wire \cpu.genblk1.mmu.r_vtop_d[3][10] ;
 wire \cpu.genblk1.mmu.r_vtop_d[3][11] ;
 wire \cpu.genblk1.mmu.r_vtop_d[3][1] ;
 wire \cpu.genblk1.mmu.r_vtop_d[3][2] ;
 wire \cpu.genblk1.mmu.r_vtop_d[3][3] ;
 wire \cpu.genblk1.mmu.r_vtop_d[3][4] ;
 wire \cpu.genblk1.mmu.r_vtop_d[3][5] ;
 wire \cpu.genblk1.mmu.r_vtop_d[3][6] ;
 wire \cpu.genblk1.mmu.r_vtop_d[3][7] ;
 wire \cpu.genblk1.mmu.r_vtop_d[3][8] ;
 wire \cpu.genblk1.mmu.r_vtop_d[3][9] ;
 wire \cpu.genblk1.mmu.r_vtop_d[4][0] ;
 wire \cpu.genblk1.mmu.r_vtop_d[4][10] ;
 wire \cpu.genblk1.mmu.r_vtop_d[4][11] ;
 wire \cpu.genblk1.mmu.r_vtop_d[4][1] ;
 wire \cpu.genblk1.mmu.r_vtop_d[4][2] ;
 wire \cpu.genblk1.mmu.r_vtop_d[4][3] ;
 wire \cpu.genblk1.mmu.r_vtop_d[4][4] ;
 wire \cpu.genblk1.mmu.r_vtop_d[4][5] ;
 wire \cpu.genblk1.mmu.r_vtop_d[4][6] ;
 wire \cpu.genblk1.mmu.r_vtop_d[4][7] ;
 wire \cpu.genblk1.mmu.r_vtop_d[4][8] ;
 wire \cpu.genblk1.mmu.r_vtop_d[4][9] ;
 wire \cpu.genblk1.mmu.r_vtop_d[5][0] ;
 wire \cpu.genblk1.mmu.r_vtop_d[5][10] ;
 wire \cpu.genblk1.mmu.r_vtop_d[5][11] ;
 wire \cpu.genblk1.mmu.r_vtop_d[5][1] ;
 wire \cpu.genblk1.mmu.r_vtop_d[5][2] ;
 wire \cpu.genblk1.mmu.r_vtop_d[5][3] ;
 wire \cpu.genblk1.mmu.r_vtop_d[5][4] ;
 wire \cpu.genblk1.mmu.r_vtop_d[5][5] ;
 wire \cpu.genblk1.mmu.r_vtop_d[5][6] ;
 wire \cpu.genblk1.mmu.r_vtop_d[5][7] ;
 wire \cpu.genblk1.mmu.r_vtop_d[5][8] ;
 wire \cpu.genblk1.mmu.r_vtop_d[5][9] ;
 wire \cpu.genblk1.mmu.r_vtop_d[6][0] ;
 wire \cpu.genblk1.mmu.r_vtop_d[6][10] ;
 wire \cpu.genblk1.mmu.r_vtop_d[6][11] ;
 wire \cpu.genblk1.mmu.r_vtop_d[6][1] ;
 wire \cpu.genblk1.mmu.r_vtop_d[6][2] ;
 wire \cpu.genblk1.mmu.r_vtop_d[6][3] ;
 wire \cpu.genblk1.mmu.r_vtop_d[6][4] ;
 wire \cpu.genblk1.mmu.r_vtop_d[6][5] ;
 wire \cpu.genblk1.mmu.r_vtop_d[6][6] ;
 wire \cpu.genblk1.mmu.r_vtop_d[6][7] ;
 wire \cpu.genblk1.mmu.r_vtop_d[6][8] ;
 wire \cpu.genblk1.mmu.r_vtop_d[6][9] ;
 wire \cpu.genblk1.mmu.r_vtop_d[7][0] ;
 wire \cpu.genblk1.mmu.r_vtop_d[7][10] ;
 wire \cpu.genblk1.mmu.r_vtop_d[7][11] ;
 wire \cpu.genblk1.mmu.r_vtop_d[7][1] ;
 wire \cpu.genblk1.mmu.r_vtop_d[7][2] ;
 wire \cpu.genblk1.mmu.r_vtop_d[7][3] ;
 wire \cpu.genblk1.mmu.r_vtop_d[7][4] ;
 wire \cpu.genblk1.mmu.r_vtop_d[7][5] ;
 wire \cpu.genblk1.mmu.r_vtop_d[7][6] ;
 wire \cpu.genblk1.mmu.r_vtop_d[7][7] ;
 wire \cpu.genblk1.mmu.r_vtop_d[7][8] ;
 wire \cpu.genblk1.mmu.r_vtop_d[7][9] ;
 wire \cpu.genblk1.mmu.r_vtop_d[8][0] ;
 wire \cpu.genblk1.mmu.r_vtop_d[8][10] ;
 wire \cpu.genblk1.mmu.r_vtop_d[8][11] ;
 wire \cpu.genblk1.mmu.r_vtop_d[8][1] ;
 wire \cpu.genblk1.mmu.r_vtop_d[8][2] ;
 wire \cpu.genblk1.mmu.r_vtop_d[8][3] ;
 wire \cpu.genblk1.mmu.r_vtop_d[8][4] ;
 wire \cpu.genblk1.mmu.r_vtop_d[8][5] ;
 wire \cpu.genblk1.mmu.r_vtop_d[8][6] ;
 wire \cpu.genblk1.mmu.r_vtop_d[8][7] ;
 wire \cpu.genblk1.mmu.r_vtop_d[8][8] ;
 wire \cpu.genblk1.mmu.r_vtop_d[8][9] ;
 wire \cpu.genblk1.mmu.r_vtop_d[9][0] ;
 wire \cpu.genblk1.mmu.r_vtop_d[9][10] ;
 wire \cpu.genblk1.mmu.r_vtop_d[9][11] ;
 wire \cpu.genblk1.mmu.r_vtop_d[9][1] ;
 wire \cpu.genblk1.mmu.r_vtop_d[9][2] ;
 wire \cpu.genblk1.mmu.r_vtop_d[9][3] ;
 wire \cpu.genblk1.mmu.r_vtop_d[9][4] ;
 wire \cpu.genblk1.mmu.r_vtop_d[9][5] ;
 wire \cpu.genblk1.mmu.r_vtop_d[9][6] ;
 wire \cpu.genblk1.mmu.r_vtop_d[9][7] ;
 wire \cpu.genblk1.mmu.r_vtop_d[9][8] ;
 wire \cpu.genblk1.mmu.r_vtop_d[9][9] ;
 wire \cpu.genblk1.mmu.r_vtop_i[0][0] ;
 wire \cpu.genblk1.mmu.r_vtop_i[0][10] ;
 wire \cpu.genblk1.mmu.r_vtop_i[0][11] ;
 wire \cpu.genblk1.mmu.r_vtop_i[0][1] ;
 wire \cpu.genblk1.mmu.r_vtop_i[0][2] ;
 wire \cpu.genblk1.mmu.r_vtop_i[0][3] ;
 wire \cpu.genblk1.mmu.r_vtop_i[0][4] ;
 wire \cpu.genblk1.mmu.r_vtop_i[0][5] ;
 wire \cpu.genblk1.mmu.r_vtop_i[0][6] ;
 wire \cpu.genblk1.mmu.r_vtop_i[0][7] ;
 wire \cpu.genblk1.mmu.r_vtop_i[0][8] ;
 wire \cpu.genblk1.mmu.r_vtop_i[0][9] ;
 wire \cpu.genblk1.mmu.r_vtop_i[10][0] ;
 wire \cpu.genblk1.mmu.r_vtop_i[10][10] ;
 wire \cpu.genblk1.mmu.r_vtop_i[10][11] ;
 wire \cpu.genblk1.mmu.r_vtop_i[10][1] ;
 wire \cpu.genblk1.mmu.r_vtop_i[10][2] ;
 wire \cpu.genblk1.mmu.r_vtop_i[10][3] ;
 wire \cpu.genblk1.mmu.r_vtop_i[10][4] ;
 wire \cpu.genblk1.mmu.r_vtop_i[10][5] ;
 wire \cpu.genblk1.mmu.r_vtop_i[10][6] ;
 wire \cpu.genblk1.mmu.r_vtop_i[10][7] ;
 wire \cpu.genblk1.mmu.r_vtop_i[10][8] ;
 wire \cpu.genblk1.mmu.r_vtop_i[10][9] ;
 wire \cpu.genblk1.mmu.r_vtop_i[11][0] ;
 wire \cpu.genblk1.mmu.r_vtop_i[11][10] ;
 wire \cpu.genblk1.mmu.r_vtop_i[11][11] ;
 wire \cpu.genblk1.mmu.r_vtop_i[11][1] ;
 wire \cpu.genblk1.mmu.r_vtop_i[11][2] ;
 wire \cpu.genblk1.mmu.r_vtop_i[11][3] ;
 wire \cpu.genblk1.mmu.r_vtop_i[11][4] ;
 wire \cpu.genblk1.mmu.r_vtop_i[11][5] ;
 wire \cpu.genblk1.mmu.r_vtop_i[11][6] ;
 wire \cpu.genblk1.mmu.r_vtop_i[11][7] ;
 wire \cpu.genblk1.mmu.r_vtop_i[11][8] ;
 wire \cpu.genblk1.mmu.r_vtop_i[11][9] ;
 wire \cpu.genblk1.mmu.r_vtop_i[12][0] ;
 wire \cpu.genblk1.mmu.r_vtop_i[12][10] ;
 wire \cpu.genblk1.mmu.r_vtop_i[12][11] ;
 wire \cpu.genblk1.mmu.r_vtop_i[12][1] ;
 wire \cpu.genblk1.mmu.r_vtop_i[12][2] ;
 wire \cpu.genblk1.mmu.r_vtop_i[12][3] ;
 wire \cpu.genblk1.mmu.r_vtop_i[12][4] ;
 wire \cpu.genblk1.mmu.r_vtop_i[12][5] ;
 wire \cpu.genblk1.mmu.r_vtop_i[12][6] ;
 wire \cpu.genblk1.mmu.r_vtop_i[12][7] ;
 wire \cpu.genblk1.mmu.r_vtop_i[12][8] ;
 wire \cpu.genblk1.mmu.r_vtop_i[12][9] ;
 wire \cpu.genblk1.mmu.r_vtop_i[13][0] ;
 wire \cpu.genblk1.mmu.r_vtop_i[13][10] ;
 wire \cpu.genblk1.mmu.r_vtop_i[13][11] ;
 wire \cpu.genblk1.mmu.r_vtop_i[13][1] ;
 wire \cpu.genblk1.mmu.r_vtop_i[13][2] ;
 wire \cpu.genblk1.mmu.r_vtop_i[13][3] ;
 wire \cpu.genblk1.mmu.r_vtop_i[13][4] ;
 wire \cpu.genblk1.mmu.r_vtop_i[13][5] ;
 wire \cpu.genblk1.mmu.r_vtop_i[13][6] ;
 wire \cpu.genblk1.mmu.r_vtop_i[13][7] ;
 wire \cpu.genblk1.mmu.r_vtop_i[13][8] ;
 wire \cpu.genblk1.mmu.r_vtop_i[13][9] ;
 wire \cpu.genblk1.mmu.r_vtop_i[14][0] ;
 wire \cpu.genblk1.mmu.r_vtop_i[14][10] ;
 wire \cpu.genblk1.mmu.r_vtop_i[14][11] ;
 wire \cpu.genblk1.mmu.r_vtop_i[14][1] ;
 wire \cpu.genblk1.mmu.r_vtop_i[14][2] ;
 wire \cpu.genblk1.mmu.r_vtop_i[14][3] ;
 wire \cpu.genblk1.mmu.r_vtop_i[14][4] ;
 wire \cpu.genblk1.mmu.r_vtop_i[14][5] ;
 wire \cpu.genblk1.mmu.r_vtop_i[14][6] ;
 wire \cpu.genblk1.mmu.r_vtop_i[14][7] ;
 wire \cpu.genblk1.mmu.r_vtop_i[14][8] ;
 wire \cpu.genblk1.mmu.r_vtop_i[14][9] ;
 wire \cpu.genblk1.mmu.r_vtop_i[15][0] ;
 wire \cpu.genblk1.mmu.r_vtop_i[15][10] ;
 wire \cpu.genblk1.mmu.r_vtop_i[15][11] ;
 wire \cpu.genblk1.mmu.r_vtop_i[15][1] ;
 wire \cpu.genblk1.mmu.r_vtop_i[15][2] ;
 wire \cpu.genblk1.mmu.r_vtop_i[15][3] ;
 wire \cpu.genblk1.mmu.r_vtop_i[15][4] ;
 wire \cpu.genblk1.mmu.r_vtop_i[15][5] ;
 wire \cpu.genblk1.mmu.r_vtop_i[15][6] ;
 wire \cpu.genblk1.mmu.r_vtop_i[15][7] ;
 wire \cpu.genblk1.mmu.r_vtop_i[15][8] ;
 wire \cpu.genblk1.mmu.r_vtop_i[15][9] ;
 wire \cpu.genblk1.mmu.r_vtop_i[16][0] ;
 wire \cpu.genblk1.mmu.r_vtop_i[16][10] ;
 wire \cpu.genblk1.mmu.r_vtop_i[16][11] ;
 wire \cpu.genblk1.mmu.r_vtop_i[16][1] ;
 wire \cpu.genblk1.mmu.r_vtop_i[16][2] ;
 wire \cpu.genblk1.mmu.r_vtop_i[16][3] ;
 wire \cpu.genblk1.mmu.r_vtop_i[16][4] ;
 wire \cpu.genblk1.mmu.r_vtop_i[16][5] ;
 wire \cpu.genblk1.mmu.r_vtop_i[16][6] ;
 wire \cpu.genblk1.mmu.r_vtop_i[16][7] ;
 wire \cpu.genblk1.mmu.r_vtop_i[16][8] ;
 wire \cpu.genblk1.mmu.r_vtop_i[16][9] ;
 wire \cpu.genblk1.mmu.r_vtop_i[17][0] ;
 wire \cpu.genblk1.mmu.r_vtop_i[17][10] ;
 wire \cpu.genblk1.mmu.r_vtop_i[17][11] ;
 wire \cpu.genblk1.mmu.r_vtop_i[17][1] ;
 wire \cpu.genblk1.mmu.r_vtop_i[17][2] ;
 wire \cpu.genblk1.mmu.r_vtop_i[17][3] ;
 wire \cpu.genblk1.mmu.r_vtop_i[17][4] ;
 wire \cpu.genblk1.mmu.r_vtop_i[17][5] ;
 wire \cpu.genblk1.mmu.r_vtop_i[17][6] ;
 wire \cpu.genblk1.mmu.r_vtop_i[17][7] ;
 wire \cpu.genblk1.mmu.r_vtop_i[17][8] ;
 wire \cpu.genblk1.mmu.r_vtop_i[17][9] ;
 wire \cpu.genblk1.mmu.r_vtop_i[18][0] ;
 wire \cpu.genblk1.mmu.r_vtop_i[18][10] ;
 wire \cpu.genblk1.mmu.r_vtop_i[18][11] ;
 wire \cpu.genblk1.mmu.r_vtop_i[18][1] ;
 wire \cpu.genblk1.mmu.r_vtop_i[18][2] ;
 wire \cpu.genblk1.mmu.r_vtop_i[18][3] ;
 wire \cpu.genblk1.mmu.r_vtop_i[18][4] ;
 wire \cpu.genblk1.mmu.r_vtop_i[18][5] ;
 wire \cpu.genblk1.mmu.r_vtop_i[18][6] ;
 wire \cpu.genblk1.mmu.r_vtop_i[18][7] ;
 wire \cpu.genblk1.mmu.r_vtop_i[18][8] ;
 wire \cpu.genblk1.mmu.r_vtop_i[18][9] ;
 wire \cpu.genblk1.mmu.r_vtop_i[19][0] ;
 wire \cpu.genblk1.mmu.r_vtop_i[19][10] ;
 wire \cpu.genblk1.mmu.r_vtop_i[19][11] ;
 wire \cpu.genblk1.mmu.r_vtop_i[19][1] ;
 wire \cpu.genblk1.mmu.r_vtop_i[19][2] ;
 wire \cpu.genblk1.mmu.r_vtop_i[19][3] ;
 wire \cpu.genblk1.mmu.r_vtop_i[19][4] ;
 wire \cpu.genblk1.mmu.r_vtop_i[19][5] ;
 wire \cpu.genblk1.mmu.r_vtop_i[19][6] ;
 wire \cpu.genblk1.mmu.r_vtop_i[19][7] ;
 wire \cpu.genblk1.mmu.r_vtop_i[19][8] ;
 wire \cpu.genblk1.mmu.r_vtop_i[19][9] ;
 wire \cpu.genblk1.mmu.r_vtop_i[1][0] ;
 wire \cpu.genblk1.mmu.r_vtop_i[1][10] ;
 wire \cpu.genblk1.mmu.r_vtop_i[1][11] ;
 wire \cpu.genblk1.mmu.r_vtop_i[1][1] ;
 wire \cpu.genblk1.mmu.r_vtop_i[1][2] ;
 wire \cpu.genblk1.mmu.r_vtop_i[1][3] ;
 wire \cpu.genblk1.mmu.r_vtop_i[1][4] ;
 wire \cpu.genblk1.mmu.r_vtop_i[1][5] ;
 wire \cpu.genblk1.mmu.r_vtop_i[1][6] ;
 wire \cpu.genblk1.mmu.r_vtop_i[1][7] ;
 wire \cpu.genblk1.mmu.r_vtop_i[1][8] ;
 wire \cpu.genblk1.mmu.r_vtop_i[1][9] ;
 wire \cpu.genblk1.mmu.r_vtop_i[20][0] ;
 wire \cpu.genblk1.mmu.r_vtop_i[20][10] ;
 wire \cpu.genblk1.mmu.r_vtop_i[20][11] ;
 wire \cpu.genblk1.mmu.r_vtop_i[20][1] ;
 wire \cpu.genblk1.mmu.r_vtop_i[20][2] ;
 wire \cpu.genblk1.mmu.r_vtop_i[20][3] ;
 wire \cpu.genblk1.mmu.r_vtop_i[20][4] ;
 wire \cpu.genblk1.mmu.r_vtop_i[20][5] ;
 wire \cpu.genblk1.mmu.r_vtop_i[20][6] ;
 wire \cpu.genblk1.mmu.r_vtop_i[20][7] ;
 wire \cpu.genblk1.mmu.r_vtop_i[20][8] ;
 wire \cpu.genblk1.mmu.r_vtop_i[20][9] ;
 wire \cpu.genblk1.mmu.r_vtop_i[21][0] ;
 wire \cpu.genblk1.mmu.r_vtop_i[21][10] ;
 wire \cpu.genblk1.mmu.r_vtop_i[21][11] ;
 wire \cpu.genblk1.mmu.r_vtop_i[21][1] ;
 wire \cpu.genblk1.mmu.r_vtop_i[21][2] ;
 wire \cpu.genblk1.mmu.r_vtop_i[21][3] ;
 wire \cpu.genblk1.mmu.r_vtop_i[21][4] ;
 wire \cpu.genblk1.mmu.r_vtop_i[21][5] ;
 wire \cpu.genblk1.mmu.r_vtop_i[21][6] ;
 wire \cpu.genblk1.mmu.r_vtop_i[21][7] ;
 wire \cpu.genblk1.mmu.r_vtop_i[21][8] ;
 wire \cpu.genblk1.mmu.r_vtop_i[21][9] ;
 wire \cpu.genblk1.mmu.r_vtop_i[22][0] ;
 wire \cpu.genblk1.mmu.r_vtop_i[22][10] ;
 wire \cpu.genblk1.mmu.r_vtop_i[22][11] ;
 wire \cpu.genblk1.mmu.r_vtop_i[22][1] ;
 wire \cpu.genblk1.mmu.r_vtop_i[22][2] ;
 wire \cpu.genblk1.mmu.r_vtop_i[22][3] ;
 wire \cpu.genblk1.mmu.r_vtop_i[22][4] ;
 wire \cpu.genblk1.mmu.r_vtop_i[22][5] ;
 wire \cpu.genblk1.mmu.r_vtop_i[22][6] ;
 wire \cpu.genblk1.mmu.r_vtop_i[22][7] ;
 wire \cpu.genblk1.mmu.r_vtop_i[22][8] ;
 wire \cpu.genblk1.mmu.r_vtop_i[22][9] ;
 wire \cpu.genblk1.mmu.r_vtop_i[23][0] ;
 wire \cpu.genblk1.mmu.r_vtop_i[23][10] ;
 wire \cpu.genblk1.mmu.r_vtop_i[23][11] ;
 wire \cpu.genblk1.mmu.r_vtop_i[23][1] ;
 wire \cpu.genblk1.mmu.r_vtop_i[23][2] ;
 wire \cpu.genblk1.mmu.r_vtop_i[23][3] ;
 wire \cpu.genblk1.mmu.r_vtop_i[23][4] ;
 wire \cpu.genblk1.mmu.r_vtop_i[23][5] ;
 wire \cpu.genblk1.mmu.r_vtop_i[23][6] ;
 wire \cpu.genblk1.mmu.r_vtop_i[23][7] ;
 wire \cpu.genblk1.mmu.r_vtop_i[23][8] ;
 wire \cpu.genblk1.mmu.r_vtop_i[23][9] ;
 wire \cpu.genblk1.mmu.r_vtop_i[24][0] ;
 wire \cpu.genblk1.mmu.r_vtop_i[24][10] ;
 wire \cpu.genblk1.mmu.r_vtop_i[24][11] ;
 wire \cpu.genblk1.mmu.r_vtop_i[24][1] ;
 wire \cpu.genblk1.mmu.r_vtop_i[24][2] ;
 wire \cpu.genblk1.mmu.r_vtop_i[24][3] ;
 wire \cpu.genblk1.mmu.r_vtop_i[24][4] ;
 wire \cpu.genblk1.mmu.r_vtop_i[24][5] ;
 wire \cpu.genblk1.mmu.r_vtop_i[24][6] ;
 wire \cpu.genblk1.mmu.r_vtop_i[24][7] ;
 wire \cpu.genblk1.mmu.r_vtop_i[24][8] ;
 wire \cpu.genblk1.mmu.r_vtop_i[24][9] ;
 wire \cpu.genblk1.mmu.r_vtop_i[25][0] ;
 wire \cpu.genblk1.mmu.r_vtop_i[25][10] ;
 wire \cpu.genblk1.mmu.r_vtop_i[25][11] ;
 wire \cpu.genblk1.mmu.r_vtop_i[25][1] ;
 wire \cpu.genblk1.mmu.r_vtop_i[25][2] ;
 wire \cpu.genblk1.mmu.r_vtop_i[25][3] ;
 wire \cpu.genblk1.mmu.r_vtop_i[25][4] ;
 wire \cpu.genblk1.mmu.r_vtop_i[25][5] ;
 wire \cpu.genblk1.mmu.r_vtop_i[25][6] ;
 wire \cpu.genblk1.mmu.r_vtop_i[25][7] ;
 wire \cpu.genblk1.mmu.r_vtop_i[25][8] ;
 wire \cpu.genblk1.mmu.r_vtop_i[25][9] ;
 wire \cpu.genblk1.mmu.r_vtop_i[26][0] ;
 wire \cpu.genblk1.mmu.r_vtop_i[26][10] ;
 wire \cpu.genblk1.mmu.r_vtop_i[26][11] ;
 wire \cpu.genblk1.mmu.r_vtop_i[26][1] ;
 wire \cpu.genblk1.mmu.r_vtop_i[26][2] ;
 wire \cpu.genblk1.mmu.r_vtop_i[26][3] ;
 wire \cpu.genblk1.mmu.r_vtop_i[26][4] ;
 wire \cpu.genblk1.mmu.r_vtop_i[26][5] ;
 wire \cpu.genblk1.mmu.r_vtop_i[26][6] ;
 wire \cpu.genblk1.mmu.r_vtop_i[26][7] ;
 wire \cpu.genblk1.mmu.r_vtop_i[26][8] ;
 wire \cpu.genblk1.mmu.r_vtop_i[26][9] ;
 wire \cpu.genblk1.mmu.r_vtop_i[27][0] ;
 wire \cpu.genblk1.mmu.r_vtop_i[27][10] ;
 wire \cpu.genblk1.mmu.r_vtop_i[27][11] ;
 wire \cpu.genblk1.mmu.r_vtop_i[27][1] ;
 wire \cpu.genblk1.mmu.r_vtop_i[27][2] ;
 wire \cpu.genblk1.mmu.r_vtop_i[27][3] ;
 wire \cpu.genblk1.mmu.r_vtop_i[27][4] ;
 wire \cpu.genblk1.mmu.r_vtop_i[27][5] ;
 wire \cpu.genblk1.mmu.r_vtop_i[27][6] ;
 wire \cpu.genblk1.mmu.r_vtop_i[27][7] ;
 wire \cpu.genblk1.mmu.r_vtop_i[27][8] ;
 wire \cpu.genblk1.mmu.r_vtop_i[27][9] ;
 wire \cpu.genblk1.mmu.r_vtop_i[28][0] ;
 wire \cpu.genblk1.mmu.r_vtop_i[28][10] ;
 wire \cpu.genblk1.mmu.r_vtop_i[28][11] ;
 wire \cpu.genblk1.mmu.r_vtop_i[28][1] ;
 wire \cpu.genblk1.mmu.r_vtop_i[28][2] ;
 wire \cpu.genblk1.mmu.r_vtop_i[28][3] ;
 wire \cpu.genblk1.mmu.r_vtop_i[28][4] ;
 wire \cpu.genblk1.mmu.r_vtop_i[28][5] ;
 wire \cpu.genblk1.mmu.r_vtop_i[28][6] ;
 wire \cpu.genblk1.mmu.r_vtop_i[28][7] ;
 wire \cpu.genblk1.mmu.r_vtop_i[28][8] ;
 wire \cpu.genblk1.mmu.r_vtop_i[28][9] ;
 wire \cpu.genblk1.mmu.r_vtop_i[29][0] ;
 wire \cpu.genblk1.mmu.r_vtop_i[29][10] ;
 wire \cpu.genblk1.mmu.r_vtop_i[29][11] ;
 wire \cpu.genblk1.mmu.r_vtop_i[29][1] ;
 wire \cpu.genblk1.mmu.r_vtop_i[29][2] ;
 wire \cpu.genblk1.mmu.r_vtop_i[29][3] ;
 wire \cpu.genblk1.mmu.r_vtop_i[29][4] ;
 wire \cpu.genblk1.mmu.r_vtop_i[29][5] ;
 wire \cpu.genblk1.mmu.r_vtop_i[29][6] ;
 wire \cpu.genblk1.mmu.r_vtop_i[29][7] ;
 wire \cpu.genblk1.mmu.r_vtop_i[29][8] ;
 wire \cpu.genblk1.mmu.r_vtop_i[29][9] ;
 wire \cpu.genblk1.mmu.r_vtop_i[2][0] ;
 wire \cpu.genblk1.mmu.r_vtop_i[2][10] ;
 wire \cpu.genblk1.mmu.r_vtop_i[2][11] ;
 wire \cpu.genblk1.mmu.r_vtop_i[2][1] ;
 wire \cpu.genblk1.mmu.r_vtop_i[2][2] ;
 wire \cpu.genblk1.mmu.r_vtop_i[2][3] ;
 wire \cpu.genblk1.mmu.r_vtop_i[2][4] ;
 wire \cpu.genblk1.mmu.r_vtop_i[2][5] ;
 wire \cpu.genblk1.mmu.r_vtop_i[2][6] ;
 wire \cpu.genblk1.mmu.r_vtop_i[2][7] ;
 wire \cpu.genblk1.mmu.r_vtop_i[2][8] ;
 wire \cpu.genblk1.mmu.r_vtop_i[2][9] ;
 wire \cpu.genblk1.mmu.r_vtop_i[30][0] ;
 wire \cpu.genblk1.mmu.r_vtop_i[30][10] ;
 wire \cpu.genblk1.mmu.r_vtop_i[30][11] ;
 wire \cpu.genblk1.mmu.r_vtop_i[30][1] ;
 wire \cpu.genblk1.mmu.r_vtop_i[30][2] ;
 wire \cpu.genblk1.mmu.r_vtop_i[30][3] ;
 wire \cpu.genblk1.mmu.r_vtop_i[30][4] ;
 wire \cpu.genblk1.mmu.r_vtop_i[30][5] ;
 wire \cpu.genblk1.mmu.r_vtop_i[30][6] ;
 wire \cpu.genblk1.mmu.r_vtop_i[30][7] ;
 wire \cpu.genblk1.mmu.r_vtop_i[30][8] ;
 wire \cpu.genblk1.mmu.r_vtop_i[30][9] ;
 wire \cpu.genblk1.mmu.r_vtop_i[31][0] ;
 wire \cpu.genblk1.mmu.r_vtop_i[31][10] ;
 wire \cpu.genblk1.mmu.r_vtop_i[31][11] ;
 wire \cpu.genblk1.mmu.r_vtop_i[31][1] ;
 wire \cpu.genblk1.mmu.r_vtop_i[31][2] ;
 wire \cpu.genblk1.mmu.r_vtop_i[31][3] ;
 wire \cpu.genblk1.mmu.r_vtop_i[31][4] ;
 wire \cpu.genblk1.mmu.r_vtop_i[31][5] ;
 wire \cpu.genblk1.mmu.r_vtop_i[31][6] ;
 wire \cpu.genblk1.mmu.r_vtop_i[31][7] ;
 wire \cpu.genblk1.mmu.r_vtop_i[31][8] ;
 wire \cpu.genblk1.mmu.r_vtop_i[31][9] ;
 wire \cpu.genblk1.mmu.r_vtop_i[3][0] ;
 wire \cpu.genblk1.mmu.r_vtop_i[3][10] ;
 wire \cpu.genblk1.mmu.r_vtop_i[3][11] ;
 wire \cpu.genblk1.mmu.r_vtop_i[3][1] ;
 wire \cpu.genblk1.mmu.r_vtop_i[3][2] ;
 wire \cpu.genblk1.mmu.r_vtop_i[3][3] ;
 wire \cpu.genblk1.mmu.r_vtop_i[3][4] ;
 wire \cpu.genblk1.mmu.r_vtop_i[3][5] ;
 wire \cpu.genblk1.mmu.r_vtop_i[3][6] ;
 wire \cpu.genblk1.mmu.r_vtop_i[3][7] ;
 wire \cpu.genblk1.mmu.r_vtop_i[3][8] ;
 wire \cpu.genblk1.mmu.r_vtop_i[3][9] ;
 wire \cpu.genblk1.mmu.r_vtop_i[4][0] ;
 wire \cpu.genblk1.mmu.r_vtop_i[4][10] ;
 wire \cpu.genblk1.mmu.r_vtop_i[4][11] ;
 wire \cpu.genblk1.mmu.r_vtop_i[4][1] ;
 wire \cpu.genblk1.mmu.r_vtop_i[4][2] ;
 wire \cpu.genblk1.mmu.r_vtop_i[4][3] ;
 wire \cpu.genblk1.mmu.r_vtop_i[4][4] ;
 wire \cpu.genblk1.mmu.r_vtop_i[4][5] ;
 wire \cpu.genblk1.mmu.r_vtop_i[4][6] ;
 wire \cpu.genblk1.mmu.r_vtop_i[4][7] ;
 wire \cpu.genblk1.mmu.r_vtop_i[4][8] ;
 wire \cpu.genblk1.mmu.r_vtop_i[4][9] ;
 wire \cpu.genblk1.mmu.r_vtop_i[5][0] ;
 wire \cpu.genblk1.mmu.r_vtop_i[5][10] ;
 wire \cpu.genblk1.mmu.r_vtop_i[5][11] ;
 wire \cpu.genblk1.mmu.r_vtop_i[5][1] ;
 wire \cpu.genblk1.mmu.r_vtop_i[5][2] ;
 wire \cpu.genblk1.mmu.r_vtop_i[5][3] ;
 wire \cpu.genblk1.mmu.r_vtop_i[5][4] ;
 wire \cpu.genblk1.mmu.r_vtop_i[5][5] ;
 wire \cpu.genblk1.mmu.r_vtop_i[5][6] ;
 wire \cpu.genblk1.mmu.r_vtop_i[5][7] ;
 wire \cpu.genblk1.mmu.r_vtop_i[5][8] ;
 wire \cpu.genblk1.mmu.r_vtop_i[5][9] ;
 wire \cpu.genblk1.mmu.r_vtop_i[6][0] ;
 wire \cpu.genblk1.mmu.r_vtop_i[6][10] ;
 wire \cpu.genblk1.mmu.r_vtop_i[6][11] ;
 wire \cpu.genblk1.mmu.r_vtop_i[6][1] ;
 wire \cpu.genblk1.mmu.r_vtop_i[6][2] ;
 wire \cpu.genblk1.mmu.r_vtop_i[6][3] ;
 wire \cpu.genblk1.mmu.r_vtop_i[6][4] ;
 wire \cpu.genblk1.mmu.r_vtop_i[6][5] ;
 wire \cpu.genblk1.mmu.r_vtop_i[6][6] ;
 wire \cpu.genblk1.mmu.r_vtop_i[6][7] ;
 wire \cpu.genblk1.mmu.r_vtop_i[6][8] ;
 wire \cpu.genblk1.mmu.r_vtop_i[6][9] ;
 wire \cpu.genblk1.mmu.r_vtop_i[7][0] ;
 wire \cpu.genblk1.mmu.r_vtop_i[7][10] ;
 wire \cpu.genblk1.mmu.r_vtop_i[7][11] ;
 wire \cpu.genblk1.mmu.r_vtop_i[7][1] ;
 wire \cpu.genblk1.mmu.r_vtop_i[7][2] ;
 wire \cpu.genblk1.mmu.r_vtop_i[7][3] ;
 wire \cpu.genblk1.mmu.r_vtop_i[7][4] ;
 wire \cpu.genblk1.mmu.r_vtop_i[7][5] ;
 wire \cpu.genblk1.mmu.r_vtop_i[7][6] ;
 wire \cpu.genblk1.mmu.r_vtop_i[7][7] ;
 wire \cpu.genblk1.mmu.r_vtop_i[7][8] ;
 wire \cpu.genblk1.mmu.r_vtop_i[7][9] ;
 wire \cpu.genblk1.mmu.r_vtop_i[8][0] ;
 wire \cpu.genblk1.mmu.r_vtop_i[8][10] ;
 wire \cpu.genblk1.mmu.r_vtop_i[8][11] ;
 wire \cpu.genblk1.mmu.r_vtop_i[8][1] ;
 wire \cpu.genblk1.mmu.r_vtop_i[8][2] ;
 wire \cpu.genblk1.mmu.r_vtop_i[8][3] ;
 wire \cpu.genblk1.mmu.r_vtop_i[8][4] ;
 wire \cpu.genblk1.mmu.r_vtop_i[8][5] ;
 wire \cpu.genblk1.mmu.r_vtop_i[8][6] ;
 wire \cpu.genblk1.mmu.r_vtop_i[8][7] ;
 wire \cpu.genblk1.mmu.r_vtop_i[8][8] ;
 wire \cpu.genblk1.mmu.r_vtop_i[8][9] ;
 wire \cpu.genblk1.mmu.r_vtop_i[9][0] ;
 wire \cpu.genblk1.mmu.r_vtop_i[9][10] ;
 wire \cpu.genblk1.mmu.r_vtop_i[9][11] ;
 wire \cpu.genblk1.mmu.r_vtop_i[9][1] ;
 wire \cpu.genblk1.mmu.r_vtop_i[9][2] ;
 wire \cpu.genblk1.mmu.r_vtop_i[9][3] ;
 wire \cpu.genblk1.mmu.r_vtop_i[9][4] ;
 wire \cpu.genblk1.mmu.r_vtop_i[9][5] ;
 wire \cpu.genblk1.mmu.r_vtop_i[9][6] ;
 wire \cpu.genblk1.mmu.r_vtop_i[9][7] ;
 wire \cpu.genblk1.mmu.r_vtop_i[9][8] ;
 wire \cpu.genblk1.mmu.r_vtop_i[9][9] ;
 wire \cpu.genblk1.mmu.r_writeable_d[0] ;
 wire \cpu.genblk1.mmu.r_writeable_d[10] ;
 wire \cpu.genblk1.mmu.r_writeable_d[11] ;
 wire \cpu.genblk1.mmu.r_writeable_d[12] ;
 wire \cpu.genblk1.mmu.r_writeable_d[13] ;
 wire \cpu.genblk1.mmu.r_writeable_d[14] ;
 wire \cpu.genblk1.mmu.r_writeable_d[15] ;
 wire \cpu.genblk1.mmu.r_writeable_d[16] ;
 wire \cpu.genblk1.mmu.r_writeable_d[17] ;
 wire \cpu.genblk1.mmu.r_writeable_d[18] ;
 wire \cpu.genblk1.mmu.r_writeable_d[19] ;
 wire \cpu.genblk1.mmu.r_writeable_d[1] ;
 wire \cpu.genblk1.mmu.r_writeable_d[20] ;
 wire \cpu.genblk1.mmu.r_writeable_d[21] ;
 wire \cpu.genblk1.mmu.r_writeable_d[22] ;
 wire \cpu.genblk1.mmu.r_writeable_d[23] ;
 wire \cpu.genblk1.mmu.r_writeable_d[24] ;
 wire \cpu.genblk1.mmu.r_writeable_d[25] ;
 wire \cpu.genblk1.mmu.r_writeable_d[26] ;
 wire \cpu.genblk1.mmu.r_writeable_d[27] ;
 wire \cpu.genblk1.mmu.r_writeable_d[28] ;
 wire \cpu.genblk1.mmu.r_writeable_d[29] ;
 wire \cpu.genblk1.mmu.r_writeable_d[2] ;
 wire \cpu.genblk1.mmu.r_writeable_d[30] ;
 wire \cpu.genblk1.mmu.r_writeable_d[31] ;
 wire \cpu.genblk1.mmu.r_writeable_d[3] ;
 wire \cpu.genblk1.mmu.r_writeable_d[4] ;
 wire \cpu.genblk1.mmu.r_writeable_d[5] ;
 wire \cpu.genblk1.mmu.r_writeable_d[6] ;
 wire \cpu.genblk1.mmu.r_writeable_d[7] ;
 wire \cpu.genblk1.mmu.r_writeable_d[8] ;
 wire \cpu.genblk1.mmu.r_writeable_d[9] ;
 wire \cpu.gpio.genblk1[3].srcs_o[0] ;
 wire \cpu.gpio.genblk1[3].srcs_o[11] ;
 wire \cpu.gpio.genblk1[3].srcs_o[1] ;
 wire \cpu.gpio.genblk1[3].srcs_o[2] ;
 wire \cpu.gpio.genblk1[3].srcs_o[3] ;
 wire \cpu.gpio.genblk1[3].srcs_o[4] ;
 wire \cpu.gpio.genblk1[3].srcs_o[5] ;
 wire \cpu.gpio.genblk1[3].srcs_o[6] ;
 wire \cpu.gpio.genblk1[3].srcs_o[7] ;
 wire \cpu.gpio.genblk1[3].srcs_o[8] ;
 wire \cpu.gpio.genblk1[4].srcs_o[0] ;
 wire \cpu.gpio.genblk1[5].srcs_o[0] ;
 wire \cpu.gpio.genblk1[6].srcs_o[0] ;
 wire \cpu.gpio.genblk1[7].srcs_o[0] ;
 wire \cpu.gpio.genblk2[4].srcs_io[0] ;
 wire \cpu.gpio.genblk2[5].srcs_io[0] ;
 wire \cpu.gpio.genblk2[6].srcs_io[0] ;
 wire \cpu.gpio.genblk2[7].srcs_io[0] ;
 wire \cpu.gpio.r_enable_in[0] ;
 wire \cpu.gpio.r_enable_in[1] ;
 wire \cpu.gpio.r_enable_in[2] ;
 wire \cpu.gpio.r_enable_in[3] ;
 wire \cpu.gpio.r_enable_in[4] ;
 wire \cpu.gpio.r_enable_in[5] ;
 wire \cpu.gpio.r_enable_in[6] ;
 wire \cpu.gpio.r_enable_in[7] ;
 wire \cpu.gpio.r_enable_io[4] ;
 wire \cpu.gpio.r_enable_io[5] ;
 wire \cpu.gpio.r_enable_io[6] ;
 wire \cpu.gpio.r_enable_io[7] ;
 wire \cpu.gpio.r_spi_miso_src[0][0] ;
 wire \cpu.gpio.r_spi_miso_src[0][1] ;
 wire \cpu.gpio.r_spi_miso_src[0][2] ;
 wire \cpu.gpio.r_spi_miso_src[0][3] ;
 wire \cpu.gpio.r_spi_miso_src[1][0] ;
 wire \cpu.gpio.r_spi_miso_src[1][1] ;
 wire \cpu.gpio.r_spi_miso_src[1][2] ;
 wire \cpu.gpio.r_spi_miso_src[1][3] ;
 wire \cpu.gpio.r_src_io[4][0] ;
 wire \cpu.gpio.r_src_io[4][1] ;
 wire \cpu.gpio.r_src_io[4][2] ;
 wire \cpu.gpio.r_src_io[4][3] ;
 wire \cpu.gpio.r_src_io[5][0] ;
 wire \cpu.gpio.r_src_io[5][1] ;
 wire \cpu.gpio.r_src_io[5][2] ;
 wire \cpu.gpio.r_src_io[5][3] ;
 wire \cpu.gpio.r_src_io[6][0] ;
 wire \cpu.gpio.r_src_io[6][1] ;
 wire \cpu.gpio.r_src_io[6][2] ;
 wire \cpu.gpio.r_src_io[6][3] ;
 wire \cpu.gpio.r_src_io[7][0] ;
 wire \cpu.gpio.r_src_io[7][1] ;
 wire \cpu.gpio.r_src_io[7][2] ;
 wire \cpu.gpio.r_src_io[7][3] ;
 wire \cpu.gpio.r_src_o[3][0] ;
 wire \cpu.gpio.r_src_o[3][1] ;
 wire \cpu.gpio.r_src_o[3][2] ;
 wire \cpu.gpio.r_src_o[3][3] ;
 wire \cpu.gpio.r_src_o[4][0] ;
 wire \cpu.gpio.r_src_o[4][1] ;
 wire \cpu.gpio.r_src_o[4][2] ;
 wire \cpu.gpio.r_src_o[4][3] ;
 wire \cpu.gpio.r_src_o[5][0] ;
 wire \cpu.gpio.r_src_o[5][1] ;
 wire \cpu.gpio.r_src_o[5][2] ;
 wire \cpu.gpio.r_src_o[5][3] ;
 wire \cpu.gpio.r_src_o[6][0] ;
 wire \cpu.gpio.r_src_o[6][1] ;
 wire \cpu.gpio.r_src_o[6][2] ;
 wire \cpu.gpio.r_src_o[6][3] ;
 wire \cpu.gpio.r_src_o[7][0] ;
 wire \cpu.gpio.r_src_o[7][1] ;
 wire \cpu.gpio.r_src_o[7][2] ;
 wire \cpu.gpio.r_src_o[7][3] ;
 wire \cpu.gpio.r_uart_rx_src[0] ;
 wire \cpu.gpio.r_uart_rx_src[1] ;
 wire \cpu.gpio.r_uart_rx_src[2] ;
 wire \cpu.gpio.uart_rx ;
 wire \cpu.i_wstrobe_d ;
 wire \cpu.icache.r_data[0][0] ;
 wire \cpu.icache.r_data[0][10] ;
 wire \cpu.icache.r_data[0][11] ;
 wire \cpu.icache.r_data[0][12] ;
 wire \cpu.icache.r_data[0][13] ;
 wire \cpu.icache.r_data[0][14] ;
 wire \cpu.icache.r_data[0][15] ;
 wire \cpu.icache.r_data[0][16] ;
 wire \cpu.icache.r_data[0][17] ;
 wire \cpu.icache.r_data[0][18] ;
 wire \cpu.icache.r_data[0][19] ;
 wire \cpu.icache.r_data[0][1] ;
 wire \cpu.icache.r_data[0][20] ;
 wire \cpu.icache.r_data[0][21] ;
 wire \cpu.icache.r_data[0][22] ;
 wire \cpu.icache.r_data[0][23] ;
 wire \cpu.icache.r_data[0][24] ;
 wire \cpu.icache.r_data[0][25] ;
 wire \cpu.icache.r_data[0][26] ;
 wire \cpu.icache.r_data[0][27] ;
 wire \cpu.icache.r_data[0][28] ;
 wire \cpu.icache.r_data[0][29] ;
 wire \cpu.icache.r_data[0][2] ;
 wire \cpu.icache.r_data[0][30] ;
 wire \cpu.icache.r_data[0][31] ;
 wire \cpu.icache.r_data[0][3] ;
 wire \cpu.icache.r_data[0][4] ;
 wire \cpu.icache.r_data[0][5] ;
 wire \cpu.icache.r_data[0][6] ;
 wire \cpu.icache.r_data[0][7] ;
 wire \cpu.icache.r_data[0][8] ;
 wire \cpu.icache.r_data[0][9] ;
 wire \cpu.icache.r_data[1][0] ;
 wire \cpu.icache.r_data[1][10] ;
 wire \cpu.icache.r_data[1][11] ;
 wire \cpu.icache.r_data[1][12] ;
 wire \cpu.icache.r_data[1][13] ;
 wire \cpu.icache.r_data[1][14] ;
 wire \cpu.icache.r_data[1][15] ;
 wire \cpu.icache.r_data[1][16] ;
 wire \cpu.icache.r_data[1][17] ;
 wire \cpu.icache.r_data[1][18] ;
 wire \cpu.icache.r_data[1][19] ;
 wire \cpu.icache.r_data[1][1] ;
 wire \cpu.icache.r_data[1][20] ;
 wire \cpu.icache.r_data[1][21] ;
 wire \cpu.icache.r_data[1][22] ;
 wire \cpu.icache.r_data[1][23] ;
 wire \cpu.icache.r_data[1][24] ;
 wire \cpu.icache.r_data[1][25] ;
 wire \cpu.icache.r_data[1][26] ;
 wire \cpu.icache.r_data[1][27] ;
 wire \cpu.icache.r_data[1][28] ;
 wire \cpu.icache.r_data[1][29] ;
 wire \cpu.icache.r_data[1][2] ;
 wire \cpu.icache.r_data[1][30] ;
 wire \cpu.icache.r_data[1][31] ;
 wire \cpu.icache.r_data[1][3] ;
 wire \cpu.icache.r_data[1][4] ;
 wire \cpu.icache.r_data[1][5] ;
 wire \cpu.icache.r_data[1][6] ;
 wire \cpu.icache.r_data[1][7] ;
 wire \cpu.icache.r_data[1][8] ;
 wire \cpu.icache.r_data[1][9] ;
 wire \cpu.icache.r_data[2][0] ;
 wire \cpu.icache.r_data[2][10] ;
 wire \cpu.icache.r_data[2][11] ;
 wire \cpu.icache.r_data[2][12] ;
 wire \cpu.icache.r_data[2][13] ;
 wire \cpu.icache.r_data[2][14] ;
 wire \cpu.icache.r_data[2][15] ;
 wire \cpu.icache.r_data[2][16] ;
 wire \cpu.icache.r_data[2][17] ;
 wire \cpu.icache.r_data[2][18] ;
 wire \cpu.icache.r_data[2][19] ;
 wire \cpu.icache.r_data[2][1] ;
 wire \cpu.icache.r_data[2][20] ;
 wire \cpu.icache.r_data[2][21] ;
 wire \cpu.icache.r_data[2][22] ;
 wire \cpu.icache.r_data[2][23] ;
 wire \cpu.icache.r_data[2][24] ;
 wire \cpu.icache.r_data[2][25] ;
 wire \cpu.icache.r_data[2][26] ;
 wire \cpu.icache.r_data[2][27] ;
 wire \cpu.icache.r_data[2][28] ;
 wire \cpu.icache.r_data[2][29] ;
 wire \cpu.icache.r_data[2][2] ;
 wire \cpu.icache.r_data[2][30] ;
 wire \cpu.icache.r_data[2][31] ;
 wire \cpu.icache.r_data[2][3] ;
 wire \cpu.icache.r_data[2][4] ;
 wire \cpu.icache.r_data[2][5] ;
 wire \cpu.icache.r_data[2][6] ;
 wire \cpu.icache.r_data[2][7] ;
 wire \cpu.icache.r_data[2][8] ;
 wire \cpu.icache.r_data[2][9] ;
 wire \cpu.icache.r_data[3][0] ;
 wire \cpu.icache.r_data[3][10] ;
 wire \cpu.icache.r_data[3][11] ;
 wire \cpu.icache.r_data[3][12] ;
 wire \cpu.icache.r_data[3][13] ;
 wire \cpu.icache.r_data[3][14] ;
 wire \cpu.icache.r_data[3][15] ;
 wire \cpu.icache.r_data[3][16] ;
 wire \cpu.icache.r_data[3][17] ;
 wire \cpu.icache.r_data[3][18] ;
 wire \cpu.icache.r_data[3][19] ;
 wire \cpu.icache.r_data[3][1] ;
 wire \cpu.icache.r_data[3][20] ;
 wire \cpu.icache.r_data[3][21] ;
 wire \cpu.icache.r_data[3][22] ;
 wire \cpu.icache.r_data[3][23] ;
 wire \cpu.icache.r_data[3][24] ;
 wire \cpu.icache.r_data[3][25] ;
 wire \cpu.icache.r_data[3][26] ;
 wire \cpu.icache.r_data[3][27] ;
 wire \cpu.icache.r_data[3][28] ;
 wire \cpu.icache.r_data[3][29] ;
 wire \cpu.icache.r_data[3][2] ;
 wire \cpu.icache.r_data[3][30] ;
 wire \cpu.icache.r_data[3][31] ;
 wire \cpu.icache.r_data[3][3] ;
 wire \cpu.icache.r_data[3][4] ;
 wire \cpu.icache.r_data[3][5] ;
 wire \cpu.icache.r_data[3][6] ;
 wire \cpu.icache.r_data[3][7] ;
 wire \cpu.icache.r_data[3][8] ;
 wire \cpu.icache.r_data[3][9] ;
 wire \cpu.icache.r_data[4][0] ;
 wire \cpu.icache.r_data[4][10] ;
 wire \cpu.icache.r_data[4][11] ;
 wire \cpu.icache.r_data[4][12] ;
 wire \cpu.icache.r_data[4][13] ;
 wire \cpu.icache.r_data[4][14] ;
 wire \cpu.icache.r_data[4][15] ;
 wire \cpu.icache.r_data[4][16] ;
 wire \cpu.icache.r_data[4][17] ;
 wire \cpu.icache.r_data[4][18] ;
 wire \cpu.icache.r_data[4][19] ;
 wire \cpu.icache.r_data[4][1] ;
 wire \cpu.icache.r_data[4][20] ;
 wire \cpu.icache.r_data[4][21] ;
 wire \cpu.icache.r_data[4][22] ;
 wire \cpu.icache.r_data[4][23] ;
 wire \cpu.icache.r_data[4][24] ;
 wire \cpu.icache.r_data[4][25] ;
 wire \cpu.icache.r_data[4][26] ;
 wire \cpu.icache.r_data[4][27] ;
 wire \cpu.icache.r_data[4][28] ;
 wire \cpu.icache.r_data[4][29] ;
 wire \cpu.icache.r_data[4][2] ;
 wire \cpu.icache.r_data[4][30] ;
 wire \cpu.icache.r_data[4][31] ;
 wire \cpu.icache.r_data[4][3] ;
 wire \cpu.icache.r_data[4][4] ;
 wire \cpu.icache.r_data[4][5] ;
 wire \cpu.icache.r_data[4][6] ;
 wire \cpu.icache.r_data[4][7] ;
 wire \cpu.icache.r_data[4][8] ;
 wire \cpu.icache.r_data[4][9] ;
 wire \cpu.icache.r_data[5][0] ;
 wire \cpu.icache.r_data[5][10] ;
 wire \cpu.icache.r_data[5][11] ;
 wire \cpu.icache.r_data[5][12] ;
 wire \cpu.icache.r_data[5][13] ;
 wire \cpu.icache.r_data[5][14] ;
 wire \cpu.icache.r_data[5][15] ;
 wire \cpu.icache.r_data[5][16] ;
 wire \cpu.icache.r_data[5][17] ;
 wire \cpu.icache.r_data[5][18] ;
 wire \cpu.icache.r_data[5][19] ;
 wire \cpu.icache.r_data[5][1] ;
 wire \cpu.icache.r_data[5][20] ;
 wire \cpu.icache.r_data[5][21] ;
 wire \cpu.icache.r_data[5][22] ;
 wire \cpu.icache.r_data[5][23] ;
 wire \cpu.icache.r_data[5][24] ;
 wire \cpu.icache.r_data[5][25] ;
 wire \cpu.icache.r_data[5][26] ;
 wire \cpu.icache.r_data[5][27] ;
 wire \cpu.icache.r_data[5][28] ;
 wire \cpu.icache.r_data[5][29] ;
 wire \cpu.icache.r_data[5][2] ;
 wire \cpu.icache.r_data[5][30] ;
 wire \cpu.icache.r_data[5][31] ;
 wire \cpu.icache.r_data[5][3] ;
 wire \cpu.icache.r_data[5][4] ;
 wire \cpu.icache.r_data[5][5] ;
 wire \cpu.icache.r_data[5][6] ;
 wire \cpu.icache.r_data[5][7] ;
 wire \cpu.icache.r_data[5][8] ;
 wire \cpu.icache.r_data[5][9] ;
 wire \cpu.icache.r_data[6][0] ;
 wire \cpu.icache.r_data[6][10] ;
 wire \cpu.icache.r_data[6][11] ;
 wire \cpu.icache.r_data[6][12] ;
 wire \cpu.icache.r_data[6][13] ;
 wire \cpu.icache.r_data[6][14] ;
 wire \cpu.icache.r_data[6][15] ;
 wire \cpu.icache.r_data[6][16] ;
 wire \cpu.icache.r_data[6][17] ;
 wire \cpu.icache.r_data[6][18] ;
 wire \cpu.icache.r_data[6][19] ;
 wire \cpu.icache.r_data[6][1] ;
 wire \cpu.icache.r_data[6][20] ;
 wire \cpu.icache.r_data[6][21] ;
 wire \cpu.icache.r_data[6][22] ;
 wire \cpu.icache.r_data[6][23] ;
 wire \cpu.icache.r_data[6][24] ;
 wire \cpu.icache.r_data[6][25] ;
 wire \cpu.icache.r_data[6][26] ;
 wire \cpu.icache.r_data[6][27] ;
 wire \cpu.icache.r_data[6][28] ;
 wire \cpu.icache.r_data[6][29] ;
 wire \cpu.icache.r_data[6][2] ;
 wire \cpu.icache.r_data[6][30] ;
 wire \cpu.icache.r_data[6][31] ;
 wire \cpu.icache.r_data[6][3] ;
 wire \cpu.icache.r_data[6][4] ;
 wire \cpu.icache.r_data[6][5] ;
 wire \cpu.icache.r_data[6][6] ;
 wire \cpu.icache.r_data[6][7] ;
 wire \cpu.icache.r_data[6][8] ;
 wire \cpu.icache.r_data[6][9] ;
 wire \cpu.icache.r_data[7][0] ;
 wire \cpu.icache.r_data[7][10] ;
 wire \cpu.icache.r_data[7][11] ;
 wire \cpu.icache.r_data[7][12] ;
 wire \cpu.icache.r_data[7][13] ;
 wire \cpu.icache.r_data[7][14] ;
 wire \cpu.icache.r_data[7][15] ;
 wire \cpu.icache.r_data[7][16] ;
 wire \cpu.icache.r_data[7][17] ;
 wire \cpu.icache.r_data[7][18] ;
 wire \cpu.icache.r_data[7][19] ;
 wire \cpu.icache.r_data[7][1] ;
 wire \cpu.icache.r_data[7][20] ;
 wire \cpu.icache.r_data[7][21] ;
 wire \cpu.icache.r_data[7][22] ;
 wire \cpu.icache.r_data[7][23] ;
 wire \cpu.icache.r_data[7][24] ;
 wire \cpu.icache.r_data[7][25] ;
 wire \cpu.icache.r_data[7][26] ;
 wire \cpu.icache.r_data[7][27] ;
 wire \cpu.icache.r_data[7][28] ;
 wire \cpu.icache.r_data[7][29] ;
 wire \cpu.icache.r_data[7][2] ;
 wire \cpu.icache.r_data[7][30] ;
 wire \cpu.icache.r_data[7][31] ;
 wire \cpu.icache.r_data[7][3] ;
 wire \cpu.icache.r_data[7][4] ;
 wire \cpu.icache.r_data[7][5] ;
 wire \cpu.icache.r_data[7][6] ;
 wire \cpu.icache.r_data[7][7] ;
 wire \cpu.icache.r_data[7][8] ;
 wire \cpu.icache.r_data[7][9] ;
 wire \cpu.icache.r_offset[0] ;
 wire \cpu.icache.r_offset[1] ;
 wire \cpu.icache.r_offset[2] ;
 wire \cpu.icache.r_tag[0][10] ;
 wire \cpu.icache.r_tag[0][11] ;
 wire \cpu.icache.r_tag[0][12] ;
 wire \cpu.icache.r_tag[0][13] ;
 wire \cpu.icache.r_tag[0][14] ;
 wire \cpu.icache.r_tag[0][15] ;
 wire \cpu.icache.r_tag[0][16] ;
 wire \cpu.icache.r_tag[0][17] ;
 wire \cpu.icache.r_tag[0][18] ;
 wire \cpu.icache.r_tag[0][19] ;
 wire \cpu.icache.r_tag[0][20] ;
 wire \cpu.icache.r_tag[0][21] ;
 wire \cpu.icache.r_tag[0][22] ;
 wire \cpu.icache.r_tag[0][23] ;
 wire \cpu.icache.r_tag[0][5] ;
 wire \cpu.icache.r_tag[0][6] ;
 wire \cpu.icache.r_tag[0][7] ;
 wire \cpu.icache.r_tag[0][8] ;
 wire \cpu.icache.r_tag[0][9] ;
 wire \cpu.icache.r_tag[1][10] ;
 wire \cpu.icache.r_tag[1][11] ;
 wire \cpu.icache.r_tag[1][12] ;
 wire \cpu.icache.r_tag[1][13] ;
 wire \cpu.icache.r_tag[1][14] ;
 wire \cpu.icache.r_tag[1][15] ;
 wire \cpu.icache.r_tag[1][16] ;
 wire \cpu.icache.r_tag[1][17] ;
 wire \cpu.icache.r_tag[1][18] ;
 wire \cpu.icache.r_tag[1][19] ;
 wire \cpu.icache.r_tag[1][20] ;
 wire \cpu.icache.r_tag[1][21] ;
 wire \cpu.icache.r_tag[1][22] ;
 wire \cpu.icache.r_tag[1][23] ;
 wire \cpu.icache.r_tag[1][5] ;
 wire \cpu.icache.r_tag[1][6] ;
 wire \cpu.icache.r_tag[1][7] ;
 wire \cpu.icache.r_tag[1][8] ;
 wire \cpu.icache.r_tag[1][9] ;
 wire \cpu.icache.r_tag[2][10] ;
 wire \cpu.icache.r_tag[2][11] ;
 wire \cpu.icache.r_tag[2][12] ;
 wire \cpu.icache.r_tag[2][13] ;
 wire \cpu.icache.r_tag[2][14] ;
 wire \cpu.icache.r_tag[2][15] ;
 wire \cpu.icache.r_tag[2][16] ;
 wire \cpu.icache.r_tag[2][17] ;
 wire \cpu.icache.r_tag[2][18] ;
 wire \cpu.icache.r_tag[2][19] ;
 wire \cpu.icache.r_tag[2][20] ;
 wire \cpu.icache.r_tag[2][21] ;
 wire \cpu.icache.r_tag[2][22] ;
 wire \cpu.icache.r_tag[2][23] ;
 wire \cpu.icache.r_tag[2][5] ;
 wire \cpu.icache.r_tag[2][6] ;
 wire \cpu.icache.r_tag[2][7] ;
 wire \cpu.icache.r_tag[2][8] ;
 wire \cpu.icache.r_tag[2][9] ;
 wire \cpu.icache.r_tag[3][10] ;
 wire \cpu.icache.r_tag[3][11] ;
 wire \cpu.icache.r_tag[3][12] ;
 wire \cpu.icache.r_tag[3][13] ;
 wire \cpu.icache.r_tag[3][14] ;
 wire \cpu.icache.r_tag[3][15] ;
 wire \cpu.icache.r_tag[3][16] ;
 wire \cpu.icache.r_tag[3][17] ;
 wire \cpu.icache.r_tag[3][18] ;
 wire \cpu.icache.r_tag[3][19] ;
 wire \cpu.icache.r_tag[3][20] ;
 wire \cpu.icache.r_tag[3][21] ;
 wire \cpu.icache.r_tag[3][22] ;
 wire \cpu.icache.r_tag[3][23] ;
 wire \cpu.icache.r_tag[3][5] ;
 wire \cpu.icache.r_tag[3][6] ;
 wire \cpu.icache.r_tag[3][7] ;
 wire \cpu.icache.r_tag[3][8] ;
 wire \cpu.icache.r_tag[3][9] ;
 wire \cpu.icache.r_tag[4][10] ;
 wire \cpu.icache.r_tag[4][11] ;
 wire \cpu.icache.r_tag[4][12] ;
 wire \cpu.icache.r_tag[4][13] ;
 wire \cpu.icache.r_tag[4][14] ;
 wire \cpu.icache.r_tag[4][15] ;
 wire \cpu.icache.r_tag[4][16] ;
 wire \cpu.icache.r_tag[4][17] ;
 wire \cpu.icache.r_tag[4][18] ;
 wire \cpu.icache.r_tag[4][19] ;
 wire \cpu.icache.r_tag[4][20] ;
 wire \cpu.icache.r_tag[4][21] ;
 wire \cpu.icache.r_tag[4][22] ;
 wire \cpu.icache.r_tag[4][23] ;
 wire \cpu.icache.r_tag[4][5] ;
 wire \cpu.icache.r_tag[4][6] ;
 wire \cpu.icache.r_tag[4][7] ;
 wire \cpu.icache.r_tag[4][8] ;
 wire \cpu.icache.r_tag[4][9] ;
 wire \cpu.icache.r_tag[5][10] ;
 wire \cpu.icache.r_tag[5][11] ;
 wire \cpu.icache.r_tag[5][12] ;
 wire \cpu.icache.r_tag[5][13] ;
 wire \cpu.icache.r_tag[5][14] ;
 wire \cpu.icache.r_tag[5][15] ;
 wire \cpu.icache.r_tag[5][16] ;
 wire \cpu.icache.r_tag[5][17] ;
 wire \cpu.icache.r_tag[5][18] ;
 wire \cpu.icache.r_tag[5][19] ;
 wire \cpu.icache.r_tag[5][20] ;
 wire \cpu.icache.r_tag[5][21] ;
 wire \cpu.icache.r_tag[5][22] ;
 wire \cpu.icache.r_tag[5][23] ;
 wire \cpu.icache.r_tag[5][5] ;
 wire \cpu.icache.r_tag[5][6] ;
 wire \cpu.icache.r_tag[5][7] ;
 wire \cpu.icache.r_tag[5][8] ;
 wire \cpu.icache.r_tag[5][9] ;
 wire \cpu.icache.r_tag[6][10] ;
 wire \cpu.icache.r_tag[6][11] ;
 wire \cpu.icache.r_tag[6][12] ;
 wire \cpu.icache.r_tag[6][13] ;
 wire \cpu.icache.r_tag[6][14] ;
 wire \cpu.icache.r_tag[6][15] ;
 wire \cpu.icache.r_tag[6][16] ;
 wire \cpu.icache.r_tag[6][17] ;
 wire \cpu.icache.r_tag[6][18] ;
 wire \cpu.icache.r_tag[6][19] ;
 wire \cpu.icache.r_tag[6][20] ;
 wire \cpu.icache.r_tag[6][21] ;
 wire \cpu.icache.r_tag[6][22] ;
 wire \cpu.icache.r_tag[6][23] ;
 wire \cpu.icache.r_tag[6][5] ;
 wire \cpu.icache.r_tag[6][6] ;
 wire \cpu.icache.r_tag[6][7] ;
 wire \cpu.icache.r_tag[6][8] ;
 wire \cpu.icache.r_tag[6][9] ;
 wire \cpu.icache.r_tag[7][10] ;
 wire \cpu.icache.r_tag[7][11] ;
 wire \cpu.icache.r_tag[7][12] ;
 wire \cpu.icache.r_tag[7][13] ;
 wire \cpu.icache.r_tag[7][14] ;
 wire \cpu.icache.r_tag[7][15] ;
 wire \cpu.icache.r_tag[7][16] ;
 wire \cpu.icache.r_tag[7][17] ;
 wire \cpu.icache.r_tag[7][18] ;
 wire \cpu.icache.r_tag[7][19] ;
 wire \cpu.icache.r_tag[7][20] ;
 wire \cpu.icache.r_tag[7][21] ;
 wire \cpu.icache.r_tag[7][22] ;
 wire \cpu.icache.r_tag[7][23] ;
 wire \cpu.icache.r_tag[7][5] ;
 wire \cpu.icache.r_tag[7][6] ;
 wire \cpu.icache.r_tag[7][7] ;
 wire \cpu.icache.r_tag[7][8] ;
 wire \cpu.icache.r_tag[7][9] ;
 wire \cpu.icache.r_valid[0] ;
 wire \cpu.icache.r_valid[1] ;
 wire \cpu.icache.r_valid[2] ;
 wire \cpu.icache.r_valid[3] ;
 wire \cpu.icache.r_valid[4] ;
 wire \cpu.icache.r_valid[5] ;
 wire \cpu.icache.r_valid[6] ;
 wire \cpu.icache.r_valid[7] ;
 wire \cpu.intr.r_clock ;
 wire \cpu.intr.r_clock_cmp[0] ;
 wire \cpu.intr.r_clock_cmp[10] ;
 wire \cpu.intr.r_clock_cmp[11] ;
 wire \cpu.intr.r_clock_cmp[12] ;
 wire \cpu.intr.r_clock_cmp[13] ;
 wire \cpu.intr.r_clock_cmp[14] ;
 wire \cpu.intr.r_clock_cmp[15] ;
 wire \cpu.intr.r_clock_cmp[16] ;
 wire \cpu.intr.r_clock_cmp[17] ;
 wire \cpu.intr.r_clock_cmp[18] ;
 wire \cpu.intr.r_clock_cmp[19] ;
 wire \cpu.intr.r_clock_cmp[1] ;
 wire \cpu.intr.r_clock_cmp[20] ;
 wire \cpu.intr.r_clock_cmp[21] ;
 wire \cpu.intr.r_clock_cmp[22] ;
 wire \cpu.intr.r_clock_cmp[23] ;
 wire \cpu.intr.r_clock_cmp[24] ;
 wire \cpu.intr.r_clock_cmp[25] ;
 wire \cpu.intr.r_clock_cmp[26] ;
 wire \cpu.intr.r_clock_cmp[27] ;
 wire \cpu.intr.r_clock_cmp[28] ;
 wire \cpu.intr.r_clock_cmp[29] ;
 wire \cpu.intr.r_clock_cmp[2] ;
 wire \cpu.intr.r_clock_cmp[30] ;
 wire \cpu.intr.r_clock_cmp[31] ;
 wire \cpu.intr.r_clock_cmp[3] ;
 wire \cpu.intr.r_clock_cmp[4] ;
 wire \cpu.intr.r_clock_cmp[5] ;
 wire \cpu.intr.r_clock_cmp[6] ;
 wire \cpu.intr.r_clock_cmp[7] ;
 wire \cpu.intr.r_clock_cmp[8] ;
 wire \cpu.intr.r_clock_cmp[9] ;
 wire \cpu.intr.r_clock_count[0] ;
 wire \cpu.intr.r_clock_count[10] ;
 wire \cpu.intr.r_clock_count[11] ;
 wire \cpu.intr.r_clock_count[12] ;
 wire \cpu.intr.r_clock_count[13] ;
 wire \cpu.intr.r_clock_count[14] ;
 wire \cpu.intr.r_clock_count[15] ;
 wire \cpu.intr.r_clock_count[16] ;
 wire \cpu.intr.r_clock_count[17] ;
 wire \cpu.intr.r_clock_count[18] ;
 wire \cpu.intr.r_clock_count[19] ;
 wire \cpu.intr.r_clock_count[1] ;
 wire \cpu.intr.r_clock_count[20] ;
 wire \cpu.intr.r_clock_count[21] ;
 wire \cpu.intr.r_clock_count[22] ;
 wire \cpu.intr.r_clock_count[23] ;
 wire \cpu.intr.r_clock_count[24] ;
 wire \cpu.intr.r_clock_count[25] ;
 wire \cpu.intr.r_clock_count[26] ;
 wire \cpu.intr.r_clock_count[27] ;
 wire \cpu.intr.r_clock_count[28] ;
 wire \cpu.intr.r_clock_count[29] ;
 wire \cpu.intr.r_clock_count[2] ;
 wire \cpu.intr.r_clock_count[30] ;
 wire \cpu.intr.r_clock_count[31] ;
 wire \cpu.intr.r_clock_count[3] ;
 wire \cpu.intr.r_clock_count[4] ;
 wire \cpu.intr.r_clock_count[5] ;
 wire \cpu.intr.r_clock_count[6] ;
 wire \cpu.intr.r_clock_count[7] ;
 wire \cpu.intr.r_clock_count[8] ;
 wire \cpu.intr.r_clock_count[9] ;
 wire \cpu.intr.r_enable[0] ;
 wire \cpu.intr.r_enable[1] ;
 wire \cpu.intr.r_enable[2] ;
 wire \cpu.intr.r_enable[3] ;
 wire \cpu.intr.r_enable[4] ;
 wire \cpu.intr.r_enable[5] ;
 wire \cpu.intr.r_swi ;
 wire \cpu.intr.r_timer ;
 wire \cpu.intr.r_timer_count[0] ;
 wire \cpu.intr.r_timer_count[10] ;
 wire \cpu.intr.r_timer_count[11] ;
 wire \cpu.intr.r_timer_count[12] ;
 wire \cpu.intr.r_timer_count[13] ;
 wire \cpu.intr.r_timer_count[14] ;
 wire \cpu.intr.r_timer_count[15] ;
 wire \cpu.intr.r_timer_count[16] ;
 wire \cpu.intr.r_timer_count[17] ;
 wire \cpu.intr.r_timer_count[18] ;
 wire \cpu.intr.r_timer_count[19] ;
 wire \cpu.intr.r_timer_count[1] ;
 wire \cpu.intr.r_timer_count[20] ;
 wire \cpu.intr.r_timer_count[21] ;
 wire \cpu.intr.r_timer_count[22] ;
 wire \cpu.intr.r_timer_count[23] ;
 wire \cpu.intr.r_timer_count[2] ;
 wire \cpu.intr.r_timer_count[3] ;
 wire \cpu.intr.r_timer_count[4] ;
 wire \cpu.intr.r_timer_count[5] ;
 wire \cpu.intr.r_timer_count[6] ;
 wire \cpu.intr.r_timer_count[7] ;
 wire \cpu.intr.r_timer_count[8] ;
 wire \cpu.intr.r_timer_count[9] ;
 wire \cpu.intr.r_timer_reload[0] ;
 wire \cpu.intr.r_timer_reload[10] ;
 wire \cpu.intr.r_timer_reload[11] ;
 wire \cpu.intr.r_timer_reload[12] ;
 wire \cpu.intr.r_timer_reload[13] ;
 wire \cpu.intr.r_timer_reload[14] ;
 wire \cpu.intr.r_timer_reload[15] ;
 wire \cpu.intr.r_timer_reload[16] ;
 wire \cpu.intr.r_timer_reload[17] ;
 wire \cpu.intr.r_timer_reload[18] ;
 wire \cpu.intr.r_timer_reload[19] ;
 wire \cpu.intr.r_timer_reload[1] ;
 wire \cpu.intr.r_timer_reload[20] ;
 wire \cpu.intr.r_timer_reload[21] ;
 wire \cpu.intr.r_timer_reload[22] ;
 wire \cpu.intr.r_timer_reload[23] ;
 wire \cpu.intr.r_timer_reload[2] ;
 wire \cpu.intr.r_timer_reload[3] ;
 wire \cpu.intr.r_timer_reload[4] ;
 wire \cpu.intr.r_timer_reload[5] ;
 wire \cpu.intr.r_timer_reload[6] ;
 wire \cpu.intr.r_timer_reload[7] ;
 wire \cpu.intr.r_timer_reload[8] ;
 wire \cpu.intr.r_timer_reload[9] ;
 wire \cpu.intr.spi_intr ;
 wire \cpu.qspi.c_rstrobe_d ;
 wire \cpu.qspi.c_wstrobe_d ;
 wire \cpu.qspi.c_wstrobe_i ;
 wire \cpu.qspi.r_count[0] ;
 wire \cpu.qspi.r_count[1] ;
 wire \cpu.qspi.r_count[2] ;
 wire \cpu.qspi.r_count[3] ;
 wire \cpu.qspi.r_count[4] ;
 wire \cpu.qspi.r_ind ;
 wire \cpu.qspi.r_mask[0] ;
 wire \cpu.qspi.r_mask[1] ;
 wire \cpu.qspi.r_mask[2] ;
 wire \cpu.qspi.r_quad[0] ;
 wire \cpu.qspi.r_quad[1] ;
 wire \cpu.qspi.r_quad[2] ;
 wire \cpu.qspi.r_read_delay[0][0] ;
 wire \cpu.qspi.r_read_delay[0][1] ;
 wire \cpu.qspi.r_read_delay[0][2] ;
 wire \cpu.qspi.r_read_delay[0][3] ;
 wire \cpu.qspi.r_read_delay[1][0] ;
 wire \cpu.qspi.r_read_delay[1][1] ;
 wire \cpu.qspi.r_read_delay[1][2] ;
 wire \cpu.qspi.r_read_delay[1][3] ;
 wire \cpu.qspi.r_read_delay[2][0] ;
 wire \cpu.qspi.r_read_delay[2][1] ;
 wire \cpu.qspi.r_read_delay[2][2] ;
 wire \cpu.qspi.r_read_delay[2][3] ;
 wire \cpu.qspi.r_rom_mode[0] ;
 wire \cpu.qspi.r_rom_mode[1] ;
 wire \cpu.qspi.r_state[0] ;
 wire \cpu.qspi.r_state[10] ;
 wire \cpu.qspi.r_state[11] ;
 wire \cpu.qspi.r_state[12] ;
 wire \cpu.qspi.r_state[13] ;
 wire \cpu.qspi.r_state[14] ;
 wire \cpu.qspi.r_state[15] ;
 wire \cpu.qspi.r_state[16] ;
 wire \cpu.qspi.r_state[17] ;
 wire \cpu.qspi.r_state[1] ;
 wire \cpu.qspi.r_state[2] ;
 wire \cpu.qspi.r_state[3] ;
 wire \cpu.qspi.r_state[4] ;
 wire \cpu.qspi.r_state[5] ;
 wire \cpu.qspi.r_state[6] ;
 wire \cpu.qspi.r_state[7] ;
 wire \cpu.qspi.r_state[8] ;
 wire \cpu.qspi.r_state[9] ;
 wire \cpu.r_clk_invert ;
 wire \cpu.spi.r_bits[0] ;
 wire \cpu.spi.r_bits[1] ;
 wire \cpu.spi.r_bits[2] ;
 wire \cpu.spi.r_clk_count[0][0] ;
 wire \cpu.spi.r_clk_count[0][1] ;
 wire \cpu.spi.r_clk_count[0][2] ;
 wire \cpu.spi.r_clk_count[0][3] ;
 wire \cpu.spi.r_clk_count[0][4] ;
 wire \cpu.spi.r_clk_count[0][5] ;
 wire \cpu.spi.r_clk_count[0][6] ;
 wire \cpu.spi.r_clk_count[0][7] ;
 wire \cpu.spi.r_clk_count[1][0] ;
 wire \cpu.spi.r_clk_count[1][1] ;
 wire \cpu.spi.r_clk_count[1][2] ;
 wire \cpu.spi.r_clk_count[1][3] ;
 wire \cpu.spi.r_clk_count[1][4] ;
 wire \cpu.spi.r_clk_count[1][5] ;
 wire \cpu.spi.r_clk_count[1][6] ;
 wire \cpu.spi.r_clk_count[1][7] ;
 wire \cpu.spi.r_clk_count[2][0] ;
 wire \cpu.spi.r_clk_count[2][1] ;
 wire \cpu.spi.r_clk_count[2][2] ;
 wire \cpu.spi.r_clk_count[2][3] ;
 wire \cpu.spi.r_clk_count[2][4] ;
 wire \cpu.spi.r_clk_count[2][5] ;
 wire \cpu.spi.r_clk_count[2][6] ;
 wire \cpu.spi.r_clk_count[2][7] ;
 wire \cpu.spi.r_count[0] ;
 wire \cpu.spi.r_count[1] ;
 wire \cpu.spi.r_count[2] ;
 wire \cpu.spi.r_count[3] ;
 wire \cpu.spi.r_count[4] ;
 wire \cpu.spi.r_count[5] ;
 wire \cpu.spi.r_count[6] ;
 wire \cpu.spi.r_count[7] ;
 wire \cpu.spi.r_in[0] ;
 wire \cpu.spi.r_in[1] ;
 wire \cpu.spi.r_in[2] ;
 wire \cpu.spi.r_in[3] ;
 wire \cpu.spi.r_in[4] ;
 wire \cpu.spi.r_in[5] ;
 wire \cpu.spi.r_in[6] ;
 wire \cpu.spi.r_in[7] ;
 wire \cpu.spi.r_mode[0][0] ;
 wire \cpu.spi.r_mode[0][1] ;
 wire \cpu.spi.r_mode[1][0] ;
 wire \cpu.spi.r_mode[1][1] ;
 wire \cpu.spi.r_mode[2][0] ;
 wire \cpu.spi.r_mode[2][1] ;
 wire \cpu.spi.r_out[0] ;
 wire \cpu.spi.r_out[1] ;
 wire \cpu.spi.r_out[2] ;
 wire \cpu.spi.r_out[3] ;
 wire \cpu.spi.r_out[4] ;
 wire \cpu.spi.r_out[5] ;
 wire \cpu.spi.r_out[6] ;
 wire \cpu.spi.r_out[7] ;
 wire \cpu.spi.r_ready ;
 wire \cpu.spi.r_searching ;
 wire \cpu.spi.r_sel[0] ;
 wire \cpu.spi.r_sel[1] ;
 wire \cpu.spi.r_src[0] ;
 wire \cpu.spi.r_src[1] ;
 wire \cpu.spi.r_src[2] ;
 wire \cpu.spi.r_state[0] ;
 wire \cpu.spi.r_state[1] ;
 wire \cpu.spi.r_state[2] ;
 wire \cpu.spi.r_state[3] ;
 wire \cpu.spi.r_state[4] ;
 wire \cpu.spi.r_state[5] ;
 wire \cpu.spi.r_state[6] ;
 wire \cpu.spi.r_timeout[0] ;
 wire \cpu.spi.r_timeout[1] ;
 wire \cpu.spi.r_timeout[2] ;
 wire \cpu.spi.r_timeout[3] ;
 wire \cpu.spi.r_timeout[4] ;
 wire \cpu.spi.r_timeout[5] ;
 wire \cpu.spi.r_timeout[6] ;
 wire \cpu.spi.r_timeout[7] ;
 wire \cpu.spi.r_timeout_count[0] ;
 wire \cpu.spi.r_timeout_count[1] ;
 wire \cpu.spi.r_timeout_count[2] ;
 wire \cpu.spi.r_timeout_count[3] ;
 wire \cpu.spi.r_timeout_count[4] ;
 wire \cpu.spi.r_timeout_count[5] ;
 wire \cpu.spi.r_timeout_count[6] ;
 wire \cpu.spi.r_timeout_count[7] ;
 wire \cpu.uart.r_div[0] ;
 wire \cpu.uart.r_div[10] ;
 wire \cpu.uart.r_div[11] ;
 wire \cpu.uart.r_div[1] ;
 wire \cpu.uart.r_div[2] ;
 wire \cpu.uart.r_div[3] ;
 wire \cpu.uart.r_div[4] ;
 wire \cpu.uart.r_div[5] ;
 wire \cpu.uart.r_div[6] ;
 wire \cpu.uart.r_div[7] ;
 wire \cpu.uart.r_div[8] ;
 wire \cpu.uart.r_div[9] ;
 wire \cpu.uart.r_div_value[0] ;
 wire \cpu.uart.r_div_value[10] ;
 wire \cpu.uart.r_div_value[11] ;
 wire \cpu.uart.r_div_value[1] ;
 wire \cpu.uart.r_div_value[2] ;
 wire \cpu.uart.r_div_value[3] ;
 wire \cpu.uart.r_div_value[4] ;
 wire \cpu.uart.r_div_value[5] ;
 wire \cpu.uart.r_div_value[6] ;
 wire \cpu.uart.r_div_value[7] ;
 wire \cpu.uart.r_div_value[8] ;
 wire \cpu.uart.r_div_value[9] ;
 wire \cpu.uart.r_ib[0] ;
 wire \cpu.uart.r_ib[1] ;
 wire \cpu.uart.r_ib[2] ;
 wire \cpu.uart.r_ib[3] ;
 wire \cpu.uart.r_ib[4] ;
 wire \cpu.uart.r_ib[5] ;
 wire \cpu.uart.r_ib[6] ;
 wire \cpu.uart.r_in[0] ;
 wire \cpu.uart.r_in[1] ;
 wire \cpu.uart.r_in[2] ;
 wire \cpu.uart.r_in[3] ;
 wire \cpu.uart.r_in[4] ;
 wire \cpu.uart.r_in[5] ;
 wire \cpu.uart.r_in[6] ;
 wire \cpu.uart.r_in[7] ;
 wire \cpu.uart.r_out[0] ;
 wire \cpu.uart.r_out[1] ;
 wire \cpu.uart.r_out[2] ;
 wire \cpu.uart.r_out[3] ;
 wire \cpu.uart.r_out[4] ;
 wire \cpu.uart.r_out[5] ;
 wire \cpu.uart.r_out[6] ;
 wire \cpu.uart.r_out[7] ;
 wire \cpu.uart.r_r ;
 wire \cpu.uart.r_r_int ;
 wire \cpu.uart.r_r_invert ;
 wire \cpu.uart.r_rcnt[0] ;
 wire \cpu.uart.r_rcnt[1] ;
 wire \cpu.uart.r_rstate[0] ;
 wire \cpu.uart.r_rstate[1] ;
 wire \cpu.uart.r_rstate[2] ;
 wire \cpu.uart.r_rstate[3] ;
 wire \cpu.uart.r_x_int ;
 wire \cpu.uart.r_x_invert ;
 wire \cpu.uart.r_xcnt[0] ;
 wire \cpu.uart.r_xcnt[1] ;
 wire \cpu.uart.r_xstate[0] ;
 wire \cpu.uart.r_xstate[1] ;
 wire \cpu.uart.r_xstate[2] ;
 wire \cpu.uart.r_xstate[3] ;
 wire r_reset;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net180;
 wire net181;
 wire net182;
 wire net183;
 wire net184;
 wire net185;
 wire net186;
 wire net187;
 wire net188;
 wire net189;
 wire net190;
 wire net191;
 wire net192;
 wire net193;
 wire net194;
 wire net195;
 wire net196;
 wire net197;
 wire net198;
 wire net199;
 wire net200;
 wire net201;
 wire net202;
 wire net203;
 wire net204;
 wire net205;
 wire net206;
 wire net207;
 wire net208;
 wire net209;
 wire net210;
 wire net211;
 wire net212;
 wire net213;
 wire net214;
 wire net215;
 wire net216;
 wire net217;
 wire net218;
 wire net219;
 wire net220;
 wire net221;
 wire net222;
 wire net223;
 wire net224;
 wire net225;
 wire net226;
 wire net227;
 wire net228;
 wire net229;
 wire net230;
 wire net231;
 wire net232;
 wire net233;
 wire net234;
 wire net235;
 wire net236;
 wire net237;
 wire net238;
 wire net239;
 wire net240;
 wire net241;
 wire net242;
 wire net243;
 wire net244;
 wire net245;
 wire net246;
 wire net247;
 wire net248;
 wire net249;
 wire net250;
 wire net251;
 wire net252;
 wire net253;
 wire net254;
 wire net255;
 wire net256;
 wire net257;
 wire net258;
 wire net259;
 wire net260;
 wire net261;
 wire net262;
 wire net263;
 wire net264;
 wire net265;
 wire net266;
 wire net267;
 wire net268;
 wire net269;
 wire net270;
 wire net271;
 wire net272;
 wire net273;
 wire net274;
 wire net275;
 wire net276;
 wire net277;
 wire net278;
 wire net279;
 wire net280;
 wire net281;
 wire net282;
 wire net283;
 wire net284;
 wire net285;
 wire net286;
 wire net287;
 wire net288;
 wire net289;
 wire net290;
 wire net291;
 wire net292;
 wire net293;
 wire net294;
 wire net295;
 wire net296;
 wire net297;
 wire net298;
 wire net299;
 wire net300;
 wire net301;
 wire net302;
 wire net303;
 wire net304;
 wire net305;
 wire net306;
 wire net307;
 wire net308;
 wire net309;
 wire net310;
 wire net311;
 wire net312;
 wire net313;
 wire net314;
 wire net315;
 wire net316;
 wire net317;
 wire net318;
 wire net319;
 wire net320;
 wire net321;
 wire net322;
 wire net323;
 wire net324;
 wire net325;
 wire net326;
 wire net327;
 wire net328;
 wire net329;
 wire net330;
 wire net331;
 wire net332;
 wire net333;
 wire net334;
 wire net335;
 wire net336;
 wire net337;
 wire net338;
 wire net339;
 wire net340;
 wire net341;
 wire net342;
 wire net343;
 wire net344;
 wire net345;
 wire net346;
 wire net347;
 wire net348;
 wire net349;
 wire net350;
 wire net351;
 wire net352;
 wire net353;
 wire net354;
 wire net355;
 wire net356;
 wire net357;
 wire net358;
 wire net359;
 wire net360;
 wire net361;
 wire net362;
 wire net363;
 wire net364;
 wire net365;
 wire net366;
 wire net367;
 wire net368;
 wire net369;
 wire net370;
 wire net371;
 wire net372;
 wire net373;
 wire net374;
 wire net375;
 wire net376;
 wire net377;
 wire net378;
 wire net379;
 wire net380;
 wire net381;
 wire net382;
 wire net383;
 wire net384;
 wire net385;
 wire net386;
 wire net387;
 wire net388;
 wire net389;
 wire net390;
 wire net391;
 wire net392;
 wire net393;
 wire net394;
 wire net395;
 wire net396;
 wire net397;
 wire net398;
 wire net399;
 wire net400;
 wire net401;
 wire net402;
 wire net403;
 wire net404;
 wire net405;
 wire net406;
 wire net407;
 wire net408;
 wire net409;
 wire net410;
 wire net411;
 wire net412;
 wire net413;
 wire net414;
 wire net415;
 wire net416;
 wire net417;
 wire net418;
 wire net419;
 wire net420;
 wire net421;
 wire net422;
 wire net423;
 wire net424;
 wire net425;
 wire net426;
 wire net427;
 wire net428;
 wire net429;
 wire net430;
 wire net431;
 wire net432;
 wire net433;
 wire net434;
 wire net435;
 wire net436;
 wire net437;
 wire net438;
 wire net439;
 wire net440;
 wire net441;
 wire net442;
 wire net443;
 wire net444;
 wire net445;
 wire net446;
 wire net447;
 wire net448;
 wire net449;
 wire net450;
 wire net451;
 wire net452;
 wire net453;
 wire net454;
 wire net455;
 wire net456;
 wire net457;
 wire net458;
 wire net459;
 wire net460;
 wire net461;
 wire net462;
 wire net463;
 wire net464;
 wire net465;
 wire net466;
 wire net467;
 wire net468;
 wire net469;
 wire net470;
 wire net471;
 wire net472;
 wire net473;
 wire net474;
 wire net475;
 wire net476;
 wire net477;
 wire net478;
 wire net479;
 wire net480;
 wire net481;
 wire net482;
 wire net483;
 wire net484;
 wire net485;
 wire net486;
 wire net487;
 wire net488;
 wire net489;
 wire net490;
 wire net491;
 wire net492;
 wire net493;
 wire net494;
 wire net495;
 wire net496;
 wire net497;
 wire net498;
 wire net499;
 wire net500;
 wire net501;
 wire net502;
 wire net503;
 wire net504;
 wire net505;
 wire net506;
 wire net507;
 wire net508;
 wire net509;
 wire net510;
 wire net511;
 wire net512;
 wire net513;
 wire net514;
 wire net515;
 wire net516;
 wire net517;
 wire net518;
 wire net519;
 wire net520;
 wire net521;
 wire net522;
 wire net523;
 wire net524;
 wire net525;
 wire net526;
 wire net527;
 wire net528;
 wire net529;
 wire net530;
 wire net531;
 wire net532;
 wire net533;
 wire net534;
 wire net535;
 wire net536;
 wire net537;
 wire net538;
 wire net539;
 wire net540;
 wire net541;
 wire net542;
 wire net543;
 wire net544;
 wire net545;
 wire net546;
 wire net547;
 wire net548;
 wire net549;
 wire net550;
 wire net551;
 wire net552;
 wire net553;
 wire net554;
 wire net555;
 wire net556;
 wire net557;
 wire net558;
 wire net559;
 wire net560;
 wire net561;
 wire net562;
 wire net563;
 wire net564;
 wire net565;
 wire net566;
 wire net567;
 wire net568;
 wire net569;
 wire net570;
 wire net571;
 wire net572;
 wire net573;
 wire net574;
 wire net575;
 wire net576;
 wire net577;
 wire net578;
 wire net579;
 wire net580;
 wire net581;
 wire net582;
 wire net583;
 wire net584;
 wire net585;
 wire net586;
 wire net587;
 wire net588;
 wire net589;
 wire net590;
 wire net591;
 wire net592;
 wire net593;
 wire net594;
 wire net595;
 wire net596;
 wire net597;
 wire net598;
 wire net599;
 wire net600;
 wire net601;
 wire net602;
 wire net603;
 wire net604;
 wire net605;
 wire net606;
 wire net607;
 wire net608;
 wire net609;
 wire net610;
 wire net611;
 wire net612;
 wire net613;
 wire net614;
 wire net615;
 wire net616;
 wire net617;
 wire net618;
 wire net619;
 wire net620;
 wire net621;
 wire net622;
 wire net623;
 wire net624;
 wire net625;
 wire net626;
 wire net627;
 wire net628;
 wire net629;
 wire net630;
 wire net631;
 wire net632;
 wire net633;
 wire net634;
 wire net635;
 wire net636;
 wire net637;
 wire net638;
 wire net639;
 wire net640;
 wire net641;
 wire net642;
 wire net643;
 wire net644;
 wire net645;
 wire net646;
 wire net647;
 wire net648;
 wire net649;
 wire net650;
 wire net651;
 wire net652;
 wire net653;
 wire net654;
 wire net655;
 wire net656;
 wire net657;
 wire net658;
 wire net659;
 wire net660;
 wire net661;
 wire net662;
 wire net663;
 wire net664;
 wire net665;
 wire net666;
 wire net667;
 wire net668;
 wire net669;
 wire net670;
 wire net671;
 wire net672;
 wire net673;
 wire net674;
 wire net675;
 wire net676;
 wire net677;
 wire net678;
 wire net679;
 wire net680;
 wire net681;
 wire net682;
 wire net683;
 wire net684;
 wire net685;
 wire net686;
 wire net687;
 wire net688;
 wire net689;
 wire net690;
 wire net691;
 wire net692;
 wire net693;
 wire net694;
 wire net695;
 wire net696;
 wire net697;
 wire net698;
 wire net699;
 wire net700;
 wire net701;
 wire net702;
 wire net703;
 wire net704;
 wire net705;
 wire net706;
 wire net707;
 wire net708;
 wire net709;
 wire net710;
 wire net711;
 wire net712;
 wire net713;
 wire net714;
 wire net715;
 wire net716;
 wire net717;
 wire net718;
 wire net719;
 wire net720;
 wire net721;
 wire net722;
 wire net723;
 wire net724;
 wire net725;
 wire net726;
 wire net727;
 wire net728;
 wire net729;
 wire net730;
 wire net731;
 wire net732;
 wire net733;
 wire net734;
 wire net735;
 wire net736;
 wire net737;
 wire net738;
 wire net739;
 wire net740;
 wire net741;
 wire net742;
 wire net743;
 wire net744;
 wire net745;
 wire net746;
 wire net747;
 wire net748;
 wire net749;
 wire net750;
 wire net751;
 wire net752;
 wire net753;
 wire net754;
 wire net755;
 wire net756;
 wire net757;
 wire net758;
 wire net759;
 wire net760;
 wire net761;
 wire net762;
 wire net763;
 wire net764;
 wire net765;
 wire net766;
 wire net767;
 wire net768;
 wire net769;
 wire net770;
 wire net771;
 wire net772;
 wire net773;
 wire net774;
 wire net775;
 wire net776;
 wire net777;
 wire net778;
 wire net779;
 wire net780;
 wire net781;
 wire net782;
 wire net783;
 wire net784;
 wire net785;
 wire net786;
 wire net787;
 wire net788;
 wire net789;
 wire net790;
 wire net791;
 wire net792;
 wire net793;
 wire net794;
 wire net795;
 wire net796;
 wire net797;
 wire net798;
 wire net799;
 wire net800;
 wire net801;
 wire net802;
 wire net803;
 wire net804;
 wire net805;
 wire net806;
 wire net807;
 wire net808;
 wire net809;
 wire net810;
 wire net811;
 wire net812;
 wire net813;
 wire net814;
 wire net815;
 wire net816;
 wire net817;
 wire net818;
 wire net819;
 wire net820;
 wire net821;
 wire net822;
 wire net823;
 wire net824;
 wire net825;
 wire net826;
 wire net827;
 wire net828;
 wire net829;
 wire net830;
 wire net831;
 wire net832;
 wire net833;
 wire net834;
 wire net835;
 wire net836;
 wire net837;
 wire net838;
 wire net839;
 wire net840;
 wire net841;
 wire net842;
 wire net843;
 wire net844;
 wire net845;
 wire net846;
 wire net847;
 wire net848;
 wire net849;
 wire net850;
 wire net851;
 wire net852;
 wire net853;
 wire net854;
 wire net855;
 wire net856;
 wire net857;
 wire net858;
 wire net859;
 wire net860;
 wire net861;
 wire net862;
 wire net863;
 wire net864;
 wire net865;
 wire net866;
 wire net867;
 wire net868;
 wire net869;
 wire net870;
 wire net871;
 wire net872;
 wire net873;
 wire net874;
 wire net875;
 wire net876;
 wire net877;
 wire net878;
 wire net879;
 wire net880;
 wire net881;
 wire net882;
 wire net883;
 wire net884;
 wire net885;
 wire net886;
 wire net887;
 wire net888;
 wire net889;
 wire net890;
 wire net891;
 wire net892;
 wire net893;
 wire net894;
 wire net895;
 wire net896;
 wire net897;
 wire net898;
 wire net899;
 wire net900;
 wire net901;
 wire net902;
 wire net903;
 wire net904;
 wire net905;
 wire net906;
 wire net907;
 wire net908;
 wire net909;
 wire net910;
 wire net911;
 wire net912;
 wire net913;
 wire net914;
 wire net915;
 wire net916;
 wire net917;
 wire net918;
 wire net919;
 wire net920;
 wire net921;
 wire net922;
 wire net923;
 wire net924;
 wire net925;
 wire net926;
 wire net927;
 wire net928;
 wire net929;
 wire net930;
 wire net931;
 wire net932;
 wire net933;
 wire net934;
 wire net935;
 wire net936;
 wire net937;
 wire net938;
 wire net939;
 wire net940;
 wire net941;
 wire net942;
 wire net943;
 wire net944;
 wire net945;
 wire net946;
 wire net947;
 wire net948;
 wire net949;
 wire net950;
 wire net951;
 wire net952;
 wire net953;
 wire net954;
 wire net955;
 wire net956;
 wire net957;
 wire net958;
 wire net959;
 wire net960;
 wire net961;
 wire net962;
 wire net963;
 wire net964;
 wire net965;
 wire net966;
 wire net967;
 wire net968;
 wire net969;
 wire net970;
 wire net971;
 wire net972;
 wire net973;
 wire net974;
 wire net975;
 wire net976;
 wire net977;
 wire net978;
 wire net979;
 wire net980;
 wire net981;
 wire net982;
 wire net983;
 wire net984;
 wire net985;
 wire net986;
 wire net987;
 wire net988;
 wire net989;
 wire net990;
 wire net991;
 wire net992;
 wire net993;
 wire net994;
 wire net995;
 wire net996;
 wire net997;
 wire net998;
 wire net999;
 wire net1000;
 wire net1001;
 wire net1002;
 wire net1003;
 wire net1004;
 wire net1005;
 wire net1006;
 wire net1007;
 wire net1008;
 wire net1009;
 wire net1010;
 wire net1011;
 wire net1012;
 wire net1013;
 wire net1014;
 wire net1015;
 wire net1016;
 wire net1017;
 wire net1018;
 wire net1019;
 wire net1020;
 wire net1021;
 wire net1022;
 wire net1023;
 wire net1024;
 wire net1025;
 wire net1026;
 wire net1027;
 wire net1028;
 wire net1029;
 wire net1030;
 wire net1031;
 wire net1032;
 wire net1033;
 wire net1034;
 wire net1035;
 wire net1036;
 wire net1037;
 wire net1038;
 wire net1039;
 wire net1040;
 wire net1041;
 wire net1042;
 wire net1043;
 wire net1044;
 wire net1045;
 wire net1046;
 wire net1047;
 wire net1048;
 wire net1049;
 wire net1050;
 wire net1051;
 wire net1052;
 wire net1053;
 wire net1054;
 wire net1055;
 wire net1056;
 wire net1057;
 wire net1058;
 wire net1059;
 wire net1060;
 wire net1061;
 wire net1062;
 wire net1063;
 wire net1064;
 wire net1065;
 wire net1066;
 wire net1067;
 wire net1068;
 wire net1069;
 wire net1070;
 wire net1071;
 wire net1072;
 wire net1073;
 wire net1074;
 wire net1075;
 wire net1076;
 wire net1077;
 wire net1078;
 wire net1079;
 wire net1080;
 wire net1081;
 wire net1082;
 wire net1083;
 wire net1084;
 wire net1085;
 wire net1086;
 wire net1087;
 wire net1088;
 wire net1089;
 wire net1090;
 wire net1091;
 wire net1092;
 wire net1093;
 wire net1094;
 wire net1095;
 wire net1096;
 wire net1097;
 wire net1098;
 wire net1099;
 wire net1100;
 wire net1101;
 wire net1102;
 wire net1103;
 wire net1104;
 wire net1105;
 wire net1106;
 wire net1107;
 wire net1108;
 wire net1109;
 wire net1110;
 wire net1111;
 wire net1112;
 wire net1113;
 wire net1114;
 wire net1115;
 wire net1116;
 wire net1117;
 wire net1118;
 wire net1119;
 wire net1120;
 wire net1121;
 wire net1122;
 wire net1123;
 wire net1124;
 wire net1125;
 wire net1126;
 wire net1127;
 wire net1128;
 wire net1129;
 wire net1130;
 wire net1131;
 wire net1132;
 wire net1133;
 wire net1134;
 wire net1135;
 wire net1136;
 wire net1137;
 wire net1138;
 wire net1139;
 wire net1140;
 wire net1141;
 wire net1142;
 wire net1143;
 wire net1144;
 wire net1145;
 wire net1146;
 wire net1147;
 wire net1148;
 wire net1149;
 wire net1150;
 wire net1151;
 wire net1152;
 wire net1153;
 wire net1154;
 wire net1155;
 wire net1156;
 wire net1157;
 wire net1158;
 wire net1159;
 wire net1160;
 wire net1161;
 wire net1162;
 wire net1163;
 wire net1164;
 wire net1165;
 wire net1166;
 wire net1167;
 wire net1168;
 wire net1169;
 wire net1170;
 wire net1171;
 wire net1172;
 wire net1173;
 wire net1174;
 wire net1175;
 wire net1176;
 wire net1177;
 wire net1178;
 wire net1179;
 wire net1180;
 wire net1181;
 wire net1182;
 wire net1183;
 wire net1184;
 wire net1185;
 wire net1186;
 wire net1187;
 wire net1188;
 wire net1189;
 wire net1190;
 wire net1191;
 wire net1192;
 wire net1193;
 wire net1194;
 wire net1195;
 wire net1196;
 wire net1197;
 wire net1198;
 wire net1199;
 wire net1200;
 wire net1201;
 wire net1202;
 wire net1203;
 wire net1204;
 wire net1205;
 wire net1206;
 wire net1207;
 wire net1208;
 wire net1209;
 wire net1210;
 wire net1211;
 wire net1212;
 wire net1213;
 wire net1214;
 wire net1215;
 wire net1216;
 wire net1217;
 wire net1218;
 wire net1219;
 wire net1220;
 wire net1221;
 wire net1222;
 wire net1223;
 wire net1224;
 wire net1225;
 wire net1226;
 wire net1227;
 wire net1228;
 wire net1229;
 wire net1230;
 wire net1231;
 wire net1232;
 wire net1233;
 wire net1234;
 wire net1235;
 wire net1236;
 wire net1237;
 wire net1238;
 wire net1239;
 wire net1240;
 wire net1241;
 wire net1242;
 wire net1243;
 wire net1244;
 wire net1245;
 wire net1246;
 wire net1247;
 wire net1248;
 wire net1249;
 wire net1250;
 wire net1251;
 wire net1252;
 wire net1253;
 wire net1254;
 wire net1255;
 wire net1256;
 wire net1257;
 wire net1258;
 wire net1259;
 wire net1260;
 wire net1261;
 wire net1262;
 wire net1263;
 wire net1264;
 wire net1265;
 wire net1266;
 wire net1267;
 wire net1268;
 wire net1269;
 wire net1270;
 wire net1271;
 wire net1272;
 wire net1273;
 wire net1274;
 wire net1275;
 wire net1276;
 wire net1277;
 wire net1278;
 wire net1279;
 wire net1280;
 wire net1281;
 wire net1282;
 wire net1283;
 wire net1284;
 wire net1285;
 wire net1286;
 wire net1287;
 wire net1288;
 wire net1289;
 wire net1290;
 wire net1291;
 wire net1292;
 wire net1293;
 wire net1294;
 wire net1295;
 wire net1296;
 wire net1297;
 wire net1298;
 wire net1299;
 wire net1300;
 wire net1301;
 wire net1302;
 wire net1303;
 wire net1304;
 wire net1305;
 wire net1306;
 wire net1307;
 wire net1308;
 wire net1309;
 wire net1310;
 wire net1311;
 wire net1312;
 wire net1313;
 wire net1314;
 wire net1315;
 wire net1316;
 wire net1317;
 wire net1318;
 wire net1319;
 wire net1320;
 wire net1321;
 wire net1322;
 wire net1323;
 wire net1324;
 wire net1325;
 wire net1326;
 wire net1327;
 wire net1328;
 wire net1329;
 wire net1330;
 wire net1331;
 wire net1332;
 wire net1333;
 wire net1334;
 wire net1335;
 wire net1336;
 wire net1337;
 wire net1338;
 wire net1339;
 wire net1340;
 wire net1341;
 wire net1342;
 wire net1343;
 wire net1344;
 wire net1345;
 wire net1346;
 wire net1347;
 wire net1348;
 wire net1349;
 wire net1350;
 wire net1351;
 wire net1352;
 wire net1353;
 wire net1354;
 wire net1355;
 wire net1356;
 wire net1357;
 wire net1358;
 wire net1359;
 wire net1360;
 wire net1361;
 wire net1362;
 wire net1363;
 wire net1364;
 wire net1365;
 wire net1366;
 wire net1367;
 wire net1368;
 wire net1369;
 wire net1370;
 wire net1371;
 wire net1372;
 wire net1373;
 wire net1374;
 wire net1375;
 wire net1376;
 wire net1377;
 wire net1378;
 wire net1379;
 wire net1380;
 wire net1381;
 wire net1382;
 wire net1383;
 wire net1384;
 wire net1385;
 wire net1386;
 wire net1387;
 wire net1388;
 wire net1389;
 wire net1390;
 wire net1391;
 wire net1392;
 wire net1393;
 wire net1394;
 wire net1395;
 wire net1396;
 wire net1397;
 wire net1398;
 wire net1399;
 wire net1400;
 wire net1401;
 wire net1402;
 wire net1403;
 wire net1404;
 wire net1405;
 wire net1406;
 wire net1407;
 wire net1408;
 wire net1409;
 wire net1410;
 wire net1411;
 wire net1412;
 wire net1413;
 wire net1414;
 wire net1415;
 wire net1416;
 wire net1417;
 wire net1418;
 wire net1419;
 wire net1420;
 wire net1421;
 wire net1422;
 wire net1423;
 wire net1424;
 wire net1425;
 wire net1426;
 wire net1427;
 wire net1428;
 wire net1429;
 wire net1430;
 wire net1431;
 wire net1432;
 wire net1433;
 wire net1434;
 wire net1435;
 wire net1436;
 wire net1437;
 wire net1438;
 wire net1439;
 wire net1440;
 wire net1441;
 wire net1442;
 wire net1443;
 wire net1444;
 wire net1445;
 wire net1446;
 wire net1447;
 wire net1448;
 wire net1449;
 wire net1450;
 wire net1451;
 wire net1452;
 wire net1453;
 wire net1454;
 wire net1455;
 wire net1456;
 wire net1457;
 wire net1458;
 wire net1459;
 wire net1460;
 wire net1461;
 wire net1462;
 wire net1463;
 wire net1464;
 wire net1465;
 wire net1466;
 wire net1467;
 wire net1468;
 wire net1469;
 wire net1470;
 wire net1471;
 wire net1472;
 wire net1473;
 wire net1474;
 wire net1475;
 wire net1476;
 wire net1477;
 wire net1478;
 wire net1479;
 wire net1480;
 wire net1481;
 wire net1482;
 wire net1483;
 wire net1484;
 wire net1485;
 wire net1486;
 wire net1487;
 wire net1488;
 wire net1489;
 wire net1490;
 wire net1491;
 wire net1492;
 wire net1493;
 wire net1494;
 wire net1495;
 wire net1496;
 wire net1497;
 wire net1498;
 wire net1499;
 wire net1500;
 wire net1501;
 wire net1502;
 wire net1503;
 wire net1504;
 wire net1505;
 wire net1506;
 wire net1507;
 wire net1508;
 wire net1509;
 wire net1510;
 wire net1511;
 wire net1512;
 wire net1513;
 wire net1514;
 wire net1515;
 wire net1516;
 wire net1517;
 wire net1518;
 wire net1519;
 wire net1520;
 wire net1521;
 wire net1522;
 wire net1523;
 wire net1524;
 wire net1525;
 wire net1526;
 wire net1527;
 wire net1528;
 wire net1529;
 wire net1530;
 wire net1531;
 wire net1532;
 wire net1533;
 wire net1534;
 wire net1535;
 wire net1536;
 wire net1537;
 wire net1538;
 wire net1539;
 wire net1540;
 wire net1541;
 wire net1542;
 wire net1543;
 wire net1544;
 wire net1545;
 wire net1546;
 wire net1547;
 wire net1548;
 wire net1549;
 wire net1550;
 wire net1551;
 wire net1552;
 wire net1553;
 wire net1554;
 wire net1555;
 wire net1556;
 wire net1557;
 wire net1558;
 wire net1559;
 wire net1560;
 wire net1561;
 wire net1562;
 wire net1563;
 wire net1564;
 wire net1565;
 wire net1566;
 wire net1567;
 wire net1568;
 wire net1569;
 wire net1570;
 wire net1571;
 wire net1572;
 wire net1573;
 wire net1574;
 wire net1575;
 wire net1576;
 wire net1577;
 wire net1578;
 wire net1579;
 wire net1580;
 wire net1581;
 wire net1582;
 wire net1583;
 wire net1584;
 wire net1585;
 wire net1586;
 wire net1587;
 wire net1588;
 wire net1589;
 wire net1590;
 wire net1591;
 wire net1592;
 wire net1593;
 wire net1594;
 wire net1595;
 wire net1596;
 wire net1597;
 wire net1598;
 wire net1599;
 wire net1600;
 wire net1601;
 wire net1602;
 wire net1603;
 wire net1604;
 wire net1605;
 wire net1606;
 wire net1607;
 wire net1608;
 wire net1609;
 wire net1610;
 wire net1611;
 wire net1612;
 wire net1613;
 wire net1614;
 wire net1615;
 wire net1616;
 wire net1617;
 wire net1618;
 wire net1619;
 wire net1620;
 wire net1621;
 wire net1622;
 wire net1623;
 wire net1624;
 wire net1625;
 wire net1626;
 wire net1627;
 wire net1628;
 wire net1629;
 wire net1630;
 wire net1631;
 wire net1632;
 wire net1633;
 wire net1634;
 wire net1635;
 wire net1636;
 wire net1637;
 wire net1638;
 wire net1639;
 wire net1640;
 wire net1641;
 wire net1642;
 wire net1643;
 wire net1644;
 wire net1645;
 wire net1646;
 wire net1647;
 wire net1648;
 wire net1649;
 wire net1650;
 wire net1651;
 wire net1652;
 wire net1653;
 wire net1654;
 wire net1655;
 wire net1656;
 wire net1657;
 wire net1658;
 wire net1659;
 wire net1660;
 wire net1661;
 wire net1662;
 wire net1663;
 wire net1664;
 wire net1665;
 wire net1666;
 wire net1667;
 wire net1668;
 wire net1669;
 wire net1670;
 wire net1671;
 wire net1672;
 wire net1673;
 wire net1674;
 wire net1675;
 wire net1676;
 wire net1677;
 wire net1678;
 wire net1679;
 wire net1680;
 wire net1681;
 wire net1682;
 wire net1683;
 wire net1684;
 wire net1685;
 wire net1686;
 wire net1687;
 wire net1688;
 wire net1689;
 wire net1690;
 wire net1691;
 wire net1692;
 wire net1693;
 wire net1694;
 wire net1695;
 wire net1696;
 wire net1697;
 wire net1698;
 wire net1699;
 wire net1700;
 wire net1701;
 wire net1702;
 wire net1703;
 wire net1704;
 wire net1705;
 wire net1706;
 wire net1707;
 wire net1708;
 wire net1709;
 wire net1710;
 wire net1711;
 wire net1712;
 wire net1713;
 wire net1714;
 wire net1715;
 wire net1716;
 wire net1717;
 wire net1718;
 wire net1719;
 wire net1720;
 wire net1721;
 wire net1722;
 wire net1723;
 wire net1724;
 wire net1725;
 wire net1726;
 wire net1727;
 wire net1728;
 wire net1729;
 wire net1730;
 wire net1731;
 wire net1732;
 wire net1733;
 wire net1734;
 wire net1735;
 wire net1736;
 wire net1737;
 wire net1738;
 wire net1739;
 wire net1740;
 wire net1741;
 wire net1742;
 wire net1743;
 wire net1744;
 wire net1745;
 wire net1746;
 wire net1747;
 wire net1748;
 wire net1749;
 wire net1750;
 wire net1751;
 wire net1752;
 wire net1753;
 wire net1754;
 wire net1755;
 wire net1756;
 wire net1757;
 wire net1758;
 wire net1759;
 wire net1760;
 wire net1761;
 wire net1762;
 wire net1763;
 wire net1764;
 wire net1765;
 wire net1766;
 wire net1767;
 wire net1768;
 wire net1769;
 wire net1770;
 wire net1771;
 wire net1772;
 wire net1773;
 wire net1774;
 wire net1775;
 wire net1776;
 wire net1777;
 wire net1778;
 wire net1779;
 wire net1780;
 wire net1781;
 wire net1782;
 wire net1783;
 wire net1784;
 wire net1785;
 wire net1786;
 wire net1787;
 wire net1788;
 wire net1789;
 wire net1790;
 wire net1791;
 wire net1792;
 wire net1793;
 wire net1794;
 wire net1795;
 wire net1796;
 wire net1797;
 wire net1798;
 wire net1799;
 wire net1800;
 wire net1801;
 wire net1802;
 wire net1803;
 wire net1804;
 wire net1805;
 wire net1806;
 wire net1807;
 wire net1808;
 wire net1809;
 wire net1810;
 wire net1811;
 wire net1812;
 wire net1813;
 wire net1814;
 wire net1815;
 wire net1816;
 wire net1817;
 wire net1818;
 wire net1819;
 wire net1820;
 wire net1821;
 wire net1822;
 wire net1823;
 wire net1824;
 wire net1825;
 wire net1826;
 wire net1827;
 wire net1828;
 wire net1829;
 wire net1830;
 wire net1831;
 wire net1832;
 wire net1833;
 wire net1834;
 wire net1835;
 wire net1836;
 wire net1837;
 wire net1838;
 wire net1839;
 wire net1840;
 wire net1841;
 wire net1842;
 wire net1843;
 wire net1844;
 wire net1845;
 wire net1846;
 wire net1847;
 wire net1848;
 wire net1849;
 wire net1850;
 wire net1851;
 wire net1852;
 wire net1853;
 wire net1854;
 wire net1855;
 wire net1856;
 wire net1857;
 wire net1858;
 wire net1859;
 wire net1860;
 wire net1861;
 wire net1862;
 wire net1863;
 wire net1864;
 wire net1865;
 wire net1866;
 wire net1867;
 wire net1868;
 wire net1869;
 wire net1870;
 wire net1871;
 wire net1872;
 wire net1873;
 wire net1874;
 wire net1875;
 wire net1876;
 wire net1877;
 wire net1878;
 wire net1879;
 wire net1880;
 wire net1881;
 wire net1882;
 wire net1883;
 wire net1884;
 wire net1885;
 wire net1886;
 wire net1887;
 wire net1888;
 wire net1889;
 wire net1890;
 wire net1891;
 wire net1892;
 wire net1893;
 wire net1894;
 wire net1895;
 wire net1896;
 wire net1897;
 wire net1898;
 wire net1899;
 wire net1900;
 wire net1901;
 wire net1902;
 wire net1903;
 wire net1904;
 wire net1905;
 wire net1906;
 wire net1907;
 wire net1908;
 wire net1909;
 wire net1910;
 wire net1911;
 wire net1912;
 wire net1913;
 wire net1914;
 wire net1915;
 wire net1916;
 wire net1917;
 wire net1918;
 wire net1919;
 wire net1920;
 wire net1921;
 wire net1922;
 wire net1923;
 wire net1924;
 wire net1925;
 wire net1926;
 wire net1927;
 wire net1928;
 wire net1929;
 wire net1930;
 wire net1931;
 wire net1932;
 wire net1933;
 wire net1934;
 wire net1935;
 wire net1936;
 wire net1937;
 wire net1938;
 wire net1939;
 wire net1940;
 wire net1941;
 wire net1942;
 wire net1943;
 wire net1944;
 wire net1945;
 wire net1946;
 wire net1947;
 wire net1948;
 wire net1949;
 wire net1950;
 wire net1951;
 wire net1952;
 wire net1953;
 wire net1954;
 wire net1955;
 wire net1956;
 wire net1957;
 wire net1958;
 wire net1959;
 wire net1960;
 wire net1961;
 wire net1962;
 wire net1963;
 wire net1964;
 wire net1965;
 wire net1966;
 wire net1967;
 wire net1968;
 wire net1969;
 wire net1970;
 wire net1971;
 wire net1972;
 wire net1973;
 wire net1974;
 wire net1975;
 wire net1976;
 wire net1977;
 wire net1978;
 wire net1979;
 wire net1980;
 wire net1981;
 wire net1982;
 wire net1983;
 wire net1984;
 wire net1985;
 wire net1986;
 wire net1987;
 wire net1988;
 wire net1989;
 wire net1990;
 wire net1991;
 wire net1992;
 wire net1993;
 wire net1994;
 wire net1995;
 wire net1996;
 wire net1997;
 wire net1998;
 wire net1999;
 wire net2000;
 wire net2001;
 wire net2002;
 wire net2003;
 wire net2004;
 wire net2005;
 wire net2006;
 wire net2007;
 wire net2008;
 wire net2009;
 wire net2010;
 wire net2011;
 wire net2012;
 wire net2013;
 wire net2014;
 wire net2015;
 wire net2016;
 wire net2017;
 wire net2018;
 wire net2019;
 wire net2020;
 wire net2021;
 wire net2022;
 wire net2023;
 wire net2024;
 wire net2025;
 wire net2026;
 wire net2027;
 wire net2028;
 wire net2029;
 wire net2030;
 wire net2031;
 wire net2032;
 wire net2033;
 wire net2034;
 wire net2035;
 wire net2036;
 wire net2037;
 wire net2038;
 wire net2039;
 wire net2040;
 wire net2041;
 wire net2042;
 wire net2043;
 wire net2044;
 wire net2045;
 wire net2046;
 wire net2047;
 wire net2048;
 wire net2049;
 wire net2050;
 wire net2051;
 wire net2052;
 wire net2053;
 wire net2054;
 wire net2055;
 wire net2056;
 wire net2057;
 wire net2058;
 wire net2059;
 wire net2060;
 wire net2061;
 wire net2062;
 wire net2063;
 wire net2064;
 wire net2065;
 wire net2066;
 wire net2067;
 wire net2068;
 wire net2069;
 wire net2070;
 wire net2071;
 wire net2072;
 wire net2073;
 wire net2074;
 wire net2075;
 wire net2076;
 wire net2077;
 wire net2078;
 wire net2079;
 wire net2080;
 wire net2081;
 wire net2082;
 wire net2083;
 wire net2084;
 wire net2085;
 wire net2086;
 wire net2087;
 wire net2088;
 wire net2089;
 wire net2090;
 wire net2091;
 wire net2092;
 wire net2093;
 wire net2094;
 wire net2095;
 wire net2096;
 wire net2097;
 wire net2098;
 wire net2099;
 wire net2100;
 wire net2101;
 wire net2102;
 wire net2103;
 wire net2104;
 wire net2105;
 wire net2106;
 wire net2107;
 wire net2108;
 wire net2109;
 wire net2110;
 wire net2111;
 wire net2112;
 wire net2113;
 wire net2114;
 wire net2115;
 wire net2116;
 wire net2117;
 wire net2118;
 wire net2119;
 wire net2120;
 wire net2121;
 wire net2122;
 wire net2123;
 wire net2124;
 wire net2125;
 wire net2126;
 wire net2127;
 wire net2128;
 wire net2129;
 wire net2130;
 wire net2131;
 wire net2132;
 wire net2133;
 wire net2134;
 wire net2135;
 wire net2136;
 wire net2137;
 wire net2138;
 wire net2139;
 wire net2140;
 wire net2141;
 wire net2142;
 wire net2143;
 wire net2144;
 wire net2145;
 wire net2146;
 wire net2147;
 wire net2148;
 wire net2149;
 wire net2150;
 wire net2151;
 wire net2152;
 wire net2153;
 wire net2154;
 wire net2155;
 wire net2156;
 wire net2157;
 wire net2158;
 wire net2159;
 wire net2160;
 wire net2161;
 wire net2162;
 wire net2163;
 wire net2164;
 wire net2165;
 wire net2166;
 wire net2167;
 wire net2168;
 wire net2169;
 wire net2170;
 wire net2171;
 wire net2172;
 wire net2173;
 wire net2174;
 wire net2175;
 wire net2176;
 wire net2177;
 wire net2178;
 wire net2179;
 wire net2180;
 wire net2181;
 wire net2182;
 wire net2183;
 wire net2184;
 wire net2185;
 wire net2186;
 wire net2187;
 wire net2188;
 wire net2189;
 wire net2190;
 wire net2191;
 wire net2192;
 wire net2193;
 wire net2194;
 wire net2195;
 wire net2196;
 wire net2197;
 wire net2198;
 wire net2199;
 wire net2200;
 wire net2201;
 wire net2202;
 wire net2203;
 wire net2204;
 wire net2205;
 wire net2206;
 wire net2207;
 wire net2208;
 wire net2209;
 wire net2210;
 wire net2211;
 wire net2212;
 wire net2213;
 wire net2214;
 wire net2215;
 wire net2216;
 wire net2217;
 wire net2218;
 wire net2219;
 wire net2220;
 wire net2221;
 wire net2222;
 wire net2223;
 wire net2224;
 wire net2225;
 wire net2226;
 wire net2227;
 wire net2228;
 wire net2229;
 wire net2230;
 wire net2231;
 wire net2232;
 wire net2233;
 wire net2234;
 wire net2235;
 wire net2236;
 wire net2237;
 wire net2238;
 wire net2239;
 wire net2240;
 wire net2241;
 wire net2242;
 wire net2243;
 wire net2244;
 wire net2245;
 wire net2246;
 wire net2247;
 wire net2248;
 wire net2249;
 wire net2250;
 wire net2251;
 wire net2252;
 wire net2253;
 wire net2254;
 wire net2255;
 wire net2256;
 wire net2257;
 wire net2258;
 wire net2259;
 wire net2260;
 wire net2261;
 wire net2262;
 wire net2263;
 wire net2264;
 wire net2265;
 wire net2266;
 wire net2267;
 wire net2268;
 wire net2269;
 wire net2270;
 wire net2271;
 wire net2272;
 wire net2273;
 wire net2274;
 wire net2275;
 wire net2276;
 wire net2277;
 wire net2278;
 wire net2279;
 wire net2280;
 wire net2281;
 wire net2282;
 wire net2283;
 wire net2284;
 wire net2285;
 wire net2286;
 wire net2287;
 wire net2288;
 wire net2289;
 wire net2290;
 wire net2291;
 wire net2292;
 wire net2293;
 wire net2294;
 wire net2295;
 wire net2296;
 wire net2297;
 wire net2298;
 wire net2299;
 wire net2300;
 wire net2301;
 wire net2302;
 wire net2303;
 wire net2304;
 wire net2305;
 wire net2306;
 wire net2307;
 wire net2308;
 wire net2309;
 wire net2310;
 wire net2311;
 wire net2312;
 wire net2313;
 wire net2314;
 wire net2315;
 wire net2316;
 wire net2317;
 wire net2318;
 wire net2319;
 wire net2320;
 wire net2321;
 wire net2322;
 wire net2323;
 wire net2324;
 wire net2325;
 wire net2326;
 wire net2327;
 wire net2328;
 wire net2329;
 wire net2330;
 wire net2331;
 wire net2332;
 wire net2333;
 wire net2334;
 wire net2335;
 wire net2336;
 wire net2337;
 wire net2338;
 wire net2339;
 wire net2340;
 wire net2341;
 wire net2342;
 wire net2343;
 wire net2344;
 wire net2345;
 wire net2346;
 wire net2347;
 wire net2348;
 wire net2349;
 wire net2350;
 wire net2351;
 wire net2352;
 wire net2353;
 wire net2354;
 wire net2355;
 wire net2356;
 wire net2357;
 wire net2358;
 wire net2359;
 wire net2360;
 wire net2361;
 wire net2362;
 wire net2363;
 wire net2364;
 wire net2365;
 wire net2366;
 wire net2367;
 wire net2368;
 wire net2369;
 wire net2370;
 wire net2371;
 wire net2372;
 wire net2373;
 wire net2374;
 wire net2375;
 wire net2376;
 wire net2377;
 wire net2378;
 wire net2379;
 wire net2380;
 wire net2381;
 wire net2382;
 wire net2383;
 wire net2384;
 wire net2385;
 wire net2386;
 wire net2387;
 wire net2388;
 wire net2389;
 wire net2390;
 wire net2391;
 wire net2392;
 wire net2393;
 wire net2394;
 wire net2395;
 wire net2396;
 wire net2397;
 wire net2398;
 wire net2399;
 wire net2400;
 wire net2401;
 wire net2402;
 wire net2403;
 wire net2404;
 wire net2405;
 wire net2406;
 wire net2407;
 wire net2408;
 wire net2409;
 wire net2410;
 wire net2411;
 wire net2412;
 wire net2413;
 wire net2414;
 wire net2415;
 wire net2416;
 wire net2417;
 wire net2418;
 wire net2419;
 wire net2420;
 wire net2421;
 wire net2422;
 wire net2423;
 wire net2424;
 wire net2425;
 wire net2426;
 wire net2427;
 wire net2428;
 wire net2429;
 wire net2430;
 wire net2431;
 wire net2432;
 wire net2433;
 wire net2434;
 wire net2435;
 wire net2436;
 wire net2437;
 wire net2438;
 wire net2439;
 wire net2440;
 wire net2441;
 wire net2442;
 wire net2443;
 wire net2444;
 wire net2445;
 wire net2446;
 wire net2447;
 wire net2448;
 wire net2449;
 wire net2450;
 wire net2451;
 wire net2452;
 wire net2453;
 wire net2454;
 wire net2455;
 wire net2456;
 wire net2457;
 wire net2458;
 wire net2459;
 wire net2460;
 wire net2461;
 wire net2462;
 wire net2463;
 wire net2464;
 wire net2465;
 wire net2466;
 wire net2467;
 wire net2468;
 wire net2469;
 wire net2470;
 wire net2471;
 wire net2472;
 wire net2473;
 wire net2474;
 wire net2475;
 wire net2476;
 wire net2477;
 wire net2478;
 wire net2479;
 wire net2480;
 wire net2481;
 wire net2482;
 wire net2483;
 wire net2484;
 wire net2485;
 wire net2486;
 wire net2487;
 wire net2488;
 wire net2489;
 wire net2490;
 wire net2491;
 wire net2492;
 wire net2493;
 wire net2494;
 wire net2495;
 wire net2496;
 wire net2497;
 wire net2498;
 wire net2499;
 wire net2500;
 wire net2501;
 wire net2502;
 wire net2503;
 wire net2504;
 wire net2505;
 wire net2506;
 wire net2507;
 wire net2508;
 wire net2509;
 wire net2510;
 wire net2511;
 wire net2512;
 wire net2513;
 wire net2514;
 wire net2515;
 wire net2516;
 wire net2517;
 wire net2518;
 wire net2519;
 wire net2520;
 wire net2521;
 wire net2522;
 wire net2523;
 wire net2524;
 wire net2525;
 wire net2526;
 wire net2527;
 wire net2528;
 wire net2529;
 wire net2530;
 wire net2531;
 wire net2532;
 wire net2533;
 wire net2534;
 wire net2535;
 wire net2536;
 wire net2537;
 wire net2538;
 wire net2539;
 wire net2540;
 wire net2541;
 wire net2542;
 wire net2543;
 wire net2544;
 wire net2545;
 wire net2546;
 wire net2547;
 wire net2548;
 wire net2549;
 wire net2550;
 wire net2551;
 wire net2552;
 wire net2553;
 wire net2554;
 wire net2555;
 wire net2556;
 wire net2557;
 wire net2558;
 wire net2559;
 wire net2560;
 wire net2561;
 wire net2562;
 wire net2563;
 wire net2564;
 wire net2565;
 wire net2566;
 wire net2567;
 wire net2568;
 wire net2569;
 wire net2570;
 wire net2571;
 wire net2572;
 wire net2573;
 wire net2574;
 wire net2575;
 wire net2576;
 wire net2577;
 wire net2578;
 wire net2579;
 wire net2580;
 wire net2581;
 wire net2582;
 wire net2583;
 wire net2584;
 wire net2585;
 wire net2586;
 wire net2587;
 wire net2588;
 wire net2589;
 wire net2590;
 wire net2591;
 wire net2592;
 wire net2593;
 wire net2594;
 wire net2595;
 wire net2596;
 wire net2597;
 wire net2598;
 wire net2599;
 wire net2600;
 wire net2601;
 wire net2602;
 wire net2603;
 wire net2604;
 wire net2605;
 wire net2606;
 wire net2607;
 wire net2608;
 wire net2609;
 wire net2610;
 wire net2611;
 wire net2612;
 wire net2613;
 wire net2614;
 wire net2615;
 wire net2616;
 wire net2617;
 wire net2618;
 wire net2619;
 wire net2620;
 wire net2621;
 wire net2622;
 wire net2623;
 wire net2624;
 wire net2625;
 wire net2626;
 wire net2627;
 wire net2628;
 wire net2629;
 wire net2630;
 wire net2631;
 wire net2632;
 wire net2633;
 wire net2634;
 wire net2635;
 wire net2636;
 wire net2637;
 wire net2638;
 wire net2639;
 wire net2640;
 wire net2641;
 wire net2642;
 wire net2643;
 wire net2644;
 wire net2645;
 wire net2646;
 wire net2647;
 wire net2648;
 wire net2649;
 wire net2650;
 wire net2651;
 wire net2652;
 wire net2653;
 wire net2654;
 wire net2655;
 wire net2656;
 wire net2657;
 wire net2658;
 wire net2659;
 wire net2660;
 wire net2661;
 wire net2662;
 wire net2663;
 wire net2664;
 wire net2665;
 wire net2666;
 wire net2667;
 wire net2668;
 wire net2669;
 wire net2670;
 wire net2671;
 wire net2672;
 wire net2673;
 wire net2674;
 wire net2675;
 wire net2676;
 wire net2677;
 wire net2678;
 wire net2679;
 wire net2680;
 wire net2681;
 wire net2682;
 wire net2683;
 wire net2684;
 wire net2685;
 wire net2686;
 wire net2687;
 wire net2688;
 wire net2689;
 wire net2690;
 wire net2691;
 wire net2692;
 wire net2693;
 wire net2694;
 wire net2695;
 wire net2696;
 wire net2697;
 wire net2698;
 wire net2699;
 wire net2700;
 wire net2701;
 wire net2702;
 wire net2703;
 wire net2704;
 wire net2705;
 wire net2706;
 wire net2707;
 wire net2708;
 wire net2709;
 wire net2710;
 wire net2711;
 wire net2712;
 wire net2713;
 wire net2714;
 wire net2715;
 wire net2716;
 wire net2717;
 wire net2718;
 wire net2719;
 wire net2720;
 wire net2721;
 wire net2722;
 wire net2723;
 wire net2724;
 wire net2725;
 wire net2726;
 wire net2727;
 wire net2728;
 wire net2729;
 wire net2730;
 wire net2731;
 wire net2732;
 wire net2733;
 wire net2734;
 wire net2735;
 wire net2736;
 wire net2737;
 wire net2738;
 wire net2739;
 wire net2740;
 wire net2741;
 wire net2742;
 wire net2743;
 wire net2744;
 wire net2745;
 wire net2746;
 wire net2747;
 wire net2748;
 wire net2749;
 wire net2750;
 wire net2751;
 wire net2752;
 wire net2753;
 wire net2754;
 wire net2755;
 wire net2756;
 wire net2757;
 wire net2758;
 wire net2759;
 wire net2760;
 wire net2761;
 wire net2762;
 wire net2763;
 wire net2764;
 wire net2765;
 wire net2766;
 wire net2767;
 wire net2768;
 wire net2769;
 wire net2770;
 wire net2771;
 wire net2772;
 wire net2773;
 wire net2774;
 wire net2775;
 wire net2776;
 wire net2777;
 wire net2778;
 wire net2779;
 wire net2780;
 wire net2781;
 wire net2782;
 wire net2783;
 wire net2784;
 wire net2785;
 wire net2786;
 wire net2787;
 wire net2788;
 wire net2789;
 wire net2790;
 wire net2791;
 wire net2792;
 wire net2793;
 wire net2794;
 wire net2795;
 wire net2796;
 wire net2797;
 wire net2798;
 wire net2799;
 wire net2800;
 wire net2801;
 wire net2802;
 wire net2803;
 wire net2804;
 wire net2805;
 wire net2806;
 wire net2807;
 wire net2808;
 wire net2809;
 wire net2810;
 wire net2811;
 wire net2812;
 wire net2813;
 wire net2814;
 wire net2815;
 wire net2816;
 wire net2817;
 wire net2818;
 wire net2819;
 wire net2820;
 wire net2821;
 wire net2822;
 wire net2823;
 wire net2824;
 wire net2825;
 wire net2826;
 wire net2827;
 wire net2828;
 wire net2829;
 wire net2830;
 wire net2831;
 wire net2832;
 wire net2833;
 wire net2834;
 wire net2835;
 wire net2836;
 wire net2837;
 wire net2838;
 wire net2839;
 wire net2840;
 wire net2841;
 wire net2842;
 wire net2843;
 wire net2844;
 wire net2845;
 wire net2846;
 wire net2847;
 wire net2848;
 wire net2849;
 wire net2850;
 wire net2851;
 wire net2852;
 wire net2853;
 wire net2854;
 wire net2855;
 wire net2856;
 wire net2857;
 wire net2858;
 wire net2859;
 wire net2860;
 wire net2861;
 wire net2862;
 wire net2863;
 wire net2864;
 wire net2865;
 wire net2866;
 wire net2867;
 wire net2868;
 wire net2869;
 wire net2870;
 wire net2871;
 wire net2872;
 wire net2873;
 wire net2874;
 wire net2875;
 wire net2876;
 wire net2877;
 wire net2878;
 wire net2879;
 wire net2880;
 wire net2881;
 wire net2882;
 wire net2883;
 wire net2884;
 wire net2885;
 wire net2886;
 wire net2887;
 wire net2888;
 wire net2889;
 wire net2890;
 wire net2891;
 wire net2892;
 wire net2893;
 wire net2894;
 wire net2895;
 wire net2896;
 wire net2897;
 wire net2898;
 wire net2899;
 wire net2900;
 wire net2901;
 wire net2902;
 wire net2903;
 wire net2904;
 wire net2905;
 wire net2906;
 wire net2907;
 wire net2908;
 wire net2909;
 wire net2910;
 wire net2911;
 wire net2912;
 wire net2913;
 wire net2914;
 wire net2915;
 wire net2916;
 wire net2917;
 wire net2918;
 wire net2919;
 wire net2920;
 wire net2921;
 wire net2922;
 wire net2923;
 wire net2924;
 wire net2925;
 wire net2926;
 wire net2927;
 wire net2928;
 wire net2929;
 wire net2930;
 wire net2931;
 wire net2932;
 wire net2933;
 wire net2934;
 wire net2935;
 wire net2936;
 wire net2937;
 wire net2938;
 wire net2939;
 wire net2940;
 wire net2941;
 wire net2942;
 wire net2943;
 wire net2944;
 wire net2945;
 wire net2946;
 wire net2947;
 wire net2948;
 wire net2949;
 wire net2950;
 wire net2951;
 wire net2952;
 wire net2953;
 wire net2954;
 wire net2955;
 wire net2956;
 wire net2957;
 wire net2958;
 wire net2959;
 wire net2960;
 wire net2961;
 wire net2962;
 wire net2963;
 wire net2964;
 wire net2965;
 wire net2966;
 wire net2967;
 wire net2968;
 wire net2969;
 wire net2970;
 wire net2971;
 wire net2972;
 wire net2973;
 wire net2974;
 wire net2975;
 wire net2976;
 wire net2977;
 wire net2978;
 wire net2979;
 wire net2980;
 wire net2981;
 wire net2982;
 wire net2983;
 wire net2984;
 wire net2985;
 wire net2986;
 wire net2987;
 wire net2988;
 wire net2989;
 wire net2990;
 wire net2991;
 wire net2992;
 wire net2993;
 wire net2994;
 wire net2995;
 wire net2996;
 wire net2997;
 wire net2998;
 wire net2999;
 wire net3000;
 wire net3001;
 wire net3002;
 wire net3003;
 wire net3004;
 wire net3005;
 wire net3006;
 wire net3007;
 wire net3008;
 wire net3009;
 wire net3010;
 wire net3011;
 wire net3012;
 wire net3013;
 wire net3014;
 wire net3015;
 wire net3016;
 wire net3017;
 wire net3018;
 wire net3019;
 wire net3020;
 wire net3021;
 wire net3022;
 wire net3023;
 wire net3024;
 wire net3025;
 wire net3026;
 wire net3027;
 wire net3028;
 wire net3029;
 wire net3030;
 wire net3031;
 wire net3032;
 wire net3033;
 wire net3034;
 wire net3035;
 wire net3036;
 wire net3037;
 wire net3038;
 wire net3039;
 wire net3040;
 wire net3041;
 wire net3042;
 wire net3043;
 wire net3044;
 wire net3045;
 wire net3046;
 wire net3047;
 wire net3048;
 wire net3049;
 wire net3050;
 wire net3051;
 wire net3052;
 wire net3053;
 wire net3054;
 wire net3055;
 wire net3056;
 wire net3057;
 wire net3058;
 wire net3059;
 wire net3060;
 wire net3061;
 wire net3062;
 wire net3063;
 wire net3064;
 wire net3065;
 wire net3066;
 wire net3067;
 wire net3068;
 wire net3069;
 wire net3070;
 wire net3071;
 wire net3072;
 wire net3073;
 wire net3074;
 wire net3075;
 wire net3076;
 wire net3077;
 wire net3078;
 wire net3079;
 wire net3080;
 wire net3081;
 wire net3082;
 wire net3083;
 wire net3084;
 wire net3085;
 wire net3086;
 wire net3087;
 wire net3088;
 wire net3089;
 wire net3090;
 wire net3091;
 wire net3092;
 wire net3093;
 wire net3094;
 wire net3095;
 wire net3096;
 wire net3097;
 wire net3098;
 wire net3099;
 wire net3100;
 wire net3101;
 wire net3102;
 wire net3103;
 wire net3104;
 wire net3105;
 wire net3106;
 wire net3107;
 wire net3108;
 wire net3109;
 wire net3110;
 wire net3111;
 wire net3112;
 wire net3113;
 wire net3114;
 wire net3115;
 wire net3116;
 wire net3117;
 wire net3118;
 wire net3119;
 wire net3120;
 wire net3121;
 wire net3122;
 wire net3123;
 wire net3124;
 wire net3125;
 wire net3126;
 wire net3127;
 wire net3128;
 wire net3129;
 wire net3130;
 wire net3131;
 wire net3132;
 wire net3133;
 wire net3134;
 wire net3135;
 wire net3136;
 wire net3137;
 wire net3138;
 wire net3139;
 wire net3140;
 wire net3141;
 wire net3142;
 wire net3143;
 wire net3144;
 wire net3145;
 wire net3146;
 wire net3147;
 wire net3148;
 wire net3149;
 wire net3150;
 wire net3151;
 wire net3152;
 wire net3153;
 wire net3154;
 wire net3155;
 wire net3156;
 wire net3157;
 wire net3158;
 wire net3159;
 wire net3160;
 wire net3161;
 wire net3162;
 wire net3163;
 wire net3164;
 wire net3165;
 wire net3166;
 wire net3167;
 wire net3168;
 wire net3169;
 wire net3170;
 wire net3171;
 wire net3172;
 wire net3173;
 wire net3174;
 wire net3175;
 wire net3176;
 wire net3177;
 wire net3178;
 wire net3179;
 wire net3180;
 wire net3181;
 wire net3182;
 wire net3183;
 wire net3184;
 wire net3185;
 wire net3186;
 wire net3187;
 wire net3188;
 wire net3189;
 wire net3190;
 wire net3191;
 wire net3192;
 wire net3193;
 wire net3194;
 wire net3195;
 wire net3196;
 wire net3197;
 wire net3198;
 wire net3199;
 wire net3200;
 wire net3201;
 wire net3202;
 wire net3203;
 wire net3204;
 wire net3205;
 wire net3206;
 wire net3207;
 wire net3208;
 wire net3209;
 wire net3210;
 wire net3211;
 wire net3212;
 wire net3213;
 wire net3214;
 wire net3215;
 wire net3216;
 wire net3217;
 wire net3218;
 wire net3219;
 wire net3220;
 wire net3221;
 wire net3222;
 wire net3223;
 wire net3224;
 wire net3225;
 wire net3226;
 wire net3227;
 wire net3228;
 wire net3229;
 wire net3230;
 wire net3231;
 wire net3232;
 wire net3233;
 wire net3234;
 wire net3235;
 wire net3236;
 wire net3237;
 wire net3238;
 wire net3239;
 wire net3240;
 wire net3241;
 wire net3242;
 wire net3243;
 wire net3244;
 wire net3245;
 wire net3246;
 wire net3247;
 wire net3248;
 wire net3249;
 wire net3250;
 wire net3251;
 wire net3252;
 wire net3253;
 wire net3254;
 wire net3255;
 wire net3256;
 wire net3257;
 wire net3258;
 wire net3259;
 wire net3260;
 wire net3261;
 wire net3262;
 wire net3263;
 wire net3264;
 wire net3265;
 wire net3266;
 wire net3267;
 wire net3268;
 wire net3269;
 wire net3270;
 wire net3271;
 wire net3272;
 wire net3273;
 wire net3274;
 wire net3275;
 wire net3276;
 wire net3277;
 wire net3278;
 wire net3279;
 wire net3280;
 wire net3281;
 wire net3282;
 wire net3283;
 wire net3284;
 wire net3285;
 wire net3286;
 wire net3287;
 wire net3288;
 wire net3289;
 wire net3290;
 wire net3291;
 wire net3292;
 wire net3293;
 wire net3294;
 wire net3295;
 wire net3296;
 wire net3297;
 wire net3298;
 wire net3299;
 wire net3300;
 wire net3301;
 wire net3302;
 wire net3303;
 wire net3304;
 wire net3305;
 wire net3306;
 wire net3307;
 wire net3308;
 wire net3309;
 wire net3310;
 wire net3311;
 wire net3312;
 wire net3313;
 wire net3314;
 wire net3315;
 wire net3316;
 wire net3317;
 wire net3318;
 wire net3319;
 wire net3320;
 wire net3321;
 wire net3322;
 wire net3323;
 wire net3324;
 wire net3325;
 wire net3326;
 wire net3327;
 wire net3328;
 wire net3329;
 wire net3330;
 wire net3331;
 wire net3332;
 wire net3333;
 wire net3334;
 wire net3335;
 wire net3336;
 wire net3337;
 wire net3338;
 wire net3339;
 wire net3340;
 wire net3341;
 wire net3342;
 wire net3343;
 wire net3344;
 wire net3345;
 wire net3346;
 wire net3347;
 wire net3348;
 wire net3349;
 wire net3350;
 wire net3351;
 wire net3352;
 wire net3353;
 wire net3354;
 wire net3355;
 wire net3356;
 wire net3357;
 wire net3358;
 wire net3359;
 wire net3360;
 wire net3361;
 wire net3362;
 wire net3363;
 wire net3364;
 wire net3365;
 wire net3366;
 wire net3367;
 wire net3368;
 wire net3369;
 wire net3370;
 wire net3371;
 wire net3372;
 wire net3373;
 wire net3374;
 wire net3375;
 wire net3376;
 wire net3377;
 wire net3378;
 wire net3379;
 wire net3380;
 wire net3381;
 wire net3382;
 wire net3383;
 wire net3384;
 wire net3385;
 wire net3386;
 wire net3387;
 wire net3388;
 wire net3389;
 wire net3390;
 wire net3391;
 wire net3392;
 wire net3393;
 wire net3394;
 wire net3395;
 wire net3396;
 wire net3397;
 wire net3398;
 wire net3399;
 wire net3400;
 wire net3401;
 wire net3402;
 wire net3403;
 wire net3404;
 wire net3405;
 wire net3406;
 wire net3407;
 wire net3408;
 wire net3409;
 wire net3410;
 wire net3411;
 wire net3412;
 wire net3413;
 wire net3414;
 wire net3415;
 wire net3416;
 wire net3417;
 wire net3418;
 wire net3419;
 wire net3420;
 wire net3421;
 wire net3422;
 wire net3423;
 wire net3424;
 wire net3425;
 wire net3426;
 wire net3427;
 wire net3428;
 wire net3429;
 wire net3430;
 wire net3431;
 wire net3432;
 wire net3433;
 wire net3434;
 wire net3435;
 wire net3436;
 wire net3437;
 wire net3438;
 wire net3439;
 wire net3440;
 wire net3441;
 wire net3442;
 wire net3443;
 wire net3444;
 wire net3445;
 wire net3446;
 wire net3447;
 wire net3448;
 wire net3449;
 wire net3450;
 wire net3451;
 wire net3452;
 wire net3453;
 wire net3454;
 wire net3455;
 wire net3456;
 wire net3457;
 wire net3458;
 wire net3459;
 wire net3460;
 wire net3461;
 wire net3462;
 wire net3463;
 wire net3464;
 wire net3465;
 wire net3466;
 wire net3467;
 wire net3468;
 wire net3469;
 wire net3470;
 wire net3471;
 wire net3472;
 wire net3473;
 wire net3474;
 wire net3475;
 wire net3476;
 wire net3477;
 wire net3478;
 wire net3479;
 wire net3480;
 wire net3481;
 wire net3482;
 wire net3483;
 wire net3484;
 wire net3485;
 wire net3486;
 wire net3487;
 wire net3488;
 wire net3489;
 wire net3490;
 wire net3491;
 wire net3492;
 wire net3493;
 wire net3494;
 wire net3495;
 wire net3496;
 wire net3497;
 wire net3498;
 wire net3499;
 wire net3500;
 wire net3501;
 wire net3502;
 wire net3503;
 wire net3504;
 wire net3505;
 wire net3506;
 wire net3507;
 wire net3508;
 wire net3509;
 wire net3510;
 wire net3511;
 wire net3512;
 wire net3513;
 wire net3514;
 wire net3515;
 wire net3516;
 wire net3517;
 wire net3518;
 wire net3519;
 wire net3520;
 wire net3521;
 wire net3522;
 wire net3523;
 wire net3524;
 wire net3525;
 wire net3526;
 wire net3527;
 wire net3528;
 wire net3529;
 wire net3530;
 wire net3531;
 wire net3532;
 wire net3533;
 wire net3534;
 wire net3535;
 wire net3536;
 wire net3537;
 wire net3538;
 wire net3539;
 wire net3540;
 wire net3541;
 wire net3542;
 wire net3543;
 wire net3544;
 wire net3545;
 wire net3546;
 wire net3547;
 wire net3548;
 wire net3549;
 wire net3550;
 wire net3551;
 wire net3552;
 wire net3553;
 wire net3554;
 wire net3555;
 wire net3556;
 wire net3557;
 wire net3558;
 wire net3559;
 wire net3560;
 wire net3561;
 wire net3562;
 wire net3563;
 wire net3564;
 wire net3565;
 wire net3566;
 wire net3567;
 wire net3568;
 wire net3569;
 wire net3570;
 wire net3571;
 wire net3572;
 wire net3573;
 wire net3574;
 wire net3575;
 wire net3576;
 wire net3577;
 wire net3578;
 wire net3579;
 wire net3580;
 wire net3581;
 wire net3582;
 wire net3583;
 wire net3584;
 wire net3585;
 wire net3586;
 wire net3587;
 wire net3588;
 wire net3589;
 wire net3590;
 wire net3591;
 wire net3592;
 wire net3593;
 wire net3594;
 wire net3595;
 wire net3596;
 wire net3597;
 wire net3598;
 wire net3599;
 wire net3600;
 wire net3601;
 wire net3602;
 wire net3603;
 wire net3604;
 wire net3605;
 wire net3606;
 wire net3607;
 wire net3608;
 wire net3609;
 wire net3610;
 wire net3611;
 wire net3612;
 wire net3613;
 wire net3614;
 wire net3615;
 wire net3616;
 wire net3617;
 wire net3618;
 wire net3619;
 wire net3620;
 wire net3621;
 wire net3622;
 wire net3623;
 wire net3624;
 wire net3625;
 wire net3626;
 wire net3627;
 wire net3628;
 wire net3629;
 wire net3630;
 wire net3631;
 wire net3632;
 wire net3633;
 wire clknet_leaf_1_clk;
 wire clknet_leaf_2_clk;
 wire clknet_leaf_3_clk;
 wire clknet_leaf_4_clk;
 wire clknet_leaf_5_clk;
 wire clknet_leaf_6_clk;
 wire clknet_leaf_7_clk;
 wire clknet_leaf_8_clk;
 wire clknet_leaf_9_clk;
 wire clknet_leaf_10_clk;
 wire clknet_leaf_11_clk;
 wire clknet_leaf_12_clk;
 wire clknet_leaf_13_clk;
 wire clknet_leaf_14_clk;
 wire clknet_leaf_15_clk;
 wire clknet_leaf_16_clk;
 wire clknet_leaf_17_clk;
 wire clknet_leaf_18_clk;
 wire clknet_leaf_19_clk;
 wire clknet_leaf_20_clk;
 wire clknet_leaf_21_clk;
 wire clknet_leaf_22_clk;
 wire clknet_leaf_23_clk;
 wire clknet_leaf_24_clk;
 wire clknet_leaf_25_clk;
 wire clknet_leaf_26_clk;
 wire clknet_leaf_27_clk;
 wire clknet_leaf_28_clk;
 wire clknet_leaf_29_clk;
 wire clknet_leaf_30_clk;
 wire clknet_leaf_31_clk;
 wire clknet_leaf_32_clk;
 wire clknet_leaf_33_clk;
 wire clknet_leaf_34_clk;
 wire clknet_leaf_35_clk;
 wire clknet_leaf_36_clk;
 wire clknet_leaf_37_clk;
 wire clknet_leaf_38_clk;
 wire clknet_leaf_39_clk;
 wire clknet_leaf_40_clk;
 wire clknet_leaf_41_clk;
 wire clknet_leaf_42_clk;
 wire clknet_leaf_43_clk;
 wire clknet_leaf_44_clk;
 wire clknet_leaf_45_clk;
 wire clknet_leaf_46_clk;
 wire clknet_leaf_47_clk;
 wire clknet_leaf_48_clk;
 wire clknet_leaf_49_clk;
 wire clknet_leaf_50_clk;
 wire clknet_leaf_51_clk;
 wire clknet_leaf_52_clk;
 wire clknet_leaf_53_clk;
 wire clknet_leaf_54_clk;
 wire clknet_leaf_55_clk;
 wire clknet_leaf_56_clk;
 wire clknet_leaf_57_clk;
 wire clknet_leaf_58_clk;
 wire clknet_leaf_59_clk;
 wire clknet_leaf_60_clk;
 wire clknet_leaf_61_clk;
 wire clknet_leaf_62_clk;
 wire clknet_leaf_63_clk;
 wire clknet_leaf_64_clk;
 wire clknet_leaf_65_clk;
 wire clknet_leaf_66_clk;
 wire clknet_leaf_67_clk;
 wire clknet_leaf_68_clk;
 wire clknet_leaf_69_clk;
 wire clknet_leaf_70_clk;
 wire clknet_leaf_71_clk;
 wire clknet_leaf_72_clk;
 wire clknet_leaf_73_clk;
 wire clknet_leaf_74_clk;
 wire clknet_leaf_75_clk;
 wire clknet_leaf_76_clk;
 wire clknet_leaf_77_clk;
 wire clknet_leaf_78_clk;
 wire clknet_leaf_79_clk;
 wire clknet_leaf_80_clk;
 wire clknet_leaf_81_clk;
 wire clknet_leaf_82_clk;
 wire clknet_leaf_83_clk;
 wire clknet_leaf_84_clk;
 wire clknet_leaf_85_clk;
 wire clknet_leaf_86_clk;
 wire clknet_leaf_87_clk;
 wire clknet_leaf_88_clk;
 wire clknet_leaf_89_clk;
 wire clknet_leaf_90_clk;
 wire clknet_leaf_91_clk;
 wire clknet_leaf_92_clk;
 wire clknet_leaf_93_clk;
 wire clknet_leaf_94_clk;
 wire clknet_leaf_95_clk;
 wire clknet_leaf_96_clk;
 wire clknet_leaf_97_clk;
 wire clknet_leaf_98_clk;
 wire clknet_leaf_99_clk;
 wire clknet_leaf_100_clk;
 wire clknet_leaf_101_clk;
 wire clknet_leaf_102_clk;
 wire clknet_leaf_103_clk;
 wire clknet_leaf_104_clk;
 wire clknet_leaf_105_clk;
 wire clknet_leaf_106_clk;
 wire clknet_leaf_107_clk;
 wire clknet_leaf_108_clk;
 wire clknet_leaf_109_clk;
 wire clknet_leaf_110_clk;
 wire clknet_leaf_111_clk;
 wire clknet_leaf_112_clk;
 wire clknet_leaf_113_clk;
 wire clknet_leaf_114_clk;
 wire clknet_leaf_115_clk;
 wire clknet_leaf_116_clk;
 wire clknet_leaf_117_clk;
 wire clknet_leaf_118_clk;
 wire clknet_leaf_119_clk;
 wire clknet_leaf_120_clk;
 wire clknet_leaf_121_clk;
 wire clknet_leaf_122_clk;
 wire clknet_leaf_123_clk;
 wire clknet_leaf_124_clk;
 wire clknet_leaf_125_clk;
 wire clknet_leaf_126_clk;
 wire clknet_leaf_127_clk;
 wire clknet_leaf_128_clk;
 wire clknet_leaf_129_clk;
 wire clknet_leaf_130_clk;
 wire clknet_leaf_131_clk;
 wire clknet_leaf_132_clk;
 wire clknet_leaf_133_clk;
 wire clknet_leaf_134_clk;
 wire clknet_leaf_135_clk;
 wire clknet_leaf_136_clk;
 wire clknet_leaf_137_clk;
 wire clknet_leaf_138_clk;
 wire clknet_leaf_139_clk;
 wire clknet_leaf_140_clk;
 wire clknet_leaf_141_clk;
 wire clknet_leaf_142_clk;
 wire clknet_leaf_143_clk;
 wire clknet_leaf_144_clk;
 wire clknet_leaf_145_clk;
 wire clknet_leaf_146_clk;
 wire clknet_leaf_147_clk;
 wire clknet_leaf_148_clk;
 wire clknet_leaf_149_clk;
 wire clknet_leaf_150_clk;
 wire clknet_leaf_151_clk;
 wire clknet_leaf_152_clk;
 wire clknet_leaf_153_clk;
 wire clknet_leaf_154_clk;
 wire clknet_leaf_155_clk;
 wire clknet_leaf_156_clk;
 wire clknet_leaf_157_clk;
 wire clknet_leaf_158_clk;
 wire clknet_leaf_159_clk;
 wire clknet_leaf_160_clk;
 wire clknet_leaf_161_clk;
 wire clknet_leaf_162_clk;
 wire clknet_leaf_163_clk;
 wire clknet_leaf_164_clk;
 wire clknet_leaf_165_clk;
 wire clknet_leaf_166_clk;
 wire clknet_leaf_167_clk;
 wire clknet_leaf_168_clk;
 wire clknet_leaf_169_clk;
 wire clknet_leaf_170_clk;
 wire clknet_leaf_171_clk;
 wire clknet_leaf_172_clk;
 wire clknet_leaf_173_clk;
 wire clknet_leaf_174_clk;
 wire clknet_leaf_175_clk;
 wire clknet_leaf_176_clk;
 wire clknet_leaf_177_clk;
 wire clknet_leaf_178_clk;
 wire clknet_leaf_179_clk;
 wire clknet_leaf_180_clk;
 wire clknet_leaf_181_clk;
 wire clknet_leaf_182_clk;
 wire clknet_leaf_183_clk;
 wire clknet_leaf_184_clk;
 wire clknet_leaf_185_clk;
 wire clknet_leaf_186_clk;
 wire clknet_leaf_187_clk;
 wire clknet_leaf_188_clk;
 wire clknet_leaf_189_clk;
 wire clknet_leaf_190_clk;
 wire clknet_leaf_191_clk;
 wire clknet_leaf_192_clk;
 wire clknet_leaf_193_clk;
 wire clknet_leaf_194_clk;
 wire clknet_leaf_195_clk;
 wire clknet_leaf_196_clk;
 wire clknet_leaf_197_clk;
 wire clknet_leaf_198_clk;
 wire clknet_leaf_199_clk;
 wire clknet_leaf_200_clk;
 wire clknet_leaf_201_clk;
 wire clknet_leaf_202_clk;
 wire clknet_leaf_203_clk;
 wire clknet_leaf_204_clk;
 wire clknet_leaf_205_clk;
 wire clknet_leaf_206_clk;
 wire clknet_leaf_207_clk;
 wire clknet_leaf_208_clk;
 wire clknet_leaf_209_clk;
 wire clknet_leaf_210_clk;
 wire clknet_leaf_211_clk;
 wire clknet_leaf_212_clk;
 wire clknet_leaf_213_clk;
 wire clknet_leaf_214_clk;
 wire clknet_leaf_215_clk;
 wire clknet_leaf_216_clk;
 wire clknet_leaf_217_clk;
 wire clknet_leaf_218_clk;
 wire clknet_leaf_219_clk;
 wire clknet_leaf_220_clk;
 wire clknet_leaf_221_clk;
 wire clknet_leaf_222_clk;
 wire clknet_leaf_223_clk;
 wire clknet_leaf_224_clk;
 wire clknet_leaf_225_clk;
 wire clknet_leaf_226_clk;
 wire clknet_leaf_227_clk;
 wire clknet_leaf_228_clk;
 wire clknet_leaf_229_clk;
 wire clknet_leaf_230_clk;
 wire clknet_leaf_231_clk;
 wire clknet_leaf_232_clk;
 wire clknet_leaf_233_clk;
 wire clknet_leaf_234_clk;
 wire clknet_leaf_235_clk;
 wire clknet_leaf_236_clk;
 wire clknet_leaf_237_clk;
 wire clknet_leaf_238_clk;
 wire clknet_leaf_239_clk;
 wire clknet_leaf_240_clk;
 wire clknet_leaf_241_clk;
 wire clknet_leaf_242_clk;
 wire clknet_leaf_243_clk;
 wire clknet_leaf_244_clk;
 wire clknet_leaf_245_clk;
 wire clknet_leaf_246_clk;
 wire clknet_leaf_247_clk;
 wire clknet_leaf_248_clk;
 wire clknet_leaf_249_clk;
 wire clknet_leaf_250_clk;
 wire clknet_leaf_251_clk;
 wire clknet_leaf_252_clk;
 wire clknet_leaf_253_clk;
 wire clknet_leaf_254_clk;
 wire clknet_leaf_255_clk;
 wire clknet_leaf_256_clk;
 wire clknet_leaf_257_clk;
 wire clknet_leaf_258_clk;
 wire clknet_leaf_259_clk;
 wire clknet_leaf_260_clk;
 wire clknet_leaf_261_clk;
 wire clknet_leaf_262_clk;
 wire clknet_leaf_263_clk;
 wire clknet_leaf_264_clk;
 wire clknet_leaf_265_clk;
 wire clknet_leaf_266_clk;
 wire clknet_leaf_267_clk;
 wire clknet_leaf_268_clk;
 wire clknet_leaf_269_clk;
 wire clknet_leaf_270_clk;
 wire clknet_leaf_271_clk;
 wire clknet_leaf_272_clk;
 wire clknet_leaf_273_clk;
 wire clknet_leaf_274_clk;
 wire clknet_leaf_275_clk;
 wire clknet_leaf_276_clk;
 wire clknet_leaf_277_clk;
 wire clknet_leaf_278_clk;
 wire clknet_leaf_279_clk;
 wire clknet_leaf_280_clk;
 wire clknet_leaf_281_clk;
 wire clknet_leaf_282_clk;
 wire clknet_leaf_283_clk;
 wire clknet_leaf_284_clk;
 wire clknet_leaf_285_clk;
 wire clknet_leaf_286_clk;
 wire clknet_leaf_287_clk;
 wire clknet_leaf_288_clk;
 wire clknet_leaf_289_clk;
 wire clknet_leaf_290_clk;
 wire clknet_leaf_291_clk;
 wire clknet_leaf_292_clk;
 wire clknet_leaf_293_clk;
 wire clknet_leaf_294_clk;
 wire clknet_leaf_295_clk;
 wire clknet_leaf_296_clk;
 wire clknet_leaf_297_clk;
 wire clknet_leaf_298_clk;
 wire clknet_leaf_299_clk;
 wire clknet_leaf_300_clk;
 wire clknet_leaf_301_clk;
 wire clknet_leaf_302_clk;
 wire clknet_leaf_303_clk;
 wire clknet_leaf_304_clk;
 wire clknet_leaf_305_clk;
 wire clknet_leaf_306_clk;
 wire clknet_leaf_307_clk;
 wire clknet_leaf_308_clk;
 wire clknet_leaf_309_clk;
 wire clknet_leaf_310_clk;
 wire clknet_leaf_311_clk;
 wire clknet_leaf_312_clk;
 wire clknet_0_clk;
 wire clknet_3_0_0_clk;
 wire clknet_3_1_0_clk;
 wire clknet_3_2_0_clk;
 wire clknet_3_3_0_clk;
 wire clknet_3_4_0_clk;
 wire clknet_3_5_0_clk;
 wire clknet_3_6_0_clk;
 wire clknet_3_7_0_clk;
 wire clknet_6_0__leaf_clk;
 wire clknet_6_1__leaf_clk;
 wire clknet_6_2__leaf_clk;
 wire clknet_6_3__leaf_clk;
 wire clknet_6_4__leaf_clk;
 wire clknet_6_5__leaf_clk;
 wire clknet_6_6__leaf_clk;
 wire clknet_6_7__leaf_clk;
 wire clknet_6_8__leaf_clk;
 wire clknet_6_9__leaf_clk;
 wire clknet_6_10__leaf_clk;
 wire clknet_6_11__leaf_clk;
 wire clknet_6_12__leaf_clk;
 wire clknet_6_13__leaf_clk;
 wire clknet_6_14__leaf_clk;
 wire clknet_6_15__leaf_clk;
 wire clknet_6_16__leaf_clk;
 wire clknet_6_17__leaf_clk;
 wire clknet_6_18__leaf_clk;
 wire clknet_6_19__leaf_clk;
 wire clknet_6_20__leaf_clk;
 wire clknet_6_21__leaf_clk;
 wire clknet_6_22__leaf_clk;
 wire clknet_6_23__leaf_clk;
 wire clknet_6_24__leaf_clk;
 wire clknet_6_25__leaf_clk;
 wire clknet_6_26__leaf_clk;
 wire clknet_6_27__leaf_clk;
 wire clknet_6_28__leaf_clk;
 wire clknet_6_29__leaf_clk;
 wire clknet_6_30__leaf_clk;
 wire clknet_6_31__leaf_clk;
 wire clknet_6_32__leaf_clk;
 wire clknet_6_33__leaf_clk;
 wire clknet_6_34__leaf_clk;
 wire clknet_6_35__leaf_clk;
 wire clknet_6_36__leaf_clk;
 wire clknet_6_37__leaf_clk;
 wire clknet_6_38__leaf_clk;
 wire clknet_6_39__leaf_clk;
 wire clknet_6_40__leaf_clk;
 wire clknet_6_41__leaf_clk;
 wire clknet_6_42__leaf_clk;
 wire clknet_6_43__leaf_clk;
 wire clknet_6_44__leaf_clk;
 wire clknet_6_45__leaf_clk;
 wire clknet_6_46__leaf_clk;
 wire clknet_6_47__leaf_clk;
 wire clknet_6_48__leaf_clk;
 wire clknet_6_49__leaf_clk;
 wire clknet_6_50__leaf_clk;
 wire clknet_6_51__leaf_clk;
 wire clknet_6_52__leaf_clk;
 wire clknet_6_53__leaf_clk;
 wire clknet_6_54__leaf_clk;
 wire clknet_6_55__leaf_clk;
 wire clknet_6_56__leaf_clk;
 wire clknet_6_57__leaf_clk;
 wire clknet_6_58__leaf_clk;
 wire clknet_6_59__leaf_clk;
 wire clknet_6_60__leaf_clk;
 wire clknet_6_61__leaf_clk;
 wire clknet_6_62__leaf_clk;
 wire clknet_6_63__leaf_clk;

 sg13g2_buf_2 _15084_ (.A(\cpu.dec.r_op[6] ),
    .X(_08335_));
 sg13g2_buf_1 _15085_ (.A(_08335_),
    .X(_08336_));
 sg13g2_buf_1 _15086_ (.A(net1090),
    .X(_08337_));
 sg13g2_buf_8 _15087_ (.A(\cpu.ex.genblk3.r_mmu_enable ),
    .X(_08338_));
 sg13g2_inv_2 _15088_ (.Y(_08339_),
    .A(net1149));
 sg13g2_buf_2 _15089_ (.A(\cpu.ex.io_access ),
    .X(_08340_));
 sg13g2_buf_8 _15090_ (.A(\cpu.ex.r_wmask[0] ),
    .X(_08341_));
 sg13g2_nor2_1 _15091_ (.A(\cpu.ex.r_wmask[1] ),
    .B(_08341_),
    .Y(_08342_));
 sg13g2_buf_2 _15092_ (.A(_08342_),
    .X(_08343_));
 sg13g2_nor3_2 _15093_ (.A(_08339_),
    .B(_08340_),
    .C(_08343_),
    .Y(_08344_));
 sg13g2_buf_8 _15094_ (.A(\cpu.ex.ifetch ),
    .X(_08345_));
 sg13g2_inv_4 _15095_ (.A(_08345_),
    .Y(_08346_));
 sg13g2_buf_2 _15096_ (.A(\cpu.ex.genblk3.r_mmu_d_proxy ),
    .X(_08347_));
 sg13g2_buf_2 _15097_ (.A(_00183_),
    .X(_08348_));
 sg13g2_a21oi_2 _15098_ (.B1(_08348_),
    .Y(_08349_),
    .A2(_08347_),
    .A1(_08346_));
 sg13g2_buf_8 _15099_ (.A(\cpu.addr[13] ),
    .X(_08350_));
 sg13g2_buf_8 _15100_ (.A(_08350_),
    .X(_08351_));
 sg13g2_buf_8 _15101_ (.A(\cpu.addr[12] ),
    .X(_08352_));
 sg13g2_buf_1 _15102_ (.A(\cpu.addr[15] ),
    .X(_08353_));
 sg13g2_nor2_1 _15103_ (.A(_08352_),
    .B(_08353_),
    .Y(_08354_));
 sg13g2_buf_8 _15104_ (.A(\cpu.addr[14] ),
    .X(_08355_));
 sg13g2_mux2_1 _15105_ (.A0(\cpu.genblk1.mmu.r_writeable_d[18] ),
    .A1(\cpu.genblk1.mmu.r_writeable_d[22] ),
    .S(net1148),
    .X(_08356_));
 sg13g2_nand3_1 _15106_ (.B(_08354_),
    .C(_08356_),
    .A(_08351_),
    .Y(_08357_));
 sg13g2_nor2b_1 _15107_ (.A(_08353_),
    .B_N(_08352_),
    .Y(_08358_));
 sg13g2_mux4_1 _15108_ (.S0(_08350_),
    .A0(\cpu.genblk1.mmu.r_writeable_d[17] ),
    .A1(\cpu.genblk1.mmu.r_writeable_d[19] ),
    .A2(\cpu.genblk1.mmu.r_writeable_d[21] ),
    .A3(\cpu.genblk1.mmu.r_writeable_d[23] ),
    .S1(net1148),
    .X(_08359_));
 sg13g2_nor3_1 _15109_ (.A(_08352_),
    .B(_08351_),
    .C(_08353_),
    .Y(_08360_));
 sg13g2_mux2_1 _15110_ (.A0(\cpu.genblk1.mmu.r_writeable_d[16] ),
    .A1(\cpu.genblk1.mmu.r_writeable_d[20] ),
    .S(net1148),
    .X(_08361_));
 sg13g2_a22oi_1 _15111_ (.Y(_08362_),
    .B1(_08360_),
    .B2(_08361_),
    .A2(_08359_),
    .A1(_08358_));
 sg13g2_and4_1 _15112_ (.A(_08344_),
    .B(_08349_),
    .C(_08357_),
    .D(_08362_),
    .X(_08363_));
 sg13g2_buf_8 _15113_ (.A(net1089),
    .X(_08364_));
 sg13g2_buf_8 _15114_ (.A(_08352_),
    .X(_08365_));
 sg13g2_buf_8 _15115_ (.A(_08355_),
    .X(_08366_));
 sg13g2_mux4_1 _15116_ (.S0(net1088),
    .A0(\cpu.genblk1.mmu.r_writeable_d[26] ),
    .A1(\cpu.genblk1.mmu.r_writeable_d[27] ),
    .A2(\cpu.genblk1.mmu.r_writeable_d[30] ),
    .A3(\cpu.genblk1.mmu.r_writeable_d[31] ),
    .S1(net1087),
    .X(_08367_));
 sg13g2_mux4_1 _15117_ (.S0(_08352_),
    .A0(\cpu.genblk1.mmu.r_writeable_d[24] ),
    .A1(\cpu.genblk1.mmu.r_writeable_d[25] ),
    .A2(\cpu.genblk1.mmu.r_writeable_d[28] ),
    .A3(\cpu.genblk1.mmu.r_writeable_d[29] ),
    .S1(_08355_),
    .X(_08368_));
 sg13g2_nor2b_1 _15118_ (.A(net947),
    .B_N(_08368_),
    .Y(_08369_));
 sg13g2_a21oi_1 _15119_ (.A1(net947),
    .A2(_08367_),
    .Y(_08370_),
    .B1(_08369_));
 sg13g2_a21o_1 _15120_ (.A2(_08347_),
    .A1(_08346_),
    .B1(_08348_),
    .X(_08371_));
 sg13g2_buf_2 _15121_ (.A(_08371_),
    .X(_08372_));
 sg13g2_mux2_1 _15122_ (.A0(\cpu.genblk1.mmu.r_writeable_d[2] ),
    .A1(\cpu.genblk1.mmu.r_writeable_d[6] ),
    .S(net1148),
    .X(_08373_));
 sg13g2_nand3_1 _15123_ (.B(_08354_),
    .C(_08373_),
    .A(net947),
    .Y(_08374_));
 sg13g2_mux4_1 _15124_ (.S0(net1089),
    .A0(\cpu.genblk1.mmu.r_writeable_d[1] ),
    .A1(\cpu.genblk1.mmu.r_writeable_d[3] ),
    .A2(\cpu.genblk1.mmu.r_writeable_d[5] ),
    .A3(\cpu.genblk1.mmu.r_writeable_d[7] ),
    .S1(net1148),
    .X(_08375_));
 sg13g2_mux2_1 _15125_ (.A0(\cpu.genblk1.mmu.r_writeable_d[0] ),
    .A1(\cpu.genblk1.mmu.r_writeable_d[4] ),
    .S(net1148),
    .X(_08376_));
 sg13g2_a22oi_1 _15126_ (.Y(_08377_),
    .B1(_08376_),
    .B2(_08360_),
    .A2(_08375_),
    .A1(_08358_));
 sg13g2_and4_1 _15127_ (.A(_08344_),
    .B(net826),
    .C(_08374_),
    .D(_08377_),
    .X(_08378_));
 sg13g2_mux4_1 _15128_ (.S0(net1088),
    .A0(\cpu.genblk1.mmu.r_writeable_d[8] ),
    .A1(\cpu.genblk1.mmu.r_writeable_d[9] ),
    .A2(\cpu.genblk1.mmu.r_writeable_d[12] ),
    .A3(\cpu.genblk1.mmu.r_writeable_d[13] ),
    .S1(net1087),
    .X(_08379_));
 sg13g2_mux4_1 _15129_ (.S0(_08352_),
    .A0(\cpu.genblk1.mmu.r_writeable_d[10] ),
    .A1(\cpu.genblk1.mmu.r_writeable_d[11] ),
    .A2(\cpu.genblk1.mmu.r_writeable_d[14] ),
    .A3(\cpu.genblk1.mmu.r_writeable_d[15] ),
    .S1(_08366_),
    .X(_08380_));
 sg13g2_nand2b_1 _15130_ (.Y(_08381_),
    .B(_08364_),
    .A_N(_08380_));
 sg13g2_o21ai_1 _15131_ (.B1(_08381_),
    .Y(_08382_),
    .A1(net947),
    .A2(_08379_));
 sg13g2_a22oi_1 _15132_ (.Y(_08383_),
    .B1(_08378_),
    .B2(_08382_),
    .A2(_08370_),
    .A1(_08363_));
 sg13g2_buf_1 _15133_ (.A(_08353_),
    .X(_08384_));
 sg13g2_inv_2 _15134_ (.Y(_08385_),
    .A(_08384_));
 sg13g2_o21ai_1 _15135_ (.B1(_08385_),
    .Y(_08386_),
    .A1(_08363_),
    .A2(_08378_));
 sg13g2_and2_1 _15136_ (.A(_08383_),
    .B(_08386_),
    .X(_08387_));
 sg13g2_buf_1 _15137_ (.A(_08387_),
    .X(_08388_));
 sg13g2_buf_8 _15138_ (.A(\cpu.ex.pc[13] ),
    .X(_08389_));
 sg13g2_buf_8 _15139_ (.A(_08389_),
    .X(_08390_));
 sg13g2_buf_8 _15140_ (.A(\cpu.ex.pc[14] ),
    .X(_08391_));
 sg13g2_buf_1 _15141_ (.A(_08391_),
    .X(_08392_));
 sg13g2_mux4_1 _15142_ (.S0(net1085),
    .A0(\cpu.genblk1.mmu.r_valid_i[0] ),
    .A1(\cpu.genblk1.mmu.r_valid_i[2] ),
    .A2(\cpu.genblk1.mmu.r_valid_i[4] ),
    .A3(\cpu.genblk1.mmu.r_valid_i[6] ),
    .S1(_08392_),
    .X(_08393_));
 sg13g2_mux4_1 _15143_ (.S0(net1085),
    .A0(\cpu.genblk1.mmu.r_valid_i[1] ),
    .A1(\cpu.genblk1.mmu.r_valid_i[3] ),
    .A2(\cpu.genblk1.mmu.r_valid_i[5] ),
    .A3(\cpu.genblk1.mmu.r_valid_i[7] ),
    .S1(net1084),
    .X(_08394_));
 sg13g2_buf_1 _15144_ (.A(\cpu.ex.pc[12] ),
    .X(_08395_));
 sg13g2_mux2_1 _15145_ (.A0(_08393_),
    .A1(_08394_),
    .S(net1147),
    .X(_08396_));
 sg13g2_buf_2 _15146_ (.A(\cpu.ex.pc[15] ),
    .X(_08397_));
 sg13g2_mux2_1 _15147_ (.A0(\cpu.genblk1.mmu.r_valid_i[8] ),
    .A1(\cpu.genblk1.mmu.r_valid_i[12] ),
    .S(_08391_),
    .X(_08398_));
 sg13g2_mux2_1 _15148_ (.A0(\cpu.genblk1.mmu.r_valid_i[9] ),
    .A1(\cpu.genblk1.mmu.r_valid_i[13] ),
    .S(_08391_),
    .X(_08399_));
 sg13g2_mux2_1 _15149_ (.A0(\cpu.genblk1.mmu.r_valid_i[10] ),
    .A1(\cpu.genblk1.mmu.r_valid_i[14] ),
    .S(_08391_),
    .X(_08400_));
 sg13g2_mux2_1 _15150_ (.A0(\cpu.genblk1.mmu.r_valid_i[11] ),
    .A1(\cpu.genblk1.mmu.r_valid_i[15] ),
    .S(_08391_),
    .X(_08401_));
 sg13g2_mux4_1 _15151_ (.S0(net1147),
    .A0(_08398_),
    .A1(_08399_),
    .A2(_08400_),
    .A3(_08401_),
    .S1(net1085),
    .X(_08402_));
 sg13g2_buf_8 _15152_ (.A(\cpu.dec.supmode ),
    .X(_08403_));
 sg13g2_inv_2 _15153_ (.Y(_08404_),
    .A(net1146));
 sg13g2_buf_1 _15154_ (.A(_08404_),
    .X(_08405_));
 sg13g2_nand3_1 _15155_ (.B(net1149),
    .C(_08345_),
    .A(net946),
    .Y(_08406_));
 sg13g2_a21o_1 _15156_ (.A2(_08402_),
    .A1(_08397_),
    .B1(_08406_),
    .X(_08407_));
 sg13g2_mux4_1 _15157_ (.S0(net1085),
    .A0(\cpu.genblk1.mmu.r_valid_i[16] ),
    .A1(\cpu.genblk1.mmu.r_valid_i[18] ),
    .A2(\cpu.genblk1.mmu.r_valid_i[20] ),
    .A3(\cpu.genblk1.mmu.r_valid_i[22] ),
    .S1(_08391_),
    .X(_08408_));
 sg13g2_mux4_1 _15158_ (.S0(_08389_),
    .A0(\cpu.genblk1.mmu.r_valid_i[17] ),
    .A1(\cpu.genblk1.mmu.r_valid_i[19] ),
    .A2(\cpu.genblk1.mmu.r_valid_i[21] ),
    .A3(\cpu.genblk1.mmu.r_valid_i[23] ),
    .S1(_08391_),
    .X(_08409_));
 sg13g2_mux2_1 _15159_ (.A0(_08408_),
    .A1(_08409_),
    .S(_08395_),
    .X(_08410_));
 sg13g2_nand3_1 _15160_ (.B(net1149),
    .C(_08345_),
    .A(net1146),
    .Y(_08411_));
 sg13g2_or3_1 _15161_ (.A(_08397_),
    .B(_08410_),
    .C(_08411_),
    .X(_08412_));
 sg13g2_o21ai_1 _15162_ (.B1(_08412_),
    .Y(_08413_),
    .A1(_08396_),
    .A2(_08407_));
 sg13g2_mux4_1 _15163_ (.S0(_08390_),
    .A0(\cpu.genblk1.mmu.r_valid_i[24] ),
    .A1(\cpu.genblk1.mmu.r_valid_i[26] ),
    .A2(\cpu.genblk1.mmu.r_valid_i[28] ),
    .A3(\cpu.genblk1.mmu.r_valid_i[30] ),
    .S1(_08392_),
    .X(_08414_));
 sg13g2_mux4_1 _15164_ (.S0(_08390_),
    .A0(\cpu.genblk1.mmu.r_valid_i[25] ),
    .A1(\cpu.genblk1.mmu.r_valid_i[27] ),
    .A2(\cpu.genblk1.mmu.r_valid_i[29] ),
    .A3(\cpu.genblk1.mmu.r_valid_i[31] ),
    .S1(_08391_),
    .X(_08415_));
 sg13g2_mux2_1 _15165_ (.A0(_08414_),
    .A1(_08415_),
    .S(_08395_),
    .X(_08416_));
 sg13g2_or2_1 _15166_ (.X(_08417_),
    .B(_08416_),
    .A(_08411_));
 sg13g2_inv_2 _15167_ (.Y(_08418_),
    .A(_08397_));
 sg13g2_a21oi_2 _15168_ (.B1(_08418_),
    .Y(_08419_),
    .A2(_08417_),
    .A1(_08407_));
 sg13g2_buf_1 _15169_ (.A(\cpu.ex.r_read_stall ),
    .X(_08420_));
 sg13g2_nand3b_1 _15170_ (.B(_08343_),
    .C(_00179_),
    .Y(_08421_),
    .A_N(_08420_));
 sg13g2_o21ai_1 _15171_ (.B1(_08421_),
    .Y(_08422_),
    .A1(_08413_),
    .A2(_08419_));
 sg13g2_buf_1 _15172_ (.A(_08422_),
    .X(_08423_));
 sg13g2_nand2b_1 _15173_ (.Y(_08424_),
    .B(net1086),
    .A_N(net1088));
 sg13g2_mux2_1 _15174_ (.A0(\cpu.genblk1.mmu.r_valid_d[24] ),
    .A1(\cpu.genblk1.mmu.r_valid_d[28] ),
    .S(net1148),
    .X(_08425_));
 sg13g2_nor2_1 _15175_ (.A(_08424_),
    .B(_08425_),
    .Y(_08426_));
 sg13g2_nor3_1 _15176_ (.A(net947),
    .B(net826),
    .C(_08426_),
    .Y(_08427_));
 sg13g2_nand2b_1 _15177_ (.Y(_08428_),
    .B(net1087),
    .A_N(\cpu.genblk1.mmu.r_valid_d[20] ));
 sg13g2_o21ai_1 _15178_ (.B1(_08428_),
    .Y(_08429_),
    .A1(net1087),
    .A2(\cpu.genblk1.mmu.r_valid_d[16] ));
 sg13g2_nand2b_1 _15179_ (.Y(_08430_),
    .B(net1087),
    .A_N(\cpu.genblk1.mmu.r_valid_d[21] ));
 sg13g2_o21ai_1 _15180_ (.B1(_08430_),
    .Y(_08431_),
    .A1(net1087),
    .A2(\cpu.genblk1.mmu.r_valid_d[17] ));
 sg13g2_nand2_1 _15181_ (.Y(_08432_),
    .A(net1088),
    .B(net1086));
 sg13g2_mux2_1 _15182_ (.A0(\cpu.genblk1.mmu.r_valid_d[25] ),
    .A1(\cpu.genblk1.mmu.r_valid_d[29] ),
    .S(net1148),
    .X(_08433_));
 sg13g2_nor2_1 _15183_ (.A(_08432_),
    .B(_08433_),
    .Y(_08434_));
 sg13g2_a221oi_1 _15184_ (.B2(_08358_),
    .C1(_08434_),
    .B1(_08431_),
    .A1(_08354_),
    .Y(_08435_),
    .A2(_08429_));
 sg13g2_buf_2 _15185_ (.A(_08366_),
    .X(_08436_));
 sg13g2_mux2_1 _15186_ (.A0(\cpu.genblk1.mmu.r_valid_d[8] ),
    .A1(\cpu.genblk1.mmu.r_valid_d[10] ),
    .S(net1089),
    .X(_08437_));
 sg13g2_nor2_1 _15187_ (.A(_08424_),
    .B(_08437_),
    .Y(_08438_));
 sg13g2_nor3_1 _15188_ (.A(net945),
    .B(_08349_),
    .C(_08438_),
    .Y(_08439_));
 sg13g2_nand2b_1 _15189_ (.Y(_08440_),
    .B(net1089),
    .A_N(\cpu.genblk1.mmu.r_valid_d[2] ));
 sg13g2_o21ai_1 _15190_ (.B1(_08440_),
    .Y(_08441_),
    .A1(\cpu.genblk1.mmu.r_valid_d[0] ),
    .A2(net947));
 sg13g2_nand2b_1 _15191_ (.Y(_08442_),
    .B(net1089),
    .A_N(\cpu.genblk1.mmu.r_valid_d[3] ));
 sg13g2_o21ai_1 _15192_ (.B1(_08442_),
    .Y(_08443_),
    .A1(\cpu.genblk1.mmu.r_valid_d[1] ),
    .A2(net947));
 sg13g2_mux2_1 _15193_ (.A0(\cpu.genblk1.mmu.r_valid_d[9] ),
    .A1(\cpu.genblk1.mmu.r_valid_d[11] ),
    .S(net1089),
    .X(_08444_));
 sg13g2_nor2_1 _15194_ (.A(_08432_),
    .B(_08444_),
    .Y(_08445_));
 sg13g2_a221oi_1 _15195_ (.B2(_08358_),
    .C1(_08445_),
    .B1(_08443_),
    .A1(_08354_),
    .Y(_08446_),
    .A2(_08441_));
 sg13g2_a22oi_1 _15196_ (.Y(_08447_),
    .B1(_08439_),
    .B2(_08446_),
    .A2(_08435_),
    .A1(_08427_));
 sg13g2_mux4_1 _15197_ (.S0(net1088),
    .A0(\cpu.genblk1.mmu.r_valid_d[26] ),
    .A1(\cpu.genblk1.mmu.r_valid_d[27] ),
    .A2(\cpu.genblk1.mmu.r_valid_d[30] ),
    .A3(\cpu.genblk1.mmu.r_valid_d[31] ),
    .S1(net1087),
    .X(_08448_));
 sg13g2_mux4_1 _15198_ (.S0(net1088),
    .A0(\cpu.genblk1.mmu.r_valid_d[18] ),
    .A1(\cpu.genblk1.mmu.r_valid_d[19] ),
    .A2(\cpu.genblk1.mmu.r_valid_d[22] ),
    .A3(\cpu.genblk1.mmu.r_valid_d[23] ),
    .S1(net1087),
    .X(_08449_));
 sg13g2_mux2_1 _15199_ (.A0(_08448_),
    .A1(_08449_),
    .S(_08385_),
    .X(_08450_));
 sg13g2_nand3_1 _15200_ (.B(_08349_),
    .C(_08450_),
    .A(net947),
    .Y(_08451_));
 sg13g2_buf_1 _15201_ (.A(\cpu.ex.mmu_reg_data[0] ),
    .X(_08452_));
 sg13g2_buf_1 _15202_ (.A(\cpu.cond[0] ),
    .X(_08453_));
 sg13g2_buf_1 _15203_ (.A(_00188_),
    .X(_08454_));
 sg13g2_a21oi_2 _15204_ (.B1(net1143),
    .Y(_08455_),
    .A2(net1144),
    .A1(net1145));
 sg13g2_or2_1 _15205_ (.X(_08456_),
    .B(_08455_),
    .A(_08420_));
 sg13g2_nor2b_1 _15206_ (.A(net1145),
    .B_N(net1144),
    .Y(_08457_));
 sg13g2_nand2_1 _15207_ (.Y(_08458_),
    .A(net1149),
    .B(_00187_));
 sg13g2_a21oi_1 _15208_ (.A1(net1143),
    .A2(_08457_),
    .Y(_08459_),
    .B1(_08458_));
 sg13g2_a21o_1 _15209_ (.A2(_08459_),
    .A1(_08456_),
    .B1(_08344_),
    .X(_08460_));
 sg13g2_mux4_1 _15210_ (.S0(net1088),
    .A0(\cpu.genblk1.mmu.r_valid_d[4] ),
    .A1(\cpu.genblk1.mmu.r_valid_d[5] ),
    .A2(\cpu.genblk1.mmu.r_valid_d[6] ),
    .A3(\cpu.genblk1.mmu.r_valid_d[7] ),
    .S1(net1089),
    .X(_08461_));
 sg13g2_nand4_1 _15211_ (.B(_08385_),
    .C(net826),
    .A(net945),
    .Y(_08462_),
    .D(_08461_));
 sg13g2_mux4_1 _15212_ (.S0(net1088),
    .A0(\cpu.genblk1.mmu.r_valid_d[12] ),
    .A1(\cpu.genblk1.mmu.r_valid_d[13] ),
    .A2(\cpu.genblk1.mmu.r_valid_d[14] ),
    .A3(\cpu.genblk1.mmu.r_valid_d[15] ),
    .S1(net1089),
    .X(_08463_));
 sg13g2_nand4_1 _15213_ (.B(net1086),
    .C(net826),
    .A(net945),
    .Y(_08464_),
    .D(_08463_));
 sg13g2_and4_1 _15214_ (.A(_08421_),
    .B(_08460_),
    .C(_08462_),
    .D(_08464_),
    .X(_08465_));
 sg13g2_nand3_1 _15215_ (.B(_08451_),
    .C(_08465_),
    .A(_08447_),
    .Y(_08466_));
 sg13g2_buf_1 _15216_ (.A(_08466_),
    .X(_08467_));
 sg13g2_nand3_1 _15217_ (.B(_08423_),
    .C(_08467_),
    .A(_08388_),
    .Y(_08468_));
 sg13g2_buf_1 _15218_ (.A(_08468_),
    .X(_08469_));
 sg13g2_buf_8 _15219_ (.A(_08469_),
    .X(_08470_));
 sg13g2_nor2_1 _15220_ (.A(_00179_),
    .B(_08470_),
    .Y(_08471_));
 sg13g2_buf_1 _15221_ (.A(net1085),
    .X(_08472_));
 sg13g2_buf_1 _15222_ (.A(net944),
    .X(_08473_));
 sg13g2_buf_1 _15223_ (.A(net825),
    .X(_08474_));
 sg13g2_buf_1 _15224_ (.A(net1149),
    .X(_08475_));
 sg13g2_buf_4 _15225_ (.X(_08476_),
    .A(net1147));
 sg13g2_buf_2 _15226_ (.A(_08476_),
    .X(_08477_));
 sg13g2_buf_1 _15227_ (.A(net944),
    .X(_08478_));
 sg13g2_mux4_1 _15228_ (.S0(net943),
    .A0(\cpu.genblk1.mmu.r_vtop_i[24][1] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[25][1] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[26][1] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[27][1] ),
    .S1(net824),
    .X(_08479_));
 sg13g2_mux4_1 _15229_ (.S0(net943),
    .A0(\cpu.genblk1.mmu.r_vtop_i[16][1] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[17][1] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[18][1] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[19][1] ),
    .S1(net824),
    .X(_08480_));
 sg13g2_buf_2 _15230_ (.A(_08476_),
    .X(_08481_));
 sg13g2_mux4_1 _15231_ (.S0(net942),
    .A0(\cpu.genblk1.mmu.r_vtop_i[28][1] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[29][1] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[30][1] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[31][1] ),
    .S1(net825),
    .X(_08482_));
 sg13g2_mux4_1 _15232_ (.S0(net942),
    .A0(\cpu.genblk1.mmu.r_vtop_i[20][1] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[21][1] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[22][1] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[23][1] ),
    .S1(net824),
    .X(_08483_));
 sg13g2_buf_2 _15233_ (.A(_08418_),
    .X(_08484_));
 sg13g2_buf_1 _15234_ (.A(net1084),
    .X(_08485_));
 sg13g2_mux4_1 _15235_ (.S0(net941),
    .A0(_08479_),
    .A1(_08480_),
    .A2(_08482_),
    .A3(_08483_),
    .S1(net940),
    .X(_08486_));
 sg13g2_nand2_1 _15236_ (.Y(_08487_),
    .A(net1146),
    .B(_08486_));
 sg13g2_buf_1 _15237_ (.A(_08405_),
    .X(_08488_));
 sg13g2_mux4_1 _15238_ (.S0(net943),
    .A0(\cpu.genblk1.mmu.r_vtop_i[8][1] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[9][1] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[10][1] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[11][1] ),
    .S1(net824),
    .X(_08489_));
 sg13g2_mux4_1 _15239_ (.S0(net943),
    .A0(\cpu.genblk1.mmu.r_vtop_i[0][1] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[1][1] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[2][1] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[3][1] ),
    .S1(net824),
    .X(_08490_));
 sg13g2_mux4_1 _15240_ (.S0(net942),
    .A0(\cpu.genblk1.mmu.r_vtop_i[12][1] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[13][1] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[14][1] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[15][1] ),
    .S1(net825),
    .X(_08491_));
 sg13g2_mux4_1 _15241_ (.S0(net942),
    .A0(\cpu.genblk1.mmu.r_vtop_i[4][1] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[5][1] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[6][1] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[7][1] ),
    .S1(net825),
    .X(_08492_));
 sg13g2_mux4_1 _15242_ (.S0(net941),
    .A0(_08489_),
    .A1(_08490_),
    .A2(_08491_),
    .A3(_08492_),
    .S1(net940),
    .X(_08493_));
 sg13g2_nand2_1 _15243_ (.Y(_08494_),
    .A(net823),
    .B(_08493_));
 sg13g2_nand3_1 _15244_ (.B(_08487_),
    .C(_08494_),
    .A(net1083),
    .Y(_08495_));
 sg13g2_o21ai_1 _15245_ (.B1(_08495_),
    .Y(_08496_),
    .A1(net726),
    .A2(net1083));
 sg13g2_buf_2 _15246_ (.A(_08496_),
    .X(_08497_));
 sg13g2_buf_2 _15247_ (.A(_00180_),
    .X(_08498_));
 sg13g2_buf_2 _15248_ (.A(\cpu.ex.pc[2] ),
    .X(_08499_));
 sg13g2_buf_2 _15249_ (.A(\cpu.ex.pc[3] ),
    .X(_08500_));
 sg13g2_nor2b_1 _15250_ (.A(\cpu.ex.pc[4] ),
    .B_N(_08500_),
    .Y(_08501_));
 sg13g2_buf_1 _15251_ (.A(\cpu.ex.pc[4] ),
    .X(_08502_));
 sg13g2_nand2b_1 _15252_ (.Y(_08503_),
    .B(net1141),
    .A_N(_08500_));
 sg13g2_o21ai_1 _15253_ (.B1(_08503_),
    .Y(_08504_),
    .A1(net1142),
    .A2(_08501_));
 sg13g2_nand2_1 _15254_ (.Y(_08505_),
    .A(_08498_),
    .B(_08504_));
 sg13g2_buf_1 _15255_ (.A(_08505_),
    .X(_08506_));
 sg13g2_buf_1 _15256_ (.A(_08506_),
    .X(_08507_));
 sg13g2_buf_1 _15257_ (.A(_08507_),
    .X(_08508_));
 sg13g2_buf_1 _15258_ (.A(net584),
    .X(_08509_));
 sg13g2_nor2b_1 _15259_ (.A(net1142),
    .B_N(_08500_),
    .Y(_08510_));
 sg13g2_nor2b_1 _15260_ (.A(net1141),
    .B_N(_08510_),
    .Y(_08511_));
 sg13g2_buf_2 _15261_ (.A(_08511_),
    .X(_08512_));
 sg13g2_buf_1 _15262_ (.A(_08512_),
    .X(_08513_));
 sg13g2_buf_1 _15263_ (.A(net725),
    .X(_08514_));
 sg13g2_inv_2 _15264_ (.Y(_08515_),
    .A(_08499_));
 sg13g2_nor3_1 _15265_ (.A(_08515_),
    .B(_08500_),
    .C(_08498_),
    .Y(_08516_));
 sg13g2_buf_1 _15266_ (.A(_08516_),
    .X(_08517_));
 sg13g2_buf_1 _15267_ (.A(net822),
    .X(_08518_));
 sg13g2_a22oi_1 _15268_ (.Y(_08519_),
    .B1(net724),
    .B2(\cpu.icache.r_tag[5][13] ),
    .A2(net643),
    .A1(\cpu.icache.r_tag[2][13] ));
 sg13g2_nor3_1 _15269_ (.A(_08515_),
    .B(_08500_),
    .C(net1141),
    .Y(_08520_));
 sg13g2_buf_2 _15270_ (.A(_08520_),
    .X(_08521_));
 sg13g2_buf_1 _15271_ (.A(_08521_),
    .X(_08522_));
 sg13g2_buf_1 _15272_ (.A(_08522_),
    .X(_08523_));
 sg13g2_inv_1 _15273_ (.Y(_08524_),
    .A(_08498_));
 sg13g2_buf_1 _15274_ (.A(_08524_),
    .X(_08525_));
 sg13g2_nand2_1 _15275_ (.Y(_08526_),
    .A(net1142),
    .B(_08500_));
 sg13g2_buf_2 _15276_ (.A(_08526_),
    .X(_08527_));
 sg13g2_nor2_1 _15277_ (.A(net939),
    .B(_08527_),
    .Y(_08528_));
 sg13g2_buf_1 _15278_ (.A(_08528_),
    .X(_08529_));
 sg13g2_buf_2 _15279_ (.A(net722),
    .X(_08530_));
 sg13g2_buf_1 _15280_ (.A(net641),
    .X(_08531_));
 sg13g2_a22oi_1 _15281_ (.Y(_08532_),
    .B1(_08531_),
    .B2(\cpu.icache.r_tag[3][13] ),
    .A2(net642),
    .A1(\cpu.icache.r_tag[1][13] ));
 sg13g2_buf_1 _15282_ (.A(_08498_),
    .X(_08533_));
 sg13g2_buf_1 _15283_ (.A(net1082),
    .X(_08534_));
 sg13g2_buf_1 _15284_ (.A(net938),
    .X(_08535_));
 sg13g2_buf_1 _15285_ (.A(net821),
    .X(_08536_));
 sg13g2_and2_1 _15286_ (.A(net1142),
    .B(_08500_),
    .X(_08537_));
 sg13g2_buf_1 _15287_ (.A(_08537_),
    .X(_08538_));
 sg13g2_buf_1 _15288_ (.A(net937),
    .X(_08539_));
 sg13g2_buf_1 _15289_ (.A(_08500_),
    .X(_08540_));
 sg13g2_buf_1 _15290_ (.A(net1081),
    .X(_08541_));
 sg13g2_buf_1 _15291_ (.A(net936),
    .X(_08542_));
 sg13g2_mux2_1 _15292_ (.A0(\cpu.icache.r_tag[4][13] ),
    .A1(\cpu.icache.r_tag[6][13] ),
    .S(net819),
    .X(_08543_));
 sg13g2_buf_1 _15293_ (.A(_08515_),
    .X(_08544_));
 sg13g2_a22oi_1 _15294_ (.Y(_08545_),
    .B1(_08543_),
    .B2(_08544_),
    .A2(_08539_),
    .A1(\cpu.icache.r_tag[7][13] ));
 sg13g2_or2_1 _15295_ (.X(_08546_),
    .B(_08545_),
    .A(_08536_));
 sg13g2_nand4_1 _15296_ (.B(_08519_),
    .C(_08532_),
    .A(net584),
    .Y(_08547_),
    .D(_08546_));
 sg13g2_o21ai_1 _15297_ (.B1(_08547_),
    .Y(_08548_),
    .A1(\cpu.icache.r_tag[0][13] ),
    .A2(net521));
 sg13g2_xnor2_1 _15298_ (.Y(_08549_),
    .A(net431),
    .B(_08548_));
 sg13g2_buf_1 _15299_ (.A(net942),
    .X(_08550_));
 sg13g2_mux4_1 _15300_ (.S0(net943),
    .A0(\cpu.genblk1.mmu.r_vtop_i[24][0] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[25][0] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[26][0] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[27][0] ),
    .S1(net824),
    .X(_08551_));
 sg13g2_mux4_1 _15301_ (.S0(net943),
    .A0(\cpu.genblk1.mmu.r_vtop_i[16][0] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[17][0] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[18][0] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[19][0] ),
    .S1(net824),
    .X(_08552_));
 sg13g2_mux4_1 _15302_ (.S0(net942),
    .A0(\cpu.genblk1.mmu.r_vtop_i[28][0] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[29][0] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[30][0] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[31][0] ),
    .S1(net825),
    .X(_08553_));
 sg13g2_mux4_1 _15303_ (.S0(net942),
    .A0(\cpu.genblk1.mmu.r_vtop_i[20][0] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[21][0] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[22][0] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[23][0] ),
    .S1(net825),
    .X(_08554_));
 sg13g2_mux4_1 _15304_ (.S0(net941),
    .A0(_08551_),
    .A1(_08552_),
    .A2(_08553_),
    .A3(_08554_),
    .S1(net940),
    .X(_08555_));
 sg13g2_nand2_1 _15305_ (.Y(_08556_),
    .A(net1146),
    .B(_08555_));
 sg13g2_mux4_1 _15306_ (.S0(net943),
    .A0(\cpu.genblk1.mmu.r_vtop_i[8][0] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[9][0] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[10][0] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[11][0] ),
    .S1(_08478_),
    .X(_08557_));
 sg13g2_mux4_1 _15307_ (.S0(_08477_),
    .A0(\cpu.genblk1.mmu.r_vtop_i[0][0] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[1][0] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[2][0] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[3][0] ),
    .S1(_08478_),
    .X(_08558_));
 sg13g2_mux4_1 _15308_ (.S0(_08481_),
    .A0(\cpu.genblk1.mmu.r_vtop_i[12][0] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[13][0] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[14][0] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[15][0] ),
    .S1(net825),
    .X(_08559_));
 sg13g2_mux4_1 _15309_ (.S0(_08481_),
    .A0(\cpu.genblk1.mmu.r_vtop_i[4][0] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[5][0] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[6][0] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[7][0] ),
    .S1(net825),
    .X(_08560_));
 sg13g2_mux4_1 _15310_ (.S0(net941),
    .A0(_08557_),
    .A1(_08558_),
    .A2(_08559_),
    .A3(_08560_),
    .S1(net940),
    .X(_08561_));
 sg13g2_nand2_1 _15311_ (.Y(_08562_),
    .A(net946),
    .B(_08561_));
 sg13g2_nand3_1 _15312_ (.B(_08556_),
    .C(_08562_),
    .A(net1083),
    .Y(_08563_));
 sg13g2_o21ai_1 _15313_ (.B1(_08563_),
    .Y(_08564_),
    .A1(net818),
    .A2(net1083));
 sg13g2_buf_2 _15314_ (.A(_08564_),
    .X(_08565_));
 sg13g2_nor2_2 _15315_ (.A(net1142),
    .B(_08498_),
    .Y(_08566_));
 sg13g2_and2_1 _15316_ (.A(net1081),
    .B(_08566_),
    .X(_08567_));
 sg13g2_buf_1 _15317_ (.A(_08567_),
    .X(_08568_));
 sg13g2_buf_1 _15318_ (.A(_08568_),
    .X(_08569_));
 sg13g2_a22oi_1 _15319_ (.Y(_08570_),
    .B1(net720),
    .B2(\cpu.icache.r_tag[6][12] ),
    .A2(net642),
    .A1(\cpu.icache.r_tag[1][12] ));
 sg13g2_a22oi_1 _15320_ (.Y(_08571_),
    .B1(net724),
    .B2(\cpu.icache.r_tag[5][12] ),
    .A2(net643),
    .A1(\cpu.icache.r_tag[2][12] ));
 sg13g2_nor3_1 _15321_ (.A(net1142),
    .B(_08540_),
    .C(net1082),
    .Y(_08572_));
 sg13g2_buf_1 _15322_ (.A(_08572_),
    .X(_08573_));
 sg13g2_buf_1 _15323_ (.A(_08573_),
    .X(_08574_));
 sg13g2_buf_2 _15324_ (.A(net938),
    .X(_08575_));
 sg13g2_mux2_1 _15325_ (.A0(\cpu.icache.r_tag[7][12] ),
    .A1(\cpu.icache.r_tag[3][12] ),
    .S(net817),
    .X(_08576_));
 sg13g2_a22oi_1 _15326_ (.Y(_08577_),
    .B1(_08576_),
    .B2(_08539_),
    .A2(net719),
    .A1(\cpu.icache.r_tag[4][12] ));
 sg13g2_nand4_1 _15327_ (.B(_08570_),
    .C(_08571_),
    .A(net584),
    .Y(_08578_),
    .D(_08577_));
 sg13g2_o21ai_1 _15328_ (.B1(_08578_),
    .Y(_08579_),
    .A1(\cpu.icache.r_tag[0][12] ),
    .A2(net521));
 sg13g2_xnor2_1 _15329_ (.Y(_08580_),
    .A(net430),
    .B(_08579_));
 sg13g2_nand2_1 _15330_ (.Y(_08581_),
    .A(_08549_),
    .B(_08580_));
 sg13g2_buf_2 _15331_ (.A(_00182_),
    .X(_08582_));
 sg13g2_buf_1 _15332_ (.A(_08582_),
    .X(_08583_));
 sg13g2_buf_1 _15333_ (.A(_08476_),
    .X(_08584_));
 sg13g2_buf_2 _15334_ (.A(net934),
    .X(_08585_));
 sg13g2_buf_1 _15335_ (.A(_08472_),
    .X(_08586_));
 sg13g2_buf_1 _15336_ (.A(net815),
    .X(_08587_));
 sg13g2_mux4_1 _15337_ (.S0(net816),
    .A0(\cpu.genblk1.mmu.r_vtop_i[24][6] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[25][6] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[26][6] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[27][6] ),
    .S1(net718),
    .X(_08588_));
 sg13g2_mux4_1 _15338_ (.S0(net816),
    .A0(\cpu.genblk1.mmu.r_vtop_i[16][6] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[17][6] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[18][6] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[19][6] ),
    .S1(net718),
    .X(_08589_));
 sg13g2_buf_2 _15339_ (.A(_08476_),
    .X(_08590_));
 sg13g2_buf_1 _15340_ (.A(net815),
    .X(_08591_));
 sg13g2_mux4_1 _15341_ (.S0(net933),
    .A0(\cpu.genblk1.mmu.r_vtop_i[28][6] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[29][6] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[30][6] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[31][6] ),
    .S1(net717),
    .X(_08592_));
 sg13g2_mux4_1 _15342_ (.S0(net933),
    .A0(\cpu.genblk1.mmu.r_vtop_i[20][6] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[21][6] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[22][6] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[23][6] ),
    .S1(net717),
    .X(_08593_));
 sg13g2_buf_2 _15343_ (.A(_08484_),
    .X(_08594_));
 sg13g2_mux4_1 _15344_ (.S0(net814),
    .A0(_08588_),
    .A1(_08589_),
    .A2(_08592_),
    .A3(_08593_),
    .S1(net940),
    .X(_08595_));
 sg13g2_mux4_1 _15345_ (.S0(net933),
    .A0(\cpu.genblk1.mmu.r_vtop_i[8][6] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[9][6] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[10][6] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[11][6] ),
    .S1(net717),
    .X(_08596_));
 sg13g2_mux4_1 _15346_ (.S0(net933),
    .A0(\cpu.genblk1.mmu.r_vtop_i[0][6] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[1][6] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[2][6] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[3][6] ),
    .S1(net717),
    .X(_08597_));
 sg13g2_mux4_1 _15347_ (.S0(_08590_),
    .A0(\cpu.genblk1.mmu.r_vtop_i[12][6] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[13][6] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[14][6] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[15][6] ),
    .S1(_08591_),
    .X(_08598_));
 sg13g2_mux4_1 _15348_ (.S0(_08590_),
    .A0(\cpu.genblk1.mmu.r_vtop_i[4][6] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[5][6] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[6][6] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[7][6] ),
    .S1(_08591_),
    .X(_08599_));
 sg13g2_mux4_1 _15349_ (.S0(net941),
    .A0(_08596_),
    .A1(_08597_),
    .A2(_08598_),
    .A3(_08599_),
    .S1(net940),
    .X(_08600_));
 sg13g2_mux2_1 _15350_ (.A0(_08595_),
    .A1(_08600_),
    .S(net823),
    .X(_08601_));
 sg13g2_nand2b_1 _15351_ (.Y(_08602_),
    .B(_08601_),
    .A_N(net1080));
 sg13g2_buf_2 _15352_ (.A(_08602_),
    .X(_08603_));
 sg13g2_buf_1 _15353_ (.A(_08506_),
    .X(_08604_));
 sg13g2_buf_1 _15354_ (.A(net640),
    .X(_08605_));
 sg13g2_buf_1 _15355_ (.A(net582),
    .X(_08606_));
 sg13g2_a22oi_1 _15356_ (.Y(_08607_),
    .B1(net642),
    .B2(\cpu.icache.r_tag[1][18] ),
    .A2(net643),
    .A1(\cpu.icache.r_tag[2][18] ));
 sg13g2_buf_1 _15357_ (.A(net1142),
    .X(_08608_));
 sg13g2_buf_2 _15358_ (.A(net1079),
    .X(_08609_));
 sg13g2_buf_1 _15359_ (.A(net936),
    .X(_08610_));
 sg13g2_buf_1 _15360_ (.A(_08610_),
    .X(_08611_));
 sg13g2_mux4_1 _15361_ (.S0(net932),
    .A0(\cpu.icache.r_tag[4][18] ),
    .A1(\cpu.icache.r_tag[5][18] ),
    .A2(\cpu.icache.r_tag[6][18] ),
    .A3(\cpu.icache.r_tag[7][18] ),
    .S1(net716),
    .X(_08612_));
 sg13g2_buf_1 _15362_ (.A(net939),
    .X(_08613_));
 sg13g2_buf_1 _15363_ (.A(net812),
    .X(_08614_));
 sg13g2_a22oi_1 _15364_ (.Y(_08615_),
    .B1(_08612_),
    .B2(_08614_),
    .A2(net583),
    .A1(\cpu.icache.r_tag[3][18] ));
 sg13g2_nand3_1 _15365_ (.B(_08607_),
    .C(_08615_),
    .A(net584),
    .Y(_08616_));
 sg13g2_o21ai_1 _15366_ (.B1(_08616_),
    .Y(_08617_),
    .A1(\cpu.icache.r_tag[0][18] ),
    .A2(net520));
 sg13g2_xnor2_1 _15367_ (.Y(_08618_),
    .A(net429),
    .B(_08617_));
 sg13g2_mux4_1 _15368_ (.S0(net818),
    .A0(\cpu.genblk1.mmu.r_vtop_i[24][5] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[25][5] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[26][5] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[27][5] ),
    .S1(net726),
    .X(_08619_));
 sg13g2_mux4_1 _15369_ (.S0(net818),
    .A0(\cpu.genblk1.mmu.r_vtop_i[16][5] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[17][5] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[18][5] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[19][5] ),
    .S1(net726),
    .X(_08620_));
 sg13g2_buf_2 _15370_ (.A(net934),
    .X(_08621_));
 sg13g2_buf_2 _15371_ (.A(net815),
    .X(_08622_));
 sg13g2_mux4_1 _15372_ (.S0(_08621_),
    .A0(\cpu.genblk1.mmu.r_vtop_i[28][5] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[29][5] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[30][5] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[31][5] ),
    .S1(_08622_),
    .X(_08623_));
 sg13g2_mux4_1 _15373_ (.S0(net811),
    .A0(\cpu.genblk1.mmu.r_vtop_i[20][5] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[21][5] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[22][5] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[23][5] ),
    .S1(net726),
    .X(_08624_));
 sg13g2_buf_1 _15374_ (.A(net1084),
    .X(_08625_));
 sg13g2_mux4_1 _15375_ (.S0(_08594_),
    .A0(_08619_),
    .A1(_08620_),
    .A2(_08623_),
    .A3(_08624_),
    .S1(net931),
    .X(_08626_));
 sg13g2_mux4_1 _15376_ (.S0(net818),
    .A0(\cpu.genblk1.mmu.r_vtop_i[8][5] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[9][5] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[10][5] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[11][5] ),
    .S1(net726),
    .X(_08627_));
 sg13g2_mux4_1 _15377_ (.S0(net818),
    .A0(\cpu.genblk1.mmu.r_vtop_i[0][5] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[1][5] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[2][5] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[3][5] ),
    .S1(net726),
    .X(_08628_));
 sg13g2_mux4_1 _15378_ (.S0(net811),
    .A0(\cpu.genblk1.mmu.r_vtop_i[12][5] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[13][5] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[14][5] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[15][5] ),
    .S1(net714),
    .X(_08629_));
 sg13g2_mux4_1 _15379_ (.S0(_08621_),
    .A0(\cpu.genblk1.mmu.r_vtop_i[4][5] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[5][5] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[6][5] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[7][5] ),
    .S1(_08622_),
    .X(_08630_));
 sg13g2_mux4_1 _15380_ (.S0(_08594_),
    .A0(_08627_),
    .A1(_08628_),
    .A2(_08629_),
    .A3(_08630_),
    .S1(net931),
    .X(_08631_));
 sg13g2_mux2_1 _15381_ (.A0(_08626_),
    .A1(_08631_),
    .S(net823),
    .X(_08632_));
 sg13g2_nand2b_1 _15382_ (.Y(_08633_),
    .B(_08632_),
    .A_N(net1080));
 sg13g2_buf_1 _15383_ (.A(_08633_),
    .X(_08634_));
 sg13g2_nand2_1 _15384_ (.Y(_08635_),
    .A(\cpu.icache.r_tag[4][17] ),
    .B(net719));
 sg13g2_buf_1 _15385_ (.A(_08521_),
    .X(_08636_));
 sg13g2_buf_1 _15386_ (.A(net713),
    .X(_08637_));
 sg13g2_nor2_1 _15387_ (.A(net1082),
    .B(_08527_),
    .Y(_08638_));
 sg13g2_buf_2 _15388_ (.A(_08638_),
    .X(_08639_));
 sg13g2_a22oi_1 _15389_ (.Y(_08640_),
    .B1(_08639_),
    .B2(\cpu.icache.r_tag[7][17] ),
    .A2(net639),
    .A1(\cpu.icache.r_tag[1][17] ));
 sg13g2_buf_1 _15390_ (.A(_08512_),
    .X(_08641_));
 sg13g2_buf_1 _15391_ (.A(net712),
    .X(_08642_));
 sg13g2_a22oi_1 _15392_ (.Y(_08643_),
    .B1(net724),
    .B2(\cpu.icache.r_tag[5][17] ),
    .A2(net638),
    .A1(\cpu.icache.r_tag[2][17] ));
 sg13g2_a22oi_1 _15393_ (.Y(_08644_),
    .B1(net720),
    .B2(\cpu.icache.r_tag[6][17] ),
    .A2(net641),
    .A1(\cpu.icache.r_tag[3][17] ));
 sg13g2_nand4_1 _15394_ (.B(_08640_),
    .C(_08643_),
    .A(_08635_),
    .Y(_08645_),
    .D(_08644_));
 sg13g2_mux2_1 _15395_ (.A0(\cpu.icache.r_tag[0][17] ),
    .A1(_08645_),
    .S(net520),
    .X(_08646_));
 sg13g2_xor2_1 _15396_ (.B(_08646_),
    .A(_08634_),
    .X(_08647_));
 sg13g2_mux4_1 _15397_ (.S0(net933),
    .A0(\cpu.genblk1.mmu.r_vtop_i[16][3] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[17][3] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[18][3] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[19][3] ),
    .S1(net717),
    .X(_08648_));
 sg13g2_mux4_1 _15398_ (.S0(net933),
    .A0(\cpu.genblk1.mmu.r_vtop_i[0][3] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[1][3] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[2][3] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[3][3] ),
    .S1(net717),
    .X(_08649_));
 sg13g2_mux4_1 _15399_ (.S0(net943),
    .A0(\cpu.genblk1.mmu.r_vtop_i[20][3] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[21][3] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[22][3] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[23][3] ),
    .S1(net824),
    .X(_08650_));
 sg13g2_mux4_1 _15400_ (.S0(_08477_),
    .A0(\cpu.genblk1.mmu.r_vtop_i[4][3] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[5][3] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[6][3] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[7][3] ),
    .S1(net717),
    .X(_08651_));
 sg13g2_mux4_1 _15401_ (.S0(net946),
    .A0(_08648_),
    .A1(_08649_),
    .A2(_08650_),
    .A3(_08651_),
    .S1(_08485_),
    .X(_08652_));
 sg13g2_a21oi_1 _15402_ (.A1(net1083),
    .A2(_08652_),
    .Y(_08653_),
    .B1(_08397_));
 sg13g2_mux4_1 _15403_ (.S0(net816),
    .A0(\cpu.genblk1.mmu.r_vtop_i[24][3] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[25][3] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[26][3] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[27][3] ),
    .S1(net718),
    .X(_08654_));
 sg13g2_buf_2 _15404_ (.A(_08584_),
    .X(_08655_));
 sg13g2_buf_1 _15405_ (.A(net815),
    .X(_08656_));
 sg13g2_mux4_1 _15406_ (.S0(net810),
    .A0(\cpu.genblk1.mmu.r_vtop_i[8][3] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[9][3] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[10][3] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[11][3] ),
    .S1(net711),
    .X(_08657_));
 sg13g2_mux4_1 _15407_ (.S0(net816),
    .A0(\cpu.genblk1.mmu.r_vtop_i[28][3] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[29][3] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[30][3] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[31][3] ),
    .S1(net718),
    .X(_08658_));
 sg13g2_mux4_1 _15408_ (.S0(_08585_),
    .A0(\cpu.genblk1.mmu.r_vtop_i[12][3] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[13][3] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[14][3] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[15][3] ),
    .S1(net718),
    .X(_08659_));
 sg13g2_mux4_1 _15409_ (.S0(net946),
    .A0(_08654_),
    .A1(_08657_),
    .A2(_08658_),
    .A3(_08659_),
    .S1(net940),
    .X(_08660_));
 sg13g2_nor3_1 _15410_ (.A(net814),
    .B(_08339_),
    .C(_08660_),
    .Y(_08661_));
 sg13g2_or2_1 _15411_ (.X(_08662_),
    .B(_08661_),
    .A(_08653_));
 sg13g2_buf_2 _15412_ (.A(_08662_),
    .X(_08663_));
 sg13g2_and2_1 _15413_ (.A(\cpu.icache.r_tag[7][15] ),
    .B(_08639_),
    .X(_08664_));
 sg13g2_a221oi_1 _15414_ (.B2(\cpu.icache.r_tag[5][15] ),
    .C1(_08664_),
    .B1(net822),
    .A1(\cpu.icache.r_tag[2][15] ),
    .Y(_08665_),
    .A2(net638));
 sg13g2_a22oi_1 _15415_ (.Y(_08666_),
    .B1(net719),
    .B2(\cpu.icache.r_tag[4][15] ),
    .A2(net639),
    .A1(\cpu.icache.r_tag[1][15] ));
 sg13g2_a22oi_1 _15416_ (.Y(_08667_),
    .B1(net720),
    .B2(\cpu.icache.r_tag[6][15] ),
    .A2(_08531_),
    .A1(\cpu.icache.r_tag[3][15] ));
 sg13g2_nand4_1 _15417_ (.B(_08665_),
    .C(_08666_),
    .A(net584),
    .Y(_08668_),
    .D(_08667_));
 sg13g2_o21ai_1 _15418_ (.B1(_08668_),
    .Y(_08669_),
    .A1(\cpu.icache.r_tag[0][15] ),
    .A2(net520));
 sg13g2_xnor2_1 _15419_ (.Y(_08670_),
    .A(net428),
    .B(_08669_));
 sg13g2_buf_2 _15420_ (.A(\cpu.ex.pc[5] ),
    .X(_08671_));
 sg13g2_mux4_1 _15421_ (.S0(net1079),
    .A0(\cpu.icache.r_tag[4][5] ),
    .A1(\cpu.icache.r_tag[5][5] ),
    .A2(\cpu.icache.r_tag[6][5] ),
    .A3(\cpu.icache.r_tag[7][5] ),
    .S1(net819),
    .X(_08672_));
 sg13g2_nand2_1 _15422_ (.Y(_08673_),
    .A(_08613_),
    .B(_08672_));
 sg13g2_nand2_1 _15423_ (.Y(_08674_),
    .A(\cpu.icache.r_tag[1][5] ),
    .B(net713));
 sg13g2_a22oi_1 _15424_ (.Y(_08675_),
    .B1(net722),
    .B2(\cpu.icache.r_tag[3][5] ),
    .A2(net712),
    .A1(\cpu.icache.r_tag[2][5] ));
 sg13g2_nand4_1 _15425_ (.B(_08673_),
    .C(_08674_),
    .A(net640),
    .Y(_08676_),
    .D(_08675_));
 sg13g2_o21ai_1 _15426_ (.B1(_08676_),
    .Y(_08677_),
    .A1(\cpu.icache.r_tag[0][5] ),
    .A2(net644));
 sg13g2_xor2_1 _15427_ (.B(_08677_),
    .A(_08671_),
    .X(_08678_));
 sg13g2_buf_1 _15428_ (.A(\cpu.ex.pc[9] ),
    .X(_08679_));
 sg13g2_mux4_1 _15429_ (.S0(net1079),
    .A0(\cpu.icache.r_tag[4][9] ),
    .A1(\cpu.icache.r_tag[5][9] ),
    .A2(\cpu.icache.r_tag[6][9] ),
    .A3(\cpu.icache.r_tag[7][9] ),
    .S1(net819),
    .X(_08680_));
 sg13g2_nand2_1 _15430_ (.Y(_08681_),
    .A(net939),
    .B(_08680_));
 sg13g2_nand2_1 _15431_ (.Y(_08682_),
    .A(\cpu.icache.r_tag[1][9] ),
    .B(net713));
 sg13g2_a22oi_1 _15432_ (.Y(_08683_),
    .B1(net722),
    .B2(\cpu.icache.r_tag[3][9] ),
    .A2(_08512_),
    .A1(\cpu.icache.r_tag[2][9] ));
 sg13g2_nand4_1 _15433_ (.B(_08681_),
    .C(_08682_),
    .A(net640),
    .Y(_08684_),
    .D(_08683_));
 sg13g2_o21ai_1 _15434_ (.B1(_08684_),
    .Y(_08685_),
    .A1(\cpu.icache.r_tag[0][9] ),
    .A2(net644));
 sg13g2_xor2_1 _15435_ (.B(_08685_),
    .A(_08679_),
    .X(_08686_));
 sg13g2_nand2_1 _15436_ (.Y(_08687_),
    .A(_08678_),
    .B(_08686_));
 sg13g2_buf_1 _15437_ (.A(\cpu.ex.pc[10] ),
    .X(_08688_));
 sg13g2_nand2_1 _15438_ (.Y(_08689_),
    .A(\cpu.icache.r_tag[2][10] ),
    .B(_08513_));
 sg13g2_a22oi_1 _15439_ (.Y(_08690_),
    .B1(_08639_),
    .B2(\cpu.icache.r_tag[7][10] ),
    .A2(_08573_),
    .A1(\cpu.icache.r_tag[4][10] ));
 sg13g2_nand3_1 _15440_ (.B(net1082),
    .C(\cpu.icache.r_tag[3][10] ),
    .A(_08542_),
    .Y(_08691_));
 sg13g2_nor2_2 _15441_ (.A(net1081),
    .B(net1082),
    .Y(_08692_));
 sg13g2_nand2_1 _15442_ (.Y(_08693_),
    .A(\cpu.icache.r_tag[5][10] ),
    .B(_08692_));
 sg13g2_a21oi_1 _15443_ (.A1(_08691_),
    .A2(_08693_),
    .Y(_08694_),
    .B1(_08544_));
 sg13g2_a221oi_1 _15444_ (.B2(\cpu.icache.r_tag[6][10] ),
    .C1(_08694_),
    .B1(_08568_),
    .A1(\cpu.icache.r_tag[1][10] ),
    .Y(_08695_),
    .A2(_08636_));
 sg13g2_nand4_1 _15445_ (.B(_08689_),
    .C(_08690_),
    .A(_08507_),
    .Y(_08696_),
    .D(_08695_));
 sg13g2_o21ai_1 _15446_ (.B1(_08696_),
    .Y(_08697_),
    .A1(\cpu.icache.r_tag[0][10] ),
    .A2(net582));
 sg13g2_xnor2_1 _15447_ (.Y(_08698_),
    .A(_08688_),
    .B(_08697_));
 sg13g2_buf_1 _15448_ (.A(\cpu.ex.pc[7] ),
    .X(_08699_));
 sg13g2_a22oi_1 _15449_ (.Y(_08700_),
    .B1(_08573_),
    .B2(\cpu.icache.r_tag[4][7] ),
    .A2(net725),
    .A1(\cpu.icache.r_tag[2][7] ));
 sg13g2_a22oi_1 _15450_ (.Y(_08701_),
    .B1(net722),
    .B2(\cpu.icache.r_tag[3][7] ),
    .A2(_08522_),
    .A1(\cpu.icache.r_tag[1][7] ));
 sg13g2_mux2_1 _15451_ (.A0(\cpu.icache.r_tag[5][7] ),
    .A1(\cpu.icache.r_tag[7][7] ),
    .S(net936),
    .X(_08702_));
 sg13g2_a22oi_1 _15452_ (.Y(_08703_),
    .B1(_08702_),
    .B2(_08608_),
    .A2(_08510_),
    .A1(\cpu.icache.r_tag[6][7] ));
 sg13g2_or2_1 _15453_ (.X(_08704_),
    .B(_08703_),
    .A(net817));
 sg13g2_nand3_1 _15454_ (.B(_08701_),
    .C(_08704_),
    .A(_08700_),
    .Y(_08705_));
 sg13g2_mux2_1 _15455_ (.A0(\cpu.icache.r_tag[0][7] ),
    .A1(_08705_),
    .S(_08605_),
    .X(_08706_));
 sg13g2_xor2_1 _15456_ (.B(_08706_),
    .A(_08699_),
    .X(_08707_));
 sg13g2_inv_1 _15457_ (.Y(_08708_),
    .A(\cpu.ex.pc[8] ));
 sg13g2_buf_1 _15458_ (.A(_08708_),
    .X(_08709_));
 sg13g2_a22oi_1 _15459_ (.Y(_08710_),
    .B1(_08517_),
    .B2(\cpu.icache.r_tag[5][8] ),
    .A2(net712),
    .A1(\cpu.icache.r_tag[2][8] ));
 sg13g2_a22oi_1 _15460_ (.Y(_08711_),
    .B1(_08529_),
    .B2(\cpu.icache.r_tag[3][8] ),
    .A2(net713),
    .A1(\cpu.icache.r_tag[1][8] ));
 sg13g2_mux2_1 _15461_ (.A0(\cpu.icache.r_tag[4][8] ),
    .A1(\cpu.icache.r_tag[6][8] ),
    .S(net1081),
    .X(_08712_));
 sg13g2_a22oi_1 _15462_ (.Y(_08713_),
    .B1(_08712_),
    .B2(_08515_),
    .A2(_08538_),
    .A1(\cpu.icache.r_tag[7][8] ));
 sg13g2_or2_1 _15463_ (.X(_08714_),
    .B(_08713_),
    .A(_08534_));
 sg13g2_nand4_1 _15464_ (.B(_08710_),
    .C(_08711_),
    .A(net644),
    .Y(_08715_),
    .D(_08714_));
 sg13g2_o21ai_1 _15465_ (.B1(_08715_),
    .Y(_08716_),
    .A1(\cpu.icache.r_tag[0][8] ),
    .A2(net644));
 sg13g2_xnor2_1 _15466_ (.Y(_08717_),
    .A(net1078),
    .B(_08716_));
 sg13g2_buf_1 _15467_ (.A(\cpu.ex.pc[6] ),
    .X(_08718_));
 sg13g2_a22oi_1 _15468_ (.Y(_08719_),
    .B1(_08568_),
    .B2(\cpu.icache.r_tag[6][6] ),
    .A2(_08636_),
    .A1(\cpu.icache.r_tag[1][6] ));
 sg13g2_a22oi_1 _15469_ (.Y(_08720_),
    .B1(_08573_),
    .B2(\cpu.icache.r_tag[4][6] ),
    .A2(_08641_),
    .A1(\cpu.icache.r_tag[2][6] ));
 sg13g2_mux2_1 _15470_ (.A0(\cpu.icache.r_tag[7][6] ),
    .A1(\cpu.icache.r_tag[3][6] ),
    .S(net1082),
    .X(_08721_));
 sg13g2_a22oi_1 _15471_ (.Y(_08722_),
    .B1(_08721_),
    .B2(_08542_),
    .A2(_08692_),
    .A1(\cpu.icache.r_tag[5][6] ));
 sg13g2_nand2b_1 _15472_ (.Y(_08723_),
    .B(net932),
    .A_N(_08722_));
 sg13g2_nand4_1 _15473_ (.B(_08719_),
    .C(_08720_),
    .A(_08604_),
    .Y(_08724_),
    .D(_08723_));
 sg13g2_o21ai_1 _15474_ (.B1(_08724_),
    .Y(_08725_),
    .A1(\cpu.icache.r_tag[0][6] ),
    .A2(net644));
 sg13g2_xor2_1 _15475_ (.B(_08725_),
    .A(_08718_),
    .X(_08726_));
 sg13g2_mux4_1 _15476_ (.S0(net932),
    .A0(\cpu.icache.r_valid[0] ),
    .A1(\cpu.icache.r_valid[1] ),
    .A2(\cpu.icache.r_valid[2] ),
    .A3(\cpu.icache.r_valid[3] ),
    .S1(net716),
    .X(_08727_));
 sg13g2_mux4_1 _15477_ (.S0(net932),
    .A0(\cpu.icache.r_valid[4] ),
    .A1(\cpu.icache.r_valid[5] ),
    .A2(\cpu.icache.r_valid[6] ),
    .A3(\cpu.icache.r_valid[7] ),
    .S1(net716),
    .X(_08728_));
 sg13g2_mux2_1 _15478_ (.A0(_08727_),
    .A1(_08728_),
    .S(_08502_),
    .X(_08729_));
 sg13g2_inv_1 _15479_ (.Y(_08730_),
    .A(\cpu.ex.pc[11] ));
 sg13g2_buf_1 _15480_ (.A(_08730_),
    .X(_08731_));
 sg13g2_a22oi_1 _15481_ (.Y(_08732_),
    .B1(_08568_),
    .B2(\cpu.icache.r_tag[6][11] ),
    .A2(_08641_),
    .A1(\cpu.icache.r_tag[2][11] ));
 sg13g2_a22oi_1 _15482_ (.Y(_08733_),
    .B1(_08529_),
    .B2(\cpu.icache.r_tag[3][11] ),
    .A2(_08521_),
    .A1(\cpu.icache.r_tag[1][11] ));
 sg13g2_nor2_2 _15483_ (.A(net1142),
    .B(net1081),
    .Y(_08734_));
 sg13g2_mux2_1 _15484_ (.A0(\cpu.icache.r_tag[5][11] ),
    .A1(\cpu.icache.r_tag[7][11] ),
    .S(_08540_),
    .X(_08735_));
 sg13g2_a22oi_1 _15485_ (.Y(_08736_),
    .B1(_08735_),
    .B2(net1079),
    .A2(_08734_),
    .A1(\cpu.icache.r_tag[4][11] ));
 sg13g2_or2_1 _15486_ (.X(_08737_),
    .B(_08736_),
    .A(_08534_));
 sg13g2_nand4_1 _15487_ (.B(_08732_),
    .C(_08733_),
    .A(_08604_),
    .Y(_08738_),
    .D(_08737_));
 sg13g2_o21ai_1 _15488_ (.B1(_08738_),
    .Y(_08739_),
    .A1(\cpu.icache.r_tag[0][11] ),
    .A2(net644));
 sg13g2_xnor2_1 _15489_ (.Y(_08740_),
    .A(net1077),
    .B(_08739_));
 sg13g2_nand4_1 _15490_ (.B(_08726_),
    .C(_08729_),
    .A(_08717_),
    .Y(_08741_),
    .D(_08740_));
 sg13g2_nor4_1 _15491_ (.A(_08687_),
    .B(_08698_),
    .C(_08707_),
    .D(_08741_),
    .Y(_08742_));
 sg13g2_nand4_1 _15492_ (.B(_08647_),
    .C(_08670_),
    .A(_08618_),
    .Y(_08743_),
    .D(_08742_));
 sg13g2_buf_2 _15493_ (.A(_08476_),
    .X(_08744_));
 sg13g2_buf_1 _15494_ (.A(net944),
    .X(_08745_));
 sg13g2_mux4_1 _15495_ (.S0(net930),
    .A0(\cpu.genblk1.mmu.r_vtop_i[24][4] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[25][4] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[26][4] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[27][4] ),
    .S1(net809),
    .X(_08746_));
 sg13g2_mux4_1 _15496_ (.S0(net930),
    .A0(\cpu.genblk1.mmu.r_vtop_i[16][4] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[17][4] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[18][4] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[19][4] ),
    .S1(net809),
    .X(_08747_));
 sg13g2_mux4_1 _15497_ (.S0(net934),
    .A0(\cpu.genblk1.mmu.r_vtop_i[28][4] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[29][4] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[30][4] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[31][4] ),
    .S1(net815),
    .X(_08748_));
 sg13g2_mux4_1 _15498_ (.S0(net934),
    .A0(\cpu.genblk1.mmu.r_vtop_i[20][4] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[21][4] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[22][4] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[23][4] ),
    .S1(net815),
    .X(_08749_));
 sg13g2_mux4_1 _15499_ (.S0(net941),
    .A0(_08746_),
    .A1(_08747_),
    .A2(_08748_),
    .A3(_08749_),
    .S1(net1084),
    .X(_08750_));
 sg13g2_mux4_1 _15500_ (.S0(net934),
    .A0(\cpu.genblk1.mmu.r_vtop_i[8][4] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[9][4] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[10][4] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[11][4] ),
    .S1(net809),
    .X(_08751_));
 sg13g2_mux4_1 _15501_ (.S0(net930),
    .A0(\cpu.genblk1.mmu.r_vtop_i[0][4] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[1][4] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[2][4] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[3][4] ),
    .S1(net809),
    .X(_08752_));
 sg13g2_mux4_1 _15502_ (.S0(net934),
    .A0(\cpu.genblk1.mmu.r_vtop_i[12][4] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[13][4] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[14][4] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[15][4] ),
    .S1(net815),
    .X(_08753_));
 sg13g2_mux4_1 _15503_ (.S0(net934),
    .A0(\cpu.genblk1.mmu.r_vtop_i[4][4] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[5][4] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[6][4] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[7][4] ),
    .S1(_08586_),
    .X(_08754_));
 sg13g2_mux4_1 _15504_ (.S0(_08484_),
    .A0(_08751_),
    .A1(_08752_),
    .A2(_08753_),
    .A3(_08754_),
    .S1(net1084),
    .X(_08755_));
 sg13g2_mux2_1 _15505_ (.A0(_08750_),
    .A1(_08755_),
    .S(net946),
    .X(_08756_));
 sg13g2_nand2b_1 _15506_ (.Y(_08757_),
    .B(_08756_),
    .A_N(net1080));
 sg13g2_buf_2 _15507_ (.A(_08757_),
    .X(_08758_));
 sg13g2_mux4_1 _15508_ (.S0(_08609_),
    .A0(\cpu.icache.r_tag[4][16] ),
    .A1(\cpu.icache.r_tag[5][16] ),
    .A2(\cpu.icache.r_tag[6][16] ),
    .A3(\cpu.icache.r_tag[7][16] ),
    .S1(net813),
    .X(_08759_));
 sg13g2_nand2_1 _15509_ (.Y(_08760_),
    .A(_08613_),
    .B(_08759_));
 sg13g2_nand2_1 _15510_ (.Y(_08761_),
    .A(\cpu.icache.r_tag[1][16] ),
    .B(net639));
 sg13g2_a22oi_1 _15511_ (.Y(_08762_),
    .B1(net641),
    .B2(\cpu.icache.r_tag[3][16] ),
    .A2(net638),
    .A1(\cpu.icache.r_tag[2][16] ));
 sg13g2_nand4_1 _15512_ (.B(_08760_),
    .C(_08761_),
    .A(_08605_),
    .Y(_08763_),
    .D(_08762_));
 sg13g2_o21ai_1 _15513_ (.B1(_08763_),
    .Y(_08764_),
    .A1(\cpu.icache.r_tag[0][16] ),
    .A2(net584));
 sg13g2_xor2_1 _15514_ (.B(_08764_),
    .A(_08758_),
    .X(_08765_));
 sg13g2_mux4_1 _15515_ (.S0(net930),
    .A0(\cpu.genblk1.mmu.r_vtop_i[24][9] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[25][9] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[26][9] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[27][9] ),
    .S1(_08473_),
    .X(_08766_));
 sg13g2_mux4_1 _15516_ (.S0(net942),
    .A0(\cpu.genblk1.mmu.r_vtop_i[16][9] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[17][9] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[18][9] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[19][9] ),
    .S1(_08473_),
    .X(_08767_));
 sg13g2_mux4_1 _15517_ (.S0(net930),
    .A0(\cpu.genblk1.mmu.r_vtop_i[28][9] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[29][9] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[30][9] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[31][9] ),
    .S1(net809),
    .X(_08768_));
 sg13g2_mux4_1 _15518_ (.S0(net930),
    .A0(\cpu.genblk1.mmu.r_vtop_i[20][9] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[21][9] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[22][9] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[23][9] ),
    .S1(net809),
    .X(_08769_));
 sg13g2_mux4_1 _15519_ (.S0(net941),
    .A0(_08766_),
    .A1(_08767_),
    .A2(_08768_),
    .A3(_08769_),
    .S1(_08485_),
    .X(_08770_));
 sg13g2_mux4_1 _15520_ (.S0(net930),
    .A0(\cpu.genblk1.mmu.r_vtop_i[8][9] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[9][9] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[10][9] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[11][9] ),
    .S1(_08745_),
    .X(_08771_));
 sg13g2_mux4_1 _15521_ (.S0(_08744_),
    .A0(\cpu.genblk1.mmu.r_vtop_i[0][9] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[1][9] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[2][9] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[3][9] ),
    .S1(net809),
    .X(_08772_));
 sg13g2_mux4_1 _15522_ (.S0(net930),
    .A0(\cpu.genblk1.mmu.r_vtop_i[12][9] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[13][9] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[14][9] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[15][9] ),
    .S1(net809),
    .X(_08773_));
 sg13g2_mux4_1 _15523_ (.S0(_08744_),
    .A0(\cpu.genblk1.mmu.r_vtop_i[4][9] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[5][9] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[6][9] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[7][9] ),
    .S1(_08745_),
    .X(_08774_));
 sg13g2_mux4_1 _15524_ (.S0(net941),
    .A0(_08771_),
    .A1(_08772_),
    .A2(_08773_),
    .A3(_08774_),
    .S1(net1084),
    .X(_08775_));
 sg13g2_mux2_1 _15525_ (.A0(_08770_),
    .A1(_08775_),
    .S(net946),
    .X(_08776_));
 sg13g2_nand2b_1 _15526_ (.Y(_08777_),
    .B(_08776_),
    .A_N(net1080));
 sg13g2_buf_1 _15527_ (.A(_08777_),
    .X(_08778_));
 sg13g2_a22oi_1 _15528_ (.Y(_08779_),
    .B1(_08637_),
    .B2(\cpu.icache.r_tag[1][21] ),
    .A2(_08642_),
    .A1(\cpu.icache.r_tag[2][21] ));
 sg13g2_mux2_1 _15529_ (.A0(\cpu.icache.r_tag[4][21] ),
    .A1(\cpu.icache.r_tag[6][21] ),
    .S(net813),
    .X(_08780_));
 sg13g2_a22oi_1 _15530_ (.Y(_08781_),
    .B1(_08566_),
    .B2(_08780_),
    .A2(net641),
    .A1(\cpu.icache.r_tag[3][21] ));
 sg13g2_a22oi_1 _15531_ (.Y(_08782_),
    .B1(_08639_),
    .B2(\cpu.icache.r_tag[7][21] ),
    .A2(_08517_),
    .A1(\cpu.icache.r_tag[5][21] ));
 sg13g2_nand4_1 _15532_ (.B(_08779_),
    .C(_08781_),
    .A(_08508_),
    .Y(_08783_),
    .D(_08782_));
 sg13g2_o21ai_1 _15533_ (.B1(_08783_),
    .Y(_08784_),
    .A1(\cpu.icache.r_tag[0][21] ),
    .A2(_08508_));
 sg13g2_xor2_1 _15534_ (.B(_08784_),
    .A(net464),
    .X(_08785_));
 sg13g2_nor2_1 _15535_ (.A(_08765_),
    .B(_08785_),
    .Y(_08786_));
 sg13g2_mux4_1 _15536_ (.S0(_08476_),
    .A0(\cpu.genblk1.mmu.r_vtop_i[24][11] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[25][11] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[26][11] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[27][11] ),
    .S1(net944),
    .X(_08787_));
 sg13g2_mux4_1 _15537_ (.S0(_08476_),
    .A0(\cpu.genblk1.mmu.r_vtop_i[16][11] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[17][11] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[18][11] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[19][11] ),
    .S1(net944),
    .X(_08788_));
 sg13g2_mux4_1 _15538_ (.S0(net1147),
    .A0(\cpu.genblk1.mmu.r_vtop_i[28][11] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[29][11] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[30][11] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[31][11] ),
    .S1(net1085),
    .X(_08789_));
 sg13g2_mux4_1 _15539_ (.S0(net1147),
    .A0(\cpu.genblk1.mmu.r_vtop_i[20][11] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[21][11] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[22][11] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[23][11] ),
    .S1(net944),
    .X(_08790_));
 sg13g2_mux4_1 _15540_ (.S0(_08418_),
    .A0(_08787_),
    .A1(_08788_),
    .A2(_08789_),
    .A3(_08790_),
    .S1(net1084),
    .X(_08791_));
 sg13g2_mux4_1 _15541_ (.S0(net1147),
    .A0(\cpu.genblk1.mmu.r_vtop_i[8][11] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[9][11] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[10][11] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[11][11] ),
    .S1(net944),
    .X(_08792_));
 sg13g2_mux4_1 _15542_ (.S0(_08476_),
    .A0(\cpu.genblk1.mmu.r_vtop_i[0][11] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[1][11] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[2][11] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[3][11] ),
    .S1(net944),
    .X(_08793_));
 sg13g2_mux4_1 _15543_ (.S0(net1147),
    .A0(\cpu.genblk1.mmu.r_vtop_i[12][11] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[13][11] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[14][11] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[15][11] ),
    .S1(net1085),
    .X(_08794_));
 sg13g2_mux4_1 _15544_ (.S0(net1147),
    .A0(\cpu.genblk1.mmu.r_vtop_i[4][11] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[5][11] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[6][11] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[7][11] ),
    .S1(net1085),
    .X(_08795_));
 sg13g2_mux4_1 _15545_ (.S0(_08418_),
    .A0(_08792_),
    .A1(_08793_),
    .A2(_08794_),
    .A3(_08795_),
    .S1(net1084),
    .X(_08796_));
 sg13g2_mux2_1 _15546_ (.A0(_08791_),
    .A1(_08796_),
    .S(_08405_),
    .X(_08797_));
 sg13g2_nand2b_1 _15547_ (.Y(_08798_),
    .B(_08797_),
    .A_N(net1080));
 sg13g2_buf_2 _15548_ (.A(_08798_),
    .X(_08799_));
 sg13g2_buf_1 _15549_ (.A(net638),
    .X(_08800_));
 sg13g2_mux4_1 _15550_ (.S0(_08609_),
    .A0(\cpu.icache.r_tag[4][23] ),
    .A1(\cpu.icache.r_tag[5][23] ),
    .A2(\cpu.icache.r_tag[6][23] ),
    .A3(\cpu.icache.r_tag[7][23] ),
    .S1(net716),
    .X(_08801_));
 sg13g2_a22oi_1 _15551_ (.Y(_08802_),
    .B1(_08530_),
    .B2(\cpu.icache.r_tag[3][23] ),
    .A2(_08637_),
    .A1(\cpu.icache.r_tag[1][23] ));
 sg13g2_inv_1 _15552_ (.Y(_08803_),
    .A(_08802_));
 sg13g2_a221oi_1 _15553_ (.B2(_08614_),
    .C1(_08803_),
    .B1(_08801_),
    .A1(\cpu.icache.r_tag[2][23] ),
    .Y(_08804_),
    .A2(_08800_));
 sg13g2_nor2_1 _15554_ (.A(\cpu.icache.r_tag[0][23] ),
    .B(net520),
    .Y(_08805_));
 sg13g2_a21oi_1 _15555_ (.A1(net521),
    .A2(_08804_),
    .Y(_08806_),
    .B1(_08805_));
 sg13g2_xor2_1 _15556_ (.B(_08806_),
    .A(net519),
    .X(_08807_));
 sg13g2_mux4_1 _15557_ (.S0(net816),
    .A0(\cpu.genblk1.mmu.r_vtop_i[24][7] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[25][7] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[26][7] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[27][7] ),
    .S1(net711),
    .X(_08808_));
 sg13g2_mux4_1 _15558_ (.S0(net810),
    .A0(\cpu.genblk1.mmu.r_vtop_i[16][7] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[17][7] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[18][7] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[19][7] ),
    .S1(net711),
    .X(_08809_));
 sg13g2_mux4_1 _15559_ (.S0(net816),
    .A0(\cpu.genblk1.mmu.r_vtop_i[28][7] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[29][7] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[30][7] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[31][7] ),
    .S1(net718),
    .X(_08810_));
 sg13g2_mux4_1 _15560_ (.S0(net816),
    .A0(\cpu.genblk1.mmu.r_vtop_i[20][7] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[21][7] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[22][7] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[23][7] ),
    .S1(net718),
    .X(_08811_));
 sg13g2_mux4_1 _15561_ (.S0(net814),
    .A0(_08808_),
    .A1(_08809_),
    .A2(_08810_),
    .A3(_08811_),
    .S1(net931),
    .X(_08812_));
 sg13g2_mux4_1 _15562_ (.S0(_08585_),
    .A0(\cpu.genblk1.mmu.r_vtop_i[8][7] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[9][7] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[10][7] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[11][7] ),
    .S1(_08587_),
    .X(_08813_));
 sg13g2_mux4_1 _15563_ (.S0(net816),
    .A0(\cpu.genblk1.mmu.r_vtop_i[0][7] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[1][7] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[2][7] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[3][7] ),
    .S1(net718),
    .X(_08814_));
 sg13g2_mux4_1 _15564_ (.S0(net933),
    .A0(\cpu.genblk1.mmu.r_vtop_i[12][7] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[13][7] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[14][7] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[15][7] ),
    .S1(net717),
    .X(_08815_));
 sg13g2_mux4_1 _15565_ (.S0(net933),
    .A0(\cpu.genblk1.mmu.r_vtop_i[4][7] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[5][7] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[6][7] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[7][7] ),
    .S1(_08587_),
    .X(_08816_));
 sg13g2_mux4_1 _15566_ (.S0(net814),
    .A0(_08813_),
    .A1(_08814_),
    .A2(_08815_),
    .A3(_08816_),
    .S1(net940),
    .X(_08817_));
 sg13g2_mux2_1 _15567_ (.A0(_08812_),
    .A1(_08817_),
    .S(net823),
    .X(_08818_));
 sg13g2_nand2b_1 _15568_ (.Y(_08819_),
    .B(_08818_),
    .A_N(net1080));
 sg13g2_buf_2 _15569_ (.A(_08819_),
    .X(_08820_));
 sg13g2_a22oi_1 _15570_ (.Y(_08821_),
    .B1(net719),
    .B2(\cpu.icache.r_tag[4][19] ),
    .A2(_08642_),
    .A1(\cpu.icache.r_tag[2][19] ));
 sg13g2_a22oi_1 _15571_ (.Y(_08822_),
    .B1(net642),
    .B2(\cpu.icache.r_tag[1][19] ),
    .A2(net724),
    .A1(\cpu.icache.r_tag[5][19] ));
 sg13g2_mux2_1 _15572_ (.A0(\cpu.icache.r_tag[7][19] ),
    .A1(\cpu.icache.r_tag[3][19] ),
    .S(net938),
    .X(_08823_));
 sg13g2_buf_2 _15573_ (.A(net932),
    .X(_08824_));
 sg13g2_a22oi_1 _15574_ (.Y(_08825_),
    .B1(_08823_),
    .B2(net808),
    .A2(_08566_),
    .A1(\cpu.icache.r_tag[6][19] ));
 sg13g2_buf_2 _15575_ (.A(_08610_),
    .X(_08826_));
 sg13g2_nand2b_1 _15576_ (.Y(_08827_),
    .B(net710),
    .A_N(_08825_));
 sg13g2_nand3_1 _15577_ (.B(_08822_),
    .C(_08827_),
    .A(_08821_),
    .Y(_08828_));
 sg13g2_mux2_1 _15578_ (.A0(\cpu.icache.r_tag[0][19] ),
    .A1(_08828_),
    .S(net520),
    .X(_08829_));
 sg13g2_xor2_1 _15579_ (.B(_08829_),
    .A(net427),
    .X(_08830_));
 sg13g2_nand3_1 _15580_ (.B(_08807_),
    .C(_08830_),
    .A(_08786_),
    .Y(_08831_));
 sg13g2_mux4_1 _15581_ (.S0(net811),
    .A0(\cpu.genblk1.mmu.r_vtop_i[16][2] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[17][2] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[18][2] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[19][2] ),
    .S1(net714),
    .X(_08832_));
 sg13g2_mux4_1 _15582_ (.S0(net811),
    .A0(\cpu.genblk1.mmu.r_vtop_i[0][2] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[1][2] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[2][2] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[3][2] ),
    .S1(net714),
    .X(_08833_));
 sg13g2_buf_2 _15583_ (.A(net934),
    .X(_08834_));
 sg13g2_buf_2 _15584_ (.A(net815),
    .X(_08835_));
 sg13g2_mux4_1 _15585_ (.S0(net807),
    .A0(\cpu.genblk1.mmu.r_vtop_i[24][2] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[25][2] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[26][2] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[27][2] ),
    .S1(net709),
    .X(_08836_));
 sg13g2_mux4_1 _15586_ (.S0(net807),
    .A0(\cpu.genblk1.mmu.r_vtop_i[8][2] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[9][2] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[10][2] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[11][2] ),
    .S1(net714),
    .X(_08837_));
 sg13g2_mux4_1 _15587_ (.S0(net946),
    .A0(_08832_),
    .A1(_08833_),
    .A2(_08836_),
    .A3(_08837_),
    .S1(_08397_),
    .X(_08838_));
 sg13g2_a21oi_1 _15588_ (.A1(net1083),
    .A2(_08838_),
    .Y(_08839_),
    .B1(net931));
 sg13g2_inv_1 _15589_ (.Y(_08840_),
    .A(net931));
 sg13g2_mux4_1 _15590_ (.S0(net811),
    .A0(\cpu.genblk1.mmu.r_vtop_i[20][2] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[21][2] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[22][2] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[23][2] ),
    .S1(net714),
    .X(_08841_));
 sg13g2_mux4_1 _15591_ (.S0(net811),
    .A0(\cpu.genblk1.mmu.r_vtop_i[4][2] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[5][2] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[6][2] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[7][2] ),
    .S1(net714),
    .X(_08842_));
 sg13g2_mux4_1 _15592_ (.S0(net811),
    .A0(\cpu.genblk1.mmu.r_vtop_i[28][2] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[29][2] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[30][2] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[31][2] ),
    .S1(net714),
    .X(_08843_));
 sg13g2_mux4_1 _15593_ (.S0(net811),
    .A0(\cpu.genblk1.mmu.r_vtop_i[12][2] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[13][2] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[14][2] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[15][2] ),
    .S1(net714),
    .X(_08844_));
 sg13g2_mux4_1 _15594_ (.S0(net946),
    .A0(_08841_),
    .A1(_08842_),
    .A2(_08843_),
    .A3(_08844_),
    .S1(_08397_),
    .X(_08845_));
 sg13g2_nor3_1 _15595_ (.A(_08840_),
    .B(_08339_),
    .C(_08845_),
    .Y(_08846_));
 sg13g2_or2_1 _15596_ (.X(_08847_),
    .B(_08846_),
    .A(_08839_));
 sg13g2_buf_2 _15597_ (.A(_08847_),
    .X(_08848_));
 sg13g2_a22oi_1 _15598_ (.Y(_08849_),
    .B1(net719),
    .B2(\cpu.icache.r_tag[4][14] ),
    .A2(net642),
    .A1(\cpu.icache.r_tag[1][14] ));
 sg13g2_a22oi_1 _15599_ (.Y(_08850_),
    .B1(_08518_),
    .B2(\cpu.icache.r_tag[5][14] ),
    .A2(net643),
    .A1(\cpu.icache.r_tag[2][14] ));
 sg13g2_mux2_1 _15600_ (.A0(\cpu.icache.r_tag[7][14] ),
    .A1(\cpu.icache.r_tag[3][14] ),
    .S(net817),
    .X(_08851_));
 sg13g2_a22oi_1 _15601_ (.Y(_08852_),
    .B1(_08851_),
    .B2(net808),
    .A2(_08566_),
    .A1(\cpu.icache.r_tag[6][14] ));
 sg13g2_nand2b_1 _15602_ (.Y(_08853_),
    .B(net710),
    .A_N(_08852_));
 sg13g2_nand4_1 _15603_ (.B(_08849_),
    .C(_08850_),
    .A(net520),
    .Y(_08854_),
    .D(_08853_));
 sg13g2_o21ai_1 _15604_ (.B1(_08854_),
    .Y(_08855_),
    .A1(\cpu.icache.r_tag[0][14] ),
    .A2(net521));
 sg13g2_xnor2_1 _15605_ (.Y(_08856_),
    .A(net426),
    .B(_08855_));
 sg13g2_mux4_1 _15606_ (.S0(_08834_),
    .A0(\cpu.genblk1.mmu.r_vtop_i[24][8] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[25][8] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[26][8] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[27][8] ),
    .S1(net709),
    .X(_08857_));
 sg13g2_mux4_1 _15607_ (.S0(_08834_),
    .A0(\cpu.genblk1.mmu.r_vtop_i[16][8] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[17][8] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[18][8] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[19][8] ),
    .S1(_08835_),
    .X(_08858_));
 sg13g2_mux4_1 _15608_ (.S0(_08655_),
    .A0(\cpu.genblk1.mmu.r_vtop_i[28][8] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[29][8] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[30][8] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[31][8] ),
    .S1(_08656_),
    .X(_08859_));
 sg13g2_mux4_1 _15609_ (.S0(_08655_),
    .A0(\cpu.genblk1.mmu.r_vtop_i[20][8] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[21][8] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[22][8] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[23][8] ),
    .S1(_08835_),
    .X(_08860_));
 sg13g2_mux4_1 _15610_ (.S0(net814),
    .A0(_08857_),
    .A1(_08858_),
    .A2(_08859_),
    .A3(_08860_),
    .S1(_08625_),
    .X(_08861_));
 sg13g2_mux4_1 _15611_ (.S0(net807),
    .A0(\cpu.genblk1.mmu.r_vtop_i[8][8] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[9][8] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[10][8] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[11][8] ),
    .S1(net709),
    .X(_08862_));
 sg13g2_mux4_1 _15612_ (.S0(net807),
    .A0(\cpu.genblk1.mmu.r_vtop_i[0][8] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[1][8] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[2][8] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[3][8] ),
    .S1(net709),
    .X(_08863_));
 sg13g2_mux4_1 _15613_ (.S0(net810),
    .A0(\cpu.genblk1.mmu.r_vtop_i[12][8] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[13][8] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[14][8] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[15][8] ),
    .S1(_08656_),
    .X(_08864_));
 sg13g2_mux4_1 _15614_ (.S0(net810),
    .A0(\cpu.genblk1.mmu.r_vtop_i[4][8] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[5][8] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[6][8] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[7][8] ),
    .S1(net711),
    .X(_08865_));
 sg13g2_mux4_1 _15615_ (.S0(net814),
    .A0(_08862_),
    .A1(_08863_),
    .A2(_08864_),
    .A3(_08865_),
    .S1(_08625_),
    .X(_08866_));
 sg13g2_mux2_1 _15616_ (.A0(_08861_),
    .A1(_08866_),
    .S(net823),
    .X(_08867_));
 sg13g2_nand2b_1 _15617_ (.Y(_08868_),
    .B(_08867_),
    .A_N(net1080));
 sg13g2_buf_1 _15618_ (.A(_08868_),
    .X(_08869_));
 sg13g2_a22oi_1 _15619_ (.Y(_08870_),
    .B1(_08569_),
    .B2(\cpu.icache.r_tag[6][20] ),
    .A2(_08523_),
    .A1(\cpu.icache.r_tag[1][20] ));
 sg13g2_a22oi_1 _15620_ (.Y(_08871_),
    .B1(_08574_),
    .B2(\cpu.icache.r_tag[4][20] ),
    .A2(_08514_),
    .A1(\cpu.icache.r_tag[2][20] ));
 sg13g2_mux2_1 _15621_ (.A0(\cpu.icache.r_tag[7][20] ),
    .A1(\cpu.icache.r_tag[3][20] ),
    .S(_08575_),
    .X(_08872_));
 sg13g2_a22oi_1 _15622_ (.Y(_08873_),
    .B1(_08872_),
    .B2(_08611_),
    .A2(_08692_),
    .A1(\cpu.icache.r_tag[5][20] ));
 sg13g2_nand2b_1 _15623_ (.Y(_08874_),
    .B(net808),
    .A_N(_08873_));
 sg13g2_nand4_1 _15624_ (.B(_08870_),
    .C(_08871_),
    .A(_08606_),
    .Y(_08875_),
    .D(_08874_));
 sg13g2_o21ai_1 _15625_ (.B1(_08875_),
    .Y(_08876_),
    .A1(\cpu.icache.r_tag[0][20] ),
    .A2(_08509_));
 sg13g2_xnor2_1 _15626_ (.Y(_08877_),
    .A(net425),
    .B(_08876_));
 sg13g2_mux4_1 _15627_ (.S0(net807),
    .A0(\cpu.genblk1.mmu.r_vtop_i[24][10] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[25][10] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[26][10] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[27][10] ),
    .S1(net709),
    .X(_08878_));
 sg13g2_mux4_1 _15628_ (.S0(net807),
    .A0(\cpu.genblk1.mmu.r_vtop_i[16][10] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[17][10] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[18][10] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[19][10] ),
    .S1(net709),
    .X(_08879_));
 sg13g2_mux4_1 _15629_ (.S0(net810),
    .A0(\cpu.genblk1.mmu.r_vtop_i[28][10] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[29][10] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[30][10] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[31][10] ),
    .S1(net711),
    .X(_08880_));
 sg13g2_mux4_1 _15630_ (.S0(net810),
    .A0(\cpu.genblk1.mmu.r_vtop_i[20][10] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[21][10] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[22][10] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[23][10] ),
    .S1(net711),
    .X(_08881_));
 sg13g2_mux4_1 _15631_ (.S0(net814),
    .A0(_08878_),
    .A1(_08879_),
    .A2(_08880_),
    .A3(_08881_),
    .S1(net931),
    .X(_08882_));
 sg13g2_mux4_1 _15632_ (.S0(net807),
    .A0(\cpu.genblk1.mmu.r_vtop_i[8][10] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[9][10] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[10][10] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[11][10] ),
    .S1(net709),
    .X(_08883_));
 sg13g2_mux4_1 _15633_ (.S0(net807),
    .A0(\cpu.genblk1.mmu.r_vtop_i[0][10] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[1][10] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[2][10] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[3][10] ),
    .S1(net709),
    .X(_08884_));
 sg13g2_mux4_1 _15634_ (.S0(net810),
    .A0(\cpu.genblk1.mmu.r_vtop_i[12][10] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[13][10] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[14][10] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[15][10] ),
    .S1(net711),
    .X(_08885_));
 sg13g2_mux4_1 _15635_ (.S0(net810),
    .A0(\cpu.genblk1.mmu.r_vtop_i[4][10] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[5][10] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[6][10] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[7][10] ),
    .S1(net711),
    .X(_08886_));
 sg13g2_mux4_1 _15636_ (.S0(net814),
    .A0(_08883_),
    .A1(_08884_),
    .A2(_08885_),
    .A3(_08886_),
    .S1(net931),
    .X(_08887_));
 sg13g2_mux2_1 _15637_ (.A0(_08882_),
    .A1(_08887_),
    .S(net823),
    .X(_08888_));
 sg13g2_nand2b_2 _15638_ (.Y(_08889_),
    .B(_08888_),
    .A_N(net1080));
 sg13g2_buf_1 _15639_ (.A(_08889_),
    .X(_08890_));
 sg13g2_a22oi_1 _15640_ (.Y(_08891_),
    .B1(_08569_),
    .B2(\cpu.icache.r_tag[6][22] ),
    .A2(_08523_),
    .A1(\cpu.icache.r_tag[1][22] ));
 sg13g2_a22oi_1 _15641_ (.Y(_08892_),
    .B1(_08574_),
    .B2(\cpu.icache.r_tag[4][22] ),
    .A2(_08514_),
    .A1(\cpu.icache.r_tag[2][22] ));
 sg13g2_mux2_1 _15642_ (.A0(\cpu.icache.r_tag[7][22] ),
    .A1(\cpu.icache.r_tag[3][22] ),
    .S(_08575_),
    .X(_08893_));
 sg13g2_a22oi_1 _15643_ (.Y(_08894_),
    .B1(_08893_),
    .B2(_08611_),
    .A2(_08692_),
    .A1(\cpu.icache.r_tag[5][22] ));
 sg13g2_nand2b_1 _15644_ (.Y(_08895_),
    .B(net808),
    .A_N(_08894_));
 sg13g2_nand4_1 _15645_ (.B(_08891_),
    .C(_08892_),
    .A(_08606_),
    .Y(_08896_),
    .D(_08895_));
 sg13g2_o21ai_1 _15646_ (.B1(_08896_),
    .Y(_08897_),
    .A1(\cpu.icache.r_tag[0][22] ),
    .A2(_08509_));
 sg13g2_xnor2_1 _15647_ (.Y(_08898_),
    .A(net424),
    .B(_08897_));
 sg13g2_nand3_1 _15648_ (.B(_08877_),
    .C(_08898_),
    .A(_08856_),
    .Y(_08899_));
 sg13g2_nor4_2 _15649_ (.A(_08581_),
    .B(_08743_),
    .C(_08831_),
    .Y(_08900_),
    .D(_08899_));
 sg13g2_nand2_1 _15650_ (.Y(_08901_),
    .A(_08471_),
    .B(_08900_));
 sg13g2_buf_2 _15651_ (.A(_08901_),
    .X(_08902_));
 sg13g2_buf_1 _15652_ (.A(_08902_),
    .X(_08903_));
 sg13g2_buf_1 _15653_ (.A(net173),
    .X(_08904_));
 sg13g2_buf_1 _15654_ (.A(_08902_),
    .X(_08905_));
 sg13g2_buf_1 _15655_ (.A(\cpu.ex.pc[1] ),
    .X(_08906_));
 sg13g2_mux4_1 _15656_ (.S0(net1079),
    .A0(\cpu.icache.r_data[4][22] ),
    .A1(\cpu.icache.r_data[5][22] ),
    .A2(\cpu.icache.r_data[6][22] ),
    .A3(\cpu.icache.r_data[7][22] ),
    .S1(net813),
    .X(_08907_));
 sg13g2_and2_1 _15657_ (.A(\cpu.icache.r_data[3][22] ),
    .B(_08528_),
    .X(_08908_));
 sg13g2_a221oi_1 _15658_ (.B2(\cpu.icache.r_data[1][22] ),
    .C1(_08908_),
    .B1(_08521_),
    .A1(\cpu.icache.r_data[2][22] ),
    .Y(_08909_),
    .A2(_08512_));
 sg13g2_o21ai_1 _15659_ (.B1(_08909_),
    .Y(_08910_),
    .A1(_00202_),
    .A2(net640));
 sg13g2_a21oi_1 _15660_ (.A1(net812),
    .A2(_08907_),
    .Y(_08911_),
    .B1(_08910_));
 sg13g2_and2_1 _15661_ (.A(net1082),
    .B(_08504_),
    .X(_08912_));
 sg13g2_buf_1 _15662_ (.A(_08912_),
    .X(_08913_));
 sg13g2_nand2_1 _15663_ (.Y(_08914_),
    .A(_00201_),
    .B(_08913_));
 sg13g2_a22oi_1 _15664_ (.Y(_08915_),
    .B1(_08521_),
    .B2(\cpu.icache.r_data[1][6] ),
    .A2(_08512_),
    .A1(\cpu.icache.r_data[2][6] ));
 sg13g2_mux4_1 _15665_ (.S0(_08499_),
    .A0(\cpu.icache.r_data[4][6] ),
    .A1(\cpu.icache.r_data[5][6] ),
    .A2(\cpu.icache.r_data[6][6] ),
    .A3(\cpu.icache.r_data[7][6] ),
    .S1(net936),
    .X(_08916_));
 sg13g2_a22oi_1 _15666_ (.Y(_08917_),
    .B1(_08916_),
    .B2(net939),
    .A2(_08528_),
    .A1(\cpu.icache.r_data[3][6] ));
 sg13g2_nand3_1 _15667_ (.B(_08915_),
    .C(_08917_),
    .A(net640),
    .Y(_08918_));
 sg13g2_a21oi_1 _15668_ (.A1(_08914_),
    .A2(_08918_),
    .Y(_08919_),
    .B1(_08906_));
 sg13g2_a21oi_1 _15669_ (.A1(_08906_),
    .A2(_08911_),
    .Y(_08920_),
    .B1(_08919_));
 sg13g2_buf_2 _15670_ (.A(_08920_),
    .X(_08921_));
 sg13g2_inv_2 _15671_ (.Y(_08922_),
    .A(_08921_));
 sg13g2_nor2_1 _15672_ (.A(_00200_),
    .B(_08506_),
    .Y(_08923_));
 sg13g2_nor2_1 _15673_ (.A(_08515_),
    .B(net1081),
    .Y(_08924_));
 sg13g2_mux2_1 _15674_ (.A0(\cpu.icache.r_data[4][21] ),
    .A1(\cpu.icache.r_data[6][21] ),
    .S(net936),
    .X(_08925_));
 sg13g2_a22oi_1 _15675_ (.Y(_08926_),
    .B1(_08925_),
    .B2(_08515_),
    .A2(_08924_),
    .A1(\cpu.icache.r_data[5][21] ));
 sg13g2_nor2_1 _15676_ (.A(net817),
    .B(_08926_),
    .Y(_08927_));
 sg13g2_and2_1 _15677_ (.A(_08533_),
    .B(\cpu.icache.r_data[3][21] ),
    .X(_08928_));
 sg13g2_a21oi_1 _15678_ (.A1(net939),
    .A2(\cpu.icache.r_data[7][21] ),
    .Y(_08929_),
    .B1(_08928_));
 sg13g2_a22oi_1 _15679_ (.Y(_08930_),
    .B1(_08521_),
    .B2(\cpu.icache.r_data[1][21] ),
    .A2(_08512_),
    .A1(\cpu.icache.r_data[2][21] ));
 sg13g2_o21ai_1 _15680_ (.B1(_08930_),
    .Y(_08931_),
    .A1(_08527_),
    .A2(_08929_));
 sg13g2_nor3_1 _15681_ (.A(_08923_),
    .B(_08927_),
    .C(_08931_),
    .Y(_08932_));
 sg13g2_nand2_1 _15682_ (.Y(_08933_),
    .A(_00199_),
    .B(_08913_));
 sg13g2_a22oi_1 _15683_ (.Y(_08934_),
    .B1(_08521_),
    .B2(\cpu.icache.r_data[1][5] ),
    .A2(_08512_),
    .A1(\cpu.icache.r_data[2][5] ));
 sg13g2_a22oi_1 _15684_ (.Y(_08935_),
    .B1(_08528_),
    .B2(\cpu.icache.r_data[3][5] ),
    .A2(net822),
    .A1(\cpu.icache.r_data[5][5] ));
 sg13g2_mux2_1 _15685_ (.A0(\cpu.icache.r_data[4][5] ),
    .A1(\cpu.icache.r_data[6][5] ),
    .S(net1081),
    .X(_08936_));
 sg13g2_a22oi_1 _15686_ (.Y(_08937_),
    .B1(_08936_),
    .B2(_08515_),
    .A2(net937),
    .A1(\cpu.icache.r_data[7][5] ));
 sg13g2_or2_1 _15687_ (.X(_08938_),
    .B(_08937_),
    .A(net938));
 sg13g2_nand4_1 _15688_ (.B(_08934_),
    .C(_08935_),
    .A(net640),
    .Y(_08939_),
    .D(_08938_));
 sg13g2_a21oi_1 _15689_ (.A1(_08933_),
    .A2(_08939_),
    .Y(_08940_),
    .B1(_08906_));
 sg13g2_a21oi_1 _15690_ (.A1(_08906_),
    .A2(_08932_),
    .Y(_08941_),
    .B1(_08940_));
 sg13g2_buf_2 _15691_ (.A(_08941_),
    .X(_08942_));
 sg13g2_inv_2 _15692_ (.Y(_08943_),
    .A(_08942_));
 sg13g2_nand2_1 _15693_ (.Y(_08944_),
    .A(_08922_),
    .B(_08943_));
 sg13g2_buf_1 _15694_ (.A(_08944_),
    .X(_08945_));
 sg13g2_inv_1 _15695_ (.Y(_08946_),
    .A(_08906_));
 sg13g2_nor2_1 _15696_ (.A(_00198_),
    .B(net584),
    .Y(_08947_));
 sg13g2_buf_1 _15697_ (.A(_08924_),
    .X(_08948_));
 sg13g2_mux2_1 _15698_ (.A0(\cpu.icache.r_data[4][31] ),
    .A1(\cpu.icache.r_data[6][31] ),
    .S(net813),
    .X(_08949_));
 sg13g2_buf_2 _15699_ (.A(net935),
    .X(_08950_));
 sg13g2_a22oi_1 _15700_ (.Y(_08951_),
    .B1(_08949_),
    .B2(net805),
    .A2(net806),
    .A1(\cpu.icache.r_data[5][31] ));
 sg13g2_nor2_1 _15701_ (.A(net721),
    .B(_08951_),
    .Y(_08952_));
 sg13g2_and2_1 _15702_ (.A(net817),
    .B(\cpu.icache.r_data[3][31] ),
    .X(_08953_));
 sg13g2_a21oi_1 _15703_ (.A1(net812),
    .A2(\cpu.icache.r_data[7][31] ),
    .Y(_08954_),
    .B1(_08953_));
 sg13g2_a22oi_1 _15704_ (.Y(_08955_),
    .B1(net639),
    .B2(\cpu.icache.r_data[1][31] ),
    .A2(net638),
    .A1(\cpu.icache.r_data[2][31] ));
 sg13g2_o21ai_1 _15705_ (.B1(_08955_),
    .Y(_08956_),
    .A1(_08527_),
    .A2(_08954_));
 sg13g2_nor4_1 _15706_ (.A(net1076),
    .B(_08947_),
    .C(_08952_),
    .D(_08956_),
    .Y(_08957_));
 sg13g2_buf_1 _15707_ (.A(_08913_),
    .X(_08958_));
 sg13g2_buf_1 _15708_ (.A(_08958_),
    .X(_08959_));
 sg13g2_nand2_1 _15709_ (.Y(_08960_),
    .A(_00197_),
    .B(net580));
 sg13g2_a22oi_1 _15710_ (.Y(_08961_),
    .B1(net639),
    .B2(\cpu.icache.r_data[1][15] ),
    .A2(net638),
    .A1(\cpu.icache.r_data[2][15] ));
 sg13g2_a22oi_1 _15711_ (.Y(_08962_),
    .B1(net720),
    .B2(\cpu.icache.r_data[6][15] ),
    .A2(net583),
    .A1(\cpu.icache.r_data[3][15] ));
 sg13g2_mux2_1 _15712_ (.A0(\cpu.icache.r_data[5][15] ),
    .A1(\cpu.icache.r_data[7][15] ),
    .S(net819),
    .X(_08963_));
 sg13g2_a22oi_1 _15713_ (.Y(_08964_),
    .B1(_08963_),
    .B2(net932),
    .A2(_08734_),
    .A1(\cpu.icache.r_data[4][15] ));
 sg13g2_or2_1 _15714_ (.X(_08965_),
    .B(_08964_),
    .A(net821));
 sg13g2_nand4_1 _15715_ (.B(_08961_),
    .C(_08962_),
    .A(net584),
    .Y(_08966_),
    .D(_08965_));
 sg13g2_buf_1 _15716_ (.A(_08906_),
    .X(_08967_));
 sg13g2_buf_1 _15717_ (.A(net1075),
    .X(_08968_));
 sg13g2_a21oi_1 _15718_ (.A1(_08960_),
    .A2(_08966_),
    .Y(_08969_),
    .B1(net929));
 sg13g2_or2_1 _15719_ (.X(_08970_),
    .B(_08969_),
    .A(_08957_));
 sg13g2_buf_2 _15720_ (.A(_08970_),
    .X(_08971_));
 sg13g2_nand2_1 _15721_ (.Y(_08972_),
    .A(\cpu.icache.r_data[0][13] ),
    .B(net637));
 sg13g2_mux4_1 _15722_ (.S0(net932),
    .A0(\cpu.icache.r_data[4][13] ),
    .A1(\cpu.icache.r_data[5][13] ),
    .A2(\cpu.icache.r_data[6][13] ),
    .A3(\cpu.icache.r_data[7][13] ),
    .S1(net716),
    .X(_08973_));
 sg13g2_nand2_1 _15723_ (.Y(_08974_),
    .A(net715),
    .B(_08973_));
 sg13g2_nand2_1 _15724_ (.Y(_08975_),
    .A(\cpu.icache.r_data[3][13] ),
    .B(net583));
 sg13g2_a22oi_1 _15725_ (.Y(_08976_),
    .B1(net642),
    .B2(\cpu.icache.r_data[1][13] ),
    .A2(net638),
    .A1(\cpu.icache.r_data[2][13] ));
 sg13g2_nand4_1 _15726_ (.B(_08974_),
    .C(_08975_),
    .A(_08972_),
    .Y(_08977_),
    .D(_08976_));
 sg13g2_mux2_1 _15727_ (.A0(\cpu.icache.r_data[4][29] ),
    .A1(\cpu.icache.r_data[6][29] ),
    .S(net936),
    .X(_08978_));
 sg13g2_a22oi_1 _15728_ (.Y(_08979_),
    .B1(_08978_),
    .B2(net935),
    .A2(net937),
    .A1(\cpu.icache.r_data[7][29] ));
 sg13g2_or2_1 _15729_ (.X(_08980_),
    .B(_08979_),
    .A(net821));
 sg13g2_a22oi_1 _15730_ (.Y(_08981_),
    .B1(net723),
    .B2(\cpu.icache.r_data[1][29] ),
    .A2(net725),
    .A1(\cpu.icache.r_data[2][29] ));
 sg13g2_a22oi_1 _15731_ (.Y(_08982_),
    .B1(net641),
    .B2(\cpu.icache.r_data[3][29] ),
    .A2(net822),
    .A1(\cpu.icache.r_data[5][29] ));
 sg13g2_nand3_1 _15732_ (.B(_08981_),
    .C(_08982_),
    .A(_08980_),
    .Y(_08983_));
 sg13g2_a21oi_1 _15733_ (.A1(\cpu.icache.r_data[0][29] ),
    .A2(net637),
    .Y(_08984_),
    .B1(_08983_));
 sg13g2_nand2_1 _15734_ (.Y(_08985_),
    .A(net1075),
    .B(_08984_));
 sg13g2_o21ai_1 _15735_ (.B1(_08985_),
    .Y(_08986_),
    .A1(net929),
    .A2(_08977_));
 sg13g2_buf_1 _15736_ (.A(_08986_),
    .X(_08987_));
 sg13g2_inv_1 _15737_ (.Y(_08988_),
    .A(_00196_));
 sg13g2_a22oi_1 _15738_ (.Y(_08989_),
    .B1(_08573_),
    .B2(\cpu.icache.r_data[4][30] ),
    .A2(net723),
    .A1(\cpu.icache.r_data[1][30] ));
 sg13g2_mux2_1 _15739_ (.A0(\cpu.icache.r_data[7][30] ),
    .A1(\cpu.icache.r_data[3][30] ),
    .S(net938),
    .X(_08990_));
 sg13g2_a22oi_1 _15740_ (.Y(_08991_),
    .B1(net937),
    .B2(_08990_),
    .A2(net822),
    .A1(\cpu.icache.r_data[5][30] ));
 sg13g2_a22oi_1 _15741_ (.Y(_08992_),
    .B1(net720),
    .B2(\cpu.icache.r_data[6][30] ),
    .A2(net712),
    .A1(\cpu.icache.r_data[2][30] ));
 sg13g2_nand3_1 _15742_ (.B(_08991_),
    .C(_08992_),
    .A(_08989_),
    .Y(_08993_));
 sg13g2_a21oi_1 _15743_ (.A1(_08988_),
    .A2(net637),
    .Y(_08994_),
    .B1(_08993_));
 sg13g2_nand2_1 _15744_ (.Y(_08995_),
    .A(_00195_),
    .B(net637));
 sg13g2_mux4_1 _15745_ (.S0(net1079),
    .A0(\cpu.icache.r_data[4][14] ),
    .A1(\cpu.icache.r_data[5][14] ),
    .A2(\cpu.icache.r_data[6][14] ),
    .A3(\cpu.icache.r_data[7][14] ),
    .S1(net819),
    .X(_08996_));
 sg13g2_nand2_1 _15746_ (.Y(_08997_),
    .A(net812),
    .B(_08996_));
 sg13g2_nand2_1 _15747_ (.Y(_08998_),
    .A(\cpu.icache.r_data[1][14] ),
    .B(net723));
 sg13g2_a22oi_1 _15748_ (.Y(_08999_),
    .B1(net722),
    .B2(\cpu.icache.r_data[3][14] ),
    .A2(net712),
    .A1(\cpu.icache.r_data[2][14] ));
 sg13g2_nand4_1 _15749_ (.B(_08997_),
    .C(_08998_),
    .A(net644),
    .Y(_09000_),
    .D(_08999_));
 sg13g2_nand3_1 _15750_ (.B(_08995_),
    .C(_09000_),
    .A(net1076),
    .Y(_09001_));
 sg13g2_o21ai_1 _15751_ (.B1(_09001_),
    .Y(_09002_),
    .A1(net1076),
    .A2(_08994_));
 sg13g2_buf_1 _15752_ (.A(_09002_),
    .X(_09003_));
 sg13g2_inv_1 _15753_ (.Y(_09004_),
    .A(_09003_));
 sg13g2_nand2_1 _15754_ (.Y(_09005_),
    .A(net293),
    .B(_09004_));
 sg13g2_buf_2 _15755_ (.A(_09005_),
    .X(_09006_));
 sg13g2_nor2_1 _15756_ (.A(_08971_),
    .B(_09006_),
    .Y(_09007_));
 sg13g2_buf_1 _15757_ (.A(_09007_),
    .X(_09008_));
 sg13g2_buf_1 _15758_ (.A(net929),
    .X(_09009_));
 sg13g2_buf_1 _15759_ (.A(net639),
    .X(_09010_));
 sg13g2_nand2_1 _15760_ (.Y(_09011_),
    .A(\cpu.icache.r_data[1][0] ),
    .B(net579));
 sg13g2_a22oi_1 _15761_ (.Y(_09012_),
    .B1(_08639_),
    .B2(\cpu.icache.r_data[7][0] ),
    .A2(net720),
    .A1(\cpu.icache.r_data[6][0] ));
 sg13g2_a22oi_1 _15762_ (.Y(_09013_),
    .B1(net719),
    .B2(\cpu.icache.r_data[4][0] ),
    .A2(net581),
    .A1(\cpu.icache.r_data[2][0] ));
 sg13g2_a22oi_1 _15763_ (.Y(_09014_),
    .B1(net583),
    .B2(\cpu.icache.r_data[3][0] ),
    .A2(net724),
    .A1(\cpu.icache.r_data[5][0] ));
 sg13g2_nand4_1 _15764_ (.B(_09012_),
    .C(_09013_),
    .A(_09011_),
    .Y(_09015_),
    .D(_09014_));
 sg13g2_mux2_1 _15765_ (.A0(\cpu.icache.r_data[0][0] ),
    .A1(_09015_),
    .S(net521),
    .X(_09016_));
 sg13g2_mux2_1 _15766_ (.A0(\cpu.icache.r_data[4][16] ),
    .A1(\cpu.icache.r_data[6][16] ),
    .S(net716),
    .X(_09017_));
 sg13g2_a22oi_1 _15767_ (.Y(_09018_),
    .B1(_09017_),
    .B2(net805),
    .A2(net820),
    .A1(\cpu.icache.r_data[7][16] ));
 sg13g2_or2_1 _15768_ (.X(_09019_),
    .B(_09018_),
    .A(net721));
 sg13g2_a22oi_1 _15769_ (.Y(_09020_),
    .B1(net579),
    .B2(\cpu.icache.r_data[1][16] ),
    .A2(net724),
    .A1(\cpu.icache.r_data[5][16] ));
 sg13g2_a22oi_1 _15770_ (.Y(_09021_),
    .B1(net583),
    .B2(\cpu.icache.r_data[3][16] ),
    .A2(net581),
    .A1(\cpu.icache.r_data[2][16] ));
 sg13g2_nand3_1 _15771_ (.B(_09020_),
    .C(_09021_),
    .A(_09019_),
    .Y(_09022_));
 sg13g2_a21oi_1 _15772_ (.A1(\cpu.icache.r_data[0][16] ),
    .A2(net580),
    .Y(_09023_),
    .B1(_09022_));
 sg13g2_nand2_1 _15773_ (.Y(_09024_),
    .A(net929),
    .B(_09023_));
 sg13g2_o21ai_1 _15774_ (.B1(_09024_),
    .Y(_09025_),
    .A1(net804),
    .A2(_09016_));
 sg13g2_buf_1 _15775_ (.A(_09025_),
    .X(_09026_));
 sg13g2_buf_1 _15776_ (.A(_09026_),
    .X(_09027_));
 sg13g2_mux4_1 _15777_ (.S0(net808),
    .A0(\cpu.icache.r_data[4][1] ),
    .A1(\cpu.icache.r_data[5][1] ),
    .A2(\cpu.icache.r_data[6][1] ),
    .A3(\cpu.icache.r_data[7][1] ),
    .S1(net710),
    .X(_09028_));
 sg13g2_nand2_1 _15778_ (.Y(_09029_),
    .A(net715),
    .B(_09028_));
 sg13g2_nand2_1 _15779_ (.Y(_09030_),
    .A(\cpu.icache.r_data[1][1] ),
    .B(net579));
 sg13g2_buf_2 _15780_ (.A(net583),
    .X(_09031_));
 sg13g2_a22oi_1 _15781_ (.Y(_09032_),
    .B1(net518),
    .B2(\cpu.icache.r_data[3][1] ),
    .A2(net581),
    .A1(\cpu.icache.r_data[2][1] ));
 sg13g2_nand4_1 _15782_ (.B(_09029_),
    .C(_09030_),
    .A(net521),
    .Y(_09033_),
    .D(_09032_));
 sg13g2_o21ai_1 _15783_ (.B1(_09033_),
    .Y(_09034_),
    .A1(\cpu.icache.r_data[0][1] ),
    .A2(net521));
 sg13g2_buf_1 _15784_ (.A(net719),
    .X(_09035_));
 sg13g2_a22oi_1 _15785_ (.Y(_09036_),
    .B1(net636),
    .B2(\cpu.icache.r_data[4][17] ),
    .A2(net579),
    .A1(\cpu.icache.r_data[1][17] ));
 sg13g2_buf_1 _15786_ (.A(net720),
    .X(_09037_));
 sg13g2_mux2_1 _15787_ (.A0(\cpu.icache.r_data[7][17] ),
    .A1(\cpu.icache.r_data[3][17] ),
    .S(net721),
    .X(_09038_));
 sg13g2_a22oi_1 _15788_ (.Y(_09039_),
    .B1(_09038_),
    .B2(net820),
    .A2(net635),
    .A1(\cpu.icache.r_data[6][17] ));
 sg13g2_a22oi_1 _15789_ (.Y(_09040_),
    .B1(net724),
    .B2(\cpu.icache.r_data[5][17] ),
    .A2(net581),
    .A1(\cpu.icache.r_data[2][17] ));
 sg13g2_nand2_1 _15790_ (.Y(_09041_),
    .A(\cpu.icache.r_data[0][17] ),
    .B(net580));
 sg13g2_nand4_1 _15791_ (.B(_09039_),
    .C(_09040_),
    .A(_09036_),
    .Y(_09042_),
    .D(_09041_));
 sg13g2_nand2_1 _15792_ (.Y(_09043_),
    .A(net804),
    .B(_09042_));
 sg13g2_o21ai_1 _15793_ (.B1(_09043_),
    .Y(_09044_),
    .A1(net804),
    .A2(_09034_));
 sg13g2_buf_2 _15794_ (.A(_09044_),
    .X(_09045_));
 sg13g2_nor2_1 _15795_ (.A(net225),
    .B(_09045_),
    .Y(_09046_));
 sg13g2_buf_1 _15796_ (.A(_09046_),
    .X(_09047_));
 sg13g2_nor2_1 _15797_ (.A(_00194_),
    .B(net640),
    .Y(_09048_));
 sg13g2_mux2_1 _15798_ (.A0(\cpu.icache.r_data[4][27] ),
    .A1(\cpu.icache.r_data[6][27] ),
    .S(_08541_),
    .X(_09049_));
 sg13g2_a22oi_1 _15799_ (.Y(_09050_),
    .B1(_09049_),
    .B2(net935),
    .A2(_08924_),
    .A1(\cpu.icache.r_data[5][27] ));
 sg13g2_nor2_1 _15800_ (.A(net821),
    .B(_09050_),
    .Y(_09051_));
 sg13g2_and2_1 _15801_ (.A(net1082),
    .B(\cpu.icache.r_data[3][27] ),
    .X(_09052_));
 sg13g2_a21oi_1 _15802_ (.A1(_08525_),
    .A2(\cpu.icache.r_data[7][27] ),
    .Y(_09053_),
    .B1(_09052_));
 sg13g2_a22oi_1 _15803_ (.Y(_09054_),
    .B1(net713),
    .B2(\cpu.icache.r_data[1][27] ),
    .A2(net712),
    .A1(\cpu.icache.r_data[2][27] ));
 sg13g2_o21ai_1 _15804_ (.B1(_09054_),
    .Y(_09055_),
    .A1(_08527_),
    .A2(_09053_));
 sg13g2_nor3_1 _15805_ (.A(_09048_),
    .B(_09051_),
    .C(_09055_),
    .Y(_09056_));
 sg13g2_nand2_1 _15806_ (.Y(_09057_),
    .A(_00193_),
    .B(_08913_));
 sg13g2_a22oi_1 _15807_ (.Y(_09058_),
    .B1(net713),
    .B2(\cpu.icache.r_data[1][11] ),
    .A2(net712),
    .A1(\cpu.icache.r_data[2][11] ));
 sg13g2_a22oi_1 _15808_ (.Y(_09059_),
    .B1(net722),
    .B2(\cpu.icache.r_data[3][11] ),
    .A2(net822),
    .A1(\cpu.icache.r_data[5][11] ));
 sg13g2_mux2_1 _15809_ (.A0(\cpu.icache.r_data[4][11] ),
    .A1(\cpu.icache.r_data[6][11] ),
    .S(net1081),
    .X(_09060_));
 sg13g2_a22oi_1 _15810_ (.Y(_09061_),
    .B1(_09060_),
    .B2(_08515_),
    .A2(net937),
    .A1(\cpu.icache.r_data[7][11] ));
 sg13g2_or2_1 _15811_ (.X(_09062_),
    .B(_09061_),
    .A(net938));
 sg13g2_nand4_1 _15812_ (.B(_09058_),
    .C(_09059_),
    .A(net640),
    .Y(_09063_),
    .D(_09062_));
 sg13g2_a21oi_1 _15813_ (.A1(_09057_),
    .A2(_09063_),
    .Y(_09064_),
    .B1(_08906_));
 sg13g2_a21oi_1 _15814_ (.A1(_08967_),
    .A2(_09056_),
    .Y(_09065_),
    .B1(_09064_));
 sg13g2_buf_1 _15815_ (.A(_09065_),
    .X(_09066_));
 sg13g2_inv_2 _15816_ (.Y(_09067_),
    .A(net423));
 sg13g2_mux4_1 _15817_ (.S0(net1079),
    .A0(\cpu.icache.r_data[4][10] ),
    .A1(\cpu.icache.r_data[5][10] ),
    .A2(\cpu.icache.r_data[6][10] ),
    .A3(\cpu.icache.r_data[7][10] ),
    .S1(net813),
    .X(_09068_));
 sg13g2_nand2_1 _15818_ (.Y(_09069_),
    .A(net812),
    .B(_09068_));
 sg13g2_nand2_1 _15819_ (.Y(_09070_),
    .A(\cpu.icache.r_data[1][10] ),
    .B(net723));
 sg13g2_a22oi_1 _15820_ (.Y(_09071_),
    .B1(net641),
    .B2(\cpu.icache.r_data[3][10] ),
    .A2(_08513_),
    .A1(\cpu.icache.r_data[2][10] ));
 sg13g2_and4_1 _15821_ (.A(net582),
    .B(_09069_),
    .C(_09070_),
    .D(_09071_),
    .X(_09072_));
 sg13g2_a21oi_1 _15822_ (.A1(_00191_),
    .A2(_08959_),
    .Y(_09073_),
    .B1(_09072_));
 sg13g2_inv_1 _15823_ (.Y(_09074_),
    .A(_00192_));
 sg13g2_a22oi_1 _15824_ (.Y(_09075_),
    .B1(net643),
    .B2(\cpu.icache.r_data[2][26] ),
    .A2(_08958_),
    .A1(_09074_));
 sg13g2_mux2_1 _15825_ (.A0(\cpu.icache.r_data[4][26] ),
    .A1(\cpu.icache.r_data[6][26] ),
    .S(net813),
    .X(_09076_));
 sg13g2_a22oi_1 _15826_ (.Y(_09077_),
    .B1(_09076_),
    .B2(net805),
    .A2(net806),
    .A1(\cpu.icache.r_data[5][26] ));
 sg13g2_or2_1 _15827_ (.X(_09078_),
    .B(_09077_),
    .A(net721));
 sg13g2_mux2_1 _15828_ (.A0(\cpu.icache.r_data[7][26] ),
    .A1(\cpu.icache.r_data[3][26] ),
    .S(net821),
    .X(_09079_));
 sg13g2_a22oi_1 _15829_ (.Y(_09080_),
    .B1(net820),
    .B2(_09079_),
    .A2(net642),
    .A1(\cpu.icache.r_data[1][26] ));
 sg13g2_nand4_1 _15830_ (.B(_09075_),
    .C(_09078_),
    .A(net1075),
    .Y(_09081_),
    .D(_09080_));
 sg13g2_o21ai_1 _15831_ (.B1(_09081_),
    .Y(_09082_),
    .A1(net929),
    .A2(_09073_));
 sg13g2_buf_1 _15832_ (.A(_09082_),
    .X(_09083_));
 sg13g2_buf_1 _15833_ (.A(_09083_),
    .X(_09084_));
 sg13g2_nor2_2 _15834_ (.A(_09067_),
    .B(_09084_),
    .Y(_09085_));
 sg13g2_nand3_1 _15835_ (.B(_09047_),
    .C(_09085_),
    .A(_09008_),
    .Y(_09086_));
 sg13g2_nor3_1 _15836_ (.A(_08905_),
    .B(_08945_),
    .C(_09086_),
    .Y(_09087_));
 sg13g2_a21o_1 _15837_ (.A2(_08904_),
    .A1(net948),
    .B1(_09087_),
    .X(_00017_));
 sg13g2_buf_2 _15838_ (.A(\cpu.dec.r_op[4] ),
    .X(_09088_));
 sg13g2_inv_1 _15839_ (.Y(_09089_),
    .A(_09088_));
 sg13g2_nand4_1 _15840_ (.B(_08670_),
    .C(_08807_),
    .A(_08618_),
    .Y(_09090_),
    .D(_08877_));
 sg13g2_buf_2 _15841_ (.A(_08634_),
    .X(_09091_));
 sg13g2_xnor2_1 _15842_ (.Y(_09092_),
    .A(net370),
    .B(_08646_));
 sg13g2_or3_1 _15843_ (.A(_09092_),
    .B(_08765_),
    .C(_08785_),
    .X(_09093_));
 sg13g2_nand2b_1 _15844_ (.Y(_09094_),
    .B(_08729_),
    .A_N(_08698_));
 sg13g2_and2_1 _15845_ (.A(_08717_),
    .B(_08740_),
    .X(_09095_));
 sg13g2_nand3b_1 _15846_ (.B(_08726_),
    .C(_09095_),
    .Y(_09096_),
    .A_N(_08707_));
 sg13g2_nor3_1 _15847_ (.A(_08687_),
    .B(_09094_),
    .C(_09096_),
    .Y(_09097_));
 sg13g2_nand4_1 _15848_ (.B(_08856_),
    .C(_08898_),
    .A(_08830_),
    .Y(_09098_),
    .D(_09097_));
 sg13g2_nor4_2 _15849_ (.A(_08581_),
    .B(_09090_),
    .C(_09093_),
    .Y(_09099_),
    .D(_09098_));
 sg13g2_and2_1 _15850_ (.A(_08471_),
    .B(_09099_),
    .X(_09100_));
 sg13g2_buf_1 _15851_ (.A(_09100_),
    .X(_09101_));
 sg13g2_buf_1 _15852_ (.A(_09101_),
    .X(_09102_));
 sg13g2_nor2_1 _15853_ (.A(_00204_),
    .B(net582),
    .Y(_09103_));
 sg13g2_mux2_1 _15854_ (.A0(\cpu.icache.r_data[4][28] ),
    .A1(\cpu.icache.r_data[6][28] ),
    .S(net819),
    .X(_09104_));
 sg13g2_a22oi_1 _15855_ (.Y(_09105_),
    .B1(_09104_),
    .B2(net935),
    .A2(net806),
    .A1(\cpu.icache.r_data[5][28] ));
 sg13g2_nor2_1 _15856_ (.A(net821),
    .B(_09105_),
    .Y(_09106_));
 sg13g2_and2_1 _15857_ (.A(net817),
    .B(\cpu.icache.r_data[3][28] ),
    .X(_09107_));
 sg13g2_a21oi_1 _15858_ (.A1(net812),
    .A2(\cpu.icache.r_data[7][28] ),
    .Y(_09108_),
    .B1(_09107_));
 sg13g2_a22oi_1 _15859_ (.Y(_09109_),
    .B1(net723),
    .B2(\cpu.icache.r_data[1][28] ),
    .A2(net725),
    .A1(\cpu.icache.r_data[2][28] ));
 sg13g2_o21ai_1 _15860_ (.B1(_09109_),
    .Y(_09110_),
    .A1(_08527_),
    .A2(_09108_));
 sg13g2_nor4_1 _15861_ (.A(net1076),
    .B(_09103_),
    .C(_09106_),
    .D(_09110_),
    .Y(_09111_));
 sg13g2_nand2_1 _15862_ (.Y(_09112_),
    .A(_00203_),
    .B(net637));
 sg13g2_a22oi_1 _15863_ (.Y(_09113_),
    .B1(net723),
    .B2(\cpu.icache.r_data[1][12] ),
    .A2(net725),
    .A1(\cpu.icache.r_data[2][12] ));
 sg13g2_a22oi_1 _15864_ (.Y(_09114_),
    .B1(net641),
    .B2(\cpu.icache.r_data[3][12] ),
    .A2(net822),
    .A1(\cpu.icache.r_data[5][12] ));
 sg13g2_mux2_1 _15865_ (.A0(\cpu.icache.r_data[4][12] ),
    .A1(\cpu.icache.r_data[6][12] ),
    .S(net936),
    .X(_09115_));
 sg13g2_a22oi_1 _15866_ (.Y(_09116_),
    .B1(_09115_),
    .B2(net935),
    .A2(net937),
    .A1(\cpu.icache.r_data[7][12] ));
 sg13g2_or2_1 _15867_ (.X(_09117_),
    .B(_09116_),
    .A(net817));
 sg13g2_nand4_1 _15868_ (.B(_09113_),
    .C(_09114_),
    .A(net582),
    .Y(_09118_),
    .D(_09117_));
 sg13g2_a21oi_1 _15869_ (.A1(_09112_),
    .A2(_09118_),
    .Y(_09119_),
    .B1(net1075));
 sg13g2_or2_1 _15870_ (.X(_09120_),
    .B(_09119_),
    .A(_09111_));
 sg13g2_buf_2 _15871_ (.A(_09120_),
    .X(_09121_));
 sg13g2_buf_1 _15872_ (.A(_09121_),
    .X(_09122_));
 sg13g2_buf_1 _15873_ (.A(_09008_),
    .X(_09123_));
 sg13g2_nor2b_1 _15874_ (.A(_09026_),
    .B_N(_09045_),
    .Y(_09124_));
 sg13g2_buf_1 _15875_ (.A(_09124_),
    .X(_09125_));
 sg13g2_buf_1 _15876_ (.A(_09125_),
    .X(_09126_));
 sg13g2_nand3_1 _15877_ (.B(_09085_),
    .C(net170),
    .A(net149),
    .Y(_09127_));
 sg13g2_buf_1 _15878_ (.A(_09127_),
    .X(_09128_));
 sg13g2_or4_1 _15879_ (.A(_08902_),
    .B(_08945_),
    .C(net291),
    .D(_09128_),
    .X(_09129_));
 sg13g2_o21ai_1 _15880_ (.B1(_09129_),
    .Y(_00015_),
    .A1(_09089_),
    .A2(net150));
 sg13g2_buf_2 _15881_ (.A(\cpu.dec.r_op[5] ),
    .X(_09130_));
 sg13g2_nand2_1 _15882_ (.Y(_09131_),
    .A(_09123_),
    .B(_09047_));
 sg13g2_nor4_1 _15883_ (.A(net173),
    .B(_09131_),
    .C(net423),
    .D(net292),
    .Y(_09132_));
 sg13g2_a21o_1 _15884_ (.A2(_08904_),
    .A1(_09130_),
    .B1(_09132_),
    .X(_00016_));
 sg13g2_buf_1 _15885_ (.A(\cpu.dec.r_op[7] ),
    .X(_09133_));
 sg13g2_buf_1 _15886_ (.A(_08903_),
    .X(_09134_));
 sg13g2_nor4_1 _15887_ (.A(net173),
    .B(_08922_),
    .C(_08943_),
    .D(_09128_),
    .Y(_09135_));
 sg13g2_a21o_1 _15888_ (.A2(_09134_),
    .A1(_09133_),
    .B1(_09135_),
    .X(_00018_));
 sg13g2_buf_1 _15889_ (.A(\cpu.dec.r_op[3] ),
    .X(_09136_));
 sg13g2_inv_2 _15890_ (.Y(_09137_),
    .A(net1140));
 sg13g2_buf_1 _15891_ (.A(_09101_),
    .X(_09138_));
 sg13g2_inv_1 _15892_ (.Y(_09139_),
    .A(_09121_));
 sg13g2_buf_1 _15893_ (.A(net149),
    .X(_09140_));
 sg13g2_nand2_1 _15894_ (.Y(_09141_),
    .A(net126),
    .B(_09085_));
 sg13g2_buf_1 _15895_ (.A(_08942_),
    .X(_09142_));
 sg13g2_nand2_1 _15896_ (.Y(_09143_),
    .A(_08922_),
    .B(net369));
 sg13g2_nor3_1 _15897_ (.A(net290),
    .B(_09141_),
    .C(_09143_),
    .Y(_09144_));
 sg13g2_nand3_1 _15898_ (.B(net171),
    .C(_09144_),
    .A(net147),
    .Y(_09145_));
 sg13g2_o21ai_1 _15899_ (.B1(_09145_),
    .Y(_00014_),
    .A1(_09137_),
    .A2(net150));
 sg13g2_buf_1 _15900_ (.A(\cpu.dec.r_op[2] ),
    .X(_09146_));
 sg13g2_inv_2 _15901_ (.Y(_09147_),
    .A(_09146_));
 sg13g2_buf_1 _15902_ (.A(_09101_),
    .X(_09148_));
 sg13g2_or3_1 _15903_ (.A(_08922_),
    .B(_09086_),
    .C(net290),
    .X(_09149_));
 sg13g2_nand2_1 _15904_ (.Y(_09150_),
    .A(net423),
    .B(net292));
 sg13g2_or2_1 _15905_ (.X(_09151_),
    .B(_09150_),
    .A(_09131_));
 sg13g2_o21ai_1 _15906_ (.B1(_09151_),
    .Y(_09152_),
    .A1(_08943_),
    .A2(_09149_));
 sg13g2_nand2_1 _15907_ (.Y(_09153_),
    .A(net146),
    .B(_09152_));
 sg13g2_o21ai_1 _15908_ (.B1(_09153_),
    .Y(_00013_),
    .A1(_09147_),
    .A2(_09102_));
 sg13g2_nor2b_1 _15909_ (.A(r_reset),
    .B_N(net1),
    .Y(_09154_));
 sg13g2_buf_2 _15910_ (.A(_09154_),
    .X(_09155_));
 sg13g2_buf_1 _15911_ (.A(_09155_),
    .X(_09156_));
 sg13g2_buf_1 _15912_ (.A(net928),
    .X(_09157_));
 sg13g2_buf_1 _15913_ (.A(net803),
    .X(_09158_));
 sg13g2_buf_1 _15914_ (.A(net708),
    .X(_09159_));
 sg13g2_buf_2 _15915_ (.A(\cpu.ex.r_ie ),
    .X(_09160_));
 sg13g2_buf_1 _15916_ (.A(\cpu.intr.r_timer ),
    .X(_09161_));
 sg13g2_buf_1 _15917_ (.A(\cpu.intr.r_enable[2] ),
    .X(_09162_));
 sg13g2_buf_1 _15918_ (.A(\cpu.intr.r_swi ),
    .X(_09163_));
 sg13g2_a22oi_1 _15919_ (.Y(_09164_),
    .B1(\cpu.intr.r_enable[3] ),
    .B2(_09163_),
    .A2(_09162_),
    .A1(_09161_));
 sg13g2_buf_2 _15920_ (.A(\cpu.uart.r_x_int ),
    .X(_09165_));
 sg13g2_buf_2 _15921_ (.A(\cpu.uart.r_r_int ),
    .X(_09166_));
 sg13g2_buf_1 _15922_ (.A(\cpu.intr.r_enable[0] ),
    .X(_09167_));
 sg13g2_o21ai_1 _15923_ (.B1(_09167_),
    .Y(_09168_),
    .A1(_09165_),
    .A2(_09166_));
 sg13g2_buf_1 _15924_ (.A(\cpu.intr.r_enable[1] ),
    .X(_09169_));
 sg13g2_buf_2 _15925_ (.A(\cpu.intr.spi_intr ),
    .X(_09170_));
 sg13g2_a22oi_1 _15926_ (.Y(_09171_),
    .B1(_09170_),
    .B2(\cpu.intr.r_enable[5] ),
    .A2(_09169_),
    .A1(\cpu.intr.r_clock ));
 sg13g2_nand3_1 _15927_ (.B(_09168_),
    .C(_09171_),
    .A(_09164_),
    .Y(_09172_));
 sg13g2_and2_1 _15928_ (.A(_09160_),
    .B(_09172_),
    .X(_09173_));
 sg13g2_buf_1 _15929_ (.A(_09173_),
    .X(_09174_));
 sg13g2_buf_2 _15930_ (.A(ui_in[6]),
    .X(_09175_));
 sg13g2_nand2_1 _15931_ (.Y(_09176_),
    .A(\cpu.gpio.r_enable_in[6] ),
    .B(_09175_));
 sg13g2_buf_2 _15932_ (.A(ui_in[4]),
    .X(_09177_));
 sg13g2_nand2_1 _15933_ (.Y(_09178_),
    .A(\cpu.gpio.r_enable_in[4] ),
    .B(_09177_));
 sg13g2_buf_2 _15934_ (.A(\cpu.gpio.r_enable_in[0] ),
    .X(_09179_));
 sg13g2_buf_2 _15935_ (.A(ui_in[0]),
    .X(_09180_));
 sg13g2_buf_1 _15936_ (.A(\cpu.gpio.r_enable_in[1] ),
    .X(_09181_));
 sg13g2_buf_2 _15937_ (.A(ui_in[1]),
    .X(_09182_));
 sg13g2_a22oi_1 _15938_ (.Y(_09183_),
    .B1(_09181_),
    .B2(_09182_),
    .A2(_09180_),
    .A1(_09179_));
 sg13g2_and3_1 _15939_ (.X(_09184_),
    .A(_09176_),
    .B(_09178_),
    .C(_09183_));
 sg13g2_buf_1 _15940_ (.A(\cpu.gpio.r_enable_in[7] ),
    .X(_09185_));
 sg13g2_buf_2 _15941_ (.A(ui_in[7]),
    .X(_09186_));
 sg13g2_buf_2 _15942_ (.A(\cpu.gpio.r_enable_io[6] ),
    .X(_09187_));
 sg13g2_buf_1 _15943_ (.A(uio_in[6]),
    .X(_09188_));
 sg13g2_a22oi_1 _15944_ (.Y(_09189_),
    .B1(_09187_),
    .B2(_09188_),
    .A2(_09186_),
    .A1(_09185_));
 sg13g2_buf_2 _15945_ (.A(ui_in[2]),
    .X(_09190_));
 sg13g2_buf_2 _15946_ (.A(uio_in[7]),
    .X(_09191_));
 sg13g2_a22oi_1 _15947_ (.Y(_09192_),
    .B1(\cpu.gpio.r_enable_io[7] ),
    .B2(_09191_),
    .A2(_09190_),
    .A1(\cpu.gpio.r_enable_in[2] ));
 sg13g2_buf_2 _15948_ (.A(ui_in[5]),
    .X(_09193_));
 sg13g2_buf_1 _15949_ (.A(\cpu.gpio.r_enable_io[5] ),
    .X(_09194_));
 sg13g2_buf_2 _15950_ (.A(uio_in[5]),
    .X(_09195_));
 sg13g2_a22oi_1 _15951_ (.Y(_09196_),
    .B1(_09194_),
    .B2(_09195_),
    .A2(_09193_),
    .A1(\cpu.gpio.r_enable_in[5] ));
 sg13g2_buf_1 _15952_ (.A(\cpu.gpio.r_enable_in[3] ),
    .X(_09197_));
 sg13g2_buf_2 _15953_ (.A(ui_in[3]),
    .X(_09198_));
 sg13g2_buf_2 _15954_ (.A(\cpu.gpio.r_enable_io[4] ),
    .X(_09199_));
 sg13g2_buf_2 _15955_ (.A(uio_in[4]),
    .X(_09200_));
 sg13g2_a22oi_1 _15956_ (.Y(_09201_),
    .B1(_09199_),
    .B2(_09200_),
    .A2(_09198_),
    .A1(_09197_));
 sg13g2_and4_1 _15957_ (.A(_09189_),
    .B(_09192_),
    .C(_09196_),
    .D(_09201_),
    .X(_09202_));
 sg13g2_buf_1 _15958_ (.A(\cpu.intr.r_enable[4] ),
    .X(_09203_));
 sg13g2_nand2_1 _15959_ (.Y(_09204_),
    .A(_09203_),
    .B(_09160_));
 sg13g2_a21oi_2 _15960_ (.B1(_09204_),
    .Y(_09205_),
    .A2(_09202_),
    .A1(_09184_));
 sg13g2_or2_1 _15961_ (.X(_09206_),
    .B(_09205_),
    .A(_09174_));
 sg13g2_buf_1 _15962_ (.A(_09206_),
    .X(_09207_));
 sg13g2_buf_1 _15963_ (.A(\cpu.dec.r_trap ),
    .X(_09208_));
 sg13g2_or2_1 _15964_ (.X(_09209_),
    .B(net371),
    .A(_09208_));
 sg13g2_buf_1 _15965_ (.A(_09209_),
    .X(_09210_));
 sg13g2_a21oi_2 _15966_ (.B1(_09210_),
    .Y(_09211_),
    .A2(_09207_),
    .A1(_08403_));
 sg13g2_nand2b_2 _15967_ (.Y(_09212_),
    .B(_09211_),
    .A_N(_00187_));
 sg13g2_inv_2 _15968_ (.Y(_09213_),
    .A(net1144));
 sg13g2_buf_1 _15969_ (.A(_08420_),
    .X(_09214_));
 sg13g2_nand2_1 _15970_ (.Y(_09215_),
    .A(net1145),
    .B(net1074));
 sg13g2_o21ai_1 _15971_ (.B1(_09215_),
    .Y(_09216_),
    .A1(net1145),
    .A2(net1143));
 sg13g2_nand2b_1 _15972_ (.Y(_09217_),
    .B(net1143),
    .A_N(net1074));
 sg13g2_o21ai_1 _15973_ (.B1(_09217_),
    .Y(_09218_),
    .A1(_09213_),
    .A2(_09216_));
 sg13g2_buf_1 _15974_ (.A(_09218_),
    .X(_09219_));
 sg13g2_buf_2 _15975_ (.A(\cpu.addr[6] ),
    .X(_09220_));
 sg13g2_buf_1 _15976_ (.A(\cpu.addr[8] ),
    .X(_09221_));
 sg13g2_buf_1 _15977_ (.A(\cpu.addr[7] ),
    .X(_09222_));
 sg13g2_inv_2 _15978_ (.Y(_09223_),
    .A(net1138));
 sg13g2_nor2_2 _15979_ (.A(net1139),
    .B(_09223_),
    .Y(_09224_));
 sg13g2_nand2_2 _15980_ (.Y(_09225_),
    .A(_09220_),
    .B(_09224_));
 sg13g2_buf_1 _15981_ (.A(_00207_),
    .X(_09226_));
 sg13g2_buf_2 _15982_ (.A(\cpu.addr[1] ),
    .X(_09227_));
 sg13g2_buf_1 _15983_ (.A(_09227_),
    .X(_09228_));
 sg13g2_buf_2 _15984_ (.A(\cpu.addr[2] ),
    .X(_09229_));
 sg13g2_buf_1 _15985_ (.A(_09229_),
    .X(_09230_));
 sg13g2_buf_2 _15986_ (.A(_09230_),
    .X(_09231_));
 sg13g2_buf_1 _15987_ (.A(net927),
    .X(_09232_));
 sg13g2_buf_2 _15988_ (.A(net802),
    .X(_09233_));
 sg13g2_buf_1 _15989_ (.A(net707),
    .X(_09234_));
 sg13g2_nor2_2 _15990_ (.A(net1073),
    .B(net633),
    .Y(_09235_));
 sg13g2_nand2_2 _15991_ (.Y(_09236_),
    .A(_09226_),
    .B(_09235_));
 sg13g2_nor4_2 _15992_ (.A(_09212_),
    .B(_09219_),
    .C(_09225_),
    .Y(_09237_),
    .D(_09236_));
 sg13g2_buf_1 _15993_ (.A(\cpu.spi.r_state[1] ),
    .X(_09238_));
 sg13g2_buf_8 _15994_ (.A(\cpu.addr[3] ),
    .X(_09239_));
 sg13g2_inv_2 _15995_ (.Y(_09240_),
    .A(net1136));
 sg13g2_buf_1 _15996_ (.A(_09240_),
    .X(_09241_));
 sg13g2_inv_1 _15997_ (.Y(_09242_),
    .A(\cpu.ex.r_wmask[1] ));
 sg13g2_inv_1 _15998_ (.Y(_09243_),
    .A(_08341_));
 sg13g2_nand2_1 _15999_ (.Y(_09244_),
    .A(_09242_),
    .B(_09243_));
 sg13g2_nand3_1 _16000_ (.B(_09244_),
    .C(_09211_),
    .A(_08340_),
    .Y(_09245_));
 sg13g2_buf_2 _16001_ (.A(_09245_),
    .X(_09246_));
 sg13g2_nor2_1 _16002_ (.A(_09225_),
    .B(_09246_),
    .Y(_09247_));
 sg13g2_buf_1 _16003_ (.A(_09247_),
    .X(_09248_));
 sg13g2_nand2_2 _16004_ (.Y(_09249_),
    .A(net926),
    .B(_09248_));
 sg13g2_nand2_1 _16005_ (.Y(_09250_),
    .A(net1137),
    .B(_09249_));
 sg13g2_buf_1 _16006_ (.A(\cpu.spi.r_state[6] ),
    .X(_09251_));
 sg13g2_buf_1 _16007_ (.A(_09251_),
    .X(_09252_));
 sg13g2_buf_1 _16008_ (.A(\cpu.spi.r_bits[0] ),
    .X(_09253_));
 sg13g2_buf_1 _16009_ (.A(\cpu.spi.r_bits[1] ),
    .X(_09254_));
 sg13g2_nor3_1 _16010_ (.A(_09253_),
    .B(_09254_),
    .C(\cpu.spi.r_bits[2] ),
    .Y(_09255_));
 sg13g2_nor3_2 _16011_ (.A(\cpu.spi.r_timeout_count[0] ),
    .B(\cpu.spi.r_timeout_count[1] ),
    .C(\cpu.spi.r_timeout_count[2] ),
    .Y(_09256_));
 sg13g2_nor2b_1 _16012_ (.A(\cpu.spi.r_timeout_count[3] ),
    .B_N(_09256_),
    .Y(_09257_));
 sg13g2_nand2b_1 _16013_ (.Y(_09258_),
    .B(_09257_),
    .A_N(\cpu.spi.r_timeout_count[4] ));
 sg13g2_nor2_1 _16014_ (.A(\cpu.spi.r_timeout_count[5] ),
    .B(_09258_),
    .Y(_09259_));
 sg13g2_nand2b_1 _16015_ (.Y(_09260_),
    .B(_09259_),
    .A_N(\cpu.spi.r_timeout_count[6] ));
 sg13g2_buf_1 _16016_ (.A(_09260_),
    .X(_09261_));
 sg13g2_o21ai_1 _16017_ (.B1(\cpu.spi.r_searching ),
    .Y(_09262_),
    .A1(\cpu.spi.r_timeout_count[7] ),
    .A2(_09261_));
 sg13g2_nand2_1 _16018_ (.Y(_09263_),
    .A(_09255_),
    .B(_09262_));
 sg13g2_buf_1 _16019_ (.A(\cpu.spi.r_in[3] ),
    .X(_09264_));
 sg13g2_buf_1 _16020_ (.A(\cpu.spi.r_in[6] ),
    .X(_09265_));
 sg13g2_buf_1 _16021_ (.A(\cpu.spi.r_in[1] ),
    .X(_09266_));
 sg13g2_buf_1 _16022_ (.A(\cpu.spi.r_in[0] ),
    .X(_09267_));
 sg13g2_nand2_1 _16023_ (.Y(_09268_),
    .A(_09266_),
    .B(_09267_));
 sg13g2_nand3_1 _16024_ (.B(_09265_),
    .C(_09268_),
    .A(_09264_),
    .Y(_09269_));
 sg13g2_buf_1 _16025_ (.A(\cpu.spi.r_in[2] ),
    .X(_09270_));
 sg13g2_buf_1 _16026_ (.A(\cpu.spi.r_in[5] ),
    .X(_09271_));
 sg13g2_buf_1 _16027_ (.A(\cpu.spi.r_in[4] ),
    .X(_09272_));
 sg13g2_nand4_1 _16028_ (.B(_09271_),
    .C(_09272_),
    .A(_09270_),
    .Y(_09273_),
    .D(\cpu.spi.r_in[7] ));
 sg13g2_nor2_1 _16029_ (.A(_09269_),
    .B(_09273_),
    .Y(_09274_));
 sg13g2_o21ai_1 _16030_ (.B1(\cpu.spi.r_searching ),
    .Y(_09275_),
    .A1(_00206_),
    .A2(_09274_));
 sg13g2_nand2_2 _16031_ (.Y(_09276_),
    .A(_09263_),
    .B(_09275_));
 sg13g2_buf_1 _16032_ (.A(\cpu.spi.r_count[7] ),
    .X(_09277_));
 sg13g2_buf_1 _16033_ (.A(\cpu.spi.r_count[3] ),
    .X(_09278_));
 sg13g2_buf_1 _16034_ (.A(\cpu.spi.r_count[0] ),
    .X(_09279_));
 sg13g2_nor2_1 _16035_ (.A(_09279_),
    .B(\cpu.spi.r_count[1] ),
    .Y(_09280_));
 sg13g2_nand2b_1 _16036_ (.Y(_09281_),
    .B(_09280_),
    .A_N(\cpu.spi.r_count[2] ));
 sg13g2_nor3_1 _16037_ (.A(_09278_),
    .B(\cpu.spi.r_count[4] ),
    .C(_09281_),
    .Y(_09282_));
 sg13g2_nor2b_1 _16038_ (.A(\cpu.spi.r_count[5] ),
    .B_N(_09282_),
    .Y(_09283_));
 sg13g2_nor2b_1 _16039_ (.A(\cpu.spi.r_count[6] ),
    .B_N(_09283_),
    .Y(_09284_));
 sg13g2_nor2b_1 _16040_ (.A(_09277_),
    .B_N(_09284_),
    .Y(_09285_));
 sg13g2_buf_1 _16041_ (.A(_09285_),
    .X(_09286_));
 sg13g2_nand3_1 _16042_ (.B(_09276_),
    .C(net517),
    .A(net1071),
    .Y(_09287_));
 sg13g2_o21ai_1 _16043_ (.B1(_09287_),
    .Y(_09288_),
    .A1(_09237_),
    .A2(_09250_));
 sg13g2_and2_1 _16044_ (.A(net634),
    .B(_09288_),
    .X(_00030_));
 sg13g2_buf_1 _16045_ (.A(net1137),
    .X(_09289_));
 sg13g2_buf_1 _16046_ (.A(net1070),
    .X(_09290_));
 sg13g2_buf_1 _16047_ (.A(net1136),
    .X(_09291_));
 sg13g2_buf_1 _16048_ (.A(net1069),
    .X(_09292_));
 sg13g2_buf_1 _16049_ (.A(net924),
    .X(_09293_));
 sg13g2_buf_1 _16050_ (.A(net801),
    .X(_09294_));
 sg13g2_buf_1 _16051_ (.A(net706),
    .X(_09295_));
 sg13g2_buf_2 _16052_ (.A(net632),
    .X(_09296_));
 sg13g2_buf_2 _16053_ (.A(net578),
    .X(_09297_));
 sg13g2_buf_2 _16054_ (.A(net516),
    .X(_09298_));
 sg13g2_or2_1 _16055_ (.X(_09299_),
    .B(_09246_),
    .A(_09225_));
 sg13g2_buf_1 _16056_ (.A(_09299_),
    .X(_09300_));
 sg13g2_nor2_1 _16057_ (.A(net463),
    .B(_09300_),
    .Y(_09301_));
 sg13g2_buf_1 _16058_ (.A(_09301_),
    .X(_09302_));
 sg13g2_buf_1 _16059_ (.A(net100),
    .X(_09303_));
 sg13g2_inv_1 _16060_ (.Y(_09304_),
    .A(_09251_));
 sg13g2_buf_1 _16061_ (.A(\cpu.spi.r_state[4] ),
    .X(_09305_));
 sg13g2_nand2b_1 _16062_ (.Y(_09306_),
    .B(_09284_),
    .A_N(_09277_));
 sg13g2_buf_1 _16063_ (.A(_09306_),
    .X(_09307_));
 sg13g2_buf_1 _16064_ (.A(_09307_),
    .X(_09308_));
 sg13g2_buf_1 _16065_ (.A(net462),
    .X(_09309_));
 sg13g2_nor3_1 _16066_ (.A(\cpu.spi.r_state[5] ),
    .B(net1135),
    .C(net422),
    .Y(_09310_));
 sg13g2_o21ai_1 _16067_ (.B1(_09310_),
    .Y(_09311_),
    .A1(_09304_),
    .A2(_09276_));
 sg13g2_a21oi_1 _16068_ (.A1(_09290_),
    .A2(net91),
    .Y(_09312_),
    .B1(_09311_));
 sg13g2_buf_1 _16069_ (.A(\cpu.spi.r_state[2] ),
    .X(_09313_));
 sg13g2_o21ai_1 _16070_ (.B1(net708),
    .Y(_09314_),
    .A1(net1134),
    .A2(_09286_));
 sg13g2_nor2_1 _16071_ (.A(_09312_),
    .B(_09314_),
    .Y(_00031_));
 sg13g2_nand2b_1 _16072_ (.Y(_09315_),
    .B(net1),
    .A_N(r_reset));
 sg13g2_buf_2 _16073_ (.A(_09315_),
    .X(_09316_));
 sg13g2_buf_2 _16074_ (.A(_09316_),
    .X(_09317_));
 sg13g2_buf_1 _16075_ (.A(net923),
    .X(_09318_));
 sg13g2_inv_2 _16076_ (.Y(_09319_),
    .A(net1137));
 sg13g2_nor2_1 _16077_ (.A(_09319_),
    .B(_09301_),
    .Y(_09320_));
 sg13g2_buf_2 _16078_ (.A(\cpu.spi.r_state[3] ),
    .X(_09321_));
 sg13g2_a21oi_1 _16079_ (.A1(_09237_),
    .A2(_09320_),
    .Y(_09322_),
    .B1(_09321_));
 sg13g2_nor3_1 _16080_ (.A(net800),
    .B(net517),
    .C(_09322_),
    .Y(_00032_));
 sg13g2_buf_1 _16081_ (.A(net800),
    .X(_09323_));
 sg13g2_nor2_1 _16082_ (.A(_09236_),
    .B(_09300_),
    .Y(_09324_));
 sg13g2_buf_2 _16083_ (.A(\cpu.spi.r_state[0] ),
    .X(_09325_));
 sg13g2_a22oi_1 _16084_ (.Y(_09326_),
    .B1(_09324_),
    .B2(_09325_),
    .A2(net422),
    .A1(net1135));
 sg13g2_nor2_1 _16085_ (.A(net705),
    .B(_09326_),
    .Y(_00033_));
 sg13g2_a21oi_1 _16086_ (.A1(_09290_),
    .A2(_09303_),
    .Y(_09327_),
    .B1(\cpu.spi.r_state[5] ));
 sg13g2_nor3_1 _16087_ (.A(net800),
    .B(_09286_),
    .C(_09327_),
    .Y(_00034_));
 sg13g2_nand2_1 _16088_ (.Y(_09328_),
    .A(net1071),
    .B(net422));
 sg13g2_nand2_1 _16089_ (.Y(_09329_),
    .A(net1134),
    .B(net517));
 sg13g2_buf_2 _16090_ (.A(net923),
    .X(_09330_));
 sg13g2_buf_1 _16091_ (.A(_09330_),
    .X(_09331_));
 sg13g2_a21oi_1 _16092_ (.A1(_09328_),
    .A2(_09329_),
    .Y(_00035_),
    .B1(net704));
 sg13g2_buf_1 _16093_ (.A(\cpu.ex.r_mult_off[0] ),
    .X(_09332_));
 sg13g2_buf_2 _16094_ (.A(\cpu.dec.mult ),
    .X(_09333_));
 sg13g2_inv_1 _16095_ (.Y(_09334_),
    .A(_09333_));
 sg13g2_nand3b_1 _16096_ (.B(\cpu.dec.iready ),
    .C(_00189_),
    .Y(_09335_),
    .A_N(\cpu.ex.r_branch_stall ));
 sg13g2_buf_2 _16097_ (.A(_09335_),
    .X(_09336_));
 sg13g2_nor3_1 _16098_ (.A(_09334_),
    .B(_09316_),
    .C(_09336_),
    .Y(_09337_));
 sg13g2_buf_2 _16099_ (.A(_09337_),
    .X(_09338_));
 sg13g2_inv_1 _16100_ (.Y(_09339_),
    .A(\cpu.dec.div ));
 sg13g2_nor3_1 _16101_ (.A(_09339_),
    .B(_09316_),
    .C(_09336_),
    .Y(_09340_));
 sg13g2_nor2_1 _16102_ (.A(_09338_),
    .B(_09340_),
    .Y(_09341_));
 sg13g2_buf_2 _16103_ (.A(_09341_),
    .X(_09342_));
 sg13g2_and2_1 _16104_ (.A(_09332_),
    .B(_09342_),
    .X(_09343_));
 sg13g2_buf_2 _16105_ (.A(_09343_),
    .X(_09344_));
 sg13g2_inv_4 _16106_ (.A(_09344_),
    .Y(\cpu.ex.c_mult_off[0] ));
 sg13g2_buf_1 _16107_ (.A(\cpu.ex.r_div_running ),
    .X(_09345_));
 sg13g2_buf_1 _16108_ (.A(\cpu.ex.r_mult_off[1] ),
    .X(_09346_));
 sg13g2_buf_1 _16109_ (.A(_09346_),
    .X(_09347_));
 sg13g2_buf_1 _16110_ (.A(\cpu.ex.r_mult_off[2] ),
    .X(_09348_));
 sg13g2_buf_1 _16111_ (.A(\cpu.ex.r_mult_off[3] ),
    .X(_09349_));
 sg13g2_nor4_2 _16112_ (.A(net1068),
    .B(_09348_),
    .C(_09349_),
    .Y(_09350_),
    .D(\cpu.ex.c_mult_off[0] ));
 sg13g2_buf_1 _16113_ (.A(_09340_),
    .X(_09351_));
 sg13g2_o21ai_1 _16114_ (.B1(_09155_),
    .Y(_09352_),
    .A1(_09345_),
    .A2(net799));
 sg13g2_a21oi_1 _16115_ (.A1(_09345_),
    .A2(_09350_),
    .Y(\cpu.ex.c_div_running ),
    .B1(_09352_));
 sg13g2_buf_1 _16116_ (.A(\cpu.ex.r_mult_running ),
    .X(_09353_));
 sg13g2_buf_1 _16117_ (.A(_09338_),
    .X(_09354_));
 sg13g2_o21ai_1 _16118_ (.B1(_09155_),
    .Y(_09355_),
    .A1(net1133),
    .A2(net703));
 sg13g2_a21oi_1 _16119_ (.A1(net1133),
    .A2(_09350_),
    .Y(\cpu.ex.c_mult_running ),
    .B1(_09355_));
 sg13g2_o21ai_1 _16120_ (.B1(_09325_),
    .Y(_09356_),
    .A1(_09236_),
    .A2(_09300_));
 sg13g2_buf_1 _16121_ (.A(_09356_),
    .X(_09357_));
 sg13g2_and2_1 _16122_ (.A(_09155_),
    .B(_09357_),
    .X(_09358_));
 sg13g2_buf_1 _16123_ (.A(_09358_),
    .X(_09359_));
 sg13g2_o21ai_1 _16124_ (.B1(_09359_),
    .Y(_00029_),
    .A1(net422),
    .A2(_09322_));
 sg13g2_inv_1 _16125_ (.Y(_09360_),
    .A(\cpu.qspi.r_state[17] ));
 sg13g2_buf_2 _16126_ (.A(\cpu.dcache.flush_write ),
    .X(_09361_));
 sg13g2_inv_1 _16127_ (.Y(_09362_),
    .A(_09361_));
 sg13g2_buf_2 _16128_ (.A(net826),
    .X(_09363_));
 sg13g2_buf_8 _16129_ (.A(_08365_),
    .X(_09364_));
 sg13g2_buf_8 _16130_ (.A(_09364_),
    .X(_09365_));
 sg13g2_buf_2 _16131_ (.A(_09365_),
    .X(_09366_));
 sg13g2_buf_8 _16132_ (.A(_08364_),
    .X(_09367_));
 sg13g2_buf_1 _16133_ (.A(_09367_),
    .X(_09368_));
 sg13g2_buf_8 _16134_ (.A(net700),
    .X(_09369_));
 sg13g2_mux4_1 _16135_ (.S0(net701),
    .A0(\cpu.genblk1.mmu.r_vtop_d[8][0] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[9][0] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[10][0] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[11][0] ),
    .S1(net631),
    .X(_09370_));
 sg13g2_mux4_1 _16136_ (.S0(net701),
    .A0(\cpu.genblk1.mmu.r_vtop_d[0][0] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[1][0] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[2][0] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[3][0] ),
    .S1(_09369_),
    .X(_09371_));
 sg13g2_mux4_1 _16137_ (.S0(net701),
    .A0(\cpu.genblk1.mmu.r_vtop_d[12][0] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[13][0] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[14][0] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[15][0] ),
    .S1(net631),
    .X(_09372_));
 sg13g2_mux4_1 _16138_ (.S0(net701),
    .A0(\cpu.genblk1.mmu.r_vtop_d[4][0] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[5][0] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[6][0] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[7][0] ),
    .S1(net631),
    .X(_09373_));
 sg13g2_buf_8 _16139_ (.A(_08385_),
    .X(_09374_));
 sg13g2_buf_2 _16140_ (.A(net797),
    .X(_09375_));
 sg13g2_buf_2 _16141_ (.A(net945),
    .X(_09376_));
 sg13g2_mux4_1 _16142_ (.S0(net699),
    .A0(_09370_),
    .A1(_09371_),
    .A2(_09372_),
    .A3(_09373_),
    .S1(_09376_),
    .X(_09377_));
 sg13g2_buf_1 _16143_ (.A(_08349_),
    .X(_09378_));
 sg13g2_buf_2 _16144_ (.A(_08365_),
    .X(_09379_));
 sg13g2_buf_2 _16145_ (.A(net922),
    .X(_09380_));
 sg13g2_buf_8 _16146_ (.A(_09367_),
    .X(_09381_));
 sg13g2_buf_2 _16147_ (.A(net698),
    .X(_09382_));
 sg13g2_mux4_1 _16148_ (.S0(net794),
    .A0(\cpu.genblk1.mmu.r_vtop_d[24][0] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[25][0] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[26][0] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[27][0] ),
    .S1(net630),
    .X(_09383_));
 sg13g2_buf_8 _16149_ (.A(_09364_),
    .X(_09384_));
 sg13g2_buf_8 _16150_ (.A(net793),
    .X(_09385_));
 sg13g2_mux4_1 _16151_ (.S0(net697),
    .A0(\cpu.genblk1.mmu.r_vtop_d[16][0] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[17][0] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[18][0] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[19][0] ),
    .S1(net630),
    .X(_09386_));
 sg13g2_buf_1 _16152_ (.A(_09367_),
    .X(_09387_));
 sg13g2_buf_1 _16153_ (.A(net696),
    .X(_09388_));
 sg13g2_mux4_1 _16154_ (.S0(_09380_),
    .A0(\cpu.genblk1.mmu.r_vtop_d[28][0] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[29][0] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[30][0] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[31][0] ),
    .S1(net629),
    .X(_09389_));
 sg13g2_mux4_1 _16155_ (.S0(_09380_),
    .A0(\cpu.genblk1.mmu.r_vtop_d[20][0] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[21][0] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[22][0] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[23][0] ),
    .S1(net629),
    .X(_09390_));
 sg13g2_buf_2 _16156_ (.A(net797),
    .X(_09391_));
 sg13g2_mux4_1 _16157_ (.S0(_09391_),
    .A0(_09383_),
    .A1(_09386_),
    .A2(_09389_),
    .A3(_09390_),
    .S1(net796),
    .X(_09392_));
 sg13g2_and2_1 _16158_ (.A(net795),
    .B(_09392_),
    .X(_09393_));
 sg13g2_a21oi_1 _16159_ (.A1(net702),
    .A2(_09377_),
    .Y(_09394_),
    .B1(_09393_));
 sg13g2_nor2_1 _16160_ (.A(_08475_),
    .B(net701),
    .Y(_09395_));
 sg13g2_a21oi_1 _16161_ (.A1(_08475_),
    .A2(_09394_),
    .Y(_09396_),
    .B1(_09395_));
 sg13g2_buf_1 _16162_ (.A(_09396_),
    .X(_09397_));
 sg13g2_inv_1 _16163_ (.Y(_09398_),
    .A(_00227_));
 sg13g2_buf_2 _16164_ (.A(_00212_),
    .X(_09399_));
 sg13g2_inv_1 _16165_ (.Y(_09400_),
    .A(_09399_));
 sg13g2_nor2_1 _16166_ (.A(_09229_),
    .B(net1136),
    .Y(_09401_));
 sg13g2_buf_1 _16167_ (.A(_09401_),
    .X(_09402_));
 sg13g2_buf_2 _16168_ (.A(\cpu.addr[4] ),
    .X(_09403_));
 sg13g2_inv_1 _16169_ (.Y(_09404_),
    .A(_09403_));
 sg13g2_buf_1 _16170_ (.A(_09404_),
    .X(_09405_));
 sg13g2_o21ai_1 _16171_ (.B1(_09405_),
    .Y(_09406_),
    .A1(_09400_),
    .A2(_09402_));
 sg13g2_buf_2 _16172_ (.A(_09406_),
    .X(_09407_));
 sg13g2_buf_1 _16173_ (.A(_09407_),
    .X(_09408_));
 sg13g2_inv_1 _16174_ (.Y(_09409_),
    .A(net1072));
 sg13g2_and2_1 _16175_ (.A(net1136),
    .B(_09399_),
    .X(_09410_));
 sg13g2_buf_1 _16176_ (.A(_09410_),
    .X(_09411_));
 sg13g2_and2_1 _16177_ (.A(_09409_),
    .B(net919),
    .X(_09412_));
 sg13g2_buf_2 _16178_ (.A(_09412_),
    .X(_09413_));
 sg13g2_buf_1 _16179_ (.A(_09399_),
    .X(_09414_));
 sg13g2_nor2b_1 _16180_ (.A(\cpu.addr[3] ),
    .B_N(_09229_),
    .Y(_09415_));
 sg13g2_buf_1 _16181_ (.A(_09415_),
    .X(_09416_));
 sg13g2_and2_1 _16182_ (.A(_09414_),
    .B(net918),
    .X(_09417_));
 sg13g2_buf_2 _16183_ (.A(_09417_),
    .X(_09418_));
 sg13g2_buf_1 _16184_ (.A(_09418_),
    .X(_09419_));
 sg13g2_a22oi_1 _16185_ (.Y(_09420_),
    .B1(net627),
    .B2(\cpu.dcache.r_tag[1][12] ),
    .A2(_09413_),
    .A1(\cpu.dcache.r_tag[2][12] ));
 sg13g2_buf_1 _16186_ (.A(_09409_),
    .X(_09421_));
 sg13g2_nor3_1 _16187_ (.A(net792),
    .B(net920),
    .C(_09240_),
    .Y(_09422_));
 sg13g2_buf_2 _16188_ (.A(_09422_),
    .X(_09423_));
 sg13g2_and2_1 _16189_ (.A(net1072),
    .B(net919),
    .X(_09424_));
 sg13g2_buf_2 _16190_ (.A(_09424_),
    .X(_09425_));
 sg13g2_a22oi_1 _16191_ (.Y(_09426_),
    .B1(_09425_),
    .B2(\cpu.dcache.r_tag[3][12] ),
    .A2(_09423_),
    .A1(\cpu.dcache.r_tag[7][12] ));
 sg13g2_mux2_1 _16192_ (.A0(\cpu.dcache.r_tag[4][12] ),
    .A1(\cpu.dcache.r_tag[6][12] ),
    .S(net801),
    .X(_09427_));
 sg13g2_buf_1 _16193_ (.A(net792),
    .X(_09428_));
 sg13g2_a22oi_1 _16194_ (.Y(_09429_),
    .B1(_09427_),
    .B2(net694),
    .A2(net918),
    .A1(\cpu.dcache.r_tag[5][12] ));
 sg13g2_buf_1 _16195_ (.A(_09403_),
    .X(_09430_));
 sg13g2_buf_1 _16196_ (.A(net1066),
    .X(_09431_));
 sg13g2_nand2b_1 _16197_ (.Y(_09432_),
    .B(net917),
    .A_N(_09429_));
 sg13g2_nand4_1 _16198_ (.B(_09420_),
    .C(_09426_),
    .A(net628),
    .Y(_09433_),
    .D(_09432_));
 sg13g2_o21ai_1 _16199_ (.B1(_09433_),
    .Y(_09434_),
    .A1(_09398_),
    .A2(net628));
 sg13g2_xor2_1 _16200_ (.B(_09434_),
    .A(_09397_),
    .X(_09435_));
 sg13g2_mux4_1 _16201_ (.S0(net701),
    .A0(\cpu.genblk1.mmu.r_vtop_d[8][1] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[9][1] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[10][1] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[11][1] ),
    .S1(net631),
    .X(_09436_));
 sg13g2_mux4_1 _16202_ (.S0(_09366_),
    .A0(\cpu.genblk1.mmu.r_vtop_d[0][1] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[1][1] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[2][1] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[3][1] ),
    .S1(net631),
    .X(_09437_));
 sg13g2_mux4_1 _16203_ (.S0(net697),
    .A0(\cpu.genblk1.mmu.r_vtop_d[12][1] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[13][1] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[14][1] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[15][1] ),
    .S1(net631),
    .X(_09438_));
 sg13g2_mux4_1 _16204_ (.S0(_09366_),
    .A0(\cpu.genblk1.mmu.r_vtop_d[4][1] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[5][1] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[6][1] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[7][1] ),
    .S1(net631),
    .X(_09439_));
 sg13g2_mux4_1 _16205_ (.S0(_09375_),
    .A0(_09436_),
    .A1(_09437_),
    .A2(_09438_),
    .A3(_09439_),
    .S1(_09376_),
    .X(_09440_));
 sg13g2_mux4_1 _16206_ (.S0(net794),
    .A0(\cpu.genblk1.mmu.r_vtop_d[24][1] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[25][1] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[26][1] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[27][1] ),
    .S1(net629),
    .X(_09441_));
 sg13g2_mux4_1 _16207_ (.S0(net794),
    .A0(\cpu.genblk1.mmu.r_vtop_d[16][1] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[17][1] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[18][1] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[19][1] ),
    .S1(net629),
    .X(_09442_));
 sg13g2_mux4_1 _16208_ (.S0(net794),
    .A0(\cpu.genblk1.mmu.r_vtop_d[28][1] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[29][1] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[30][1] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[31][1] ),
    .S1(_09388_),
    .X(_09443_));
 sg13g2_mux4_1 _16209_ (.S0(net794),
    .A0(\cpu.genblk1.mmu.r_vtop_d[20][1] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[21][1] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[22][1] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[23][1] ),
    .S1(_09388_),
    .X(_09444_));
 sg13g2_mux4_1 _16210_ (.S0(net695),
    .A0(_09441_),
    .A1(_09442_),
    .A2(_09443_),
    .A3(_09444_),
    .S1(net796),
    .X(_09445_));
 sg13g2_and2_1 _16211_ (.A(net795),
    .B(_09445_),
    .X(_09446_));
 sg13g2_a21oi_1 _16212_ (.A1(net702),
    .A2(_09440_),
    .Y(_09447_),
    .B1(_09446_));
 sg13g2_buf_1 _16213_ (.A(net631),
    .X(_09448_));
 sg13g2_nor2_1 _16214_ (.A(net1149),
    .B(net577),
    .Y(_09449_));
 sg13g2_a21oi_1 _16215_ (.A1(net1083),
    .A2(_09447_),
    .Y(_09450_),
    .B1(_09449_));
 sg13g2_buf_1 _16216_ (.A(_09450_),
    .X(_09451_));
 sg13g2_and2_1 _16217_ (.A(net1072),
    .B(net1136),
    .X(_09452_));
 sg13g2_buf_2 _16218_ (.A(_09452_),
    .X(_09453_));
 sg13g2_mux2_1 _16219_ (.A0(\cpu.dcache.r_tag[4][13] ),
    .A1(\cpu.dcache.r_tag[6][13] ),
    .S(net801),
    .X(_09454_));
 sg13g2_a22oi_1 _16220_ (.Y(_09455_),
    .B1(_09454_),
    .B2(net694),
    .A2(_09453_),
    .A1(\cpu.dcache.r_tag[7][13] ));
 sg13g2_buf_1 _16221_ (.A(net917),
    .X(_09456_));
 sg13g2_nand2b_1 _16222_ (.Y(_09457_),
    .B(net791),
    .A_N(_09455_));
 sg13g2_buf_1 _16223_ (.A(net1136),
    .X(_09458_));
 sg13g2_nor3_1 _16224_ (.A(_09409_),
    .B(_09404_),
    .C(net1065),
    .Y(_09459_));
 sg13g2_buf_2 _16225_ (.A(_09459_),
    .X(_09460_));
 sg13g2_mux2_1 _16226_ (.A0(\cpu.dcache.r_tag[2][13] ),
    .A1(\cpu.dcache.r_tag[3][13] ),
    .S(net707),
    .X(_09461_));
 sg13g2_buf_1 _16227_ (.A(_09411_),
    .X(_09462_));
 sg13g2_a22oi_1 _16228_ (.Y(_09463_),
    .B1(_09461_),
    .B2(net790),
    .A2(_09460_),
    .A1(\cpu.dcache.r_tag[5][13] ));
 sg13g2_nand2_1 _16229_ (.Y(_09464_),
    .A(\cpu.dcache.r_tag[1][13] ),
    .B(net627));
 sg13g2_or2_1 _16230_ (.X(_09465_),
    .B(_09239_),
    .A(_09229_));
 sg13g2_a21oi_1 _16231_ (.A1(_09399_),
    .A2(_09465_),
    .Y(_09466_),
    .B1(_09403_));
 sg13g2_buf_2 _16232_ (.A(_09466_),
    .X(_09467_));
 sg13g2_buf_1 _16233_ (.A(_09467_),
    .X(_09468_));
 sg13g2_nand2b_1 _16234_ (.Y(_09469_),
    .B(_09468_),
    .A_N(_00228_));
 sg13g2_nand4_1 _16235_ (.B(_09463_),
    .C(_09464_),
    .A(_09457_),
    .Y(_09470_),
    .D(_09469_));
 sg13g2_xnor2_1 _16236_ (.Y(_09471_),
    .A(_09451_),
    .B(_09470_));
 sg13g2_buf_2 _16237_ (.A(_09364_),
    .X(_09472_));
 sg13g2_buf_2 _16238_ (.A(_09367_),
    .X(_09473_));
 sg13g2_mux4_1 _16239_ (.S0(net789),
    .A0(\cpu.genblk1.mmu.r_vtop_d[24][8] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[25][8] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[26][8] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[27][8] ),
    .S1(net692),
    .X(_09474_));
 sg13g2_buf_2 _16240_ (.A(_09364_),
    .X(_09475_));
 sg13g2_buf_1 _16241_ (.A(net696),
    .X(_09476_));
 sg13g2_mux4_1 _16242_ (.S0(net788),
    .A0(\cpu.genblk1.mmu.r_vtop_d[16][8] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[17][8] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[18][8] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[19][8] ),
    .S1(net626),
    .X(_09477_));
 sg13g2_buf_2 _16243_ (.A(_09367_),
    .X(_09478_));
 sg13g2_mux4_1 _16244_ (.S0(net798),
    .A0(\cpu.genblk1.mmu.r_vtop_d[28][8] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[29][8] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[30][8] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[31][8] ),
    .S1(net691),
    .X(_09479_));
 sg13g2_buf_2 _16245_ (.A(_09364_),
    .X(_09480_));
 sg13g2_mux4_1 _16246_ (.S0(net787),
    .A0(\cpu.genblk1.mmu.r_vtop_d[20][8] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[21][8] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[22][8] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[23][8] ),
    .S1(net691),
    .X(_09481_));
 sg13g2_buf_2 _16247_ (.A(net945),
    .X(_09482_));
 sg13g2_mux4_1 _16248_ (.S0(net695),
    .A0(_09474_),
    .A1(_09477_),
    .A2(_09479_),
    .A3(_09481_),
    .S1(net786),
    .X(_09483_));
 sg13g2_nand2_1 _16249_ (.Y(_09484_),
    .A(net795),
    .B(_09483_));
 sg13g2_mux4_1 _16250_ (.S0(net787),
    .A0(\cpu.genblk1.mmu.r_vtop_d[8][8] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[9][8] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[10][8] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[11][8] ),
    .S1(net691),
    .X(_09485_));
 sg13g2_mux4_1 _16251_ (.S0(net789),
    .A0(\cpu.genblk1.mmu.r_vtop_d[0][8] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[1][8] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[2][8] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[3][8] ),
    .S1(net692),
    .X(_09486_));
 sg13g2_buf_1 _16252_ (.A(_09367_),
    .X(_09487_));
 sg13g2_mux4_1 _16253_ (.S0(_09365_),
    .A0(\cpu.genblk1.mmu.r_vtop_d[12][8] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[13][8] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[14][8] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[15][8] ),
    .S1(net690),
    .X(_09488_));
 sg13g2_mux4_1 _16254_ (.S0(net798),
    .A0(\cpu.genblk1.mmu.r_vtop_d[4][8] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[5][8] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[6][8] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[7][8] ),
    .S1(net690),
    .X(_09489_));
 sg13g2_mux4_1 _16255_ (.S0(net797),
    .A0(_09485_),
    .A1(_09486_),
    .A2(_09488_),
    .A3(_09489_),
    .S1(net786),
    .X(_09490_));
 sg13g2_nand2_1 _16256_ (.Y(_09491_),
    .A(net702),
    .B(_09490_));
 sg13g2_a21oi_2 _16257_ (.B1(_08582_),
    .Y(_09492_),
    .A2(_09491_),
    .A1(_09484_));
 sg13g2_buf_1 _16258_ (.A(_09492_),
    .X(_09493_));
 sg13g2_buf_1 _16259_ (.A(net1067),
    .X(_09494_));
 sg13g2_a22oi_1 _16260_ (.Y(_09495_),
    .B1(\cpu.dcache.r_tag[1][20] ),
    .B2(net916),
    .A2(\cpu.dcache.r_tag[5][20] ),
    .A1(net1066));
 sg13g2_inv_1 _16261_ (.Y(_09496_),
    .A(_09495_));
 sg13g2_nor2b_1 _16262_ (.A(_09229_),
    .B_N(_09403_),
    .Y(_09497_));
 sg13g2_buf_1 _16263_ (.A(_09497_),
    .X(_09498_));
 sg13g2_a22oi_1 _16264_ (.Y(_09499_),
    .B1(net915),
    .B2(\cpu.dcache.r_tag[4][20] ),
    .A2(_09496_),
    .A1(net802));
 sg13g2_or2_1 _16265_ (.X(_09500_),
    .B(_09499_),
    .A(net801));
 sg13g2_nand2_1 _16266_ (.Y(_09501_),
    .A(\cpu.dcache.r_tag[7][20] ),
    .B(_09423_));
 sg13g2_and2_1 _16267_ (.A(net1069),
    .B(net915),
    .X(_09502_));
 sg13g2_buf_1 _16268_ (.A(_09502_),
    .X(_09503_));
 sg13g2_mux2_1 _16269_ (.A0(\cpu.dcache.r_tag[2][20] ),
    .A1(\cpu.dcache.r_tag[3][20] ),
    .S(net802),
    .X(_09504_));
 sg13g2_a22oi_1 _16270_ (.Y(_09505_),
    .B1(net790),
    .B2(_09504_),
    .A2(_09503_),
    .A1(\cpu.dcache.r_tag[6][20] ));
 sg13g2_nand4_1 _16271_ (.B(_09500_),
    .C(_09501_),
    .A(net628),
    .Y(_09506_),
    .D(_09505_));
 sg13g2_o21ai_1 _16272_ (.B1(_09506_),
    .Y(_09507_),
    .A1(\cpu.dcache.r_tag[0][20] ),
    .A2(net628));
 sg13g2_xnor2_1 _16273_ (.Y(_09508_),
    .A(net368),
    .B(_09507_));
 sg13g2_mux4_1 _16274_ (.S0(net789),
    .A0(\cpu.genblk1.mmu.r_vtop_d[24][7] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[25][7] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[26][7] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[27][7] ),
    .S1(net626),
    .X(_09509_));
 sg13g2_mux4_1 _16275_ (.S0(net788),
    .A0(\cpu.genblk1.mmu.r_vtop_d[16][7] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[17][7] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[18][7] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[19][7] ),
    .S1(net626),
    .X(_09510_));
 sg13g2_mux4_1 _16276_ (.S0(_09480_),
    .A0(\cpu.genblk1.mmu.r_vtop_d[28][7] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[29][7] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[30][7] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[31][7] ),
    .S1(_09478_),
    .X(_09511_));
 sg13g2_mux4_1 _16277_ (.S0(net787),
    .A0(\cpu.genblk1.mmu.r_vtop_d[20][7] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[21][7] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[22][7] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[23][7] ),
    .S1(net691),
    .X(_09512_));
 sg13g2_mux4_1 _16278_ (.S0(net695),
    .A0(_09509_),
    .A1(_09510_),
    .A2(_09511_),
    .A3(_09512_),
    .S1(net786),
    .X(_09513_));
 sg13g2_nand2_1 _16279_ (.Y(_09514_),
    .A(net795),
    .B(_09513_));
 sg13g2_mux4_1 _16280_ (.S0(net789),
    .A0(\cpu.genblk1.mmu.r_vtop_d[8][7] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[9][7] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[10][7] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[11][7] ),
    .S1(net692),
    .X(_09515_));
 sg13g2_mux4_1 _16281_ (.S0(_09472_),
    .A0(\cpu.genblk1.mmu.r_vtop_d[0][7] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[1][7] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[2][7] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[3][7] ),
    .S1(_09473_),
    .X(_09516_));
 sg13g2_mux4_1 _16282_ (.S0(net798),
    .A0(\cpu.genblk1.mmu.r_vtop_d[12][7] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[13][7] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[14][7] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[15][7] ),
    .S1(net690),
    .X(_09517_));
 sg13g2_mux4_1 _16283_ (.S0(net798),
    .A0(\cpu.genblk1.mmu.r_vtop_d[4][7] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[5][7] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[6][7] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[7][7] ),
    .S1(net690),
    .X(_09518_));
 sg13g2_mux4_1 _16284_ (.S0(_09374_),
    .A0(_09515_),
    .A1(_09516_),
    .A2(_09517_),
    .A3(_09518_),
    .S1(net786),
    .X(_09519_));
 sg13g2_nand2_1 _16285_ (.Y(_09520_),
    .A(net702),
    .B(_09519_));
 sg13g2_a21oi_2 _16286_ (.B1(_08582_),
    .Y(_09521_),
    .A2(_09520_),
    .A1(_09514_));
 sg13g2_buf_1 _16287_ (.A(_09521_),
    .X(_09522_));
 sg13g2_inv_1 _16288_ (.Y(_09523_),
    .A(_00234_));
 sg13g2_a22oi_1 _16289_ (.Y(_09524_),
    .B1(_09413_),
    .B2(\cpu.dcache.r_tag[2][19] ),
    .A2(_09425_),
    .A1(\cpu.dcache.r_tag[3][19] ));
 sg13g2_a22oi_1 _16290_ (.Y(_09525_),
    .B1(net627),
    .B2(\cpu.dcache.r_tag[1][19] ),
    .A2(_09460_),
    .A1(\cpu.dcache.r_tag[5][19] ));
 sg13g2_mux2_1 _16291_ (.A0(\cpu.dcache.r_tag[4][19] ),
    .A1(\cpu.dcache.r_tag[6][19] ),
    .S(net1065),
    .X(_09526_));
 sg13g2_a22oi_1 _16292_ (.Y(_09527_),
    .B1(_09453_),
    .B2(\cpu.dcache.r_tag[7][19] ),
    .A2(_09526_),
    .A1(net792));
 sg13g2_nand2b_1 _16293_ (.Y(_09528_),
    .B(net917),
    .A_N(_09527_));
 sg13g2_nand4_1 _16294_ (.B(_09524_),
    .C(_09525_),
    .A(net628),
    .Y(_09529_),
    .D(_09528_));
 sg13g2_o21ai_1 _16295_ (.B1(_09529_),
    .Y(_09530_),
    .A1(_09523_),
    .A2(net628));
 sg13g2_xnor2_1 _16296_ (.Y(_09531_),
    .A(net367),
    .B(_09530_));
 sg13g2_mux4_1 _16297_ (.S0(net788),
    .A0(\cpu.genblk1.mmu.r_vtop_d[24][6] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[25][6] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[26][6] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[27][6] ),
    .S1(net626),
    .X(_09532_));
 sg13g2_mux4_1 _16298_ (.S0(net788),
    .A0(\cpu.genblk1.mmu.r_vtop_d[16][6] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[17][6] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[18][6] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[19][6] ),
    .S1(net626),
    .X(_09533_));
 sg13g2_mux4_1 _16299_ (.S0(net787),
    .A0(\cpu.genblk1.mmu.r_vtop_d[28][6] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[29][6] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[30][6] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[31][6] ),
    .S1(net692),
    .X(_09534_));
 sg13g2_mux4_1 _16300_ (.S0(net789),
    .A0(\cpu.genblk1.mmu.r_vtop_d[20][6] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[21][6] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[22][6] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[23][6] ),
    .S1(net692),
    .X(_09535_));
 sg13g2_mux4_1 _16301_ (.S0(net695),
    .A0(_09532_),
    .A1(_09533_),
    .A2(_09534_),
    .A3(_09535_),
    .S1(net786),
    .X(_09536_));
 sg13g2_nand2_1 _16302_ (.Y(_09537_),
    .A(_09378_),
    .B(_09536_));
 sg13g2_mux4_1 _16303_ (.S0(_09475_),
    .A0(\cpu.genblk1.mmu.r_vtop_d[8][6] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[9][6] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[10][6] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[11][6] ),
    .S1(_09476_),
    .X(_09538_));
 sg13g2_mux4_1 _16304_ (.S0(_09475_),
    .A0(\cpu.genblk1.mmu.r_vtop_d[0][6] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[1][6] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[2][6] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[3][6] ),
    .S1(_09476_),
    .X(_09539_));
 sg13g2_mux4_1 _16305_ (.S0(_09480_),
    .A0(\cpu.genblk1.mmu.r_vtop_d[12][6] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[13][6] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[14][6] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[15][6] ),
    .S1(_09478_),
    .X(_09540_));
 sg13g2_mux4_1 _16306_ (.S0(net787),
    .A0(\cpu.genblk1.mmu.r_vtop_d[4][6] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[5][6] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[6][6] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[7][6] ),
    .S1(net691),
    .X(_09541_));
 sg13g2_mux4_1 _16307_ (.S0(net695),
    .A0(_09538_),
    .A1(_09539_),
    .A2(_09540_),
    .A3(_09541_),
    .S1(net786),
    .X(_09542_));
 sg13g2_nand2_1 _16308_ (.Y(_09543_),
    .A(net702),
    .B(_09542_));
 sg13g2_a21oi_2 _16309_ (.B1(_08582_),
    .Y(_09544_),
    .A2(_09543_),
    .A1(_09537_));
 sg13g2_buf_1 _16310_ (.A(_09544_),
    .X(_09545_));
 sg13g2_nor2b_1 _16311_ (.A(net1072),
    .B_N(net1136),
    .Y(_09546_));
 sg13g2_buf_1 _16312_ (.A(_09546_),
    .X(_09547_));
 sg13g2_mux2_1 _16313_ (.A0(\cpu.dcache.r_tag[5][18] ),
    .A1(\cpu.dcache.r_tag[7][18] ),
    .S(net924),
    .X(_09548_));
 sg13g2_a22oi_1 _16314_ (.Y(_09549_),
    .B1(_09548_),
    .B2(net802),
    .A2(net785),
    .A1(\cpu.dcache.r_tag[6][18] ));
 sg13g2_nand2b_1 _16315_ (.Y(_09550_),
    .B(net917),
    .A_N(_09549_));
 sg13g2_and2_1 _16316_ (.A(_09240_),
    .B(_09498_),
    .X(_09551_));
 sg13g2_buf_2 _16317_ (.A(_09551_),
    .X(_09552_));
 sg13g2_mux2_1 _16318_ (.A0(\cpu.dcache.r_tag[2][18] ),
    .A1(\cpu.dcache.r_tag[3][18] ),
    .S(net802),
    .X(_09553_));
 sg13g2_a22oi_1 _16319_ (.Y(_09554_),
    .B1(_09553_),
    .B2(_09462_),
    .A2(_09552_),
    .A1(\cpu.dcache.r_tag[4][18] ));
 sg13g2_nand2_1 _16320_ (.Y(_09555_),
    .A(\cpu.dcache.r_tag[1][18] ),
    .B(net627));
 sg13g2_nand2b_1 _16321_ (.Y(_09556_),
    .B(net693),
    .A_N(_00233_));
 sg13g2_nand4_1 _16322_ (.B(_09554_),
    .C(_09555_),
    .A(_09550_),
    .Y(_09557_),
    .D(_09556_));
 sg13g2_xor2_1 _16323_ (.B(_09557_),
    .A(net366),
    .X(_09558_));
 sg13g2_nor2_1 _16324_ (.A(_09409_),
    .B(net920),
    .Y(_09559_));
 sg13g2_buf_1 _16325_ (.A(_09559_),
    .X(_09560_));
 sg13g2_mux2_1 _16326_ (.A0(\cpu.dcache.r_tag[5][10] ),
    .A1(\cpu.dcache.r_tag[7][10] ),
    .S(net924),
    .X(_09561_));
 sg13g2_a22oi_1 _16327_ (.Y(_09562_),
    .B1(\cpu.dcache.r_tag[2][10] ),
    .B2(net916),
    .A2(\cpu.dcache.r_tag[6][10] ),
    .A1(net1066));
 sg13g2_nand3_1 _16328_ (.B(net916),
    .C(\cpu.dcache.r_tag[3][10] ),
    .A(net927),
    .Y(_09563_));
 sg13g2_o21ai_1 _16329_ (.B1(_09563_),
    .Y(_09564_),
    .A1(net802),
    .A2(_09562_));
 sg13g2_and2_1 _16330_ (.A(net1072),
    .B(net916),
    .X(_09565_));
 sg13g2_a22oi_1 _16331_ (.Y(_09566_),
    .B1(_09565_),
    .B2(\cpu.dcache.r_tag[1][10] ),
    .A2(net915),
    .A1(\cpu.dcache.r_tag[4][10] ));
 sg13g2_nor2_1 _16332_ (.A(_09293_),
    .B(_09566_),
    .Y(_09567_));
 sg13g2_a221oi_1 _16333_ (.B2(_09293_),
    .C1(_09567_),
    .B1(_09564_),
    .A1(net689),
    .Y(_09568_),
    .A2(_09561_));
 sg13g2_mux2_1 _16334_ (.A0(_00224_),
    .A1(_09568_),
    .S(_09407_),
    .X(_09569_));
 sg13g2_xnor2_1 _16335_ (.Y(_09570_),
    .A(_00223_),
    .B(_09569_));
 sg13g2_inv_1 _16336_ (.Y(_09571_),
    .A(_00215_));
 sg13g2_and2_1 _16337_ (.A(net1065),
    .B(\cpu.dcache.r_tag[6][6] ),
    .X(_09572_));
 sg13g2_a21oi_1 _16338_ (.A1(_09240_),
    .A2(\cpu.dcache.r_tag[4][6] ),
    .Y(_09573_),
    .B1(_09572_));
 sg13g2_nand2_1 _16339_ (.Y(_09574_),
    .A(\cpu.dcache.r_tag[7][6] ),
    .B(_09453_));
 sg13g2_o21ai_1 _16340_ (.B1(_09574_),
    .Y(_09575_),
    .A1(net802),
    .A2(_09573_));
 sg13g2_a22oi_1 _16341_ (.Y(_09576_),
    .B1(\cpu.dcache.r_tag[1][6] ),
    .B2(net916),
    .A2(\cpu.dcache.r_tag[5][6] ),
    .A1(net1066));
 sg13g2_nand2_1 _16342_ (.Y(_09577_),
    .A(\cpu.dcache.r_tag[3][6] ),
    .B(net919));
 sg13g2_o21ai_1 _16343_ (.B1(_09577_),
    .Y(_09578_),
    .A1(net801),
    .A2(_09576_));
 sg13g2_a22oi_1 _16344_ (.Y(_09579_),
    .B1(_09578_),
    .B2(_09232_),
    .A2(_09575_),
    .A1(_09431_));
 sg13g2_nor2_1 _16345_ (.A(_09430_),
    .B(net1065),
    .Y(_09580_));
 sg13g2_buf_2 _16346_ (.A(_09580_),
    .X(_09581_));
 sg13g2_a21o_1 _16347_ (.A2(net919),
    .A1(\cpu.dcache.r_tag[2][6] ),
    .B1(_09581_),
    .X(_09582_));
 sg13g2_a22oi_1 _16348_ (.Y(_09583_),
    .B1(_09582_),
    .B2(net694),
    .A2(_09400_),
    .A1(_09405_));
 sg13g2_a22oi_1 _16349_ (.Y(_09584_),
    .B1(_09579_),
    .B2(_09583_),
    .A2(net693),
    .A1(_00216_));
 sg13g2_xnor2_1 _16350_ (.Y(_09585_),
    .A(_09571_),
    .B(_09584_));
 sg13g2_a22oi_1 _16351_ (.Y(_09586_),
    .B1(\cpu.dcache.r_tag[1][11] ),
    .B2(_09494_),
    .A2(\cpu.dcache.r_tag[5][11] ),
    .A1(net1066));
 sg13g2_nand2_1 _16352_ (.Y(_09587_),
    .A(\cpu.dcache.r_tag[4][11] ),
    .B(_09498_));
 sg13g2_o21ai_1 _16353_ (.B1(_09587_),
    .Y(_09588_),
    .A1(net792),
    .A2(_09586_));
 sg13g2_mux2_1 _16354_ (.A0(\cpu.dcache.r_tag[2][11] ),
    .A1(\cpu.dcache.r_tag[3][11] ),
    .S(net1072),
    .X(_09589_));
 sg13g2_and4_1 _16355_ (.A(net927),
    .B(net1066),
    .C(_09458_),
    .D(\cpu.dcache.r_tag[7][11] ),
    .X(_09590_));
 sg13g2_a21o_1 _16356_ (.A2(_09589_),
    .A1(net919),
    .B1(_09590_),
    .X(_09591_));
 sg13g2_a221oi_1 _16357_ (.B2(_09240_),
    .C1(_09591_),
    .B1(_09588_),
    .A1(\cpu.dcache.r_tag[6][11] ),
    .Y(_09592_),
    .A2(_09503_));
 sg13g2_mux2_1 _16358_ (.A0(_00226_),
    .A1(_09592_),
    .S(_09407_),
    .X(_09593_));
 sg13g2_xnor2_1 _16359_ (.Y(_09594_),
    .A(_00225_),
    .B(_09593_));
 sg13g2_a22oi_1 _16360_ (.Y(_09595_),
    .B1(\cpu.dcache.r_tag[3][9] ),
    .B2(net1067),
    .A2(\cpu.dcache.r_tag[7][9] ),
    .A1(_09403_));
 sg13g2_a221oi_1 _16361_ (.B2(net1067),
    .C1(_09230_),
    .B1(\cpu.dcache.r_tag[2][9] ),
    .A1(_09403_),
    .Y(_09596_),
    .A2(\cpu.dcache.r_tag[6][9] ));
 sg13g2_a21oi_1 _16362_ (.A1(net927),
    .A2(_09595_),
    .Y(_09597_),
    .B1(_09596_));
 sg13g2_nor2b_1 _16363_ (.A(net1069),
    .B_N(_09403_),
    .Y(_09598_));
 sg13g2_mux2_1 _16364_ (.A0(\cpu.dcache.r_tag[4][9] ),
    .A1(\cpu.dcache.r_tag[5][9] ),
    .S(net1072),
    .X(_09599_));
 sg13g2_and2_1 _16365_ (.A(_09598_),
    .B(_09599_),
    .X(_09600_));
 sg13g2_a221oi_1 _16366_ (.B2(net924),
    .C1(_09600_),
    .B1(_09597_),
    .A1(\cpu.dcache.r_tag[1][9] ),
    .Y(_09601_),
    .A2(_09418_));
 sg13g2_mux2_1 _16367_ (.A0(_00222_),
    .A1(_09601_),
    .S(_09407_),
    .X(_09602_));
 sg13g2_xor2_1 _16368_ (.B(_09602_),
    .A(_00221_),
    .X(_09603_));
 sg13g2_buf_1 _16369_ (.A(_00213_),
    .X(_09604_));
 sg13g2_mux2_1 _16370_ (.A0(\cpu.dcache.r_tag[4][5] ),
    .A1(\cpu.dcache.r_tag[6][5] ),
    .S(net1065),
    .X(_09605_));
 sg13g2_a22oi_1 _16371_ (.Y(_09606_),
    .B1(_09605_),
    .B2(_09421_),
    .A2(_09453_),
    .A1(\cpu.dcache.r_tag[7][5] ));
 sg13g2_inv_1 _16372_ (.Y(_09607_),
    .A(_00214_));
 sg13g2_a22oi_1 _16373_ (.Y(_09608_),
    .B1(\cpu.dcache.r_tag[1][5] ),
    .B2(net1067),
    .A2(\cpu.dcache.r_tag[5][5] ),
    .A1(net1066));
 sg13g2_nand3_1 _16374_ (.B(net1067),
    .C(\cpu.dcache.r_tag[3][5] ),
    .A(net1069),
    .Y(_09609_));
 sg13g2_o21ai_1 _16375_ (.B1(_09609_),
    .Y(_09610_),
    .A1(net924),
    .A2(_09608_));
 sg13g2_inv_1 _16376_ (.Y(_09611_),
    .A(\cpu.dcache.r_tag[2][5] ));
 sg13g2_nand3b_1 _16377_ (.B(_09239_),
    .C(_09399_),
    .Y(_09612_),
    .A_N(net1072));
 sg13g2_buf_1 _16378_ (.A(_09612_),
    .X(_09613_));
 sg13g2_nor2_1 _16379_ (.A(_09611_),
    .B(_09613_),
    .Y(_09614_));
 sg13g2_a221oi_1 _16380_ (.B2(net927),
    .C1(_09614_),
    .B1(_09610_),
    .A1(_09607_),
    .Y(_09615_),
    .A2(_09467_));
 sg13g2_o21ai_1 _16381_ (.B1(_09615_),
    .Y(_09616_),
    .A1(net920),
    .A2(_09606_));
 sg13g2_xnor2_1 _16382_ (.Y(_09617_),
    .A(_09604_),
    .B(_09616_));
 sg13g2_mux2_1 _16383_ (.A0(\cpu.dcache.r_tag[4][8] ),
    .A1(\cpu.dcache.r_tag[6][8] ),
    .S(net1065),
    .X(_09618_));
 sg13g2_a22oi_1 _16384_ (.Y(_09619_),
    .B1(_09618_),
    .B2(net792),
    .A2(_09453_),
    .A1(\cpu.dcache.r_tag[7][8] ));
 sg13g2_inv_1 _16385_ (.Y(_09620_),
    .A(_00220_));
 sg13g2_a22oi_1 _16386_ (.Y(_09621_),
    .B1(\cpu.dcache.r_tag[1][8] ),
    .B2(net1067),
    .A2(\cpu.dcache.r_tag[5][8] ),
    .A1(_09430_));
 sg13g2_nand3_1 _16387_ (.B(net1067),
    .C(\cpu.dcache.r_tag[3][8] ),
    .A(net1069),
    .Y(_09622_));
 sg13g2_o21ai_1 _16388_ (.B1(_09622_),
    .Y(_09623_),
    .A1(_09292_),
    .A2(_09621_));
 sg13g2_inv_1 _16389_ (.Y(_09624_),
    .A(\cpu.dcache.r_tag[2][8] ));
 sg13g2_nor2_1 _16390_ (.A(_09624_),
    .B(_09613_),
    .Y(_09625_));
 sg13g2_a221oi_1 _16391_ (.B2(net927),
    .C1(_09625_),
    .B1(_09623_),
    .A1(_09620_),
    .Y(_09626_),
    .A2(_09467_));
 sg13g2_o21ai_1 _16392_ (.B1(_09626_),
    .Y(_09627_),
    .A1(net920),
    .A2(_09619_));
 sg13g2_xnor2_1 _16393_ (.Y(_09628_),
    .A(_00219_),
    .B(_09627_));
 sg13g2_mux2_1 _16394_ (.A0(\cpu.dcache.r_tag[4][7] ),
    .A1(\cpu.dcache.r_tag[6][7] ),
    .S(net1065),
    .X(_09629_));
 sg13g2_a22oi_1 _16395_ (.Y(_09630_),
    .B1(_09629_),
    .B2(net792),
    .A2(_09453_),
    .A1(\cpu.dcache.r_tag[7][7] ));
 sg13g2_inv_1 _16396_ (.Y(_09631_),
    .A(_00218_));
 sg13g2_a22oi_1 _16397_ (.Y(_09632_),
    .B1(\cpu.dcache.r_tag[1][7] ),
    .B2(_09414_),
    .A2(\cpu.dcache.r_tag[5][7] ),
    .A1(net1066));
 sg13g2_nand3_1 _16398_ (.B(net1067),
    .C(\cpu.dcache.r_tag[3][7] ),
    .A(net1065),
    .Y(_09633_));
 sg13g2_o21ai_1 _16399_ (.B1(_09633_),
    .Y(_09634_),
    .A1(_09292_),
    .A2(_09632_));
 sg13g2_inv_1 _16400_ (.Y(_09635_),
    .A(\cpu.dcache.r_tag[2][7] ));
 sg13g2_nor2_1 _16401_ (.A(_09635_),
    .B(_09613_),
    .Y(_09636_));
 sg13g2_a221oi_1 _16402_ (.B2(_09232_),
    .C1(_09636_),
    .B1(_09634_),
    .A1(_09631_),
    .Y(_09637_),
    .A2(_09467_));
 sg13g2_o21ai_1 _16403_ (.B1(_09637_),
    .Y(_09638_),
    .A1(net920),
    .A2(_09630_));
 sg13g2_xnor2_1 _16404_ (.Y(_09639_),
    .A(_00217_),
    .B(_09638_));
 sg13g2_nor4_1 _16405_ (.A(_09603_),
    .B(_09617_),
    .C(_09628_),
    .D(_09639_),
    .Y(_09640_));
 sg13g2_nand4_1 _16406_ (.B(_09585_),
    .C(_09594_),
    .A(_09570_),
    .Y(_09641_),
    .D(_09640_));
 sg13g2_nor4_1 _16407_ (.A(_09508_),
    .B(_09531_),
    .C(_09558_),
    .D(_09641_),
    .Y(_09642_));
 sg13g2_buf_1 _16408_ (.A(net796),
    .X(_09643_));
 sg13g2_buf_8 _16409_ (.A(_09364_),
    .X(_09644_));
 sg13g2_mux4_1 _16410_ (.S0(net784),
    .A0(\cpu.genblk1.mmu.r_vtop_d[16][2] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[17][2] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[18][2] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[19][2] ),
    .S1(net700),
    .X(_09645_));
 sg13g2_mux4_1 _16411_ (.S0(net784),
    .A0(\cpu.genblk1.mmu.r_vtop_d[0][2] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[1][2] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[2][2] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[3][2] ),
    .S1(_09487_),
    .X(_09646_));
 sg13g2_mux4_1 _16412_ (.S0(net784),
    .A0(\cpu.genblk1.mmu.r_vtop_d[24][2] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[25][2] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[26][2] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[27][2] ),
    .S1(net700),
    .X(_09647_));
 sg13g2_mux4_1 _16413_ (.S0(net784),
    .A0(\cpu.genblk1.mmu.r_vtop_d[8][2] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[9][2] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[10][2] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[11][2] ),
    .S1(net700),
    .X(_09648_));
 sg13g2_mux4_1 _16414_ (.S0(net826),
    .A0(_09645_),
    .A1(_09646_),
    .A2(_09647_),
    .A3(_09648_),
    .S1(net1086),
    .X(_09649_));
 sg13g2_nand2_1 _16415_ (.Y(_09650_),
    .A(_08338_),
    .B(_09649_));
 sg13g2_mux4_1 _16416_ (.S0(net798),
    .A0(\cpu.genblk1.mmu.r_vtop_d[20][2] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[21][2] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[22][2] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[23][2] ),
    .S1(net690),
    .X(_09651_));
 sg13g2_mux4_1 _16417_ (.S0(net798),
    .A0(\cpu.genblk1.mmu.r_vtop_d[4][2] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[5][2] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[6][2] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[7][2] ),
    .S1(net690),
    .X(_09652_));
 sg13g2_mux4_1 _16418_ (.S0(net784),
    .A0(\cpu.genblk1.mmu.r_vtop_d[28][2] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[29][2] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[30][2] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[31][2] ),
    .S1(net700),
    .X(_09653_));
 sg13g2_mux4_1 _16419_ (.S0(net784),
    .A0(\cpu.genblk1.mmu.r_vtop_d[12][2] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[13][2] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[14][2] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[15][2] ),
    .S1(_09487_),
    .X(_09654_));
 sg13g2_mux4_1 _16420_ (.S0(net826),
    .A0(_09651_),
    .A1(_09652_),
    .A2(_09653_),
    .A3(_09654_),
    .S1(net1086),
    .X(_09655_));
 sg13g2_o21ai_1 _16421_ (.B1(net796),
    .Y(_09656_),
    .A1(_08339_),
    .A2(_09655_));
 sg13g2_o21ai_1 _16422_ (.B1(_09656_),
    .Y(_09657_),
    .A1(_09643_),
    .A2(_09650_));
 sg13g2_buf_1 _16423_ (.A(_09657_),
    .X(_09658_));
 sg13g2_a22oi_1 _16424_ (.Y(_09659_),
    .B1(_09552_),
    .B2(\cpu.dcache.r_tag[4][14] ),
    .A2(_09418_),
    .A1(\cpu.dcache.r_tag[1][14] ));
 sg13g2_a22oi_1 _16425_ (.Y(_09660_),
    .B1(_09413_),
    .B2(\cpu.dcache.r_tag[2][14] ),
    .A2(_09503_),
    .A1(\cpu.dcache.r_tag[6][14] ));
 sg13g2_mux2_1 _16426_ (.A0(\cpu.dcache.r_tag[5][14] ),
    .A1(\cpu.dcache.r_tag[7][14] ),
    .S(net924),
    .X(_09661_));
 sg13g2_a22oi_1 _16427_ (.Y(_09662_),
    .B1(_09661_),
    .B2(_09559_),
    .A2(_09425_),
    .A1(\cpu.dcache.r_tag[3][14] ));
 sg13g2_and4_1 _16428_ (.A(_09407_),
    .B(_09659_),
    .C(_09660_),
    .D(_09662_),
    .X(_09663_));
 sg13g2_a21oi_1 _16429_ (.A1(_00229_),
    .A2(net693),
    .Y(_09664_),
    .B1(_09663_));
 sg13g2_xor2_1 _16430_ (.B(_09664_),
    .A(_09658_),
    .X(_09665_));
 sg13g2_mux4_1 _16431_ (.S0(_09472_),
    .A0(\cpu.genblk1.mmu.r_vtop_d[24][10] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[25][10] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[26][10] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[27][10] ),
    .S1(_09473_),
    .X(_09666_));
 sg13g2_mux4_1 _16432_ (.S0(net788),
    .A0(\cpu.genblk1.mmu.r_vtop_d[16][10] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[17][10] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[18][10] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[19][10] ),
    .S1(net626),
    .X(_09667_));
 sg13g2_mux4_1 _16433_ (.S0(net787),
    .A0(\cpu.genblk1.mmu.r_vtop_d[28][10] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[29][10] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[30][10] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[31][10] ),
    .S1(net691),
    .X(_09668_));
 sg13g2_mux4_1 _16434_ (.S0(net787),
    .A0(\cpu.genblk1.mmu.r_vtop_d[20][10] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[21][10] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[22][10] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[23][10] ),
    .S1(net691),
    .X(_09669_));
 sg13g2_mux4_1 _16435_ (.S0(net695),
    .A0(_09666_),
    .A1(_09667_),
    .A2(_09668_),
    .A3(_09669_),
    .S1(net786),
    .X(_09670_));
 sg13g2_nand2_1 _16436_ (.Y(_09671_),
    .A(_09378_),
    .B(_09670_));
 sg13g2_mux4_1 _16437_ (.S0(net787),
    .A0(\cpu.genblk1.mmu.r_vtop_d[8][10] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[9][10] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[10][10] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[11][10] ),
    .S1(net691),
    .X(_09672_));
 sg13g2_mux4_1 _16438_ (.S0(net789),
    .A0(\cpu.genblk1.mmu.r_vtop_d[0][10] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[1][10] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[2][10] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[3][10] ),
    .S1(net692),
    .X(_09673_));
 sg13g2_mux4_1 _16439_ (.S0(net798),
    .A0(\cpu.genblk1.mmu.r_vtop_d[12][10] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[13][10] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[14][10] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[15][10] ),
    .S1(net690),
    .X(_09674_));
 sg13g2_mux4_1 _16440_ (.S0(net798),
    .A0(\cpu.genblk1.mmu.r_vtop_d[4][10] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[5][10] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[6][10] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[7][10] ),
    .S1(net690),
    .X(_09675_));
 sg13g2_mux4_1 _16441_ (.S0(_09374_),
    .A0(_09672_),
    .A1(_09673_),
    .A2(_09674_),
    .A3(_09675_),
    .S1(net786),
    .X(_09676_));
 sg13g2_nand2_1 _16442_ (.Y(_09677_),
    .A(net702),
    .B(_09676_));
 sg13g2_a21oi_2 _16443_ (.B1(_08582_),
    .Y(_09678_),
    .A2(_09677_),
    .A1(_09671_));
 sg13g2_buf_1 _16444_ (.A(_09678_),
    .X(_09679_));
 sg13g2_mux2_1 _16445_ (.A0(\cpu.dcache.r_tag[4][22] ),
    .A1(\cpu.dcache.r_tag[6][22] ),
    .S(net801),
    .X(_09680_));
 sg13g2_a22oi_1 _16446_ (.Y(_09681_),
    .B1(_09680_),
    .B2(net917),
    .A2(_09462_),
    .A1(\cpu.dcache.r_tag[2][22] ));
 sg13g2_mux2_1 _16447_ (.A0(\cpu.dcache.r_tag[1][22] ),
    .A1(\cpu.dcache.r_tag[3][22] ),
    .S(net924),
    .X(_09682_));
 sg13g2_mux2_1 _16448_ (.A0(\cpu.dcache.r_tag[5][22] ),
    .A1(\cpu.dcache.r_tag[7][22] ),
    .S(net801),
    .X(_09683_));
 sg13g2_a221oi_1 _16449_ (.B2(net917),
    .C1(net694),
    .B1(_09683_),
    .A1(net916),
    .Y(_09684_),
    .A2(_09682_));
 sg13g2_a21oi_1 _16450_ (.A1(_09428_),
    .A2(_09681_),
    .Y(_09685_),
    .B1(_09684_));
 sg13g2_a21oi_1 _16451_ (.A1(\cpu.dcache.r_tag[0][22] ),
    .A2(net693),
    .Y(_09686_),
    .B1(_09685_));
 sg13g2_xnor2_1 _16452_ (.Y(_09687_),
    .A(net365),
    .B(_09686_));
 sg13g2_mux4_1 _16453_ (.S0(net794),
    .A0(\cpu.genblk1.mmu.r_vtop_d[24][9] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[25][9] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[26][9] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[27][9] ),
    .S1(net629),
    .X(_09688_));
 sg13g2_mux4_1 _16454_ (.S0(net794),
    .A0(\cpu.genblk1.mmu.r_vtop_d[16][9] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[17][9] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[18][9] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[19][9] ),
    .S1(net629),
    .X(_09689_));
 sg13g2_mux4_1 _16455_ (.S0(net788),
    .A0(\cpu.genblk1.mmu.r_vtop_d[28][9] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[29][9] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[30][9] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[31][9] ),
    .S1(net626),
    .X(_09690_));
 sg13g2_mux4_1 _16456_ (.S0(net788),
    .A0(\cpu.genblk1.mmu.r_vtop_d[20][9] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[21][9] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[22][9] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[23][9] ),
    .S1(net626),
    .X(_09691_));
 sg13g2_mux4_1 _16457_ (.S0(net695),
    .A0(_09688_),
    .A1(_09689_),
    .A2(_09690_),
    .A3(_09691_),
    .S1(net796),
    .X(_09692_));
 sg13g2_nand2_1 _16458_ (.Y(_09693_),
    .A(net795),
    .B(_09692_));
 sg13g2_mux4_1 _16459_ (.S0(net788),
    .A0(\cpu.genblk1.mmu.r_vtop_d[8][9] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[9][9] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[10][9] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[11][9] ),
    .S1(net629),
    .X(_09694_));
 sg13g2_mux4_1 _16460_ (.S0(net794),
    .A0(\cpu.genblk1.mmu.r_vtop_d[0][9] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[1][9] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[2][9] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[3][9] ),
    .S1(net629),
    .X(_09695_));
 sg13g2_mux4_1 _16461_ (.S0(net789),
    .A0(\cpu.genblk1.mmu.r_vtop_d[12][9] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[13][9] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[14][9] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[15][9] ),
    .S1(net692),
    .X(_09696_));
 sg13g2_mux4_1 _16462_ (.S0(net789),
    .A0(\cpu.genblk1.mmu.r_vtop_d[4][9] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[5][9] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[6][9] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[7][9] ),
    .S1(net692),
    .X(_09697_));
 sg13g2_mux4_1 _16463_ (.S0(net695),
    .A0(_09694_),
    .A1(_09695_),
    .A2(_09696_),
    .A3(_09697_),
    .S1(net796),
    .X(_09698_));
 sg13g2_nand2_1 _16464_ (.Y(_09699_),
    .A(net702),
    .B(_09698_));
 sg13g2_a21oi_2 _16465_ (.B1(_08583_),
    .Y(_09700_),
    .A2(_09699_),
    .A1(_09693_));
 sg13g2_buf_1 _16466_ (.A(_09700_),
    .X(_09701_));
 sg13g2_and2_1 _16467_ (.A(\cpu.dcache.r_tag[1][21] ),
    .B(_09418_),
    .X(_09702_));
 sg13g2_a221oi_1 _16468_ (.B2(\cpu.dcache.r_tag[4][21] ),
    .C1(_09702_),
    .B1(_09552_),
    .A1(\cpu.dcache.r_tag[2][21] ),
    .Y(_09703_),
    .A2(_09413_));
 sg13g2_a22oi_1 _16469_ (.Y(_09704_),
    .B1(_09460_),
    .B2(\cpu.dcache.r_tag[5][21] ),
    .A2(_09425_),
    .A1(\cpu.dcache.r_tag[3][21] ));
 sg13g2_buf_1 _16470_ (.A(_09503_),
    .X(_09705_));
 sg13g2_a22oi_1 _16471_ (.Y(_09706_),
    .B1(net625),
    .B2(\cpu.dcache.r_tag[6][21] ),
    .A2(_09423_),
    .A1(\cpu.dcache.r_tag[7][21] ));
 sg13g2_nand4_1 _16472_ (.B(_09703_),
    .C(_09704_),
    .A(_09408_),
    .Y(_09707_),
    .D(_09706_));
 sg13g2_o21ai_1 _16473_ (.B1(_09707_),
    .Y(_09708_),
    .A1(\cpu.dcache.r_tag[0][21] ),
    .A2(_09408_));
 sg13g2_xnor2_1 _16474_ (.Y(_09709_),
    .A(net364),
    .B(_09708_));
 sg13g2_mux4_1 _16475_ (.S0(net784),
    .A0(\cpu.genblk1.mmu.r_vtop_d[24][5] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[25][5] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[26][5] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[27][5] ),
    .S1(net700),
    .X(_09710_));
 sg13g2_mux4_1 _16476_ (.S0(net784),
    .A0(\cpu.genblk1.mmu.r_vtop_d[16][5] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[17][5] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[18][5] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[19][5] ),
    .S1(net700),
    .X(_09711_));
 sg13g2_mux4_1 _16477_ (.S0(net793),
    .A0(\cpu.genblk1.mmu.r_vtop_d[28][5] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[29][5] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[30][5] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[31][5] ),
    .S1(net698),
    .X(_09712_));
 sg13g2_mux4_1 _16478_ (.S0(net793),
    .A0(\cpu.genblk1.mmu.r_vtop_d[20][5] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[21][5] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[22][5] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[23][5] ),
    .S1(net700),
    .X(_09713_));
 sg13g2_mux4_1 _16479_ (.S0(net797),
    .A0(_09710_),
    .A1(_09711_),
    .A2(_09712_),
    .A3(_09713_),
    .S1(_09482_),
    .X(_09714_));
 sg13g2_nand2_1 _16480_ (.Y(_09715_),
    .A(net795),
    .B(_09714_));
 sg13g2_mux4_1 _16481_ (.S0(_09644_),
    .A0(\cpu.genblk1.mmu.r_vtop_d[8][5] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[9][5] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[10][5] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[11][5] ),
    .S1(_09368_),
    .X(_09716_));
 sg13g2_mux4_1 _16482_ (.S0(_09644_),
    .A0(\cpu.genblk1.mmu.r_vtop_d[0][5] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[1][5] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[2][5] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[3][5] ),
    .S1(_09368_),
    .X(_09717_));
 sg13g2_mux4_1 _16483_ (.S0(_09384_),
    .A0(\cpu.genblk1.mmu.r_vtop_d[12][5] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[13][5] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[14][5] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[15][5] ),
    .S1(_09381_),
    .X(_09718_));
 sg13g2_mux4_1 _16484_ (.S0(_09384_),
    .A0(\cpu.genblk1.mmu.r_vtop_d[4][5] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[5][5] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[6][5] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[7][5] ),
    .S1(_09381_),
    .X(_09719_));
 sg13g2_mux4_1 _16485_ (.S0(net797),
    .A0(_09716_),
    .A1(_09717_),
    .A2(_09718_),
    .A3(_09719_),
    .S1(_09482_),
    .X(_09720_));
 sg13g2_nand2_1 _16486_ (.Y(_09721_),
    .A(_09363_),
    .B(_09720_));
 sg13g2_a21oi_2 _16487_ (.B1(_08582_),
    .Y(_09722_),
    .A2(_09721_),
    .A1(_09715_));
 sg13g2_buf_1 _16488_ (.A(_09722_),
    .X(_09723_));
 sg13g2_a22oi_1 _16489_ (.Y(_09724_),
    .B1(_09598_),
    .B2(\cpu.dcache.r_tag[4][17] ),
    .A2(net919),
    .A1(\cpu.dcache.r_tag[2][17] ));
 sg13g2_mux2_1 _16490_ (.A0(\cpu.dcache.r_tag[1][17] ),
    .A1(\cpu.dcache.r_tag[3][17] ),
    .S(net1069),
    .X(_09725_));
 sg13g2_a21oi_1 _16491_ (.A1(_09494_),
    .A2(_09725_),
    .Y(_09726_),
    .B1(net792));
 sg13g2_a21oi_1 _16492_ (.A1(net792),
    .A2(_09724_),
    .Y(_09727_),
    .B1(_09726_));
 sg13g2_mux2_1 _16493_ (.A0(\cpu.dcache.r_tag[5][17] ),
    .A1(\cpu.dcache.r_tag[7][17] ),
    .S(net1069),
    .X(_09728_));
 sg13g2_a22oi_1 _16494_ (.Y(_09729_),
    .B1(net785),
    .B2(\cpu.dcache.r_tag[6][17] ),
    .A2(_09728_),
    .A1(net927));
 sg13g2_nor2_1 _16495_ (.A(net920),
    .B(_09729_),
    .Y(_09730_));
 sg13g2_nor3_1 _16496_ (.A(_09467_),
    .B(_09727_),
    .C(_09730_),
    .Y(_09731_));
 sg13g2_a21oi_1 _16497_ (.A1(_00232_),
    .A2(net693),
    .Y(_09732_),
    .B1(_09731_));
 sg13g2_xnor2_1 _16498_ (.Y(_09733_),
    .A(net420),
    .B(_09732_));
 sg13g2_mux4_1 _16499_ (.S0(net697),
    .A0(\cpu.genblk1.mmu.r_vtop_d[24][11] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[25][11] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[26][11] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[27][11] ),
    .S1(net630),
    .X(_09734_));
 sg13g2_mux4_1 _16500_ (.S0(net697),
    .A0(\cpu.genblk1.mmu.r_vtop_d[16][11] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[17][11] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[18][11] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[19][11] ),
    .S1(_09369_),
    .X(_09735_));
 sg13g2_mux4_1 _16501_ (.S0(net697),
    .A0(\cpu.genblk1.mmu.r_vtop_d[28][11] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[29][11] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[30][11] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[31][11] ),
    .S1(net630),
    .X(_09736_));
 sg13g2_mux4_1 _16502_ (.S0(net697),
    .A0(\cpu.genblk1.mmu.r_vtop_d[20][11] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[21][11] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[22][11] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[23][11] ),
    .S1(net630),
    .X(_09737_));
 sg13g2_mux4_1 _16503_ (.S0(_09375_),
    .A0(_09734_),
    .A1(_09735_),
    .A2(_09736_),
    .A3(_09737_),
    .S1(net796),
    .X(_09738_));
 sg13g2_nand2_1 _16504_ (.Y(_09739_),
    .A(net795),
    .B(_09738_));
 sg13g2_mux4_1 _16505_ (.S0(net697),
    .A0(\cpu.genblk1.mmu.r_vtop_d[8][11] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[9][11] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[10][11] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[11][11] ),
    .S1(_09382_),
    .X(_09740_));
 sg13g2_mux4_1 _16506_ (.S0(net697),
    .A0(\cpu.genblk1.mmu.r_vtop_d[0][11] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[1][11] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[2][11] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[3][11] ),
    .S1(net630),
    .X(_09741_));
 sg13g2_mux4_1 _16507_ (.S0(_09385_),
    .A0(\cpu.genblk1.mmu.r_vtop_d[12][11] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[13][11] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[14][11] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[15][11] ),
    .S1(net630),
    .X(_09742_));
 sg13g2_mux4_1 _16508_ (.S0(_09385_),
    .A0(\cpu.genblk1.mmu.r_vtop_d[4][11] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[5][11] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[6][11] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[7][11] ),
    .S1(net630),
    .X(_09743_));
 sg13g2_mux4_1 _16509_ (.S0(_09391_),
    .A0(_09740_),
    .A1(_09741_),
    .A2(_09742_),
    .A3(_09743_),
    .S1(net796),
    .X(_09744_));
 sg13g2_nand2_1 _16510_ (.Y(_09745_),
    .A(net702),
    .B(_09744_));
 sg13g2_a21oi_2 _16511_ (.B1(_08583_),
    .Y(_09746_),
    .A2(_09745_),
    .A1(_09739_));
 sg13g2_a22oi_1 _16512_ (.Y(_09747_),
    .B1(_09416_),
    .B2(\cpu.dcache.r_tag[1][23] ),
    .A2(net785),
    .A1(\cpu.dcache.r_tag[2][23] ));
 sg13g2_mux2_1 _16513_ (.A0(\cpu.dcache.r_tag[4][23] ),
    .A1(\cpu.dcache.r_tag[6][23] ),
    .S(net1069),
    .X(_09748_));
 sg13g2_nand2_1 _16514_ (.Y(_09749_),
    .A(net915),
    .B(_09748_));
 sg13g2_o21ai_1 _16515_ (.B1(_09749_),
    .Y(_09750_),
    .A1(_09400_),
    .A2(_09747_));
 sg13g2_mux2_1 _16516_ (.A0(\cpu.dcache.r_tag[5][23] ),
    .A1(\cpu.dcache.r_tag[7][23] ),
    .S(_09291_),
    .X(_09751_));
 sg13g2_a22oi_1 _16517_ (.Y(_09752_),
    .B1(_09751_),
    .B2(net917),
    .A2(net919),
    .A1(\cpu.dcache.r_tag[3][23] ));
 sg13g2_nor2_1 _16518_ (.A(_09428_),
    .B(_09752_),
    .Y(_09753_));
 sg13g2_nor3_1 _16519_ (.A(_09467_),
    .B(_09750_),
    .C(_09753_),
    .Y(_09754_));
 sg13g2_a21o_1 _16520_ (.A2(_09468_),
    .A1(_00235_),
    .B1(_09754_),
    .X(_09755_));
 sg13g2_xor2_1 _16521_ (.B(_09755_),
    .A(_09746_),
    .X(_09756_));
 sg13g2_mux4_1 _16522_ (.S0(net922),
    .A0(\cpu.genblk1.mmu.r_vtop_d[16][3] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[17][3] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[18][3] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[19][3] ),
    .S1(net696),
    .X(_09757_));
 sg13g2_mux4_1 _16523_ (.S0(net922),
    .A0(\cpu.genblk1.mmu.r_vtop_d[0][3] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[1][3] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[2][3] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[3][3] ),
    .S1(net696),
    .X(_09758_));
 sg13g2_mux4_1 _16524_ (.S0(_09364_),
    .A0(\cpu.genblk1.mmu.r_vtop_d[20][3] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[21][3] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[22][3] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[23][3] ),
    .S1(_09367_),
    .X(_09759_));
 sg13g2_mux4_1 _16525_ (.S0(_09364_),
    .A0(\cpu.genblk1.mmu.r_vtop_d[4][3] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[5][3] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[6][3] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[7][3] ),
    .S1(_09367_),
    .X(_09760_));
 sg13g2_mux4_1 _16526_ (.S0(net826),
    .A0(_09757_),
    .A1(_09758_),
    .A2(_09759_),
    .A3(_09760_),
    .S1(net945),
    .X(_09761_));
 sg13g2_nand2_1 _16527_ (.Y(_09762_),
    .A(_08338_),
    .B(_09761_));
 sg13g2_mux4_1 _16528_ (.S0(net922),
    .A0(\cpu.genblk1.mmu.r_vtop_d[24][3] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[25][3] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[26][3] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[27][3] ),
    .S1(net698),
    .X(_09763_));
 sg13g2_mux4_1 _16529_ (.S0(net793),
    .A0(\cpu.genblk1.mmu.r_vtop_d[8][3] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[9][3] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[10][3] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[11][3] ),
    .S1(net698),
    .X(_09764_));
 sg13g2_mux4_1 _16530_ (.S0(net922),
    .A0(\cpu.genblk1.mmu.r_vtop_d[28][3] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[29][3] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[30][3] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[31][3] ),
    .S1(net696),
    .X(_09765_));
 sg13g2_mux4_1 _16531_ (.S0(net922),
    .A0(\cpu.genblk1.mmu.r_vtop_d[12][3] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[13][3] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[14][3] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[15][3] ),
    .S1(net696),
    .X(_09766_));
 sg13g2_mux4_1 _16532_ (.S0(_08372_),
    .A0(_09763_),
    .A1(_09764_),
    .A2(_09765_),
    .A3(_09766_),
    .S1(net945),
    .X(_09767_));
 sg13g2_o21ai_1 _16533_ (.B1(net1086),
    .Y(_09768_),
    .A1(_08339_),
    .A2(_09767_));
 sg13g2_o21ai_1 _16534_ (.B1(_09768_),
    .Y(_09769_),
    .A1(_08384_),
    .A2(_09762_));
 sg13g2_buf_1 _16535_ (.A(_09769_),
    .X(_09770_));
 sg13g2_a22oi_1 _16536_ (.Y(_09771_),
    .B1(_09425_),
    .B2(\cpu.dcache.r_tag[3][15] ),
    .A2(_09503_),
    .A1(\cpu.dcache.r_tag[6][15] ));
 sg13g2_a22oi_1 _16537_ (.Y(_09772_),
    .B1(_09418_),
    .B2(\cpu.dcache.r_tag[1][15] ),
    .A2(_09413_),
    .A1(\cpu.dcache.r_tag[2][15] ));
 sg13g2_mux2_1 _16538_ (.A0(\cpu.dcache.r_tag[5][15] ),
    .A1(\cpu.dcache.r_tag[7][15] ),
    .S(net1136),
    .X(_09773_));
 sg13g2_a22oi_1 _16539_ (.Y(_09774_),
    .B1(_09773_),
    .B2(net927),
    .A2(_09402_),
    .A1(\cpu.dcache.r_tag[4][15] ));
 sg13g2_nand2b_1 _16540_ (.Y(_09775_),
    .B(net917),
    .A_N(_09774_));
 sg13g2_and4_1 _16541_ (.A(_09407_),
    .B(_09771_),
    .C(_09772_),
    .D(_09775_),
    .X(_09776_));
 sg13g2_a21oi_1 _16542_ (.A1(_00230_),
    .A2(net693),
    .Y(_09777_),
    .B1(_09776_));
 sg13g2_xnor2_1 _16543_ (.Y(_09778_),
    .A(_09770_),
    .B(_09777_));
 sg13g2_mux4_1 _16544_ (.S0(net793),
    .A0(\cpu.genblk1.mmu.r_vtop_d[24][4] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[25][4] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[26][4] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[27][4] ),
    .S1(net698),
    .X(_09779_));
 sg13g2_mux4_1 _16545_ (.S0(net793),
    .A0(\cpu.genblk1.mmu.r_vtop_d[16][4] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[17][4] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[18][4] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[19][4] ),
    .S1(net698),
    .X(_09780_));
 sg13g2_mux4_1 _16546_ (.S0(net922),
    .A0(\cpu.genblk1.mmu.r_vtop_d[28][4] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[29][4] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[30][4] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[31][4] ),
    .S1(net696),
    .X(_09781_));
 sg13g2_mux4_1 _16547_ (.S0(net922),
    .A0(\cpu.genblk1.mmu.r_vtop_d[20][4] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[21][4] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[22][4] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[23][4] ),
    .S1(net696),
    .X(_09782_));
 sg13g2_mux4_1 _16548_ (.S0(net797),
    .A0(_09779_),
    .A1(_09780_),
    .A2(_09781_),
    .A3(_09782_),
    .S1(_08436_),
    .X(_09783_));
 sg13g2_nand2_1 _16549_ (.Y(_09784_),
    .A(net795),
    .B(_09783_));
 sg13g2_mux4_1 _16550_ (.S0(net793),
    .A0(\cpu.genblk1.mmu.r_vtop_d[8][4] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[9][4] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[10][4] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[11][4] ),
    .S1(net698),
    .X(_09785_));
 sg13g2_mux4_1 _16551_ (.S0(net793),
    .A0(\cpu.genblk1.mmu.r_vtop_d[0][4] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[1][4] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[2][4] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[3][4] ),
    .S1(net698),
    .X(_09786_));
 sg13g2_mux4_1 _16552_ (.S0(_09379_),
    .A0(\cpu.genblk1.mmu.r_vtop_d[12][4] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[13][4] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[14][4] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[15][4] ),
    .S1(_09387_),
    .X(_09787_));
 sg13g2_mux4_1 _16553_ (.S0(_09379_),
    .A0(\cpu.genblk1.mmu.r_vtop_d[4][4] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[5][4] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[6][4] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[7][4] ),
    .S1(_09387_),
    .X(_09788_));
 sg13g2_mux4_1 _16554_ (.S0(net797),
    .A0(_09785_),
    .A1(_09786_),
    .A2(_09787_),
    .A3(_09788_),
    .S1(_08436_),
    .X(_09789_));
 sg13g2_nand2_1 _16555_ (.Y(_09790_),
    .A(_08372_),
    .B(_09789_));
 sg13g2_a21oi_2 _16556_ (.B1(_08582_),
    .Y(_09791_),
    .A2(_09790_),
    .A1(_09784_));
 sg13g2_buf_1 _16557_ (.A(_09791_),
    .X(_09792_));
 sg13g2_mux2_1 _16558_ (.A0(\cpu.dcache.r_tag[5][16] ),
    .A1(\cpu.dcache.r_tag[7][16] ),
    .S(net924),
    .X(_09793_));
 sg13g2_a22oi_1 _16559_ (.Y(_09794_),
    .B1(_09793_),
    .B2(net802),
    .A2(_09547_),
    .A1(\cpu.dcache.r_tag[6][16] ));
 sg13g2_nand2b_1 _16560_ (.Y(_09795_),
    .B(_09431_),
    .A_N(_09794_));
 sg13g2_mux2_1 _16561_ (.A0(\cpu.dcache.r_tag[2][16] ),
    .A1(\cpu.dcache.r_tag[3][16] ),
    .S(_09231_),
    .X(_09796_));
 sg13g2_a22oi_1 _16562_ (.Y(_09797_),
    .B1(_09796_),
    .B2(net919),
    .A2(_09552_),
    .A1(\cpu.dcache.r_tag[4][16] ));
 sg13g2_nand2_1 _16563_ (.Y(_09798_),
    .A(\cpu.dcache.r_tag[1][16] ),
    .B(_09419_));
 sg13g2_nand2b_1 _16564_ (.Y(_09799_),
    .B(_09467_),
    .A_N(_00231_));
 sg13g2_nand4_1 _16565_ (.B(_09797_),
    .C(_09798_),
    .A(_09795_),
    .Y(_09800_),
    .D(_09799_));
 sg13g2_xnor2_1 _16566_ (.Y(_09801_),
    .A(net418),
    .B(_09800_));
 sg13g2_nand4_1 _16567_ (.B(_09756_),
    .C(_09778_),
    .A(_09733_),
    .Y(_09802_),
    .D(_09801_));
 sg13g2_nor4_1 _16568_ (.A(_09665_),
    .B(_09687_),
    .C(_09709_),
    .D(_09802_),
    .Y(_09803_));
 sg13g2_and4_1 _16569_ (.A(_09435_),
    .B(_09471_),
    .C(_09642_),
    .D(_09803_),
    .X(_09804_));
 sg13g2_mux4_1 _16570_ (.S0(_09233_),
    .A0(\cpu.dcache.r_valid[4] ),
    .A1(\cpu.dcache.r_valid[5] ),
    .A2(\cpu.dcache.r_valid[6] ),
    .A3(\cpu.dcache.r_valid[7] ),
    .S1(_09294_),
    .X(_09805_));
 sg13g2_mux4_1 _16571_ (.S0(_09233_),
    .A0(\cpu.dcache.r_valid[0] ),
    .A1(\cpu.dcache.r_valid[1] ),
    .A2(\cpu.dcache.r_valid[2] ),
    .A3(\cpu.dcache.r_valid[3] ),
    .S1(net801),
    .X(_09806_));
 sg13g2_mux2_1 _16572_ (.A0(_09805_),
    .A1(_09806_),
    .S(net920),
    .X(_09807_));
 sg13g2_mux4_1 _16573_ (.S0(net707),
    .A0(\cpu.dcache.r_dirty[4] ),
    .A1(\cpu.dcache.r_dirty[5] ),
    .A2(\cpu.dcache.r_dirty[6] ),
    .A3(\cpu.dcache.r_dirty[7] ),
    .S1(_09294_),
    .X(_09808_));
 sg13g2_mux4_1 _16574_ (.S0(net707),
    .A0(\cpu.dcache.r_dirty[0] ),
    .A1(\cpu.dcache.r_dirty[1] ),
    .A2(\cpu.dcache.r_dirty[2] ),
    .A3(\cpu.dcache.r_dirty[3] ),
    .S1(net706),
    .X(_09809_));
 sg13g2_buf_1 _16575_ (.A(net920),
    .X(_09810_));
 sg13g2_mux2_1 _16576_ (.A0(_09808_),
    .A1(_09809_),
    .S(net783),
    .X(_09811_));
 sg13g2_nand3_1 _16577_ (.B(_09807_),
    .C(_09811_),
    .A(_09211_),
    .Y(_09812_));
 sg13g2_buf_1 _16578_ (.A(_09812_),
    .X(_09813_));
 sg13g2_a21oi_1 _16579_ (.A1(_09362_),
    .A2(_09804_),
    .Y(_09814_),
    .B1(_09813_));
 sg13g2_inv_1 _16580_ (.Y(_09815_),
    .A(_09813_));
 sg13g2_and2_1 _16581_ (.A(_09807_),
    .B(_09804_),
    .X(_09816_));
 sg13g2_buf_1 _16582_ (.A(_09816_),
    .X(_09817_));
 sg13g2_nor3_1 _16583_ (.A(_09361_),
    .B(_09815_),
    .C(_09817_),
    .Y(_09818_));
 sg13g2_buf_1 _16584_ (.A(_09818_),
    .X(_09819_));
 sg13g2_or2_1 _16585_ (.X(_09820_),
    .B(_09819_),
    .A(_09814_));
 sg13g2_nor2b_1 _16586_ (.A(_08340_),
    .B_N(_09211_),
    .Y(_09821_));
 sg13g2_nand2_1 _16587_ (.Y(_09822_),
    .A(_08343_),
    .B(_09219_));
 sg13g2_nand3_1 _16588_ (.B(_09821_),
    .C(_09822_),
    .A(_09820_),
    .Y(_09823_));
 sg13g2_o21ai_1 _16589_ (.B1(_09823_),
    .Y(_09824_),
    .A1(_08346_),
    .A2(_08900_));
 sg13g2_nor2_1 _16590_ (.A(_09360_),
    .B(_09824_),
    .Y(_09825_));
 sg13g2_inv_1 _16591_ (.Y(_09826_),
    .A(_09825_));
 sg13g2_buf_2 _16592_ (.A(\cpu.qspi.r_state[7] ),
    .X(_09827_));
 sg13g2_buf_1 _16593_ (.A(\cpu.qspi.r_ind ),
    .X(_09828_));
 sg13g2_buf_1 _16594_ (.A(_00236_),
    .X(_09829_));
 sg13g2_buf_1 _16595_ (.A(\cpu.qspi.r_count[0] ),
    .X(_09830_));
 sg13g2_buf_2 _16596_ (.A(\cpu.qspi.r_count[1] ),
    .X(_09831_));
 sg13g2_buf_1 _16597_ (.A(\cpu.qspi.r_count[2] ),
    .X(_09832_));
 sg13g2_nor3_1 _16598_ (.A(_09830_),
    .B(_09831_),
    .C(_09832_),
    .Y(_09833_));
 sg13g2_nor2b_1 _16599_ (.A(\cpu.qspi.r_count[3] ),
    .B_N(_09833_),
    .Y(_09834_));
 sg13g2_buf_1 _16600_ (.A(_09834_),
    .X(_09835_));
 sg13g2_and2_1 _16601_ (.A(_09829_),
    .B(_09835_),
    .X(_09836_));
 sg13g2_buf_1 _16602_ (.A(_09836_),
    .X(_09837_));
 sg13g2_buf_2 _16603_ (.A(\cpu.qspi.r_state[2] ),
    .X(_09838_));
 sg13g2_buf_1 _16604_ (.A(\cpu.qspi.r_state[1] ),
    .X(_09839_));
 sg13g2_a221oi_1 _16605_ (.B2(_09838_),
    .C1(_09839_),
    .B1(_09837_),
    .A1(_09827_),
    .Y(_09840_),
    .A2(_09828_));
 sg13g2_a21oi_1 _16606_ (.A1(_09826_),
    .A2(_09840_),
    .Y(_00026_),
    .B1(net704));
 sg13g2_buf_2 _16607_ (.A(\cpu.qspi.r_state[16] ),
    .X(_09841_));
 sg13g2_nand2_1 _16608_ (.Y(_09842_),
    .A(_09829_),
    .B(_09835_));
 sg13g2_buf_1 _16609_ (.A(_09842_),
    .X(_09843_));
 sg13g2_and2_1 _16610_ (.A(_08346_),
    .B(_09814_),
    .X(_09844_));
 sg13g2_buf_1 _16611_ (.A(_09844_),
    .X(_09845_));
 sg13g2_buf_2 _16612_ (.A(\cpu.qspi.r_state[8] ),
    .X(_09846_));
 sg13g2_a22oi_1 _16613_ (.Y(_09847_),
    .B1(net111),
    .B2(_09846_),
    .A2(net624),
    .A1(_09841_));
 sg13g2_nor2_1 _16614_ (.A(net705),
    .B(_09847_),
    .Y(_00025_));
 sg13g2_buf_1 _16615_ (.A(_00261_),
    .X(_09848_));
 sg13g2_buf_1 _16616_ (.A(\cpu.qspi.r_state[12] ),
    .X(_09849_));
 sg13g2_buf_1 _16617_ (.A(_09849_),
    .X(_09850_));
 sg13g2_nand2_1 _16618_ (.Y(_09851_),
    .A(net1064),
    .B(net624));
 sg13g2_buf_2 _16619_ (.A(net923),
    .X(_09852_));
 sg13g2_buf_1 _16620_ (.A(_09852_),
    .X(_09853_));
 sg13g2_a21oi_1 _16621_ (.A1(_09848_),
    .A2(_09851_),
    .Y(_00023_),
    .B1(net687));
 sg13g2_buf_1 _16622_ (.A(\cpu.qspi.r_state[4] ),
    .X(_09854_));
 sg13g2_buf_1 _16623_ (.A(\cpu.qspi.r_rom_mode[1] ),
    .X(_09855_));
 sg13g2_buf_1 _16624_ (.A(\cpu.qspi.r_rom_mode[0] ),
    .X(_09856_));
 sg13g2_buf_1 _16625_ (.A(_09746_),
    .X(_09857_));
 sg13g2_nor2_1 _16626_ (.A(_08346_),
    .B(_08799_),
    .Y(_09858_));
 sg13g2_a21oi_1 _16627_ (.A1(_08346_),
    .A2(net363),
    .Y(_09859_),
    .B1(_09858_));
 sg13g2_nor2b_1 _16628_ (.A(_09856_),
    .B_N(_09859_),
    .Y(_09860_));
 sg13g2_a21oi_1 _16629_ (.A1(_09856_),
    .A2(net111),
    .Y(_09861_),
    .B1(_09860_));
 sg13g2_and2_1 _16630_ (.A(_09855_),
    .B(_09861_),
    .X(_09862_));
 sg13g2_buf_1 _16631_ (.A(_09862_),
    .X(_09863_));
 sg13g2_nor3_1 _16632_ (.A(_09856_),
    .B(_09855_),
    .C(_09859_),
    .Y(_09864_));
 sg13g2_buf_1 _16633_ (.A(_09864_),
    .X(_09865_));
 sg13g2_nor2_2 _16634_ (.A(net224),
    .B(net81),
    .Y(_09866_));
 sg13g2_and2_1 _16635_ (.A(\cpu.qspi.r_quad[2] ),
    .B(net224),
    .X(_09867_));
 sg13g2_a221oi_1 _16636_ (.B2(\cpu.qspi.r_quad[0] ),
    .C1(_09867_),
    .B1(_09866_),
    .A1(\cpu.qspi.r_quad[1] ),
    .Y(_09868_),
    .A2(net81));
 sg13g2_buf_2 _16637_ (.A(_09868_),
    .X(_09869_));
 sg13g2_and2_1 _16638_ (.A(\cpu.qspi.r_state[17] ),
    .B(_09824_),
    .X(_09870_));
 sg13g2_a22oi_1 _16639_ (.Y(_09871_),
    .B1(_09869_),
    .B2(_09870_),
    .A2(net624),
    .A1(_09854_));
 sg13g2_nor2_1 _16640_ (.A(net705),
    .B(_09871_),
    .Y(_00028_));
 sg13g2_nand2_1 _16641_ (.Y(_09872_),
    .A(_09838_),
    .B(net624));
 sg13g2_buf_2 _16642_ (.A(\cpu.qspi.r_state[14] ),
    .X(_09873_));
 sg13g2_nand2_1 _16643_ (.Y(_09874_),
    .A(_09873_),
    .B(_09837_));
 sg13g2_a21oi_1 _16644_ (.A1(_09872_),
    .A2(_09874_),
    .Y(_00027_),
    .B1(_09853_));
 sg13g2_inv_1 _16645_ (.Y(_09875_),
    .A(_09828_));
 sg13g2_buf_1 _16646_ (.A(net923),
    .X(_09876_));
 sg13g2_a21o_1 _16647_ (.A2(_09875_),
    .A1(_09827_),
    .B1(_09876_),
    .X(_00021_));
 sg13g2_buf_2 _16648_ (.A(\cpu.dec.r_op[1] ),
    .X(_09877_));
 sg13g2_nor4_1 _16649_ (.A(net173),
    .B(_08922_),
    .C(_09142_),
    .D(_09128_),
    .Y(_09878_));
 sg13g2_a21o_1 _16650_ (.A2(_09134_),
    .A1(_09877_),
    .B1(_09878_),
    .X(_00012_));
 sg13g2_buf_2 _16651_ (.A(\cpu.dec.r_op[10] ),
    .X(_09879_));
 sg13g2_nand2_1 _16652_ (.Y(_09880_),
    .A(_09067_),
    .B(_09084_));
 sg13g2_nor3_1 _16653_ (.A(net172),
    .B(_09131_),
    .C(_09880_),
    .Y(_09881_));
 sg13g2_a21o_1 _16654_ (.A2(net148),
    .A1(_09879_),
    .B1(_09881_),
    .X(_00011_));
 sg13g2_buf_1 _16655_ (.A(\cpu.dec.r_op[9] ),
    .X(_09882_));
 sg13g2_buf_1 _16656_ (.A(net1131),
    .X(_09883_));
 sg13g2_nand4_1 _16657_ (.B(net423),
    .C(net292),
    .A(net126),
    .Y(_09884_),
    .D(net170));
 sg13g2_o21ai_1 _16658_ (.B1(_09884_),
    .Y(_09885_),
    .A1(_09142_),
    .A2(_09149_));
 sg13g2_mux2_1 _16659_ (.A0(net1063),
    .A1(_09885_),
    .S(net146),
    .X(_00020_));
 sg13g2_buf_1 _16660_ (.A(\cpu.qspi.r_state[9] ),
    .X(_09886_));
 sg13g2_a21oi_1 _16661_ (.A1(_09854_),
    .A2(_09837_),
    .Y(_09887_),
    .B1(_09886_));
 sg13g2_nor2_1 _16662_ (.A(net705),
    .B(_09887_),
    .Y(_00022_));
 sg13g2_buf_1 _16663_ (.A(\cpu.qspi.r_state[5] ),
    .X(_09888_));
 sg13g2_inv_1 _16664_ (.Y(_09889_),
    .A(_09888_));
 sg13g2_nand2_1 _16665_ (.Y(_09890_),
    .A(_09873_),
    .B(net624));
 sg13g2_a21oi_1 _16666_ (.A1(_09889_),
    .A2(_09890_),
    .Y(_00024_),
    .B1(_09853_));
 sg13g2_buf_1 _16667_ (.A(\cpu.dec.r_op[8] ),
    .X(_09891_));
 sg13g2_inv_2 _16668_ (.Y(_09892_),
    .A(net1130));
 sg13g2_nand2_2 _16669_ (.Y(_09893_),
    .A(_08971_),
    .B(net293));
 sg13g2_buf_1 _16670_ (.A(_09004_),
    .X(_09894_));
 sg13g2_and2_1 _16671_ (.A(_09027_),
    .B(_09045_),
    .X(_09895_));
 sg13g2_buf_1 _16672_ (.A(_09895_),
    .X(_09896_));
 sg13g2_buf_1 _16673_ (.A(_09896_),
    .X(_09897_));
 sg13g2_nand2_1 _16674_ (.Y(_09898_),
    .A(net287),
    .B(net145));
 sg13g2_or3_1 _16675_ (.A(_08903_),
    .B(_09893_),
    .C(_09898_),
    .X(_09899_));
 sg13g2_o21ai_1 _16676_ (.B1(_09899_),
    .Y(_00019_),
    .A1(_09892_),
    .A2(_09102_));
 sg13g2_buf_1 _16677_ (.A(\cpu.uart.r_div[11] ),
    .X(_09900_));
 sg13g2_nor3_1 _16678_ (.A(\cpu.uart.r_div[0] ),
    .B(\cpu.uart.r_div[1] ),
    .C(\cpu.uart.r_div[2] ),
    .Y(_09901_));
 sg13g2_nor2b_1 _16679_ (.A(\cpu.uart.r_div[3] ),
    .B_N(_09901_),
    .Y(_09902_));
 sg13g2_nor2b_1 _16680_ (.A(\cpu.uart.r_div[4] ),
    .B_N(_09902_),
    .Y(_09903_));
 sg13g2_nor2b_1 _16681_ (.A(\cpu.uart.r_div[5] ),
    .B_N(_09903_),
    .Y(_09904_));
 sg13g2_nor2b_1 _16682_ (.A(\cpu.uart.r_div[6] ),
    .B_N(_09904_),
    .Y(_09905_));
 sg13g2_nand2b_1 _16683_ (.Y(_09906_),
    .B(_09905_),
    .A_N(\cpu.uart.r_div[7] ));
 sg13g2_nor2_1 _16684_ (.A(\cpu.uart.r_div[8] ),
    .B(_09906_),
    .Y(_09907_));
 sg13g2_nand2b_1 _16685_ (.Y(_09908_),
    .B(_09907_),
    .A_N(\cpu.uart.r_div[9] ));
 sg13g2_buf_1 _16686_ (.A(_09908_),
    .X(_09909_));
 sg13g2_nor3_1 _16687_ (.A(_09900_),
    .B(\cpu.uart.r_div[10] ),
    .C(_09909_),
    .Y(_09910_));
 sg13g2_buf_2 _16688_ (.A(_09910_),
    .X(_09911_));
 sg13g2_nor2_1 _16689_ (.A(net923),
    .B(_09911_),
    .Y(_09912_));
 sg13g2_buf_1 _16690_ (.A(_09912_),
    .X(_09913_));
 sg13g2_buf_1 _16691_ (.A(net243),
    .X(_09914_));
 sg13g2_mux2_1 _16692_ (.A0(\cpu.uart.r_div_value[0] ),
    .A1(_00263_),
    .S(_09914_),
    .X(_00079_));
 sg13g2_xnor2_1 _16693_ (.Y(_09915_),
    .A(\cpu.uart.r_div[0] ),
    .B(\cpu.uart.r_div[1] ));
 sg13g2_mux2_1 _16694_ (.A0(\cpu.uart.r_div_value[1] ),
    .A1(_09915_),
    .S(_09914_),
    .X(_00082_));
 sg13g2_o21ai_1 _16695_ (.B1(\cpu.uart.r_div[2] ),
    .Y(_09916_),
    .A1(\cpu.uart.r_div[0] ),
    .A2(\cpu.uart.r_div[1] ));
 sg13g2_nor2b_1 _16696_ (.A(_09901_),
    .B_N(_09916_),
    .Y(_09917_));
 sg13g2_nor2_1 _16697_ (.A(\cpu.uart.r_div_value[2] ),
    .B(net243),
    .Y(_09918_));
 sg13g2_a21oi_1 _16698_ (.A1(net223),
    .A2(_09917_),
    .Y(_00083_),
    .B1(_09918_));
 sg13g2_xnor2_1 _16699_ (.Y(_09919_),
    .A(\cpu.uart.r_div[3] ),
    .B(_09901_));
 sg13g2_nor2_1 _16700_ (.A(\cpu.uart.r_div_value[3] ),
    .B(net243),
    .Y(_09920_));
 sg13g2_a21oi_1 _16701_ (.A1(net223),
    .A2(_09919_),
    .Y(_00084_),
    .B1(_09920_));
 sg13g2_xnor2_1 _16702_ (.Y(_09921_),
    .A(\cpu.uart.r_div[4] ),
    .B(_09902_));
 sg13g2_nor2_1 _16703_ (.A(\cpu.uart.r_div_value[4] ),
    .B(net243),
    .Y(_09922_));
 sg13g2_a21oi_1 _16704_ (.A1(net223),
    .A2(_09921_),
    .Y(_00085_),
    .B1(_09922_));
 sg13g2_xnor2_1 _16705_ (.Y(_09923_),
    .A(\cpu.uart.r_div[5] ),
    .B(_09903_));
 sg13g2_nor2_1 _16706_ (.A(\cpu.uart.r_div_value[5] ),
    .B(net243),
    .Y(_09924_));
 sg13g2_a21oi_1 _16707_ (.A1(net223),
    .A2(_09923_),
    .Y(_00086_),
    .B1(_09924_));
 sg13g2_xnor2_1 _16708_ (.Y(_09925_),
    .A(\cpu.uart.r_div[6] ),
    .B(_09904_));
 sg13g2_nor2_1 _16709_ (.A(\cpu.uart.r_div_value[6] ),
    .B(net243),
    .Y(_09926_));
 sg13g2_a21oi_1 _16710_ (.A1(net223),
    .A2(_09925_),
    .Y(_00087_),
    .B1(_09926_));
 sg13g2_xnor2_1 _16711_ (.Y(_09927_),
    .A(\cpu.uart.r_div[7] ),
    .B(_09905_));
 sg13g2_nor2_1 _16712_ (.A(\cpu.uart.r_div_value[7] ),
    .B(net243),
    .Y(_09928_));
 sg13g2_a21oi_1 _16713_ (.A1(net223),
    .A2(_09927_),
    .Y(_00088_),
    .B1(_09928_));
 sg13g2_xor2_1 _16714_ (.B(_09906_),
    .A(\cpu.uart.r_div[8] ),
    .X(_09929_));
 sg13g2_nor2_1 _16715_ (.A(\cpu.uart.r_div_value[8] ),
    .B(net243),
    .Y(_09930_));
 sg13g2_a21oi_1 _16716_ (.A1(net223),
    .A2(_09929_),
    .Y(_00089_),
    .B1(_09930_));
 sg13g2_xnor2_1 _16717_ (.Y(_09931_),
    .A(\cpu.uart.r_div[9] ),
    .B(_09907_));
 sg13g2_nor2_1 _16718_ (.A(\cpu.uart.r_div_value[9] ),
    .B(_09913_),
    .Y(_09932_));
 sg13g2_a21oi_1 _16719_ (.A1(net223),
    .A2(_09931_),
    .Y(_00090_),
    .B1(_09932_));
 sg13g2_buf_1 _16720_ (.A(\cpu.uart.r_div_value[10] ),
    .X(_09933_));
 sg13g2_inv_1 _16721_ (.Y(_09934_),
    .A(_09933_));
 sg13g2_nand2_1 _16722_ (.Y(_09935_),
    .A(net803),
    .B(_09909_));
 sg13g2_o21ai_1 _16723_ (.B1(_09935_),
    .Y(_09936_),
    .A1(_09900_),
    .A2(_09933_));
 sg13g2_inv_1 _16724_ (.Y(_09937_),
    .A(\cpu.uart.r_div[10] ));
 sg13g2_nor3_1 _16725_ (.A(_09937_),
    .B(_09330_),
    .C(_09909_),
    .Y(_09938_));
 sg13g2_a221oi_1 _16726_ (.B2(_09937_),
    .C1(_09938_),
    .B1(_09936_),
    .A1(_09934_),
    .Y(_00080_),
    .A2(net800));
 sg13g2_nor2_1 _16727_ (.A(\cpu.uart.r_div[10] ),
    .B(_09909_),
    .Y(_09939_));
 sg13g2_nand2_1 _16728_ (.Y(_09940_),
    .A(_09900_),
    .B(net708));
 sg13g2_o21ai_1 _16729_ (.B1(\cpu.uart.r_div_value[11] ),
    .Y(_09941_),
    .A1(_09330_),
    .A2(_09911_));
 sg13g2_o21ai_1 _16730_ (.B1(_09941_),
    .Y(_00081_),
    .A1(_09939_),
    .A2(_09940_));
 sg13g2_buf_1 _16731_ (.A(_09228_),
    .X(_09942_));
 sg13g2_buf_1 _16732_ (.A(net914),
    .X(_09943_));
 sg13g2_buf_1 _16733_ (.A(_09943_),
    .X(_09944_));
 sg13g2_buf_1 _16734_ (.A(net686),
    .X(_09945_));
 sg13g2_buf_1 _16735_ (.A(_09423_),
    .X(_09946_));
 sg13g2_buf_1 _16736_ (.A(net576),
    .X(_09947_));
 sg13g2_buf_1 _16737_ (.A(\cpu.addr[5] ),
    .X(_09948_));
 sg13g2_nor3_2 _16738_ (.A(net1129),
    .B(net1139),
    .C(net1138),
    .Y(_09949_));
 sg13g2_nand2_1 _16739_ (.Y(_09950_),
    .A(_09220_),
    .B(_09949_));
 sg13g2_buf_2 _16740_ (.A(_09950_),
    .X(_09951_));
 sg13g2_nor2_1 _16741_ (.A(_09246_),
    .B(_09951_),
    .Y(_09952_));
 sg13g2_buf_1 _16742_ (.A(_09952_),
    .X(_09953_));
 sg13g2_nand3_1 _16743_ (.B(net515),
    .C(_09953_),
    .A(net623),
    .Y(_09954_));
 sg13g2_buf_1 _16744_ (.A(_09954_),
    .X(_09955_));
 sg13g2_buf_1 _16745_ (.A(\cpu.intr.r_timer_count[19] ),
    .X(_09956_));
 sg13g2_buf_1 _16746_ (.A(\cpu.intr.r_timer_count[18] ),
    .X(_09957_));
 sg13g2_buf_1 _16747_ (.A(\cpu.intr.r_timer_count[17] ),
    .X(_09958_));
 sg13g2_buf_1 _16748_ (.A(\cpu.intr.r_timer_count[16] ),
    .X(_09959_));
 sg13g2_buf_1 _16749_ (.A(\cpu.intr.r_timer_count[14] ),
    .X(_09960_));
 sg13g2_buf_1 _16750_ (.A(\cpu.intr.r_timer_count[12] ),
    .X(_09961_));
 sg13g2_buf_1 _16751_ (.A(\cpu.intr.r_timer_count[8] ),
    .X(_09962_));
 sg13g2_buf_1 _16752_ (.A(\cpu.intr.r_timer_count[4] ),
    .X(_09963_));
 sg13g2_buf_2 _16753_ (.A(\cpu.intr.r_timer_count[1] ),
    .X(_09964_));
 sg13g2_buf_2 _16754_ (.A(\cpu.intr.r_timer_count[0] ),
    .X(_09965_));
 sg13g2_buf_1 _16755_ (.A(\cpu.intr.r_timer_count[2] ),
    .X(_09966_));
 sg13g2_or4_1 _16756_ (.A(_09964_),
    .B(_09965_),
    .C(_09966_),
    .D(\cpu.intr.r_timer_count[3] ),
    .X(_09967_));
 sg13g2_buf_1 _16757_ (.A(_09967_),
    .X(_09968_));
 sg13g2_nor3_1 _16758_ (.A(_09963_),
    .B(\cpu.intr.r_timer_count[5] ),
    .C(_09968_),
    .Y(_09969_));
 sg13g2_nor2b_1 _16759_ (.A(\cpu.intr.r_timer_count[6] ),
    .B_N(_09969_),
    .Y(_09970_));
 sg13g2_nor2b_1 _16760_ (.A(\cpu.intr.r_timer_count[7] ),
    .B_N(_09970_),
    .Y(_09971_));
 sg13g2_inv_1 _16761_ (.Y(_09972_),
    .A(_09971_));
 sg13g2_nor3_1 _16762_ (.A(_09962_),
    .B(\cpu.intr.r_timer_count[9] ),
    .C(_09972_),
    .Y(_09973_));
 sg13g2_nor2b_1 _16763_ (.A(\cpu.intr.r_timer_count[10] ),
    .B_N(_09973_),
    .Y(_09974_));
 sg13g2_nand2b_1 _16764_ (.Y(_09975_),
    .B(_09974_),
    .A_N(\cpu.intr.r_timer_count[11] ));
 sg13g2_nor3_2 _16765_ (.A(_09961_),
    .B(\cpu.intr.r_timer_count[13] ),
    .C(_09975_),
    .Y(_09976_));
 sg13g2_inv_1 _16766_ (.Y(_09977_),
    .A(_09976_));
 sg13g2_nor3_2 _16767_ (.A(_09960_),
    .B(\cpu.intr.r_timer_count[15] ),
    .C(_09977_),
    .Y(_09978_));
 sg13g2_nor2b_1 _16768_ (.A(_09959_),
    .B_N(_09978_),
    .Y(_09979_));
 sg13g2_nor2b_1 _16769_ (.A(_09958_),
    .B_N(_09979_),
    .Y(_09980_));
 sg13g2_nand2b_1 _16770_ (.Y(_09981_),
    .B(_09980_),
    .A_N(_09957_));
 sg13g2_or2_1 _16771_ (.X(_09982_),
    .B(_09981_),
    .A(_09956_));
 sg13g2_buf_1 _16772_ (.A(_09982_),
    .X(_09983_));
 sg13g2_buf_1 _16773_ (.A(\cpu.intr.r_timer_count[23] ),
    .X(_09984_));
 sg13g2_buf_1 _16774_ (.A(\cpu.intr.r_timer_count[20] ),
    .X(_09985_));
 sg13g2_buf_1 _16775_ (.A(\cpu.intr.r_timer_count[21] ),
    .X(_09986_));
 sg13g2_nor3_1 _16776_ (.A(_09985_),
    .B(_09986_),
    .C(\cpu.intr.r_timer_count[22] ),
    .Y(_09987_));
 sg13g2_nor2b_1 _16777_ (.A(_09984_),
    .B_N(_09987_),
    .Y(_09988_));
 sg13g2_nand2b_1 _16778_ (.Y(_09989_),
    .B(_09988_),
    .A_N(_09983_));
 sg13g2_buf_2 _16779_ (.A(_09989_),
    .X(_09990_));
 sg13g2_nand2_1 _16780_ (.Y(_09991_),
    .A(_09955_),
    .B(_09990_));
 sg13g2_buf_2 _16781_ (.A(_09991_),
    .X(_09992_));
 sg13g2_buf_8 _16782_ (.A(_09992_),
    .X(_09993_));
 sg13g2_mux2_1 _16783_ (.A0(_00269_),
    .A1(\cpu.intr.r_timer_reload[0] ),
    .S(net66),
    .X(_00055_));
 sg13g2_buf_1 _16784_ (.A(_09992_),
    .X(_09994_));
 sg13g2_xor2_1 _16785_ (.B(_09965_),
    .A(_09964_),
    .X(_09995_));
 sg13g2_nand2_1 _16786_ (.Y(_09996_),
    .A(\cpu.intr.r_timer_reload[1] ),
    .B(net66));
 sg13g2_o21ai_1 _16787_ (.B1(_09996_),
    .Y(_00066_),
    .A1(net65),
    .A2(_09995_));
 sg13g2_nor3_1 _16788_ (.A(_09964_),
    .B(_09965_),
    .C(_09966_),
    .Y(_09997_));
 sg13g2_o21ai_1 _16789_ (.B1(_09966_),
    .Y(_09998_),
    .A1(_09964_),
    .A2(_09965_));
 sg13g2_nor2b_1 _16790_ (.A(_09997_),
    .B_N(_09998_),
    .Y(_09999_));
 sg13g2_nand2_1 _16791_ (.Y(_10000_),
    .A(\cpu.intr.r_timer_reload[2] ),
    .B(net66));
 sg13g2_o21ai_1 _16792_ (.B1(_10000_),
    .Y(_00071_),
    .A1(net65),
    .A2(_09999_));
 sg13g2_xnor2_1 _16793_ (.Y(_10001_),
    .A(\cpu.intr.r_timer_count[3] ),
    .B(_09997_));
 sg13g2_nand2_1 _16794_ (.Y(_10002_),
    .A(\cpu.intr.r_timer_reload[3] ),
    .B(_09993_));
 sg13g2_o21ai_1 _16795_ (.B1(_10002_),
    .Y(_00072_),
    .A1(net65),
    .A2(_10001_));
 sg13g2_xor2_1 _16796_ (.B(_09968_),
    .A(_09963_),
    .X(_10003_));
 sg13g2_nand2_1 _16797_ (.Y(_10004_),
    .A(\cpu.intr.r_timer_reload[4] ),
    .B(_09993_));
 sg13g2_o21ai_1 _16798_ (.B1(_10004_),
    .Y(_00073_),
    .A1(net65),
    .A2(_10003_));
 sg13g2_o21ai_1 _16799_ (.B1(\cpu.intr.r_timer_count[5] ),
    .Y(_10005_),
    .A1(_09963_),
    .A2(_09968_));
 sg13g2_nor2b_1 _16800_ (.A(_09969_),
    .B_N(_10005_),
    .Y(_10006_));
 sg13g2_buf_8 _16801_ (.A(_09992_),
    .X(_10007_));
 sg13g2_nand2_1 _16802_ (.Y(_10008_),
    .A(\cpu.intr.r_timer_reload[5] ),
    .B(_10007_));
 sg13g2_o21ai_1 _16803_ (.B1(_10008_),
    .Y(_00074_),
    .A1(net65),
    .A2(_10006_));
 sg13g2_xnor2_1 _16804_ (.Y(_10009_),
    .A(\cpu.intr.r_timer_count[6] ),
    .B(_09969_));
 sg13g2_nand2_1 _16805_ (.Y(_10010_),
    .A(\cpu.intr.r_timer_reload[6] ),
    .B(_10007_));
 sg13g2_o21ai_1 _16806_ (.B1(_10010_),
    .Y(_00075_),
    .A1(_09994_),
    .A2(_10009_));
 sg13g2_xnor2_1 _16807_ (.Y(_10011_),
    .A(\cpu.intr.r_timer_count[7] ),
    .B(_09970_));
 sg13g2_nand2_1 _16808_ (.Y(_10012_),
    .A(\cpu.intr.r_timer_reload[7] ),
    .B(net64));
 sg13g2_o21ai_1 _16809_ (.B1(_10012_),
    .Y(_00076_),
    .A1(_09994_),
    .A2(_10011_));
 sg13g2_xnor2_1 _16810_ (.Y(_10013_),
    .A(_09962_),
    .B(_09971_));
 sg13g2_nand2_1 _16811_ (.Y(_10014_),
    .A(\cpu.intr.r_timer_reload[8] ),
    .B(net64));
 sg13g2_o21ai_1 _16812_ (.B1(_10014_),
    .Y(_00077_),
    .A1(net65),
    .A2(_10013_));
 sg13g2_o21ai_1 _16813_ (.B1(\cpu.intr.r_timer_count[9] ),
    .Y(_10015_),
    .A1(_09962_),
    .A2(_09972_));
 sg13g2_nor2b_1 _16814_ (.A(_09973_),
    .B_N(_10015_),
    .Y(_10016_));
 sg13g2_nand2_1 _16815_ (.Y(_10017_),
    .A(\cpu.intr.r_timer_reload[9] ),
    .B(net64));
 sg13g2_o21ai_1 _16816_ (.B1(_10017_),
    .Y(_00078_),
    .A1(net65),
    .A2(_10016_));
 sg13g2_xnor2_1 _16817_ (.Y(_10018_),
    .A(\cpu.intr.r_timer_count[10] ),
    .B(_09973_));
 sg13g2_nand2_1 _16818_ (.Y(_10019_),
    .A(\cpu.intr.r_timer_reload[10] ),
    .B(net64));
 sg13g2_o21ai_1 _16819_ (.B1(_10019_),
    .Y(_00056_),
    .A1(net65),
    .A2(_10018_));
 sg13g2_xnor2_1 _16820_ (.Y(_10020_),
    .A(\cpu.intr.r_timer_count[11] ),
    .B(_09974_));
 sg13g2_nand2_1 _16821_ (.Y(_10021_),
    .A(\cpu.intr.r_timer_reload[11] ),
    .B(net64));
 sg13g2_o21ai_1 _16822_ (.B1(_10021_),
    .Y(_00057_),
    .A1(net66),
    .A2(_10020_));
 sg13g2_xor2_1 _16823_ (.B(_09975_),
    .A(_09961_),
    .X(_10022_));
 sg13g2_nand2_1 _16824_ (.Y(_10023_),
    .A(\cpu.intr.r_timer_reload[12] ),
    .B(net64));
 sg13g2_o21ai_1 _16825_ (.B1(_10023_),
    .Y(_00058_),
    .A1(net66),
    .A2(_10022_));
 sg13g2_o21ai_1 _16826_ (.B1(\cpu.intr.r_timer_count[13] ),
    .Y(_10024_),
    .A1(_09961_),
    .A2(_09975_));
 sg13g2_nor2b_1 _16827_ (.A(_09976_),
    .B_N(_10024_),
    .Y(_10025_));
 sg13g2_nand2_1 _16828_ (.Y(_10026_),
    .A(\cpu.intr.r_timer_reload[13] ),
    .B(net64));
 sg13g2_o21ai_1 _16829_ (.B1(_10026_),
    .Y(_00059_),
    .A1(net66),
    .A2(_10025_));
 sg13g2_xnor2_1 _16830_ (.Y(_10027_),
    .A(_09960_),
    .B(_09976_));
 sg13g2_nand2_1 _16831_ (.Y(_10028_),
    .A(\cpu.intr.r_timer_reload[14] ),
    .B(net64));
 sg13g2_o21ai_1 _16832_ (.B1(_10028_),
    .Y(_00060_),
    .A1(net66),
    .A2(_10027_));
 sg13g2_o21ai_1 _16833_ (.B1(\cpu.intr.r_timer_count[15] ),
    .Y(_10029_),
    .A1(_09960_),
    .A2(_09977_));
 sg13g2_nor2b_1 _16834_ (.A(_09978_),
    .B_N(_10029_),
    .Y(_10030_));
 sg13g2_nand2_1 _16835_ (.Y(_10031_),
    .A(\cpu.intr.r_timer_reload[15] ),
    .B(_09992_));
 sg13g2_o21ai_1 _16836_ (.B1(_10031_),
    .Y(_00061_),
    .A1(net66),
    .A2(_10030_));
 sg13g2_buf_1 _16837_ (.A(\cpu.dcache.wdata[0] ),
    .X(_10032_));
 sg13g2_buf_1 _16838_ (.A(_10032_),
    .X(_10033_));
 sg13g2_buf_1 _16839_ (.A(_10033_),
    .X(_10034_));
 sg13g2_nor4_1 _16840_ (.A(_09958_),
    .B(_09957_),
    .C(_09956_),
    .D(\cpu.intr.r_timer_reload[16] ),
    .Y(_10035_));
 sg13g2_a21oi_1 _16841_ (.A1(_09988_),
    .A2(_10035_),
    .Y(_10036_),
    .B1(_09959_));
 sg13g2_mux2_1 _16842_ (.A0(_09959_),
    .A1(_10036_),
    .S(_09978_),
    .X(_10037_));
 sg13g2_mux2_1 _16843_ (.A0(net913),
    .A1(_10037_),
    .S(_09955_),
    .X(_00062_));
 sg13g2_inv_1 _16844_ (.Y(_10038_),
    .A(_09227_));
 sg13g2_buf_1 _16845_ (.A(_10038_),
    .X(_10039_));
 sg13g2_buf_1 _16846_ (.A(_10039_),
    .X(_10040_));
 sg13g2_buf_1 _16847_ (.A(_10040_),
    .X(_10041_));
 sg13g2_buf_1 _16848_ (.A(_10041_),
    .X(_10042_));
 sg13g2_nand2_1 _16849_ (.Y(_10043_),
    .A(net706),
    .B(net689));
 sg13g2_buf_1 _16850_ (.A(_10043_),
    .X(_10044_));
 sg13g2_nor4_1 _16851_ (.A(net622),
    .B(_09246_),
    .C(net575),
    .D(_09951_),
    .Y(_10045_));
 sg13g2_buf_1 _16852_ (.A(_10045_),
    .X(_10046_));
 sg13g2_buf_1 _16853_ (.A(net125),
    .X(_10047_));
 sg13g2_xor2_1 _16854_ (.B(_09979_),
    .A(_09958_),
    .X(_10048_));
 sg13g2_o21ai_1 _16855_ (.B1(_10048_),
    .Y(_10049_),
    .A1(\cpu.intr.r_timer_reload[17] ),
    .A2(_09990_));
 sg13g2_buf_2 _16856_ (.A(\cpu.dcache.wdata[1] ),
    .X(_10050_));
 sg13g2_buf_1 _16857_ (.A(_10050_),
    .X(_10051_));
 sg13g2_nand2_1 _16858_ (.Y(_10052_),
    .A(net1061),
    .B(net125));
 sg13g2_o21ai_1 _16859_ (.B1(_10052_),
    .Y(_00063_),
    .A1(net110),
    .A2(_10049_));
 sg13g2_xor2_1 _16860_ (.B(_09980_),
    .A(_09957_),
    .X(_10053_));
 sg13g2_o21ai_1 _16861_ (.B1(_10053_),
    .Y(_10054_),
    .A1(\cpu.intr.r_timer_reload[18] ),
    .A2(_09990_));
 sg13g2_buf_1 _16862_ (.A(\cpu.dcache.wdata[2] ),
    .X(_10055_));
 sg13g2_buf_1 _16863_ (.A(_10055_),
    .X(_10056_));
 sg13g2_nand2_1 _16864_ (.Y(_10057_),
    .A(net1060),
    .B(net125));
 sg13g2_o21ai_1 _16865_ (.B1(_10057_),
    .Y(_00064_),
    .A1(net110),
    .A2(_10054_));
 sg13g2_xnor2_1 _16866_ (.Y(_10058_),
    .A(_09956_),
    .B(_09981_));
 sg13g2_o21ai_1 _16867_ (.B1(_10058_),
    .Y(_10059_),
    .A1(\cpu.intr.r_timer_reload[19] ),
    .A2(_09990_));
 sg13g2_buf_1 _16868_ (.A(\cpu.dcache.wdata[3] ),
    .X(_10060_));
 sg13g2_nand2_1 _16869_ (.Y(_10061_),
    .A(net1128),
    .B(net125));
 sg13g2_o21ai_1 _16870_ (.B1(_10061_),
    .Y(_00065_),
    .A1(_10047_),
    .A2(_10059_));
 sg13g2_inv_1 _16871_ (.Y(_10062_),
    .A(\cpu.intr.r_timer_reload[20] ));
 sg13g2_a21oi_1 _16872_ (.A1(_10062_),
    .A2(_09988_),
    .Y(_10063_),
    .B1(_09985_));
 sg13g2_nor2b_1 _16873_ (.A(_09983_),
    .B_N(_10063_),
    .Y(_10064_));
 sg13g2_a21oi_1 _16874_ (.A1(_09985_),
    .A2(_09983_),
    .Y(_10065_),
    .B1(_10064_));
 sg13g2_buf_1 _16875_ (.A(\cpu.dcache.wdata[4] ),
    .X(_10066_));
 sg13g2_buf_1 _16876_ (.A(_10066_),
    .X(_10067_));
 sg13g2_nand2_1 _16877_ (.Y(_10068_),
    .A(net1059),
    .B(net125));
 sg13g2_o21ai_1 _16878_ (.B1(_10068_),
    .Y(_00067_),
    .A1(net110),
    .A2(_10065_));
 sg13g2_o21ai_1 _16879_ (.B1(_09955_),
    .Y(_10069_),
    .A1(\cpu.intr.r_timer_reload[21] ),
    .A2(_09990_));
 sg13g2_nor2_1 _16880_ (.A(_09985_),
    .B(_09983_),
    .Y(_10070_));
 sg13g2_xnor2_1 _16881_ (.Y(_10071_),
    .A(_09986_),
    .B(_10070_));
 sg13g2_buf_1 _16882_ (.A(\cpu.dcache.wdata[5] ),
    .X(_10072_));
 sg13g2_buf_1 _16883_ (.A(_10072_),
    .X(_10073_));
 sg13g2_nand2_1 _16884_ (.Y(_10074_),
    .A(net1058),
    .B(net125));
 sg13g2_o21ai_1 _16885_ (.B1(_10074_),
    .Y(_00068_),
    .A1(_10069_),
    .A2(_10071_));
 sg13g2_o21ai_1 _16886_ (.B1(_09955_),
    .Y(_10075_),
    .A1(\cpu.intr.r_timer_reload[22] ),
    .A2(_09990_));
 sg13g2_nor3_1 _16887_ (.A(_09985_),
    .B(_09986_),
    .C(_09983_),
    .Y(_10076_));
 sg13g2_xnor2_1 _16888_ (.Y(_10077_),
    .A(\cpu.intr.r_timer_count[22] ),
    .B(_10076_));
 sg13g2_buf_1 _16889_ (.A(\cpu.dcache.wdata[6] ),
    .X(_10078_));
 sg13g2_buf_1 _16890_ (.A(_10078_),
    .X(_10079_));
 sg13g2_nand2_1 _16891_ (.Y(_10080_),
    .A(net1057),
    .B(net125));
 sg13g2_o21ai_1 _16892_ (.B1(_10080_),
    .Y(_00069_),
    .A1(_10075_),
    .A2(_10077_));
 sg13g2_buf_2 _16893_ (.A(\cpu.dcache.wdata[7] ),
    .X(_10081_));
 sg13g2_buf_1 _16894_ (.A(_10081_),
    .X(_10082_));
 sg13g2_nor2b_1 _16895_ (.A(_09984_),
    .B_N(\cpu.intr.r_timer_reload[23] ),
    .Y(_10083_));
 sg13g2_nor2b_1 _16896_ (.A(_09983_),
    .B_N(_09987_),
    .Y(_10084_));
 sg13g2_mux2_1 _16897_ (.A0(_09984_),
    .A1(_10083_),
    .S(_10084_),
    .X(_10085_));
 sg13g2_mux2_1 _16898_ (.A0(net1056),
    .A1(_10085_),
    .S(_09955_),
    .X(_00070_));
 sg13g2_buf_1 _16899_ (.A(_09552_),
    .X(_10086_));
 sg13g2_buf_1 _16900_ (.A(net621),
    .X(_10087_));
 sg13g2_nand2_1 _16901_ (.Y(_10088_),
    .A(net574),
    .B(_09953_));
 sg13g2_buf_1 _16902_ (.A(_10088_),
    .X(_10089_));
 sg13g2_buf_1 _16903_ (.A(_10089_),
    .X(_10090_));
 sg13g2_nand2_1 _16904_ (.Y(_10091_),
    .A(net926),
    .B(net915));
 sg13g2_buf_1 _16905_ (.A(_10091_),
    .X(_10092_));
 sg13g2_nor2_1 _16906_ (.A(net1073),
    .B(net684),
    .Y(_10093_));
 sg13g2_buf_1 _16907_ (.A(_10093_),
    .X(_10094_));
 sg13g2_buf_1 _16908_ (.A(_10094_),
    .X(_10095_));
 sg13g2_and2_1 _16909_ (.A(_09953_),
    .B(net514),
    .X(_10096_));
 sg13g2_buf_1 _16910_ (.A(_10096_),
    .X(_10097_));
 sg13g2_buf_1 _16911_ (.A(_10097_),
    .X(_10098_));
 sg13g2_buf_1 _16912_ (.A(net1062),
    .X(_10099_));
 sg13g2_a22oi_1 _16913_ (.Y(_10100_),
    .B1(net89),
    .B2(net911),
    .A2(_10090_),
    .A1(_00270_));
 sg13g2_inv_1 _16914_ (.Y(_00036_),
    .A(_10100_));
 sg13g2_buf_1 _16915_ (.A(_10050_),
    .X(_10101_));
 sg13g2_buf_1 _16916_ (.A(\cpu.intr.r_clock_count[0] ),
    .X(_10102_));
 sg13g2_buf_2 _16917_ (.A(\cpu.intr.r_clock_count[1] ),
    .X(_10103_));
 sg13g2_xor2_1 _16918_ (.B(_10103_),
    .A(_10102_),
    .X(_10104_));
 sg13g2_buf_1 _16919_ (.A(net90),
    .X(_10105_));
 sg13g2_a22oi_1 _16920_ (.Y(_10106_),
    .B1(_10104_),
    .B2(net80),
    .A2(net89),
    .A1(net1055));
 sg13g2_inv_1 _16921_ (.Y(_00043_),
    .A(_10106_));
 sg13g2_buf_1 _16922_ (.A(net1060),
    .X(_10107_));
 sg13g2_buf_2 _16923_ (.A(\cpu.intr.r_clock_count[2] ),
    .X(_10108_));
 sg13g2_nand2_1 _16924_ (.Y(_10109_),
    .A(_10102_),
    .B(_10103_));
 sg13g2_xnor2_1 _16925_ (.Y(_10110_),
    .A(_10108_),
    .B(_10109_));
 sg13g2_nor2_1 _16926_ (.A(_10038_),
    .B(net707),
    .Y(_10111_));
 sg13g2_buf_2 _16927_ (.A(_10111_),
    .X(_10112_));
 sg13g2_and2_1 _16928_ (.A(_09598_),
    .B(_10112_),
    .X(_10113_));
 sg13g2_buf_1 _16929_ (.A(_10113_),
    .X(_10114_));
 sg13g2_buf_1 _16930_ (.A(_10114_),
    .X(_10115_));
 sg13g2_buf_1 _16931_ (.A(net417),
    .X(_10116_));
 sg13g2_and2_1 _16932_ (.A(_09953_),
    .B(_10116_),
    .X(_10117_));
 sg13g2_buf_1 _16933_ (.A(_10117_),
    .X(_10118_));
 sg13g2_nor2_1 _16934_ (.A(_10097_),
    .B(_10118_),
    .Y(_10119_));
 sg13g2_a22oi_1 _16935_ (.Y(_10120_),
    .B1(_10110_),
    .B2(_10119_),
    .A2(net89),
    .A1(net910));
 sg13g2_inv_1 _16936_ (.Y(_00044_),
    .A(_10120_));
 sg13g2_buf_1 _16937_ (.A(net1128),
    .X(_10121_));
 sg13g2_buf_2 _16938_ (.A(\cpu.intr.r_clock_count[3] ),
    .X(_10122_));
 sg13g2_nand2_1 _16939_ (.Y(_10123_),
    .A(_10103_),
    .B(_10108_));
 sg13g2_nor2_1 _16940_ (.A(_00270_),
    .B(_10123_),
    .Y(_10124_));
 sg13g2_xor2_1 _16941_ (.B(_10124_),
    .A(_10122_),
    .X(_10125_));
 sg13g2_a22oi_1 _16942_ (.Y(_10126_),
    .B1(_10125_),
    .B2(net80),
    .A2(net89),
    .A1(net1054));
 sg13g2_inv_1 _16943_ (.Y(_00045_),
    .A(_10126_));
 sg13g2_buf_2 _16944_ (.A(\cpu.intr.r_clock_count[4] ),
    .X(_10127_));
 sg13g2_and4_1 _16945_ (.A(_10102_),
    .B(_10103_),
    .C(_10108_),
    .D(_10122_),
    .X(_10128_));
 sg13g2_buf_1 _16946_ (.A(_10128_),
    .X(_10129_));
 sg13g2_xor2_1 _16947_ (.B(_10129_),
    .A(_10127_),
    .X(_10130_));
 sg13g2_a22oi_1 _16948_ (.Y(_10131_),
    .B1(_10130_),
    .B2(net80),
    .A2(_10098_),
    .A1(net1059));
 sg13g2_inv_1 _16949_ (.Y(_00046_),
    .A(_10131_));
 sg13g2_buf_2 _16950_ (.A(\cpu.intr.r_clock_count[5] ),
    .X(_10132_));
 sg13g2_nand3_1 _16951_ (.B(_10127_),
    .C(_10124_),
    .A(_10122_),
    .Y(_10133_));
 sg13g2_xnor2_1 _16952_ (.Y(_10134_),
    .A(_10132_),
    .B(_10133_));
 sg13g2_a22oi_1 _16953_ (.Y(_10135_),
    .B1(_10134_),
    .B2(_10105_),
    .A2(net89),
    .A1(net1058));
 sg13g2_inv_1 _16954_ (.Y(_00047_),
    .A(_10135_));
 sg13g2_buf_2 _16955_ (.A(\cpu.intr.r_clock_count[6] ),
    .X(_10136_));
 sg13g2_nand3_1 _16956_ (.B(_10132_),
    .C(_10129_),
    .A(_10127_),
    .Y(_10137_));
 sg13g2_xnor2_1 _16957_ (.Y(_10138_),
    .A(_10136_),
    .B(_10137_));
 sg13g2_a22oi_1 _16958_ (.Y(_10139_),
    .B1(_10119_),
    .B2(_10138_),
    .A2(_10098_),
    .A1(net1057));
 sg13g2_inv_1 _16959_ (.Y(_00048_),
    .A(_10139_));
 sg13g2_buf_1 _16960_ (.A(_10081_),
    .X(_10140_));
 sg13g2_buf_1 _16961_ (.A(\cpu.intr.r_clock_count[7] ),
    .X(_10141_));
 sg13g2_and3_1 _16962_ (.X(_10142_),
    .A(_10122_),
    .B(_10127_),
    .C(_10124_));
 sg13g2_nand3_1 _16963_ (.B(_10136_),
    .C(_10142_),
    .A(_10132_),
    .Y(_10143_));
 sg13g2_xnor2_1 _16964_ (.Y(_10144_),
    .A(_10141_),
    .B(_10143_));
 sg13g2_a22oi_1 _16965_ (.Y(_10145_),
    .B1(_10144_),
    .B2(_10105_),
    .A2(net89),
    .A1(net1053));
 sg13g2_inv_1 _16966_ (.Y(_00049_),
    .A(_10145_));
 sg13g2_buf_2 _16967_ (.A(\cpu.dcache.wdata[8] ),
    .X(_10146_));
 sg13g2_buf_2 _16968_ (.A(\cpu.intr.r_clock_count[8] ),
    .X(_10147_));
 sg13g2_nand2_1 _16969_ (.Y(_10148_),
    .A(_10127_),
    .B(_10129_));
 sg13g2_nand3_1 _16970_ (.B(_10136_),
    .C(_10141_),
    .A(_10132_),
    .Y(_10149_));
 sg13g2_nor2_1 _16971_ (.A(_10148_),
    .B(_10149_),
    .Y(_10150_));
 sg13g2_xor2_1 _16972_ (.B(_10150_),
    .A(_10147_),
    .X(_10151_));
 sg13g2_a22oi_1 _16973_ (.Y(_10152_),
    .B1(_10151_),
    .B2(net80),
    .A2(net89),
    .A1(_10146_));
 sg13g2_inv_1 _16974_ (.Y(_00050_),
    .A(_10152_));
 sg13g2_buf_2 _16975_ (.A(\cpu.intr.r_clock_count[9] ),
    .X(_10153_));
 sg13g2_nand2_1 _16976_ (.Y(_10154_),
    .A(_10147_),
    .B(_10150_));
 sg13g2_xnor2_1 _16977_ (.Y(_10155_),
    .A(_10153_),
    .B(_10154_));
 sg13g2_a22oi_1 _16978_ (.Y(_10156_),
    .B1(_10155_),
    .B2(net80),
    .A2(net89),
    .A1(\cpu.dcache.wdata[9] ));
 sg13g2_inv_1 _16979_ (.Y(_00051_),
    .A(_10156_));
 sg13g2_buf_1 _16980_ (.A(_10097_),
    .X(_10157_));
 sg13g2_buf_1 _16981_ (.A(\cpu.intr.r_clock_count[10] ),
    .X(_10158_));
 sg13g2_nand3_1 _16982_ (.B(_10153_),
    .C(_10150_),
    .A(_10147_),
    .Y(_10159_));
 sg13g2_xnor2_1 _16983_ (.Y(_10160_),
    .A(_10158_),
    .B(_10159_));
 sg13g2_a22oi_1 _16984_ (.Y(_10161_),
    .B1(_10160_),
    .B2(net80),
    .A2(net88),
    .A1(\cpu.dcache.wdata[10] ));
 sg13g2_inv_1 _16985_ (.Y(_00037_),
    .A(_10161_));
 sg13g2_buf_2 _16986_ (.A(\cpu.dcache.wdata[11] ),
    .X(_10162_));
 sg13g2_buf_1 _16987_ (.A(\cpu.intr.r_clock_count[11] ),
    .X(_10163_));
 sg13g2_nand3_1 _16988_ (.B(_10153_),
    .C(_10158_),
    .A(_10147_),
    .Y(_10164_));
 sg13g2_nor2_1 _16989_ (.A(_10149_),
    .B(_10164_),
    .Y(_10165_));
 sg13g2_nand2_1 _16990_ (.Y(_10166_),
    .A(_10142_),
    .B(_10165_));
 sg13g2_xnor2_1 _16991_ (.Y(_10167_),
    .A(_10163_),
    .B(_10166_));
 sg13g2_a22oi_1 _16992_ (.Y(_10168_),
    .B1(_10167_),
    .B2(net80),
    .A2(net88),
    .A1(_10162_));
 sg13g2_inv_1 _16993_ (.Y(_00038_),
    .A(_10168_));
 sg13g2_buf_1 _16994_ (.A(\cpu.intr.r_clock_count[12] ),
    .X(_10169_));
 sg13g2_nand4_1 _16995_ (.B(_10163_),
    .C(_10129_),
    .A(_10127_),
    .Y(_10170_),
    .D(_10165_));
 sg13g2_xnor2_1 _16996_ (.Y(_10171_),
    .A(_10169_),
    .B(_10170_));
 sg13g2_a22oi_1 _16997_ (.Y(_10172_),
    .B1(_10171_),
    .B2(net80),
    .A2(net88),
    .A1(\cpu.dcache.wdata[12] ));
 sg13g2_inv_1 _16998_ (.Y(_00039_),
    .A(_10172_));
 sg13g2_buf_2 _16999_ (.A(\cpu.intr.r_clock_count[13] ),
    .X(_10173_));
 sg13g2_nand3_1 _17000_ (.B(_10169_),
    .C(_10165_),
    .A(_10163_),
    .Y(_10174_));
 sg13g2_buf_1 _17001_ (.A(_10174_),
    .X(_10175_));
 sg13g2_nor2_1 _17002_ (.A(_10133_),
    .B(_10175_),
    .Y(_10176_));
 sg13g2_xor2_1 _17003_ (.B(_10176_),
    .A(_10173_),
    .X(_10177_));
 sg13g2_a22oi_1 _17004_ (.Y(_10178_),
    .B1(_10177_),
    .B2(net90),
    .A2(net88),
    .A1(\cpu.dcache.wdata[13] ));
 sg13g2_inv_1 _17005_ (.Y(_00040_),
    .A(_10178_));
 sg13g2_buf_1 _17006_ (.A(\cpu.intr.r_clock_count[14] ),
    .X(_10179_));
 sg13g2_nor2_1 _17007_ (.A(_10148_),
    .B(_10175_),
    .Y(_10180_));
 sg13g2_nand2_1 _17008_ (.Y(_10181_),
    .A(_10173_),
    .B(_10180_));
 sg13g2_xnor2_1 _17009_ (.Y(_10182_),
    .A(_10179_),
    .B(_10181_));
 sg13g2_a22oi_1 _17010_ (.Y(_10183_),
    .B1(_10182_),
    .B2(net90),
    .A2(_10157_),
    .A1(\cpu.dcache.wdata[14] ));
 sg13g2_inv_1 _17011_ (.Y(_00041_),
    .A(_10183_));
 sg13g2_buf_1 _17012_ (.A(\cpu.intr.r_clock_count[15] ),
    .X(_10184_));
 sg13g2_nand3_1 _17013_ (.B(_10179_),
    .C(_10176_),
    .A(_10173_),
    .Y(_10185_));
 sg13g2_xnor2_1 _17014_ (.Y(_10186_),
    .A(_10184_),
    .B(_10185_));
 sg13g2_a22oi_1 _17015_ (.Y(_10187_),
    .B1(_10186_),
    .B2(net90),
    .A2(_10157_),
    .A1(\cpu.dcache.wdata[15] ));
 sg13g2_inv_1 _17016_ (.Y(_00042_),
    .A(_10187_));
 sg13g2_buf_1 _17017_ (.A(\cpu.ex.r_wb_valid ),
    .X(_10188_));
 sg13g2_inv_1 _17018_ (.Y(_10189_),
    .A(net1127));
 sg13g2_buf_8 _17019_ (.A(\cpu.ex.r_wb_addr[3] ),
    .X(_10190_));
 sg13g2_buf_1 _17020_ (.A(\cpu.ex.r_wb_addr[2] ),
    .X(_10191_));
 sg13g2_buf_8 _17021_ (.A(_10191_),
    .X(_10192_));
 sg13g2_nand2b_1 _17022_ (.Y(_10193_),
    .B(net1052),
    .A_N(net1126));
 sg13g2_buf_1 _17023_ (.A(_10193_),
    .X(_10194_));
 sg13g2_buf_8 _17024_ (.A(\cpu.ex.r_wb_addr[1] ),
    .X(_10195_));
 sg13g2_buf_8 _17025_ (.A(\cpu.ex.r_wb_addr[0] ),
    .X(_10196_));
 sg13g2_nand2_1 _17026_ (.Y(_10197_),
    .A(net1125),
    .B(net1124));
 sg13g2_or3_1 _17027_ (.A(_10189_),
    .B(_10194_),
    .C(_10197_),
    .X(_10198_));
 sg13g2_buf_1 _17028_ (.A(_10198_),
    .X(_10199_));
 sg13g2_buf_1 _17029_ (.A(\cpu.ex.r_set_cc ),
    .X(_10200_));
 sg13g2_nand2_2 _17030_ (.Y(_10201_),
    .A(net1127),
    .B(_10200_));
 sg13g2_nand2_1 _17031_ (.Y(_10202_),
    .A(_10199_),
    .B(_10201_));
 sg13g2_buf_2 _17032_ (.A(_10202_),
    .X(_10203_));
 sg13g2_buf_2 _17033_ (.A(\cpu.dec.r_rs2_pc ),
    .X(_10204_));
 sg13g2_inv_2 _17034_ (.Y(_10205_),
    .A(_10204_));
 sg13g2_buf_1 _17035_ (.A(_10205_),
    .X(_10206_));
 sg13g2_buf_8 _17036_ (.A(\cpu.dec.r_rs2[2] ),
    .X(_10207_));
 sg13g2_xnor2_1 _17037_ (.Y(_10208_),
    .A(_10191_),
    .B(_10207_));
 sg13g2_buf_8 _17038_ (.A(\cpu.dec.r_rs2[1] ),
    .X(_10209_));
 sg13g2_xnor2_1 _17039_ (.Y(_10210_),
    .A(net1125),
    .B(_10209_));
 sg13g2_nand2_2 _17040_ (.Y(_10211_),
    .A(_10208_),
    .B(_10210_));
 sg13g2_buf_8 _17041_ (.A(\cpu.dec.r_rs2[3] ),
    .X(_10212_));
 sg13g2_xnor2_1 _17042_ (.Y(_10213_),
    .A(net1126),
    .B(_10212_));
 sg13g2_buf_8 _17043_ (.A(\cpu.dec.r_rs2[0] ),
    .X(_10214_));
 sg13g2_xnor2_1 _17044_ (.Y(_10215_),
    .A(net1124),
    .B(_10214_));
 sg13g2_or4_1 _17045_ (.A(net1125),
    .B(net1124),
    .C(\cpu.ex.r_wb_addr[3] ),
    .D(_10191_),
    .X(_10216_));
 sg13g2_buf_1 _17046_ (.A(_10216_),
    .X(_10217_));
 sg13g2_nand4_1 _17047_ (.B(_10213_),
    .C(_10215_),
    .A(net1127),
    .Y(_10218_),
    .D(_10217_));
 sg13g2_buf_1 _17048_ (.A(_10218_),
    .X(_10219_));
 sg13g2_nor2_1 _17049_ (.A(net1123),
    .B(_10209_),
    .Y(_10220_));
 sg13g2_buf_2 _17050_ (.A(_10220_),
    .X(_10221_));
 sg13g2_buf_2 _17051_ (.A(_10212_),
    .X(_10222_));
 sg13g2_buf_8 _17052_ (.A(net1051),
    .X(_10223_));
 sg13g2_buf_8 _17053_ (.A(_10207_),
    .X(_10224_));
 sg13g2_buf_8 _17054_ (.A(_10224_),
    .X(_10225_));
 sg13g2_nor2_2 _17055_ (.A(net908),
    .B(_10225_),
    .Y(_10226_));
 sg13g2_nand2_1 _17056_ (.Y(_10227_),
    .A(_10221_),
    .B(_10226_));
 sg13g2_o21ai_1 _17057_ (.B1(_10227_),
    .Y(_10228_),
    .A1(_10211_),
    .A2(_10219_));
 sg13g2_buf_1 _17058_ (.A(_10228_),
    .X(_10229_));
 sg13g2_inv_1 _17059_ (.Y(_10230_),
    .A(net1123));
 sg13g2_buf_1 _17060_ (.A(_10230_),
    .X(_10231_));
 sg13g2_buf_1 _17061_ (.A(net906),
    .X(_10232_));
 sg13g2_inv_1 _17062_ (.Y(_10233_),
    .A(net908));
 sg13g2_buf_1 _17063_ (.A(_10233_),
    .X(_10234_));
 sg13g2_buf_8 _17064_ (.A(_10209_),
    .X(_10235_));
 sg13g2_and2_1 _17065_ (.A(net1049),
    .B(net907),
    .X(_10236_));
 sg13g2_buf_2 _17066_ (.A(_10236_),
    .X(_10237_));
 sg13g2_nor2_1 _17067_ (.A(net1049),
    .B(net907),
    .Y(_10238_));
 sg13g2_buf_2 _17068_ (.A(_10238_),
    .X(_10239_));
 sg13g2_a22oi_1 _17069_ (.Y(_10240_),
    .B1(_10239_),
    .B2(\cpu.ex.r_8[13] ),
    .A2(_10237_),
    .A1(\cpu.ex.r_14[13] ));
 sg13g2_buf_2 _17070_ (.A(net1050),
    .X(_10241_));
 sg13g2_buf_8 _17071_ (.A(net905),
    .X(_10242_));
 sg13g2_buf_8 _17072_ (.A(net778),
    .X(_10243_));
 sg13g2_buf_8 _17073_ (.A(net682),
    .X(_10244_));
 sg13g2_buf_1 _17074_ (.A(net620),
    .X(_10245_));
 sg13g2_nor2b_1 _17075_ (.A(_10209_),
    .B_N(_10212_),
    .Y(_10246_));
 sg13g2_buf_2 _17076_ (.A(_10246_),
    .X(_10247_));
 sg13g2_buf_1 _17077_ (.A(_10247_),
    .X(_10248_));
 sg13g2_nand3_1 _17078_ (.B(net571),
    .C(net777),
    .A(\cpu.ex.r_12[13] ),
    .Y(_10249_));
 sg13g2_o21ai_1 _17079_ (.B1(_10249_),
    .Y(_10250_),
    .A1(net683),
    .A2(_10240_));
 sg13g2_buf_8 _17080_ (.A(net1049),
    .X(_10251_));
 sg13g2_buf_1 _17081_ (.A(net904),
    .X(_10252_));
 sg13g2_buf_1 _17082_ (.A(_10252_),
    .X(_10253_));
 sg13g2_and2_1 _17083_ (.A(net908),
    .B(net907),
    .X(_10254_));
 sg13g2_buf_2 _17084_ (.A(_10254_),
    .X(_10255_));
 sg13g2_inv_1 _17085_ (.Y(_10256_),
    .A(_00255_));
 sg13g2_a22oi_1 _17086_ (.Y(_10257_),
    .B1(_10255_),
    .B2(_10256_),
    .A2(_10226_),
    .A1(\cpu.ex.r_epc[13] ));
 sg13g2_nor2b_1 _17087_ (.A(_10207_),
    .B_N(_10222_),
    .Y(_10258_));
 sg13g2_buf_2 _17088_ (.A(_10258_),
    .X(_10259_));
 sg13g2_buf_8 _17089_ (.A(_10259_),
    .X(_10260_));
 sg13g2_nor2b_1 _17090_ (.A(net1051),
    .B_N(net1050),
    .Y(_10261_));
 sg13g2_buf_2 _17091_ (.A(_10261_),
    .X(_10262_));
 sg13g2_buf_2 _17092_ (.A(\cpu.ex.r_mult[29] ),
    .X(_10263_));
 sg13g2_a22oi_1 _17093_ (.Y(_10264_),
    .B1(_10262_),
    .B2(_10263_),
    .A2(net680),
    .A1(\cpu.ex.r_11[13] ));
 sg13g2_nand3_1 _17094_ (.B(_10257_),
    .C(_10264_),
    .A(net681),
    .Y(_10265_));
 sg13g2_buf_1 _17095_ (.A(\cpu.ex.mmu_read[13] ),
    .X(_10266_));
 sg13g2_a22oi_1 _17096_ (.Y(_10267_),
    .B1(_10262_),
    .B2(_10266_),
    .A2(net680),
    .A1(\cpu.ex.r_9[13] ));
 sg13g2_a21oi_1 _17097_ (.A1(\cpu.ex.r_lr[13] ),
    .A2(_10226_),
    .Y(_10268_),
    .B1(net681));
 sg13g2_a21oi_1 _17098_ (.A1(_10267_),
    .A2(_10268_),
    .Y(_10269_),
    .B1(net779));
 sg13g2_nor2b_1 _17099_ (.A(net1123),
    .B_N(_10209_),
    .Y(_10270_));
 sg13g2_buf_1 _17100_ (.A(_10270_),
    .X(_10271_));
 sg13g2_buf_1 _17101_ (.A(_10271_),
    .X(_10272_));
 sg13g2_inv_1 _17102_ (.Y(_10273_),
    .A(net775));
 sg13g2_mux2_1 _17103_ (.A0(\cpu.ex.r_sp[13] ),
    .A1(\cpu.ex.r_stmp[13] ),
    .S(net620),
    .X(_10274_));
 sg13g2_a22oi_1 _17104_ (.Y(_10275_),
    .B1(_10274_),
    .B2(net683),
    .A2(net680),
    .A1(\cpu.ex.r_10[13] ));
 sg13g2_buf_8 _17105_ (.A(net1123),
    .X(_10276_));
 sg13g2_buf_8 _17106_ (.A(_10276_),
    .X(_10277_));
 sg13g2_buf_8 _17107_ (.A(net903),
    .X(_10278_));
 sg13g2_buf_8 _17108_ (.A(net774),
    .X(_10279_));
 sg13g2_buf_8 _17109_ (.A(net679),
    .X(_10280_));
 sg13g2_buf_1 _17110_ (.A(net619),
    .X(_10281_));
 sg13g2_nand4_1 _17111_ (.B(net570),
    .C(net571),
    .A(\cpu.ex.r_13[13] ),
    .Y(_10282_),
    .D(net777));
 sg13g2_o21ai_1 _17112_ (.B1(_10282_),
    .Y(_10283_),
    .A1(_10273_),
    .A2(_10275_));
 sg13g2_a221oi_1 _17113_ (.B2(_10269_),
    .C1(_10283_),
    .B1(_10265_),
    .A1(net779),
    .Y(_10284_),
    .A2(_10250_));
 sg13g2_nor2_1 _17114_ (.A(_10211_),
    .B(_10219_),
    .Y(_10285_));
 sg13g2_buf_1 _17115_ (.A(_10285_),
    .X(_10286_));
 sg13g2_nand2_1 _17116_ (.Y(_10287_),
    .A(net577),
    .B(net569));
 sg13g2_o21ai_1 _17117_ (.B1(_10287_),
    .Y(_10288_),
    .A1(net572),
    .A2(_10284_));
 sg13g2_buf_1 _17118_ (.A(\cpu.dec.needs_rs2 ),
    .X(_10289_));
 sg13g2_buf_1 _17119_ (.A(_10289_),
    .X(_10290_));
 sg13g2_buf_1 _17120_ (.A(net1047),
    .X(_10291_));
 sg13g2_mux2_1 _17121_ (.A0(\cpu.dec.imm[13] ),
    .A1(_10288_),
    .S(_10291_),
    .X(_10292_));
 sg13g2_nor2_1 _17122_ (.A(net909),
    .B(_00186_),
    .Y(_10293_));
 sg13g2_a21o_1 _17123_ (.A2(_10292_),
    .A1(net909),
    .B1(_10293_),
    .X(_10294_));
 sg13g2_buf_1 _17124_ (.A(_10294_),
    .X(_10295_));
 sg13g2_buf_1 _17125_ (.A(_00273_),
    .X(_10296_));
 sg13g2_buf_1 _17126_ (.A(_10204_),
    .X(_10297_));
 sg13g2_buf_1 _17127_ (.A(_10297_),
    .X(_10298_));
 sg13g2_nand2b_1 _17128_ (.Y(_10299_),
    .B(net901),
    .A_N(_10296_));
 sg13g2_buf_2 _17129_ (.A(_10299_),
    .X(_10300_));
 sg13g2_inv_2 _17130_ (.Y(_10301_),
    .A(_10289_));
 sg13g2_inv_1 _17131_ (.Y(_10302_),
    .A(\cpu.dec.imm[12] ));
 sg13g2_nand2_1 _17132_ (.Y(_10303_),
    .A(_10301_),
    .B(_10302_));
 sg13g2_nand2_1 _17133_ (.Y(_10304_),
    .A(net1051),
    .B(_10224_));
 sg13g2_nor2_2 _17134_ (.A(net1049),
    .B(_10304_),
    .Y(_10305_));
 sg13g2_buf_8 _17135_ (.A(net908),
    .X(_10306_));
 sg13g2_buf_1 _17136_ (.A(net773),
    .X(_10307_));
 sg13g2_buf_8 _17137_ (.A(net678),
    .X(_10308_));
 sg13g2_mux2_1 _17138_ (.A0(\cpu.ex.r_epc[12] ),
    .A1(\cpu.ex.r_11[12] ),
    .S(net618),
    .X(_10309_));
 sg13g2_nor2b_1 _17139_ (.A(net907),
    .B_N(net1049),
    .Y(_10310_));
 sg13g2_buf_2 _17140_ (.A(_10310_),
    .X(_10311_));
 sg13g2_a22oi_1 _17141_ (.Y(_10312_),
    .B1(_10309_),
    .B2(_10311_),
    .A2(_10305_),
    .A1(\cpu.ex.r_13[12] ));
 sg13g2_buf_1 _17142_ (.A(\cpu.ex.mmu_read[12] ),
    .X(_10313_));
 sg13g2_mux2_1 _17143_ (.A0(\cpu.ex.r_lr[12] ),
    .A1(_10313_),
    .S(net620),
    .X(_10314_));
 sg13g2_a22oi_1 _17144_ (.Y(_10315_),
    .B1(_10314_),
    .B2(net683),
    .A2(net680),
    .A1(\cpu.ex.r_9[12] ));
 sg13g2_or2_1 _17145_ (.X(_10316_),
    .B(_10315_),
    .A(net681));
 sg13g2_a21oi_1 _17146_ (.A1(_10312_),
    .A2(_10316_),
    .Y(_10317_),
    .B1(net779));
 sg13g2_nor2b_1 _17147_ (.A(_00254_),
    .B_N(net619),
    .Y(_10318_));
 sg13g2_nor2b_1 _17148_ (.A(net619),
    .B_N(\cpu.ex.r_8[12] ),
    .Y(_10319_));
 sg13g2_a22oi_1 _17149_ (.Y(_10320_),
    .B1(_10319_),
    .B2(_10239_),
    .A2(_10318_),
    .A1(_10237_));
 sg13g2_nand2b_1 _17150_ (.Y(_10321_),
    .B(net618),
    .A_N(_10320_));
 sg13g2_buf_2 _17151_ (.A(\cpu.ex.r_mult[28] ),
    .X(_10322_));
 sg13g2_inv_1 _17152_ (.Y(_10323_),
    .A(_10322_));
 sg13g2_nand2b_1 _17153_ (.Y(_10324_),
    .B(_10235_),
    .A_N(_10222_));
 sg13g2_buf_2 _17154_ (.A(_10324_),
    .X(_10325_));
 sg13g2_nor3_1 _17155_ (.A(_10323_),
    .B(net779),
    .C(_10325_),
    .Y(_10326_));
 sg13g2_and3_1 _17156_ (.X(_10327_),
    .A(\cpu.ex.r_12[12] ),
    .B(net779),
    .C(net777));
 sg13g2_o21ai_1 _17157_ (.B1(net571),
    .Y(_10328_),
    .A1(_10326_),
    .A2(_10327_));
 sg13g2_buf_1 _17158_ (.A(\cpu.ex.r_sp[12] ),
    .X(_10329_));
 sg13g2_mux4_1 _17159_ (.S0(net620),
    .A0(_10329_),
    .A1(\cpu.ex.r_stmp[12] ),
    .A2(\cpu.ex.r_10[12] ),
    .A3(\cpu.ex.r_14[12] ),
    .S1(net618),
    .X(_10330_));
 sg13g2_nand2_1 _17160_ (.Y(_10331_),
    .A(net775),
    .B(_10330_));
 sg13g2_nand3_1 _17161_ (.B(_10328_),
    .C(_10331_),
    .A(_10321_),
    .Y(_10332_));
 sg13g2_and2_1 _17162_ (.A(_10208_),
    .B(_10210_),
    .X(_10333_));
 sg13g2_buf_1 _17163_ (.A(_10333_),
    .X(_10334_));
 sg13g2_and4_1 _17164_ (.A(net1127),
    .B(_10213_),
    .C(_10215_),
    .D(_10217_),
    .X(_10335_));
 sg13g2_buf_1 _17165_ (.A(_10335_),
    .X(_10336_));
 sg13g2_a22oi_1 _17166_ (.Y(_10337_),
    .B1(_10221_),
    .B2(_10226_),
    .A2(_10336_),
    .A1(_10334_));
 sg13g2_buf_1 _17167_ (.A(_10337_),
    .X(_10338_));
 sg13g2_buf_1 _17168_ (.A(_10338_),
    .X(_10339_));
 sg13g2_o21ai_1 _17169_ (.B1(net513),
    .Y(_10340_),
    .A1(_10317_),
    .A2(_10332_));
 sg13g2_buf_1 _17170_ (.A(net701),
    .X(_10341_));
 sg13g2_buf_1 _17171_ (.A(net569),
    .X(_10342_));
 sg13g2_nand2_1 _17172_ (.Y(_10343_),
    .A(net617),
    .B(_10342_));
 sg13g2_nand3_1 _17173_ (.B(_10340_),
    .C(_10343_),
    .A(_10291_),
    .Y(_10344_));
 sg13g2_nand3_1 _17174_ (.B(_10303_),
    .C(_10344_),
    .A(net909),
    .Y(_10345_));
 sg13g2_buf_2 _17175_ (.A(_10345_),
    .X(_10346_));
 sg13g2_nand2_1 _17176_ (.Y(_10347_),
    .A(_10300_),
    .B(_10346_));
 sg13g2_buf_1 _17177_ (.A(_10347_),
    .X(_10348_));
 sg13g2_nor2_1 _17178_ (.A(net222),
    .B(_10348_),
    .Y(_10349_));
 sg13g2_inv_1 _17179_ (.Y(_10350_),
    .A(_10207_));
 sg13g2_buf_1 _17180_ (.A(_10350_),
    .X(_10351_));
 sg13g2_buf_1 _17181_ (.A(net900),
    .X(_10352_));
 sg13g2_nor2b_1 _17182_ (.A(net1048),
    .B_N(net908),
    .Y(_10353_));
 sg13g2_buf_2 _17183_ (.A(_10353_),
    .X(_10354_));
 sg13g2_nor2b_1 _17184_ (.A(net908),
    .B_N(net1048),
    .Y(_10355_));
 sg13g2_buf_1 _17185_ (.A(_10355_),
    .X(_10356_));
 sg13g2_and3_1 _17186_ (.X(_10357_),
    .A(\cpu.ex.r_9[11] ),
    .B(net619),
    .C(net678));
 sg13g2_a221oi_1 _17187_ (.B2(\cpu.ex.r_lr[11] ),
    .C1(_10357_),
    .B1(_10356_),
    .A1(\cpu.ex.r_8[11] ),
    .Y(_10358_),
    .A2(_10354_));
 sg13g2_buf_1 _17188_ (.A(\cpu.ex.r_sp[11] ),
    .X(_10359_));
 sg13g2_nor2b_1 _17189_ (.A(_10212_),
    .B_N(_10209_),
    .Y(_10360_));
 sg13g2_buf_1 _17190_ (.A(_10360_),
    .X(_10361_));
 sg13g2_buf_1 _17191_ (.A(_10361_),
    .X(_10362_));
 sg13g2_nand3_1 _17192_ (.B(_10232_),
    .C(net771),
    .A(_10359_),
    .Y(_10363_));
 sg13g2_o21ai_1 _17193_ (.B1(_10363_),
    .Y(_10364_),
    .A1(net776),
    .A2(_10358_));
 sg13g2_mux2_1 _17194_ (.A0(\cpu.ex.r_10[11] ),
    .A1(\cpu.ex.r_11[11] ),
    .S(net619),
    .X(_10365_));
 sg13g2_mux2_1 _17195_ (.A0(\cpu.ex.r_12[11] ),
    .A1(\cpu.ex.r_13[11] ),
    .S(net619),
    .X(_10366_));
 sg13g2_nor2b_1 _17196_ (.A(net1049),
    .B_N(_10225_),
    .Y(_10367_));
 sg13g2_buf_2 _17197_ (.A(_10367_),
    .X(_10368_));
 sg13g2_a22oi_1 _17198_ (.Y(_10369_),
    .B1(_10366_),
    .B2(_10368_),
    .A2(_10365_),
    .A1(_10311_));
 sg13g2_inv_1 _17199_ (.Y(_10370_),
    .A(_10369_));
 sg13g2_nand2_1 _17200_ (.Y(_10371_),
    .A(net619),
    .B(net776));
 sg13g2_inv_1 _17201_ (.Y(_10372_),
    .A(_00253_));
 sg13g2_mux2_1 _17202_ (.A0(\cpu.ex.r_epc[11] ),
    .A1(\cpu.ex.r_mult[27] ),
    .S(net682),
    .X(_10373_));
 sg13g2_a22oi_1 _17203_ (.Y(_10374_),
    .B1(_10373_),
    .B2(net683),
    .A2(_10255_),
    .A1(_10372_));
 sg13g2_mux2_1 _17204_ (.A0(\cpu.ex.r_stmp[11] ),
    .A1(\cpu.ex.r_14[11] ),
    .S(net618),
    .X(_10375_));
 sg13g2_nand3_1 _17205_ (.B(net775),
    .C(_10375_),
    .A(net571),
    .Y(_10376_));
 sg13g2_o21ai_1 _17206_ (.B1(_10376_),
    .Y(_10377_),
    .A1(_10371_),
    .A2(_10374_));
 sg13g2_a221oi_1 _17207_ (.B2(_10308_),
    .C1(_10377_),
    .B1(_10370_),
    .A1(_10352_),
    .Y(_10378_),
    .A2(_10364_));
 sg13g2_buf_1 _17208_ (.A(\cpu.addr[11] ),
    .X(_10379_));
 sg13g2_nand2_1 _17209_ (.Y(_10380_),
    .A(net1122),
    .B(net569));
 sg13g2_o21ai_1 _17210_ (.B1(_10380_),
    .Y(_10381_),
    .A1(net572),
    .A2(_10378_));
 sg13g2_inv_1 _17211_ (.Y(_10382_),
    .A(\cpu.dec.imm[11] ));
 sg13g2_nor2_1 _17212_ (.A(net902),
    .B(_10382_),
    .Y(_10383_));
 sg13g2_a21oi_1 _17213_ (.A1(net902),
    .A2(_10381_),
    .Y(_10384_),
    .B1(_10383_));
 sg13g2_inv_2 _17214_ (.Y(_10385_),
    .A(_00274_));
 sg13g2_nand2_1 _17215_ (.Y(_10386_),
    .A(net901),
    .B(_10385_));
 sg13g2_o21ai_1 _17216_ (.B1(_10386_),
    .Y(_10387_),
    .A1(net901),
    .A2(_10384_));
 sg13g2_buf_2 _17217_ (.A(_10387_),
    .X(_10388_));
 sg13g2_inv_2 _17218_ (.Y(_10389_),
    .A(_00275_));
 sg13g2_nand2_1 _17219_ (.Y(_10390_),
    .A(_10298_),
    .B(_10389_));
 sg13g2_nor2_1 _17220_ (.A(net902),
    .B(\cpu.dec.imm[10] ),
    .Y(_10391_));
 sg13g2_buf_2 _17221_ (.A(\cpu.addr[10] ),
    .X(_10392_));
 sg13g2_nand3_1 _17222_ (.B(net570),
    .C(net771),
    .A(\cpu.ex.r_epc[10] ),
    .Y(_10393_));
 sg13g2_nand3_1 _17223_ (.B(net779),
    .C(net777),
    .A(\cpu.ex.r_8[10] ),
    .Y(_10394_));
 sg13g2_a21o_1 _17224_ (.A2(_10394_),
    .A1(_10393_),
    .B1(_10245_),
    .X(_10395_));
 sg13g2_buf_1 _17225_ (.A(net1123),
    .X(_10396_));
 sg13g2_and2_1 _17226_ (.A(net1045),
    .B(net908),
    .X(_10397_));
 sg13g2_buf_2 _17227_ (.A(_10397_),
    .X(_10398_));
 sg13g2_inv_1 _17228_ (.Y(_10399_),
    .A(_00252_));
 sg13g2_inv_2 _17229_ (.Y(_10400_),
    .A(net904));
 sg13g2_mux4_1 _17230_ (.S0(_10400_),
    .A0(_10399_),
    .A1(\cpu.ex.r_13[10] ),
    .A2(\cpu.ex.r_11[10] ),
    .A3(\cpu.ex.r_9[10] ),
    .S1(net772),
    .X(_10401_));
 sg13g2_nand2_1 _17231_ (.Y(_10402_),
    .A(_10398_),
    .B(_10401_));
 sg13g2_buf_1 _17232_ (.A(\cpu.ex.r_sp[10] ),
    .X(_10403_));
 sg13g2_mux2_1 _17233_ (.A0(_10403_),
    .A1(\cpu.ex.r_stmp[10] ),
    .S(net620),
    .X(_10404_));
 sg13g2_a22oi_1 _17234_ (.Y(_10405_),
    .B1(_10404_),
    .B2(net683),
    .A2(_10255_),
    .A1(\cpu.ex.r_14[10] ));
 sg13g2_nand2b_1 _17235_ (.Y(_10406_),
    .B(net775),
    .A_N(_10405_));
 sg13g2_inv_1 _17236_ (.Y(_10407_),
    .A(\cpu.ex.r_lr[10] ));
 sg13g2_or2_1 _17237_ (.X(_10408_),
    .B(_10241_),
    .A(net904));
 sg13g2_buf_1 _17238_ (.A(_10408_),
    .X(_10409_));
 sg13g2_buf_1 _17239_ (.A(\cpu.ex.r_mult[26] ),
    .X(_10410_));
 sg13g2_nand3_1 _17240_ (.B(net776),
    .C(net620),
    .A(_10410_),
    .Y(_10411_));
 sg13g2_o21ai_1 _17241_ (.B1(_10411_),
    .Y(_10412_),
    .A1(_10407_),
    .A2(_10409_));
 sg13g2_inv_1 _17242_ (.Y(_10413_),
    .A(\cpu.ex.r_10[10] ));
 sg13g2_nand2b_1 _17243_ (.Y(_10414_),
    .B(net904),
    .A_N(net778));
 sg13g2_nand3b_1 _17244_ (.B(_10244_),
    .C(\cpu.ex.r_12[10] ),
    .Y(_10415_),
    .A_N(net776));
 sg13g2_o21ai_1 _17245_ (.B1(_10415_),
    .Y(_10416_),
    .A1(_10413_),
    .A2(_10414_));
 sg13g2_a22oi_1 _17246_ (.Y(_10417_),
    .B1(_10416_),
    .B2(_10354_),
    .A2(_10412_),
    .A1(_10356_));
 sg13g2_nand4_1 _17247_ (.B(_10402_),
    .C(_10406_),
    .A(_10395_),
    .Y(_10418_),
    .D(_10417_));
 sg13g2_a221oi_1 _17248_ (.B2(_10418_),
    .C1(_10301_),
    .B1(net513),
    .A1(_10392_),
    .Y(_10419_),
    .A2(net512));
 sg13g2_or3_1 _17249_ (.A(net901),
    .B(_10391_),
    .C(_10419_),
    .X(_10420_));
 sg13g2_nand2_1 _17250_ (.Y(_10421_),
    .A(_10390_),
    .B(_10420_));
 sg13g2_buf_1 _17251_ (.A(_10421_),
    .X(_10422_));
 sg13g2_nor2_1 _17252_ (.A(_10388_),
    .B(net221),
    .Y(_10423_));
 sg13g2_buf_1 _17253_ (.A(net909),
    .X(_10424_));
 sg13g2_nor2_1 _17254_ (.A(net906),
    .B(net682),
    .Y(_10425_));
 sg13g2_nor2_1 _17255_ (.A(net570),
    .B(net772),
    .Y(_10426_));
 sg13g2_a22oi_1 _17256_ (.Y(_10427_),
    .B1(_10426_),
    .B2(\cpu.ex.r_stmp[15] ),
    .A2(_10425_),
    .A1(\cpu.ex.r_epc[15] ));
 sg13g2_and2_1 _17257_ (.A(net1048),
    .B(net1049),
    .X(_10428_));
 sg13g2_a22oi_1 _17258_ (.Y(_10429_),
    .B1(_10428_),
    .B2(\cpu.ex.r_15[15] ),
    .A2(_10221_),
    .A1(\cpu.ex.r_12[15] ));
 sg13g2_nand2b_1 _17259_ (.Y(_10430_),
    .B(_10255_),
    .A_N(_10429_));
 sg13g2_o21ai_1 _17260_ (.B1(_10430_),
    .Y(_10431_),
    .A1(_10325_),
    .A2(_10427_));
 sg13g2_nor2b_1 _17261_ (.A(_10252_),
    .B_N(net679),
    .Y(_10432_));
 sg13g2_mux2_1 _17262_ (.A0(\cpu.ex.r_lr[15] ),
    .A1(\cpu.ex.r_9[15] ),
    .S(net618),
    .X(_10433_));
 sg13g2_nand2_1 _17263_ (.Y(_10434_),
    .A(_10432_),
    .B(_10433_));
 sg13g2_nand3_1 _17264_ (.B(net618),
    .C(net775),
    .A(\cpu.ex.r_10[15] ),
    .Y(_10435_));
 sg13g2_a21oi_1 _17265_ (.A1(_10434_),
    .A2(_10435_),
    .Y(_10436_),
    .B1(net571));
 sg13g2_a221oi_1 _17266_ (.B2(\cpu.ex.r_8[15] ),
    .C1(net570),
    .B1(_10239_),
    .A1(\cpu.ex.r_14[15] ),
    .Y(_10437_),
    .A2(_10237_));
 sg13g2_a221oi_1 _17267_ (.B2(\cpu.ex.r_13[15] ),
    .C1(net779),
    .B1(_10368_),
    .A1(\cpu.ex.r_11[15] ),
    .Y(_10438_),
    .A2(_10311_));
 sg13g2_nor3_1 _17268_ (.A(net683),
    .B(_10437_),
    .C(_10438_),
    .Y(_10439_));
 sg13g2_buf_1 _17269_ (.A(\cpu.ex.r_sp[15] ),
    .X(_10440_));
 sg13g2_nor2_1 _17270_ (.A(net570),
    .B(_10414_),
    .Y(_10441_));
 sg13g2_nor2_1 _17271_ (.A(net779),
    .B(net772),
    .Y(_10442_));
 sg13g2_buf_1 _17272_ (.A(\cpu.ex.mmu_read[15] ),
    .X(_10443_));
 sg13g2_inv_1 _17273_ (.Y(_10444_),
    .A(_10443_));
 sg13g2_nand2_1 _17274_ (.Y(_10445_),
    .A(\cpu.ex.r_mult[31] ),
    .B(_10253_));
 sg13g2_o21ai_1 _17275_ (.B1(_10445_),
    .Y(_10446_),
    .A1(net1044),
    .A2(_10253_));
 sg13g2_a22oi_1 _17276_ (.Y(_10447_),
    .B1(_10442_),
    .B2(_10446_),
    .A2(_10441_),
    .A1(_10440_));
 sg13g2_nor2_1 _17277_ (.A(net618),
    .B(_10447_),
    .Y(_10448_));
 sg13g2_or4_1 _17278_ (.A(_10431_),
    .B(_10436_),
    .C(_10439_),
    .D(_10448_),
    .X(_10449_));
 sg13g2_a22oi_1 _17279_ (.Y(_10450_),
    .B1(net513),
    .B2(_10449_),
    .A2(_10342_),
    .A1(net1086));
 sg13g2_nor2_1 _17280_ (.A(net902),
    .B(\cpu.dec.imm[15] ),
    .Y(_10451_));
 sg13g2_a21oi_1 _17281_ (.A1(net902),
    .A2(_10450_),
    .Y(_10452_),
    .B1(_10451_));
 sg13g2_nor2_1 _17282_ (.A(_00184_),
    .B(net770),
    .Y(_10453_));
 sg13g2_a21o_1 _17283_ (.A2(_10452_),
    .A1(net770),
    .B1(_10453_),
    .X(_10454_));
 sg13g2_buf_1 _17284_ (.A(_10454_),
    .X(_10455_));
 sg13g2_buf_1 _17285_ (.A(\cpu.ex.r_sp[14] ),
    .X(_10456_));
 sg13g2_nor3_1 _17286_ (.A(_10276_),
    .B(_10223_),
    .C(_10241_),
    .Y(_10457_));
 sg13g2_and3_1 _17287_ (.X(_10458_),
    .A(net1045),
    .B(_10223_),
    .C(net905));
 sg13g2_inv_1 _17288_ (.Y(_10459_),
    .A(_00256_));
 sg13g2_a22oi_1 _17289_ (.Y(_10460_),
    .B1(_10458_),
    .B2(_10459_),
    .A2(_10457_),
    .A1(_10456_));
 sg13g2_nand2b_1 _17290_ (.Y(_10461_),
    .B(net681),
    .A_N(_10460_));
 sg13g2_a22oi_1 _17291_ (.Y(_10462_),
    .B1(net775),
    .B2(\cpu.ex.r_10[14] ),
    .A2(_10432_),
    .A1(\cpu.ex.r_9[14] ));
 sg13g2_nand2b_1 _17292_ (.Y(_10463_),
    .B(net680),
    .A_N(_10462_));
 sg13g2_mux2_1 _17293_ (.A0(\cpu.ex.r_epc[14] ),
    .A1(\cpu.ex.r_11[14] ),
    .S(net618),
    .X(_10464_));
 sg13g2_nor2_1 _17294_ (.A(net571),
    .B(_10371_),
    .Y(_10465_));
 sg13g2_mux2_1 _17295_ (.A0(\cpu.ex.r_12[14] ),
    .A1(\cpu.ex.r_13[14] ),
    .S(net570),
    .X(_10466_));
 sg13g2_a22oi_1 _17296_ (.Y(_10467_),
    .B1(_10466_),
    .B2(_10305_),
    .A2(_10465_),
    .A1(_10464_));
 sg13g2_inv_1 _17297_ (.Y(_10468_),
    .A(\cpu.ex.r_8[14] ));
 sg13g2_nand3_1 _17298_ (.B(net776),
    .C(_10245_),
    .A(\cpu.ex.r_14[14] ),
    .Y(_10469_));
 sg13g2_o21ai_1 _17299_ (.B1(_10469_),
    .Y(_10470_),
    .A1(_10468_),
    .A2(_10409_));
 sg13g2_inv_1 _17300_ (.Y(_10471_),
    .A(\cpu.ex.r_lr[14] ));
 sg13g2_nand3_1 _17301_ (.B(net681),
    .C(net571),
    .A(\cpu.ex.r_mult[30] ),
    .Y(_10472_));
 sg13g2_o21ai_1 _17302_ (.B1(_10472_),
    .Y(_10473_),
    .A1(_10471_),
    .A2(_10409_));
 sg13g2_buf_2 _17303_ (.A(\cpu.ex.mmu_read[14] ),
    .X(_10474_));
 sg13g2_nand3b_1 _17304_ (.B(net570),
    .C(_10474_),
    .Y(_10475_),
    .A_N(net776));
 sg13g2_nand3b_1 _17305_ (.B(net681),
    .C(\cpu.ex.r_stmp[14] ),
    .Y(_10476_),
    .A_N(net570));
 sg13g2_nand2b_1 _17306_ (.Y(_10477_),
    .B(net571),
    .A_N(_10308_));
 sg13g2_a21oi_1 _17307_ (.A1(_10475_),
    .A2(_10476_),
    .Y(_10478_),
    .B1(_10477_));
 sg13g2_a221oi_1 _17308_ (.B2(_10356_),
    .C1(_10478_),
    .B1(_10473_),
    .A1(_10354_),
    .Y(_10479_),
    .A2(_10470_));
 sg13g2_nand4_1 _17309_ (.B(_10463_),
    .C(_10467_),
    .A(_10461_),
    .Y(_10480_),
    .D(_10479_));
 sg13g2_a22oi_1 _17310_ (.Y(_10481_),
    .B1(net513),
    .B2(_10480_),
    .A2(net512),
    .A1(net688));
 sg13g2_nor2_1 _17311_ (.A(net902),
    .B(\cpu.dec.imm[14] ),
    .Y(_10482_));
 sg13g2_a21oi_1 _17312_ (.A1(net902),
    .A2(_10481_),
    .Y(_10483_),
    .B1(_10482_));
 sg13g2_nor2_1 _17313_ (.A(net909),
    .B(_00185_),
    .Y(_10484_));
 sg13g2_a21o_1 _17314_ (.A2(_10483_),
    .A1(net770),
    .B1(_10484_),
    .X(_10485_));
 sg13g2_buf_1 _17315_ (.A(_10485_),
    .X(_10486_));
 sg13g2_buf_2 _17316_ (.A(_00277_),
    .X(_10487_));
 sg13g2_inv_1 _17317_ (.Y(_10488_),
    .A(_10487_));
 sg13g2_nand2_1 _17318_ (.Y(_10489_),
    .A(net901),
    .B(_10488_));
 sg13g2_nand2_1 _17319_ (.Y(_10490_),
    .A(net904),
    .B(net682));
 sg13g2_nand2_1 _17320_ (.Y(_10491_),
    .A(\cpu.ex.r_9[8] ),
    .B(_10239_));
 sg13g2_o21ai_1 _17321_ (.B1(_10491_),
    .Y(_10492_),
    .A1(_00250_),
    .A2(_10490_));
 sg13g2_nand2_1 _17322_ (.Y(_10493_),
    .A(_10230_),
    .B(net773));
 sg13g2_and2_1 _17323_ (.A(\cpu.ex.r_14[8] ),
    .B(net682),
    .X(_10494_));
 sg13g2_a21oi_1 _17324_ (.A1(\cpu.ex.r_10[8] ),
    .A2(net772),
    .Y(_10495_),
    .B1(_10494_));
 sg13g2_nand3_1 _17325_ (.B(net619),
    .C(_10262_),
    .A(\cpu.ex.r_mult[24] ),
    .Y(_10496_));
 sg13g2_o21ai_1 _17326_ (.B1(_10496_),
    .Y(_10497_),
    .A1(_10493_),
    .A2(_10495_));
 sg13g2_nand2_1 _17327_ (.Y(_10498_),
    .A(net1048),
    .B(_10350_));
 sg13g2_and2_1 _17328_ (.A(_10209_),
    .B(_10212_),
    .X(_10499_));
 sg13g2_buf_1 _17329_ (.A(_10499_),
    .X(_10500_));
 sg13g2_nor2_2 _17330_ (.A(_10235_),
    .B(net1051),
    .Y(_10501_));
 sg13g2_a22oi_1 _17331_ (.Y(_10502_),
    .B1(_10501_),
    .B2(\cpu.ex.r_lr[8] ),
    .A2(_10500_),
    .A1(\cpu.ex.r_11[8] ));
 sg13g2_nor2_1 _17332_ (.A(_10498_),
    .B(_10502_),
    .Y(_10503_));
 sg13g2_a221oi_1 _17333_ (.B2(net681),
    .C1(_10503_),
    .B1(_10497_),
    .A1(_10398_),
    .Y(_10504_),
    .A2(_10492_));
 sg13g2_buf_1 _17334_ (.A(\cpu.ex.r_sp[8] ),
    .X(_10505_));
 sg13g2_nand3_1 _17335_ (.B(net772),
    .C(net771),
    .A(_10505_),
    .Y(_10506_));
 sg13g2_nand3_1 _17336_ (.B(net620),
    .C(net777),
    .A(\cpu.ex.r_12[8] ),
    .Y(_10507_));
 sg13g2_nand3_1 _17337_ (.B(net776),
    .C(_10262_),
    .A(\cpu.ex.r_stmp[8] ),
    .Y(_10508_));
 sg13g2_nand3_1 _17338_ (.B(_10400_),
    .C(net680),
    .A(\cpu.ex.r_8[8] ),
    .Y(_10509_));
 sg13g2_nand4_1 _17339_ (.B(_10507_),
    .C(_10508_),
    .A(_10506_),
    .Y(_10510_),
    .D(_10509_));
 sg13g2_nand3_1 _17340_ (.B(net620),
    .C(net777),
    .A(\cpu.ex.r_13[8] ),
    .Y(_10511_));
 sg13g2_nand3_1 _17341_ (.B(_10352_),
    .C(net771),
    .A(\cpu.ex.r_epc[8] ),
    .Y(_10512_));
 sg13g2_nand3_1 _17342_ (.B(_10511_),
    .C(_10512_),
    .A(_10280_),
    .Y(_10513_));
 sg13g2_o21ai_1 _17343_ (.B1(_10513_),
    .Y(_10514_),
    .A1(_10281_),
    .A2(_10510_));
 sg13g2_a21o_1 _17344_ (.A2(_10514_),
    .A1(_10504_),
    .B1(net572),
    .X(_10515_));
 sg13g2_buf_2 _17345_ (.A(_10515_),
    .X(_10516_));
 sg13g2_a21oi_1 _17346_ (.A1(net1139),
    .A2(_10286_),
    .Y(_10517_),
    .B1(_10301_));
 sg13g2_o21ai_1 _17347_ (.B1(_10206_),
    .Y(_10518_),
    .A1(net902),
    .A2(\cpu.dec.imm[8] ));
 sg13g2_a21o_1 _17348_ (.A2(_10517_),
    .A1(_10516_),
    .B1(_10518_),
    .X(_10519_));
 sg13g2_buf_1 _17349_ (.A(_10519_),
    .X(_10520_));
 sg13g2_nand2_1 _17350_ (.Y(_10521_),
    .A(_10489_),
    .B(_10520_));
 sg13g2_buf_2 _17351_ (.A(_10521_),
    .X(_10522_));
 sg13g2_buf_1 _17352_ (.A(_10522_),
    .X(_10523_));
 sg13g2_buf_2 _17353_ (.A(\cpu.addr[9] ),
    .X(_10524_));
 sg13g2_a22oi_1 _17354_ (.Y(_10525_),
    .B1(_10262_),
    .B2(\cpu.ex.r_mult[25] ),
    .A2(net680),
    .A1(\cpu.ex.r_11[9] ));
 sg13g2_nand3b_1 _17355_ (.B(net679),
    .C(\cpu.ex.r_epc[9] ),
    .Y(_10526_),
    .A_N(net682));
 sg13g2_nand3b_1 _17356_ (.B(net682),
    .C(\cpu.ex.r_stmp[9] ),
    .Y(_10527_),
    .A_N(net679));
 sg13g2_a21o_1 _17357_ (.A2(_10527_),
    .A1(_10526_),
    .B1(_10325_),
    .X(_10528_));
 sg13g2_o21ai_1 _17358_ (.B1(_10528_),
    .Y(_10529_),
    .A1(_10371_),
    .A2(_10525_));
 sg13g2_buf_1 _17359_ (.A(\cpu.ex.r_sp[9] ),
    .X(_10530_));
 sg13g2_mux2_1 _17360_ (.A0(_10530_),
    .A1(\cpu.ex.r_10[9] ),
    .S(_10307_),
    .X(_10531_));
 sg13g2_mux2_1 _17361_ (.A0(\cpu.ex.r_lr[9] ),
    .A1(\cpu.ex.r_9[9] ),
    .S(_10307_),
    .X(_10532_));
 sg13g2_a22oi_1 _17362_ (.Y(_10533_),
    .B1(_10532_),
    .B2(_10432_),
    .A2(_10531_),
    .A1(_10272_));
 sg13g2_nor2_1 _17363_ (.A(_10244_),
    .B(_10533_),
    .Y(_10534_));
 sg13g2_nand2_1 _17364_ (.Y(_10535_),
    .A(_10242_),
    .B(_10247_));
 sg13g2_and2_1 _17365_ (.A(\cpu.ex.r_13[9] ),
    .B(net679),
    .X(_10536_));
 sg13g2_a21oi_1 _17366_ (.A1(\cpu.ex.r_12[9] ),
    .A2(_10231_),
    .Y(_10537_),
    .B1(_10536_));
 sg13g2_nand3_1 _17367_ (.B(_10221_),
    .C(_10260_),
    .A(\cpu.ex.r_8[9] ),
    .Y(_10538_));
 sg13g2_o21ai_1 _17368_ (.B1(_10538_),
    .Y(_10539_),
    .A1(_10535_),
    .A2(_10537_));
 sg13g2_nand2_1 _17369_ (.Y(_10540_),
    .A(net1049),
    .B(net908));
 sg13g2_nor2b_1 _17370_ (.A(_00251_),
    .B_N(_10280_),
    .Y(_10541_));
 sg13g2_a21oi_1 _17371_ (.A1(\cpu.ex.r_14[9] ),
    .A2(_10232_),
    .Y(_10542_),
    .B1(_10541_));
 sg13g2_nor3_1 _17372_ (.A(net772),
    .B(_10540_),
    .C(_10542_),
    .Y(_10543_));
 sg13g2_or4_1 _17373_ (.A(_10529_),
    .B(_10534_),
    .C(_10539_),
    .D(_10543_),
    .X(_10544_));
 sg13g2_a221oi_1 _17374_ (.B2(_10544_),
    .C1(_10301_),
    .B1(_10339_),
    .A1(_10524_),
    .Y(_10545_),
    .A2(net569));
 sg13g2_o21ai_1 _17375_ (.B1(_10205_),
    .Y(_10546_),
    .A1(net1047),
    .A2(\cpu.dec.imm[9] ));
 sg13g2_buf_1 _17376_ (.A(_00276_),
    .X(_10547_));
 sg13g2_inv_1 _17377_ (.Y(_10548_),
    .A(_10547_));
 sg13g2_nand2_1 _17378_ (.Y(_10549_),
    .A(net901),
    .B(_10548_));
 sg13g2_o21ai_1 _17379_ (.B1(_10549_),
    .Y(_10550_),
    .A1(_10545_),
    .A2(_10546_));
 sg13g2_buf_1 _17380_ (.A(_10550_),
    .X(_10551_));
 sg13g2_buf_1 _17381_ (.A(net242),
    .X(_10552_));
 sg13g2_nor4_1 _17382_ (.A(_10455_),
    .B(net201),
    .C(net169),
    .D(net220),
    .Y(_10553_));
 sg13g2_and2_1 _17383_ (.A(\cpu.ex.r_stmp[2] ),
    .B(net1050),
    .X(_10554_));
 sg13g2_nor2b_1 _17384_ (.A(net1050),
    .B_N(\cpu.ex.r_8[2] ),
    .Y(_10555_));
 sg13g2_a22oi_1 _17385_ (.Y(_10556_),
    .B1(_10555_),
    .B2(_10247_),
    .A2(_10554_),
    .A1(_10361_));
 sg13g2_nand3b_1 _17386_ (.B(net1051),
    .C(\cpu.ex.r_9[2] ),
    .Y(_10557_),
    .A_N(net1050));
 sg13g2_buf_1 _17387_ (.A(\cpu.ex.mmu_read[2] ),
    .X(_10558_));
 sg13g2_nand3b_1 _17388_ (.B(net1050),
    .C(net1121),
    .Y(_10559_),
    .A_N(net1051));
 sg13g2_nand2b_1 _17389_ (.Y(_10560_),
    .B(net1123),
    .A_N(_10209_));
 sg13g2_a21o_1 _17390_ (.A2(_10559_),
    .A1(_10557_),
    .B1(_10560_),
    .X(_10561_));
 sg13g2_o21ai_1 _17391_ (.B1(_10561_),
    .Y(_10562_),
    .A1(net1045),
    .A2(_10556_));
 sg13g2_a22oi_1 _17392_ (.Y(_10563_),
    .B1(_10501_),
    .B2(\cpu.ex.r_lr[2] ),
    .A2(_10500_),
    .A1(\cpu.ex.r_11[2] ));
 sg13g2_nor2_1 _17393_ (.A(_10498_),
    .B(_10563_),
    .Y(_10564_));
 sg13g2_mux2_1 _17394_ (.A0(net1146),
    .A1(\cpu.ex.r_12[2] ),
    .S(net1051),
    .X(_10565_));
 sg13g2_nand2_1 _17395_ (.Y(_10566_),
    .A(_10221_),
    .B(_10565_));
 sg13g2_nor2b_1 _17396_ (.A(_00244_),
    .B_N(net1123),
    .Y(_10567_));
 sg13g2_nor2b_1 _17397_ (.A(net1123),
    .B_N(\cpu.ex.r_14[2] ),
    .Y(_10568_));
 sg13g2_o21ai_1 _17398_ (.B1(_10500_),
    .Y(_10569_),
    .A1(_10567_),
    .A2(_10568_));
 sg13g2_a21oi_1 _17399_ (.A1(_10566_),
    .A2(_10569_),
    .Y(_10570_),
    .B1(net900));
 sg13g2_nand4_1 _17400_ (.B(net1048),
    .C(net907),
    .A(\cpu.ex.r_13[2] ),
    .Y(_10571_),
    .D(_10247_));
 sg13g2_mux2_1 _17401_ (.A0(\cpu.ex.r_epc[2] ),
    .A1(\cpu.ex.r_mult[18] ),
    .S(net1050),
    .X(_10572_));
 sg13g2_nand3_1 _17402_ (.B(_10361_),
    .C(_10572_),
    .A(net1048),
    .Y(_10573_));
 sg13g2_buf_1 _17403_ (.A(\cpu.ex.r_sp[2] ),
    .X(_10574_));
 sg13g2_mux2_1 _17404_ (.A0(_10574_),
    .A1(\cpu.ex.r_10[2] ),
    .S(net1051),
    .X(_10575_));
 sg13g2_nand3_1 _17405_ (.B(_10271_),
    .C(_10575_),
    .A(net900),
    .Y(_10576_));
 sg13g2_nand3_1 _17406_ (.B(_10573_),
    .C(_10576_),
    .A(_10571_),
    .Y(_10577_));
 sg13g2_or4_1 _17407_ (.A(_10562_),
    .B(_10564_),
    .C(_10570_),
    .D(_10577_),
    .X(_10578_));
 sg13g2_nand2_2 _17408_ (.Y(_10579_),
    .A(_10205_),
    .B(_10289_));
 sg13g2_a221oi_1 _17409_ (.B2(_10578_),
    .C1(_10579_),
    .B1(_10338_),
    .A1(_09229_),
    .Y(_10580_),
    .A2(net569));
 sg13g2_buf_1 _17410_ (.A(_10580_),
    .X(_10581_));
 sg13g2_buf_1 _17411_ (.A(_00281_),
    .X(_10582_));
 sg13g2_buf_1 _17412_ (.A(\cpu.dec.imm[2] ),
    .X(_10583_));
 sg13g2_nor3_1 _17413_ (.A(_10583_),
    .B(_10204_),
    .C(net1047),
    .Y(_10584_));
 sg13g2_a21o_1 _17414_ (.A2(_10582_),
    .A1(_10204_),
    .B1(_10584_),
    .X(_10585_));
 sg13g2_buf_1 _17415_ (.A(_10585_),
    .X(_10586_));
 sg13g2_or2_1 _17416_ (.X(_10587_),
    .B(_10586_),
    .A(_10581_));
 sg13g2_buf_1 _17417_ (.A(_10587_),
    .X(_10588_));
 sg13g2_buf_1 _17418_ (.A(_10588_),
    .X(_10589_));
 sg13g2_nand2b_1 _17419_ (.Y(_10590_),
    .B(net773),
    .A_N(_00245_));
 sg13g2_nand2b_1 _17420_ (.Y(_10591_),
    .B(\cpu.ex.r_mult[19] ),
    .A_N(net773));
 sg13g2_nand2_1 _17421_ (.Y(_10592_),
    .A(net1048),
    .B(net907));
 sg13g2_a21oi_1 _17422_ (.A1(_10590_),
    .A2(_10591_),
    .Y(_10593_),
    .B1(_10592_));
 sg13g2_buf_1 _17423_ (.A(\cpu.ex.r_sp[3] ),
    .X(_10594_));
 sg13g2_mux4_1 _17424_ (.S0(net905),
    .A0(_10594_),
    .A1(\cpu.ex.r_stmp[3] ),
    .A2(\cpu.ex.r_10[3] ),
    .A3(\cpu.ex.r_14[3] ),
    .S1(net773),
    .X(_10595_));
 sg13g2_and2_1 _17425_ (.A(net906),
    .B(_10595_),
    .X(_10596_));
 sg13g2_o21ai_1 _17426_ (.B1(net776),
    .Y(_10597_),
    .A1(_10593_),
    .A2(_10596_));
 sg13g2_mux4_1 _17427_ (.S0(net904),
    .A0(\cpu.ex.r_lr[3] ),
    .A1(\cpu.ex.r_epc[3] ),
    .A2(\cpu.ex.r_9[3] ),
    .A3(\cpu.ex.r_11[3] ),
    .S1(net678),
    .X(_10598_));
 sg13g2_nand2_1 _17428_ (.Y(_10599_),
    .A(_10425_),
    .B(_10598_));
 sg13g2_nand2b_1 _17429_ (.Y(_10600_),
    .B(\cpu.ex.r_8[3] ),
    .A_N(net903));
 sg13g2_nand3_1 _17430_ (.B(net903),
    .C(net778),
    .A(\cpu.ex.r_13[3] ),
    .Y(_10601_));
 sg13g2_o21ai_1 _17431_ (.B1(_10601_),
    .Y(_10602_),
    .A1(net778),
    .A2(_10600_));
 sg13g2_nor2b_1 _17432_ (.A(net774),
    .B_N(\cpu.ex.r_12[3] ),
    .Y(_10603_));
 sg13g2_buf_1 _17433_ (.A(\cpu.ex.mmu_read[3] ),
    .X(_10604_));
 sg13g2_mux2_1 _17434_ (.A0(net1149),
    .A1(_10604_),
    .S(net903),
    .X(_10605_));
 sg13g2_and3_1 _17435_ (.X(_10606_),
    .A(_10242_),
    .B(_10501_),
    .C(_10605_));
 sg13g2_a221oi_1 _17436_ (.B2(_10305_),
    .C1(_10606_),
    .B1(_10603_),
    .A1(net777),
    .Y(_10607_),
    .A2(_10602_));
 sg13g2_and3_1 _17437_ (.X(_10608_),
    .A(_10597_),
    .B(_10599_),
    .C(_10607_));
 sg13g2_a21oi_1 _17438_ (.A1(_09291_),
    .A2(net569),
    .Y(_10609_),
    .B1(_10579_));
 sg13g2_o21ai_1 _17439_ (.B1(_10609_),
    .Y(_10610_),
    .A1(net572),
    .A2(_10608_));
 sg13g2_buf_2 _17440_ (.A(_10610_),
    .X(_10611_));
 sg13g2_buf_2 _17441_ (.A(_00181_),
    .X(_10612_));
 sg13g2_buf_1 _17442_ (.A(\cpu.dec.imm[3] ),
    .X(_10613_));
 sg13g2_nor2_1 _17443_ (.A(_10613_),
    .B(_10297_),
    .Y(_10614_));
 sg13g2_a22oi_1 _17444_ (.Y(_10615_),
    .B1(_10614_),
    .B2(_10301_),
    .A2(_10612_),
    .A1(net1046));
 sg13g2_buf_1 _17445_ (.A(_10615_),
    .X(_10616_));
 sg13g2_nand2_1 _17446_ (.Y(_10617_),
    .A(_10611_),
    .B(_10616_));
 sg13g2_buf_1 _17447_ (.A(_10617_),
    .X(_10618_));
 sg13g2_nand2_1 _17448_ (.Y(_10619_),
    .A(net286),
    .B(_10618_));
 sg13g2_buf_1 _17449_ (.A(_10619_),
    .X(_10620_));
 sg13g2_nor2_1 _17450_ (.A(_10204_),
    .B(_10301_),
    .Y(_10621_));
 sg13g2_buf_2 _17451_ (.A(_10621_),
    .X(_10622_));
 sg13g2_mux2_1 _17452_ (.A0(\cpu.ex.r_lr[1] ),
    .A1(\cpu.ex.mmu_read[1] ),
    .S(net1050),
    .X(_10623_));
 sg13g2_a221oi_1 _17453_ (.B2(_10233_),
    .C1(_10230_),
    .B1(_10623_),
    .A1(\cpu.ex.r_9[1] ),
    .Y(_10624_),
    .A2(_10259_));
 sg13g2_buf_1 _17454_ (.A(\cpu.ex.r_prev_ie ),
    .X(_10625_));
 sg13g2_a21oi_1 _17455_ (.A1(_10625_),
    .A2(_10262_),
    .Y(_10626_),
    .B1(net1045));
 sg13g2_or3_1 _17456_ (.A(net904),
    .B(_10624_),
    .C(_10626_),
    .X(_10627_));
 sg13g2_buf_1 _17457_ (.A(\cpu.ex.r_sp[1] ),
    .X(_10628_));
 sg13g2_mux4_1 _17458_ (.S0(net907),
    .A0(_10628_),
    .A1(\cpu.ex.r_stmp[1] ),
    .A2(\cpu.ex.r_10[1] ),
    .A3(\cpu.ex.r_14[1] ),
    .S1(net773),
    .X(_10629_));
 sg13g2_nand2_1 _17459_ (.Y(_10630_),
    .A(net775),
    .B(_10629_));
 sg13g2_mux2_1 _17460_ (.A0(\cpu.ex.r_12[1] ),
    .A1(\cpu.ex.r_13[1] ),
    .S(net1048),
    .X(_10631_));
 sg13g2_mux2_1 _17461_ (.A0(\cpu.ex.r_epc[1] ),
    .A1(\cpu.ex.r_mult[17] ),
    .S(net907),
    .X(_10632_));
 sg13g2_nor2_1 _17462_ (.A(_10230_),
    .B(_10325_),
    .Y(_10633_));
 sg13g2_nor3_1 _17463_ (.A(_00243_),
    .B(_10540_),
    .C(_10592_),
    .Y(_10634_));
 sg13g2_a221oi_1 _17464_ (.B2(_10633_),
    .C1(_10634_),
    .B1(_10632_),
    .A1(_10305_),
    .Y(_10635_),
    .A2(_10631_));
 sg13g2_a22oi_1 _17465_ (.Y(_10636_),
    .B1(_10428_),
    .B2(\cpu.ex.r_11[1] ),
    .A2(_10221_),
    .A1(\cpu.ex.r_8[1] ));
 sg13g2_nand2b_1 _17466_ (.Y(_10637_),
    .B(_10259_),
    .A_N(_10636_));
 sg13g2_nand4_1 _17467_ (.B(_10630_),
    .C(_10635_),
    .A(_10627_),
    .Y(_10638_),
    .D(_10637_));
 sg13g2_buf_1 _17468_ (.A(_10638_),
    .X(_10639_));
 sg13g2_nor3_1 _17469_ (.A(_10038_),
    .B(_10211_),
    .C(_10219_),
    .Y(_10640_));
 sg13g2_a21o_1 _17470_ (.A2(_10639_),
    .A1(_10338_),
    .B1(_10640_),
    .X(_10641_));
 sg13g2_buf_2 _17471_ (.A(_10641_),
    .X(_10642_));
 sg13g2_buf_1 _17472_ (.A(_00190_),
    .X(_10643_));
 sg13g2_inv_1 _17473_ (.Y(_10644_),
    .A(_10643_));
 sg13g2_buf_1 _17474_ (.A(\cpu.dec.imm[1] ),
    .X(_10645_));
 sg13g2_nor2b_1 _17475_ (.A(_10204_),
    .B_N(_10645_),
    .Y(_10646_));
 sg13g2_a22oi_1 _17476_ (.Y(_10647_),
    .B1(_10646_),
    .B2(_10301_),
    .A2(_10644_),
    .A1(net1046));
 sg13g2_inv_1 _17477_ (.Y(_10648_),
    .A(_10647_));
 sg13g2_a21oi_1 _17478_ (.A1(_10622_),
    .A2(_10642_),
    .Y(_10649_),
    .B1(_10648_));
 sg13g2_buf_1 _17479_ (.A(_10649_),
    .X(_10650_));
 sg13g2_buf_1 _17480_ (.A(\cpu.dec.imm[0] ),
    .X(_10651_));
 sg13g2_or2_1 _17481_ (.X(_10652_),
    .B(net1047),
    .A(_10651_));
 sg13g2_mux2_1 _17482_ (.A0(\cpu.ex.r_9[0] ),
    .A1(\cpu.ex.r_11[0] ),
    .S(_10251_),
    .X(_10653_));
 sg13g2_a22oi_1 _17483_ (.Y(_10654_),
    .B1(_10653_),
    .B2(_10278_),
    .A2(_10221_),
    .A1(\cpu.ex.r_8[0] ));
 sg13g2_inv_1 _17484_ (.Y(_10655_),
    .A(_10654_));
 sg13g2_inv_1 _17485_ (.Y(_10656_),
    .A(\cpu.ex.r_13[0] ));
 sg13g2_buf_1 _17486_ (.A(\cpu.ex.genblk3.r_prev_supmode ),
    .X(_10657_));
 sg13g2_nand3_1 _17487_ (.B(net900),
    .C(_10362_),
    .A(_10657_),
    .Y(_10658_));
 sg13g2_o21ai_1 _17488_ (.B1(_10658_),
    .Y(_10659_),
    .A1(_10656_),
    .A2(_10535_));
 sg13g2_a22oi_1 _17489_ (.Y(_10660_),
    .B1(_10368_),
    .B2(\cpu.ex.r_12[0] ),
    .A2(_10311_),
    .A1(\cpu.ex.r_10[0] ));
 sg13g2_nand4_1 _17490_ (.B(_10231_),
    .C(net682),
    .A(\cpu.ex.r_stmp[0] ),
    .Y(_10661_),
    .D(net771));
 sg13g2_o21ai_1 _17491_ (.B1(_10661_),
    .Y(_10662_),
    .A1(_10493_),
    .A2(_10660_));
 sg13g2_a221oi_1 _17492_ (.B2(_10279_),
    .C1(_10662_),
    .B1(_10659_),
    .A1(net680),
    .Y(_10663_),
    .A2(_10655_));
 sg13g2_mux2_1 _17493_ (.A0(\cpu.ex.r_mult[16] ),
    .A1(\cpu.ex.r_15[0] ),
    .S(_10306_),
    .X(_10664_));
 sg13g2_a22oi_1 _17494_ (.Y(_10665_),
    .B1(_10664_),
    .B2(_10278_),
    .A2(_10354_),
    .A1(\cpu.ex.r_14[0] ));
 sg13g2_nor2_1 _17495_ (.A(_10277_),
    .B(_10306_),
    .Y(_10666_));
 sg13g2_nand3_1 _17496_ (.B(_10400_),
    .C(_10666_),
    .A(_09160_),
    .Y(_10667_));
 sg13g2_o21ai_1 _17497_ (.B1(_10667_),
    .Y(_10668_),
    .A1(_10400_),
    .A2(_10665_));
 sg13g2_nand2_1 _17498_ (.Y(_10669_),
    .A(_10243_),
    .B(_10668_));
 sg13g2_a21o_1 _17499_ (.A2(_10669_),
    .A1(_10663_),
    .B1(net572),
    .X(_10670_));
 sg13g2_nand2_1 _17500_ (.Y(_10671_),
    .A(_08452_),
    .B(net569));
 sg13g2_nand3_1 _17501_ (.B(_10670_),
    .C(_10671_),
    .A(net1047),
    .Y(_10672_));
 sg13g2_nand3_1 _17502_ (.B(_10652_),
    .C(_10672_),
    .A(net770),
    .Y(_10673_));
 sg13g2_buf_1 _17503_ (.A(_10673_),
    .X(_10674_));
 sg13g2_nand2_1 _17504_ (.Y(_10675_),
    .A(net284),
    .B(_10674_));
 sg13g2_nor2_1 _17505_ (.A(_10620_),
    .B(_10675_),
    .Y(_10676_));
 sg13g2_buf_2 _17506_ (.A(_10676_),
    .X(_10677_));
 sg13g2_and4_1 _17507_ (.A(_10349_),
    .B(_10423_),
    .C(_10553_),
    .D(_10677_),
    .X(_10678_));
 sg13g2_buf_1 _17508_ (.A(_00279_),
    .X(_10679_));
 sg13g2_a22oi_1 _17509_ (.Y(_10680_),
    .B1(_10247_),
    .B2(\cpu.ex.r_9[6] ),
    .A2(_10361_),
    .A1(\cpu.ex.r_epc[6] ));
 sg13g2_nand3b_1 _17510_ (.B(net905),
    .C(\cpu.ex.r_14[6] ),
    .Y(_10681_),
    .A_N(net1045));
 sg13g2_nand3b_1 _17511_ (.B(net1045),
    .C(\cpu.ex.r_11[6] ),
    .Y(_10682_),
    .A_N(net905));
 sg13g2_a21o_1 _17512_ (.A2(_10682_),
    .A1(_10681_),
    .B1(_10540_),
    .X(_10683_));
 sg13g2_o21ai_1 _17513_ (.B1(_10683_),
    .Y(_10684_),
    .A1(_10498_),
    .A2(_10680_));
 sg13g2_buf_1 _17514_ (.A(\cpu.ex.r_sp[6] ),
    .X(_10685_));
 sg13g2_inv_1 _17515_ (.Y(_10686_),
    .A(_00248_));
 sg13g2_a22oi_1 _17516_ (.Y(_10687_),
    .B1(_10458_),
    .B2(_10686_),
    .A2(_10457_),
    .A1(_10685_));
 sg13g2_nor2_1 _17517_ (.A(_10400_),
    .B(_10687_),
    .Y(_10688_));
 sg13g2_a22oi_1 _17518_ (.Y(_10689_),
    .B1(_10356_),
    .B2(\cpu.ex.r_lr[6] ),
    .A2(_10354_),
    .A1(\cpu.ex.r_8[6] ));
 sg13g2_nand3_1 _17519_ (.B(_10271_),
    .C(_10259_),
    .A(\cpu.ex.r_10[6] ),
    .Y(_10690_));
 sg13g2_o21ai_1 _17520_ (.B1(_10690_),
    .Y(_10691_),
    .A1(_10409_),
    .A2(_10689_));
 sg13g2_nor2b_1 _17521_ (.A(_10277_),
    .B_N(\cpu.ex.r_stmp[6] ),
    .Y(_10692_));
 sg13g2_and2_1 _17522_ (.A(\cpu.ex.r_mult[22] ),
    .B(net1045),
    .X(_10693_));
 sg13g2_o21ai_1 _17523_ (.B1(net771),
    .Y(_10694_),
    .A1(_10692_),
    .A2(_10693_));
 sg13g2_mux2_1 _17524_ (.A0(\cpu.ex.r_12[6] ),
    .A1(\cpu.ex.r_13[6] ),
    .S(net1045),
    .X(_10695_));
 sg13g2_nand2_1 _17525_ (.Y(_10696_),
    .A(_10247_),
    .B(_10695_));
 sg13g2_a21oi_1 _17526_ (.A1(_10694_),
    .A2(_10696_),
    .Y(_10697_),
    .B1(net900));
 sg13g2_or4_1 _17527_ (.A(_10684_),
    .B(_10688_),
    .C(_10691_),
    .D(_10697_),
    .X(_10698_));
 sg13g2_buf_1 _17528_ (.A(_10698_),
    .X(_10699_));
 sg13g2_nor2_1 _17529_ (.A(net572),
    .B(_10579_),
    .Y(_10700_));
 sg13g2_and3_1 _17530_ (.X(_10701_),
    .A(_09220_),
    .B(_10334_),
    .C(_10336_));
 sg13g2_nor2_1 _17531_ (.A(_10204_),
    .B(net1047),
    .Y(_10702_));
 sg13g2_and2_1 _17532_ (.A(\cpu.dec.imm[6] ),
    .B(_10702_),
    .X(_10703_));
 sg13g2_a21o_1 _17533_ (.A2(_10701_),
    .A1(_10622_),
    .B1(_10703_),
    .X(_10704_));
 sg13g2_a21oi_1 _17534_ (.A1(_10699_),
    .A2(_10700_),
    .Y(_10705_),
    .B1(_10704_));
 sg13g2_o21ai_1 _17535_ (.B1(_10705_),
    .Y(_10706_),
    .A1(_10205_),
    .A2(_10679_));
 sg13g2_buf_1 _17536_ (.A(_10706_),
    .X(_10707_));
 sg13g2_inv_1 _17537_ (.Y(_10708_),
    .A(_00249_));
 sg13g2_a22oi_1 _17538_ (.Y(_10709_),
    .B1(_10239_),
    .B2(\cpu.ex.r_9[7] ),
    .A2(_10237_),
    .A1(_10708_));
 sg13g2_a221oi_1 _17539_ (.B2(\cpu.ex.r_lr[7] ),
    .C1(net773),
    .B1(_10239_),
    .A1(\cpu.ex.r_mult[23] ),
    .Y(_10710_),
    .A2(_10237_));
 sg13g2_a21oi_1 _17540_ (.A1(net678),
    .A2(_10709_),
    .Y(_10711_),
    .B1(_10710_));
 sg13g2_nand3_1 _17541_ (.B(net904),
    .C(_10262_),
    .A(\cpu.ex.r_stmp[7] ),
    .Y(_10712_));
 sg13g2_nand3_1 _17542_ (.B(_10400_),
    .C(_10259_),
    .A(\cpu.ex.r_8[7] ),
    .Y(_10713_));
 sg13g2_a21oi_1 _17543_ (.A1(_10712_),
    .A2(_10713_),
    .Y(_10714_),
    .B1(net679));
 sg13g2_a21oi_1 _17544_ (.A1(net679),
    .A2(_10711_),
    .Y(_10715_),
    .B1(_10714_));
 sg13g2_nand3b_1 _17545_ (.B(_10396_),
    .C(\cpu.ex.r_11[7] ),
    .Y(_10716_),
    .A_N(net905));
 sg13g2_nand3b_1 _17546_ (.B(net905),
    .C(\cpu.ex.r_14[7] ),
    .Y(_10717_),
    .A_N(_10396_));
 sg13g2_a21o_1 _17547_ (.A2(_10717_),
    .A1(_10716_),
    .B1(_10400_),
    .X(_10718_));
 sg13g2_nand3_1 _17548_ (.B(net903),
    .C(_10368_),
    .A(\cpu.ex.r_13[7] ),
    .Y(_10719_));
 sg13g2_nand3_1 _17549_ (.B(_10351_),
    .C(net775),
    .A(\cpu.ex.r_10[7] ),
    .Y(_10720_));
 sg13g2_nand4_1 _17550_ (.B(_10718_),
    .C(_10719_),
    .A(net678),
    .Y(_10721_),
    .D(_10720_));
 sg13g2_buf_1 _17551_ (.A(\cpu.ex.r_sp[7] ),
    .X(_10722_));
 sg13g2_buf_1 _17552_ (.A(\cpu.dec.user_io ),
    .X(_10723_));
 sg13g2_a22oi_1 _17553_ (.Y(_10724_),
    .B1(_10368_),
    .B2(_10723_),
    .A2(_10311_),
    .A1(_10722_));
 sg13g2_o21ai_1 _17554_ (.B1(net683),
    .Y(_10725_),
    .A1(net774),
    .A2(_10724_));
 sg13g2_nand3_1 _17555_ (.B(net778),
    .C(net777),
    .A(\cpu.ex.r_12[7] ),
    .Y(_10726_));
 sg13g2_nand4_1 _17556_ (.B(net774),
    .C(net900),
    .A(\cpu.ex.r_epc[7] ),
    .Y(_10727_),
    .D(net771));
 sg13g2_o21ai_1 _17557_ (.B1(_10727_),
    .Y(_10728_),
    .A1(net774),
    .A2(_10726_));
 sg13g2_a21oi_1 _17558_ (.A1(_10721_),
    .A2(_10725_),
    .Y(_10729_),
    .B1(_10728_));
 sg13g2_a21o_1 _17559_ (.A2(_10729_),
    .A1(_10715_),
    .B1(net572),
    .X(_10730_));
 sg13g2_buf_1 _17560_ (.A(_10730_),
    .X(_10731_));
 sg13g2_a21oi_1 _17561_ (.A1(\cpu.addr[7] ),
    .A2(_10286_),
    .Y(_10732_),
    .B1(_10579_));
 sg13g2_buf_1 _17562_ (.A(_00278_),
    .X(_10733_));
 sg13g2_inv_1 _17563_ (.Y(_10734_),
    .A(\cpu.dec.imm[7] ));
 sg13g2_a22oi_1 _17564_ (.Y(_10735_),
    .B1(_10734_),
    .B2(_10702_),
    .A2(_10733_),
    .A1(net1046));
 sg13g2_inv_1 _17565_ (.Y(_10736_),
    .A(_10735_));
 sg13g2_a21oi_1 _17566_ (.A1(_10731_),
    .A2(_10732_),
    .Y(_10737_),
    .B1(_10736_));
 sg13g2_buf_1 _17567_ (.A(_10737_),
    .X(_10738_));
 sg13g2_nor2_1 _17568_ (.A(_10707_),
    .B(net283),
    .Y(_10739_));
 sg13g2_inv_2 _17569_ (.Y(_10740_),
    .A(_00280_));
 sg13g2_a22oi_1 _17570_ (.Y(_10741_),
    .B1(\cpu.dec.imm[5] ),
    .B2(_10702_),
    .A2(_10740_),
    .A1(net1046));
 sg13g2_buf_1 _17571_ (.A(_10741_),
    .X(_10742_));
 sg13g2_inv_1 _17572_ (.Y(_10743_),
    .A(\cpu.addr[5] ));
 sg13g2_buf_1 _17573_ (.A(_10743_),
    .X(_10744_));
 sg13g2_nor3_2 _17574_ (.A(net1043),
    .B(_10211_),
    .C(_10219_),
    .Y(_10745_));
 sg13g2_a221oi_1 _17575_ (.B2(\cpu.ex.r_lr[5] ),
    .C1(net678),
    .B1(_10239_),
    .A1(\cpu.ex.r_mult[21] ),
    .Y(_10746_),
    .A2(_10237_));
 sg13g2_a221oi_1 _17576_ (.B2(\cpu.ex.r_13[5] ),
    .C1(_10234_),
    .B1(_10368_),
    .A1(\cpu.ex.r_11[5] ),
    .Y(_10747_),
    .A2(_10311_));
 sg13g2_nor3_1 _17577_ (.A(net906),
    .B(_10746_),
    .C(_10747_),
    .Y(_10748_));
 sg13g2_nand3b_1 _17578_ (.B(net778),
    .C(\cpu.ex.r_stmp[5] ),
    .Y(_10749_),
    .A_N(net903));
 sg13g2_nand3b_1 _17579_ (.B(net903),
    .C(\cpu.ex.r_epc[5] ),
    .Y(_10750_),
    .A_N(net778));
 sg13g2_a21o_1 _17580_ (.A2(_10750_),
    .A1(_10749_),
    .B1(_10325_),
    .X(_10751_));
 sg13g2_nand4_1 _17581_ (.B(net774),
    .C(net900),
    .A(\cpu.ex.r_9[5] ),
    .Y(_10752_),
    .D(_10248_));
 sg13g2_buf_1 _17582_ (.A(\cpu.ex.r_sp[5] ),
    .X(_10753_));
 sg13g2_nand4_1 _17583_ (.B(net906),
    .C(net900),
    .A(_10753_),
    .Y(_10754_),
    .D(net771));
 sg13g2_nand3_1 _17584_ (.B(_10752_),
    .C(_10754_),
    .A(_10751_),
    .Y(_10755_));
 sg13g2_nand3b_1 _17585_ (.B(_10237_),
    .C(_10398_),
    .Y(_10756_),
    .A_N(_00247_));
 sg13g2_mux2_1 _17586_ (.A0(\cpu.ex.r_8[5] ),
    .A1(\cpu.ex.r_12[5] ),
    .S(net778),
    .X(_10757_));
 sg13g2_nand3_1 _17587_ (.B(_10248_),
    .C(_10757_),
    .A(net906),
    .Y(_10758_));
 sg13g2_mux2_1 _17588_ (.A0(\cpu.ex.r_10[5] ),
    .A1(\cpu.ex.r_14[5] ),
    .S(net905),
    .X(_10759_));
 sg13g2_nand3_1 _17589_ (.B(_10272_),
    .C(_10759_),
    .A(net678),
    .Y(_10760_));
 sg13g2_nand3_1 _17590_ (.B(_10758_),
    .C(_10760_),
    .A(_10756_),
    .Y(_10761_));
 sg13g2_nor4_2 _17591_ (.A(_10745_),
    .B(_10748_),
    .C(_10755_),
    .Y(_10762_),
    .D(_10761_));
 sg13g2_nor2_1 _17592_ (.A(_10338_),
    .B(_10745_),
    .Y(_10763_));
 sg13g2_or3_1 _17593_ (.A(_10579_),
    .B(_10762_),
    .C(_10763_),
    .X(_10764_));
 sg13g2_buf_2 _17594_ (.A(_10764_),
    .X(_10765_));
 sg13g2_nand2_1 _17595_ (.Y(_10766_),
    .A(_10742_),
    .B(_10765_));
 sg13g2_buf_8 _17596_ (.A(_10766_),
    .X(_10767_));
 sg13g2_buf_1 _17597_ (.A(\cpu.ex.r_sp[4] ),
    .X(_10768_));
 sg13g2_a22oi_1 _17598_ (.Y(_10769_),
    .B1(_10666_),
    .B2(_10768_),
    .A2(_10398_),
    .A1(\cpu.ex.r_11[4] ));
 sg13g2_nand3_1 _17599_ (.B(net774),
    .C(_10362_),
    .A(\cpu.ex.r_epc[4] ),
    .Y(_10770_));
 sg13g2_o21ai_1 _17600_ (.B1(_10770_),
    .Y(_10771_),
    .A1(_10400_),
    .A2(_10769_));
 sg13g2_mux2_1 _17601_ (.A0(\cpu.ex.r_stmp[4] ),
    .A1(\cpu.ex.r_14[4] ),
    .S(net773),
    .X(_10772_));
 sg13g2_a22oi_1 _17602_ (.Y(_10773_),
    .B1(_10772_),
    .B2(net906),
    .A2(_10356_),
    .A1(\cpu.ex.r_mult[20] ));
 sg13g2_nor2_1 _17603_ (.A(_10490_),
    .B(_10773_),
    .Y(_10774_));
 sg13g2_a21oi_2 _17604_ (.B1(_10774_),
    .Y(_10775_),
    .A2(_10771_),
    .A1(net772));
 sg13g2_nand3b_1 _17605_ (.B(_10243_),
    .C(_10500_),
    .Y(_10776_),
    .A_N(_00246_));
 sg13g2_nand3_1 _17606_ (.B(_10351_),
    .C(_10501_),
    .A(\cpu.ex.r_lr[4] ),
    .Y(_10777_));
 sg13g2_a21oi_1 _17607_ (.A1(_10776_),
    .A2(_10777_),
    .Y(_10778_),
    .B1(net906));
 sg13g2_and4_1 _17608_ (.A(\cpu.ex.r_13[4] ),
    .B(net774),
    .C(net678),
    .D(_10368_),
    .X(_10779_));
 sg13g2_inv_1 _17609_ (.Y(_10780_),
    .A(\cpu.ex.r_10[4] ));
 sg13g2_nor4_1 _17610_ (.A(_10780_),
    .B(net679),
    .C(_10234_),
    .D(_10414_),
    .Y(_10781_));
 sg13g2_and2_1 _17611_ (.A(\cpu.ex.r_9[4] ),
    .B(net903),
    .X(_10782_));
 sg13g2_nand2_1 _17612_ (.Y(_10783_),
    .A(_10259_),
    .B(_10782_));
 sg13g2_o21ai_1 _17613_ (.B1(_10260_),
    .Y(_10784_),
    .A1(\cpu.ex.r_8[4] ),
    .A2(_10782_));
 sg13g2_a22oi_1 _17614_ (.Y(_10785_),
    .B1(_10262_),
    .B2(_08347_),
    .A2(_10255_),
    .A1(\cpu.ex.r_12[4] ));
 sg13g2_a221oi_1 _17615_ (.B2(_10785_),
    .C1(_10251_),
    .B1(_10784_),
    .A1(_10279_),
    .Y(_10786_),
    .A2(_10783_));
 sg13g2_nor4_2 _17616_ (.A(_10778_),
    .B(_10779_),
    .C(_10781_),
    .Y(_10787_),
    .D(_10786_));
 sg13g2_nand2_1 _17617_ (.Y(_10788_),
    .A(_10338_),
    .B(_10622_));
 sg13g2_a21o_1 _17618_ (.A2(_10787_),
    .A1(_10775_),
    .B1(_10788_),
    .X(_10789_));
 sg13g2_buf_2 _17619_ (.A(_10789_),
    .X(_10790_));
 sg13g2_inv_1 _17620_ (.Y(_10791_),
    .A(\cpu.dec.imm[4] ));
 sg13g2_nand4_1 _17621_ (.B(net1047),
    .C(_10334_),
    .A(_09403_),
    .Y(_10792_),
    .D(_10336_));
 sg13g2_o21ai_1 _17622_ (.B1(_10792_),
    .Y(_10793_),
    .A1(_10290_),
    .A2(_10791_));
 sg13g2_nand2_1 _17623_ (.Y(_10794_),
    .A(_08498_),
    .B(net1046));
 sg13g2_o21ai_1 _17624_ (.B1(_10794_),
    .Y(_10795_),
    .A1(net1046),
    .A2(_10793_));
 sg13g2_buf_2 _17625_ (.A(_10795_),
    .X(_10796_));
 sg13g2_nand2_1 _17626_ (.Y(_10797_),
    .A(_10790_),
    .B(_10796_));
 sg13g2_buf_8 _17627_ (.A(_10797_),
    .X(_10798_));
 sg13g2_nor2_1 _17628_ (.A(net282),
    .B(net281),
    .Y(_10799_));
 sg13g2_and2_1 _17629_ (.A(_10739_),
    .B(_10799_),
    .X(_10800_));
 sg13g2_buf_1 _17630_ (.A(net703),
    .X(_10801_));
 sg13g2_nor2_2 _17631_ (.A(net1133),
    .B(net616),
    .Y(_10802_));
 sg13g2_o21ai_1 _17632_ (.B1(_10802_),
    .Y(_10803_),
    .A1(_09345_),
    .A2(_09351_));
 sg13g2_a21oi_1 _17633_ (.A1(_10678_),
    .A2(_10800_),
    .Y(_10804_),
    .B1(_10803_));
 sg13g2_buf_1 _17634_ (.A(_10804_),
    .X(_10805_));
 sg13g2_buf_1 _17635_ (.A(_10805_),
    .X(_10806_));
 sg13g2_buf_1 _17636_ (.A(_10422_),
    .X(_10807_));
 sg13g2_buf_1 _17637_ (.A(_00286_),
    .X(_10808_));
 sg13g2_inv_1 _17638_ (.Y(_10809_),
    .A(_10808_));
 sg13g2_buf_1 _17639_ (.A(\cpu.ex.r_mult[22] ),
    .X(_10810_));
 sg13g2_inv_1 _17640_ (.Y(_10811_),
    .A(net1120));
 sg13g2_buf_1 _17641_ (.A(_00288_),
    .X(_10812_));
 sg13g2_buf_1 _17642_ (.A(_10812_),
    .X(_10813_));
 sg13g2_a21oi_1 _17643_ (.A1(_10811_),
    .A2(net1042),
    .Y(_10814_),
    .B1(net799));
 sg13g2_nand2b_1 _17644_ (.Y(_10815_),
    .B(_10739_),
    .A_N(_10814_));
 sg13g2_inv_1 _17645_ (.Y(_10816_),
    .A(_10679_));
 sg13g2_a221oi_1 _17646_ (.B2(_10700_),
    .C1(_10704_),
    .B1(_10699_),
    .A1(net1046),
    .Y(_10817_),
    .A2(_10816_));
 sg13g2_buf_8 _17647_ (.A(_10817_),
    .X(_10818_));
 sg13g2_or4_1 _17648_ (.A(net1120),
    .B(_10812_),
    .C(net361),
    .D(net283),
    .X(_10819_));
 sg13g2_xnor2_1 _17649_ (.Y(_10820_),
    .A(_10812_),
    .B(net361));
 sg13g2_nand3_1 _17650_ (.B(net283),
    .C(_10820_),
    .A(net1120),
    .Y(_10821_));
 sg13g2_a21o_1 _17651_ (.A2(_10821_),
    .A1(_10819_),
    .B1(net799),
    .X(_10822_));
 sg13g2_buf_2 _17652_ (.A(_00290_),
    .X(_10823_));
 sg13g2_nand3_1 _17653_ (.B(_10790_),
    .C(_10796_),
    .A(_10823_),
    .Y(_10824_));
 sg13g2_a21oi_2 _17654_ (.B1(_10788_),
    .Y(_10825_),
    .A2(_10787_),
    .A1(_10775_));
 sg13g2_mux2_1 _17655_ (.A0(net939),
    .A1(_10793_),
    .S(_10205_),
    .X(_10826_));
 sg13g2_buf_1 _17656_ (.A(_10826_),
    .X(_10827_));
 sg13g2_nor2_1 _17657_ (.A(_10823_),
    .B(net799),
    .Y(_10828_));
 sg13g2_o21ai_1 _17658_ (.B1(_10828_),
    .Y(_10829_),
    .A1(_10825_),
    .A2(_10827_));
 sg13g2_buf_2 _17659_ (.A(_00289_),
    .X(_10830_));
 sg13g2_inv_1 _17660_ (.Y(_10831_),
    .A(_10830_));
 sg13g2_a21oi_1 _17661_ (.A1(_10824_),
    .A2(_10829_),
    .Y(_10832_),
    .B1(_10831_));
 sg13g2_nor2_1 _17662_ (.A(_09316_),
    .B(_09336_),
    .Y(_10833_));
 sg13g2_buf_1 _17663_ (.A(_10833_),
    .X(_10834_));
 sg13g2_nand2_1 _17664_ (.Y(_10835_),
    .A(\cpu.dec.div ),
    .B(_10834_));
 sg13g2_buf_1 _17665_ (.A(_10835_),
    .X(_10836_));
 sg13g2_nor2_1 _17666_ (.A(_10836_),
    .B(net281),
    .Y(_10837_));
 sg13g2_and2_1 _17667_ (.A(_10742_),
    .B(_10765_),
    .X(_10838_));
 sg13g2_buf_2 _17668_ (.A(_10838_),
    .X(_10839_));
 sg13g2_o21ai_1 _17669_ (.B1(_10839_),
    .Y(_10840_),
    .A1(_10832_),
    .A2(_10837_));
 sg13g2_nor2_1 _17670_ (.A(_10825_),
    .B(_10827_),
    .Y(_10841_));
 sg13g2_buf_2 _17671_ (.A(_10841_),
    .X(_10842_));
 sg13g2_xnor2_1 _17672_ (.Y(_10843_),
    .A(_10823_),
    .B(_10842_));
 sg13g2_nor2_1 _17673_ (.A(_10830_),
    .B(net799),
    .Y(_10844_));
 sg13g2_nand3_1 _17674_ (.B(_10843_),
    .C(_10844_),
    .A(net282),
    .Y(_10845_));
 sg13g2_a22oi_1 _17675_ (.Y(_10846_),
    .B1(_10840_),
    .B2(_10845_),
    .A2(_10822_),
    .A1(_10815_));
 sg13g2_buf_1 _17676_ (.A(_00293_),
    .X(_10847_));
 sg13g2_a21o_1 _17677_ (.A2(_10642_),
    .A1(_10622_),
    .B1(_10648_),
    .X(_10848_));
 sg13g2_buf_1 _17678_ (.A(_10848_),
    .X(_10849_));
 sg13g2_nor2_1 _17679_ (.A(_10581_),
    .B(_10586_),
    .Y(_10850_));
 sg13g2_buf_8 _17680_ (.A(_10850_),
    .X(_10851_));
 sg13g2_buf_1 _17681_ (.A(_00292_),
    .X(_10852_));
 sg13g2_or2_1 _17682_ (.X(_10853_),
    .B(_09340_),
    .A(_10852_));
 sg13g2_buf_1 _17683_ (.A(_10853_),
    .X(_10854_));
 sg13g2_or2_1 _17684_ (.X(_10855_),
    .B(_10854_),
    .A(net360));
 sg13g2_buf_1 _17685_ (.A(_10855_),
    .X(_10856_));
 sg13g2_nand3_1 _17686_ (.B(net280),
    .C(_10856_),
    .A(_10847_),
    .Y(_10857_));
 sg13g2_or2_1 _17687_ (.X(_10858_),
    .B(net799),
    .A(_00291_));
 sg13g2_buf_1 _17688_ (.A(_10858_),
    .X(_10859_));
 sg13g2_a21oi_1 _17689_ (.A1(net360),
    .A2(_10854_),
    .Y(_10860_),
    .B1(_10859_));
 sg13g2_or2_1 _17690_ (.X(_10861_),
    .B(_09340_),
    .A(_10847_));
 sg13g2_buf_1 _17691_ (.A(_10861_),
    .X(_10862_));
 sg13g2_and2_1 _17692_ (.A(_10611_),
    .B(_10616_),
    .X(_10863_));
 sg13g2_buf_1 _17693_ (.A(_10863_),
    .X(_10864_));
 sg13g2_a221oi_1 _17694_ (.B2(net360),
    .C1(_10864_),
    .B1(_10854_),
    .A1(net280),
    .Y(_10865_),
    .A2(_10862_));
 sg13g2_a21o_1 _17695_ (.A2(_10860_),
    .A1(_10857_),
    .B1(_10865_),
    .X(_10866_));
 sg13g2_buf_1 _17696_ (.A(_10866_),
    .X(_10867_));
 sg13g2_and3_1 _17697_ (.X(_10868_),
    .A(_10205_),
    .B(_10652_),
    .C(_10672_));
 sg13g2_buf_2 _17698_ (.A(_10868_),
    .X(_10869_));
 sg13g2_o21ai_1 _17699_ (.B1(_10869_),
    .Y(_10870_),
    .A1(net280),
    .A2(_10862_));
 sg13g2_nor3_1 _17700_ (.A(net360),
    .B(_10859_),
    .C(_10854_),
    .Y(_10871_));
 sg13g2_a21oi_1 _17701_ (.A1(_10859_),
    .A2(_10856_),
    .Y(_10872_),
    .B1(_10864_));
 sg13g2_or2_1 _17702_ (.X(_10873_),
    .B(_10872_),
    .A(_10871_));
 sg13g2_a21o_1 _17703_ (.A2(_10870_),
    .A1(_10867_),
    .B1(_10873_),
    .X(_10874_));
 sg13g2_or2_1 _17704_ (.X(_10875_),
    .B(_10612_),
    .A(net1068));
 sg13g2_nand3_1 _17705_ (.B(_10644_),
    .C(_09342_),
    .A(net1068),
    .Y(_10876_));
 sg13g2_a21oi_1 _17706_ (.A1(_10875_),
    .A2(_10876_),
    .Y(_10877_),
    .B1(_09332_));
 sg13g2_nand3b_1 _17707_ (.B(_09344_),
    .C(net1068),
    .Y(_10878_),
    .A_N(_10582_));
 sg13g2_o21ai_1 _17708_ (.B1(_10878_),
    .Y(_10879_),
    .A1(_10612_),
    .A2(_09342_));
 sg13g2_or2_1 _17709_ (.X(_10880_),
    .B(_10879_),
    .A(_10877_));
 sg13g2_and2_1 _17710_ (.A(net1127),
    .B(_10217_),
    .X(_10881_));
 sg13g2_buf_8 _17711_ (.A(\cpu.dec.r_rs1[3] ),
    .X(_10882_));
 sg13g2_xor2_1 _17712_ (.B(_10882_),
    .A(_10190_),
    .X(_10883_));
 sg13g2_buf_2 _17713_ (.A(\cpu.dec.r_rs1[0] ),
    .X(_10884_));
 sg13g2_xor2_1 _17714_ (.B(_10884_),
    .A(_10196_),
    .X(_10885_));
 sg13g2_buf_8 _17715_ (.A(\cpu.dec.r_rs1[2] ),
    .X(_10886_));
 sg13g2_xor2_1 _17716_ (.B(net1119),
    .A(net1052),
    .X(_10887_));
 sg13g2_buf_8 _17717_ (.A(\cpu.dec.r_rs1[1] ),
    .X(_10888_));
 sg13g2_xor2_1 _17718_ (.B(_10888_),
    .A(_10195_),
    .X(_10889_));
 sg13g2_nor4_1 _17719_ (.A(_10883_),
    .B(_10885_),
    .C(_10887_),
    .D(_10889_),
    .Y(_10890_));
 sg13g2_and2_1 _17720_ (.A(_10881_),
    .B(_10890_),
    .X(_10891_));
 sg13g2_buf_8 _17721_ (.A(_10891_),
    .X(_10892_));
 sg13g2_buf_1 _17722_ (.A(_10892_),
    .X(_10893_));
 sg13g2_nor2_2 _17723_ (.A(net1118),
    .B(_10882_),
    .Y(_10894_));
 sg13g2_buf_8 _17724_ (.A(net1118),
    .X(_10895_));
 sg13g2_buf_8 _17725_ (.A(_10882_),
    .X(_10896_));
 sg13g2_and2_1 _17726_ (.A(net1041),
    .B(_10896_),
    .X(_10897_));
 sg13g2_buf_1 _17727_ (.A(_10897_),
    .X(_10898_));
 sg13g2_a22oi_1 _17728_ (.Y(_10899_),
    .B1(_10898_),
    .B2(\cpu.ex.r_11[2] ),
    .A2(_10894_),
    .A1(\cpu.ex.r_lr[2] ));
 sg13g2_buf_8 _17729_ (.A(_10884_),
    .X(_10900_));
 sg13g2_buf_8 _17730_ (.A(_10900_),
    .X(_10901_));
 sg13g2_buf_8 _17731_ (.A(net899),
    .X(_10902_));
 sg13g2_buf_1 _17732_ (.A(net769),
    .X(_10903_));
 sg13g2_nand2b_1 _17733_ (.Y(_10904_),
    .B(net677),
    .A_N(_10899_));
 sg13g2_buf_1 _17734_ (.A(net1040),
    .X(_10905_));
 sg13g2_nand2b_1 _17735_ (.Y(_10906_),
    .B(net1041),
    .A_N(net1039));
 sg13g2_buf_2 _17736_ (.A(_10906_),
    .X(_10907_));
 sg13g2_nor2_2 _17737_ (.A(net898),
    .B(_10907_),
    .Y(_10908_));
 sg13g2_nor2b_1 _17738_ (.A(net1118),
    .B_N(_10884_),
    .Y(_10909_));
 sg13g2_buf_1 _17739_ (.A(_10909_),
    .X(_10910_));
 sg13g2_buf_1 _17740_ (.A(_10910_),
    .X(_10911_));
 sg13g2_and2_1 _17741_ (.A(net898),
    .B(net768),
    .X(_10912_));
 sg13g2_buf_1 _17742_ (.A(_10912_),
    .X(_10913_));
 sg13g2_a22oi_1 _17743_ (.Y(_10914_),
    .B1(_10913_),
    .B2(\cpu.ex.r_9[2] ),
    .A2(_10908_),
    .A1(_10574_));
 sg13g2_buf_8 _17744_ (.A(net1119),
    .X(_10915_));
 sg13g2_buf_1 _17745_ (.A(net1038),
    .X(_10916_));
 sg13g2_buf_1 _17746_ (.A(net897),
    .X(_10917_));
 sg13g2_a21oi_1 _17747_ (.A1(_10904_),
    .A2(_10914_),
    .Y(_10918_),
    .B1(net767));
 sg13g2_inv_2 _17748_ (.Y(_10919_),
    .A(net1119));
 sg13g2_buf_1 _17749_ (.A(_10919_),
    .X(_10920_));
 sg13g2_a22oi_1 _17750_ (.Y(_10921_),
    .B1(_10913_),
    .B2(\cpu.ex.r_13[2] ),
    .A2(_10908_),
    .A1(\cpu.ex.r_stmp[2] ));
 sg13g2_and3_1 _17751_ (.X(_10922_),
    .A(net899),
    .B(net1041),
    .C(net1119));
 sg13g2_buf_2 _17752_ (.A(_10922_),
    .X(_10923_));
 sg13g2_inv_2 _17753_ (.Y(_10924_),
    .A(net1040));
 sg13g2_nand2b_1 _17754_ (.Y(_10925_),
    .B(\cpu.ex.r_mult[18] ),
    .A_N(net898));
 sg13g2_o21ai_1 _17755_ (.B1(_10925_),
    .Y(_10926_),
    .A1(_10924_),
    .A2(_00244_));
 sg13g2_and2_1 _17756_ (.A(net1039),
    .B(net1118),
    .X(_10927_));
 sg13g2_buf_2 _17757_ (.A(_10927_),
    .X(_10928_));
 sg13g2_nor2_1 _17758_ (.A(_10882_),
    .B(net1119),
    .Y(_10929_));
 sg13g2_buf_2 _17759_ (.A(_10929_),
    .X(_10930_));
 sg13g2_and2_1 _17760_ (.A(_10928_),
    .B(_10930_),
    .X(_10931_));
 sg13g2_buf_2 _17761_ (.A(_10931_),
    .X(_10932_));
 sg13g2_buf_1 _17762_ (.A(net898),
    .X(_10933_));
 sg13g2_nor2b_1 _17763_ (.A(net1039),
    .B_N(net1118),
    .Y(_10934_));
 sg13g2_buf_1 _17764_ (.A(_10934_),
    .X(_10935_));
 sg13g2_mux2_1 _17765_ (.A0(\cpu.ex.r_10[2] ),
    .A1(\cpu.ex.r_14[2] ),
    .S(net1038),
    .X(_10936_));
 sg13g2_and3_1 _17766_ (.X(_10937_),
    .A(net766),
    .B(_10935_),
    .C(_10936_));
 sg13g2_a221oi_1 _17767_ (.B2(\cpu.ex.r_epc[2] ),
    .C1(_10937_),
    .B1(_10932_),
    .A1(_10923_),
    .Y(_10938_),
    .A2(_10926_));
 sg13g2_o21ai_1 _17768_ (.B1(_10938_),
    .Y(_10939_),
    .A1(net896),
    .A2(_10921_));
 sg13g2_inv_2 _17769_ (.Y(_10940_),
    .A(net1041));
 sg13g2_nor2b_1 _17770_ (.A(_10882_),
    .B_N(net1119),
    .Y(_10941_));
 sg13g2_buf_2 _17771_ (.A(_10941_),
    .X(_10942_));
 sg13g2_mux2_1 _17772_ (.A0(\cpu.ex.r_8[2] ),
    .A1(\cpu.ex.r_12[2] ),
    .S(net1038),
    .X(_10943_));
 sg13g2_a22oi_1 _17773_ (.Y(_10944_),
    .B1(_10943_),
    .B2(net766),
    .A2(_10942_),
    .A1(net1146));
 sg13g2_buf_8 _17774_ (.A(_10942_),
    .X(_10945_));
 sg13g2_nand3_1 _17775_ (.B(net1121),
    .C(net765),
    .A(net769),
    .Y(_10946_));
 sg13g2_o21ai_1 _17776_ (.B1(_10946_),
    .Y(_10947_),
    .A1(net677),
    .A2(_10944_));
 sg13g2_and2_1 _17777_ (.A(net895),
    .B(_10947_),
    .X(_10948_));
 sg13g2_or4_1 _17778_ (.A(net568),
    .B(_10918_),
    .C(_10939_),
    .D(_10948_),
    .X(_10949_));
 sg13g2_buf_1 _17779_ (.A(_10949_),
    .X(_10950_));
 sg13g2_nand2_1 _17780_ (.Y(_10951_),
    .A(_09421_),
    .B(net568));
 sg13g2_nand4_1 _17781_ (.B(_09344_),
    .C(_10950_),
    .A(_09347_),
    .Y(_10952_),
    .D(_10951_));
 sg13g2_nand2_1 _17782_ (.Y(_10953_),
    .A(_09333_),
    .B(_10834_));
 sg13g2_nand2_1 _17783_ (.Y(_10954_),
    .A(_10953_),
    .B(_10836_));
 sg13g2_nand2_1 _17784_ (.Y(_10955_),
    .A(_10881_),
    .B(_10890_));
 sg13g2_buf_2 _17785_ (.A(_10955_),
    .X(_10956_));
 sg13g2_buf_1 _17786_ (.A(_10956_),
    .X(_10957_));
 sg13g2_inv_1 _17787_ (.Y(_10958_),
    .A(net1039));
 sg13g2_buf_1 _17788_ (.A(_10958_),
    .X(_10959_));
 sg13g2_nand3_1 _17789_ (.B(net895),
    .C(_10945_),
    .A(net1149),
    .Y(_10960_));
 sg13g2_buf_8 _17790_ (.A(net1041),
    .X(_10961_));
 sg13g2_buf_1 _17791_ (.A(net894),
    .X(_10962_));
 sg13g2_nor2b_1 _17792_ (.A(net1119),
    .B_N(_10882_),
    .Y(_10963_));
 sg13g2_buf_1 _17793_ (.A(_10963_),
    .X(_10964_));
 sg13g2_buf_1 _17794_ (.A(_10964_),
    .X(_10965_));
 sg13g2_nand3_1 _17795_ (.B(\cpu.ex.r_10[3] ),
    .C(_10965_),
    .A(_10962_),
    .Y(_10966_));
 sg13g2_nand3_1 _17796_ (.B(_10960_),
    .C(_10966_),
    .A(net764),
    .Y(_10967_));
 sg13g2_nand4_1 _17797_ (.B(_10924_),
    .C(net896),
    .A(_10962_),
    .Y(_10968_),
    .D(\cpu.ex.r_epc[3] ));
 sg13g2_nand3_1 _17798_ (.B(_10604_),
    .C(_10894_),
    .A(net897),
    .Y(_10969_));
 sg13g2_buf_8 _17799_ (.A(net1038),
    .X(_10970_));
 sg13g2_nor2b_1 _17800_ (.A(net893),
    .B_N(\cpu.ex.r_lr[3] ),
    .Y(_10971_));
 sg13g2_nor2b_1 _17801_ (.A(net897),
    .B_N(\cpu.ex.r_11[3] ),
    .Y(_10972_));
 sg13g2_a22oi_1 _17802_ (.Y(_10973_),
    .B1(_10972_),
    .B2(_10898_),
    .A2(_10971_),
    .A1(_10894_));
 sg13g2_and2_1 _17803_ (.A(net894),
    .B(\cpu.ex.r_mult[19] ),
    .X(_10974_));
 sg13g2_nor2b_1 _17804_ (.A(net893),
    .B_N(\cpu.ex.r_9[3] ),
    .Y(_10975_));
 sg13g2_nor2b_1 _17805_ (.A(net1041),
    .B_N(net1040),
    .Y(_10976_));
 sg13g2_a221oi_1 _17806_ (.B2(_10976_),
    .C1(net764),
    .B1(_10975_),
    .A1(net765),
    .Y(_10977_),
    .A2(_10974_));
 sg13g2_nand4_1 _17807_ (.B(_10969_),
    .C(_10973_),
    .A(_10968_),
    .Y(_10978_),
    .D(_10977_));
 sg13g2_and2_1 _17808_ (.A(_10882_),
    .B(net1119),
    .X(_10979_));
 sg13g2_buf_1 _17809_ (.A(_10979_),
    .X(_10980_));
 sg13g2_nand2_1 _17810_ (.Y(_10981_),
    .A(_10902_),
    .B(_10961_));
 sg13g2_nor2_1 _17811_ (.A(_10900_),
    .B(net1118),
    .Y(_10982_));
 sg13g2_buf_1 _17812_ (.A(_10982_),
    .X(_10983_));
 sg13g2_nand2_1 _17813_ (.Y(_10984_),
    .A(\cpu.ex.r_12[3] ),
    .B(net761));
 sg13g2_o21ai_1 _17814_ (.B1(_10984_),
    .Y(_10985_),
    .A1(_00245_),
    .A2(_10981_));
 sg13g2_buf_1 _17815_ (.A(net897),
    .X(_10986_));
 sg13g2_buf_1 _17816_ (.A(_10935_),
    .X(_10987_));
 sg13g2_buf_1 _17817_ (.A(net1040),
    .X(_10988_));
 sg13g2_mux2_1 _17818_ (.A0(\cpu.ex.r_stmp[3] ),
    .A1(\cpu.ex.r_14[3] ),
    .S(_10988_),
    .X(_10989_));
 sg13g2_nand3_1 _17819_ (.B(net676),
    .C(_10989_),
    .A(net760),
    .Y(_10990_));
 sg13g2_nand3_1 _17820_ (.B(net762),
    .C(net761),
    .A(\cpu.ex.r_8[3] ),
    .Y(_10991_));
 sg13g2_nand4_1 _17821_ (.B(net760),
    .C(\cpu.ex.r_13[3] ),
    .A(net766),
    .Y(_10992_),
    .D(net768));
 sg13g2_buf_1 _17822_ (.A(_10924_),
    .X(_10993_));
 sg13g2_nand4_1 _17823_ (.B(net896),
    .C(_10594_),
    .A(_10993_),
    .Y(_10994_),
    .D(net676));
 sg13g2_nand4_1 _17824_ (.B(_10991_),
    .C(_10992_),
    .A(_10990_),
    .Y(_10995_),
    .D(_10994_));
 sg13g2_a221oi_1 _17825_ (.B2(_10985_),
    .C1(_10995_),
    .B1(_10980_),
    .A1(_10967_),
    .Y(_10996_),
    .A2(_10978_));
 sg13g2_nor2_1 _17826_ (.A(_09458_),
    .B(_10956_),
    .Y(_10997_));
 sg13g2_a21oi_2 _17827_ (.B1(_10997_),
    .Y(_10998_),
    .A2(_10996_),
    .A1(net567));
 sg13g2_nand2_1 _17828_ (.Y(_10999_),
    .A(_10954_),
    .B(_10998_));
 sg13g2_nor2_1 _17829_ (.A(net899),
    .B(net898),
    .Y(_11000_));
 sg13g2_buf_8 _17830_ (.A(net1041),
    .X(_11001_));
 sg13g2_mux2_1 _17831_ (.A0(_10625_),
    .A1(\cpu.ex.r_stmp[1] ),
    .S(net891),
    .X(_11002_));
 sg13g2_nand2_1 _17832_ (.Y(_11003_),
    .A(_11000_),
    .B(_11002_));
 sg13g2_nor2b_1 _17833_ (.A(_00243_),
    .B_N(net891),
    .Y(_11004_));
 sg13g2_nor2b_1 _17834_ (.A(net891),
    .B_N(\cpu.ex.r_13[1] ),
    .Y(_11005_));
 sg13g2_and2_1 _17835_ (.A(net1039),
    .B(net1040),
    .X(_11006_));
 sg13g2_buf_1 _17836_ (.A(_11006_),
    .X(_11007_));
 sg13g2_o21ai_1 _17837_ (.B1(_11007_),
    .Y(_11008_),
    .A1(_11004_),
    .A2(_11005_));
 sg13g2_a21o_1 _17838_ (.A2(_11008_),
    .A1(_11003_),
    .B1(net896),
    .X(_11009_));
 sg13g2_and2_1 _17839_ (.A(_10919_),
    .B(_10910_),
    .X(_11010_));
 sg13g2_buf_1 _17840_ (.A(_11010_),
    .X(_11011_));
 sg13g2_mux2_1 _17841_ (.A0(\cpu.ex.r_lr[1] ),
    .A1(\cpu.ex.r_9[1] ),
    .S(net892),
    .X(_11012_));
 sg13g2_nand2_1 _17842_ (.Y(_11013_),
    .A(_11011_),
    .B(_11012_));
 sg13g2_and2_1 _17843_ (.A(net761),
    .B(_10980_),
    .X(_11014_));
 sg13g2_mux2_1 _17844_ (.A0(\cpu.ex.r_10[1] ),
    .A1(\cpu.ex.r_11[1] ),
    .S(net769),
    .X(_11015_));
 sg13g2_nand2_1 _17845_ (.Y(_11016_),
    .A(_10895_),
    .B(_10896_));
 sg13g2_nor2_1 _17846_ (.A(_10970_),
    .B(_11016_),
    .Y(_11017_));
 sg13g2_a22oi_1 _17847_ (.Y(_11018_),
    .B1(_11015_),
    .B2(_11017_),
    .A2(_11014_),
    .A1(\cpu.ex.r_12[1] ));
 sg13g2_nor2_2 _17848_ (.A(net1039),
    .B(_10886_),
    .Y(_11019_));
 sg13g2_nand2b_1 _17849_ (.Y(_11020_),
    .B(_10628_),
    .A_N(net1040));
 sg13g2_nand3b_1 _17850_ (.B(net898),
    .C(\cpu.ex.r_8[1] ),
    .Y(_11021_),
    .A_N(net891));
 sg13g2_o21ai_1 _17851_ (.B1(_11021_),
    .Y(_11022_),
    .A1(net895),
    .A2(_11020_));
 sg13g2_and2_1 _17852_ (.A(net1041),
    .B(net1038),
    .X(_11023_));
 sg13g2_buf_2 _17853_ (.A(_11023_),
    .X(_11024_));
 sg13g2_inv_1 _17854_ (.Y(_11025_),
    .A(\cpu.ex.r_mult[17] ));
 sg13g2_nand2b_1 _17855_ (.Y(_11026_),
    .B(net1039),
    .A_N(_10882_));
 sg13g2_buf_2 _17856_ (.A(_11026_),
    .X(_11027_));
 sg13g2_nand3b_1 _17857_ (.B(net898),
    .C(\cpu.ex.r_14[1] ),
    .Y(_11028_),
    .A_N(net899));
 sg13g2_o21ai_1 _17858_ (.B1(_11028_),
    .Y(_11029_),
    .A1(_11025_),
    .A2(_11027_));
 sg13g2_nand3b_1 _17859_ (.B(net893),
    .C(\cpu.ex.mmu_read[1] ),
    .Y(_11030_),
    .A_N(net891));
 sg13g2_nand3b_1 _17860_ (.B(\cpu.ex.r_epc[1] ),
    .C(net891),
    .Y(_11031_),
    .A_N(net1038));
 sg13g2_a21oi_1 _17861_ (.A1(_11030_),
    .A2(_11031_),
    .Y(_11032_),
    .B1(_11027_));
 sg13g2_a221oi_1 _17862_ (.B2(_11029_),
    .C1(_11032_),
    .B1(_11024_),
    .A1(_11019_),
    .Y(_11033_),
    .A2(_11022_));
 sg13g2_nand4_1 _17863_ (.B(_11013_),
    .C(_11018_),
    .A(_11009_),
    .Y(_11034_),
    .D(_11033_));
 sg13g2_nand2_1 _17864_ (.Y(_11035_),
    .A(_10038_),
    .B(_10892_));
 sg13g2_o21ai_1 _17865_ (.B1(_11035_),
    .Y(_11036_),
    .A1(net568),
    .A2(_11034_));
 sg13g2_buf_2 _17866_ (.A(_11036_),
    .X(_11037_));
 sg13g2_nand2b_1 _17867_ (.Y(_11038_),
    .B(net1068),
    .A_N(_09332_));
 sg13g2_or3_1 _17868_ (.A(_10954_),
    .B(_11037_),
    .C(_11038_),
    .X(_11039_));
 sg13g2_nor2_1 _17869_ (.A(_09332_),
    .B(net1068),
    .Y(_11040_));
 sg13g2_nand2_1 _17870_ (.Y(_11041_),
    .A(_10998_),
    .B(_11040_));
 sg13g2_nand4_1 _17871_ (.B(_10999_),
    .C(_11039_),
    .A(_10952_),
    .Y(_11042_),
    .D(_11041_));
 sg13g2_buf_1 _17872_ (.A(\cpu.br ),
    .X(_11043_));
 sg13g2_a21o_1 _17873_ (.A2(_11019_),
    .A1(_10894_),
    .B1(_00257_),
    .X(_11044_));
 sg13g2_nor4_1 _17874_ (.A(_09208_),
    .B(_09174_),
    .C(_09205_),
    .D(_11044_),
    .Y(_11045_));
 sg13g2_and3_1 _17875_ (.X(_11046_),
    .A(_08383_),
    .B(_08386_),
    .C(_11045_));
 sg13g2_nand3_1 _17876_ (.B(_08467_),
    .C(_11046_),
    .A(_08423_),
    .Y(_11047_));
 sg13g2_buf_8 _17877_ (.A(_11047_),
    .X(_11048_));
 sg13g2_nand2_1 _17878_ (.Y(_11049_),
    .A(net1117),
    .B(_11048_));
 sg13g2_buf_8 _17879_ (.A(_11049_),
    .X(_11050_));
 sg13g2_mux2_1 _17880_ (.A0(_10880_),
    .A1(_11042_),
    .S(_11050_),
    .X(_11051_));
 sg13g2_inv_1 _17881_ (.Y(_11052_),
    .A(net1117));
 sg13g2_buf_1 _17882_ (.A(_11052_),
    .X(_11053_));
 sg13g2_nor2_1 _17883_ (.A(_08348_),
    .B(net890),
    .Y(_11054_));
 sg13g2_or3_1 _17884_ (.A(_09208_),
    .B(_09174_),
    .C(_09205_),
    .X(_11055_));
 sg13g2_inv_2 _17885_ (.Y(_11056_),
    .A(net1145));
 sg13g2_a21oi_1 _17886_ (.A1(_11056_),
    .A2(_10892_),
    .Y(_11057_),
    .B1(net1117));
 sg13g2_mux2_1 _17887_ (.A0(\cpu.ex.r_9[0] ),
    .A1(\cpu.ex.r_11[0] ),
    .S(net1118),
    .X(_11058_));
 sg13g2_a221oi_1 _17888_ (.B2(_10901_),
    .C1(net1038),
    .B1(_11058_),
    .A1(\cpu.ex.r_8[0] ),
    .Y(_11059_),
    .A2(_10982_));
 sg13g2_mux2_1 _17889_ (.A0(\cpu.ex.r_12[0] ),
    .A1(\cpu.ex.r_14[0] ),
    .S(net1118),
    .X(_11060_));
 sg13g2_a221oi_1 _17890_ (.B2(net764),
    .C1(_10919_),
    .B1(_11060_),
    .A1(\cpu.ex.r_13[0] ),
    .Y(_11061_),
    .A2(_10910_));
 sg13g2_nor3_1 _17891_ (.A(_10924_),
    .B(_11059_),
    .C(_11061_),
    .Y(_11062_));
 sg13g2_mux2_1 _17892_ (.A0(_09160_),
    .A1(\cpu.ex.r_stmp[0] ),
    .S(_10895_),
    .X(_11063_));
 sg13g2_a22oi_1 _17893_ (.Y(_11064_),
    .B1(_11063_),
    .B2(net764),
    .A2(_10928_),
    .A1(\cpu.ex.r_mult[16] ));
 sg13g2_nor2b_1 _17894_ (.A(_11064_),
    .B_N(_10942_),
    .Y(_11065_));
 sg13g2_and2_1 _17895_ (.A(net1039),
    .B(_10886_),
    .X(_11066_));
 sg13g2_a22oi_1 _17896_ (.Y(_11067_),
    .B1(_11066_),
    .B2(\cpu.ex.r_15[0] ),
    .A2(_11019_),
    .A1(\cpu.ex.r_10[0] ));
 sg13g2_nand3_1 _17897_ (.B(_10928_),
    .C(_10930_),
    .A(_10657_),
    .Y(_11068_));
 sg13g2_o21ai_1 _17898_ (.B1(_11068_),
    .Y(_11069_),
    .A1(_11016_),
    .A2(_11067_));
 sg13g2_or4_1 _17899_ (.A(_10892_),
    .B(_11062_),
    .C(_11065_),
    .D(_11069_),
    .X(_11070_));
 sg13g2_buf_1 _17900_ (.A(_11070_),
    .X(_11071_));
 sg13g2_a22oi_1 _17901_ (.Y(_11072_),
    .B1(_11057_),
    .B2(_11071_),
    .A2(_11055_),
    .A1(_11054_));
 sg13g2_nand2_1 _17902_ (.Y(_11073_),
    .A(_11056_),
    .B(_10892_));
 sg13g2_nand3_1 _17903_ (.B(_11071_),
    .C(_11073_),
    .A(_11045_),
    .Y(_11074_));
 sg13g2_and2_1 _17904_ (.A(_11072_),
    .B(_11074_),
    .X(_11075_));
 sg13g2_a21oi_1 _17905_ (.A1(_11071_),
    .A2(_11057_),
    .Y(_11076_),
    .B1(_11054_));
 sg13g2_mux2_1 _17906_ (.A0(_11075_),
    .A1(_11076_),
    .S(_08469_),
    .X(_11077_));
 sg13g2_buf_8 _17907_ (.A(_11077_),
    .X(_11078_));
 sg13g2_nor3_1 _17908_ (.A(_09347_),
    .B(\cpu.ex.c_mult_off[0] ),
    .C(_11078_),
    .Y(_11079_));
 sg13g2_xnor2_1 _17909_ (.Y(_11080_),
    .A(_09348_),
    .B(_11040_));
 sg13g2_and2_1 _17910_ (.A(_09342_),
    .B(_11080_),
    .X(_11081_));
 sg13g2_buf_1 _17911_ (.A(_11081_),
    .X(_11082_));
 sg13g2_inv_1 _17912_ (.Y(\cpu.ex.c_mult_off[2] ),
    .A(_11082_));
 sg13g2_nor3_1 _17913_ (.A(_09332_),
    .B(net1068),
    .C(_09348_),
    .Y(_11083_));
 sg13g2_xnor2_1 _17914_ (.Y(_11084_),
    .A(_09349_),
    .B(_11083_));
 sg13g2_nand2_1 _17915_ (.Y(\cpu.ex.c_mult_off[3] ),
    .A(_09342_),
    .B(_11084_));
 sg13g2_nor2_1 _17916_ (.A(\cpu.ex.c_mult_off[2] ),
    .B(\cpu.ex.c_mult_off[3] ),
    .Y(_11085_));
 sg13g2_o21ai_1 _17917_ (.B1(_11085_),
    .Y(_11086_),
    .A1(_11051_),
    .A2(_11079_));
 sg13g2_inv_1 _17918_ (.Y(_11087_),
    .A(_00184_));
 sg13g2_inv_1 _17919_ (.Y(_11088_),
    .A(_00186_));
 sg13g2_xor2_1 _17920_ (.B(_09346_),
    .A(_09332_),
    .X(_11089_));
 sg13g2_and2_1 _17921_ (.A(_09342_),
    .B(_11089_),
    .X(_11090_));
 sg13g2_buf_1 _17922_ (.A(_11090_),
    .X(_11091_));
 sg13g2_mux2_1 _17923_ (.A0(_11087_),
    .A1(_11088_),
    .S(net511),
    .X(_11092_));
 sg13g2_inv_1 _17924_ (.Y(_11093_),
    .A(_00185_));
 sg13g2_nor2_1 _17925_ (.A(_11093_),
    .B(net511),
    .Y(_11094_));
 sg13g2_a21oi_1 _17926_ (.A1(_10296_),
    .A2(net511),
    .Y(_11095_),
    .B1(_11094_));
 sg13g2_nor3_2 _17927_ (.A(net899),
    .B(net891),
    .C(net1038),
    .Y(_11096_));
 sg13g2_a22oi_1 _17928_ (.Y(_11097_),
    .B1(_11096_),
    .B2(\cpu.ex.r_8[15] ),
    .A2(_10923_),
    .A1(\cpu.ex.r_15[15] ));
 sg13g2_buf_8 _17929_ (.A(net766),
    .X(_11098_));
 sg13g2_nand2b_1 _17930_ (.Y(_11099_),
    .B(net675),
    .A_N(_11097_));
 sg13g2_and2_1 _17931_ (.A(net893),
    .B(_10976_),
    .X(_11100_));
 sg13g2_buf_1 _17932_ (.A(_11100_),
    .X(_11101_));
 sg13g2_mux2_1 _17933_ (.A0(\cpu.ex.r_12[15] ),
    .A1(\cpu.ex.r_13[15] ),
    .S(net769),
    .X(_11102_));
 sg13g2_nor2b_2 _17934_ (.A(net893),
    .B_N(net894),
    .Y(_11103_));
 sg13g2_and2_1 _17935_ (.A(_10924_),
    .B(_11103_),
    .X(_11104_));
 sg13g2_mux2_1 _17936_ (.A0(_10440_),
    .A1(\cpu.ex.r_epc[15] ),
    .S(net769),
    .X(_11105_));
 sg13g2_a22oi_1 _17937_ (.Y(_11106_),
    .B1(_11104_),
    .B2(_11105_),
    .A2(_11102_),
    .A1(_11101_));
 sg13g2_nor2_2 _17938_ (.A(_10919_),
    .B(_10907_),
    .Y(_11107_));
 sg13g2_mux2_1 _17939_ (.A0(\cpu.ex.r_stmp[15] ),
    .A1(\cpu.ex.r_14[15] ),
    .S(net766),
    .X(_11108_));
 sg13g2_mux2_1 _17940_ (.A0(\cpu.ex.r_10[15] ),
    .A1(\cpu.ex.r_11[15] ),
    .S(net769),
    .X(_11109_));
 sg13g2_a22oi_1 _17941_ (.Y(_11110_),
    .B1(_11109_),
    .B2(_11017_),
    .A2(_11108_),
    .A1(_11107_));
 sg13g2_a22oi_1 _17942_ (.Y(_11111_),
    .B1(_10964_),
    .B2(\cpu.ex.r_9[15] ),
    .A2(_10942_),
    .A1(_10443_));
 sg13g2_nor2b_1 _17943_ (.A(_11111_),
    .B_N(net768),
    .Y(_11112_));
 sg13g2_nor2_2 _17944_ (.A(_11001_),
    .B(_10915_),
    .Y(_11113_));
 sg13g2_a22oi_1 _17945_ (.Y(_11114_),
    .B1(_11024_),
    .B2(\cpu.ex.r_mult[31] ),
    .A2(_11113_),
    .A1(\cpu.ex.r_lr[15] ));
 sg13g2_nor2_1 _17946_ (.A(_11027_),
    .B(_11114_),
    .Y(_11115_));
 sg13g2_nor2_1 _17947_ (.A(_11112_),
    .B(_11115_),
    .Y(_11116_));
 sg13g2_and4_1 _17948_ (.A(_11099_),
    .B(_11106_),
    .C(_11110_),
    .D(_11116_),
    .X(_11117_));
 sg13g2_mux2_1 _17949_ (.A0(net797),
    .A1(_11117_),
    .S(_10956_),
    .X(_11118_));
 sg13g2_buf_1 _17950_ (.A(_11118_),
    .X(_11119_));
 sg13g2_and2_1 _17951_ (.A(_10935_),
    .B(_10942_),
    .X(_11120_));
 sg13g2_mux2_1 _17952_ (.A0(\cpu.ex.r_12[13] ),
    .A1(\cpu.ex.r_13[13] ),
    .S(net769),
    .X(_11121_));
 sg13g2_a22oi_1 _17953_ (.Y(_11122_),
    .B1(_11101_),
    .B2(_11121_),
    .A2(_11120_),
    .A1(\cpu.ex.r_stmp[13] ));
 sg13g2_mux2_1 _17954_ (.A0(\cpu.ex.r_9[13] ),
    .A1(\cpu.ex.r_11[13] ),
    .S(net891),
    .X(_11123_));
 sg13g2_mux2_1 _17955_ (.A0(_10266_),
    .A1(_10263_),
    .S(net894),
    .X(_11124_));
 sg13g2_a22oi_1 _17956_ (.Y(_11125_),
    .B1(_11124_),
    .B2(net765),
    .A2(_11123_),
    .A1(net762));
 sg13g2_nand2b_1 _17957_ (.Y(_11126_),
    .B(net677),
    .A_N(_11125_));
 sg13g2_a22oi_1 _17958_ (.Y(_11127_),
    .B1(_11096_),
    .B2(\cpu.ex.r_8[13] ),
    .A2(_10923_),
    .A1(_10256_));
 sg13g2_nand2b_1 _17959_ (.Y(_11128_),
    .B(net675),
    .A_N(_11127_));
 sg13g2_nor2_1 _17960_ (.A(net897),
    .B(_11027_),
    .Y(_11129_));
 sg13g2_mux2_1 _17961_ (.A0(\cpu.ex.r_lr[13] ),
    .A1(\cpu.ex.r_epc[13] ),
    .S(net894),
    .X(_11130_));
 sg13g2_mux2_1 _17962_ (.A0(\cpu.ex.r_sp[13] ),
    .A1(\cpu.ex.r_10[13] ),
    .S(net898),
    .X(_11131_));
 sg13g2_and3_1 _17963_ (.X(_11132_),
    .A(net892),
    .B(_10970_),
    .C(\cpu.ex.r_14[13] ));
 sg13g2_a21o_1 _17964_ (.A2(_11131_),
    .A1(_10919_),
    .B1(_11132_),
    .X(_11133_));
 sg13g2_a22oi_1 _17965_ (.Y(_11134_),
    .B1(_11133_),
    .B2(_10987_),
    .A2(_11130_),
    .A1(_11129_));
 sg13g2_nand4_1 _17966_ (.B(_11126_),
    .C(_11128_),
    .A(_11122_),
    .Y(_11135_),
    .D(_11134_));
 sg13g2_mux2_1 _17967_ (.A0(_09382_),
    .A1(_11135_),
    .S(_10956_),
    .X(_11136_));
 sg13g2_buf_1 _17968_ (.A(_11136_),
    .X(_11137_));
 sg13g2_nand2_1 _17969_ (.Y(_11138_),
    .A(_11091_),
    .B(_11137_));
 sg13g2_o21ai_1 _17970_ (.B1(_11138_),
    .Y(_11139_),
    .A1(net511),
    .A2(_11119_));
 sg13g2_and3_1 _17971_ (.X(_11140_),
    .A(net892),
    .B(\cpu.ex.r_13[14] ),
    .C(net768));
 sg13g2_a21o_1 _17972_ (.A2(_10908_),
    .A1(\cpu.ex.r_stmp[14] ),
    .B1(_11140_),
    .X(_11141_));
 sg13g2_inv_1 _17973_ (.Y(_11142_),
    .A(\cpu.ex.r_11[14] ));
 sg13g2_nand2_1 _17974_ (.Y(_11143_),
    .A(_10919_),
    .B(_10898_));
 sg13g2_nand3_1 _17975_ (.B(_10474_),
    .C(_10942_),
    .A(net895),
    .Y(_11144_));
 sg13g2_o21ai_1 _17976_ (.B1(_11144_),
    .Y(_11145_),
    .A1(_11142_),
    .A2(_11143_));
 sg13g2_a22oi_1 _17977_ (.Y(_11146_),
    .B1(_11096_),
    .B2(\cpu.ex.r_8[14] ),
    .A2(_10923_),
    .A1(_10459_));
 sg13g2_nor2_1 _17978_ (.A(net759),
    .B(_11146_),
    .Y(_11147_));
 sg13g2_a221oi_1 _17979_ (.B2(net677),
    .C1(_11147_),
    .B1(_11145_),
    .A1(net760),
    .Y(_11148_),
    .A2(_11141_));
 sg13g2_nor2b_1 _17980_ (.A(net899),
    .B_N(net1040),
    .Y(_11149_));
 sg13g2_buf_2 _17981_ (.A(_11149_),
    .X(_11150_));
 sg13g2_nor2_1 _17982_ (.A(_10959_),
    .B(net892),
    .Y(_11151_));
 sg13g2_a22oi_1 _17983_ (.Y(_11152_),
    .B1(_11151_),
    .B2(\cpu.ex.r_mult[30] ),
    .A2(_11150_),
    .A1(\cpu.ex.r_14[14] ));
 sg13g2_nand2b_1 _17984_ (.Y(_11153_),
    .B(_11024_),
    .A_N(_11152_));
 sg13g2_nand2_1 _17985_ (.Y(_11154_),
    .A(net892),
    .B(\cpu.ex.r_9[14] ));
 sg13g2_o21ai_1 _17986_ (.B1(_11154_),
    .Y(_11155_),
    .A1(net892),
    .A2(_10471_));
 sg13g2_a22oi_1 _17987_ (.Y(_11156_),
    .B1(_11011_),
    .B2(_11155_),
    .A2(_11014_),
    .A1(\cpu.ex.r_12[14] ));
 sg13g2_nor2_1 _17988_ (.A(net893),
    .B(_10907_),
    .Y(_11157_));
 sg13g2_mux2_1 _17989_ (.A0(_10456_),
    .A1(\cpu.ex.r_10[14] ),
    .S(_10988_),
    .X(_11158_));
 sg13g2_a22oi_1 _17990_ (.Y(_11159_),
    .B1(_11157_),
    .B2(_11158_),
    .A2(_10932_),
    .A1(\cpu.ex.r_epc[14] ));
 sg13g2_and2_1 _17991_ (.A(_11156_),
    .B(_11159_),
    .X(_11160_));
 sg13g2_nand4_1 _17992_ (.B(_11148_),
    .C(_11153_),
    .A(_10956_),
    .Y(_11161_),
    .D(_11160_));
 sg13g2_nand2b_1 _17993_ (.Y(_11162_),
    .B(_10893_),
    .A_N(net945));
 sg13g2_and2_1 _17994_ (.A(_11161_),
    .B(_11162_),
    .X(_11163_));
 sg13g2_buf_1 _17995_ (.A(_11163_),
    .X(_11164_));
 sg13g2_a22oi_1 _17996_ (.Y(_11165_),
    .B1(_11011_),
    .B2(\cpu.ex.r_lr[12] ),
    .A2(_11107_),
    .A1(\cpu.ex.r_stmp[12] ));
 sg13g2_a221oi_1 _17997_ (.B2(\cpu.ex.r_9[12] ),
    .C1(net759),
    .B1(_11011_),
    .A1(\cpu.ex.r_14[12] ),
    .Y(_11166_),
    .A2(_11107_));
 sg13g2_a21oi_1 _17998_ (.A1(net759),
    .A2(_11165_),
    .Y(_11167_),
    .B1(_11166_));
 sg13g2_mux2_1 _17999_ (.A0(\cpu.ex.r_8[12] ),
    .A1(\cpu.ex.r_10[12] ),
    .S(net894),
    .X(_11168_));
 sg13g2_a22oi_1 _18000_ (.Y(_11169_),
    .B1(_11168_),
    .B2(net764),
    .A2(_10928_),
    .A1(\cpu.ex.r_11[12] ));
 sg13g2_nor2b_1 _18001_ (.A(_11169_),
    .B_N(net762),
    .Y(_11170_));
 sg13g2_nor2_1 _18002_ (.A(net763),
    .B(net896),
    .Y(_11171_));
 sg13g2_a22oi_1 _18003_ (.Y(_11172_),
    .B1(_11103_),
    .B2(\cpu.ex.r_epc[12] ),
    .A2(_11171_),
    .A1(_10313_));
 sg13g2_and2_1 _18004_ (.A(_10910_),
    .B(_10980_),
    .X(_11173_));
 sg13g2_buf_1 _18005_ (.A(_11173_),
    .X(_11174_));
 sg13g2_nand2b_1 _18006_ (.Y(_11175_),
    .B(net766),
    .A_N(_00254_));
 sg13g2_o21ai_1 _18007_ (.B1(_11175_),
    .Y(_11176_),
    .A1(net766),
    .A2(_10323_));
 sg13g2_a22oi_1 _18008_ (.Y(_11177_),
    .B1(_11176_),
    .B2(_10923_),
    .A2(_11174_),
    .A1(\cpu.ex.r_13[12] ));
 sg13g2_o21ai_1 _18009_ (.B1(_11177_),
    .Y(_11178_),
    .A1(_11027_),
    .A2(_11172_));
 sg13g2_nand2_1 _18010_ (.Y(_11179_),
    .A(\cpu.ex.r_12[12] ),
    .B(_11101_));
 sg13g2_nand3_1 _18011_ (.B(_10329_),
    .C(_10930_),
    .A(net763),
    .Y(_11180_));
 sg13g2_a21oi_1 _18012_ (.A1(_11179_),
    .A2(_11180_),
    .Y(_11181_),
    .B1(net677));
 sg13g2_nor4_2 _18013_ (.A(_11167_),
    .B(_11170_),
    .C(_11178_),
    .Y(_11182_),
    .D(_11181_));
 sg13g2_nor2_1 _18014_ (.A(net701),
    .B(net567),
    .Y(_11183_));
 sg13g2_a21oi_2 _18015_ (.B1(_11183_),
    .Y(_11184_),
    .A2(_11182_),
    .A1(net567));
 sg13g2_mux2_1 _18016_ (.A0(_11164_),
    .A1(_11184_),
    .S(_11091_),
    .X(_11185_));
 sg13g2_buf_8 _18017_ (.A(_11050_),
    .X(_11186_));
 sg13g2_mux4_1 _18018_ (.S0(_09344_),
    .A0(_11092_),
    .A1(_11095_),
    .A2(_11139_),
    .A3(_11185_),
    .S1(net241),
    .X(_11187_));
 sg13g2_nand3_1 _18019_ (.B(\cpu.ex.c_mult_off[3] ),
    .C(_11187_),
    .A(\cpu.ex.c_mult_off[2] ),
    .Y(_11188_));
 sg13g2_inv_1 _18020_ (.Y(_11189_),
    .A(\cpu.ex.r_stmp[11] ));
 sg13g2_nor3_1 _18021_ (.A(net675),
    .B(_11189_),
    .C(_10907_),
    .Y(_11190_));
 sg13g2_a21o_1 _18022_ (.A2(_10913_),
    .A1(\cpu.ex.r_13[11] ),
    .B1(_11190_),
    .X(_11191_));
 sg13g2_mux2_1 _18023_ (.A0(\cpu.ex.r_12[11] ),
    .A1(\cpu.ex.r_14[11] ),
    .S(net763),
    .X(_11192_));
 sg13g2_a22oi_1 _18024_ (.Y(_11193_),
    .B1(_11192_),
    .B2(net764),
    .A2(_10928_),
    .A1(_10372_));
 sg13g2_mux2_1 _18025_ (.A0(\cpu.ex.r_9[11] ),
    .A1(\cpu.ex.r_11[11] ),
    .S(net894),
    .X(_11194_));
 sg13g2_a221oi_1 _18026_ (.B2(net677),
    .C1(net767),
    .B1(_11194_),
    .A1(\cpu.ex.r_8[11] ),
    .Y(_11195_),
    .A2(net761));
 sg13g2_a21oi_1 _18027_ (.A1(net767),
    .A2(_11193_),
    .Y(_11196_),
    .B1(_11195_));
 sg13g2_a22oi_1 _18028_ (.Y(_11197_),
    .B1(_11024_),
    .B2(\cpu.ex.r_mult[27] ),
    .A2(_11113_),
    .A1(\cpu.ex.r_lr[11] ));
 sg13g2_mux2_1 _18029_ (.A0(_10359_),
    .A1(\cpu.ex.r_10[11] ),
    .S(net766),
    .X(_11198_));
 sg13g2_a22oi_1 _18030_ (.Y(_11199_),
    .B1(_11157_),
    .B2(_11198_),
    .A2(_10932_),
    .A1(\cpu.ex.r_epc[11] ));
 sg13g2_o21ai_1 _18031_ (.B1(_11199_),
    .Y(_11200_),
    .A1(_11027_),
    .A2(_11197_));
 sg13g2_a221oi_1 _18032_ (.B2(net675),
    .C1(_11200_),
    .B1(_11196_),
    .A1(net767),
    .Y(_11201_),
    .A2(_11191_));
 sg13g2_nor2_1 _18033_ (.A(net1122),
    .B(net567),
    .Y(_11202_));
 sg13g2_a21oi_1 _18034_ (.A1(_10957_),
    .A2(_11201_),
    .Y(_11203_),
    .B1(_11202_));
 sg13g2_a221oi_1 _18035_ (.B2(\cpu.ex.r_mult[25] ),
    .C1(net675),
    .B1(_11024_),
    .A1(\cpu.ex.r_lr[9] ),
    .Y(_11204_),
    .A2(_11113_));
 sg13g2_inv_1 _18036_ (.Y(_11205_),
    .A(_00251_));
 sg13g2_a221oi_1 _18037_ (.B2(_11205_),
    .C1(net759),
    .B1(_11024_),
    .A1(\cpu.ex.r_9[9] ),
    .Y(_11206_),
    .A2(_11113_));
 sg13g2_or3_1 _18038_ (.A(_10959_),
    .B(_11204_),
    .C(_11206_),
    .X(_11207_));
 sg13g2_mux2_1 _18039_ (.A0(\cpu.ex.r_stmp[9] ),
    .A1(\cpu.ex.r_14[9] ),
    .S(net675),
    .X(_11208_));
 sg13g2_mux2_1 _18040_ (.A0(\cpu.ex.r_epc[9] ),
    .A1(\cpu.ex.r_11[9] ),
    .S(net675),
    .X(_11209_));
 sg13g2_nor2_1 _18041_ (.A(net767),
    .B(_10981_),
    .Y(_11210_));
 sg13g2_a22oi_1 _18042_ (.Y(_11211_),
    .B1(_11209_),
    .B2(_11210_),
    .A2(_11208_),
    .A1(_11107_));
 sg13g2_nand3_1 _18043_ (.B(_10930_),
    .C(_10987_),
    .A(_10530_),
    .Y(_11212_));
 sg13g2_nand2_1 _18044_ (.Y(_11213_),
    .A(_10986_),
    .B(\cpu.ex.r_12[9] ));
 sg13g2_nand3b_1 _18045_ (.B(\cpu.ex.r_10[9] ),
    .C(net763),
    .Y(_11214_),
    .A_N(_10986_));
 sg13g2_o21ai_1 _18046_ (.B1(_11214_),
    .Y(_11215_),
    .A1(net763),
    .A2(_11213_));
 sg13g2_and3_1 _18047_ (.X(_11216_),
    .A(\cpu.ex.r_8[9] ),
    .B(_10965_),
    .C(_10983_));
 sg13g2_a221oi_1 _18048_ (.B2(_11150_),
    .C1(_11216_),
    .B1(_11215_),
    .A1(\cpu.ex.r_13[9] ),
    .Y(_11217_),
    .A2(_11174_));
 sg13g2_nand4_1 _18049_ (.B(_11211_),
    .C(_11212_),
    .A(_11207_),
    .Y(_11218_),
    .D(_11217_));
 sg13g2_mux2_1 _18050_ (.A0(_10524_),
    .A1(_11218_),
    .S(net567),
    .X(_11219_));
 sg13g2_mux4_1 _18051_ (.S0(net511),
    .A0(_10385_),
    .A1(_10548_),
    .A2(_11203_),
    .A3(_11219_),
    .S1(_11050_),
    .X(_11220_));
 sg13g2_nand4_1 _18052_ (.B(_11082_),
    .C(\cpu.ex.c_mult_off[3] ),
    .A(\cpu.ex.c_mult_off[0] ),
    .Y(_11221_),
    .D(_11220_));
 sg13g2_nand3_1 _18053_ (.B(_11082_),
    .C(\cpu.ex.c_mult_off[3] ),
    .A(_09344_),
    .Y(_11222_));
 sg13g2_nor2_1 _18054_ (.A(net511),
    .B(_11222_),
    .Y(_11223_));
 sg13g2_inv_1 _18055_ (.Y(_11224_),
    .A(_10392_));
 sg13g2_buf_1 _18056_ (.A(_11224_),
    .X(_11225_));
 sg13g2_a22oi_1 _18057_ (.Y(_11226_),
    .B1(_10913_),
    .B2(\cpu.ex.r_9[10] ),
    .A2(_10908_),
    .A1(_10403_));
 sg13g2_a22oi_1 _18058_ (.Y(_11227_),
    .B1(_11096_),
    .B2(\cpu.ex.r_8[10] ),
    .A2(_10923_),
    .A1(_10399_));
 sg13g2_nor2_1 _18059_ (.A(net759),
    .B(_11227_),
    .Y(_11228_));
 sg13g2_a221oi_1 _18060_ (.B2(\cpu.ex.r_13[10] ),
    .C1(_11228_),
    .B1(_11174_),
    .A1(\cpu.ex.r_epc[10] ),
    .Y(_11229_),
    .A2(_10932_));
 sg13g2_o21ai_1 _18061_ (.B1(_11229_),
    .Y(_11230_),
    .A1(net767),
    .A2(_11226_));
 sg13g2_inv_1 _18062_ (.Y(_11231_),
    .A(_10410_));
 sg13g2_nor2_1 _18063_ (.A(net896),
    .B(_11231_),
    .Y(_11232_));
 sg13g2_nand2_1 _18064_ (.Y(_11233_),
    .A(net897),
    .B(\cpu.ex.r_14[10] ));
 sg13g2_o21ai_1 _18065_ (.B1(_11233_),
    .Y(_11234_),
    .A1(net760),
    .A2(_10413_));
 sg13g2_a22oi_1 _18066_ (.Y(_11235_),
    .B1(_11234_),
    .B2(_11150_),
    .A2(_11232_),
    .A1(_11151_));
 sg13g2_nor2b_1 _18067_ (.A(net677),
    .B_N(\cpu.ex.r_stmp[10] ),
    .Y(_11236_));
 sg13g2_nor2b_1 _18068_ (.A(net760),
    .B_N(\cpu.ex.r_11[10] ),
    .Y(_11237_));
 sg13g2_a221oi_1 _18069_ (.B2(_11007_),
    .C1(net895),
    .B1(_11237_),
    .A1(net765),
    .Y(_11238_),
    .A2(_11236_));
 sg13g2_and2_1 _18070_ (.A(net760),
    .B(_11150_),
    .X(_11239_));
 sg13g2_a221oi_1 _18071_ (.B2(\cpu.ex.r_12[10] ),
    .C1(net763),
    .B1(_11239_),
    .A1(\cpu.ex.r_lr[10] ),
    .Y(_11240_),
    .A2(_11129_));
 sg13g2_a21oi_1 _18072_ (.A1(_11235_),
    .A2(_11238_),
    .Y(_11241_),
    .B1(_11240_));
 sg13g2_nor3_1 _18073_ (.A(net568),
    .B(_11230_),
    .C(_11241_),
    .Y(_11242_));
 sg13g2_a21oi_1 _18074_ (.A1(_11225_),
    .A2(net568),
    .Y(_11243_),
    .B1(_11242_));
 sg13g2_mux2_1 _18075_ (.A0(_10389_),
    .A1(_11243_),
    .S(_11050_),
    .X(_11244_));
 sg13g2_buf_8 _18076_ (.A(_11244_),
    .X(_11245_));
 sg13g2_inv_1 _18077_ (.Y(_11246_),
    .A(_09349_));
 sg13g2_nand2_1 _18078_ (.Y(_11247_),
    .A(_09348_),
    .B(_11246_));
 sg13g2_or2_1 _18079_ (.X(_11248_),
    .B(_11247_),
    .A(\cpu.ex.c_mult_off[0] ));
 sg13g2_buf_1 _18080_ (.A(_11248_),
    .X(_11249_));
 sg13g2_inv_4 _18081_ (.A(net511),
    .Y(\cpu.ex.c_mult_off[1] ));
 sg13g2_nor2_1 _18082_ (.A(_08498_),
    .B(\cpu.ex.c_mult_off[1] ),
    .Y(_11250_));
 sg13g2_a21oi_1 _18083_ (.A1(_10816_),
    .A2(\cpu.ex.c_mult_off[1] ),
    .Y(_11251_),
    .B1(_11250_));
 sg13g2_nand3_1 _18084_ (.B(_09342_),
    .C(_11083_),
    .A(_09349_),
    .Y(_11252_));
 sg13g2_inv_1 _18085_ (.Y(_11253_),
    .A(_10733_));
 sg13g2_nand2b_1 _18086_ (.Y(_11254_),
    .B(_11253_),
    .A_N(_11252_));
 sg13g2_o21ai_1 _18087_ (.B1(_11254_),
    .Y(_11255_),
    .A1(_11249_),
    .A2(_11251_));
 sg13g2_nor3_1 _18088_ (.A(_10487_),
    .B(\cpu.ex.c_mult_off[1] ),
    .C(_11222_),
    .Y(_11256_));
 sg13g2_nor3_1 _18089_ (.A(_10954_),
    .B(_11038_),
    .C(_11247_),
    .Y(_11257_));
 sg13g2_and2_1 _18090_ (.A(_10740_),
    .B(_11257_),
    .X(_11258_));
 sg13g2_or4_1 _18091_ (.A(_11050_),
    .B(_11255_),
    .C(_11256_),
    .D(_11258_),
    .X(_11259_));
 sg13g2_nand3b_1 _18092_ (.B(_10905_),
    .C(\cpu.ex.r_14[6] ),
    .Y(_11260_),
    .A_N(net899));
 sg13g2_nand3b_1 _18093_ (.B(_10810_),
    .C(_10902_),
    .Y(_11261_),
    .A_N(_10905_));
 sg13g2_a21o_1 _18094_ (.A2(_11261_),
    .A1(_11260_),
    .B1(_10919_),
    .X(_11262_));
 sg13g2_mux2_1 _18095_ (.A0(_10685_),
    .A1(\cpu.ex.r_10[6] ),
    .S(net1040),
    .X(_11263_));
 sg13g2_nor2b_1 _18096_ (.A(_00248_),
    .B_N(net893),
    .Y(_11264_));
 sg13g2_a22oi_1 _18097_ (.Y(_11265_),
    .B1(_11264_),
    .B2(_11007_),
    .A2(_11263_),
    .A1(_11019_));
 sg13g2_a21oi_1 _18098_ (.A1(_11262_),
    .A2(_11265_),
    .Y(_11266_),
    .B1(net895));
 sg13g2_mux4_1 _18099_ (.S0(_11001_),
    .A0(\cpu.ex.r_lr[6] ),
    .A1(\cpu.ex.r_epc[6] ),
    .A2(\cpu.ex.r_9[6] ),
    .A3(\cpu.ex.r_11[6] ),
    .S1(net892),
    .X(_11267_));
 sg13g2_nor2b_1 _18100_ (.A(net893),
    .B_N(net769),
    .Y(_11268_));
 sg13g2_nand2_1 _18101_ (.Y(_11269_),
    .A(_11267_),
    .B(_11268_));
 sg13g2_nand3_1 _18102_ (.B(net676),
    .C(net765),
    .A(\cpu.ex.r_stmp[6] ),
    .Y(_11270_));
 sg13g2_nand3_1 _18103_ (.B(_10964_),
    .C(net761),
    .A(\cpu.ex.r_8[6] ),
    .Y(_11271_));
 sg13g2_mux2_1 _18104_ (.A0(\cpu.ex.r_12[6] ),
    .A1(\cpu.ex.r_13[6] ),
    .S(net899),
    .X(_11272_));
 sg13g2_nand3_1 _18105_ (.B(_10976_),
    .C(_11272_),
    .A(net897),
    .Y(_11273_));
 sg13g2_nand4_1 _18106_ (.B(_11270_),
    .C(_11271_),
    .A(_11269_),
    .Y(_11274_),
    .D(_11273_));
 sg13g2_or3_1 _18107_ (.A(_10892_),
    .B(_11266_),
    .C(_11274_),
    .X(_11275_));
 sg13g2_o21ai_1 _18108_ (.B1(_11275_),
    .Y(_11276_),
    .A1(_09220_),
    .A2(_10956_));
 sg13g2_buf_1 _18109_ (.A(_11276_),
    .X(_11277_));
 sg13g2_or3_1 _18110_ (.A(net511),
    .B(_11249_),
    .C(_11277_),
    .X(_11278_));
 sg13g2_a22oi_1 _18111_ (.Y(_11279_),
    .B1(net768),
    .B2(\cpu.ex.r_9[4] ),
    .A2(_10935_),
    .A1(\cpu.ex.r_10[4] ));
 sg13g2_nand2b_1 _18112_ (.Y(_11280_),
    .B(net762),
    .A_N(_11279_));
 sg13g2_a22oi_1 _18113_ (.Y(_11281_),
    .B1(_11007_),
    .B2(\cpu.ex.r_11[4] ),
    .A2(_11000_),
    .A1(_10768_));
 sg13g2_nand2b_1 _18114_ (.Y(_11282_),
    .B(_11103_),
    .A_N(_11281_));
 sg13g2_mux2_1 _18115_ (.A0(\cpu.ex.r_lr[4] ),
    .A1(\cpu.ex.r_epc[4] ),
    .S(net894),
    .X(_11283_));
 sg13g2_mux2_1 _18116_ (.A0(\cpu.ex.r_8[4] ),
    .A1(\cpu.ex.r_12[4] ),
    .S(_10915_),
    .X(_11284_));
 sg13g2_and3_1 _18117_ (.X(_11285_),
    .A(_10933_),
    .B(_10983_),
    .C(_11284_));
 sg13g2_a221oi_1 _18118_ (.B2(_11129_),
    .C1(_11285_),
    .B1(_11283_),
    .A1(\cpu.ex.r_13[4] ),
    .Y(_11286_),
    .A2(_11174_));
 sg13g2_nand3_1 _18119_ (.B(_11282_),
    .C(_11286_),
    .A(_11280_),
    .Y(_11287_));
 sg13g2_nor3_1 _18120_ (.A(_10924_),
    .B(_00246_),
    .C(_10981_),
    .Y(_11288_));
 sg13g2_and3_1 _18121_ (.X(_11289_),
    .A(_08347_),
    .B(net764),
    .C(_10894_));
 sg13g2_o21ai_1 _18122_ (.B1(net760),
    .Y(_11290_),
    .A1(_11288_),
    .A2(_11289_));
 sg13g2_and2_1 _18123_ (.A(_10928_),
    .B(_10942_),
    .X(_11291_));
 sg13g2_mux2_1 _18124_ (.A0(\cpu.ex.r_stmp[4] ),
    .A1(\cpu.ex.r_14[4] ),
    .S(net892),
    .X(_11292_));
 sg13g2_a22oi_1 _18125_ (.Y(_11293_),
    .B1(_11292_),
    .B2(_11107_),
    .A2(_11291_),
    .A1(\cpu.ex.r_mult[20] ));
 sg13g2_nand3_1 _18126_ (.B(_11290_),
    .C(_11293_),
    .A(_10956_),
    .Y(_11294_));
 sg13g2_nand2_1 _18127_ (.Y(_11295_),
    .A(_09404_),
    .B(_10892_));
 sg13g2_o21ai_1 _18128_ (.B1(_11295_),
    .Y(_11296_),
    .A1(_11287_),
    .A2(_11294_));
 sg13g2_buf_1 _18129_ (.A(_11296_),
    .X(_11297_));
 sg13g2_or3_1 _18130_ (.A(\cpu.ex.c_mult_off[1] ),
    .B(_11249_),
    .C(_11297_),
    .X(_11298_));
 sg13g2_inv_1 _18131_ (.Y(_11299_),
    .A(\cpu.addr[8] ));
 sg13g2_buf_1 _18132_ (.A(_11299_),
    .X(_11300_));
 sg13g2_nand3_1 _18133_ (.B(net768),
    .C(net762),
    .A(\cpu.ex.r_9[8] ),
    .Y(_11301_));
 sg13g2_nand3_1 _18134_ (.B(net676),
    .C(_10945_),
    .A(\cpu.ex.r_stmp[8] ),
    .Y(_11302_));
 sg13g2_mux2_1 _18135_ (.A0(_10505_),
    .A1(\cpu.ex.r_epc[8] ),
    .S(_10901_),
    .X(_11303_));
 sg13g2_nand3_1 _18136_ (.B(_11103_),
    .C(_11303_),
    .A(_10924_),
    .Y(_11304_));
 sg13g2_nand3_1 _18137_ (.B(_11302_),
    .C(_11304_),
    .A(_11301_),
    .Y(_11305_));
 sg13g2_nand3_1 _18138_ (.B(\cpu.ex.r_10[8] ),
    .C(net676),
    .A(_10933_),
    .Y(_11306_));
 sg13g2_nand3_1 _18139_ (.B(\cpu.ex.r_lr[8] ),
    .C(net768),
    .A(_10924_),
    .Y(_11307_));
 sg13g2_a21oi_1 _18140_ (.A1(_11306_),
    .A2(_11307_),
    .Y(_11308_),
    .B1(net767));
 sg13g2_inv_1 _18141_ (.Y(_11309_),
    .A(_00250_));
 sg13g2_a22oi_1 _18142_ (.Y(_11310_),
    .B1(net761),
    .B2(\cpu.ex.r_12[8] ),
    .A2(_10928_),
    .A1(_11309_));
 sg13g2_nor2b_1 _18143_ (.A(_11310_),
    .B_N(_10980_),
    .Y(_11311_));
 sg13g2_a22oi_1 _18144_ (.Y(_11312_),
    .B1(_11024_),
    .B2(\cpu.ex.r_14[8] ),
    .A2(_11113_),
    .A1(\cpu.ex.r_8[8] ));
 sg13g2_nor2b_1 _18145_ (.A(_11312_),
    .B_N(_11150_),
    .Y(_11313_));
 sg13g2_nor4_1 _18146_ (.A(_11305_),
    .B(_11308_),
    .C(_11311_),
    .D(_11313_),
    .Y(_11314_));
 sg13g2_a22oi_1 _18147_ (.Y(_11315_),
    .B1(net762),
    .B2(\cpu.ex.r_11[8] ),
    .A2(net765),
    .A1(\cpu.ex.r_mult[24] ));
 sg13g2_nand3_1 _18148_ (.B(\cpu.ex.r_13[8] ),
    .C(_10976_),
    .A(net760),
    .Y(_11316_));
 sg13g2_o21ai_1 _18149_ (.B1(_11316_),
    .Y(_11317_),
    .A1(net895),
    .A2(_11315_));
 sg13g2_a21oi_1 _18150_ (.A1(_10903_),
    .A2(_11317_),
    .Y(_11318_),
    .B1(net568));
 sg13g2_a22oi_1 _18151_ (.Y(_11319_),
    .B1(_11314_),
    .B2(_11318_),
    .A2(net568),
    .A1(_11300_));
 sg13g2_buf_1 _18152_ (.A(_11319_),
    .X(_11320_));
 sg13g2_nor4_1 _18153_ (.A(net1068),
    .B(_09348_),
    .C(_11246_),
    .D(\cpu.ex.c_mult_off[0] ),
    .Y(_11321_));
 sg13g2_a22oi_1 _18154_ (.Y(_11322_),
    .B1(_11007_),
    .B2(_10708_),
    .A2(_11000_),
    .A1(\cpu.ex.r_stmp[7] ));
 sg13g2_nor2_1 _18155_ (.A(net896),
    .B(_11322_),
    .Y(_11323_));
 sg13g2_nor2b_1 _18156_ (.A(_10903_),
    .B_N(_10916_),
    .Y(_11324_));
 sg13g2_a22oi_1 _18157_ (.Y(_11325_),
    .B1(_11324_),
    .B2(\cpu.ex.r_14[7] ),
    .A2(_11268_),
    .A1(\cpu.ex.r_11[7] ));
 sg13g2_nor2_1 _18158_ (.A(net759),
    .B(_11325_),
    .Y(_11326_));
 sg13g2_o21ai_1 _18159_ (.B1(net763),
    .Y(_11327_),
    .A1(_11323_),
    .A2(_11326_));
 sg13g2_a22oi_1 _18160_ (.Y(_11328_),
    .B1(_11066_),
    .B2(\cpu.ex.r_13[7] ),
    .A2(_11019_),
    .A1(\cpu.ex.r_8[7] ));
 sg13g2_a22oi_1 _18161_ (.Y(_11329_),
    .B1(_11324_),
    .B2(\cpu.ex.r_12[7] ),
    .A2(_11268_),
    .A1(\cpu.ex.r_9[7] ));
 sg13g2_a21oi_1 _18162_ (.A1(_11328_),
    .A2(_11329_),
    .Y(_11330_),
    .B1(_10993_));
 sg13g2_nand2_1 _18163_ (.Y(_11331_),
    .A(_10940_),
    .B(_11330_));
 sg13g2_nand3_1 _18164_ (.B(\cpu.ex.r_mult[23] ),
    .C(net765),
    .A(net677),
    .Y(_11332_));
 sg13g2_nand3_1 _18165_ (.B(\cpu.ex.r_10[7] ),
    .C(_11150_),
    .A(_10920_),
    .Y(_11333_));
 sg13g2_nand2_1 _18166_ (.Y(_11334_),
    .A(_11332_),
    .B(_11333_));
 sg13g2_nand3_1 _18167_ (.B(_10723_),
    .C(net761),
    .A(net767),
    .Y(_11335_));
 sg13g2_nand3_1 _18168_ (.B(\cpu.ex.r_epc[7] ),
    .C(_10928_),
    .A(_10920_),
    .Y(_11336_));
 sg13g2_nand2_1 _18169_ (.Y(_11337_),
    .A(_11335_),
    .B(_11336_));
 sg13g2_a22oi_1 _18170_ (.Y(_11338_),
    .B1(_10911_),
    .B2(\cpu.ex.r_lr[7] ),
    .A2(net676),
    .A1(_10722_));
 sg13g2_nor2b_1 _18171_ (.A(_11338_),
    .B_N(_10930_),
    .Y(_11339_));
 sg13g2_a221oi_1 _18172_ (.B2(net759),
    .C1(_11339_),
    .B1(_11337_),
    .A1(net763),
    .Y(_11340_),
    .A2(_11334_));
 sg13g2_nand4_1 _18173_ (.B(_11327_),
    .C(_11331_),
    .A(net567),
    .Y(_11341_),
    .D(_11340_));
 sg13g2_a21oi_1 _18174_ (.A1(_09223_),
    .A2(_10893_),
    .Y(_11342_),
    .B1(_11252_));
 sg13g2_a22oi_1 _18175_ (.Y(_11343_),
    .B1(_11341_),
    .B2(_11342_),
    .A2(_11321_),
    .A1(_11320_));
 sg13g2_nand2_1 _18176_ (.Y(_11344_),
    .A(_10744_),
    .B(net568));
 sg13g2_nand2_1 _18177_ (.Y(_11345_),
    .A(\cpu.ex.r_stmp[5] ),
    .B(_11120_));
 sg13g2_nand3_1 _18178_ (.B(\cpu.ex.r_10[5] ),
    .C(net676),
    .A(net675),
    .Y(_11346_));
 sg13g2_nand3_1 _18179_ (.B(\cpu.ex.r_lr[5] ),
    .C(_10911_),
    .A(net759),
    .Y(_11347_));
 sg13g2_a21o_1 _18180_ (.A2(_11347_),
    .A1(_11346_),
    .B1(_10917_),
    .X(_11348_));
 sg13g2_a22oi_1 _18181_ (.Y(_11349_),
    .B1(_11174_),
    .B2(\cpu.ex.r_13[5] ),
    .A2(_10932_),
    .A1(\cpu.ex.r_epc[5] ));
 sg13g2_nand3_1 _18182_ (.B(_10930_),
    .C(net676),
    .A(_10753_),
    .Y(_11350_));
 sg13g2_and3_1 _18183_ (.X(_11351_),
    .A(_11348_),
    .B(_11349_),
    .C(_11350_));
 sg13g2_mux2_1 _18184_ (.A0(\cpu.ex.r_12[5] ),
    .A1(\cpu.ex.r_14[5] ),
    .S(_10961_),
    .X(_11352_));
 sg13g2_nand3_1 _18185_ (.B(_11150_),
    .C(_11352_),
    .A(_10917_),
    .Y(_11353_));
 sg13g2_nand3_1 _18186_ (.B(net768),
    .C(net762),
    .A(\cpu.ex.r_9[5] ),
    .Y(_11354_));
 sg13g2_nand3_1 _18187_ (.B(net762),
    .C(net761),
    .A(\cpu.ex.r_8[5] ),
    .Y(_11355_));
 sg13g2_nand3_1 _18188_ (.B(_11354_),
    .C(_11355_),
    .A(_11353_),
    .Y(_11356_));
 sg13g2_nor2b_1 _18189_ (.A(_00247_),
    .B_N(_10916_),
    .Y(_11357_));
 sg13g2_nor2b_1 _18190_ (.A(net897),
    .B_N(\cpu.ex.r_11[5] ),
    .Y(_11358_));
 sg13g2_o21ai_1 _18191_ (.B1(_11098_),
    .Y(_11359_),
    .A1(_11357_),
    .A2(_11358_));
 sg13g2_nand2_1 _18192_ (.Y(_11360_),
    .A(\cpu.ex.r_mult[21] ),
    .B(net765));
 sg13g2_a21oi_1 _18193_ (.A1(_11359_),
    .A2(_11360_),
    .Y(_11361_),
    .B1(_10981_));
 sg13g2_nor2_1 _18194_ (.A(_11356_),
    .B(_11361_),
    .Y(_11362_));
 sg13g2_nand4_1 _18195_ (.B(_11345_),
    .C(_11351_),
    .A(net567),
    .Y(_11363_),
    .D(_11362_));
 sg13g2_nand3_1 _18196_ (.B(_11344_),
    .C(_11363_),
    .A(_11257_),
    .Y(_11364_));
 sg13g2_and4_1 _18197_ (.A(_11278_),
    .B(_11298_),
    .C(_11343_),
    .D(_11364_),
    .X(_11365_));
 sg13g2_nand2_1 _18198_ (.Y(_11366_),
    .A(net241),
    .B(_11365_));
 sg13g2_a22oi_1 _18199_ (.Y(_11367_),
    .B1(_11259_),
    .B2(_11366_),
    .A2(_11245_),
    .A1(_11223_));
 sg13g2_nand4_1 _18200_ (.B(_11188_),
    .C(_11221_),
    .A(_11086_),
    .Y(_11368_),
    .D(_11367_));
 sg13g2_buf_1 _18201_ (.A(_11368_),
    .X(_11369_));
 sg13g2_and2_1 _18202_ (.A(_10846_),
    .B(_10867_),
    .X(_11370_));
 sg13g2_a21o_1 _18203_ (.A2(_10732_),
    .A1(_10731_),
    .B1(_10736_),
    .X(_11371_));
 sg13g2_buf_1 _18204_ (.A(_11371_),
    .X(_11372_));
 sg13g2_nor2_1 _18205_ (.A(net1120),
    .B(_11372_),
    .Y(_11373_));
 sg13g2_nor2_1 _18206_ (.A(_10707_),
    .B(_11373_),
    .Y(_11374_));
 sg13g2_nor2_1 _18207_ (.A(net1042),
    .B(_11373_),
    .Y(_11375_));
 sg13g2_inv_1 _18208_ (.Y(_11376_),
    .A(_10823_));
 sg13g2_a21oi_1 _18209_ (.A1(_11376_),
    .A2(_10842_),
    .Y(_11377_),
    .B1(_10839_));
 sg13g2_nand3_1 _18210_ (.B(_10839_),
    .C(_10842_),
    .A(_11376_),
    .Y(_11378_));
 sg13g2_o21ai_1 _18211_ (.B1(_11378_),
    .Y(_11379_),
    .A1(_10830_),
    .A2(_11377_));
 sg13g2_o21ai_1 _18212_ (.B1(_11379_),
    .Y(_11380_),
    .A1(_11374_),
    .A2(_11375_));
 sg13g2_nor3_1 _18213_ (.A(net1042),
    .B(_10707_),
    .C(_11373_),
    .Y(_11381_));
 sg13g2_a21oi_1 _18214_ (.A1(net1120),
    .A2(_11372_),
    .Y(_11382_),
    .B1(_11381_));
 sg13g2_a21oi_1 _18215_ (.A1(_11380_),
    .A2(_11382_),
    .Y(_11383_),
    .B1(net799));
 sg13g2_a221oi_1 _18216_ (.B2(_11370_),
    .C1(_11383_),
    .B1(_11369_),
    .A1(_10846_),
    .Y(_11384_),
    .A2(_10874_));
 sg13g2_buf_1 _18217_ (.A(_11384_),
    .X(_11385_));
 sg13g2_o21ai_1 _18218_ (.B1(net242),
    .Y(_11386_),
    .A1(_10522_),
    .A2(_11385_));
 sg13g2_o21ai_1 _18219_ (.B1(_10808_),
    .Y(_11387_),
    .A1(_09351_),
    .A2(net220));
 sg13g2_buf_1 _18220_ (.A(_00287_),
    .X(_11388_));
 sg13g2_a21oi_1 _18221_ (.A1(net169),
    .A2(_11385_),
    .Y(_11389_),
    .B1(_11388_));
 sg13g2_nor3_1 _18222_ (.A(_10522_),
    .B(_11385_),
    .C(net242),
    .Y(_11390_));
 sg13g2_a221oi_1 _18223_ (.B2(_11389_),
    .C1(_11390_),
    .B1(_11387_),
    .A1(_10809_),
    .Y(_11391_),
    .A2(_11386_));
 sg13g2_buf_1 _18224_ (.A(_11391_),
    .X(_11392_));
 sg13g2_buf_1 _18225_ (.A(_00285_),
    .X(_11393_));
 sg13g2_o21ai_1 _18226_ (.B1(_11393_),
    .Y(_11394_),
    .A1(net200),
    .A2(_11392_));
 sg13g2_buf_1 _18227_ (.A(_11394_),
    .X(_11395_));
 sg13g2_nand2_1 _18228_ (.Y(_11396_),
    .A(_10410_),
    .B(_10836_));
 sg13g2_buf_2 _18229_ (.A(_11396_),
    .X(_11397_));
 sg13g2_buf_1 _18230_ (.A(_10388_),
    .X(_11398_));
 sg13g2_nor2_1 _18231_ (.A(net909),
    .B(_00275_),
    .Y(_11399_));
 sg13g2_nor3_2 _18232_ (.A(net901),
    .B(_10391_),
    .C(_10419_),
    .Y(_11400_));
 sg13g2_nor2_2 _18233_ (.A(_11399_),
    .B(_11400_),
    .Y(_11401_));
 sg13g2_buf_1 _18234_ (.A(_10836_),
    .X(_11402_));
 sg13g2_a21oi_1 _18235_ (.A1(_11401_),
    .A2(_11390_),
    .Y(_11403_),
    .B1(net566));
 sg13g2_a221oi_1 _18236_ (.B2(net199),
    .C1(_11403_),
    .B1(_11397_),
    .A1(net200),
    .Y(_11404_),
    .A2(_11392_));
 sg13g2_buf_1 _18237_ (.A(_11404_),
    .X(_11405_));
 sg13g2_buf_1 _18238_ (.A(net799),
    .X(_11406_));
 sg13g2_or2_1 _18239_ (.X(_11407_),
    .B(net674),
    .A(_00283_));
 sg13g2_buf_1 _18240_ (.A(_11407_),
    .X(_11408_));
 sg13g2_inv_1 _18241_ (.Y(_11409_),
    .A(_10263_));
 sg13g2_buf_2 _18242_ (.A(_00284_),
    .X(_11410_));
 sg13g2_inv_1 _18243_ (.Y(_11411_),
    .A(_11410_));
 sg13g2_o21ai_1 _18244_ (.B1(net222),
    .Y(_11412_),
    .A1(_11410_),
    .A2(_10348_));
 sg13g2_a22oi_1 _18245_ (.Y(_11413_),
    .B1(_11412_),
    .B2(_10322_),
    .A2(_10349_),
    .A1(_11411_));
 sg13g2_a21oi_1 _18246_ (.A1(_11409_),
    .A2(_11413_),
    .Y(_11414_),
    .B1(net674));
 sg13g2_a21oi_1 _18247_ (.A1(net770),
    .A2(_10483_),
    .Y(_11415_),
    .B1(_10484_));
 sg13g2_buf_2 _18248_ (.A(_11415_),
    .X(_11416_));
 sg13g2_buf_1 _18249_ (.A(_11416_),
    .X(_11417_));
 sg13g2_nor3_1 _18250_ (.A(_11409_),
    .B(net674),
    .C(_11413_),
    .Y(_11418_));
 sg13g2_a21oi_2 _18251_ (.B1(_11418_),
    .Y(_11419_),
    .A2(net168),
    .A1(_11414_));
 sg13g2_or2_1 _18252_ (.X(_11420_),
    .B(_11397_),
    .A(net199));
 sg13g2_nand3_1 _18253_ (.B(_11419_),
    .C(_11420_),
    .A(_11408_),
    .Y(_11421_));
 sg13g2_buf_1 _18254_ (.A(_10455_),
    .X(_11422_));
 sg13g2_nand3_1 _18255_ (.B(_11419_),
    .C(_11420_),
    .A(net167),
    .Y(_11423_));
 sg13g2_a22oi_1 _18256_ (.Y(_11424_),
    .B1(_11421_),
    .B2(_11423_),
    .A2(_11405_),
    .A1(_11395_));
 sg13g2_buf_1 _18257_ (.A(_11424_),
    .X(_11425_));
 sg13g2_nand2_1 _18258_ (.Y(_11426_),
    .A(_11408_),
    .B(net167));
 sg13g2_a21oi_1 _18259_ (.A1(net770),
    .A2(_10292_),
    .Y(_11427_),
    .B1(_10293_));
 sg13g2_buf_1 _18260_ (.A(_11427_),
    .X(_11428_));
 sg13g2_and2_1 _18261_ (.A(_10300_),
    .B(_10346_),
    .X(_11429_));
 sg13g2_buf_2 _18262_ (.A(_11429_),
    .X(_11430_));
 sg13g2_nor3_1 _18263_ (.A(_10322_),
    .B(_11410_),
    .C(_11430_),
    .Y(_11431_));
 sg13g2_xnor2_1 _18264_ (.Y(_11432_),
    .A(_11410_),
    .B(_11430_));
 sg13g2_nor2_1 _18265_ (.A(_10323_),
    .B(net219),
    .Y(_11433_));
 sg13g2_a22oi_1 _18266_ (.Y(_11434_),
    .B1(_11432_),
    .B2(_11433_),
    .A2(_11431_),
    .A1(net219));
 sg13g2_o21ai_1 _18267_ (.B1(_10836_),
    .Y(_11435_),
    .A1(_10322_),
    .A2(_11411_));
 sg13g2_nand2_1 _18268_ (.Y(_11436_),
    .A(_10349_),
    .B(_11435_));
 sg13g2_o21ai_1 _18269_ (.B1(_11436_),
    .Y(_11437_),
    .A1(net674),
    .A2(_11434_));
 sg13g2_nand2_1 _18270_ (.Y(_11438_),
    .A(_10263_),
    .B(net566));
 sg13g2_xnor2_1 _18271_ (.Y(_11439_),
    .A(_11438_),
    .B(_11416_));
 sg13g2_nand2_1 _18272_ (.Y(_11440_),
    .A(_11437_),
    .B(_11439_));
 sg13g2_nand3_1 _18273_ (.B(_11419_),
    .C(_11440_),
    .A(_11408_),
    .Y(_11441_));
 sg13g2_nand3_1 _18274_ (.B(_11419_),
    .C(_11440_),
    .A(net167),
    .Y(_11442_));
 sg13g2_nand3_1 _18275_ (.B(_11441_),
    .C(_11442_),
    .A(_11426_),
    .Y(_11443_));
 sg13g2_buf_1 _18276_ (.A(_11443_),
    .X(_11444_));
 sg13g2_nor2_1 _18277_ (.A(_11425_),
    .B(_11444_),
    .Y(_11445_));
 sg13g2_buf_2 _18278_ (.A(_11445_),
    .X(_11446_));
 sg13g2_buf_1 _18279_ (.A(_10674_),
    .X(_11447_));
 sg13g2_buf_1 _18280_ (.A(net240),
    .X(_11448_));
 sg13g2_buf_1 _18281_ (.A(net218),
    .X(_11449_));
 sg13g2_and4_1 _18282_ (.A(_11086_),
    .B(_11188_),
    .C(_11221_),
    .D(_11367_),
    .X(_11450_));
 sg13g2_buf_2 _18283_ (.A(_11450_),
    .X(_11451_));
 sg13g2_buf_1 _18284_ (.A(_11451_),
    .X(_11452_));
 sg13g2_buf_1 _18285_ (.A(net124),
    .X(_11453_));
 sg13g2_nor3_1 _18286_ (.A(_10802_),
    .B(net198),
    .C(net109),
    .Y(_11454_));
 sg13g2_a21oi_1 _18287_ (.A1(net87),
    .A2(_11446_),
    .Y(_11455_),
    .B1(_11454_));
 sg13g2_buf_1 _18288_ (.A(\cpu.ex.r_mult[0] ),
    .X(_11456_));
 sg13g2_nor2_1 _18289_ (.A(_09345_),
    .B(net1133),
    .Y(_11457_));
 sg13g2_and2_1 _18290_ (.A(_09342_),
    .B(_11457_),
    .X(_11458_));
 sg13g2_buf_1 _18291_ (.A(_11458_),
    .X(_11459_));
 sg13g2_and2_1 _18292_ (.A(_10199_),
    .B(_10201_),
    .X(_11460_));
 sg13g2_buf_1 _18293_ (.A(_11460_),
    .X(_11461_));
 sg13g2_nand2b_1 _18294_ (.Y(_11462_),
    .B(_11461_),
    .A_N(_11459_));
 sg13g2_buf_2 _18295_ (.A(_11462_),
    .X(_11463_));
 sg13g2_nand2_1 _18296_ (.Y(_11464_),
    .A(_11456_),
    .B(_11463_));
 sg13g2_o21ai_1 _18297_ (.B1(_11464_),
    .Y(\cpu.ex.c_mult[0] ),
    .A1(_10203_),
    .A2(_11455_));
 sg13g2_buf_1 _18298_ (.A(\cpu.dec.load ),
    .X(_11465_));
 sg13g2_nand2_1 _18299_ (.Y(_11466_),
    .A(_08345_),
    .B(net371));
 sg13g2_nand2b_1 _18300_ (.Y(_11467_),
    .B(_09155_),
    .A_N(_09350_));
 sg13g2_nand2b_1 _18301_ (.Y(_11468_),
    .B(_11467_),
    .A_N(_11457_));
 sg13g2_buf_1 _18302_ (.A(_11468_),
    .X(_11469_));
 sg13g2_nor2_1 _18303_ (.A(\cpu.ex.c_div_running ),
    .B(\cpu.ex.c_mult_running ),
    .Y(_11470_));
 sg13g2_nand2_1 _18304_ (.Y(_11471_),
    .A(_10657_),
    .B(\cpu.dec.r_swapsp ));
 sg13g2_nand2_1 _18305_ (.Y(_11472_),
    .A(\cpu.dec.iready ),
    .B(_00189_));
 sg13g2_nor2_1 _18306_ (.A(\cpu.ex.r_branch_stall ),
    .B(_11472_),
    .Y(_11473_));
 sg13g2_buf_2 _18307_ (.A(_11473_),
    .X(_11474_));
 sg13g2_nand2_2 _18308_ (.Y(_11475_),
    .A(_09155_),
    .B(_11474_));
 sg13g2_nor2_1 _18309_ (.A(net1074),
    .B(_11475_),
    .Y(_11476_));
 sg13g2_buf_1 _18310_ (.A(net1117),
    .X(_11477_));
 sg13g2_nand2_1 _18311_ (.Y(_11478_),
    .A(net1036),
    .B(\cpu.cond[2] ));
 sg13g2_nand2_1 _18312_ (.Y(_11479_),
    .A(_00242_),
    .B(_11478_));
 sg13g2_nand2_1 _18313_ (.Y(_11480_),
    .A(net1144),
    .B(_11479_));
 sg13g2_buf_1 _18314_ (.A(_11480_),
    .X(_11481_));
 sg13g2_o21ai_1 _18315_ (.B1(_11481_),
    .Y(_11482_),
    .A1(net1036),
    .A2(\cpu.dec.jmp ));
 sg13g2_nand4_1 _18316_ (.B(_11471_),
    .C(_11476_),
    .A(_11470_),
    .Y(_11483_),
    .D(_11482_));
 sg13g2_nand3_1 _18317_ (.B(net239),
    .C(_11483_),
    .A(_11466_),
    .Y(_11484_));
 sg13g2_buf_1 _18318_ (.A(_11484_),
    .X(_11485_));
 sg13g2_and2_1 _18319_ (.A(net928),
    .B(_11485_),
    .X(_11486_));
 sg13g2_buf_1 _18320_ (.A(_11486_),
    .X(_11487_));
 sg13g2_nand2_1 _18321_ (.Y(_11488_),
    .A(_00294_),
    .B(_11487_));
 sg13g2_inv_1 _18322_ (.Y(_11489_),
    .A(_09817_));
 sg13g2_o21ai_1 _18323_ (.B1(_09821_),
    .Y(_11490_),
    .A1(_09814_),
    .A2(_11489_));
 sg13g2_nor2b_2 _18324_ (.A(_09219_),
    .B_N(_11490_),
    .Y(_11491_));
 sg13g2_inv_1 _18325_ (.Y(_11492_),
    .A(_11491_));
 sg13g2_o21ai_1 _18326_ (.B1(_11488_),
    .Y(_11493_),
    .A1(_11487_),
    .A2(_11492_));
 sg13g2_nand2_1 _18327_ (.Y(_11494_),
    .A(_09214_),
    .B(_11493_));
 sg13g2_o21ai_1 _18328_ (.B1(_11494_),
    .Y(_00054_),
    .A1(_11465_),
    .A2(_11488_));
 sg13g2_buf_1 _18329_ (.A(\cpu.ex.r_mult[1] ),
    .X(_11495_));
 sg13g2_buf_1 _18330_ (.A(_11463_),
    .X(_11496_));
 sg13g2_buf_1 _18331_ (.A(_11461_),
    .X(_11497_));
 sg13g2_inv_1 _18332_ (.Y(_11498_),
    .A(net1133));
 sg13g2_buf_1 _18333_ (.A(_10953_),
    .X(_11499_));
 sg13g2_buf_1 _18334_ (.A(_11499_),
    .X(_11500_));
 sg13g2_buf_1 _18335_ (.A(_11500_),
    .X(_11501_));
 sg13g2_buf_1 _18336_ (.A(_11501_),
    .X(_11502_));
 sg13g2_nand2_1 _18337_ (.Y(_11503_),
    .A(_11456_),
    .B(net460));
 sg13g2_buf_1 _18338_ (.A(net284),
    .X(_11504_));
 sg13g2_nor2_1 _18339_ (.A(_11504_),
    .B(_11451_),
    .Y(_11505_));
 sg13g2_mux2_1 _18340_ (.A0(_11503_),
    .A1(_11456_),
    .S(_11505_),
    .X(_11506_));
 sg13g2_buf_1 _18341_ (.A(net616),
    .X(_11507_));
 sg13g2_a22oi_1 _18342_ (.Y(_11508_),
    .B1(_11505_),
    .B2(net564),
    .A2(net99),
    .A1(_11456_));
 sg13g2_o21ai_1 _18343_ (.B1(_11508_),
    .Y(_11509_),
    .A1(net1035),
    .A2(_11506_));
 sg13g2_and2_1 _18344_ (.A(_11497_),
    .B(_11509_),
    .X(_11510_));
 sg13g2_a21oi_1 _18345_ (.A1(_11495_),
    .A2(net359),
    .Y(_11511_),
    .B1(_11510_));
 sg13g2_inv_1 _18346_ (.Y(\cpu.ex.c_mult[1] ),
    .A(_11511_));
 sg13g2_buf_2 _18347_ (.A(\cpu.ex.r_mult[2] ),
    .X(_11512_));
 sg13g2_and3_1 _18348_ (.X(_11513_),
    .A(_11456_),
    .B(_10339_),
    .C(_10622_));
 sg13g2_a21o_1 _18349_ (.A2(_10640_),
    .A1(_10622_),
    .B1(_10648_),
    .X(_11514_));
 sg13g2_a22oi_1 _18350_ (.Y(_11515_),
    .B1(_11514_),
    .B2(_11456_),
    .A2(_11513_),
    .A1(_10639_));
 sg13g2_buf_1 _18351_ (.A(_11369_),
    .X(_11516_));
 sg13g2_buf_1 _18352_ (.A(net123),
    .X(_11517_));
 sg13g2_buf_1 _18353_ (.A(net360),
    .X(_11518_));
 sg13g2_nor2_1 _18354_ (.A(_11495_),
    .B(net278),
    .Y(_11519_));
 sg13g2_inv_1 _18355_ (.Y(_11520_),
    .A(_11495_));
 sg13g2_nor2_1 _18356_ (.A(_11520_),
    .B(net286),
    .Y(_11521_));
 sg13g2_a21oi_1 _18357_ (.A1(net108),
    .A2(_11519_),
    .Y(_11522_),
    .B1(_11521_));
 sg13g2_and2_1 _18358_ (.A(net286),
    .B(_11515_),
    .X(_11523_));
 sg13g2_o21ai_1 _18359_ (.B1(_11495_),
    .Y(_11524_),
    .A1(net124),
    .A2(_11523_));
 sg13g2_o21ai_1 _18360_ (.B1(_11524_),
    .Y(_11525_),
    .A1(_11515_),
    .A2(_11522_));
 sg13g2_buf_1 _18361_ (.A(net108),
    .X(_11526_));
 sg13g2_a221oi_1 _18362_ (.B2(_11456_),
    .C1(_11495_),
    .B1(_11514_),
    .A1(_10639_),
    .Y(_11527_),
    .A2(_11513_));
 sg13g2_and3_1 _18363_ (.X(_11528_),
    .A(net278),
    .B(net98),
    .C(_11527_));
 sg13g2_a21oi_1 _18364_ (.A1(net460),
    .A2(_11525_),
    .Y(_11529_),
    .B1(_11528_));
 sg13g2_nor2_2 _18365_ (.A(net460),
    .B(_11452_),
    .Y(_11530_));
 sg13g2_a22oi_1 _18366_ (.Y(_11531_),
    .B1(_11530_),
    .B2(net278),
    .A2(net99),
    .A1(_11495_));
 sg13g2_o21ai_1 _18367_ (.B1(_11531_),
    .Y(_11532_),
    .A1(net1035),
    .A2(_11529_));
 sg13g2_a22oi_1 _18368_ (.Y(_11533_),
    .B1(_11532_),
    .B2(net461),
    .A2(_11463_),
    .A1(_11512_));
 sg13g2_inv_1 _18369_ (.Y(\cpu.ex.c_mult[2] ),
    .A(_11533_));
 sg13g2_buf_2 _18370_ (.A(\cpu.ex.r_mult[3] ),
    .X(_11534_));
 sg13g2_or3_1 _18371_ (.A(_10581_),
    .B(_10586_),
    .C(_11527_),
    .X(_11535_));
 sg13g2_or2_1 _18372_ (.X(_11536_),
    .B(_11515_),
    .A(_11520_));
 sg13g2_nand2_1 _18373_ (.Y(_11537_),
    .A(_11535_),
    .B(_11536_));
 sg13g2_inv_1 _18374_ (.Y(_11538_),
    .A(_11537_));
 sg13g2_buf_1 _18375_ (.A(_10864_),
    .X(_11539_));
 sg13g2_buf_1 _18376_ (.A(net237),
    .X(_11540_));
 sg13g2_nor2_1 _18377_ (.A(_11512_),
    .B(net217),
    .Y(_11541_));
 sg13g2_and2_1 _18378_ (.A(_11512_),
    .B(net237),
    .X(_11542_));
 sg13g2_a21oi_1 _18379_ (.A1(net108),
    .A2(_11541_),
    .Y(_11543_),
    .B1(_11542_));
 sg13g2_nor2_1 _18380_ (.A(_11540_),
    .B(_11537_),
    .Y(_11544_));
 sg13g2_o21ai_1 _18381_ (.B1(_11512_),
    .Y(_11545_),
    .A1(_11452_),
    .A2(_11544_));
 sg13g2_o21ai_1 _18382_ (.B1(_11545_),
    .Y(_11546_),
    .A1(_11538_),
    .A2(_11543_));
 sg13g2_buf_1 _18383_ (.A(net285),
    .X(_11547_));
 sg13g2_nor4_1 _18384_ (.A(_11512_),
    .B(net236),
    .C(net109),
    .D(_11537_),
    .Y(_11548_));
 sg13g2_a21oi_1 _18385_ (.A1(net460),
    .A2(_11546_),
    .Y(_11549_),
    .B1(_11548_));
 sg13g2_a22oi_1 _18386_ (.Y(_11550_),
    .B1(_11530_),
    .B2(_11540_),
    .A2(net99),
    .A1(_11512_));
 sg13g2_o21ai_1 _18387_ (.B1(_11550_),
    .Y(_11551_),
    .A1(_11498_),
    .A2(_11549_));
 sg13g2_a22oi_1 _18388_ (.Y(_11552_),
    .B1(_11551_),
    .B2(net461),
    .A2(net359),
    .A1(_11534_));
 sg13g2_inv_1 _18389_ (.Y(\cpu.ex.c_mult[3] ),
    .A(_11552_));
 sg13g2_buf_1 _18390_ (.A(\cpu.ex.r_mult[4] ),
    .X(_11553_));
 sg13g2_buf_1 _18391_ (.A(_10842_),
    .X(_11554_));
 sg13g2_nor2_1 _18392_ (.A(_11534_),
    .B(net277),
    .Y(_11555_));
 sg13g2_nand2b_1 _18393_ (.Y(_11556_),
    .B(net285),
    .A_N(_11512_));
 sg13g2_nand3_1 _18394_ (.B(_10611_),
    .C(_10616_),
    .A(_11512_),
    .Y(_11557_));
 sg13g2_nand3_1 _18395_ (.B(_11536_),
    .C(_11557_),
    .A(_11535_),
    .Y(_11558_));
 sg13g2_nand2_1 _18396_ (.Y(_11559_),
    .A(_11556_),
    .B(_11558_));
 sg13g2_buf_1 _18397_ (.A(_11559_),
    .X(_11560_));
 sg13g2_inv_1 _18398_ (.Y(_11561_),
    .A(_11560_));
 sg13g2_inv_1 _18399_ (.Y(_11562_),
    .A(_11534_));
 sg13g2_nand2_1 _18400_ (.Y(_11563_),
    .A(_11562_),
    .B(net277));
 sg13g2_o21ai_1 _18401_ (.B1(_11534_),
    .Y(_11564_),
    .A1(_10825_),
    .A2(_10827_));
 sg13g2_o21ai_1 _18402_ (.B1(_11564_),
    .Y(_11565_),
    .A1(net124),
    .A2(_11563_));
 sg13g2_nor2_1 _18403_ (.A(_11562_),
    .B(net108),
    .Y(_11566_));
 sg13g2_a21o_1 _18404_ (.A2(_11565_),
    .A1(_11561_),
    .B1(_11566_),
    .X(_11567_));
 sg13g2_nand3_1 _18405_ (.B(net460),
    .C(net277),
    .A(_11534_),
    .Y(_11568_));
 sg13g2_nand2_1 _18406_ (.Y(_11569_),
    .A(net108),
    .B(_11555_));
 sg13g2_a21oi_1 _18407_ (.A1(_11568_),
    .A2(_11569_),
    .Y(_11570_),
    .B1(_11561_));
 sg13g2_a221oi_1 _18408_ (.B2(net460),
    .C1(_11570_),
    .B1(_11567_),
    .A1(_11530_),
    .Y(_11571_),
    .A2(_11555_));
 sg13g2_a22oi_1 _18409_ (.Y(_11572_),
    .B1(_11530_),
    .B2(_10798_),
    .A2(net99),
    .A1(_11534_));
 sg13g2_o21ai_1 _18410_ (.B1(_11572_),
    .Y(_11573_),
    .A1(net1035),
    .A2(_11571_));
 sg13g2_a22oi_1 _18411_ (.Y(_11574_),
    .B1(_11573_),
    .B2(net461),
    .A2(net359),
    .A1(_11553_));
 sg13g2_inv_1 _18412_ (.Y(\cpu.ex.c_mult[4] ),
    .A(_11574_));
 sg13g2_buf_2 _18413_ (.A(\cpu.ex.r_mult[5] ),
    .X(_11575_));
 sg13g2_nand2_1 _18414_ (.Y(_11576_),
    .A(_11553_),
    .B(_11502_));
 sg13g2_buf_8 _18415_ (.A(_10839_),
    .X(_11577_));
 sg13g2_a21oi_1 _18416_ (.A1(_11554_),
    .A2(_11560_),
    .Y(_11578_),
    .B1(_11562_));
 sg13g2_nor2_1 _18417_ (.A(_11554_),
    .B(_11560_),
    .Y(_11579_));
 sg13g2_o21ai_1 _18418_ (.B1(net510),
    .Y(_11580_),
    .A1(_11578_),
    .A2(_11579_));
 sg13g2_xnor2_1 _18419_ (.Y(_11581_),
    .A(_11577_),
    .B(_11580_));
 sg13g2_nor2_1 _18420_ (.A(net124),
    .B(_11581_),
    .Y(_11582_));
 sg13g2_mux2_1 _18421_ (.A0(_11576_),
    .A1(_11553_),
    .S(_11582_),
    .X(_11583_));
 sg13g2_a22oi_1 _18422_ (.Y(_11584_),
    .B1(_11582_),
    .B2(net564),
    .A2(net99),
    .A1(_11553_));
 sg13g2_o21ai_1 _18423_ (.B1(_11584_),
    .Y(_11585_),
    .A1(net1035),
    .A2(_11583_));
 sg13g2_a22oi_1 _18424_ (.Y(_11586_),
    .B1(_11585_),
    .B2(net461),
    .A2(_11496_),
    .A1(_11575_));
 sg13g2_inv_1 _18425_ (.Y(\cpu.ex.c_mult[5] ),
    .A(_11586_));
 sg13g2_buf_2 _18426_ (.A(\cpu.ex.r_mult[6] ),
    .X(_11587_));
 sg13g2_nand2_1 _18427_ (.Y(_11588_),
    .A(_11575_),
    .B(net615));
 sg13g2_buf_1 _18428_ (.A(net361),
    .X(_11589_));
 sg13g2_inv_1 _18429_ (.Y(_11590_),
    .A(_11553_));
 sg13g2_a22oi_1 _18430_ (.Y(_11591_),
    .B1(_10798_),
    .B2(_11534_),
    .A2(_10767_),
    .A1(_11553_));
 sg13g2_a21o_1 _18431_ (.A2(net235),
    .A1(_11590_),
    .B1(_11591_),
    .X(_11592_));
 sg13g2_a22oi_1 _18432_ (.Y(_11593_),
    .B1(_10842_),
    .B2(_11562_),
    .A2(net235),
    .A1(_11590_));
 sg13g2_nand3_1 _18433_ (.B(_11558_),
    .C(_11593_),
    .A(_11556_),
    .Y(_11594_));
 sg13g2_a21oi_1 _18434_ (.A1(_11592_),
    .A2(_11594_),
    .Y(_11595_),
    .B1(net616));
 sg13g2_xnor2_1 _18435_ (.Y(_11596_),
    .A(net276),
    .B(_11595_));
 sg13g2_nand2_1 _18436_ (.Y(_11597_),
    .A(net108),
    .B(_11596_));
 sg13g2_mux2_1 _18437_ (.A0(_11575_),
    .A1(_11588_),
    .S(_11597_),
    .X(_11598_));
 sg13g2_nor3_1 _18438_ (.A(net460),
    .B(net276),
    .C(net124),
    .Y(_11599_));
 sg13g2_a21oi_1 _18439_ (.A1(_11575_),
    .A2(net99),
    .Y(_11600_),
    .B1(_11599_));
 sg13g2_o21ai_1 _18440_ (.B1(_11600_),
    .Y(_11601_),
    .A1(net1035),
    .A2(_11598_));
 sg13g2_and2_1 _18441_ (.A(_11497_),
    .B(_11601_),
    .X(_11602_));
 sg13g2_a21oi_1 _18442_ (.A1(_11587_),
    .A2(_11463_),
    .Y(_11603_),
    .B1(_11602_));
 sg13g2_inv_1 _18443_ (.Y(\cpu.ex.c_mult[6] ),
    .A(_11603_));
 sg13g2_buf_2 _18444_ (.A(\cpu.ex.r_mult[7] ),
    .X(_11604_));
 sg13g2_inv_1 _18445_ (.Y(_11605_),
    .A(_11575_));
 sg13g2_nor2_1 _18446_ (.A(_11605_),
    .B(net361),
    .Y(_11606_));
 sg13g2_a221oi_1 _18447_ (.B2(_10765_),
    .C1(_11590_),
    .B1(_10742_),
    .A1(_11605_),
    .Y(_11607_),
    .A2(net361));
 sg13g2_or2_1 _18448_ (.X(_11608_),
    .B(_11607_),
    .A(_11606_));
 sg13g2_buf_1 _18449_ (.A(_11608_),
    .X(_11609_));
 sg13g2_a22oi_1 _18450_ (.Y(_11610_),
    .B1(net235),
    .B2(_11590_),
    .A2(net361),
    .A1(_11605_));
 sg13g2_a21o_1 _18451_ (.A2(_10765_),
    .A1(_10742_),
    .B1(_10818_),
    .X(_11611_));
 sg13g2_a21oi_1 _18452_ (.A1(_09338_),
    .A2(_11611_),
    .Y(_11612_),
    .B1(_11564_));
 sg13g2_nand2_1 _18453_ (.Y(_11613_),
    .A(_11610_),
    .B(_11612_));
 sg13g2_nor3_1 _18454_ (.A(_11534_),
    .B(_10825_),
    .C(_10827_),
    .Y(_11614_));
 sg13g2_a221oi_1 _18455_ (.B2(_11590_),
    .C1(_11614_),
    .B1(_11577_),
    .A1(_11605_),
    .Y(_11615_),
    .A2(_10818_));
 sg13g2_nand3_1 _18456_ (.B(net616),
    .C(_11611_),
    .A(_11562_),
    .Y(_11616_));
 sg13g2_nand2_1 _18457_ (.Y(_11617_),
    .A(_11615_),
    .B(_11616_));
 sg13g2_a21oi_1 _18458_ (.A1(_11560_),
    .A2(_11613_),
    .Y(_11618_),
    .B1(_11617_));
 sg13g2_buf_1 _18459_ (.A(_11372_),
    .X(_11619_));
 sg13g2_o21ai_1 _18460_ (.B1(net234),
    .Y(_11620_),
    .A1(_11609_),
    .A2(_11618_));
 sg13g2_or3_1 _18461_ (.A(net234),
    .B(_11609_),
    .C(_11618_),
    .X(_11621_));
 sg13g2_nand2_1 _18462_ (.Y(_11622_),
    .A(_11620_),
    .B(_11621_));
 sg13g2_inv_2 _18463_ (.Y(_11623_),
    .A(_11587_));
 sg13g2_a221oi_1 _18464_ (.B2(_11622_),
    .C1(_11623_),
    .B1(net98),
    .A1(_09333_),
    .Y(_11624_),
    .A2(_10834_));
 sg13g2_buf_1 _18465_ (.A(net283),
    .X(_11625_));
 sg13g2_a21oi_1 _18466_ (.A1(_11610_),
    .A2(_11612_),
    .Y(_11626_),
    .B1(_11609_));
 sg13g2_and2_1 _18467_ (.A(_11560_),
    .B(_11626_),
    .X(_11627_));
 sg13g2_o21ai_1 _18468_ (.B1(net565),
    .Y(_11628_),
    .A1(_11609_),
    .A2(_11615_));
 sg13g2_or3_1 _18469_ (.A(net233),
    .B(_11627_),
    .C(_11628_),
    .X(_11629_));
 sg13g2_nand2_1 _18470_ (.Y(_11630_),
    .A(_11623_),
    .B(net98));
 sg13g2_a21oi_1 _18471_ (.A1(_11621_),
    .A2(_11629_),
    .Y(_11631_),
    .B1(_11630_));
 sg13g2_o21ai_1 _18472_ (.B1(net1133),
    .Y(_11632_),
    .A1(_11624_),
    .A2(_11631_));
 sg13g2_a22oi_1 _18473_ (.Y(_11633_),
    .B1(_11530_),
    .B2(net233),
    .A2(net99),
    .A1(_11587_));
 sg13g2_a21oi_1 _18474_ (.A1(_11632_),
    .A2(_11633_),
    .Y(_11634_),
    .B1(_10203_));
 sg13g2_a21oi_1 _18475_ (.A1(_11604_),
    .A2(net359),
    .Y(_11635_),
    .B1(_11634_));
 sg13g2_inv_1 _18476_ (.Y(\cpu.ex.c_mult[7] ),
    .A(_11635_));
 sg13g2_a21o_1 _18477_ (.A2(_11594_),
    .A1(_11592_),
    .B1(_09354_),
    .X(_11636_));
 sg13g2_buf_1 _18478_ (.A(_11636_),
    .X(_11637_));
 sg13g2_nand2_2 _18479_ (.Y(_11638_),
    .A(_11587_),
    .B(net283));
 sg13g2_o21ai_1 _18480_ (.B1(_11606_),
    .Y(_11639_),
    .A1(_11587_),
    .A2(net283));
 sg13g2_buf_1 _18481_ (.A(_11639_),
    .X(_11640_));
 sg13g2_nand2_1 _18482_ (.Y(_11641_),
    .A(_11638_),
    .B(_11640_));
 sg13g2_nand2_1 _18483_ (.Y(_11642_),
    .A(net565),
    .B(_11641_));
 sg13g2_buf_1 _18484_ (.A(_10707_),
    .X(_11643_));
 sg13g2_nor3_1 _18485_ (.A(_11623_),
    .B(_09338_),
    .C(net361),
    .Y(_11644_));
 sg13g2_a21oi_1 _18486_ (.A1(_11623_),
    .A2(net234),
    .Y(_11645_),
    .B1(_11588_));
 sg13g2_or2_1 _18487_ (.X(_11646_),
    .B(_11645_),
    .A(_11644_));
 sg13g2_buf_1 _18488_ (.A(_11646_),
    .X(_11647_));
 sg13g2_a221oi_1 _18489_ (.B2(net510),
    .C1(_11647_),
    .B1(_11641_),
    .A1(net232),
    .Y(_11648_),
    .A2(_11625_));
 sg13g2_a221oi_1 _18490_ (.B2(_11642_),
    .C1(_11648_),
    .B1(_11637_),
    .A1(_10489_),
    .Y(_11649_),
    .A2(_10520_));
 sg13g2_nand2_1 _18491_ (.Y(_11650_),
    .A(_11643_),
    .B(net283));
 sg13g2_nand2b_1 _18492_ (.Y(_11651_),
    .B(_11650_),
    .A_N(_11647_));
 sg13g2_a221oi_1 _18493_ (.B2(_11595_),
    .C1(_10523_),
    .B1(_11651_),
    .A1(net510),
    .Y(_11652_),
    .A2(_11641_));
 sg13g2_nor3_1 _18494_ (.A(_11451_),
    .B(_11649_),
    .C(_11652_),
    .Y(_11653_));
 sg13g2_inv_1 _18495_ (.Y(_11654_),
    .A(_11604_));
 sg13g2_nand2_1 _18496_ (.Y(_11655_),
    .A(_11604_),
    .B(net615));
 sg13g2_buf_1 _18497_ (.A(_11655_),
    .X(_11656_));
 sg13g2_nor2_1 _18498_ (.A(_11653_),
    .B(_11656_),
    .Y(_11657_));
 sg13g2_a21oi_1 _18499_ (.A1(_11654_),
    .A2(_11653_),
    .Y(_11658_),
    .B1(_11657_));
 sg13g2_nor2_1 _18500_ (.A(net1035),
    .B(_11658_),
    .Y(_11659_));
 sg13g2_a221oi_1 _18501_ (.B2(net564),
    .C1(_11659_),
    .B1(_11653_),
    .A1(_11604_),
    .Y(_11660_),
    .A2(_10806_));
 sg13g2_buf_1 _18502_ (.A(\cpu.ex.r_mult[8] ),
    .X(_11661_));
 sg13g2_buf_1 _18503_ (.A(_11661_),
    .X(_11662_));
 sg13g2_nand2_1 _18504_ (.Y(_11663_),
    .A(net1034),
    .B(_11463_));
 sg13g2_o21ai_1 _18505_ (.B1(_11663_),
    .Y(\cpu.ex.c_mult[8] ),
    .A1(_10203_),
    .A2(_11660_));
 sg13g2_buf_2 _18506_ (.A(\cpu.ex.r_mult[9] ),
    .X(_11664_));
 sg13g2_and2_1 _18507_ (.A(_11664_),
    .B(net359),
    .X(_11665_));
 sg13g2_nand2_1 _18508_ (.Y(_11666_),
    .A(_11661_),
    .B(net615));
 sg13g2_nor2_1 _18509_ (.A(_10545_),
    .B(_10546_),
    .Y(_11667_));
 sg13g2_a21oi_1 _18510_ (.A1(net901),
    .A2(_10548_),
    .Y(_11668_),
    .B1(_11667_));
 sg13g2_buf_2 _18511_ (.A(_11668_),
    .X(_11669_));
 sg13g2_nand3_1 _18512_ (.B(_11642_),
    .C(_11656_),
    .A(_11637_),
    .Y(_11670_));
 sg13g2_nor2_1 _18513_ (.A(_10206_),
    .B(_10487_),
    .Y(_11671_));
 sg13g2_a21oi_2 _18514_ (.B1(_10518_),
    .Y(_11672_),
    .A2(_10517_),
    .A1(_10516_));
 sg13g2_nor2_1 _18515_ (.A(_11671_),
    .B(_11672_),
    .Y(_11673_));
 sg13g2_buf_1 _18516_ (.A(_11673_),
    .X(_11674_));
 sg13g2_nand3_1 _18517_ (.B(_11637_),
    .C(_11642_),
    .A(net216),
    .Y(_11675_));
 sg13g2_nand2_1 _18518_ (.Y(_11676_),
    .A(_11650_),
    .B(_11656_));
 sg13g2_nand2_1 _18519_ (.Y(_11677_),
    .A(net216),
    .B(_11650_));
 sg13g2_a221oi_1 _18520_ (.B2(_11677_),
    .C1(_11647_),
    .B1(_11676_),
    .A1(net565),
    .Y(_11678_),
    .A2(_11641_));
 sg13g2_a21oi_1 _18521_ (.A1(net216),
    .A2(_11656_),
    .Y(_11679_),
    .B1(_11678_));
 sg13g2_and3_1 _18522_ (.X(_11680_),
    .A(_11670_),
    .B(_11675_),
    .C(_11679_));
 sg13g2_xnor2_1 _18523_ (.Y(_11681_),
    .A(_11669_),
    .B(_11680_));
 sg13g2_nand2_1 _18524_ (.Y(_11682_),
    .A(_11526_),
    .B(_11681_));
 sg13g2_mux2_1 _18525_ (.A0(_11662_),
    .A1(_11666_),
    .S(_11682_),
    .X(_11683_));
 sg13g2_nor3_1 _18526_ (.A(net1035),
    .B(_10203_),
    .C(_11683_),
    .Y(_11684_));
 sg13g2_nand3_1 _18527_ (.B(_11526_),
    .C(_11681_),
    .A(net564),
    .Y(_11685_));
 sg13g2_nand2_1 _18528_ (.Y(_11686_),
    .A(_11662_),
    .B(net87));
 sg13g2_a21oi_1 _18529_ (.A1(_11685_),
    .A2(_11686_),
    .Y(_11687_),
    .B1(_10203_));
 sg13g2_or3_1 _18530_ (.A(_11665_),
    .B(_11684_),
    .C(_11687_),
    .X(\cpu.ex.c_mult[9] ));
 sg13g2_inv_1 _18531_ (.Y(_11688_),
    .A(_11664_));
 sg13g2_nor2_1 _18532_ (.A(_11688_),
    .B(net703),
    .Y(_11689_));
 sg13g2_nor2_1 _18533_ (.A(net1034),
    .B(net242),
    .Y(_11690_));
 sg13g2_nand3_1 _18534_ (.B(_11638_),
    .C(_11640_),
    .A(_11674_),
    .Y(_11691_));
 sg13g2_a21oi_1 _18535_ (.A1(_11638_),
    .A2(_11640_),
    .Y(_11692_),
    .B1(_11674_));
 sg13g2_a21oi_1 _18536_ (.A1(_11604_),
    .A2(_11691_),
    .Y(_11693_),
    .B1(_11692_));
 sg13g2_nand2_1 _18537_ (.Y(_11694_),
    .A(net1034),
    .B(net220));
 sg13g2_o21ai_1 _18538_ (.B1(_11694_),
    .Y(_11695_),
    .A1(_11690_),
    .A2(_11693_));
 sg13g2_nand2_1 _18539_ (.Y(_11696_),
    .A(_11623_),
    .B(net234));
 sg13g2_nand4_1 _18540_ (.B(_11589_),
    .C(_11638_),
    .A(_11575_),
    .Y(_11697_),
    .D(_11696_));
 sg13g2_nand4_1 _18541_ (.B(_11587_),
    .C(_10707_),
    .A(_11605_),
    .Y(_11698_),
    .D(net234));
 sg13g2_a21o_1 _18542_ (.A2(_11698_),
    .A1(_11697_),
    .B1(net616),
    .X(_11699_));
 sg13g2_o21ai_1 _18543_ (.B1(_11500_),
    .Y(_11700_),
    .A1(_11575_),
    .A2(_11587_));
 sg13g2_nand3_1 _18544_ (.B(_11625_),
    .C(_11700_),
    .A(_11643_),
    .Y(_11701_));
 sg13g2_mux2_1 _18545_ (.A0(_11666_),
    .A1(_11661_),
    .S(net242),
    .X(_11702_));
 sg13g2_nand2_1 _18546_ (.Y(_11703_),
    .A(net703),
    .B(_10551_));
 sg13g2_o21ai_1 _18547_ (.B1(_11703_),
    .Y(_11704_),
    .A1(_11604_),
    .A2(_11702_));
 sg13g2_nor4_1 _18548_ (.A(_11661_),
    .B(_10522_),
    .C(_11669_),
    .D(_11656_),
    .Y(_11705_));
 sg13g2_a21oi_1 _18549_ (.A1(_10522_),
    .A2(_11704_),
    .Y(_11706_),
    .B1(_11705_));
 sg13g2_nor2_1 _18550_ (.A(_10522_),
    .B(net242),
    .Y(_11707_));
 sg13g2_inv_1 _18551_ (.Y(_11708_),
    .A(_11661_));
 sg13g2_nor2_1 _18552_ (.A(_11708_),
    .B(_11656_),
    .Y(_11709_));
 sg13g2_nand2_1 _18553_ (.Y(_11710_),
    .A(_11707_),
    .B(_11709_));
 sg13g2_a221oi_1 _18554_ (.B2(_11710_),
    .C1(_11637_),
    .B1(_11706_),
    .A1(_11699_),
    .Y(_11711_),
    .A2(_11701_));
 sg13g2_a21o_1 _18555_ (.A2(_11695_),
    .A1(net510),
    .B1(_11711_),
    .X(_11712_));
 sg13g2_buf_1 _18556_ (.A(_11712_),
    .X(_11713_));
 sg13g2_xnor2_1 _18557_ (.Y(_11714_),
    .A(net200),
    .B(_11713_));
 sg13g2_nor2_1 _18558_ (.A(net124),
    .B(_11714_),
    .Y(_11715_));
 sg13g2_mux2_1 _18559_ (.A0(_11689_),
    .A1(_11688_),
    .S(_11715_),
    .X(_11716_));
 sg13g2_nor3_1 _18560_ (.A(_11502_),
    .B(_11453_),
    .C(_11714_),
    .Y(_11717_));
 sg13g2_a221oi_1 _18561_ (.B2(net1133),
    .C1(_11717_),
    .B1(_11716_),
    .A1(_11664_),
    .Y(_11718_),
    .A2(_10806_));
 sg13g2_buf_1 _18562_ (.A(\cpu.ex.r_mult[10] ),
    .X(_11719_));
 sg13g2_nand2_1 _18563_ (.Y(_11720_),
    .A(_11719_),
    .B(net359));
 sg13g2_o21ai_1 _18564_ (.B1(_11720_),
    .Y(\cpu.ex.c_mult[10] ),
    .A1(_10203_),
    .A2(_11718_));
 sg13g2_buf_2 _18565_ (.A(\cpu.ex.r_mult[11] ),
    .X(_11721_));
 sg13g2_nor2_2 _18566_ (.A(_10802_),
    .B(_10203_),
    .Y(_11722_));
 sg13g2_nand2_1 _18567_ (.Y(_11723_),
    .A(net1116),
    .B(net615));
 sg13g2_nor4_1 _18568_ (.A(_11587_),
    .B(_11654_),
    .C(_11671_),
    .D(_11672_),
    .Y(_11724_));
 sg13g2_nor2_1 _18569_ (.A(_09338_),
    .B(_11619_),
    .Y(_11725_));
 sg13g2_nand2_1 _18570_ (.Y(_11726_),
    .A(_11623_),
    .B(_11654_));
 sg13g2_a221oi_1 _18571_ (.B2(_11499_),
    .C1(_11619_),
    .B1(_11726_),
    .A1(_10489_),
    .Y(_11727_),
    .A2(_10520_));
 sg13g2_a21oi_1 _18572_ (.A1(_11724_),
    .A2(_11725_),
    .Y(_11728_),
    .B1(_11727_));
 sg13g2_nor3_1 _18573_ (.A(_11604_),
    .B(_11671_),
    .C(_11672_),
    .Y(_11729_));
 sg13g2_o21ai_1 _18574_ (.B1(_11604_),
    .Y(_11730_),
    .A1(_11671_),
    .A2(_11672_));
 sg13g2_nor3_1 _18575_ (.A(_11623_),
    .B(_09338_),
    .C(_10738_),
    .Y(_11731_));
 sg13g2_nand3b_1 _18576_ (.B(_11730_),
    .C(_11731_),
    .Y(_11732_),
    .A_N(_11729_));
 sg13g2_a221oi_1 _18577_ (.B2(_11732_),
    .C1(_11628_),
    .B1(_11728_),
    .A1(_11560_),
    .Y(_11733_),
    .A2(_11626_));
 sg13g2_nand2_1 _18578_ (.Y(_11734_),
    .A(_11664_),
    .B(net615));
 sg13g2_nor3_1 _18579_ (.A(_11399_),
    .B(_11400_),
    .C(_11734_),
    .Y(_11735_));
 sg13g2_a21oi_1 _18580_ (.A1(_10390_),
    .A2(_10420_),
    .Y(_11736_),
    .B1(_11664_));
 sg13g2_o21ai_1 _18581_ (.B1(_11708_),
    .Y(_11737_),
    .A1(_11735_),
    .A2(_11736_));
 sg13g2_nand2_1 _18582_ (.Y(_11738_),
    .A(net703),
    .B(net221));
 sg13g2_nand3_1 _18583_ (.B(_11737_),
    .C(_11738_),
    .A(_10551_),
    .Y(_11739_));
 sg13g2_nand4_1 _18584_ (.B(_11688_),
    .C(net565),
    .A(net1034),
    .Y(_11740_),
    .D(net221));
 sg13g2_nand2_1 _18585_ (.Y(_11741_),
    .A(_11669_),
    .B(_11740_));
 sg13g2_and3_1 _18586_ (.X(_11742_),
    .A(_11733_),
    .B(_11739_),
    .C(_11741_));
 sg13g2_nand2_1 _18587_ (.Y(_11743_),
    .A(_11688_),
    .B(_11401_));
 sg13g2_o21ai_1 _18588_ (.B1(_11730_),
    .Y(_11744_),
    .A1(_11638_),
    .A2(_11729_));
 sg13g2_nand4_1 _18589_ (.B(net565),
    .C(_11743_),
    .A(net1034),
    .Y(_11745_),
    .D(_11744_));
 sg13g2_nand4_1 _18590_ (.B(net565),
    .C(_10552_),
    .A(net1034),
    .Y(_11746_),
    .D(_11743_));
 sg13g2_nand4_1 _18591_ (.B(net221),
    .C(_10552_),
    .A(net565),
    .Y(_11747_),
    .D(_11744_));
 sg13g2_nor2_1 _18592_ (.A(_11669_),
    .B(_11734_),
    .Y(_11748_));
 sg13g2_a22oi_1 _18593_ (.Y(_11749_),
    .B1(_11744_),
    .B2(_11748_),
    .A2(_11689_),
    .A1(net221));
 sg13g2_nand4_1 _18594_ (.B(_11746_),
    .C(_11747_),
    .A(_11745_),
    .Y(_11750_),
    .D(_11749_));
 sg13g2_a21oi_1 _18595_ (.A1(net123),
    .A2(_11742_),
    .Y(_11751_),
    .B1(_11750_));
 sg13g2_nand2_1 _18596_ (.Y(_11752_),
    .A(_11401_),
    .B(_11669_));
 sg13g2_nand3_1 _18597_ (.B(_11689_),
    .C(_11733_),
    .A(net1034),
    .Y(_11753_));
 sg13g2_a21o_1 _18598_ (.A2(_11752_),
    .A1(net123),
    .B1(_11753_),
    .X(_11754_));
 sg13g2_buf_1 _18599_ (.A(_11754_),
    .X(_11755_));
 sg13g2_a21o_1 _18600_ (.A2(_11755_),
    .A1(_11751_),
    .B1(net199),
    .X(_11756_));
 sg13g2_nand3_1 _18601_ (.B(_11751_),
    .C(_11755_),
    .A(net199),
    .Y(_11757_));
 sg13g2_a21oi_1 _18602_ (.A1(_11756_),
    .A2(_11757_),
    .Y(_11758_),
    .B1(_11453_));
 sg13g2_xnor2_1 _18603_ (.Y(_11759_),
    .A(_11723_),
    .B(_11758_));
 sg13g2_inv_1 _18604_ (.Y(_11760_),
    .A(net1116));
 sg13g2_nand2_1 _18605_ (.Y(_11761_),
    .A(_11461_),
    .B(net99));
 sg13g2_nor2_1 _18606_ (.A(_11760_),
    .B(_11761_),
    .Y(_11762_));
 sg13g2_a221oi_1 _18607_ (.B2(_11759_),
    .C1(_11762_),
    .B1(_11722_),
    .A1(_11721_),
    .Y(_11763_),
    .A2(_11463_));
 sg13g2_inv_1 _18608_ (.Y(\cpu.ex.c_mult[11] ),
    .A(_11763_));
 sg13g2_nor2_1 _18609_ (.A(_11760_),
    .B(_11734_),
    .Y(_11764_));
 sg13g2_o21ai_1 _18610_ (.B1(_11764_),
    .Y(_11765_),
    .A1(_11451_),
    .A2(_10423_));
 sg13g2_mux2_1 _18611_ (.A0(_00274_),
    .A1(_10384_),
    .S(net909),
    .X(_11766_));
 sg13g2_buf_8 _18612_ (.A(_11766_),
    .X(_11767_));
 sg13g2_mux2_1 _18613_ (.A0(net1116),
    .A1(_11723_),
    .S(net215),
    .X(_11768_));
 sg13g2_nand2_1 _18614_ (.Y(_11769_),
    .A(_09338_),
    .B(_10388_));
 sg13g2_o21ai_1 _18615_ (.B1(_11769_),
    .Y(_11770_),
    .A1(_11664_),
    .A2(_11768_));
 sg13g2_nor3_1 _18616_ (.A(net1116),
    .B(net221),
    .C(_11734_),
    .Y(_11771_));
 sg13g2_a22oi_1 _18617_ (.Y(_11772_),
    .B1(_11771_),
    .B2(_10388_),
    .A2(_11770_),
    .A1(net221));
 sg13g2_nand2b_1 _18618_ (.Y(_11773_),
    .B(_11369_),
    .A_N(_11772_));
 sg13g2_nand2_1 _18619_ (.Y(_11774_),
    .A(_11765_),
    .B(_11773_));
 sg13g2_o21ai_1 _18620_ (.B1(_11694_),
    .Y(_11775_),
    .A1(_11690_),
    .A2(_11730_));
 sg13g2_o21ai_1 _18621_ (.B1(_11664_),
    .Y(_11776_),
    .A1(_11399_),
    .A2(_11400_));
 sg13g2_a21oi_2 _18622_ (.B1(_11776_),
    .Y(_11777_),
    .A2(_11767_),
    .A1(_11760_));
 sg13g2_a221oi_1 _18623_ (.B2(_11775_),
    .C1(_11777_),
    .B1(_11774_),
    .A1(net1116),
    .Y(_11778_),
    .A2(net199));
 sg13g2_a21oi_1 _18624_ (.A1(_11637_),
    .A2(_11642_),
    .Y(_11779_),
    .B1(_11648_));
 sg13g2_o21ai_1 _18625_ (.B1(_11709_),
    .Y(_11780_),
    .A1(_11451_),
    .A2(_11707_));
 sg13g2_nand2_1 _18626_ (.Y(_11781_),
    .A(_11706_),
    .B(_11780_));
 sg13g2_nand3_1 _18627_ (.B(_11774_),
    .C(_11781_),
    .A(_11779_),
    .Y(_11782_));
 sg13g2_o21ai_1 _18628_ (.B1(_11782_),
    .Y(_11783_),
    .A1(_11507_),
    .A2(_11778_));
 sg13g2_xnor2_1 _18629_ (.Y(_11784_),
    .A(_11430_),
    .B(_11783_));
 sg13g2_nand2b_1 _18630_ (.Y(_11785_),
    .B(_11461_),
    .A_N(_10802_));
 sg13g2_buf_1 _18631_ (.A(_11785_),
    .X(_11786_));
 sg13g2_nand2_2 _18632_ (.Y(_11787_),
    .A(_11721_),
    .B(net565));
 sg13g2_or2_1 _18633_ (.X(_11788_),
    .B(_11787_),
    .A(_11786_));
 sg13g2_a21oi_1 _18634_ (.A1(net98),
    .A2(_11784_),
    .Y(_11789_),
    .B1(_11788_));
 sg13g2_nand4_1 _18635_ (.B(_11722_),
    .C(_11784_),
    .A(net98),
    .Y(_11790_),
    .D(_11787_));
 sg13g2_buf_1 _18636_ (.A(\cpu.ex.r_mult[12] ),
    .X(_11791_));
 sg13g2_and2_1 _18637_ (.A(_11461_),
    .B(net87),
    .X(_11792_));
 sg13g2_buf_1 _18638_ (.A(_11792_),
    .X(_11793_));
 sg13g2_a22oi_1 _18639_ (.Y(_11794_),
    .B1(_11793_),
    .B2(_11721_),
    .A2(net359),
    .A1(_11791_));
 sg13g2_nand3b_1 _18640_ (.B(_11790_),
    .C(_11794_),
    .Y(\cpu.ex.c_mult[12] ),
    .A_N(_11789_));
 sg13g2_buf_1 _18641_ (.A(net222),
    .X(_11795_));
 sg13g2_and3_1 _18642_ (.X(_11796_),
    .A(_10424_),
    .B(_10303_),
    .C(_10344_));
 sg13g2_inv_1 _18643_ (.Y(_11797_),
    .A(_11721_));
 sg13g2_nand2_1 _18644_ (.Y(_11798_),
    .A(_11797_),
    .B(_10300_));
 sg13g2_nand2_1 _18645_ (.Y(_11799_),
    .A(net909),
    .B(net1116));
 sg13g2_nand3_1 _18646_ (.B(_10385_),
    .C(net1116),
    .A(_10298_),
    .Y(_11800_));
 sg13g2_o21ai_1 _18647_ (.B1(_11800_),
    .Y(_11801_),
    .A1(_10384_),
    .A2(_11799_));
 sg13g2_buf_1 _18648_ (.A(_11801_),
    .X(_11802_));
 sg13g2_o21ai_1 _18649_ (.B1(_11802_),
    .Y(_11803_),
    .A1(_11796_),
    .A2(_11798_));
 sg13g2_a21o_1 _18650_ (.A2(_10346_),
    .A1(_10300_),
    .B1(_11797_),
    .X(_11804_));
 sg13g2_a21oi_1 _18651_ (.A1(_11803_),
    .A2(_11804_),
    .Y(_11805_),
    .B1(_10801_));
 sg13g2_nand2_1 _18652_ (.Y(_11806_),
    .A(_11760_),
    .B(net199));
 sg13g2_mux2_1 _18653_ (.A0(_11721_),
    .A1(_11787_),
    .S(_11430_),
    .X(_11807_));
 sg13g2_buf_1 _18654_ (.A(_10348_),
    .X(_11808_));
 sg13g2_nor3_1 _18655_ (.A(_11721_),
    .B(_10388_),
    .C(_11723_),
    .Y(_11809_));
 sg13g2_a21oi_1 _18656_ (.A1(_10300_),
    .A2(_10346_),
    .Y(_11810_),
    .B1(net215));
 sg13g2_a22oi_1 _18657_ (.Y(_11811_),
    .B1(_11810_),
    .B2(_10801_),
    .A2(_11809_),
    .A1(net144));
 sg13g2_o21ai_1 _18658_ (.B1(_11811_),
    .Y(_11812_),
    .A1(_11806_),
    .A2(_11807_));
 sg13g2_nand2_1 _18659_ (.Y(_11813_),
    .A(net108),
    .B(_11812_));
 sg13g2_nand2_1 _18660_ (.Y(_11814_),
    .A(_11430_),
    .B(net215));
 sg13g2_nand3_1 _18661_ (.B(_11721_),
    .C(_11501_),
    .A(net1116),
    .Y(_11815_));
 sg13g2_a21o_1 _18662_ (.A2(_11814_),
    .A1(net123),
    .B1(_11815_),
    .X(_11816_));
 sg13g2_nand2_1 _18663_ (.Y(_11817_),
    .A(net1034),
    .B(_11689_));
 sg13g2_a21oi_1 _18664_ (.A1(net108),
    .A2(_11752_),
    .Y(_11818_),
    .B1(_11817_));
 sg13g2_and3_1 _18665_ (.X(_11819_),
    .A(net123),
    .B(_11739_),
    .C(_11741_));
 sg13g2_o21ai_1 _18666_ (.B1(_11680_),
    .Y(_11820_),
    .A1(_11818_),
    .A2(_11819_));
 sg13g2_nor2_1 _18667_ (.A(_11664_),
    .B(_10807_),
    .Y(_11821_));
 sg13g2_o21ai_1 _18668_ (.B1(_11776_),
    .Y(_11822_),
    .A1(_11694_),
    .A2(_11821_));
 sg13g2_nand2_1 _18669_ (.Y(_11823_),
    .A(net510),
    .B(_11822_));
 sg13g2_a22oi_1 _18670_ (.Y(_11824_),
    .B1(_11820_),
    .B2(_11823_),
    .A2(_11816_),
    .A1(_11813_));
 sg13g2_nor2_1 _18671_ (.A(_11805_),
    .B(_11824_),
    .Y(_11825_));
 sg13g2_xnor2_1 _18672_ (.Y(_11826_),
    .A(net197),
    .B(_11825_));
 sg13g2_inv_1 _18673_ (.Y(_11827_),
    .A(_11791_));
 sg13g2_nor2_2 _18674_ (.A(_11827_),
    .B(_09338_),
    .Y(_11828_));
 sg13g2_nor3_1 _18675_ (.A(net109),
    .B(_11786_),
    .C(_11828_),
    .Y(_11829_));
 sg13g2_nor3_1 _18676_ (.A(net219),
    .B(net124),
    .C(_11805_),
    .Y(_11830_));
 sg13g2_nor2_1 _18677_ (.A(net197),
    .B(net109),
    .Y(_11831_));
 sg13g2_mux2_1 _18678_ (.A0(_11830_),
    .A1(_11831_),
    .S(_11824_),
    .X(_11832_));
 sg13g2_nand2_1 _18679_ (.Y(_11833_),
    .A(net219),
    .B(_11805_));
 sg13g2_nor2_1 _18680_ (.A(net616),
    .B(_11786_),
    .Y(_11834_));
 sg13g2_buf_1 _18681_ (.A(_11834_),
    .X(_11835_));
 sg13g2_o21ai_1 _18682_ (.B1(_11835_),
    .Y(_11836_),
    .A1(net109),
    .A2(_11833_));
 sg13g2_o21ai_1 _18683_ (.B1(_11761_),
    .Y(_11837_),
    .A1(_11832_),
    .A2(_11836_));
 sg13g2_buf_1 _18684_ (.A(\cpu.ex.r_mult[13] ),
    .X(_11838_));
 sg13g2_and2_1 _18685_ (.A(_11838_),
    .B(_11463_),
    .X(_11839_));
 sg13g2_a221oi_1 _18686_ (.B2(_11791_),
    .C1(_11839_),
    .B1(_11837_),
    .A1(_11826_),
    .Y(_11840_),
    .A2(_11829_));
 sg13g2_buf_1 _18687_ (.A(_11840_),
    .X(_11841_));
 sg13g2_inv_1 _18688_ (.Y(\cpu.ex.c_mult[13] ),
    .A(_11841_));
 sg13g2_nand2_1 _18689_ (.Y(_11842_),
    .A(_11838_),
    .B(net615));
 sg13g2_buf_2 _18690_ (.A(_11842_),
    .X(_11843_));
 sg13g2_nor2_1 _18691_ (.A(_11827_),
    .B(_11787_),
    .Y(_11844_));
 sg13g2_o21ai_1 _18692_ (.B1(_11844_),
    .Y(_11845_),
    .A1(_10349_),
    .A2(_11451_));
 sg13g2_nand2_1 _18693_ (.Y(_11846_),
    .A(_11791_),
    .B(net615));
 sg13g2_nor2_1 _18694_ (.A(net222),
    .B(_11846_),
    .Y(_11847_));
 sg13g2_a21oi_1 _18695_ (.A1(_11827_),
    .A2(net222),
    .Y(_11848_),
    .B1(_11847_));
 sg13g2_nand2_1 _18696_ (.Y(_11849_),
    .A(_09354_),
    .B(net222));
 sg13g2_o21ai_1 _18697_ (.B1(_11849_),
    .Y(_11850_),
    .A1(_11721_),
    .A2(_11848_));
 sg13g2_nor3_1 _18698_ (.A(_11791_),
    .B(_10348_),
    .C(_11787_),
    .Y(_11851_));
 sg13g2_a22oi_1 _18699_ (.Y(_11852_),
    .B1(_11851_),
    .B2(net222),
    .A2(_11850_),
    .A1(net144));
 sg13g2_a221oi_1 _18700_ (.B2(_11852_),
    .C1(_11451_),
    .B1(_11845_),
    .A1(_11765_),
    .Y(_11853_),
    .A2(_11773_));
 sg13g2_buf_1 _18701_ (.A(_11853_),
    .X(_11854_));
 sg13g2_and2_1 _18702_ (.A(_11713_),
    .B(_11854_),
    .X(_11855_));
 sg13g2_a221oi_1 _18703_ (.B2(_11827_),
    .C1(_11797_),
    .B1(_11427_),
    .A1(_09333_),
    .Y(_11856_),
    .A2(_10834_));
 sg13g2_o21ai_1 _18704_ (.B1(_11856_),
    .Y(_11857_),
    .A1(_11777_),
    .A2(_11802_));
 sg13g2_a221oi_1 _18705_ (.B2(_10346_),
    .C1(_11427_),
    .B1(_10300_),
    .A1(_09333_),
    .Y(_11858_),
    .A2(_10834_));
 sg13g2_o21ai_1 _18706_ (.B1(_11858_),
    .Y(_11859_),
    .A1(_11777_),
    .A2(_11802_));
 sg13g2_a21oi_1 _18707_ (.A1(_10300_),
    .A2(_10346_),
    .Y(_11860_),
    .B1(_11846_));
 sg13g2_o21ai_1 _18708_ (.B1(_11860_),
    .Y(_11861_),
    .A1(_11777_),
    .A2(_11802_));
 sg13g2_a21oi_1 _18709_ (.A1(_11827_),
    .A2(_11427_),
    .Y(_11862_),
    .B1(_11797_));
 sg13g2_a21oi_1 _18710_ (.A1(_10300_),
    .A2(_10346_),
    .Y(_11863_),
    .B1(net703));
 sg13g2_a22oi_1 _18711_ (.Y(_11864_),
    .B1(_11862_),
    .B2(_11863_),
    .A2(_11828_),
    .A1(net222));
 sg13g2_nand4_1 _18712_ (.B(_11859_),
    .C(_11861_),
    .A(_11857_),
    .Y(_11865_),
    .D(_11864_));
 sg13g2_buf_1 _18713_ (.A(_11865_),
    .X(_11866_));
 sg13g2_a21oi_1 _18714_ (.A1(_11713_),
    .A2(_11854_),
    .Y(_11867_),
    .B1(_11866_));
 sg13g2_nor2_1 _18715_ (.A(net168),
    .B(net109),
    .Y(_11868_));
 sg13g2_and3_1 _18716_ (.X(_11869_),
    .A(net168),
    .B(net98),
    .C(_11866_));
 sg13g2_a221oi_1 _18717_ (.B2(_11868_),
    .C1(_11869_),
    .B1(_11867_),
    .A1(net168),
    .Y(_11870_),
    .A2(_11855_));
 sg13g2_xnor2_1 _18718_ (.Y(_11871_),
    .A(_11843_),
    .B(_11870_));
 sg13g2_nor2_1 _18719_ (.A(_11786_),
    .B(_11871_),
    .Y(_11872_));
 sg13g2_a221oi_1 _18720_ (.B2(_11838_),
    .C1(_11872_),
    .B1(_11793_),
    .A1(\cpu.ex.r_mult[14] ),
    .Y(_11873_),
    .A2(net359));
 sg13g2_buf_1 _18721_ (.A(_11873_),
    .X(_11874_));
 sg13g2_inv_1 _18722_ (.Y(\cpu.ex.c_mult[14] ),
    .A(_11874_));
 sg13g2_a21oi_2 _18723_ (.B1(_10453_),
    .Y(_11875_),
    .A2(_10452_),
    .A1(net770));
 sg13g2_nor2_1 _18724_ (.A(net197),
    .B(net201),
    .Y(_11876_));
 sg13g2_and2_1 _18725_ (.A(_11838_),
    .B(_11828_),
    .X(_11877_));
 sg13g2_o21ai_1 _18726_ (.B1(_11877_),
    .Y(_11878_),
    .A1(_11451_),
    .A2(_11876_));
 sg13g2_mux2_1 _18727_ (.A0(_11838_),
    .A1(_11843_),
    .S(_11416_),
    .X(_11879_));
 sg13g2_nand2_1 _18728_ (.Y(_11880_),
    .A(net703),
    .B(net201));
 sg13g2_o21ai_1 _18729_ (.B1(_11880_),
    .Y(_11881_),
    .A1(_11791_),
    .A2(_11879_));
 sg13g2_nor4_1 _18730_ (.A(_11838_),
    .B(_10295_),
    .C(_11416_),
    .D(_11846_),
    .Y(_11882_));
 sg13g2_a21o_1 _18731_ (.A2(_11881_),
    .A1(net197),
    .B1(_11882_),
    .X(_11883_));
 sg13g2_a221oi_1 _18732_ (.B2(_10424_),
    .C1(_10484_),
    .B1(_10483_),
    .A1(_11838_),
    .Y(_11884_),
    .A2(net615));
 sg13g2_buf_1 _18733_ (.A(_11884_),
    .X(_11885_));
 sg13g2_nand2b_1 _18734_ (.Y(_11886_),
    .B(_11828_),
    .A_N(_11885_));
 sg13g2_or3_1 _18735_ (.A(net703),
    .B(net219),
    .C(_11885_),
    .X(_11887_));
 sg13g2_a22oi_1 _18736_ (.Y(_11888_),
    .B1(_11886_),
    .B2(_11887_),
    .A2(_11804_),
    .A1(_11803_));
 sg13g2_nor2_1 _18737_ (.A(net219),
    .B(_11885_),
    .Y(_11889_));
 sg13g2_nor2_1 _18738_ (.A(_11416_),
    .B(_11843_),
    .Y(_11890_));
 sg13g2_a21oi_1 _18739_ (.A1(_11828_),
    .A2(_11889_),
    .Y(_11891_),
    .B1(_11890_));
 sg13g2_nand2b_1 _18740_ (.Y(_11892_),
    .B(_11891_),
    .A_N(_11888_));
 sg13g2_a21oi_1 _18741_ (.A1(_11516_),
    .A2(_11883_),
    .Y(_11893_),
    .B1(_11892_));
 sg13g2_a21oi_1 _18742_ (.A1(_11516_),
    .A2(_11812_),
    .Y(_11894_),
    .B1(_11892_));
 sg13g2_a22oi_1 _18743_ (.Y(_11895_),
    .B1(_11894_),
    .B2(_11816_),
    .A2(_11893_),
    .A1(_11878_));
 sg13g2_nand3b_1 _18744_ (.B(_11751_),
    .C(_11755_),
    .Y(_11896_),
    .A_N(_11892_));
 sg13g2_nand4_1 _18745_ (.B(_11517_),
    .C(_11895_),
    .A(_11875_),
    .Y(_11897_),
    .D(_11896_));
 sg13g2_nand2_1 _18746_ (.Y(_11898_),
    .A(_10455_),
    .B(_11517_));
 sg13g2_a21o_1 _18747_ (.A2(_11896_),
    .A1(_11895_),
    .B1(_11898_),
    .X(_11899_));
 sg13g2_buf_1 _18748_ (.A(_00155_),
    .X(_11900_));
 sg13g2_nor3_1 _18749_ (.A(net1035),
    .B(_11900_),
    .C(_11507_),
    .Y(_11901_));
 sg13g2_and3_1 _18750_ (.X(_11902_),
    .A(_11897_),
    .B(_11899_),
    .C(_11901_));
 sg13g2_nand2_1 _18751_ (.Y(_11903_),
    .A(_09353_),
    .B(_11900_));
 sg13g2_a21oi_1 _18752_ (.A1(_11897_),
    .A2(_11899_),
    .Y(_11904_),
    .B1(_11903_));
 sg13g2_nand2_1 _18753_ (.Y(_11905_),
    .A(net564),
    .B(_11422_));
 sg13g2_inv_1 _18754_ (.Y(_11906_),
    .A(_11900_));
 sg13g2_nand2_1 _18755_ (.Y(_11907_),
    .A(_11906_),
    .B(_10805_));
 sg13g2_o21ai_1 _18756_ (.B1(_11907_),
    .Y(_11908_),
    .A1(net124),
    .A2(_11905_));
 sg13g2_nor3_1 _18757_ (.A(_11902_),
    .B(_11904_),
    .C(_11908_),
    .Y(_11909_));
 sg13g2_buf_1 _18758_ (.A(\cpu.ex.r_mult[15] ),
    .X(_11910_));
 sg13g2_nand2_1 _18759_ (.Y(_11911_),
    .A(_11910_),
    .B(_11496_));
 sg13g2_o21ai_1 _18760_ (.B1(_11911_),
    .Y(\cpu.ex.c_mult[15] ),
    .A1(_10203_),
    .A2(_11909_));
 sg13g2_inv_1 _18761_ (.Y(_00000_),
    .A(net2));
 sg13g2_inv_1 _18762_ (.Y(_11912_),
    .A(_09846_));
 sg13g2_nor3_1 _18763_ (.A(_11912_),
    .B(net782),
    .C(net111),
    .Y(_00008_));
 sg13g2_buf_1 _18764_ (.A(_09158_),
    .X(_11913_));
 sg13g2_and3_1 _18765_ (.X(_00005_),
    .A(net1064),
    .B(net614),
    .C(_09837_));
 sg13g2_buf_1 _18766_ (.A(\cpu.qspi.r_state[11] ),
    .X(_11914_));
 sg13g2_inv_1 _18767_ (.Y(_11915_),
    .A(_11914_));
 sg13g2_nor2_1 _18768_ (.A(_11915_),
    .B(net705),
    .Y(_00004_));
 sg13g2_buf_2 _18769_ (.A(\cpu.qspi.r_state[10] ),
    .X(_11916_));
 sg13g2_inv_1 _18770_ (.Y(_11917_),
    .A(_11916_));
 sg13g2_nor2_1 _18771_ (.A(_11917_),
    .B(net705),
    .Y(_00003_));
 sg13g2_buf_1 _18772_ (.A(\cpu.qspi.r_state[15] ),
    .X(_11918_));
 sg13g2_and2_1 _18773_ (.A(_11918_),
    .B(net614),
    .X(_00002_));
 sg13g2_inv_1 _18774_ (.Y(_11919_),
    .A(_09841_));
 sg13g2_nor3_1 _18775_ (.A(_11919_),
    .B(net782),
    .C(_09843_),
    .Y(_00001_));
 sg13g2_and2_1 _18776_ (.A(_10950_),
    .B(_10951_),
    .X(_11920_));
 sg13g2_a21o_1 _18777_ (.A2(_10996_),
    .A1(_10957_),
    .B1(_10997_),
    .X(_11921_));
 sg13g2_buf_1 _18778_ (.A(_11921_),
    .X(_11922_));
 sg13g2_nand2_1 _18779_ (.Y(_11923_),
    .A(_11922_),
    .B(_11297_));
 sg13g2_and2_1 _18780_ (.A(_11344_),
    .B(_11363_),
    .X(_11924_));
 sg13g2_buf_1 _18781_ (.A(_11924_),
    .X(_11925_));
 sg13g2_or4_1 _18782_ (.A(_11137_),
    .B(_11184_),
    .C(_11320_),
    .D(_11925_),
    .X(_11926_));
 sg13g2_or4_1 _18783_ (.A(_11243_),
    .B(_11219_),
    .C(_11203_),
    .D(_11926_),
    .X(_11927_));
 sg13g2_nand2_1 _18784_ (.Y(_11928_),
    .A(_11071_),
    .B(_11073_));
 sg13g2_o21ai_1 _18785_ (.B1(_11341_),
    .Y(_11929_),
    .A1(net1138),
    .A2(net567));
 sg13g2_nor2b_1 _18786_ (.A(_11164_),
    .B_N(_11929_),
    .Y(_11930_));
 sg13g2_nand4_1 _18787_ (.B(_11928_),
    .C(_11277_),
    .A(_11037_),
    .Y(_11931_),
    .D(_11930_));
 sg13g2_nor4_1 _18788_ (.A(_11920_),
    .B(_11923_),
    .C(_11927_),
    .D(_11931_),
    .Y(_11932_));
 sg13g2_o21ai_1 _18789_ (.B1(_11119_),
    .Y(_11933_),
    .A1(\cpu.cond[1] ),
    .A2(_11932_));
 sg13g2_xnor2_1 _18790_ (.Y(_11934_),
    .A(_09213_),
    .B(_11933_));
 sg13g2_buf_1 _18791_ (.A(net890),
    .X(_11935_));
 sg13g2_a21o_1 _18792_ (.A2(_11934_),
    .A1(_00257_),
    .B1(_11935_),
    .X(_11936_));
 sg13g2_nor2b_1 _18793_ (.A(\cpu.dec.jmp ),
    .B_N(_11936_),
    .Y(_11937_));
 sg13g2_nor2_1 _18794_ (.A(_11475_),
    .B(_11937_),
    .Y(_00053_));
 sg13g2_buf_2 _18795_ (.A(\cpu.qspi.r_state[3] ),
    .X(_11938_));
 sg13g2_and2_1 _18796_ (.A(_11938_),
    .B(net614),
    .X(_00009_));
 sg13g2_buf_1 _18797_ (.A(\cpu.qspi.r_state[13] ),
    .X(_11939_));
 sg13g2_inv_1 _18798_ (.Y(_11940_),
    .A(_11939_));
 sg13g2_nor2_1 _18799_ (.A(_11940_),
    .B(net705),
    .Y(_00006_));
 sg13g2_nand2_1 _18800_ (.Y(_11941_),
    .A(net708),
    .B(_09870_));
 sg13g2_nor2_1 _18801_ (.A(_09869_),
    .B(_11941_),
    .Y(_00007_));
 sg13g2_buf_1 _18802_ (.A(\cpu.qspi.r_state[6] ),
    .X(_11942_));
 sg13g2_and2_1 _18803_ (.A(_11942_),
    .B(_11913_),
    .X(_00010_));
 sg13g2_buf_1 _18804_ (.A(net172),
    .X(_11943_));
 sg13g2_nor2_1 _18805_ (.A(net143),
    .B(_09323_),
    .Y(_00052_));
 sg13g2_or2_1 _18806_ (.X(_11944_),
    .B(net1134),
    .A(_09251_));
 sg13g2_buf_1 _18807_ (.A(_11944_),
    .X(_11945_));
 sg13g2_nor3_1 _18808_ (.A(net1135),
    .B(_09325_),
    .C(_11945_),
    .Y(_11946_));
 sg13g2_a21oi_1 _18809_ (.A1(_09309_),
    .A2(_11945_),
    .Y(_11947_),
    .B1(_11946_));
 sg13g2_nand2_1 _18810_ (.Y(_11948_),
    .A(_09359_),
    .B(_11947_));
 sg13g2_inv_1 _18811_ (.Y(_11949_),
    .A(_00211_));
 sg13g2_nor3_1 _18812_ (.A(_09313_),
    .B(net1135),
    .C(_11949_),
    .Y(_11950_));
 sg13g2_buf_1 _18813_ (.A(\cpu.spi.r_sel[1] ),
    .X(_11951_));
 sg13g2_buf_1 _18814_ (.A(_11951_),
    .X(_11952_));
 sg13g2_buf_1 _18815_ (.A(\cpu.spi.r_src[2] ),
    .X(_11953_));
 sg13g2_inv_1 _18816_ (.Y(_11954_),
    .A(_00266_));
 sg13g2_buf_1 _18817_ (.A(\cpu.spi.r_sel[0] ),
    .X(_11955_));
 sg13g2_buf_1 _18818_ (.A(net1115),
    .X(_11956_));
 sg13g2_mux2_1 _18819_ (.A0(_11953_),
    .A1(_11954_),
    .S(_11956_),
    .X(_11957_));
 sg13g2_nand2_1 _18820_ (.Y(_11958_),
    .A(net1115),
    .B(_00267_));
 sg13g2_o21ai_1 _18821_ (.B1(_11958_),
    .Y(_11959_),
    .A1(_11956_),
    .A2(_11954_));
 sg13g2_nor2_1 _18822_ (.A(_11951_),
    .B(_11959_),
    .Y(_11960_));
 sg13g2_a21oi_2 _18823_ (.B1(_11960_),
    .Y(_11961_),
    .A2(_11957_),
    .A1(net1033));
 sg13g2_nor2_1 _18824_ (.A(_11950_),
    .B(_11961_),
    .Y(_11962_));
 sg13g2_nor2_1 _18825_ (.A(net1071),
    .B(_09305_),
    .Y(_11963_));
 sg13g2_inv_1 _18826_ (.Y(_11964_),
    .A(_11951_));
 sg13g2_buf_1 _18827_ (.A(\cpu.spi.r_mode[0][1] ),
    .X(_11965_));
 sg13g2_buf_1 _18828_ (.A(\cpu.spi.r_mode[1][1] ),
    .X(_11966_));
 sg13g2_buf_1 _18829_ (.A(net1115),
    .X(_11967_));
 sg13g2_mux2_1 _18830_ (.A0(_11965_),
    .A1(_11966_),
    .S(net1031),
    .X(_11968_));
 sg13g2_nor2_1 _18831_ (.A(_11964_),
    .B(net1115),
    .Y(_11969_));
 sg13g2_buf_1 _18832_ (.A(\cpu.spi.r_mode[2][1] ),
    .X(_11970_));
 sg13g2_a22oi_1 _18833_ (.Y(_11971_),
    .B1(_11969_),
    .B2(_11970_),
    .A2(_11968_),
    .A1(_11964_));
 sg13g2_xnor2_1 _18834_ (.Y(_11972_),
    .A(_11963_),
    .B(_11971_));
 sg13g2_buf_1 _18835_ (.A(net1129),
    .X(_11973_));
 sg13g2_buf_1 _18836_ (.A(net1030),
    .X(_11974_));
 sg13g2_buf_1 _18837_ (.A(_09456_),
    .X(_11975_));
 sg13g2_buf_1 _18838_ (.A(_11975_),
    .X(_11976_));
 sg13g2_buf_1 _18839_ (.A(net613),
    .X(_11977_));
 sg13g2_nand2_1 _18840_ (.Y(_11978_),
    .A(net613),
    .B(_00267_));
 sg13g2_o21ai_1 _18841_ (.B1(_11978_),
    .Y(_11979_),
    .A1(net563),
    .A2(_11954_));
 sg13g2_nand3_1 _18842_ (.B(net783),
    .C(_11953_),
    .A(_11974_),
    .Y(_11980_));
 sg13g2_o21ai_1 _18843_ (.B1(_11980_),
    .Y(_11981_),
    .A1(_11974_),
    .A2(_11979_));
 sg13g2_and2_1 _18844_ (.A(_11950_),
    .B(_11981_),
    .X(_11982_));
 sg13g2_nand2b_1 _18845_ (.Y(_11983_),
    .B(net563),
    .A_N(_11965_));
 sg13g2_o21ai_1 _18846_ (.B1(_11983_),
    .Y(_11984_),
    .A1(_11977_),
    .A2(_11970_));
 sg13g2_mux2_1 _18847_ (.A0(_11965_),
    .A1(_11966_),
    .S(_11977_),
    .X(_11985_));
 sg13g2_nor2_1 _18848_ (.A(net888),
    .B(_11985_),
    .Y(_11986_));
 sg13g2_a21oi_1 _18849_ (.A1(net888),
    .A2(_11984_),
    .Y(_11987_),
    .B1(_11986_));
 sg13g2_a22oi_1 _18850_ (.Y(_11988_),
    .B1(_11982_),
    .B2(_11987_),
    .A2(_11972_),
    .A1(_11962_));
 sg13g2_nor2_1 _18851_ (.A(_11962_),
    .B(_11982_),
    .Y(_11989_));
 sg13g2_buf_1 _18852_ (.A(\cpu.gpio.genblk1[3].srcs_o[5] ),
    .X(_11990_));
 sg13g2_o21ai_1 _18853_ (.B1(net1114),
    .Y(_11991_),
    .A1(_11948_),
    .A2(_11989_));
 sg13g2_o21ai_1 _18854_ (.B1(_11991_),
    .Y(_00306_),
    .A1(_11948_),
    .A2(_11988_));
 sg13g2_nor2b_1 _18855_ (.A(_11948_),
    .B_N(_11989_),
    .Y(_11992_));
 sg13g2_or3_1 _18856_ (.A(net1134),
    .B(net1135),
    .C(_11949_),
    .X(_11993_));
 sg13g2_buf_1 _18857_ (.A(_11993_),
    .X(_11994_));
 sg13g2_and2_1 _18858_ (.A(_11950_),
    .B(_11987_),
    .X(_11995_));
 sg13g2_a21oi_1 _18859_ (.A1(net887),
    .A2(_11972_),
    .Y(_11996_),
    .B1(_11995_));
 sg13g2_buf_1 _18860_ (.A(\cpu.gpio.genblk1[3].srcs_o[4] ),
    .X(_11997_));
 sg13g2_nor2_1 _18861_ (.A(net1113),
    .B(_11992_),
    .Y(_11998_));
 sg13g2_a21oi_1 _18862_ (.A1(_11992_),
    .A2(_11996_),
    .Y(_00307_),
    .B1(_11998_));
 sg13g2_buf_1 _18863_ (.A(\cpu.gpio.genblk1[3].srcs_o[3] ),
    .X(_11999_));
 sg13g2_buf_1 _18864_ (.A(net1070),
    .X(_12000_));
 sg13g2_mux2_1 _18865_ (.A0(\cpu.spi.r_out[7] ),
    .A1(_10081_),
    .S(_12000_),
    .X(_12001_));
 sg13g2_nor2_1 _18866_ (.A(net1135),
    .B(_11945_),
    .Y(_12002_));
 sg13g2_buf_1 _18867_ (.A(\cpu.spi.r_mode[2][0] ),
    .X(_12003_));
 sg13g2_nor2b_1 _18868_ (.A(\cpu.spi.r_mode[1][0] ),
    .B_N(_11955_),
    .Y(_12004_));
 sg13g2_nor2b_1 _18869_ (.A(_11955_),
    .B_N(_00209_),
    .Y(_12005_));
 sg13g2_nor3_1 _18870_ (.A(_11951_),
    .B(_12004_),
    .C(_12005_),
    .Y(_12006_));
 sg13g2_a21oi_1 _18871_ (.A1(_12003_),
    .A2(_11969_),
    .Y(_12007_),
    .B1(_12006_));
 sg13g2_buf_1 _18872_ (.A(_12007_),
    .X(_12008_));
 sg13g2_nor2_1 _18873_ (.A(_09319_),
    .B(net672),
    .Y(_12009_));
 sg13g2_nand2_1 _18874_ (.Y(_12010_),
    .A(_09285_),
    .B(net672));
 sg13g2_a21o_1 _18875_ (.A2(_09255_),
    .A1(_00205_),
    .B1(net1134),
    .X(_12011_));
 sg13g2_o21ai_1 _18876_ (.B1(net1134),
    .Y(_12012_),
    .A1(_09307_),
    .A2(net672));
 sg13g2_nand2_1 _18877_ (.Y(_12013_),
    .A(_09304_),
    .B(_12012_));
 sg13g2_o21ai_1 _18878_ (.B1(_12013_),
    .Y(_12014_),
    .A1(_12010_),
    .A2(_12011_));
 sg13g2_nand3_1 _18879_ (.B(_09250_),
    .C(_12014_),
    .A(net928),
    .Y(_12015_));
 sg13g2_a221oi_1 _18880_ (.B2(net91),
    .C1(_12015_),
    .B1(_12009_),
    .A1(_09319_),
    .Y(_12016_),
    .A2(_12002_));
 sg13g2_nor2b_1 _18881_ (.A(_11961_),
    .B_N(_12016_),
    .Y(_12017_));
 sg13g2_mux2_1 _18882_ (.A0(net1112),
    .A1(_12001_),
    .S(_12017_),
    .X(_00308_));
 sg13g2_buf_1 _18883_ (.A(\cpu.gpio.genblk1[3].srcs_o[2] ),
    .X(_12018_));
 sg13g2_nand2_1 _18884_ (.Y(_12019_),
    .A(_11961_),
    .B(_12016_));
 sg13g2_mux2_1 _18885_ (.A0(_12001_),
    .A1(net1111),
    .S(_12019_),
    .X(_00309_));
 sg13g2_buf_1 _18886_ (.A(uio_in[0]),
    .X(_12020_));
 sg13g2_buf_1 _18887_ (.A(_12020_),
    .X(_12021_));
 sg13g2_nand2_1 _18888_ (.Y(_12022_),
    .A(net916),
    .B(net921));
 sg13g2_buf_1 _18889_ (.A(_12022_),
    .X(_12023_));
 sg13g2_buf_2 _18890_ (.A(\cpu.dcache.r_offset[1] ),
    .X(_12024_));
 sg13g2_buf_1 _18891_ (.A(_12024_),
    .X(_12025_));
 sg13g2_buf_2 _18892_ (.A(\cpu.dcache.r_offset[0] ),
    .X(_12026_));
 sg13g2_buf_1 _18893_ (.A(_12026_),
    .X(_12027_));
 sg13g2_nand2b_1 _18894_ (.Y(_12028_),
    .B(net1028),
    .A_N(net1029));
 sg13g2_buf_1 _18895_ (.A(\cpu.d_wstrobe_d ),
    .X(_12029_));
 sg13g2_buf_1 _18896_ (.A(_00260_),
    .X(_12030_));
 sg13g2_buf_1 _18897_ (.A(_12030_),
    .X(_12031_));
 sg13g2_nand2_2 _18898_ (.Y(_12032_),
    .A(_12029_),
    .B(net1027));
 sg13g2_or2_1 _18899_ (.X(_12033_),
    .B(_12032_),
    .A(_12028_));
 sg13g2_buf_2 _18900_ (.A(_12033_),
    .X(_12034_));
 sg13g2_or2_1 _18901_ (.X(_12035_),
    .B(_12034_),
    .A(_12023_));
 sg13g2_buf_1 _18902_ (.A(_12035_),
    .X(_12036_));
 sg13g2_mux2_1 _18903_ (.A0(net1110),
    .A1(\cpu.dcache.r_data[0][0] ),
    .S(_12036_),
    .X(_12037_));
 sg13g2_buf_1 _18904_ (.A(_08340_),
    .X(_12038_));
 sg13g2_nand2b_1 _18905_ (.Y(_12039_),
    .B(\cpu.ex.r_wmask[1] ),
    .A_N(net1026));
 sg13g2_buf_2 _18906_ (.A(_00259_),
    .X(_12040_));
 sg13g2_buf_1 _18907_ (.A(_12040_),
    .X(_12041_));
 sg13g2_o21ai_1 _18908_ (.B1(net1025),
    .Y(_12042_),
    .A1(_08341_),
    .A2(_12039_));
 sg13g2_buf_2 _18909_ (.A(_12042_),
    .X(_12043_));
 sg13g2_nor2_1 _18910_ (.A(_09400_),
    .B(_09465_),
    .Y(_12044_));
 sg13g2_buf_2 _18911_ (.A(_12044_),
    .X(_12045_));
 sg13g2_nand2_1 _18912_ (.Y(_12046_),
    .A(_12024_),
    .B(_12026_));
 sg13g2_buf_1 _18913_ (.A(\cpu.dcache.r_offset[2] ),
    .X(_12047_));
 sg13g2_nand2_1 _18914_ (.Y(_12048_),
    .A(_12047_),
    .B(_12029_));
 sg13g2_buf_1 _18915_ (.A(_12048_),
    .X(_12049_));
 sg13g2_or2_1 _18916_ (.X(_12050_),
    .B(_12049_),
    .A(_12046_));
 sg13g2_buf_2 _18917_ (.A(_12050_),
    .X(_12051_));
 sg13g2_nor2_1 _18918_ (.A(_09361_),
    .B(_08343_),
    .Y(_12052_));
 sg13g2_nand2_1 _18919_ (.Y(_12053_),
    .A(_09821_),
    .B(_12052_));
 sg13g2_a21oi_1 _18920_ (.A1(_11489_),
    .A2(_12051_),
    .Y(_12054_),
    .B1(_12053_));
 sg13g2_buf_2 _18921_ (.A(_12054_),
    .X(_12055_));
 sg13g2_nand2_1 _18922_ (.Y(_12056_),
    .A(_12045_),
    .B(_12055_));
 sg13g2_nor2_1 _18923_ (.A(_12043_),
    .B(_12056_),
    .Y(_12057_));
 sg13g2_buf_1 _18924_ (.A(_12057_),
    .X(_12058_));
 sg13g2_mux2_1 _18925_ (.A0(_12037_),
    .A1(net911),
    .S(_12058_),
    .X(_00310_));
 sg13g2_buf_1 _18926_ (.A(uio_in[2]),
    .X(_12059_));
 sg13g2_buf_1 _18927_ (.A(_12059_),
    .X(_12060_));
 sg13g2_or2_1 _18928_ (.X(_12061_),
    .B(_12032_),
    .A(_12046_));
 sg13g2_buf_2 _18929_ (.A(_12061_),
    .X(_12062_));
 sg13g2_or2_1 _18930_ (.X(_12063_),
    .B(_12062_),
    .A(_12023_));
 sg13g2_buf_1 _18931_ (.A(_12063_),
    .X(_12064_));
 sg13g2_mux2_1 _18932_ (.A0(net1109),
    .A1(\cpu.dcache.r_data[0][10] ),
    .S(_12064_),
    .X(_12065_));
 sg13g2_inv_1 _18933_ (.Y(_12066_),
    .A(\cpu.dcache.wdata[10] ));
 sg13g2_nor2_1 _18934_ (.A(_09242_),
    .B(_08340_),
    .Y(_12067_));
 sg13g2_nand2_1 _18935_ (.Y(_12068_),
    .A(_08341_),
    .B(_12067_));
 sg13g2_buf_1 _18936_ (.A(_12068_),
    .X(_12069_));
 sg13g2_buf_1 _18937_ (.A(_12069_),
    .X(_12070_));
 sg13g2_nand2_1 _18938_ (.Y(_12071_),
    .A(_10055_),
    .B(net671));
 sg13g2_o21ai_1 _18939_ (.B1(_12071_),
    .Y(_12072_),
    .A1(_12066_),
    .A2(net671));
 sg13g2_buf_2 _18940_ (.A(_12072_),
    .X(_12073_));
 sg13g2_buf_1 _18941_ (.A(_12073_),
    .X(_12074_));
 sg13g2_mux2_1 _18942_ (.A0(net685),
    .A1(_12040_),
    .S(_09243_),
    .X(_12075_));
 sg13g2_nand2_1 _18943_ (.Y(_12076_),
    .A(_12067_),
    .B(_12075_));
 sg13g2_buf_2 _18944_ (.A(_12076_),
    .X(_12077_));
 sg13g2_nor2_1 _18945_ (.A(_12056_),
    .B(_12077_),
    .Y(_12078_));
 sg13g2_buf_4 _18946_ (.X(_12079_),
    .A(_12078_));
 sg13g2_mux2_1 _18947_ (.A0(_12065_),
    .A1(net459),
    .S(_12079_),
    .X(_00311_));
 sg13g2_buf_1 _18948_ (.A(uio_in[3]),
    .X(_12080_));
 sg13g2_buf_1 _18949_ (.A(_12080_),
    .X(_12081_));
 sg13g2_mux2_1 _18950_ (.A0(net1108),
    .A1(\cpu.dcache.r_data[0][11] ),
    .S(_12064_),
    .X(_12082_));
 sg13g2_mux2_1 _18951_ (.A0(_10162_),
    .A1(net1128),
    .S(net671),
    .X(_12083_));
 sg13g2_buf_2 _18952_ (.A(_12083_),
    .X(_12084_));
 sg13g2_buf_1 _18953_ (.A(_12084_),
    .X(_12085_));
 sg13g2_mux2_1 _18954_ (.A0(_12082_),
    .A1(net509),
    .S(_12079_),
    .X(_00312_));
 sg13g2_nand2b_1 _18955_ (.Y(_12086_),
    .B(_12024_),
    .A_N(_12026_));
 sg13g2_buf_1 _18956_ (.A(_12086_),
    .X(_12087_));
 sg13g2_or2_1 _18957_ (.X(_12088_),
    .B(_12087_),
    .A(_12032_));
 sg13g2_buf_2 _18958_ (.A(_12088_),
    .X(_12089_));
 sg13g2_or2_1 _18959_ (.X(_12090_),
    .B(_12089_),
    .A(_12023_));
 sg13g2_buf_1 _18960_ (.A(_12090_),
    .X(_12091_));
 sg13g2_mux2_1 _18961_ (.A0(net1110),
    .A1(\cpu.dcache.r_data[0][12] ),
    .S(_12091_),
    .X(_12092_));
 sg13g2_inv_1 _18962_ (.Y(_12093_),
    .A(\cpu.dcache.wdata[12] ));
 sg13g2_nand2_1 _18963_ (.Y(_12094_),
    .A(_10066_),
    .B(_12069_));
 sg13g2_o21ai_1 _18964_ (.B1(_12094_),
    .Y(_12095_),
    .A1(_12093_),
    .A2(net671));
 sg13g2_buf_2 _18965_ (.A(_12095_),
    .X(_12096_));
 sg13g2_buf_1 _18966_ (.A(_12096_),
    .X(_12097_));
 sg13g2_mux2_1 _18967_ (.A0(_12092_),
    .A1(net508),
    .S(_12079_),
    .X(_00313_));
 sg13g2_buf_1 _18968_ (.A(uio_in[1]),
    .X(_12098_));
 sg13g2_buf_1 _18969_ (.A(_12098_),
    .X(_12099_));
 sg13g2_mux2_1 _18970_ (.A0(net1107),
    .A1(\cpu.dcache.r_data[0][13] ),
    .S(_12091_),
    .X(_12100_));
 sg13g2_inv_2 _18971_ (.Y(_12101_),
    .A(\cpu.dcache.wdata[13] ));
 sg13g2_nand2_1 _18972_ (.Y(_12102_),
    .A(_10072_),
    .B(_12069_));
 sg13g2_o21ai_1 _18973_ (.B1(_12102_),
    .Y(_12103_),
    .A1(_12101_),
    .A2(_12070_));
 sg13g2_buf_2 _18974_ (.A(_12103_),
    .X(_12104_));
 sg13g2_buf_1 _18975_ (.A(_12104_),
    .X(_12105_));
 sg13g2_mux2_1 _18976_ (.A0(_12100_),
    .A1(net507),
    .S(_12079_),
    .X(_00314_));
 sg13g2_mux2_1 _18977_ (.A0(net1109),
    .A1(\cpu.dcache.r_data[0][14] ),
    .S(_12091_),
    .X(_12106_));
 sg13g2_inv_2 _18978_ (.Y(_12107_),
    .A(\cpu.dcache.wdata[14] ));
 sg13g2_nand2_1 _18979_ (.Y(_12108_),
    .A(_10078_),
    .B(_12069_));
 sg13g2_o21ai_1 _18980_ (.B1(_12108_),
    .Y(_12109_),
    .A1(_12107_),
    .A2(_12070_));
 sg13g2_buf_2 _18981_ (.A(_12109_),
    .X(_12110_));
 sg13g2_buf_1 _18982_ (.A(_12110_),
    .X(_12111_));
 sg13g2_mux2_1 _18983_ (.A0(_12106_),
    .A1(net506),
    .S(_12079_),
    .X(_00315_));
 sg13g2_mux2_1 _18984_ (.A0(net1108),
    .A1(\cpu.dcache.r_data[0][15] ),
    .S(_12091_),
    .X(_12112_));
 sg13g2_inv_1 _18985_ (.Y(_12113_),
    .A(\cpu.dcache.wdata[15] ));
 sg13g2_nand2_1 _18986_ (.Y(_12114_),
    .A(_10081_),
    .B(_12069_));
 sg13g2_o21ai_1 _18987_ (.B1(_12114_),
    .Y(_12115_),
    .A1(_12113_),
    .A2(net671));
 sg13g2_buf_2 _18988_ (.A(_12115_),
    .X(_12116_));
 sg13g2_buf_1 _18989_ (.A(_12116_),
    .X(_12117_));
 sg13g2_mux2_1 _18990_ (.A0(_12112_),
    .A1(net505),
    .S(_12079_),
    .X(_00316_));
 sg13g2_nor2b_1 _18991_ (.A(_12024_),
    .B_N(_12026_),
    .Y(_12118_));
 sg13g2_nand2b_1 _18992_ (.Y(_12119_),
    .B(_12118_),
    .A_N(_12049_));
 sg13g2_buf_2 _18993_ (.A(_12119_),
    .X(_12120_));
 sg13g2_or2_1 _18994_ (.X(_12121_),
    .B(_12120_),
    .A(_12023_));
 sg13g2_buf_1 _18995_ (.A(_12121_),
    .X(_12122_));
 sg13g2_mux2_1 _18996_ (.A0(net1110),
    .A1(\cpu.dcache.r_data[0][16] ),
    .S(_12122_),
    .X(_12123_));
 sg13g2_buf_1 _18997_ (.A(net686),
    .X(_12124_));
 sg13g2_o21ai_1 _18998_ (.B1(net612),
    .Y(_12125_),
    .A1(_08341_),
    .A2(_12039_));
 sg13g2_buf_2 _18999_ (.A(_12125_),
    .X(_12126_));
 sg13g2_nor2_1 _19000_ (.A(_12056_),
    .B(_12126_),
    .Y(_12127_));
 sg13g2_buf_1 _19001_ (.A(_12127_),
    .X(_12128_));
 sg13g2_mux2_1 _19002_ (.A0(_12123_),
    .A1(_10099_),
    .S(_12128_),
    .X(_00317_));
 sg13g2_mux2_1 _19003_ (.A0(net1107),
    .A1(\cpu.dcache.r_data[0][17] ),
    .S(_12122_),
    .X(_12129_));
 sg13g2_buf_1 _19004_ (.A(net1061),
    .X(_12130_));
 sg13g2_mux2_1 _19005_ (.A0(_12129_),
    .A1(net885),
    .S(net78),
    .X(_00318_));
 sg13g2_mux2_1 _19006_ (.A0(net1109),
    .A1(\cpu.dcache.r_data[0][18] ),
    .S(_12122_),
    .X(_12131_));
 sg13g2_buf_1 _19007_ (.A(_10056_),
    .X(_12132_));
 sg13g2_mux2_1 _19008_ (.A0(_12131_),
    .A1(net884),
    .S(net78),
    .X(_00319_));
 sg13g2_mux2_1 _19009_ (.A0(net1108),
    .A1(\cpu.dcache.r_data[0][19] ),
    .S(_12122_),
    .X(_12133_));
 sg13g2_buf_1 _19010_ (.A(net1128),
    .X(_12134_));
 sg13g2_mux2_1 _19011_ (.A0(_12133_),
    .A1(net1024),
    .S(net78),
    .X(_00320_));
 sg13g2_mux2_1 _19012_ (.A0(net1107),
    .A1(\cpu.dcache.r_data[0][1] ),
    .S(_12036_),
    .X(_12135_));
 sg13g2_mux2_1 _19013_ (.A0(_12135_),
    .A1(net885),
    .S(net79),
    .X(_00321_));
 sg13g2_inv_1 _19014_ (.Y(_12136_),
    .A(_10066_));
 sg13g2_buf_1 _19015_ (.A(_12136_),
    .X(_12137_));
 sg13g2_buf_1 _19016_ (.A(net883),
    .X(_12138_));
 sg13g2_nor2_2 _19017_ (.A(_12024_),
    .B(_12026_),
    .Y(_12139_));
 sg13g2_nor2b_2 _19018_ (.A(_12049_),
    .B_N(_12139_),
    .Y(_12140_));
 sg13g2_nand2_2 _19019_ (.Y(_12141_),
    .A(_12045_),
    .B(_12140_));
 sg13g2_mux2_1 _19020_ (.A0(net1110),
    .A1(\cpu.dcache.r_data[0][20] ),
    .S(_12141_),
    .X(_12142_));
 sg13g2_nor2_1 _19021_ (.A(net78),
    .B(_12142_),
    .Y(_12143_));
 sg13g2_a21oi_1 _19022_ (.A1(net757),
    .A2(net78),
    .Y(_00322_),
    .B1(_12143_));
 sg13g2_inv_1 _19023_ (.Y(_12144_),
    .A(_10072_));
 sg13g2_buf_1 _19024_ (.A(_12144_),
    .X(_12145_));
 sg13g2_buf_1 _19025_ (.A(net882),
    .X(_12146_));
 sg13g2_mux2_1 _19026_ (.A0(net1107),
    .A1(\cpu.dcache.r_data[0][21] ),
    .S(_12141_),
    .X(_12147_));
 sg13g2_nor2_1 _19027_ (.A(net78),
    .B(_12147_),
    .Y(_12148_));
 sg13g2_a21oi_1 _19028_ (.A1(_12146_),
    .A2(net78),
    .Y(_00323_),
    .B1(_12148_));
 sg13g2_inv_1 _19029_ (.Y(_12149_),
    .A(_10078_));
 sg13g2_buf_1 _19030_ (.A(_12149_),
    .X(_12150_));
 sg13g2_buf_1 _19031_ (.A(net881),
    .X(_12151_));
 sg13g2_mux2_1 _19032_ (.A0(net1109),
    .A1(\cpu.dcache.r_data[0][22] ),
    .S(_12141_),
    .X(_12152_));
 sg13g2_nor2_1 _19033_ (.A(_12127_),
    .B(_12152_),
    .Y(_12153_));
 sg13g2_a21oi_1 _19034_ (.A1(net755),
    .A2(net78),
    .Y(_00324_),
    .B1(_12153_));
 sg13g2_mux2_1 _19035_ (.A0(net1108),
    .A1(\cpu.dcache.r_data[0][23] ),
    .S(_12141_),
    .X(_12154_));
 sg13g2_buf_1 _19036_ (.A(_10081_),
    .X(_12155_));
 sg13g2_mux2_1 _19037_ (.A0(_12154_),
    .A1(net1023),
    .S(_12128_),
    .X(_00325_));
 sg13g2_nor2_1 _19038_ (.A(_12046_),
    .B(_12049_),
    .Y(_12156_));
 sg13g2_nand2_1 _19039_ (.Y(_12157_),
    .A(_12045_),
    .B(_12156_));
 sg13g2_buf_1 _19040_ (.A(_12157_),
    .X(_12158_));
 sg13g2_mux2_1 _19041_ (.A0(_12021_),
    .A1(\cpu.dcache.r_data[0][24] ),
    .S(net611),
    .X(_12159_));
 sg13g2_mux2_1 _19042_ (.A0(_10146_),
    .A1(_10032_),
    .S(net671),
    .X(_12160_));
 sg13g2_buf_2 _19043_ (.A(_12160_),
    .X(_12161_));
 sg13g2_buf_1 _19044_ (.A(_12161_),
    .X(_12162_));
 sg13g2_nor2_1 _19045_ (.A(_08341_),
    .B(net686),
    .Y(_12163_));
 sg13g2_a21oi_1 _19046_ (.A1(_08341_),
    .A2(_12040_),
    .Y(_12164_),
    .B1(_12163_));
 sg13g2_nand2_1 _19047_ (.Y(_12165_),
    .A(_12067_),
    .B(_12164_));
 sg13g2_buf_2 _19048_ (.A(_12165_),
    .X(_12166_));
 sg13g2_nor2_1 _19049_ (.A(_12056_),
    .B(_12166_),
    .Y(_12167_));
 sg13g2_buf_4 _19050_ (.X(_12168_),
    .A(_12167_));
 sg13g2_mux2_1 _19051_ (.A0(_12159_),
    .A1(net504),
    .S(_12168_),
    .X(_00326_));
 sg13g2_mux2_1 _19052_ (.A0(_12099_),
    .A1(\cpu.dcache.r_data[0][25] ),
    .S(net611),
    .X(_12169_));
 sg13g2_inv_1 _19053_ (.Y(_12170_),
    .A(\cpu.dcache.wdata[9] ));
 sg13g2_nand2_1 _19054_ (.Y(_12171_),
    .A(_10050_),
    .B(net671));
 sg13g2_o21ai_1 _19055_ (.B1(_12171_),
    .Y(_12172_),
    .A1(_12170_),
    .A2(net671));
 sg13g2_buf_2 _19056_ (.A(_12172_),
    .X(_12173_));
 sg13g2_buf_1 _19057_ (.A(_12173_),
    .X(_12174_));
 sg13g2_mux2_1 _19058_ (.A0(_12169_),
    .A1(net458),
    .S(_12168_),
    .X(_00327_));
 sg13g2_mux2_1 _19059_ (.A0(_12060_),
    .A1(\cpu.dcache.r_data[0][26] ),
    .S(net611),
    .X(_12175_));
 sg13g2_mux2_1 _19060_ (.A0(_12175_),
    .A1(net459),
    .S(_12168_),
    .X(_00328_));
 sg13g2_mux2_1 _19061_ (.A0(_12081_),
    .A1(\cpu.dcache.r_data[0][27] ),
    .S(_12157_),
    .X(_12176_));
 sg13g2_mux2_1 _19062_ (.A0(_12176_),
    .A1(net509),
    .S(_12168_),
    .X(_00329_));
 sg13g2_or2_1 _19063_ (.X(_12177_),
    .B(_12087_),
    .A(_12049_));
 sg13g2_buf_2 _19064_ (.A(_12177_),
    .X(_12178_));
 sg13g2_or2_1 _19065_ (.X(_12179_),
    .B(_12178_),
    .A(_12023_));
 sg13g2_buf_1 _19066_ (.A(_12179_),
    .X(_12180_));
 sg13g2_mux2_1 _19067_ (.A0(net1110),
    .A1(\cpu.dcache.r_data[0][28] ),
    .S(_12180_),
    .X(_12181_));
 sg13g2_mux2_1 _19068_ (.A0(_12181_),
    .A1(net508),
    .S(_12168_),
    .X(_00330_));
 sg13g2_mux2_1 _19069_ (.A0(_12099_),
    .A1(\cpu.dcache.r_data[0][29] ),
    .S(_12180_),
    .X(_12182_));
 sg13g2_mux2_1 _19070_ (.A0(_12182_),
    .A1(net507),
    .S(_12168_),
    .X(_00331_));
 sg13g2_mux2_1 _19071_ (.A0(net1109),
    .A1(\cpu.dcache.r_data[0][2] ),
    .S(_12036_),
    .X(_12183_));
 sg13g2_mux2_1 _19072_ (.A0(_12183_),
    .A1(net884),
    .S(_12058_),
    .X(_00332_));
 sg13g2_mux2_1 _19073_ (.A0(net1109),
    .A1(\cpu.dcache.r_data[0][30] ),
    .S(_12180_),
    .X(_12184_));
 sg13g2_mux2_1 _19074_ (.A0(_12184_),
    .A1(net506),
    .S(_12168_),
    .X(_00333_));
 sg13g2_mux2_1 _19075_ (.A0(_12081_),
    .A1(\cpu.dcache.r_data[0][31] ),
    .S(_12180_),
    .X(_12185_));
 sg13g2_mux2_1 _19076_ (.A0(_12185_),
    .A1(_12117_),
    .S(_12168_),
    .X(_00334_));
 sg13g2_mux2_1 _19077_ (.A0(net1108),
    .A1(\cpu.dcache.r_data[0][3] ),
    .S(_12036_),
    .X(_12186_));
 sg13g2_mux2_1 _19078_ (.A0(_12186_),
    .A1(net1024),
    .S(net79),
    .X(_00335_));
 sg13g2_nor2b_2 _19079_ (.A(_12032_),
    .B_N(_12139_),
    .Y(_12187_));
 sg13g2_nand2_2 _19080_ (.Y(_12188_),
    .A(_12045_),
    .B(_12187_));
 sg13g2_mux2_1 _19081_ (.A0(net1110),
    .A1(\cpu.dcache.r_data[0][4] ),
    .S(_12188_),
    .X(_12189_));
 sg13g2_nor2_1 _19082_ (.A(net79),
    .B(_12189_),
    .Y(_12190_));
 sg13g2_a21oi_1 _19083_ (.A1(_12138_),
    .A2(net79),
    .Y(_00336_),
    .B1(_12190_));
 sg13g2_mux2_1 _19084_ (.A0(net1107),
    .A1(\cpu.dcache.r_data[0][5] ),
    .S(_12188_),
    .X(_12191_));
 sg13g2_nor2_1 _19085_ (.A(net79),
    .B(_12191_),
    .Y(_12192_));
 sg13g2_a21oi_1 _19086_ (.A1(_12146_),
    .A2(net79),
    .Y(_00337_),
    .B1(_12192_));
 sg13g2_mux2_1 _19087_ (.A0(net1109),
    .A1(\cpu.dcache.r_data[0][6] ),
    .S(_12188_),
    .X(_12193_));
 sg13g2_nor2_1 _19088_ (.A(_12057_),
    .B(_12193_),
    .Y(_12194_));
 sg13g2_a21oi_1 _19089_ (.A1(net755),
    .A2(net79),
    .Y(_00338_),
    .B1(_12194_));
 sg13g2_mux2_1 _19090_ (.A0(net1108),
    .A1(\cpu.dcache.r_data[0][7] ),
    .S(_12188_),
    .X(_12195_));
 sg13g2_mux2_1 _19091_ (.A0(_12195_),
    .A1(net1023),
    .S(net79),
    .X(_00339_));
 sg13g2_mux2_1 _19092_ (.A0(net1110),
    .A1(\cpu.dcache.r_data[0][8] ),
    .S(_12064_),
    .X(_12196_));
 sg13g2_mux2_1 _19093_ (.A0(_12196_),
    .A1(net504),
    .S(_12079_),
    .X(_00340_));
 sg13g2_mux2_1 _19094_ (.A0(net1107),
    .A1(\cpu.dcache.r_data[0][9] ),
    .S(_12064_),
    .X(_12197_));
 sg13g2_mux2_1 _19095_ (.A0(_12197_),
    .A1(net458),
    .S(_12079_),
    .X(_00341_));
 sg13g2_buf_1 _19096_ (.A(net627),
    .X(_12198_));
 sg13g2_buf_1 _19097_ (.A(net562),
    .X(_12199_));
 sg13g2_nand2_1 _19098_ (.Y(_12200_),
    .A(net503),
    .B(_12055_));
 sg13g2_nor2_1 _19099_ (.A(_12043_),
    .B(_12200_),
    .Y(_12201_));
 sg13g2_buf_1 _19100_ (.A(_12201_),
    .X(_12202_));
 sg13g2_buf_1 _19101_ (.A(_12202_),
    .X(_12203_));
 sg13g2_buf_1 _19102_ (.A(_12020_),
    .X(_12204_));
 sg13g2_buf_2 _19103_ (.A(net1106),
    .X(_12205_));
 sg13g2_nand2_1 _19104_ (.Y(_12206_),
    .A(net916),
    .B(_09416_));
 sg13g2_buf_1 _19105_ (.A(_12206_),
    .X(_12207_));
 sg13g2_nor2_1 _19106_ (.A(net670),
    .B(_12034_),
    .Y(_12208_));
 sg13g2_buf_2 _19107_ (.A(_12208_),
    .X(_12209_));
 sg13g2_nor2b_1 _19108_ (.A(_12209_),
    .B_N(\cpu.dcache.r_data[1][0] ),
    .Y(_12210_));
 sg13g2_a21oi_1 _19109_ (.A1(net1022),
    .A2(_12209_),
    .Y(_12211_),
    .B1(_12210_));
 sg13g2_buf_1 _19110_ (.A(_10033_),
    .X(_12212_));
 sg13g2_nand2_1 _19111_ (.Y(_12213_),
    .A(net880),
    .B(net63));
 sg13g2_o21ai_1 _19112_ (.B1(_12213_),
    .Y(_00342_),
    .A1(net63),
    .A2(_12211_));
 sg13g2_nor2_1 _19113_ (.A(_12077_),
    .B(_12200_),
    .Y(_12214_));
 sg13g2_buf_2 _19114_ (.A(_12214_),
    .X(_12215_));
 sg13g2_buf_1 _19115_ (.A(_12215_),
    .X(_12216_));
 sg13g2_buf_1 _19116_ (.A(_12059_),
    .X(_12217_));
 sg13g2_buf_2 _19117_ (.A(net1105),
    .X(_12218_));
 sg13g2_nor2_1 _19118_ (.A(net670),
    .B(_12062_),
    .Y(_12219_));
 sg13g2_buf_2 _19119_ (.A(_12219_),
    .X(_12220_));
 sg13g2_nor2b_1 _19120_ (.A(_12220_),
    .B_N(\cpu.dcache.r_data[1][10] ),
    .Y(_12221_));
 sg13g2_a21oi_1 _19121_ (.A1(net1021),
    .A2(_12220_),
    .Y(_12222_),
    .B1(_12221_));
 sg13g2_nand2_1 _19122_ (.Y(_12223_),
    .A(net459),
    .B(net62));
 sg13g2_o21ai_1 _19123_ (.B1(_12223_),
    .Y(_00343_),
    .A1(net62),
    .A2(_12222_));
 sg13g2_buf_1 _19124_ (.A(_12080_),
    .X(_12224_));
 sg13g2_buf_2 _19125_ (.A(net1104),
    .X(_12225_));
 sg13g2_nor2b_1 _19126_ (.A(_12220_),
    .B_N(\cpu.dcache.r_data[1][11] ),
    .Y(_12226_));
 sg13g2_a21oi_1 _19127_ (.A1(net1020),
    .A2(_12220_),
    .Y(_12227_),
    .B1(_12226_));
 sg13g2_nand2_1 _19128_ (.Y(_12228_),
    .A(_12085_),
    .B(net62));
 sg13g2_o21ai_1 _19129_ (.B1(_12228_),
    .Y(_00344_),
    .A1(net62),
    .A2(_12227_));
 sg13g2_nor2_1 _19130_ (.A(net670),
    .B(_12089_),
    .Y(_12229_));
 sg13g2_buf_2 _19131_ (.A(_12229_),
    .X(_12230_));
 sg13g2_inv_1 _19132_ (.Y(_12231_),
    .A(\cpu.dcache.r_data[1][12] ));
 sg13g2_nor2_1 _19133_ (.A(_12231_),
    .B(_12230_),
    .Y(_12232_));
 sg13g2_a21oi_1 _19134_ (.A1(net1022),
    .A2(_12230_),
    .Y(_12233_),
    .B1(_12232_));
 sg13g2_nand2_1 _19135_ (.Y(_12234_),
    .A(_12097_),
    .B(_12215_));
 sg13g2_o21ai_1 _19136_ (.B1(_12234_),
    .Y(_00345_),
    .A1(_12216_),
    .A2(_12233_));
 sg13g2_buf_1 _19137_ (.A(_12098_),
    .X(_12235_));
 sg13g2_buf_2 _19138_ (.A(net1103),
    .X(_12236_));
 sg13g2_nor2b_1 _19139_ (.A(_12230_),
    .B_N(\cpu.dcache.r_data[1][13] ),
    .Y(_12237_));
 sg13g2_a21oi_1 _19140_ (.A1(net1019),
    .A2(_12230_),
    .Y(_12238_),
    .B1(_12237_));
 sg13g2_nand2_1 _19141_ (.Y(_12239_),
    .A(_12105_),
    .B(_12215_));
 sg13g2_o21ai_1 _19142_ (.B1(_12239_),
    .Y(_00346_),
    .A1(_12216_),
    .A2(_12238_));
 sg13g2_nor2b_1 _19143_ (.A(_12230_),
    .B_N(\cpu.dcache.r_data[1][14] ),
    .Y(_12240_));
 sg13g2_a21oi_1 _19144_ (.A1(net1021),
    .A2(_12230_),
    .Y(_12241_),
    .B1(_12240_));
 sg13g2_nand2_1 _19145_ (.Y(_12242_),
    .A(_12111_),
    .B(_12215_));
 sg13g2_o21ai_1 _19146_ (.B1(_12242_),
    .Y(_00347_),
    .A1(net62),
    .A2(_12241_));
 sg13g2_nor2b_1 _19147_ (.A(_12230_),
    .B_N(\cpu.dcache.r_data[1][15] ),
    .Y(_12243_));
 sg13g2_a21oi_1 _19148_ (.A1(net1020),
    .A2(_12230_),
    .Y(_12244_),
    .B1(_12243_));
 sg13g2_nand2_1 _19149_ (.Y(_12245_),
    .A(_12117_),
    .B(_12215_));
 sg13g2_o21ai_1 _19150_ (.B1(_12245_),
    .Y(_00348_),
    .A1(net62),
    .A2(_12244_));
 sg13g2_nor2_1 _19151_ (.A(_12126_),
    .B(_12200_),
    .Y(_12246_));
 sg13g2_buf_2 _19152_ (.A(_12246_),
    .X(_12247_));
 sg13g2_buf_1 _19153_ (.A(_12247_),
    .X(_12248_));
 sg13g2_nor2_1 _19154_ (.A(net670),
    .B(_12120_),
    .Y(_12249_));
 sg13g2_buf_2 _19155_ (.A(_12249_),
    .X(_12250_));
 sg13g2_nor2b_1 _19156_ (.A(_12250_),
    .B_N(\cpu.dcache.r_data[1][16] ),
    .Y(_12251_));
 sg13g2_a21oi_1 _19157_ (.A1(net1022),
    .A2(_12250_),
    .Y(_12252_),
    .B1(_12251_));
 sg13g2_nand2_1 _19158_ (.Y(_12253_),
    .A(net880),
    .B(_12248_));
 sg13g2_o21ai_1 _19159_ (.B1(_12253_),
    .Y(_00349_),
    .A1(net61),
    .A2(_12252_));
 sg13g2_nor2b_1 _19160_ (.A(_12250_),
    .B_N(\cpu.dcache.r_data[1][17] ),
    .Y(_12254_));
 sg13g2_a21oi_1 _19161_ (.A1(net1019),
    .A2(_12250_),
    .Y(_12255_),
    .B1(_12254_));
 sg13g2_nand2_1 _19162_ (.Y(_12256_),
    .A(net885),
    .B(net61));
 sg13g2_o21ai_1 _19163_ (.B1(_12256_),
    .Y(_00350_),
    .A1(net61),
    .A2(_12255_));
 sg13g2_nor2b_1 _19164_ (.A(_12250_),
    .B_N(\cpu.dcache.r_data[1][18] ),
    .Y(_12257_));
 sg13g2_a21oi_1 _19165_ (.A1(net1021),
    .A2(_12250_),
    .Y(_12258_),
    .B1(_12257_));
 sg13g2_nand2_1 _19166_ (.Y(_12259_),
    .A(net884),
    .B(_12247_));
 sg13g2_o21ai_1 _19167_ (.B1(_12259_),
    .Y(_00351_),
    .A1(net61),
    .A2(_12258_));
 sg13g2_nor2b_1 _19168_ (.A(_12250_),
    .B_N(\cpu.dcache.r_data[1][19] ),
    .Y(_12260_));
 sg13g2_a21oi_1 _19169_ (.A1(net1020),
    .A2(_12250_),
    .Y(_12261_),
    .B1(_12260_));
 sg13g2_nand2_1 _19170_ (.Y(_12262_),
    .A(net1024),
    .B(_12247_));
 sg13g2_o21ai_1 _19171_ (.B1(_12262_),
    .Y(_00352_),
    .A1(_12248_),
    .A2(_12261_));
 sg13g2_nor2b_1 _19172_ (.A(_12209_),
    .B_N(\cpu.dcache.r_data[1][1] ),
    .Y(_12263_));
 sg13g2_a21oi_1 _19173_ (.A1(net1019),
    .A2(_12209_),
    .Y(_12264_),
    .B1(_12263_));
 sg13g2_nand2_1 _19174_ (.Y(_12265_),
    .A(_12130_),
    .B(_12203_));
 sg13g2_o21ai_1 _19175_ (.B1(_12265_),
    .Y(_00353_),
    .A1(_12203_),
    .A2(_12264_));
 sg13g2_buf_1 _19176_ (.A(_12020_),
    .X(_12266_));
 sg13g2_nand2b_1 _19177_ (.Y(_12267_),
    .B(_12139_),
    .A_N(_12049_));
 sg13g2_buf_1 _19178_ (.A(_12267_),
    .X(_12268_));
 sg13g2_nor2_1 _19179_ (.A(net670),
    .B(_12268_),
    .Y(_12269_));
 sg13g2_buf_2 _19180_ (.A(_12269_),
    .X(_12270_));
 sg13g2_mux2_1 _19181_ (.A0(\cpu.dcache.r_data[1][20] ),
    .A1(_12266_),
    .S(_12270_),
    .X(_12271_));
 sg13g2_nor2_1 _19182_ (.A(_12247_),
    .B(_12271_),
    .Y(_12272_));
 sg13g2_a21oi_1 _19183_ (.A1(net757),
    .A2(net61),
    .Y(_00354_),
    .B1(_12272_));
 sg13g2_buf_1 _19184_ (.A(_12098_),
    .X(_12273_));
 sg13g2_mux2_1 _19185_ (.A0(\cpu.dcache.r_data[1][21] ),
    .A1(_12273_),
    .S(_12270_),
    .X(_12274_));
 sg13g2_nor2_1 _19186_ (.A(_12247_),
    .B(_12274_),
    .Y(_12275_));
 sg13g2_a21oi_1 _19187_ (.A1(net756),
    .A2(net61),
    .Y(_00355_),
    .B1(_12275_));
 sg13g2_buf_1 _19188_ (.A(_12059_),
    .X(_12276_));
 sg13g2_mux2_1 _19189_ (.A0(\cpu.dcache.r_data[1][22] ),
    .A1(_12276_),
    .S(_12270_),
    .X(_12277_));
 sg13g2_nor2_1 _19190_ (.A(_12247_),
    .B(_12277_),
    .Y(_12278_));
 sg13g2_a21oi_1 _19191_ (.A1(net755),
    .A2(net61),
    .Y(_00356_),
    .B1(_12278_));
 sg13g2_nor2b_1 _19192_ (.A(_12270_),
    .B_N(\cpu.dcache.r_data[1][23] ),
    .Y(_12279_));
 sg13g2_a21oi_1 _19193_ (.A1(net1020),
    .A2(_12270_),
    .Y(_12280_),
    .B1(_12279_));
 sg13g2_buf_1 _19194_ (.A(_10081_),
    .X(_12281_));
 sg13g2_nand2_1 _19195_ (.Y(_12282_),
    .A(net1018),
    .B(_12247_));
 sg13g2_o21ai_1 _19196_ (.B1(_12282_),
    .Y(_00357_),
    .A1(net61),
    .A2(_12280_));
 sg13g2_nor2_1 _19197_ (.A(_12166_),
    .B(_12200_),
    .Y(_12283_));
 sg13g2_buf_2 _19198_ (.A(_12283_),
    .X(_12284_));
 sg13g2_buf_1 _19199_ (.A(_12284_),
    .X(_12285_));
 sg13g2_nor2_1 _19200_ (.A(net670),
    .B(_12051_),
    .Y(_12286_));
 sg13g2_buf_1 _19201_ (.A(_12286_),
    .X(_12287_));
 sg13g2_nor2b_1 _19202_ (.A(net561),
    .B_N(\cpu.dcache.r_data[1][24] ),
    .Y(_12288_));
 sg13g2_a21oi_1 _19203_ (.A1(net1022),
    .A2(net561),
    .Y(_12289_),
    .B1(_12288_));
 sg13g2_nand2_1 _19204_ (.Y(_12290_),
    .A(net504),
    .B(net60));
 sg13g2_o21ai_1 _19205_ (.B1(_12290_),
    .Y(_00358_),
    .A1(net60),
    .A2(_12289_));
 sg13g2_nor2b_1 _19206_ (.A(net561),
    .B_N(\cpu.dcache.r_data[1][25] ),
    .Y(_12291_));
 sg13g2_a21oi_1 _19207_ (.A1(net1019),
    .A2(net561),
    .Y(_12292_),
    .B1(_12291_));
 sg13g2_nand2_1 _19208_ (.Y(_12293_),
    .A(_12174_),
    .B(net60));
 sg13g2_o21ai_1 _19209_ (.B1(_12293_),
    .Y(_00359_),
    .A1(net60),
    .A2(_12292_));
 sg13g2_nor2b_1 _19210_ (.A(net561),
    .B_N(\cpu.dcache.r_data[1][26] ),
    .Y(_12294_));
 sg13g2_a21oi_1 _19211_ (.A1(net1021),
    .A2(net561),
    .Y(_12295_),
    .B1(_12294_));
 sg13g2_nand2_1 _19212_ (.Y(_12296_),
    .A(_12074_),
    .B(_12284_));
 sg13g2_o21ai_1 _19213_ (.B1(_12296_),
    .Y(_00360_),
    .A1(net60),
    .A2(_12295_));
 sg13g2_nor2b_1 _19214_ (.A(net561),
    .B_N(\cpu.dcache.r_data[1][27] ),
    .Y(_12297_));
 sg13g2_a21oi_1 _19215_ (.A1(net1020),
    .A2(net561),
    .Y(_12298_),
    .B1(_12297_));
 sg13g2_nand2_1 _19216_ (.Y(_12299_),
    .A(net509),
    .B(_12284_));
 sg13g2_o21ai_1 _19217_ (.B1(_12299_),
    .Y(_00361_),
    .A1(net60),
    .A2(_12298_));
 sg13g2_nor2_1 _19218_ (.A(net670),
    .B(_12178_),
    .Y(_12300_));
 sg13g2_buf_2 _19219_ (.A(_12300_),
    .X(_12301_));
 sg13g2_nor2b_1 _19220_ (.A(_12301_),
    .B_N(\cpu.dcache.r_data[1][28] ),
    .Y(_12302_));
 sg13g2_a21oi_1 _19221_ (.A1(net1022),
    .A2(_12301_),
    .Y(_12303_),
    .B1(_12302_));
 sg13g2_nand2_1 _19222_ (.Y(_12304_),
    .A(_12097_),
    .B(_12284_));
 sg13g2_o21ai_1 _19223_ (.B1(_12304_),
    .Y(_00362_),
    .A1(_12285_),
    .A2(_12303_));
 sg13g2_nor2b_1 _19224_ (.A(_12301_),
    .B_N(\cpu.dcache.r_data[1][29] ),
    .Y(_12305_));
 sg13g2_a21oi_1 _19225_ (.A1(net1019),
    .A2(_12301_),
    .Y(_12306_),
    .B1(_12305_));
 sg13g2_nand2_1 _19226_ (.Y(_12307_),
    .A(net507),
    .B(_12284_));
 sg13g2_o21ai_1 _19227_ (.B1(_12307_),
    .Y(_00363_),
    .A1(net60),
    .A2(_12306_));
 sg13g2_nor2b_1 _19228_ (.A(_12209_),
    .B_N(\cpu.dcache.r_data[1][2] ),
    .Y(_12308_));
 sg13g2_a21oi_1 _19229_ (.A1(net1021),
    .A2(_12209_),
    .Y(_12309_),
    .B1(_12308_));
 sg13g2_nand2_1 _19230_ (.Y(_12310_),
    .A(_12132_),
    .B(_12202_));
 sg13g2_o21ai_1 _19231_ (.B1(_12310_),
    .Y(_00364_),
    .A1(net63),
    .A2(_12309_));
 sg13g2_nor2b_1 _19232_ (.A(_12301_),
    .B_N(\cpu.dcache.r_data[1][30] ),
    .Y(_12311_));
 sg13g2_a21oi_1 _19233_ (.A1(net1021),
    .A2(_12301_),
    .Y(_12312_),
    .B1(_12311_));
 sg13g2_nand2_1 _19234_ (.Y(_12313_),
    .A(_12111_),
    .B(_12284_));
 sg13g2_o21ai_1 _19235_ (.B1(_12313_),
    .Y(_00365_),
    .A1(_12285_),
    .A2(_12312_));
 sg13g2_nor2b_1 _19236_ (.A(_12301_),
    .B_N(\cpu.dcache.r_data[1][31] ),
    .Y(_12314_));
 sg13g2_a21oi_1 _19237_ (.A1(net1020),
    .A2(_12301_),
    .Y(_12315_),
    .B1(_12314_));
 sg13g2_nand2_1 _19238_ (.Y(_12316_),
    .A(net505),
    .B(_12284_));
 sg13g2_o21ai_1 _19239_ (.B1(_12316_),
    .Y(_00366_),
    .A1(net60),
    .A2(_12315_));
 sg13g2_buf_1 _19240_ (.A(_12224_),
    .X(_12317_));
 sg13g2_nor2b_1 _19241_ (.A(_12209_),
    .B_N(\cpu.dcache.r_data[1][3] ),
    .Y(_12318_));
 sg13g2_a21oi_1 _19242_ (.A1(net1017),
    .A2(_12209_),
    .Y(_12319_),
    .B1(_12318_));
 sg13g2_nand2_1 _19243_ (.Y(_12320_),
    .A(net1024),
    .B(_12202_));
 sg13g2_o21ai_1 _19244_ (.B1(_12320_),
    .Y(_00367_),
    .A1(net63),
    .A2(_12319_));
 sg13g2_nand2b_1 _19245_ (.Y(_12321_),
    .B(_12139_),
    .A_N(_12032_));
 sg13g2_buf_1 _19246_ (.A(_12321_),
    .X(_12322_));
 sg13g2_nor2_1 _19247_ (.A(net670),
    .B(_12322_),
    .Y(_12323_));
 sg13g2_buf_1 _19248_ (.A(_12323_),
    .X(_12324_));
 sg13g2_mux2_1 _19249_ (.A0(\cpu.dcache.r_data[1][4] ),
    .A1(_12266_),
    .S(_12324_),
    .X(_12325_));
 sg13g2_nor2_1 _19250_ (.A(_12202_),
    .B(_12325_),
    .Y(_12326_));
 sg13g2_a21oi_1 _19251_ (.A1(net757),
    .A2(net63),
    .Y(_00368_),
    .B1(_12326_));
 sg13g2_mux2_1 _19252_ (.A0(\cpu.dcache.r_data[1][5] ),
    .A1(net1101),
    .S(_12324_),
    .X(_12327_));
 sg13g2_nor2_1 _19253_ (.A(_12202_),
    .B(_12327_),
    .Y(_12328_));
 sg13g2_a21oi_1 _19254_ (.A1(net756),
    .A2(net63),
    .Y(_00369_),
    .B1(_12328_));
 sg13g2_mux2_1 _19255_ (.A0(\cpu.dcache.r_data[1][6] ),
    .A1(net1100),
    .S(_12324_),
    .X(_12329_));
 sg13g2_nor2_1 _19256_ (.A(_12202_),
    .B(_12329_),
    .Y(_12330_));
 sg13g2_a21oi_1 _19257_ (.A1(_12151_),
    .A2(net63),
    .Y(_00370_),
    .B1(_12330_));
 sg13g2_nor2b_1 _19258_ (.A(_12324_),
    .B_N(\cpu.dcache.r_data[1][7] ),
    .Y(_12331_));
 sg13g2_a21oi_1 _19259_ (.A1(net1017),
    .A2(_12324_),
    .Y(_12332_),
    .B1(_12331_));
 sg13g2_nand2_1 _19260_ (.Y(_12333_),
    .A(net1018),
    .B(_12202_));
 sg13g2_o21ai_1 _19261_ (.B1(_12333_),
    .Y(_00371_),
    .A1(net63),
    .A2(_12332_));
 sg13g2_nor2b_1 _19262_ (.A(_12220_),
    .B_N(\cpu.dcache.r_data[1][8] ),
    .Y(_12334_));
 sg13g2_a21oi_1 _19263_ (.A1(net1022),
    .A2(_12220_),
    .Y(_12335_),
    .B1(_12334_));
 sg13g2_nand2_1 _19264_ (.Y(_12336_),
    .A(_12162_),
    .B(_12215_));
 sg13g2_o21ai_1 _19265_ (.B1(_12336_),
    .Y(_00372_),
    .A1(net62),
    .A2(_12335_));
 sg13g2_nor2b_1 _19266_ (.A(_12220_),
    .B_N(\cpu.dcache.r_data[1][9] ),
    .Y(_12337_));
 sg13g2_a21oi_1 _19267_ (.A1(net1019),
    .A2(_12220_),
    .Y(_12338_),
    .B1(_12337_));
 sg13g2_nand2_1 _19268_ (.Y(_12339_),
    .A(net458),
    .B(_12215_));
 sg13g2_o21ai_1 _19269_ (.B1(_12339_),
    .Y(_00373_),
    .A1(net62),
    .A2(_12338_));
 sg13g2_buf_1 _19270_ (.A(_09413_),
    .X(_12340_));
 sg13g2_buf_1 _19271_ (.A(net610),
    .X(_12341_));
 sg13g2_buf_1 _19272_ (.A(net560),
    .X(_12342_));
 sg13g2_nand2_1 _19273_ (.Y(_12343_),
    .A(net502),
    .B(_12055_));
 sg13g2_nor2_1 _19274_ (.A(_12043_),
    .B(_12343_),
    .Y(_12344_));
 sg13g2_buf_2 _19275_ (.A(_12344_),
    .X(_12345_));
 sg13g2_buf_1 _19276_ (.A(_12345_),
    .X(_12346_));
 sg13g2_buf_1 _19277_ (.A(net1106),
    .X(_12347_));
 sg13g2_buf_1 _19278_ (.A(_09613_),
    .X(_12348_));
 sg13g2_nor2_1 _19279_ (.A(net669),
    .B(_12034_),
    .Y(_12349_));
 sg13g2_buf_2 _19280_ (.A(_12349_),
    .X(_12350_));
 sg13g2_nor2b_1 _19281_ (.A(_12350_),
    .B_N(\cpu.dcache.r_data[2][0] ),
    .Y(_12351_));
 sg13g2_a21oi_1 _19282_ (.A1(net1016),
    .A2(_12350_),
    .Y(_12352_),
    .B1(_12351_));
 sg13g2_nand2_1 _19283_ (.Y(_12353_),
    .A(net880),
    .B(net59));
 sg13g2_o21ai_1 _19284_ (.B1(_12353_),
    .Y(_00374_),
    .A1(net59),
    .A2(_12352_));
 sg13g2_nor2_1 _19285_ (.A(_12077_),
    .B(_12343_),
    .Y(_12354_));
 sg13g2_buf_2 _19286_ (.A(_12354_),
    .X(_12355_));
 sg13g2_buf_1 _19287_ (.A(_12355_),
    .X(_12356_));
 sg13g2_buf_1 _19288_ (.A(net1105),
    .X(_12357_));
 sg13g2_nor2_1 _19289_ (.A(net669),
    .B(_12062_),
    .Y(_12358_));
 sg13g2_buf_2 _19290_ (.A(_12358_),
    .X(_12359_));
 sg13g2_nor2b_1 _19291_ (.A(_12359_),
    .B_N(\cpu.dcache.r_data[2][10] ),
    .Y(_12360_));
 sg13g2_a21oi_1 _19292_ (.A1(net1015),
    .A2(_12359_),
    .Y(_12361_),
    .B1(_12360_));
 sg13g2_nand2_1 _19293_ (.Y(_12362_),
    .A(net459),
    .B(net58));
 sg13g2_o21ai_1 _19294_ (.B1(_12362_),
    .Y(_00375_),
    .A1(net58),
    .A2(_12361_));
 sg13g2_nor2b_1 _19295_ (.A(_12359_),
    .B_N(\cpu.dcache.r_data[2][11] ),
    .Y(_12363_));
 sg13g2_a21oi_1 _19296_ (.A1(net1017),
    .A2(_12359_),
    .Y(_12364_),
    .B1(_12363_));
 sg13g2_nand2_1 _19297_ (.Y(_12365_),
    .A(_12085_),
    .B(net58));
 sg13g2_o21ai_1 _19298_ (.B1(_12365_),
    .Y(_00376_),
    .A1(net58),
    .A2(_12364_));
 sg13g2_nor2_1 _19299_ (.A(net669),
    .B(_12089_),
    .Y(_12366_));
 sg13g2_buf_2 _19300_ (.A(_12366_),
    .X(_12367_));
 sg13g2_nor2b_1 _19301_ (.A(_12367_),
    .B_N(\cpu.dcache.r_data[2][12] ),
    .Y(_12368_));
 sg13g2_a21oi_1 _19302_ (.A1(_12347_),
    .A2(_12367_),
    .Y(_12369_),
    .B1(_12368_));
 sg13g2_nand2_1 _19303_ (.Y(_12370_),
    .A(net508),
    .B(_12355_));
 sg13g2_o21ai_1 _19304_ (.B1(_12370_),
    .Y(_00377_),
    .A1(net58),
    .A2(_12369_));
 sg13g2_buf_1 _19305_ (.A(net1103),
    .X(_12371_));
 sg13g2_nor2b_1 _19306_ (.A(_12367_),
    .B_N(\cpu.dcache.r_data[2][13] ),
    .Y(_12372_));
 sg13g2_a21oi_1 _19307_ (.A1(net1014),
    .A2(_12367_),
    .Y(_12373_),
    .B1(_12372_));
 sg13g2_nand2_1 _19308_ (.Y(_12374_),
    .A(net507),
    .B(_12355_));
 sg13g2_o21ai_1 _19309_ (.B1(_12374_),
    .Y(_00378_),
    .A1(net58),
    .A2(_12373_));
 sg13g2_nor2b_1 _19310_ (.A(_12367_),
    .B_N(\cpu.dcache.r_data[2][14] ),
    .Y(_12375_));
 sg13g2_a21oi_1 _19311_ (.A1(net1015),
    .A2(_12367_),
    .Y(_12376_),
    .B1(_12375_));
 sg13g2_nand2_1 _19312_ (.Y(_12377_),
    .A(net506),
    .B(_12355_));
 sg13g2_o21ai_1 _19313_ (.B1(_12377_),
    .Y(_00379_),
    .A1(_12356_),
    .A2(_12376_));
 sg13g2_nor2b_1 _19314_ (.A(_12367_),
    .B_N(\cpu.dcache.r_data[2][15] ),
    .Y(_12378_));
 sg13g2_a21oi_1 _19315_ (.A1(net1017),
    .A2(_12367_),
    .Y(_12379_),
    .B1(_12378_));
 sg13g2_nand2_1 _19316_ (.Y(_12380_),
    .A(net505),
    .B(_12355_));
 sg13g2_o21ai_1 _19317_ (.B1(_12380_),
    .Y(_00380_),
    .A1(net58),
    .A2(_12379_));
 sg13g2_nor2_1 _19318_ (.A(_12126_),
    .B(_12343_),
    .Y(_12381_));
 sg13g2_buf_2 _19319_ (.A(_12381_),
    .X(_12382_));
 sg13g2_buf_1 _19320_ (.A(_12382_),
    .X(_12383_));
 sg13g2_nor2_1 _19321_ (.A(net669),
    .B(_12120_),
    .Y(_12384_));
 sg13g2_buf_2 _19322_ (.A(_12384_),
    .X(_12385_));
 sg13g2_nor2b_1 _19323_ (.A(_12385_),
    .B_N(\cpu.dcache.r_data[2][16] ),
    .Y(_12386_));
 sg13g2_a21oi_1 _19324_ (.A1(net1016),
    .A2(_12385_),
    .Y(_12387_),
    .B1(_12386_));
 sg13g2_nand2_1 _19325_ (.Y(_12388_),
    .A(net880),
    .B(net57));
 sg13g2_o21ai_1 _19326_ (.B1(_12388_),
    .Y(_00381_),
    .A1(_12383_),
    .A2(_12387_));
 sg13g2_nor2b_1 _19327_ (.A(_12385_),
    .B_N(\cpu.dcache.r_data[2][17] ),
    .Y(_12389_));
 sg13g2_a21oi_1 _19328_ (.A1(net1014),
    .A2(_12385_),
    .Y(_12390_),
    .B1(_12389_));
 sg13g2_nand2_1 _19329_ (.Y(_12391_),
    .A(_12130_),
    .B(net57));
 sg13g2_o21ai_1 _19330_ (.B1(_12391_),
    .Y(_00382_),
    .A1(net57),
    .A2(_12390_));
 sg13g2_nor2b_1 _19331_ (.A(_12385_),
    .B_N(\cpu.dcache.r_data[2][18] ),
    .Y(_12392_));
 sg13g2_a21oi_1 _19332_ (.A1(net1015),
    .A2(_12385_),
    .Y(_12393_),
    .B1(_12392_));
 sg13g2_nand2_1 _19333_ (.Y(_12394_),
    .A(_12132_),
    .B(_12382_));
 sg13g2_o21ai_1 _19334_ (.B1(_12394_),
    .Y(_00383_),
    .A1(_12383_),
    .A2(_12393_));
 sg13g2_nor2b_1 _19335_ (.A(_12385_),
    .B_N(\cpu.dcache.r_data[2][19] ),
    .Y(_12395_));
 sg13g2_a21oi_1 _19336_ (.A1(net1017),
    .A2(_12385_),
    .Y(_12396_),
    .B1(_12395_));
 sg13g2_nand2_1 _19337_ (.Y(_12397_),
    .A(net1024),
    .B(_12382_));
 sg13g2_o21ai_1 _19338_ (.B1(_12397_),
    .Y(_00384_),
    .A1(net57),
    .A2(_12396_));
 sg13g2_nor2b_1 _19339_ (.A(_12350_),
    .B_N(\cpu.dcache.r_data[2][1] ),
    .Y(_12398_));
 sg13g2_a21oi_1 _19340_ (.A1(net1014),
    .A2(_12350_),
    .Y(_12399_),
    .B1(_12398_));
 sg13g2_buf_1 _19341_ (.A(net1061),
    .X(_12400_));
 sg13g2_nand2_1 _19342_ (.Y(_12401_),
    .A(net879),
    .B(net59));
 sg13g2_o21ai_1 _19343_ (.B1(_12401_),
    .Y(_00385_),
    .A1(_12346_),
    .A2(_12399_));
 sg13g2_nor2_1 _19344_ (.A(net669),
    .B(_12268_),
    .Y(_12402_));
 sg13g2_buf_2 _19345_ (.A(_12402_),
    .X(_12403_));
 sg13g2_mux2_1 _19346_ (.A0(\cpu.dcache.r_data[2][20] ),
    .A1(net1102),
    .S(_12403_),
    .X(_12404_));
 sg13g2_nor2_1 _19347_ (.A(_12382_),
    .B(_12404_),
    .Y(_12405_));
 sg13g2_a21oi_1 _19348_ (.A1(_12138_),
    .A2(net57),
    .Y(_00386_),
    .B1(_12405_));
 sg13g2_mux2_1 _19349_ (.A0(\cpu.dcache.r_data[2][21] ),
    .A1(net1101),
    .S(_12403_),
    .X(_12406_));
 sg13g2_nor2_1 _19350_ (.A(_12382_),
    .B(_12406_),
    .Y(_12407_));
 sg13g2_a21oi_1 _19351_ (.A1(net756),
    .A2(net57),
    .Y(_00387_),
    .B1(_12407_));
 sg13g2_mux2_1 _19352_ (.A0(\cpu.dcache.r_data[2][22] ),
    .A1(_12276_),
    .S(_12403_),
    .X(_12408_));
 sg13g2_nor2_1 _19353_ (.A(_12382_),
    .B(_12408_),
    .Y(_12409_));
 sg13g2_a21oi_1 _19354_ (.A1(net755),
    .A2(net57),
    .Y(_00388_),
    .B1(_12409_));
 sg13g2_nor2b_1 _19355_ (.A(_12403_),
    .B_N(\cpu.dcache.r_data[2][23] ),
    .Y(_12410_));
 sg13g2_a21oi_1 _19356_ (.A1(net1017),
    .A2(_12403_),
    .Y(_12411_),
    .B1(_12410_));
 sg13g2_nand2_1 _19357_ (.Y(_12412_),
    .A(net1018),
    .B(_12382_));
 sg13g2_o21ai_1 _19358_ (.B1(_12412_),
    .Y(_00389_),
    .A1(net57),
    .A2(_12411_));
 sg13g2_nor2_1 _19359_ (.A(_12166_),
    .B(_12343_),
    .Y(_12413_));
 sg13g2_buf_2 _19360_ (.A(_12413_),
    .X(_12414_));
 sg13g2_buf_1 _19361_ (.A(_12414_),
    .X(_12415_));
 sg13g2_nor2_1 _19362_ (.A(_12348_),
    .B(_12051_),
    .Y(_12416_));
 sg13g2_buf_1 _19363_ (.A(_12416_),
    .X(_12417_));
 sg13g2_buf_1 _19364_ (.A(_12417_),
    .X(_12418_));
 sg13g2_nor2b_1 _19365_ (.A(net501),
    .B_N(\cpu.dcache.r_data[2][24] ),
    .Y(_12419_));
 sg13g2_a21oi_1 _19366_ (.A1(net1016),
    .A2(net501),
    .Y(_12420_),
    .B1(_12419_));
 sg13g2_nand2_1 _19367_ (.Y(_12421_),
    .A(net504),
    .B(net56));
 sg13g2_o21ai_1 _19368_ (.B1(_12421_),
    .Y(_00390_),
    .A1(net56),
    .A2(_12420_));
 sg13g2_nor2b_1 _19369_ (.A(net501),
    .B_N(\cpu.dcache.r_data[2][25] ),
    .Y(_12422_));
 sg13g2_a21oi_1 _19370_ (.A1(net1014),
    .A2(net501),
    .Y(_12423_),
    .B1(_12422_));
 sg13g2_nand2_1 _19371_ (.Y(_12424_),
    .A(net458),
    .B(_12415_));
 sg13g2_o21ai_1 _19372_ (.B1(_12424_),
    .Y(_00391_),
    .A1(_12415_),
    .A2(_12423_));
 sg13g2_nor2b_1 _19373_ (.A(_12417_),
    .B_N(\cpu.dcache.r_data[2][26] ),
    .Y(_12425_));
 sg13g2_a21oi_1 _19374_ (.A1(net1015),
    .A2(net501),
    .Y(_12426_),
    .B1(_12425_));
 sg13g2_nand2_1 _19375_ (.Y(_12427_),
    .A(_12074_),
    .B(_12414_));
 sg13g2_o21ai_1 _19376_ (.B1(_12427_),
    .Y(_00392_),
    .A1(net56),
    .A2(_12426_));
 sg13g2_nor2b_1 _19377_ (.A(_12417_),
    .B_N(\cpu.dcache.r_data[2][27] ),
    .Y(_12428_));
 sg13g2_a21oi_1 _19378_ (.A1(_12317_),
    .A2(net501),
    .Y(_12429_),
    .B1(_12428_));
 sg13g2_nand2_1 _19379_ (.Y(_12430_),
    .A(net509),
    .B(_12414_));
 sg13g2_o21ai_1 _19380_ (.B1(_12430_),
    .Y(_00393_),
    .A1(net56),
    .A2(_12429_));
 sg13g2_nor2_1 _19381_ (.A(net669),
    .B(_12178_),
    .Y(_12431_));
 sg13g2_buf_2 _19382_ (.A(_12431_),
    .X(_12432_));
 sg13g2_nor2b_1 _19383_ (.A(_12432_),
    .B_N(\cpu.dcache.r_data[2][28] ),
    .Y(_12433_));
 sg13g2_a21oi_1 _19384_ (.A1(_12347_),
    .A2(_12432_),
    .Y(_12434_),
    .B1(_12433_));
 sg13g2_nand2_1 _19385_ (.Y(_12435_),
    .A(net508),
    .B(_12414_));
 sg13g2_o21ai_1 _19386_ (.B1(_12435_),
    .Y(_00394_),
    .A1(net56),
    .A2(_12434_));
 sg13g2_nor2b_1 _19387_ (.A(_12432_),
    .B_N(\cpu.dcache.r_data[2][29] ),
    .Y(_12436_));
 sg13g2_a21oi_1 _19388_ (.A1(_12371_),
    .A2(_12432_),
    .Y(_12437_),
    .B1(_12436_));
 sg13g2_nand2_1 _19389_ (.Y(_12438_),
    .A(_12105_),
    .B(_12414_));
 sg13g2_o21ai_1 _19390_ (.B1(_12438_),
    .Y(_00395_),
    .A1(net56),
    .A2(_12437_));
 sg13g2_nor2b_1 _19391_ (.A(_12350_),
    .B_N(\cpu.dcache.r_data[2][2] ),
    .Y(_12439_));
 sg13g2_a21oi_1 _19392_ (.A1(net1015),
    .A2(_12350_),
    .Y(_12440_),
    .B1(_12439_));
 sg13g2_buf_1 _19393_ (.A(net1060),
    .X(_12441_));
 sg13g2_nand2_1 _19394_ (.Y(_12442_),
    .A(net878),
    .B(_12345_));
 sg13g2_o21ai_1 _19395_ (.B1(_12442_),
    .Y(_00396_),
    .A1(_12346_),
    .A2(_12440_));
 sg13g2_nor2b_1 _19396_ (.A(_12432_),
    .B_N(\cpu.dcache.r_data[2][30] ),
    .Y(_12443_));
 sg13g2_a21oi_1 _19397_ (.A1(_12357_),
    .A2(_12432_),
    .Y(_12444_),
    .B1(_12443_));
 sg13g2_nand2_1 _19398_ (.Y(_12445_),
    .A(net506),
    .B(_12414_));
 sg13g2_o21ai_1 _19399_ (.B1(_12445_),
    .Y(_00397_),
    .A1(net56),
    .A2(_12444_));
 sg13g2_nor2b_1 _19400_ (.A(_12432_),
    .B_N(\cpu.dcache.r_data[2][31] ),
    .Y(_12446_));
 sg13g2_a21oi_1 _19401_ (.A1(_12317_),
    .A2(_12432_),
    .Y(_12447_),
    .B1(_12446_));
 sg13g2_nand2_1 _19402_ (.Y(_12448_),
    .A(net505),
    .B(_12414_));
 sg13g2_o21ai_1 _19403_ (.B1(_12448_),
    .Y(_00398_),
    .A1(net56),
    .A2(_12447_));
 sg13g2_nor2b_1 _19404_ (.A(_12350_),
    .B_N(\cpu.dcache.r_data[2][3] ),
    .Y(_12449_));
 sg13g2_a21oi_1 _19405_ (.A1(net1017),
    .A2(_12350_),
    .Y(_12450_),
    .B1(_12449_));
 sg13g2_nand2_1 _19406_ (.Y(_12451_),
    .A(net1024),
    .B(_12345_));
 sg13g2_o21ai_1 _19407_ (.B1(_12451_),
    .Y(_00399_),
    .A1(net59),
    .A2(_12450_));
 sg13g2_nor2_1 _19408_ (.A(net669),
    .B(_12322_),
    .Y(_12452_));
 sg13g2_buf_2 _19409_ (.A(_12452_),
    .X(_12453_));
 sg13g2_mux2_1 _19410_ (.A0(\cpu.dcache.r_data[2][4] ),
    .A1(net1102),
    .S(_12453_),
    .X(_12454_));
 sg13g2_nor2_1 _19411_ (.A(_12345_),
    .B(_12454_),
    .Y(_12455_));
 sg13g2_a21oi_1 _19412_ (.A1(net757),
    .A2(net59),
    .Y(_00400_),
    .B1(_12455_));
 sg13g2_mux2_1 _19413_ (.A0(\cpu.dcache.r_data[2][5] ),
    .A1(net1101),
    .S(_12453_),
    .X(_12456_));
 sg13g2_nor2_1 _19414_ (.A(_12345_),
    .B(_12456_),
    .Y(_12457_));
 sg13g2_a21oi_1 _19415_ (.A1(net756),
    .A2(net59),
    .Y(_00401_),
    .B1(_12457_));
 sg13g2_mux2_1 _19416_ (.A0(\cpu.dcache.r_data[2][6] ),
    .A1(net1100),
    .S(_12453_),
    .X(_12458_));
 sg13g2_nor2_1 _19417_ (.A(_12345_),
    .B(_12458_),
    .Y(_12459_));
 sg13g2_a21oi_1 _19418_ (.A1(net755),
    .A2(net59),
    .Y(_00402_),
    .B1(_12459_));
 sg13g2_nor2b_1 _19419_ (.A(_12453_),
    .B_N(\cpu.dcache.r_data[2][7] ),
    .Y(_12460_));
 sg13g2_a21oi_1 _19420_ (.A1(net1017),
    .A2(_12453_),
    .Y(_12461_),
    .B1(_12460_));
 sg13g2_nand2_1 _19421_ (.Y(_12462_),
    .A(net1018),
    .B(_12345_));
 sg13g2_o21ai_1 _19422_ (.B1(_12462_),
    .Y(_00403_),
    .A1(net59),
    .A2(_12461_));
 sg13g2_nor2b_1 _19423_ (.A(_12359_),
    .B_N(\cpu.dcache.r_data[2][8] ),
    .Y(_12463_));
 sg13g2_a21oi_1 _19424_ (.A1(net1016),
    .A2(_12359_),
    .Y(_12464_),
    .B1(_12463_));
 sg13g2_nand2_1 _19425_ (.Y(_12465_),
    .A(_12162_),
    .B(_12355_));
 sg13g2_o21ai_1 _19426_ (.B1(_12465_),
    .Y(_00404_),
    .A1(_12356_),
    .A2(_12464_));
 sg13g2_nor2b_1 _19427_ (.A(_12359_),
    .B_N(\cpu.dcache.r_data[2][9] ),
    .Y(_12466_));
 sg13g2_a21oi_1 _19428_ (.A1(net1014),
    .A2(_12359_),
    .Y(_12467_),
    .B1(_12466_));
 sg13g2_nand2_1 _19429_ (.Y(_12468_),
    .A(_12174_),
    .B(_12355_));
 sg13g2_o21ai_1 _19430_ (.B1(_12468_),
    .Y(_00405_),
    .A1(net58),
    .A2(_12467_));
 sg13g2_buf_1 _19431_ (.A(_09425_),
    .X(_12469_));
 sg13g2_buf_1 _19432_ (.A(net609),
    .X(_12470_));
 sg13g2_nand2_1 _19433_ (.Y(_12471_),
    .A(_12470_),
    .B(_12055_));
 sg13g2_nor2_1 _19434_ (.A(_12043_),
    .B(_12471_),
    .Y(_12472_));
 sg13g2_buf_1 _19435_ (.A(_12472_),
    .X(_12473_));
 sg13g2_buf_1 _19436_ (.A(_12473_),
    .X(_12474_));
 sg13g2_buf_1 _19437_ (.A(_09234_),
    .X(_12475_));
 sg13g2_nand2_1 _19438_ (.Y(_12476_),
    .A(net558),
    .B(net790));
 sg13g2_buf_2 _19439_ (.A(_12476_),
    .X(_12477_));
 sg13g2_nor2_1 _19440_ (.A(_12477_),
    .B(_12034_),
    .Y(_12478_));
 sg13g2_buf_2 _19441_ (.A(_12478_),
    .X(_12479_));
 sg13g2_nor2b_1 _19442_ (.A(_12479_),
    .B_N(\cpu.dcache.r_data[3][0] ),
    .Y(_12480_));
 sg13g2_a21oi_1 _19443_ (.A1(net1016),
    .A2(_12479_),
    .Y(_12481_),
    .B1(_12480_));
 sg13g2_nand2_1 _19444_ (.Y(_12482_),
    .A(_12212_),
    .B(net55));
 sg13g2_o21ai_1 _19445_ (.B1(_12482_),
    .Y(_00406_),
    .A1(net55),
    .A2(_12481_));
 sg13g2_nor2_1 _19446_ (.A(_12077_),
    .B(_12471_),
    .Y(_12483_));
 sg13g2_buf_2 _19447_ (.A(_12483_),
    .X(_12484_));
 sg13g2_buf_1 _19448_ (.A(_12484_),
    .X(_12485_));
 sg13g2_nor2_1 _19449_ (.A(_12477_),
    .B(_12062_),
    .Y(_12486_));
 sg13g2_buf_2 _19450_ (.A(_12486_),
    .X(_12487_));
 sg13g2_nor2b_1 _19451_ (.A(_12487_),
    .B_N(\cpu.dcache.r_data[3][10] ),
    .Y(_12488_));
 sg13g2_a21oi_1 _19452_ (.A1(net1015),
    .A2(_12487_),
    .Y(_12489_),
    .B1(_12488_));
 sg13g2_nand2_1 _19453_ (.Y(_12490_),
    .A(net459),
    .B(net54));
 sg13g2_o21ai_1 _19454_ (.B1(_12490_),
    .Y(_00407_),
    .A1(net54),
    .A2(_12489_));
 sg13g2_buf_1 _19455_ (.A(net1104),
    .X(_12491_));
 sg13g2_nor2b_1 _19456_ (.A(_12487_),
    .B_N(\cpu.dcache.r_data[3][11] ),
    .Y(_12492_));
 sg13g2_a21oi_1 _19457_ (.A1(net1013),
    .A2(_12487_),
    .Y(_12493_),
    .B1(_12492_));
 sg13g2_nand2_1 _19458_ (.Y(_12494_),
    .A(net509),
    .B(_12485_));
 sg13g2_o21ai_1 _19459_ (.B1(_12494_),
    .Y(_00408_),
    .A1(_12485_),
    .A2(_12493_));
 sg13g2_nor2_1 _19460_ (.A(_12477_),
    .B(_12089_),
    .Y(_12495_));
 sg13g2_buf_2 _19461_ (.A(_12495_),
    .X(_12496_));
 sg13g2_nor2b_1 _19462_ (.A(_12496_),
    .B_N(\cpu.dcache.r_data[3][12] ),
    .Y(_12497_));
 sg13g2_a21oi_1 _19463_ (.A1(net1016),
    .A2(_12496_),
    .Y(_12498_),
    .B1(_12497_));
 sg13g2_nand2_1 _19464_ (.Y(_12499_),
    .A(net508),
    .B(_12484_));
 sg13g2_o21ai_1 _19465_ (.B1(_12499_),
    .Y(_00409_),
    .A1(net54),
    .A2(_12498_));
 sg13g2_nor2b_1 _19466_ (.A(_12496_),
    .B_N(\cpu.dcache.r_data[3][13] ),
    .Y(_12500_));
 sg13g2_a21oi_1 _19467_ (.A1(net1014),
    .A2(_12496_),
    .Y(_12501_),
    .B1(_12500_));
 sg13g2_nand2_1 _19468_ (.Y(_12502_),
    .A(net507),
    .B(_12484_));
 sg13g2_o21ai_1 _19469_ (.B1(_12502_),
    .Y(_00410_),
    .A1(net54),
    .A2(_12501_));
 sg13g2_nor2b_1 _19470_ (.A(_12496_),
    .B_N(\cpu.dcache.r_data[3][14] ),
    .Y(_12503_));
 sg13g2_a21oi_1 _19471_ (.A1(net1015),
    .A2(_12496_),
    .Y(_12504_),
    .B1(_12503_));
 sg13g2_nand2_1 _19472_ (.Y(_12505_),
    .A(net506),
    .B(_12484_));
 sg13g2_o21ai_1 _19473_ (.B1(_12505_),
    .Y(_00411_),
    .A1(net54),
    .A2(_12504_));
 sg13g2_nor2b_1 _19474_ (.A(_12496_),
    .B_N(\cpu.dcache.r_data[3][15] ),
    .Y(_12506_));
 sg13g2_a21oi_1 _19475_ (.A1(net1013),
    .A2(_12496_),
    .Y(_12507_),
    .B1(_12506_));
 sg13g2_nand2_1 _19476_ (.Y(_12508_),
    .A(net505),
    .B(_12484_));
 sg13g2_o21ai_1 _19477_ (.B1(_12508_),
    .Y(_00412_),
    .A1(net54),
    .A2(_12507_));
 sg13g2_nor2_1 _19478_ (.A(_12126_),
    .B(_12471_),
    .Y(_12509_));
 sg13g2_buf_1 _19479_ (.A(_12509_),
    .X(_12510_));
 sg13g2_buf_1 _19480_ (.A(_12510_),
    .X(_12511_));
 sg13g2_nor2_1 _19481_ (.A(_12477_),
    .B(_12120_),
    .Y(_12512_));
 sg13g2_buf_2 _19482_ (.A(_12512_),
    .X(_12513_));
 sg13g2_nor2b_1 _19483_ (.A(_12513_),
    .B_N(\cpu.dcache.r_data[3][16] ),
    .Y(_12514_));
 sg13g2_a21oi_1 _19484_ (.A1(net1016),
    .A2(_12513_),
    .Y(_12515_),
    .B1(_12514_));
 sg13g2_nand2_1 _19485_ (.Y(_12516_),
    .A(_12212_),
    .B(net53));
 sg13g2_o21ai_1 _19486_ (.B1(_12516_),
    .Y(_00413_),
    .A1(net53),
    .A2(_12515_));
 sg13g2_nor2b_1 _19487_ (.A(_12513_),
    .B_N(\cpu.dcache.r_data[3][17] ),
    .Y(_12517_));
 sg13g2_a21oi_1 _19488_ (.A1(net1014),
    .A2(_12513_),
    .Y(_12518_),
    .B1(_12517_));
 sg13g2_nand2_1 _19489_ (.Y(_12519_),
    .A(_12400_),
    .B(net53));
 sg13g2_o21ai_1 _19490_ (.B1(_12519_),
    .Y(_00414_),
    .A1(net53),
    .A2(_12518_));
 sg13g2_nor2b_1 _19491_ (.A(_12513_),
    .B_N(\cpu.dcache.r_data[3][18] ),
    .Y(_12520_));
 sg13g2_a21oi_1 _19492_ (.A1(net1015),
    .A2(_12513_),
    .Y(_12521_),
    .B1(_12520_));
 sg13g2_nand2_1 _19493_ (.Y(_12522_),
    .A(_12441_),
    .B(_12510_));
 sg13g2_o21ai_1 _19494_ (.B1(_12522_),
    .Y(_00415_),
    .A1(net53),
    .A2(_12521_));
 sg13g2_nor2b_1 _19495_ (.A(_12513_),
    .B_N(\cpu.dcache.r_data[3][19] ),
    .Y(_12523_));
 sg13g2_a21oi_1 _19496_ (.A1(net1013),
    .A2(_12513_),
    .Y(_12524_),
    .B1(_12523_));
 sg13g2_nand2_1 _19497_ (.Y(_12525_),
    .A(_12134_),
    .B(_12510_));
 sg13g2_o21ai_1 _19498_ (.B1(_12525_),
    .Y(_00416_),
    .A1(net53),
    .A2(_12524_));
 sg13g2_nor2b_1 _19499_ (.A(_12479_),
    .B_N(\cpu.dcache.r_data[3][1] ),
    .Y(_12526_));
 sg13g2_a21oi_1 _19500_ (.A1(net1014),
    .A2(_12479_),
    .Y(_12527_),
    .B1(_12526_));
 sg13g2_nand2_1 _19501_ (.Y(_12528_),
    .A(_12400_),
    .B(net55));
 sg13g2_o21ai_1 _19502_ (.B1(_12528_),
    .Y(_00417_),
    .A1(_12474_),
    .A2(_12527_));
 sg13g2_nand2_2 _19503_ (.Y(_12529_),
    .A(net559),
    .B(_12140_));
 sg13g2_mux2_1 _19504_ (.A0(net1102),
    .A1(\cpu.dcache.r_data[3][20] ),
    .S(_12529_),
    .X(_12530_));
 sg13g2_nor2_1 _19505_ (.A(_12510_),
    .B(_12530_),
    .Y(_12531_));
 sg13g2_a21oi_1 _19506_ (.A1(net757),
    .A2(_12511_),
    .Y(_00418_),
    .B1(_12531_));
 sg13g2_mux2_1 _19507_ (.A0(_12273_),
    .A1(\cpu.dcache.r_data[3][21] ),
    .S(_12529_),
    .X(_12532_));
 sg13g2_nor2_1 _19508_ (.A(_12510_),
    .B(_12532_),
    .Y(_12533_));
 sg13g2_a21oi_1 _19509_ (.A1(net756),
    .A2(net53),
    .Y(_00419_),
    .B1(_12533_));
 sg13g2_mux2_1 _19510_ (.A0(net1100),
    .A1(\cpu.dcache.r_data[3][22] ),
    .S(_12529_),
    .X(_12534_));
 sg13g2_nor2_1 _19511_ (.A(_12510_),
    .B(_12534_),
    .Y(_12535_));
 sg13g2_a21oi_1 _19512_ (.A1(net755),
    .A2(net53),
    .Y(_00420_),
    .B1(_12535_));
 sg13g2_mux2_1 _19513_ (.A0(net1108),
    .A1(\cpu.dcache.r_data[3][23] ),
    .S(_12529_),
    .X(_12536_));
 sg13g2_mux2_1 _19514_ (.A0(_12536_),
    .A1(net1023),
    .S(_12511_),
    .X(_00421_));
 sg13g2_nor2_1 _19515_ (.A(_12166_),
    .B(_12471_),
    .Y(_12537_));
 sg13g2_buf_2 _19516_ (.A(_12537_),
    .X(_12538_));
 sg13g2_buf_1 _19517_ (.A(_12538_),
    .X(_12539_));
 sg13g2_nor2_1 _19518_ (.A(_12477_),
    .B(_12051_),
    .Y(_12540_));
 sg13g2_buf_1 _19519_ (.A(_12540_),
    .X(_12541_));
 sg13g2_nor2b_1 _19520_ (.A(net358),
    .B_N(\cpu.dcache.r_data[3][24] ),
    .Y(_12542_));
 sg13g2_a21oi_1 _19521_ (.A1(net1016),
    .A2(net358),
    .Y(_12543_),
    .B1(_12542_));
 sg13g2_nand2_1 _19522_ (.Y(_12544_),
    .A(net504),
    .B(_12539_));
 sg13g2_o21ai_1 _19523_ (.B1(_12544_),
    .Y(_00422_),
    .A1(_12539_),
    .A2(_12543_));
 sg13g2_nor2b_1 _19524_ (.A(net358),
    .B_N(\cpu.dcache.r_data[3][25] ),
    .Y(_12545_));
 sg13g2_a21oi_1 _19525_ (.A1(_12371_),
    .A2(net358),
    .Y(_12546_),
    .B1(_12545_));
 sg13g2_nand2_1 _19526_ (.Y(_12547_),
    .A(net458),
    .B(net52));
 sg13g2_o21ai_1 _19527_ (.B1(_12547_),
    .Y(_00423_),
    .A1(net52),
    .A2(_12546_));
 sg13g2_nor2b_1 _19528_ (.A(net358),
    .B_N(\cpu.dcache.r_data[3][26] ),
    .Y(_12548_));
 sg13g2_a21oi_1 _19529_ (.A1(_12357_),
    .A2(net358),
    .Y(_12549_),
    .B1(_12548_));
 sg13g2_nand2_1 _19530_ (.Y(_12550_),
    .A(net459),
    .B(_12538_));
 sg13g2_o21ai_1 _19531_ (.B1(_12550_),
    .Y(_00424_),
    .A1(net52),
    .A2(_12549_));
 sg13g2_nor2b_1 _19532_ (.A(net358),
    .B_N(\cpu.dcache.r_data[3][27] ),
    .Y(_12551_));
 sg13g2_a21oi_1 _19533_ (.A1(net1013),
    .A2(net358),
    .Y(_12552_),
    .B1(_12551_));
 sg13g2_nand2_1 _19534_ (.Y(_12553_),
    .A(net509),
    .B(_12538_));
 sg13g2_o21ai_1 _19535_ (.B1(_12553_),
    .Y(_00425_),
    .A1(net52),
    .A2(_12552_));
 sg13g2_buf_1 _19536_ (.A(net1106),
    .X(_12554_));
 sg13g2_nor2_1 _19537_ (.A(_12477_),
    .B(_12178_),
    .Y(_12555_));
 sg13g2_buf_2 _19538_ (.A(_12555_),
    .X(_12556_));
 sg13g2_nor2b_1 _19539_ (.A(_12556_),
    .B_N(\cpu.dcache.r_data[3][28] ),
    .Y(_12557_));
 sg13g2_a21oi_1 _19540_ (.A1(net1012),
    .A2(_12556_),
    .Y(_12558_),
    .B1(_12557_));
 sg13g2_nand2_1 _19541_ (.Y(_12559_),
    .A(net508),
    .B(_12538_));
 sg13g2_o21ai_1 _19542_ (.B1(_12559_),
    .Y(_00426_),
    .A1(net52),
    .A2(_12558_));
 sg13g2_buf_1 _19543_ (.A(net1103),
    .X(_12560_));
 sg13g2_nor2b_1 _19544_ (.A(_12556_),
    .B_N(\cpu.dcache.r_data[3][29] ),
    .Y(_12561_));
 sg13g2_a21oi_1 _19545_ (.A1(net1011),
    .A2(_12556_),
    .Y(_12562_),
    .B1(_12561_));
 sg13g2_nand2_1 _19546_ (.Y(_12563_),
    .A(net507),
    .B(_12538_));
 sg13g2_o21ai_1 _19547_ (.B1(_12563_),
    .Y(_00427_),
    .A1(net52),
    .A2(_12562_));
 sg13g2_buf_1 _19548_ (.A(_12217_),
    .X(_12564_));
 sg13g2_nor2b_1 _19549_ (.A(_12479_),
    .B_N(\cpu.dcache.r_data[3][2] ),
    .Y(_12565_));
 sg13g2_a21oi_1 _19550_ (.A1(net1010),
    .A2(_12479_),
    .Y(_12566_),
    .B1(_12565_));
 sg13g2_nand2_1 _19551_ (.Y(_12567_),
    .A(_12441_),
    .B(_12473_));
 sg13g2_o21ai_1 _19552_ (.B1(_12567_),
    .Y(_00428_),
    .A1(_12474_),
    .A2(_12566_));
 sg13g2_nor2b_1 _19553_ (.A(_12556_),
    .B_N(\cpu.dcache.r_data[3][30] ),
    .Y(_12568_));
 sg13g2_a21oi_1 _19554_ (.A1(net1010),
    .A2(_12556_),
    .Y(_12569_),
    .B1(_12568_));
 sg13g2_nand2_1 _19555_ (.Y(_12570_),
    .A(net506),
    .B(_12538_));
 sg13g2_o21ai_1 _19556_ (.B1(_12570_),
    .Y(_00429_),
    .A1(net52),
    .A2(_12569_));
 sg13g2_nor2b_1 _19557_ (.A(_12556_),
    .B_N(\cpu.dcache.r_data[3][31] ),
    .Y(_12571_));
 sg13g2_a21oi_1 _19558_ (.A1(net1013),
    .A2(_12556_),
    .Y(_12572_),
    .B1(_12571_));
 sg13g2_nand2_1 _19559_ (.Y(_12573_),
    .A(net505),
    .B(_12538_));
 sg13g2_o21ai_1 _19560_ (.B1(_12573_),
    .Y(_00430_),
    .A1(net52),
    .A2(_12572_));
 sg13g2_nor2b_1 _19561_ (.A(_12479_),
    .B_N(\cpu.dcache.r_data[3][3] ),
    .Y(_12574_));
 sg13g2_a21oi_1 _19562_ (.A1(net1013),
    .A2(_12479_),
    .Y(_12575_),
    .B1(_12574_));
 sg13g2_nand2_1 _19563_ (.Y(_12576_),
    .A(_12134_),
    .B(_12473_));
 sg13g2_o21ai_1 _19564_ (.B1(_12576_),
    .Y(_00431_),
    .A1(net55),
    .A2(_12575_));
 sg13g2_nand2_2 _19565_ (.Y(_12577_),
    .A(net559),
    .B(_12187_));
 sg13g2_mux2_1 _19566_ (.A0(net1102),
    .A1(\cpu.dcache.r_data[3][4] ),
    .S(_12577_),
    .X(_12578_));
 sg13g2_nor2_1 _19567_ (.A(_12473_),
    .B(_12578_),
    .Y(_12579_));
 sg13g2_a21oi_1 _19568_ (.A1(net757),
    .A2(net55),
    .Y(_00432_),
    .B1(_12579_));
 sg13g2_mux2_1 _19569_ (.A0(net1101),
    .A1(\cpu.dcache.r_data[3][5] ),
    .S(_12577_),
    .X(_12580_));
 sg13g2_nor2_1 _19570_ (.A(_12473_),
    .B(_12580_),
    .Y(_12581_));
 sg13g2_a21oi_1 _19571_ (.A1(net756),
    .A2(net55),
    .Y(_00433_),
    .B1(_12581_));
 sg13g2_mux2_1 _19572_ (.A0(net1100),
    .A1(\cpu.dcache.r_data[3][6] ),
    .S(_12577_),
    .X(_12582_));
 sg13g2_nor2_1 _19573_ (.A(_12473_),
    .B(_12582_),
    .Y(_12583_));
 sg13g2_a21oi_1 _19574_ (.A1(net755),
    .A2(net55),
    .Y(_00434_),
    .B1(_12583_));
 sg13g2_mux2_1 _19575_ (.A0(net1104),
    .A1(\cpu.dcache.r_data[3][7] ),
    .S(_12577_),
    .X(_12584_));
 sg13g2_mux2_1 _19576_ (.A0(_12584_),
    .A1(net1023),
    .S(net55),
    .X(_00435_));
 sg13g2_nor2b_1 _19577_ (.A(_12487_),
    .B_N(\cpu.dcache.r_data[3][8] ),
    .Y(_12585_));
 sg13g2_a21oi_1 _19578_ (.A1(net1012),
    .A2(_12487_),
    .Y(_12586_),
    .B1(_12585_));
 sg13g2_nand2_1 _19579_ (.Y(_12587_),
    .A(net504),
    .B(_12484_));
 sg13g2_o21ai_1 _19580_ (.B1(_12587_),
    .Y(_00436_),
    .A1(net54),
    .A2(_12586_));
 sg13g2_nor2b_1 _19581_ (.A(_12487_),
    .B_N(\cpu.dcache.r_data[3][9] ),
    .Y(_12588_));
 sg13g2_a21oi_1 _19582_ (.A1(net1011),
    .A2(_12487_),
    .Y(_12589_),
    .B1(_12588_));
 sg13g2_nand2_1 _19583_ (.Y(_12590_),
    .A(net458),
    .B(_12484_));
 sg13g2_o21ai_1 _19584_ (.B1(_12590_),
    .Y(_00437_),
    .A1(net54),
    .A2(_12589_));
 sg13g2_nand2_1 _19585_ (.Y(_12591_),
    .A(net574),
    .B(_12055_));
 sg13g2_nor2_1 _19586_ (.A(_12043_),
    .B(_12591_),
    .Y(_12592_));
 sg13g2_buf_2 _19587_ (.A(_12592_),
    .X(_12593_));
 sg13g2_buf_1 _19588_ (.A(_12593_),
    .X(_12594_));
 sg13g2_nor2_1 _19589_ (.A(_10092_),
    .B(_12034_),
    .Y(_12595_));
 sg13g2_buf_2 _19590_ (.A(_12595_),
    .X(_12596_));
 sg13g2_nor2b_1 _19591_ (.A(_12596_),
    .B_N(\cpu.dcache.r_data[4][0] ),
    .Y(_12597_));
 sg13g2_a21oi_1 _19592_ (.A1(net1012),
    .A2(_12596_),
    .Y(_12598_),
    .B1(_12597_));
 sg13g2_nand2_1 _19593_ (.Y(_12599_),
    .A(net880),
    .B(net51));
 sg13g2_o21ai_1 _19594_ (.B1(_12599_),
    .Y(_00438_),
    .A1(net51),
    .A2(_12598_));
 sg13g2_nor2_1 _19595_ (.A(_12077_),
    .B(_12591_),
    .Y(_12600_));
 sg13g2_buf_1 _19596_ (.A(_12600_),
    .X(_12601_));
 sg13g2_buf_1 _19597_ (.A(_12601_),
    .X(_12602_));
 sg13g2_nor2_1 _19598_ (.A(net684),
    .B(_12062_),
    .Y(_12603_));
 sg13g2_buf_2 _19599_ (.A(_12603_),
    .X(_12604_));
 sg13g2_nor2b_1 _19600_ (.A(_12604_),
    .B_N(\cpu.dcache.r_data[4][10] ),
    .Y(_12605_));
 sg13g2_a21oi_1 _19601_ (.A1(net1010),
    .A2(_12604_),
    .Y(_12606_),
    .B1(_12605_));
 sg13g2_nand2_1 _19602_ (.Y(_12607_),
    .A(net459),
    .B(net50));
 sg13g2_o21ai_1 _19603_ (.B1(_12607_),
    .Y(_00439_),
    .A1(net50),
    .A2(_12606_));
 sg13g2_nor2b_1 _19604_ (.A(_12604_),
    .B_N(\cpu.dcache.r_data[4][11] ),
    .Y(_12608_));
 sg13g2_a21oi_1 _19605_ (.A1(_12491_),
    .A2(_12604_),
    .Y(_12609_),
    .B1(_12608_));
 sg13g2_nand2_1 _19606_ (.Y(_12610_),
    .A(net509),
    .B(_12602_));
 sg13g2_o21ai_1 _19607_ (.B1(_12610_),
    .Y(_00440_),
    .A1(net50),
    .A2(_12609_));
 sg13g2_nor2_1 _19608_ (.A(net684),
    .B(_12089_),
    .Y(_12611_));
 sg13g2_buf_2 _19609_ (.A(_12611_),
    .X(_12612_));
 sg13g2_nor2b_1 _19610_ (.A(_12612_),
    .B_N(\cpu.dcache.r_data[4][12] ),
    .Y(_12613_));
 sg13g2_a21oi_1 _19611_ (.A1(_12554_),
    .A2(_12612_),
    .Y(_12614_),
    .B1(_12613_));
 sg13g2_nand2_1 _19612_ (.Y(_12615_),
    .A(net508),
    .B(_12601_));
 sg13g2_o21ai_1 _19613_ (.B1(_12615_),
    .Y(_00441_),
    .A1(net50),
    .A2(_12614_));
 sg13g2_nor2b_1 _19614_ (.A(_12612_),
    .B_N(\cpu.dcache.r_data[4][13] ),
    .Y(_12616_));
 sg13g2_a21oi_1 _19615_ (.A1(_12560_),
    .A2(_12612_),
    .Y(_12617_),
    .B1(_12616_));
 sg13g2_nand2_1 _19616_ (.Y(_12618_),
    .A(net507),
    .B(_12601_));
 sg13g2_o21ai_1 _19617_ (.B1(_12618_),
    .Y(_00442_),
    .A1(net50),
    .A2(_12617_));
 sg13g2_nor2b_1 _19618_ (.A(_12612_),
    .B_N(\cpu.dcache.r_data[4][14] ),
    .Y(_12619_));
 sg13g2_a21oi_1 _19619_ (.A1(_12564_),
    .A2(_12612_),
    .Y(_12620_),
    .B1(_12619_));
 sg13g2_nand2_1 _19620_ (.Y(_12621_),
    .A(net506),
    .B(_12601_));
 sg13g2_o21ai_1 _19621_ (.B1(_12621_),
    .Y(_00443_),
    .A1(net50),
    .A2(_12620_));
 sg13g2_nor2b_1 _19622_ (.A(_12612_),
    .B_N(\cpu.dcache.r_data[4][15] ),
    .Y(_12622_));
 sg13g2_a21oi_1 _19623_ (.A1(_12491_),
    .A2(_12612_),
    .Y(_12623_),
    .B1(_12622_));
 sg13g2_nand2_1 _19624_ (.Y(_12624_),
    .A(net505),
    .B(_12601_));
 sg13g2_o21ai_1 _19625_ (.B1(_12624_),
    .Y(_00444_),
    .A1(net50),
    .A2(_12623_));
 sg13g2_nor2_1 _19626_ (.A(_12126_),
    .B(_12591_),
    .Y(_12625_));
 sg13g2_buf_2 _19627_ (.A(_12625_),
    .X(_12626_));
 sg13g2_buf_1 _19628_ (.A(_12626_),
    .X(_12627_));
 sg13g2_nor2_1 _19629_ (.A(net684),
    .B(_12120_),
    .Y(_12628_));
 sg13g2_buf_2 _19630_ (.A(_12628_),
    .X(_12629_));
 sg13g2_nor2b_1 _19631_ (.A(_12629_),
    .B_N(\cpu.dcache.r_data[4][16] ),
    .Y(_12630_));
 sg13g2_a21oi_1 _19632_ (.A1(net1012),
    .A2(_12629_),
    .Y(_12631_),
    .B1(_12630_));
 sg13g2_nand2_1 _19633_ (.Y(_12632_),
    .A(net880),
    .B(net49));
 sg13g2_o21ai_1 _19634_ (.B1(_12632_),
    .Y(_00445_),
    .A1(net49),
    .A2(_12631_));
 sg13g2_nor2b_1 _19635_ (.A(_12629_),
    .B_N(\cpu.dcache.r_data[4][17] ),
    .Y(_12633_));
 sg13g2_a21oi_1 _19636_ (.A1(net1011),
    .A2(_12629_),
    .Y(_12634_),
    .B1(_12633_));
 sg13g2_nand2_1 _19637_ (.Y(_12635_),
    .A(net879),
    .B(net49));
 sg13g2_o21ai_1 _19638_ (.B1(_12635_),
    .Y(_00446_),
    .A1(net49),
    .A2(_12634_));
 sg13g2_nor2b_1 _19639_ (.A(_12629_),
    .B_N(\cpu.dcache.r_data[4][18] ),
    .Y(_12636_));
 sg13g2_a21oi_1 _19640_ (.A1(net1010),
    .A2(_12629_),
    .Y(_12637_),
    .B1(_12636_));
 sg13g2_nand2_1 _19641_ (.Y(_12638_),
    .A(net878),
    .B(_12626_));
 sg13g2_o21ai_1 _19642_ (.B1(_12638_),
    .Y(_00447_),
    .A1(net49),
    .A2(_12637_));
 sg13g2_nor2b_1 _19643_ (.A(_12629_),
    .B_N(\cpu.dcache.r_data[4][19] ),
    .Y(_12639_));
 sg13g2_a21oi_1 _19644_ (.A1(net1013),
    .A2(_12629_),
    .Y(_12640_),
    .B1(_12639_));
 sg13g2_nand2_1 _19645_ (.Y(_12641_),
    .A(net1054),
    .B(_12626_));
 sg13g2_o21ai_1 _19646_ (.B1(_12641_),
    .Y(_00448_),
    .A1(net49),
    .A2(_12640_));
 sg13g2_nor2b_1 _19647_ (.A(_12596_),
    .B_N(\cpu.dcache.r_data[4][1] ),
    .Y(_12642_));
 sg13g2_a21oi_1 _19648_ (.A1(net1011),
    .A2(_12596_),
    .Y(_12643_),
    .B1(_12642_));
 sg13g2_nand2_1 _19649_ (.Y(_12644_),
    .A(net879),
    .B(net51));
 sg13g2_o21ai_1 _19650_ (.B1(_12644_),
    .Y(_00449_),
    .A1(net51),
    .A2(_12643_));
 sg13g2_nor2_1 _19651_ (.A(net684),
    .B(_12268_),
    .Y(_12645_));
 sg13g2_buf_2 _19652_ (.A(_12645_),
    .X(_12646_));
 sg13g2_mux2_1 _19653_ (.A0(\cpu.dcache.r_data[4][20] ),
    .A1(net1102),
    .S(_12646_),
    .X(_12647_));
 sg13g2_nor2_1 _19654_ (.A(_12626_),
    .B(_12647_),
    .Y(_12648_));
 sg13g2_a21oi_1 _19655_ (.A1(net757),
    .A2(net49),
    .Y(_00450_),
    .B1(_12648_));
 sg13g2_mux2_1 _19656_ (.A0(\cpu.dcache.r_data[4][21] ),
    .A1(net1101),
    .S(_12646_),
    .X(_12649_));
 sg13g2_nor2_1 _19657_ (.A(_12626_),
    .B(_12649_),
    .Y(_12650_));
 sg13g2_a21oi_1 _19658_ (.A1(net756),
    .A2(net49),
    .Y(_00451_),
    .B1(_12650_));
 sg13g2_mux2_1 _19659_ (.A0(\cpu.dcache.r_data[4][22] ),
    .A1(net1100),
    .S(_12646_),
    .X(_12651_));
 sg13g2_nor2_1 _19660_ (.A(_12626_),
    .B(_12651_),
    .Y(_12652_));
 sg13g2_a21oi_1 _19661_ (.A1(_12151_),
    .A2(_12627_),
    .Y(_00452_),
    .B1(_12652_));
 sg13g2_nor2b_1 _19662_ (.A(_12646_),
    .B_N(\cpu.dcache.r_data[4][23] ),
    .Y(_12653_));
 sg13g2_a21oi_1 _19663_ (.A1(net1013),
    .A2(_12646_),
    .Y(_12654_),
    .B1(_12653_));
 sg13g2_nand2_1 _19664_ (.Y(_12655_),
    .A(_12281_),
    .B(_12626_));
 sg13g2_o21ai_1 _19665_ (.B1(_12655_),
    .Y(_00453_),
    .A1(_12627_),
    .A2(_12654_));
 sg13g2_nand2_1 _19666_ (.Y(_12656_),
    .A(net574),
    .B(_12156_));
 sg13g2_buf_1 _19667_ (.A(_12656_),
    .X(_12657_));
 sg13g2_mux2_1 _19668_ (.A0(_12021_),
    .A1(\cpu.dcache.r_data[4][24] ),
    .S(net457),
    .X(_12658_));
 sg13g2_nor2_1 _19669_ (.A(_12166_),
    .B(_12591_),
    .Y(_12659_));
 sg13g2_buf_1 _19670_ (.A(_12659_),
    .X(_12660_));
 sg13g2_mux2_1 _19671_ (.A0(_12658_),
    .A1(net504),
    .S(net77),
    .X(_00454_));
 sg13g2_mux2_1 _19672_ (.A0(net1107),
    .A1(\cpu.dcache.r_data[4][25] ),
    .S(net457),
    .X(_12661_));
 sg13g2_mux2_1 _19673_ (.A0(_12661_),
    .A1(net458),
    .S(net77),
    .X(_00455_));
 sg13g2_mux2_1 _19674_ (.A0(_12060_),
    .A1(\cpu.dcache.r_data[4][26] ),
    .S(net457),
    .X(_12662_));
 sg13g2_mux2_1 _19675_ (.A0(_12662_),
    .A1(net459),
    .S(_12660_),
    .X(_00456_));
 sg13g2_mux2_1 _19676_ (.A0(net1104),
    .A1(\cpu.dcache.r_data[4][27] ),
    .S(_12656_),
    .X(_12663_));
 sg13g2_mux2_1 _19677_ (.A0(_12663_),
    .A1(net509),
    .S(_12660_),
    .X(_00457_));
 sg13g2_nor2_1 _19678_ (.A(_10092_),
    .B(_12178_),
    .Y(_12664_));
 sg13g2_buf_2 _19679_ (.A(_12664_),
    .X(_12665_));
 sg13g2_nor2b_1 _19680_ (.A(_12665_),
    .B_N(\cpu.dcache.r_data[4][28] ),
    .Y(_12666_));
 sg13g2_a21oi_1 _19681_ (.A1(net1012),
    .A2(_12665_),
    .Y(_12667_),
    .B1(_12666_));
 sg13g2_nand2_1 _19682_ (.Y(_12668_),
    .A(net508),
    .B(net77));
 sg13g2_o21ai_1 _19683_ (.B1(_12668_),
    .Y(_00458_),
    .A1(net77),
    .A2(_12667_));
 sg13g2_nor2b_1 _19684_ (.A(_12665_),
    .B_N(\cpu.dcache.r_data[4][29] ),
    .Y(_12669_));
 sg13g2_a21oi_1 _19685_ (.A1(net1011),
    .A2(_12665_),
    .Y(_12670_),
    .B1(_12669_));
 sg13g2_nand2_1 _19686_ (.Y(_12671_),
    .A(net507),
    .B(net77));
 sg13g2_o21ai_1 _19687_ (.B1(_12671_),
    .Y(_00459_),
    .A1(net77),
    .A2(_12670_));
 sg13g2_nor2b_1 _19688_ (.A(_12596_),
    .B_N(\cpu.dcache.r_data[4][2] ),
    .Y(_12672_));
 sg13g2_a21oi_1 _19689_ (.A1(net1010),
    .A2(_12596_),
    .Y(_12673_),
    .B1(_12672_));
 sg13g2_nand2_1 _19690_ (.Y(_12674_),
    .A(net878),
    .B(_12593_));
 sg13g2_o21ai_1 _19691_ (.B1(_12674_),
    .Y(_00460_),
    .A1(_12594_),
    .A2(_12673_));
 sg13g2_nor2b_1 _19692_ (.A(_12665_),
    .B_N(\cpu.dcache.r_data[4][30] ),
    .Y(_12675_));
 sg13g2_a21oi_1 _19693_ (.A1(net1010),
    .A2(_12665_),
    .Y(_12676_),
    .B1(_12675_));
 sg13g2_nand2_1 _19694_ (.Y(_12677_),
    .A(net506),
    .B(_12659_));
 sg13g2_o21ai_1 _19695_ (.B1(_12677_),
    .Y(_00461_),
    .A1(net77),
    .A2(_12676_));
 sg13g2_buf_1 _19696_ (.A(net1104),
    .X(_12678_));
 sg13g2_nor2b_1 _19697_ (.A(_12665_),
    .B_N(\cpu.dcache.r_data[4][31] ),
    .Y(_12679_));
 sg13g2_a21oi_1 _19698_ (.A1(net1009),
    .A2(_12665_),
    .Y(_12680_),
    .B1(_12679_));
 sg13g2_nand2_1 _19699_ (.Y(_12681_),
    .A(net505),
    .B(_12659_));
 sg13g2_o21ai_1 _19700_ (.B1(_12681_),
    .Y(_00462_),
    .A1(net77),
    .A2(_12680_));
 sg13g2_nor2b_1 _19701_ (.A(_12596_),
    .B_N(\cpu.dcache.r_data[4][3] ),
    .Y(_12682_));
 sg13g2_a21oi_1 _19702_ (.A1(_12678_),
    .A2(_12596_),
    .Y(_12683_),
    .B1(_12682_));
 sg13g2_nand2_1 _19703_ (.Y(_12684_),
    .A(_10121_),
    .B(_12593_));
 sg13g2_o21ai_1 _19704_ (.B1(_12684_),
    .Y(_00463_),
    .A1(_12594_),
    .A2(_12683_));
 sg13g2_nor2_1 _19705_ (.A(net684),
    .B(_12322_),
    .Y(_12685_));
 sg13g2_buf_2 _19706_ (.A(_12685_),
    .X(_12686_));
 sg13g2_mux2_1 _19707_ (.A0(\cpu.dcache.r_data[4][4] ),
    .A1(net1102),
    .S(_12686_),
    .X(_12687_));
 sg13g2_nor2_1 _19708_ (.A(_12593_),
    .B(_12687_),
    .Y(_12688_));
 sg13g2_a21oi_1 _19709_ (.A1(net757),
    .A2(net51),
    .Y(_00464_),
    .B1(_12688_));
 sg13g2_mux2_1 _19710_ (.A0(\cpu.dcache.r_data[4][5] ),
    .A1(net1101),
    .S(_12686_),
    .X(_12689_));
 sg13g2_nor2_1 _19711_ (.A(_12593_),
    .B(_12689_),
    .Y(_12690_));
 sg13g2_a21oi_1 _19712_ (.A1(net756),
    .A2(net51),
    .Y(_00465_),
    .B1(_12690_));
 sg13g2_mux2_1 _19713_ (.A0(\cpu.dcache.r_data[4][6] ),
    .A1(net1100),
    .S(_12686_),
    .X(_12691_));
 sg13g2_nor2_1 _19714_ (.A(_12593_),
    .B(_12691_),
    .Y(_12692_));
 sg13g2_a21oi_1 _19715_ (.A1(net755),
    .A2(net51),
    .Y(_00466_),
    .B1(_12692_));
 sg13g2_nor2b_1 _19716_ (.A(_12686_),
    .B_N(\cpu.dcache.r_data[4][7] ),
    .Y(_12693_));
 sg13g2_a21oi_1 _19717_ (.A1(net1009),
    .A2(_12686_),
    .Y(_12694_),
    .B1(_12693_));
 sg13g2_nand2_1 _19718_ (.Y(_12695_),
    .A(_12281_),
    .B(_12593_));
 sg13g2_o21ai_1 _19719_ (.B1(_12695_),
    .Y(_00467_),
    .A1(net51),
    .A2(_12694_));
 sg13g2_nor2b_1 _19720_ (.A(_12604_),
    .B_N(\cpu.dcache.r_data[4][8] ),
    .Y(_12696_));
 sg13g2_a21oi_1 _19721_ (.A1(net1012),
    .A2(_12604_),
    .Y(_12697_),
    .B1(_12696_));
 sg13g2_nand2_1 _19722_ (.Y(_12698_),
    .A(net504),
    .B(_12601_));
 sg13g2_o21ai_1 _19723_ (.B1(_12698_),
    .Y(_00468_),
    .A1(net50),
    .A2(_12697_));
 sg13g2_nor2b_1 _19724_ (.A(_12604_),
    .B_N(\cpu.dcache.r_data[4][9] ),
    .Y(_12699_));
 sg13g2_a21oi_1 _19725_ (.A1(net1011),
    .A2(_12604_),
    .Y(_12700_),
    .B1(_12699_));
 sg13g2_nand2_1 _19726_ (.Y(_12701_),
    .A(net458),
    .B(_12601_));
 sg13g2_o21ai_1 _19727_ (.B1(_12701_),
    .Y(_00469_),
    .A1(_12602_),
    .A2(_12700_));
 sg13g2_buf_1 _19728_ (.A(_09460_),
    .X(_12702_));
 sg13g2_buf_1 _19729_ (.A(net608),
    .X(_12703_));
 sg13g2_nand2_1 _19730_ (.Y(_12704_),
    .A(net557),
    .B(_12055_));
 sg13g2_nor2_1 _19731_ (.A(_12043_),
    .B(_12704_),
    .Y(_12705_));
 sg13g2_buf_2 _19732_ (.A(_12705_),
    .X(_12706_));
 sg13g2_buf_1 _19733_ (.A(_12706_),
    .X(_12707_));
 sg13g2_nand2_1 _19734_ (.Y(_12708_),
    .A(net926),
    .B(net689));
 sg13g2_buf_2 _19735_ (.A(_12708_),
    .X(_12709_));
 sg13g2_buf_1 _19736_ (.A(_12709_),
    .X(_12710_));
 sg13g2_nor2_1 _19737_ (.A(net500),
    .B(_12034_),
    .Y(_12711_));
 sg13g2_buf_2 _19738_ (.A(_12711_),
    .X(_12712_));
 sg13g2_nor2b_1 _19739_ (.A(_12712_),
    .B_N(\cpu.dcache.r_data[5][0] ),
    .Y(_12713_));
 sg13g2_a21oi_1 _19740_ (.A1(net1012),
    .A2(_12712_),
    .Y(_12714_),
    .B1(_12713_));
 sg13g2_nand2_1 _19741_ (.Y(_12715_),
    .A(net880),
    .B(net48));
 sg13g2_o21ai_1 _19742_ (.B1(_12715_),
    .Y(_00470_),
    .A1(net48),
    .A2(_12714_));
 sg13g2_nor2_1 _19743_ (.A(_12077_),
    .B(_12704_),
    .Y(_12716_));
 sg13g2_buf_2 _19744_ (.A(_12716_),
    .X(_12717_));
 sg13g2_buf_1 _19745_ (.A(_12717_),
    .X(_12718_));
 sg13g2_nor2_1 _19746_ (.A(net500),
    .B(_12062_),
    .Y(_12719_));
 sg13g2_buf_2 _19747_ (.A(_12719_),
    .X(_12720_));
 sg13g2_nor2b_1 _19748_ (.A(_12720_),
    .B_N(\cpu.dcache.r_data[5][10] ),
    .Y(_12721_));
 sg13g2_a21oi_1 _19749_ (.A1(net1010),
    .A2(_12720_),
    .Y(_12722_),
    .B1(_12721_));
 sg13g2_nand2_1 _19750_ (.Y(_12723_),
    .A(_12073_),
    .B(net47));
 sg13g2_o21ai_1 _19751_ (.B1(_12723_),
    .Y(_00471_),
    .A1(net47),
    .A2(_12722_));
 sg13g2_nor2b_1 _19752_ (.A(_12720_),
    .B_N(\cpu.dcache.r_data[5][11] ),
    .Y(_12724_));
 sg13g2_a21oi_1 _19753_ (.A1(net1009),
    .A2(_12720_),
    .Y(_12725_),
    .B1(_12724_));
 sg13g2_nand2_1 _19754_ (.Y(_12726_),
    .A(_12084_),
    .B(net47));
 sg13g2_o21ai_1 _19755_ (.B1(_12726_),
    .Y(_00472_),
    .A1(net47),
    .A2(_12725_));
 sg13g2_nor2_1 _19756_ (.A(net500),
    .B(_12089_),
    .Y(_12727_));
 sg13g2_buf_2 _19757_ (.A(_12727_),
    .X(_12728_));
 sg13g2_nor2b_1 _19758_ (.A(_12728_),
    .B_N(\cpu.dcache.r_data[5][12] ),
    .Y(_12729_));
 sg13g2_a21oi_1 _19759_ (.A1(_12554_),
    .A2(_12728_),
    .Y(_12730_),
    .B1(_12729_));
 sg13g2_nand2_1 _19760_ (.Y(_12731_),
    .A(_12096_),
    .B(_12717_));
 sg13g2_o21ai_1 _19761_ (.B1(_12731_),
    .Y(_00473_),
    .A1(net47),
    .A2(_12730_));
 sg13g2_nor2b_1 _19762_ (.A(_12728_),
    .B_N(\cpu.dcache.r_data[5][13] ),
    .Y(_12732_));
 sg13g2_a21oi_1 _19763_ (.A1(_12560_),
    .A2(_12728_),
    .Y(_12733_),
    .B1(_12732_));
 sg13g2_nand2_1 _19764_ (.Y(_12734_),
    .A(_12104_),
    .B(_12717_));
 sg13g2_o21ai_1 _19765_ (.B1(_12734_),
    .Y(_00474_),
    .A1(net47),
    .A2(_12733_));
 sg13g2_nor2b_1 _19766_ (.A(_12728_),
    .B_N(\cpu.dcache.r_data[5][14] ),
    .Y(_12735_));
 sg13g2_a21oi_1 _19767_ (.A1(_12564_),
    .A2(_12728_),
    .Y(_12736_),
    .B1(_12735_));
 sg13g2_nand2_1 _19768_ (.Y(_12737_),
    .A(_12110_),
    .B(_12717_));
 sg13g2_o21ai_1 _19769_ (.B1(_12737_),
    .Y(_00475_),
    .A1(_12718_),
    .A2(_12736_));
 sg13g2_nor2b_1 _19770_ (.A(_12728_),
    .B_N(\cpu.dcache.r_data[5][15] ),
    .Y(_12738_));
 sg13g2_a21oi_1 _19771_ (.A1(net1009),
    .A2(_12728_),
    .Y(_12739_),
    .B1(_12738_));
 sg13g2_nand2_1 _19772_ (.Y(_12740_),
    .A(_12116_),
    .B(_12717_));
 sg13g2_o21ai_1 _19773_ (.B1(_12740_),
    .Y(_00476_),
    .A1(net47),
    .A2(_12739_));
 sg13g2_nor2_1 _19774_ (.A(_12126_),
    .B(_12704_),
    .Y(_12741_));
 sg13g2_buf_2 _19775_ (.A(_12741_),
    .X(_12742_));
 sg13g2_buf_1 _19776_ (.A(_12742_),
    .X(_12743_));
 sg13g2_nor2_1 _19777_ (.A(net500),
    .B(_12120_),
    .Y(_12744_));
 sg13g2_buf_2 _19778_ (.A(_12744_),
    .X(_12745_));
 sg13g2_nor2b_1 _19779_ (.A(_12745_),
    .B_N(\cpu.dcache.r_data[5][16] ),
    .Y(_12746_));
 sg13g2_a21oi_1 _19780_ (.A1(net1012),
    .A2(_12745_),
    .Y(_12747_),
    .B1(_12746_));
 sg13g2_nand2_1 _19781_ (.Y(_12748_),
    .A(net880),
    .B(net46));
 sg13g2_o21ai_1 _19782_ (.B1(_12748_),
    .Y(_00477_),
    .A1(net46),
    .A2(_12747_));
 sg13g2_nor2b_1 _19783_ (.A(_12745_),
    .B_N(\cpu.dcache.r_data[5][17] ),
    .Y(_12749_));
 sg13g2_a21oi_1 _19784_ (.A1(net1011),
    .A2(_12745_),
    .Y(_12750_),
    .B1(_12749_));
 sg13g2_nand2_1 _19785_ (.Y(_12751_),
    .A(net879),
    .B(net46));
 sg13g2_o21ai_1 _19786_ (.B1(_12751_),
    .Y(_00478_),
    .A1(net46),
    .A2(_12750_));
 sg13g2_nor2b_1 _19787_ (.A(_12745_),
    .B_N(\cpu.dcache.r_data[5][18] ),
    .Y(_12752_));
 sg13g2_a21oi_1 _19788_ (.A1(net1010),
    .A2(_12745_),
    .Y(_12753_),
    .B1(_12752_));
 sg13g2_nand2_1 _19789_ (.Y(_12754_),
    .A(net878),
    .B(_12742_));
 sg13g2_o21ai_1 _19790_ (.B1(_12754_),
    .Y(_00479_),
    .A1(net46),
    .A2(_12753_));
 sg13g2_nor2b_1 _19791_ (.A(_12745_),
    .B_N(\cpu.dcache.r_data[5][19] ),
    .Y(_12755_));
 sg13g2_a21oi_1 _19792_ (.A1(net1009),
    .A2(_12745_),
    .Y(_12756_),
    .B1(_12755_));
 sg13g2_nand2_1 _19793_ (.Y(_12757_),
    .A(net1054),
    .B(_12742_));
 sg13g2_o21ai_1 _19794_ (.B1(_12757_),
    .Y(_00480_),
    .A1(net46),
    .A2(_12756_));
 sg13g2_nor2b_1 _19795_ (.A(_12712_),
    .B_N(\cpu.dcache.r_data[5][1] ),
    .Y(_12758_));
 sg13g2_a21oi_1 _19796_ (.A1(net1011),
    .A2(_12712_),
    .Y(_12759_),
    .B1(_12758_));
 sg13g2_nand2_1 _19797_ (.Y(_12760_),
    .A(net879),
    .B(net48));
 sg13g2_o21ai_1 _19798_ (.B1(_12760_),
    .Y(_00481_),
    .A1(net48),
    .A2(_12759_));
 sg13g2_buf_1 _19799_ (.A(_12136_),
    .X(_12761_));
 sg13g2_nor2_1 _19800_ (.A(net500),
    .B(_12268_),
    .Y(_12762_));
 sg13g2_buf_2 _19801_ (.A(_12762_),
    .X(_12763_));
 sg13g2_mux2_1 _19802_ (.A0(\cpu.dcache.r_data[5][20] ),
    .A1(net1106),
    .S(_12763_),
    .X(_12764_));
 sg13g2_nor2_1 _19803_ (.A(_12742_),
    .B(_12764_),
    .Y(_12765_));
 sg13g2_a21oi_1 _19804_ (.A1(net877),
    .A2(net46),
    .Y(_00482_),
    .B1(_12765_));
 sg13g2_buf_1 _19805_ (.A(_12144_),
    .X(_12766_));
 sg13g2_mux2_1 _19806_ (.A0(\cpu.dcache.r_data[5][21] ),
    .A1(net1103),
    .S(_12763_),
    .X(_12767_));
 sg13g2_nor2_1 _19807_ (.A(_12742_),
    .B(_12767_),
    .Y(_12768_));
 sg13g2_a21oi_1 _19808_ (.A1(net876),
    .A2(net46),
    .Y(_00483_),
    .B1(_12768_));
 sg13g2_buf_1 _19809_ (.A(_12149_),
    .X(_12769_));
 sg13g2_mux2_1 _19810_ (.A0(\cpu.dcache.r_data[5][22] ),
    .A1(net1105),
    .S(_12763_),
    .X(_12770_));
 sg13g2_nor2_1 _19811_ (.A(_12742_),
    .B(_12770_),
    .Y(_12771_));
 sg13g2_a21oi_1 _19812_ (.A1(net875),
    .A2(_12743_),
    .Y(_00484_),
    .B1(_12771_));
 sg13g2_nor2b_1 _19813_ (.A(_12763_),
    .B_N(\cpu.dcache.r_data[5][23] ),
    .Y(_12772_));
 sg13g2_a21oi_1 _19814_ (.A1(net1009),
    .A2(_12763_),
    .Y(_12773_),
    .B1(_12772_));
 sg13g2_nand2_1 _19815_ (.Y(_12774_),
    .A(net1053),
    .B(_12742_));
 sg13g2_o21ai_1 _19816_ (.B1(_12774_),
    .Y(_00485_),
    .A1(_12743_),
    .A2(_12773_));
 sg13g2_nor2_1 _19817_ (.A(_12166_),
    .B(_12704_),
    .Y(_12775_));
 sg13g2_buf_2 _19818_ (.A(_12775_),
    .X(_12776_));
 sg13g2_buf_1 _19819_ (.A(_12776_),
    .X(_12777_));
 sg13g2_buf_1 _19820_ (.A(net1106),
    .X(_12778_));
 sg13g2_nor2_1 _19821_ (.A(_12710_),
    .B(_12051_),
    .Y(_12779_));
 sg13g2_buf_1 _19822_ (.A(_12779_),
    .X(_12780_));
 sg13g2_nor2b_1 _19823_ (.A(net416),
    .B_N(\cpu.dcache.r_data[5][24] ),
    .Y(_12781_));
 sg13g2_a21oi_1 _19824_ (.A1(net1008),
    .A2(net416),
    .Y(_12782_),
    .B1(_12781_));
 sg13g2_nand2_1 _19825_ (.Y(_12783_),
    .A(_12161_),
    .B(net45));
 sg13g2_o21ai_1 _19826_ (.B1(_12783_),
    .Y(_00486_),
    .A1(net45),
    .A2(_12782_));
 sg13g2_buf_1 _19827_ (.A(net1103),
    .X(_12784_));
 sg13g2_nor2b_1 _19828_ (.A(net416),
    .B_N(\cpu.dcache.r_data[5][25] ),
    .Y(_12785_));
 sg13g2_a21oi_1 _19829_ (.A1(net1007),
    .A2(net416),
    .Y(_12786_),
    .B1(_12785_));
 sg13g2_nand2_1 _19830_ (.Y(_12787_),
    .A(_12173_),
    .B(_12777_));
 sg13g2_o21ai_1 _19831_ (.B1(_12787_),
    .Y(_00487_),
    .A1(_12777_),
    .A2(_12786_));
 sg13g2_buf_1 _19832_ (.A(net1105),
    .X(_12788_));
 sg13g2_nor2b_1 _19833_ (.A(net416),
    .B_N(\cpu.dcache.r_data[5][26] ),
    .Y(_12789_));
 sg13g2_a21oi_1 _19834_ (.A1(net1006),
    .A2(net416),
    .Y(_12790_),
    .B1(_12789_));
 sg13g2_nand2_1 _19835_ (.Y(_12791_),
    .A(_12073_),
    .B(_12776_));
 sg13g2_o21ai_1 _19836_ (.B1(_12791_),
    .Y(_00488_),
    .A1(net45),
    .A2(_12790_));
 sg13g2_nor2b_1 _19837_ (.A(net416),
    .B_N(\cpu.dcache.r_data[5][27] ),
    .Y(_12792_));
 sg13g2_a21oi_1 _19838_ (.A1(net1009),
    .A2(net416),
    .Y(_12793_),
    .B1(_12792_));
 sg13g2_nand2_1 _19839_ (.Y(_12794_),
    .A(_12084_),
    .B(_12776_));
 sg13g2_o21ai_1 _19840_ (.B1(_12794_),
    .Y(_00489_),
    .A1(net45),
    .A2(_12793_));
 sg13g2_nor2_1 _19841_ (.A(net500),
    .B(_12178_),
    .Y(_12795_));
 sg13g2_buf_2 _19842_ (.A(_12795_),
    .X(_12796_));
 sg13g2_nor2b_1 _19843_ (.A(_12796_),
    .B_N(\cpu.dcache.r_data[5][28] ),
    .Y(_12797_));
 sg13g2_a21oi_1 _19844_ (.A1(net1008),
    .A2(_12796_),
    .Y(_12798_),
    .B1(_12797_));
 sg13g2_nand2_1 _19845_ (.Y(_12799_),
    .A(_12096_),
    .B(_12776_));
 sg13g2_o21ai_1 _19846_ (.B1(_12799_),
    .Y(_00490_),
    .A1(net45),
    .A2(_12798_));
 sg13g2_nor2b_1 _19847_ (.A(_12796_),
    .B_N(\cpu.dcache.r_data[5][29] ),
    .Y(_12800_));
 sg13g2_a21oi_1 _19848_ (.A1(net1007),
    .A2(_12796_),
    .Y(_12801_),
    .B1(_12800_));
 sg13g2_nand2_1 _19849_ (.Y(_12802_),
    .A(_12104_),
    .B(_12776_));
 sg13g2_o21ai_1 _19850_ (.B1(_12802_),
    .Y(_00491_),
    .A1(net45),
    .A2(_12801_));
 sg13g2_nor2b_1 _19851_ (.A(_12712_),
    .B_N(\cpu.dcache.r_data[5][2] ),
    .Y(_12803_));
 sg13g2_a21oi_1 _19852_ (.A1(net1006),
    .A2(_12712_),
    .Y(_12804_),
    .B1(_12803_));
 sg13g2_nand2_1 _19853_ (.Y(_12805_),
    .A(net878),
    .B(_12706_));
 sg13g2_o21ai_1 _19854_ (.B1(_12805_),
    .Y(_00492_),
    .A1(net48),
    .A2(_12804_));
 sg13g2_nor2b_1 _19855_ (.A(_12796_),
    .B_N(\cpu.dcache.r_data[5][30] ),
    .Y(_12806_));
 sg13g2_a21oi_1 _19856_ (.A1(net1006),
    .A2(_12796_),
    .Y(_12807_),
    .B1(_12806_));
 sg13g2_nand2_1 _19857_ (.Y(_12808_),
    .A(_12110_),
    .B(_12776_));
 sg13g2_o21ai_1 _19858_ (.B1(_12808_),
    .Y(_00493_),
    .A1(net45),
    .A2(_12807_));
 sg13g2_nor2b_1 _19859_ (.A(_12796_),
    .B_N(\cpu.dcache.r_data[5][31] ),
    .Y(_12809_));
 sg13g2_a21oi_1 _19860_ (.A1(_12678_),
    .A2(_12796_),
    .Y(_12810_),
    .B1(_12809_));
 sg13g2_nand2_1 _19861_ (.Y(_12811_),
    .A(_12116_),
    .B(_12776_));
 sg13g2_o21ai_1 _19862_ (.B1(_12811_),
    .Y(_00494_),
    .A1(net45),
    .A2(_12810_));
 sg13g2_nor2b_1 _19863_ (.A(_12712_),
    .B_N(\cpu.dcache.r_data[5][3] ),
    .Y(_12812_));
 sg13g2_a21oi_1 _19864_ (.A1(net1009),
    .A2(_12712_),
    .Y(_02671_),
    .B1(_12812_));
 sg13g2_nand2_1 _19865_ (.Y(_02672_),
    .A(net1054),
    .B(_12706_));
 sg13g2_o21ai_1 _19866_ (.B1(_02672_),
    .Y(_00495_),
    .A1(net48),
    .A2(_02671_));
 sg13g2_nor2_1 _19867_ (.A(net500),
    .B(_12322_),
    .Y(_02673_));
 sg13g2_buf_2 _19868_ (.A(_02673_),
    .X(_02674_));
 sg13g2_mux2_1 _19869_ (.A0(\cpu.dcache.r_data[5][4] ),
    .A1(net1106),
    .S(_02674_),
    .X(_02675_));
 sg13g2_nor2_1 _19870_ (.A(_12706_),
    .B(_02675_),
    .Y(_02676_));
 sg13g2_a21oi_1 _19871_ (.A1(net877),
    .A2(net48),
    .Y(_00496_),
    .B1(_02676_));
 sg13g2_mux2_1 _19872_ (.A0(\cpu.dcache.r_data[5][5] ),
    .A1(net1103),
    .S(_02674_),
    .X(_02677_));
 sg13g2_nor2_1 _19873_ (.A(_12706_),
    .B(_02677_),
    .Y(_02678_));
 sg13g2_a21oi_1 _19874_ (.A1(net876),
    .A2(net48),
    .Y(_00497_),
    .B1(_02678_));
 sg13g2_mux2_1 _19875_ (.A0(\cpu.dcache.r_data[5][6] ),
    .A1(net1105),
    .S(_02674_),
    .X(_02679_));
 sg13g2_nor2_1 _19876_ (.A(_12706_),
    .B(_02679_),
    .Y(_02680_));
 sg13g2_a21oi_1 _19877_ (.A1(net875),
    .A2(_12707_),
    .Y(_00498_),
    .B1(_02680_));
 sg13g2_buf_1 _19878_ (.A(net1104),
    .X(_02681_));
 sg13g2_nor2b_1 _19879_ (.A(_02674_),
    .B_N(\cpu.dcache.r_data[5][7] ),
    .Y(_02682_));
 sg13g2_a21oi_1 _19880_ (.A1(net1005),
    .A2(_02674_),
    .Y(_02683_),
    .B1(_02682_));
 sg13g2_nand2_1 _19881_ (.Y(_02684_),
    .A(net1053),
    .B(_12706_));
 sg13g2_o21ai_1 _19882_ (.B1(_02684_),
    .Y(_00499_),
    .A1(_12707_),
    .A2(_02683_));
 sg13g2_nor2b_1 _19883_ (.A(_12720_),
    .B_N(\cpu.dcache.r_data[5][8] ),
    .Y(_02685_));
 sg13g2_a21oi_1 _19884_ (.A1(net1008),
    .A2(_12720_),
    .Y(_02686_),
    .B1(_02685_));
 sg13g2_nand2_1 _19885_ (.Y(_02687_),
    .A(_12161_),
    .B(_12717_));
 sg13g2_o21ai_1 _19886_ (.B1(_02687_),
    .Y(_00500_),
    .A1(net47),
    .A2(_02686_));
 sg13g2_nor2b_1 _19887_ (.A(_12720_),
    .B_N(\cpu.dcache.r_data[5][9] ),
    .Y(_02688_));
 sg13g2_a21oi_1 _19888_ (.A1(_12784_),
    .A2(_12720_),
    .Y(_02689_),
    .B1(_02688_));
 sg13g2_nand2_1 _19889_ (.Y(_02690_),
    .A(_12173_),
    .B(_12717_));
 sg13g2_o21ai_1 _19890_ (.B1(_02690_),
    .Y(_00501_),
    .A1(_12718_),
    .A2(_02689_));
 sg13g2_buf_1 _19891_ (.A(net625),
    .X(_02691_));
 sg13g2_buf_1 _19892_ (.A(net556),
    .X(_02692_));
 sg13g2_nand2_1 _19893_ (.Y(_02693_),
    .A(net499),
    .B(_12055_));
 sg13g2_nor2_1 _19894_ (.A(_12043_),
    .B(_02693_),
    .Y(_02694_));
 sg13g2_buf_2 _19895_ (.A(_02694_),
    .X(_02695_));
 sg13g2_buf_1 _19896_ (.A(_02695_),
    .X(_02696_));
 sg13g2_nand2_1 _19897_ (.Y(_02697_),
    .A(net706),
    .B(net915));
 sg13g2_buf_1 _19898_ (.A(_02697_),
    .X(_02698_));
 sg13g2_buf_1 _19899_ (.A(_02698_),
    .X(_02699_));
 sg13g2_nor2_1 _19900_ (.A(net498),
    .B(_12034_),
    .Y(_02700_));
 sg13g2_buf_2 _19901_ (.A(_02700_),
    .X(_02701_));
 sg13g2_nor2b_1 _19902_ (.A(_02701_),
    .B_N(\cpu.dcache.r_data[6][0] ),
    .Y(_02702_));
 sg13g2_a21oi_1 _19903_ (.A1(net1008),
    .A2(_02701_),
    .Y(_02703_),
    .B1(_02702_));
 sg13g2_buf_1 _19904_ (.A(net1062),
    .X(_02704_));
 sg13g2_nand2_1 _19905_ (.Y(_02705_),
    .A(net874),
    .B(_02696_));
 sg13g2_o21ai_1 _19906_ (.B1(_02705_),
    .Y(_00502_),
    .A1(net44),
    .A2(_02703_));
 sg13g2_nor2_1 _19907_ (.A(_12077_),
    .B(_02693_),
    .Y(_02706_));
 sg13g2_buf_2 _19908_ (.A(_02706_),
    .X(_02707_));
 sg13g2_buf_1 _19909_ (.A(_02707_),
    .X(_02708_));
 sg13g2_nor2_1 _19910_ (.A(net498),
    .B(_12062_),
    .Y(_02709_));
 sg13g2_buf_2 _19911_ (.A(_02709_),
    .X(_02710_));
 sg13g2_nor2b_1 _19912_ (.A(_02710_),
    .B_N(\cpu.dcache.r_data[6][10] ),
    .Y(_02711_));
 sg13g2_a21oi_1 _19913_ (.A1(net1006),
    .A2(_02710_),
    .Y(_02712_),
    .B1(_02711_));
 sg13g2_nand2_1 _19914_ (.Y(_02713_),
    .A(_12073_),
    .B(_02708_));
 sg13g2_o21ai_1 _19915_ (.B1(_02713_),
    .Y(_00503_),
    .A1(_02708_),
    .A2(_02712_));
 sg13g2_nor2b_1 _19916_ (.A(_02710_),
    .B_N(\cpu.dcache.r_data[6][11] ),
    .Y(_02714_));
 sg13g2_a21oi_1 _19917_ (.A1(net1005),
    .A2(_02710_),
    .Y(_02715_),
    .B1(_02714_));
 sg13g2_nand2_1 _19918_ (.Y(_02716_),
    .A(_12084_),
    .B(net43));
 sg13g2_o21ai_1 _19919_ (.B1(_02716_),
    .Y(_00504_),
    .A1(net43),
    .A2(_02715_));
 sg13g2_nor2_1 _19920_ (.A(net498),
    .B(_12089_),
    .Y(_02717_));
 sg13g2_buf_2 _19921_ (.A(_02717_),
    .X(_02718_));
 sg13g2_nor2b_1 _19922_ (.A(_02718_),
    .B_N(\cpu.dcache.r_data[6][12] ),
    .Y(_02719_));
 sg13g2_a21oi_1 _19923_ (.A1(net1008),
    .A2(_02718_),
    .Y(_02720_),
    .B1(_02719_));
 sg13g2_nand2_1 _19924_ (.Y(_02721_),
    .A(_12096_),
    .B(_02707_));
 sg13g2_o21ai_1 _19925_ (.B1(_02721_),
    .Y(_00505_),
    .A1(net43),
    .A2(_02720_));
 sg13g2_nor2b_1 _19926_ (.A(_02718_),
    .B_N(\cpu.dcache.r_data[6][13] ),
    .Y(_02722_));
 sg13g2_a21oi_1 _19927_ (.A1(_12784_),
    .A2(_02718_),
    .Y(_02723_),
    .B1(_02722_));
 sg13g2_nand2_1 _19928_ (.Y(_02724_),
    .A(_12104_),
    .B(_02707_));
 sg13g2_o21ai_1 _19929_ (.B1(_02724_),
    .Y(_00506_),
    .A1(net43),
    .A2(_02723_));
 sg13g2_nor2b_1 _19930_ (.A(_02718_),
    .B_N(\cpu.dcache.r_data[6][14] ),
    .Y(_02725_));
 sg13g2_a21oi_1 _19931_ (.A1(_12788_),
    .A2(_02718_),
    .Y(_02726_),
    .B1(_02725_));
 sg13g2_nand2_1 _19932_ (.Y(_02727_),
    .A(_12110_),
    .B(_02707_));
 sg13g2_o21ai_1 _19933_ (.B1(_02727_),
    .Y(_00507_),
    .A1(net43),
    .A2(_02726_));
 sg13g2_nor2b_1 _19934_ (.A(_02718_),
    .B_N(\cpu.dcache.r_data[6][15] ),
    .Y(_02728_));
 sg13g2_a21oi_1 _19935_ (.A1(net1005),
    .A2(_02718_),
    .Y(_02729_),
    .B1(_02728_));
 sg13g2_nand2_1 _19936_ (.Y(_02730_),
    .A(_12116_),
    .B(_02707_));
 sg13g2_o21ai_1 _19937_ (.B1(_02730_),
    .Y(_00508_),
    .A1(net43),
    .A2(_02729_));
 sg13g2_nor2_1 _19938_ (.A(_12126_),
    .B(_02693_),
    .Y(_02731_));
 sg13g2_buf_2 _19939_ (.A(_02731_),
    .X(_02732_));
 sg13g2_buf_1 _19940_ (.A(_02732_),
    .X(_02733_));
 sg13g2_nor2_1 _19941_ (.A(net498),
    .B(_12120_),
    .Y(_02734_));
 sg13g2_buf_2 _19942_ (.A(_02734_),
    .X(_02735_));
 sg13g2_nor2b_1 _19943_ (.A(_02735_),
    .B_N(\cpu.dcache.r_data[6][16] ),
    .Y(_02736_));
 sg13g2_a21oi_1 _19944_ (.A1(net1008),
    .A2(_02735_),
    .Y(_02737_),
    .B1(_02736_));
 sg13g2_nand2_1 _19945_ (.Y(_02738_),
    .A(net874),
    .B(net42));
 sg13g2_o21ai_1 _19946_ (.B1(_02738_),
    .Y(_00509_),
    .A1(net42),
    .A2(_02737_));
 sg13g2_nor2b_1 _19947_ (.A(_02735_),
    .B_N(\cpu.dcache.r_data[6][17] ),
    .Y(_02739_));
 sg13g2_a21oi_1 _19948_ (.A1(net1007),
    .A2(_02735_),
    .Y(_02740_),
    .B1(_02739_));
 sg13g2_nand2_1 _19949_ (.Y(_02741_),
    .A(net879),
    .B(net42));
 sg13g2_o21ai_1 _19950_ (.B1(_02741_),
    .Y(_00510_),
    .A1(net42),
    .A2(_02740_));
 sg13g2_nor2b_1 _19951_ (.A(_02735_),
    .B_N(\cpu.dcache.r_data[6][18] ),
    .Y(_02742_));
 sg13g2_a21oi_1 _19952_ (.A1(net1006),
    .A2(_02735_),
    .Y(_02743_),
    .B1(_02742_));
 sg13g2_nand2_1 _19953_ (.Y(_02744_),
    .A(net878),
    .B(_02732_));
 sg13g2_o21ai_1 _19954_ (.B1(_02744_),
    .Y(_00511_),
    .A1(net42),
    .A2(_02743_));
 sg13g2_nor2b_1 _19955_ (.A(_02735_),
    .B_N(\cpu.dcache.r_data[6][19] ),
    .Y(_02745_));
 sg13g2_a21oi_1 _19956_ (.A1(net1005),
    .A2(_02735_),
    .Y(_02746_),
    .B1(_02745_));
 sg13g2_nand2_1 _19957_ (.Y(_02747_),
    .A(net1054),
    .B(_02732_));
 sg13g2_o21ai_1 _19958_ (.B1(_02747_),
    .Y(_00512_),
    .A1(net42),
    .A2(_02746_));
 sg13g2_nor2b_1 _19959_ (.A(_02701_),
    .B_N(\cpu.dcache.r_data[6][1] ),
    .Y(_02748_));
 sg13g2_a21oi_1 _19960_ (.A1(net1007),
    .A2(_02701_),
    .Y(_02749_),
    .B1(_02748_));
 sg13g2_nand2_1 _19961_ (.Y(_02750_),
    .A(net879),
    .B(net44));
 sg13g2_o21ai_1 _19962_ (.B1(_02750_),
    .Y(_00513_),
    .A1(net44),
    .A2(_02749_));
 sg13g2_nor2_1 _19963_ (.A(net498),
    .B(_12268_),
    .Y(_02751_));
 sg13g2_buf_2 _19964_ (.A(_02751_),
    .X(_02752_));
 sg13g2_mux2_1 _19965_ (.A0(\cpu.dcache.r_data[6][20] ),
    .A1(net1106),
    .S(_02752_),
    .X(_02753_));
 sg13g2_nor2_1 _19966_ (.A(_02732_),
    .B(_02753_),
    .Y(_02754_));
 sg13g2_a21oi_1 _19967_ (.A1(net877),
    .A2(net42),
    .Y(_00514_),
    .B1(_02754_));
 sg13g2_mux2_1 _19968_ (.A0(\cpu.dcache.r_data[6][21] ),
    .A1(net1103),
    .S(_02752_),
    .X(_02755_));
 sg13g2_nor2_1 _19969_ (.A(_02732_),
    .B(_02755_),
    .Y(_02756_));
 sg13g2_a21oi_1 _19970_ (.A1(net876),
    .A2(net42),
    .Y(_00515_),
    .B1(_02756_));
 sg13g2_mux2_1 _19971_ (.A0(\cpu.dcache.r_data[6][22] ),
    .A1(net1105),
    .S(_02752_),
    .X(_02757_));
 sg13g2_nor2_1 _19972_ (.A(_02732_),
    .B(_02757_),
    .Y(_02758_));
 sg13g2_a21oi_1 _19973_ (.A1(net875),
    .A2(_02733_),
    .Y(_00516_),
    .B1(_02758_));
 sg13g2_nor2b_1 _19974_ (.A(_02752_),
    .B_N(\cpu.dcache.r_data[6][23] ),
    .Y(_02759_));
 sg13g2_a21oi_1 _19975_ (.A1(net1005),
    .A2(_02752_),
    .Y(_02760_),
    .B1(_02759_));
 sg13g2_nand2_1 _19976_ (.Y(_02761_),
    .A(net1053),
    .B(_02732_));
 sg13g2_o21ai_1 _19977_ (.B1(_02761_),
    .Y(_00517_),
    .A1(_02733_),
    .A2(_02760_));
 sg13g2_nor2_1 _19978_ (.A(_12166_),
    .B(_02693_),
    .Y(_02762_));
 sg13g2_buf_2 _19979_ (.A(_02762_),
    .X(_02763_));
 sg13g2_buf_1 _19980_ (.A(_02763_),
    .X(_02764_));
 sg13g2_nor2_1 _19981_ (.A(_02699_),
    .B(_12051_),
    .Y(_02765_));
 sg13g2_buf_1 _19982_ (.A(_02765_),
    .X(_02766_));
 sg13g2_nor2b_1 _19983_ (.A(net415),
    .B_N(\cpu.dcache.r_data[6][24] ),
    .Y(_02767_));
 sg13g2_a21oi_1 _19984_ (.A1(_12778_),
    .A2(net415),
    .Y(_02768_),
    .B1(_02767_));
 sg13g2_nand2_1 _19985_ (.Y(_02769_),
    .A(_12161_),
    .B(net41));
 sg13g2_o21ai_1 _19986_ (.B1(_02769_),
    .Y(_00518_),
    .A1(net41),
    .A2(_02768_));
 sg13g2_nor2b_1 _19987_ (.A(net415),
    .B_N(\cpu.dcache.r_data[6][25] ),
    .Y(_02770_));
 sg13g2_a21oi_1 _19988_ (.A1(net1007),
    .A2(net415),
    .Y(_02771_),
    .B1(_02770_));
 sg13g2_nand2_1 _19989_ (.Y(_02772_),
    .A(_12173_),
    .B(net41));
 sg13g2_o21ai_1 _19990_ (.B1(_02772_),
    .Y(_00519_),
    .A1(_02764_),
    .A2(_02771_));
 sg13g2_nor2b_1 _19991_ (.A(net415),
    .B_N(\cpu.dcache.r_data[6][26] ),
    .Y(_02773_));
 sg13g2_a21oi_1 _19992_ (.A1(net1006),
    .A2(net415),
    .Y(_02774_),
    .B1(_02773_));
 sg13g2_nand2_1 _19993_ (.Y(_02775_),
    .A(_12073_),
    .B(_02763_));
 sg13g2_o21ai_1 _19994_ (.B1(_02775_),
    .Y(_00520_),
    .A1(_02764_),
    .A2(_02774_));
 sg13g2_nor2b_1 _19995_ (.A(net415),
    .B_N(\cpu.dcache.r_data[6][27] ),
    .Y(_02776_));
 sg13g2_a21oi_1 _19996_ (.A1(net1005),
    .A2(net415),
    .Y(_02777_),
    .B1(_02776_));
 sg13g2_nand2_1 _19997_ (.Y(_02778_),
    .A(_12084_),
    .B(_02763_));
 sg13g2_o21ai_1 _19998_ (.B1(_02778_),
    .Y(_00521_),
    .A1(net41),
    .A2(_02777_));
 sg13g2_nor2_1 _19999_ (.A(net498),
    .B(_12178_),
    .Y(_02779_));
 sg13g2_buf_2 _20000_ (.A(_02779_),
    .X(_02780_));
 sg13g2_nor2b_1 _20001_ (.A(_02780_),
    .B_N(\cpu.dcache.r_data[6][28] ),
    .Y(_02781_));
 sg13g2_a21oi_1 _20002_ (.A1(_12778_),
    .A2(_02780_),
    .Y(_02782_),
    .B1(_02781_));
 sg13g2_nand2_1 _20003_ (.Y(_02783_),
    .A(_12096_),
    .B(_02763_));
 sg13g2_o21ai_1 _20004_ (.B1(_02783_),
    .Y(_00522_),
    .A1(net41),
    .A2(_02782_));
 sg13g2_nor2b_1 _20005_ (.A(_02780_),
    .B_N(\cpu.dcache.r_data[6][29] ),
    .Y(_02784_));
 sg13g2_a21oi_1 _20006_ (.A1(net1007),
    .A2(_02780_),
    .Y(_02785_),
    .B1(_02784_));
 sg13g2_nand2_1 _20007_ (.Y(_02786_),
    .A(_12104_),
    .B(_02763_));
 sg13g2_o21ai_1 _20008_ (.B1(_02786_),
    .Y(_00523_),
    .A1(net41),
    .A2(_02785_));
 sg13g2_nor2b_1 _20009_ (.A(_02701_),
    .B_N(\cpu.dcache.r_data[6][2] ),
    .Y(_02787_));
 sg13g2_a21oi_1 _20010_ (.A1(net1006),
    .A2(_02701_),
    .Y(_02788_),
    .B1(_02787_));
 sg13g2_nand2_1 _20011_ (.Y(_02789_),
    .A(net878),
    .B(_02695_));
 sg13g2_o21ai_1 _20012_ (.B1(_02789_),
    .Y(_00524_),
    .A1(net44),
    .A2(_02788_));
 sg13g2_nor2b_1 _20013_ (.A(_02780_),
    .B_N(\cpu.dcache.r_data[6][30] ),
    .Y(_02790_));
 sg13g2_a21oi_1 _20014_ (.A1(_12788_),
    .A2(_02780_),
    .Y(_02791_),
    .B1(_02790_));
 sg13g2_nand2_1 _20015_ (.Y(_02792_),
    .A(_12110_),
    .B(_02763_));
 sg13g2_o21ai_1 _20016_ (.B1(_02792_),
    .Y(_00525_),
    .A1(net41),
    .A2(_02791_));
 sg13g2_nor2b_1 _20017_ (.A(_02780_),
    .B_N(\cpu.dcache.r_data[6][31] ),
    .Y(_02793_));
 sg13g2_a21oi_1 _20018_ (.A1(_02681_),
    .A2(_02780_),
    .Y(_02794_),
    .B1(_02793_));
 sg13g2_nand2_1 _20019_ (.Y(_02795_),
    .A(_12116_),
    .B(_02763_));
 sg13g2_o21ai_1 _20020_ (.B1(_02795_),
    .Y(_00526_),
    .A1(net41),
    .A2(_02794_));
 sg13g2_nor2b_1 _20021_ (.A(_02701_),
    .B_N(\cpu.dcache.r_data[6][3] ),
    .Y(_02796_));
 sg13g2_a21oi_1 _20022_ (.A1(net1005),
    .A2(_02701_),
    .Y(_02797_),
    .B1(_02796_));
 sg13g2_nand2_1 _20023_ (.Y(_02798_),
    .A(net1054),
    .B(_02695_));
 sg13g2_o21ai_1 _20024_ (.B1(_02798_),
    .Y(_00527_),
    .A1(_02696_),
    .A2(_02797_));
 sg13g2_nor2_1 _20025_ (.A(net498),
    .B(_12322_),
    .Y(_02799_));
 sg13g2_buf_2 _20026_ (.A(_02799_),
    .X(_02800_));
 sg13g2_mux2_1 _20027_ (.A0(\cpu.dcache.r_data[6][4] ),
    .A1(net1106),
    .S(_02800_),
    .X(_02801_));
 sg13g2_nor2_1 _20028_ (.A(_02695_),
    .B(_02801_),
    .Y(_02802_));
 sg13g2_a21oi_1 _20029_ (.A1(net877),
    .A2(net44),
    .Y(_00528_),
    .B1(_02802_));
 sg13g2_mux2_1 _20030_ (.A0(\cpu.dcache.r_data[6][5] ),
    .A1(net1103),
    .S(_02800_),
    .X(_02803_));
 sg13g2_nor2_1 _20031_ (.A(_02695_),
    .B(_02803_),
    .Y(_02804_));
 sg13g2_a21oi_1 _20032_ (.A1(net876),
    .A2(net44),
    .Y(_00529_),
    .B1(_02804_));
 sg13g2_mux2_1 _20033_ (.A0(\cpu.dcache.r_data[6][6] ),
    .A1(net1105),
    .S(_02800_),
    .X(_02805_));
 sg13g2_nor2_1 _20034_ (.A(_02695_),
    .B(_02805_),
    .Y(_02806_));
 sg13g2_a21oi_1 _20035_ (.A1(net875),
    .A2(net44),
    .Y(_00530_),
    .B1(_02806_));
 sg13g2_nor2b_1 _20036_ (.A(_02800_),
    .B_N(\cpu.dcache.r_data[6][7] ),
    .Y(_02807_));
 sg13g2_a21oi_1 _20037_ (.A1(net1005),
    .A2(_02800_),
    .Y(_02808_),
    .B1(_02807_));
 sg13g2_nand2_1 _20038_ (.Y(_02809_),
    .A(net1053),
    .B(_02695_));
 sg13g2_o21ai_1 _20039_ (.B1(_02809_),
    .Y(_00531_),
    .A1(net44),
    .A2(_02808_));
 sg13g2_nor2b_1 _20040_ (.A(_02710_),
    .B_N(\cpu.dcache.r_data[6][8] ),
    .Y(_02810_));
 sg13g2_a21oi_1 _20041_ (.A1(net1008),
    .A2(_02710_),
    .Y(_02811_),
    .B1(_02810_));
 sg13g2_nand2_1 _20042_ (.Y(_02812_),
    .A(_12161_),
    .B(_02707_));
 sg13g2_o21ai_1 _20043_ (.B1(_02812_),
    .Y(_00532_),
    .A1(net43),
    .A2(_02811_));
 sg13g2_nor2b_1 _20044_ (.A(_02710_),
    .B_N(\cpu.dcache.r_data[6][9] ),
    .Y(_02813_));
 sg13g2_a21oi_1 _20045_ (.A1(net1007),
    .A2(_02710_),
    .Y(_02814_),
    .B1(_02813_));
 sg13g2_nand2_1 _20046_ (.Y(_02815_),
    .A(_12173_),
    .B(_02707_));
 sg13g2_o21ai_1 _20047_ (.B1(_02815_),
    .Y(_00533_),
    .A1(net43),
    .A2(_02814_));
 sg13g2_nand2_1 _20048_ (.Y(_02816_),
    .A(net515),
    .B(_12055_));
 sg13g2_nor2_1 _20049_ (.A(_12043_),
    .B(_02816_),
    .Y(_02817_));
 sg13g2_buf_1 _20050_ (.A(_02817_),
    .X(_02818_));
 sg13g2_buf_1 _20051_ (.A(_02818_),
    .X(_02819_));
 sg13g2_nor2_1 _20052_ (.A(net575),
    .B(_12034_),
    .Y(_02820_));
 sg13g2_buf_2 _20053_ (.A(_02820_),
    .X(_02821_));
 sg13g2_nor2b_1 _20054_ (.A(_02821_),
    .B_N(\cpu.dcache.r_data[7][0] ),
    .Y(_02822_));
 sg13g2_a21oi_1 _20055_ (.A1(net1008),
    .A2(_02821_),
    .Y(_02823_),
    .B1(_02822_));
 sg13g2_nand2_1 _20056_ (.Y(_02824_),
    .A(net874),
    .B(_02819_));
 sg13g2_o21ai_1 _20057_ (.B1(_02824_),
    .Y(_00534_),
    .A1(_02819_),
    .A2(_02823_));
 sg13g2_nor2_1 _20058_ (.A(_12077_),
    .B(_02816_),
    .Y(_02825_));
 sg13g2_buf_2 _20059_ (.A(_02825_),
    .X(_02826_));
 sg13g2_buf_1 _20060_ (.A(_02826_),
    .X(_02827_));
 sg13g2_nor2_1 _20061_ (.A(net575),
    .B(_12062_),
    .Y(_02828_));
 sg13g2_buf_2 _20062_ (.A(_02828_),
    .X(_02829_));
 sg13g2_nor2b_1 _20063_ (.A(_02829_),
    .B_N(\cpu.dcache.r_data[7][10] ),
    .Y(_02830_));
 sg13g2_a21oi_1 _20064_ (.A1(net1006),
    .A2(_02829_),
    .Y(_02831_),
    .B1(_02830_));
 sg13g2_nand2_1 _20065_ (.Y(_02832_),
    .A(_12073_),
    .B(net39));
 sg13g2_o21ai_1 _20066_ (.B1(_02832_),
    .Y(_00535_),
    .A1(net39),
    .A2(_02831_));
 sg13g2_nor2b_1 _20067_ (.A(_02829_),
    .B_N(\cpu.dcache.r_data[7][11] ),
    .Y(_02833_));
 sg13g2_a21oi_1 _20068_ (.A1(_02681_),
    .A2(_02829_),
    .Y(_02834_),
    .B1(_02833_));
 sg13g2_nand2_1 _20069_ (.Y(_02835_),
    .A(_12084_),
    .B(_02827_));
 sg13g2_o21ai_1 _20070_ (.B1(_02835_),
    .Y(_00536_),
    .A1(net39),
    .A2(_02834_));
 sg13g2_buf_2 _20071_ (.A(_12204_),
    .X(_02836_));
 sg13g2_nor2_1 _20072_ (.A(net575),
    .B(_12089_),
    .Y(_02837_));
 sg13g2_buf_2 _20073_ (.A(_02837_),
    .X(_02838_));
 sg13g2_nor2b_1 _20074_ (.A(_02838_),
    .B_N(\cpu.dcache.r_data[7][12] ),
    .Y(_02839_));
 sg13g2_a21oi_1 _20075_ (.A1(net1004),
    .A2(_02838_),
    .Y(_02840_),
    .B1(_02839_));
 sg13g2_nand2_1 _20076_ (.Y(_02841_),
    .A(_12096_),
    .B(_02826_));
 sg13g2_o21ai_1 _20077_ (.B1(_02841_),
    .Y(_00537_),
    .A1(_02827_),
    .A2(_02840_));
 sg13g2_nor2b_1 _20078_ (.A(_02838_),
    .B_N(\cpu.dcache.r_data[7][13] ),
    .Y(_02842_));
 sg13g2_a21oi_1 _20079_ (.A1(net1007),
    .A2(_02838_),
    .Y(_02843_),
    .B1(_02842_));
 sg13g2_nand2_1 _20080_ (.Y(_02844_),
    .A(_12104_),
    .B(_02826_));
 sg13g2_o21ai_1 _20081_ (.B1(_02844_),
    .Y(_00538_),
    .A1(net39),
    .A2(_02843_));
 sg13g2_buf_2 _20082_ (.A(net1105),
    .X(_02845_));
 sg13g2_nor2b_1 _20083_ (.A(_02838_),
    .B_N(\cpu.dcache.r_data[7][14] ),
    .Y(_02846_));
 sg13g2_a21oi_1 _20084_ (.A1(net1003),
    .A2(_02838_),
    .Y(_02847_),
    .B1(_02846_));
 sg13g2_nand2_1 _20085_ (.Y(_02848_),
    .A(_12110_),
    .B(_02826_));
 sg13g2_o21ai_1 _20086_ (.B1(_02848_),
    .Y(_00539_),
    .A1(net39),
    .A2(_02847_));
 sg13g2_buf_2 _20087_ (.A(_12080_),
    .X(_02849_));
 sg13g2_nor2b_1 _20088_ (.A(_02838_),
    .B_N(\cpu.dcache.r_data[7][15] ),
    .Y(_02850_));
 sg13g2_a21oi_1 _20089_ (.A1(net1099),
    .A2(_02838_),
    .Y(_02851_),
    .B1(_02850_));
 sg13g2_nand2_1 _20090_ (.Y(_02852_),
    .A(_12116_),
    .B(_02826_));
 sg13g2_o21ai_1 _20091_ (.B1(_02852_),
    .Y(_00540_),
    .A1(net39),
    .A2(_02851_));
 sg13g2_nor2_1 _20092_ (.A(_12126_),
    .B(_02816_),
    .Y(_02853_));
 sg13g2_buf_1 _20093_ (.A(_02853_),
    .X(_02854_));
 sg13g2_buf_1 _20094_ (.A(_02854_),
    .X(_02855_));
 sg13g2_nor2_1 _20095_ (.A(net575),
    .B(_12120_),
    .Y(_02856_));
 sg13g2_buf_2 _20096_ (.A(_02856_),
    .X(_02857_));
 sg13g2_nor2b_1 _20097_ (.A(_02857_),
    .B_N(\cpu.dcache.r_data[7][16] ),
    .Y(_02858_));
 sg13g2_a21oi_1 _20098_ (.A1(net1004),
    .A2(_02857_),
    .Y(_02859_),
    .B1(_02858_));
 sg13g2_nand2_1 _20099_ (.Y(_02860_),
    .A(net874),
    .B(net38));
 sg13g2_o21ai_1 _20100_ (.B1(_02860_),
    .Y(_00541_),
    .A1(net38),
    .A2(_02859_));
 sg13g2_buf_2 _20101_ (.A(_12235_),
    .X(_02861_));
 sg13g2_nor2b_1 _20102_ (.A(_02857_),
    .B_N(\cpu.dcache.r_data[7][17] ),
    .Y(_02862_));
 sg13g2_a21oi_1 _20103_ (.A1(net1002),
    .A2(_02857_),
    .Y(_02863_),
    .B1(_02862_));
 sg13g2_nand2_1 _20104_ (.Y(_02864_),
    .A(net879),
    .B(net38));
 sg13g2_o21ai_1 _20105_ (.B1(_02864_),
    .Y(_00542_),
    .A1(net38),
    .A2(_02863_));
 sg13g2_nor2b_1 _20106_ (.A(_02857_),
    .B_N(\cpu.dcache.r_data[7][18] ),
    .Y(_02865_));
 sg13g2_a21oi_1 _20107_ (.A1(net1003),
    .A2(_02857_),
    .Y(_02866_),
    .B1(_02865_));
 sg13g2_nand2_1 _20108_ (.Y(_02867_),
    .A(net878),
    .B(_02854_));
 sg13g2_o21ai_1 _20109_ (.B1(_02867_),
    .Y(_00543_),
    .A1(net38),
    .A2(_02866_));
 sg13g2_nor2b_1 _20110_ (.A(_02857_),
    .B_N(\cpu.dcache.r_data[7][19] ),
    .Y(_02868_));
 sg13g2_a21oi_1 _20111_ (.A1(net1099),
    .A2(_02857_),
    .Y(_02869_),
    .B1(_02868_));
 sg13g2_nand2_1 _20112_ (.Y(_02870_),
    .A(net1054),
    .B(_02854_));
 sg13g2_o21ai_1 _20113_ (.B1(_02870_),
    .Y(_00544_),
    .A1(net38),
    .A2(_02869_));
 sg13g2_nor2b_1 _20114_ (.A(_02821_),
    .B_N(\cpu.dcache.r_data[7][1] ),
    .Y(_02871_));
 sg13g2_a21oi_1 _20115_ (.A1(net1002),
    .A2(_02821_),
    .Y(_02872_),
    .B1(_02871_));
 sg13g2_nand2_1 _20116_ (.Y(_02873_),
    .A(net1055),
    .B(net40));
 sg13g2_o21ai_1 _20117_ (.B1(_02873_),
    .Y(_00545_),
    .A1(net40),
    .A2(_02872_));
 sg13g2_nand2_2 _20118_ (.Y(_02874_),
    .A(_09947_),
    .B(_12140_));
 sg13g2_mux2_1 _20119_ (.A0(net1102),
    .A1(\cpu.dcache.r_data[7][20] ),
    .S(_02874_),
    .X(_02875_));
 sg13g2_nor2_1 _20120_ (.A(_02854_),
    .B(_02875_),
    .Y(_02876_));
 sg13g2_a21oi_1 _20121_ (.A1(net877),
    .A2(net38),
    .Y(_00546_),
    .B1(_02876_));
 sg13g2_mux2_1 _20122_ (.A0(net1101),
    .A1(\cpu.dcache.r_data[7][21] ),
    .S(_02874_),
    .X(_02877_));
 sg13g2_nor2_1 _20123_ (.A(_02854_),
    .B(_02877_),
    .Y(_02878_));
 sg13g2_a21oi_1 _20124_ (.A1(net876),
    .A2(net38),
    .Y(_00547_),
    .B1(_02878_));
 sg13g2_mux2_1 _20125_ (.A0(net1100),
    .A1(\cpu.dcache.r_data[7][22] ),
    .S(_02874_),
    .X(_02879_));
 sg13g2_nor2_1 _20126_ (.A(_02854_),
    .B(_02879_),
    .Y(_02880_));
 sg13g2_a21oi_1 _20127_ (.A1(net875),
    .A2(_02855_),
    .Y(_00548_),
    .B1(_02880_));
 sg13g2_mux2_1 _20128_ (.A0(net1104),
    .A1(\cpu.dcache.r_data[7][23] ),
    .S(_02874_),
    .X(_02881_));
 sg13g2_mux2_1 _20129_ (.A0(_02881_),
    .A1(_12155_),
    .S(_02855_),
    .X(_00549_));
 sg13g2_nor2_1 _20130_ (.A(_12166_),
    .B(_02816_),
    .Y(_02882_));
 sg13g2_buf_2 _20131_ (.A(_02882_),
    .X(_02883_));
 sg13g2_buf_1 _20132_ (.A(_02883_),
    .X(_02884_));
 sg13g2_nor2_1 _20133_ (.A(_10044_),
    .B(_12051_),
    .Y(_02885_));
 sg13g2_buf_1 _20134_ (.A(_02885_),
    .X(_02886_));
 sg13g2_nor2b_1 _20135_ (.A(net456),
    .B_N(\cpu.dcache.r_data[7][24] ),
    .Y(_02887_));
 sg13g2_a21oi_1 _20136_ (.A1(net1004),
    .A2(net456),
    .Y(_02888_),
    .B1(_02887_));
 sg13g2_nand2_1 _20137_ (.Y(_02889_),
    .A(_12161_),
    .B(net37));
 sg13g2_o21ai_1 _20138_ (.B1(_02889_),
    .Y(_00550_),
    .A1(net37),
    .A2(_02888_));
 sg13g2_nor2b_1 _20139_ (.A(net456),
    .B_N(\cpu.dcache.r_data[7][25] ),
    .Y(_02890_));
 sg13g2_a21oi_1 _20140_ (.A1(net1002),
    .A2(net456),
    .Y(_02891_),
    .B1(_02890_));
 sg13g2_nand2_1 _20141_ (.Y(_02892_),
    .A(_12173_),
    .B(_02884_));
 sg13g2_o21ai_1 _20142_ (.B1(_02892_),
    .Y(_00551_),
    .A1(net37),
    .A2(_02891_));
 sg13g2_nor2b_1 _20143_ (.A(net456),
    .B_N(\cpu.dcache.r_data[7][26] ),
    .Y(_02893_));
 sg13g2_a21oi_1 _20144_ (.A1(net1003),
    .A2(net456),
    .Y(_02894_),
    .B1(_02893_));
 sg13g2_nand2_1 _20145_ (.Y(_02895_),
    .A(_12073_),
    .B(_02883_));
 sg13g2_o21ai_1 _20146_ (.B1(_02895_),
    .Y(_00552_),
    .A1(_02884_),
    .A2(_02894_));
 sg13g2_nor2b_1 _20147_ (.A(net456),
    .B_N(\cpu.dcache.r_data[7][27] ),
    .Y(_02896_));
 sg13g2_a21oi_1 _20148_ (.A1(net1099),
    .A2(net456),
    .Y(_02897_),
    .B1(_02896_));
 sg13g2_nand2_1 _20149_ (.Y(_02898_),
    .A(_12084_),
    .B(_02883_));
 sg13g2_o21ai_1 _20150_ (.B1(_02898_),
    .Y(_00553_),
    .A1(net37),
    .A2(_02897_));
 sg13g2_nor2_1 _20151_ (.A(net575),
    .B(_12178_),
    .Y(_02899_));
 sg13g2_buf_2 _20152_ (.A(_02899_),
    .X(_02900_));
 sg13g2_nor2b_1 _20153_ (.A(_02900_),
    .B_N(\cpu.dcache.r_data[7][28] ),
    .Y(_02901_));
 sg13g2_a21oi_1 _20154_ (.A1(net1004),
    .A2(_02900_),
    .Y(_02902_),
    .B1(_02901_));
 sg13g2_nand2_1 _20155_ (.Y(_02903_),
    .A(_12096_),
    .B(_02883_));
 sg13g2_o21ai_1 _20156_ (.B1(_02903_),
    .Y(_00554_),
    .A1(net37),
    .A2(_02902_));
 sg13g2_nor2b_1 _20157_ (.A(_02900_),
    .B_N(\cpu.dcache.r_data[7][29] ),
    .Y(_02904_));
 sg13g2_a21oi_1 _20158_ (.A1(net1002),
    .A2(_02900_),
    .Y(_02905_),
    .B1(_02904_));
 sg13g2_nand2_1 _20159_ (.Y(_02906_),
    .A(_12104_),
    .B(_02883_));
 sg13g2_o21ai_1 _20160_ (.B1(_02906_),
    .Y(_00555_),
    .A1(net37),
    .A2(_02905_));
 sg13g2_nor2b_1 _20161_ (.A(_02821_),
    .B_N(\cpu.dcache.r_data[7][2] ),
    .Y(_02907_));
 sg13g2_a21oi_1 _20162_ (.A1(net1003),
    .A2(_02821_),
    .Y(_02908_),
    .B1(_02907_));
 sg13g2_nand2_1 _20163_ (.Y(_02909_),
    .A(net910),
    .B(_02818_));
 sg13g2_o21ai_1 _20164_ (.B1(_02909_),
    .Y(_00556_),
    .A1(net40),
    .A2(_02908_));
 sg13g2_nor2b_1 _20165_ (.A(_02900_),
    .B_N(\cpu.dcache.r_data[7][30] ),
    .Y(_02910_));
 sg13g2_a21oi_1 _20166_ (.A1(net1003),
    .A2(_02900_),
    .Y(_02911_),
    .B1(_02910_));
 sg13g2_nand2_1 _20167_ (.Y(_02912_),
    .A(_12110_),
    .B(_02883_));
 sg13g2_o21ai_1 _20168_ (.B1(_02912_),
    .Y(_00557_),
    .A1(net37),
    .A2(_02911_));
 sg13g2_nor2b_1 _20169_ (.A(_02900_),
    .B_N(\cpu.dcache.r_data[7][31] ),
    .Y(_02913_));
 sg13g2_a21oi_1 _20170_ (.A1(net1099),
    .A2(_02900_),
    .Y(_02914_),
    .B1(_02913_));
 sg13g2_nand2_1 _20171_ (.Y(_02915_),
    .A(_12116_),
    .B(_02883_));
 sg13g2_o21ai_1 _20172_ (.B1(_02915_),
    .Y(_00558_),
    .A1(net37),
    .A2(_02914_));
 sg13g2_nor2b_1 _20173_ (.A(_02821_),
    .B_N(\cpu.dcache.r_data[7][3] ),
    .Y(_02916_));
 sg13g2_a21oi_1 _20174_ (.A1(net1099),
    .A2(_02821_),
    .Y(_02917_),
    .B1(_02916_));
 sg13g2_nand2_1 _20175_ (.Y(_02918_),
    .A(net1054),
    .B(_02818_));
 sg13g2_o21ai_1 _20176_ (.B1(_02918_),
    .Y(_00559_),
    .A1(net40),
    .A2(_02917_));
 sg13g2_nand2_2 _20177_ (.Y(_02919_),
    .A(_09947_),
    .B(_12187_));
 sg13g2_mux2_1 _20178_ (.A0(net1102),
    .A1(\cpu.dcache.r_data[7][4] ),
    .S(_02919_),
    .X(_02920_));
 sg13g2_nor2_1 _20179_ (.A(_02818_),
    .B(_02920_),
    .Y(_02921_));
 sg13g2_a21oi_1 _20180_ (.A1(net877),
    .A2(net40),
    .Y(_00560_),
    .B1(_02921_));
 sg13g2_mux2_1 _20181_ (.A0(net1101),
    .A1(\cpu.dcache.r_data[7][5] ),
    .S(_02919_),
    .X(_02922_));
 sg13g2_nor2_1 _20182_ (.A(_02818_),
    .B(_02922_),
    .Y(_02923_));
 sg13g2_a21oi_1 _20183_ (.A1(net876),
    .A2(net40),
    .Y(_00561_),
    .B1(_02923_));
 sg13g2_mux2_1 _20184_ (.A0(net1100),
    .A1(\cpu.dcache.r_data[7][6] ),
    .S(_02919_),
    .X(_02924_));
 sg13g2_nor2_1 _20185_ (.A(_02818_),
    .B(_02924_),
    .Y(_02925_));
 sg13g2_a21oi_1 _20186_ (.A1(net875),
    .A2(net40),
    .Y(_00562_),
    .B1(_02925_));
 sg13g2_mux2_1 _20187_ (.A0(net1104),
    .A1(\cpu.dcache.r_data[7][7] ),
    .S(_02919_),
    .X(_02926_));
 sg13g2_mux2_1 _20188_ (.A0(_02926_),
    .A1(_12155_),
    .S(net40),
    .X(_00563_));
 sg13g2_nor2b_1 _20189_ (.A(_02829_),
    .B_N(\cpu.dcache.r_data[7][8] ),
    .Y(_02927_));
 sg13g2_a21oi_1 _20190_ (.A1(net1004),
    .A2(_02829_),
    .Y(_02928_),
    .B1(_02927_));
 sg13g2_nand2_1 _20191_ (.Y(_02929_),
    .A(_12161_),
    .B(_02826_));
 sg13g2_o21ai_1 _20192_ (.B1(_02929_),
    .Y(_00564_),
    .A1(net39),
    .A2(_02928_));
 sg13g2_nor2b_1 _20193_ (.A(_02829_),
    .B_N(\cpu.dcache.r_data[7][9] ),
    .Y(_02930_));
 sg13g2_a21oi_1 _20194_ (.A1(net1002),
    .A2(_02829_),
    .Y(_02931_),
    .B1(_02930_));
 sg13g2_nand2_1 _20195_ (.Y(_02932_),
    .A(_12173_),
    .B(_02826_));
 sg13g2_o21ai_1 _20196_ (.B1(_02932_),
    .Y(_00565_),
    .A1(net39),
    .A2(_02931_));
 sg13g2_nand3_1 _20197_ (.B(_09821_),
    .C(_12052_),
    .A(_09817_),
    .Y(_02933_));
 sg13g2_buf_1 _20198_ (.A(\cpu.d_rstrobe_d ),
    .X(_02934_));
 sg13g2_nor2_1 _20199_ (.A(net1026),
    .B(_02934_),
    .Y(_02935_));
 sg13g2_nand3_1 _20200_ (.B(_12052_),
    .C(_02935_),
    .A(_12029_),
    .Y(_02936_));
 sg13g2_nand2_1 _20201_ (.Y(_02937_),
    .A(_02933_),
    .B(_02936_));
 sg13g2_buf_2 _20202_ (.A(_02937_),
    .X(_02938_));
 sg13g2_buf_1 _20203_ (.A(_12047_),
    .X(_02939_));
 sg13g2_and2_1 _20204_ (.A(_12024_),
    .B(_12026_),
    .X(_02940_));
 sg13g2_buf_1 _20205_ (.A(_02940_),
    .X(_02941_));
 sg13g2_xor2_1 _20206_ (.B(_12029_),
    .A(_02934_),
    .X(_02942_));
 sg13g2_nand3_1 _20207_ (.B(_02941_),
    .C(_02942_),
    .A(net1001),
    .Y(_02943_));
 sg13g2_and2_1 _20208_ (.A(_02943_),
    .B(_02933_),
    .X(_02944_));
 sg13g2_buf_2 _20209_ (.A(_02944_),
    .X(_02945_));
 sg13g2_nor2_1 _20210_ (.A(_12023_),
    .B(_02945_),
    .Y(_02946_));
 sg13g2_mux2_1 _20211_ (.A0(\cpu.dcache.r_dirty[0] ),
    .A1(_02938_),
    .S(_02946_),
    .X(_00566_));
 sg13g2_nor2_1 _20212_ (.A(_12207_),
    .B(_02945_),
    .Y(_02947_));
 sg13g2_mux2_1 _20213_ (.A0(\cpu.dcache.r_dirty[1] ),
    .A1(_02938_),
    .S(_02947_),
    .X(_00567_));
 sg13g2_nor2_1 _20214_ (.A(_12348_),
    .B(_02945_),
    .Y(_02948_));
 sg13g2_mux2_1 _20215_ (.A0(\cpu.dcache.r_dirty[2] ),
    .A1(_02938_),
    .S(_02948_),
    .X(_00568_));
 sg13g2_nor2_1 _20216_ (.A(_12477_),
    .B(_02945_),
    .Y(_02949_));
 sg13g2_mux2_1 _20217_ (.A0(\cpu.dcache.r_dirty[3] ),
    .A1(_02938_),
    .S(_02949_),
    .X(_00569_));
 sg13g2_nor2_1 _20218_ (.A(net684),
    .B(_02945_),
    .Y(_02950_));
 sg13g2_mux2_1 _20219_ (.A0(\cpu.dcache.r_dirty[4] ),
    .A1(_02938_),
    .S(_02950_),
    .X(_00570_));
 sg13g2_nor2_1 _20220_ (.A(_12710_),
    .B(_02945_),
    .Y(_02951_));
 sg13g2_mux2_1 _20221_ (.A0(\cpu.dcache.r_dirty[5] ),
    .A1(_02938_),
    .S(_02951_),
    .X(_00571_));
 sg13g2_nor2_1 _20222_ (.A(_02699_),
    .B(_02945_),
    .Y(_02952_));
 sg13g2_mux2_1 _20223_ (.A0(\cpu.dcache.r_dirty[6] ),
    .A1(_02938_),
    .S(_02952_),
    .X(_00572_));
 sg13g2_nor2_1 _20224_ (.A(net575),
    .B(_02945_),
    .Y(_02953_));
 sg13g2_mux2_1 _20225_ (.A0(\cpu.dcache.r_dirty[7] ),
    .A1(_02938_),
    .S(_02953_),
    .X(_00573_));
 sg13g2_buf_1 _20226_ (.A(net1043),
    .X(_02954_));
 sg13g2_buf_1 _20227_ (.A(_02954_),
    .X(_02955_));
 sg13g2_buf_1 _20228_ (.A(net611),
    .X(_02956_));
 sg13g2_nand2_1 _20229_ (.Y(_02957_),
    .A(\cpu.dcache.r_tag[0][5] ),
    .B(net611));
 sg13g2_o21ai_1 _20230_ (.B1(_02957_),
    .Y(_00577_),
    .A1(_02955_),
    .A2(net555));
 sg13g2_mux2_1 _20231_ (.A0(_09770_),
    .A1(\cpu.dcache.r_tag[0][15] ),
    .S(net555),
    .X(_00578_));
 sg13g2_mux2_1 _20232_ (.A0(net418),
    .A1(\cpu.dcache.r_tag[0][16] ),
    .S(net555),
    .X(_00579_));
 sg13g2_mux2_1 _20233_ (.A0(net420),
    .A1(\cpu.dcache.r_tag[0][17] ),
    .S(net555),
    .X(_00580_));
 sg13g2_mux2_1 _20234_ (.A0(net366),
    .A1(\cpu.dcache.r_tag[0][18] ),
    .S(net555),
    .X(_00581_));
 sg13g2_buf_1 _20235_ (.A(net611),
    .X(_02958_));
 sg13g2_mux2_1 _20236_ (.A0(net367),
    .A1(\cpu.dcache.r_tag[0][19] ),
    .S(net554),
    .X(_00582_));
 sg13g2_mux2_1 _20237_ (.A0(net368),
    .A1(\cpu.dcache.r_tag[0][20] ),
    .S(net554),
    .X(_00583_));
 sg13g2_mux2_1 _20238_ (.A0(net364),
    .A1(\cpu.dcache.r_tag[0][21] ),
    .S(net554),
    .X(_00584_));
 sg13g2_mux2_1 _20239_ (.A0(net365),
    .A1(\cpu.dcache.r_tag[0][22] ),
    .S(net554),
    .X(_00585_));
 sg13g2_mux2_1 _20240_ (.A0(net363),
    .A1(\cpu.dcache.r_tag[0][23] ),
    .S(net554),
    .X(_00586_));
 sg13g2_buf_2 _20241_ (.A(_09220_),
    .X(_02959_));
 sg13g2_buf_1 _20242_ (.A(net1000),
    .X(_02960_));
 sg13g2_buf_1 _20243_ (.A(net872),
    .X(_02961_));
 sg13g2_mux2_1 _20244_ (.A0(_02961_),
    .A1(\cpu.dcache.r_tag[0][6] ),
    .S(_02958_),
    .X(_00587_));
 sg13g2_buf_1 _20245_ (.A(_09223_),
    .X(_02962_));
 sg13g2_buf_1 _20246_ (.A(_02962_),
    .X(_02963_));
 sg13g2_nand2_1 _20247_ (.Y(_02964_),
    .A(\cpu.dcache.r_tag[0][7] ),
    .B(net611));
 sg13g2_o21ai_1 _20248_ (.B1(_02964_),
    .Y(_00588_),
    .A1(_02963_),
    .A2(net555));
 sg13g2_buf_1 _20249_ (.A(net1037),
    .X(_02965_));
 sg13g2_nand2_1 _20250_ (.Y(_02966_),
    .A(\cpu.dcache.r_tag[0][8] ),
    .B(net611));
 sg13g2_o21ai_1 _20251_ (.B1(_02966_),
    .Y(_00589_),
    .A1(_02965_),
    .A2(net555));
 sg13g2_inv_1 _20252_ (.Y(_02967_),
    .A(_10524_));
 sg13g2_buf_1 _20253_ (.A(_02967_),
    .X(_02968_));
 sg13g2_buf_1 _20254_ (.A(_02968_),
    .X(_02969_));
 sg13g2_nand2_1 _20255_ (.Y(_02970_),
    .A(\cpu.dcache.r_tag[0][9] ),
    .B(_12158_));
 sg13g2_o21ai_1 _20256_ (.B1(_02970_),
    .Y(_00590_),
    .A1(_02969_),
    .A2(_02956_));
 sg13g2_buf_1 _20257_ (.A(net889),
    .X(_02971_));
 sg13g2_nand2_1 _20258_ (.Y(_02972_),
    .A(\cpu.dcache.r_tag[0][10] ),
    .B(_12158_));
 sg13g2_o21ai_1 _20259_ (.B1(_02972_),
    .Y(_00591_),
    .A1(_02971_),
    .A2(_02956_));
 sg13g2_buf_1 _20260_ (.A(net1122),
    .X(_02973_));
 sg13g2_buf_1 _20261_ (.A(net999),
    .X(_02974_));
 sg13g2_mux2_1 _20262_ (.A0(_02974_),
    .A1(\cpu.dcache.r_tag[0][11] ),
    .S(_02958_),
    .X(_00592_));
 sg13g2_mux2_1 _20263_ (.A0(net289),
    .A1(\cpu.dcache.r_tag[0][12] ),
    .S(net554),
    .X(_00593_));
 sg13g2_mux2_1 _20264_ (.A0(net288),
    .A1(\cpu.dcache.r_tag[0][13] ),
    .S(net554),
    .X(_00594_));
 sg13g2_mux2_1 _20265_ (.A0(net421),
    .A1(\cpu.dcache.r_tag[0][14] ),
    .S(net554),
    .X(_00595_));
 sg13g2_buf_1 _20266_ (.A(net888),
    .X(_02975_));
 sg13g2_buf_2 _20267_ (.A(_02975_),
    .X(_02976_));
 sg13g2_buf_1 _20268_ (.A(net668),
    .X(_02977_));
 sg13g2_buf_1 _20269_ (.A(_12287_),
    .X(_02978_));
 sg13g2_mux2_1 _20270_ (.A0(\cpu.dcache.r_tag[1][5] ),
    .A1(net607),
    .S(net497),
    .X(_00596_));
 sg13g2_mux2_1 _20271_ (.A0(\cpu.dcache.r_tag[1][15] ),
    .A1(net419),
    .S(_02978_),
    .X(_00597_));
 sg13g2_mux2_1 _20272_ (.A0(\cpu.dcache.r_tag[1][16] ),
    .A1(_09792_),
    .S(net497),
    .X(_00598_));
 sg13g2_mux2_1 _20273_ (.A0(\cpu.dcache.r_tag[1][17] ),
    .A1(net420),
    .S(net497),
    .X(_00599_));
 sg13g2_mux2_1 _20274_ (.A0(\cpu.dcache.r_tag[1][18] ),
    .A1(_09545_),
    .S(net497),
    .X(_00600_));
 sg13g2_mux2_1 _20275_ (.A0(\cpu.dcache.r_tag[1][19] ),
    .A1(net367),
    .S(_02978_),
    .X(_00601_));
 sg13g2_mux2_1 _20276_ (.A0(\cpu.dcache.r_tag[1][20] ),
    .A1(net368),
    .S(net497),
    .X(_00602_));
 sg13g2_mux2_1 _20277_ (.A0(\cpu.dcache.r_tag[1][21] ),
    .A1(net364),
    .S(net497),
    .X(_00603_));
 sg13g2_mux2_1 _20278_ (.A0(\cpu.dcache.r_tag[1][22] ),
    .A1(net365),
    .S(net497),
    .X(_00604_));
 sg13g2_mux2_1 _20279_ (.A0(\cpu.dcache.r_tag[1][23] ),
    .A1(net363),
    .S(net497),
    .X(_00605_));
 sg13g2_buf_1 _20280_ (.A(net872),
    .X(_02979_));
 sg13g2_buf_1 _20281_ (.A(_12287_),
    .X(_02980_));
 sg13g2_mux2_1 _20282_ (.A0(\cpu.dcache.r_tag[1][6] ),
    .A1(net748),
    .S(_02980_),
    .X(_00606_));
 sg13g2_buf_1 _20283_ (.A(net1138),
    .X(_02981_));
 sg13g2_buf_1 _20284_ (.A(net998),
    .X(_02982_));
 sg13g2_mux2_1 _20285_ (.A0(\cpu.dcache.r_tag[1][7] ),
    .A1(net867),
    .S(net496),
    .X(_00607_));
 sg13g2_buf_1 _20286_ (.A(net1139),
    .X(_02983_));
 sg13g2_buf_1 _20287_ (.A(net997),
    .X(_02984_));
 sg13g2_mux2_1 _20288_ (.A0(\cpu.dcache.r_tag[1][8] ),
    .A1(net866),
    .S(net496),
    .X(_00608_));
 sg13g2_buf_1 _20289_ (.A(_10524_),
    .X(_02985_));
 sg13g2_buf_1 _20290_ (.A(net996),
    .X(_02986_));
 sg13g2_mux2_1 _20291_ (.A0(\cpu.dcache.r_tag[1][9] ),
    .A1(net865),
    .S(net496),
    .X(_00609_));
 sg13g2_buf_1 _20292_ (.A(_10392_),
    .X(_02987_));
 sg13g2_buf_1 _20293_ (.A(net995),
    .X(_02988_));
 sg13g2_mux2_1 _20294_ (.A0(\cpu.dcache.r_tag[1][10] ),
    .A1(net864),
    .S(net496),
    .X(_00610_));
 sg13g2_buf_1 _20295_ (.A(net999),
    .X(_02989_));
 sg13g2_mux2_1 _20296_ (.A0(\cpu.dcache.r_tag[1][11] ),
    .A1(net863),
    .S(_02980_),
    .X(_00611_));
 sg13g2_mux2_1 _20297_ (.A0(\cpu.dcache.r_tag[1][12] ),
    .A1(net289),
    .S(net496),
    .X(_00612_));
 sg13g2_mux2_1 _20298_ (.A0(\cpu.dcache.r_tag[1][13] ),
    .A1(net288),
    .S(net496),
    .X(_00613_));
 sg13g2_mux2_1 _20299_ (.A0(\cpu.dcache.r_tag[1][14] ),
    .A1(net421),
    .S(net496),
    .X(_00614_));
 sg13g2_buf_1 _20300_ (.A(_12418_),
    .X(_02990_));
 sg13g2_buf_1 _20301_ (.A(_12417_),
    .X(_02991_));
 sg13g2_nand2_1 _20302_ (.Y(_02992_),
    .A(net668),
    .B(_02991_));
 sg13g2_o21ai_1 _20303_ (.B1(_02992_),
    .Y(_00615_),
    .A1(_09611_),
    .A2(_02990_));
 sg13g2_mux2_1 _20304_ (.A0(\cpu.dcache.r_tag[2][15] ),
    .A1(net419),
    .S(net455),
    .X(_00616_));
 sg13g2_mux2_1 _20305_ (.A0(\cpu.dcache.r_tag[2][16] ),
    .A1(net418),
    .S(net455),
    .X(_00617_));
 sg13g2_mux2_1 _20306_ (.A0(\cpu.dcache.r_tag[2][17] ),
    .A1(net420),
    .S(_02990_),
    .X(_00618_));
 sg13g2_mux2_1 _20307_ (.A0(\cpu.dcache.r_tag[2][18] ),
    .A1(net366),
    .S(net455),
    .X(_00619_));
 sg13g2_mux2_1 _20308_ (.A0(\cpu.dcache.r_tag[2][19] ),
    .A1(net367),
    .S(net455),
    .X(_00620_));
 sg13g2_mux2_1 _20309_ (.A0(\cpu.dcache.r_tag[2][20] ),
    .A1(net368),
    .S(net455),
    .X(_00621_));
 sg13g2_mux2_1 _20310_ (.A0(\cpu.dcache.r_tag[2][21] ),
    .A1(net364),
    .S(net455),
    .X(_00622_));
 sg13g2_mux2_1 _20311_ (.A0(\cpu.dcache.r_tag[2][22] ),
    .A1(_09679_),
    .S(net495),
    .X(_00623_));
 sg13g2_mux2_1 _20312_ (.A0(\cpu.dcache.r_tag[2][23] ),
    .A1(net363),
    .S(net495),
    .X(_00624_));
 sg13g2_mux2_1 _20313_ (.A0(\cpu.dcache.r_tag[2][6] ),
    .A1(net748),
    .S(net495),
    .X(_00625_));
 sg13g2_nand2_1 _20314_ (.Y(_02993_),
    .A(net998),
    .B(net501));
 sg13g2_o21ai_1 _20315_ (.B1(_02993_),
    .Y(_00626_),
    .A1(_09635_),
    .A2(net455));
 sg13g2_nand2_1 _20316_ (.Y(_02994_),
    .A(net997),
    .B(_12418_));
 sg13g2_o21ai_1 _20317_ (.B1(_02994_),
    .Y(_00627_),
    .A1(_09624_),
    .A2(net455));
 sg13g2_mux2_1 _20318_ (.A0(\cpu.dcache.r_tag[2][9] ),
    .A1(net865),
    .S(net495),
    .X(_00628_));
 sg13g2_mux2_1 _20319_ (.A0(\cpu.dcache.r_tag[2][10] ),
    .A1(net864),
    .S(_02991_),
    .X(_00629_));
 sg13g2_mux2_1 _20320_ (.A0(\cpu.dcache.r_tag[2][11] ),
    .A1(net863),
    .S(net495),
    .X(_00630_));
 sg13g2_mux2_1 _20321_ (.A0(\cpu.dcache.r_tag[2][12] ),
    .A1(net289),
    .S(net495),
    .X(_00631_));
 sg13g2_mux2_1 _20322_ (.A0(\cpu.dcache.r_tag[2][13] ),
    .A1(net288),
    .S(net495),
    .X(_00632_));
 sg13g2_mux2_1 _20323_ (.A0(\cpu.dcache.r_tag[2][14] ),
    .A1(net421),
    .S(net495),
    .X(_00633_));
 sg13g2_buf_1 _20324_ (.A(_12541_),
    .X(_02995_));
 sg13g2_mux2_1 _20325_ (.A0(\cpu.dcache.r_tag[3][5] ),
    .A1(net607),
    .S(net274),
    .X(_00634_));
 sg13g2_mux2_1 _20326_ (.A0(\cpu.dcache.r_tag[3][15] ),
    .A1(net419),
    .S(_02995_),
    .X(_00635_));
 sg13g2_mux2_1 _20327_ (.A0(\cpu.dcache.r_tag[3][16] ),
    .A1(net418),
    .S(net274),
    .X(_00636_));
 sg13g2_mux2_1 _20328_ (.A0(\cpu.dcache.r_tag[3][17] ),
    .A1(net420),
    .S(_02995_),
    .X(_00637_));
 sg13g2_mux2_1 _20329_ (.A0(\cpu.dcache.r_tag[3][18] ),
    .A1(net366),
    .S(net274),
    .X(_00638_));
 sg13g2_mux2_1 _20330_ (.A0(\cpu.dcache.r_tag[3][19] ),
    .A1(net367),
    .S(net274),
    .X(_00639_));
 sg13g2_mux2_1 _20331_ (.A0(\cpu.dcache.r_tag[3][20] ),
    .A1(net368),
    .S(net274),
    .X(_00640_));
 sg13g2_mux2_1 _20332_ (.A0(\cpu.dcache.r_tag[3][21] ),
    .A1(net364),
    .S(net274),
    .X(_00641_));
 sg13g2_mux2_1 _20333_ (.A0(\cpu.dcache.r_tag[3][22] ),
    .A1(net365),
    .S(net274),
    .X(_00642_));
 sg13g2_mux2_1 _20334_ (.A0(\cpu.dcache.r_tag[3][23] ),
    .A1(net363),
    .S(net274),
    .X(_00643_));
 sg13g2_buf_1 _20335_ (.A(_12541_),
    .X(_02996_));
 sg13g2_mux2_1 _20336_ (.A0(\cpu.dcache.r_tag[3][6] ),
    .A1(net748),
    .S(net273),
    .X(_00644_));
 sg13g2_mux2_1 _20337_ (.A0(\cpu.dcache.r_tag[3][7] ),
    .A1(net867),
    .S(net273),
    .X(_00645_));
 sg13g2_mux2_1 _20338_ (.A0(\cpu.dcache.r_tag[3][8] ),
    .A1(net866),
    .S(net273),
    .X(_00646_));
 sg13g2_mux2_1 _20339_ (.A0(\cpu.dcache.r_tag[3][9] ),
    .A1(net865),
    .S(net273),
    .X(_00647_));
 sg13g2_mux2_1 _20340_ (.A0(\cpu.dcache.r_tag[3][10] ),
    .A1(net864),
    .S(_02996_),
    .X(_00648_));
 sg13g2_mux2_1 _20341_ (.A0(\cpu.dcache.r_tag[3][11] ),
    .A1(net863),
    .S(_02996_),
    .X(_00649_));
 sg13g2_mux2_1 _20342_ (.A0(\cpu.dcache.r_tag[3][12] ),
    .A1(net289),
    .S(net273),
    .X(_00650_));
 sg13g2_mux2_1 _20343_ (.A0(\cpu.dcache.r_tag[3][13] ),
    .A1(net288),
    .S(net273),
    .X(_00651_));
 sg13g2_mux2_1 _20344_ (.A0(\cpu.dcache.r_tag[3][14] ),
    .A1(net421),
    .S(net273),
    .X(_00652_));
 sg13g2_buf_1 _20345_ (.A(net457),
    .X(_02997_));
 sg13g2_nand2_1 _20346_ (.Y(_02998_),
    .A(\cpu.dcache.r_tag[4][5] ),
    .B(net457));
 sg13g2_o21ai_1 _20347_ (.B1(_02998_),
    .Y(_00653_),
    .A1(_02955_),
    .A2(net414));
 sg13g2_mux2_1 _20348_ (.A0(net419),
    .A1(\cpu.dcache.r_tag[4][15] ),
    .S(net414),
    .X(_00654_));
 sg13g2_mux2_1 _20349_ (.A0(net418),
    .A1(\cpu.dcache.r_tag[4][16] ),
    .S(net414),
    .X(_00655_));
 sg13g2_mux2_1 _20350_ (.A0(net420),
    .A1(\cpu.dcache.r_tag[4][17] ),
    .S(_02997_),
    .X(_00656_));
 sg13g2_mux2_1 _20351_ (.A0(net366),
    .A1(\cpu.dcache.r_tag[4][18] ),
    .S(net414),
    .X(_00657_));
 sg13g2_buf_1 _20352_ (.A(net457),
    .X(_02999_));
 sg13g2_mux2_1 _20353_ (.A0(net367),
    .A1(\cpu.dcache.r_tag[4][19] ),
    .S(net413),
    .X(_00658_));
 sg13g2_mux2_1 _20354_ (.A0(net368),
    .A1(\cpu.dcache.r_tag[4][20] ),
    .S(net413),
    .X(_00659_));
 sg13g2_mux2_1 _20355_ (.A0(net364),
    .A1(\cpu.dcache.r_tag[4][21] ),
    .S(net413),
    .X(_00660_));
 sg13g2_mux2_1 _20356_ (.A0(net365),
    .A1(\cpu.dcache.r_tag[4][22] ),
    .S(net413),
    .X(_00661_));
 sg13g2_mux2_1 _20357_ (.A0(net363),
    .A1(\cpu.dcache.r_tag[4][23] ),
    .S(net413),
    .X(_00662_));
 sg13g2_mux2_1 _20358_ (.A0(_02961_),
    .A1(\cpu.dcache.r_tag[4][6] ),
    .S(_02999_),
    .X(_00663_));
 sg13g2_nand2_1 _20359_ (.Y(_03000_),
    .A(\cpu.dcache.r_tag[4][7] ),
    .B(net457));
 sg13g2_o21ai_1 _20360_ (.B1(_03000_),
    .Y(_00664_),
    .A1(_02963_),
    .A2(net414));
 sg13g2_nand2_1 _20361_ (.Y(_03001_),
    .A(\cpu.dcache.r_tag[4][8] ),
    .B(net457));
 sg13g2_o21ai_1 _20362_ (.B1(_03001_),
    .Y(_00665_),
    .A1(_02965_),
    .A2(net414));
 sg13g2_nand2_1 _20363_ (.Y(_03002_),
    .A(\cpu.dcache.r_tag[4][9] ),
    .B(_12657_));
 sg13g2_o21ai_1 _20364_ (.B1(_03002_),
    .Y(_00666_),
    .A1(_02969_),
    .A2(net414));
 sg13g2_nand2_1 _20365_ (.Y(_03003_),
    .A(\cpu.dcache.r_tag[4][10] ),
    .B(_12657_));
 sg13g2_o21ai_1 _20366_ (.B1(_03003_),
    .Y(_00667_),
    .A1(net750),
    .A2(_02997_));
 sg13g2_mux2_1 _20367_ (.A0(net868),
    .A1(\cpu.dcache.r_tag[4][11] ),
    .S(_02999_),
    .X(_00668_));
 sg13g2_mux2_1 _20368_ (.A0(net289),
    .A1(\cpu.dcache.r_tag[4][12] ),
    .S(net413),
    .X(_00669_));
 sg13g2_mux2_1 _20369_ (.A0(net288),
    .A1(\cpu.dcache.r_tag[4][13] ),
    .S(net413),
    .X(_00670_));
 sg13g2_mux2_1 _20370_ (.A0(net421),
    .A1(\cpu.dcache.r_tag[4][14] ),
    .S(net413),
    .X(_00671_));
 sg13g2_buf_1 _20371_ (.A(_12780_),
    .X(_03004_));
 sg13g2_mux2_1 _20372_ (.A0(\cpu.dcache.r_tag[5][5] ),
    .A1(net607),
    .S(net357),
    .X(_00672_));
 sg13g2_mux2_1 _20373_ (.A0(\cpu.dcache.r_tag[5][15] ),
    .A1(net419),
    .S(net357),
    .X(_00673_));
 sg13g2_mux2_1 _20374_ (.A0(\cpu.dcache.r_tag[5][16] ),
    .A1(net418),
    .S(net357),
    .X(_00674_));
 sg13g2_mux2_1 _20375_ (.A0(\cpu.dcache.r_tag[5][17] ),
    .A1(net420),
    .S(net357),
    .X(_00675_));
 sg13g2_mux2_1 _20376_ (.A0(\cpu.dcache.r_tag[5][18] ),
    .A1(net366),
    .S(_03004_),
    .X(_00676_));
 sg13g2_mux2_1 _20377_ (.A0(\cpu.dcache.r_tag[5][19] ),
    .A1(net367),
    .S(net357),
    .X(_00677_));
 sg13g2_mux2_1 _20378_ (.A0(\cpu.dcache.r_tag[5][20] ),
    .A1(net368),
    .S(net357),
    .X(_00678_));
 sg13g2_mux2_1 _20379_ (.A0(\cpu.dcache.r_tag[5][21] ),
    .A1(_09701_),
    .S(net357),
    .X(_00679_));
 sg13g2_mux2_1 _20380_ (.A0(\cpu.dcache.r_tag[5][22] ),
    .A1(net365),
    .S(_03004_),
    .X(_00680_));
 sg13g2_mux2_1 _20381_ (.A0(\cpu.dcache.r_tag[5][23] ),
    .A1(net363),
    .S(net357),
    .X(_00681_));
 sg13g2_buf_1 _20382_ (.A(_12780_),
    .X(_03005_));
 sg13g2_mux2_1 _20383_ (.A0(\cpu.dcache.r_tag[5][6] ),
    .A1(_02979_),
    .S(net356),
    .X(_00682_));
 sg13g2_mux2_1 _20384_ (.A0(\cpu.dcache.r_tag[5][7] ),
    .A1(net867),
    .S(net356),
    .X(_00683_));
 sg13g2_mux2_1 _20385_ (.A0(\cpu.dcache.r_tag[5][8] ),
    .A1(net866),
    .S(net356),
    .X(_00684_));
 sg13g2_mux2_1 _20386_ (.A0(\cpu.dcache.r_tag[5][9] ),
    .A1(net865),
    .S(_03005_),
    .X(_00685_));
 sg13g2_mux2_1 _20387_ (.A0(\cpu.dcache.r_tag[5][10] ),
    .A1(net864),
    .S(net356),
    .X(_00686_));
 sg13g2_mux2_1 _20388_ (.A0(\cpu.dcache.r_tag[5][11] ),
    .A1(_02989_),
    .S(_03005_),
    .X(_00687_));
 sg13g2_mux2_1 _20389_ (.A0(\cpu.dcache.r_tag[5][12] ),
    .A1(net289),
    .S(net356),
    .X(_00688_));
 sg13g2_mux2_1 _20390_ (.A0(\cpu.dcache.r_tag[5][13] ),
    .A1(net288),
    .S(net356),
    .X(_00689_));
 sg13g2_mux2_1 _20391_ (.A0(\cpu.dcache.r_tag[5][14] ),
    .A1(net421),
    .S(net356),
    .X(_00690_));
 sg13g2_buf_1 _20392_ (.A(_02766_),
    .X(_03006_));
 sg13g2_mux2_1 _20393_ (.A0(\cpu.dcache.r_tag[6][5] ),
    .A1(net607),
    .S(net355),
    .X(_00691_));
 sg13g2_mux2_1 _20394_ (.A0(\cpu.dcache.r_tag[6][15] ),
    .A1(net419),
    .S(net355),
    .X(_00692_));
 sg13g2_mux2_1 _20395_ (.A0(\cpu.dcache.r_tag[6][16] ),
    .A1(_09792_),
    .S(net355),
    .X(_00693_));
 sg13g2_mux2_1 _20396_ (.A0(\cpu.dcache.r_tag[6][17] ),
    .A1(_09723_),
    .S(_03006_),
    .X(_00694_));
 sg13g2_mux2_1 _20397_ (.A0(\cpu.dcache.r_tag[6][18] ),
    .A1(_09545_),
    .S(net355),
    .X(_00695_));
 sg13g2_mux2_1 _20398_ (.A0(\cpu.dcache.r_tag[6][19] ),
    .A1(_09522_),
    .S(_03006_),
    .X(_00696_));
 sg13g2_mux2_1 _20399_ (.A0(\cpu.dcache.r_tag[6][20] ),
    .A1(_09493_),
    .S(net355),
    .X(_00697_));
 sg13g2_mux2_1 _20400_ (.A0(\cpu.dcache.r_tag[6][21] ),
    .A1(net364),
    .S(net355),
    .X(_00698_));
 sg13g2_mux2_1 _20401_ (.A0(\cpu.dcache.r_tag[6][22] ),
    .A1(net365),
    .S(net355),
    .X(_00699_));
 sg13g2_mux2_1 _20402_ (.A0(\cpu.dcache.r_tag[6][23] ),
    .A1(_09857_),
    .S(net355),
    .X(_00700_));
 sg13g2_buf_1 _20403_ (.A(_02766_),
    .X(_03007_));
 sg13g2_mux2_1 _20404_ (.A0(\cpu.dcache.r_tag[6][6] ),
    .A1(_02979_),
    .S(net354),
    .X(_00701_));
 sg13g2_mux2_1 _20405_ (.A0(\cpu.dcache.r_tag[6][7] ),
    .A1(net867),
    .S(net354),
    .X(_00702_));
 sg13g2_mux2_1 _20406_ (.A0(\cpu.dcache.r_tag[6][8] ),
    .A1(net866),
    .S(net354),
    .X(_00703_));
 sg13g2_mux2_1 _20407_ (.A0(\cpu.dcache.r_tag[6][9] ),
    .A1(net865),
    .S(net354),
    .X(_00704_));
 sg13g2_mux2_1 _20408_ (.A0(\cpu.dcache.r_tag[6][10] ),
    .A1(net864),
    .S(_03007_),
    .X(_00705_));
 sg13g2_mux2_1 _20409_ (.A0(\cpu.dcache.r_tag[6][11] ),
    .A1(_02989_),
    .S(_03007_),
    .X(_00706_));
 sg13g2_mux2_1 _20410_ (.A0(\cpu.dcache.r_tag[6][12] ),
    .A1(net289),
    .S(net354),
    .X(_00707_));
 sg13g2_mux2_1 _20411_ (.A0(\cpu.dcache.r_tag[6][13] ),
    .A1(net288),
    .S(net354),
    .X(_00708_));
 sg13g2_mux2_1 _20412_ (.A0(\cpu.dcache.r_tag[6][14] ),
    .A1(net421),
    .S(net354),
    .X(_00709_));
 sg13g2_buf_1 _20413_ (.A(_02886_),
    .X(_03008_));
 sg13g2_mux2_1 _20414_ (.A0(\cpu.dcache.r_tag[7][5] ),
    .A1(net607),
    .S(net412),
    .X(_00710_));
 sg13g2_mux2_1 _20415_ (.A0(\cpu.dcache.r_tag[7][15] ),
    .A1(net419),
    .S(net412),
    .X(_00711_));
 sg13g2_mux2_1 _20416_ (.A0(\cpu.dcache.r_tag[7][16] ),
    .A1(net418),
    .S(_03008_),
    .X(_00712_));
 sg13g2_mux2_1 _20417_ (.A0(\cpu.dcache.r_tag[7][17] ),
    .A1(_09723_),
    .S(net412),
    .X(_00713_));
 sg13g2_mux2_1 _20418_ (.A0(\cpu.dcache.r_tag[7][18] ),
    .A1(net366),
    .S(net412),
    .X(_00714_));
 sg13g2_mux2_1 _20419_ (.A0(\cpu.dcache.r_tag[7][19] ),
    .A1(_09522_),
    .S(_03008_),
    .X(_00715_));
 sg13g2_mux2_1 _20420_ (.A0(\cpu.dcache.r_tag[7][20] ),
    .A1(net368),
    .S(net412),
    .X(_00716_));
 sg13g2_mux2_1 _20421_ (.A0(\cpu.dcache.r_tag[7][21] ),
    .A1(net364),
    .S(net412),
    .X(_00717_));
 sg13g2_mux2_1 _20422_ (.A0(\cpu.dcache.r_tag[7][22] ),
    .A1(net365),
    .S(net412),
    .X(_00718_));
 sg13g2_mux2_1 _20423_ (.A0(\cpu.dcache.r_tag[7][23] ),
    .A1(_09857_),
    .S(net412),
    .X(_00719_));
 sg13g2_buf_1 _20424_ (.A(net872),
    .X(_03009_));
 sg13g2_buf_1 _20425_ (.A(_02886_),
    .X(_03010_));
 sg13g2_mux2_1 _20426_ (.A0(\cpu.dcache.r_tag[7][6] ),
    .A1(net747),
    .S(net411),
    .X(_00720_));
 sg13g2_mux2_1 _20427_ (.A0(\cpu.dcache.r_tag[7][7] ),
    .A1(net867),
    .S(net411),
    .X(_00721_));
 sg13g2_mux2_1 _20428_ (.A0(\cpu.dcache.r_tag[7][8] ),
    .A1(net866),
    .S(net411),
    .X(_00722_));
 sg13g2_mux2_1 _20429_ (.A0(\cpu.dcache.r_tag[7][9] ),
    .A1(net865),
    .S(_03010_),
    .X(_00723_));
 sg13g2_mux2_1 _20430_ (.A0(\cpu.dcache.r_tag[7][10] ),
    .A1(net864),
    .S(net411),
    .X(_00724_));
 sg13g2_buf_1 _20431_ (.A(net999),
    .X(_03011_));
 sg13g2_mux2_1 _20432_ (.A0(\cpu.dcache.r_tag[7][11] ),
    .A1(net862),
    .S(_03010_),
    .X(_00725_));
 sg13g2_mux2_1 _20433_ (.A0(\cpu.dcache.r_tag[7][12] ),
    .A1(net289),
    .S(net411),
    .X(_00726_));
 sg13g2_mux2_1 _20434_ (.A0(\cpu.dcache.r_tag[7][13] ),
    .A1(net288),
    .S(net411),
    .X(_00727_));
 sg13g2_mux2_1 _20435_ (.A0(\cpu.dcache.r_tag[7][14] ),
    .A1(net421),
    .S(net411),
    .X(_00728_));
 sg13g2_inv_1 _20436_ (.Y(_03012_),
    .A(_09026_));
 sg13g2_buf_1 _20437_ (.A(_03012_),
    .X(_03013_));
 sg13g2_inv_1 _20438_ (.Y(_03014_),
    .A(net293));
 sg13g2_nand2_2 _20439_ (.Y(_03015_),
    .A(net231),
    .B(_09894_));
 sg13g2_inv_1 _20440_ (.Y(_03016_),
    .A(_08971_));
 sg13g2_nand2_1 _20441_ (.Y(_03017_),
    .A(_03016_),
    .B(_09003_));
 sg13g2_buf_1 _20442_ (.A(_03017_),
    .X(_03018_));
 sg13g2_o21ai_1 _20443_ (.B1(_03018_),
    .Y(_03019_),
    .A1(_09045_),
    .A2(_03015_));
 sg13g2_buf_1 _20444_ (.A(_03019_),
    .X(_03020_));
 sg13g2_buf_1 _20445_ (.A(_09045_),
    .X(_03021_));
 sg13g2_nor2_1 _20446_ (.A(_03012_),
    .B(_03021_),
    .Y(_03022_));
 sg13g2_buf_1 _20447_ (.A(_03022_),
    .X(_03023_));
 sg13g2_buf_1 _20448_ (.A(_08902_),
    .X(_03024_));
 sg13g2_a221oi_1 _20449_ (.B2(net126),
    .C1(net166),
    .B1(_03023_),
    .A1(net196),
    .Y(_03025_),
    .A2(_03020_));
 sg13g2_a21oi_1 _20450_ (.A1(net758),
    .A2(net143),
    .Y(_00737_),
    .B1(_03025_));
 sg13g2_buf_1 _20451_ (.A(_09003_),
    .X(_03026_));
 sg13g2_buf_1 _20452_ (.A(net353),
    .X(_03027_));
 sg13g2_buf_1 _20453_ (.A(net214),
    .X(_03028_));
 sg13g2_a21oi_1 _20454_ (.A1(net195),
    .A2(net291),
    .Y(_03029_),
    .B1(net196));
 sg13g2_nor2_1 _20455_ (.A(net231),
    .B(net214),
    .Y(_03030_));
 sg13g2_nor2_1 _20456_ (.A(_03029_),
    .B(_03030_),
    .Y(_03031_));
 sg13g2_buf_1 _20457_ (.A(_08971_),
    .X(_03032_));
 sg13g2_buf_1 _20458_ (.A(net230),
    .X(_03033_));
 sg13g2_nand2_1 _20459_ (.Y(_03034_),
    .A(net230),
    .B(net196));
 sg13g2_nor2_1 _20460_ (.A(_08987_),
    .B(_09004_),
    .Y(_03035_));
 sg13g2_buf_2 _20461_ (.A(_03035_),
    .X(_03036_));
 sg13g2_a22oi_1 _20462_ (.Y(_03037_),
    .B1(_03034_),
    .B2(_03036_),
    .A2(net171),
    .A1(net213));
 sg13g2_o21ai_1 _20463_ (.B1(_03037_),
    .Y(_03038_),
    .A1(net272),
    .A2(_03031_));
 sg13g2_nor2_1 _20464_ (.A(net166),
    .B(_03038_),
    .Y(_03039_));
 sg13g2_a21oi_1 _20465_ (.A1(_09213_),
    .A2(net143),
    .Y(_00738_),
    .B1(_03039_));
 sg13g2_nand2_1 _20466_ (.Y(_03040_),
    .A(_03012_),
    .B(_09045_));
 sg13g2_buf_2 _20467_ (.A(_03040_),
    .X(_03041_));
 sg13g2_buf_1 _20468_ (.A(_03018_),
    .X(_03042_));
 sg13g2_nor3_1 _20469_ (.A(net172),
    .B(_03041_),
    .C(net165),
    .Y(_03043_));
 sg13g2_a21o_1 _20470_ (.A2(net148),
    .A1(\cpu.cond[1] ),
    .B1(_03043_),
    .X(_00739_));
 sg13g2_a21oi_1 _20471_ (.A1(_03027_),
    .A2(_03034_),
    .Y(_03044_),
    .B1(net195));
 sg13g2_buf_1 _20472_ (.A(_08902_),
    .X(_03045_));
 sg13g2_mux2_1 _20473_ (.A0(_03044_),
    .A1(\cpu.cond[2] ),
    .S(_03045_),
    .X(_00740_));
 sg13g2_nand3_1 _20474_ (.B(net170),
    .C(_09144_),
    .A(_09138_),
    .Y(_03046_));
 sg13g2_o21ai_1 _20475_ (.B1(_03046_),
    .Y(_00741_),
    .A1(_09339_),
    .A2(net150));
 sg13g2_nor2_1 _20476_ (.A(_03016_),
    .B(_09006_),
    .Y(_03047_));
 sg13g2_buf_2 _20477_ (.A(_03047_),
    .X(_03048_));
 sg13g2_nand2_1 _20478_ (.Y(_03049_),
    .A(_09125_),
    .B(_03048_));
 sg13g2_buf_1 _20479_ (.A(_03049_),
    .X(_03050_));
 sg13g2_inv_1 _20480_ (.Y(_03051_),
    .A(_00159_));
 sg13g2_mux2_1 _20481_ (.A0(\cpu.icache.r_data[4][24] ),
    .A1(\cpu.icache.r_data[6][24] ),
    .S(net819),
    .X(_03052_));
 sg13g2_a22oi_1 _20482_ (.Y(_03053_),
    .B1(_03052_),
    .B2(net935),
    .A2(_08948_),
    .A1(\cpu.icache.r_data[5][24] ));
 sg13g2_mux2_1 _20483_ (.A0(\cpu.icache.r_data[7][24] ),
    .A1(\cpu.icache.r_data[3][24] ),
    .S(net938),
    .X(_03054_));
 sg13g2_a22oi_1 _20484_ (.Y(_03055_),
    .B1(net820),
    .B2(_03054_),
    .A2(net723),
    .A1(\cpu.icache.r_data[1][24] ));
 sg13g2_o21ai_1 _20485_ (.B1(_03055_),
    .Y(_03056_),
    .A1(_08535_),
    .A2(_03053_));
 sg13g2_a221oi_1 _20486_ (.B2(\cpu.icache.r_data[2][24] ),
    .C1(_03056_),
    .B1(net643),
    .A1(_03051_),
    .Y(_03057_),
    .A2(net637));
 sg13g2_nand2_1 _20487_ (.Y(_03058_),
    .A(_00158_),
    .B(net637));
 sg13g2_mux4_1 _20488_ (.S0(_08608_),
    .A0(\cpu.icache.r_data[4][8] ),
    .A1(\cpu.icache.r_data[5][8] ),
    .A2(\cpu.icache.r_data[6][8] ),
    .A3(\cpu.icache.r_data[7][8] ),
    .S1(net813),
    .X(_03059_));
 sg13g2_nand2_1 _20489_ (.Y(_03060_),
    .A(net812),
    .B(_03059_));
 sg13g2_nand2_1 _20490_ (.Y(_03061_),
    .A(\cpu.icache.r_data[1][8] ),
    .B(net639));
 sg13g2_a22oi_1 _20491_ (.Y(_03062_),
    .B1(_08530_),
    .B2(\cpu.icache.r_data[3][8] ),
    .A2(net725),
    .A1(\cpu.icache.r_data[2][8] ));
 sg13g2_nand4_1 _20492_ (.B(_03060_),
    .C(_03061_),
    .A(net582),
    .Y(_03063_),
    .D(_03062_));
 sg13g2_a21oi_1 _20493_ (.A1(_03058_),
    .A2(_03063_),
    .Y(_03064_),
    .B1(net1075));
 sg13g2_a21o_1 _20494_ (.A2(_03057_),
    .A1(_08968_),
    .B1(_03064_),
    .X(_03065_));
 sg13g2_buf_2 _20495_ (.A(_03065_),
    .X(_03066_));
 sg13g2_inv_1 _20496_ (.Y(_03067_),
    .A(_00161_));
 sg13g2_mux2_1 _20497_ (.A0(\cpu.icache.r_data[4][25] ),
    .A1(\cpu.icache.r_data[6][25] ),
    .S(_08541_),
    .X(_03068_));
 sg13g2_a22oi_1 _20498_ (.Y(_03069_),
    .B1(_03068_),
    .B2(net935),
    .A2(_08948_),
    .A1(\cpu.icache.r_data[5][25] ));
 sg13g2_mux2_1 _20499_ (.A0(\cpu.icache.r_data[7][25] ),
    .A1(\cpu.icache.r_data[3][25] ),
    .S(net938),
    .X(_03070_));
 sg13g2_a22oi_1 _20500_ (.Y(_03071_),
    .B1(net937),
    .B2(_03070_),
    .A2(net713),
    .A1(\cpu.icache.r_data[1][25] ));
 sg13g2_o21ai_1 _20501_ (.B1(_03071_),
    .Y(_03072_),
    .A1(_08535_),
    .A2(_03069_));
 sg13g2_a221oi_1 _20502_ (.B2(\cpu.icache.r_data[2][25] ),
    .C1(_03072_),
    .B1(net638),
    .A1(_03067_),
    .Y(_03073_),
    .A2(_08913_));
 sg13g2_nand2_1 _20503_ (.Y(_03074_),
    .A(_00160_),
    .B(_08913_));
 sg13g2_mux4_1 _20504_ (.S0(net1079),
    .A0(\cpu.icache.r_data[4][9] ),
    .A1(\cpu.icache.r_data[5][9] ),
    .A2(\cpu.icache.r_data[6][9] ),
    .A3(\cpu.icache.r_data[7][9] ),
    .S1(net819),
    .X(_03075_));
 sg13g2_nand2_1 _20505_ (.Y(_03076_),
    .A(net812),
    .B(_03075_));
 sg13g2_nand2_1 _20506_ (.Y(_03077_),
    .A(\cpu.icache.r_data[1][9] ),
    .B(net713));
 sg13g2_a22oi_1 _20507_ (.Y(_03078_),
    .B1(net722),
    .B2(\cpu.icache.r_data[3][9] ),
    .A2(net712),
    .A1(\cpu.icache.r_data[2][9] ));
 sg13g2_nand4_1 _20508_ (.B(_03076_),
    .C(_03077_),
    .A(net644),
    .Y(_03079_),
    .D(_03078_));
 sg13g2_a21oi_1 _20509_ (.A1(_03074_),
    .A2(_03079_),
    .Y(_03080_),
    .B1(net1075));
 sg13g2_a21oi_1 _20510_ (.A1(_08967_),
    .A2(_03073_),
    .Y(_03081_),
    .B1(_03080_));
 sg13g2_buf_2 _20511_ (.A(_03081_),
    .X(_03082_));
 sg13g2_mux4_1 _20512_ (.S0(_08824_),
    .A0(\cpu.icache.r_data[4][23] ),
    .A1(\cpu.icache.r_data[5][23] ),
    .A2(\cpu.icache.r_data[6][23] ),
    .A3(\cpu.icache.r_data[7][23] ),
    .S1(net710),
    .X(_03083_));
 sg13g2_and2_1 _20513_ (.A(\cpu.icache.r_data[3][23] ),
    .B(net722),
    .X(_03084_));
 sg13g2_a221oi_1 _20514_ (.B2(\cpu.icache.r_data[1][23] ),
    .C1(_03084_),
    .B1(net723),
    .A1(\cpu.icache.r_data[2][23] ),
    .Y(_03085_),
    .A2(net725));
 sg13g2_o21ai_1 _20515_ (.B1(_03085_),
    .Y(_03086_),
    .A1(_00157_),
    .A2(net582));
 sg13g2_a21oi_1 _20516_ (.A1(net715),
    .A2(_03083_),
    .Y(_03087_),
    .B1(_03086_));
 sg13g2_nand2_1 _20517_ (.Y(_03088_),
    .A(_00156_),
    .B(net637));
 sg13g2_a22oi_1 _20518_ (.Y(_03089_),
    .B1(net639),
    .B2(\cpu.icache.r_data[1][7] ),
    .A2(net725),
    .A1(\cpu.icache.r_data[2][7] ));
 sg13g2_a22oi_1 _20519_ (.Y(_03090_),
    .B1(net641),
    .B2(\cpu.icache.r_data[3][7] ),
    .A2(net822),
    .A1(\cpu.icache.r_data[5][7] ));
 sg13g2_mux2_1 _20520_ (.A0(\cpu.icache.r_data[4][7] ),
    .A1(\cpu.icache.r_data[6][7] ),
    .S(net936),
    .X(_03091_));
 sg13g2_a22oi_1 _20521_ (.Y(_03092_),
    .B1(_03091_),
    .B2(net935),
    .A2(net937),
    .A1(\cpu.icache.r_data[7][7] ));
 sg13g2_or2_1 _20522_ (.X(_03093_),
    .B(_03092_),
    .A(net817));
 sg13g2_nand4_1 _20523_ (.B(_03089_),
    .C(_03090_),
    .A(net582),
    .Y(_03094_),
    .D(_03093_));
 sg13g2_a21oi_1 _20524_ (.A1(_03088_),
    .A2(_03094_),
    .Y(_03095_),
    .B1(net1075));
 sg13g2_a21oi_1 _20525_ (.A1(net1075),
    .A2(_03087_),
    .Y(_03096_),
    .B1(_03095_));
 sg13g2_nor2_1 _20526_ (.A(_03082_),
    .B(_03096_),
    .Y(_03097_));
 sg13g2_nand2_1 _20527_ (.Y(_03098_),
    .A(_03066_),
    .B(_03097_));
 sg13g2_nand3_1 _20528_ (.B(_09083_),
    .C(_09121_),
    .A(_09067_),
    .Y(_03099_));
 sg13g2_or2_1 _20529_ (.X(_03100_),
    .B(_03099_),
    .A(_03098_));
 sg13g2_buf_1 _20530_ (.A(_03100_),
    .X(_03101_));
 sg13g2_inv_1 _20531_ (.Y(_03102_),
    .A(_00167_));
 sg13g2_mux2_1 _20532_ (.A0(\cpu.icache.r_data[4][20] ),
    .A1(\cpu.icache.r_data[6][20] ),
    .S(net813),
    .X(_03103_));
 sg13g2_a22oi_1 _20533_ (.Y(_03104_),
    .B1(_03103_),
    .B2(net805),
    .A2(net806),
    .A1(\cpu.icache.r_data[5][20] ));
 sg13g2_mux2_1 _20534_ (.A0(\cpu.icache.r_data[7][20] ),
    .A1(\cpu.icache.r_data[3][20] ),
    .S(net821),
    .X(_03105_));
 sg13g2_a22oi_1 _20535_ (.Y(_03106_),
    .B1(net820),
    .B2(_03105_),
    .A2(net579),
    .A1(\cpu.icache.r_data[1][20] ));
 sg13g2_o21ai_1 _20536_ (.B1(_03106_),
    .Y(_03107_),
    .A1(net721),
    .A2(_03104_));
 sg13g2_a221oi_1 _20537_ (.B2(\cpu.icache.r_data[2][20] ),
    .C1(_03107_),
    .B1(net581),
    .A1(_03102_),
    .Y(_03108_),
    .A2(net580));
 sg13g2_nand2_1 _20538_ (.Y(_03109_),
    .A(_00166_),
    .B(_08959_));
 sg13g2_mux4_1 _20539_ (.S0(net932),
    .A0(\cpu.icache.r_data[4][4] ),
    .A1(\cpu.icache.r_data[5][4] ),
    .A2(\cpu.icache.r_data[6][4] ),
    .A3(\cpu.icache.r_data[7][4] ),
    .S1(net716),
    .X(_03110_));
 sg13g2_nand2_1 _20540_ (.Y(_03111_),
    .A(net715),
    .B(_03110_));
 sg13g2_nand2_1 _20541_ (.Y(_03112_),
    .A(\cpu.icache.r_data[1][4] ),
    .B(_09010_));
 sg13g2_a22oi_1 _20542_ (.Y(_03113_),
    .B1(net583),
    .B2(\cpu.icache.r_data[3][4] ),
    .A2(net643),
    .A1(\cpu.icache.r_data[2][4] ));
 sg13g2_nand4_1 _20543_ (.B(_03111_),
    .C(_03112_),
    .A(net520),
    .Y(_03114_),
    .D(_03113_));
 sg13g2_a21oi_1 _20544_ (.A1(_03109_),
    .A2(_03114_),
    .Y(_03115_),
    .B1(net929));
 sg13g2_a21oi_1 _20545_ (.A1(net929),
    .A2(_03108_),
    .Y(_03116_),
    .B1(_03115_));
 sg13g2_buf_2 _20546_ (.A(_03116_),
    .X(_03117_));
 sg13g2_nor4_1 _20547_ (.A(_09143_),
    .B(_03050_),
    .C(_03101_),
    .D(_03117_),
    .Y(_03118_));
 sg13g2_mux2_1 _20548_ (.A0(_03118_),
    .A1(\cpu.dec.do_flush_all ),
    .S(net164),
    .X(_00742_));
 sg13g2_buf_1 _20549_ (.A(_03016_),
    .X(_03119_));
 sg13g2_nor2_1 _20550_ (.A(_08987_),
    .B(_09003_),
    .Y(_03120_));
 sg13g2_nand2_1 _20551_ (.Y(_03121_),
    .A(_03119_),
    .B(_03120_));
 sg13g2_nor3_1 _20552_ (.A(net172),
    .B(_03041_),
    .C(_03121_),
    .Y(_03122_));
 sg13g2_a21o_1 _20553_ (.A2(net148),
    .A1(\cpu.dec.do_flush_write ),
    .B1(_03122_),
    .X(_00743_));
 sg13g2_nand2_1 _20554_ (.Y(_03123_),
    .A(net225),
    .B(net214));
 sg13g2_buf_1 _20555_ (.A(_03123_),
    .X(_03124_));
 sg13g2_nand2_1 _20556_ (.Y(_03125_),
    .A(net293),
    .B(net171));
 sg13g2_a21oi_1 _20557_ (.A1(net163),
    .A2(_03125_),
    .Y(_03126_),
    .B1(net272));
 sg13g2_buf_1 _20558_ (.A(net225),
    .X(_03127_));
 sg13g2_nor2_1 _20559_ (.A(net231),
    .B(net225),
    .Y(_03128_));
 sg13g2_a22oi_1 _20560_ (.Y(_03129_),
    .B1(_03128_),
    .B2(net230),
    .A2(_03036_),
    .A1(net194));
 sg13g2_nor2_1 _20561_ (.A(net195),
    .B(_03129_),
    .Y(_03130_));
 sg13g2_o21ai_1 _20562_ (.B1(net369),
    .Y(_03131_),
    .A1(_03126_),
    .A2(_03130_));
 sg13g2_nand2_1 _20563_ (.Y(_03132_),
    .A(\cpu.icache.r_data[5][2] ),
    .B(net724));
 sg13g2_a22oi_1 _20564_ (.Y(_03133_),
    .B1(_08639_),
    .B2(\cpu.icache.r_data[7][2] ),
    .A2(net719),
    .A1(\cpu.icache.r_data[4][2] ));
 sg13g2_a22oi_1 _20565_ (.Y(_03134_),
    .B1(net720),
    .B2(\cpu.icache.r_data[6][2] ),
    .A2(net643),
    .A1(\cpu.icache.r_data[2][2] ));
 sg13g2_a22oi_1 _20566_ (.Y(_03135_),
    .B1(net583),
    .B2(\cpu.icache.r_data[3][2] ),
    .A2(net642),
    .A1(\cpu.icache.r_data[1][2] ));
 sg13g2_nand4_1 _20567_ (.B(_03133_),
    .C(_03134_),
    .A(_03132_),
    .Y(_03136_),
    .D(_03135_));
 sg13g2_nand2_1 _20568_ (.Y(_03137_),
    .A(_00162_),
    .B(net580));
 sg13g2_o21ai_1 _20569_ (.B1(_03137_),
    .Y(_03138_),
    .A1(net580),
    .A2(_03136_));
 sg13g2_nor2_1 _20570_ (.A(_00163_),
    .B(net520),
    .Y(_03139_));
 sg13g2_mux2_1 _20571_ (.A0(\cpu.icache.r_data[4][18] ),
    .A1(\cpu.icache.r_data[6][18] ),
    .S(net716),
    .X(_03140_));
 sg13g2_a22oi_1 _20572_ (.Y(_03141_),
    .B1(_03140_),
    .B2(net805),
    .A2(net806),
    .A1(\cpu.icache.r_data[5][18] ));
 sg13g2_nor2_1 _20573_ (.A(net721),
    .B(_03141_),
    .Y(_03142_));
 sg13g2_and2_1 _20574_ (.A(net821),
    .B(\cpu.icache.r_data[3][18] ),
    .X(_03143_));
 sg13g2_a21oi_1 _20575_ (.A1(net715),
    .A2(\cpu.icache.r_data[7][18] ),
    .Y(_03144_),
    .B1(_03143_));
 sg13g2_a22oi_1 _20576_ (.Y(_03145_),
    .B1(net579),
    .B2(\cpu.icache.r_data[1][18] ),
    .A2(net581),
    .A1(\cpu.icache.r_data[2][18] ));
 sg13g2_o21ai_1 _20577_ (.B1(_03145_),
    .Y(_03146_),
    .A1(_08527_),
    .A2(_03144_));
 sg13g2_nor4_1 _20578_ (.A(net1076),
    .B(_03139_),
    .C(_03142_),
    .D(_03146_),
    .Y(_03147_));
 sg13g2_a21oi_1 _20579_ (.A1(net1076),
    .A2(_03138_),
    .Y(_03148_),
    .B1(_03147_));
 sg13g2_buf_2 _20580_ (.A(_03148_),
    .X(_03149_));
 sg13g2_nor2_1 _20581_ (.A(net212),
    .B(_03149_),
    .Y(_03150_));
 sg13g2_o21ai_1 _20582_ (.B1(_03012_),
    .Y(_03151_),
    .A1(net369),
    .A2(_03032_));
 sg13g2_nor3_1 _20583_ (.A(_09006_),
    .B(_03150_),
    .C(_03151_),
    .Y(_03152_));
 sg13g2_inv_1 _20584_ (.Y(_03153_),
    .A(_03117_));
 sg13g2_buf_1 _20585_ (.A(_03153_),
    .X(_03154_));
 sg13g2_nor2_1 _20586_ (.A(_03012_),
    .B(_03154_),
    .Y(_03155_));
 sg13g2_and2_1 _20587_ (.A(_03036_),
    .B(_03155_),
    .X(_03156_));
 sg13g2_o21ai_1 _20588_ (.B1(net195),
    .Y(_03157_),
    .A1(_03152_),
    .A2(_03156_));
 sg13g2_a21oi_1 _20589_ (.A1(_03131_),
    .A2(_03157_),
    .Y(_03158_),
    .B1(net166));
 sg13g2_a21o_1 _20590_ (.A2(net148),
    .A1(_10651_),
    .B1(_03158_),
    .X(_00744_));
 sg13g2_inv_1 _20591_ (.Y(_03159_),
    .A(\cpu.dec.imm[10] ));
 sg13g2_nor2_1 _20592_ (.A(_03016_),
    .B(net231),
    .Y(_03160_));
 sg13g2_or2_1 _20593_ (.X(_03161_),
    .B(_09045_),
    .A(net225));
 sg13g2_buf_1 _20594_ (.A(_03161_),
    .X(_03162_));
 sg13g2_a21oi_1 _20595_ (.A1(_03160_),
    .A2(net211),
    .Y(_03163_),
    .B1(_03162_));
 sg13g2_buf_2 _20596_ (.A(_03163_),
    .X(_03164_));
 sg13g2_buf_1 _20597_ (.A(_03120_),
    .X(_03165_));
 sg13g2_a21oi_1 _20598_ (.A1(_08968_),
    .A2(_03057_),
    .Y(_03166_),
    .B1(_03064_));
 sg13g2_buf_2 _20599_ (.A(_03166_),
    .X(_03167_));
 sg13g2_inv_1 _20600_ (.Y(_03168_),
    .A(_03018_));
 sg13g2_nand2_1 _20601_ (.Y(_03169_),
    .A(net290),
    .B(_03168_));
 sg13g2_buf_2 _20602_ (.A(_03169_),
    .X(_03170_));
 sg13g2_nand2_1 _20603_ (.Y(_03171_),
    .A(_09893_),
    .B(_03170_));
 sg13g2_a21o_1 _20604_ (.A2(_03167_),
    .A1(net210),
    .B1(_03171_),
    .X(_03172_));
 sg13g2_nand2_1 _20605_ (.Y(_03173_),
    .A(_08971_),
    .B(_03036_));
 sg13g2_buf_1 _20606_ (.A(_03173_),
    .X(_03174_));
 sg13g2_buf_1 _20607_ (.A(_03174_),
    .X(_03175_));
 sg13g2_nor2_1 _20608_ (.A(_03041_),
    .B(_03048_),
    .Y(_03176_));
 sg13g2_buf_2 _20609_ (.A(_03176_),
    .X(_03177_));
 sg13g2_nand2b_1 _20610_ (.Y(_03178_),
    .B(_03177_),
    .A_N(_03170_));
 sg13g2_o21ai_1 _20611_ (.B1(_03178_),
    .Y(_03179_),
    .A1(net211),
    .A2(net142));
 sg13g2_o21ai_1 _20612_ (.B1(_03162_),
    .Y(_03180_),
    .A1(_03041_),
    .A2(_03048_));
 sg13g2_a22oi_1 _20613_ (.Y(_03181_),
    .B1(_03179_),
    .B2(_03180_),
    .A2(_03172_),
    .A1(_03164_));
 sg13g2_nor2_1 _20614_ (.A(_03016_),
    .B(_03015_),
    .Y(_03182_));
 sg13g2_mux2_1 _20615_ (.A0(_09008_),
    .A1(_03182_),
    .S(_03021_),
    .X(_03183_));
 sg13g2_a21oi_1 _20616_ (.A1(_03155_),
    .A2(_03183_),
    .Y(_03184_),
    .B1(_08902_));
 sg13g2_buf_2 _20617_ (.A(_03184_),
    .X(_03185_));
 sg13g2_a22oi_1 _20618_ (.Y(_00745_),
    .B1(_03181_),
    .B2(_03185_),
    .A2(net143),
    .A1(_03159_));
 sg13g2_nand2_1 _20619_ (.Y(_03186_),
    .A(_08971_),
    .B(_09003_));
 sg13g2_a21oi_1 _20620_ (.A1(net290),
    .A2(_03186_),
    .Y(_03187_),
    .B1(net293));
 sg13g2_a21oi_1 _20621_ (.A1(_09006_),
    .A2(_09139_),
    .Y(_03188_),
    .B1(net230));
 sg13g2_nor2_1 _20622_ (.A(_03187_),
    .B(_03188_),
    .Y(_03189_));
 sg13g2_nand3_1 _20623_ (.B(_03167_),
    .C(_03097_),
    .A(net292),
    .Y(_03190_));
 sg13g2_buf_2 _20624_ (.A(_03190_),
    .X(_03191_));
 sg13g2_inv_1 _20625_ (.Y(_03192_),
    .A(_03191_));
 sg13g2_a21o_1 _20626_ (.A2(_03192_),
    .A1(_03153_),
    .B1(_03174_),
    .X(_03193_));
 sg13g2_buf_1 _20627_ (.A(_03193_),
    .X(_03194_));
 sg13g2_a21oi_1 _20628_ (.A1(_08943_),
    .A2(_03191_),
    .Y(_03195_),
    .B1(_03194_));
 sg13g2_or2_1 _20629_ (.X(_03196_),
    .B(_03195_),
    .A(_03189_));
 sg13g2_o21ai_1 _20630_ (.B1(_03170_),
    .Y(_03197_),
    .A1(_08943_),
    .A2(net142));
 sg13g2_a22oi_1 _20631_ (.Y(_03198_),
    .B1(_03197_),
    .B2(_03177_),
    .A2(_03196_),
    .A1(_03164_));
 sg13g2_a22oi_1 _20632_ (.Y(_00746_),
    .B1(_03185_),
    .B2(_03198_),
    .A2(net143),
    .A1(_10382_));
 sg13g2_a21oi_1 _20633_ (.A1(_08922_),
    .A2(_03191_),
    .Y(_03199_),
    .B1(_03194_));
 sg13g2_or2_1 _20634_ (.X(_03200_),
    .B(_03199_),
    .A(_03189_));
 sg13g2_o21ai_1 _20635_ (.B1(_03170_),
    .Y(_03201_),
    .A1(_08922_),
    .A2(net142));
 sg13g2_a22oi_1 _20636_ (.Y(_03202_),
    .B1(_03201_),
    .B2(_03177_),
    .A2(_03200_),
    .A1(_03164_));
 sg13g2_a22oi_1 _20637_ (.Y(_00747_),
    .B1(_03185_),
    .B2(_03202_),
    .A2(net143),
    .A1(_10302_));
 sg13g2_a21oi_1 _20638_ (.A1(net291),
    .A2(_03191_),
    .Y(_03203_),
    .B1(_03194_));
 sg13g2_o21ai_1 _20639_ (.B1(_03164_),
    .Y(_03204_),
    .A1(_03189_),
    .A2(_03203_));
 sg13g2_nand4_1 _20640_ (.B(net290),
    .C(_09126_),
    .A(net272),
    .Y(_03205_),
    .D(_09893_));
 sg13g2_nand3_1 _20641_ (.B(_03204_),
    .C(_03205_),
    .A(_03185_),
    .Y(_03206_));
 sg13g2_o21ai_1 _20642_ (.B1(_03206_),
    .Y(_03207_),
    .A1(\cpu.dec.imm[13] ),
    .A2(net147));
 sg13g2_inv_1 _20643_ (.Y(_00748_),
    .A(_03207_));
 sg13g2_inv_1 _20644_ (.Y(_03208_),
    .A(\cpu.dec.imm[14] ));
 sg13g2_o21ai_1 _20645_ (.B1(_03170_),
    .Y(_03209_),
    .A1(_09067_),
    .A2(net142));
 sg13g2_nand2_1 _20646_ (.Y(_03210_),
    .A(_03177_),
    .B(_03209_));
 sg13g2_a21oi_1 _20647_ (.A1(_09067_),
    .A2(_03191_),
    .Y(_03211_),
    .B1(_03194_));
 sg13g2_o21ai_1 _20648_ (.B1(_03164_),
    .Y(_03212_),
    .A1(_03189_),
    .A2(_03211_));
 sg13g2_and2_1 _20649_ (.A(_03185_),
    .B(_03212_),
    .X(_03213_));
 sg13g2_a22oi_1 _20650_ (.Y(_00749_),
    .B1(_03210_),
    .B2(_03213_),
    .A2(_11943_),
    .A1(_03208_));
 sg13g2_inv_1 _20651_ (.Y(_03214_),
    .A(\cpu.dec.imm[15] ));
 sg13g2_o21ai_1 _20652_ (.B1(_03170_),
    .Y(_03215_),
    .A1(net423),
    .A2(net142));
 sg13g2_nand2_1 _20653_ (.Y(_03216_),
    .A(_03177_),
    .B(_03215_));
 sg13g2_a22oi_1 _20654_ (.Y(_00750_),
    .B1(_03213_),
    .B2(_03216_),
    .A2(net151),
    .A1(_03214_));
 sg13g2_o21ai_1 _20655_ (.B1(net231),
    .Y(_03217_),
    .A1(net214),
    .A2(_03191_));
 sg13g2_a221oi_1 _20656_ (.B2(net353),
    .C1(_03030_),
    .B1(_03217_),
    .A1(net195),
    .Y(_03218_),
    .A2(net210));
 sg13g2_nor2_1 _20657_ (.A(net126),
    .B(net194),
    .Y(_03219_));
 sg13g2_o21ai_1 _20658_ (.B1(_03219_),
    .Y(_03220_),
    .A1(net212),
    .A2(_03218_));
 sg13g2_nand2_1 _20659_ (.Y(_03221_),
    .A(net196),
    .B(_03020_));
 sg13g2_nand2_1 _20660_ (.Y(_03222_),
    .A(_03221_),
    .B(_03050_));
 sg13g2_inv_1 _20661_ (.Y(_03223_),
    .A(_00165_));
 sg13g2_mux2_1 _20662_ (.A0(\cpu.icache.r_data[4][19] ),
    .A1(\cpu.icache.r_data[6][19] ),
    .S(net710),
    .X(_03224_));
 sg13g2_a22oi_1 _20663_ (.Y(_03225_),
    .B1(_03224_),
    .B2(net805),
    .A2(net806),
    .A1(\cpu.icache.r_data[5][19] ));
 sg13g2_mux2_1 _20664_ (.A0(\cpu.icache.r_data[7][19] ),
    .A1(\cpu.icache.r_data[3][19] ),
    .S(net721),
    .X(_03226_));
 sg13g2_a22oi_1 _20665_ (.Y(_03227_),
    .B1(net820),
    .B2(_03226_),
    .A2(net579),
    .A1(\cpu.icache.r_data[1][19] ));
 sg13g2_o21ai_1 _20666_ (.B1(_03227_),
    .Y(_03228_),
    .A1(net721),
    .A2(_03225_));
 sg13g2_a221oi_1 _20667_ (.B2(\cpu.icache.r_data[2][19] ),
    .C1(_03228_),
    .B1(net581),
    .A1(_03223_),
    .Y(_03229_),
    .A2(net580));
 sg13g2_nand2_1 _20668_ (.Y(_03230_),
    .A(_00164_),
    .B(net580));
 sg13g2_mux4_1 _20669_ (.S0(_08824_),
    .A0(\cpu.icache.r_data[4][3] ),
    .A1(\cpu.icache.r_data[5][3] ),
    .A2(\cpu.icache.r_data[6][3] ),
    .A3(\cpu.icache.r_data[7][3] ),
    .S1(_08826_),
    .X(_03231_));
 sg13g2_nand2_1 _20670_ (.Y(_03232_),
    .A(net715),
    .B(_03231_));
 sg13g2_nand2_1 _20671_ (.Y(_03233_),
    .A(\cpu.icache.r_data[1][3] ),
    .B(net579));
 sg13g2_a22oi_1 _20672_ (.Y(_03234_),
    .B1(net518),
    .B2(\cpu.icache.r_data[3][3] ),
    .A2(net581),
    .A1(\cpu.icache.r_data[2][3] ));
 sg13g2_nand4_1 _20673_ (.B(_03232_),
    .C(_03233_),
    .A(net521),
    .Y(_03235_),
    .D(_03234_));
 sg13g2_a21oi_1 _20674_ (.A1(_03230_),
    .A2(_03235_),
    .Y(_03236_),
    .B1(net929));
 sg13g2_a21oi_1 _20675_ (.A1(_09009_),
    .A2(_03229_),
    .Y(_03237_),
    .B1(_03236_));
 sg13g2_buf_1 _20676_ (.A(_03237_),
    .X(_03238_));
 sg13g2_inv_1 _20677_ (.Y(_03239_),
    .A(net229));
 sg13g2_nor2_1 _20678_ (.A(_03023_),
    .B(_03239_),
    .Y(_03240_));
 sg13g2_a22oi_1 _20679_ (.Y(_03241_),
    .B1(_03222_),
    .B2(_03240_),
    .A2(_03220_),
    .A1(_08921_));
 sg13g2_nand2_1 _20680_ (.Y(_03242_),
    .A(_10645_),
    .B(net164));
 sg13g2_o21ai_1 _20681_ (.B1(_03242_),
    .Y(_00751_),
    .A1(net151),
    .A2(_03241_));
 sg13g2_inv_1 _20682_ (.Y(_03243_),
    .A(net292));
 sg13g2_o21ai_1 _20683_ (.B1(net214),
    .Y(_03244_),
    .A1(net287),
    .A2(net225));
 sg13g2_buf_1 _20684_ (.A(net293),
    .X(_03245_));
 sg13g2_a22oi_1 _20685_ (.Y(_03246_),
    .B1(_03244_),
    .B2(net228),
    .A2(net210),
    .A1(net170));
 sg13g2_nand2b_1 _20686_ (.Y(_03247_),
    .B(_09027_),
    .A_N(_09045_));
 sg13g2_buf_1 _20687_ (.A(_03247_),
    .X(_03248_));
 sg13g2_o21ai_1 _20688_ (.B1(net162),
    .Y(_03249_),
    .A1(net212),
    .A2(_03246_));
 sg13g2_nand2_1 _20689_ (.Y(_03250_),
    .A(_03243_),
    .B(_03249_));
 sg13g2_nand2_1 _20690_ (.Y(_03251_),
    .A(_03117_),
    .B(_03222_));
 sg13g2_nor2_1 _20691_ (.A(net142),
    .B(_03191_),
    .Y(_03252_));
 sg13g2_nand4_1 _20692_ (.B(net171),
    .C(_09893_),
    .A(net369),
    .Y(_03253_),
    .D(_03252_));
 sg13g2_nand2_2 _20693_ (.Y(_03254_),
    .A(_03032_),
    .B(_03120_));
 sg13g2_nor2_1 _20694_ (.A(_09003_),
    .B(_03238_),
    .Y(_03255_));
 sg13g2_a21oi_1 _20695_ (.A1(_08943_),
    .A2(net353),
    .Y(_03256_),
    .B1(_03255_));
 sg13g2_nand2_1 _20696_ (.Y(_03257_),
    .A(_03254_),
    .B(_03256_));
 sg13g2_o21ai_1 _20697_ (.B1(_03257_),
    .Y(_03258_),
    .A1(net292),
    .A2(_03254_));
 sg13g2_nor4_1 _20698_ (.A(net213),
    .B(_09006_),
    .C(net194),
    .D(_03239_),
    .Y(_03259_));
 sg13g2_a21oi_1 _20699_ (.A1(net145),
    .A2(_03258_),
    .Y(_03260_),
    .B1(_03259_));
 sg13g2_nand4_1 _20700_ (.B(_03251_),
    .C(_03253_),
    .A(_03250_),
    .Y(_03261_),
    .D(_03260_));
 sg13g2_mux2_1 _20701_ (.A0(_10583_),
    .A1(_03261_),
    .S(net146),
    .X(_00752_));
 sg13g2_nor2_1 _20702_ (.A(net292),
    .B(_03018_),
    .Y(_03262_));
 sg13g2_a21oi_1 _20703_ (.A1(_09008_),
    .A2(_03117_),
    .Y(_03263_),
    .B1(_03262_));
 sg13g2_inv_1 _20704_ (.Y(_03264_),
    .A(_03263_));
 sg13g2_a221oi_1 _20705_ (.B2(net423),
    .C1(_03264_),
    .B1(_03252_),
    .A1(_08942_),
    .Y(_03265_),
    .A2(net210));
 sg13g2_nor3_1 _20706_ (.A(_03162_),
    .B(_03160_),
    .C(_03265_),
    .Y(_03266_));
 sg13g2_nand2_1 _20707_ (.Y(_03267_),
    .A(net369),
    .B(_03048_));
 sg13g2_a21oi_1 _20708_ (.A1(_03263_),
    .A2(_03267_),
    .Y(_03268_),
    .B1(_03041_));
 sg13g2_nor3_1 _20709_ (.A(_09898_),
    .B(net211),
    .C(_03182_),
    .Y(_03269_));
 sg13g2_nor3_1 _20710_ (.A(_03266_),
    .B(_03268_),
    .C(_03269_),
    .Y(_03270_));
 sg13g2_a21oi_1 _20711_ (.A1(net287),
    .A2(_03254_),
    .Y(_03271_),
    .B1(net163));
 sg13g2_o21ai_1 _20712_ (.B1(net423),
    .Y(_03272_),
    .A1(_03249_),
    .A2(_03271_));
 sg13g2_a21oi_1 _20713_ (.A1(_03270_),
    .A2(_03272_),
    .Y(_03273_),
    .B1(net172));
 sg13g2_a21o_1 _20714_ (.A2(net148),
    .A1(_10613_),
    .B1(_03273_),
    .X(_00753_));
 sg13g2_a21oi_1 _20715_ (.A1(net353),
    .A2(_03192_),
    .Y(_03274_),
    .B1(net228));
 sg13g2_nor3_1 _20716_ (.A(net212),
    .B(net214),
    .C(_03274_),
    .Y(_03275_));
 sg13g2_nor3_1 _20717_ (.A(net126),
    .B(net194),
    .C(_03275_),
    .Y(_03276_));
 sg13g2_nand3_1 _20718_ (.B(net423),
    .C(_03020_),
    .A(net196),
    .Y(_03277_));
 sg13g2_o21ai_1 _20719_ (.B1(_03277_),
    .Y(_03278_),
    .A1(net291),
    .A2(_03276_));
 sg13g2_nand2_1 _20720_ (.Y(_03279_),
    .A(net147),
    .B(_03278_));
 sg13g2_o21ai_1 _20721_ (.B1(_03279_),
    .Y(_00754_),
    .A1(_10791_),
    .A2(net150));
 sg13g2_o21ai_1 _20722_ (.B1(_03149_),
    .Y(_03280_),
    .A1(_09140_),
    .A2(_03248_));
 sg13g2_or4_1 _20723_ (.A(_08943_),
    .B(net149),
    .C(net162),
    .D(_03036_),
    .X(_03281_));
 sg13g2_o21ai_1 _20724_ (.B1(_09046_),
    .Y(_03282_),
    .A1(_03174_),
    .A2(_03192_));
 sg13g2_nor2_1 _20725_ (.A(_03014_),
    .B(_09003_),
    .Y(_03283_));
 sg13g2_buf_2 _20726_ (.A(_03283_),
    .X(_03284_));
 sg13g2_nand2_1 _20727_ (.Y(_03285_),
    .A(_03016_),
    .B(_03284_));
 sg13g2_buf_2 _20728_ (.A(_03285_),
    .X(_03286_));
 sg13g2_nand2_1 _20729_ (.Y(_03287_),
    .A(_03286_),
    .B(_03042_));
 sg13g2_a21oi_1 _20730_ (.A1(_03028_),
    .A2(_03287_),
    .Y(_03288_),
    .B1(net194));
 sg13g2_a221oi_1 _20731_ (.B2(_03288_),
    .C1(_08905_),
    .B1(_03282_),
    .A1(_03280_),
    .Y(_03289_),
    .A2(_03281_));
 sg13g2_a21o_1 _20732_ (.A2(net148),
    .A1(\cpu.dec.imm[5] ),
    .B1(_03289_),
    .X(_00755_));
 sg13g2_buf_1 _20733_ (.A(_03096_),
    .X(_03290_));
 sg13g2_inv_1 _20734_ (.Y(_03291_),
    .A(net352));
 sg13g2_o21ai_1 _20735_ (.B1(_03238_),
    .Y(_03292_),
    .A1(_03160_),
    .A2(_03252_));
 sg13g2_o21ai_1 _20736_ (.B1(_03292_),
    .Y(_03293_),
    .A1(_03015_),
    .A2(_03291_));
 sg13g2_nand2_1 _20737_ (.Y(_03294_),
    .A(net369),
    .B(net196));
 sg13g2_o21ai_1 _20738_ (.B1(net162),
    .Y(_03295_),
    .A1(net165),
    .A2(_03294_));
 sg13g2_a221oi_1 _20739_ (.B2(net171),
    .C1(_03295_),
    .B1(_03293_),
    .A1(net229),
    .Y(_03296_),
    .A2(_03271_));
 sg13g2_nor2_1 _20740_ (.A(net353),
    .B(net126),
    .Y(_03297_));
 sg13g2_a221oi_1 _20741_ (.B2(net352),
    .C1(net162),
    .B1(_03297_),
    .A1(net126),
    .Y(_03298_),
    .A2(net229));
 sg13g2_nor3_1 _20742_ (.A(net172),
    .B(_03296_),
    .C(_03298_),
    .Y(_03299_));
 sg13g2_a21o_1 _20743_ (.A2(net148),
    .A1(\cpu.dec.imm[6] ),
    .B1(_03299_),
    .X(_00756_));
 sg13g2_o21ai_1 _20744_ (.B1(_03125_),
    .Y(_03300_),
    .A1(_03123_),
    .A2(_03015_));
 sg13g2_nand3_1 _20745_ (.B(net171),
    .C(_03192_),
    .A(net230),
    .Y(_03301_));
 sg13g2_o21ai_1 _20746_ (.B1(_03301_),
    .Y(_03302_),
    .A1(net231),
    .A2(net163));
 sg13g2_a22oi_1 _20747_ (.Y(_03303_),
    .B1(_03302_),
    .B2(net272),
    .A2(_03300_),
    .A1(_03033_));
 sg13g2_and2_1 _20748_ (.A(net196),
    .B(_03020_),
    .X(_03304_));
 sg13g2_nand2_1 _20749_ (.Y(_03305_),
    .A(net287),
    .B(_03286_));
 sg13g2_nand2_1 _20750_ (.Y(_03306_),
    .A(net149),
    .B(_03117_));
 sg13g2_o21ai_1 _20751_ (.B1(_03306_),
    .Y(_03307_),
    .A1(_03066_),
    .A2(_03305_));
 sg13g2_a22oi_1 _20752_ (.Y(_03308_),
    .B1(_03023_),
    .B2(_03307_),
    .A2(_03304_),
    .A1(_08921_));
 sg13g2_o21ai_1 _20753_ (.B1(_03308_),
    .Y(_03309_),
    .A1(net211),
    .A2(_03303_));
 sg13g2_nand2_1 _20754_ (.Y(_03310_),
    .A(net147),
    .B(_03309_));
 sg13g2_o21ai_1 _20755_ (.B1(_03310_),
    .Y(_00757_),
    .A1(_10734_),
    .A2(net150));
 sg13g2_inv_1 _20756_ (.Y(_03311_),
    .A(\cpu.dec.imm[8] ));
 sg13g2_inv_2 _20757_ (.Y(_03312_),
    .A(_03149_));
 sg13g2_o21ai_1 _20758_ (.B1(_03170_),
    .Y(_03313_),
    .A1(_03312_),
    .A2(_03175_));
 sg13g2_nor2_1 _20759_ (.A(_03149_),
    .B(_03192_),
    .Y(_03314_));
 sg13g2_a21oi_1 _20760_ (.A1(net210),
    .A2(_03082_),
    .Y(_03315_),
    .B1(_03171_));
 sg13g2_o21ai_1 _20761_ (.B1(_03315_),
    .Y(_03316_),
    .A1(_03194_),
    .A2(_03314_));
 sg13g2_inv_1 _20762_ (.Y(_03317_),
    .A(_03082_));
 sg13g2_nor2_1 _20763_ (.A(net162),
    .B(_03317_),
    .Y(_03318_));
 sg13g2_nor2b_1 _20764_ (.A(_03305_),
    .B_N(_03318_),
    .Y(_03319_));
 sg13g2_a221oi_1 _20765_ (.B2(_03164_),
    .C1(_03319_),
    .B1(_03316_),
    .A1(_03177_),
    .Y(_03320_),
    .A2(_03313_));
 sg13g2_a22oi_1 _20766_ (.Y(_00758_),
    .B1(_03185_),
    .B2(_03320_),
    .A2(net151),
    .A1(_03311_));
 sg13g2_inv_1 _20767_ (.Y(_03321_),
    .A(\cpu.dec.imm[9] ));
 sg13g2_nor2_1 _20768_ (.A(_03192_),
    .B(net229),
    .Y(_03322_));
 sg13g2_a21oi_1 _20769_ (.A1(_03243_),
    .A2(net210),
    .Y(_03323_),
    .B1(_03171_));
 sg13g2_o21ai_1 _20770_ (.B1(_03323_),
    .Y(_03324_),
    .A1(_03194_),
    .A2(_03322_));
 sg13g2_o21ai_1 _20771_ (.B1(_03170_),
    .Y(_03325_),
    .A1(_03175_),
    .A2(_03239_));
 sg13g2_a22oi_1 _20772_ (.Y(_03326_),
    .B1(_03325_),
    .B2(_03177_),
    .A2(_03324_),
    .A1(_03164_));
 sg13g2_a22oi_1 _20773_ (.Y(_00759_),
    .B1(_03185_),
    .B2(_03326_),
    .A2(net151),
    .A1(_03321_));
 sg13g2_nor4_1 _20774_ (.A(_08488_),
    .B(_08922_),
    .C(_03050_),
    .D(_03101_),
    .Y(_03327_));
 sg13g2_buf_1 _20775_ (.A(\cpu.dec.do_inv_mmu ),
    .X(_03328_));
 sg13g2_mux2_1 _20776_ (.A0(_03327_),
    .A1(_03328_),
    .S(_03045_),
    .X(_00760_));
 sg13g2_nand2_1 _20777_ (.Y(_03329_),
    .A(net213),
    .B(net170));
 sg13g2_nor4_1 _20778_ (.A(net173),
    .B(_03284_),
    .C(_03036_),
    .D(_03329_),
    .Y(_03330_));
 sg13g2_a21o_1 _20779_ (.A2(net148),
    .A1(\cpu.dec.io ),
    .B1(_03330_),
    .X(_00761_));
 sg13g2_or4_1 _20780_ (.A(_08945_),
    .B(_03117_),
    .C(_03149_),
    .D(_03237_),
    .X(_03331_));
 sg13g2_buf_2 _20781_ (.A(_03331_),
    .X(_03332_));
 sg13g2_nor4_1 _20782_ (.A(net173),
    .B(_03286_),
    .C(net163),
    .D(_03332_),
    .Y(_03333_));
 sg13g2_a21o_1 _20783_ (.A2(net164),
    .A1(\cpu.dec.jmp ),
    .B1(_03333_),
    .X(_00762_));
 sg13g2_a21oi_1 _20784_ (.A1(net228),
    .A2(net195),
    .Y(_03334_),
    .B1(net194));
 sg13g2_nor3_1 _20785_ (.A(net172),
    .B(_03186_),
    .C(_03334_),
    .Y(_03335_));
 sg13g2_a21o_1 _20786_ (.A2(net164),
    .A1(_11465_),
    .B1(_03335_),
    .X(_00763_));
 sg13g2_nor4_1 _20787_ (.A(net173),
    .B(_08945_),
    .C(net290),
    .D(_09128_),
    .Y(_03336_));
 sg13g2_a21o_1 _20788_ (.A2(net164),
    .A1(_09333_),
    .B1(_03336_),
    .X(_00764_));
 sg13g2_o21ai_1 _20789_ (.B1(_09150_),
    .Y(_03337_),
    .A1(_09066_),
    .A2(net290));
 sg13g2_nand3_1 _20790_ (.B(_03127_),
    .C(net291),
    .A(net213),
    .Y(_03338_));
 sg13g2_nand3b_1 _20791_ (.B(_03013_),
    .C(_03119_),
    .Y(_03339_),
    .A_N(_09085_));
 sg13g2_nand4_1 _20792_ (.B(_03028_),
    .C(_03338_),
    .A(_03284_),
    .Y(_03340_),
    .D(_03339_));
 sg13g2_o21ai_1 _20793_ (.B1(_03340_),
    .Y(_03341_),
    .A1(_09131_),
    .A2(_03337_));
 sg13g2_nor2_1 _20794_ (.A(net166),
    .B(_03341_),
    .Y(_03342_));
 sg13g2_a21oi_1 _20795_ (.A1(_10301_),
    .A2(_11943_),
    .Y(_00765_),
    .B1(_03342_));
 sg13g2_inv_1 _20796_ (.Y(_03343_),
    .A(\cpu.dec.r_rd[0] ));
 sg13g2_nor3_1 _20797_ (.A(net230),
    .B(_09121_),
    .C(_03332_),
    .Y(_03344_));
 sg13g2_a21oi_1 _20798_ (.A1(_03290_),
    .A2(_03332_),
    .Y(_03345_),
    .B1(_03344_));
 sg13g2_nor2_1 _20799_ (.A(_09006_),
    .B(_03345_),
    .Y(_03346_));
 sg13g2_a21oi_1 _20800_ (.A1(net213),
    .A2(net352),
    .Y(_03347_),
    .B1(_03346_));
 sg13g2_o21ai_1 _20801_ (.B1(net194),
    .Y(_03348_),
    .A1(_03165_),
    .A2(_03150_));
 sg13g2_inv_1 _20802_ (.Y(_03349_),
    .A(_03121_));
 sg13g2_nor3_1 _20803_ (.A(net225),
    .B(_03165_),
    .C(net352),
    .Y(_03350_));
 sg13g2_nor4_1 _20804_ (.A(net214),
    .B(_03168_),
    .C(_03349_),
    .D(_03350_),
    .Y(_03351_));
 sg13g2_nor2_2 _20805_ (.A(net212),
    .B(net287),
    .Y(_03352_));
 sg13g2_nor2_1 _20806_ (.A(net293),
    .B(net352),
    .Y(_03353_));
 sg13g2_a21oi_1 _20807_ (.A1(net293),
    .A2(_03312_),
    .Y(_03354_),
    .B1(_03353_));
 sg13g2_a22oi_1 _20808_ (.Y(_03355_),
    .B1(_03352_),
    .B2(_03354_),
    .A2(net352),
    .A1(net149));
 sg13g2_inv_1 _20809_ (.Y(_03356_),
    .A(_03355_));
 sg13g2_a22oi_1 _20810_ (.Y(_03357_),
    .B1(_03356_),
    .B2(net170),
    .A2(_03351_),
    .A1(_03348_));
 sg13g2_o21ai_1 _20811_ (.B1(_03357_),
    .Y(_03358_),
    .A1(net163),
    .A2(_03347_));
 sg13g2_nand2_1 _20812_ (.Y(_03359_),
    .A(net147),
    .B(_03358_));
 sg13g2_o21ai_1 _20813_ (.B1(_03359_),
    .Y(_00766_),
    .A1(_03343_),
    .A2(net150));
 sg13g2_a21o_1 _20814_ (.A2(_03332_),
    .A1(_09896_),
    .B1(net171),
    .X(_03360_));
 sg13g2_o21ai_1 _20815_ (.B1(_03123_),
    .Y(_03361_),
    .A1(net287),
    .A2(_03162_));
 sg13g2_a22oi_1 _20816_ (.Y(_03362_),
    .B1(_03361_),
    .B2(_03033_),
    .A2(_03360_),
    .A1(_03284_));
 sg13g2_nor3_1 _20817_ (.A(net212),
    .B(net210),
    .C(net162),
    .Y(_03363_));
 sg13g2_a21oi_1 _20818_ (.A1(net353),
    .A2(_03239_),
    .Y(_03364_),
    .B1(net212));
 sg13g2_nor2_1 _20819_ (.A(net353),
    .B(_03066_),
    .Y(_03365_));
 sg13g2_o21ai_1 _20820_ (.B1(net228),
    .Y(_03366_),
    .A1(_03364_),
    .A2(_03365_));
 sg13g2_nand3_1 _20821_ (.B(_03167_),
    .C(_03352_),
    .A(net231),
    .Y(_03367_));
 sg13g2_nor3_1 _20822_ (.A(_08945_),
    .B(_03101_),
    .C(_03153_),
    .Y(_03368_));
 sg13g2_nand3_1 _20823_ (.B(net229),
    .C(_03368_),
    .A(_03312_),
    .Y(_03369_));
 sg13g2_buf_1 _20824_ (.A(_03369_),
    .X(_03370_));
 sg13g2_a221oi_1 _20825_ (.B2(_03048_),
    .C1(_03041_),
    .B1(_03370_),
    .A1(_03366_),
    .Y(_03371_),
    .A2(_03367_));
 sg13g2_a21oi_1 _20826_ (.A1(net229),
    .A2(_03363_),
    .Y(_03372_),
    .B1(_03371_));
 sg13g2_o21ai_1 _20827_ (.B1(_03372_),
    .Y(_03373_),
    .A1(_03066_),
    .A2(_03362_));
 sg13g2_mux2_1 _20828_ (.A0(\cpu.dec.r_rd[1] ),
    .A1(_03373_),
    .S(net146),
    .X(_00767_));
 sg13g2_inv_1 _20829_ (.Y(_03374_),
    .A(\cpu.dec.r_rd[2] ));
 sg13g2_nor2_1 _20830_ (.A(_03317_),
    .B(_03362_),
    .Y(_03375_));
 sg13g2_nor2_1 _20831_ (.A(_03245_),
    .B(_03082_),
    .Y(_03376_));
 sg13g2_a21oi_1 _20832_ (.A1(_03245_),
    .A2(net211),
    .Y(_03377_),
    .B1(_03376_));
 sg13g2_a22oi_1 _20833_ (.Y(_03378_),
    .B1(_03352_),
    .B2(_03377_),
    .A2(_03082_),
    .A1(net126));
 sg13g2_nand2_1 _20834_ (.Y(_03379_),
    .A(_03117_),
    .B(_03363_));
 sg13g2_o21ai_1 _20835_ (.B1(_03379_),
    .Y(_03380_),
    .A1(_03041_),
    .A2(_03378_));
 sg13g2_o21ai_1 _20836_ (.B1(_09138_),
    .Y(_03381_),
    .A1(_03375_),
    .A2(_03380_));
 sg13g2_o21ai_1 _20837_ (.B1(_03381_),
    .Y(_00768_),
    .A1(_03374_),
    .A2(net150));
 sg13g2_o21ai_1 _20838_ (.B1(net212),
    .Y(_03382_),
    .A1(net353),
    .A2(net194));
 sg13g2_nor3_1 _20839_ (.A(net228),
    .B(net225),
    .C(_03243_),
    .Y(_03383_));
 sg13g2_a21oi_1 _20840_ (.A1(net272),
    .A2(net145),
    .Y(_03384_),
    .B1(_03383_));
 sg13g2_nand2_1 _20841_ (.Y(_03385_),
    .A(_03382_),
    .B(_03384_));
 sg13g2_a21oi_1 _20842_ (.A1(net228),
    .A2(_03329_),
    .Y(_03386_),
    .B1(net272));
 sg13g2_a21o_1 _20843_ (.A2(_03332_),
    .A1(net149),
    .B1(_03352_),
    .X(_03387_));
 sg13g2_nand3_1 _20844_ (.B(net145),
    .C(_03387_),
    .A(_03243_),
    .Y(_03388_));
 sg13g2_o21ai_1 _20845_ (.B1(_03388_),
    .Y(_03389_),
    .A1(_03385_),
    .A2(_03386_));
 sg13g2_mux2_1 _20846_ (.A0(\cpu.dec.r_rd[3] ),
    .A1(_03389_),
    .S(_09148_),
    .X(_00769_));
 sg13g2_o21ai_1 _20847_ (.B1(_03286_),
    .Y(_03390_),
    .A1(net287),
    .A2(_03291_));
 sg13g2_nand2_1 _20848_ (.Y(_03391_),
    .A(_09126_),
    .B(net142));
 sg13g2_nand2_1 _20849_ (.Y(_03392_),
    .A(_09006_),
    .B(_03042_));
 sg13g2_nand2_1 _20850_ (.Y(_03393_),
    .A(_09121_),
    .B(_03332_));
 sg13g2_nand2_1 _20851_ (.Y(_03394_),
    .A(_09008_),
    .B(_03393_));
 sg13g2_nand2_1 _20852_ (.Y(_03395_),
    .A(_03305_),
    .B(_03394_));
 sg13g2_a22oi_1 _20853_ (.Y(_03396_),
    .B1(_03395_),
    .B2(_09897_),
    .A2(_03392_),
    .A1(net171));
 sg13g2_o21ai_1 _20854_ (.B1(_03396_),
    .Y(_03397_),
    .A1(_03048_),
    .A2(_03391_));
 sg13g2_a221oi_1 _20855_ (.B2(net352),
    .C1(_03024_),
    .B1(_03397_),
    .A1(_03023_),
    .Y(_03398_),
    .A2(_03390_));
 sg13g2_a21oi_1 _20856_ (.A1(net764),
    .A2(net143),
    .Y(_00770_),
    .B1(_03398_));
 sg13g2_nand3_1 _20857_ (.B(_09125_),
    .C(net142),
    .A(net230),
    .Y(_03399_));
 sg13g2_o21ai_1 _20858_ (.B1(_03399_),
    .Y(_03400_),
    .A1(_03066_),
    .A2(_03282_));
 sg13g2_nand2_1 _20859_ (.Y(_03401_),
    .A(_03026_),
    .B(_09893_));
 sg13g2_o21ai_1 _20860_ (.B1(_03391_),
    .Y(_03402_),
    .A1(_03401_),
    .A2(_03282_));
 sg13g2_o21ai_1 _20861_ (.B1(_03167_),
    .Y(_03403_),
    .A1(_03286_),
    .A2(_03393_));
 sg13g2_a21oi_1 _20862_ (.A1(net287),
    .A2(_03403_),
    .Y(_03404_),
    .B1(_03013_));
 sg13g2_a221oi_1 _20863_ (.B2(_03167_),
    .C1(_03404_),
    .B1(_03402_),
    .A1(_03284_),
    .Y(_03405_),
    .A2(_03400_));
 sg13g2_nand2_1 _20864_ (.Y(_03406_),
    .A(_03026_),
    .B(_03066_));
 sg13g2_a21oi_1 _20865_ (.A1(_03286_),
    .A2(_03406_),
    .Y(_03407_),
    .B1(net162));
 sg13g2_a21oi_1 _20866_ (.A1(net162),
    .A2(_03405_),
    .Y(_03408_),
    .B1(_03407_));
 sg13g2_nand2_1 _20867_ (.Y(_03409_),
    .A(net147),
    .B(_03408_));
 sg13g2_o21ai_1 _20868_ (.B1(_03409_),
    .Y(_00771_),
    .A1(net895),
    .A2(net150));
 sg13g2_nand2_1 _20869_ (.Y(_03410_),
    .A(_03396_),
    .B(_03391_));
 sg13g2_a21oi_1 _20870_ (.A1(_03050_),
    .A2(_03317_),
    .Y(_03411_),
    .B1(_03023_));
 sg13g2_a221oi_1 _20871_ (.B2(_03411_),
    .C1(_03024_),
    .B1(_03410_),
    .A1(_03027_),
    .Y(_03412_),
    .A2(_03318_));
 sg13g2_a21oi_1 _20872_ (.A1(net896),
    .A2(net143),
    .Y(_00772_),
    .B1(_03412_));
 sg13g2_nor2_1 _20873_ (.A(net292),
    .B(_03394_),
    .Y(_03413_));
 sg13g2_nor2_1 _20874_ (.A(net163),
    .B(_03413_),
    .Y(_03414_));
 sg13g2_a21oi_1 _20875_ (.A1(net213),
    .A2(_03334_),
    .Y(_03415_),
    .B1(_03414_));
 sg13g2_nand2_1 _20876_ (.Y(_03416_),
    .A(net228),
    .B(net170));
 sg13g2_o21ai_1 _20877_ (.B1(_03416_),
    .Y(_03417_),
    .A1(net228),
    .A2(net196));
 sg13g2_o21ai_1 _20878_ (.B1(net195),
    .Y(_03418_),
    .A1(net213),
    .A2(_03413_));
 sg13g2_a21oi_1 _20879_ (.A1(net231),
    .A2(net195),
    .Y(_03419_),
    .B1(_03128_));
 sg13g2_a221oi_1 _20880_ (.B2(_03419_),
    .C1(net272),
    .B1(_03418_),
    .A1(net213),
    .Y(_03420_),
    .A2(_03417_));
 sg13g2_a21oi_1 _20881_ (.A1(net272),
    .A2(_03415_),
    .Y(_03421_),
    .B1(_03420_));
 sg13g2_nand2_1 _20882_ (.Y(_03422_),
    .A(_11098_),
    .B(net164));
 sg13g2_o21ai_1 _20883_ (.B1(_03422_),
    .Y(_00773_),
    .A1(net151),
    .A2(_03421_));
 sg13g2_nor2_1 _20884_ (.A(net165),
    .B(net352),
    .Y(_03423_));
 sg13g2_a21oi_1 _20885_ (.A1(net165),
    .A2(_03312_),
    .Y(_03424_),
    .B1(_03423_));
 sg13g2_nand3_1 _20886_ (.B(_09085_),
    .C(net290),
    .A(_08921_),
    .Y(_03425_));
 sg13g2_nand2_1 _20887_ (.Y(_03426_),
    .A(net214),
    .B(_03254_));
 sg13g2_a21oi_2 _20888_ (.B1(_03426_),
    .Y(_03427_),
    .A2(_03425_),
    .A1(net149));
 sg13g2_nor3_1 _20889_ (.A(net145),
    .B(_03312_),
    .C(_03427_),
    .Y(_03428_));
 sg13g2_a21oi_1 _20890_ (.A1(net145),
    .A2(_03424_),
    .Y(_03429_),
    .B1(_03428_));
 sg13g2_nand2_1 _20891_ (.Y(_03430_),
    .A(_10281_),
    .B(net166));
 sg13g2_o21ai_1 _20892_ (.B1(_03430_),
    .Y(_00774_),
    .A1(net151),
    .A2(_03429_));
 sg13g2_nor2_1 _20893_ (.A(net165),
    .B(_03167_),
    .Y(_03431_));
 sg13g2_a21oi_1 _20894_ (.A1(net165),
    .A2(_03239_),
    .Y(_03432_),
    .B1(_03431_));
 sg13g2_o21ai_1 _20895_ (.B1(net163),
    .Y(_03433_),
    .A1(_03239_),
    .A2(_03427_));
 sg13g2_o21ai_1 _20896_ (.B1(_03433_),
    .Y(_03434_),
    .A1(net163),
    .A2(_03432_));
 sg13g2_nand2_1 _20897_ (.Y(_03435_),
    .A(net681),
    .B(net166));
 sg13g2_o21ai_1 _20898_ (.B1(_03435_),
    .Y(_00775_),
    .A1(net151),
    .A2(_03434_));
 sg13g2_nand2_1 _20899_ (.Y(_03436_),
    .A(net165),
    .B(net211));
 sg13g2_o21ai_1 _20900_ (.B1(_03436_),
    .Y(_03437_),
    .A1(net165),
    .A2(_03082_));
 sg13g2_nor2_1 _20901_ (.A(_03124_),
    .B(_03437_),
    .Y(_03438_));
 sg13g2_nor3_1 _20902_ (.A(net145),
    .B(net211),
    .C(_03427_),
    .Y(_03439_));
 sg13g2_o21ai_1 _20903_ (.B1(net147),
    .Y(_03440_),
    .A1(_03438_),
    .A2(_03439_));
 sg13g2_o21ai_1 _20904_ (.B1(_03440_),
    .Y(_00776_),
    .A1(net772),
    .A2(net146));
 sg13g2_nand2_1 _20905_ (.Y(_03441_),
    .A(_03124_),
    .B(_03427_));
 sg13g2_a21oi_1 _20906_ (.A1(net369),
    .A2(_09140_),
    .Y(_03442_),
    .B1(_03262_));
 sg13g2_nand3_1 _20907_ (.B(_03287_),
    .C(_03442_),
    .A(_09897_),
    .Y(_03443_));
 sg13g2_nand3_1 _20908_ (.B(_03441_),
    .C(_03443_),
    .A(net147),
    .Y(_03444_));
 sg13g2_o21ai_1 _20909_ (.B1(_03444_),
    .Y(_00777_),
    .A1(net683),
    .A2(net146));
 sg13g2_or4_1 _20910_ (.A(_08902_),
    .B(net291),
    .C(_09128_),
    .D(_09143_),
    .X(_03445_));
 sg13g2_o21ai_1 _20911_ (.B1(_03445_),
    .Y(_00778_),
    .A1(net770),
    .A2(_09148_));
 sg13g2_nor4_1 _20912_ (.A(net173),
    .B(_08921_),
    .C(_09086_),
    .D(net291),
    .Y(_03446_));
 sg13g2_a21o_1 _20913_ (.A2(net164),
    .A1(\cpu.dec.r_set_cc ),
    .B1(_03446_),
    .X(_00779_));
 sg13g2_a22oi_1 _20914_ (.Y(_03447_),
    .B1(net210),
    .B2(net170),
    .A2(_03168_),
    .A1(_03127_));
 sg13g2_buf_1 _20915_ (.A(\cpu.dec.r_store ),
    .X(_03448_));
 sg13g2_nand2_1 _20916_ (.Y(_03449_),
    .A(_03448_),
    .B(net166));
 sg13g2_o21ai_1 _20917_ (.B1(_03449_),
    .Y(_00780_),
    .A1(net151),
    .A2(_03447_));
 sg13g2_nor3_1 _20918_ (.A(net172),
    .B(_03050_),
    .C(_03370_),
    .Y(_03450_));
 sg13g2_a21o_1 _20919_ (.A2(net164),
    .A1(\cpu.dec.r_swapsp ),
    .B1(_03450_),
    .X(_00781_));
 sg13g2_nor3_1 _20920_ (.A(_03050_),
    .B(_03312_),
    .C(net229),
    .Y(_03451_));
 sg13g2_and2_1 _20921_ (.A(_03368_),
    .B(_03451_),
    .X(_03452_));
 sg13g2_mux2_1 _20922_ (.A0(\cpu.dec.r_sys_call ),
    .A1(_03452_),
    .S(net146),
    .X(_00782_));
 sg13g2_a21o_1 _20923_ (.A2(_03394_),
    .A1(_09894_),
    .B1(_03243_),
    .X(_03453_));
 sg13g2_nand2_1 _20924_ (.Y(_03454_),
    .A(_03167_),
    .B(_03290_));
 sg13g2_xnor2_1 _20925_ (.Y(_03455_),
    .A(_03082_),
    .B(_03454_));
 sg13g2_nand2_1 _20926_ (.Y(_03456_),
    .A(_08488_),
    .B(_03455_));
 sg13g2_a21oi_1 _20927_ (.A1(_03254_),
    .A2(_03453_),
    .Y(_03457_),
    .B1(_03456_));
 sg13g2_nand2_1 _20928_ (.Y(_03458_),
    .A(_08971_),
    .B(_03284_));
 sg13g2_a21oi_1 _20929_ (.A1(_09121_),
    .A2(_03312_),
    .Y(_03459_),
    .B1(_03458_));
 sg13g2_o21ai_1 _20930_ (.B1(_03459_),
    .Y(_03460_),
    .A1(_08945_),
    .A2(_09122_));
 sg13g2_nand3_1 _20931_ (.B(_03121_),
    .C(_03460_),
    .A(net145),
    .Y(_03461_));
 sg13g2_nand2_1 _20932_ (.Y(_03462_),
    .A(_03149_),
    .B(net229));
 sg13g2_xnor2_1 _20933_ (.Y(_03463_),
    .A(net211),
    .B(_03462_));
 sg13g2_buf_1 _20934_ (.A(net1146),
    .X(_03464_));
 sg13g2_nor2_1 _20935_ (.A(_03464_),
    .B(_09121_),
    .Y(_03465_));
 sg13g2_a21oi_1 _20936_ (.A1(_08348_),
    .A2(net291),
    .Y(_03466_),
    .B1(_03465_));
 sg13g2_nor4_1 _20937_ (.A(net369),
    .B(_03286_),
    .C(_03463_),
    .D(_03466_),
    .Y(_03467_));
 sg13g2_nor3_1 _20938_ (.A(_03457_),
    .B(_03461_),
    .C(_03467_),
    .Y(_03468_));
 sg13g2_o21ai_1 _20939_ (.B1(_09123_),
    .Y(_03469_),
    .A1(_08942_),
    .A2(_03098_));
 sg13g2_nand3_1 _20940_ (.B(_03023_),
    .C(_03469_),
    .A(_03015_),
    .Y(_03470_));
 sg13g2_nor4_1 _20941_ (.A(_09880_),
    .B(_03458_),
    .C(_03098_),
    .D(_03332_),
    .Y(_03471_));
 sg13g2_nor2_1 _20942_ (.A(_03470_),
    .B(_03471_),
    .Y(_03472_));
 sg13g2_a22oi_1 _20943_ (.Y(_03473_),
    .B1(_09150_),
    .B2(_08921_),
    .A2(_09067_),
    .A1(_08942_));
 sg13g2_nand3_1 _20944_ (.B(_09121_),
    .C(_03149_),
    .A(_09067_),
    .Y(_03474_));
 sg13g2_o21ai_1 _20945_ (.B1(_03474_),
    .Y(_03475_),
    .A1(_09122_),
    .A2(_03473_));
 sg13g2_and2_1 _20946_ (.A(net149),
    .B(_03475_),
    .X(_03476_));
 sg13g2_nor3_1 _20947_ (.A(_03243_),
    .B(_03174_),
    .C(_03456_),
    .Y(_03477_));
 sg13g2_nor3_1 _20948_ (.A(_03162_),
    .B(_03476_),
    .C(_03477_),
    .Y(_03478_));
 sg13g2_nor3_1 _20949_ (.A(net823),
    .B(_03099_),
    .C(_03332_),
    .Y(_03479_));
 sg13g2_or2_1 _20950_ (.X(_03480_),
    .B(_10723_),
    .A(net1146));
 sg13g2_o21ai_1 _20951_ (.B1(_09006_),
    .Y(_03481_),
    .A1(_03036_),
    .A2(_03480_));
 sg13g2_a221oi_1 _20952_ (.B2(net230),
    .C1(_03477_),
    .B1(_03481_),
    .A1(_03284_),
    .Y(_03482_),
    .A2(_09067_));
 sg13g2_o21ai_1 _20953_ (.B1(_03482_),
    .Y(_03483_),
    .A1(_03121_),
    .A2(_03479_));
 sg13g2_a21oi_1 _20954_ (.A1(_08942_),
    .A2(_03154_),
    .Y(_03484_),
    .B1(_08921_));
 sg13g2_o21ai_1 _20955_ (.B1(_03370_),
    .Y(_03485_),
    .A1(_03101_),
    .A2(_03484_));
 sg13g2_nand3_1 _20956_ (.B(_03048_),
    .C(_03485_),
    .A(_03464_),
    .Y(_03486_));
 sg13g2_a21oi_1 _20957_ (.A1(_03483_),
    .A2(_03486_),
    .Y(_03487_),
    .B1(_03041_));
 sg13g2_nor4_1 _20958_ (.A(_03468_),
    .B(_03472_),
    .C(_03478_),
    .D(_03487_),
    .Y(_03488_));
 sg13g2_mux2_1 _20959_ (.A0(_09208_),
    .A1(_03488_),
    .S(net146),
    .X(_00783_));
 sg13g2_buf_1 _20960_ (.A(net1145),
    .X(_03489_));
 sg13g2_buf_1 _20961_ (.A(_03489_),
    .X(_03490_));
 sg13g2_nand2b_1 _20962_ (.Y(_03491_),
    .B(net1125),
    .A_N(net1124));
 sg13g2_buf_1 _20963_ (.A(_03491_),
    .X(_03492_));
 sg13g2_nand3b_1 _20964_ (.B(net1127),
    .C(net1126),
    .Y(_03493_),
    .A_N(net1052));
 sg13g2_buf_1 _20965_ (.A(_03493_),
    .X(_03494_));
 sg13g2_nor2_1 _20966_ (.A(_03492_),
    .B(_03494_),
    .Y(_03495_));
 sg13g2_buf_1 _20967_ (.A(_03495_),
    .X(_03496_));
 sg13g2_buf_1 _20968_ (.A(net606),
    .X(_03497_));
 sg13g2_mux2_1 _20969_ (.A0(\cpu.ex.r_10[0] ),
    .A1(net861),
    .S(net553),
    .X(_00788_));
 sg13g2_nand2_1 _20970_ (.Y(_03498_),
    .A(net995),
    .B(net606));
 sg13g2_o21ai_1 _20971_ (.B1(_03498_),
    .Y(_00789_),
    .A1(_10413_),
    .A2(net553));
 sg13g2_mux2_1 _20972_ (.A0(\cpu.ex.r_10[11] ),
    .A1(net862),
    .S(net553),
    .X(_00790_));
 sg13g2_buf_1 _20973_ (.A(net617),
    .X(_03499_));
 sg13g2_buf_1 _20974_ (.A(net552),
    .X(_03500_));
 sg13g2_mux2_1 _20975_ (.A0(\cpu.ex.r_10[12] ),
    .A1(net494),
    .S(net553),
    .X(_00791_));
 sg13g2_buf_1 _20976_ (.A(net577),
    .X(_03501_));
 sg13g2_buf_1 _20977_ (.A(net493),
    .X(_03502_));
 sg13g2_mux2_1 _20978_ (.A0(\cpu.ex.r_10[13] ),
    .A1(net454),
    .S(_03497_),
    .X(_00792_));
 sg13g2_buf_1 _20979_ (.A(net688),
    .X(_03503_));
 sg13g2_buf_1 _20980_ (.A(net605),
    .X(_03504_));
 sg13g2_mux2_1 _20981_ (.A0(\cpu.ex.r_10[14] ),
    .A1(net551),
    .S(net553),
    .X(_00793_));
 sg13g2_buf_1 _20982_ (.A(net1086),
    .X(_03505_));
 sg13g2_buf_1 _20983_ (.A(net860),
    .X(_03506_));
 sg13g2_mux2_1 _20984_ (.A0(\cpu.ex.r_10[15] ),
    .A1(net746),
    .S(net553),
    .X(_00794_));
 sg13g2_buf_2 _20985_ (.A(net623),
    .X(_03507_));
 sg13g2_buf_1 _20986_ (.A(net550),
    .X(_03508_));
 sg13g2_mux2_1 _20987_ (.A0(\cpu.ex.r_10[1] ),
    .A1(net492),
    .S(net553),
    .X(_00795_));
 sg13g2_buf_1 _20988_ (.A(_12475_),
    .X(_03509_));
 sg13g2_buf_1 _20989_ (.A(net491),
    .X(_03510_));
 sg13g2_mux2_1 _20990_ (.A0(\cpu.ex.r_10[2] ),
    .A1(net453),
    .S(_03497_),
    .X(_00796_));
 sg13g2_buf_1 _20991_ (.A(net463),
    .X(_03511_));
 sg13g2_mux2_1 _20992_ (.A0(\cpu.ex.r_10[3] ),
    .A1(net410),
    .S(net606),
    .X(_00797_));
 sg13g2_buf_1 _20993_ (.A(net563),
    .X(_03512_));
 sg13g2_buf_2 _20994_ (.A(net490),
    .X(_03513_));
 sg13g2_nand2_1 _20995_ (.Y(_03514_),
    .A(net452),
    .B(_03496_));
 sg13g2_o21ai_1 _20996_ (.B1(_03514_),
    .Y(_00798_),
    .A1(_10780_),
    .A2(net553));
 sg13g2_mux2_1 _20997_ (.A0(\cpu.ex.r_10[5] ),
    .A1(net607),
    .S(net606),
    .X(_00799_));
 sg13g2_mux2_1 _20998_ (.A0(\cpu.ex.r_10[6] ),
    .A1(net747),
    .S(net606),
    .X(_00800_));
 sg13g2_mux2_1 _20999_ (.A0(\cpu.ex.r_10[7] ),
    .A1(_02982_),
    .S(net606),
    .X(_00801_));
 sg13g2_mux2_1 _21000_ (.A0(\cpu.ex.r_10[8] ),
    .A1(_02984_),
    .S(net606),
    .X(_00802_));
 sg13g2_mux2_1 _21001_ (.A0(\cpu.ex.r_10[9] ),
    .A1(net865),
    .S(net606),
    .X(_00803_));
 sg13g2_nor2_1 _21002_ (.A(_10197_),
    .B(_03494_),
    .Y(_03515_));
 sg13g2_buf_4 _21003_ (.X(_03516_),
    .A(_03515_));
 sg13g2_buf_1 _21004_ (.A(_03516_),
    .X(_03517_));
 sg13g2_mux2_1 _21005_ (.A0(\cpu.ex.r_11[0] ),
    .A1(net861),
    .S(_03517_),
    .X(_00804_));
 sg13g2_mux2_1 _21006_ (.A0(\cpu.ex.r_11[10] ),
    .A1(net864),
    .S(net549),
    .X(_00805_));
 sg13g2_mux2_1 _21007_ (.A0(\cpu.ex.r_11[11] ),
    .A1(net862),
    .S(net549),
    .X(_00806_));
 sg13g2_mux2_1 _21008_ (.A0(\cpu.ex.r_11[12] ),
    .A1(net494),
    .S(net549),
    .X(_00807_));
 sg13g2_mux2_1 _21009_ (.A0(\cpu.ex.r_11[13] ),
    .A1(net454),
    .S(net549),
    .X(_00808_));
 sg13g2_nand2_1 _21010_ (.Y(_03518_),
    .A(net605),
    .B(_03516_));
 sg13g2_o21ai_1 _21011_ (.B1(_03518_),
    .Y(_00809_),
    .A1(_11142_),
    .A2(net549));
 sg13g2_mux2_1 _21012_ (.A0(\cpu.ex.r_11[15] ),
    .A1(net746),
    .S(net549),
    .X(_00810_));
 sg13g2_mux2_1 _21013_ (.A0(\cpu.ex.r_11[1] ),
    .A1(_03508_),
    .S(net549),
    .X(_00811_));
 sg13g2_mux2_1 _21014_ (.A0(\cpu.ex.r_11[2] ),
    .A1(net453),
    .S(_03517_),
    .X(_00812_));
 sg13g2_mux2_1 _21015_ (.A0(\cpu.ex.r_11[3] ),
    .A1(_03511_),
    .S(net549),
    .X(_00813_));
 sg13g2_buf_1 _21016_ (.A(net452),
    .X(_03519_));
 sg13g2_mux2_1 _21017_ (.A0(\cpu.ex.r_11[4] ),
    .A1(net409),
    .S(_03516_),
    .X(_00814_));
 sg13g2_mux2_1 _21018_ (.A0(\cpu.ex.r_11[5] ),
    .A1(net607),
    .S(_03516_),
    .X(_00815_));
 sg13g2_mux2_1 _21019_ (.A0(\cpu.ex.r_11[6] ),
    .A1(net747),
    .S(_03516_),
    .X(_00816_));
 sg13g2_mux2_1 _21020_ (.A0(\cpu.ex.r_11[7] ),
    .A1(net867),
    .S(_03516_),
    .X(_00817_));
 sg13g2_mux2_1 _21021_ (.A0(\cpu.ex.r_11[8] ),
    .A1(net866),
    .S(_03516_),
    .X(_00818_));
 sg13g2_mux2_1 _21022_ (.A0(\cpu.ex.r_11[9] ),
    .A1(_02986_),
    .S(_03516_),
    .X(_00819_));
 sg13g2_nand3_1 _21023_ (.B(net1052),
    .C(_10188_),
    .A(net1126),
    .Y(_03520_));
 sg13g2_buf_1 _21024_ (.A(_03520_),
    .X(_03521_));
 sg13g2_nor3_1 _21025_ (.A(net1125),
    .B(_10196_),
    .C(_03521_),
    .Y(_03522_));
 sg13g2_buf_2 _21026_ (.A(_03522_),
    .X(_03523_));
 sg13g2_buf_1 _21027_ (.A(_03523_),
    .X(_03524_));
 sg13g2_mux2_1 _21028_ (.A0(\cpu.ex.r_12[0] ),
    .A1(net861),
    .S(_03524_),
    .X(_00820_));
 sg13g2_mux2_1 _21029_ (.A0(\cpu.ex.r_12[10] ),
    .A1(net864),
    .S(net548),
    .X(_00821_));
 sg13g2_mux2_1 _21030_ (.A0(\cpu.ex.r_12[11] ),
    .A1(net862),
    .S(net548),
    .X(_00822_));
 sg13g2_mux2_1 _21031_ (.A0(\cpu.ex.r_12[12] ),
    .A1(net494),
    .S(net548),
    .X(_00823_));
 sg13g2_mux2_1 _21032_ (.A0(\cpu.ex.r_12[13] ),
    .A1(net454),
    .S(_03524_),
    .X(_00824_));
 sg13g2_mux2_1 _21033_ (.A0(\cpu.ex.r_12[14] ),
    .A1(net551),
    .S(net548),
    .X(_00825_));
 sg13g2_mux2_1 _21034_ (.A0(\cpu.ex.r_12[15] ),
    .A1(net746),
    .S(net548),
    .X(_00826_));
 sg13g2_mux2_1 _21035_ (.A0(\cpu.ex.r_12[1] ),
    .A1(net492),
    .S(net548),
    .X(_00827_));
 sg13g2_mux2_1 _21036_ (.A0(\cpu.ex.r_12[2] ),
    .A1(net453),
    .S(net548),
    .X(_00828_));
 sg13g2_mux2_1 _21037_ (.A0(\cpu.ex.r_12[3] ),
    .A1(net410),
    .S(net548),
    .X(_00829_));
 sg13g2_mux2_1 _21038_ (.A0(\cpu.ex.r_12[4] ),
    .A1(_03519_),
    .S(_03523_),
    .X(_00830_));
 sg13g2_mux2_1 _21039_ (.A0(\cpu.ex.r_12[5] ),
    .A1(net607),
    .S(_03523_),
    .X(_00831_));
 sg13g2_mux2_1 _21040_ (.A0(\cpu.ex.r_12[6] ),
    .A1(_03009_),
    .S(_03523_),
    .X(_00832_));
 sg13g2_mux2_1 _21041_ (.A0(\cpu.ex.r_12[7] ),
    .A1(net867),
    .S(_03523_),
    .X(_00833_));
 sg13g2_mux2_1 _21042_ (.A0(\cpu.ex.r_12[8] ),
    .A1(net866),
    .S(_03523_),
    .X(_00834_));
 sg13g2_mux2_1 _21043_ (.A0(\cpu.ex.r_12[9] ),
    .A1(_02986_),
    .S(_03523_),
    .X(_00835_));
 sg13g2_nand2b_1 _21044_ (.Y(_03525_),
    .B(net1124),
    .A_N(_10195_));
 sg13g2_buf_1 _21045_ (.A(_03525_),
    .X(_03526_));
 sg13g2_nor2_1 _21046_ (.A(_03521_),
    .B(_03526_),
    .Y(_03527_));
 sg13g2_buf_2 _21047_ (.A(_03527_),
    .X(_03528_));
 sg13g2_buf_1 _21048_ (.A(_03528_),
    .X(_03529_));
 sg13g2_nand2_1 _21049_ (.Y(_03530_),
    .A(_03490_),
    .B(_03528_));
 sg13g2_o21ai_1 _21050_ (.B1(_03530_),
    .Y(_00836_),
    .A1(_10656_),
    .A2(_03529_));
 sg13g2_mux2_1 _21051_ (.A0(\cpu.ex.r_13[10] ),
    .A1(_02988_),
    .S(net547),
    .X(_00837_));
 sg13g2_mux2_1 _21052_ (.A0(\cpu.ex.r_13[11] ),
    .A1(net862),
    .S(net547),
    .X(_00838_));
 sg13g2_mux2_1 _21053_ (.A0(\cpu.ex.r_13[12] ),
    .A1(net494),
    .S(net547),
    .X(_00839_));
 sg13g2_mux2_1 _21054_ (.A0(\cpu.ex.r_13[13] ),
    .A1(net454),
    .S(net547),
    .X(_00840_));
 sg13g2_mux2_1 _21055_ (.A0(\cpu.ex.r_13[14] ),
    .A1(net551),
    .S(net547),
    .X(_00841_));
 sg13g2_mux2_1 _21056_ (.A0(\cpu.ex.r_13[15] ),
    .A1(_03506_),
    .S(_03529_),
    .X(_00842_));
 sg13g2_mux2_1 _21057_ (.A0(\cpu.ex.r_13[1] ),
    .A1(net492),
    .S(net547),
    .X(_00843_));
 sg13g2_mux2_1 _21058_ (.A0(\cpu.ex.r_13[2] ),
    .A1(net453),
    .S(net547),
    .X(_00844_));
 sg13g2_mux2_1 _21059_ (.A0(\cpu.ex.r_13[3] ),
    .A1(net410),
    .S(net547),
    .X(_00845_));
 sg13g2_mux2_1 _21060_ (.A0(\cpu.ex.r_13[4] ),
    .A1(net409),
    .S(_03528_),
    .X(_00846_));
 sg13g2_mux2_1 _21061_ (.A0(\cpu.ex.r_13[5] ),
    .A1(_02977_),
    .S(_03528_),
    .X(_00847_));
 sg13g2_mux2_1 _21062_ (.A0(\cpu.ex.r_13[6] ),
    .A1(_03009_),
    .S(_03528_),
    .X(_00848_));
 sg13g2_mux2_1 _21063_ (.A0(\cpu.ex.r_13[7] ),
    .A1(_02982_),
    .S(_03528_),
    .X(_00849_));
 sg13g2_mux2_1 _21064_ (.A0(\cpu.ex.r_13[8] ),
    .A1(_02984_),
    .S(_03528_),
    .X(_00850_));
 sg13g2_mux2_1 _21065_ (.A0(\cpu.ex.r_13[9] ),
    .A1(net865),
    .S(_03528_),
    .X(_00851_));
 sg13g2_nor2_1 _21066_ (.A(_03492_),
    .B(_03521_),
    .Y(_03531_));
 sg13g2_buf_2 _21067_ (.A(_03531_),
    .X(_03532_));
 sg13g2_buf_1 _21068_ (.A(_03532_),
    .X(_03533_));
 sg13g2_mux2_1 _21069_ (.A0(\cpu.ex.r_14[0] ),
    .A1(net861),
    .S(_03533_),
    .X(_00852_));
 sg13g2_mux2_1 _21070_ (.A0(\cpu.ex.r_14[10] ),
    .A1(_02988_),
    .S(net546),
    .X(_00853_));
 sg13g2_mux2_1 _21071_ (.A0(\cpu.ex.r_14[11] ),
    .A1(_03011_),
    .S(net546),
    .X(_00854_));
 sg13g2_mux2_1 _21072_ (.A0(\cpu.ex.r_14[12] ),
    .A1(net494),
    .S(net546),
    .X(_00855_));
 sg13g2_mux2_1 _21073_ (.A0(\cpu.ex.r_14[13] ),
    .A1(_03502_),
    .S(_03533_),
    .X(_00856_));
 sg13g2_mux2_1 _21074_ (.A0(\cpu.ex.r_14[14] ),
    .A1(net551),
    .S(net546),
    .X(_00857_));
 sg13g2_mux2_1 _21075_ (.A0(\cpu.ex.r_14[15] ),
    .A1(net746),
    .S(net546),
    .X(_00858_));
 sg13g2_mux2_1 _21076_ (.A0(\cpu.ex.r_14[1] ),
    .A1(net492),
    .S(net546),
    .X(_00859_));
 sg13g2_mux2_1 _21077_ (.A0(\cpu.ex.r_14[2] ),
    .A1(_03510_),
    .S(net546),
    .X(_00860_));
 sg13g2_mux2_1 _21078_ (.A0(\cpu.ex.r_14[3] ),
    .A1(net410),
    .S(net546),
    .X(_00861_));
 sg13g2_mux2_1 _21079_ (.A0(\cpu.ex.r_14[4] ),
    .A1(net409),
    .S(_03532_),
    .X(_00862_));
 sg13g2_mux2_1 _21080_ (.A0(\cpu.ex.r_14[5] ),
    .A1(_02977_),
    .S(_03532_),
    .X(_00863_));
 sg13g2_mux2_1 _21081_ (.A0(\cpu.ex.r_14[6] ),
    .A1(net747),
    .S(_03532_),
    .X(_00864_));
 sg13g2_mux2_1 _21082_ (.A0(\cpu.ex.r_14[7] ),
    .A1(net867),
    .S(_03532_),
    .X(_00865_));
 sg13g2_mux2_1 _21083_ (.A0(\cpu.ex.r_14[8] ),
    .A1(net866),
    .S(_03532_),
    .X(_00866_));
 sg13g2_buf_1 _21084_ (.A(_02985_),
    .X(_03534_));
 sg13g2_mux2_1 _21085_ (.A0(\cpu.ex.r_14[9] ),
    .A1(net859),
    .S(_03532_),
    .X(_00867_));
 sg13g2_nor2_1 _21086_ (.A(_10197_),
    .B(_03521_),
    .Y(_03535_));
 sg13g2_buf_2 _21087_ (.A(_03535_),
    .X(_03536_));
 sg13g2_buf_1 _21088_ (.A(_03536_),
    .X(_03537_));
 sg13g2_mux2_1 _21089_ (.A0(\cpu.ex.r_15[0] ),
    .A1(net861),
    .S(_03537_),
    .X(_00868_));
 sg13g2_buf_1 _21090_ (.A(net995),
    .X(_03538_));
 sg13g2_mux2_1 _21091_ (.A0(\cpu.ex.r_15[10] ),
    .A1(net858),
    .S(net545),
    .X(_00869_));
 sg13g2_mux2_1 _21092_ (.A0(\cpu.ex.r_15[11] ),
    .A1(net862),
    .S(net545),
    .X(_00870_));
 sg13g2_mux2_1 _21093_ (.A0(\cpu.ex.r_15[12] ),
    .A1(net494),
    .S(net545),
    .X(_00871_));
 sg13g2_mux2_1 _21094_ (.A0(\cpu.ex.r_15[13] ),
    .A1(_03502_),
    .S(_03537_),
    .X(_00872_));
 sg13g2_mux2_1 _21095_ (.A0(\cpu.ex.r_15[14] ),
    .A1(net551),
    .S(net545),
    .X(_00873_));
 sg13g2_mux2_1 _21096_ (.A0(\cpu.ex.r_15[15] ),
    .A1(net746),
    .S(net545),
    .X(_00874_));
 sg13g2_mux2_1 _21097_ (.A0(\cpu.ex.r_15[1] ),
    .A1(net492),
    .S(net545),
    .X(_00875_));
 sg13g2_mux2_1 _21098_ (.A0(\cpu.ex.r_15[2] ),
    .A1(_03510_),
    .S(net545),
    .X(_00876_));
 sg13g2_mux2_1 _21099_ (.A0(\cpu.ex.r_15[3] ),
    .A1(net410),
    .S(net545),
    .X(_00877_));
 sg13g2_mux2_1 _21100_ (.A0(\cpu.ex.r_15[4] ),
    .A1(net409),
    .S(_03536_),
    .X(_00878_));
 sg13g2_buf_2 _21101_ (.A(net888),
    .X(_03539_));
 sg13g2_buf_1 _21102_ (.A(net745),
    .X(_03540_));
 sg13g2_mux2_1 _21103_ (.A0(\cpu.ex.r_15[5] ),
    .A1(net667),
    .S(_03536_),
    .X(_00879_));
 sg13g2_mux2_1 _21104_ (.A0(\cpu.ex.r_15[6] ),
    .A1(net747),
    .S(_03536_),
    .X(_00880_));
 sg13g2_buf_1 _21105_ (.A(net1138),
    .X(_03541_));
 sg13g2_mux2_1 _21106_ (.A0(\cpu.ex.r_15[7] ),
    .A1(net992),
    .S(_03536_),
    .X(_00881_));
 sg13g2_buf_1 _21107_ (.A(net997),
    .X(_03542_));
 sg13g2_mux2_1 _21108_ (.A0(\cpu.ex.r_15[8] ),
    .A1(net857),
    .S(_03536_),
    .X(_00882_));
 sg13g2_mux2_1 _21109_ (.A0(\cpu.ex.r_15[9] ),
    .A1(net859),
    .S(_03536_),
    .X(_00883_));
 sg13g2_nor3_1 _21110_ (.A(net1125),
    .B(net1124),
    .C(_03494_),
    .Y(_03543_));
 sg13g2_buf_4 _21111_ (.X(_03544_),
    .A(_03543_));
 sg13g2_buf_1 _21112_ (.A(_03544_),
    .X(_03545_));
 sg13g2_mux2_1 _21113_ (.A0(\cpu.ex.r_8[0] ),
    .A1(net861),
    .S(_03545_),
    .X(_00884_));
 sg13g2_mux2_1 _21114_ (.A0(\cpu.ex.r_8[10] ),
    .A1(net858),
    .S(net544),
    .X(_00885_));
 sg13g2_mux2_1 _21115_ (.A0(\cpu.ex.r_8[11] ),
    .A1(net862),
    .S(net544),
    .X(_00886_));
 sg13g2_mux2_1 _21116_ (.A0(\cpu.ex.r_8[12] ),
    .A1(net494),
    .S(net544),
    .X(_00887_));
 sg13g2_mux2_1 _21117_ (.A0(\cpu.ex.r_8[13] ),
    .A1(net454),
    .S(_03545_),
    .X(_00888_));
 sg13g2_nand2_1 _21118_ (.Y(_03546_),
    .A(net605),
    .B(_03544_));
 sg13g2_o21ai_1 _21119_ (.B1(_03546_),
    .Y(_00889_),
    .A1(_10468_),
    .A2(net544));
 sg13g2_mux2_1 _21120_ (.A0(\cpu.ex.r_8[15] ),
    .A1(net746),
    .S(net544),
    .X(_00890_));
 sg13g2_mux2_1 _21121_ (.A0(\cpu.ex.r_8[1] ),
    .A1(net492),
    .S(net544),
    .X(_00891_));
 sg13g2_mux2_1 _21122_ (.A0(\cpu.ex.r_8[2] ),
    .A1(net453),
    .S(net544),
    .X(_00892_));
 sg13g2_mux2_1 _21123_ (.A0(\cpu.ex.r_8[3] ),
    .A1(net410),
    .S(net544),
    .X(_00893_));
 sg13g2_mux2_1 _21124_ (.A0(\cpu.ex.r_8[4] ),
    .A1(net409),
    .S(_03544_),
    .X(_00894_));
 sg13g2_mux2_1 _21125_ (.A0(\cpu.ex.r_8[5] ),
    .A1(net667),
    .S(_03544_),
    .X(_00895_));
 sg13g2_mux2_1 _21126_ (.A0(\cpu.ex.r_8[6] ),
    .A1(net747),
    .S(_03544_),
    .X(_00896_));
 sg13g2_mux2_1 _21127_ (.A0(\cpu.ex.r_8[7] ),
    .A1(net992),
    .S(_03544_),
    .X(_00897_));
 sg13g2_mux2_1 _21128_ (.A0(\cpu.ex.r_8[8] ),
    .A1(net857),
    .S(_03544_),
    .X(_00898_));
 sg13g2_mux2_1 _21129_ (.A0(\cpu.ex.r_8[9] ),
    .A1(net859),
    .S(_03544_),
    .X(_00899_));
 sg13g2_nor2_1 _21130_ (.A(_03494_),
    .B(_03526_),
    .Y(_03547_));
 sg13g2_buf_2 _21131_ (.A(_03547_),
    .X(_03548_));
 sg13g2_buf_1 _21132_ (.A(_03548_),
    .X(_03549_));
 sg13g2_mux2_1 _21133_ (.A0(\cpu.ex.r_9[0] ),
    .A1(net861),
    .S(net543),
    .X(_00900_));
 sg13g2_mux2_1 _21134_ (.A0(\cpu.ex.r_9[10] ),
    .A1(net858),
    .S(net543),
    .X(_00901_));
 sg13g2_mux2_1 _21135_ (.A0(\cpu.ex.r_9[11] ),
    .A1(net862),
    .S(_03549_),
    .X(_00902_));
 sg13g2_buf_1 _21136_ (.A(_10341_),
    .X(_03550_));
 sg13g2_mux2_1 _21137_ (.A0(\cpu.ex.r_9[12] ),
    .A1(net542),
    .S(net543),
    .X(_00903_));
 sg13g2_buf_1 _21138_ (.A(net577),
    .X(_03551_));
 sg13g2_mux2_1 _21139_ (.A0(\cpu.ex.r_9[13] ),
    .A1(net489),
    .S(net543),
    .X(_00904_));
 sg13g2_mux2_1 _21140_ (.A0(\cpu.ex.r_9[14] ),
    .A1(_03504_),
    .S(net543),
    .X(_00905_));
 sg13g2_mux2_1 _21141_ (.A0(\cpu.ex.r_9[15] ),
    .A1(_03506_),
    .S(net543),
    .X(_00906_));
 sg13g2_mux2_1 _21142_ (.A0(\cpu.ex.r_9[1] ),
    .A1(net492),
    .S(net543),
    .X(_00907_));
 sg13g2_mux2_1 _21143_ (.A0(\cpu.ex.r_9[2] ),
    .A1(net453),
    .S(net543),
    .X(_00908_));
 sg13g2_mux2_1 _21144_ (.A0(\cpu.ex.r_9[3] ),
    .A1(net410),
    .S(_03549_),
    .X(_00909_));
 sg13g2_mux2_1 _21145_ (.A0(\cpu.ex.r_9[4] ),
    .A1(net409),
    .S(_03548_),
    .X(_00910_));
 sg13g2_mux2_1 _21146_ (.A0(\cpu.ex.r_9[5] ),
    .A1(net667),
    .S(_03548_),
    .X(_00911_));
 sg13g2_mux2_1 _21147_ (.A0(\cpu.ex.r_9[6] ),
    .A1(net747),
    .S(_03548_),
    .X(_00912_));
 sg13g2_mux2_1 _21148_ (.A0(\cpu.ex.r_9[7] ),
    .A1(net992),
    .S(_03548_),
    .X(_00913_));
 sg13g2_mux2_1 _21149_ (.A0(\cpu.ex.r_9[8] ),
    .A1(net857),
    .S(_03548_),
    .X(_00914_));
 sg13g2_mux2_1 _21150_ (.A0(\cpu.ex.r_9[9] ),
    .A1(net859),
    .S(_03548_),
    .X(_00915_));
 sg13g2_nand2_1 _21151_ (.Y(_03552_),
    .A(_09155_),
    .B(_11485_));
 sg13g2_buf_1 _21152_ (.A(_03552_),
    .X(_03553_));
 sg13g2_nand2_1 _21153_ (.Y(_03554_),
    .A(net1074),
    .B(_11491_));
 sg13g2_buf_1 _21154_ (.A(_03554_),
    .X(_03555_));
 sg13g2_nand2_1 _21155_ (.Y(_03556_),
    .A(net141),
    .B(_03555_));
 sg13g2_buf_2 _21156_ (.A(_03556_),
    .X(_03557_));
 sg13g2_and3_1 _21157_ (.X(_03558_),
    .A(_08423_),
    .B(_08467_),
    .C(_11046_));
 sg13g2_buf_2 _21158_ (.A(_03558_),
    .X(_03559_));
 sg13g2_buf_8 _21159_ (.A(_03559_),
    .X(_03560_));
 sg13g2_nor2_2 _21160_ (.A(net758),
    .B(_03560_),
    .Y(_03561_));
 sg13g2_buf_8 _21161_ (.A(_11048_),
    .X(_03562_));
 sg13g2_a21oi_1 _21162_ (.A1(net1036),
    .A2(net350),
    .Y(_03563_),
    .B1(_11119_));
 sg13g2_a21o_1 _21163_ (.A2(_03561_),
    .A1(_11087_),
    .B1(_03563_),
    .X(_03564_));
 sg13g2_buf_2 _21164_ (.A(_03564_),
    .X(_03565_));
 sg13g2_buf_1 _21165_ (.A(_03565_),
    .X(_03566_));
 sg13g2_buf_1 _21166_ (.A(_03566_),
    .X(_03567_));
 sg13g2_buf_1 _21167_ (.A(_11186_),
    .X(_03568_));
 sg13g2_mux2_1 _21168_ (.A0(_10385_),
    .A1(_11203_),
    .S(net209),
    .X(_03569_));
 sg13g2_buf_2 _21169_ (.A(_03569_),
    .X(_03570_));
 sg13g2_inv_1 _21170_ (.Y(_03571_),
    .A(_03570_));
 sg13g2_nand2_1 _21171_ (.Y(_03572_),
    .A(_11398_),
    .B(_03571_));
 sg13g2_nand3_1 _21172_ (.B(_10740_),
    .C(net350),
    .A(net1117),
    .Y(_03573_));
 sg13g2_buf_1 _21173_ (.A(_03573_),
    .X(_03574_));
 sg13g2_o21ai_1 _21174_ (.B1(_11925_),
    .Y(_03575_),
    .A1(net890),
    .A2(_03559_));
 sg13g2_nand2_1 _21175_ (.Y(_03576_),
    .A(_03574_),
    .B(_03575_));
 sg13g2_buf_2 _21176_ (.A(_03576_),
    .X(_03577_));
 sg13g2_nand2_1 _21177_ (.Y(_03578_),
    .A(net235),
    .B(_03577_));
 sg13g2_nand3_1 _21178_ (.B(net1036),
    .C(net350),
    .A(net939),
    .Y(_03579_));
 sg13g2_buf_1 _21179_ (.A(_03579_),
    .X(_03580_));
 sg13g2_inv_1 _21180_ (.Y(_03581_),
    .A(_11297_));
 sg13g2_o21ai_1 _21181_ (.B1(_03581_),
    .Y(_03582_),
    .A1(net890),
    .A2(net351));
 sg13g2_nor2_1 _21182_ (.A(net285),
    .B(_10998_),
    .Y(_03583_));
 sg13g2_inv_1 _21183_ (.Y(_03584_),
    .A(_10612_));
 sg13g2_nor4_1 _21184_ (.A(net758),
    .B(_03584_),
    .C(net285),
    .D(net351),
    .Y(_03585_));
 sg13g2_a221oi_1 _21185_ (.B2(_03568_),
    .C1(_03585_),
    .B1(_03583_),
    .A1(_03580_),
    .Y(_03586_),
    .A2(_03582_));
 sg13g2_nand4_1 _21186_ (.B(_10616_),
    .C(_11922_),
    .A(_10611_),
    .Y(_03587_),
    .D(_11297_));
 sg13g2_a21oi_1 _21187_ (.A1(net1036),
    .A2(net350),
    .Y(_03588_),
    .B1(_03587_));
 sg13g2_nor2_1 _21188_ (.A(net939),
    .B(_03584_),
    .Y(_03589_));
 sg13g2_and4_1 _21189_ (.A(net1036),
    .B(net237),
    .C(_03562_),
    .D(_03589_),
    .X(_03590_));
 sg13g2_nor3_1 _21190_ (.A(net281),
    .B(_03588_),
    .C(_03590_),
    .Y(_03591_));
 sg13g2_nand3_1 _21191_ (.B(_03574_),
    .C(_03575_),
    .A(net282),
    .Y(_03592_));
 sg13g2_o21ai_1 _21192_ (.B1(_03592_),
    .Y(_03593_),
    .A1(_03586_),
    .A2(_03591_));
 sg13g2_nand2_1 _21193_ (.Y(_03594_),
    .A(_03578_),
    .B(_03593_));
 sg13g2_nand3b_1 _21194_ (.B(_11048_),
    .C(net1117),
    .Y(_03595_),
    .A_N(_10582_));
 sg13g2_buf_1 _21195_ (.A(_03595_),
    .X(_03596_));
 sg13g2_o21ai_1 _21196_ (.B1(_11920_),
    .Y(_03597_),
    .A1(net890),
    .A2(_03559_));
 sg13g2_nand2_1 _21197_ (.Y(_03598_),
    .A(_03596_),
    .B(_03597_));
 sg13g2_buf_2 _21198_ (.A(_03598_),
    .X(_03599_));
 sg13g2_nand2_1 _21199_ (.Y(_03600_),
    .A(net286),
    .B(_03599_));
 sg13g2_and2_1 _21200_ (.A(net280),
    .B(_11037_),
    .X(_03601_));
 sg13g2_nor4_1 _21201_ (.A(net758),
    .B(_10644_),
    .C(net284),
    .D(net351),
    .Y(_03602_));
 sg13g2_a221oi_1 _21202_ (.B2(net241),
    .C1(_03602_),
    .B1(_03601_),
    .A1(_10869_),
    .Y(_03603_),
    .A2(net279));
 sg13g2_nor2_1 _21203_ (.A(net280),
    .B(_11037_),
    .Y(_03604_));
 sg13g2_nor4_1 _21204_ (.A(net758),
    .B(_10643_),
    .C(net280),
    .D(net351),
    .Y(_03605_));
 sg13g2_a21o_1 _21205_ (.A2(_03604_),
    .A1(net241),
    .B1(_03605_),
    .X(_03606_));
 sg13g2_nand3_1 _21206_ (.B(_03596_),
    .C(_03597_),
    .A(net360),
    .Y(_03607_));
 sg13g2_o21ai_1 _21207_ (.B1(_03607_),
    .Y(_03608_),
    .A1(_03603_),
    .A2(_03606_));
 sg13g2_nand2_1 _21208_ (.Y(_03609_),
    .A(_03580_),
    .B(_03582_));
 sg13g2_buf_2 _21209_ (.A(_03609_),
    .X(_03610_));
 sg13g2_nand2_1 _21210_ (.Y(_03611_),
    .A(net277),
    .B(_03610_));
 sg13g2_nor3_2 _21211_ (.A(net890),
    .B(_10612_),
    .C(_03559_),
    .Y(_03612_));
 sg13g2_a21oi_2 _21212_ (.B1(_11922_),
    .Y(_03613_),
    .A2(_11048_),
    .A1(net1117));
 sg13g2_or2_1 _21213_ (.X(_03614_),
    .B(_03613_),
    .A(_03612_));
 sg13g2_buf_1 _21214_ (.A(_03614_),
    .X(_03615_));
 sg13g2_buf_1 _21215_ (.A(_03615_),
    .X(_03616_));
 sg13g2_a22oi_1 _21216_ (.Y(_03617_),
    .B1(net208),
    .B2(net285),
    .A2(_03577_),
    .A1(net235));
 sg13g2_nand4_1 _21217_ (.B(_03608_),
    .C(_03611_),
    .A(_03600_),
    .Y(_03618_),
    .D(_03617_));
 sg13g2_buf_1 _21218_ (.A(_03618_),
    .X(_03619_));
 sg13g2_nand3_1 _21219_ (.B(_10816_),
    .C(net350),
    .A(net1036),
    .Y(_03620_));
 sg13g2_o21ai_1 _21220_ (.B1(_03620_),
    .Y(_03621_),
    .A1(_03561_),
    .A2(_11277_));
 sg13g2_buf_2 _21221_ (.A(_03621_),
    .X(_03622_));
 sg13g2_nor3_1 _21222_ (.A(_11935_),
    .B(_10487_),
    .C(net351),
    .Y(_03623_));
 sg13g2_a21oi_2 _21223_ (.B1(_03623_),
    .Y(_03624_),
    .A2(_11320_),
    .A1(net209));
 sg13g2_nor3_1 _21224_ (.A(net758),
    .B(_10733_),
    .C(net351),
    .Y(_03625_));
 sg13g2_a21oi_1 _21225_ (.A1(net1036),
    .A2(net350),
    .Y(_03626_),
    .B1(_11929_));
 sg13g2_nor2_1 _21226_ (.A(_03625_),
    .B(_03626_),
    .Y(_03627_));
 sg13g2_buf_2 _21227_ (.A(_03627_),
    .X(_03628_));
 sg13g2_nor3_2 _21228_ (.A(net758),
    .B(_10547_),
    .C(_03560_),
    .Y(_03629_));
 sg13g2_inv_1 _21229_ (.Y(_03630_),
    .A(_11219_));
 sg13g2_a21oi_1 _21230_ (.A1(_11477_),
    .A2(net350),
    .Y(_03631_),
    .B1(_03630_));
 sg13g2_nor3_1 _21231_ (.A(_11669_),
    .B(_03629_),
    .C(_03631_),
    .Y(_03632_));
 sg13g2_a221oi_1 _21232_ (.B2(net283),
    .C1(_03632_),
    .B1(_03628_),
    .A1(_10522_),
    .Y(_03633_),
    .A2(_03624_));
 sg13g2_buf_1 _21233_ (.A(_03633_),
    .X(_03634_));
 sg13g2_and2_1 _21234_ (.A(_11245_),
    .B(_03634_),
    .X(_03635_));
 sg13g2_nand4_1 _21235_ (.B(_03619_),
    .C(_03622_),
    .A(_03594_),
    .Y(_03636_),
    .D(_03635_));
 sg13g2_nor2_2 _21236_ (.A(_03629_),
    .B(_03631_),
    .Y(_03637_));
 sg13g2_nor2_1 _21237_ (.A(net242),
    .B(_03637_),
    .Y(_03638_));
 sg13g2_o21ai_1 _21238_ (.B1(_11372_),
    .Y(_03639_),
    .A1(_03625_),
    .A2(_03626_));
 sg13g2_buf_1 _21239_ (.A(_03639_),
    .X(_03640_));
 sg13g2_buf_8 _21240_ (.A(_03624_),
    .X(_03641_));
 sg13g2_a221oi_1 _21241_ (.B2(net160),
    .C1(_10522_),
    .B1(_03640_),
    .A1(net242),
    .Y(_03642_),
    .A2(_03637_));
 sg13g2_nor3_1 _21242_ (.A(net160),
    .B(_03632_),
    .C(_03640_),
    .Y(_03643_));
 sg13g2_nor3_1 _21243_ (.A(_03638_),
    .B(_03642_),
    .C(_03643_),
    .Y(_03644_));
 sg13g2_nand2b_1 _21244_ (.Y(_03645_),
    .B(_11245_),
    .A_N(_03644_));
 sg13g2_a21oi_1 _21245_ (.A1(net277),
    .A2(_03610_),
    .Y(_03646_),
    .B1(_03622_));
 sg13g2_nand4_1 _21246_ (.B(_03608_),
    .C(_03617_),
    .A(_03600_),
    .Y(_03647_),
    .D(_03646_));
 sg13g2_mux2_1 _21247_ (.A0(_10679_),
    .A1(_11277_),
    .S(net241),
    .X(_03648_));
 sg13g2_buf_2 _21248_ (.A(_03648_),
    .X(_03649_));
 sg13g2_nand3_1 _21249_ (.B(_03593_),
    .C(_03649_),
    .A(_03578_),
    .Y(_03650_));
 sg13g2_inv_1 _21250_ (.Y(_03651_),
    .A(_11245_));
 sg13g2_nor2_1 _21251_ (.A(net232),
    .B(_03651_),
    .Y(_03652_));
 sg13g2_nand4_1 _21252_ (.B(_03650_),
    .C(_03634_),
    .A(_03647_),
    .Y(_03653_),
    .D(_03652_));
 sg13g2_and4_1 _21253_ (.A(net221),
    .B(_03636_),
    .C(_03645_),
    .D(_03653_),
    .X(_03654_));
 sg13g2_nand4_1 _21254_ (.B(_03647_),
    .C(_03650_),
    .A(_11589_),
    .Y(_03655_),
    .D(_03634_));
 sg13g2_nand4_1 _21255_ (.B(_03619_),
    .C(_03622_),
    .A(_03594_),
    .Y(_03656_),
    .D(_03634_));
 sg13g2_and4_1 _21256_ (.A(_03651_),
    .B(_03655_),
    .C(_03644_),
    .D(_03656_),
    .X(_03657_));
 sg13g2_nand2_1 _21257_ (.Y(_03658_),
    .A(net215),
    .B(_03570_));
 sg13g2_o21ai_1 _21258_ (.B1(_03658_),
    .Y(_03659_),
    .A1(_03654_),
    .A2(_03657_));
 sg13g2_mux2_1 _21259_ (.A0(_11093_),
    .A1(_11164_),
    .S(net209),
    .X(_03660_));
 sg13g2_buf_1 _21260_ (.A(_03660_),
    .X(_03661_));
 sg13g2_buf_1 _21261_ (.A(_03661_),
    .X(_03662_));
 sg13g2_nand2_1 _21262_ (.Y(_03663_),
    .A(net168),
    .B(_03662_));
 sg13g2_nor2_1 _21263_ (.A(_00186_),
    .B(net209),
    .Y(_03664_));
 sg13g2_a21oi_1 _21264_ (.A1(_03568_),
    .A2(_11137_),
    .Y(_03665_),
    .B1(_03664_));
 sg13g2_buf_2 _21265_ (.A(_03665_),
    .X(_03666_));
 sg13g2_nand2_1 _21266_ (.Y(_03667_),
    .A(net209),
    .B(_11184_));
 sg13g2_o21ai_1 _21267_ (.B1(_03667_),
    .Y(_03668_),
    .A1(_10296_),
    .A2(net209));
 sg13g2_buf_1 _21268_ (.A(_03668_),
    .X(_03669_));
 sg13g2_buf_1 _21269_ (.A(_03669_),
    .X(_03670_));
 sg13g2_nand2_1 _21270_ (.Y(_03671_),
    .A(_11430_),
    .B(net122));
 sg13g2_nand3_1 _21271_ (.B(_03666_),
    .C(_03671_),
    .A(_03663_),
    .Y(_03672_));
 sg13g2_nand3_1 _21272_ (.B(_03663_),
    .C(_03671_),
    .A(net197),
    .Y(_03673_));
 sg13g2_a22oi_1 _21273_ (.Y(_03674_),
    .B1(_03672_),
    .B2(_03673_),
    .A2(_03659_),
    .A1(_03572_));
 sg13g2_inv_1 _21274_ (.Y(_03675_),
    .A(_03661_));
 sg13g2_nor2_1 _21275_ (.A(net201),
    .B(_03675_),
    .Y(_03676_));
 sg13g2_nand2_2 _21276_ (.Y(_03677_),
    .A(net197),
    .B(_03666_));
 sg13g2_nand2b_1 _21277_ (.Y(_03678_),
    .B(net144),
    .A_N(_03669_));
 sg13g2_buf_1 _21278_ (.A(_03678_),
    .X(_03679_));
 sg13g2_nor2_1 _21279_ (.A(_03676_),
    .B(_03679_),
    .Y(_03680_));
 sg13g2_o21ai_1 _21280_ (.B1(_03680_),
    .Y(_03681_),
    .A1(net197),
    .A2(_03666_));
 sg13g2_o21ai_1 _21281_ (.B1(_03681_),
    .Y(_03682_),
    .A1(_03676_),
    .A2(_03677_));
 sg13g2_nor2_1 _21282_ (.A(net168),
    .B(_03661_),
    .Y(_03683_));
 sg13g2_nor3_1 _21283_ (.A(_03674_),
    .B(_03682_),
    .C(_03683_),
    .Y(_03684_));
 sg13g2_a21o_1 _21284_ (.A2(_03684_),
    .A1(net161),
    .B1(_11875_),
    .X(_03685_));
 sg13g2_or2_1 _21285_ (.X(_03686_),
    .B(_03684_),
    .A(net161));
 sg13g2_nand4_1 _21286_ (.B(_03557_),
    .C(_03685_),
    .A(net948),
    .Y(_03687_),
    .D(_03686_));
 sg13g2_o21ai_1 _21287_ (.B1(_03687_),
    .Y(_03688_),
    .A1(\cpu.ex.r_cc ),
    .A2(_03557_));
 sg13g2_buf_1 _21288_ (.A(net141),
    .X(_03689_));
 sg13g2_buf_1 _21289_ (.A(_03555_),
    .X(_03690_));
 sg13g2_buf_1 _21290_ (.A(net76),
    .X(_03691_));
 sg13g2_or2_1 _21291_ (.X(_03692_),
    .B(net161),
    .A(net167));
 sg13g2_nand2_1 _21292_ (.Y(_03693_),
    .A(net215),
    .B(_03571_));
 sg13g2_buf_1 _21293_ (.A(_03693_),
    .X(_03694_));
 sg13g2_nand3_1 _21294_ (.B(net122),
    .C(_03694_),
    .A(net200),
    .Y(_03695_));
 sg13g2_buf_1 _21295_ (.A(_11245_),
    .X(_03696_));
 sg13g2_nand3_1 _21296_ (.B(_03669_),
    .C(_03694_),
    .A(net192),
    .Y(_03697_));
 sg13g2_nand3_1 _21297_ (.B(_03580_),
    .C(_03582_),
    .A(_10842_),
    .Y(_03698_));
 sg13g2_buf_1 _21298_ (.A(_03698_),
    .X(_03699_));
 sg13g2_o21ai_1 _21299_ (.B1(net282),
    .Y(_03700_),
    .A1(_03577_),
    .A2(_03699_));
 sg13g2_nand2_1 _21300_ (.Y(_03701_),
    .A(_03577_),
    .B(_03699_));
 sg13g2_nand2_1 _21301_ (.Y(_03702_),
    .A(_03700_),
    .B(_03701_));
 sg13g2_a22oi_1 _21302_ (.Y(_03703_),
    .B1(_11925_),
    .B2(net282),
    .A2(_03581_),
    .A1(net281));
 sg13g2_a21oi_1 _21303_ (.A1(_10742_),
    .A2(_10765_),
    .Y(_03704_),
    .B1(_00280_));
 sg13g2_a21oi_1 _21304_ (.A1(_10790_),
    .A2(_10796_),
    .Y(_03705_),
    .B1(_08498_));
 sg13g2_nor4_1 _21305_ (.A(_11053_),
    .B(net351),
    .C(_03704_),
    .D(_03705_),
    .Y(_03706_));
 sg13g2_a21o_1 _21306_ (.A2(_03703_),
    .A1(net241),
    .B1(_03706_),
    .X(_03707_));
 sg13g2_buf_1 _21307_ (.A(_03707_),
    .X(_03708_));
 sg13g2_nand3_1 _21308_ (.B(_03596_),
    .C(_03597_),
    .A(net286),
    .Y(_03709_));
 sg13g2_buf_2 _21309_ (.A(_03709_),
    .X(_03710_));
 sg13g2_nor2_1 _21310_ (.A(net208),
    .B(_03710_),
    .Y(_03711_));
 sg13g2_a22oi_1 _21311_ (.Y(_03712_),
    .B1(net513),
    .B2(_10578_),
    .A2(net569),
    .A1(_09231_));
 sg13g2_o21ai_1 _21312_ (.B1(_10205_),
    .Y(_03713_),
    .A1(_10583_),
    .A2(_10290_));
 sg13g2_a21o_1 _21313_ (.A2(_03712_),
    .A1(net1047),
    .B1(_03713_),
    .X(_03714_));
 sg13g2_nand2b_1 _21314_ (.Y(_03715_),
    .B(net1046),
    .A_N(_10582_));
 sg13g2_nand2_1 _21315_ (.Y(_03716_),
    .A(_10950_),
    .B(_10951_));
 sg13g2_a221oi_1 _21316_ (.B2(net1117),
    .C1(_03716_),
    .B1(net350),
    .A1(_03714_),
    .Y(_03717_),
    .A2(_03715_));
 sg13g2_buf_2 _21317_ (.A(_03717_),
    .X(_03718_));
 sg13g2_nor4_2 _21318_ (.A(net758),
    .B(_10582_),
    .C(_10588_),
    .Y(_03719_),
    .D(net351));
 sg13g2_a21oi_1 _21319_ (.A1(net241),
    .A2(_03703_),
    .Y(_03720_),
    .B1(_03706_));
 sg13g2_nor4_1 _21320_ (.A(_03615_),
    .B(_03718_),
    .C(_03719_),
    .D(_03720_),
    .Y(_03721_));
 sg13g2_nor3_2 _21321_ (.A(net890),
    .B(_10643_),
    .C(_03559_),
    .Y(_03722_));
 sg13g2_a21oi_1 _21322_ (.A1(_11043_),
    .A2(_11048_),
    .Y(_03723_),
    .B1(_11037_));
 sg13g2_nor3_1 _21323_ (.A(net280),
    .B(_03722_),
    .C(_03723_),
    .Y(_03724_));
 sg13g2_nand2_1 _21324_ (.Y(_03725_),
    .A(_11072_),
    .B(_11074_));
 sg13g2_nand2b_1 _21325_ (.Y(_03726_),
    .B(_11072_),
    .A_N(_11054_));
 sg13g2_mux2_1 _21326_ (.A0(_03725_),
    .A1(_03726_),
    .S(_08470_),
    .X(_03727_));
 sg13g2_buf_1 _21327_ (.A(_03727_),
    .X(_03728_));
 sg13g2_nor2_1 _21328_ (.A(net284),
    .B(_11037_),
    .Y(_03729_));
 sg13g2_nor4_1 _21329_ (.A(net890),
    .B(_10643_),
    .C(net284),
    .D(_03559_),
    .Y(_03730_));
 sg13g2_a221oi_1 _21330_ (.B2(net241),
    .C1(_03730_),
    .B1(_03729_),
    .A1(_10869_),
    .Y(_03731_),
    .A2(_03728_));
 sg13g2_or2_1 _21331_ (.X(_03732_),
    .B(_03731_),
    .A(_03724_));
 sg13g2_buf_1 _21332_ (.A(_03732_),
    .X(_03733_));
 sg13g2_nor3_1 _21333_ (.A(net237),
    .B(_03710_),
    .C(_03720_),
    .Y(_03734_));
 sg13g2_a221oi_1 _21334_ (.B2(_03733_),
    .C1(_03734_),
    .B1(_03721_),
    .A1(_03708_),
    .Y(_03735_),
    .A2(_03711_));
 sg13g2_nor2_1 _21335_ (.A(net237),
    .B(net208),
    .Y(_03736_));
 sg13g2_nor4_1 _21336_ (.A(net237),
    .B(_03718_),
    .C(_03719_),
    .D(_03720_),
    .Y(_03737_));
 sg13g2_a22oi_1 _21337_ (.Y(_03738_),
    .B1(_03737_),
    .B2(_03733_),
    .A2(_03736_),
    .A1(_03708_));
 sg13g2_a21oi_1 _21338_ (.A1(net234),
    .A2(_03628_),
    .Y(_03739_),
    .B1(_03649_));
 sg13g2_nand4_1 _21339_ (.B(_03735_),
    .C(_03738_),
    .A(_03702_),
    .Y(_03740_),
    .D(_03739_));
 sg13g2_buf_1 _21340_ (.A(_03740_),
    .X(_03741_));
 sg13g2_or2_1 _21341_ (.X(_03742_),
    .B(_03626_),
    .A(_03625_));
 sg13g2_buf_1 _21342_ (.A(_03742_),
    .X(_03743_));
 sg13g2_nand2_2 _21343_ (.Y(_03744_),
    .A(net233),
    .B(_03743_));
 sg13g2_nor2_1 _21344_ (.A(_03718_),
    .B(_03719_),
    .Y(_03745_));
 sg13g2_o21ai_1 _21345_ (.B1(_03745_),
    .Y(_03746_),
    .A1(_03724_),
    .A2(_03731_));
 sg13g2_buf_1 _21346_ (.A(_03746_),
    .X(_03747_));
 sg13g2_o21ai_1 _21347_ (.B1(net237),
    .Y(_03748_),
    .A1(_03612_),
    .A2(_03613_));
 sg13g2_nand3_1 _21348_ (.B(_03708_),
    .C(_03748_),
    .A(_03649_),
    .Y(_03749_));
 sg13g2_a21o_1 _21349_ (.A2(_03710_),
    .A1(_03747_),
    .B1(_03749_),
    .X(_03750_));
 sg13g2_buf_1 _21350_ (.A(_03750_),
    .X(_03751_));
 sg13g2_nand2_1 _21351_ (.Y(_03752_),
    .A(net282),
    .B(_11925_));
 sg13g2_nand2_1 _21352_ (.Y(_03753_),
    .A(_10740_),
    .B(_10767_));
 sg13g2_mux2_1 _21353_ (.A0(_03752_),
    .A1(_03753_),
    .S(_03561_),
    .X(_03754_));
 sg13g2_and2_1 _21354_ (.A(_03649_),
    .B(_03754_),
    .X(_03755_));
 sg13g2_a21oi_1 _21355_ (.A1(net285),
    .A2(_11922_),
    .Y(_03756_),
    .B1(_11297_));
 sg13g2_a21oi_1 _21356_ (.A1(_10612_),
    .A2(net285),
    .Y(_03757_),
    .B1(_08533_));
 sg13g2_mux2_1 _21357_ (.A0(_03756_),
    .A1(_03757_),
    .S(_03561_),
    .X(_03758_));
 sg13g2_nor2_1 _21358_ (.A(_10864_),
    .B(_11923_),
    .Y(_03759_));
 sg13g2_and4_1 _21359_ (.A(_11477_),
    .B(net285),
    .C(_03562_),
    .D(_03589_),
    .X(_03760_));
 sg13g2_a221oi_1 _21360_ (.B2(_03759_),
    .C1(_03760_),
    .B1(_11186_),
    .A1(_10790_),
    .Y(_03761_),
    .A2(_10796_));
 sg13g2_nand3_1 _21361_ (.B(_03574_),
    .C(_03575_),
    .A(_10839_),
    .Y(_03762_));
 sg13g2_o21ai_1 _21362_ (.B1(_03762_),
    .Y(_03763_),
    .A1(_03758_),
    .A2(_03761_));
 sg13g2_a221oi_1 _21363_ (.B2(_03763_),
    .C1(net361),
    .B1(_03755_),
    .A1(net234),
    .Y(_03764_),
    .A2(_03628_));
 sg13g2_buf_1 _21364_ (.A(_03764_),
    .X(_03765_));
 sg13g2_a21o_1 _21365_ (.A2(_11320_),
    .A1(net209),
    .B1(_03623_),
    .X(_03766_));
 sg13g2_buf_1 _21366_ (.A(_03766_),
    .X(_03767_));
 sg13g2_a21oi_1 _21367_ (.A1(_03751_),
    .A2(_03765_),
    .Y(_03768_),
    .B1(_03767_));
 sg13g2_or2_1 _21368_ (.X(_03769_),
    .B(_03631_),
    .A(_03629_));
 sg13g2_buf_2 _21369_ (.A(_03769_),
    .X(_03770_));
 sg13g2_nand2_1 _21370_ (.Y(_03771_),
    .A(net220),
    .B(_03770_));
 sg13g2_nand4_1 _21371_ (.B(_03744_),
    .C(_03768_),
    .A(_03741_),
    .Y(_03772_),
    .D(_03771_));
 sg13g2_nand2_1 _21372_ (.Y(_03773_),
    .A(_03751_),
    .B(_03765_));
 sg13g2_nor2_1 _21373_ (.A(net169),
    .B(_03770_),
    .Y(_03774_));
 sg13g2_nand4_1 _21374_ (.B(_03741_),
    .C(_03744_),
    .A(_03773_),
    .Y(_03775_),
    .D(_03774_));
 sg13g2_nand4_1 _21375_ (.B(_03773_),
    .C(_03741_),
    .A(_11707_),
    .Y(_03776_),
    .D(_03744_));
 sg13g2_nor3_1 _21376_ (.A(net169),
    .B(_03767_),
    .C(_03770_),
    .Y(_03777_));
 sg13g2_a221oi_1 _21377_ (.B2(_11669_),
    .C1(_03777_),
    .B1(_03637_),
    .A1(_11707_),
    .Y(_03778_),
    .A2(net160));
 sg13g2_nand4_1 _21378_ (.B(_03775_),
    .C(_03776_),
    .A(_03772_),
    .Y(_03779_),
    .D(_03778_));
 sg13g2_buf_1 _21379_ (.A(_03779_),
    .X(_03780_));
 sg13g2_a21o_1 _21380_ (.A2(_03697_),
    .A1(_03695_),
    .B1(_03780_),
    .X(_03781_));
 sg13g2_buf_1 _21381_ (.A(_03781_),
    .X(_03782_));
 sg13g2_nor2_1 _21382_ (.A(_11767_),
    .B(_03571_),
    .Y(_03783_));
 sg13g2_buf_1 _21383_ (.A(_03783_),
    .X(_03784_));
 sg13g2_and3_1 _21384_ (.X(_03785_),
    .A(_11245_),
    .B(_03669_),
    .C(_03694_));
 sg13g2_a221oi_1 _21385_ (.B2(net200),
    .C1(net144),
    .B1(_03785_),
    .A1(net122),
    .Y(_03786_),
    .A2(_03784_));
 sg13g2_buf_1 _21386_ (.A(_03786_),
    .X(_03787_));
 sg13g2_nor2_1 _21387_ (.A(_03651_),
    .B(_11401_),
    .Y(_03788_));
 sg13g2_nor2_1 _21388_ (.A(_11245_),
    .B(_10422_),
    .Y(_03789_));
 sg13g2_inv_1 _21389_ (.Y(_03790_),
    .A(_03789_));
 sg13g2_and3_1 _21390_ (.X(_03791_),
    .A(_03772_),
    .B(_03790_),
    .C(_03694_));
 sg13g2_nor2_1 _21391_ (.A(_11669_),
    .B(_03777_),
    .Y(_03792_));
 sg13g2_buf_1 _21392_ (.A(_03743_),
    .X(_03793_));
 sg13g2_a221oi_1 _21393_ (.B2(_03765_),
    .C1(net169),
    .B1(_03751_),
    .A1(net233),
    .Y(_03794_),
    .A2(net191));
 sg13g2_a221oi_1 _21394_ (.B2(_03794_),
    .C1(_03637_),
    .B1(_03741_),
    .A1(net216),
    .Y(_03795_),
    .A2(net160));
 sg13g2_a21o_1 _21395_ (.A2(_03792_),
    .A1(_03775_),
    .B1(_03795_),
    .X(_03796_));
 sg13g2_a22oi_1 _21396_ (.Y(_03797_),
    .B1(_03791_),
    .B2(_03796_),
    .A2(_03694_),
    .A1(_03788_));
 sg13g2_buf_1 _21397_ (.A(_03797_),
    .X(_03798_));
 sg13g2_buf_1 _21398_ (.A(_03670_),
    .X(_03799_));
 sg13g2_nor2_1 _21399_ (.A(net107),
    .B(_03784_),
    .Y(_03800_));
 sg13g2_buf_1 _21400_ (.A(net140),
    .X(_03801_));
 sg13g2_a21o_1 _21401_ (.A2(_11137_),
    .A1(net209),
    .B1(_03664_),
    .X(_03802_));
 sg13g2_buf_1 _21402_ (.A(_03802_),
    .X(_03803_));
 sg13g2_buf_1 _21403_ (.A(_03803_),
    .X(_03804_));
 sg13g2_nand2_1 _21404_ (.Y(_03805_),
    .A(_03801_),
    .B(_03804_));
 sg13g2_a221oi_1 _21405_ (.B2(_03800_),
    .C1(_03805_),
    .B1(_03798_),
    .A1(_03782_),
    .Y(_03806_),
    .A2(_03787_));
 sg13g2_nand2_1 _21406_ (.Y(_03807_),
    .A(_11795_),
    .B(net120));
 sg13g2_a221oi_1 _21407_ (.B2(_03800_),
    .C1(_03807_),
    .B1(_03798_),
    .A1(_03782_),
    .Y(_03808_),
    .A2(_03787_));
 sg13g2_nor2_1 _21408_ (.A(_03666_),
    .B(_03807_),
    .Y(_03809_));
 sg13g2_nor4_2 _21409_ (.A(net201),
    .B(_03806_),
    .C(_03808_),
    .Y(_03810_),
    .D(_03809_));
 sg13g2_nand2_1 _21410_ (.Y(_03811_),
    .A(_11428_),
    .B(_03666_));
 sg13g2_inv_1 _21411_ (.Y(_03812_),
    .A(_03811_));
 sg13g2_a221oi_1 _21412_ (.B2(_03800_),
    .C1(_03812_),
    .B1(_03798_),
    .A1(_03782_),
    .Y(_03813_),
    .A2(_03787_));
 sg13g2_buf_1 _21413_ (.A(_03813_),
    .X(_03814_));
 sg13g2_nor2_2 _21414_ (.A(_11428_),
    .B(_03666_),
    .Y(_03815_));
 sg13g2_nor3_1 _21415_ (.A(net120),
    .B(_03814_),
    .C(_03815_),
    .Y(_03816_));
 sg13g2_nand2_1 _21416_ (.Y(_03817_),
    .A(net167),
    .B(net193));
 sg13g2_o21ai_1 _21417_ (.B1(_03817_),
    .Y(_03818_),
    .A1(_03810_),
    .A2(_03816_));
 sg13g2_a221oi_1 _21418_ (.B2(_03818_),
    .C1(net948),
    .B1(_03692_),
    .A1(net121),
    .Y(_03819_),
    .A2(net36));
 sg13g2_nor2_1 _21419_ (.A(_03688_),
    .B(_03819_),
    .Y(_00916_));
 sg13g2_or4_1 _21420_ (.A(net1126),
    .B(net1052),
    .C(_10189_),
    .D(_10197_),
    .X(_03820_));
 sg13g2_nor2_1 _21421_ (.A(_08348_),
    .B(_03820_),
    .Y(_03821_));
 sg13g2_buf_2 _21422_ (.A(_03821_),
    .X(_03822_));
 sg13g2_buf_1 _21423_ (.A(_03822_),
    .X(_03823_));
 sg13g2_mux2_1 _21424_ (.A0(\cpu.ex.r_epc[1] ),
    .A1(net492),
    .S(net604),
    .X(_00918_));
 sg13g2_mux2_1 _21425_ (.A0(\cpu.ex.r_epc[11] ),
    .A1(_03011_),
    .S(net604),
    .X(_00919_));
 sg13g2_mux2_1 _21426_ (.A0(\cpu.ex.r_epc[12] ),
    .A1(net542),
    .S(net604),
    .X(_00920_));
 sg13g2_mux2_1 _21427_ (.A0(\cpu.ex.r_epc[13] ),
    .A1(net489),
    .S(net604),
    .X(_00921_));
 sg13g2_mux2_1 _21428_ (.A0(\cpu.ex.r_epc[14] ),
    .A1(_03504_),
    .S(net604),
    .X(_00922_));
 sg13g2_mux2_1 _21429_ (.A0(\cpu.ex.r_epc[15] ),
    .A1(net746),
    .S(net604),
    .X(_00923_));
 sg13g2_mux2_1 _21430_ (.A0(\cpu.ex.r_epc[2] ),
    .A1(net453),
    .S(net604),
    .X(_00924_));
 sg13g2_mux2_1 _21431_ (.A0(\cpu.ex.r_epc[3] ),
    .A1(net410),
    .S(_03823_),
    .X(_00925_));
 sg13g2_mux2_1 _21432_ (.A0(\cpu.ex.r_epc[4] ),
    .A1(net409),
    .S(_03823_),
    .X(_00926_));
 sg13g2_mux2_1 _21433_ (.A0(\cpu.ex.r_epc[5] ),
    .A1(net667),
    .S(net604),
    .X(_00927_));
 sg13g2_mux2_1 _21434_ (.A0(\cpu.ex.r_epc[6] ),
    .A1(net747),
    .S(_03822_),
    .X(_00928_));
 sg13g2_mux2_1 _21435_ (.A0(\cpu.ex.r_epc[7] ),
    .A1(net992),
    .S(_03822_),
    .X(_00929_));
 sg13g2_mux2_1 _21436_ (.A0(\cpu.ex.r_epc[8] ),
    .A1(net857),
    .S(_03822_),
    .X(_00930_));
 sg13g2_mux2_1 _21437_ (.A0(\cpu.ex.r_epc[9] ),
    .A1(net859),
    .S(_03822_),
    .X(_00931_));
 sg13g2_mux2_1 _21438_ (.A0(\cpu.ex.r_epc[10] ),
    .A1(net858),
    .S(_03822_),
    .X(_00932_));
 sg13g2_or4_1 _21439_ (.A(net1126),
    .B(_10192_),
    .C(_10189_),
    .D(_03526_),
    .X(_03824_));
 sg13g2_buf_1 _21440_ (.A(_03824_),
    .X(_03825_));
 sg13g2_buf_1 _21441_ (.A(_03825_),
    .X(_03826_));
 sg13g2_buf_1 _21442_ (.A(_03825_),
    .X(_03827_));
 sg13g2_nand2_1 _21443_ (.Y(_03828_),
    .A(\cpu.ex.r_lr[1] ),
    .B(net602));
 sg13g2_o21ai_1 _21444_ (.B1(_03828_),
    .Y(_00938_),
    .A1(net622),
    .A2(net603));
 sg13g2_mux2_1 _21445_ (.A0(_02974_),
    .A1(\cpu.ex.r_lr[11] ),
    .S(net602),
    .X(_00939_));
 sg13g2_buf_1 _21446_ (.A(net552),
    .X(_03829_));
 sg13g2_mux2_1 _21447_ (.A0(net488),
    .A1(\cpu.ex.r_lr[12] ),
    .S(_03827_),
    .X(_00940_));
 sg13g2_buf_1 _21448_ (.A(net493),
    .X(_03830_));
 sg13g2_mux2_1 _21449_ (.A0(net451),
    .A1(\cpu.ex.r_lr[13] ),
    .S(_03827_),
    .X(_00941_));
 sg13g2_buf_1 _21450_ (.A(net605),
    .X(_03831_));
 sg13g2_mux2_1 _21451_ (.A0(net541),
    .A1(\cpu.ex.r_lr[14] ),
    .S(net602),
    .X(_00942_));
 sg13g2_buf_1 _21452_ (.A(net699),
    .X(_03832_));
 sg13g2_nand2_1 _21453_ (.Y(_03833_),
    .A(\cpu.ex.r_lr[15] ),
    .B(net602));
 sg13g2_o21ai_1 _21454_ (.B1(_03833_),
    .Y(_00943_),
    .A1(_03832_),
    .A2(net603));
 sg13g2_buf_1 _21455_ (.A(net694),
    .X(_03834_));
 sg13g2_buf_1 _21456_ (.A(net600),
    .X(_03835_));
 sg13g2_nand2_1 _21457_ (.Y(_03836_),
    .A(\cpu.ex.r_lr[2] ),
    .B(net602));
 sg13g2_o21ai_1 _21458_ (.B1(_03836_),
    .Y(_00944_),
    .A1(_03835_),
    .A2(net603));
 sg13g2_nand2_1 _21459_ (.Y(_03837_),
    .A(\cpu.ex.r_lr[3] ),
    .B(net602));
 sg13g2_o21ai_1 _21460_ (.B1(_03837_),
    .Y(_00945_),
    .A1(net926),
    .A2(net603));
 sg13g2_buf_1 _21461_ (.A(_09810_),
    .X(_03838_));
 sg13g2_buf_1 _21462_ (.A(net666),
    .X(_03839_));
 sg13g2_nand2_1 _21463_ (.Y(_03840_),
    .A(\cpu.ex.r_lr[4] ),
    .B(net602));
 sg13g2_o21ai_1 _21464_ (.B1(_03840_),
    .Y(_00946_),
    .A1(net599),
    .A2(net603));
 sg13g2_nand2_1 _21465_ (.Y(_03841_),
    .A(\cpu.ex.r_lr[5] ),
    .B(_03825_));
 sg13g2_o21ai_1 _21466_ (.B1(_03841_),
    .Y(_00947_),
    .A1(net754),
    .A2(net603));
 sg13g2_mux2_1 _21467_ (.A0(net753),
    .A1(\cpu.ex.r_lr[6] ),
    .S(net602),
    .X(_00948_));
 sg13g2_nand2_1 _21468_ (.Y(_03842_),
    .A(\cpu.ex.r_lr[7] ),
    .B(_03825_));
 sg13g2_o21ai_1 _21469_ (.B1(_03842_),
    .Y(_00949_),
    .A1(net752),
    .A2(net603));
 sg13g2_nand2_1 _21470_ (.Y(_03843_),
    .A(\cpu.ex.r_lr[8] ),
    .B(_03825_));
 sg13g2_o21ai_1 _21471_ (.B1(_03843_),
    .Y(_00950_),
    .A1(net870),
    .A2(net603));
 sg13g2_nand2_1 _21472_ (.Y(_03844_),
    .A(\cpu.ex.r_lr[9] ),
    .B(_03825_));
 sg13g2_o21ai_1 _21473_ (.B1(_03844_),
    .Y(_00951_),
    .A1(net751),
    .A2(_03826_));
 sg13g2_nand2_1 _21474_ (.Y(_03845_),
    .A(\cpu.ex.r_lr[10] ),
    .B(_03825_));
 sg13g2_o21ai_1 _21475_ (.B1(_03845_),
    .Y(_00952_),
    .A1(_02971_),
    .A2(_03826_));
 sg13g2_nor2_1 _21476_ (.A(_11843_),
    .B(_11867_),
    .Y(_03846_));
 sg13g2_a21oi_1 _21477_ (.A1(_11843_),
    .A2(_11867_),
    .Y(_03847_),
    .B1(net168));
 sg13g2_nor2_1 _21478_ (.A(_03846_),
    .B(_03847_),
    .Y(_03848_));
 sg13g2_nand3_1 _21479_ (.B(net510),
    .C(_10455_),
    .A(_11906_),
    .Y(_03849_));
 sg13g2_a21oi_1 _21480_ (.A1(_03848_),
    .A2(_03849_),
    .Y(_03850_),
    .B1(net109));
 sg13g2_nand2_1 _21481_ (.Y(_03851_),
    .A(_11900_),
    .B(_11875_));
 sg13g2_nand2_1 _21482_ (.Y(_03852_),
    .A(_11910_),
    .B(net510));
 sg13g2_a21oi_1 _21483_ (.A1(_03850_),
    .A2(_03851_),
    .Y(_03853_),
    .B1(_03852_));
 sg13g2_and2_1 _21484_ (.A(net167),
    .B(_03852_),
    .X(_03854_));
 sg13g2_nor3_1 _21485_ (.A(_11900_),
    .B(_11910_),
    .C(net564),
    .Y(_03855_));
 sg13g2_o21ai_1 _21486_ (.B1(_03850_),
    .Y(_03856_),
    .A1(_03854_),
    .A2(_03855_));
 sg13g2_nor2b_1 _21487_ (.A(_03853_),
    .B_N(_03856_),
    .Y(_03857_));
 sg13g2_nor3_1 _21488_ (.A(_10189_),
    .B(_10194_),
    .C(_10197_),
    .Y(_03858_));
 sg13g2_buf_1 _21489_ (.A(_03858_),
    .X(_03859_));
 sg13g2_buf_1 _21490_ (.A(net598),
    .X(_03860_));
 sg13g2_buf_8 _21491_ (.A(_11425_),
    .X(_03861_));
 sg13g2_buf_1 _21492_ (.A(_11444_),
    .X(_03862_));
 sg13g2_nor3_1 _21493_ (.A(net198),
    .B(net28),
    .C(net32),
    .Y(_03863_));
 sg13g2_xnor2_1 _21494_ (.Y(_03864_),
    .A(net109),
    .B(_03863_));
 sg13g2_nand3_1 _21495_ (.B(_10200_),
    .C(\cpu.ex.r_cc ),
    .A(net1127),
    .Y(_03865_));
 sg13g2_nand3_1 _21496_ (.B(_10201_),
    .C(_11459_),
    .A(\cpu.ex.r_mult[16] ),
    .Y(_03866_));
 sg13g2_a21oi_1 _21497_ (.A1(_03865_),
    .A2(_03866_),
    .Y(_03867_),
    .B1(_03859_));
 sg13g2_a221oi_1 _21498_ (.B2(_03864_),
    .C1(_03867_),
    .B1(_11793_),
    .A1(_03490_),
    .Y(_03868_),
    .A2(net539));
 sg13g2_o21ai_1 _21499_ (.B1(_03868_),
    .Y(_00953_),
    .A1(_11786_),
    .A2(_03857_));
 sg13g2_nand2_1 _21500_ (.Y(_03869_),
    .A(_11416_),
    .B(_11843_));
 sg13g2_a21oi_1 _21501_ (.A1(_10455_),
    .A2(_03869_),
    .Y(_03870_),
    .B1(_11906_));
 sg13g2_nor2_1 _21502_ (.A(_10455_),
    .B(_03869_),
    .Y(_03871_));
 sg13g2_nor2_1 _21503_ (.A(_11900_),
    .B(_11843_),
    .Y(_03872_));
 sg13g2_nor2_1 _21504_ (.A(net123),
    .B(_03872_),
    .Y(_03873_));
 sg13g2_nor4_2 _21505_ (.A(_03852_),
    .B(_03870_),
    .C(_03871_),
    .Y(_03874_),
    .D(_03873_));
 sg13g2_o21ai_1 _21506_ (.B1(_03869_),
    .Y(_03875_),
    .A1(_11866_),
    .A2(_11890_));
 sg13g2_nand4_1 _21507_ (.B(net510),
    .C(net123),
    .A(_11910_),
    .Y(_03876_),
    .D(_03851_));
 sg13g2_a21oi_1 _21508_ (.A1(_03849_),
    .A2(_03875_),
    .Y(_03877_),
    .B1(_03876_));
 sg13g2_a21oi_2 _21509_ (.B1(_03877_),
    .Y(_03878_),
    .A2(_03874_),
    .A1(_11855_));
 sg13g2_nor2_1 _21510_ (.A(_10847_),
    .B(net564),
    .Y(_03879_));
 sg13g2_xnor2_1 _21511_ (.Y(_03880_),
    .A(_03878_),
    .B(_03879_));
 sg13g2_nand2_2 _21512_ (.Y(_03881_),
    .A(_10201_),
    .B(_11459_));
 sg13g2_nand4_1 _21513_ (.B(net1127),
    .C(_10200_),
    .A(_08335_),
    .Y(_03882_),
    .D(\cpu.ex.r_cc ));
 sg13g2_a21oi_1 _21514_ (.A1(_03881_),
    .A2(_03882_),
    .Y(_03883_),
    .B1(_03859_));
 sg13g2_buf_1 _21515_ (.A(_03883_),
    .X(_03884_));
 sg13g2_buf_1 _21516_ (.A(_03884_),
    .X(_03885_));
 sg13g2_a221oi_1 _21517_ (.B2(_03880_),
    .C1(net271),
    .B1(_11722_),
    .A1(net550),
    .Y(_03886_),
    .A2(net539));
 sg13g2_buf_1 _21518_ (.A(_11793_),
    .X(_03887_));
 sg13g2_buf_1 _21519_ (.A(net280),
    .X(_03888_));
 sg13g2_buf_1 _21520_ (.A(net227),
    .X(_03889_));
 sg13g2_nor2_1 _21521_ (.A(net198),
    .B(net98),
    .Y(_03890_));
 sg13g2_xnor2_1 _21522_ (.Y(_03891_),
    .A(net207),
    .B(_03890_));
 sg13g2_nor3_1 _21523_ (.A(_03861_),
    .B(_03862_),
    .C(_03891_),
    .Y(_03892_));
 sg13g2_xnor2_1 _21524_ (.Y(_03893_),
    .A(_10862_),
    .B(_03892_));
 sg13g2_nand2_1 _21525_ (.Y(_03894_),
    .A(net31),
    .B(_03893_));
 sg13g2_nand2_1 _21526_ (.Y(_03895_),
    .A(net461),
    .B(_11459_));
 sg13g2_buf_1 _21527_ (.A(_03895_),
    .X(_03896_));
 sg13g2_nor2_1 _21528_ (.A(\cpu.ex.r_mult[17] ),
    .B(net349),
    .Y(_03897_));
 sg13g2_a21oi_1 _21529_ (.A1(_03886_),
    .A2(_03894_),
    .Y(_00954_),
    .B1(_03897_));
 sg13g2_nor2_1 _21530_ (.A(_10870_),
    .B(net98),
    .Y(_03898_));
 sg13g2_a21oi_1 _21531_ (.A1(net207),
    .A2(_10862_),
    .Y(_03899_),
    .B1(_03898_));
 sg13g2_xnor2_1 _21532_ (.Y(_03900_),
    .A(net286),
    .B(_03899_));
 sg13g2_nor3_1 _21533_ (.A(_03861_),
    .B(_03862_),
    .C(_03900_),
    .Y(_03901_));
 sg13g2_xnor2_1 _21534_ (.Y(_03902_),
    .A(_10854_),
    .B(_03901_));
 sg13g2_nand2_1 _21535_ (.Y(_03903_),
    .A(net31),
    .B(_03902_));
 sg13g2_nor3_1 _21536_ (.A(_10852_),
    .B(_10847_),
    .C(_03878_),
    .Y(_03904_));
 sg13g2_o21ai_1 _21537_ (.B1(_10852_),
    .Y(_03905_),
    .A1(_10847_),
    .A2(_03878_));
 sg13g2_nor2b_1 _21538_ (.A(_03904_),
    .B_N(_03905_),
    .Y(_03906_));
 sg13g2_a221oi_1 _21539_ (.B2(_03906_),
    .C1(net271),
    .B1(net275),
    .A1(net491),
    .Y(_03907_),
    .A2(net598));
 sg13g2_nor2_1 _21540_ (.A(\cpu.ex.r_mult[18] ),
    .B(net349),
    .Y(_03908_));
 sg13g2_a21oi_1 _21541_ (.A1(_03903_),
    .A2(_03907_),
    .Y(_00955_),
    .B1(_03908_));
 sg13g2_xnor2_1 _21542_ (.Y(_03909_),
    .A(_00291_),
    .B(_03904_));
 sg13g2_a221oi_1 _21543_ (.B2(_03909_),
    .C1(net271),
    .B1(net275),
    .A1(net463),
    .Y(_03910_),
    .A2(_03860_));
 sg13g2_nor2b_1 _21544_ (.A(_03899_),
    .B_N(_10856_),
    .Y(_03911_));
 sg13g2_a21oi_1 _21545_ (.A1(net278),
    .A2(_10854_),
    .Y(_03912_),
    .B1(_03911_));
 sg13g2_xnor2_1 _21546_ (.Y(_03913_),
    .A(net236),
    .B(_03912_));
 sg13g2_nor3_1 _21547_ (.A(net28),
    .B(net32),
    .C(_03913_),
    .Y(_03914_));
 sg13g2_xnor2_1 _21548_ (.Y(_03915_),
    .A(_10859_),
    .B(_03914_));
 sg13g2_nand2_1 _21549_ (.Y(_03916_),
    .A(net31),
    .B(_03915_));
 sg13g2_nor2_1 _21550_ (.A(\cpu.ex.r_mult[19] ),
    .B(net349),
    .Y(_03917_));
 sg13g2_a21oi_1 _21551_ (.A1(_03910_),
    .A2(_03916_),
    .Y(_00956_),
    .B1(_03917_));
 sg13g2_nor4_1 _21552_ (.A(_00291_),
    .B(_10852_),
    .C(_10847_),
    .D(net616),
    .Y(_03918_));
 sg13g2_and4_1 _21553_ (.A(_11713_),
    .B(_11854_),
    .C(_03874_),
    .D(_03918_),
    .X(_03919_));
 sg13g2_and2_1 _21554_ (.A(_03877_),
    .B(_03918_),
    .X(_03920_));
 sg13g2_nor2_1 _21555_ (.A(_03919_),
    .B(_03920_),
    .Y(_03921_));
 sg13g2_buf_2 _21556_ (.A(_03921_),
    .X(_03922_));
 sg13g2_xnor2_1 _21557_ (.Y(_03923_),
    .A(_11376_),
    .B(_03922_));
 sg13g2_a221oi_1 _21558_ (.B2(_03923_),
    .C1(net271),
    .B1(net275),
    .A1(net452),
    .Y(_03924_),
    .A2(net539));
 sg13g2_a21o_1 _21559_ (.A2(net123),
    .A1(_10867_),
    .B1(_10874_),
    .X(_03925_));
 sg13g2_buf_1 _21560_ (.A(_03925_),
    .X(_03926_));
 sg13g2_nand2b_1 _21561_ (.Y(_03927_),
    .B(net281),
    .A_N(_03926_));
 sg13g2_buf_1 _21562_ (.A(_03927_),
    .X(_03928_));
 sg13g2_inv_1 _21563_ (.Y(_03929_),
    .A(_03928_));
 sg13g2_and2_1 _21564_ (.A(net277),
    .B(_03926_),
    .X(_03930_));
 sg13g2_nor4_1 _21565_ (.A(net28),
    .B(net32),
    .C(_03929_),
    .D(_03930_),
    .Y(_03931_));
 sg13g2_xor2_1 _21566_ (.B(_03931_),
    .A(_10828_),
    .X(_03932_));
 sg13g2_nand2_1 _21567_ (.Y(_03933_),
    .A(net31),
    .B(_03932_));
 sg13g2_nor2_1 _21568_ (.A(\cpu.ex.r_mult[20] ),
    .B(net349),
    .Y(_03934_));
 sg13g2_a21oi_1 _21569_ (.A1(_03924_),
    .A2(_03933_),
    .Y(_00957_),
    .B1(_03934_));
 sg13g2_nor3_2 _21570_ (.A(_10830_),
    .B(_10823_),
    .C(_03922_),
    .Y(_03935_));
 sg13g2_o21ai_1 _21571_ (.B1(_10830_),
    .Y(_03936_),
    .A1(_10823_),
    .A2(_03922_));
 sg13g2_nor2b_1 _21572_ (.A(_03935_),
    .B_N(_03936_),
    .Y(_03937_));
 sg13g2_a221oi_1 _21573_ (.B2(_03937_),
    .C1(net271),
    .B1(net275),
    .A1(net745),
    .Y(_03938_),
    .A2(net539));
 sg13g2_a21o_1 _21574_ (.A2(_03926_),
    .A1(net277),
    .B1(_10828_),
    .X(_03939_));
 sg13g2_a21oi_1 _21575_ (.A1(_03928_),
    .A2(_03939_),
    .Y(_03940_),
    .B1(net235));
 sg13g2_nand3_1 _21576_ (.B(_03928_),
    .C(_03939_),
    .A(net235),
    .Y(_03941_));
 sg13g2_inv_1 _21577_ (.Y(_03942_),
    .A(_03941_));
 sg13g2_nor4_1 _21578_ (.A(net28),
    .B(net32),
    .C(_03940_),
    .D(_03942_),
    .Y(_03943_));
 sg13g2_xor2_1 _21579_ (.B(_03943_),
    .A(_10844_),
    .X(_03944_));
 sg13g2_nand2_1 _21580_ (.Y(_03945_),
    .A(net31),
    .B(_03944_));
 sg13g2_nor2_1 _21581_ (.A(\cpu.ex.r_mult[21] ),
    .B(net349),
    .Y(_03946_));
 sg13g2_a21oi_1 _21582_ (.A1(_03938_),
    .A2(_03945_),
    .Y(_00958_),
    .B1(_03946_));
 sg13g2_nor2_1 _21583_ (.A(net1042),
    .B(net564),
    .Y(_03947_));
 sg13g2_xor2_1 _21584_ (.B(_03947_),
    .A(_03935_),
    .X(_03948_));
 sg13g2_a221oi_1 _21585_ (.B2(_03948_),
    .C1(net271),
    .B1(_11722_),
    .A1(net1000),
    .Y(_03949_),
    .A2(_03860_));
 sg13g2_buf_1 _21586_ (.A(_10834_),
    .X(_03950_));
 sg13g2_and2_1 _21587_ (.A(_10799_),
    .B(_03926_),
    .X(_03951_));
 sg13g2_nand3_1 _21588_ (.B(net235),
    .C(_03928_),
    .A(_11376_),
    .Y(_03952_));
 sg13g2_o21ai_1 _21589_ (.B1(_03928_),
    .Y(_03953_),
    .A1(_11376_),
    .A2(_03930_));
 sg13g2_a22oi_1 _21590_ (.Y(_03954_),
    .B1(_03953_),
    .B2(net282),
    .A2(_03952_),
    .A1(_10830_));
 sg13g2_nor2_1 _21591_ (.A(_03951_),
    .B(_03954_),
    .Y(_03955_));
 sg13g2_xnor2_1 _21592_ (.Y(_03956_),
    .A(net276),
    .B(_03955_));
 sg13g2_a221oi_1 _21593_ (.B2(_03956_),
    .C1(net1042),
    .B1(_11446_),
    .A1(\cpu.dec.div ),
    .Y(_03957_),
    .A2(_03950_));
 sg13g2_or2_1 _21594_ (.X(_03958_),
    .B(_11444_),
    .A(_11425_));
 sg13g2_buf_1 _21595_ (.A(_03958_),
    .X(_03959_));
 sg13g2_nand2_1 _21596_ (.Y(_03960_),
    .A(net276),
    .B(_03954_));
 sg13g2_a21oi_1 _21597_ (.A1(net1042),
    .A2(_03960_),
    .Y(_03961_),
    .B1(_11406_));
 sg13g2_a221oi_1 _21598_ (.B2(net566),
    .C1(net276),
    .B1(_03954_),
    .A1(_10799_),
    .Y(_03962_),
    .A2(_03926_));
 sg13g2_and2_1 _21599_ (.A(net276),
    .B(_03951_),
    .X(_03963_));
 sg13g2_nor4_1 _21600_ (.A(_03959_),
    .B(_03961_),
    .C(_03962_),
    .D(_03963_),
    .Y(_03964_));
 sg13g2_o21ai_1 _21601_ (.B1(net31),
    .Y(_03965_),
    .A1(_03957_),
    .A2(_03964_));
 sg13g2_nor2_1 _21602_ (.A(net1120),
    .B(net349),
    .Y(_03966_));
 sg13g2_a21oi_1 _21603_ (.A1(_03949_),
    .A2(_03965_),
    .Y(_00959_),
    .B1(_03966_));
 sg13g2_a21oi_1 _21604_ (.A1(_10813_),
    .A2(net232),
    .Y(_03967_),
    .B1(_10830_));
 sg13g2_nor2b_1 _21605_ (.A(_03940_),
    .B_N(_03967_),
    .Y(_03968_));
 sg13g2_a21oi_1 _21606_ (.A1(net232),
    .A2(_03941_),
    .Y(_03969_),
    .B1(_10813_));
 sg13g2_o21ai_1 _21607_ (.B1(net566),
    .Y(_03970_),
    .A1(_03968_),
    .A2(_03969_));
 sg13g2_nand2_1 _21608_ (.Y(_03971_),
    .A(net276),
    .B(_03942_));
 sg13g2_and3_1 _21609_ (.X(_03972_),
    .A(net233),
    .B(_03970_),
    .C(_03971_));
 sg13g2_a21oi_1 _21610_ (.A1(_03970_),
    .A2(_03971_),
    .Y(_03973_),
    .B1(net233));
 sg13g2_nor3_1 _21611_ (.A(_03959_),
    .B(_03972_),
    .C(_03973_),
    .Y(_03974_));
 sg13g2_nand2_1 _21612_ (.Y(_03975_),
    .A(_10810_),
    .B(net566));
 sg13g2_xor2_1 _21613_ (.B(_03975_),
    .A(_03974_),
    .X(_03976_));
 sg13g2_or2_1 _21614_ (.X(_03977_),
    .B(_03884_),
    .A(_10201_));
 sg13g2_nand2_1 _21615_ (.Y(_03978_),
    .A(_10199_),
    .B(_03977_));
 sg13g2_nor2_1 _21616_ (.A(\cpu.ex.r_mult[23] ),
    .B(_03881_),
    .Y(_03979_));
 sg13g2_nor2_1 _21617_ (.A(_03978_),
    .B(_03979_),
    .Y(_03980_));
 sg13g2_nand2_1 _21618_ (.Y(_03981_),
    .A(net87),
    .B(_03980_));
 sg13g2_nand2_1 _21619_ (.Y(_03982_),
    .A(_09353_),
    .B(net460));
 sg13g2_inv_1 _21620_ (.Y(_03983_),
    .A(_03982_));
 sg13g2_nor3_1 _21621_ (.A(net1042),
    .B(_10830_),
    .C(_10823_),
    .Y(_03984_));
 sg13g2_nor2b_1 _21622_ (.A(_03922_),
    .B_N(_03984_),
    .Y(_03985_));
 sg13g2_xnor2_1 _21623_ (.Y(_03986_),
    .A(_10811_),
    .B(_03985_));
 sg13g2_a21o_1 _21624_ (.A2(_03986_),
    .A1(_03983_),
    .B1(_03884_),
    .X(_03987_));
 sg13g2_a22oi_1 _21625_ (.Y(_03988_),
    .B1(_03980_),
    .B2(_03987_),
    .A2(net539),
    .A1(net998));
 sg13g2_o21ai_1 _21626_ (.B1(_03988_),
    .Y(_00960_),
    .A1(_03976_),
    .A2(_03981_));
 sg13g2_nand2_1 _21627_ (.Y(_03989_),
    .A(net1120),
    .B(_03985_));
 sg13g2_xor2_1 _21628_ (.B(_03989_),
    .A(_11388_),
    .X(_03990_));
 sg13g2_a221oi_1 _21629_ (.B2(_03990_),
    .C1(net271),
    .B1(net275),
    .A1(net1139),
    .Y(_03991_),
    .A2(net598));
 sg13g2_nor2_1 _21630_ (.A(_11388_),
    .B(net674),
    .Y(_03992_));
 sg13g2_nor2_1 _21631_ (.A(net169),
    .B(_11385_),
    .Y(_03993_));
 sg13g2_and2_1 _21632_ (.A(net169),
    .B(_11385_),
    .X(_03994_));
 sg13g2_nor4_1 _21633_ (.A(_03993_),
    .B(_03994_),
    .C(net28),
    .D(net32),
    .Y(_03995_));
 sg13g2_xor2_1 _21634_ (.B(_03995_),
    .A(_03992_),
    .X(_03996_));
 sg13g2_nand2_1 _21635_ (.Y(_03997_),
    .A(net31),
    .B(_03996_));
 sg13g2_nor2_1 _21636_ (.A(\cpu.ex.r_mult[24] ),
    .B(net349),
    .Y(_03998_));
 sg13g2_a21oi_1 _21637_ (.A1(_03991_),
    .A2(_03997_),
    .Y(_00961_),
    .B1(_03998_));
 sg13g2_nand3b_1 _21638_ (.B(_03985_),
    .C(net1120),
    .Y(_03999_),
    .A_N(_11388_));
 sg13g2_xnor2_1 _21639_ (.Y(_04000_),
    .A(_10809_),
    .B(_03999_));
 sg13g2_a221oi_1 _21640_ (.B2(_04000_),
    .C1(net271),
    .B1(net275),
    .A1(_10524_),
    .Y(_04001_),
    .A2(net598));
 sg13g2_a21oi_1 _21641_ (.A1(net566),
    .A2(_11389_),
    .Y(_04002_),
    .B1(_03993_));
 sg13g2_xnor2_1 _21642_ (.Y(_04003_),
    .A(net220),
    .B(_04002_));
 sg13g2_nor3_1 _21643_ (.A(net28),
    .B(net32),
    .C(_04003_),
    .Y(_04004_));
 sg13g2_nor2_1 _21644_ (.A(_10808_),
    .B(net674),
    .Y(_04005_));
 sg13g2_xor2_1 _21645_ (.B(_04005_),
    .A(_04004_),
    .X(_04006_));
 sg13g2_nand2_1 _21646_ (.Y(_04007_),
    .A(net31),
    .B(_04006_));
 sg13g2_nor2_1 _21647_ (.A(\cpu.ex.r_mult[25] ),
    .B(net349),
    .Y(_04008_));
 sg13g2_a21oi_1 _21648_ (.A1(_04001_),
    .A2(_04007_),
    .Y(_00962_),
    .B1(_04008_));
 sg13g2_nor3_1 _21649_ (.A(_10811_),
    .B(_10808_),
    .C(_11388_),
    .Y(_04009_));
 sg13g2_nand3b_1 _21650_ (.B(_03935_),
    .C(_04009_),
    .Y(_04010_),
    .A_N(net1042));
 sg13g2_xor2_1 _21651_ (.B(_04010_),
    .A(_11393_),
    .X(_04011_));
 sg13g2_a221oi_1 _21652_ (.B2(_04011_),
    .C1(_03885_),
    .B1(net275),
    .A1(_10392_),
    .Y(_04012_),
    .A2(net598));
 sg13g2_nand2_1 _21653_ (.Y(_04013_),
    .A(_10808_),
    .B(net220));
 sg13g2_a22oi_1 _21654_ (.Y(_04014_),
    .B1(_11386_),
    .B2(_10809_),
    .A2(_04013_),
    .A1(_11389_));
 sg13g2_inv_1 _21655_ (.Y(_04015_),
    .A(_11390_));
 sg13g2_o21ai_1 _21656_ (.B1(_04015_),
    .Y(_04016_),
    .A1(_11406_),
    .A2(_04014_));
 sg13g2_xnor2_1 _21657_ (.Y(_04017_),
    .A(_11401_),
    .B(_04016_));
 sg13g2_nor3_1 _21658_ (.A(net28),
    .B(net32),
    .C(_04017_),
    .Y(_04018_));
 sg13g2_nor2_1 _21659_ (.A(_11393_),
    .B(net674),
    .Y(_04019_));
 sg13g2_xor2_1 _21660_ (.B(_04019_),
    .A(_04018_),
    .X(_04020_));
 sg13g2_nand2_1 _21661_ (.Y(_04021_),
    .A(_03887_),
    .B(_04020_));
 sg13g2_nor2_1 _21662_ (.A(_10410_),
    .B(_03896_),
    .Y(_04022_));
 sg13g2_a21oi_1 _21663_ (.A1(_04012_),
    .A2(_04021_),
    .Y(_00963_),
    .B1(_04022_));
 sg13g2_o21ai_1 _21664_ (.B1(_03977_),
    .Y(_04023_),
    .A1(\cpu.ex.r_mult[27] ),
    .A2(_03881_));
 sg13g2_nand2_1 _21665_ (.Y(_04024_),
    .A(_03984_),
    .B(_04009_));
 sg13g2_nor2_1 _21666_ (.A(_11393_),
    .B(_04024_),
    .Y(_04025_));
 sg13g2_o21ai_1 _21667_ (.B1(_04025_),
    .Y(_04026_),
    .A1(_03919_),
    .A2(_03920_));
 sg13g2_buf_2 _21668_ (.A(_04026_),
    .X(_04027_));
 sg13g2_nor2_1 _21669_ (.A(_11231_),
    .B(net616),
    .Y(_04028_));
 sg13g2_nand2_1 _21670_ (.Y(_04029_),
    .A(_04028_),
    .B(_04027_));
 sg13g2_o21ai_1 _21671_ (.B1(_04029_),
    .Y(_04030_),
    .A1(_10410_),
    .A2(_04027_));
 sg13g2_a221oi_1 _21672_ (.B2(net1133),
    .C1(_03884_),
    .B1(_04030_),
    .A1(net1122),
    .Y(_04031_),
    .A2(net598));
 sg13g2_a21oi_1 _21673_ (.A1(net200),
    .A2(_11392_),
    .Y(_04032_),
    .B1(_11403_));
 sg13g2_nand2_1 _21674_ (.Y(_04033_),
    .A(_04032_),
    .B(_11395_));
 sg13g2_xnor2_1 _21675_ (.Y(_04034_),
    .A(net215),
    .B(_04033_));
 sg13g2_a21oi_1 _21676_ (.A1(_11446_),
    .A2(_04034_),
    .Y(_04035_),
    .B1(_11397_));
 sg13g2_and3_1 _21677_ (.X(_04036_),
    .A(_11397_),
    .B(_11446_),
    .C(_04034_));
 sg13g2_o21ai_1 _21678_ (.B1(net87),
    .Y(_04037_),
    .A1(_04035_),
    .A2(_04036_));
 sg13g2_nor2_1 _21679_ (.A(net999),
    .B(_10199_),
    .Y(_04038_));
 sg13g2_a221oi_1 _21680_ (.B2(_04037_),
    .C1(_04038_),
    .B1(_04031_),
    .A1(_10199_),
    .Y(_00964_),
    .A2(_04023_));
 sg13g2_nand2_1 _21681_ (.Y(_04039_),
    .A(_03499_),
    .B(net539));
 sg13g2_inv_1 _21682_ (.Y(_04040_),
    .A(_03978_));
 sg13g2_o21ai_1 _21683_ (.B1(_04040_),
    .Y(_04041_),
    .A1(_10322_),
    .A2(_03881_));
 sg13g2_nor2_1 _21684_ (.A(net199),
    .B(_11397_),
    .Y(_04042_));
 sg13g2_a21o_1 _21685_ (.A2(_11405_),
    .A1(_11395_),
    .B1(_04042_),
    .X(_04043_));
 sg13g2_xnor2_1 _21686_ (.Y(_04044_),
    .A(net144),
    .B(_04043_));
 sg13g2_nand2_1 _21687_ (.Y(_04045_),
    .A(_11411_),
    .B(net566));
 sg13g2_a21oi_1 _21688_ (.A1(_11446_),
    .A2(_04044_),
    .Y(_04046_),
    .B1(_04045_));
 sg13g2_and3_1 _21689_ (.X(_04047_),
    .A(_11446_),
    .B(_04045_),
    .C(_04044_));
 sg13g2_o21ai_1 _21690_ (.B1(net87),
    .Y(_04048_),
    .A1(_04046_),
    .A2(_04047_));
 sg13g2_nor2_1 _21691_ (.A(_11231_),
    .B(_04027_),
    .Y(_04049_));
 sg13g2_xnor2_1 _21692_ (.Y(_04050_),
    .A(_11410_),
    .B(_04049_));
 sg13g2_a221oi_1 _21693_ (.B2(_04050_),
    .C1(_03885_),
    .B1(_03983_),
    .A1(net617),
    .Y(_04051_),
    .A2(net539));
 sg13g2_a22oi_1 _21694_ (.Y(_00965_),
    .B1(_04048_),
    .B2(_04051_),
    .A2(_04041_),
    .A1(_04039_));
 sg13g2_nand2_1 _21695_ (.Y(_04052_),
    .A(_11411_),
    .B(_04028_));
 sg13g2_inv_1 _21696_ (.Y(_04053_),
    .A(net275));
 sg13g2_nor2_1 _21697_ (.A(_10323_),
    .B(_04053_),
    .Y(_04054_));
 sg13g2_o21ai_1 _21698_ (.B1(_04054_),
    .Y(_04055_),
    .A1(_04027_),
    .A2(_04052_));
 sg13g2_or4_1 _21699_ (.A(_10322_),
    .B(_04053_),
    .C(_04027_),
    .D(_04052_),
    .X(_04056_));
 sg13g2_a21oi_1 _21700_ (.A1(net577),
    .A2(net598),
    .Y(_04057_),
    .B1(_03884_));
 sg13g2_and3_1 _21701_ (.X(_04058_),
    .A(_04055_),
    .B(_04056_),
    .C(_04057_));
 sg13g2_buf_1 _21702_ (.A(_04058_),
    .X(_04059_));
 sg13g2_nor2_1 _21703_ (.A(_11397_),
    .B(_04045_),
    .Y(_04060_));
 sg13g2_nor2_1 _21704_ (.A(net144),
    .B(_04045_),
    .Y(_04061_));
 sg13g2_a21oi_1 _21705_ (.A1(net215),
    .A2(_04060_),
    .Y(_04062_),
    .B1(_04061_));
 sg13g2_o21ai_1 _21706_ (.B1(_04062_),
    .Y(_04063_),
    .A1(_11397_),
    .A2(_11814_));
 sg13g2_a221oi_1 _21707_ (.B2(net144),
    .C1(_04033_),
    .B1(_04045_),
    .A1(net199),
    .Y(_04064_),
    .A2(_11397_));
 sg13g2_nor3_1 _21708_ (.A(net219),
    .B(net28),
    .C(net32),
    .Y(_04065_));
 sg13g2_o21ai_1 _21709_ (.B1(_04065_),
    .Y(_04066_),
    .A1(_04063_),
    .A2(_04064_));
 sg13g2_or4_1 _21710_ (.A(net197),
    .B(_03959_),
    .C(_04063_),
    .D(_04064_),
    .X(_04067_));
 sg13g2_nand2_1 _21711_ (.Y(_04068_),
    .A(_10322_),
    .B(net566));
 sg13g2_and4_1 _21712_ (.A(_04059_),
    .B(_04066_),
    .C(_04067_),
    .D(_04068_),
    .X(_04069_));
 sg13g2_nand3_1 _21713_ (.B(_11402_),
    .C(_04059_),
    .A(_10322_),
    .Y(_04070_));
 sg13g2_a21oi_1 _21714_ (.A1(_04066_),
    .A2(_04067_),
    .Y(_04071_),
    .B1(_04070_));
 sg13g2_nand2_1 _21715_ (.Y(_04072_),
    .A(_11761_),
    .B(_04059_));
 sg13g2_o21ai_1 _21716_ (.B1(_04072_),
    .Y(_04073_),
    .A1(_10263_),
    .A2(_03896_));
 sg13g2_nor3_1 _21717_ (.A(_04069_),
    .B(_04071_),
    .C(_04073_),
    .Y(_00966_));
 sg13g2_nor2_1 _21718_ (.A(\cpu.ex.r_mult[30] ),
    .B(_03895_),
    .Y(_04074_));
 sg13g2_nor2_1 _21719_ (.A(net674),
    .B(_11413_),
    .Y(_04075_));
 sg13g2_a21oi_1 _21720_ (.A1(_11437_),
    .A2(_04043_),
    .Y(_04076_),
    .B1(_04075_));
 sg13g2_xnor2_1 _21721_ (.Y(_04077_),
    .A(net168),
    .B(_04076_));
 sg13g2_or4_1 _21722_ (.A(_10323_),
    .B(_11393_),
    .C(_04024_),
    .D(_04052_),
    .X(_04078_));
 sg13g2_nor2_1 _21723_ (.A(_03922_),
    .B(_04078_),
    .Y(_04079_));
 sg13g2_xnor2_1 _21724_ (.Y(_04080_),
    .A(_10263_),
    .B(_04079_));
 sg13g2_a21oi_1 _21725_ (.A1(net688),
    .A2(net598),
    .Y(_04081_),
    .B1(_03884_));
 sg13g2_o21ai_1 _21726_ (.B1(_04081_),
    .Y(_04082_),
    .A1(_04053_),
    .A2(_04080_));
 sg13g2_a221oi_1 _21727_ (.B2(_04077_),
    .C1(_04082_),
    .B1(_11446_),
    .A1(_10263_),
    .Y(_04083_),
    .A2(_11402_));
 sg13g2_xnor2_1 _21728_ (.Y(_04084_),
    .A(net201),
    .B(_04076_));
 sg13g2_nor4_1 _21729_ (.A(_11438_),
    .B(_03959_),
    .C(_04082_),
    .D(_04084_),
    .Y(_04085_));
 sg13g2_nor2_1 _21730_ (.A(_03887_),
    .B(_04082_),
    .Y(_04086_));
 sg13g2_nor4_1 _21731_ (.A(_04074_),
    .B(_04083_),
    .C(_04085_),
    .D(_04086_),
    .Y(_00967_));
 sg13g2_nor3_1 _21732_ (.A(_11409_),
    .B(_03922_),
    .C(_04078_),
    .Y(_04087_));
 sg13g2_xnor2_1 _21733_ (.Y(_04088_),
    .A(_00283_),
    .B(_04087_));
 sg13g2_a21oi_1 _21734_ (.A1(_11395_),
    .A2(_11405_),
    .Y(_04089_),
    .B1(_04042_));
 sg13g2_o21ai_1 _21735_ (.B1(_11419_),
    .Y(_04090_),
    .A1(_11440_),
    .A2(_04089_));
 sg13g2_xnor2_1 _21736_ (.Y(_04091_),
    .A(_11875_),
    .B(_04090_));
 sg13g2_nor2b_1 _21737_ (.A(_11408_),
    .B_N(net87),
    .Y(_04092_));
 sg13g2_a221oi_1 _21738_ (.B2(_04092_),
    .C1(_03884_),
    .B1(_04091_),
    .A1(_03983_),
    .Y(_04093_),
    .A2(_04088_));
 sg13g2_o21ai_1 _21739_ (.B1(_04040_),
    .Y(_04094_),
    .A1(\cpu.ex.r_mult[31] ),
    .A2(_03881_));
 sg13g2_nand2_1 _21740_ (.Y(_04095_),
    .A(net860),
    .B(net539));
 sg13g2_o21ai_1 _21741_ (.B1(_04095_),
    .Y(_00968_),
    .A1(_04093_),
    .A2(_04094_));
 sg13g2_inv_1 _21742_ (.Y(_04096_),
    .A(_00242_));
 sg13g2_nand2_1 _21743_ (.Y(_04097_),
    .A(net1143),
    .B(_04096_));
 sg13g2_mux2_1 _21744_ (.A0(net1074),
    .A1(_04097_),
    .S(_11936_),
    .X(_04098_));
 sg13g2_nor2_1 _21745_ (.A(_09210_),
    .B(_09207_),
    .Y(_04099_));
 sg13g2_buf_2 _21746_ (.A(_04099_),
    .X(_04100_));
 sg13g2_nand3b_1 _21747_ (.B(_04100_),
    .C(net665),
    .Y(_04101_),
    .A_N(_04098_));
 sg13g2_buf_1 _21748_ (.A(_04101_),
    .X(_04102_));
 sg13g2_buf_1 _21749_ (.A(_04102_),
    .X(_04103_));
 sg13g2_nor2b_1 _21750_ (.A(_11457_),
    .B_N(_11467_),
    .Y(_04104_));
 sg13g2_buf_2 _21751_ (.A(_04104_),
    .X(_04105_));
 sg13g2_buf_1 _21752_ (.A(_04105_),
    .X(_04106_));
 sg13g2_buf_1 _21753_ (.A(net206),
    .X(_04107_));
 sg13g2_nor2_2 _21754_ (.A(_03722_),
    .B(_03723_),
    .Y(_04108_));
 sg13g2_xnor2_1 _21755_ (.Y(_04109_),
    .A(net227),
    .B(_04108_));
 sg13g2_buf_1 _21756_ (.A(_10869_),
    .X(_04110_));
 sg13g2_nor2_1 _21757_ (.A(_09130_),
    .B(_09879_),
    .Y(_04111_));
 sg13g2_nor4_1 _21758_ (.A(_09088_),
    .B(_09146_),
    .C(net1131),
    .D(\cpu.dec.r_op[8] ),
    .Y(_04112_));
 sg13g2_nor4_1 _21759_ (.A(_08335_),
    .B(_09133_),
    .C(\cpu.dec.r_op[3] ),
    .D(_09877_),
    .Y(_04113_));
 sg13g2_and3_1 _21760_ (.X(_04114_),
    .A(_04111_),
    .B(_04112_),
    .C(_04113_));
 sg13g2_buf_1 _21761_ (.A(_04114_),
    .X(_04115_));
 sg13g2_nor3_1 _21762_ (.A(_09133_),
    .B(_09877_),
    .C(net744),
    .Y(_04116_));
 sg13g2_nand3_1 _21763_ (.B(_04109_),
    .C(_04116_),
    .A(net226),
    .Y(_04117_));
 sg13g2_o21ai_1 _21764_ (.B1(_04117_),
    .Y(_04118_),
    .A1(_08335_),
    .A2(_04109_));
 sg13g2_nor2_1 _21765_ (.A(net218),
    .B(net279),
    .Y(_04119_));
 sg13g2_a21oi_1 _21766_ (.A1(_04119_),
    .A2(_04109_),
    .Y(_04120_),
    .B1(_04116_));
 sg13g2_or3_1 _21767_ (.A(_09133_),
    .B(_09877_),
    .C(net744),
    .X(_04121_));
 sg13g2_buf_1 _21768_ (.A(_04121_),
    .X(_04122_));
 sg13g2_o21ai_1 _21769_ (.B1(net226),
    .Y(_04123_),
    .A1(net279),
    .A2(_04122_));
 sg13g2_nand2b_1 _21770_ (.Y(_04124_),
    .B(_04123_),
    .A_N(_04109_));
 sg13g2_o21ai_1 _21771_ (.B1(_04124_),
    .Y(_04125_),
    .A1(_08335_),
    .A2(_04120_));
 sg13g2_a21oi_1 _21772_ (.A1(_11078_),
    .A2(_04118_),
    .Y(_04126_),
    .B1(_04125_));
 sg13g2_nor2_1 _21773_ (.A(net238),
    .B(_04108_),
    .Y(_04127_));
 sg13g2_nor2_1 _21774_ (.A(net1140),
    .B(_04127_),
    .Y(_04128_));
 sg13g2_a21oi_1 _21775_ (.A1(_09147_),
    .A2(_04127_),
    .Y(_04129_),
    .B1(_04128_));
 sg13g2_nor2_1 _21776_ (.A(net1063),
    .B(_04129_),
    .Y(_04130_));
 sg13g2_buf_1 _21777_ (.A(_09088_),
    .X(_04131_));
 sg13g2_buf_1 _21778_ (.A(_10620_),
    .X(_04132_));
 sg13g2_nor3_1 _21779_ (.A(net227),
    .B(net240),
    .C(net189),
    .Y(_04133_));
 sg13g2_buf_2 _21780_ (.A(_04133_),
    .X(_04134_));
 sg13g2_buf_1 _21781_ (.A(_04134_),
    .X(_04135_));
 sg13g2_buf_1 _21782_ (.A(net118),
    .X(_04136_));
 sg13g2_nor2_1 _21783_ (.A(_09892_),
    .B(net279),
    .Y(_04137_));
 sg13g2_a221oi_1 _21784_ (.B2(_04137_),
    .C1(net206),
    .B1(net106),
    .A1(net991),
    .Y(_04138_),
    .A2(net220));
 sg13g2_o21ai_1 _21785_ (.B1(_04138_),
    .Y(_04139_),
    .A1(_03724_),
    .A2(_04130_));
 sg13g2_nor2_1 _21786_ (.A(_04126_),
    .B(_04139_),
    .Y(_04140_));
 sg13g2_buf_1 _21787_ (.A(_04111_),
    .X(_04141_));
 sg13g2_and2_1 _21788_ (.A(_09130_),
    .B(_03565_),
    .X(_04142_));
 sg13g2_buf_1 _21789_ (.A(_04142_),
    .X(_04143_));
 sg13g2_buf_1 _21790_ (.A(net238),
    .X(_04144_));
 sg13g2_o21ai_1 _21791_ (.B1(net205),
    .Y(_04145_),
    .A1(_04110_),
    .A2(net159));
 sg13g2_buf_1 _21792_ (.A(net208),
    .X(_04146_));
 sg13g2_nor2_1 _21793_ (.A(net238),
    .B(net226),
    .Y(_04147_));
 sg13g2_buf_2 _21794_ (.A(_04147_),
    .X(_04148_));
 sg13g2_nand2_1 _21795_ (.Y(_04149_),
    .A(net188),
    .B(_04148_));
 sg13g2_a21oi_1 _21796_ (.A1(_04145_),
    .A2(_04149_),
    .Y(_04150_),
    .B1(net189));
 sg13g2_nor2_1 _21797_ (.A(net286),
    .B(net236),
    .Y(_04151_));
 sg13g2_buf_1 _21798_ (.A(_04151_),
    .X(_04152_));
 sg13g2_nand3_1 _21799_ (.B(net120),
    .C(net187),
    .A(net226),
    .Y(_04153_));
 sg13g2_buf_1 _21800_ (.A(_03770_),
    .X(_04154_));
 sg13g2_nor2_1 _21801_ (.A(net360),
    .B(net236),
    .Y(_04155_));
 sg13g2_nand3_1 _21802_ (.B(net186),
    .C(_04155_),
    .A(_11448_),
    .Y(_04156_));
 sg13g2_a21oi_1 _21803_ (.A1(_04153_),
    .A2(_04156_),
    .Y(_04157_),
    .B1(net207));
 sg13g2_nand2_1 _21804_ (.Y(_04158_),
    .A(net286),
    .B(_11539_));
 sg13g2_buf_2 _21805_ (.A(_04158_),
    .X(_04159_));
 sg13g2_nor3_1 _21806_ (.A(net238),
    .B(net240),
    .C(_04159_),
    .Y(_04160_));
 sg13g2_buf_2 _21807_ (.A(_04160_),
    .X(_04161_));
 sg13g2_nand2_1 _21808_ (.Y(_04162_),
    .A(net107),
    .B(_04161_));
 sg13g2_buf_1 _21809_ (.A(_03610_),
    .X(_04163_));
 sg13g2_nor3_1 _21810_ (.A(net284),
    .B(net240),
    .C(_10620_),
    .Y(_04164_));
 sg13g2_buf_2 _21811_ (.A(_04164_),
    .X(_04165_));
 sg13g2_buf_1 _21812_ (.A(_04165_),
    .X(_04166_));
 sg13g2_nand2_1 _21813_ (.Y(_04167_),
    .A(net158),
    .B(net139));
 sg13g2_nor3_1 _21814_ (.A(net227),
    .B(_11447_),
    .C(_04159_),
    .Y(_04168_));
 sg13g2_buf_1 _21815_ (.A(_04168_),
    .X(_04169_));
 sg13g2_nand2_2 _21816_ (.Y(_04170_),
    .A(net360),
    .B(net236));
 sg13g2_nor3_1 _21817_ (.A(_10849_),
    .B(net240),
    .C(_04170_),
    .Y(_04171_));
 sg13g2_buf_1 _21818_ (.A(_04171_),
    .X(_04172_));
 sg13g2_buf_1 _21819_ (.A(net157),
    .X(_04173_));
 sg13g2_buf_1 _21820_ (.A(_03622_),
    .X(_04174_));
 sg13g2_a22oi_1 _21821_ (.Y(_04175_),
    .B1(net137),
    .B2(net185),
    .A2(net138),
    .A1(net192));
 sg13g2_nor2_1 _21822_ (.A(net238),
    .B(net240),
    .Y(_04176_));
 sg13g2_nand3_1 _21823_ (.B(_04176_),
    .C(net187),
    .A(net159),
    .Y(_04177_));
 sg13g2_nand4_1 _21824_ (.B(_04167_),
    .C(_04175_),
    .A(_04162_),
    .Y(_04178_),
    .D(_04177_));
 sg13g2_nor3_1 _21825_ (.A(net284),
    .B(_10674_),
    .C(_04170_),
    .Y(_04179_));
 sg13g2_buf_2 _21826_ (.A(_04179_),
    .X(_04180_));
 sg13g2_nand2_1 _21827_ (.Y(_04181_),
    .A(_03767_),
    .B(_04180_));
 sg13g2_nor3_1 _21828_ (.A(net284),
    .B(_10869_),
    .C(_04170_),
    .Y(_04182_));
 sg13g2_buf_1 _21829_ (.A(_04182_),
    .X(_04183_));
 sg13g2_buf_1 _21830_ (.A(net156),
    .X(_04184_));
 sg13g2_nor3_2 _21831_ (.A(_10849_),
    .B(_10869_),
    .C(_04170_),
    .Y(_04185_));
 sg13g2_buf_1 _21832_ (.A(_04185_),
    .X(_04186_));
 sg13g2_buf_1 _21833_ (.A(net155),
    .X(_04187_));
 sg13g2_buf_1 _21834_ (.A(_03577_),
    .X(_04188_));
 sg13g2_a22oi_1 _21835_ (.Y(_04189_),
    .B1(net135),
    .B2(net154),
    .A2(net136),
    .A1(net191));
 sg13g2_nand3_1 _21836_ (.B(_04148_),
    .C(net187),
    .A(net193),
    .Y(_04190_));
 sg13g2_nand2_1 _21837_ (.Y(_04191_),
    .A(_10851_),
    .B(net237));
 sg13g2_nor2_1 _21838_ (.A(_10675_),
    .B(_04191_),
    .Y(_04192_));
 sg13g2_buf_1 _21839_ (.A(_04192_),
    .X(_04193_));
 sg13g2_nor3_1 _21840_ (.A(net238),
    .B(net226),
    .C(_04159_),
    .Y(_04194_));
 sg13g2_buf_2 _21841_ (.A(_04194_),
    .X(_04195_));
 sg13g2_buf_1 _21842_ (.A(_03570_),
    .X(_04196_));
 sg13g2_a22oi_1 _21843_ (.Y(_04197_),
    .B1(_04195_),
    .B2(net134),
    .A2(_04193_),
    .A1(net119));
 sg13g2_nand4_1 _21844_ (.B(_04189_),
    .C(_04190_),
    .A(_04181_),
    .Y(_04198_),
    .D(_04197_));
 sg13g2_nor4_1 _21845_ (.A(_04150_),
    .B(_04157_),
    .C(_04178_),
    .D(_04198_),
    .Y(_04199_));
 sg13g2_buf_1 _21846_ (.A(_03599_),
    .X(_04200_));
 sg13g2_nor2_1 _21847_ (.A(net227),
    .B(net240),
    .Y(_04201_));
 sg13g2_nand2b_1 _21848_ (.Y(_04202_),
    .B(_04201_),
    .A_N(net189));
 sg13g2_buf_2 _21849_ (.A(_04202_),
    .X(_04203_));
 sg13g2_nor2_1 _21850_ (.A(net184),
    .B(_04203_),
    .Y(_04204_));
 sg13g2_or3_1 _21851_ (.A(net856),
    .B(_04199_),
    .C(_04204_),
    .X(_04205_));
 sg13g2_a22oi_1 _21852_ (.Y(_04206_),
    .B1(_04140_),
    .B2(_04205_),
    .A2(_11511_),
    .A1(net190));
 sg13g2_inv_1 _21853_ (.Y(_04207_),
    .A(_04206_));
 sg13g2_and4_1 _21854_ (.A(net1143),
    .B(net665),
    .C(_04100_),
    .D(_11937_),
    .X(_04208_));
 sg13g2_buf_1 _21855_ (.A(_04208_),
    .X(_04209_));
 sg13g2_or2_1 _21856_ (.X(_04210_),
    .B(_09207_),
    .A(_09210_));
 sg13g2_buf_1 _21857_ (.A(_04210_),
    .X(_04211_));
 sg13g2_nor3_2 _21858_ (.A(_11475_),
    .B(_04211_),
    .C(_04098_),
    .Y(_04212_));
 sg13g2_nand2_1 _21859_ (.Y(_04213_),
    .A(_09208_),
    .B(_11474_));
 sg13g2_mux2_1 _21860_ (.A0(_04213_),
    .A1(_11474_),
    .S(net371),
    .X(_04214_));
 sg13g2_nor2_1 _21861_ (.A(net1074),
    .B(_04214_),
    .Y(_04215_));
 sg13g2_inv_1 _21862_ (.Y(_04216_),
    .A(_09210_));
 sg13g2_nand4_1 _21863_ (.B(_04216_),
    .C(_09207_),
    .A(_08454_),
    .Y(_04217_),
    .D(net665));
 sg13g2_nand2_1 _21864_ (.Y(_04218_),
    .A(_09156_),
    .B(_04217_));
 sg13g2_nor4_1 _21865_ (.A(_04212_),
    .B(_04209_),
    .C(_04215_),
    .D(_04218_),
    .Y(_04219_));
 sg13g2_buf_1 _21866_ (.A(_04219_),
    .X(_04220_));
 sg13g2_buf_1 _21867_ (.A(_04220_),
    .X(_04221_));
 sg13g2_a22oi_1 _21868_ (.Y(_04222_),
    .B1(_04221_),
    .B2(net804),
    .A2(net97),
    .A1(_10643_));
 sg13g2_o21ai_1 _21869_ (.B1(_04222_),
    .Y(_00969_),
    .A1(net86),
    .A2(_04207_));
 sg13g2_nand2_1 _21870_ (.Y(_04223_),
    .A(net233),
    .B(_03628_));
 sg13g2_and2_1 _21871_ (.A(_04223_),
    .B(_03640_),
    .X(_04224_));
 sg13g2_buf_1 _21872_ (.A(_04224_),
    .X(_04225_));
 sg13g2_nand3_1 _21873_ (.B(_03735_),
    .C(_03738_),
    .A(_03702_),
    .Y(_04226_));
 sg13g2_nand2_1 _21874_ (.Y(_04227_),
    .A(net232),
    .B(_03622_));
 sg13g2_nor2_1 _21875_ (.A(net232),
    .B(_03622_),
    .Y(_04228_));
 sg13g2_a21oi_1 _21876_ (.A1(_04226_),
    .A2(_04227_),
    .Y(_04229_),
    .B1(_04228_));
 sg13g2_xnor2_1 _21877_ (.Y(_04230_),
    .A(_04225_),
    .B(_04229_));
 sg13g2_a21oi_1 _21878_ (.A1(_09877_),
    .A2(_04230_),
    .Y(_04231_),
    .B1(_04115_));
 sg13g2_or2_1 _21879_ (.X(_04232_),
    .B(_03657_),
    .A(_03654_));
 sg13g2_and2_1 _21880_ (.A(_03572_),
    .B(_03658_),
    .X(_04233_));
 sg13g2_xnor2_1 _21881_ (.Y(_04234_),
    .A(_04232_),
    .B(_04233_));
 sg13g2_nand2b_1 _21882_ (.Y(_04235_),
    .B(net106),
    .A_N(_03799_));
 sg13g2_nand3_1 _21883_ (.B(net161),
    .C(_04187_),
    .A(_09879_),
    .Y(_04236_));
 sg13g2_nor2_1 _21884_ (.A(net227),
    .B(_04143_),
    .Y(_04237_));
 sg13g2_nor3_1 _21885_ (.A(net205),
    .B(_04132_),
    .C(net119),
    .Y(_04238_));
 sg13g2_o21ai_1 _21886_ (.B1(net218),
    .Y(_04239_),
    .A1(_04237_),
    .A2(_04238_));
 sg13g2_nand2_2 _21887_ (.Y(_04240_),
    .A(_09130_),
    .B(_03565_));
 sg13g2_a21oi_1 _21888_ (.A1(net189),
    .A2(_04240_),
    .Y(_04241_),
    .B1(_04141_));
 sg13g2_nand2_1 _21889_ (.Y(_04242_),
    .A(_03675_),
    .B(_04166_));
 sg13g2_nand3_1 _21890_ (.B(_04241_),
    .C(_04242_),
    .A(_04239_),
    .Y(_04243_));
 sg13g2_nand2_1 _21891_ (.Y(_04244_),
    .A(_04236_),
    .B(_04243_));
 sg13g2_buf_1 _21892_ (.A(_03728_),
    .X(_04245_));
 sg13g2_nor3_1 _21893_ (.A(_10650_),
    .B(_10869_),
    .C(_10620_),
    .Y(_04246_));
 sg13g2_buf_1 _21894_ (.A(_04246_),
    .X(_04247_));
 sg13g2_buf_1 _21895_ (.A(_04247_),
    .X(_04248_));
 sg13g2_a221oi_1 _21896_ (.B2(net186),
    .C1(net118),
    .B1(net133),
    .A1(_04245_),
    .Y(_04249_),
    .A2(_04161_));
 sg13g2_buf_1 _21897_ (.A(_03767_),
    .X(_04250_));
 sg13g2_nor2_1 _21898_ (.A(_10675_),
    .B(_04159_),
    .Y(_04251_));
 sg13g2_buf_1 _21899_ (.A(_04251_),
    .X(_04252_));
 sg13g2_buf_1 _21900_ (.A(_04252_),
    .X(_04253_));
 sg13g2_a22oi_1 _21901_ (.Y(_04254_),
    .B1(net117),
    .B2(net188),
    .A2(net139),
    .A1(net132));
 sg13g2_a22oi_1 _21902_ (.Y(_04255_),
    .B1(net136),
    .B2(_04188_),
    .A2(net138),
    .A1(_03599_));
 sg13g2_or2_1 _21903_ (.X(_04256_),
    .B(_03723_),
    .A(_03722_));
 sg13g2_buf_1 _21904_ (.A(_04256_),
    .X(_04257_));
 sg13g2_nand2_1 _21905_ (.Y(_04258_),
    .A(net185),
    .B(net157));
 sg13g2_nand2_1 _21906_ (.Y(_04259_),
    .A(net191),
    .B(_04185_));
 sg13g2_nand2_1 _21907_ (.Y(_04260_),
    .A(_04258_),
    .B(_04259_));
 sg13g2_a221oi_1 _21908_ (.B2(_04257_),
    .C1(_04260_),
    .B1(_04195_),
    .A1(_03610_),
    .Y(_04261_),
    .A2(_04180_));
 sg13g2_nand4_1 _21909_ (.B(_04254_),
    .C(_04255_),
    .A(_04249_),
    .Y(_04262_),
    .D(_04261_));
 sg13g2_nand2_1 _21910_ (.Y(_04263_),
    .A(_03651_),
    .B(net118));
 sg13g2_nand3_1 _21911_ (.B(_04262_),
    .C(_04263_),
    .A(_09891_),
    .Y(_04264_));
 sg13g2_nor2_1 _21912_ (.A(_09136_),
    .B(_03784_),
    .Y(_04265_));
 sg13g2_a21oi_1 _21913_ (.A1(_09147_),
    .A2(_03784_),
    .Y(_04266_),
    .B1(_04265_));
 sg13g2_o21ai_1 _21914_ (.B1(_03694_),
    .Y(_04267_),
    .A1(net1063),
    .A2(_04266_));
 sg13g2_nand2_1 _21915_ (.Y(_04268_),
    .A(net991),
    .B(net217));
 sg13g2_nand3_1 _21916_ (.B(_04267_),
    .C(_04268_),
    .A(_04264_),
    .Y(_04269_));
 sg13g2_a221oi_1 _21917_ (.B2(_04244_),
    .C1(_04269_),
    .B1(_04235_),
    .A1(_08336_),
    .Y(_04270_),
    .A2(_04234_));
 sg13g2_nand2_1 _21918_ (.Y(_04271_),
    .A(_03696_),
    .B(net200));
 sg13g2_a21oi_1 _21919_ (.A1(_03780_),
    .A2(_04271_),
    .Y(_04272_),
    .B1(_03789_));
 sg13g2_xor2_1 _21920_ (.B(_04233_),
    .A(_04272_),
    .X(_04273_));
 sg13g2_a22oi_1 _21921_ (.Y(_04274_),
    .B1(_04273_),
    .B2(net744),
    .A2(_04270_),
    .A1(_04231_));
 sg13g2_nor2_1 _21922_ (.A(net239),
    .B(_11763_),
    .Y(_04275_));
 sg13g2_a21oi_1 _21923_ (.A1(net239),
    .A2(_04274_),
    .Y(_04276_),
    .B1(_04275_));
 sg13g2_nor2_1 _21924_ (.A(_08946_),
    .B(_08527_),
    .Y(_04277_));
 sg13g2_and2_1 _21925_ (.A(net1141),
    .B(_04277_),
    .X(_04278_));
 sg13g2_buf_1 _21926_ (.A(_04278_),
    .X(_04279_));
 sg13g2_nand4_1 _21927_ (.B(_08718_),
    .C(_08699_),
    .A(_08671_),
    .Y(_04280_),
    .D(_04279_));
 sg13g2_nor2_1 _21928_ (.A(_08709_),
    .B(_04280_),
    .Y(_04281_));
 sg13g2_nand3_1 _21929_ (.B(_08688_),
    .C(_04281_),
    .A(_08679_),
    .Y(_04282_));
 sg13g2_xnor2_1 _21930_ (.Y(_04283_),
    .A(_10385_),
    .B(_04282_));
 sg13g2_buf_1 _21931_ (.A(net97),
    .X(_04284_));
 sg13g2_a22oi_1 _21932_ (.Y(_04285_),
    .B1(_04283_),
    .B2(net85),
    .A2(net35),
    .A1(\cpu.ex.pc[11] ));
 sg13g2_o21ai_1 _21933_ (.B1(_04285_),
    .Y(_00970_),
    .A1(net86),
    .A2(_04276_));
 sg13g2_o21ai_1 _21934_ (.B1(net215),
    .Y(_04286_),
    .A1(_03571_),
    .A2(_03789_));
 sg13g2_o21ai_1 _21935_ (.B1(_04286_),
    .Y(_04287_),
    .A1(_04196_),
    .A2(_03790_));
 sg13g2_and2_1 _21936_ (.A(_03679_),
    .B(_03671_),
    .X(_04288_));
 sg13g2_buf_1 _21937_ (.A(_04288_),
    .X(_04289_));
 sg13g2_mux2_1 _21938_ (.A0(_04287_),
    .A1(_03784_),
    .S(_04289_),
    .X(_04290_));
 sg13g2_nor2b_1 _21939_ (.A(_03798_),
    .B_N(_04289_),
    .Y(_04291_));
 sg13g2_o21ai_1 _21940_ (.B1(net744),
    .Y(_04292_),
    .A1(_04290_),
    .A2(_04291_));
 sg13g2_nand3_1 _21941_ (.B(_04112_),
    .C(_04113_),
    .A(net856),
    .Y(_04293_));
 sg13g2_buf_1 _21942_ (.A(_04293_),
    .X(_04294_));
 sg13g2_nor4_1 _21943_ (.A(_03784_),
    .B(_03788_),
    .C(_04294_),
    .D(_04289_),
    .Y(_04295_));
 sg13g2_nand2_1 _21944_ (.Y(_04296_),
    .A(net204),
    .B(_04193_));
 sg13g2_a21oi_1 _21945_ (.A1(net186),
    .A2(_04165_),
    .Y(_04297_),
    .B1(_04135_));
 sg13g2_a22oi_1 _21946_ (.Y(_04298_),
    .B1(_04195_),
    .B2(net184),
    .A2(net137),
    .A1(net191));
 sg13g2_nand2b_1 _21947_ (.Y(_04299_),
    .B(_04148_),
    .A_N(net189));
 sg13g2_nor2_1 _21948_ (.A(_03651_),
    .B(_04299_),
    .Y(_04300_));
 sg13g2_a21oi_1 _21949_ (.A1(net132),
    .A2(_04186_),
    .Y(_04301_),
    .B1(_04300_));
 sg13g2_buf_1 _21950_ (.A(_04180_),
    .X(_04302_));
 sg13g2_a22oi_1 _21951_ (.Y(_04303_),
    .B1(net131),
    .B2(_04188_),
    .A2(net138),
    .A1(net208));
 sg13g2_buf_1 _21952_ (.A(_04257_),
    .X(_04304_));
 sg13g2_nand2_1 _21953_ (.Y(_04305_),
    .A(net203),
    .B(_04161_));
 sg13g2_a22oi_1 _21954_ (.Y(_04306_),
    .B1(net117),
    .B2(_03610_),
    .A2(net156),
    .A1(net185));
 sg13g2_and4_1 _21955_ (.A(_04301_),
    .B(_04303_),
    .C(_04305_),
    .D(_04306_),
    .X(_04307_));
 sg13g2_nand4_1 _21956_ (.B(_04297_),
    .C(_04298_),
    .A(_04296_),
    .Y(_04308_),
    .D(_04307_));
 sg13g2_nand2_1 _21957_ (.Y(_04309_),
    .A(_03571_),
    .B(net106));
 sg13g2_nand3_1 _21958_ (.B(_04308_),
    .C(_04309_),
    .A(net1130),
    .Y(_04310_));
 sg13g2_nand2_1 _21959_ (.Y(_04311_),
    .A(_04131_),
    .B(net281));
 sg13g2_nand2_1 _21960_ (.Y(_04312_),
    .A(_03666_),
    .B(net106));
 sg13g2_nand2b_1 _21961_ (.Y(_04313_),
    .B(net139),
    .A_N(net161));
 sg13g2_nor3_1 _21962_ (.A(net205),
    .B(_04132_),
    .C(net120),
    .Y(_04314_));
 sg13g2_o21ai_1 _21963_ (.B1(net198),
    .Y(_04315_),
    .A1(_04237_),
    .A2(_04314_));
 sg13g2_nand4_1 _21964_ (.B(_04312_),
    .C(_04313_),
    .A(_04241_),
    .Y(_04316_),
    .D(_04315_));
 sg13g2_nand2_1 _21965_ (.Y(_04317_),
    .A(net144),
    .B(net107));
 sg13g2_buf_1 _21966_ (.A(_09146_),
    .X(_04318_));
 sg13g2_nor2_1 _21967_ (.A(net990),
    .B(_04317_),
    .Y(_04319_));
 sg13g2_a21oi_1 _21968_ (.A1(_09137_),
    .A2(_04317_),
    .Y(_04320_),
    .B1(_04319_));
 sg13g2_or2_1 _21969_ (.X(_04321_),
    .B(net107),
    .A(_11808_));
 sg13g2_o21ai_1 _21970_ (.B1(_04321_),
    .Y(_04322_),
    .A1(_09883_),
    .A2(_04320_));
 sg13g2_nand4_1 _21971_ (.B(_04311_),
    .C(_04316_),
    .A(_04310_),
    .Y(_04323_),
    .D(_04322_));
 sg13g2_a21oi_1 _21972_ (.A1(_03780_),
    .A2(_04295_),
    .Y(_04324_),
    .B1(_04323_));
 sg13g2_and2_1 _21973_ (.A(_03572_),
    .B(_03659_),
    .X(_04325_));
 sg13g2_buf_1 _21974_ (.A(_04325_),
    .X(_04326_));
 sg13g2_xor2_1 _21975_ (.B(_04289_),
    .A(_04326_),
    .X(_04327_));
 sg13g2_nand2_1 _21976_ (.Y(_04328_),
    .A(_08337_),
    .B(_04327_));
 sg13g2_a21oi_2 _21977_ (.B1(_04105_),
    .Y(_04329_),
    .A2(_04230_),
    .A1(_09877_));
 sg13g2_nand4_1 _21978_ (.B(_04324_),
    .C(_04328_),
    .A(_04292_),
    .Y(_04330_),
    .D(_04329_));
 sg13g2_o21ai_1 _21979_ (.B1(_04330_),
    .Y(_04331_),
    .A1(net239),
    .A2(\cpu.ex.c_mult[12] ));
 sg13g2_nor2_1 _21980_ (.A(_08731_),
    .B(_04282_),
    .Y(_04332_));
 sg13g2_xnor2_1 _21981_ (.Y(_04333_),
    .A(_10296_),
    .B(_04332_));
 sg13g2_a22oi_1 _21982_ (.Y(_04334_),
    .B1(_04333_),
    .B2(net85),
    .A2(net35),
    .A1(net818));
 sg13g2_o21ai_1 _21983_ (.B1(_04334_),
    .Y(_00971_),
    .A1(net86),
    .A2(_04331_));
 sg13g2_and2_1 _21984_ (.A(_11430_),
    .B(_03799_),
    .X(_04335_));
 sg13g2_o21ai_1 _21985_ (.B1(_03679_),
    .Y(_04336_),
    .A1(_04326_),
    .A2(_04335_));
 sg13g2_nand2_1 _21986_ (.Y(_04337_),
    .A(net219),
    .B(_03804_));
 sg13g2_nand2_1 _21987_ (.Y(_04338_),
    .A(_03677_),
    .B(_04337_));
 sg13g2_xor2_1 _21988_ (.B(_04338_),
    .A(_04336_),
    .X(_04339_));
 sg13g2_a22oi_1 _21989_ (.Y(_04340_),
    .B1(_03798_),
    .B2(_03800_),
    .A2(_03787_),
    .A1(_03782_));
 sg13g2_xor2_1 _21990_ (.B(_04338_),
    .A(_04340_),
    .X(_04341_));
 sg13g2_nor2_2 _21991_ (.A(_03612_),
    .B(_03613_),
    .Y(_04342_));
 sg13g2_nor2_1 _21992_ (.A(net207),
    .B(net154),
    .Y(_04343_));
 sg13g2_a21oi_1 _21993_ (.A1(net207),
    .A2(_04342_),
    .Y(_04344_),
    .B1(_04343_));
 sg13g2_a22oi_1 _21994_ (.Y(_04345_),
    .B1(_04344_),
    .B2(net198),
    .A2(_04201_),
    .A1(net158));
 sg13g2_nand2_1 _21995_ (.Y(_04346_),
    .A(net226),
    .B(net279));
 sg13g2_nand3_1 _21996_ (.B(_04346_),
    .C(net187),
    .A(net205),
    .Y(_04347_));
 sg13g2_a21oi_1 _21997_ (.A1(net198),
    .A2(_04108_),
    .Y(_04348_),
    .B1(_04347_));
 sg13g2_a22oi_1 _21998_ (.Y(_04349_),
    .B1(net137),
    .B2(net132),
    .A2(net131),
    .A1(net185));
 sg13g2_a22oi_1 _21999_ (.Y(_04350_),
    .B1(_04161_),
    .B2(net184),
    .A2(net136),
    .A1(_03793_));
 sg13g2_a21oi_1 _22000_ (.A1(_03570_),
    .A2(_04247_),
    .Y(_04351_),
    .B1(_04134_));
 sg13g2_and2_1 _22001_ (.A(_11245_),
    .B(_04165_),
    .X(_04352_));
 sg13g2_a21oi_1 _22002_ (.A1(_04154_),
    .A2(net155),
    .Y(_04353_),
    .B1(_04352_));
 sg13g2_nand4_1 _22003_ (.B(_04350_),
    .C(_04351_),
    .A(_04349_),
    .Y(_04354_),
    .D(_04353_));
 sg13g2_nor2_1 _22004_ (.A(_04348_),
    .B(_04354_),
    .Y(_04355_));
 sg13g2_o21ai_1 _22005_ (.B1(_04355_),
    .Y(_04356_),
    .A1(_04159_),
    .A2(_04345_));
 sg13g2_nand3_1 _22006_ (.B(_04235_),
    .C(_04356_),
    .A(net1130),
    .Y(_04357_));
 sg13g2_mux2_1 _22007_ (.A0(net1140),
    .A1(net990),
    .S(_03815_),
    .X(_04358_));
 sg13g2_o21ai_1 _22008_ (.B1(_03811_),
    .Y(_04359_),
    .A1(net1063),
    .A2(_04358_));
 sg13g2_buf_1 _22009_ (.A(_04135_),
    .X(_04360_));
 sg13g2_a22oi_1 _22010_ (.Y(_04361_),
    .B1(net133),
    .B2(net161),
    .A2(_04360_),
    .A1(net120));
 sg13g2_inv_1 _22011_ (.Y(_04362_),
    .A(_04361_));
 sg13g2_o21ai_1 _22012_ (.B1(_09130_),
    .Y(_04363_),
    .A1(net161),
    .A2(_04136_));
 sg13g2_a21oi_1 _22013_ (.A1(_03675_),
    .A2(_04136_),
    .Y(_04364_),
    .B1(_04363_));
 sg13g2_a221oi_1 _22014_ (.B2(_09879_),
    .C1(_04364_),
    .B1(_04362_),
    .A1(_04131_),
    .Y(_04365_),
    .A2(net282));
 sg13g2_nand4_1 _22015_ (.B(_04357_),
    .C(_04359_),
    .A(_04329_),
    .Y(_04366_),
    .D(_04365_));
 sg13g2_a221oi_1 _22016_ (.B2(net744),
    .C1(_04366_),
    .B1(_04341_),
    .A1(net948),
    .Y(_04367_),
    .A2(_04339_));
 sg13g2_a21o_1 _22017_ (.A2(_11841_),
    .A1(net190),
    .B1(_04367_),
    .X(_04368_));
 sg13g2_nand2_1 _22018_ (.Y(_04369_),
    .A(net818),
    .B(_04332_));
 sg13g2_xnor2_1 _22019_ (.Y(_04370_),
    .A(_11088_),
    .B(_04369_));
 sg13g2_a22oi_1 _22020_ (.Y(_04371_),
    .B1(_04370_),
    .B2(net85),
    .A2(net35),
    .A1(net726));
 sg13g2_o21ai_1 _22021_ (.B1(_04371_),
    .Y(_00972_),
    .A1(net86),
    .A2(_04368_));
 sg13g2_nor2_1 _22022_ (.A(net218),
    .B(_04108_),
    .Y(_04372_));
 sg13g2_a21oi_1 _22023_ (.A1(net198),
    .A2(net184),
    .Y(_04373_),
    .B1(_04372_));
 sg13g2_nor3_1 _22024_ (.A(net207),
    .B(_04191_),
    .C(_04373_),
    .Y(_04374_));
 sg13g2_a22oi_1 _22025_ (.Y(_04375_),
    .B1(_04253_),
    .B2(_04174_),
    .A2(net138),
    .A1(net154));
 sg13g2_nand2_1 _22026_ (.Y(_04376_),
    .A(net122),
    .B(_04248_));
 sg13g2_nand2_1 _22027_ (.Y(_04377_),
    .A(_03770_),
    .B(net157));
 sg13g2_and2_1 _22028_ (.A(net191),
    .B(_04180_),
    .X(_04378_));
 sg13g2_a221oi_1 _22029_ (.B2(net158),
    .C1(_04378_),
    .B1(_04195_),
    .A1(net188),
    .Y(_04379_),
    .A2(_04161_));
 sg13g2_nand4_1 _22030_ (.B(_04376_),
    .C(_04377_),
    .A(_04375_),
    .Y(_04380_),
    .D(_04379_));
 sg13g2_nand3_1 _22031_ (.B(_04148_),
    .C(net187),
    .A(net204),
    .Y(_04381_));
 sg13g2_a21oi_1 _22032_ (.A1(_04196_),
    .A2(_04166_),
    .Y(_04382_),
    .B1(net118));
 sg13g2_nand2_1 _22033_ (.Y(_04383_),
    .A(net192),
    .B(net155));
 sg13g2_nand2_1 _22034_ (.Y(_04384_),
    .A(net132),
    .B(net136));
 sg13g2_nand4_1 _22035_ (.B(_04382_),
    .C(_04383_),
    .A(_04381_),
    .Y(_04385_),
    .D(_04384_));
 sg13g2_nor3_1 _22036_ (.A(_04374_),
    .B(_04380_),
    .C(_04385_),
    .Y(_04386_));
 sg13g2_nand2_1 _22037_ (.Y(_04387_),
    .A(net1130),
    .B(_04312_));
 sg13g2_nor2_1 _22038_ (.A(_03676_),
    .B(_03683_),
    .Y(_04388_));
 sg13g2_buf_1 _22039_ (.A(_04388_),
    .X(_04389_));
 sg13g2_a21oi_1 _22040_ (.A1(_03677_),
    .A2(_04335_),
    .Y(_04390_),
    .B1(_04389_));
 sg13g2_a22oi_1 _22041_ (.Y(_04391_),
    .B1(_04390_),
    .B2(_04337_),
    .A2(_04389_),
    .A1(_03677_));
 sg13g2_nand3_1 _22042_ (.B(net161),
    .C(net105),
    .A(_09879_),
    .Y(_04392_));
 sg13g2_nand2_1 _22043_ (.Y(_04393_),
    .A(_09088_),
    .B(net232));
 sg13g2_o21ai_1 _22044_ (.B1(_09136_),
    .Y(_04394_),
    .A1(_11417_),
    .A2(_03675_));
 sg13g2_nand3_1 _22045_ (.B(net201),
    .C(net140),
    .A(net990),
    .Y(_04395_));
 sg13g2_nand3b_1 _22046_ (.B(_04394_),
    .C(_04395_),
    .Y(_04396_),
    .A_N(net1131));
 sg13g2_o21ai_1 _22047_ (.B1(_04396_),
    .Y(_04397_),
    .A1(net201),
    .A2(net120));
 sg13g2_nand3_1 _22048_ (.B(_04393_),
    .C(_04397_),
    .A(_04392_),
    .Y(_04398_));
 sg13g2_a21oi_1 _22049_ (.A1(net1090),
    .A2(_04391_),
    .Y(_04399_),
    .B1(_04398_));
 sg13g2_o21ai_1 _22050_ (.B1(_04399_),
    .Y(_04400_),
    .A1(_04386_),
    .A2(_04387_));
 sg13g2_nor2_1 _22051_ (.A(_04143_),
    .B(_04400_),
    .Y(_04401_));
 sg13g2_nor2b_1 _22052_ (.A(_04389_),
    .B_N(net1090),
    .Y(_04402_));
 sg13g2_nand4_1 _22053_ (.B(_03677_),
    .C(_03679_),
    .A(_04326_),
    .Y(_04403_),
    .D(_04402_));
 sg13g2_nand4_1 _22054_ (.B(_04336_),
    .C(_04337_),
    .A(net948),
    .Y(_04404_),
    .D(_04389_));
 sg13g2_and4_1 _22055_ (.A(_04329_),
    .B(_04401_),
    .C(_04403_),
    .D(_04404_),
    .X(_04405_));
 sg13g2_o21ai_1 _22056_ (.B1(_04389_),
    .Y(_04406_),
    .A1(_03814_),
    .A2(_03815_));
 sg13g2_or3_1 _22057_ (.A(_03814_),
    .B(_03815_),
    .C(_04389_),
    .X(_04407_));
 sg13g2_a21o_1 _22058_ (.A2(_04407_),
    .A1(_04406_),
    .B1(_04294_),
    .X(_04408_));
 sg13g2_a221oi_1 _22059_ (.B2(_04408_),
    .C1(_04102_),
    .B1(_04405_),
    .A1(net190),
    .Y(_04409_),
    .A2(_11874_));
 sg13g2_nand3_1 _22060_ (.B(net726),
    .C(_04332_),
    .A(net818),
    .Y(_04410_));
 sg13g2_xnor2_1 _22061_ (.Y(_04411_),
    .A(_11093_),
    .B(_04410_));
 sg13g2_a22oi_1 _22062_ (.Y(_04412_),
    .B1(_04411_),
    .B2(net85),
    .A2(net35),
    .A1(net931));
 sg13g2_nand2b_1 _22063_ (.Y(_00973_),
    .B(_04412_),
    .A_N(_04409_));
 sg13g2_xnor2_1 _22064_ (.Y(_04413_),
    .A(net167),
    .B(net193));
 sg13g2_nand3_1 _22065_ (.B(_03683_),
    .C(_04413_),
    .A(_08337_),
    .Y(_04414_));
 sg13g2_nand2_1 _22066_ (.Y(_04415_),
    .A(_03675_),
    .B(net106));
 sg13g2_inv_1 _22067_ (.Y(_04416_),
    .A(_03577_));
 sg13g2_nor2_1 _22068_ (.A(net227),
    .B(net191),
    .Y(_04417_));
 sg13g2_a21oi_1 _22069_ (.A1(_03888_),
    .A2(_04416_),
    .Y(_04418_),
    .B1(_04417_));
 sg13g2_a22oi_1 _22070_ (.Y(_04419_),
    .B1(_04418_),
    .B2(_11448_),
    .A2(_04176_),
    .A1(net158));
 sg13g2_nand2_1 _22071_ (.Y(_04420_),
    .A(net134),
    .B(net155));
 sg13g2_a21oi_1 _22072_ (.A1(net208),
    .A2(_04193_),
    .Y(_04421_),
    .B1(_04134_));
 sg13g2_nand3_1 _22073_ (.B(_04420_),
    .C(_04421_),
    .A(_04181_),
    .Y(_04422_));
 sg13g2_nand2_1 _22074_ (.Y(_04423_),
    .A(net122),
    .B(_04165_));
 sg13g2_nand2_1 _22075_ (.Y(_04424_),
    .A(net192),
    .B(_04172_));
 sg13g2_a22oi_1 _22076_ (.Y(_04425_),
    .B1(_04247_),
    .B2(_03803_),
    .A2(net156),
    .A1(_03770_));
 sg13g2_nand3_1 _22077_ (.B(_04424_),
    .C(_04425_),
    .A(_04423_),
    .Y(_04426_));
 sg13g2_nor2_1 _22078_ (.A(_03888_),
    .B(net278),
    .Y(_04427_));
 sg13g2_nor2_1 _22079_ (.A(net238),
    .B(net279),
    .Y(_04428_));
 sg13g2_a22oi_1 _22080_ (.Y(_04429_),
    .B1(_04428_),
    .B2(net278),
    .A2(net185),
    .A1(_04427_));
 sg13g2_nor3_1 _22081_ (.A(net236),
    .B(net218),
    .C(_04429_),
    .Y(_04430_));
 sg13g2_nand2_1 _22082_ (.Y(_04431_),
    .A(net240),
    .B(_04127_));
 sg13g2_nand2_1 _22083_ (.Y(_04432_),
    .A(_03599_),
    .B(_04201_));
 sg13g2_a21oi_1 _22084_ (.A1(_04431_),
    .A2(_04432_),
    .Y(_04433_),
    .B1(_04191_));
 sg13g2_nor4_1 _22085_ (.A(_04422_),
    .B(_04426_),
    .C(_04430_),
    .D(_04433_),
    .Y(_04434_));
 sg13g2_o21ai_1 _22086_ (.B1(_04434_),
    .Y(_04435_),
    .A1(_04159_),
    .A2(_04419_));
 sg13g2_nand3_1 _22087_ (.B(_04415_),
    .C(_04435_),
    .A(_09891_),
    .Y(_04436_));
 sg13g2_nand2_1 _22088_ (.Y(_04437_),
    .A(net1140),
    .B(_03817_));
 sg13g2_nand3_1 _22089_ (.B(_11422_),
    .C(_03566_),
    .A(_04318_),
    .Y(_04438_));
 sg13g2_nand3b_1 _22090_ (.B(_04437_),
    .C(_04438_),
    .Y(_04439_),
    .A_N(_09883_));
 sg13g2_a22oi_1 _22091_ (.Y(_04440_),
    .B1(_03692_),
    .B2(_04439_),
    .A2(net233),
    .A1(net991));
 sg13g2_and4_1 _22092_ (.A(_04240_),
    .B(_04329_),
    .C(_04436_),
    .D(_04440_),
    .X(_04441_));
 sg13g2_o21ai_1 _22093_ (.B1(_08335_),
    .Y(_04442_),
    .A1(_11417_),
    .A2(_03801_));
 sg13g2_or4_1 _22094_ (.A(_03674_),
    .B(_03682_),
    .C(_04413_),
    .D(_04442_),
    .X(_04443_));
 sg13g2_and2_1 _22095_ (.A(net1090),
    .B(_04413_),
    .X(_04444_));
 sg13g2_o21ai_1 _22096_ (.B1(_04444_),
    .Y(_04445_),
    .A1(_03674_),
    .A2(_03682_));
 sg13g2_nand4_1 _22097_ (.B(_04441_),
    .C(_04443_),
    .A(_04414_),
    .Y(_04446_),
    .D(_04445_));
 sg13g2_o21ai_1 _22098_ (.B1(net461),
    .Y(_04447_),
    .A1(_11902_),
    .A2(_11904_));
 sg13g2_a221oi_1 _22099_ (.B2(_11461_),
    .C1(net239),
    .B1(_11908_),
    .A1(_11910_),
    .Y(_04448_),
    .A2(_11463_));
 sg13g2_buf_1 _22100_ (.A(_04448_),
    .X(_04449_));
 sg13g2_nand2_1 _22101_ (.Y(_04450_),
    .A(_04447_),
    .B(_04449_));
 sg13g2_nand2b_1 _22102_ (.Y(_04451_),
    .B(_04115_),
    .A_N(_04413_));
 sg13g2_a21oi_1 _22103_ (.A1(_04447_),
    .A2(_04449_),
    .Y(_04452_),
    .B1(_04451_));
 sg13g2_a22oi_1 _22104_ (.Y(_04453_),
    .B1(_04452_),
    .B2(_03810_),
    .A2(_04450_),
    .A1(_04446_));
 sg13g2_nand2_1 _22105_ (.Y(_04454_),
    .A(_03816_),
    .B(_04452_));
 sg13g2_and2_1 _22106_ (.A(_04447_),
    .B(_04449_),
    .X(_04455_));
 sg13g2_nand2_1 _22107_ (.Y(_04456_),
    .A(net744),
    .B(_04413_));
 sg13g2_or4_1 _22108_ (.A(_03810_),
    .B(_03816_),
    .C(_04455_),
    .D(_04456_),
    .X(_04457_));
 sg13g2_and3_1 _22109_ (.X(_04458_),
    .A(_04453_),
    .B(_04454_),
    .C(_04457_));
 sg13g2_or2_1 _22110_ (.X(_04459_),
    .B(_04410_),
    .A(_08840_));
 sg13g2_xnor2_1 _22111_ (.Y(_04460_),
    .A(_11087_),
    .B(_04459_));
 sg13g2_a22oi_1 _22112_ (.Y(_04461_),
    .B1(_04460_),
    .B2(net85),
    .A2(net35),
    .A1(_08397_));
 sg13g2_o21ai_1 _22113_ (.B1(_04461_),
    .Y(_00974_),
    .A1(net86),
    .A2(_04458_));
 sg13g2_and2_1 _22114_ (.A(_08423_),
    .B(_08467_),
    .X(_04462_));
 sg13g2_nand4_1 _22115_ (.B(_08388_),
    .C(_04462_),
    .A(_09208_),
    .Y(_04463_),
    .D(_11476_));
 sg13g2_and2_1 _22116_ (.A(net1076),
    .B(net97),
    .X(_04464_));
 sg13g2_o21ai_1 _22117_ (.B1(net808),
    .Y(_04465_),
    .A1(_04220_),
    .A2(_04464_));
 sg13g2_nand3_1 _22118_ (.B(net804),
    .C(net97),
    .A(net805),
    .Y(_04466_));
 sg13g2_nor2_1 _22119_ (.A(_03603_),
    .B(_03606_),
    .Y(_04467_));
 sg13g2_nand2_1 _22120_ (.Y(_04468_),
    .A(_03600_),
    .B(_03607_));
 sg13g2_xor2_1 _22121_ (.B(_04468_),
    .A(_04467_),
    .X(_04469_));
 sg13g2_xor2_1 _22122_ (.B(_04468_),
    .A(_03733_),
    .X(_04470_));
 sg13g2_nand2_1 _22123_ (.Y(_04471_),
    .A(net203),
    .B(net118));
 sg13g2_o21ai_1 _22124_ (.B1(_04471_),
    .Y(_04472_),
    .A1(net279),
    .A2(_04299_));
 sg13g2_o21ai_1 _22125_ (.B1(net990),
    .Y(_04473_),
    .A1(_03718_),
    .A2(_03719_));
 sg13g2_a21oi_1 _22126_ (.A1(_09088_),
    .A2(net200),
    .Y(_04474_),
    .B1(_04105_));
 sg13g2_nor3_1 _22127_ (.A(_09137_),
    .B(_03718_),
    .C(_03719_),
    .Y(_04475_));
 sg13g2_o21ai_1 _22128_ (.B1(_03710_),
    .Y(_04476_),
    .A1(net1131),
    .A2(_04475_));
 sg13g2_nand3_1 _22129_ (.B(_04474_),
    .C(_04476_),
    .A(_04473_),
    .Y(_04477_));
 sg13g2_a21oi_1 _22130_ (.A1(net1130),
    .A2(_04472_),
    .Y(_04478_),
    .B1(_04477_));
 sg13g2_o21ai_1 _22131_ (.B1(_04478_),
    .Y(_04479_),
    .A1(_04116_),
    .A2(_04470_));
 sg13g2_a21oi_1 _22132_ (.A1(net948),
    .A2(_04469_),
    .Y(_04480_),
    .B1(_04479_));
 sg13g2_nand2_1 _22133_ (.Y(_04481_),
    .A(net158),
    .B(_04148_));
 sg13g2_a21oi_1 _22134_ (.A1(_04145_),
    .A2(_04481_),
    .Y(_04482_),
    .B1(net189));
 sg13g2_nand3_1 _22135_ (.B(net217),
    .C(net193),
    .A(net205),
    .Y(_04483_));
 sg13g2_nand3_1 _22136_ (.B(net236),
    .C(net186),
    .A(net207),
    .Y(_04484_));
 sg13g2_a221oi_1 _22137_ (.B2(_04484_),
    .C1(_11449_),
    .B1(_04483_),
    .A1(_03714_),
    .Y(_04485_),
    .A2(_03715_));
 sg13g2_nand2_1 _22138_ (.Y(_04486_),
    .A(_03793_),
    .B(net137));
 sg13g2_nand2_1 _22139_ (.Y(_04487_),
    .A(_03577_),
    .B(_04165_));
 sg13g2_nand3_1 _22140_ (.B(net159),
    .C(net187),
    .A(net207),
    .Y(_04488_));
 sg13g2_nand2_1 _22141_ (.Y(_04489_),
    .A(net134),
    .B(net138));
 sg13g2_nand4_1 _22142_ (.B(_04487_),
    .C(_04488_),
    .A(_04486_),
    .Y(_04490_),
    .D(_04489_));
 sg13g2_nand2_1 _22143_ (.Y(_04491_),
    .A(net185),
    .B(net135));
 sg13g2_a22oi_1 _22144_ (.Y(_04492_),
    .B1(_04193_),
    .B2(net120),
    .A2(_04161_),
    .A1(net119));
 sg13g2_a22oi_1 _22145_ (.Y(_04493_),
    .B1(net117),
    .B2(net192),
    .A2(_04195_),
    .A1(net107));
 sg13g2_nand4_1 _22146_ (.B(_04491_),
    .C(_04492_),
    .A(_04384_),
    .Y(_04494_),
    .D(_04493_));
 sg13g2_nor4_1 _22147_ (.A(_04482_),
    .B(_04485_),
    .C(_04490_),
    .D(_04494_),
    .Y(_04495_));
 sg13g2_nor2_1 _22148_ (.A(net188),
    .B(_04203_),
    .Y(_04496_));
 sg13g2_nor3_1 _22149_ (.A(net856),
    .B(_04495_),
    .C(_04496_),
    .Y(_04497_));
 sg13g2_inv_1 _22150_ (.Y(_04498_),
    .A(_04497_));
 sg13g2_a22oi_1 _22151_ (.Y(_04499_),
    .B1(_04480_),
    .B2(_04498_),
    .A2(_11533_),
    .A1(net206));
 sg13g2_nand2_1 _22152_ (.Y(_04500_),
    .A(_04212_),
    .B(_04499_));
 sg13g2_nand4_1 _22153_ (.B(_04465_),
    .C(_04466_),
    .A(_04463_),
    .Y(_00975_),
    .D(_04500_));
 sg13g2_nand2_1 _22154_ (.Y(_04501_),
    .A(_03747_),
    .B(_03710_));
 sg13g2_xnor2_1 _22155_ (.Y(_04502_),
    .A(net217),
    .B(_04342_));
 sg13g2_xnor2_1 _22156_ (.Y(_04503_),
    .A(_04501_),
    .B(_04502_));
 sg13g2_and2_1 _22157_ (.A(_03600_),
    .B(_03608_),
    .X(_04504_));
 sg13g2_buf_1 _22158_ (.A(_04504_),
    .X(_04505_));
 sg13g2_xor2_1 _22159_ (.B(_04502_),
    .A(_04505_),
    .X(_04506_));
 sg13g2_nand2_1 _22160_ (.Y(_04507_),
    .A(net1140),
    .B(_03748_));
 sg13g2_o21ai_1 _22161_ (.B1(_04507_),
    .Y(_04508_),
    .A1(_09147_),
    .A2(_03748_));
 sg13g2_nand2_1 _22162_ (.Y(_04509_),
    .A(net236),
    .B(_04342_));
 sg13g2_o21ai_1 _22163_ (.B1(_04509_),
    .Y(_04510_),
    .A1(net1063),
    .A2(_04508_));
 sg13g2_a21oi_1 _22164_ (.A1(net205),
    .A2(net184),
    .Y(_04511_),
    .B1(_04428_));
 sg13g2_o21ai_1 _22165_ (.B1(_04431_),
    .Y(_04512_),
    .A1(net218),
    .A2(_04511_));
 sg13g2_nor2_1 _22166_ (.A(_09892_),
    .B(net189),
    .Y(_04513_));
 sg13g2_a221oi_1 _22167_ (.B2(_04513_),
    .C1(_04105_),
    .B1(_04512_),
    .A1(net991),
    .Y(_04514_),
    .A2(_11398_));
 sg13g2_a22oi_1 _22168_ (.Y(_04515_),
    .B1(net137),
    .B2(net132),
    .A2(net136),
    .A1(net186));
 sg13g2_a22oi_1 _22169_ (.Y(_04516_),
    .B1(_04161_),
    .B2(net140),
    .A2(_04169_),
    .A1(net107));
 sg13g2_a22oi_1 _22170_ (.Y(_04517_),
    .B1(_04195_),
    .B2(net119),
    .A2(_04193_),
    .A1(net193));
 sg13g2_a22oi_1 _22171_ (.Y(_04518_),
    .B1(net117),
    .B2(net134),
    .A2(net133),
    .A1(net154));
 sg13g2_nand4_1 _22172_ (.B(_04516_),
    .C(_04517_),
    .A(_04515_),
    .Y(_04519_),
    .D(_04518_));
 sg13g2_nand2_1 _22173_ (.Y(_04520_),
    .A(net192),
    .B(net131));
 sg13g2_a21oi_1 _22174_ (.A1(net185),
    .A2(net139),
    .Y(_04521_),
    .B1(net118));
 sg13g2_a21oi_1 _22175_ (.A1(net205),
    .A2(net218),
    .Y(_04522_),
    .B1(_04191_));
 sg13g2_o21ai_1 _22176_ (.B1(net159),
    .Y(_04523_),
    .A1(_10677_),
    .A2(_04522_));
 sg13g2_nand4_1 _22177_ (.B(_04520_),
    .C(_04521_),
    .A(_04259_),
    .Y(_04524_),
    .D(_04523_));
 sg13g2_inv_1 _22178_ (.Y(_04525_),
    .A(_03610_));
 sg13g2_a21oi_1 _22179_ (.A1(_04525_),
    .A2(net105),
    .Y(_04526_),
    .B1(net856));
 sg13g2_o21ai_1 _22180_ (.B1(_04526_),
    .Y(_04527_),
    .A1(_04519_),
    .A2(_04524_));
 sg13g2_nand3_1 _22181_ (.B(_04514_),
    .C(_04527_),
    .A(_04510_),
    .Y(_04528_));
 sg13g2_a221oi_1 _22182_ (.B2(net1090),
    .C1(_04528_),
    .B1(_04506_),
    .A1(_04122_),
    .Y(_04529_),
    .A2(_04503_));
 sg13g2_a21o_1 _22183_ (.A2(_11552_),
    .A1(_04107_),
    .B1(_04529_),
    .X(_04530_));
 sg13g2_nand2_1 _22184_ (.Y(_04531_),
    .A(net808),
    .B(net804));
 sg13g2_a21o_1 _22185_ (.A2(_04531_),
    .A1(net97),
    .B1(_04220_),
    .X(_04532_));
 sg13g2_nor2_1 _22186_ (.A(net710),
    .B(_04531_),
    .Y(_04533_));
 sg13g2_o21ai_1 _22187_ (.B1(_04217_),
    .Y(_04534_),
    .A1(_00258_),
    .A2(_04463_));
 sg13g2_a221oi_1 _22188_ (.B2(net97),
    .C1(_04534_),
    .B1(_04533_),
    .A1(net710),
    .Y(_04535_),
    .A2(_04532_));
 sg13g2_o21ai_1 _22189_ (.B1(_04535_),
    .Y(_00976_),
    .A1(net86),
    .A2(_04530_));
 sg13g2_a21oi_1 _22190_ (.A1(_03747_),
    .A2(_03710_),
    .Y(_04536_),
    .B1(net208));
 sg13g2_nand3_1 _22191_ (.B(_03747_),
    .C(_03710_),
    .A(net208),
    .Y(_04537_));
 sg13g2_o21ai_1 _22192_ (.B1(_04537_),
    .Y(_04538_),
    .A1(_11547_),
    .A2(_04536_));
 sg13g2_xnor2_1 _22193_ (.Y(_04539_),
    .A(net281),
    .B(net158));
 sg13g2_xnor2_1 _22194_ (.Y(_04540_),
    .A(_04538_),
    .B(_04539_));
 sg13g2_inv_1 _22195_ (.Y(_04541_),
    .A(_04505_));
 sg13g2_a21oi_1 _22196_ (.A1(_04342_),
    .A2(_04505_),
    .Y(_04542_),
    .B1(net217));
 sg13g2_a21oi_1 _22197_ (.A1(net188),
    .A2(_04541_),
    .Y(_04543_),
    .B1(_04542_));
 sg13g2_xnor2_1 _22198_ (.Y(_04544_),
    .A(_04539_),
    .B(_04543_));
 sg13g2_nand2_1 _22199_ (.Y(_04545_),
    .A(net281),
    .B(_03610_));
 sg13g2_nor2_1 _22200_ (.A(net990),
    .B(_04545_),
    .Y(_04546_));
 sg13g2_a21oi_1 _22201_ (.A1(_09137_),
    .A2(_04545_),
    .Y(_04547_),
    .B1(_04546_));
 sg13g2_o21ai_1 _22202_ (.B1(_03699_),
    .Y(_04548_),
    .A1(net1063),
    .A2(_04547_));
 sg13g2_a21oi_1 _22203_ (.A1(_03599_),
    .A2(_04247_),
    .Y(_04549_),
    .B1(_04134_));
 sg13g2_a22oi_1 _22204_ (.Y(_04550_),
    .B1(net139),
    .B2(net203),
    .A2(net135),
    .A1(net204));
 sg13g2_nand2_1 _22205_ (.Y(_04551_),
    .A(_04549_),
    .B(_04550_));
 sg13g2_nor2_1 _22206_ (.A(_09892_),
    .B(_04496_),
    .Y(_04552_));
 sg13g2_a221oi_1 _22207_ (.B2(_04552_),
    .C1(net206),
    .B1(_04551_),
    .A1(net991),
    .Y(_04553_),
    .A2(_11808_));
 sg13g2_nor2_1 _22208_ (.A(_11504_),
    .B(_03565_),
    .Y(_04554_));
 sg13g2_a21oi_1 _22209_ (.A1(net238),
    .A2(_03666_),
    .Y(_04555_),
    .B1(_04554_));
 sg13g2_a22oi_1 _22210_ (.Y(_04556_),
    .B1(_04555_),
    .B2(_04110_),
    .A2(_04148_),
    .A1(net120));
 sg13g2_nor2_1 _22211_ (.A(_04159_),
    .B(_04556_),
    .Y(_04557_));
 sg13g2_o21ai_1 _22212_ (.B1(net159),
    .Y(_04558_),
    .A1(_10677_),
    .A2(_04152_));
 sg13g2_a21oi_1 _22213_ (.A1(net191),
    .A2(_04165_),
    .Y(_04559_),
    .B1(_04134_));
 sg13g2_nand2_1 _22214_ (.Y(_04560_),
    .A(net185),
    .B(_04247_));
 sg13g2_and3_1 _22215_ (.X(_04561_),
    .A(_04377_),
    .B(_04559_),
    .C(_04560_));
 sg13g2_a22oi_1 _22216_ (.Y(_04562_),
    .B1(net117),
    .B2(net107),
    .A2(net136),
    .A1(net192));
 sg13g2_a22oi_1 _22217_ (.Y(_04563_),
    .B1(net135),
    .B2(net132),
    .A2(net131),
    .A1(net134));
 sg13g2_nand4_1 _22218_ (.B(_04561_),
    .C(_04562_),
    .A(_04558_),
    .Y(_04564_),
    .D(_04563_));
 sg13g2_a21oi_1 _22219_ (.A1(_04416_),
    .A2(net105),
    .Y(_04565_),
    .B1(_04141_));
 sg13g2_o21ai_1 _22220_ (.B1(_04565_),
    .Y(_04566_),
    .A1(_04557_),
    .A2(_04564_));
 sg13g2_nand3_1 _22221_ (.B(_04553_),
    .C(_04566_),
    .A(_04548_),
    .Y(_04567_));
 sg13g2_a221oi_1 _22222_ (.B2(net948),
    .C1(_04567_),
    .B1(_04544_),
    .A1(_04122_),
    .Y(_04568_),
    .A2(_04540_));
 sg13g2_a21o_1 _22223_ (.A2(_11574_),
    .A1(net190),
    .B1(_04568_),
    .X(_04569_));
 sg13g2_nand2_1 _22224_ (.Y(_04570_),
    .A(_09009_),
    .B(net820));
 sg13g2_nor2_1 _22225_ (.A(net1141),
    .B(_04570_),
    .Y(_04571_));
 sg13g2_nor3_1 _22226_ (.A(net1074),
    .B(_09317_),
    .C(_11474_),
    .Y(_04572_));
 sg13g2_buf_1 _22227_ (.A(net371),
    .X(_04573_));
 sg13g2_a21oi_1 _22228_ (.A1(net97),
    .A2(_04570_),
    .Y(_04574_),
    .B1(_04220_));
 sg13g2_nor2b_1 _22229_ (.A(_04574_),
    .B_N(net1141),
    .Y(_04575_));
 sg13g2_a221oi_1 _22230_ (.B2(_04573_),
    .C1(_04575_),
    .B1(_04572_),
    .A1(net97),
    .Y(_04576_),
    .A2(_04571_));
 sg13g2_o21ai_1 _22231_ (.B1(_04576_),
    .Y(_00977_),
    .A1(net86),
    .A2(_04569_));
 sg13g2_nand2_1 _22232_ (.Y(_04577_),
    .A(_03578_),
    .B(_03592_));
 sg13g2_nor2_1 _22233_ (.A(net277),
    .B(net158),
    .Y(_04578_));
 sg13g2_o21ai_1 _22234_ (.B1(_03611_),
    .Y(_04579_),
    .A1(_04578_),
    .A2(_04543_));
 sg13g2_xnor2_1 _22235_ (.Y(_04580_),
    .A(_04577_),
    .B(_04579_));
 sg13g2_nand2b_1 _22236_ (.Y(_04581_),
    .B(_04545_),
    .A_N(_04538_));
 sg13g2_nand2_1 _22237_ (.Y(_04582_),
    .A(_03699_),
    .B(_04581_));
 sg13g2_xnor2_1 _22238_ (.Y(_04583_),
    .A(_04577_),
    .B(_04582_));
 sg13g2_nand2_1 _22239_ (.Y(_04584_),
    .A(_04525_),
    .B(net105));
 sg13g2_a22oi_1 _22240_ (.Y(_04585_),
    .B1(net133),
    .B2(_04146_),
    .A2(net139),
    .A1(net184));
 sg13g2_nand2_1 _22241_ (.Y(_04586_),
    .A(net204),
    .B(net137));
 sg13g2_a21oi_1 _22242_ (.A1(net203),
    .A2(net135),
    .Y(_04587_),
    .B1(net118));
 sg13g2_nand3_1 _22243_ (.B(_04586_),
    .C(_04587_),
    .A(_04585_),
    .Y(_04588_));
 sg13g2_nand3_1 _22244_ (.B(_04584_),
    .C(_04588_),
    .A(net1130),
    .Y(_04589_));
 sg13g2_nor2_1 _22245_ (.A(net990),
    .B(_03754_),
    .Y(_04590_));
 sg13g2_a21oi_1 _22246_ (.A1(_09137_),
    .A2(_03754_),
    .Y(_04591_),
    .B1(_04590_));
 sg13g2_o21ai_1 _22247_ (.B1(_03762_),
    .Y(_04592_),
    .A1(net1063),
    .A2(_04591_));
 sg13g2_a21oi_1 _22248_ (.A1(net991),
    .A2(_11795_),
    .Y(_04593_),
    .B1(_04105_));
 sg13g2_o21ai_1 _22249_ (.B1(net217),
    .Y(_04594_),
    .A1(net278),
    .A2(_04176_));
 sg13g2_nor2_1 _22250_ (.A(_04240_),
    .B(_04594_),
    .Y(_04595_));
 sg13g2_nand2_1 _22251_ (.Y(_04596_),
    .A(_04154_),
    .B(net155));
 sg13g2_a22oi_1 _22252_ (.Y(_04597_),
    .B1(_04195_),
    .B2(_03565_),
    .A2(net138),
    .A1(net140));
 sg13g2_nand3_1 _22253_ (.B(_04424_),
    .C(_04597_),
    .A(_04596_),
    .Y(_04598_));
 sg13g2_a22oi_1 _22254_ (.Y(_04599_),
    .B1(_04252_),
    .B2(net119),
    .A2(_04180_),
    .A1(net122));
 sg13g2_nand2_1 _22255_ (.Y(_04600_),
    .A(net191),
    .B(net133));
 sg13g2_nand2_1 _22256_ (.Y(_04601_),
    .A(net134),
    .B(net156));
 sg13g2_nand3_1 _22257_ (.B(_04600_),
    .C(_04601_),
    .A(_04599_),
    .Y(_04602_));
 sg13g2_nand2_1 _22258_ (.Y(_04603_),
    .A(net227),
    .B(_03641_));
 sg13g2_a22oi_1 _22259_ (.Y(_04604_),
    .B1(_04603_),
    .B2(net226),
    .A2(net159),
    .A1(_04144_));
 sg13g2_nor2_1 _22260_ (.A(net189),
    .B(_04604_),
    .Y(_04605_));
 sg13g2_nor4_1 _22261_ (.A(_04595_),
    .B(_04598_),
    .C(_04602_),
    .D(_04605_),
    .Y(_04606_));
 sg13g2_a21oi_1 _22262_ (.A1(_03649_),
    .A2(net105),
    .Y(_04607_),
    .B1(net856));
 sg13g2_nand2b_1 _22263_ (.Y(_04608_),
    .B(_04607_),
    .A_N(_04606_));
 sg13g2_nand4_1 _22264_ (.B(_04592_),
    .C(_04593_),
    .A(_04589_),
    .Y(_04609_),
    .D(_04608_));
 sg13g2_a221oi_1 _22265_ (.B2(_04122_),
    .C1(_04609_),
    .B1(_04583_),
    .A1(net1090),
    .Y(_04610_),
    .A2(_04580_));
 sg13g2_a21o_1 _22266_ (.A2(_11586_),
    .A1(net190),
    .B1(_04610_),
    .X(_04611_));
 sg13g2_buf_1 _22267_ (.A(_08671_),
    .X(_04612_));
 sg13g2_xnor2_1 _22268_ (.Y(_04613_),
    .A(_00280_),
    .B(_04279_));
 sg13g2_a22oi_1 _22269_ (.Y(_04614_),
    .B1(_04613_),
    .B2(_04284_),
    .A2(net35),
    .A1(net989));
 sg13g2_o21ai_1 _22270_ (.B1(_04614_),
    .Y(_00978_),
    .A1(_04103_),
    .A2(_04611_));
 sg13g2_a22oi_1 _22271_ (.Y(_04615_),
    .B1(net133),
    .B2(_03767_),
    .A2(net156),
    .A1(net122));
 sg13g2_a22oi_1 _22272_ (.Y(_04616_),
    .B1(_04252_),
    .B2(net140),
    .A2(_04168_),
    .A1(_03565_));
 sg13g2_and2_1 _22273_ (.A(_04615_),
    .B(_04616_),
    .X(_04617_));
 sg13g2_a22oi_1 _22274_ (.Y(_04618_),
    .B1(net157),
    .B2(net134),
    .A2(net131),
    .A1(net119));
 sg13g2_nand4_1 _22275_ (.B(_04383_),
    .C(_04617_),
    .A(_04297_),
    .Y(_04619_),
    .D(_04618_));
 sg13g2_a21o_1 _22276_ (.A2(_04619_),
    .A1(_09879_),
    .B1(_09130_),
    .X(_04620_));
 sg13g2_a21oi_1 _22277_ (.A1(net205),
    .A2(_10589_),
    .Y(_04621_),
    .B1(_11547_));
 sg13g2_o21ai_1 _22278_ (.B1(net193),
    .Y(_04622_),
    .A1(_10677_),
    .A2(_04621_));
 sg13g2_nor2b_1 _22279_ (.A(_04619_),
    .B_N(_04622_),
    .Y(_04623_));
 sg13g2_a21oi_1 _22280_ (.A1(_03628_),
    .A2(net106),
    .Y(_04624_),
    .B1(_04623_));
 sg13g2_nand2_1 _22281_ (.Y(_04625_),
    .A(_03594_),
    .B(_03619_));
 sg13g2_nand2_1 _22282_ (.Y(_04626_),
    .A(net276),
    .B(_03622_));
 sg13g2_nand2_1 _22283_ (.Y(_04627_),
    .A(net232),
    .B(_03649_));
 sg13g2_nand2_1 _22284_ (.Y(_04628_),
    .A(_04626_),
    .B(_04627_));
 sg13g2_xor2_1 _22285_ (.B(_04628_),
    .A(_04625_),
    .X(_04629_));
 sg13g2_nor2_1 _22286_ (.A(net990),
    .B(_04227_),
    .Y(_04630_));
 sg13g2_a21oi_1 _22287_ (.A1(_09137_),
    .A2(_04227_),
    .Y(_04631_),
    .B1(_04630_));
 sg13g2_nor2_1 _22288_ (.A(net1131),
    .B(_04631_),
    .Y(_04632_));
 sg13g2_a21oi_1 _22289_ (.A1(_09088_),
    .A2(_10486_),
    .Y(_04633_),
    .B1(_04105_));
 sg13g2_o21ai_1 _22290_ (.B1(_04633_),
    .Y(_04634_),
    .A1(_04228_),
    .A2(_04632_));
 sg13g2_nor2_1 _22291_ (.A(_04525_),
    .B(_04299_),
    .Y(_04635_));
 sg13g2_a221oi_1 _22292_ (.B2(net203),
    .C1(_04635_),
    .B1(net137),
    .A1(net184),
    .Y(_04636_),
    .A2(net135));
 sg13g2_a221oi_1 _22293_ (.B2(net188),
    .C1(net105),
    .B1(net139),
    .A1(net204),
    .Y(_04637_),
    .A2(net136));
 sg13g2_o21ai_1 _22294_ (.B1(net1130),
    .Y(_04638_),
    .A1(net154),
    .A2(_04203_));
 sg13g2_a21o_1 _22295_ (.A2(_04637_),
    .A1(_04636_),
    .B1(_04638_),
    .X(_04639_));
 sg13g2_nand2b_1 _22296_ (.Y(_04640_),
    .B(_04639_),
    .A_N(_04634_));
 sg13g2_a221oi_1 _22297_ (.B2(net1090),
    .C1(_04640_),
    .B1(_04629_),
    .A1(_04620_),
    .Y(_04641_),
    .A2(_04624_));
 sg13g2_xnor2_1 _22298_ (.Y(_04642_),
    .A(_04226_),
    .B(_04628_));
 sg13g2_nand2_1 _22299_ (.Y(_04643_),
    .A(_04122_),
    .B(_04642_));
 sg13g2_a22oi_1 _22300_ (.Y(_04644_),
    .B1(_04641_),
    .B2(_04643_),
    .A2(_11603_),
    .A1(net206));
 sg13g2_inv_1 _22301_ (.Y(_04645_),
    .A(_04644_));
 sg13g2_buf_1 _22302_ (.A(_08718_),
    .X(_04646_));
 sg13g2_nand2_1 _22303_ (.Y(_04647_),
    .A(_08671_),
    .B(_04279_));
 sg13g2_xnor2_1 _22304_ (.Y(_04648_),
    .A(_10816_),
    .B(_04647_));
 sg13g2_a22oi_1 _22305_ (.Y(_04649_),
    .B1(_04648_),
    .B2(net85),
    .A2(net35),
    .A1(net988));
 sg13g2_o21ai_1 _22306_ (.B1(_04649_),
    .Y(_00979_),
    .A1(net86),
    .A2(_04645_));
 sg13g2_nand2b_1 _22307_ (.Y(_04650_),
    .B(_04294_),
    .A_N(_09133_));
 sg13g2_nand3_1 _22308_ (.B(_03619_),
    .C(_04627_),
    .A(_03594_),
    .Y(_04651_));
 sg13g2_nand2_1 _22309_ (.Y(_04652_),
    .A(_04626_),
    .B(_04651_));
 sg13g2_xor2_1 _22310_ (.B(_04652_),
    .A(_04225_),
    .X(_04653_));
 sg13g2_nor2_1 _22311_ (.A(net132),
    .B(_04203_),
    .Y(_04654_));
 sg13g2_a21oi_1 _22312_ (.A1(_03770_),
    .A2(_04248_),
    .Y(_04655_),
    .B1(_04134_));
 sg13g2_o21ai_1 _22313_ (.B1(net159),
    .Y(_04656_),
    .A1(_11539_),
    .A2(_10677_));
 sg13g2_a22oi_1 _22314_ (.Y(_04657_),
    .B1(net157),
    .B2(_03670_),
    .A2(net156),
    .A1(_03803_));
 sg13g2_a221oi_1 _22315_ (.B2(_03570_),
    .C1(_04352_),
    .B1(_04185_),
    .A1(_03661_),
    .Y(_04658_),
    .A2(_04180_));
 sg13g2_nand4_1 _22316_ (.B(_04656_),
    .C(_04657_),
    .A(_04655_),
    .Y(_04659_),
    .D(_04658_));
 sg13g2_a21o_1 _22317_ (.A2(net117),
    .A1(_03567_),
    .B1(_04659_),
    .X(_04660_));
 sg13g2_a22oi_1 _22318_ (.Y(_04661_),
    .B1(_04660_),
    .B2(_09879_),
    .A2(_04659_),
    .A1(_09130_));
 sg13g2_a22oi_1 _22319_ (.Y(_04662_),
    .B1(_04173_),
    .B2(net184),
    .A2(net135),
    .A1(net188));
 sg13g2_a21oi_1 _22320_ (.A1(net204),
    .A2(net131),
    .Y(_04663_),
    .B1(net118));
 sg13g2_a22oi_1 _22321_ (.Y(_04664_),
    .B1(net133),
    .B2(net154),
    .A2(_04184_),
    .A1(net203));
 sg13g2_nand4_1 _22322_ (.B(_04662_),
    .C(_04663_),
    .A(_04167_),
    .Y(_04665_),
    .D(_04664_));
 sg13g2_a21oi_1 _22323_ (.A1(_03649_),
    .A2(net105),
    .Y(_04666_),
    .B1(_09892_));
 sg13g2_mux2_1 _22324_ (.A0(net990),
    .A1(net1140),
    .S(_03744_),
    .X(_04667_));
 sg13g2_nor2_1 _22325_ (.A(net1131),
    .B(_04667_),
    .Y(_04668_));
 sg13g2_a21oi_1 _22326_ (.A1(net234),
    .A2(_03628_),
    .Y(_04669_),
    .B1(_04668_));
 sg13g2_a221oi_1 _22327_ (.B2(_04666_),
    .C1(_04669_),
    .B1(_04665_),
    .A1(net991),
    .Y(_04670_),
    .A2(net167));
 sg13g2_o21ai_1 _22328_ (.B1(_04670_),
    .Y(_04671_),
    .A1(_04654_),
    .A2(_04661_));
 sg13g2_a221oi_1 _22329_ (.B2(net1090),
    .C1(_04671_),
    .B1(_04653_),
    .A1(_04230_),
    .Y(_04672_),
    .A2(_04650_));
 sg13g2_a22oi_1 _22330_ (.Y(_04673_),
    .B1(_04329_),
    .B2(_04672_),
    .A2(_11635_),
    .A1(_04107_));
 sg13g2_nand2_1 _22331_ (.Y(_04674_),
    .A(_04212_),
    .B(_04673_));
 sg13g2_buf_1 _22332_ (.A(_08699_),
    .X(_04675_));
 sg13g2_nand3_1 _22333_ (.B(_08718_),
    .C(_04279_),
    .A(_08671_),
    .Y(_04676_));
 sg13g2_xnor2_1 _22334_ (.Y(_04677_),
    .A(_11253_),
    .B(_04676_));
 sg13g2_a22oi_1 _22335_ (.Y(_04678_),
    .B1(_04677_),
    .B2(_04284_),
    .A2(_04221_),
    .A1(net987));
 sg13g2_nand2_1 _22336_ (.Y(_00980_),
    .A(_04674_),
    .B(_04678_));
 sg13g2_a221oi_1 _22337_ (.B2(net119),
    .C1(_04300_),
    .B1(net157),
    .A1(net140),
    .Y(_04679_),
    .A2(_04183_));
 sg13g2_a22oi_1 _22338_ (.Y(_04680_),
    .B1(_04187_),
    .B2(net107),
    .A2(_04302_),
    .A1(net193));
 sg13g2_nand4_1 _22339_ (.B(_04656_),
    .C(_04679_),
    .A(_04382_),
    .Y(_04681_),
    .D(_04680_));
 sg13g2_a21oi_1 _22340_ (.A1(_03637_),
    .A2(_04360_),
    .Y(_04682_),
    .B1(net856));
 sg13g2_nand2_1 _22341_ (.Y(_04683_),
    .A(net204),
    .B(_04253_));
 sg13g2_a22oi_1 _22342_ (.Y(_04684_),
    .B1(_04173_),
    .B2(net188),
    .A2(net131),
    .A1(_04304_));
 sg13g2_nand2_1 _22343_ (.Y(_04685_),
    .A(_04487_),
    .B(_04560_));
 sg13g2_a221oi_1 _22344_ (.B2(_04163_),
    .C1(_04685_),
    .B1(net155),
    .A1(_04200_),
    .Y(_04686_),
    .A2(_04184_));
 sg13g2_nand4_1 _22345_ (.B(_04683_),
    .C(_04684_),
    .A(_04203_),
    .Y(_04687_),
    .D(_04686_));
 sg13g2_a21oi_1 _22346_ (.A1(_03628_),
    .A2(net105),
    .Y(_04688_),
    .B1(_09892_));
 sg13g2_nor2_1 _22347_ (.A(net216),
    .B(net160),
    .Y(_04689_));
 sg13g2_mux2_1 _22348_ (.A0(net1140),
    .A1(_09146_),
    .S(_04689_),
    .X(_04690_));
 sg13g2_nand2_1 _22349_ (.Y(_04691_),
    .A(net216),
    .B(net160));
 sg13g2_o21ai_1 _22350_ (.B1(_04691_),
    .Y(_04692_),
    .A1(_09882_),
    .A2(_04690_));
 sg13g2_o21ai_1 _22351_ (.B1(_04692_),
    .Y(_04693_),
    .A1(_09089_),
    .A2(_11449_));
 sg13g2_a221oi_1 _22352_ (.B2(_04688_),
    .C1(_04693_),
    .B1(_04687_),
    .A1(_04681_),
    .Y(_04694_),
    .A2(_04682_));
 sg13g2_xnor2_1 _22353_ (.Y(_04695_),
    .A(net216),
    .B(net160));
 sg13g2_nand3_1 _22354_ (.B(_04626_),
    .C(_04651_),
    .A(_03640_),
    .Y(_04696_));
 sg13g2_buf_1 _22355_ (.A(_04696_),
    .X(_04697_));
 sg13g2_nand3_1 _22356_ (.B(_04695_),
    .C(_04697_),
    .A(_04223_),
    .Y(_04698_));
 sg13g2_a21o_1 _22357_ (.A2(_04697_),
    .A1(_04223_),
    .B1(_04695_),
    .X(_04699_));
 sg13g2_nand3_1 _22358_ (.B(_04698_),
    .C(_04699_),
    .A(_08335_),
    .Y(_04700_));
 sg13g2_nand3_1 _22359_ (.B(_04694_),
    .C(_04700_),
    .A(_04231_),
    .Y(_04701_));
 sg13g2_nand3_1 _22360_ (.B(_03741_),
    .C(_03744_),
    .A(_03773_),
    .Y(_04702_));
 sg13g2_xnor2_1 _22361_ (.Y(_04703_),
    .A(_04702_),
    .B(_04695_));
 sg13g2_nand2b_1 _22362_ (.Y(_04704_),
    .B(net744),
    .A_N(_04703_));
 sg13g2_a21o_1 _22363_ (.A2(_04704_),
    .A1(_04701_),
    .B1(_04106_),
    .X(_04705_));
 sg13g2_o21ai_1 _22364_ (.B1(_04705_),
    .Y(_04706_),
    .A1(net239),
    .A2(\cpu.ex.c_mult[8] ));
 sg13g2_xnor2_1 _22365_ (.Y(_04707_),
    .A(_10488_),
    .B(_04280_));
 sg13g2_a22oi_1 _22366_ (.Y(_04708_),
    .B1(_04707_),
    .B2(net85),
    .A2(_04220_),
    .A1(\cpu.ex.pc[8] ));
 sg13g2_o21ai_1 _22367_ (.B1(_04708_),
    .Y(_00981_),
    .A1(_04103_),
    .A2(_04706_));
 sg13g2_or2_1 _22368_ (.X(_04709_),
    .B(_03638_),
    .A(_03632_));
 sg13g2_buf_1 _22369_ (.A(_04709_),
    .X(_04710_));
 sg13g2_a22oi_1 _22370_ (.Y(_04711_),
    .B1(_04223_),
    .B2(_04697_),
    .A2(net132),
    .A1(net216));
 sg13g2_a21oi_1 _22371_ (.A1(net169),
    .A2(net160),
    .Y(_04712_),
    .B1(_04711_));
 sg13g2_xnor2_1 _22372_ (.Y(_04713_),
    .A(_04710_),
    .B(_04712_));
 sg13g2_a21oi_1 _22373_ (.A1(_04702_),
    .A2(_04691_),
    .Y(_04714_),
    .B1(_04689_));
 sg13g2_xor2_1 _22374_ (.B(_04710_),
    .A(_04714_),
    .X(_04715_));
 sg13g2_nand2_1 _22375_ (.Y(_04716_),
    .A(_04245_),
    .B(_04169_));
 sg13g2_a22oi_1 _22376_ (.Y(_04717_),
    .B1(net117),
    .B2(net203),
    .A2(net135),
    .A1(net154));
 sg13g2_nand2_1 _22377_ (.Y(_04718_),
    .A(_03599_),
    .B(_04180_));
 sg13g2_nand2_1 _22378_ (.Y(_04719_),
    .A(_04600_),
    .B(_04718_));
 sg13g2_a221oi_1 _22379_ (.B2(net158),
    .C1(_04719_),
    .B1(net137),
    .A1(_04146_),
    .Y(_04720_),
    .A2(net136));
 sg13g2_nand4_1 _22380_ (.B(_04716_),
    .C(_04717_),
    .A(_04521_),
    .Y(_04721_),
    .D(_04720_));
 sg13g2_a21oi_1 _22381_ (.A1(_03641_),
    .A2(net106),
    .Y(_04722_),
    .B1(_09892_));
 sg13g2_nand2_1 _22382_ (.Y(_04723_),
    .A(_03662_),
    .B(_04172_));
 sg13g2_a22oi_1 _22383_ (.Y(_04724_),
    .B1(net155),
    .B2(_03803_),
    .A2(_04183_),
    .A1(_03565_));
 sg13g2_nand4_1 _22384_ (.B(_04423_),
    .C(_04723_),
    .A(_04351_),
    .Y(_04725_),
    .D(_04724_));
 sg13g2_a21oi_1 _22385_ (.A1(_09879_),
    .A2(_04725_),
    .Y(_04726_),
    .B1(_09130_));
 sg13g2_a21oi_1 _22386_ (.A1(_03567_),
    .A2(_04302_),
    .Y(_04727_),
    .B1(_04725_));
 sg13g2_o21ai_1 _22387_ (.B1(_04656_),
    .Y(_04728_),
    .A1(_04726_),
    .A2(_04727_));
 sg13g2_nor2_1 _22388_ (.A(net220),
    .B(net186),
    .Y(_04729_));
 sg13g2_nor2_1 _22389_ (.A(_04318_),
    .B(_03771_),
    .Y(_04730_));
 sg13g2_a21oi_1 _22390_ (.A1(_09137_),
    .A2(_03771_),
    .Y(_04731_),
    .B1(_04730_));
 sg13g2_nor2_1 _22391_ (.A(net1131),
    .B(_04731_),
    .Y(_04732_));
 sg13g2_nand2_1 _22392_ (.Y(_04733_),
    .A(_09088_),
    .B(_03889_));
 sg13g2_o21ai_1 _22393_ (.B1(_04733_),
    .Y(_04734_),
    .A1(_04729_),
    .A2(_04732_));
 sg13g2_a221oi_1 _22394_ (.B2(_04263_),
    .C1(_04734_),
    .B1(_04728_),
    .A1(_04721_),
    .Y(_04735_),
    .A2(_04722_));
 sg13g2_o21ai_1 _22395_ (.B1(_04735_),
    .Y(_04736_),
    .A1(_04294_),
    .A2(_04715_));
 sg13g2_a221oi_1 _22396_ (.B2(net948),
    .C1(_04736_),
    .B1(_04713_),
    .A1(_09877_),
    .Y(_04737_),
    .A2(_04230_));
 sg13g2_nor4_1 _22397_ (.A(_11469_),
    .B(_11665_),
    .C(_11684_),
    .D(_11687_),
    .Y(_04738_));
 sg13g2_a21oi_1 _22398_ (.A1(_11469_),
    .A2(_04737_),
    .Y(_04739_),
    .B1(_04738_));
 sg13g2_nand2_1 _22399_ (.Y(_04740_),
    .A(_04212_),
    .B(_04739_));
 sg13g2_buf_1 _22400_ (.A(_08679_),
    .X(_04741_));
 sg13g2_xnor2_1 _22401_ (.Y(_04742_),
    .A(_10547_),
    .B(_04281_));
 sg13g2_a22oi_1 _22402_ (.Y(_04743_),
    .B1(_04742_),
    .B2(net85),
    .A2(net35),
    .A1(net986));
 sg13g2_nand2_1 _22403_ (.Y(_00982_),
    .A(_04740_),
    .B(_04743_));
 sg13g2_a21oi_1 _22404_ (.A1(_03889_),
    .A2(net278),
    .Y(_04744_),
    .B1(net217));
 sg13g2_nor2_1 _22405_ (.A(net217),
    .B(_11447_),
    .Y(_04745_));
 sg13g2_o21ai_1 _22406_ (.B1(_04745_),
    .Y(_04746_),
    .A1(_10589_),
    .A2(net193));
 sg13g2_o21ai_1 _22407_ (.B1(_04746_),
    .Y(_04747_),
    .A1(_11518_),
    .A2(_04240_));
 sg13g2_nand2_1 _22408_ (.Y(_04748_),
    .A(net140),
    .B(net155));
 sg13g2_nand2_1 _22409_ (.Y(_04749_),
    .A(_04376_),
    .B(_04748_));
 sg13g2_a221oi_1 _22410_ (.B2(_04144_),
    .C1(_04749_),
    .B1(_04747_),
    .A1(net119),
    .Y(_04750_),
    .A2(net139));
 sg13g2_o21ai_1 _22411_ (.B1(_04750_),
    .Y(_04751_),
    .A1(_04240_),
    .A2(_04744_));
 sg13g2_a21oi_1 _22412_ (.A1(_03571_),
    .A2(net106),
    .Y(_04752_),
    .B1(net856));
 sg13g2_nand3_1 _22413_ (.B(_03644_),
    .C(_03656_),
    .A(_03655_),
    .Y(_04753_));
 sg13g2_xnor2_1 _22414_ (.Y(_04754_),
    .A(_03696_),
    .B(_10807_));
 sg13g2_xor2_1 _22415_ (.B(_04754_),
    .A(_04753_),
    .X(_04755_));
 sg13g2_nand2_1 _22416_ (.Y(_04756_),
    .A(net204),
    .B(_04195_));
 sg13g2_nand2_1 _22417_ (.Y(_04757_),
    .A(_04559_),
    .B(_04756_));
 sg13g2_nand2_1 _22418_ (.Y(_04758_),
    .A(_04250_),
    .B(net133));
 sg13g2_a22oi_1 _22419_ (.Y(_04759_),
    .B1(net156),
    .B2(_04163_),
    .A2(net131),
    .A1(_03616_));
 sg13g2_a22oi_1 _22420_ (.Y(_04760_),
    .B1(net117),
    .B2(_04200_),
    .A2(net157),
    .A1(net154));
 sg13g2_a22oi_1 _22421_ (.Y(_04761_),
    .B1(_04186_),
    .B2(_04174_),
    .A2(net138),
    .A1(_04304_));
 sg13g2_nand4_1 _22422_ (.B(_04759_),
    .C(_04760_),
    .A(_04758_),
    .Y(_04762_),
    .D(_04761_));
 sg13g2_nor2_1 _22423_ (.A(_04757_),
    .B(_04762_),
    .Y(_04763_));
 sg13g2_o21ai_1 _22424_ (.B1(net1130),
    .Y(_04764_),
    .A1(net186),
    .A2(_04203_));
 sg13g2_mux2_1 _22425_ (.A0(_09147_),
    .A1(_09137_),
    .S(_04271_),
    .X(_04765_));
 sg13g2_nand2b_1 _22426_ (.Y(_04766_),
    .B(_04765_),
    .A_N(_09882_));
 sg13g2_a22oi_1 _22427_ (.Y(_04767_),
    .B1(_03790_),
    .B2(_04766_),
    .A2(_11518_),
    .A1(_09088_));
 sg13g2_o21ai_1 _22428_ (.B1(_04767_),
    .Y(_04768_),
    .A1(_04763_),
    .A2(_04764_));
 sg13g2_a221oi_1 _22429_ (.B2(_08336_),
    .C1(_04768_),
    .B1(_04755_),
    .A1(_04751_),
    .Y(_04769_),
    .A2(_04752_));
 sg13g2_xnor2_1 _22430_ (.Y(_04770_),
    .A(_03780_),
    .B(_04754_));
 sg13g2_a221oi_1 _22431_ (.B2(net744),
    .C1(net190),
    .B1(_04770_),
    .A1(_04231_),
    .Y(_04771_),
    .A2(_04769_));
 sg13g2_a21o_1 _22432_ (.A2(\cpu.ex.c_mult[10] ),
    .A1(net190),
    .B1(_04771_),
    .X(_04772_));
 sg13g2_inv_1 _22433_ (.Y(_04773_),
    .A(_04772_));
 sg13g2_buf_1 _22434_ (.A(_08688_),
    .X(_04774_));
 sg13g2_nand2_1 _22435_ (.Y(_04775_),
    .A(_08679_),
    .B(_04281_));
 sg13g2_xnor2_1 _22436_ (.Y(_04776_),
    .A(_10389_),
    .B(_04775_));
 sg13g2_a22oi_1 _22437_ (.Y(_04777_),
    .B1(_04776_),
    .B2(_04209_),
    .A2(_04220_),
    .A1(net985));
 sg13g2_o21ai_1 _22438_ (.B1(_04777_),
    .Y(_00983_),
    .A1(_04102_),
    .A2(_04773_));
 sg13g2_mux2_1 _22439_ (.A0(_10200_),
    .A1(\cpu.dec.r_set_cc ),
    .S(_03557_),
    .X(_00986_));
 sg13g2_buf_1 _22440_ (.A(_00240_),
    .X(_04778_));
 sg13g2_nor4_1 _22441_ (.A(net1126),
    .B(_10192_),
    .C(_04778_),
    .D(_03492_),
    .Y(_04779_));
 sg13g2_buf_2 _22442_ (.A(_04779_),
    .X(_04780_));
 sg13g2_buf_1 _22443_ (.A(_04780_),
    .X(_04781_));
 sg13g2_mux2_1 _22444_ (.A0(_10628_),
    .A1(_03508_),
    .S(net597),
    .X(_00987_));
 sg13g2_buf_1 _22445_ (.A(net1122),
    .X(_04782_));
 sg13g2_mux2_1 _22446_ (.A0(_10359_),
    .A1(_04782_),
    .S(_04781_),
    .X(_00988_));
 sg13g2_mux2_1 _22447_ (.A0(_10329_),
    .A1(net542),
    .S(net597),
    .X(_00989_));
 sg13g2_mux2_1 _22448_ (.A0(\cpu.ex.r_sp[13] ),
    .A1(net489),
    .S(net597),
    .X(_00990_));
 sg13g2_buf_1 _22449_ (.A(net605),
    .X(_04783_));
 sg13g2_mux2_1 _22450_ (.A0(_10456_),
    .A1(_04783_),
    .S(_04781_),
    .X(_00991_));
 sg13g2_mux2_1 _22451_ (.A0(_10440_),
    .A1(net746),
    .S(net597),
    .X(_00992_));
 sg13g2_mux2_1 _22452_ (.A0(_10574_),
    .A1(net453),
    .S(net597),
    .X(_00993_));
 sg13g2_mux2_1 _22453_ (.A0(_10594_),
    .A1(_03511_),
    .S(net597),
    .X(_00994_));
 sg13g2_mux2_1 _22454_ (.A0(_10768_),
    .A1(net409),
    .S(net597),
    .X(_00995_));
 sg13g2_mux2_1 _22455_ (.A0(_10753_),
    .A1(net667),
    .S(net597),
    .X(_00996_));
 sg13g2_buf_1 _22456_ (.A(net872),
    .X(_04784_));
 sg13g2_mux2_1 _22457_ (.A0(_10685_),
    .A1(_04784_),
    .S(_04780_),
    .X(_00997_));
 sg13g2_mux2_1 _22458_ (.A0(_10722_),
    .A1(net992),
    .S(_04780_),
    .X(_00998_));
 sg13g2_mux2_1 _22459_ (.A0(_10505_),
    .A1(net857),
    .S(_04780_),
    .X(_00999_));
 sg13g2_mux2_1 _22460_ (.A0(_10530_),
    .A1(net859),
    .S(_04780_),
    .X(_01000_));
 sg13g2_mux2_1 _22461_ (.A0(_10403_),
    .A1(net858),
    .S(_04780_),
    .X(_01001_));
 sg13g2_or2_1 _22462_ (.X(_04785_),
    .B(_03492_),
    .A(_10194_));
 sg13g2_buf_2 _22463_ (.A(_04785_),
    .X(_04786_));
 sg13g2_buf_1 _22464_ (.A(_04786_),
    .X(_04787_));
 sg13g2_nor2_1 _22465_ (.A(net823),
    .B(_04778_),
    .Y(_04788_));
 sg13g2_nand2_1 _22466_ (.Y(_04789_),
    .A(net861),
    .B(_04788_));
 sg13g2_nor2b_1 _22467_ (.A(net1052),
    .B_N(\cpu.ex.r_wb_swapsp ),
    .Y(_04790_));
 sg13g2_a21oi_1 _22468_ (.A1(net994),
    .A2(net1052),
    .Y(_04791_),
    .B1(_04790_));
 sg13g2_or4_1 _22469_ (.A(_10190_),
    .B(_04778_),
    .C(_03492_),
    .D(_04791_),
    .X(_04792_));
 sg13g2_buf_1 _22470_ (.A(_04792_),
    .X(_04793_));
 sg13g2_buf_1 _22471_ (.A(net596),
    .X(_04794_));
 sg13g2_nand2_1 _22472_ (.Y(_04795_),
    .A(\cpu.ex.r_stmp[0] ),
    .B(_04794_));
 sg13g2_o21ai_1 _22473_ (.B1(_04795_),
    .Y(_01002_),
    .A1(_04787_),
    .A2(_04789_));
 sg13g2_buf_1 _22474_ (.A(net596),
    .X(_04796_));
 sg13g2_buf_1 _22475_ (.A(_04786_),
    .X(_04797_));
 sg13g2_nor2_1 _22476_ (.A(_11225_),
    .B(net534),
    .Y(_04798_));
 sg13g2_a21oi_1 _22477_ (.A1(_10403_),
    .A2(net537),
    .Y(_04799_),
    .B1(_04798_));
 sg13g2_nand2_1 _22478_ (.Y(_04800_),
    .A(\cpu.ex.r_stmp[10] ),
    .B(net536));
 sg13g2_o21ai_1 _22479_ (.B1(_04800_),
    .Y(_01003_),
    .A1(net535),
    .A2(_04799_));
 sg13g2_mux2_1 _22480_ (.A0(net1122),
    .A1(_10359_),
    .S(_04786_),
    .X(_04801_));
 sg13g2_nor2_1 _22481_ (.A(net596),
    .B(_04801_),
    .Y(_04802_));
 sg13g2_a21oi_1 _22482_ (.A1(_11189_),
    .A2(net535),
    .Y(_01004_),
    .B1(_04802_));
 sg13g2_mux2_1 _22483_ (.A0(net617),
    .A1(_10329_),
    .S(net534),
    .X(_04803_));
 sg13g2_mux2_1 _22484_ (.A0(_04803_),
    .A1(\cpu.ex.r_stmp[12] ),
    .S(net536),
    .X(_01005_));
 sg13g2_mux2_1 _22485_ (.A0(net577),
    .A1(\cpu.ex.r_sp[13] ),
    .S(net534),
    .X(_04804_));
 sg13g2_mux2_1 _22486_ (.A0(_04804_),
    .A1(\cpu.ex.r_stmp[13] ),
    .S(net536),
    .X(_01006_));
 sg13g2_mux2_1 _22487_ (.A0(net688),
    .A1(_10456_),
    .S(_04797_),
    .X(_04805_));
 sg13g2_mux2_1 _22488_ (.A0(_04805_),
    .A1(\cpu.ex.r_stmp[14] ),
    .S(net536),
    .X(_01007_));
 sg13g2_nor2_1 _22489_ (.A(net699),
    .B(net534),
    .Y(_04806_));
 sg13g2_a21oi_1 _22490_ (.A1(_10440_),
    .A2(net537),
    .Y(_04807_),
    .B1(_04806_));
 sg13g2_nand2_1 _22491_ (.Y(_04808_),
    .A(\cpu.ex.r_stmp[15] ),
    .B(net536));
 sg13g2_o21ai_1 _22492_ (.B1(_04808_),
    .Y(_01008_),
    .A1(net535),
    .A2(_04807_));
 sg13g2_nor2_1 _22493_ (.A(net622),
    .B(net534),
    .Y(_04809_));
 sg13g2_a21oi_1 _22494_ (.A1(_10628_),
    .A2(net537),
    .Y(_04810_),
    .B1(_04809_));
 sg13g2_nand2_1 _22495_ (.Y(_04811_),
    .A(\cpu.ex.r_stmp[1] ),
    .B(net536));
 sg13g2_o21ai_1 _22496_ (.B1(_04811_),
    .Y(_01009_),
    .A1(net535),
    .A2(_04810_));
 sg13g2_nor2_1 _22497_ (.A(_03835_),
    .B(net534),
    .Y(_04812_));
 sg13g2_a21oi_1 _22498_ (.A1(_10574_),
    .A2(net537),
    .Y(_04813_),
    .B1(_04812_));
 sg13g2_nand2_1 _22499_ (.Y(_04814_),
    .A(\cpu.ex.r_stmp[2] ),
    .B(net536));
 sg13g2_o21ai_1 _22500_ (.B1(_04814_),
    .Y(_01010_),
    .A1(net535),
    .A2(_04813_));
 sg13g2_nor2_1 _22501_ (.A(_09241_),
    .B(net534),
    .Y(_04815_));
 sg13g2_a21oi_1 _22502_ (.A1(_10594_),
    .A2(net537),
    .Y(_04816_),
    .B1(_04815_));
 sg13g2_nand2_1 _22503_ (.Y(_04817_),
    .A(\cpu.ex.r_stmp[3] ),
    .B(net596));
 sg13g2_o21ai_1 _22504_ (.B1(_04817_),
    .Y(_01011_),
    .A1(_04796_),
    .A2(_04816_));
 sg13g2_nor2_1 _22505_ (.A(net666),
    .B(_04786_),
    .Y(_04818_));
 sg13g2_a21oi_1 _22506_ (.A1(_10768_),
    .A2(net537),
    .Y(_04819_),
    .B1(_04818_));
 sg13g2_nand2_1 _22507_ (.Y(_04820_),
    .A(\cpu.ex.r_stmp[4] ),
    .B(net596));
 sg13g2_o21ai_1 _22508_ (.B1(_04820_),
    .Y(_01012_),
    .A1(net535),
    .A2(_04819_));
 sg13g2_nor2_1 _22509_ (.A(net873),
    .B(_04786_),
    .Y(_04821_));
 sg13g2_a21oi_1 _22510_ (.A1(_10753_),
    .A2(net537),
    .Y(_04822_),
    .B1(_04821_));
 sg13g2_nand2_1 _22511_ (.Y(_04823_),
    .A(\cpu.ex.r_stmp[5] ),
    .B(net596));
 sg13g2_o21ai_1 _22512_ (.B1(_04823_),
    .Y(_01013_),
    .A1(net535),
    .A2(_04822_));
 sg13g2_mux2_1 _22513_ (.A0(net1000),
    .A1(_10685_),
    .S(net534),
    .X(_04824_));
 sg13g2_mux2_1 _22514_ (.A0(_04824_),
    .A1(\cpu.ex.r_stmp[6] ),
    .S(net536),
    .X(_01014_));
 sg13g2_nor2_1 _22515_ (.A(net871),
    .B(_04786_),
    .Y(_04825_));
 sg13g2_a21oi_1 _22516_ (.A1(_10722_),
    .A2(net537),
    .Y(_04826_),
    .B1(_04825_));
 sg13g2_nand2_1 _22517_ (.Y(_04827_),
    .A(\cpu.ex.r_stmp[7] ),
    .B(net596));
 sg13g2_o21ai_1 _22518_ (.B1(_04827_),
    .Y(_01015_),
    .A1(net535),
    .A2(_04826_));
 sg13g2_nor2_1 _22519_ (.A(_11300_),
    .B(_04786_),
    .Y(_04828_));
 sg13g2_a21oi_1 _22520_ (.A1(_10505_),
    .A2(_04787_),
    .Y(_04829_),
    .B1(_04828_));
 sg13g2_nand2_1 _22521_ (.Y(_04830_),
    .A(\cpu.ex.r_stmp[8] ),
    .B(net596));
 sg13g2_o21ai_1 _22522_ (.B1(_04830_),
    .Y(_01016_),
    .A1(_04796_),
    .A2(_04829_));
 sg13g2_nor2_1 _22523_ (.A(_02968_),
    .B(_04786_),
    .Y(_04831_));
 sg13g2_a21oi_1 _22524_ (.A1(_10530_),
    .A2(_04797_),
    .Y(_04832_),
    .B1(_04831_));
 sg13g2_nand2_1 _22525_ (.Y(_04833_),
    .A(\cpu.ex.r_stmp[9] ),
    .B(_04793_));
 sg13g2_o21ai_1 _22526_ (.B1(_04833_),
    .Y(_01017_),
    .A1(_04794_),
    .A2(_04832_));
 sg13g2_buf_1 _22527_ (.A(net1026),
    .X(_04834_));
 sg13g2_a22oi_1 _22528_ (.Y(_04835_),
    .B1(_09460_),
    .B2(\cpu.dcache.r_data[5][16] ),
    .A2(net609),
    .A1(\cpu.dcache.r_data[3][16] ));
 sg13g2_a22oi_1 _22529_ (.Y(_04836_),
    .B1(net562),
    .B2(\cpu.dcache.r_data[1][16] ),
    .A2(net610),
    .A1(\cpu.dcache.r_data[2][16] ));
 sg13g2_buf_1 _22530_ (.A(_09453_),
    .X(_04837_));
 sg13g2_mux2_1 _22531_ (.A0(\cpu.dcache.r_data[4][16] ),
    .A1(\cpu.dcache.r_data[6][16] ),
    .S(net632),
    .X(_04838_));
 sg13g2_a22oi_1 _22532_ (.Y(_04839_),
    .B1(_04838_),
    .B2(net600),
    .A2(net664),
    .A1(\cpu.dcache.r_data[7][16] ));
 sg13g2_nand2b_1 _22533_ (.Y(_04840_),
    .B(net673),
    .A_N(_04839_));
 sg13g2_nand3_1 _22534_ (.B(_04836_),
    .C(_04840_),
    .A(_04835_),
    .Y(_04841_));
 sg13g2_buf_1 _22535_ (.A(net628),
    .X(_04842_));
 sg13g2_mux2_1 _22536_ (.A0(\cpu.dcache.r_data[0][16] ),
    .A1(_04841_),
    .S(net533),
    .X(_04843_));
 sg13g2_nand2_1 _22537_ (.Y(_04844_),
    .A(net612),
    .B(_04843_));
 sg13g2_a22oi_1 _22538_ (.Y(_04845_),
    .B1(net562),
    .B2(\cpu.dcache.r_data[1][0] ),
    .A2(net610),
    .A1(\cpu.dcache.r_data[2][0] ));
 sg13g2_a22oi_1 _22539_ (.Y(_04846_),
    .B1(net609),
    .B2(\cpu.dcache.r_data[3][0] ),
    .A2(_09423_),
    .A1(\cpu.dcache.r_data[7][0] ));
 sg13g2_mux2_1 _22540_ (.A0(\cpu.dcache.r_data[4][0] ),
    .A1(\cpu.dcache.r_data[6][0] ),
    .S(net632),
    .X(_04847_));
 sg13g2_a22oi_1 _22541_ (.Y(_04848_),
    .B1(_04847_),
    .B2(net600),
    .A2(net918),
    .A1(\cpu.dcache.r_data[5][0] ));
 sg13g2_nand2b_1 _22542_ (.Y(_04849_),
    .B(net673),
    .A_N(_04848_));
 sg13g2_nand4_1 _22543_ (.B(_04845_),
    .C(_04846_),
    .A(net533),
    .Y(_04850_),
    .D(_04849_));
 sg13g2_o21ai_1 _22544_ (.B1(_04850_),
    .Y(_04851_),
    .A1(\cpu.dcache.r_data[0][0] ),
    .A2(net533));
 sg13g2_buf_1 _22545_ (.A(_12040_),
    .X(_04852_));
 sg13g2_mux2_1 _22546_ (.A0(_04844_),
    .A1(_04851_),
    .S(net983),
    .X(_04853_));
 sg13g2_nand2b_1 _22547_ (.Y(_04854_),
    .B(_08420_),
    .A_N(_08340_));
 sg13g2_or2_1 _22548_ (.X(_04855_),
    .B(_04854_),
    .A(_08457_));
 sg13g2_buf_1 _22549_ (.A(_04855_),
    .X(_04856_));
 sg13g2_buf_1 _22550_ (.A(_04856_),
    .X(_04857_));
 sg13g2_buf_1 _22551_ (.A(_04857_),
    .X(_04858_));
 sg13g2_buf_1 _22552_ (.A(net693),
    .X(_04859_));
 sg13g2_a22oi_1 _22553_ (.Y(_04860_),
    .B1(net609),
    .B2(\cpu.dcache.r_data[3][8] ),
    .A2(_09705_),
    .A1(\cpu.dcache.r_data[6][8] ));
 sg13g2_a22oi_1 _22554_ (.Y(_04861_),
    .B1(net562),
    .B2(\cpu.dcache.r_data[1][8] ),
    .A2(net610),
    .A1(\cpu.dcache.r_data[2][8] ));
 sg13g2_mux2_1 _22555_ (.A0(\cpu.dcache.r_data[5][8] ),
    .A1(\cpu.dcache.r_data[7][8] ),
    .S(net632),
    .X(_04862_));
 sg13g2_a22oi_1 _22556_ (.Y(_04863_),
    .B1(_04862_),
    .B2(net633),
    .A2(net921),
    .A1(\cpu.dcache.r_data[4][8] ));
 sg13g2_nand2b_1 _22557_ (.Y(_04864_),
    .B(_09456_),
    .A_N(_04863_));
 sg13g2_and4_1 _22558_ (.A(net533),
    .B(_04860_),
    .C(_04861_),
    .D(_04864_),
    .X(_04865_));
 sg13g2_a21oi_1 _22559_ (.A1(_00296_),
    .A2(net594),
    .Y(_04866_),
    .B1(_04865_));
 sg13g2_and2_1 _22560_ (.A(net685),
    .B(_04866_),
    .X(_04867_));
 sg13g2_a22oi_1 _22561_ (.Y(_04868_),
    .B1(_12469_),
    .B2(\cpu.dcache.r_data[3][24] ),
    .A2(net625),
    .A1(\cpu.dcache.r_data[6][24] ));
 sg13g2_a22oi_1 _22562_ (.Y(_04869_),
    .B1(net621),
    .B2(\cpu.dcache.r_data[4][24] ),
    .A2(net610),
    .A1(\cpu.dcache.r_data[2][24] ));
 sg13g2_mux2_1 _22563_ (.A0(\cpu.dcache.r_data[5][24] ),
    .A1(\cpu.dcache.r_data[7][24] ),
    .S(net632),
    .X(_04870_));
 sg13g2_a22oi_1 _22564_ (.Y(_04871_),
    .B1(_04870_),
    .B2(_09560_),
    .A2(_12198_),
    .A1(\cpu.dcache.r_data[1][24] ));
 sg13g2_and4_1 _22565_ (.A(_04842_),
    .B(_04868_),
    .C(_04869_),
    .D(_04871_),
    .X(_04872_));
 sg13g2_a21oi_1 _22566_ (.A1(_00295_),
    .A2(net594),
    .Y(_04873_),
    .B1(_04872_));
 sg13g2_nor2b_1 _22567_ (.A(net983),
    .B_N(_04873_),
    .Y(_04874_));
 sg13g2_nor3_1 _22568_ (.A(_04858_),
    .B(_04867_),
    .C(_04874_),
    .Y(_04875_));
 sg13g2_a21oi_1 _22569_ (.A1(_04853_),
    .A2(net595),
    .Y(_04876_),
    .B1(_04875_));
 sg13g2_buf_1 _22570_ (.A(net623),
    .X(_04877_));
 sg13g2_o21ai_1 _22571_ (.B1(_04844_),
    .Y(_04878_),
    .A1(net532),
    .A2(_04851_));
 sg13g2_nor3_2 _22572_ (.A(_08453_),
    .B(net1143),
    .C(_04854_),
    .Y(_04879_));
 sg13g2_buf_1 _22573_ (.A(_04879_),
    .X(_04880_));
 sg13g2_buf_1 _22574_ (.A(net742),
    .X(_04881_));
 sg13g2_mux2_1 _22575_ (.A0(_04876_),
    .A1(_04878_),
    .S(net662),
    .X(_04882_));
 sg13g2_nand2b_1 _22576_ (.Y(_04883_),
    .B(_09224_),
    .A_N(net1000));
 sg13g2_buf_2 _22577_ (.A(_04883_),
    .X(_04884_));
 sg13g2_nor2_1 _22578_ (.A(_09948_),
    .B(net1073),
    .Y(_04885_));
 sg13g2_nand2_1 _22579_ (.Y(_04886_),
    .A(_10039_),
    .B(net707));
 sg13g2_a221oi_1 _22580_ (.B2(net926),
    .C1(_09948_),
    .B1(_04886_),
    .A1(_09604_),
    .Y(_04887_),
    .A2(_04837_));
 sg13g2_nor2_1 _22581_ (.A(net694),
    .B(net1132),
    .Y(_04888_));
 sg13g2_o21ai_1 _22582_ (.B1(net1129),
    .Y(_04889_),
    .A1(net921),
    .A2(_04888_));
 sg13g2_nand2b_1 _22583_ (.Y(_04890_),
    .B(_04889_),
    .A_N(_04887_));
 sg13g2_o21ai_1 _22584_ (.B1(net1132),
    .Y(_04891_),
    .A1(_09228_),
    .A2(net791));
 sg13g2_nor2_1 _22585_ (.A(_09296_),
    .B(_04891_),
    .Y(_04892_));
 sg13g2_a221oi_1 _22586_ (.B2(net783),
    .C1(_04892_),
    .B1(_04890_),
    .A1(net785),
    .Y(_04893_),
    .A2(_04885_));
 sg13g2_buf_2 _22587_ (.A(_04893_),
    .X(_04894_));
 sg13g2_nor2_1 _22588_ (.A(_09227_),
    .B(net694),
    .Y(_04895_));
 sg13g2_and2_1 _22589_ (.A(_09581_),
    .B(_04895_),
    .X(_04896_));
 sg13g2_buf_2 _22590_ (.A(_04896_),
    .X(_04897_));
 sg13g2_and2_1 _22591_ (.A(net1043),
    .B(_04897_),
    .X(_04898_));
 sg13g2_buf_2 _22592_ (.A(_04898_),
    .X(_04899_));
 sg13g2_a21o_1 _22593_ (.A2(_04894_),
    .A1(_09179_),
    .B1(_04899_),
    .X(_04900_));
 sg13g2_buf_2 _22594_ (.A(\cpu.gpio.r_src_o[4][0] ),
    .X(_04901_));
 sg13g2_inv_2 _22595_ (.Y(_04902_),
    .A(net1132));
 sg13g2_nand2_1 _22596_ (.Y(_04903_),
    .A(_04902_),
    .B(_04897_));
 sg13g2_buf_1 _22597_ (.A(_04903_),
    .X(_04904_));
 sg13g2_inv_1 _22598_ (.Y(_04905_),
    .A(_04904_));
 sg13g2_nor4_1 _22599_ (.A(net912),
    .B(net694),
    .C(net791),
    .D(_09295_),
    .Y(_04906_));
 sg13g2_buf_1 _22600_ (.A(_04906_),
    .X(_04907_));
 sg13g2_and2_1 _22601_ (.A(net1129),
    .B(net487),
    .X(_04908_));
 sg13g2_buf_1 _22602_ (.A(_04908_),
    .X(_04909_));
 sg13g2_buf_2 _22603_ (.A(\cpu.gpio.r_src_o[6][0] ),
    .X(_04910_));
 sg13g2_a22oi_1 _22604_ (.Y(_04911_),
    .B1(net408),
    .B2(_04910_),
    .A2(_04905_),
    .A1(_04901_));
 sg13g2_nor2_1 _22605_ (.A(net791),
    .B(_09240_),
    .Y(_04912_));
 sg13g2_and2_1 _22606_ (.A(_04912_),
    .B(_04888_),
    .X(_04913_));
 sg13g2_buf_1 _22607_ (.A(_04913_),
    .X(_04914_));
 sg13g2_buf_2 _22608_ (.A(\cpu.gpio.r_src_io[4][0] ),
    .X(_04915_));
 sg13g2_buf_2 _22609_ (.A(\cpu.gpio.r_src_io[6][0] ),
    .X(_04916_));
 sg13g2_mux2_1 _22610_ (.A0(_04915_),
    .A1(_04916_),
    .S(net686),
    .X(_04917_));
 sg13g2_and2_1 _22611_ (.A(_09235_),
    .B(_04912_),
    .X(_04918_));
 sg13g2_buf_2 _22612_ (.A(_04918_),
    .X(_04919_));
 sg13g2_and2_1 _22613_ (.A(net1043),
    .B(_04919_),
    .X(_04920_));
 sg13g2_buf_1 _22614_ (.A(_04920_),
    .X(_04921_));
 sg13g2_a22oi_1 _22615_ (.Y(_04922_),
    .B1(net348),
    .B2(_09179_),
    .A2(_04917_),
    .A1(_04914_));
 sg13g2_buf_2 _22616_ (.A(\cpu.gpio.r_spi_miso_src[0][0] ),
    .X(_04923_));
 sg13g2_nor3_2 _22617_ (.A(net912),
    .B(_04902_),
    .C(_12709_),
    .Y(_04924_));
 sg13g2_nor3_1 _22618_ (.A(net1129),
    .B(_09227_),
    .C(_02698_),
    .Y(_04925_));
 sg13g2_buf_1 _22619_ (.A(_04925_),
    .X(_04926_));
 sg13g2_buf_2 _22620_ (.A(\cpu.gpio.r_uart_rx_src[0] ),
    .X(_04927_));
 sg13g2_a22oi_1 _22621_ (.Y(_04928_),
    .B1(net450),
    .B2(_04927_),
    .A2(_04924_),
    .A1(_04923_));
 sg13g2_nand3_1 _22622_ (.B(_04922_),
    .C(_04928_),
    .A(_04911_),
    .Y(_04929_));
 sg13g2_a21oi_1 _22623_ (.A1(_09180_),
    .A2(_04900_),
    .Y(_04930_),
    .B1(_04929_));
 sg13g2_and2_1 _22624_ (.A(net1000),
    .B(_09949_),
    .X(_04931_));
 sg13g2_buf_1 _22625_ (.A(_04931_),
    .X(_04932_));
 sg13g2_nor2_1 _22626_ (.A(net912),
    .B(_12709_),
    .Y(_04933_));
 sg13g2_buf_2 _22627_ (.A(_04933_),
    .X(_04934_));
 sg13g2_buf_1 _22628_ (.A(_04934_),
    .X(_04935_));
 sg13g2_a22oi_1 _22629_ (.Y(_04936_),
    .B1(_04935_),
    .B2(\cpu.intr.r_clock_cmp[16] ),
    .A2(net514),
    .A1(_10102_));
 sg13g2_nor2_1 _22630_ (.A(net1073),
    .B(net575),
    .Y(_04937_));
 sg13g2_buf_1 _22631_ (.A(_04937_),
    .X(_04938_));
 sg13g2_nor2_1 _22632_ (.A(net912),
    .B(net926),
    .Y(_04939_));
 sg13g2_nor2_2 _22633_ (.A(net1073),
    .B(net632),
    .Y(_04940_));
 sg13g2_a22oi_1 _22634_ (.Y(_04941_),
    .B1(_04940_),
    .B2(\cpu.intr.r_clock_cmp[0] ),
    .A2(_04939_),
    .A1(\cpu.intr.r_timer_reload[16] ));
 sg13g2_inv_1 _22635_ (.Y(_04942_),
    .A(_04941_));
 sg13g2_nor2_1 _22636_ (.A(net781),
    .B(_00269_),
    .Y(_04943_));
 sg13g2_a21oi_1 _22637_ (.A1(net686),
    .A2(_09959_),
    .Y(_04944_),
    .B1(_04943_));
 sg13g2_buf_2 _22638_ (.A(\cpu.intr.r_clock_count[16] ),
    .X(_04945_));
 sg13g2_buf_1 _22639_ (.A(_04897_),
    .X(_04946_));
 sg13g2_a22oi_1 _22640_ (.Y(_04947_),
    .B1(net448),
    .B2(_09167_),
    .A2(net417),
    .A1(_04945_));
 sg13g2_o21ai_1 _22641_ (.B1(_04947_),
    .Y(_04948_),
    .A1(_02698_),
    .A2(_04944_));
 sg13g2_a221oi_1 _22642_ (.B2(net689),
    .C1(_04948_),
    .B1(_04942_),
    .A1(\cpu.intr.r_timer_reload[0] ),
    .Y(_04949_),
    .A2(_04938_));
 sg13g2_nor2_1 _22643_ (.A(_10112_),
    .B(_04895_),
    .Y(_04950_));
 sg13g2_nor2_1 _22644_ (.A(net632),
    .B(_04950_),
    .Y(_04951_));
 sg13g2_nor2_1 _22645_ (.A(net791),
    .B(_04951_),
    .Y(_04952_));
 sg13g2_buf_1 _22646_ (.A(_04952_),
    .X(_04953_));
 sg13g2_and2_1 _22647_ (.A(_09581_),
    .B(_10112_),
    .X(_04954_));
 sg13g2_buf_1 _22648_ (.A(_04954_),
    .X(_04955_));
 sg13g2_a21o_1 _22649_ (.A2(net347),
    .A1(_09167_),
    .B1(net447),
    .X(_04956_));
 sg13g2_o21ai_1 _22650_ (.B1(_04956_),
    .Y(_04957_),
    .A1(_09165_),
    .A2(_09166_));
 sg13g2_nand3_1 _22651_ (.B(_04949_),
    .C(_04957_),
    .A(_04936_),
    .Y(_04958_));
 sg13g2_nor2_1 _22652_ (.A(net1073),
    .B(_02698_),
    .Y(_04959_));
 sg13g2_buf_1 _22653_ (.A(_04959_),
    .X(_04960_));
 sg13g2_nand2_1 _22654_ (.Y(_04961_),
    .A(_10112_),
    .B(_04912_));
 sg13g2_buf_1 _22655_ (.A(_04919_),
    .X(_04962_));
 sg13g2_nand2b_1 _22656_ (.Y(_04963_),
    .B(net406),
    .A_N(_00209_));
 sg13g2_o21ai_1 _22657_ (.B1(_04963_),
    .Y(_04964_),
    .A1(_00298_),
    .A2(_04961_));
 sg13g2_a21oi_1 _22658_ (.A1(\cpu.spi.r_mode[1][0] ),
    .A2(_04960_),
    .Y(_04965_),
    .B1(_04964_));
 sg13g2_o21ai_1 _22659_ (.B1(net706),
    .Y(_04966_),
    .A1(net783),
    .A2(net1132));
 sg13g2_inv_1 _22660_ (.Y(_04967_),
    .A(_09226_));
 sg13g2_nor2_1 _22661_ (.A(net707),
    .B(net791),
    .Y(_04968_));
 sg13g2_a22oi_1 _22662_ (.Y(_04969_),
    .B1(net1132),
    .B2(_04968_),
    .A2(_04967_),
    .A1(_09240_));
 sg13g2_nor3_1 _22663_ (.A(_09227_),
    .B(net915),
    .C(_04837_),
    .Y(_04970_));
 sg13g2_a21oi_1 _22664_ (.A1(_09227_),
    .A2(_04969_),
    .Y(_04971_),
    .B1(_04970_));
 sg13g2_a21oi_1 _22665_ (.A1(_03834_),
    .A2(_04966_),
    .Y(_04972_),
    .B1(_04971_));
 sg13g2_nor2_1 _22666_ (.A(net1129),
    .B(_04961_),
    .Y(_04973_));
 sg13g2_nor3_1 _22667_ (.A(net450),
    .B(_04972_),
    .C(_04973_),
    .Y(_04974_));
 sg13g2_buf_2 _22668_ (.A(_04974_),
    .X(_04975_));
 sg13g2_a22oi_1 _22669_ (.Y(_04976_),
    .B1(\cpu.spi.r_timeout[0] ),
    .B2(net463),
    .A2(_09226_),
    .A1(_09170_));
 sg13g2_inv_1 _22670_ (.Y(_04977_),
    .A(_04976_));
 sg13g2_a22oi_1 _22671_ (.Y(_04978_),
    .B1(_04977_),
    .B2(net686),
    .A2(_04940_),
    .A1(\cpu.spi.r_ready ));
 sg13g2_inv_1 _22672_ (.Y(_04979_),
    .A(_04978_));
 sg13g2_buf_1 _22673_ (.A(net1132),
    .X(_04980_));
 sg13g2_nand3_1 _22674_ (.B(net982),
    .C(net625),
    .A(net1073),
    .Y(_04981_));
 sg13g2_buf_2 _22675_ (.A(_04981_),
    .X(_04982_));
 sg13g2_buf_1 _22676_ (.A(\cpu.spi.r_clk_count[2][0] ),
    .X(_04983_));
 sg13g2_nor2_1 _22677_ (.A(net1132),
    .B(_04961_),
    .Y(_04984_));
 sg13g2_buf_2 _22678_ (.A(_04984_),
    .X(_04985_));
 sg13g2_and2_1 _22679_ (.A(net1030),
    .B(_12003_),
    .X(_04986_));
 sg13g2_a22oi_1 _22680_ (.Y(_04987_),
    .B1(_04986_),
    .B2(_04919_),
    .A2(_04985_),
    .A1(_04983_));
 sg13g2_o21ai_1 _22681_ (.B1(_04987_),
    .Y(_04988_),
    .A1(_00297_),
    .A2(_04982_));
 sg13g2_a221oi_1 _22682_ (.B2(net558),
    .C1(_04988_),
    .B1(_04979_),
    .A1(_09267_),
    .Y(_04989_),
    .A2(_04975_));
 sg13g2_o21ai_1 _22683_ (.B1(_04989_),
    .Y(_04990_),
    .A1(net888),
    .A2(_04965_));
 sg13g2_and2_1 _22684_ (.A(_09220_),
    .B(_09224_),
    .X(_04991_));
 sg13g2_buf_1 _22685_ (.A(_04991_),
    .X(_04992_));
 sg13g2_nand2b_1 _22686_ (.Y(_04993_),
    .B(_09951_),
    .A_N(_09224_));
 sg13g2_buf_1 _22687_ (.A(_04993_),
    .X(_04994_));
 sg13g2_o21ai_1 _22688_ (.B1(net783),
    .Y(_04995_),
    .A1(net785),
    .A2(net918));
 sg13g2_buf_2 _22689_ (.A(_04995_),
    .X(_04996_));
 sg13g2_and2_1 _22690_ (.A(_10112_),
    .B(_04912_),
    .X(_04997_));
 sg13g2_buf_1 _22691_ (.A(_04997_),
    .X(_04998_));
 sg13g2_a22oi_1 _22692_ (.Y(_04999_),
    .B1(net445),
    .B2(\cpu.uart.r_div_value[8] ),
    .A2(net406),
    .A1(\cpu.uart.r_div_value[0] ));
 sg13g2_a22oi_1 _22693_ (.Y(_05000_),
    .B1(net487),
    .B2(\cpu.uart.r_x_invert ),
    .A2(net448),
    .A1(_09165_));
 sg13g2_nand2_1 _22694_ (.Y(_05001_),
    .A(_04999_),
    .B(_05000_));
 sg13g2_a21oi_1 _22695_ (.A1(\cpu.uart.r_in[0] ),
    .A2(_04996_),
    .Y(_05002_),
    .B1(_05001_));
 sg13g2_o21ai_1 _22696_ (.B1(net1026),
    .Y(_05003_),
    .A1(net593),
    .A2(_05002_));
 sg13g2_a221oi_1 _22697_ (.B2(_04992_),
    .C1(_05003_),
    .B1(_04990_),
    .A1(_04932_),
    .Y(_05004_),
    .A2(_04958_));
 sg13g2_o21ai_1 _22698_ (.B1(_05004_),
    .Y(_05005_),
    .A1(_04884_),
    .A2(_04930_));
 sg13g2_o21ai_1 _22699_ (.B1(_05005_),
    .Y(_05006_),
    .A1(net855),
    .A2(_04882_));
 sg13g2_buf_1 _22700_ (.A(_03555_),
    .X(_05007_));
 sg13g2_nand2_1 _22701_ (.Y(_05008_),
    .A(_03489_),
    .B(net75));
 sg13g2_o21ai_1 _22702_ (.B1(_05008_),
    .Y(_05009_),
    .A1(net36),
    .A2(_05006_));
 sg13g2_nand2_2 _22703_ (.Y(_05010_),
    .A(_04100_),
    .B(_11481_));
 sg13g2_nand3_1 _22704_ (.B(net87),
    .C(net206),
    .A(net461),
    .Y(_05011_));
 sg13g2_nor3_1 _22705_ (.A(_11425_),
    .B(_11444_),
    .C(_05011_),
    .Y(_05012_));
 sg13g2_nand3_1 _22706_ (.B(net187),
    .C(_04555_),
    .A(net226),
    .Y(_05013_));
 sg13g2_and2_1 _22707_ (.A(net134),
    .B(_04161_),
    .X(_05014_));
 sg13g2_a221oi_1 _22708_ (.B2(_04250_),
    .C1(_05014_),
    .B1(_04252_),
    .A1(net186),
    .Y(_05015_),
    .A2(net138));
 sg13g2_a22oi_1 _22709_ (.Y(_05016_),
    .B1(net187),
    .B2(net140),
    .A2(_04155_),
    .A1(net192));
 sg13g2_nand2b_1 _22710_ (.Y(_05017_),
    .B(_04148_),
    .A_N(_05016_));
 sg13g2_a22oi_1 _22711_ (.Y(_05018_),
    .B1(_04165_),
    .B2(_03616_),
    .A2(_04185_),
    .A1(_03610_));
 sg13g2_a21oi_1 _22712_ (.A1(net122),
    .A2(_04193_),
    .Y(_05019_),
    .B1(_04378_));
 sg13g2_a22oi_1 _22713_ (.Y(_05020_),
    .B1(net157),
    .B2(_03577_),
    .A2(net156),
    .A1(_03622_));
 sg13g2_and4_1 _22714_ (.A(_04549_),
    .B(_05018_),
    .C(_05019_),
    .D(_05020_),
    .X(_05021_));
 sg13g2_and4_1 _22715_ (.A(_05013_),
    .B(_05015_),
    .C(_05017_),
    .D(_05021_),
    .X(_05022_));
 sg13g2_nand2_1 _22716_ (.Y(_05023_),
    .A(_10677_),
    .B(net159));
 sg13g2_o21ai_1 _22717_ (.B1(_05023_),
    .Y(_05024_),
    .A1(net856),
    .A2(_05022_));
 sg13g2_o21ai_1 _22718_ (.B1(_05024_),
    .Y(_05025_),
    .A1(net203),
    .A2(_04203_));
 sg13g2_nor3_1 _22719_ (.A(_08335_),
    .B(net1140),
    .C(_04122_),
    .Y(_05026_));
 sg13g2_a22oi_1 _22720_ (.Y(_05027_),
    .B1(_05026_),
    .B2(net218),
    .A2(_04119_),
    .A1(_09147_));
 sg13g2_or2_1 _22721_ (.X(_05028_),
    .B(_05027_),
    .A(net1063));
 sg13g2_nor2b_1 _22722_ (.A(net1131),
    .B_N(_05026_),
    .Y(_05029_));
 sg13g2_o21ai_1 _22723_ (.B1(net279),
    .Y(_05030_),
    .A1(net198),
    .A2(_05029_));
 sg13g2_a221oi_1 _22724_ (.B2(_05030_),
    .C1(net206),
    .B1(_05028_),
    .A1(net991),
    .Y(_05031_),
    .A2(_10523_));
 sg13g2_a22oi_1 _22725_ (.Y(_05032_),
    .B1(_05025_),
    .B2(_05031_),
    .A2(_04106_),
    .A1(_11464_));
 sg13g2_nand3_1 _22726_ (.B(_11454_),
    .C(net206),
    .A(net461),
    .Y(_05033_));
 sg13g2_nand2b_1 _22727_ (.Y(_05034_),
    .B(_05033_),
    .A_N(_05032_));
 sg13g2_nor2_1 _22728_ (.A(_05012_),
    .B(_05034_),
    .Y(_05035_));
 sg13g2_nand2_1 _22729_ (.Y(_05036_),
    .A(net994),
    .B(_05010_));
 sg13g2_o21ai_1 _22730_ (.B1(_05036_),
    .Y(_05037_),
    .A1(_05010_),
    .A2(_05035_));
 sg13g2_buf_2 _22731_ (.A(_11487_),
    .X(_05038_));
 sg13g2_mux2_1 _22732_ (.A0(_05009_),
    .A1(_05037_),
    .S(_05038_),
    .X(_01018_));
 sg13g2_buf_1 _22733_ (.A(net141),
    .X(_05039_));
 sg13g2_a22oi_1 _22734_ (.Y(_05040_),
    .B1(net609),
    .B2(\cpu.dcache.r_data[3][7] ),
    .A2(net625),
    .A1(\cpu.dcache.r_data[6][7] ));
 sg13g2_a22oi_1 _22735_ (.Y(_05041_),
    .B1(net627),
    .B2(\cpu.dcache.r_data[1][7] ),
    .A2(net610),
    .A1(\cpu.dcache.r_data[2][7] ));
 sg13g2_mux2_1 _22736_ (.A0(\cpu.dcache.r_data[5][7] ),
    .A1(\cpu.dcache.r_data[7][7] ),
    .S(net706),
    .X(_05042_));
 sg13g2_a22oi_1 _22737_ (.Y(_05043_),
    .B1(_05042_),
    .B2(net633),
    .A2(net921),
    .A1(\cpu.dcache.r_data[4][7] ));
 sg13g2_nand2b_1 _22738_ (.Y(_05044_),
    .B(net791),
    .A_N(_05043_));
 sg13g2_and4_1 _22739_ (.A(net533),
    .B(_05040_),
    .C(_05041_),
    .D(_05044_),
    .X(_05045_));
 sg13g2_a21oi_1 _22740_ (.A1(_00144_),
    .A2(net594),
    .Y(_05046_),
    .B1(_05045_));
 sg13g2_mux2_1 _22741_ (.A0(\cpu.dcache.r_data[5][23] ),
    .A1(\cpu.dcache.r_data[7][23] ),
    .S(net706),
    .X(_05047_));
 sg13g2_a22oi_1 _22742_ (.Y(_05048_),
    .B1(_05047_),
    .B2(net633),
    .A2(net785),
    .A1(\cpu.dcache.r_data[6][23] ));
 sg13g2_nand2b_1 _22743_ (.Y(_05049_),
    .B(net791),
    .A_N(_05048_));
 sg13g2_mux2_1 _22744_ (.A0(\cpu.dcache.r_data[2][23] ),
    .A1(\cpu.dcache.r_data[3][23] ),
    .S(net707),
    .X(_05050_));
 sg13g2_a22oi_1 _22745_ (.Y(_05051_),
    .B1(_05050_),
    .B2(net790),
    .A2(_09552_),
    .A1(\cpu.dcache.r_data[4][23] ));
 sg13g2_nand2_1 _22746_ (.Y(_05052_),
    .A(\cpu.dcache.r_data[1][23] ),
    .B(net627));
 sg13g2_nand2b_1 _22747_ (.Y(_05053_),
    .B(net693),
    .A_N(_00145_));
 sg13g2_nand4_1 _22748_ (.B(_05051_),
    .C(_05052_),
    .A(_05049_),
    .Y(_05054_),
    .D(_05053_));
 sg13g2_and2_1 _22749_ (.A(_09942_),
    .B(_05054_),
    .X(_05055_));
 sg13g2_a21oi_1 _22750_ (.A1(_10040_),
    .A2(_05046_),
    .Y(_05056_),
    .B1(_05055_));
 sg13g2_inv_1 _22751_ (.Y(_05057_),
    .A(_00146_));
 sg13g2_a22oi_1 _22752_ (.Y(_05058_),
    .B1(_09425_),
    .B2(\cpu.dcache.r_data[3][31] ),
    .A2(net625),
    .A1(\cpu.dcache.r_data[6][31] ));
 sg13g2_a22oi_1 _22753_ (.Y(_05059_),
    .B1(net621),
    .B2(\cpu.dcache.r_data[4][31] ),
    .A2(_12340_),
    .A1(\cpu.dcache.r_data[2][31] ));
 sg13g2_mux2_1 _22754_ (.A0(\cpu.dcache.r_data[5][31] ),
    .A1(\cpu.dcache.r_data[7][31] ),
    .S(net706),
    .X(_05060_));
 sg13g2_a22oi_1 _22755_ (.Y(_05061_),
    .B1(_05060_),
    .B2(_09560_),
    .A2(net627),
    .A1(\cpu.dcache.r_data[1][31] ));
 sg13g2_nand4_1 _22756_ (.B(_05058_),
    .C(_05059_),
    .A(net628),
    .Y(_05062_),
    .D(_05061_));
 sg13g2_o21ai_1 _22757_ (.B1(_05062_),
    .Y(_05063_),
    .A1(_05057_),
    .A2(_04842_));
 sg13g2_nand3_1 _22758_ (.B(_04856_),
    .C(_05054_),
    .A(_09942_),
    .Y(_05064_));
 sg13g2_o21ai_1 _22759_ (.B1(_05064_),
    .Y(_05065_),
    .A1(net663),
    .A2(_05063_));
 sg13g2_nor2b_1 _22760_ (.A(_12040_),
    .B_N(_05065_),
    .Y(_05066_));
 sg13g2_nand2_1 _22761_ (.Y(_05067_),
    .A(\cpu.dcache.r_data[2][15] ),
    .B(net610));
 sg13g2_a22oi_1 _22762_ (.Y(_05068_),
    .B1(_09460_),
    .B2(\cpu.dcache.r_data[5][15] ),
    .A2(_09423_),
    .A1(\cpu.dcache.r_data[7][15] ));
 sg13g2_a22oi_1 _22763_ (.Y(_05069_),
    .B1(net621),
    .B2(\cpu.dcache.r_data[4][15] ),
    .A2(_09419_),
    .A1(\cpu.dcache.r_data[1][15] ));
 sg13g2_a22oi_1 _22764_ (.Y(_05070_),
    .B1(_09425_),
    .B2(\cpu.dcache.r_data[3][15] ),
    .A2(net625),
    .A1(\cpu.dcache.r_data[6][15] ));
 sg13g2_nand4_1 _22765_ (.B(_05068_),
    .C(_05069_),
    .A(_05067_),
    .Y(_05071_),
    .D(_05070_));
 sg13g2_nand2_1 _22766_ (.Y(_05072_),
    .A(_00147_),
    .B(net594));
 sg13g2_o21ai_1 _22767_ (.B1(_05072_),
    .Y(_05073_),
    .A1(net594),
    .A2(_05071_));
 sg13g2_nor3_1 _22768_ (.A(net914),
    .B(net663),
    .C(_05073_),
    .Y(_05074_));
 sg13g2_and3_1 _22769_ (.X(_05075_),
    .A(_12040_),
    .B(net663),
    .C(_05046_));
 sg13g2_nor4_1 _22770_ (.A(_04879_),
    .B(_05066_),
    .C(_05074_),
    .D(_05075_),
    .Y(_05076_));
 sg13g2_a21oi_1 _22771_ (.A1(_04879_),
    .A2(_05056_),
    .Y(_05077_),
    .B1(_05076_));
 sg13g2_nand3_1 _22772_ (.B(_09186_),
    .C(_04894_),
    .A(_09185_),
    .Y(_05078_));
 sg13g2_nor2_1 _22773_ (.A(net1073),
    .B(_12709_),
    .Y(_05079_));
 sg13g2_buf_1 _22774_ (.A(_05079_),
    .X(_05080_));
 sg13g2_nand2_1 _22775_ (.Y(_05081_),
    .A(net10),
    .B(_05080_));
 sg13g2_a22oi_1 _22776_ (.Y(_05082_),
    .B1(_10114_),
    .B2(\cpu.gpio.genblk2[7].srcs_io[0] ),
    .A2(_10093_),
    .A1(\cpu.gpio.genblk1[7].srcs_o[0] ));
 sg13g2_a21oi_1 _22777_ (.A1(_05081_),
    .A2(_05082_),
    .Y(_05083_),
    .B1(_04902_));
 sg13g2_nand2_2 _22778_ (.Y(_05084_),
    .A(_09581_),
    .B(_10112_));
 sg13g2_nor2_1 _22779_ (.A(_00153_),
    .B(_05084_),
    .Y(_05085_));
 sg13g2_nor2b_1 _22780_ (.A(net1129),
    .B_N(_09185_),
    .Y(_05086_));
 sg13g2_a22oi_1 _22781_ (.Y(_05087_),
    .B1(_05086_),
    .B2(_04919_),
    .A2(_05085_),
    .A1(net1129));
 sg13g2_inv_1 _22782_ (.Y(_05088_),
    .A(_00154_));
 sg13g2_nand2_1 _22783_ (.Y(_05089_),
    .A(_09191_),
    .B(net1132));
 sg13g2_nand2_1 _22784_ (.Y(_05090_),
    .A(net1043),
    .B(net445));
 sg13g2_buf_2 _22785_ (.A(_05090_),
    .X(_05091_));
 sg13g2_o21ai_1 _22786_ (.B1(_05091_),
    .Y(_05092_),
    .A1(_05084_),
    .A2(_05089_));
 sg13g2_a22oi_1 _22787_ (.Y(_05093_),
    .B1(_05092_),
    .B2(\cpu.gpio.r_enable_io[7] ),
    .A2(_04924_),
    .A1(_05088_));
 sg13g2_buf_1 _22788_ (.A(\cpu.gpio.r_src_io[5][3] ),
    .X(_05094_));
 sg13g2_nand2_1 _22789_ (.Y(_05095_),
    .A(net912),
    .B(_05094_));
 sg13g2_o21ai_1 _22790_ (.B1(_05095_),
    .Y(_05096_),
    .A1(net912),
    .A2(_00150_));
 sg13g2_o21ai_1 _22791_ (.B1(_05089_),
    .Y(_05097_),
    .A1(net1043),
    .A2(_00151_));
 sg13g2_a22oi_1 _22792_ (.Y(_05098_),
    .B1(_05097_),
    .B2(_04907_),
    .A2(_05096_),
    .A1(net486));
 sg13g2_inv_1 _22793_ (.Y(_05099_),
    .A(_00152_));
 sg13g2_a22oi_1 _22794_ (.Y(_05100_),
    .B1(_04899_),
    .B2(_09186_),
    .A2(_04905_),
    .A1(_05099_));
 sg13g2_nand4_1 _22795_ (.B(_05093_),
    .C(_05098_),
    .A(_05087_),
    .Y(_05101_),
    .D(_05100_));
 sg13g2_nor2_1 _22796_ (.A(_05083_),
    .B(_05101_),
    .Y(_05102_));
 sg13g2_a21oi_1 _22797_ (.A1(_05078_),
    .A2(_05102_),
    .Y(_05103_),
    .B1(_04884_));
 sg13g2_nor2_1 _22798_ (.A(_09951_),
    .B(net347),
    .Y(_05104_));
 sg13g2_a22oi_1 _22799_ (.Y(_05105_),
    .B1(_09460_),
    .B2(\cpu.intr.r_clock_cmp[23] ),
    .A2(net625),
    .A1(_09984_));
 sg13g2_nand2b_1 _22800_ (.Y(_05106_),
    .B(net914),
    .A_N(_05105_));
 sg13g2_a22oi_1 _22801_ (.Y(_05107_),
    .B1(_04940_),
    .B2(\cpu.intr.r_clock_cmp[7] ),
    .A2(_04939_),
    .A1(\cpu.intr.r_timer_reload[23] ));
 sg13g2_nor2b_1 _22802_ (.A(_05107_),
    .B_N(net689),
    .Y(_05108_));
 sg13g2_a221oi_1 _22803_ (.B2(\cpu.intr.r_timer_reload[7] ),
    .C1(_05108_),
    .B1(_04937_),
    .A1(_10141_),
    .Y(_05109_),
    .A2(net573));
 sg13g2_buf_1 _22804_ (.A(\cpu.intr.r_clock_count[23] ),
    .X(_05110_));
 sg13g2_a22oi_1 _22805_ (.Y(_05111_),
    .B1(_04959_),
    .B2(\cpu.intr.r_timer_count[7] ),
    .A2(_10114_),
    .A1(_05110_));
 sg13g2_nand3_1 _22806_ (.B(_05109_),
    .C(_05111_),
    .A(_05106_),
    .Y(_05112_));
 sg13g2_or2_1 _22807_ (.X(_05113_),
    .B(_04982_),
    .A(_00148_));
 sg13g2_buf_1 _22808_ (.A(\cpu.spi.r_clk_count[2][7] ),
    .X(_05114_));
 sg13g2_nor3_1 _22809_ (.A(net912),
    .B(_03834_),
    .C(net926),
    .Y(_05115_));
 sg13g2_buf_2 _22810_ (.A(_05115_),
    .X(_05116_));
 sg13g2_nor2_1 _22811_ (.A(_00149_),
    .B(_05091_),
    .Y(_05117_));
 sg13g2_a221oi_1 _22812_ (.B2(\cpu.spi.r_timeout[7] ),
    .C1(_05117_),
    .B1(_05116_),
    .A1(_05114_),
    .Y(_05118_),
    .A2(_04985_));
 sg13g2_nand2b_1 _22813_ (.Y(_05119_),
    .B(_04975_),
    .A_N(_00206_));
 sg13g2_nand3_1 _22814_ (.B(_05118_),
    .C(_05119_),
    .A(_05113_),
    .Y(_05120_));
 sg13g2_a22oi_1 _22815_ (.Y(_05121_),
    .B1(_04996_),
    .B2(\cpu.uart.r_in[7] ),
    .A2(_04919_),
    .A1(\cpu.uart.r_div_value[7] ));
 sg13g2_nor2_1 _22816_ (.A(net593),
    .B(_05121_),
    .Y(_05122_));
 sg13g2_a221oi_1 _22817_ (.B2(_04992_),
    .C1(_05122_),
    .B1(_05120_),
    .A1(_05104_),
    .Y(_05123_),
    .A2(_05112_));
 sg13g2_nand3b_1 _22818_ (.B(_05123_),
    .C(_08340_),
    .Y(_05124_),
    .A_N(_05103_));
 sg13g2_o21ai_1 _22819_ (.B1(_05124_),
    .Y(_05125_),
    .A1(net1026),
    .A2(_05077_));
 sg13g2_and2_1 _22820_ (.A(_08453_),
    .B(_05125_),
    .X(_05126_));
 sg13g2_buf_1 _22821_ (.A(_05126_),
    .X(_05127_));
 sg13g2_buf_1 _22822_ (.A(net594),
    .X(_05128_));
 sg13g2_buf_1 _22823_ (.A(_05128_),
    .X(_05129_));
 sg13g2_nand2_1 _22824_ (.Y(_05130_),
    .A(\cpu.dcache.r_data[2][26] ),
    .B(net502));
 sg13g2_a22oi_1 _22825_ (.Y(_05131_),
    .B1(_12702_),
    .B2(\cpu.dcache.r_data[5][26] ),
    .A2(net576),
    .A1(\cpu.dcache.r_data[7][26] ));
 sg13g2_buf_1 _22826_ (.A(net562),
    .X(_05132_));
 sg13g2_a22oi_1 _22827_ (.Y(_05133_),
    .B1(net621),
    .B2(\cpu.dcache.r_data[4][26] ),
    .A2(net484),
    .A1(\cpu.dcache.r_data[1][26] ));
 sg13g2_buf_1 _22828_ (.A(net609),
    .X(_05134_));
 sg13g2_a22oi_1 _22829_ (.Y(_05135_),
    .B1(net530),
    .B2(\cpu.dcache.r_data[3][26] ),
    .A2(net556),
    .A1(\cpu.dcache.r_data[6][26] ));
 sg13g2_nand4_1 _22830_ (.B(_05131_),
    .C(_05133_),
    .A(_05130_),
    .Y(_05136_),
    .D(_05135_));
 sg13g2_nor2_1 _22831_ (.A(net531),
    .B(_05136_),
    .Y(_05137_));
 sg13g2_a21oi_1 _22832_ (.A1(_00098_),
    .A2(net485),
    .Y(_05138_),
    .B1(_05137_));
 sg13g2_nand2_1 _22833_ (.Y(_05139_),
    .A(\cpu.dcache.r_data[2][10] ),
    .B(net502));
 sg13g2_a22oi_1 _22834_ (.Y(_05140_),
    .B1(_12703_),
    .B2(\cpu.dcache.r_data[5][10] ),
    .A2(_09946_),
    .A1(\cpu.dcache.r_data[7][10] ));
 sg13g2_a22oi_1 _22835_ (.Y(_05141_),
    .B1(net574),
    .B2(\cpu.dcache.r_data[4][10] ),
    .A2(net503),
    .A1(\cpu.dcache.r_data[1][10] ));
 sg13g2_a22oi_1 _22836_ (.Y(_05142_),
    .B1(net559),
    .B2(\cpu.dcache.r_data[3][10] ),
    .A2(_02692_),
    .A1(\cpu.dcache.r_data[6][10] ));
 sg13g2_nand4_1 _22837_ (.B(_05140_),
    .C(_05141_),
    .A(_05139_),
    .Y(_05143_),
    .D(_05142_));
 sg13g2_nand2_1 _22838_ (.Y(_05144_),
    .A(_00099_),
    .B(net485));
 sg13g2_o21ai_1 _22839_ (.B1(_05144_),
    .Y(_05145_),
    .A1(net485),
    .A2(_05143_));
 sg13g2_nor2_1 _22840_ (.A(net612),
    .B(_05145_),
    .Y(_05146_));
 sg13g2_a21o_1 _22841_ (.A2(_05138_),
    .A1(net532),
    .B1(_05146_),
    .X(_05147_));
 sg13g2_and2_1 _22842_ (.A(net1026),
    .B(_05104_),
    .X(_05148_));
 sg13g2_buf_2 _22843_ (.A(_05148_),
    .X(_05149_));
 sg13g2_a22oi_1 _22844_ (.Y(_05150_),
    .B1(net446),
    .B2(\cpu.intr.r_timer_count[10] ),
    .A2(net407),
    .A1(\cpu.intr.r_clock_cmp[26] ));
 sg13g2_a22oi_1 _22845_ (.Y(_05151_),
    .B1(net449),
    .B2(\cpu.intr.r_timer_reload[10] ),
    .A2(net514),
    .A1(_10158_));
 sg13g2_buf_2 _22846_ (.A(\cpu.intr.r_clock_count[26] ),
    .X(_05152_));
 sg13g2_buf_1 _22847_ (.A(_05080_),
    .X(_05153_));
 sg13g2_a22oi_1 _22848_ (.Y(_05154_),
    .B1(net405),
    .B2(\cpu.intr.r_clock_cmp[10] ),
    .A2(net362),
    .A1(_05152_));
 sg13g2_nand3_1 _22849_ (.B(_05151_),
    .C(_05154_),
    .A(_05150_),
    .Y(_05155_));
 sg13g2_buf_1 _22850_ (.A(net1144),
    .X(_05156_));
 sg13g2_a221oi_1 _22851_ (.B2(_05155_),
    .C1(net981),
    .B1(_05149_),
    .A1(net662),
    .Y(_05157_),
    .A2(_05147_));
 sg13g2_nor3_1 _22852_ (.A(net76),
    .B(_05127_),
    .C(_05157_),
    .Y(_05158_));
 sg13g2_a21oi_1 _22853_ (.A1(_10392_),
    .A2(net75),
    .Y(_05159_),
    .B1(_05158_));
 sg13g2_a21oi_1 _22854_ (.A1(_00242_),
    .A2(_11478_),
    .Y(_05160_),
    .B1(_09213_));
 sg13g2_buf_1 _22855_ (.A(_05160_),
    .X(_05161_));
 sg13g2_buf_1 _22856_ (.A(net661),
    .X(_05162_));
 sg13g2_nand2b_1 _22857_ (.Y(_05163_),
    .B(_05162_),
    .A_N(_04776_));
 sg13g2_o21ai_1 _22858_ (.B1(_05163_),
    .Y(_05164_),
    .A1(net592),
    .A2(_04772_));
 sg13g2_buf_1 _22859_ (.A(_04211_),
    .X(_05165_));
 sg13g2_nor2_1 _22860_ (.A(net153),
    .B(net141),
    .Y(_05166_));
 sg13g2_buf_1 _22861_ (.A(_04100_),
    .X(_05167_));
 sg13g2_buf_1 _22862_ (.A(_05167_),
    .X(_05168_));
 sg13g2_nor3_1 _22863_ (.A(net985),
    .B(net130),
    .C(net121),
    .Y(_05169_));
 sg13g2_a221oi_1 _22864_ (.B2(_05166_),
    .C1(_05169_),
    .B1(_05164_),
    .A1(net115),
    .Y(_01019_),
    .A2(_05159_));
 sg13g2_buf_1 _22865_ (.A(_11487_),
    .X(_05170_));
 sg13g2_a221oi_1 _22866_ (.B2(net239),
    .C1(_04275_),
    .B1(_04274_),
    .A1(net981),
    .Y(_05171_),
    .A2(_11479_));
 sg13g2_buf_1 _22867_ (.A(_11481_),
    .X(_05172_));
 sg13g2_o21ai_1 _22868_ (.B1(_05167_),
    .Y(_05173_),
    .A1(net529),
    .A2(_04283_));
 sg13g2_nand2_1 _22869_ (.Y(_05174_),
    .A(\cpu.ex.pc[11] ),
    .B(net153));
 sg13g2_o21ai_1 _22870_ (.B1(_05174_),
    .Y(_05175_),
    .A1(_05171_),
    .A2(_05173_));
 sg13g2_nand2_1 _22871_ (.Y(_05176_),
    .A(\cpu.dcache.r_data[2][27] ),
    .B(net502));
 sg13g2_a22oi_1 _22872_ (.Y(_05177_),
    .B1(net608),
    .B2(\cpu.dcache.r_data[5][27] ),
    .A2(net576),
    .A1(\cpu.dcache.r_data[7][27] ));
 sg13g2_a22oi_1 _22873_ (.Y(_05178_),
    .B1(net621),
    .B2(\cpu.dcache.r_data[4][27] ),
    .A2(net484),
    .A1(\cpu.dcache.r_data[1][27] ));
 sg13g2_a22oi_1 _22874_ (.Y(_05179_),
    .B1(net530),
    .B2(\cpu.dcache.r_data[3][27] ),
    .A2(net556),
    .A1(\cpu.dcache.r_data[6][27] ));
 sg13g2_nand4_1 _22875_ (.B(_05177_),
    .C(_05178_),
    .A(_05176_),
    .Y(_05180_),
    .D(_05179_));
 sg13g2_nor2_1 _22876_ (.A(net531),
    .B(_05180_),
    .Y(_05181_));
 sg13g2_a21oi_1 _22877_ (.A1(_00108_),
    .A2(net485),
    .Y(_05182_),
    .B1(_05181_));
 sg13g2_inv_1 _22878_ (.Y(_05183_),
    .A(_00109_));
 sg13g2_buf_1 _22879_ (.A(net533),
    .X(_05184_));
 sg13g2_a22oi_1 _22880_ (.Y(_05185_),
    .B1(net502),
    .B2(\cpu.dcache.r_data[2][11] ),
    .A2(net559),
    .A1(\cpu.dcache.r_data[3][11] ));
 sg13g2_a22oi_1 _22881_ (.Y(_05186_),
    .B1(net503),
    .B2(\cpu.dcache.r_data[1][11] ),
    .A2(net608),
    .A1(\cpu.dcache.r_data[5][11] ));
 sg13g2_mux2_1 _22882_ (.A0(\cpu.dcache.r_data[4][11] ),
    .A1(\cpu.dcache.r_data[6][11] ),
    .S(_09297_),
    .X(_05187_));
 sg13g2_a22oi_1 _22883_ (.Y(_05188_),
    .B1(_05187_),
    .B2(net540),
    .A2(net664),
    .A1(\cpu.dcache.r_data[7][11] ));
 sg13g2_nand2b_1 _22884_ (.Y(_05189_),
    .B(net613),
    .A_N(_05188_));
 sg13g2_nand4_1 _22885_ (.B(_05185_),
    .C(_05186_),
    .A(_05184_),
    .Y(_05190_),
    .D(_05189_));
 sg13g2_o21ai_1 _22886_ (.B1(_05190_),
    .Y(_05191_),
    .A1(_05183_),
    .A2(net483));
 sg13g2_nor2_1 _22887_ (.A(net612),
    .B(_05191_),
    .Y(_05192_));
 sg13g2_a21o_1 _22888_ (.A2(_05182_),
    .A1(net532),
    .B1(_05192_),
    .X(_05193_));
 sg13g2_a22oi_1 _22889_ (.Y(_05194_),
    .B1(net446),
    .B2(\cpu.intr.r_timer_count[11] ),
    .A2(net514),
    .A1(_10163_));
 sg13g2_a22oi_1 _22890_ (.Y(_05195_),
    .B1(net405),
    .B2(\cpu.intr.r_clock_cmp[11] ),
    .A2(net449),
    .A1(\cpu.intr.r_timer_reload[11] ));
 sg13g2_buf_1 _22891_ (.A(\cpu.intr.r_clock_count[27] ),
    .X(_05196_));
 sg13g2_a22oi_1 _22892_ (.Y(_05197_),
    .B1(net407),
    .B2(\cpu.intr.r_clock_cmp[27] ),
    .A2(net362),
    .A1(_05196_));
 sg13g2_nand3_1 _22893_ (.B(_05195_),
    .C(_05197_),
    .A(_05194_),
    .Y(_05198_));
 sg13g2_a221oi_1 _22894_ (.B2(_05149_),
    .C1(net1144),
    .B1(_05198_),
    .A1(net662),
    .Y(_05199_),
    .A2(_05193_));
 sg13g2_nor3_1 _22895_ (.A(_03555_),
    .B(_05127_),
    .C(_05199_),
    .Y(_05200_));
 sg13g2_a21oi_1 _22896_ (.A1(net1122),
    .A2(_05007_),
    .Y(_05201_),
    .B1(_05200_));
 sg13g2_nor2_1 _22897_ (.A(_11487_),
    .B(_05201_),
    .Y(_05202_));
 sg13g2_a21o_1 _22898_ (.A2(_05175_),
    .A1(_05170_),
    .B1(_05202_),
    .X(_01020_));
 sg13g2_nand3b_1 _22899_ (.B(net592),
    .C(net152),
    .Y(_05203_),
    .A_N(_04333_));
 sg13g2_o21ai_1 _22900_ (.B1(_05203_),
    .Y(_05204_),
    .A1(_08550_),
    .A2(net152));
 sg13g2_nor2_1 _22901_ (.A(net121),
    .B(_05010_),
    .Y(_05205_));
 sg13g2_a22oi_1 _22902_ (.Y(_05206_),
    .B1(net449),
    .B2(\cpu.intr.r_timer_reload[12] ),
    .A2(net514),
    .A1(_10169_));
 sg13g2_a22oi_1 _22903_ (.Y(_05207_),
    .B1(net405),
    .B2(\cpu.intr.r_clock_cmp[12] ),
    .A2(net407),
    .A1(\cpu.intr.r_clock_cmp[28] ));
 sg13g2_buf_2 _22904_ (.A(\cpu.intr.r_clock_count[28] ),
    .X(_05208_));
 sg13g2_a22oi_1 _22905_ (.Y(_05209_),
    .B1(net446),
    .B2(_09961_),
    .A2(net362),
    .A1(_05208_));
 sg13g2_nand3_1 _22906_ (.B(_05207_),
    .C(_05209_),
    .A(_05206_),
    .Y(_05210_));
 sg13g2_mux2_1 _22907_ (.A0(\cpu.dcache.r_data[4][12] ),
    .A1(\cpu.dcache.r_data[6][12] ),
    .S(net578),
    .X(_05211_));
 sg13g2_a22oi_1 _22908_ (.Y(_05212_),
    .B1(_05211_),
    .B2(net540),
    .A2(net664),
    .A1(\cpu.dcache.r_data[7][12] ));
 sg13g2_nor2_1 _22909_ (.A(net783),
    .B(_05212_),
    .Y(_05213_));
 sg13g2_mux2_1 _22910_ (.A0(\cpu.dcache.r_data[2][12] ),
    .A1(\cpu.dcache.r_data[3][12] ),
    .S(net633),
    .X(_05214_));
 sg13g2_a22oi_1 _22911_ (.Y(_05215_),
    .B1(_05214_),
    .B2(net790),
    .A2(net608),
    .A1(\cpu.dcache.r_data[5][12] ));
 sg13g2_o21ai_1 _22912_ (.B1(_05215_),
    .Y(_05216_),
    .A1(_12231_),
    .A2(_12206_));
 sg13g2_buf_1 _22913_ (.A(net533),
    .X(_05217_));
 sg13g2_nor2_1 _22914_ (.A(_00119_),
    .B(net482),
    .Y(_05218_));
 sg13g2_nor3_2 _22915_ (.A(_05213_),
    .B(_05216_),
    .C(_05218_),
    .Y(_05219_));
 sg13g2_nand2_1 _22916_ (.Y(_05220_),
    .A(\cpu.dcache.r_data[2][28] ),
    .B(_12340_));
 sg13g2_a22oi_1 _22917_ (.Y(_05221_),
    .B1(_09460_),
    .B2(\cpu.dcache.r_data[5][28] ),
    .A2(_09423_),
    .A1(\cpu.dcache.r_data[7][28] ));
 sg13g2_a22oi_1 _22918_ (.Y(_05222_),
    .B1(_10086_),
    .B2(\cpu.dcache.r_data[4][28] ),
    .A2(_12198_),
    .A1(\cpu.dcache.r_data[1][28] ));
 sg13g2_a22oi_1 _22919_ (.Y(_05223_),
    .B1(_12469_),
    .B2(\cpu.dcache.r_data[3][28] ),
    .A2(_09705_),
    .A1(\cpu.dcache.r_data[6][28] ));
 sg13g2_nand4_1 _22920_ (.B(_05221_),
    .C(_05222_),
    .A(_05220_),
    .Y(_05224_),
    .D(_05223_));
 sg13g2_nor2_1 _22921_ (.A(net594),
    .B(_05224_),
    .Y(_05225_));
 sg13g2_a21oi_1 _22922_ (.A1(_00118_),
    .A2(_04859_),
    .Y(_05226_),
    .B1(_05225_));
 sg13g2_nand2_1 _22923_ (.Y(_05227_),
    .A(net532),
    .B(_05226_));
 sg13g2_o21ai_1 _22924_ (.B1(_05227_),
    .Y(_05228_),
    .A1(net550),
    .A2(_05219_));
 sg13g2_a221oi_1 _22925_ (.B2(net662),
    .C1(net981),
    .B1(_05228_),
    .A1(_05149_),
    .Y(_05229_),
    .A2(_05210_));
 sg13g2_nor3_1 _22926_ (.A(net76),
    .B(_05127_),
    .C(_05229_),
    .Y(_05230_));
 sg13g2_a221oi_1 _22927_ (.B2(net617),
    .C1(_05230_),
    .B1(_03691_),
    .A1(_09157_),
    .Y(_05231_),
    .A2(_11485_));
 sg13g2_a221oi_1 _22928_ (.B2(_04331_),
    .C1(_05231_),
    .B1(_05205_),
    .A1(net114),
    .Y(_01021_),
    .A2(_05204_));
 sg13g2_nor2_1 _22929_ (.A(_08474_),
    .B(net152),
    .Y(_05232_));
 sg13g2_nor2_1 _22930_ (.A(net239),
    .B(net661),
    .Y(_05233_));
 sg13g2_nor2_1 _22931_ (.A(_11481_),
    .B(_04370_),
    .Y(_05234_));
 sg13g2_a21o_1 _22932_ (.A2(_05233_),
    .A1(_11841_),
    .B1(_05234_),
    .X(_05235_));
 sg13g2_a21o_1 _22933_ (.A2(_04367_),
    .A1(_05172_),
    .B1(_05235_),
    .X(_05236_));
 sg13g2_a22oi_1 _22934_ (.Y(_05237_),
    .B1(net449),
    .B2(\cpu.intr.r_timer_reload[13] ),
    .A2(net514),
    .A1(_10173_));
 sg13g2_a22oi_1 _22935_ (.Y(_05238_),
    .B1(net405),
    .B2(\cpu.intr.r_clock_cmp[13] ),
    .A2(net407),
    .A1(\cpu.intr.r_clock_cmp[29] ));
 sg13g2_buf_2 _22936_ (.A(\cpu.intr.r_clock_count[29] ),
    .X(_05239_));
 sg13g2_a22oi_1 _22937_ (.Y(_05240_),
    .B1(net446),
    .B2(\cpu.intr.r_timer_count[13] ),
    .A2(net362),
    .A1(_05239_));
 sg13g2_nand3_1 _22938_ (.B(_05238_),
    .C(_05240_),
    .A(_05237_),
    .Y(_05241_));
 sg13g2_mux2_1 _22939_ (.A0(\cpu.dcache.r_data[4][29] ),
    .A1(\cpu.dcache.r_data[6][29] ),
    .S(net516),
    .X(_05242_));
 sg13g2_a22oi_1 _22940_ (.Y(_05243_),
    .B1(_05242_),
    .B2(net540),
    .A2(net664),
    .A1(\cpu.dcache.r_data[7][29] ));
 sg13g2_nand2b_1 _22941_ (.Y(_05244_),
    .B(net613),
    .A_N(_05243_));
 sg13g2_mux2_1 _22942_ (.A0(\cpu.dcache.r_data[2][29] ),
    .A1(\cpu.dcache.r_data[3][29] ),
    .S(net558),
    .X(_05245_));
 sg13g2_a22oi_1 _22943_ (.Y(_05246_),
    .B1(_05245_),
    .B2(net790),
    .A2(_12702_),
    .A1(\cpu.dcache.r_data[5][29] ));
 sg13g2_nand2_1 _22944_ (.Y(_05247_),
    .A(\cpu.dcache.r_data[1][29] ),
    .B(_12199_));
 sg13g2_nand2b_1 _22945_ (.Y(_05248_),
    .B(_04859_),
    .A_N(_00124_));
 sg13g2_nand4_1 _22946_ (.B(_05246_),
    .C(_05247_),
    .A(_05244_),
    .Y(_05249_),
    .D(_05248_));
 sg13g2_buf_1 _22947_ (.A(_05249_),
    .X(_05250_));
 sg13g2_a22oi_1 _22948_ (.Y(_05251_),
    .B1(net559),
    .B2(\cpu.dcache.r_data[3][13] ),
    .A2(net556),
    .A1(\cpu.dcache.r_data[6][13] ));
 sg13g2_a22oi_1 _22949_ (.Y(_05252_),
    .B1(net484),
    .B2(\cpu.dcache.r_data[1][13] ),
    .A2(net560),
    .A1(\cpu.dcache.r_data[2][13] ));
 sg13g2_mux2_1 _22950_ (.A0(\cpu.dcache.r_data[5][13] ),
    .A1(\cpu.dcache.r_data[7][13] ),
    .S(net578),
    .X(_05253_));
 sg13g2_a22oi_1 _22951_ (.Y(_05254_),
    .B1(_05253_),
    .B2(net633),
    .A2(net921),
    .A1(\cpu.dcache.r_data[4][13] ));
 sg13g2_nand2b_1 _22952_ (.Y(_05255_),
    .B(net613),
    .A_N(_05254_));
 sg13g2_and4_1 _22953_ (.A(_05217_),
    .B(_05251_),
    .C(_05252_),
    .D(_05255_),
    .X(_05256_));
 sg13g2_a21oi_1 _22954_ (.A1(_00125_),
    .A2(_05129_),
    .Y(_05257_),
    .B1(_05256_));
 sg13g2_and2_1 _22955_ (.A(net685),
    .B(_05257_),
    .X(_05258_));
 sg13g2_a21o_1 _22956_ (.A2(_05250_),
    .A1(net623),
    .B1(_05258_),
    .X(_05259_));
 sg13g2_a22oi_1 _22957_ (.Y(_05260_),
    .B1(_05259_),
    .B2(net662),
    .A2(_05241_),
    .A1(_05149_));
 sg13g2_o21ai_1 _22958_ (.B1(net141),
    .Y(_05261_),
    .A1(_09213_),
    .A2(_05125_));
 sg13g2_inv_1 _22959_ (.Y(_05262_),
    .A(_05261_));
 sg13g2_o21ai_1 _22960_ (.B1(_05262_),
    .Y(_05263_),
    .A1(_05156_),
    .A2(_05260_));
 sg13g2_or2_1 _22961_ (.X(_05264_),
    .B(_05263_),
    .A(net76));
 sg13g2_o21ai_1 _22962_ (.B1(_05264_),
    .Y(_05265_),
    .A1(net493),
    .A2(_03557_));
 sg13g2_a221oi_1 _22963_ (.B2(_05166_),
    .C1(_05265_),
    .B1(_05236_),
    .A1(_05170_),
    .Y(_01022_),
    .A2(_05232_));
 sg13g2_a22oi_1 _22964_ (.Y(_05266_),
    .B1(net446),
    .B2(_09960_),
    .A2(net573),
    .A1(_10179_));
 sg13g2_a22oi_1 _22965_ (.Y(_05267_),
    .B1(_05153_),
    .B2(\cpu.intr.r_clock_cmp[14] ),
    .A2(_04938_),
    .A1(\cpu.intr.r_timer_reload[14] ));
 sg13g2_buf_1 _22966_ (.A(\cpu.intr.r_clock_count[30] ),
    .X(_05268_));
 sg13g2_a22oi_1 _22967_ (.Y(_05269_),
    .B1(_04934_),
    .B2(\cpu.intr.r_clock_cmp[30] ),
    .A2(net417),
    .A1(_05268_));
 sg13g2_nand3_1 _22968_ (.B(_05267_),
    .C(_05269_),
    .A(_05266_),
    .Y(_05270_));
 sg13g2_nand2_1 _22969_ (.Y(_05271_),
    .A(\cpu.dcache.r_data[2][30] ),
    .B(_12342_));
 sg13g2_a22oi_1 _22970_ (.Y(_05272_),
    .B1(net608),
    .B2(\cpu.dcache.r_data[5][30] ),
    .A2(_09946_),
    .A1(\cpu.dcache.r_data[7][30] ));
 sg13g2_a22oi_1 _22971_ (.Y(_05273_),
    .B1(_10086_),
    .B2(\cpu.dcache.r_data[4][30] ),
    .A2(_05132_),
    .A1(\cpu.dcache.r_data[1][30] ));
 sg13g2_a22oi_1 _22972_ (.Y(_05274_),
    .B1(_05134_),
    .B2(\cpu.dcache.r_data[3][30] ),
    .A2(net556),
    .A1(\cpu.dcache.r_data[6][30] ));
 sg13g2_nand4_1 _22973_ (.B(_05272_),
    .C(_05273_),
    .A(_05271_),
    .Y(_05275_),
    .D(_05274_));
 sg13g2_nand2_1 _22974_ (.Y(_05276_),
    .A(_00135_),
    .B(net531));
 sg13g2_o21ai_1 _22975_ (.B1(_05276_),
    .Y(_05277_),
    .A1(_05128_),
    .A2(_05275_));
 sg13g2_nand2_1 _22976_ (.Y(_05278_),
    .A(\cpu.dcache.r_data[2][14] ),
    .B(_12341_));
 sg13g2_a22oi_1 _22977_ (.Y(_05279_),
    .B1(net608),
    .B2(\cpu.dcache.r_data[5][14] ),
    .A2(net576),
    .A1(\cpu.dcache.r_data[7][14] ));
 sg13g2_a22oi_1 _22978_ (.Y(_05280_),
    .B1(net621),
    .B2(\cpu.dcache.r_data[4][14] ),
    .A2(net562),
    .A1(\cpu.dcache.r_data[1][14] ));
 sg13g2_a22oi_1 _22979_ (.Y(_05281_),
    .B1(net609),
    .B2(\cpu.dcache.r_data[3][14] ),
    .A2(_02691_),
    .A1(\cpu.dcache.r_data[6][14] ));
 sg13g2_nand4_1 _22980_ (.B(_05279_),
    .C(_05280_),
    .A(_05278_),
    .Y(_05282_),
    .D(_05281_));
 sg13g2_nor2_1 _22981_ (.A(net531),
    .B(_05282_),
    .Y(_05283_));
 sg13g2_a21oi_1 _22982_ (.A1(_00136_),
    .A2(net531),
    .Y(_05284_),
    .B1(_05283_));
 sg13g2_nand2_1 _22983_ (.Y(_05285_),
    .A(net685),
    .B(_05284_));
 sg13g2_o21ai_1 _22984_ (.B1(_05285_),
    .Y(_05286_),
    .A1(net622),
    .A2(_05277_));
 sg13g2_a22oi_1 _22985_ (.Y(_05287_),
    .B1(_05286_),
    .B2(net742),
    .A2(_05270_),
    .A1(_05149_));
 sg13g2_o21ai_1 _22986_ (.B1(_05262_),
    .Y(_05288_),
    .A1(net1144),
    .A2(_05287_));
 sg13g2_nor2_1 _22987_ (.A(_04211_),
    .B(_04411_),
    .Y(_05289_));
 sg13g2_a22oi_1 _22988_ (.Y(_05290_),
    .B1(net661),
    .B2(_05289_),
    .A2(net153),
    .A1(_08840_));
 sg13g2_nand3_1 _22989_ (.B(_05288_),
    .C(_05290_),
    .A(_03557_),
    .Y(_05291_));
 sg13g2_a221oi_1 _22990_ (.B2(_04408_),
    .C1(_05291_),
    .B1(_04405_),
    .A1(net190),
    .Y(_05292_),
    .A2(_11874_));
 sg13g2_mux2_1 _22991_ (.A0(_05288_),
    .A1(net688),
    .S(_03690_),
    .X(_05293_));
 sg13g2_nand2_1 _22992_ (.Y(_05294_),
    .A(_05288_),
    .B(_05290_));
 sg13g2_nor2b_1 _22993_ (.A(_05294_),
    .B_N(_03557_),
    .Y(_05295_));
 sg13g2_a22oi_1 _22994_ (.Y(_05296_),
    .B1(_05295_),
    .B2(_05010_),
    .A2(_05293_),
    .A1(net121));
 sg13g2_nand2b_1 _22995_ (.Y(_01023_),
    .B(_05296_),
    .A_N(_05292_));
 sg13g2_nor3_1 _22996_ (.A(net153),
    .B(net592),
    .C(net141),
    .Y(_05297_));
 sg13g2_nor2_1 _22997_ (.A(net529),
    .B(_04460_),
    .Y(_05298_));
 sg13g2_a22oi_1 _22998_ (.Y(_05299_),
    .B1(net449),
    .B2(\cpu.intr.r_timer_reload[15] ),
    .A2(net573),
    .A1(_10184_));
 sg13g2_a22oi_1 _22999_ (.Y(_05300_),
    .B1(net405),
    .B2(\cpu.intr.r_clock_cmp[15] ),
    .A2(net407),
    .A1(\cpu.intr.r_clock_cmp[31] ));
 sg13g2_buf_1 _23000_ (.A(\cpu.intr.r_clock_count[31] ),
    .X(_05301_));
 sg13g2_a22oi_1 _23001_ (.Y(_05302_),
    .B1(net446),
    .B2(\cpu.intr.r_timer_count[15] ),
    .A2(net362),
    .A1(_05301_));
 sg13g2_nand3_1 _23002_ (.B(_05300_),
    .C(_05302_),
    .A(_05299_),
    .Y(_05303_));
 sg13g2_inv_1 _23003_ (.Y(_05304_),
    .A(_05063_));
 sg13g2_nand2_1 _23004_ (.Y(_05305_),
    .A(net623),
    .B(_05304_));
 sg13g2_o21ai_1 _23005_ (.B1(_05305_),
    .Y(_05306_),
    .A1(net623),
    .A2(_05073_));
 sg13g2_a221oi_1 _23006_ (.B2(net742),
    .C1(net1144),
    .B1(_05306_),
    .A1(_05149_),
    .Y(_05307_),
    .A2(_05303_));
 sg13g2_nor3_1 _23007_ (.A(_03555_),
    .B(_05127_),
    .C(_05307_),
    .Y(_05308_));
 sg13g2_a21oi_1 _23008_ (.A1(net860),
    .A2(_03690_),
    .Y(_05309_),
    .B1(_05308_));
 sg13g2_nor3_1 _23009_ (.A(_08397_),
    .B(net152),
    .C(_03553_),
    .Y(_05310_));
 sg13g2_a21o_1 _23010_ (.A2(_05309_),
    .A1(net121),
    .B1(_05310_),
    .X(_05311_));
 sg13g2_a221oi_1 _23011_ (.B2(_05166_),
    .C1(_05311_),
    .B1(_05298_),
    .A1(_04458_),
    .Y(_01024_),
    .A2(_05297_));
 sg13g2_nor2_1 _23012_ (.A(_10644_),
    .B(_11481_),
    .Y(_05312_));
 sg13g2_a21oi_1 _23013_ (.A1(net529),
    .A2(_04206_),
    .Y(_05313_),
    .B1(_05312_));
 sg13g2_mux2_1 _23014_ (.A0(net1076),
    .A1(_05313_),
    .S(net152),
    .X(_05314_));
 sg13g2_a22oi_1 _23015_ (.Y(_05315_),
    .B1(net562),
    .B2(\cpu.dcache.r_data[1][1] ),
    .A2(net560),
    .A1(\cpu.dcache.r_data[2][1] ));
 sg13g2_a22oi_1 _23016_ (.Y(_05316_),
    .B1(net530),
    .B2(\cpu.dcache.r_data[3][1] ),
    .A2(net576),
    .A1(\cpu.dcache.r_data[7][1] ));
 sg13g2_mux2_1 _23017_ (.A0(\cpu.dcache.r_data[4][1] ),
    .A1(\cpu.dcache.r_data[6][1] ),
    .S(net632),
    .X(_05317_));
 sg13g2_a22oi_1 _23018_ (.Y(_05318_),
    .B1(_05317_),
    .B2(net600),
    .A2(net918),
    .A1(\cpu.dcache.r_data[5][1] ));
 sg13g2_nand2b_1 _23019_ (.Y(_05319_),
    .B(net673),
    .A_N(_05318_));
 sg13g2_nand4_1 _23020_ (.B(_05315_),
    .C(_05316_),
    .A(net482),
    .Y(_05320_),
    .D(_05319_));
 sg13g2_o21ai_1 _23021_ (.B1(_05320_),
    .Y(_05321_),
    .A1(\cpu.dcache.r_data[0][1] ),
    .A2(net482));
 sg13g2_inv_1 _23022_ (.Y(_05322_),
    .A(_05321_));
 sg13g2_a22oi_1 _23023_ (.Y(_05323_),
    .B1(net560),
    .B2(\cpu.dcache.r_data[2][17] ),
    .A2(net530),
    .A1(\cpu.dcache.r_data[3][17] ));
 sg13g2_a22oi_1 _23024_ (.Y(_05324_),
    .B1(net484),
    .B2(\cpu.dcache.r_data[1][17] ),
    .A2(net608),
    .A1(\cpu.dcache.r_data[5][17] ));
 sg13g2_mux2_1 _23025_ (.A0(\cpu.dcache.r_data[4][17] ),
    .A1(\cpu.dcache.r_data[6][17] ),
    .S(net578),
    .X(_05325_));
 sg13g2_a22oi_1 _23026_ (.Y(_05326_),
    .B1(_05325_),
    .B2(net600),
    .A2(net664),
    .A1(\cpu.dcache.r_data[7][17] ));
 sg13g2_nand2b_1 _23027_ (.Y(_05327_),
    .B(net673),
    .A_N(_05326_));
 sg13g2_and4_1 _23028_ (.A(net482),
    .B(_05323_),
    .C(_05324_),
    .D(_05327_),
    .X(_05328_));
 sg13g2_a21oi_1 _23029_ (.A1(_00299_),
    .A2(net485),
    .Y(_05329_),
    .B1(_05328_));
 sg13g2_nand2_1 _23030_ (.Y(_05330_),
    .A(_09944_),
    .B(_05329_));
 sg13g2_nor2_1 _23031_ (.A(net1025),
    .B(_05330_),
    .Y(_05331_));
 sg13g2_a21oi_1 _23032_ (.A1(net983),
    .A2(_05322_),
    .Y(_05332_),
    .B1(_05331_));
 sg13g2_a22oi_1 _23033_ (.Y(_05333_),
    .B1(_05134_),
    .B2(\cpu.dcache.r_data[3][9] ),
    .A2(_02691_),
    .A1(\cpu.dcache.r_data[6][9] ));
 sg13g2_a22oi_1 _23034_ (.Y(_05334_),
    .B1(_05132_),
    .B2(\cpu.dcache.r_data[1][9] ),
    .A2(_12341_),
    .A1(\cpu.dcache.r_data[2][9] ));
 sg13g2_mux2_1 _23035_ (.A0(\cpu.dcache.r_data[5][9] ),
    .A1(\cpu.dcache.r_data[7][9] ),
    .S(net578),
    .X(_05335_));
 sg13g2_a22oi_1 _23036_ (.Y(_05336_),
    .B1(_05335_),
    .B2(_09234_),
    .A2(net921),
    .A1(\cpu.dcache.r_data[4][9] ));
 sg13g2_nand2b_1 _23037_ (.Y(_05337_),
    .B(_11975_),
    .A_N(_05336_));
 sg13g2_and4_1 _23038_ (.A(_05217_),
    .B(_05333_),
    .C(_05334_),
    .D(_05337_),
    .X(_05338_));
 sg13g2_a21oi_1 _23039_ (.A1(_00301_),
    .A2(_05129_),
    .Y(_05339_),
    .B1(_05338_));
 sg13g2_and2_1 _23040_ (.A(_10041_),
    .B(_05339_),
    .X(_05340_));
 sg13g2_a22oi_1 _23041_ (.Y(_05341_),
    .B1(_12342_),
    .B2(\cpu.dcache.r_data[2][25] ),
    .A2(_12470_),
    .A1(\cpu.dcache.r_data[3][25] ));
 sg13g2_a22oi_1 _23042_ (.Y(_05342_),
    .B1(_12199_),
    .B2(\cpu.dcache.r_data[1][25] ),
    .A2(net608),
    .A1(\cpu.dcache.r_data[5][25] ));
 sg13g2_mux2_1 _23043_ (.A0(\cpu.dcache.r_data[4][25] ),
    .A1(\cpu.dcache.r_data[6][25] ),
    .S(net578),
    .X(_05343_));
 sg13g2_a22oi_1 _23044_ (.Y(_05344_),
    .B1(_05343_),
    .B2(net600),
    .A2(net664),
    .A1(\cpu.dcache.r_data[7][25] ));
 sg13g2_nand2b_1 _23045_ (.Y(_05345_),
    .B(_11976_),
    .A_N(_05344_));
 sg13g2_and4_1 _23046_ (.A(_05184_),
    .B(_05341_),
    .C(_05342_),
    .D(_05345_),
    .X(_05346_));
 sg13g2_a21oi_1 _23047_ (.A1(_00300_),
    .A2(net485),
    .Y(_05347_),
    .B1(_05346_));
 sg13g2_nor2b_1 _23048_ (.A(net1025),
    .B_N(_05347_),
    .Y(_05348_));
 sg13g2_nor3_1 _23049_ (.A(net663),
    .B(_05340_),
    .C(_05348_),
    .Y(_05349_));
 sg13g2_a21oi_1 _23050_ (.A1(net595),
    .A2(_05332_),
    .Y(_05350_),
    .B1(_05349_));
 sg13g2_o21ai_1 _23051_ (.B1(_05330_),
    .Y(_05351_),
    .A1(net532),
    .A2(_05321_));
 sg13g2_mux2_1 _23052_ (.A0(_05350_),
    .A1(_05351_),
    .S(net662),
    .X(_05352_));
 sg13g2_nor2_1 _23053_ (.A(net780),
    .B(_00092_),
    .Y(_05353_));
 sg13g2_buf_2 _23054_ (.A(\cpu.gpio.r_src_io[4][1] ),
    .X(_05354_));
 sg13g2_nor2b_1 _23055_ (.A(net781),
    .B_N(_05354_),
    .Y(_05355_));
 sg13g2_o21ai_1 _23056_ (.B1(net486),
    .Y(_05356_),
    .A1(_05353_),
    .A2(_05355_));
 sg13g2_o21ai_1 _23057_ (.B1(_05356_),
    .Y(_05357_),
    .A1(_00094_),
    .A2(_04904_));
 sg13g2_nand2_1 _23058_ (.Y(_05358_),
    .A(_11973_),
    .B(net487));
 sg13g2_nand2_1 _23059_ (.Y(_05359_),
    .A(_09181_),
    .B(net348));
 sg13g2_o21ai_1 _23060_ (.B1(_05359_),
    .Y(_05360_),
    .A1(_00093_),
    .A2(_05358_));
 sg13g2_nor2b_1 _23061_ (.A(_00096_),
    .B_N(_04924_),
    .Y(_05361_));
 sg13g2_nor2b_1 _23062_ (.A(_00095_),
    .B_N(net450),
    .Y(_05362_));
 sg13g2_nor4_1 _23063_ (.A(_05357_),
    .B(_05360_),
    .C(_05361_),
    .D(_05362_),
    .Y(_05363_));
 sg13g2_a21oi_1 _23064_ (.A1(_09181_),
    .A2(_04894_),
    .Y(_05364_),
    .B1(_04899_));
 sg13g2_nand2b_1 _23065_ (.Y(_05365_),
    .B(_09182_),
    .A_N(_05364_));
 sg13g2_a21oi_1 _23066_ (.A1(_05363_),
    .A2(_05365_),
    .Y(_05366_),
    .B1(_04884_));
 sg13g2_mux2_1 _23067_ (.A0(_11965_),
    .A1(_11970_),
    .S(net1030),
    .X(_05367_));
 sg13g2_a22oi_1 _23068_ (.Y(_05368_),
    .B1(_05367_),
    .B2(_04919_),
    .A2(_05116_),
    .A1(\cpu.spi.r_timeout[1] ));
 sg13g2_o21ai_1 _23069_ (.B1(_05368_),
    .Y(_05369_),
    .A1(_00302_),
    .A2(_04982_));
 sg13g2_inv_1 _23070_ (.Y(_05370_),
    .A(_00091_));
 sg13g2_buf_1 _23071_ (.A(_04973_),
    .X(_05371_));
 sg13g2_buf_1 _23072_ (.A(\cpu.spi.r_clk_count[2][1] ),
    .X(_05372_));
 sg13g2_a22oi_1 _23073_ (.Y(_05373_),
    .B1(_04985_),
    .B2(_05372_),
    .A2(net404),
    .A1(_05370_));
 sg13g2_nand2b_1 _23074_ (.Y(_05374_),
    .B(_05373_),
    .A_N(_05369_));
 sg13g2_a221oi_1 _23075_ (.B2(_09266_),
    .C1(_05374_),
    .B1(_04975_),
    .A1(_11966_),
    .Y(_05375_),
    .A2(net450));
 sg13g2_nor2_1 _23076_ (.A(_09225_),
    .B(_05375_),
    .Y(_05376_));
 sg13g2_a22oi_1 _23077_ (.Y(_05377_),
    .B1(net487),
    .B2(\cpu.uart.r_r_invert ),
    .A2(net448),
    .A1(_09166_));
 sg13g2_a22oi_1 _23078_ (.Y(_05378_),
    .B1(net445),
    .B2(\cpu.uart.r_div_value[9] ),
    .A2(_04919_),
    .A1(\cpu.uart.r_div_value[1] ));
 sg13g2_nand2_1 _23079_ (.Y(_05379_),
    .A(_05377_),
    .B(_05378_));
 sg13g2_a21oi_1 _23080_ (.A1(\cpu.uart.r_in[1] ),
    .A2(_04996_),
    .Y(_05380_),
    .B1(_05379_));
 sg13g2_a22oi_1 _23081_ (.Y(_05381_),
    .B1(net499),
    .B2(_09964_),
    .A2(net515),
    .A1(\cpu.intr.r_timer_reload[1] ));
 sg13g2_a221oi_1 _23082_ (.B2(_09958_),
    .C1(net780),
    .B1(net499),
    .A1(\cpu.intr.r_timer_reload[17] ),
    .Y(_05382_),
    .A2(net515));
 sg13g2_a21o_1 _23083_ (.A2(_05381_),
    .A1(net780),
    .B1(_05382_),
    .X(_05383_));
 sg13g2_buf_1 _23084_ (.A(\cpu.intr.r_clock_count[17] ),
    .X(_05384_));
 sg13g2_a22oi_1 _23085_ (.Y(_05385_),
    .B1(_04897_),
    .B2(_09169_),
    .A2(net417),
    .A1(_05384_));
 sg13g2_nand2_1 _23086_ (.Y(_05386_),
    .A(\cpu.intr.r_clock_cmp[17] ),
    .B(_04934_));
 sg13g2_a22oi_1 _23087_ (.Y(_05387_),
    .B1(_05080_),
    .B2(\cpu.intr.r_clock_cmp[1] ),
    .A2(net573),
    .A1(_10103_));
 sg13g2_nand4_1 _23088_ (.B(_05385_),
    .C(_05386_),
    .A(_05383_),
    .Y(_05388_),
    .D(_05387_));
 sg13g2_a21oi_1 _23089_ (.A1(_09169_),
    .A2(net347),
    .Y(_05389_),
    .B1(net447));
 sg13g2_nor2b_1 _23090_ (.A(_05389_),
    .B_N(\cpu.intr.r_clock ),
    .Y(_05390_));
 sg13g2_o21ai_1 _23091_ (.B1(_04932_),
    .Y(_05391_),
    .A1(_05388_),
    .A2(_05390_));
 sg13g2_o21ai_1 _23092_ (.B1(_05391_),
    .Y(_05392_),
    .A1(net593),
    .A2(_05380_));
 sg13g2_nor3_1 _23093_ (.A(_05366_),
    .B(_05376_),
    .C(_05392_),
    .Y(_05393_));
 sg13g2_nand2_1 _23094_ (.Y(_05394_),
    .A(net855),
    .B(_05393_));
 sg13g2_o21ai_1 _23095_ (.B1(_05394_),
    .Y(_05395_),
    .A1(net855),
    .A2(_05352_));
 sg13g2_nor2_1 _23096_ (.A(net75),
    .B(_05395_),
    .Y(_05396_));
 sg13g2_a221oi_1 _23097_ (.B2(_03507_),
    .C1(_05396_),
    .B1(net36),
    .A1(net708),
    .Y(_05397_),
    .A2(_11485_));
 sg13g2_a21oi_1 _23098_ (.A1(net114),
    .A2(_05314_),
    .Y(_01025_),
    .B1(_05397_));
 sg13g2_a22oi_1 _23099_ (.Y(_05398_),
    .B1(net530),
    .B2(\cpu.dcache.r_data[3][18] ),
    .A2(net556),
    .A1(\cpu.dcache.r_data[6][18] ));
 sg13g2_a22oi_1 _23100_ (.Y(_05399_),
    .B1(net484),
    .B2(\cpu.dcache.r_data[1][18] ),
    .A2(net560),
    .A1(\cpu.dcache.r_data[2][18] ));
 sg13g2_mux2_1 _23101_ (.A0(\cpu.dcache.r_data[5][18] ),
    .A1(\cpu.dcache.r_data[7][18] ),
    .S(net578),
    .X(_05400_));
 sg13g2_a22oi_1 _23102_ (.Y(_05401_),
    .B1(_05400_),
    .B2(net633),
    .A2(net921),
    .A1(\cpu.dcache.r_data[4][18] ));
 sg13g2_nand2b_1 _23103_ (.Y(_05402_),
    .B(net673),
    .A_N(_05401_));
 sg13g2_and4_1 _23104_ (.A(net482),
    .B(_05398_),
    .C(_05399_),
    .D(_05402_),
    .X(_05403_));
 sg13g2_a21oi_1 _23105_ (.A1(_00097_),
    .A2(net531),
    .Y(_05404_),
    .B1(_05403_));
 sg13g2_nand2_1 _23106_ (.Y(_05405_),
    .A(_12124_),
    .B(_05404_));
 sg13g2_a22oi_1 _23107_ (.Y(_05406_),
    .B1(net530),
    .B2(\cpu.dcache.r_data[3][2] ),
    .A2(net556),
    .A1(\cpu.dcache.r_data[6][2] ));
 sg13g2_a22oi_1 _23108_ (.Y(_05407_),
    .B1(net621),
    .B2(\cpu.dcache.r_data[4][2] ),
    .A2(net560),
    .A1(\cpu.dcache.r_data[2][2] ));
 sg13g2_mux2_1 _23109_ (.A0(\cpu.dcache.r_data[5][2] ),
    .A1(\cpu.dcache.r_data[7][2] ),
    .S(net516),
    .X(_05408_));
 sg13g2_a22oi_1 _23110_ (.Y(_05409_),
    .B1(_05408_),
    .B2(net689),
    .A2(net484),
    .A1(\cpu.dcache.r_data[1][2] ));
 sg13g2_nand4_1 _23111_ (.B(_05406_),
    .C(_05407_),
    .A(net482),
    .Y(_05410_),
    .D(_05409_));
 sg13g2_o21ai_1 _23112_ (.B1(_05410_),
    .Y(_05411_),
    .A1(\cpu.dcache.r_data[0][2] ),
    .A2(net483));
 sg13g2_mux2_1 _23113_ (.A0(_05405_),
    .A1(_05411_),
    .S(net983),
    .X(_05412_));
 sg13g2_nor2b_1 _23114_ (.A(net1025),
    .B_N(_05138_),
    .Y(_05413_));
 sg13g2_nor3_1 _23115_ (.A(net595),
    .B(_05146_),
    .C(_05413_),
    .Y(_05414_));
 sg13g2_a21oi_1 _23116_ (.A1(net595),
    .A2(_05412_),
    .Y(_05415_),
    .B1(_05414_));
 sg13g2_o21ai_1 _23117_ (.B1(_05405_),
    .Y(_05416_),
    .A1(net532),
    .A2(_05411_));
 sg13g2_mux2_1 _23118_ (.A0(_05415_),
    .A1(_05416_),
    .S(net662),
    .X(_05417_));
 sg13g2_nand2_1 _23119_ (.Y(_05418_),
    .A(_09190_),
    .B(_04899_));
 sg13g2_o21ai_1 _23120_ (.B1(_05418_),
    .Y(_05419_),
    .A1(_00104_),
    .A2(_04904_));
 sg13g2_nor2_1 _23121_ (.A(net685),
    .B(_00102_),
    .Y(_05420_));
 sg13g2_buf_1 _23122_ (.A(\cpu.gpio.r_src_io[4][2] ),
    .X(_05421_));
 sg13g2_nor2b_1 _23123_ (.A(net612),
    .B_N(_05421_),
    .Y(_05422_));
 sg13g2_o21ai_1 _23124_ (.B1(net486),
    .Y(_05423_),
    .A1(_05420_),
    .A2(_05422_));
 sg13g2_o21ai_1 _23125_ (.B1(_05423_),
    .Y(_05424_),
    .A1(_00103_),
    .A2(_05358_));
 sg13g2_inv_1 _23126_ (.Y(_05425_),
    .A(_00106_));
 sg13g2_nor2b_1 _23127_ (.A(_00105_),
    .B_N(net450),
    .Y(_05426_));
 sg13g2_a21o_1 _23128_ (.A2(_04924_),
    .A1(_05425_),
    .B1(_05426_),
    .X(_05427_));
 sg13g2_a21oi_1 _23129_ (.A1(_09190_),
    .A2(_04894_),
    .Y(_05428_),
    .B1(net348));
 sg13g2_nor2b_1 _23130_ (.A(_05428_),
    .B_N(\cpu.gpio.r_enable_in[2] ),
    .Y(_05429_));
 sg13g2_nor4_1 _23131_ (.A(_05419_),
    .B(_05424_),
    .C(_05427_),
    .D(_05429_),
    .Y(_05430_));
 sg13g2_mux2_1 _23132_ (.A0(\cpu.intr.r_timer_reload[2] ),
    .A1(\cpu.intr.r_timer_reload[18] ),
    .S(net686),
    .X(_05431_));
 sg13g2_a22oi_1 _23133_ (.Y(_05432_),
    .B1(_05431_),
    .B2(net515),
    .A2(net448),
    .A1(_09162_));
 sg13g2_buf_1 _23134_ (.A(\cpu.intr.r_clock_count[18] ),
    .X(_05433_));
 sg13g2_a22oi_1 _23135_ (.Y(_05434_),
    .B1(net447),
    .B2(_09161_),
    .A2(_10116_),
    .A1(_05433_));
 sg13g2_a22oi_1 _23136_ (.Y(_05435_),
    .B1(_04940_),
    .B2(_10108_),
    .A2(_04939_),
    .A1(_09957_));
 sg13g2_inv_1 _23137_ (.Y(_05436_),
    .A(_05435_));
 sg13g2_a22oi_1 _23138_ (.Y(_05437_),
    .B1(_05436_),
    .B2(net915),
    .A2(_04935_),
    .A1(\cpu.intr.r_clock_cmp[18] ));
 sg13g2_a22oi_1 _23139_ (.Y(_05438_),
    .B1(net557),
    .B2(\cpu.intr.r_clock_cmp[2] ),
    .A2(net499),
    .A1(_09966_));
 sg13g2_nand3_1 _23140_ (.B(_09162_),
    .C(net347),
    .A(_09161_),
    .Y(_05439_));
 sg13g2_o21ai_1 _23141_ (.B1(_05439_),
    .Y(_05440_),
    .A1(net612),
    .A2(_05438_));
 sg13g2_inv_1 _23142_ (.Y(_05441_),
    .A(_05440_));
 sg13g2_nand4_1 _23143_ (.B(_05434_),
    .C(_05437_),
    .A(_05432_),
    .Y(_05442_),
    .D(_05441_));
 sg13g2_nand2b_1 _23144_ (.Y(_05443_),
    .B(net450),
    .A_N(_00267_));
 sg13g2_inv_1 _23145_ (.Y(_05444_),
    .A(_00101_));
 sg13g2_buf_1 _23146_ (.A(\cpu.spi.r_clk_count[2][2] ),
    .X(_05445_));
 sg13g2_nand2_1 _23147_ (.Y(_05446_),
    .A(net1030),
    .B(_11953_));
 sg13g2_o21ai_1 _23148_ (.B1(_05446_),
    .Y(_05447_),
    .A1(net1030),
    .A2(_00266_));
 sg13g2_a22oi_1 _23149_ (.Y(_05448_),
    .B1(_05447_),
    .B2(_04919_),
    .A2(_05116_),
    .A1(\cpu.spi.r_timeout[2] ));
 sg13g2_o21ai_1 _23150_ (.B1(_05448_),
    .Y(_05449_),
    .A1(_00100_),
    .A2(_04982_));
 sg13g2_a221oi_1 _23151_ (.B2(_05445_),
    .C1(_05449_),
    .B1(_04985_),
    .A1(_05444_),
    .Y(_05450_),
    .A2(net404));
 sg13g2_nand2_1 _23152_ (.Y(_05451_),
    .A(_09270_),
    .B(_04975_));
 sg13g2_nand3_1 _23153_ (.B(_05450_),
    .C(_05451_),
    .A(_05443_),
    .Y(_05452_));
 sg13g2_and2_1 _23154_ (.A(\cpu.uart.r_in[2] ),
    .B(_04996_),
    .X(_05453_));
 sg13g2_a221oi_1 _23155_ (.B2(_09933_),
    .C1(_05453_),
    .B1(net445),
    .A1(\cpu.uart.r_div_value[2] ),
    .Y(_05454_),
    .A2(net406));
 sg13g2_o21ai_1 _23156_ (.B1(net1026),
    .Y(_05455_),
    .A1(net593),
    .A2(_05454_));
 sg13g2_a221oi_1 _23157_ (.B2(_04992_),
    .C1(_05455_),
    .B1(_05452_),
    .A1(_04932_),
    .Y(_05456_),
    .A2(_05442_));
 sg13g2_o21ai_1 _23158_ (.B1(_05456_),
    .Y(_05457_),
    .A1(_04884_),
    .A2(_05430_));
 sg13g2_o21ai_1 _23159_ (.B1(_05457_),
    .Y(_05458_),
    .A1(net855),
    .A2(_05417_));
 sg13g2_nand2_1 _23160_ (.Y(_05459_),
    .A(net491),
    .B(net75));
 sg13g2_o21ai_1 _23161_ (.B1(_05459_),
    .Y(_05460_),
    .A1(net36),
    .A2(_05458_));
 sg13g2_o21ai_1 _23162_ (.B1(_04100_),
    .Y(_05461_),
    .A1(net804),
    .A2(net529));
 sg13g2_nand3_1 _23163_ (.B(net804),
    .C(net661),
    .A(net808),
    .Y(_05462_));
 sg13g2_o21ai_1 _23164_ (.B1(_05462_),
    .Y(_05463_),
    .A1(net592),
    .A2(_04499_));
 sg13g2_a221oi_1 _23165_ (.B2(net152),
    .C1(_03689_),
    .B1(_05463_),
    .A1(net805),
    .Y(_05464_),
    .A2(_05461_));
 sg13g2_a21o_1 _23166_ (.A2(_05460_),
    .A1(net115),
    .B1(_05464_),
    .X(_01026_));
 sg13g2_buf_1 _23167_ (.A(net121),
    .X(_05465_));
 sg13g2_mux2_1 _23168_ (.A0(\cpu.dcache.r_data[5][19] ),
    .A1(\cpu.dcache.r_data[7][19] ),
    .S(_09297_),
    .X(_05466_));
 sg13g2_a22oi_1 _23169_ (.Y(_05467_),
    .B1(_05466_),
    .B2(net558),
    .A2(net785),
    .A1(\cpu.dcache.r_data[6][19] ));
 sg13g2_nand2b_1 _23170_ (.Y(_05468_),
    .B(_11976_),
    .A_N(_05467_));
 sg13g2_mux2_1 _23171_ (.A0(\cpu.dcache.r_data[2][19] ),
    .A1(\cpu.dcache.r_data[3][19] ),
    .S(net558),
    .X(_05469_));
 sg13g2_a22oi_1 _23172_ (.Y(_05470_),
    .B1(_05469_),
    .B2(net790),
    .A2(net574),
    .A1(\cpu.dcache.r_data[4][19] ));
 sg13g2_nand2_1 _23173_ (.Y(_05471_),
    .A(\cpu.dcache.r_data[1][19] ),
    .B(net503));
 sg13g2_nand2b_1 _23174_ (.Y(_05472_),
    .B(net531),
    .A_N(_00107_));
 sg13g2_nand4_1 _23175_ (.B(_05470_),
    .C(_05471_),
    .A(_05468_),
    .Y(_05473_),
    .D(_05472_));
 sg13g2_nand2_1 _23176_ (.Y(_05474_),
    .A(net612),
    .B(_05473_));
 sg13g2_a22oi_1 _23177_ (.Y(_05475_),
    .B1(net503),
    .B2(\cpu.dcache.r_data[1][3] ),
    .A2(_02692_),
    .A1(\cpu.dcache.r_data[6][3] ));
 sg13g2_a22oi_1 _23178_ (.Y(_05476_),
    .B1(_10087_),
    .B2(\cpu.dcache.r_data[4][3] ),
    .A2(net559),
    .A1(\cpu.dcache.r_data[3][3] ));
 sg13g2_mux2_1 _23179_ (.A0(\cpu.dcache.r_data[5][3] ),
    .A1(\cpu.dcache.r_data[7][3] ),
    .S(net516),
    .X(_05477_));
 sg13g2_a22oi_1 _23180_ (.Y(_05478_),
    .B1(_05477_),
    .B2(net689),
    .A2(net502),
    .A1(\cpu.dcache.r_data[2][3] ));
 sg13g2_nand4_1 _23181_ (.B(_05475_),
    .C(_05476_),
    .A(net483),
    .Y(_05479_),
    .D(_05478_));
 sg13g2_o21ai_1 _23182_ (.B1(_05479_),
    .Y(_05480_),
    .A1(\cpu.dcache.r_data[0][3] ),
    .A2(net483));
 sg13g2_mux2_1 _23183_ (.A0(_05474_),
    .A1(_05480_),
    .S(net1025),
    .X(_05481_));
 sg13g2_nor2b_1 _23184_ (.A(net1025),
    .B_N(_05182_),
    .Y(_05482_));
 sg13g2_nor3_1 _23185_ (.A(_04857_),
    .B(_05192_),
    .C(_05482_),
    .Y(_05483_));
 sg13g2_a21oi_1 _23186_ (.A1(net595),
    .A2(_05481_),
    .Y(_05484_),
    .B1(_05483_));
 sg13g2_o21ai_1 _23187_ (.B1(_05474_),
    .Y(_05485_),
    .A1(net532),
    .A2(_05480_));
 sg13g2_mux2_1 _23188_ (.A0(_05484_),
    .A1(_05485_),
    .S(net742),
    .X(_05486_));
 sg13g2_buf_1 _23189_ (.A(\cpu.spi.r_clk_count[2][3] ),
    .X(_05487_));
 sg13g2_nor2_1 _23190_ (.A(_00111_),
    .B(_05091_),
    .Y(_05488_));
 sg13g2_a221oi_1 _23191_ (.B2(\cpu.spi.r_timeout[3] ),
    .C1(_05488_),
    .B1(_05116_),
    .A1(_05487_),
    .Y(_05489_),
    .A2(_04985_));
 sg13g2_o21ai_1 _23192_ (.B1(_05489_),
    .Y(_05490_),
    .A1(_00110_),
    .A2(_04982_));
 sg13g2_a21oi_1 _23193_ (.A1(_09264_),
    .A2(_04975_),
    .Y(_05491_),
    .B1(_05490_));
 sg13g2_nand3_1 _23194_ (.B(_09198_),
    .C(_04894_),
    .A(_09197_),
    .Y(_05492_));
 sg13g2_buf_1 _23195_ (.A(\cpu.gpio.r_src_io[4][3] ),
    .X(_05493_));
 sg13g2_nand2_1 _23196_ (.Y(_05494_),
    .A(net780),
    .B(_05493_));
 sg13g2_o21ai_1 _23197_ (.B1(_05494_),
    .Y(_05495_),
    .A1(net685),
    .A2(_00112_));
 sg13g2_inv_1 _23198_ (.Y(_05496_),
    .A(_00115_));
 sg13g2_a22oi_1 _23199_ (.Y(_05497_),
    .B1(_04934_),
    .B2(_05496_),
    .A2(net573),
    .A1(\cpu.gpio.genblk1[3].srcs_o[0] ));
 sg13g2_nand2b_1 _23200_ (.Y(_05498_),
    .B(net408),
    .A_N(_00113_));
 sg13g2_o21ai_1 _23201_ (.B1(_05498_),
    .Y(_05499_),
    .A1(_00114_),
    .A2(_04904_));
 sg13g2_a21oi_1 _23202_ (.A1(_09197_),
    .A2(net348),
    .Y(_05500_),
    .B1(_05499_));
 sg13g2_o21ai_1 _23203_ (.B1(_05500_),
    .Y(_05501_),
    .A1(_04902_),
    .A2(_05497_));
 sg13g2_a221oi_1 _23204_ (.B2(net486),
    .C1(_05501_),
    .B1(_05495_),
    .A1(_09198_),
    .Y(_05502_),
    .A2(_04899_));
 sg13g2_a21oi_1 _23205_ (.A1(_05492_),
    .A2(_05502_),
    .Y(_05503_),
    .B1(_04884_));
 sg13g2_mux4_1 _23206_ (.S0(net781),
    .A0(\cpu.intr.r_clock_cmp[3] ),
    .A1(\cpu.intr.r_clock_cmp[19] ),
    .A2(\cpu.intr.r_timer_reload[3] ),
    .A3(\cpu.intr.r_timer_reload[19] ),
    .S1(net463),
    .X(_05504_));
 sg13g2_inv_1 _23207_ (.Y(_05505_),
    .A(_09163_));
 sg13g2_buf_1 _23208_ (.A(\cpu.intr.r_clock_count[19] ),
    .X(_05506_));
 sg13g2_mux2_1 _23209_ (.A0(\cpu.intr.r_timer_count[3] ),
    .A1(_09956_),
    .S(net781),
    .X(_05507_));
 sg13g2_a22oi_1 _23210_ (.Y(_05508_),
    .B1(_05507_),
    .B2(net499),
    .A2(net417),
    .A1(_05506_));
 sg13g2_o21ai_1 _23211_ (.B1(_05508_),
    .Y(_05509_),
    .A1(_05505_),
    .A2(_05084_));
 sg13g2_a221oi_1 _23212_ (.B2(net689),
    .C1(_05509_),
    .B1(_05504_),
    .A1(_10122_),
    .Y(_05510_),
    .A2(net573));
 sg13g2_a21oi_1 _23213_ (.A1(_09163_),
    .A2(net347),
    .Y(_05511_),
    .B1(net448));
 sg13g2_nand2b_1 _23214_ (.Y(_05512_),
    .B(\cpu.intr.r_enable[3] ),
    .A_N(_05511_));
 sg13g2_a21oi_1 _23215_ (.A1(_05510_),
    .A2(_05512_),
    .Y(_05513_),
    .B1(_09951_));
 sg13g2_and2_1 _23216_ (.A(\cpu.uart.r_in[3] ),
    .B(_04996_),
    .X(_05514_));
 sg13g2_a221oi_1 _23217_ (.B2(\cpu.uart.r_div_value[11] ),
    .C1(_05514_),
    .B1(_04998_),
    .A1(\cpu.uart.r_div_value[3] ),
    .Y(_05515_),
    .A2(net406));
 sg13g2_o21ai_1 _23218_ (.B1(net1026),
    .Y(_05516_),
    .A1(net593),
    .A2(_05515_));
 sg13g2_nor3_1 _23219_ (.A(_05503_),
    .B(_05513_),
    .C(_05516_),
    .Y(_05517_));
 sg13g2_o21ai_1 _23220_ (.B1(_05517_),
    .Y(_05518_),
    .A1(_09225_),
    .A2(_05491_));
 sg13g2_o21ai_1 _23221_ (.B1(_05518_),
    .Y(_05519_),
    .A1(net855),
    .A2(_05486_));
 sg13g2_nor2_1 _23222_ (.A(net75),
    .B(_05519_),
    .Y(_05520_));
 sg13g2_a21oi_1 _23223_ (.A1(net463),
    .A2(net36),
    .Y(_05521_),
    .B1(_05520_));
 sg13g2_a21o_1 _23224_ (.A2(_04531_),
    .A1(net592),
    .B1(net153),
    .X(_05522_));
 sg13g2_nand2_1 _23225_ (.Y(_05523_),
    .A(net661),
    .B(_04533_));
 sg13g2_o21ai_1 _23226_ (.B1(_05523_),
    .Y(_05524_),
    .A1(net592),
    .A2(_04530_));
 sg13g2_a221oi_1 _23227_ (.B2(_05168_),
    .C1(_03689_),
    .B1(_05524_),
    .A1(net710),
    .Y(_05525_),
    .A2(_05522_));
 sg13g2_a21oi_1 _23228_ (.A1(net104),
    .A2(_05521_),
    .Y(_01027_),
    .B1(_05525_));
 sg13g2_o21ai_1 _23229_ (.B1(net152),
    .Y(_05526_),
    .A1(net529),
    .A2(_04277_));
 sg13g2_nand2_1 _23230_ (.Y(_05527_),
    .A(net661),
    .B(_04571_));
 sg13g2_o21ai_1 _23231_ (.B1(_05527_),
    .Y(_05528_),
    .A1(net592),
    .A2(_04569_));
 sg13g2_a22oi_1 _23232_ (.Y(_05529_),
    .B1(_05528_),
    .B2(net130),
    .A2(_05526_),
    .A1(net1141));
 sg13g2_buf_1 _23233_ (.A(\cpu.spi.r_clk_count[2][4] ),
    .X(_05530_));
 sg13g2_nor2_1 _23234_ (.A(_00121_),
    .B(_05091_),
    .Y(_05531_));
 sg13g2_a221oi_1 _23235_ (.B2(\cpu.spi.r_timeout[4] ),
    .C1(_05531_),
    .B1(_05116_),
    .A1(_05530_),
    .Y(_05532_),
    .A2(_04985_));
 sg13g2_o21ai_1 _23236_ (.B1(_05532_),
    .Y(_05533_),
    .A1(_00120_),
    .A2(_04982_));
 sg13g2_a21o_1 _23237_ (.A2(_04975_),
    .A1(_09272_),
    .B1(_05533_),
    .X(_05534_));
 sg13g2_inv_1 _23238_ (.Y(_05535_),
    .A(_09203_));
 sg13g2_mux2_1 _23239_ (.A0(\cpu.intr.r_clock_cmp[20] ),
    .A1(\cpu.intr.r_timer_reload[20] ),
    .S(net516),
    .X(_05536_));
 sg13g2_a22oi_1 _23240_ (.Y(_05537_),
    .B1(_05536_),
    .B2(net558),
    .A2(net785),
    .A1(_09985_));
 sg13g2_o21ai_1 _23241_ (.B1(net781),
    .Y(_05538_),
    .A1(net783),
    .A2(_05537_));
 sg13g2_a21o_1 _23242_ (.A2(net557),
    .A1(\cpu.intr.r_clock_cmp[4] ),
    .B1(net781),
    .X(_05539_));
 sg13g2_nand2_1 _23243_ (.Y(_05540_),
    .A(\cpu.intr.r_timer_reload[4] ),
    .B(_04937_));
 sg13g2_buf_2 _23244_ (.A(\cpu.intr.r_clock_count[20] ),
    .X(_05541_));
 sg13g2_a22oi_1 _23245_ (.Y(_05542_),
    .B1(_04897_),
    .B2(_09203_),
    .A2(net417),
    .A1(_05541_));
 sg13g2_a221oi_1 _23246_ (.B2(_09963_),
    .C1(net347),
    .B1(_04960_),
    .A1(_10127_),
    .Y(_05543_),
    .A2(net573));
 sg13g2_nand3_1 _23247_ (.B(_05542_),
    .C(_05543_),
    .A(_05540_),
    .Y(_05544_));
 sg13g2_a21oi_1 _23248_ (.A1(_05538_),
    .A2(_05539_),
    .Y(_05545_),
    .B1(_05544_));
 sg13g2_a221oi_1 _23249_ (.B2(_05084_),
    .C1(_09951_),
    .B1(_05545_),
    .A1(_05535_),
    .Y(_05546_),
    .A2(_04953_));
 sg13g2_and2_1 _23250_ (.A(_09184_),
    .B(_09202_),
    .X(_05547_));
 sg13g2_o21ai_1 _23251_ (.B1(_05547_),
    .Y(_05548_),
    .A1(net347),
    .A2(_05545_));
 sg13g2_nand2b_1 _23252_ (.Y(_05549_),
    .B(_04894_),
    .A_N(_09178_));
 sg13g2_buf_2 _23253_ (.A(\cpu.gpio.r_spi_miso_src[1][0] ),
    .X(_05550_));
 sg13g2_a22oi_1 _23254_ (.Y(_05551_),
    .B1(_04934_),
    .B2(_05550_),
    .A2(_10094_),
    .A1(\cpu.gpio.genblk1[4].srcs_o[0] ));
 sg13g2_a22oi_1 _23255_ (.Y(_05552_),
    .B1(_05080_),
    .B2(net7),
    .A2(net487),
    .A1(_09200_));
 sg13g2_a21oi_1 _23256_ (.A1(_05551_),
    .A2(_05552_),
    .Y(_05553_),
    .B1(_04902_));
 sg13g2_buf_2 _23257_ (.A(\cpu.gpio.r_src_io[5][0] ),
    .X(_05554_));
 sg13g2_buf_2 _23258_ (.A(\cpu.gpio.r_src_io[7][0] ),
    .X(_05555_));
 sg13g2_mux2_1 _23259_ (.A0(_05554_),
    .A1(_05555_),
    .S(net914),
    .X(_05556_));
 sg13g2_a22oi_1 _23260_ (.Y(_05557_),
    .B1(_05556_),
    .B2(net486),
    .A2(net404),
    .A1(_09199_));
 sg13g2_a22oi_1 _23261_ (.Y(_05558_),
    .B1(_04899_),
    .B2(_09177_),
    .A2(net348),
    .A1(\cpu.gpio.r_enable_in[4] ));
 sg13g2_buf_2 _23262_ (.A(\cpu.gpio.r_src_o[7][0] ),
    .X(_05559_));
 sg13g2_buf_2 _23263_ (.A(\cpu.gpio.r_src_o[3][0] ),
    .X(_05560_));
 sg13g2_inv_1 _23264_ (.Y(_05561_),
    .A(_05560_));
 sg13g2_nand3_1 _23265_ (.B(_09200_),
    .C(net982),
    .A(_09199_),
    .Y(_05562_));
 sg13g2_o21ai_1 _23266_ (.B1(_05562_),
    .Y(_05563_),
    .A1(net1043),
    .A2(_05561_));
 sg13g2_buf_2 _23267_ (.A(\cpu.gpio.r_src_o[5][0] ),
    .X(_05564_));
 sg13g2_nand2_1 _23268_ (.Y(_05565_),
    .A(_05564_),
    .B(_04897_));
 sg13g2_nand3_1 _23269_ (.B(\cpu.gpio.genblk2[4].srcs_io[0] ),
    .C(_10114_),
    .A(net982),
    .Y(_05566_));
 sg13g2_o21ai_1 _23270_ (.B1(_05566_),
    .Y(_05567_),
    .A1(net982),
    .A2(_05565_));
 sg13g2_a221oi_1 _23271_ (.B2(_05563_),
    .C1(_05567_),
    .B1(net447),
    .A1(_05559_),
    .Y(_05568_),
    .A2(net408));
 sg13g2_nand3_1 _23272_ (.B(_05558_),
    .C(_05568_),
    .A(_05557_),
    .Y(_05569_));
 sg13g2_nor2_1 _23273_ (.A(_05553_),
    .B(_05569_),
    .Y(_05570_));
 sg13g2_a21oi_1 _23274_ (.A1(_05549_),
    .A2(_05570_),
    .Y(_05571_),
    .B1(_04884_));
 sg13g2_a221oi_1 _23275_ (.B2(_05548_),
    .C1(_05571_),
    .B1(_05546_),
    .A1(_04992_),
    .Y(_05572_),
    .A2(_05534_));
 sg13g2_a221oi_1 _23276_ (.B2(\cpu.uart.r_in[4] ),
    .C1(net593),
    .B1(_04996_),
    .A1(\cpu.uart.r_div_value[4] ),
    .Y(_05573_),
    .A2(net406));
 sg13g2_a21oi_1 _23277_ (.A1(_04994_),
    .A2(_05572_),
    .Y(_05574_),
    .B1(_05573_));
 sg13g2_mux2_1 _23278_ (.A0(\cpu.dcache.r_data[4][20] ),
    .A1(\cpu.dcache.r_data[6][20] ),
    .S(net516),
    .X(_05575_));
 sg13g2_a22oi_1 _23279_ (.Y(_05576_),
    .B1(_05575_),
    .B2(net540),
    .A2(net664),
    .A1(\cpu.dcache.r_data[7][20] ));
 sg13g2_nand2b_1 _23280_ (.Y(_05577_),
    .B(net613),
    .A_N(_05576_));
 sg13g2_mux2_1 _23281_ (.A0(\cpu.dcache.r_data[2][20] ),
    .A1(\cpu.dcache.r_data[3][20] ),
    .S(net558),
    .X(_05578_));
 sg13g2_a22oi_1 _23282_ (.Y(_05579_),
    .B1(_05578_),
    .B2(net790),
    .A2(net557),
    .A1(\cpu.dcache.r_data[5][20] ));
 sg13g2_nand2_1 _23283_ (.Y(_05580_),
    .A(\cpu.dcache.r_data[1][20] ),
    .B(net503));
 sg13g2_nand2b_1 _23284_ (.Y(_05581_),
    .B(net531),
    .A_N(_00117_));
 sg13g2_nand4_1 _23285_ (.B(_05579_),
    .C(_05580_),
    .A(_05577_),
    .Y(_05582_),
    .D(_05581_));
 sg13g2_and2_1 _23286_ (.A(net622),
    .B(_04880_),
    .X(_05583_));
 sg13g2_a22oi_1 _23287_ (.Y(_05584_),
    .B1(net502),
    .B2(\cpu.dcache.r_data[2][4] ),
    .A2(net559),
    .A1(\cpu.dcache.r_data[3][4] ));
 sg13g2_a22oi_1 _23288_ (.Y(_05585_),
    .B1(net503),
    .B2(\cpu.dcache.r_data[1][4] ),
    .A2(_12703_),
    .A1(\cpu.dcache.r_data[5][4] ));
 sg13g2_mux2_1 _23289_ (.A0(\cpu.dcache.r_data[4][4] ),
    .A1(\cpu.dcache.r_data[6][4] ),
    .S(net516),
    .X(_05586_));
 sg13g2_a22oi_1 _23290_ (.Y(_05587_),
    .B1(_05586_),
    .B2(net540),
    .A2(net664),
    .A1(\cpu.dcache.r_data[7][4] ));
 sg13g2_nand2b_1 _23291_ (.Y(_05588_),
    .B(net613),
    .A_N(_05587_));
 sg13g2_and4_1 _23292_ (.A(net483),
    .B(_05584_),
    .C(_05585_),
    .D(_05588_),
    .X(_05589_));
 sg13g2_a21oi_2 _23293_ (.B1(_05589_),
    .Y(_05590_),
    .A2(net485),
    .A1(_00116_));
 sg13g2_nand2_1 _23294_ (.Y(_05591_),
    .A(_12041_),
    .B(_05590_));
 sg13g2_a21oi_1 _23295_ (.A1(_04858_),
    .A2(_05591_),
    .Y(_05592_),
    .B1(_04880_));
 sg13g2_a221oi_1 _23296_ (.B2(_05590_),
    .C1(_05592_),
    .B1(_05583_),
    .A1(_04877_),
    .Y(_05593_),
    .A2(_05582_));
 sg13g2_nor2_1 _23297_ (.A(net663),
    .B(_05226_),
    .Y(_05594_));
 sg13g2_nor2_1 _23298_ (.A(net983),
    .B(_05594_),
    .Y(_05595_));
 sg13g2_nor3_1 _23299_ (.A(net623),
    .B(net595),
    .C(_05219_),
    .Y(_05596_));
 sg13g2_and2_1 _23300_ (.A(net595),
    .B(_05590_),
    .X(_05597_));
 sg13g2_nor4_1 _23301_ (.A(net742),
    .B(_05595_),
    .C(_05596_),
    .D(_05597_),
    .Y(_05598_));
 sg13g2_nor3_1 _23302_ (.A(_12038_),
    .B(_05593_),
    .C(_05598_),
    .Y(_05599_));
 sg13g2_a21oi_1 _23303_ (.A1(_04834_),
    .A2(_05574_),
    .Y(_05600_),
    .B1(_05599_));
 sg13g2_nand2_1 _23304_ (.Y(_05601_),
    .A(net452),
    .B(net76));
 sg13g2_o21ai_1 _23305_ (.B1(_05601_),
    .Y(_05602_),
    .A1(net75),
    .A2(_05600_));
 sg13g2_nand2_1 _23306_ (.Y(_05603_),
    .A(net115),
    .B(_05602_));
 sg13g2_o21ai_1 _23307_ (.B1(_05603_),
    .Y(_01028_),
    .A1(_05465_),
    .A2(_05529_));
 sg13g2_nand2_1 _23308_ (.Y(_05604_),
    .A(net661),
    .B(_04613_));
 sg13g2_o21ai_1 _23309_ (.B1(_05604_),
    .Y(_05605_),
    .A1(net592),
    .A2(_04611_));
 sg13g2_and2_1 _23310_ (.A(net989),
    .B(net153),
    .X(_05606_));
 sg13g2_a21oi_1 _23311_ (.A1(_05168_),
    .A2(_05605_),
    .Y(_05607_),
    .B1(_05606_));
 sg13g2_a21o_1 _23312_ (.A2(_04894_),
    .A1(_09193_),
    .B1(net348),
    .X(_05608_));
 sg13g2_nor2_1 _23313_ (.A(net780),
    .B(_00132_),
    .Y(_05609_));
 sg13g2_a21oi_1 _23314_ (.A1(net780),
    .A2(net8),
    .Y(_05610_),
    .B1(_05609_));
 sg13g2_nand3_1 _23315_ (.B(_09195_),
    .C(net447),
    .A(_09194_),
    .Y(_05611_));
 sg13g2_o21ai_1 _23316_ (.B1(_05611_),
    .Y(_05612_),
    .A1(_12709_),
    .A2(_05610_));
 sg13g2_a221oi_1 _23317_ (.B2(\cpu.gpio.genblk2[5].srcs_io[0] ),
    .C1(_05612_),
    .B1(_10115_),
    .A1(\cpu.gpio.genblk1[5].srcs_o[0] ),
    .Y(_05613_),
    .A2(net573));
 sg13g2_nor2_1 _23318_ (.A(_00131_),
    .B(_05084_),
    .Y(_05614_));
 sg13g2_buf_2 _23319_ (.A(\cpu.gpio.r_src_io[5][1] ),
    .X(_05615_));
 sg13g2_nand2_1 _23320_ (.Y(_05616_),
    .A(net912),
    .B(_05615_));
 sg13g2_o21ai_1 _23321_ (.B1(_05616_),
    .Y(_05617_),
    .A1(net780),
    .A2(_00128_));
 sg13g2_inv_1 _23322_ (.Y(_05618_),
    .A(_00129_));
 sg13g2_a22oi_1 _23323_ (.Y(_05619_),
    .B1(_05618_),
    .B2(net1030),
    .A2(net982),
    .A1(_09195_));
 sg13g2_nor2b_1 _23324_ (.A(_05619_),
    .B_N(net487),
    .Y(_05620_));
 sg13g2_a221oi_1 _23325_ (.B2(_04914_),
    .C1(_05620_),
    .B1(_05617_),
    .A1(_09194_),
    .Y(_05621_),
    .A2(_04973_));
 sg13g2_o21ai_1 _23326_ (.B1(_05621_),
    .Y(_05622_),
    .A1(_00130_),
    .A2(_04904_));
 sg13g2_a221oi_1 _23327_ (.B2(net1030),
    .C1(_05622_),
    .B1(_05614_),
    .A1(_09193_),
    .Y(_05623_),
    .A2(_04899_));
 sg13g2_o21ai_1 _23328_ (.B1(_05623_),
    .Y(_05624_),
    .A1(_04902_),
    .A2(_05613_));
 sg13g2_a21oi_1 _23329_ (.A1(\cpu.gpio.r_enable_in[5] ),
    .A2(_05608_),
    .Y(_05625_),
    .B1(_05624_));
 sg13g2_buf_1 _23330_ (.A(\cpu.spi.r_clk_count[2][5] ),
    .X(_05626_));
 sg13g2_nor2_1 _23331_ (.A(_00127_),
    .B(_05091_),
    .Y(_05627_));
 sg13g2_a221oi_1 _23332_ (.B2(\cpu.spi.r_timeout[5] ),
    .C1(_05627_),
    .B1(_05116_),
    .A1(_05626_),
    .Y(_05628_),
    .A2(_04985_));
 sg13g2_o21ai_1 _23333_ (.B1(_05628_),
    .Y(_05629_),
    .A1(_00126_),
    .A2(_04982_));
 sg13g2_a21o_1 _23334_ (.A2(_04975_),
    .A1(_09271_),
    .B1(_05629_),
    .X(_05630_));
 sg13g2_a22oi_1 _23335_ (.Y(_05631_),
    .B1(_04996_),
    .B2(\cpu.uart.r_in[5] ),
    .A2(net406),
    .A1(\cpu.uart.r_div_value[5] ));
 sg13g2_mux2_1 _23336_ (.A0(\cpu.intr.r_timer_count[5] ),
    .A1(_09986_),
    .S(net914),
    .X(_05632_));
 sg13g2_a22oi_1 _23337_ (.Y(_05633_),
    .B1(_05632_),
    .B2(net499),
    .A2(net447),
    .A1(_09170_));
 sg13g2_buf_2 _23338_ (.A(\cpu.intr.r_clock_count[21] ),
    .X(_05634_));
 sg13g2_mux2_1 _23339_ (.A0(\cpu.intr.r_timer_reload[5] ),
    .A1(\cpu.intr.r_timer_reload[21] ),
    .S(net914),
    .X(_05635_));
 sg13g2_a22oi_1 _23340_ (.Y(_05636_),
    .B1(_05635_),
    .B2(net515),
    .A2(net417),
    .A1(_05634_));
 sg13g2_nand3_1 _23341_ (.B(\cpu.intr.r_clock_cmp[21] ),
    .C(net557),
    .A(net781),
    .Y(_05637_));
 sg13g2_a22oi_1 _23342_ (.Y(_05638_),
    .B1(net574),
    .B2(_10132_),
    .A2(net557),
    .A1(\cpu.intr.r_clock_cmp[5] ));
 sg13g2_or2_1 _23343_ (.X(_05639_),
    .B(_05638_),
    .A(net781));
 sg13g2_nand4_1 _23344_ (.B(_05636_),
    .C(_05637_),
    .A(_05633_),
    .Y(_05640_),
    .D(_05639_));
 sg13g2_a21oi_1 _23345_ (.A1(_09170_),
    .A2(net347),
    .Y(_05641_),
    .B1(net448));
 sg13g2_nor2b_1 _23346_ (.A(_05641_),
    .B_N(\cpu.intr.r_enable[5] ),
    .Y(_05642_));
 sg13g2_o21ai_1 _23347_ (.B1(_04932_),
    .Y(_05643_),
    .A1(_05640_),
    .A2(_05642_));
 sg13g2_o21ai_1 _23348_ (.B1(_05643_),
    .Y(_05644_),
    .A1(net593),
    .A2(_05631_));
 sg13g2_a21oi_1 _23349_ (.A1(_04992_),
    .A2(_05630_),
    .Y(_05645_),
    .B1(_05644_));
 sg13g2_o21ai_1 _23350_ (.B1(_05645_),
    .Y(_05646_),
    .A1(_04884_),
    .A2(_05625_));
 sg13g2_a22oi_1 _23351_ (.Y(_05647_),
    .B1(net530),
    .B2(\cpu.dcache.r_data[3][21] ),
    .A2(net556),
    .A1(\cpu.dcache.r_data[6][21] ));
 sg13g2_a22oi_1 _23352_ (.Y(_05648_),
    .B1(net484),
    .B2(\cpu.dcache.r_data[1][21] ),
    .A2(net560),
    .A1(\cpu.dcache.r_data[2][21] ));
 sg13g2_mux2_1 _23353_ (.A0(\cpu.dcache.r_data[5][21] ),
    .A1(\cpu.dcache.r_data[7][21] ),
    .S(_09296_),
    .X(_05649_));
 sg13g2_a22oi_1 _23354_ (.Y(_05650_),
    .B1(_05649_),
    .B2(net633),
    .A2(net921),
    .A1(\cpu.dcache.r_data[4][21] ));
 sg13g2_nand2b_1 _23355_ (.Y(_05651_),
    .B(net673),
    .A_N(_05650_));
 sg13g2_and4_1 _23356_ (.A(net482),
    .B(_05647_),
    .C(_05648_),
    .D(_05651_),
    .X(_05652_));
 sg13g2_a21oi_1 _23357_ (.A1(_00123_),
    .A2(net485),
    .Y(_05653_),
    .B1(_05652_));
 sg13g2_nand2_1 _23358_ (.Y(_05654_),
    .A(_09944_),
    .B(_05653_));
 sg13g2_inv_1 _23359_ (.Y(_05655_),
    .A(_00122_));
 sg13g2_a22oi_1 _23360_ (.Y(_05656_),
    .B1(net503),
    .B2(\cpu.dcache.r_data[1][5] ),
    .A2(net502),
    .A1(\cpu.dcache.r_data[2][5] ));
 sg13g2_a22oi_1 _23361_ (.Y(_05657_),
    .B1(net559),
    .B2(\cpu.dcache.r_data[3][5] ),
    .A2(net576),
    .A1(\cpu.dcache.r_data[7][5] ));
 sg13g2_mux2_1 _23362_ (.A0(\cpu.dcache.r_data[4][5] ),
    .A1(\cpu.dcache.r_data[6][5] ),
    .S(net516),
    .X(_05658_));
 sg13g2_a22oi_1 _23363_ (.Y(_05659_),
    .B1(_05658_),
    .B2(net540),
    .A2(net918),
    .A1(\cpu.dcache.r_data[5][5] ));
 sg13g2_nand2b_1 _23364_ (.Y(_05660_),
    .B(net613),
    .A_N(_05659_));
 sg13g2_nand4_1 _23365_ (.B(_05656_),
    .C(_05657_),
    .A(net483),
    .Y(_05661_),
    .D(_05660_));
 sg13g2_o21ai_1 _23366_ (.B1(_05661_),
    .Y(_05662_),
    .A1(_05655_),
    .A2(net483));
 sg13g2_mux2_1 _23367_ (.A0(_05654_),
    .A1(_05662_),
    .S(net1025),
    .X(_05663_));
 sg13g2_nor2b_1 _23368_ (.A(net1025),
    .B_N(_05250_),
    .Y(_05664_));
 sg13g2_nor3_1 _23369_ (.A(net663),
    .B(_05258_),
    .C(_05664_),
    .Y(_05665_));
 sg13g2_a21oi_1 _23370_ (.A1(net595),
    .A2(_05663_),
    .Y(_05666_),
    .B1(_05665_));
 sg13g2_nand2b_1 _23371_ (.Y(_05667_),
    .B(_05666_),
    .A_N(net742));
 sg13g2_o21ai_1 _23372_ (.B1(_05654_),
    .Y(_05668_),
    .A1(_09945_),
    .A2(_05662_));
 sg13g2_nand2_1 _23373_ (.Y(_05669_),
    .A(net662),
    .B(_05668_));
 sg13g2_a21oi_1 _23374_ (.A1(_05667_),
    .A2(_05669_),
    .Y(_05670_),
    .B1(net855));
 sg13g2_a21oi_1 _23375_ (.A1(net855),
    .A2(_05646_),
    .Y(_05671_),
    .B1(_05670_));
 sg13g2_nor2_1 _23376_ (.A(net75),
    .B(_05671_),
    .Y(_05672_));
 sg13g2_a221oi_1 _23377_ (.B2(net668),
    .C1(_05672_),
    .B1(net36),
    .A1(net803),
    .Y(_05673_),
    .A2(_11485_));
 sg13g2_a21oi_1 _23378_ (.A1(net114),
    .A2(_05607_),
    .Y(_01029_),
    .B1(_05673_));
 sg13g2_mux2_1 _23379_ (.A0(_04644_),
    .A1(_04648_),
    .S(net661),
    .X(_05674_));
 sg13g2_and2_1 _23380_ (.A(net988),
    .B(_05165_),
    .X(_05675_));
 sg13g2_a21oi_1 _23381_ (.A1(net130),
    .A2(_05674_),
    .Y(_05676_),
    .B1(_05675_));
 sg13g2_nor3_1 _23382_ (.A(net685),
    .B(_00143_),
    .C(_12709_),
    .Y(_05677_));
 sg13g2_a22oi_1 _23383_ (.Y(_05678_),
    .B1(net574),
    .B2(\cpu.gpio.genblk1[6].srcs_o[0] ),
    .A2(net557),
    .A1(net9));
 sg13g2_a21oi_1 _23384_ (.A1(_09187_),
    .A2(net447),
    .Y(_05679_),
    .B1(net487));
 sg13g2_nand2b_1 _23385_ (.Y(_05680_),
    .B(_09188_),
    .A_N(_05679_));
 sg13g2_o21ai_1 _23386_ (.B1(_05680_),
    .Y(_05681_),
    .A1(net612),
    .A2(_05678_));
 sg13g2_or2_1 _23387_ (.X(_05682_),
    .B(_05681_),
    .A(_05677_));
 sg13g2_buf_1 _23388_ (.A(\cpu.gpio.r_src_io[5][2] ),
    .X(_05683_));
 sg13g2_nand2_1 _23389_ (.Y(_05684_),
    .A(net780),
    .B(_05683_));
 sg13g2_o21ai_1 _23390_ (.B1(_05684_),
    .Y(_05685_),
    .A1(net685),
    .A2(_00139_));
 sg13g2_a22oi_1 _23391_ (.Y(_05686_),
    .B1(_05685_),
    .B2(net486),
    .A2(net348),
    .A1(\cpu.gpio.r_enable_in[6] ));
 sg13g2_inv_1 _23392_ (.Y(_05687_),
    .A(_00140_));
 sg13g2_a22oi_1 _23393_ (.Y(_05688_),
    .B1(net404),
    .B2(_09187_),
    .A2(_04909_),
    .A1(_05687_));
 sg13g2_and2_1 _23394_ (.A(net982),
    .B(_10115_),
    .X(_05689_));
 sg13g2_nand3b_1 _23395_ (.B(net447),
    .C(_11973_),
    .Y(_05690_),
    .A_N(_00142_));
 sg13g2_o21ai_1 _23396_ (.B1(_05690_),
    .Y(_05691_),
    .A1(_00141_),
    .A2(_04904_));
 sg13g2_a221oi_1 _23397_ (.B2(\cpu.gpio.genblk2[6].srcs_io[0] ),
    .C1(_05691_),
    .B1(_05689_),
    .A1(_09175_),
    .Y(_05692_),
    .A2(_04899_));
 sg13g2_nand2b_1 _23398_ (.Y(_05693_),
    .B(_04894_),
    .A_N(_09176_));
 sg13g2_nand4_1 _23399_ (.B(_05688_),
    .C(_05692_),
    .A(_05686_),
    .Y(_05694_),
    .D(_05693_));
 sg13g2_a21oi_1 _23400_ (.A1(net982),
    .A2(_05682_),
    .Y(_05695_),
    .B1(_05694_));
 sg13g2_buf_1 _23401_ (.A(\cpu.spi.r_clk_count[2][6] ),
    .X(_05696_));
 sg13g2_nor2_1 _23402_ (.A(_00138_),
    .B(_05091_),
    .Y(_05697_));
 sg13g2_a221oi_1 _23403_ (.B2(\cpu.spi.r_timeout[6] ),
    .C1(_05697_),
    .B1(_05116_),
    .A1(_05696_),
    .Y(_05698_),
    .A2(_04985_));
 sg13g2_o21ai_1 _23404_ (.B1(_05698_),
    .Y(_05699_),
    .A1(_00137_),
    .A2(_04982_));
 sg13g2_a21o_1 _23405_ (.A2(_04975_),
    .A1(_09265_),
    .B1(_05699_),
    .X(_05700_));
 sg13g2_a22oi_1 _23406_ (.Y(_05701_),
    .B1(net574),
    .B2(_10136_),
    .A2(net515),
    .A1(\cpu.intr.r_timer_reload[6] ));
 sg13g2_buf_1 _23407_ (.A(\cpu.intr.r_clock_count[22] ),
    .X(_05702_));
 sg13g2_nand3_1 _23408_ (.B(\cpu.intr.r_timer_reload[22] ),
    .C(net515),
    .A(net686),
    .Y(_05703_));
 sg13g2_mux2_1 _23409_ (.A0(\cpu.intr.r_clock_cmp[6] ),
    .A1(\cpu.intr.r_clock_cmp[22] ),
    .S(net914),
    .X(_05704_));
 sg13g2_mux2_1 _23410_ (.A0(\cpu.intr.r_timer_count[6] ),
    .A1(\cpu.intr.r_timer_count[22] ),
    .S(net914),
    .X(_05705_));
 sg13g2_a22oi_1 _23411_ (.Y(_05706_),
    .B1(_05705_),
    .B2(net499),
    .A2(_05704_),
    .A1(net557));
 sg13g2_nand2_1 _23412_ (.Y(_05707_),
    .A(_05703_),
    .B(_05706_));
 sg13g2_a21oi_1 _23413_ (.A1(_05702_),
    .A2(net417),
    .Y(_05708_),
    .B1(_05707_));
 sg13g2_o21ai_1 _23414_ (.B1(_05708_),
    .Y(_05709_),
    .A1(net623),
    .A2(_05701_));
 sg13g2_a22oi_1 _23415_ (.Y(_05710_),
    .B1(_04996_),
    .B2(\cpu.uart.r_in[6] ),
    .A2(net406),
    .A1(\cpu.uart.r_div_value[6] ));
 sg13g2_nor2_1 _23416_ (.A(net593),
    .B(_05710_),
    .Y(_05711_));
 sg13g2_a221oi_1 _23417_ (.B2(_05104_),
    .C1(_05711_),
    .B1(_05709_),
    .A1(_04992_),
    .Y(_05712_),
    .A2(_05700_));
 sg13g2_o21ai_1 _23418_ (.B1(_05712_),
    .Y(_05713_),
    .A1(_04884_),
    .A2(_05695_));
 sg13g2_inv_1 _23419_ (.Y(_05714_),
    .A(_00133_));
 sg13g2_a22oi_1 _23420_ (.Y(_05715_),
    .B1(net484),
    .B2(\cpu.dcache.r_data[1][6] ),
    .A2(net560),
    .A1(\cpu.dcache.r_data[2][6] ));
 sg13g2_a22oi_1 _23421_ (.Y(_05716_),
    .B1(net530),
    .B2(\cpu.dcache.r_data[3][6] ),
    .A2(net576),
    .A1(\cpu.dcache.r_data[7][6] ));
 sg13g2_mux2_1 _23422_ (.A0(\cpu.dcache.r_data[4][6] ),
    .A1(\cpu.dcache.r_data[6][6] ),
    .S(net578),
    .X(_05717_));
 sg13g2_a22oi_1 _23423_ (.Y(_05718_),
    .B1(_05717_),
    .B2(net600),
    .A2(net918),
    .A1(\cpu.dcache.r_data[5][6] ));
 sg13g2_nand2b_1 _23424_ (.Y(_05719_),
    .B(net673),
    .A_N(_05718_));
 sg13g2_nand4_1 _23425_ (.B(_05715_),
    .C(_05716_),
    .A(net482),
    .Y(_05720_),
    .D(_05719_));
 sg13g2_o21ai_1 _23426_ (.B1(_05720_),
    .Y(_05721_),
    .A1(_05714_),
    .A2(net483));
 sg13g2_a22oi_1 _23427_ (.Y(_05722_),
    .B1(net562),
    .B2(\cpu.dcache.r_data[1][22] ),
    .A2(net610),
    .A1(\cpu.dcache.r_data[2][22] ));
 sg13g2_a22oi_1 _23428_ (.Y(_05723_),
    .B1(net609),
    .B2(\cpu.dcache.r_data[3][22] ),
    .A2(net576),
    .A1(\cpu.dcache.r_data[7][22] ));
 sg13g2_mux2_1 _23429_ (.A0(\cpu.dcache.r_data[4][22] ),
    .A1(\cpu.dcache.r_data[6][22] ),
    .S(_09295_),
    .X(_05724_));
 sg13g2_a22oi_1 _23430_ (.Y(_05725_),
    .B1(_05724_),
    .B2(net600),
    .A2(net918),
    .A1(\cpu.dcache.r_data[5][22] ));
 sg13g2_nand2b_1 _23431_ (.Y(_05726_),
    .B(net673),
    .A_N(_05725_));
 sg13g2_and4_1 _23432_ (.A(net533),
    .B(_05722_),
    .C(_05723_),
    .D(_05726_),
    .X(_05727_));
 sg13g2_a21oi_1 _23433_ (.A1(_00134_),
    .A2(net594),
    .Y(_05728_),
    .B1(_05727_));
 sg13g2_nand2_1 _23434_ (.Y(_05729_),
    .A(_09943_),
    .B(_05728_));
 sg13g2_o21ai_1 _23435_ (.B1(_05729_),
    .Y(_05730_),
    .A1(_09945_),
    .A2(_05721_));
 sg13g2_o21ai_1 _23436_ (.B1(_05285_),
    .Y(_05731_),
    .A1(_12041_),
    .A2(_05277_));
 sg13g2_mux2_1 _23437_ (.A0(_05729_),
    .A1(_05721_),
    .S(_12040_),
    .X(_05732_));
 sg13g2_nand2_1 _23438_ (.Y(_05733_),
    .A(net663),
    .B(_05732_));
 sg13g2_o21ai_1 _23439_ (.B1(_05733_),
    .Y(_05734_),
    .A1(net663),
    .A2(_05731_));
 sg13g2_nor2_1 _23440_ (.A(net742),
    .B(_05734_),
    .Y(_05735_));
 sg13g2_a21oi_1 _23441_ (.A1(net742),
    .A2(_05730_),
    .Y(_05736_),
    .B1(_05735_));
 sg13g2_nor2_1 _23442_ (.A(_12038_),
    .B(_05736_),
    .Y(_05737_));
 sg13g2_a21oi_1 _23443_ (.A1(net855),
    .A2(_05713_),
    .Y(_05738_),
    .B1(_05737_));
 sg13g2_nand2_1 _23444_ (.Y(_05739_),
    .A(net1000),
    .B(net76));
 sg13g2_o21ai_1 _23445_ (.B1(_05739_),
    .Y(_05740_),
    .A1(net75),
    .A2(_05738_));
 sg13g2_nand2_1 _23446_ (.Y(_05741_),
    .A(net115),
    .B(_05740_));
 sg13g2_o21ai_1 _23447_ (.B1(_05741_),
    .Y(_01030_),
    .A1(_05465_),
    .A2(_05676_));
 sg13g2_and2_1 _23448_ (.A(_05161_),
    .B(_04677_),
    .X(_05742_));
 sg13g2_a21oi_1 _23449_ (.A1(net529),
    .A2(_04673_),
    .Y(_05743_),
    .B1(_05742_));
 sg13g2_nor2_1 _23450_ (.A(net987),
    .B(net152),
    .Y(_05744_));
 sg13g2_a21oi_1 _23451_ (.A1(net130),
    .A2(_05743_),
    .Y(_05745_),
    .B1(_05744_));
 sg13g2_nand2_1 _23452_ (.Y(_05746_),
    .A(_09222_),
    .B(_05007_));
 sg13g2_o21ai_1 _23453_ (.B1(_05746_),
    .Y(_05747_),
    .A1(net36),
    .A2(_05125_));
 sg13g2_mux2_1 _23454_ (.A0(_05745_),
    .A1(_05747_),
    .S(net115),
    .X(_01031_));
 sg13g2_nor2_1 _23455_ (.A(net529),
    .B(_04707_),
    .Y(_05748_));
 sg13g2_a21o_1 _23456_ (.A2(_04706_),
    .A1(net529),
    .B1(_05748_),
    .X(_05749_));
 sg13g2_a22oi_1 _23457_ (.Y(_05750_),
    .B1(net449),
    .B2(\cpu.intr.r_timer_reload[8] ),
    .A2(net514),
    .A1(_10147_));
 sg13g2_a22oi_1 _23458_ (.Y(_05751_),
    .B1(net405),
    .B2(\cpu.intr.r_clock_cmp[8] ),
    .A2(net407),
    .A1(\cpu.intr.r_clock_cmp[24] ));
 sg13g2_buf_1 _23459_ (.A(\cpu.intr.r_clock_count[24] ),
    .X(_05752_));
 sg13g2_a22oi_1 _23460_ (.Y(_05753_),
    .B1(net446),
    .B2(_09962_),
    .A2(net362),
    .A1(_05752_));
 sg13g2_nand3_1 _23461_ (.B(_05751_),
    .C(_05753_),
    .A(_05750_),
    .Y(_05754_));
 sg13g2_a21o_1 _23462_ (.A2(_04873_),
    .A1(_04877_),
    .B1(_04867_),
    .X(_05755_));
 sg13g2_a221oi_1 _23463_ (.B2(_04881_),
    .C1(net981),
    .B1(_05755_),
    .A1(_05149_),
    .Y(_05756_),
    .A2(_05754_));
 sg13g2_nor3_1 _23464_ (.A(net76),
    .B(_05127_),
    .C(_05756_),
    .Y(_05757_));
 sg13g2_a21oi_1 _23465_ (.A1(_09221_),
    .A2(_03691_),
    .Y(_05758_),
    .B1(_05757_));
 sg13g2_nor3_1 _23466_ (.A(\cpu.ex.pc[8] ),
    .B(net130),
    .C(net121),
    .Y(_05759_));
 sg13g2_a221oi_1 _23467_ (.B2(net115),
    .C1(_05759_),
    .B1(_05758_),
    .A1(_05166_),
    .Y(_01032_),
    .A2(_05749_));
 sg13g2_a21o_1 _23468_ (.A2(_04742_),
    .A1(_05162_),
    .B1(_05165_),
    .X(_05760_));
 sg13g2_a21oi_1 _23469_ (.A1(_05172_),
    .A2(_04739_),
    .Y(_05761_),
    .B1(_05760_));
 sg13g2_o21ai_1 _23470_ (.B1(_11487_),
    .Y(_05762_),
    .A1(net986),
    .A2(net130));
 sg13g2_a21oi_1 _23471_ (.A1(net1074),
    .A2(_11491_),
    .Y(_05763_),
    .B1(net869));
 sg13g2_a21o_1 _23472_ (.A2(_05347_),
    .A1(net532),
    .B1(_05340_),
    .X(_05764_));
 sg13g2_a22oi_1 _23473_ (.Y(_05765_),
    .B1(net446),
    .B2(\cpu.intr.r_timer_count[9] ),
    .A2(net514),
    .A1(_10153_));
 sg13g2_a22oi_1 _23474_ (.Y(_05766_),
    .B1(net449),
    .B2(\cpu.intr.r_timer_reload[9] ),
    .A2(net407),
    .A1(\cpu.intr.r_clock_cmp[25] ));
 sg13g2_buf_2 _23475_ (.A(\cpu.intr.r_clock_count[25] ),
    .X(_05767_));
 sg13g2_a22oi_1 _23476_ (.Y(_05768_),
    .B1(net405),
    .B2(\cpu.intr.r_clock_cmp[9] ),
    .A2(net362),
    .A1(_05767_));
 sg13g2_nand3_1 _23477_ (.B(_05766_),
    .C(_05768_),
    .A(_05765_),
    .Y(_05769_));
 sg13g2_a221oi_1 _23478_ (.B2(_05149_),
    .C1(net981),
    .B1(_05769_),
    .A1(_04881_),
    .Y(_05770_),
    .A2(_05764_));
 sg13g2_nor3_1 _23479_ (.A(net76),
    .B(_05127_),
    .C(_05770_),
    .Y(_05771_));
 sg13g2_buf_1 _23480_ (.A(net141),
    .X(_05772_));
 sg13g2_o21ai_1 _23481_ (.B1(_05772_),
    .Y(_05773_),
    .A1(_05763_),
    .A2(_05771_));
 sg13g2_o21ai_1 _23482_ (.B1(_05773_),
    .Y(_01033_),
    .A1(_05761_),
    .A2(_05762_));
 sg13g2_o21ai_1 _23483_ (.B1(net130),
    .Y(_05774_),
    .A1(_03448_),
    .A2(_03343_));
 sg13g2_mux2_1 _23484_ (.A0(net1124),
    .A1(_05774_),
    .S(_05038_),
    .X(_01034_));
 sg13g2_nand2b_1 _23485_ (.Y(_05775_),
    .B(\cpu.dec.r_rd[1] ),
    .A_N(_03448_));
 sg13g2_a21oi_1 _23486_ (.A1(net130),
    .A2(_05775_),
    .Y(_05776_),
    .B1(net121));
 sg13g2_a21o_1 _23487_ (.A2(_05039_),
    .A1(net1125),
    .B1(_05776_),
    .X(_01035_));
 sg13g2_nor4_2 _23488_ (.A(_03448_),
    .B(_09317_),
    .C(net153),
    .Y(_05777_),
    .D(net141));
 sg13g2_a22oi_1 _23489_ (.Y(_05778_),
    .B1(_05777_),
    .B2(\cpu.dec.r_rd[2] ),
    .A2(_05772_),
    .A1(net1052));
 sg13g2_inv_1 _23490_ (.Y(_01036_),
    .A(_05778_));
 sg13g2_a22oi_1 _23491_ (.Y(_05779_),
    .B1(_05777_),
    .B2(\cpu.dec.r_rd[3] ),
    .A2(net113),
    .A1(net1126));
 sg13g2_inv_1 _23492_ (.Y(_01037_),
    .A(_05779_));
 sg13g2_mux2_1 _23493_ (.A0(\cpu.dec.r_swapsp ),
    .A1(\cpu.ex.r_wb_swapsp ),
    .S(_05039_),
    .X(_01038_));
 sg13g2_nand2_2 _23494_ (.Y(_05780_),
    .A(_10670_),
    .B(_10671_));
 sg13g2_mux2_1 _23495_ (.A0(net913),
    .A1(_05780_),
    .S(net116),
    .X(_01039_));
 sg13g2_buf_1 _23496_ (.A(net981),
    .X(_05781_));
 sg13g2_a221oi_1 _23497_ (.B2(_10418_),
    .C1(_05156_),
    .B1(net513),
    .A1(_10392_),
    .Y(_05782_),
    .A2(net512));
 sg13g2_a21o_1 _23498_ (.A2(_03712_),
    .A1(net854),
    .B1(_05782_),
    .X(_05783_));
 sg13g2_nand2_1 _23499_ (.Y(_05784_),
    .A(\cpu.dcache.wdata[10] ),
    .B(net115));
 sg13g2_o21ai_1 _23500_ (.B1(_05784_),
    .Y(_01040_),
    .A1(net104),
    .A2(_05783_));
 sg13g2_nor2_1 _23501_ (.A(net572),
    .B(_10608_),
    .Y(_05785_));
 sg13g2_a21oi_1 _23502_ (.A1(_09298_),
    .A2(net512),
    .Y(_05786_),
    .B1(_05785_));
 sg13g2_nor2_1 _23503_ (.A(_09213_),
    .B(_05786_),
    .Y(_05787_));
 sg13g2_a21oi_1 _23504_ (.A1(_09213_),
    .A2(_10381_),
    .Y(_05788_),
    .B1(_05787_));
 sg13g2_nand2_1 _23505_ (.Y(_05789_),
    .A(_10162_),
    .B(net113));
 sg13g2_o21ai_1 _23506_ (.B1(_05789_),
    .Y(_01041_),
    .A1(net104),
    .A2(_05788_));
 sg13g2_a21oi_1 _23507_ (.A1(_10775_),
    .A2(_10787_),
    .Y(_05790_),
    .B1(_10229_));
 sg13g2_a21o_1 _23508_ (.A2(net512),
    .A1(_03513_),
    .B1(_05790_),
    .X(_05791_));
 sg13g2_a21oi_1 _23509_ (.A1(_10340_),
    .A2(_10343_),
    .Y(_05792_),
    .B1(_05781_));
 sg13g2_a21oi_1 _23510_ (.A1(net854),
    .A2(_05791_),
    .Y(_05793_),
    .B1(_05792_));
 sg13g2_nand2_1 _23511_ (.Y(_05794_),
    .A(\cpu.dcache.wdata[12] ),
    .B(net113));
 sg13g2_o21ai_1 _23512_ (.B1(_05794_),
    .Y(_01042_),
    .A1(net104),
    .A2(_05793_));
 sg13g2_nor2_2 _23513_ (.A(_10762_),
    .B(_10763_),
    .Y(_05795_));
 sg13g2_mux2_1 _23514_ (.A0(_10288_),
    .A1(_05795_),
    .S(net981),
    .X(_05796_));
 sg13g2_nand2_1 _23515_ (.Y(_05797_),
    .A(net116),
    .B(_05796_));
 sg13g2_o21ai_1 _23516_ (.B1(_05797_),
    .Y(_01043_),
    .A1(_12101_),
    .A2(net114));
 sg13g2_a21o_1 _23517_ (.A2(_10699_),
    .A1(net513),
    .B1(_10701_),
    .X(_05798_));
 sg13g2_nand2_1 _23518_ (.Y(_05799_),
    .A(net981),
    .B(_05798_));
 sg13g2_o21ai_1 _23519_ (.B1(_05799_),
    .Y(_05800_),
    .A1(net854),
    .A2(_10481_));
 sg13g2_nand2_1 _23520_ (.Y(_05801_),
    .A(net116),
    .B(_05800_));
 sg13g2_o21ai_1 _23521_ (.B1(_05801_),
    .Y(_01044_),
    .A1(_12107_),
    .A2(net114));
 sg13g2_nand2_1 _23522_ (.Y(_05802_),
    .A(net1138),
    .B(net512));
 sg13g2_nand2_1 _23523_ (.Y(_05803_),
    .A(_10731_),
    .B(_05802_));
 sg13g2_nor2_1 _23524_ (.A(net854),
    .B(_10450_),
    .Y(_05804_));
 sg13g2_a21oi_1 _23525_ (.A1(net854),
    .A2(_05803_),
    .Y(_05805_),
    .B1(_05804_));
 sg13g2_nand2_1 _23526_ (.Y(_05806_),
    .A(\cpu.dcache.wdata[15] ),
    .B(net113));
 sg13g2_o21ai_1 _23527_ (.B1(_05806_),
    .Y(_01045_),
    .A1(net104),
    .A2(_05805_));
 sg13g2_buf_1 _23528_ (.A(net1061),
    .X(_05807_));
 sg13g2_mux2_1 _23529_ (.A0(_05807_),
    .A1(_10642_),
    .S(net116),
    .X(_01046_));
 sg13g2_nand2_1 _23530_ (.Y(_05808_),
    .A(_10107_),
    .B(net113));
 sg13g2_o21ai_1 _23531_ (.B1(_05808_),
    .Y(_01047_),
    .A1(_03712_),
    .A2(net104));
 sg13g2_nand2_1 _23532_ (.Y(_05809_),
    .A(_10121_),
    .B(net113));
 sg13g2_o21ai_1 _23533_ (.B1(_05809_),
    .Y(_01048_),
    .A1(_05786_),
    .A2(net104));
 sg13g2_nand2_1 _23534_ (.Y(_05810_),
    .A(net116),
    .B(_05791_));
 sg13g2_o21ai_1 _23535_ (.B1(_05810_),
    .Y(_01049_),
    .A1(_12761_),
    .A2(net114));
 sg13g2_nand2_1 _23536_ (.Y(_05811_),
    .A(_05795_),
    .B(net116));
 sg13g2_o21ai_1 _23537_ (.B1(_05811_),
    .Y(_01050_),
    .A1(_12766_),
    .A2(net114));
 sg13g2_nand2_1 _23538_ (.Y(_05812_),
    .A(net116),
    .B(_05798_));
 sg13g2_o21ai_1 _23539_ (.B1(_05812_),
    .Y(_01051_),
    .A1(net875),
    .A2(net114));
 sg13g2_mux2_1 _23540_ (.A0(net1056),
    .A1(_05803_),
    .S(net116),
    .X(_01052_));
 sg13g2_nand2_1 _23541_ (.Y(_05813_),
    .A(net1139),
    .B(net512));
 sg13g2_a21oi_1 _23542_ (.A1(_10516_),
    .A2(_05813_),
    .Y(_05814_),
    .B1(_05781_));
 sg13g2_a21oi_1 _23543_ (.A1(net854),
    .A2(_05780_),
    .Y(_05815_),
    .B1(_05814_));
 sg13g2_nand2_1 _23544_ (.Y(_05816_),
    .A(_10146_),
    .B(net113));
 sg13g2_o21ai_1 _23545_ (.B1(_05816_),
    .Y(_01053_),
    .A1(net104),
    .A2(_05815_));
 sg13g2_a22oi_1 _23546_ (.Y(_05817_),
    .B1(net513),
    .B2(_10544_),
    .A2(net512),
    .A1(_10524_));
 sg13g2_nor2_1 _23547_ (.A(net854),
    .B(_05817_),
    .Y(_05818_));
 sg13g2_a21oi_1 _23548_ (.A1(net854),
    .A2(_10642_),
    .Y(_05819_),
    .B1(_05818_));
 sg13g2_nand2_1 _23549_ (.Y(_05820_),
    .A(\cpu.dcache.wdata[9] ),
    .B(net113));
 sg13g2_o21ai_1 _23550_ (.B1(_05820_),
    .Y(_01054_),
    .A1(net115),
    .A2(_05819_));
 sg13g2_nor2_2 _23551_ (.A(_08413_),
    .B(_08419_),
    .Y(_05821_));
 sg13g2_mux2_1 _23552_ (.A0(_08550_),
    .A1(net617),
    .S(_05821_),
    .X(_05822_));
 sg13g2_inv_1 _23553_ (.Y(_05823_),
    .A(_05822_));
 sg13g2_or3_1 _23554_ (.A(_10651_),
    .B(_10583_),
    .C(_10613_),
    .X(_05824_));
 sg13g2_o21ai_1 _23555_ (.B1(_03328_),
    .Y(_05825_),
    .A1(_10645_),
    .A2(_05824_));
 sg13g2_buf_1 _23556_ (.A(_05825_),
    .X(_05826_));
 sg13g2_buf_1 _23557_ (.A(_05826_),
    .X(_05827_));
 sg13g2_nor4_2 _23558_ (.A(_08348_),
    .B(_04778_),
    .C(_10194_),
    .Y(_05828_),
    .D(_03526_));
 sg13g2_nand2_2 _23559_ (.Y(_05829_),
    .A(net660),
    .B(_05828_));
 sg13g2_buf_2 _23560_ (.A(_00272_),
    .X(_05830_));
 sg13g2_inv_2 _23561_ (.Y(_05831_),
    .A(_05830_));
 sg13g2_nor2_1 _23562_ (.A(net993),
    .B(net617),
    .Y(_05832_));
 sg13g2_a21oi_1 _23563_ (.A1(net993),
    .A2(_05831_),
    .Y(_05833_),
    .B1(_05832_));
 sg13g2_nor3_1 _23564_ (.A(net371),
    .B(_05829_),
    .C(_05833_),
    .Y(_05834_));
 sg13g2_a21o_1 _23565_ (.A2(_05823_),
    .A1(net270),
    .B1(_05834_),
    .X(_05835_));
 sg13g2_and2_1 _23566_ (.A(net660),
    .B(_05828_),
    .X(_05836_));
 sg13g2_o21ai_1 _23567_ (.B1(_09156_),
    .Y(_05837_),
    .A1(net371),
    .A2(_05836_));
 sg13g2_buf_1 _23568_ (.A(_05837_),
    .X(_05838_));
 sg13g2_buf_1 _23569_ (.A(_10313_),
    .X(_05839_));
 sg13g2_inv_2 _23570_ (.Y(_05840_),
    .A(_05839_));
 sg13g2_a22oi_1 _23571_ (.Y(_01057_),
    .B1(_05838_),
    .B2(_05840_),
    .A2(_05835_),
    .A1(_09159_));
 sg13g2_buf_1 _23572_ (.A(_10266_),
    .X(_05841_));
 sg13g2_inv_2 _23573_ (.Y(_05842_),
    .A(net979));
 sg13g2_nor2_1 _23574_ (.A(_05840_),
    .B(_05842_),
    .Y(_05843_));
 sg13g2_buf_2 _23575_ (.A(_05843_),
    .X(_05844_));
 sg13g2_nor2_1 _23576_ (.A(net980),
    .B(net979),
    .Y(_05845_));
 sg13g2_o21ai_1 _23577_ (.B1(net993),
    .Y(_05846_),
    .A1(_05844_),
    .A2(_05845_));
 sg13g2_o21ai_1 _23578_ (.B1(_05846_),
    .Y(_05847_),
    .A1(net993),
    .A2(net577));
 sg13g2_nor2_1 _23579_ (.A(_05829_),
    .B(_05847_),
    .Y(_05848_));
 sg13g2_mux2_1 _23580_ (.A0(_08474_),
    .A1(net577),
    .S(_05821_),
    .X(_05849_));
 sg13g2_mux2_1 _23581_ (.A0(_05848_),
    .A1(_05849_),
    .S(net270),
    .X(_05850_));
 sg13g2_a22oi_1 _23582_ (.Y(_05851_),
    .B1(_05850_),
    .B2(net708),
    .A2(_05838_),
    .A1(_05841_));
 sg13g2_inv_1 _23583_ (.Y(_01058_),
    .A(_05851_));
 sg13g2_inv_1 _23584_ (.Y(_05852_),
    .A(_10474_));
 sg13g2_nand2_1 _23585_ (.Y(_05853_),
    .A(net688),
    .B(_05821_));
 sg13g2_o21ai_1 _23586_ (.B1(_05853_),
    .Y(_05854_),
    .A1(_08840_),
    .A2(_05821_));
 sg13g2_inv_1 _23587_ (.Y(_05855_),
    .A(_05854_));
 sg13g2_nand2_1 _23588_ (.Y(_05856_),
    .A(_05839_),
    .B(_05841_));
 sg13g2_buf_2 _23589_ (.A(_05856_),
    .X(_05857_));
 sg13g2_xnor2_1 _23590_ (.Y(_05858_),
    .A(net978),
    .B(_05857_));
 sg13g2_nor2_1 _23591_ (.A(net993),
    .B(net688),
    .Y(_05859_));
 sg13g2_a21oi_1 _23592_ (.A1(net993),
    .A2(_05858_),
    .Y(_05860_),
    .B1(_05859_));
 sg13g2_nor3_1 _23593_ (.A(net270),
    .B(_05829_),
    .C(_05860_),
    .Y(_05861_));
 sg13g2_a21o_1 _23594_ (.A2(_05855_),
    .A1(net270),
    .B1(_05861_),
    .X(_05862_));
 sg13g2_buf_1 _23595_ (.A(net708),
    .X(_05863_));
 sg13g2_a22oi_1 _23596_ (.Y(_01059_),
    .B1(_05862_),
    .B2(_05863_),
    .A2(_05838_),
    .A1(net978));
 sg13g2_nor2_1 _23597_ (.A(net993),
    .B(net860),
    .Y(_05864_));
 sg13g2_buf_1 _23598_ (.A(_10443_),
    .X(_05865_));
 sg13g2_buf_1 _23599_ (.A(_10474_),
    .X(_05866_));
 sg13g2_nand2_1 _23600_ (.Y(_05867_),
    .A(_05866_),
    .B(_05844_));
 sg13g2_buf_2 _23601_ (.A(_05867_),
    .X(_05868_));
 sg13g2_nor2_1 _23602_ (.A(_05865_),
    .B(_05868_),
    .Y(_05869_));
 sg13g2_buf_1 _23603_ (.A(net976),
    .X(_05870_));
 sg13g2_a21oi_1 _23604_ (.A1(net852),
    .A2(_05844_),
    .Y(_05871_),
    .B1(net1044));
 sg13g2_nor3_1 _23605_ (.A(_11056_),
    .B(_05869_),
    .C(_05871_),
    .Y(_05872_));
 sg13g2_o21ai_1 _23606_ (.B1(_05836_),
    .Y(_05873_),
    .A1(_05864_),
    .A2(_05872_));
 sg13g2_a21o_1 _23607_ (.A2(_05821_),
    .A1(net860),
    .B1(_08419_),
    .X(_05874_));
 sg13g2_mux2_1 _23608_ (.A0(_05873_),
    .A1(_05874_),
    .S(net270),
    .X(_05875_));
 sg13g2_nor2_1 _23609_ (.A(_09318_),
    .B(_05875_),
    .Y(_05876_));
 sg13g2_a21oi_1 _23610_ (.A1(_10444_),
    .A2(_05838_),
    .Y(_01060_),
    .B1(_05876_));
 sg13g2_buf_2 _23611_ (.A(_00178_),
    .X(_05877_));
 sg13g2_nor2_1 _23612_ (.A(net1121),
    .B(net977),
    .Y(_05878_));
 sg13g2_buf_1 _23613_ (.A(_05878_),
    .X(_05879_));
 sg13g2_nand2_1 _23614_ (.Y(_05880_),
    .A(_05877_),
    .B(_05879_));
 sg13g2_nand3b_1 _23615_ (.B(_05828_),
    .C(net1145),
    .Y(_05881_),
    .A_N(_10604_));
 sg13g2_buf_1 _23616_ (.A(_05881_),
    .X(_05882_));
 sg13g2_nand3b_1 _23617_ (.B(_05842_),
    .C(_05840_),
    .Y(_05883_),
    .A_N(_05882_));
 sg13g2_buf_1 _23618_ (.A(_05883_),
    .X(_05884_));
 sg13g2_nor2_1 _23619_ (.A(_05880_),
    .B(_05884_),
    .Y(_05885_));
 sg13g2_buf_1 _23620_ (.A(_05885_),
    .X(_05886_));
 sg13g2_buf_1 _23621_ (.A(_05886_),
    .X(_05887_));
 sg13g2_mux2_1 _23622_ (.A0(\cpu.genblk1.mmu.r_vtop_d[0][0] ),
    .A1(_03519_),
    .S(_05887_),
    .X(_01128_));
 sg13g2_mux2_1 _23623_ (.A0(\cpu.genblk1.mmu.r_vtop_d[0][10] ),
    .A1(net538),
    .S(net269),
    .X(_01129_));
 sg13g2_buf_1 _23624_ (.A(net860),
    .X(_05888_));
 sg13g2_mux2_1 _23625_ (.A0(\cpu.genblk1.mmu.r_vtop_d[0][11] ),
    .A1(net741),
    .S(net269),
    .X(_01130_));
 sg13g2_mux2_1 _23626_ (.A0(\cpu.genblk1.mmu.r_vtop_d[0][1] ),
    .A1(net667),
    .S(_05887_),
    .X(_01131_));
 sg13g2_mux2_1 _23627_ (.A0(\cpu.genblk1.mmu.r_vtop_d[0][2] ),
    .A1(net743),
    .S(net269),
    .X(_01132_));
 sg13g2_mux2_1 _23628_ (.A0(\cpu.genblk1.mmu.r_vtop_d[0][3] ),
    .A1(net992),
    .S(net269),
    .X(_01133_));
 sg13g2_mux2_1 _23629_ (.A0(\cpu.genblk1.mmu.r_vtop_d[0][4] ),
    .A1(net857),
    .S(net269),
    .X(_01134_));
 sg13g2_mux2_1 _23630_ (.A0(\cpu.genblk1.mmu.r_vtop_d[0][5] ),
    .A1(net859),
    .S(net269),
    .X(_01135_));
 sg13g2_mux2_1 _23631_ (.A0(\cpu.genblk1.mmu.r_vtop_d[0][6] ),
    .A1(net858),
    .S(net269),
    .X(_01136_));
 sg13g2_mux2_1 _23632_ (.A0(\cpu.genblk1.mmu.r_vtop_d[0][7] ),
    .A1(net984),
    .S(net269),
    .X(_01137_));
 sg13g2_mux2_1 _23633_ (.A0(\cpu.genblk1.mmu.r_vtop_d[0][8] ),
    .A1(net542),
    .S(_05886_),
    .X(_01138_));
 sg13g2_mux2_1 _23634_ (.A0(\cpu.genblk1.mmu.r_vtop_d[0][9] ),
    .A1(net489),
    .S(_05886_),
    .X(_01139_));
 sg13g2_buf_1 _23635_ (.A(net452),
    .X(_05889_));
 sg13g2_buf_1 _23636_ (.A(_05882_),
    .X(_05890_));
 sg13g2_nand2_1 _23637_ (.Y(_05891_),
    .A(_05840_),
    .B(net979));
 sg13g2_buf_1 _23638_ (.A(_05891_),
    .X(_05892_));
 sg13g2_nand2b_1 _23639_ (.Y(_05893_),
    .B(_10443_),
    .A_N(net1121));
 sg13g2_buf_2 _23640_ (.A(_05893_),
    .X(_05894_));
 sg13g2_nor3_2 _23641_ (.A(_05870_),
    .B(_05892_),
    .C(_05894_),
    .Y(_05895_));
 sg13g2_nor2b_1 _23642_ (.A(net481),
    .B_N(_05895_),
    .Y(_05896_));
 sg13g2_buf_1 _23643_ (.A(_05896_),
    .X(_05897_));
 sg13g2_buf_1 _23644_ (.A(_05897_),
    .X(_05898_));
 sg13g2_mux2_1 _23645_ (.A0(\cpu.genblk1.mmu.r_vtop_d[10][0] ),
    .A1(net403),
    .S(net346),
    .X(_01140_));
 sg13g2_mux2_1 _23646_ (.A0(\cpu.genblk1.mmu.r_vtop_d[10][10] ),
    .A1(_04783_),
    .S(net346),
    .X(_01141_));
 sg13g2_mux2_1 _23647_ (.A0(\cpu.genblk1.mmu.r_vtop_d[10][11] ),
    .A1(_05888_),
    .S(net346),
    .X(_01142_));
 sg13g2_mux2_1 _23648_ (.A0(\cpu.genblk1.mmu.r_vtop_d[10][1] ),
    .A1(net667),
    .S(net346),
    .X(_01143_));
 sg13g2_mux2_1 _23649_ (.A0(\cpu.genblk1.mmu.r_vtop_d[10][2] ),
    .A1(net743),
    .S(_05898_),
    .X(_01144_));
 sg13g2_mux2_1 _23650_ (.A0(\cpu.genblk1.mmu.r_vtop_d[10][3] ),
    .A1(net992),
    .S(net346),
    .X(_01145_));
 sg13g2_mux2_1 _23651_ (.A0(\cpu.genblk1.mmu.r_vtop_d[10][4] ),
    .A1(net857),
    .S(net346),
    .X(_01146_));
 sg13g2_mux2_1 _23652_ (.A0(\cpu.genblk1.mmu.r_vtop_d[10][5] ),
    .A1(net859),
    .S(_05898_),
    .X(_01147_));
 sg13g2_mux2_1 _23653_ (.A0(\cpu.genblk1.mmu.r_vtop_d[10][6] ),
    .A1(net858),
    .S(net346),
    .X(_01148_));
 sg13g2_mux2_1 _23654_ (.A0(\cpu.genblk1.mmu.r_vtop_d[10][7] ),
    .A1(net984),
    .S(net346),
    .X(_01149_));
 sg13g2_mux2_1 _23655_ (.A0(\cpu.genblk1.mmu.r_vtop_d[10][8] ),
    .A1(net542),
    .S(_05897_),
    .X(_01150_));
 sg13g2_mux2_1 _23656_ (.A0(\cpu.genblk1.mmu.r_vtop_d[10][9] ),
    .A1(net489),
    .S(_05897_),
    .X(_01151_));
 sg13g2_nor3_1 _23657_ (.A(net976),
    .B(_05857_),
    .C(_05894_),
    .Y(_05899_));
 sg13g2_buf_2 _23658_ (.A(_05899_),
    .X(_05900_));
 sg13g2_nor2b_1 _23659_ (.A(net481),
    .B_N(_05900_),
    .Y(_05901_));
 sg13g2_buf_1 _23660_ (.A(_05901_),
    .X(_05902_));
 sg13g2_buf_1 _23661_ (.A(_05902_),
    .X(_05903_));
 sg13g2_mux2_1 _23662_ (.A0(\cpu.genblk1.mmu.r_vtop_d[11][0] ),
    .A1(net403),
    .S(net345),
    .X(_01152_));
 sg13g2_mux2_1 _23663_ (.A0(\cpu.genblk1.mmu.r_vtop_d[11][10] ),
    .A1(net538),
    .S(net345),
    .X(_01153_));
 sg13g2_mux2_1 _23664_ (.A0(\cpu.genblk1.mmu.r_vtop_d[11][11] ),
    .A1(_05888_),
    .S(net345),
    .X(_01154_));
 sg13g2_mux2_1 _23665_ (.A0(\cpu.genblk1.mmu.r_vtop_d[11][1] ),
    .A1(net667),
    .S(net345),
    .X(_01155_));
 sg13g2_mux2_1 _23666_ (.A0(\cpu.genblk1.mmu.r_vtop_d[11][2] ),
    .A1(net743),
    .S(_05903_),
    .X(_01156_));
 sg13g2_mux2_1 _23667_ (.A0(\cpu.genblk1.mmu.r_vtop_d[11][3] ),
    .A1(net992),
    .S(net345),
    .X(_01157_));
 sg13g2_mux2_1 _23668_ (.A0(\cpu.genblk1.mmu.r_vtop_d[11][4] ),
    .A1(net857),
    .S(net345),
    .X(_01158_));
 sg13g2_mux2_1 _23669_ (.A0(\cpu.genblk1.mmu.r_vtop_d[11][5] ),
    .A1(_03534_),
    .S(_05903_),
    .X(_01159_));
 sg13g2_mux2_1 _23670_ (.A0(\cpu.genblk1.mmu.r_vtop_d[11][6] ),
    .A1(net858),
    .S(net345),
    .X(_01160_));
 sg13g2_mux2_1 _23671_ (.A0(\cpu.genblk1.mmu.r_vtop_d[11][7] ),
    .A1(net984),
    .S(net345),
    .X(_01161_));
 sg13g2_mux2_1 _23672_ (.A0(\cpu.genblk1.mmu.r_vtop_d[11][8] ),
    .A1(net542),
    .S(_05902_),
    .X(_01162_));
 sg13g2_mux2_1 _23673_ (.A0(\cpu.genblk1.mmu.r_vtop_d[11][9] ),
    .A1(net489),
    .S(_05902_),
    .X(_01163_));
 sg13g2_or2_1 _23674_ (.X(_05904_),
    .B(_05894_),
    .A(_05877_));
 sg13g2_buf_1 _23675_ (.A(_05904_),
    .X(_05905_));
 sg13g2_nor2_1 _23676_ (.A(_05884_),
    .B(_05905_),
    .Y(_05906_));
 sg13g2_buf_1 _23677_ (.A(_05906_),
    .X(_05907_));
 sg13g2_buf_1 _23678_ (.A(_05907_),
    .X(_05908_));
 sg13g2_mux2_1 _23679_ (.A0(\cpu.genblk1.mmu.r_vtop_d[12][0] ),
    .A1(net403),
    .S(net268),
    .X(_01164_));
 sg13g2_mux2_1 _23680_ (.A0(\cpu.genblk1.mmu.r_vtop_d[12][10] ),
    .A1(net538),
    .S(net268),
    .X(_01165_));
 sg13g2_mux2_1 _23681_ (.A0(\cpu.genblk1.mmu.r_vtop_d[12][11] ),
    .A1(net741),
    .S(net268),
    .X(_01166_));
 sg13g2_mux2_1 _23682_ (.A0(\cpu.genblk1.mmu.r_vtop_d[12][1] ),
    .A1(_03540_),
    .S(net268),
    .X(_01167_));
 sg13g2_mux2_1 _23683_ (.A0(\cpu.genblk1.mmu.r_vtop_d[12][2] ),
    .A1(net743),
    .S(_05908_),
    .X(_01168_));
 sg13g2_mux2_1 _23684_ (.A0(\cpu.genblk1.mmu.r_vtop_d[12][3] ),
    .A1(_03541_),
    .S(net268),
    .X(_01169_));
 sg13g2_mux2_1 _23685_ (.A0(\cpu.genblk1.mmu.r_vtop_d[12][4] ),
    .A1(_03542_),
    .S(net268),
    .X(_01170_));
 sg13g2_mux2_1 _23686_ (.A0(\cpu.genblk1.mmu.r_vtop_d[12][5] ),
    .A1(_03534_),
    .S(_05908_),
    .X(_01171_));
 sg13g2_mux2_1 _23687_ (.A0(\cpu.genblk1.mmu.r_vtop_d[12][6] ),
    .A1(_03538_),
    .S(net268),
    .X(_01172_));
 sg13g2_mux2_1 _23688_ (.A0(\cpu.genblk1.mmu.r_vtop_d[12][7] ),
    .A1(_04782_),
    .S(net268),
    .X(_01173_));
 sg13g2_mux2_1 _23689_ (.A0(\cpu.genblk1.mmu.r_vtop_d[12][8] ),
    .A1(net542),
    .S(_05907_),
    .X(_01174_));
 sg13g2_mux2_1 _23690_ (.A0(\cpu.genblk1.mmu.r_vtop_d[12][9] ),
    .A1(net489),
    .S(_05907_),
    .X(_01175_));
 sg13g2_nand2_2 _23691_ (.Y(_05909_),
    .A(net980),
    .B(_05842_));
 sg13g2_or2_1 _23692_ (.X(_05910_),
    .B(_05882_),
    .A(_05909_));
 sg13g2_buf_2 _23693_ (.A(_05910_),
    .X(_05911_));
 sg13g2_nor2_1 _23694_ (.A(_05905_),
    .B(_05911_),
    .Y(_05912_));
 sg13g2_buf_1 _23695_ (.A(_05912_),
    .X(_05913_));
 sg13g2_buf_1 _23696_ (.A(_05913_),
    .X(_05914_));
 sg13g2_mux2_1 _23697_ (.A0(\cpu.genblk1.mmu.r_vtop_d[13][0] ),
    .A1(net403),
    .S(net267),
    .X(_01176_));
 sg13g2_mux2_1 _23698_ (.A0(\cpu.genblk1.mmu.r_vtop_d[13][10] ),
    .A1(net538),
    .S(net267),
    .X(_01177_));
 sg13g2_mux2_1 _23699_ (.A0(\cpu.genblk1.mmu.r_vtop_d[13][11] ),
    .A1(net741),
    .S(net267),
    .X(_01178_));
 sg13g2_mux2_1 _23700_ (.A0(\cpu.genblk1.mmu.r_vtop_d[13][1] ),
    .A1(_03540_),
    .S(net267),
    .X(_01179_));
 sg13g2_mux2_1 _23701_ (.A0(\cpu.genblk1.mmu.r_vtop_d[13][2] ),
    .A1(net743),
    .S(_05914_),
    .X(_01180_));
 sg13g2_mux2_1 _23702_ (.A0(\cpu.genblk1.mmu.r_vtop_d[13][3] ),
    .A1(_03541_),
    .S(net267),
    .X(_01181_));
 sg13g2_mux2_1 _23703_ (.A0(\cpu.genblk1.mmu.r_vtop_d[13][4] ),
    .A1(_03542_),
    .S(_05914_),
    .X(_01182_));
 sg13g2_buf_1 _23704_ (.A(_10524_),
    .X(_05915_));
 sg13g2_mux2_1 _23705_ (.A0(\cpu.genblk1.mmu.r_vtop_d[13][5] ),
    .A1(net975),
    .S(net267),
    .X(_01183_));
 sg13g2_mux2_1 _23706_ (.A0(\cpu.genblk1.mmu.r_vtop_d[13][6] ),
    .A1(_03538_),
    .S(net267),
    .X(_01184_));
 sg13g2_mux2_1 _23707_ (.A0(\cpu.genblk1.mmu.r_vtop_d[13][7] ),
    .A1(net984),
    .S(net267),
    .X(_01185_));
 sg13g2_mux2_1 _23708_ (.A0(\cpu.genblk1.mmu.r_vtop_d[13][8] ),
    .A1(net542),
    .S(_05913_),
    .X(_01186_));
 sg13g2_mux2_1 _23709_ (.A0(\cpu.genblk1.mmu.r_vtop_d[13][9] ),
    .A1(net489),
    .S(_05913_),
    .X(_01187_));
 sg13g2_buf_1 _23710_ (.A(_05882_),
    .X(_05916_));
 sg13g2_nor3_1 _23711_ (.A(net659),
    .B(net480),
    .C(_05905_),
    .Y(_05917_));
 sg13g2_buf_1 _23712_ (.A(_05917_),
    .X(_05918_));
 sg13g2_buf_1 _23713_ (.A(_05918_),
    .X(_05919_));
 sg13g2_mux2_1 _23714_ (.A0(\cpu.genblk1.mmu.r_vtop_d[14][0] ),
    .A1(_05889_),
    .S(net344),
    .X(_01188_));
 sg13g2_mux2_1 _23715_ (.A0(\cpu.genblk1.mmu.r_vtop_d[14][10] ),
    .A1(net538),
    .S(net344),
    .X(_01189_));
 sg13g2_mux2_1 _23716_ (.A0(\cpu.genblk1.mmu.r_vtop_d[14][11] ),
    .A1(net741),
    .S(net344),
    .X(_01190_));
 sg13g2_buf_1 _23717_ (.A(_03539_),
    .X(_05920_));
 sg13g2_mux2_1 _23718_ (.A0(\cpu.genblk1.mmu.r_vtop_d[14][1] ),
    .A1(_05920_),
    .S(net344),
    .X(_01191_));
 sg13g2_mux2_1 _23719_ (.A0(\cpu.genblk1.mmu.r_vtop_d[14][2] ),
    .A1(net743),
    .S(_05919_),
    .X(_01192_));
 sg13g2_buf_1 _23720_ (.A(_09222_),
    .X(_05921_));
 sg13g2_mux2_1 _23721_ (.A0(\cpu.genblk1.mmu.r_vtop_d[14][3] ),
    .A1(_05921_),
    .S(_05919_),
    .X(_01193_));
 sg13g2_buf_1 _23722_ (.A(_09221_),
    .X(_05922_));
 sg13g2_mux2_1 _23723_ (.A0(\cpu.genblk1.mmu.r_vtop_d[14][4] ),
    .A1(_05922_),
    .S(net344),
    .X(_01194_));
 sg13g2_mux2_1 _23724_ (.A0(\cpu.genblk1.mmu.r_vtop_d[14][5] ),
    .A1(net975),
    .S(net344),
    .X(_01195_));
 sg13g2_buf_1 _23725_ (.A(_10392_),
    .X(_05923_));
 sg13g2_mux2_1 _23726_ (.A0(\cpu.genblk1.mmu.r_vtop_d[14][6] ),
    .A1(_05923_),
    .S(net344),
    .X(_01196_));
 sg13g2_mux2_1 _23727_ (.A0(\cpu.genblk1.mmu.r_vtop_d[14][7] ),
    .A1(net984),
    .S(net344),
    .X(_01197_));
 sg13g2_mux2_1 _23728_ (.A0(\cpu.genblk1.mmu.r_vtop_d[14][8] ),
    .A1(_03550_),
    .S(_05918_),
    .X(_01198_));
 sg13g2_mux2_1 _23729_ (.A0(\cpu.genblk1.mmu.r_vtop_d[14][9] ),
    .A1(_03551_),
    .S(_05918_),
    .X(_01199_));
 sg13g2_nor3_1 _23730_ (.A(_05857_),
    .B(_05916_),
    .C(_05905_),
    .Y(_05924_));
 sg13g2_buf_1 _23731_ (.A(_05924_),
    .X(_05925_));
 sg13g2_buf_1 _23732_ (.A(_05925_),
    .X(_05926_));
 sg13g2_mux2_1 _23733_ (.A0(\cpu.genblk1.mmu.r_vtop_d[15][0] ),
    .A1(_05889_),
    .S(net343),
    .X(_01200_));
 sg13g2_mux2_1 _23734_ (.A0(\cpu.genblk1.mmu.r_vtop_d[15][10] ),
    .A1(net538),
    .S(net343),
    .X(_01201_));
 sg13g2_mux2_1 _23735_ (.A0(\cpu.genblk1.mmu.r_vtop_d[15][11] ),
    .A1(net741),
    .S(net343),
    .X(_01202_));
 sg13g2_mux2_1 _23736_ (.A0(\cpu.genblk1.mmu.r_vtop_d[15][1] ),
    .A1(net658),
    .S(net343),
    .X(_01203_));
 sg13g2_mux2_1 _23737_ (.A0(\cpu.genblk1.mmu.r_vtop_d[15][2] ),
    .A1(_04784_),
    .S(_05926_),
    .X(_01204_));
 sg13g2_mux2_1 _23738_ (.A0(\cpu.genblk1.mmu.r_vtop_d[15][3] ),
    .A1(_05921_),
    .S(net343),
    .X(_01205_));
 sg13g2_mux2_1 _23739_ (.A0(\cpu.genblk1.mmu.r_vtop_d[15][4] ),
    .A1(_05922_),
    .S(_05926_),
    .X(_01206_));
 sg13g2_mux2_1 _23740_ (.A0(\cpu.genblk1.mmu.r_vtop_d[15][5] ),
    .A1(_05915_),
    .S(net343),
    .X(_01207_));
 sg13g2_mux2_1 _23741_ (.A0(\cpu.genblk1.mmu.r_vtop_d[15][6] ),
    .A1(net972),
    .S(net343),
    .X(_01208_));
 sg13g2_mux2_1 _23742_ (.A0(\cpu.genblk1.mmu.r_vtop_d[15][7] ),
    .A1(net984),
    .S(net343),
    .X(_01209_));
 sg13g2_mux2_1 _23743_ (.A0(\cpu.genblk1.mmu.r_vtop_d[15][8] ),
    .A1(_03550_),
    .S(_05925_),
    .X(_01210_));
 sg13g2_mux2_1 _23744_ (.A0(\cpu.genblk1.mmu.r_vtop_d[15][9] ),
    .A1(_03551_),
    .S(_05925_),
    .X(_01211_));
 sg13g2_nand2_1 _23745_ (.Y(_05927_),
    .A(net1121),
    .B(net1044));
 sg13g2_buf_2 _23746_ (.A(_05927_),
    .X(_05928_));
 sg13g2_nand2_2 _23747_ (.Y(_05929_),
    .A(net978),
    .B(_05845_));
 sg13g2_nor3_1 _23748_ (.A(net480),
    .B(_05928_),
    .C(_05929_),
    .Y(_05930_));
 sg13g2_buf_1 _23749_ (.A(_05930_),
    .X(_05931_));
 sg13g2_buf_1 _23750_ (.A(_05931_),
    .X(_05932_));
 sg13g2_mux2_1 _23751_ (.A0(\cpu.genblk1.mmu.r_vtop_d[16][0] ),
    .A1(net403),
    .S(net342),
    .X(_01212_));
 sg13g2_mux2_1 _23752_ (.A0(\cpu.genblk1.mmu.r_vtop_d[16][10] ),
    .A1(net538),
    .S(net342),
    .X(_01213_));
 sg13g2_mux2_1 _23753_ (.A0(\cpu.genblk1.mmu.r_vtop_d[16][11] ),
    .A1(net741),
    .S(net342),
    .X(_01214_));
 sg13g2_mux2_1 _23754_ (.A0(\cpu.genblk1.mmu.r_vtop_d[16][1] ),
    .A1(net658),
    .S(net342),
    .X(_01215_));
 sg13g2_mux2_1 _23755_ (.A0(\cpu.genblk1.mmu.r_vtop_d[16][2] ),
    .A1(net743),
    .S(_05932_),
    .X(_01216_));
 sg13g2_mux2_1 _23756_ (.A0(\cpu.genblk1.mmu.r_vtop_d[16][3] ),
    .A1(net974),
    .S(_05932_),
    .X(_01217_));
 sg13g2_mux2_1 _23757_ (.A0(\cpu.genblk1.mmu.r_vtop_d[16][4] ),
    .A1(net973),
    .S(net342),
    .X(_01218_));
 sg13g2_mux2_1 _23758_ (.A0(\cpu.genblk1.mmu.r_vtop_d[16][5] ),
    .A1(net975),
    .S(net342),
    .X(_01219_));
 sg13g2_mux2_1 _23759_ (.A0(\cpu.genblk1.mmu.r_vtop_d[16][6] ),
    .A1(net972),
    .S(net342),
    .X(_01220_));
 sg13g2_mux2_1 _23760_ (.A0(\cpu.genblk1.mmu.r_vtop_d[16][7] ),
    .A1(net984),
    .S(net342),
    .X(_01221_));
 sg13g2_buf_1 _23761_ (.A(net617),
    .X(_05933_));
 sg13g2_mux2_1 _23762_ (.A0(\cpu.genblk1.mmu.r_vtop_d[16][8] ),
    .A1(_05933_),
    .S(_05931_),
    .X(_01222_));
 sg13g2_buf_1 _23763_ (.A(_09448_),
    .X(_05934_));
 sg13g2_mux2_1 _23764_ (.A0(\cpu.genblk1.mmu.r_vtop_d[16][9] ),
    .A1(net479),
    .S(_05931_),
    .X(_01223_));
 sg13g2_nor3_1 _23765_ (.A(net852),
    .B(_05911_),
    .C(_05928_),
    .Y(_05935_));
 sg13g2_buf_1 _23766_ (.A(_05935_),
    .X(_05936_));
 sg13g2_buf_1 _23767_ (.A(_05936_),
    .X(_05937_));
 sg13g2_mux2_1 _23768_ (.A0(\cpu.genblk1.mmu.r_vtop_d[17][0] ),
    .A1(net403),
    .S(net266),
    .X(_01224_));
 sg13g2_mux2_1 _23769_ (.A0(\cpu.genblk1.mmu.r_vtop_d[17][10] ),
    .A1(net538),
    .S(net266),
    .X(_01225_));
 sg13g2_mux2_1 _23770_ (.A0(\cpu.genblk1.mmu.r_vtop_d[17][11] ),
    .A1(net741),
    .S(net266),
    .X(_01226_));
 sg13g2_mux2_1 _23771_ (.A0(\cpu.genblk1.mmu.r_vtop_d[17][1] ),
    .A1(net658),
    .S(net266),
    .X(_01227_));
 sg13g2_mux2_1 _23772_ (.A0(\cpu.genblk1.mmu.r_vtop_d[17][2] ),
    .A1(net743),
    .S(_05937_),
    .X(_01228_));
 sg13g2_mux2_1 _23773_ (.A0(\cpu.genblk1.mmu.r_vtop_d[17][3] ),
    .A1(net974),
    .S(_05937_),
    .X(_01229_));
 sg13g2_mux2_1 _23774_ (.A0(\cpu.genblk1.mmu.r_vtop_d[17][4] ),
    .A1(net973),
    .S(net266),
    .X(_01230_));
 sg13g2_mux2_1 _23775_ (.A0(\cpu.genblk1.mmu.r_vtop_d[17][5] ),
    .A1(net975),
    .S(net266),
    .X(_01231_));
 sg13g2_mux2_1 _23776_ (.A0(\cpu.genblk1.mmu.r_vtop_d[17][6] ),
    .A1(net972),
    .S(net266),
    .X(_01232_));
 sg13g2_mux2_1 _23777_ (.A0(\cpu.genblk1.mmu.r_vtop_d[17][7] ),
    .A1(net984),
    .S(net266),
    .X(_01233_));
 sg13g2_mux2_1 _23778_ (.A0(\cpu.genblk1.mmu.r_vtop_d[17][8] ),
    .A1(net528),
    .S(_05936_),
    .X(_01234_));
 sg13g2_mux2_1 _23779_ (.A0(\cpu.genblk1.mmu.r_vtop_d[17][9] ),
    .A1(net479),
    .S(_05936_),
    .X(_01235_));
 sg13g2_nand2_2 _23780_ (.Y(_05938_),
    .A(net1121),
    .B(_05840_));
 sg13g2_nor4_2 _23781_ (.A(_05842_),
    .B(net976),
    .C(net977),
    .Y(_05939_),
    .D(_05938_));
 sg13g2_nor2b_1 _23782_ (.A(net481),
    .B_N(_05939_),
    .Y(_05940_));
 sg13g2_buf_1 _23783_ (.A(_05940_),
    .X(_05941_));
 sg13g2_buf_1 _23784_ (.A(_05941_),
    .X(_05942_));
 sg13g2_mux2_1 _23785_ (.A0(\cpu.genblk1.mmu.r_vtop_d[18][0] ),
    .A1(net403),
    .S(net341),
    .X(_01236_));
 sg13g2_buf_1 _23786_ (.A(net688),
    .X(_05943_));
 sg13g2_mux2_1 _23787_ (.A0(\cpu.genblk1.mmu.r_vtop_d[18][10] ),
    .A1(net590),
    .S(net341),
    .X(_01237_));
 sg13g2_mux2_1 _23788_ (.A0(\cpu.genblk1.mmu.r_vtop_d[18][11] ),
    .A1(net741),
    .S(net341),
    .X(_01238_));
 sg13g2_mux2_1 _23789_ (.A0(\cpu.genblk1.mmu.r_vtop_d[18][1] ),
    .A1(net658),
    .S(net341),
    .X(_01239_));
 sg13g2_buf_1 _23790_ (.A(_02959_),
    .X(_05944_));
 sg13g2_mux2_1 _23791_ (.A0(\cpu.genblk1.mmu.r_vtop_d[18][2] ),
    .A1(net851),
    .S(net341),
    .X(_01240_));
 sg13g2_mux2_1 _23792_ (.A0(\cpu.genblk1.mmu.r_vtop_d[18][3] ),
    .A1(net974),
    .S(net341),
    .X(_01241_));
 sg13g2_mux2_1 _23793_ (.A0(\cpu.genblk1.mmu.r_vtop_d[18][4] ),
    .A1(net973),
    .S(_05942_),
    .X(_01242_));
 sg13g2_mux2_1 _23794_ (.A0(\cpu.genblk1.mmu.r_vtop_d[18][5] ),
    .A1(net975),
    .S(_05942_),
    .X(_01243_));
 sg13g2_mux2_1 _23795_ (.A0(\cpu.genblk1.mmu.r_vtop_d[18][6] ),
    .A1(net972),
    .S(net341),
    .X(_01244_));
 sg13g2_buf_1 _23796_ (.A(net1122),
    .X(_05945_));
 sg13g2_mux2_1 _23797_ (.A0(\cpu.genblk1.mmu.r_vtop_d[18][7] ),
    .A1(net971),
    .S(net341),
    .X(_01245_));
 sg13g2_mux2_1 _23798_ (.A0(\cpu.genblk1.mmu.r_vtop_d[18][8] ),
    .A1(_05933_),
    .S(_05941_),
    .X(_01246_));
 sg13g2_mux2_1 _23799_ (.A0(\cpu.genblk1.mmu.r_vtop_d[18][9] ),
    .A1(net479),
    .S(_05941_),
    .X(_01247_));
 sg13g2_nor3_1 _23800_ (.A(net976),
    .B(_05857_),
    .C(_05928_),
    .Y(_05946_));
 sg13g2_buf_1 _23801_ (.A(_05946_),
    .X(_05947_));
 sg13g2_nor2b_1 _23802_ (.A(net481),
    .B_N(_05947_),
    .Y(_05948_));
 sg13g2_buf_1 _23803_ (.A(_05948_),
    .X(_05949_));
 sg13g2_buf_1 _23804_ (.A(_05949_),
    .X(_05950_));
 sg13g2_mux2_1 _23805_ (.A0(\cpu.genblk1.mmu.r_vtop_d[19][0] ),
    .A1(net403),
    .S(net340),
    .X(_01248_));
 sg13g2_mux2_1 _23806_ (.A0(\cpu.genblk1.mmu.r_vtop_d[19][10] ),
    .A1(_05943_),
    .S(net340),
    .X(_01249_));
 sg13g2_buf_1 _23807_ (.A(net860),
    .X(_05951_));
 sg13g2_mux2_1 _23808_ (.A0(\cpu.genblk1.mmu.r_vtop_d[19][11] ),
    .A1(_05951_),
    .S(net340),
    .X(_01250_));
 sg13g2_mux2_1 _23809_ (.A0(\cpu.genblk1.mmu.r_vtop_d[19][1] ),
    .A1(net658),
    .S(net340),
    .X(_01251_));
 sg13g2_mux2_1 _23810_ (.A0(\cpu.genblk1.mmu.r_vtop_d[19][2] ),
    .A1(_05944_),
    .S(net340),
    .X(_01252_));
 sg13g2_mux2_1 _23811_ (.A0(\cpu.genblk1.mmu.r_vtop_d[19][3] ),
    .A1(net974),
    .S(net340),
    .X(_01253_));
 sg13g2_mux2_1 _23812_ (.A0(\cpu.genblk1.mmu.r_vtop_d[19][4] ),
    .A1(net973),
    .S(_05950_),
    .X(_01254_));
 sg13g2_mux2_1 _23813_ (.A0(\cpu.genblk1.mmu.r_vtop_d[19][5] ),
    .A1(net975),
    .S(_05950_),
    .X(_01255_));
 sg13g2_mux2_1 _23814_ (.A0(\cpu.genblk1.mmu.r_vtop_d[19][6] ),
    .A1(net972),
    .S(net340),
    .X(_01256_));
 sg13g2_mux2_1 _23815_ (.A0(\cpu.genblk1.mmu.r_vtop_d[19][7] ),
    .A1(_05945_),
    .S(net340),
    .X(_01257_));
 sg13g2_mux2_1 _23816_ (.A0(\cpu.genblk1.mmu.r_vtop_d[19][8] ),
    .A1(net528),
    .S(_05949_),
    .X(_01258_));
 sg13g2_mux2_1 _23817_ (.A0(\cpu.genblk1.mmu.r_vtop_d[19][9] ),
    .A1(_05934_),
    .S(_05949_),
    .X(_01259_));
 sg13g2_buf_1 _23818_ (.A(net452),
    .X(_05952_));
 sg13g2_nor2_1 _23819_ (.A(_05880_),
    .B(_05911_),
    .Y(_05953_));
 sg13g2_buf_1 _23820_ (.A(_05953_),
    .X(_05954_));
 sg13g2_buf_1 _23821_ (.A(_05954_),
    .X(_05955_));
 sg13g2_mux2_1 _23822_ (.A0(\cpu.genblk1.mmu.r_vtop_d[1][0] ),
    .A1(_05952_),
    .S(net265),
    .X(_01260_));
 sg13g2_mux2_1 _23823_ (.A0(\cpu.genblk1.mmu.r_vtop_d[1][10] ),
    .A1(net590),
    .S(net265),
    .X(_01261_));
 sg13g2_mux2_1 _23824_ (.A0(\cpu.genblk1.mmu.r_vtop_d[1][11] ),
    .A1(_05951_),
    .S(net265),
    .X(_01262_));
 sg13g2_mux2_1 _23825_ (.A0(\cpu.genblk1.mmu.r_vtop_d[1][1] ),
    .A1(_05920_),
    .S(net265),
    .X(_01263_));
 sg13g2_mux2_1 _23826_ (.A0(\cpu.genblk1.mmu.r_vtop_d[1][2] ),
    .A1(_05944_),
    .S(_05955_),
    .X(_01264_));
 sg13g2_mux2_1 _23827_ (.A0(\cpu.genblk1.mmu.r_vtop_d[1][3] ),
    .A1(net974),
    .S(net265),
    .X(_01265_));
 sg13g2_mux2_1 _23828_ (.A0(\cpu.genblk1.mmu.r_vtop_d[1][4] ),
    .A1(net973),
    .S(net265),
    .X(_01266_));
 sg13g2_mux2_1 _23829_ (.A0(\cpu.genblk1.mmu.r_vtop_d[1][5] ),
    .A1(_05915_),
    .S(_05955_),
    .X(_01267_));
 sg13g2_mux2_1 _23830_ (.A0(\cpu.genblk1.mmu.r_vtop_d[1][6] ),
    .A1(_05923_),
    .S(net265),
    .X(_01268_));
 sg13g2_mux2_1 _23831_ (.A0(\cpu.genblk1.mmu.r_vtop_d[1][7] ),
    .A1(_05945_),
    .S(net265),
    .X(_01269_));
 sg13g2_mux2_1 _23832_ (.A0(\cpu.genblk1.mmu.r_vtop_d[1][8] ),
    .A1(net528),
    .S(_05954_),
    .X(_01270_));
 sg13g2_mux2_1 _23833_ (.A0(\cpu.genblk1.mmu.r_vtop_d[1][9] ),
    .A1(_05934_),
    .S(_05954_),
    .X(_01271_));
 sg13g2_or2_1 _23834_ (.X(_05956_),
    .B(_05928_),
    .A(_05877_));
 sg13g2_buf_1 _23835_ (.A(_05956_),
    .X(_05957_));
 sg13g2_nor2_1 _23836_ (.A(_05884_),
    .B(_05957_),
    .Y(_05958_));
 sg13g2_buf_1 _23837_ (.A(_05958_),
    .X(_05959_));
 sg13g2_buf_1 _23838_ (.A(_05959_),
    .X(_05960_));
 sg13g2_mux2_1 _23839_ (.A0(\cpu.genblk1.mmu.r_vtop_d[20][0] ),
    .A1(net402),
    .S(net264),
    .X(_01272_));
 sg13g2_mux2_1 _23840_ (.A0(\cpu.genblk1.mmu.r_vtop_d[20][10] ),
    .A1(net590),
    .S(net264),
    .X(_01273_));
 sg13g2_mux2_1 _23841_ (.A0(\cpu.genblk1.mmu.r_vtop_d[20][11] ),
    .A1(net740),
    .S(net264),
    .X(_01274_));
 sg13g2_mux2_1 _23842_ (.A0(\cpu.genblk1.mmu.r_vtop_d[20][1] ),
    .A1(net658),
    .S(net264),
    .X(_01275_));
 sg13g2_mux2_1 _23843_ (.A0(\cpu.genblk1.mmu.r_vtop_d[20][2] ),
    .A1(net851),
    .S(_05960_),
    .X(_01276_));
 sg13g2_mux2_1 _23844_ (.A0(\cpu.genblk1.mmu.r_vtop_d[20][3] ),
    .A1(net974),
    .S(_05960_),
    .X(_01277_));
 sg13g2_mux2_1 _23845_ (.A0(\cpu.genblk1.mmu.r_vtop_d[20][4] ),
    .A1(net973),
    .S(net264),
    .X(_01278_));
 sg13g2_mux2_1 _23846_ (.A0(\cpu.genblk1.mmu.r_vtop_d[20][5] ),
    .A1(net975),
    .S(net264),
    .X(_01279_));
 sg13g2_mux2_1 _23847_ (.A0(\cpu.genblk1.mmu.r_vtop_d[20][6] ),
    .A1(net972),
    .S(net264),
    .X(_01280_));
 sg13g2_mux2_1 _23848_ (.A0(\cpu.genblk1.mmu.r_vtop_d[20][7] ),
    .A1(net971),
    .S(net264),
    .X(_01281_));
 sg13g2_mux2_1 _23849_ (.A0(\cpu.genblk1.mmu.r_vtop_d[20][8] ),
    .A1(net528),
    .S(_05959_),
    .X(_01282_));
 sg13g2_mux2_1 _23850_ (.A0(\cpu.genblk1.mmu.r_vtop_d[20][9] ),
    .A1(net479),
    .S(_05959_),
    .X(_01283_));
 sg13g2_nor2_1 _23851_ (.A(_05911_),
    .B(_05957_),
    .Y(_05961_));
 sg13g2_buf_1 _23852_ (.A(_05961_),
    .X(_05962_));
 sg13g2_buf_1 _23853_ (.A(_05962_),
    .X(_05963_));
 sg13g2_mux2_1 _23854_ (.A0(\cpu.genblk1.mmu.r_vtop_d[21][0] ),
    .A1(net402),
    .S(net263),
    .X(_01284_));
 sg13g2_mux2_1 _23855_ (.A0(\cpu.genblk1.mmu.r_vtop_d[21][10] ),
    .A1(net590),
    .S(net263),
    .X(_01285_));
 sg13g2_mux2_1 _23856_ (.A0(\cpu.genblk1.mmu.r_vtop_d[21][11] ),
    .A1(net740),
    .S(net263),
    .X(_01286_));
 sg13g2_mux2_1 _23857_ (.A0(\cpu.genblk1.mmu.r_vtop_d[21][1] ),
    .A1(net658),
    .S(net263),
    .X(_01287_));
 sg13g2_mux2_1 _23858_ (.A0(\cpu.genblk1.mmu.r_vtop_d[21][2] ),
    .A1(net851),
    .S(_05963_),
    .X(_01288_));
 sg13g2_mux2_1 _23859_ (.A0(\cpu.genblk1.mmu.r_vtop_d[21][3] ),
    .A1(net974),
    .S(_05963_),
    .X(_01289_));
 sg13g2_mux2_1 _23860_ (.A0(\cpu.genblk1.mmu.r_vtop_d[21][4] ),
    .A1(net973),
    .S(net263),
    .X(_01290_));
 sg13g2_mux2_1 _23861_ (.A0(\cpu.genblk1.mmu.r_vtop_d[21][5] ),
    .A1(net975),
    .S(net263),
    .X(_01291_));
 sg13g2_mux2_1 _23862_ (.A0(\cpu.genblk1.mmu.r_vtop_d[21][6] ),
    .A1(net972),
    .S(net263),
    .X(_01292_));
 sg13g2_mux2_1 _23863_ (.A0(\cpu.genblk1.mmu.r_vtop_d[21][7] ),
    .A1(net971),
    .S(net263),
    .X(_01293_));
 sg13g2_mux2_1 _23864_ (.A0(\cpu.genblk1.mmu.r_vtop_d[21][8] ),
    .A1(net528),
    .S(_05962_),
    .X(_01294_));
 sg13g2_mux2_1 _23865_ (.A0(\cpu.genblk1.mmu.r_vtop_d[21][9] ),
    .A1(net479),
    .S(_05962_),
    .X(_01295_));
 sg13g2_nor3_1 _23866_ (.A(net659),
    .B(net480),
    .C(_05957_),
    .Y(_05964_));
 sg13g2_buf_1 _23867_ (.A(_05964_),
    .X(_05965_));
 sg13g2_buf_1 _23868_ (.A(_05965_),
    .X(_05966_));
 sg13g2_mux2_1 _23869_ (.A0(\cpu.genblk1.mmu.r_vtop_d[22][0] ),
    .A1(net402),
    .S(net339),
    .X(_01296_));
 sg13g2_mux2_1 _23870_ (.A0(\cpu.genblk1.mmu.r_vtop_d[22][10] ),
    .A1(net590),
    .S(net339),
    .X(_01297_));
 sg13g2_mux2_1 _23871_ (.A0(\cpu.genblk1.mmu.r_vtop_d[22][11] ),
    .A1(net740),
    .S(net339),
    .X(_01298_));
 sg13g2_mux2_1 _23872_ (.A0(\cpu.genblk1.mmu.r_vtop_d[22][1] ),
    .A1(net658),
    .S(net339),
    .X(_01299_));
 sg13g2_mux2_1 _23873_ (.A0(\cpu.genblk1.mmu.r_vtop_d[22][2] ),
    .A1(net851),
    .S(_05966_),
    .X(_01300_));
 sg13g2_mux2_1 _23874_ (.A0(\cpu.genblk1.mmu.r_vtop_d[22][3] ),
    .A1(net974),
    .S(_05966_),
    .X(_01301_));
 sg13g2_mux2_1 _23875_ (.A0(\cpu.genblk1.mmu.r_vtop_d[22][4] ),
    .A1(net973),
    .S(net339),
    .X(_01302_));
 sg13g2_buf_1 _23876_ (.A(_10524_),
    .X(_05967_));
 sg13g2_mux2_1 _23877_ (.A0(\cpu.genblk1.mmu.r_vtop_d[22][5] ),
    .A1(net970),
    .S(net339),
    .X(_01303_));
 sg13g2_mux2_1 _23878_ (.A0(\cpu.genblk1.mmu.r_vtop_d[22][6] ),
    .A1(net972),
    .S(net339),
    .X(_01304_));
 sg13g2_mux2_1 _23879_ (.A0(\cpu.genblk1.mmu.r_vtop_d[22][7] ),
    .A1(net971),
    .S(net339),
    .X(_01305_));
 sg13g2_mux2_1 _23880_ (.A0(\cpu.genblk1.mmu.r_vtop_d[22][8] ),
    .A1(net528),
    .S(_05965_),
    .X(_01306_));
 sg13g2_mux2_1 _23881_ (.A0(\cpu.genblk1.mmu.r_vtop_d[22][9] ),
    .A1(net479),
    .S(_05965_),
    .X(_01307_));
 sg13g2_nor3_1 _23882_ (.A(_05857_),
    .B(net480),
    .C(_05957_),
    .Y(_05968_));
 sg13g2_buf_1 _23883_ (.A(_05968_),
    .X(_05969_));
 sg13g2_buf_1 _23884_ (.A(_05969_),
    .X(_05970_));
 sg13g2_mux2_1 _23885_ (.A0(\cpu.genblk1.mmu.r_vtop_d[23][0] ),
    .A1(net402),
    .S(net338),
    .X(_01308_));
 sg13g2_mux2_1 _23886_ (.A0(\cpu.genblk1.mmu.r_vtop_d[23][10] ),
    .A1(_05943_),
    .S(net338),
    .X(_01309_));
 sg13g2_mux2_1 _23887_ (.A0(\cpu.genblk1.mmu.r_vtop_d[23][11] ),
    .A1(net740),
    .S(net338),
    .X(_01310_));
 sg13g2_buf_1 _23888_ (.A(_03539_),
    .X(_05971_));
 sg13g2_mux2_1 _23889_ (.A0(\cpu.genblk1.mmu.r_vtop_d[23][1] ),
    .A1(net657),
    .S(net338),
    .X(_01311_));
 sg13g2_mux2_1 _23890_ (.A0(\cpu.genblk1.mmu.r_vtop_d[23][2] ),
    .A1(net851),
    .S(_05970_),
    .X(_01312_));
 sg13g2_buf_1 _23891_ (.A(net1138),
    .X(_05972_));
 sg13g2_mux2_1 _23892_ (.A0(\cpu.genblk1.mmu.r_vtop_d[23][3] ),
    .A1(_05972_),
    .S(_05970_),
    .X(_01313_));
 sg13g2_buf_1 _23893_ (.A(net1139),
    .X(_05973_));
 sg13g2_mux2_1 _23894_ (.A0(\cpu.genblk1.mmu.r_vtop_d[23][4] ),
    .A1(_05973_),
    .S(net338),
    .X(_01314_));
 sg13g2_mux2_1 _23895_ (.A0(\cpu.genblk1.mmu.r_vtop_d[23][5] ),
    .A1(_05967_),
    .S(net338),
    .X(_01315_));
 sg13g2_buf_1 _23896_ (.A(_10392_),
    .X(_05974_));
 sg13g2_mux2_1 _23897_ (.A0(\cpu.genblk1.mmu.r_vtop_d[23][6] ),
    .A1(net967),
    .S(net338),
    .X(_01316_));
 sg13g2_mux2_1 _23898_ (.A0(\cpu.genblk1.mmu.r_vtop_d[23][7] ),
    .A1(net971),
    .S(net338),
    .X(_01317_));
 sg13g2_mux2_1 _23899_ (.A0(\cpu.genblk1.mmu.r_vtop_d[23][8] ),
    .A1(net528),
    .S(_05969_),
    .X(_01318_));
 sg13g2_mux2_1 _23900_ (.A0(\cpu.genblk1.mmu.r_vtop_d[23][9] ),
    .A1(net479),
    .S(_05969_),
    .X(_01319_));
 sg13g2_nand2_1 _23901_ (.Y(_05975_),
    .A(net1121),
    .B(_10443_));
 sg13g2_buf_1 _23902_ (.A(_05975_),
    .X(_05976_));
 sg13g2_nor3_1 _23903_ (.A(net480),
    .B(_05929_),
    .C(_05976_),
    .Y(_05977_));
 sg13g2_buf_1 _23904_ (.A(_05977_),
    .X(_05978_));
 sg13g2_buf_1 _23905_ (.A(_05978_),
    .X(_05979_));
 sg13g2_mux2_1 _23906_ (.A0(\cpu.genblk1.mmu.r_vtop_d[24][0] ),
    .A1(_05952_),
    .S(net337),
    .X(_01320_));
 sg13g2_mux2_1 _23907_ (.A0(\cpu.genblk1.mmu.r_vtop_d[24][10] ),
    .A1(net590),
    .S(net337),
    .X(_01321_));
 sg13g2_mux2_1 _23908_ (.A0(\cpu.genblk1.mmu.r_vtop_d[24][11] ),
    .A1(net740),
    .S(net337),
    .X(_01322_));
 sg13g2_mux2_1 _23909_ (.A0(\cpu.genblk1.mmu.r_vtop_d[24][1] ),
    .A1(net657),
    .S(_05979_),
    .X(_01323_));
 sg13g2_mux2_1 _23910_ (.A0(\cpu.genblk1.mmu.r_vtop_d[24][2] ),
    .A1(net851),
    .S(net337),
    .X(_01324_));
 sg13g2_mux2_1 _23911_ (.A0(\cpu.genblk1.mmu.r_vtop_d[24][3] ),
    .A1(net969),
    .S(net337),
    .X(_01325_));
 sg13g2_mux2_1 _23912_ (.A0(\cpu.genblk1.mmu.r_vtop_d[24][4] ),
    .A1(net968),
    .S(net337),
    .X(_01326_));
 sg13g2_mux2_1 _23913_ (.A0(\cpu.genblk1.mmu.r_vtop_d[24][5] ),
    .A1(net970),
    .S(net337),
    .X(_01327_));
 sg13g2_mux2_1 _23914_ (.A0(\cpu.genblk1.mmu.r_vtop_d[24][6] ),
    .A1(net967),
    .S(_05979_),
    .X(_01328_));
 sg13g2_mux2_1 _23915_ (.A0(\cpu.genblk1.mmu.r_vtop_d[24][7] ),
    .A1(net971),
    .S(net337),
    .X(_01329_));
 sg13g2_mux2_1 _23916_ (.A0(\cpu.genblk1.mmu.r_vtop_d[24][8] ),
    .A1(net528),
    .S(_05978_),
    .X(_01330_));
 sg13g2_mux2_1 _23917_ (.A0(\cpu.genblk1.mmu.r_vtop_d[24][9] ),
    .A1(net479),
    .S(_05978_),
    .X(_01331_));
 sg13g2_nor3_1 _23918_ (.A(net852),
    .B(_05911_),
    .C(_05976_),
    .Y(_05980_));
 sg13g2_buf_1 _23919_ (.A(_05980_),
    .X(_05981_));
 sg13g2_buf_1 _23920_ (.A(_05981_),
    .X(_05982_));
 sg13g2_mux2_1 _23921_ (.A0(\cpu.genblk1.mmu.r_vtop_d[25][0] ),
    .A1(net402),
    .S(net262),
    .X(_01332_));
 sg13g2_mux2_1 _23922_ (.A0(\cpu.genblk1.mmu.r_vtop_d[25][10] ),
    .A1(net590),
    .S(net262),
    .X(_01333_));
 sg13g2_mux2_1 _23923_ (.A0(\cpu.genblk1.mmu.r_vtop_d[25][11] ),
    .A1(net740),
    .S(net262),
    .X(_01334_));
 sg13g2_mux2_1 _23924_ (.A0(\cpu.genblk1.mmu.r_vtop_d[25][1] ),
    .A1(net657),
    .S(_05982_),
    .X(_01335_));
 sg13g2_mux2_1 _23925_ (.A0(\cpu.genblk1.mmu.r_vtop_d[25][2] ),
    .A1(net851),
    .S(net262),
    .X(_01336_));
 sg13g2_mux2_1 _23926_ (.A0(\cpu.genblk1.mmu.r_vtop_d[25][3] ),
    .A1(net969),
    .S(net262),
    .X(_01337_));
 sg13g2_mux2_1 _23927_ (.A0(\cpu.genblk1.mmu.r_vtop_d[25][4] ),
    .A1(net968),
    .S(net262),
    .X(_01338_));
 sg13g2_mux2_1 _23928_ (.A0(\cpu.genblk1.mmu.r_vtop_d[25][5] ),
    .A1(net970),
    .S(net262),
    .X(_01339_));
 sg13g2_mux2_1 _23929_ (.A0(\cpu.genblk1.mmu.r_vtop_d[25][6] ),
    .A1(net967),
    .S(_05982_),
    .X(_01340_));
 sg13g2_mux2_1 _23930_ (.A0(\cpu.genblk1.mmu.r_vtop_d[25][7] ),
    .A1(net971),
    .S(net262),
    .X(_01341_));
 sg13g2_buf_1 _23931_ (.A(_10341_),
    .X(_05983_));
 sg13g2_mux2_1 _23932_ (.A0(\cpu.genblk1.mmu.r_vtop_d[25][8] ),
    .A1(net527),
    .S(_05981_),
    .X(_01342_));
 sg13g2_buf_1 _23933_ (.A(_09448_),
    .X(_05984_));
 sg13g2_mux2_1 _23934_ (.A0(\cpu.genblk1.mmu.r_vtop_d[25][9] ),
    .A1(net478),
    .S(_05981_),
    .X(_01343_));
 sg13g2_nor4_2 _23935_ (.A(_05842_),
    .B(net976),
    .C(net1044),
    .Y(_05985_),
    .D(_05938_));
 sg13g2_nor2b_1 _23936_ (.A(net481),
    .B_N(_05985_),
    .Y(_05986_));
 sg13g2_buf_1 _23937_ (.A(_05986_),
    .X(_05987_));
 sg13g2_buf_1 _23938_ (.A(_05987_),
    .X(_05988_));
 sg13g2_mux2_1 _23939_ (.A0(\cpu.genblk1.mmu.r_vtop_d[26][0] ),
    .A1(net402),
    .S(net336),
    .X(_01344_));
 sg13g2_mux2_1 _23940_ (.A0(\cpu.genblk1.mmu.r_vtop_d[26][10] ),
    .A1(net590),
    .S(net336),
    .X(_01345_));
 sg13g2_mux2_1 _23941_ (.A0(\cpu.genblk1.mmu.r_vtop_d[26][11] ),
    .A1(net740),
    .S(net336),
    .X(_01346_));
 sg13g2_mux2_1 _23942_ (.A0(\cpu.genblk1.mmu.r_vtop_d[26][1] ),
    .A1(net657),
    .S(_05988_),
    .X(_01347_));
 sg13g2_mux2_1 _23943_ (.A0(\cpu.genblk1.mmu.r_vtop_d[26][2] ),
    .A1(net851),
    .S(net336),
    .X(_01348_));
 sg13g2_mux2_1 _23944_ (.A0(\cpu.genblk1.mmu.r_vtop_d[26][3] ),
    .A1(net969),
    .S(net336),
    .X(_01349_));
 sg13g2_mux2_1 _23945_ (.A0(\cpu.genblk1.mmu.r_vtop_d[26][4] ),
    .A1(net968),
    .S(net336),
    .X(_01350_));
 sg13g2_mux2_1 _23946_ (.A0(\cpu.genblk1.mmu.r_vtop_d[26][5] ),
    .A1(net970),
    .S(net336),
    .X(_01351_));
 sg13g2_mux2_1 _23947_ (.A0(\cpu.genblk1.mmu.r_vtop_d[26][6] ),
    .A1(net967),
    .S(_05988_),
    .X(_01352_));
 sg13g2_mux2_1 _23948_ (.A0(\cpu.genblk1.mmu.r_vtop_d[26][7] ),
    .A1(net971),
    .S(net336),
    .X(_01353_));
 sg13g2_mux2_1 _23949_ (.A0(\cpu.genblk1.mmu.r_vtop_d[26][8] ),
    .A1(net527),
    .S(_05987_),
    .X(_01354_));
 sg13g2_mux2_1 _23950_ (.A0(\cpu.genblk1.mmu.r_vtop_d[26][9] ),
    .A1(net478),
    .S(_05987_),
    .X(_01355_));
 sg13g2_nor3_1 _23951_ (.A(net976),
    .B(_05857_),
    .C(_05976_),
    .Y(_05989_));
 sg13g2_buf_1 _23952_ (.A(_05989_),
    .X(_05990_));
 sg13g2_nor2b_1 _23953_ (.A(net481),
    .B_N(_05990_),
    .Y(_05991_));
 sg13g2_buf_1 _23954_ (.A(_05991_),
    .X(_05992_));
 sg13g2_buf_1 _23955_ (.A(_05992_),
    .X(_05993_));
 sg13g2_mux2_1 _23956_ (.A0(\cpu.genblk1.mmu.r_vtop_d[27][0] ),
    .A1(net402),
    .S(net335),
    .X(_01356_));
 sg13g2_buf_1 _23957_ (.A(_09643_),
    .X(_05994_));
 sg13g2_mux2_1 _23958_ (.A0(\cpu.genblk1.mmu.r_vtop_d[27][10] ),
    .A1(net589),
    .S(net335),
    .X(_01357_));
 sg13g2_mux2_1 _23959_ (.A0(\cpu.genblk1.mmu.r_vtop_d[27][11] ),
    .A1(net740),
    .S(net335),
    .X(_01358_));
 sg13g2_mux2_1 _23960_ (.A0(\cpu.genblk1.mmu.r_vtop_d[27][1] ),
    .A1(net657),
    .S(_05993_),
    .X(_01359_));
 sg13g2_buf_1 _23961_ (.A(_02959_),
    .X(_05995_));
 sg13g2_mux2_1 _23962_ (.A0(\cpu.genblk1.mmu.r_vtop_d[27][2] ),
    .A1(net850),
    .S(net335),
    .X(_01360_));
 sg13g2_mux2_1 _23963_ (.A0(\cpu.genblk1.mmu.r_vtop_d[27][3] ),
    .A1(net969),
    .S(net335),
    .X(_01361_));
 sg13g2_mux2_1 _23964_ (.A0(\cpu.genblk1.mmu.r_vtop_d[27][4] ),
    .A1(net968),
    .S(net335),
    .X(_01362_));
 sg13g2_mux2_1 _23965_ (.A0(\cpu.genblk1.mmu.r_vtop_d[27][5] ),
    .A1(net970),
    .S(net335),
    .X(_01363_));
 sg13g2_mux2_1 _23966_ (.A0(\cpu.genblk1.mmu.r_vtop_d[27][6] ),
    .A1(net967),
    .S(_05993_),
    .X(_01364_));
 sg13g2_buf_1 _23967_ (.A(_10379_),
    .X(_05996_));
 sg13g2_mux2_1 _23968_ (.A0(\cpu.genblk1.mmu.r_vtop_d[27][7] ),
    .A1(net966),
    .S(net335),
    .X(_01365_));
 sg13g2_mux2_1 _23969_ (.A0(\cpu.genblk1.mmu.r_vtop_d[27][8] ),
    .A1(net527),
    .S(_05992_),
    .X(_01366_));
 sg13g2_mux2_1 _23970_ (.A0(\cpu.genblk1.mmu.r_vtop_d[27][9] ),
    .A1(net478),
    .S(_05992_),
    .X(_01367_));
 sg13g2_or2_1 _23971_ (.X(_05997_),
    .B(_05976_),
    .A(_05877_));
 sg13g2_buf_1 _23972_ (.A(_05997_),
    .X(_05998_));
 sg13g2_nor2_1 _23973_ (.A(_05884_),
    .B(_05998_),
    .Y(_05999_));
 sg13g2_buf_1 _23974_ (.A(_05999_),
    .X(_06000_));
 sg13g2_buf_1 _23975_ (.A(_06000_),
    .X(_06001_));
 sg13g2_mux2_1 _23976_ (.A0(\cpu.genblk1.mmu.r_vtop_d[28][0] ),
    .A1(net402),
    .S(net261),
    .X(_01368_));
 sg13g2_mux2_1 _23977_ (.A0(\cpu.genblk1.mmu.r_vtop_d[28][10] ),
    .A1(net589),
    .S(net261),
    .X(_01369_));
 sg13g2_buf_1 _23978_ (.A(net860),
    .X(_06002_));
 sg13g2_mux2_1 _23979_ (.A0(\cpu.genblk1.mmu.r_vtop_d[28][11] ),
    .A1(net739),
    .S(net261),
    .X(_01370_));
 sg13g2_mux2_1 _23980_ (.A0(\cpu.genblk1.mmu.r_vtop_d[28][1] ),
    .A1(net657),
    .S(net261),
    .X(_01371_));
 sg13g2_mux2_1 _23981_ (.A0(\cpu.genblk1.mmu.r_vtop_d[28][2] ),
    .A1(net850),
    .S(net261),
    .X(_01372_));
 sg13g2_mux2_1 _23982_ (.A0(\cpu.genblk1.mmu.r_vtop_d[28][3] ),
    .A1(net969),
    .S(_06001_),
    .X(_01373_));
 sg13g2_mux2_1 _23983_ (.A0(\cpu.genblk1.mmu.r_vtop_d[28][4] ),
    .A1(net968),
    .S(_06001_),
    .X(_01374_));
 sg13g2_mux2_1 _23984_ (.A0(\cpu.genblk1.mmu.r_vtop_d[28][5] ),
    .A1(net970),
    .S(net261),
    .X(_01375_));
 sg13g2_mux2_1 _23985_ (.A0(\cpu.genblk1.mmu.r_vtop_d[28][6] ),
    .A1(net967),
    .S(net261),
    .X(_01376_));
 sg13g2_mux2_1 _23986_ (.A0(\cpu.genblk1.mmu.r_vtop_d[28][7] ),
    .A1(net966),
    .S(net261),
    .X(_01377_));
 sg13g2_mux2_1 _23987_ (.A0(\cpu.genblk1.mmu.r_vtop_d[28][8] ),
    .A1(_05983_),
    .S(_06000_),
    .X(_01378_));
 sg13g2_mux2_1 _23988_ (.A0(\cpu.genblk1.mmu.r_vtop_d[28][9] ),
    .A1(net478),
    .S(_06000_),
    .X(_01379_));
 sg13g2_buf_1 _23989_ (.A(_03513_),
    .X(_06003_));
 sg13g2_nor2_1 _23990_ (.A(_05911_),
    .B(_05998_),
    .Y(_06004_));
 sg13g2_buf_1 _23991_ (.A(_06004_),
    .X(_06005_));
 sg13g2_buf_1 _23992_ (.A(_06005_),
    .X(_06006_));
 sg13g2_mux2_1 _23993_ (.A0(\cpu.genblk1.mmu.r_vtop_d[29][0] ),
    .A1(net401),
    .S(net260),
    .X(_01380_));
 sg13g2_mux2_1 _23994_ (.A0(\cpu.genblk1.mmu.r_vtop_d[29][10] ),
    .A1(net589),
    .S(net260),
    .X(_01381_));
 sg13g2_mux2_1 _23995_ (.A0(\cpu.genblk1.mmu.r_vtop_d[29][11] ),
    .A1(net739),
    .S(net260),
    .X(_01382_));
 sg13g2_mux2_1 _23996_ (.A0(\cpu.genblk1.mmu.r_vtop_d[29][1] ),
    .A1(net657),
    .S(net260),
    .X(_01383_));
 sg13g2_mux2_1 _23997_ (.A0(\cpu.genblk1.mmu.r_vtop_d[29][2] ),
    .A1(net850),
    .S(net260),
    .X(_01384_));
 sg13g2_mux2_1 _23998_ (.A0(\cpu.genblk1.mmu.r_vtop_d[29][3] ),
    .A1(net969),
    .S(_06006_),
    .X(_01385_));
 sg13g2_mux2_1 _23999_ (.A0(\cpu.genblk1.mmu.r_vtop_d[29][4] ),
    .A1(net968),
    .S(_06006_),
    .X(_01386_));
 sg13g2_mux2_1 _24000_ (.A0(\cpu.genblk1.mmu.r_vtop_d[29][5] ),
    .A1(net970),
    .S(net260),
    .X(_01387_));
 sg13g2_mux2_1 _24001_ (.A0(\cpu.genblk1.mmu.r_vtop_d[29][6] ),
    .A1(net967),
    .S(net260),
    .X(_01388_));
 sg13g2_mux2_1 _24002_ (.A0(\cpu.genblk1.mmu.r_vtop_d[29][7] ),
    .A1(net966),
    .S(net260),
    .X(_01389_));
 sg13g2_mux2_1 _24003_ (.A0(\cpu.genblk1.mmu.r_vtop_d[29][8] ),
    .A1(net527),
    .S(_06005_),
    .X(_01390_));
 sg13g2_mux2_1 _24004_ (.A0(\cpu.genblk1.mmu.r_vtop_d[29][9] ),
    .A1(net478),
    .S(_06005_),
    .X(_01391_));
 sg13g2_nor3_1 _24005_ (.A(net659),
    .B(_05880_),
    .C(net481),
    .Y(_06007_));
 sg13g2_buf_1 _24006_ (.A(_06007_),
    .X(_06008_));
 sg13g2_buf_1 _24007_ (.A(_06008_),
    .X(_06009_));
 sg13g2_mux2_1 _24008_ (.A0(\cpu.genblk1.mmu.r_vtop_d[2][0] ),
    .A1(net401),
    .S(_06009_),
    .X(_01392_));
 sg13g2_mux2_1 _24009_ (.A0(\cpu.genblk1.mmu.r_vtop_d[2][10] ),
    .A1(net589),
    .S(net334),
    .X(_01393_));
 sg13g2_mux2_1 _24010_ (.A0(\cpu.genblk1.mmu.r_vtop_d[2][11] ),
    .A1(_06002_),
    .S(net334),
    .X(_01394_));
 sg13g2_mux2_1 _24011_ (.A0(\cpu.genblk1.mmu.r_vtop_d[2][1] ),
    .A1(_05971_),
    .S(_06009_),
    .X(_01395_));
 sg13g2_mux2_1 _24012_ (.A0(\cpu.genblk1.mmu.r_vtop_d[2][2] ),
    .A1(_05995_),
    .S(net334),
    .X(_01396_));
 sg13g2_mux2_1 _24013_ (.A0(\cpu.genblk1.mmu.r_vtop_d[2][3] ),
    .A1(_05972_),
    .S(net334),
    .X(_01397_));
 sg13g2_mux2_1 _24014_ (.A0(\cpu.genblk1.mmu.r_vtop_d[2][4] ),
    .A1(_05973_),
    .S(net334),
    .X(_01398_));
 sg13g2_mux2_1 _24015_ (.A0(\cpu.genblk1.mmu.r_vtop_d[2][5] ),
    .A1(_05967_),
    .S(net334),
    .X(_01399_));
 sg13g2_mux2_1 _24016_ (.A0(\cpu.genblk1.mmu.r_vtop_d[2][6] ),
    .A1(_05974_),
    .S(net334),
    .X(_01400_));
 sg13g2_mux2_1 _24017_ (.A0(\cpu.genblk1.mmu.r_vtop_d[2][7] ),
    .A1(_05996_),
    .S(net334),
    .X(_01401_));
 sg13g2_mux2_1 _24018_ (.A0(\cpu.genblk1.mmu.r_vtop_d[2][8] ),
    .A1(net527),
    .S(_06008_),
    .X(_01402_));
 sg13g2_mux2_1 _24019_ (.A0(\cpu.genblk1.mmu.r_vtop_d[2][9] ),
    .A1(net478),
    .S(_06008_),
    .X(_01403_));
 sg13g2_nor3_1 _24020_ (.A(net659),
    .B(net480),
    .C(_05998_),
    .Y(_06010_));
 sg13g2_buf_1 _24021_ (.A(_06010_),
    .X(_06011_));
 sg13g2_buf_1 _24022_ (.A(_06011_),
    .X(_06012_));
 sg13g2_mux2_1 _24023_ (.A0(\cpu.genblk1.mmu.r_vtop_d[30][0] ),
    .A1(net401),
    .S(net333),
    .X(_01404_));
 sg13g2_mux2_1 _24024_ (.A0(\cpu.genblk1.mmu.r_vtop_d[30][10] ),
    .A1(_05994_),
    .S(net333),
    .X(_01405_));
 sg13g2_mux2_1 _24025_ (.A0(\cpu.genblk1.mmu.r_vtop_d[30][11] ),
    .A1(net739),
    .S(net333),
    .X(_01406_));
 sg13g2_mux2_1 _24026_ (.A0(\cpu.genblk1.mmu.r_vtop_d[30][1] ),
    .A1(net657),
    .S(net333),
    .X(_01407_));
 sg13g2_mux2_1 _24027_ (.A0(\cpu.genblk1.mmu.r_vtop_d[30][2] ),
    .A1(net850),
    .S(net333),
    .X(_01408_));
 sg13g2_mux2_1 _24028_ (.A0(\cpu.genblk1.mmu.r_vtop_d[30][3] ),
    .A1(net969),
    .S(_06012_),
    .X(_01409_));
 sg13g2_mux2_1 _24029_ (.A0(\cpu.genblk1.mmu.r_vtop_d[30][4] ),
    .A1(net968),
    .S(_06012_),
    .X(_01410_));
 sg13g2_mux2_1 _24030_ (.A0(\cpu.genblk1.mmu.r_vtop_d[30][5] ),
    .A1(net970),
    .S(net333),
    .X(_01411_));
 sg13g2_mux2_1 _24031_ (.A0(\cpu.genblk1.mmu.r_vtop_d[30][6] ),
    .A1(_05974_),
    .S(net333),
    .X(_01412_));
 sg13g2_mux2_1 _24032_ (.A0(\cpu.genblk1.mmu.r_vtop_d[30][7] ),
    .A1(net966),
    .S(net333),
    .X(_01413_));
 sg13g2_mux2_1 _24033_ (.A0(\cpu.genblk1.mmu.r_vtop_d[30][8] ),
    .A1(_05983_),
    .S(_06011_),
    .X(_01414_));
 sg13g2_mux2_1 _24034_ (.A0(\cpu.genblk1.mmu.r_vtop_d[30][9] ),
    .A1(_05984_),
    .S(_06011_),
    .X(_01415_));
 sg13g2_nor3_1 _24035_ (.A(_05857_),
    .B(net480),
    .C(_05998_),
    .Y(_06013_));
 sg13g2_buf_1 _24036_ (.A(_06013_),
    .X(_06014_));
 sg13g2_buf_1 _24037_ (.A(_06014_),
    .X(_06015_));
 sg13g2_mux2_1 _24038_ (.A0(\cpu.genblk1.mmu.r_vtop_d[31][0] ),
    .A1(net401),
    .S(net332),
    .X(_01416_));
 sg13g2_mux2_1 _24039_ (.A0(\cpu.genblk1.mmu.r_vtop_d[31][10] ),
    .A1(_05994_),
    .S(net332),
    .X(_01417_));
 sg13g2_mux2_1 _24040_ (.A0(\cpu.genblk1.mmu.r_vtop_d[31][11] ),
    .A1(net739),
    .S(net332),
    .X(_01418_));
 sg13g2_mux2_1 _24041_ (.A0(\cpu.genblk1.mmu.r_vtop_d[31][1] ),
    .A1(_05971_),
    .S(net332),
    .X(_01419_));
 sg13g2_mux2_1 _24042_ (.A0(\cpu.genblk1.mmu.r_vtop_d[31][2] ),
    .A1(net850),
    .S(net332),
    .X(_01420_));
 sg13g2_mux2_1 _24043_ (.A0(\cpu.genblk1.mmu.r_vtop_d[31][3] ),
    .A1(net969),
    .S(_06015_),
    .X(_01421_));
 sg13g2_mux2_1 _24044_ (.A0(\cpu.genblk1.mmu.r_vtop_d[31][4] ),
    .A1(net968),
    .S(_06015_),
    .X(_01422_));
 sg13g2_mux2_1 _24045_ (.A0(\cpu.genblk1.mmu.r_vtop_d[31][5] ),
    .A1(_02985_),
    .S(net332),
    .X(_01423_));
 sg13g2_mux2_1 _24046_ (.A0(\cpu.genblk1.mmu.r_vtop_d[31][6] ),
    .A1(net967),
    .S(net332),
    .X(_01424_));
 sg13g2_mux2_1 _24047_ (.A0(\cpu.genblk1.mmu.r_vtop_d[31][7] ),
    .A1(net966),
    .S(net332),
    .X(_01425_));
 sg13g2_mux2_1 _24048_ (.A0(\cpu.genblk1.mmu.r_vtop_d[31][8] ),
    .A1(net527),
    .S(_06014_),
    .X(_01426_));
 sg13g2_mux2_1 _24049_ (.A0(\cpu.genblk1.mmu.r_vtop_d[31][9] ),
    .A1(net478),
    .S(_06014_),
    .X(_01427_));
 sg13g2_nor3_1 _24050_ (.A(_05857_),
    .B(_05880_),
    .C(net480),
    .Y(_06016_));
 sg13g2_buf_1 _24051_ (.A(_06016_),
    .X(_06017_));
 sg13g2_buf_1 _24052_ (.A(_06017_),
    .X(_06018_));
 sg13g2_mux2_1 _24053_ (.A0(\cpu.genblk1.mmu.r_vtop_d[3][0] ),
    .A1(net401),
    .S(net331),
    .X(_01428_));
 sg13g2_mux2_1 _24054_ (.A0(\cpu.genblk1.mmu.r_vtop_d[3][10] ),
    .A1(net589),
    .S(net331),
    .X(_01429_));
 sg13g2_mux2_1 _24055_ (.A0(\cpu.genblk1.mmu.r_vtop_d[3][11] ),
    .A1(_06002_),
    .S(net331),
    .X(_01430_));
 sg13g2_mux2_1 _24056_ (.A0(\cpu.genblk1.mmu.r_vtop_d[3][1] ),
    .A1(net668),
    .S(net331),
    .X(_01431_));
 sg13g2_mux2_1 _24057_ (.A0(\cpu.genblk1.mmu.r_vtop_d[3][2] ),
    .A1(_05995_),
    .S(_06018_),
    .X(_01432_));
 sg13g2_mux2_1 _24058_ (.A0(\cpu.genblk1.mmu.r_vtop_d[3][3] ),
    .A1(net998),
    .S(net331),
    .X(_01433_));
 sg13g2_mux2_1 _24059_ (.A0(\cpu.genblk1.mmu.r_vtop_d[3][4] ),
    .A1(net997),
    .S(net331),
    .X(_01434_));
 sg13g2_mux2_1 _24060_ (.A0(\cpu.genblk1.mmu.r_vtop_d[3][5] ),
    .A1(net996),
    .S(_06018_),
    .X(_01435_));
 sg13g2_mux2_1 _24061_ (.A0(\cpu.genblk1.mmu.r_vtop_d[3][6] ),
    .A1(net995),
    .S(net331),
    .X(_01436_));
 sg13g2_mux2_1 _24062_ (.A0(\cpu.genblk1.mmu.r_vtop_d[3][7] ),
    .A1(_05996_),
    .S(net331),
    .X(_01437_));
 sg13g2_mux2_1 _24063_ (.A0(\cpu.genblk1.mmu.r_vtop_d[3][8] ),
    .A1(net527),
    .S(_06017_),
    .X(_01438_));
 sg13g2_mux2_1 _24064_ (.A0(\cpu.genblk1.mmu.r_vtop_d[3][9] ),
    .A1(net478),
    .S(_06017_),
    .X(_01439_));
 sg13g2_nand2_1 _24065_ (.Y(_06019_),
    .A(_05866_),
    .B(_05879_));
 sg13g2_nor2_1 _24066_ (.A(_05884_),
    .B(_06019_),
    .Y(_06020_));
 sg13g2_buf_1 _24067_ (.A(_06020_),
    .X(_06021_));
 sg13g2_buf_1 _24068_ (.A(_06021_),
    .X(_06022_));
 sg13g2_mux2_1 _24069_ (.A0(\cpu.genblk1.mmu.r_vtop_d[4][0] ),
    .A1(net401),
    .S(net259),
    .X(_01440_));
 sg13g2_mux2_1 _24070_ (.A0(\cpu.genblk1.mmu.r_vtop_d[4][10] ),
    .A1(net589),
    .S(net259),
    .X(_01441_));
 sg13g2_mux2_1 _24071_ (.A0(\cpu.genblk1.mmu.r_vtop_d[4][11] ),
    .A1(net739),
    .S(net259),
    .X(_01442_));
 sg13g2_mux2_1 _24072_ (.A0(\cpu.genblk1.mmu.r_vtop_d[4][1] ),
    .A1(net668),
    .S(net259),
    .X(_01443_));
 sg13g2_mux2_1 _24073_ (.A0(\cpu.genblk1.mmu.r_vtop_d[4][2] ),
    .A1(net850),
    .S(net259),
    .X(_01444_));
 sg13g2_mux2_1 _24074_ (.A0(\cpu.genblk1.mmu.r_vtop_d[4][3] ),
    .A1(net998),
    .S(net259),
    .X(_01445_));
 sg13g2_mux2_1 _24075_ (.A0(\cpu.genblk1.mmu.r_vtop_d[4][4] ),
    .A1(net997),
    .S(_06022_),
    .X(_01446_));
 sg13g2_mux2_1 _24076_ (.A0(\cpu.genblk1.mmu.r_vtop_d[4][5] ),
    .A1(net996),
    .S(_06022_),
    .X(_01447_));
 sg13g2_mux2_1 _24077_ (.A0(\cpu.genblk1.mmu.r_vtop_d[4][6] ),
    .A1(net995),
    .S(net259),
    .X(_01448_));
 sg13g2_mux2_1 _24078_ (.A0(\cpu.genblk1.mmu.r_vtop_d[4][7] ),
    .A1(net966),
    .S(net259),
    .X(_01449_));
 sg13g2_mux2_1 _24079_ (.A0(\cpu.genblk1.mmu.r_vtop_d[4][8] ),
    .A1(net527),
    .S(_06021_),
    .X(_01450_));
 sg13g2_mux2_1 _24080_ (.A0(\cpu.genblk1.mmu.r_vtop_d[4][9] ),
    .A1(_05984_),
    .S(_06021_),
    .X(_01451_));
 sg13g2_nor2_1 _24081_ (.A(_05909_),
    .B(_06019_),
    .Y(_06023_));
 sg13g2_buf_2 _24082_ (.A(_06023_),
    .X(_06024_));
 sg13g2_nor2b_1 _24083_ (.A(net481),
    .B_N(_06024_),
    .Y(_06025_));
 sg13g2_buf_1 _24084_ (.A(_06025_),
    .X(_06026_));
 sg13g2_buf_1 _24085_ (.A(_06026_),
    .X(_06027_));
 sg13g2_mux2_1 _24086_ (.A0(\cpu.genblk1.mmu.r_vtop_d[5][0] ),
    .A1(net401),
    .S(net330),
    .X(_01452_));
 sg13g2_mux2_1 _24087_ (.A0(\cpu.genblk1.mmu.r_vtop_d[5][10] ),
    .A1(net589),
    .S(net330),
    .X(_01453_));
 sg13g2_mux2_1 _24088_ (.A0(\cpu.genblk1.mmu.r_vtop_d[5][11] ),
    .A1(net739),
    .S(net330),
    .X(_01454_));
 sg13g2_mux2_1 _24089_ (.A0(\cpu.genblk1.mmu.r_vtop_d[5][1] ),
    .A1(net668),
    .S(net330),
    .X(_01455_));
 sg13g2_mux2_1 _24090_ (.A0(\cpu.genblk1.mmu.r_vtop_d[5][2] ),
    .A1(net850),
    .S(net330),
    .X(_01456_));
 sg13g2_mux2_1 _24091_ (.A0(\cpu.genblk1.mmu.r_vtop_d[5][3] ),
    .A1(net998),
    .S(net330),
    .X(_01457_));
 sg13g2_mux2_1 _24092_ (.A0(\cpu.genblk1.mmu.r_vtop_d[5][4] ),
    .A1(net997),
    .S(_06027_),
    .X(_01458_));
 sg13g2_mux2_1 _24093_ (.A0(\cpu.genblk1.mmu.r_vtop_d[5][5] ),
    .A1(net996),
    .S(_06027_),
    .X(_01459_));
 sg13g2_mux2_1 _24094_ (.A0(\cpu.genblk1.mmu.r_vtop_d[5][6] ),
    .A1(net995),
    .S(net330),
    .X(_01460_));
 sg13g2_mux2_1 _24095_ (.A0(\cpu.genblk1.mmu.r_vtop_d[5][7] ),
    .A1(net966),
    .S(net330),
    .X(_01461_));
 sg13g2_mux2_1 _24096_ (.A0(\cpu.genblk1.mmu.r_vtop_d[5][8] ),
    .A1(net552),
    .S(_06026_),
    .X(_01462_));
 sg13g2_mux2_1 _24097_ (.A0(\cpu.genblk1.mmu.r_vtop_d[5][9] ),
    .A1(net493),
    .S(_06026_),
    .X(_01463_));
 sg13g2_nor2_1 _24098_ (.A(net978),
    .B(net659),
    .Y(_06028_));
 sg13g2_and2_1 _24099_ (.A(_05879_),
    .B(_06028_),
    .X(_06029_));
 sg13g2_buf_1 _24100_ (.A(_06029_),
    .X(_06030_));
 sg13g2_nor2b_1 _24101_ (.A(_05890_),
    .B_N(_06030_),
    .Y(_06031_));
 sg13g2_buf_1 _24102_ (.A(_06031_),
    .X(_06032_));
 sg13g2_buf_1 _24103_ (.A(_06032_),
    .X(_06033_));
 sg13g2_mux2_1 _24104_ (.A0(\cpu.genblk1.mmu.r_vtop_d[6][0] ),
    .A1(net401),
    .S(net329),
    .X(_01464_));
 sg13g2_mux2_1 _24105_ (.A0(\cpu.genblk1.mmu.r_vtop_d[6][10] ),
    .A1(net589),
    .S(net329),
    .X(_01465_));
 sg13g2_mux2_1 _24106_ (.A0(\cpu.genblk1.mmu.r_vtop_d[6][11] ),
    .A1(net739),
    .S(net329),
    .X(_01466_));
 sg13g2_mux2_1 _24107_ (.A0(\cpu.genblk1.mmu.r_vtop_d[6][1] ),
    .A1(net668),
    .S(net329),
    .X(_01467_));
 sg13g2_mux2_1 _24108_ (.A0(\cpu.genblk1.mmu.r_vtop_d[6][2] ),
    .A1(net850),
    .S(net329),
    .X(_01468_));
 sg13g2_mux2_1 _24109_ (.A0(\cpu.genblk1.mmu.r_vtop_d[6][3] ),
    .A1(net998),
    .S(net329),
    .X(_01469_));
 sg13g2_mux2_1 _24110_ (.A0(\cpu.genblk1.mmu.r_vtop_d[6][4] ),
    .A1(net997),
    .S(_06033_),
    .X(_01470_));
 sg13g2_mux2_1 _24111_ (.A0(\cpu.genblk1.mmu.r_vtop_d[6][5] ),
    .A1(net996),
    .S(_06033_),
    .X(_01471_));
 sg13g2_mux2_1 _24112_ (.A0(\cpu.genblk1.mmu.r_vtop_d[6][6] ),
    .A1(net995),
    .S(net329),
    .X(_01472_));
 sg13g2_mux2_1 _24113_ (.A0(\cpu.genblk1.mmu.r_vtop_d[6][7] ),
    .A1(net966),
    .S(net329),
    .X(_01473_));
 sg13g2_mux2_1 _24114_ (.A0(\cpu.genblk1.mmu.r_vtop_d[6][8] ),
    .A1(net552),
    .S(_06032_),
    .X(_01474_));
 sg13g2_mux2_1 _24115_ (.A0(\cpu.genblk1.mmu.r_vtop_d[6][9] ),
    .A1(net493),
    .S(_06032_),
    .X(_01475_));
 sg13g2_nor2b_1 _24116_ (.A(_05868_),
    .B_N(_05879_),
    .Y(_06034_));
 sg13g2_buf_2 _24117_ (.A(_06034_),
    .X(_06035_));
 sg13g2_nor2b_1 _24118_ (.A(_05890_),
    .B_N(_06035_),
    .Y(_06036_));
 sg13g2_buf_1 _24119_ (.A(_06036_),
    .X(_06037_));
 sg13g2_buf_1 _24120_ (.A(_06037_),
    .X(_06038_));
 sg13g2_mux2_1 _24121_ (.A0(\cpu.genblk1.mmu.r_vtop_d[7][0] ),
    .A1(_06003_),
    .S(net258),
    .X(_01476_));
 sg13g2_mux2_1 _24122_ (.A0(\cpu.genblk1.mmu.r_vtop_d[7][10] ),
    .A1(net605),
    .S(net258),
    .X(_01477_));
 sg13g2_mux2_1 _24123_ (.A0(\cpu.genblk1.mmu.r_vtop_d[7][11] ),
    .A1(net739),
    .S(net258),
    .X(_01478_));
 sg13g2_mux2_1 _24124_ (.A0(\cpu.genblk1.mmu.r_vtop_d[7][1] ),
    .A1(net668),
    .S(net258),
    .X(_01479_));
 sg13g2_mux2_1 _24125_ (.A0(\cpu.genblk1.mmu.r_vtop_d[7][2] ),
    .A1(net872),
    .S(net258),
    .X(_01480_));
 sg13g2_mux2_1 _24126_ (.A0(\cpu.genblk1.mmu.r_vtop_d[7][3] ),
    .A1(net998),
    .S(_06038_),
    .X(_01481_));
 sg13g2_mux2_1 _24127_ (.A0(\cpu.genblk1.mmu.r_vtop_d[7][4] ),
    .A1(net997),
    .S(_06038_),
    .X(_01482_));
 sg13g2_mux2_1 _24128_ (.A0(\cpu.genblk1.mmu.r_vtop_d[7][5] ),
    .A1(net996),
    .S(net258),
    .X(_01483_));
 sg13g2_mux2_1 _24129_ (.A0(\cpu.genblk1.mmu.r_vtop_d[7][6] ),
    .A1(net995),
    .S(net258),
    .X(_01484_));
 sg13g2_mux2_1 _24130_ (.A0(\cpu.genblk1.mmu.r_vtop_d[7][7] ),
    .A1(net999),
    .S(net258),
    .X(_01485_));
 sg13g2_mux2_1 _24131_ (.A0(\cpu.genblk1.mmu.r_vtop_d[7][8] ),
    .A1(net552),
    .S(_06037_),
    .X(_01486_));
 sg13g2_mux2_1 _24132_ (.A0(\cpu.genblk1.mmu.r_vtop_d[7][9] ),
    .A1(net493),
    .S(_06037_),
    .X(_01487_));
 sg13g2_nor3_1 _24133_ (.A(_05916_),
    .B(_05894_),
    .C(_05929_),
    .Y(_06039_));
 sg13g2_buf_1 _24134_ (.A(_06039_),
    .X(_06040_));
 sg13g2_buf_1 _24135_ (.A(_06040_),
    .X(_06041_));
 sg13g2_mux2_1 _24136_ (.A0(\cpu.genblk1.mmu.r_vtop_d[8][0] ),
    .A1(_06003_),
    .S(net328),
    .X(_01488_));
 sg13g2_mux2_1 _24137_ (.A0(\cpu.genblk1.mmu.r_vtop_d[8][10] ),
    .A1(_03503_),
    .S(net328),
    .X(_01489_));
 sg13g2_mux2_1 _24138_ (.A0(\cpu.genblk1.mmu.r_vtop_d[8][11] ),
    .A1(_03505_),
    .S(net328),
    .X(_01490_));
 sg13g2_mux2_1 _24139_ (.A0(\cpu.genblk1.mmu.r_vtop_d[8][1] ),
    .A1(_02976_),
    .S(_06041_),
    .X(_01491_));
 sg13g2_mux2_1 _24140_ (.A0(\cpu.genblk1.mmu.r_vtop_d[8][2] ),
    .A1(net872),
    .S(net328),
    .X(_01492_));
 sg13g2_mux2_1 _24141_ (.A0(\cpu.genblk1.mmu.r_vtop_d[8][3] ),
    .A1(_02981_),
    .S(net328),
    .X(_01493_));
 sg13g2_mux2_1 _24142_ (.A0(\cpu.genblk1.mmu.r_vtop_d[8][4] ),
    .A1(_02983_),
    .S(net328),
    .X(_01494_));
 sg13g2_mux2_1 _24143_ (.A0(\cpu.genblk1.mmu.r_vtop_d[8][5] ),
    .A1(net996),
    .S(_06041_),
    .X(_01495_));
 sg13g2_mux2_1 _24144_ (.A0(\cpu.genblk1.mmu.r_vtop_d[8][6] ),
    .A1(_02987_),
    .S(net328),
    .X(_01496_));
 sg13g2_mux2_1 _24145_ (.A0(\cpu.genblk1.mmu.r_vtop_d[8][7] ),
    .A1(net999),
    .S(net328),
    .X(_01497_));
 sg13g2_mux2_1 _24146_ (.A0(\cpu.genblk1.mmu.r_vtop_d[8][8] ),
    .A1(_03499_),
    .S(_06040_),
    .X(_01498_));
 sg13g2_mux2_1 _24147_ (.A0(\cpu.genblk1.mmu.r_vtop_d[8][9] ),
    .A1(_03501_),
    .S(_06040_),
    .X(_01499_));
 sg13g2_nor3_1 _24148_ (.A(_05870_),
    .B(_05894_),
    .C(_05911_),
    .Y(_06042_));
 sg13g2_buf_1 _24149_ (.A(_06042_),
    .X(_06043_));
 sg13g2_buf_1 _24150_ (.A(_06043_),
    .X(_06044_));
 sg13g2_mux2_1 _24151_ (.A0(\cpu.genblk1.mmu.r_vtop_d[9][0] ),
    .A1(net452),
    .S(net257),
    .X(_01500_));
 sg13g2_mux2_1 _24152_ (.A0(\cpu.genblk1.mmu.r_vtop_d[9][10] ),
    .A1(_03503_),
    .S(net257),
    .X(_01501_));
 sg13g2_mux2_1 _24153_ (.A0(\cpu.genblk1.mmu.r_vtop_d[9][11] ),
    .A1(_03505_),
    .S(net257),
    .X(_01502_));
 sg13g2_mux2_1 _24154_ (.A0(\cpu.genblk1.mmu.r_vtop_d[9][1] ),
    .A1(_02976_),
    .S(_06044_),
    .X(_01503_));
 sg13g2_mux2_1 _24155_ (.A0(\cpu.genblk1.mmu.r_vtop_d[9][2] ),
    .A1(_02960_),
    .S(net257),
    .X(_01504_));
 sg13g2_mux2_1 _24156_ (.A0(\cpu.genblk1.mmu.r_vtop_d[9][3] ),
    .A1(_02981_),
    .S(net257),
    .X(_01505_));
 sg13g2_mux2_1 _24157_ (.A0(\cpu.genblk1.mmu.r_vtop_d[9][4] ),
    .A1(_02983_),
    .S(net257),
    .X(_01506_));
 sg13g2_mux2_1 _24158_ (.A0(\cpu.genblk1.mmu.r_vtop_d[9][5] ),
    .A1(net996),
    .S(_06044_),
    .X(_01507_));
 sg13g2_mux2_1 _24159_ (.A0(\cpu.genblk1.mmu.r_vtop_d[9][6] ),
    .A1(_02987_),
    .S(net257),
    .X(_01508_));
 sg13g2_mux2_1 _24160_ (.A0(\cpu.genblk1.mmu.r_vtop_d[9][7] ),
    .A1(_02973_),
    .S(net257),
    .X(_01509_));
 sg13g2_mux2_1 _24161_ (.A0(\cpu.genblk1.mmu.r_vtop_d[9][8] ),
    .A1(net552),
    .S(_06043_),
    .X(_01510_));
 sg13g2_mux2_1 _24162_ (.A0(\cpu.genblk1.mmu.r_vtop_d[9][9] ),
    .A1(_03501_),
    .S(_06043_),
    .X(_01511_));
 sg13g2_and2_1 _24163_ (.A(_05877_),
    .B(_05879_),
    .X(_06045_));
 sg13g2_buf_1 _24164_ (.A(_06045_),
    .X(_06046_));
 sg13g2_and3_1 _24165_ (.X(_06047_),
    .A(net1145),
    .B(_10604_),
    .C(_05828_));
 sg13g2_buf_1 _24166_ (.A(_06047_),
    .X(_06048_));
 sg13g2_and2_1 _24167_ (.A(_05845_),
    .B(_06048_),
    .X(_06049_));
 sg13g2_buf_1 _24168_ (.A(_06049_),
    .X(_06050_));
 sg13g2_nand2_1 _24169_ (.Y(_06051_),
    .A(_06046_),
    .B(_06050_));
 sg13g2_buf_1 _24170_ (.A(_06051_),
    .X(_06052_));
 sg13g2_buf_1 _24171_ (.A(net327),
    .X(_06053_));
 sg13g2_nand2_1 _24172_ (.Y(_06054_),
    .A(\cpu.genblk1.mmu.r_vtop_i[0][0] ),
    .B(net327));
 sg13g2_o21ai_1 _24173_ (.B1(_06054_),
    .Y(_01512_),
    .A1(net599),
    .A2(net256));
 sg13g2_mux2_1 _24174_ (.A0(net541),
    .A1(\cpu.genblk1.mmu.r_vtop_i[0][10] ),
    .S(net256),
    .X(_01513_));
 sg13g2_nand2_1 _24175_ (.Y(_06055_),
    .A(\cpu.genblk1.mmu.r_vtop_i[0][11] ),
    .B(_06052_));
 sg13g2_o21ai_1 _24176_ (.B1(_06055_),
    .Y(_01514_),
    .A1(net601),
    .A2(net256));
 sg13g2_nand2_1 _24177_ (.Y(_06056_),
    .A(\cpu.genblk1.mmu.r_vtop_i[0][1] ),
    .B(net327));
 sg13g2_o21ai_1 _24178_ (.B1(_06056_),
    .Y(_01515_),
    .A1(net754),
    .A2(net256));
 sg13g2_mux2_1 _24179_ (.A0(net753),
    .A1(\cpu.genblk1.mmu.r_vtop_i[0][2] ),
    .S(net256),
    .X(_01516_));
 sg13g2_nand2_1 _24180_ (.Y(_06057_),
    .A(\cpu.genblk1.mmu.r_vtop_i[0][3] ),
    .B(net327));
 sg13g2_o21ai_1 _24181_ (.B1(_06057_),
    .Y(_01517_),
    .A1(net752),
    .A2(net256));
 sg13g2_nand2_1 _24182_ (.Y(_06058_),
    .A(\cpu.genblk1.mmu.r_vtop_i[0][4] ),
    .B(_06052_));
 sg13g2_o21ai_1 _24183_ (.B1(_06058_),
    .Y(_01518_),
    .A1(net870),
    .A2(_06053_));
 sg13g2_nand2_1 _24184_ (.Y(_06059_),
    .A(\cpu.genblk1.mmu.r_vtop_i[0][5] ),
    .B(net327));
 sg13g2_o21ai_1 _24185_ (.B1(_06059_),
    .Y(_01519_),
    .A1(net751),
    .A2(_06053_));
 sg13g2_nand2_1 _24186_ (.Y(_06060_),
    .A(\cpu.genblk1.mmu.r_vtop_i[0][6] ),
    .B(net327));
 sg13g2_o21ai_1 _24187_ (.B1(_06060_),
    .Y(_01520_),
    .A1(net750),
    .A2(net256));
 sg13g2_mux2_1 _24188_ (.A0(net868),
    .A1(\cpu.genblk1.mmu.r_vtop_i[0][7] ),
    .S(net256),
    .X(_01521_));
 sg13g2_mux2_1 _24189_ (.A0(net488),
    .A1(\cpu.genblk1.mmu.r_vtop_i[0][8] ),
    .S(net327),
    .X(_01522_));
 sg13g2_mux2_1 _24190_ (.A0(_03830_),
    .A1(\cpu.genblk1.mmu.r_vtop_i[0][9] ),
    .S(net327),
    .X(_01523_));
 sg13g2_buf_1 _24191_ (.A(_06048_),
    .X(_06061_));
 sg13g2_nand2_1 _24192_ (.Y(_06062_),
    .A(_05895_),
    .B(net477));
 sg13g2_buf_1 _24193_ (.A(_06062_),
    .X(_06063_));
 sg13g2_buf_1 _24194_ (.A(net400),
    .X(_06064_));
 sg13g2_nand2_1 _24195_ (.Y(_06065_),
    .A(\cpu.genblk1.mmu.r_vtop_i[10][0] ),
    .B(net400));
 sg13g2_o21ai_1 _24196_ (.B1(_06065_),
    .Y(_01524_),
    .A1(net599),
    .A2(net326));
 sg13g2_mux2_1 _24197_ (.A0(net541),
    .A1(\cpu.genblk1.mmu.r_vtop_i[10][10] ),
    .S(net326),
    .X(_01525_));
 sg13g2_nand2_1 _24198_ (.Y(_06066_),
    .A(\cpu.genblk1.mmu.r_vtop_i[10][11] ),
    .B(_06063_));
 sg13g2_o21ai_1 _24199_ (.B1(_06066_),
    .Y(_01526_),
    .A1(net601),
    .A2(net326));
 sg13g2_nand2_1 _24200_ (.Y(_06067_),
    .A(\cpu.genblk1.mmu.r_vtop_i[10][1] ),
    .B(net400));
 sg13g2_o21ai_1 _24201_ (.B1(_06067_),
    .Y(_01527_),
    .A1(net754),
    .A2(_06064_));
 sg13g2_mux2_1 _24202_ (.A0(net753),
    .A1(\cpu.genblk1.mmu.r_vtop_i[10][2] ),
    .S(net326),
    .X(_01528_));
 sg13g2_nand2_1 _24203_ (.Y(_06068_),
    .A(\cpu.genblk1.mmu.r_vtop_i[10][3] ),
    .B(net400));
 sg13g2_o21ai_1 _24204_ (.B1(_06068_),
    .Y(_01529_),
    .A1(net752),
    .A2(net326));
 sg13g2_nand2_1 _24205_ (.Y(_06069_),
    .A(\cpu.genblk1.mmu.r_vtop_i[10][4] ),
    .B(_06063_));
 sg13g2_o21ai_1 _24206_ (.B1(_06069_),
    .Y(_01530_),
    .A1(net870),
    .A2(net326));
 sg13g2_nand2_1 _24207_ (.Y(_06070_),
    .A(\cpu.genblk1.mmu.r_vtop_i[10][5] ),
    .B(net400));
 sg13g2_o21ai_1 _24208_ (.B1(_06070_),
    .Y(_01531_),
    .A1(net751),
    .A2(_06064_));
 sg13g2_nand2_1 _24209_ (.Y(_06071_),
    .A(\cpu.genblk1.mmu.r_vtop_i[10][6] ),
    .B(net400));
 sg13g2_o21ai_1 _24210_ (.B1(_06071_),
    .Y(_01532_),
    .A1(net750),
    .A2(net326));
 sg13g2_mux2_1 _24211_ (.A0(net868),
    .A1(\cpu.genblk1.mmu.r_vtop_i[10][7] ),
    .S(net326),
    .X(_01533_));
 sg13g2_mux2_1 _24212_ (.A0(net488),
    .A1(\cpu.genblk1.mmu.r_vtop_i[10][8] ),
    .S(net400),
    .X(_01534_));
 sg13g2_mux2_1 _24213_ (.A0(_03830_),
    .A1(\cpu.genblk1.mmu.r_vtop_i[10][9] ),
    .S(net400),
    .X(_01535_));
 sg13g2_nand2_1 _24214_ (.Y(_06072_),
    .A(_05900_),
    .B(net477));
 sg13g2_buf_1 _24215_ (.A(_06072_),
    .X(_06073_));
 sg13g2_buf_1 _24216_ (.A(net399),
    .X(_06074_));
 sg13g2_nand2_1 _24217_ (.Y(_06075_),
    .A(\cpu.genblk1.mmu.r_vtop_i[11][0] ),
    .B(net399));
 sg13g2_o21ai_1 _24218_ (.B1(_06075_),
    .Y(_01536_),
    .A1(net599),
    .A2(net325));
 sg13g2_mux2_1 _24219_ (.A0(net541),
    .A1(\cpu.genblk1.mmu.r_vtop_i[11][10] ),
    .S(net325),
    .X(_01537_));
 sg13g2_nand2_1 _24220_ (.Y(_06076_),
    .A(\cpu.genblk1.mmu.r_vtop_i[11][11] ),
    .B(_06073_));
 sg13g2_o21ai_1 _24221_ (.B1(_06076_),
    .Y(_01538_),
    .A1(net601),
    .A2(net325));
 sg13g2_nand2_1 _24222_ (.Y(_06077_),
    .A(\cpu.genblk1.mmu.r_vtop_i[11][1] ),
    .B(net399));
 sg13g2_o21ai_1 _24223_ (.B1(_06077_),
    .Y(_01539_),
    .A1(net754),
    .A2(net325));
 sg13g2_mux2_1 _24224_ (.A0(net753),
    .A1(\cpu.genblk1.mmu.r_vtop_i[11][2] ),
    .S(net325),
    .X(_01540_));
 sg13g2_nand2_1 _24225_ (.Y(_06078_),
    .A(\cpu.genblk1.mmu.r_vtop_i[11][3] ),
    .B(net399));
 sg13g2_o21ai_1 _24226_ (.B1(_06078_),
    .Y(_01541_),
    .A1(net752),
    .A2(net325));
 sg13g2_nand2_1 _24227_ (.Y(_06079_),
    .A(\cpu.genblk1.mmu.r_vtop_i[11][4] ),
    .B(_06073_));
 sg13g2_o21ai_1 _24228_ (.B1(_06079_),
    .Y(_01542_),
    .A1(net870),
    .A2(_06074_));
 sg13g2_nand2_1 _24229_ (.Y(_06080_),
    .A(\cpu.genblk1.mmu.r_vtop_i[11][5] ),
    .B(net399));
 sg13g2_o21ai_1 _24230_ (.B1(_06080_),
    .Y(_01543_),
    .A1(net751),
    .A2(_06074_));
 sg13g2_nand2_1 _24231_ (.Y(_06081_),
    .A(\cpu.genblk1.mmu.r_vtop_i[11][6] ),
    .B(net399));
 sg13g2_o21ai_1 _24232_ (.B1(_06081_),
    .Y(_01544_),
    .A1(net750),
    .A2(net325));
 sg13g2_mux2_1 _24233_ (.A0(net868),
    .A1(\cpu.genblk1.mmu.r_vtop_i[11][7] ),
    .S(net325),
    .X(_01545_));
 sg13g2_mux2_1 _24234_ (.A0(_03829_),
    .A1(\cpu.genblk1.mmu.r_vtop_i[11][8] ),
    .S(net399),
    .X(_01546_));
 sg13g2_mux2_1 _24235_ (.A0(net451),
    .A1(\cpu.genblk1.mmu.r_vtop_i[11][9] ),
    .S(net399),
    .X(_01547_));
 sg13g2_nor2_1 _24236_ (.A(_05877_),
    .B(_05894_),
    .Y(_06082_));
 sg13g2_nand2_1 _24237_ (.Y(_06083_),
    .A(_06082_),
    .B(_06050_));
 sg13g2_buf_1 _24238_ (.A(_06083_),
    .X(_06084_));
 sg13g2_buf_1 _24239_ (.A(net324),
    .X(_06085_));
 sg13g2_nand2_1 _24240_ (.Y(_06086_),
    .A(\cpu.genblk1.mmu.r_vtop_i[12][0] ),
    .B(net324));
 sg13g2_o21ai_1 _24241_ (.B1(_06086_),
    .Y(_01548_),
    .A1(net599),
    .A2(net255));
 sg13g2_mux2_1 _24242_ (.A0(net541),
    .A1(\cpu.genblk1.mmu.r_vtop_i[12][10] ),
    .S(net255),
    .X(_01549_));
 sg13g2_nand2_1 _24243_ (.Y(_06087_),
    .A(\cpu.genblk1.mmu.r_vtop_i[12][11] ),
    .B(net324));
 sg13g2_o21ai_1 _24244_ (.B1(_06087_),
    .Y(_01550_),
    .A1(net601),
    .A2(_06085_));
 sg13g2_nand2_1 _24245_ (.Y(_06088_),
    .A(\cpu.genblk1.mmu.r_vtop_i[12][1] ),
    .B(net324));
 sg13g2_o21ai_1 _24246_ (.B1(_06088_),
    .Y(_01551_),
    .A1(net754),
    .A2(net255));
 sg13g2_mux2_1 _24247_ (.A0(net753),
    .A1(\cpu.genblk1.mmu.r_vtop_i[12][2] ),
    .S(net255),
    .X(_01552_));
 sg13g2_nand2_1 _24248_ (.Y(_06089_),
    .A(\cpu.genblk1.mmu.r_vtop_i[12][3] ),
    .B(net324));
 sg13g2_o21ai_1 _24249_ (.B1(_06089_),
    .Y(_01553_),
    .A1(net752),
    .A2(net255));
 sg13g2_nand2_1 _24250_ (.Y(_06090_),
    .A(\cpu.genblk1.mmu.r_vtop_i[12][4] ),
    .B(net324));
 sg13g2_o21ai_1 _24251_ (.B1(_06090_),
    .Y(_01554_),
    .A1(net870),
    .A2(net255));
 sg13g2_nand2_1 _24252_ (.Y(_06091_),
    .A(\cpu.genblk1.mmu.r_vtop_i[12][5] ),
    .B(net324));
 sg13g2_o21ai_1 _24253_ (.B1(_06091_),
    .Y(_01555_),
    .A1(net751),
    .A2(net255));
 sg13g2_nand2_1 _24254_ (.Y(_06092_),
    .A(\cpu.genblk1.mmu.r_vtop_i[12][6] ),
    .B(net324));
 sg13g2_o21ai_1 _24255_ (.B1(_06092_),
    .Y(_01556_),
    .A1(net750),
    .A2(_06085_));
 sg13g2_mux2_1 _24256_ (.A0(net868),
    .A1(\cpu.genblk1.mmu.r_vtop_i[12][7] ),
    .S(net255),
    .X(_01557_));
 sg13g2_mux2_1 _24257_ (.A0(net488),
    .A1(\cpu.genblk1.mmu.r_vtop_i[12][8] ),
    .S(_06084_),
    .X(_01558_));
 sg13g2_mux2_1 _24258_ (.A0(net451),
    .A1(\cpu.genblk1.mmu.r_vtop_i[12][9] ),
    .S(_06084_),
    .X(_01559_));
 sg13g2_nor2b_1 _24259_ (.A(_05909_),
    .B_N(_06048_),
    .Y(_06093_));
 sg13g2_buf_2 _24260_ (.A(_06093_),
    .X(_06094_));
 sg13g2_nand2_1 _24261_ (.Y(_06095_),
    .A(_06082_),
    .B(_06094_));
 sg13g2_buf_1 _24262_ (.A(_06095_),
    .X(_06096_));
 sg13g2_buf_1 _24263_ (.A(net323),
    .X(_06097_));
 sg13g2_nand2_1 _24264_ (.Y(_06098_),
    .A(\cpu.genblk1.mmu.r_vtop_i[13][0] ),
    .B(net323));
 sg13g2_o21ai_1 _24265_ (.B1(_06098_),
    .Y(_01560_),
    .A1(net599),
    .A2(net254));
 sg13g2_mux2_1 _24266_ (.A0(net541),
    .A1(\cpu.genblk1.mmu.r_vtop_i[13][10] ),
    .S(net254),
    .X(_01561_));
 sg13g2_nand2_1 _24267_ (.Y(_06099_),
    .A(\cpu.genblk1.mmu.r_vtop_i[13][11] ),
    .B(net323));
 sg13g2_o21ai_1 _24268_ (.B1(_06099_),
    .Y(_01562_),
    .A1(net601),
    .A2(_06097_));
 sg13g2_nand2_1 _24269_ (.Y(_06100_),
    .A(\cpu.genblk1.mmu.r_vtop_i[13][1] ),
    .B(net323));
 sg13g2_o21ai_1 _24270_ (.B1(_06100_),
    .Y(_01563_),
    .A1(net754),
    .A2(net254));
 sg13g2_mux2_1 _24271_ (.A0(net753),
    .A1(\cpu.genblk1.mmu.r_vtop_i[13][2] ),
    .S(net254),
    .X(_01564_));
 sg13g2_nand2_1 _24272_ (.Y(_06101_),
    .A(\cpu.genblk1.mmu.r_vtop_i[13][3] ),
    .B(net323));
 sg13g2_o21ai_1 _24273_ (.B1(_06101_),
    .Y(_01565_),
    .A1(net752),
    .A2(net254));
 sg13g2_nand2_1 _24274_ (.Y(_06102_),
    .A(\cpu.genblk1.mmu.r_vtop_i[13][4] ),
    .B(net323));
 sg13g2_o21ai_1 _24275_ (.B1(_06102_),
    .Y(_01566_),
    .A1(net870),
    .A2(net254));
 sg13g2_nand2_1 _24276_ (.Y(_06103_),
    .A(\cpu.genblk1.mmu.r_vtop_i[13][5] ),
    .B(net323));
 sg13g2_o21ai_1 _24277_ (.B1(_06103_),
    .Y(_01567_),
    .A1(net751),
    .A2(net254));
 sg13g2_nand2_1 _24278_ (.Y(_06104_),
    .A(\cpu.genblk1.mmu.r_vtop_i[13][6] ),
    .B(net323));
 sg13g2_o21ai_1 _24279_ (.B1(_06104_),
    .Y(_01568_),
    .A1(net750),
    .A2(_06097_));
 sg13g2_mux2_1 _24280_ (.A0(net868),
    .A1(\cpu.genblk1.mmu.r_vtop_i[13][7] ),
    .S(net254),
    .X(_01569_));
 sg13g2_mux2_1 _24281_ (.A0(net488),
    .A1(\cpu.genblk1.mmu.r_vtop_i[13][8] ),
    .S(_06096_),
    .X(_01570_));
 sg13g2_mux2_1 _24282_ (.A0(net451),
    .A1(\cpu.genblk1.mmu.r_vtop_i[13][9] ),
    .S(_06096_),
    .X(_01571_));
 sg13g2_nor2_1 _24283_ (.A(net980),
    .B(_05842_),
    .Y(_06105_));
 sg13g2_nand3_1 _24284_ (.B(_06082_),
    .C(_06061_),
    .A(_06105_),
    .Y(_06106_));
 sg13g2_buf_1 _24285_ (.A(_06106_),
    .X(_06107_));
 sg13g2_buf_1 _24286_ (.A(net398),
    .X(_06108_));
 sg13g2_nand2_1 _24287_ (.Y(_06109_),
    .A(\cpu.genblk1.mmu.r_vtop_i[14][0] ),
    .B(net398));
 sg13g2_o21ai_1 _24288_ (.B1(_06109_),
    .Y(_01572_),
    .A1(_03839_),
    .A2(net322));
 sg13g2_mux2_1 _24289_ (.A0(_03831_),
    .A1(\cpu.genblk1.mmu.r_vtop_i[14][10] ),
    .S(net322),
    .X(_01573_));
 sg13g2_nand2_1 _24290_ (.Y(_06110_),
    .A(\cpu.genblk1.mmu.r_vtop_i[14][11] ),
    .B(net398));
 sg13g2_o21ai_1 _24291_ (.B1(_06110_),
    .Y(_01574_),
    .A1(net601),
    .A2(_06108_));
 sg13g2_nand2_1 _24292_ (.Y(_06111_),
    .A(\cpu.genblk1.mmu.r_vtop_i[14][1] ),
    .B(net398));
 sg13g2_o21ai_1 _24293_ (.B1(_06111_),
    .Y(_01575_),
    .A1(net754),
    .A2(net322));
 sg13g2_mux2_1 _24294_ (.A0(net753),
    .A1(\cpu.genblk1.mmu.r_vtop_i[14][2] ),
    .S(net322),
    .X(_01576_));
 sg13g2_nand2_1 _24295_ (.Y(_06112_),
    .A(\cpu.genblk1.mmu.r_vtop_i[14][3] ),
    .B(net398));
 sg13g2_o21ai_1 _24296_ (.B1(_06112_),
    .Y(_01577_),
    .A1(net752),
    .A2(net322));
 sg13g2_nand2_1 _24297_ (.Y(_06113_),
    .A(\cpu.genblk1.mmu.r_vtop_i[14][4] ),
    .B(net398));
 sg13g2_o21ai_1 _24298_ (.B1(_06113_),
    .Y(_01578_),
    .A1(net870),
    .A2(_06108_));
 sg13g2_nand2_1 _24299_ (.Y(_06114_),
    .A(\cpu.genblk1.mmu.r_vtop_i[14][5] ),
    .B(net398));
 sg13g2_o21ai_1 _24300_ (.B1(_06114_),
    .Y(_01579_),
    .A1(net751),
    .A2(net322));
 sg13g2_nand2_1 _24301_ (.Y(_06115_),
    .A(\cpu.genblk1.mmu.r_vtop_i[14][6] ),
    .B(net398));
 sg13g2_o21ai_1 _24302_ (.B1(_06115_),
    .Y(_01580_),
    .A1(net750),
    .A2(net322));
 sg13g2_mux2_1 _24303_ (.A0(net868),
    .A1(\cpu.genblk1.mmu.r_vtop_i[14][7] ),
    .S(net322),
    .X(_01581_));
 sg13g2_mux2_1 _24304_ (.A0(_03829_),
    .A1(\cpu.genblk1.mmu.r_vtop_i[14][8] ),
    .S(_06107_),
    .X(_01582_));
 sg13g2_mux2_1 _24305_ (.A0(net451),
    .A1(\cpu.genblk1.mmu.r_vtop_i[14][9] ),
    .S(_06107_),
    .X(_01583_));
 sg13g2_buf_1 _24306_ (.A(_06048_),
    .X(_06116_));
 sg13g2_nand3_1 _24307_ (.B(_06082_),
    .C(_06116_),
    .A(_05844_),
    .Y(_06117_));
 sg13g2_buf_1 _24308_ (.A(_06117_),
    .X(_06118_));
 sg13g2_buf_1 _24309_ (.A(net397),
    .X(_06119_));
 sg13g2_nand2_1 _24310_ (.Y(_06120_),
    .A(\cpu.genblk1.mmu.r_vtop_i[15][0] ),
    .B(net397));
 sg13g2_o21ai_1 _24311_ (.B1(_06120_),
    .Y(_01584_),
    .A1(_03839_),
    .A2(net321));
 sg13g2_mux2_1 _24312_ (.A0(_03831_),
    .A1(\cpu.genblk1.mmu.r_vtop_i[15][10] ),
    .S(net321),
    .X(_01585_));
 sg13g2_nand2_1 _24313_ (.Y(_06121_),
    .A(\cpu.genblk1.mmu.r_vtop_i[15][11] ),
    .B(net397));
 sg13g2_o21ai_1 _24314_ (.B1(_06121_),
    .Y(_01586_),
    .A1(_03832_),
    .A2(_06119_));
 sg13g2_nand2_1 _24315_ (.Y(_06122_),
    .A(\cpu.genblk1.mmu.r_vtop_i[15][1] ),
    .B(net397));
 sg13g2_o21ai_1 _24316_ (.B1(_06122_),
    .Y(_01587_),
    .A1(net754),
    .A2(net321));
 sg13g2_mux2_1 _24317_ (.A0(net753),
    .A1(\cpu.genblk1.mmu.r_vtop_i[15][2] ),
    .S(net321),
    .X(_01588_));
 sg13g2_nand2_1 _24318_ (.Y(_06123_),
    .A(\cpu.genblk1.mmu.r_vtop_i[15][3] ),
    .B(net397));
 sg13g2_o21ai_1 _24319_ (.B1(_06123_),
    .Y(_01589_),
    .A1(net752),
    .A2(net321));
 sg13g2_nand2_1 _24320_ (.Y(_06124_),
    .A(\cpu.genblk1.mmu.r_vtop_i[15][4] ),
    .B(net397));
 sg13g2_o21ai_1 _24321_ (.B1(_06124_),
    .Y(_01590_),
    .A1(net870),
    .A2(_06119_));
 sg13g2_nand2_1 _24322_ (.Y(_06125_),
    .A(\cpu.genblk1.mmu.r_vtop_i[15][5] ),
    .B(net397));
 sg13g2_o21ai_1 _24323_ (.B1(_06125_),
    .Y(_01591_),
    .A1(net751),
    .A2(net321));
 sg13g2_nand2_1 _24324_ (.Y(_06126_),
    .A(\cpu.genblk1.mmu.r_vtop_i[15][6] ),
    .B(net397));
 sg13g2_o21ai_1 _24325_ (.B1(_06126_),
    .Y(_01592_),
    .A1(net750),
    .A2(net321));
 sg13g2_mux2_1 _24326_ (.A0(net868),
    .A1(\cpu.genblk1.mmu.r_vtop_i[15][7] ),
    .S(net321),
    .X(_01593_));
 sg13g2_mux2_1 _24327_ (.A0(net488),
    .A1(\cpu.genblk1.mmu.r_vtop_i[15][8] ),
    .S(_06118_),
    .X(_01594_));
 sg13g2_mux2_1 _24328_ (.A0(net451),
    .A1(\cpu.genblk1.mmu.r_vtop_i[15][9] ),
    .S(_06118_),
    .X(_01595_));
 sg13g2_buf_1 _24329_ (.A(net1121),
    .X(_06127_));
 sg13g2_nor3_2 _24330_ (.A(net980),
    .B(net979),
    .C(net976),
    .Y(_06128_));
 sg13g2_nand4_1 _24331_ (.B(net1044),
    .C(_06128_),
    .A(net965),
    .Y(_06129_),
    .D(net476));
 sg13g2_buf_1 _24332_ (.A(_06129_),
    .X(_06130_));
 sg13g2_buf_1 _24333_ (.A(net396),
    .X(_06131_));
 sg13g2_nand2_1 _24334_ (.Y(_06132_),
    .A(\cpu.genblk1.mmu.r_vtop_i[16][0] ),
    .B(net396));
 sg13g2_o21ai_1 _24335_ (.B1(_06132_),
    .Y(_01596_),
    .A1(net599),
    .A2(net320));
 sg13g2_mux2_1 _24336_ (.A0(net541),
    .A1(\cpu.genblk1.mmu.r_vtop_i[16][10] ),
    .S(net320),
    .X(_01597_));
 sg13g2_nand2_1 _24337_ (.Y(_06133_),
    .A(\cpu.genblk1.mmu.r_vtop_i[16][11] ),
    .B(net396));
 sg13g2_o21ai_1 _24338_ (.B1(_06133_),
    .Y(_01598_),
    .A1(net601),
    .A2(net320));
 sg13g2_buf_1 _24339_ (.A(net873),
    .X(_06134_));
 sg13g2_nand2_1 _24340_ (.Y(_06135_),
    .A(\cpu.genblk1.mmu.r_vtop_i[16][1] ),
    .B(net396));
 sg13g2_o21ai_1 _24341_ (.B1(_06135_),
    .Y(_01599_),
    .A1(net738),
    .A2(_06131_));
 sg13g2_buf_1 _24342_ (.A(net872),
    .X(_06136_));
 sg13g2_mux2_1 _24343_ (.A0(net737),
    .A1(\cpu.genblk1.mmu.r_vtop_i[16][2] ),
    .S(net320),
    .X(_01600_));
 sg13g2_buf_1 _24344_ (.A(net871),
    .X(_06137_));
 sg13g2_nand2_1 _24345_ (.Y(_06138_),
    .A(\cpu.genblk1.mmu.r_vtop_i[16][3] ),
    .B(net396));
 sg13g2_o21ai_1 _24346_ (.B1(_06138_),
    .Y(_01601_),
    .A1(net736),
    .A2(net320));
 sg13g2_buf_1 _24347_ (.A(net1037),
    .X(_06139_));
 sg13g2_nand2_1 _24348_ (.Y(_06140_),
    .A(\cpu.genblk1.mmu.r_vtop_i[16][4] ),
    .B(net396));
 sg13g2_o21ai_1 _24349_ (.B1(_06140_),
    .Y(_01602_),
    .A1(net849),
    .A2(_06131_));
 sg13g2_buf_1 _24350_ (.A(net869),
    .X(_06141_));
 sg13g2_nand2_1 _24351_ (.Y(_06142_),
    .A(\cpu.genblk1.mmu.r_vtop_i[16][5] ),
    .B(net396));
 sg13g2_o21ai_1 _24352_ (.B1(_06142_),
    .Y(_01603_),
    .A1(net735),
    .A2(net320));
 sg13g2_buf_1 _24353_ (.A(net889),
    .X(_06143_));
 sg13g2_nand2_1 _24354_ (.Y(_06144_),
    .A(\cpu.genblk1.mmu.r_vtop_i[16][6] ),
    .B(net396));
 sg13g2_o21ai_1 _24355_ (.B1(_06144_),
    .Y(_01604_),
    .A1(net734),
    .A2(net320));
 sg13g2_buf_1 _24356_ (.A(net999),
    .X(_06145_));
 sg13g2_mux2_1 _24357_ (.A0(net848),
    .A1(\cpu.genblk1.mmu.r_vtop_i[16][7] ),
    .S(net320),
    .X(_01605_));
 sg13g2_mux2_1 _24358_ (.A0(net488),
    .A1(\cpu.genblk1.mmu.r_vtop_i[16][8] ),
    .S(_06130_),
    .X(_01606_));
 sg13g2_mux2_1 _24359_ (.A0(net451),
    .A1(\cpu.genblk1.mmu.r_vtop_i[16][9] ),
    .S(_06130_),
    .X(_01607_));
 sg13g2_nand4_1 _24360_ (.B(net978),
    .C(net1044),
    .A(net965),
    .Y(_06146_),
    .D(_06094_));
 sg13g2_buf_1 _24361_ (.A(_06146_),
    .X(_06147_));
 sg13g2_buf_1 _24362_ (.A(net319),
    .X(_06148_));
 sg13g2_nand2_1 _24363_ (.Y(_06149_),
    .A(\cpu.genblk1.mmu.r_vtop_i[17][0] ),
    .B(net319));
 sg13g2_o21ai_1 _24364_ (.B1(_06149_),
    .Y(_01608_),
    .A1(net599),
    .A2(net253));
 sg13g2_mux2_1 _24365_ (.A0(net541),
    .A1(\cpu.genblk1.mmu.r_vtop_i[17][10] ),
    .S(net253),
    .X(_01609_));
 sg13g2_nand2_1 _24366_ (.Y(_06150_),
    .A(\cpu.genblk1.mmu.r_vtop_i[17][11] ),
    .B(net319));
 sg13g2_o21ai_1 _24367_ (.B1(_06150_),
    .Y(_01610_),
    .A1(net601),
    .A2(net253));
 sg13g2_nand2_1 _24368_ (.Y(_06151_),
    .A(\cpu.genblk1.mmu.r_vtop_i[17][1] ),
    .B(net319));
 sg13g2_o21ai_1 _24369_ (.B1(_06151_),
    .Y(_01611_),
    .A1(net738),
    .A2(_06148_));
 sg13g2_mux2_1 _24370_ (.A0(net737),
    .A1(\cpu.genblk1.mmu.r_vtop_i[17][2] ),
    .S(net253),
    .X(_01612_));
 sg13g2_nand2_1 _24371_ (.Y(_06152_),
    .A(\cpu.genblk1.mmu.r_vtop_i[17][3] ),
    .B(net319));
 sg13g2_o21ai_1 _24372_ (.B1(_06152_),
    .Y(_01613_),
    .A1(net736),
    .A2(net253));
 sg13g2_nand2_1 _24373_ (.Y(_06153_),
    .A(\cpu.genblk1.mmu.r_vtop_i[17][4] ),
    .B(net319));
 sg13g2_o21ai_1 _24374_ (.B1(_06153_),
    .Y(_01614_),
    .A1(_06139_),
    .A2(_06148_));
 sg13g2_nand2_1 _24375_ (.Y(_06154_),
    .A(\cpu.genblk1.mmu.r_vtop_i[17][5] ),
    .B(net319));
 sg13g2_o21ai_1 _24376_ (.B1(_06154_),
    .Y(_01615_),
    .A1(net735),
    .A2(net253));
 sg13g2_nand2_1 _24377_ (.Y(_06155_),
    .A(\cpu.genblk1.mmu.r_vtop_i[17][6] ),
    .B(net319));
 sg13g2_o21ai_1 _24378_ (.B1(_06155_),
    .Y(_01616_),
    .A1(_06143_),
    .A2(net253));
 sg13g2_mux2_1 _24379_ (.A0(net848),
    .A1(\cpu.genblk1.mmu.r_vtop_i[17][7] ),
    .S(net253),
    .X(_01617_));
 sg13g2_mux2_1 _24380_ (.A0(net488),
    .A1(\cpu.genblk1.mmu.r_vtop_i[17][8] ),
    .S(_06147_),
    .X(_01618_));
 sg13g2_mux2_1 _24381_ (.A0(net451),
    .A1(\cpu.genblk1.mmu.r_vtop_i[17][9] ),
    .S(_06147_),
    .X(_01619_));
 sg13g2_buf_1 _24382_ (.A(net666),
    .X(_06156_));
 sg13g2_nand2_1 _24383_ (.Y(_06157_),
    .A(_05939_),
    .B(net477));
 sg13g2_buf_1 _24384_ (.A(_06157_),
    .X(_06158_));
 sg13g2_buf_1 _24385_ (.A(net395),
    .X(_06159_));
 sg13g2_nand2_1 _24386_ (.Y(_06160_),
    .A(\cpu.genblk1.mmu.r_vtop_i[18][0] ),
    .B(net395));
 sg13g2_o21ai_1 _24387_ (.B1(_06160_),
    .Y(_01620_),
    .A1(net588),
    .A2(net318));
 sg13g2_buf_1 _24388_ (.A(net605),
    .X(_06161_));
 sg13g2_mux2_1 _24389_ (.A0(net526),
    .A1(\cpu.genblk1.mmu.r_vtop_i[18][10] ),
    .S(net318),
    .X(_01621_));
 sg13g2_buf_1 _24390_ (.A(net699),
    .X(_06162_));
 sg13g2_nand2_1 _24391_ (.Y(_06163_),
    .A(\cpu.genblk1.mmu.r_vtop_i[18][11] ),
    .B(net395));
 sg13g2_o21ai_1 _24392_ (.B1(_06163_),
    .Y(_01622_),
    .A1(net587),
    .A2(net318));
 sg13g2_nand2_1 _24393_ (.Y(_06164_),
    .A(\cpu.genblk1.mmu.r_vtop_i[18][1] ),
    .B(net395));
 sg13g2_o21ai_1 _24394_ (.B1(_06164_),
    .Y(_01623_),
    .A1(net738),
    .A2(_06159_));
 sg13g2_mux2_1 _24395_ (.A0(net737),
    .A1(\cpu.genblk1.mmu.r_vtop_i[18][2] ),
    .S(net318),
    .X(_01624_));
 sg13g2_nand2_1 _24396_ (.Y(_06165_),
    .A(\cpu.genblk1.mmu.r_vtop_i[18][3] ),
    .B(net395));
 sg13g2_o21ai_1 _24397_ (.B1(_06165_),
    .Y(_01625_),
    .A1(net736),
    .A2(net318));
 sg13g2_nand2_1 _24398_ (.Y(_06166_),
    .A(\cpu.genblk1.mmu.r_vtop_i[18][4] ),
    .B(net395));
 sg13g2_o21ai_1 _24399_ (.B1(_06166_),
    .Y(_01626_),
    .A1(net849),
    .A2(_06159_));
 sg13g2_nand2_1 _24400_ (.Y(_06167_),
    .A(\cpu.genblk1.mmu.r_vtop_i[18][5] ),
    .B(net395));
 sg13g2_o21ai_1 _24401_ (.B1(_06167_),
    .Y(_01627_),
    .A1(net735),
    .A2(net318));
 sg13g2_nand2_1 _24402_ (.Y(_06168_),
    .A(\cpu.genblk1.mmu.r_vtop_i[18][6] ),
    .B(net395));
 sg13g2_o21ai_1 _24403_ (.B1(_06168_),
    .Y(_01628_),
    .A1(net734),
    .A2(net318));
 sg13g2_mux2_1 _24404_ (.A0(net848),
    .A1(\cpu.genblk1.mmu.r_vtop_i[18][7] ),
    .S(net318),
    .X(_01629_));
 sg13g2_buf_1 _24405_ (.A(net552),
    .X(_06169_));
 sg13g2_mux2_1 _24406_ (.A0(net475),
    .A1(\cpu.genblk1.mmu.r_vtop_i[18][8] ),
    .S(_06158_),
    .X(_01630_));
 sg13g2_buf_1 _24407_ (.A(net493),
    .X(_06170_));
 sg13g2_mux2_1 _24408_ (.A0(net444),
    .A1(\cpu.genblk1.mmu.r_vtop_i[18][9] ),
    .S(_06158_),
    .X(_01631_));
 sg13g2_nand2_1 _24409_ (.Y(_06171_),
    .A(_05947_),
    .B(net477));
 sg13g2_buf_1 _24410_ (.A(_06171_),
    .X(_06172_));
 sg13g2_buf_1 _24411_ (.A(net394),
    .X(_06173_));
 sg13g2_nand2_1 _24412_ (.Y(_06174_),
    .A(\cpu.genblk1.mmu.r_vtop_i[19][0] ),
    .B(net394));
 sg13g2_o21ai_1 _24413_ (.B1(_06174_),
    .Y(_01632_),
    .A1(net588),
    .A2(net317));
 sg13g2_mux2_1 _24414_ (.A0(net526),
    .A1(\cpu.genblk1.mmu.r_vtop_i[19][10] ),
    .S(net317),
    .X(_01633_));
 sg13g2_nand2_1 _24415_ (.Y(_06175_),
    .A(\cpu.genblk1.mmu.r_vtop_i[19][11] ),
    .B(net394));
 sg13g2_o21ai_1 _24416_ (.B1(_06175_),
    .Y(_01634_),
    .A1(net587),
    .A2(net317));
 sg13g2_nand2_1 _24417_ (.Y(_06176_),
    .A(\cpu.genblk1.mmu.r_vtop_i[19][1] ),
    .B(net394));
 sg13g2_o21ai_1 _24418_ (.B1(_06176_),
    .Y(_01635_),
    .A1(net738),
    .A2(_06173_));
 sg13g2_mux2_1 _24419_ (.A0(net737),
    .A1(\cpu.genblk1.mmu.r_vtop_i[19][2] ),
    .S(net317),
    .X(_01636_));
 sg13g2_nand2_1 _24420_ (.Y(_06177_),
    .A(\cpu.genblk1.mmu.r_vtop_i[19][3] ),
    .B(net394));
 sg13g2_o21ai_1 _24421_ (.B1(_06177_),
    .Y(_01637_),
    .A1(net736),
    .A2(net317));
 sg13g2_nand2_1 _24422_ (.Y(_06178_),
    .A(\cpu.genblk1.mmu.r_vtop_i[19][4] ),
    .B(net394));
 sg13g2_o21ai_1 _24423_ (.B1(_06178_),
    .Y(_01638_),
    .A1(net849),
    .A2(_06173_));
 sg13g2_nand2_1 _24424_ (.Y(_06179_),
    .A(\cpu.genblk1.mmu.r_vtop_i[19][5] ),
    .B(net394));
 sg13g2_o21ai_1 _24425_ (.B1(_06179_),
    .Y(_01639_),
    .A1(net735),
    .A2(net317));
 sg13g2_nand2_1 _24426_ (.Y(_06180_),
    .A(\cpu.genblk1.mmu.r_vtop_i[19][6] ),
    .B(net394));
 sg13g2_o21ai_1 _24427_ (.B1(_06180_),
    .Y(_01640_),
    .A1(net734),
    .A2(net317));
 sg13g2_mux2_1 _24428_ (.A0(net848),
    .A1(\cpu.genblk1.mmu.r_vtop_i[19][7] ),
    .S(net317),
    .X(_01641_));
 sg13g2_mux2_1 _24429_ (.A0(net475),
    .A1(\cpu.genblk1.mmu.r_vtop_i[19][8] ),
    .S(_06172_),
    .X(_01642_));
 sg13g2_mux2_1 _24430_ (.A0(net444),
    .A1(\cpu.genblk1.mmu.r_vtop_i[19][9] ),
    .S(_06172_),
    .X(_01643_));
 sg13g2_nand2_1 _24431_ (.Y(_06181_),
    .A(_06046_),
    .B(_06094_));
 sg13g2_buf_1 _24432_ (.A(_06181_),
    .X(_06182_));
 sg13g2_buf_1 _24433_ (.A(_06182_),
    .X(_06183_));
 sg13g2_nand2_1 _24434_ (.Y(_06184_),
    .A(\cpu.genblk1.mmu.r_vtop_i[1][0] ),
    .B(net316));
 sg13g2_o21ai_1 _24435_ (.B1(_06184_),
    .Y(_01644_),
    .A1(net588),
    .A2(net252));
 sg13g2_mux2_1 _24436_ (.A0(_06161_),
    .A1(\cpu.genblk1.mmu.r_vtop_i[1][10] ),
    .S(net252),
    .X(_01645_));
 sg13g2_nand2_1 _24437_ (.Y(_06185_),
    .A(\cpu.genblk1.mmu.r_vtop_i[1][11] ),
    .B(net316));
 sg13g2_o21ai_1 _24438_ (.B1(_06185_),
    .Y(_01646_),
    .A1(_06162_),
    .A2(net252));
 sg13g2_nand2_1 _24439_ (.Y(_06186_),
    .A(\cpu.genblk1.mmu.r_vtop_i[1][1] ),
    .B(net316));
 sg13g2_o21ai_1 _24440_ (.B1(_06186_),
    .Y(_01647_),
    .A1(_06134_),
    .A2(_06183_));
 sg13g2_mux2_1 _24441_ (.A0(_06136_),
    .A1(\cpu.genblk1.mmu.r_vtop_i[1][2] ),
    .S(net252),
    .X(_01648_));
 sg13g2_nand2_1 _24442_ (.Y(_06187_),
    .A(\cpu.genblk1.mmu.r_vtop_i[1][3] ),
    .B(net316));
 sg13g2_o21ai_1 _24443_ (.B1(_06187_),
    .Y(_01649_),
    .A1(_06137_),
    .A2(net252));
 sg13g2_nand2_1 _24444_ (.Y(_06188_),
    .A(\cpu.genblk1.mmu.r_vtop_i[1][4] ),
    .B(net316));
 sg13g2_o21ai_1 _24445_ (.B1(_06188_),
    .Y(_01650_),
    .A1(_06139_),
    .A2(net252));
 sg13g2_nand2_1 _24446_ (.Y(_06189_),
    .A(\cpu.genblk1.mmu.r_vtop_i[1][5] ),
    .B(net316));
 sg13g2_o21ai_1 _24447_ (.B1(_06189_),
    .Y(_01651_),
    .A1(_06141_),
    .A2(_06183_));
 sg13g2_nand2_1 _24448_ (.Y(_06190_),
    .A(\cpu.genblk1.mmu.r_vtop_i[1][6] ),
    .B(net316));
 sg13g2_o21ai_1 _24449_ (.B1(_06190_),
    .Y(_01652_),
    .A1(_06143_),
    .A2(net252));
 sg13g2_mux2_1 _24450_ (.A0(_06145_),
    .A1(\cpu.genblk1.mmu.r_vtop_i[1][7] ),
    .S(net252),
    .X(_01653_));
 sg13g2_mux2_1 _24451_ (.A0(_06169_),
    .A1(\cpu.genblk1.mmu.r_vtop_i[1][8] ),
    .S(_06182_),
    .X(_01654_));
 sg13g2_mux2_1 _24452_ (.A0(_06170_),
    .A1(\cpu.genblk1.mmu.r_vtop_i[1][9] ),
    .S(net316),
    .X(_01655_));
 sg13g2_nor2_1 _24453_ (.A(_05877_),
    .B(_05928_),
    .Y(_06191_));
 sg13g2_nand2_1 _24454_ (.Y(_06192_),
    .A(_06191_),
    .B(_06050_));
 sg13g2_buf_1 _24455_ (.A(_06192_),
    .X(_06193_));
 sg13g2_buf_1 _24456_ (.A(_06193_),
    .X(_06194_));
 sg13g2_nand2_1 _24457_ (.Y(_06195_),
    .A(\cpu.genblk1.mmu.r_vtop_i[20][0] ),
    .B(net315));
 sg13g2_o21ai_1 _24458_ (.B1(_06195_),
    .Y(_01656_),
    .A1(net588),
    .A2(net251));
 sg13g2_mux2_1 _24459_ (.A0(net526),
    .A1(\cpu.genblk1.mmu.r_vtop_i[20][10] ),
    .S(net251),
    .X(_01657_));
 sg13g2_nand2_1 _24460_ (.Y(_06196_),
    .A(\cpu.genblk1.mmu.r_vtop_i[20][11] ),
    .B(_06193_));
 sg13g2_o21ai_1 _24461_ (.B1(_06196_),
    .Y(_01658_),
    .A1(net587),
    .A2(net251));
 sg13g2_nand2_1 _24462_ (.Y(_06197_),
    .A(\cpu.genblk1.mmu.r_vtop_i[20][1] ),
    .B(net315));
 sg13g2_o21ai_1 _24463_ (.B1(_06197_),
    .Y(_01659_),
    .A1(net738),
    .A2(net251));
 sg13g2_mux2_1 _24464_ (.A0(net737),
    .A1(\cpu.genblk1.mmu.r_vtop_i[20][2] ),
    .S(net251),
    .X(_01660_));
 sg13g2_nand2_1 _24465_ (.Y(_06198_),
    .A(\cpu.genblk1.mmu.r_vtop_i[20][3] ),
    .B(net315));
 sg13g2_o21ai_1 _24466_ (.B1(_06198_),
    .Y(_01661_),
    .A1(net736),
    .A2(net251));
 sg13g2_nand2_1 _24467_ (.Y(_06199_),
    .A(\cpu.genblk1.mmu.r_vtop_i[20][4] ),
    .B(net315));
 sg13g2_o21ai_1 _24468_ (.B1(_06199_),
    .Y(_01662_),
    .A1(net849),
    .A2(_06194_));
 sg13g2_nand2_1 _24469_ (.Y(_06200_),
    .A(\cpu.genblk1.mmu.r_vtop_i[20][5] ),
    .B(net315));
 sg13g2_o21ai_1 _24470_ (.B1(_06200_),
    .Y(_01663_),
    .A1(net735),
    .A2(_06194_));
 sg13g2_nand2_1 _24471_ (.Y(_06201_),
    .A(\cpu.genblk1.mmu.r_vtop_i[20][6] ),
    .B(net315));
 sg13g2_o21ai_1 _24472_ (.B1(_06201_),
    .Y(_01664_),
    .A1(net734),
    .A2(net251));
 sg13g2_mux2_1 _24473_ (.A0(net848),
    .A1(\cpu.genblk1.mmu.r_vtop_i[20][7] ),
    .S(net251),
    .X(_01665_));
 sg13g2_mux2_1 _24474_ (.A0(net475),
    .A1(\cpu.genblk1.mmu.r_vtop_i[20][8] ),
    .S(net315),
    .X(_01666_));
 sg13g2_mux2_1 _24475_ (.A0(net444),
    .A1(\cpu.genblk1.mmu.r_vtop_i[20][9] ),
    .S(net315),
    .X(_01667_));
 sg13g2_nand2_1 _24476_ (.Y(_06202_),
    .A(_06191_),
    .B(_06094_));
 sg13g2_buf_1 _24477_ (.A(_06202_),
    .X(_06203_));
 sg13g2_buf_1 _24478_ (.A(_06203_),
    .X(_06204_));
 sg13g2_nand2_1 _24479_ (.Y(_06205_),
    .A(\cpu.genblk1.mmu.r_vtop_i[21][0] ),
    .B(net314));
 sg13g2_o21ai_1 _24480_ (.B1(_06205_),
    .Y(_01668_),
    .A1(net588),
    .A2(net250));
 sg13g2_mux2_1 _24481_ (.A0(net526),
    .A1(\cpu.genblk1.mmu.r_vtop_i[21][10] ),
    .S(net250),
    .X(_01669_));
 sg13g2_nand2_1 _24482_ (.Y(_06206_),
    .A(\cpu.genblk1.mmu.r_vtop_i[21][11] ),
    .B(_06203_));
 sg13g2_o21ai_1 _24483_ (.B1(_06206_),
    .Y(_01670_),
    .A1(net587),
    .A2(net250));
 sg13g2_nand2_1 _24484_ (.Y(_06207_),
    .A(\cpu.genblk1.mmu.r_vtop_i[21][1] ),
    .B(net314));
 sg13g2_o21ai_1 _24485_ (.B1(_06207_),
    .Y(_01671_),
    .A1(net738),
    .A2(_06204_));
 sg13g2_mux2_1 _24486_ (.A0(net737),
    .A1(\cpu.genblk1.mmu.r_vtop_i[21][2] ),
    .S(net250),
    .X(_01672_));
 sg13g2_nand2_1 _24487_ (.Y(_06208_),
    .A(\cpu.genblk1.mmu.r_vtop_i[21][3] ),
    .B(net314));
 sg13g2_o21ai_1 _24488_ (.B1(_06208_),
    .Y(_01673_),
    .A1(net736),
    .A2(net250));
 sg13g2_nand2_1 _24489_ (.Y(_06209_),
    .A(\cpu.genblk1.mmu.r_vtop_i[21][4] ),
    .B(net314));
 sg13g2_o21ai_1 _24490_ (.B1(_06209_),
    .Y(_01674_),
    .A1(net849),
    .A2(net250));
 sg13g2_nand2_1 _24491_ (.Y(_06210_),
    .A(\cpu.genblk1.mmu.r_vtop_i[21][5] ),
    .B(net314));
 sg13g2_o21ai_1 _24492_ (.B1(_06210_),
    .Y(_01675_),
    .A1(net735),
    .A2(_06204_));
 sg13g2_nand2_1 _24493_ (.Y(_06211_),
    .A(\cpu.genblk1.mmu.r_vtop_i[21][6] ),
    .B(net314));
 sg13g2_o21ai_1 _24494_ (.B1(_06211_),
    .Y(_01676_),
    .A1(net734),
    .A2(net250));
 sg13g2_mux2_1 _24495_ (.A0(net848),
    .A1(\cpu.genblk1.mmu.r_vtop_i[21][7] ),
    .S(net250),
    .X(_01677_));
 sg13g2_mux2_1 _24496_ (.A0(net475),
    .A1(\cpu.genblk1.mmu.r_vtop_i[21][8] ),
    .S(net314),
    .X(_01678_));
 sg13g2_mux2_1 _24497_ (.A0(net444),
    .A1(\cpu.genblk1.mmu.r_vtop_i[21][9] ),
    .S(net314),
    .X(_01679_));
 sg13g2_nand3_1 _24498_ (.B(_06191_),
    .C(net476),
    .A(_06105_),
    .Y(_06212_));
 sg13g2_buf_1 _24499_ (.A(_06212_),
    .X(_06213_));
 sg13g2_buf_1 _24500_ (.A(net393),
    .X(_06214_));
 sg13g2_nand2_1 _24501_ (.Y(_06215_),
    .A(\cpu.genblk1.mmu.r_vtop_i[22][0] ),
    .B(net393));
 sg13g2_o21ai_1 _24502_ (.B1(_06215_),
    .Y(_01680_),
    .A1(net588),
    .A2(net313));
 sg13g2_mux2_1 _24503_ (.A0(net526),
    .A1(\cpu.genblk1.mmu.r_vtop_i[22][10] ),
    .S(net313),
    .X(_01681_));
 sg13g2_nand2_1 _24504_ (.Y(_06216_),
    .A(\cpu.genblk1.mmu.r_vtop_i[22][11] ),
    .B(net393));
 sg13g2_o21ai_1 _24505_ (.B1(_06216_),
    .Y(_01682_),
    .A1(net587),
    .A2(net313));
 sg13g2_nand2_1 _24506_ (.Y(_06217_),
    .A(\cpu.genblk1.mmu.r_vtop_i[22][1] ),
    .B(net393));
 sg13g2_o21ai_1 _24507_ (.B1(_06217_),
    .Y(_01683_),
    .A1(net738),
    .A2(_06214_));
 sg13g2_mux2_1 _24508_ (.A0(net737),
    .A1(\cpu.genblk1.mmu.r_vtop_i[22][2] ),
    .S(net313),
    .X(_01684_));
 sg13g2_nand2_1 _24509_ (.Y(_06218_),
    .A(\cpu.genblk1.mmu.r_vtop_i[22][3] ),
    .B(net393));
 sg13g2_o21ai_1 _24510_ (.B1(_06218_),
    .Y(_01685_),
    .A1(net736),
    .A2(net313));
 sg13g2_nand2_1 _24511_ (.Y(_06219_),
    .A(\cpu.genblk1.mmu.r_vtop_i[22][4] ),
    .B(net393));
 sg13g2_o21ai_1 _24512_ (.B1(_06219_),
    .Y(_01686_),
    .A1(net849),
    .A2(net313));
 sg13g2_nand2_1 _24513_ (.Y(_06220_),
    .A(\cpu.genblk1.mmu.r_vtop_i[22][5] ),
    .B(net393));
 sg13g2_o21ai_1 _24514_ (.B1(_06220_),
    .Y(_01687_),
    .A1(net735),
    .A2(_06214_));
 sg13g2_nand2_1 _24515_ (.Y(_06221_),
    .A(\cpu.genblk1.mmu.r_vtop_i[22][6] ),
    .B(net393));
 sg13g2_o21ai_1 _24516_ (.B1(_06221_),
    .Y(_01688_),
    .A1(net734),
    .A2(net313));
 sg13g2_mux2_1 _24517_ (.A0(net848),
    .A1(\cpu.genblk1.mmu.r_vtop_i[22][7] ),
    .S(net313),
    .X(_01689_));
 sg13g2_mux2_1 _24518_ (.A0(net475),
    .A1(\cpu.genblk1.mmu.r_vtop_i[22][8] ),
    .S(_06213_),
    .X(_01690_));
 sg13g2_mux2_1 _24519_ (.A0(net444),
    .A1(\cpu.genblk1.mmu.r_vtop_i[22][9] ),
    .S(_06213_),
    .X(_01691_));
 sg13g2_nand3_1 _24520_ (.B(_06191_),
    .C(net476),
    .A(_05844_),
    .Y(_06222_));
 sg13g2_buf_1 _24521_ (.A(_06222_),
    .X(_06223_));
 sg13g2_buf_1 _24522_ (.A(net392),
    .X(_06224_));
 sg13g2_nand2_1 _24523_ (.Y(_06225_),
    .A(\cpu.genblk1.mmu.r_vtop_i[23][0] ),
    .B(net392));
 sg13g2_o21ai_1 _24524_ (.B1(_06225_),
    .Y(_01692_),
    .A1(net588),
    .A2(net312));
 sg13g2_mux2_1 _24525_ (.A0(net526),
    .A1(\cpu.genblk1.mmu.r_vtop_i[23][10] ),
    .S(net312),
    .X(_01693_));
 sg13g2_nand2_1 _24526_ (.Y(_06226_),
    .A(\cpu.genblk1.mmu.r_vtop_i[23][11] ),
    .B(net392));
 sg13g2_o21ai_1 _24527_ (.B1(_06226_),
    .Y(_01694_),
    .A1(net587),
    .A2(net312));
 sg13g2_nand2_1 _24528_ (.Y(_06227_),
    .A(\cpu.genblk1.mmu.r_vtop_i[23][1] ),
    .B(net392));
 sg13g2_o21ai_1 _24529_ (.B1(_06227_),
    .Y(_01695_),
    .A1(net738),
    .A2(net312));
 sg13g2_mux2_1 _24530_ (.A0(net737),
    .A1(\cpu.genblk1.mmu.r_vtop_i[23][2] ),
    .S(net312),
    .X(_01696_));
 sg13g2_nand2_1 _24531_ (.Y(_06228_),
    .A(\cpu.genblk1.mmu.r_vtop_i[23][3] ),
    .B(net392));
 sg13g2_o21ai_1 _24532_ (.B1(_06228_),
    .Y(_01697_),
    .A1(net736),
    .A2(net312));
 sg13g2_nand2_1 _24533_ (.Y(_06229_),
    .A(\cpu.genblk1.mmu.r_vtop_i[23][4] ),
    .B(net392));
 sg13g2_o21ai_1 _24534_ (.B1(_06229_),
    .Y(_01698_),
    .A1(net849),
    .A2(_06224_));
 sg13g2_nand2_1 _24535_ (.Y(_06230_),
    .A(\cpu.genblk1.mmu.r_vtop_i[23][5] ),
    .B(net392));
 sg13g2_o21ai_1 _24536_ (.B1(_06230_),
    .Y(_01699_),
    .A1(net735),
    .A2(_06224_));
 sg13g2_nand2_1 _24537_ (.Y(_06231_),
    .A(\cpu.genblk1.mmu.r_vtop_i[23][6] ),
    .B(net392));
 sg13g2_o21ai_1 _24538_ (.B1(_06231_),
    .Y(_01700_),
    .A1(net734),
    .A2(net312));
 sg13g2_mux2_1 _24539_ (.A0(net848),
    .A1(\cpu.genblk1.mmu.r_vtop_i[23][7] ),
    .S(net312),
    .X(_01701_));
 sg13g2_mux2_1 _24540_ (.A0(net475),
    .A1(\cpu.genblk1.mmu.r_vtop_i[23][8] ),
    .S(_06223_),
    .X(_01702_));
 sg13g2_mux2_1 _24541_ (.A0(net444),
    .A1(\cpu.genblk1.mmu.r_vtop_i[23][9] ),
    .S(_06223_),
    .X(_01703_));
 sg13g2_inv_1 _24542_ (.Y(_06232_),
    .A(_05976_));
 sg13g2_nand3_1 _24543_ (.B(_06232_),
    .C(net476),
    .A(_06128_),
    .Y(_06233_));
 sg13g2_buf_1 _24544_ (.A(_06233_),
    .X(_06234_));
 sg13g2_buf_1 _24545_ (.A(_06234_),
    .X(_06235_));
 sg13g2_nand2_1 _24546_ (.Y(_06236_),
    .A(\cpu.genblk1.mmu.r_vtop_i[24][0] ),
    .B(net391));
 sg13g2_o21ai_1 _24547_ (.B1(_06236_),
    .Y(_01704_),
    .A1(_06156_),
    .A2(net311));
 sg13g2_mux2_1 _24548_ (.A0(net526),
    .A1(\cpu.genblk1.mmu.r_vtop_i[24][10] ),
    .S(net311),
    .X(_01705_));
 sg13g2_nand2_1 _24549_ (.Y(_06237_),
    .A(\cpu.genblk1.mmu.r_vtop_i[24][11] ),
    .B(net391));
 sg13g2_o21ai_1 _24550_ (.B1(_06237_),
    .Y(_01706_),
    .A1(_06162_),
    .A2(net311));
 sg13g2_nand2_1 _24551_ (.Y(_06238_),
    .A(\cpu.genblk1.mmu.r_vtop_i[24][1] ),
    .B(net391));
 sg13g2_o21ai_1 _24552_ (.B1(_06238_),
    .Y(_01707_),
    .A1(_06134_),
    .A2(net311));
 sg13g2_mux2_1 _24553_ (.A0(_06136_),
    .A1(\cpu.genblk1.mmu.r_vtop_i[24][2] ),
    .S(net311),
    .X(_01708_));
 sg13g2_nand2_1 _24554_ (.Y(_06239_),
    .A(\cpu.genblk1.mmu.r_vtop_i[24][3] ),
    .B(net391));
 sg13g2_o21ai_1 _24555_ (.B1(_06239_),
    .Y(_01709_),
    .A1(_06137_),
    .A2(net311));
 sg13g2_nand2_1 _24556_ (.Y(_06240_),
    .A(\cpu.genblk1.mmu.r_vtop_i[24][4] ),
    .B(net391));
 sg13g2_o21ai_1 _24557_ (.B1(_06240_),
    .Y(_01710_),
    .A1(net849),
    .A2(_06235_));
 sg13g2_nand2_1 _24558_ (.Y(_06241_),
    .A(\cpu.genblk1.mmu.r_vtop_i[24][5] ),
    .B(net391));
 sg13g2_o21ai_1 _24559_ (.B1(_06241_),
    .Y(_01711_),
    .A1(_06141_),
    .A2(_06235_));
 sg13g2_nand2_1 _24560_ (.Y(_06242_),
    .A(\cpu.genblk1.mmu.r_vtop_i[24][6] ),
    .B(net391));
 sg13g2_o21ai_1 _24561_ (.B1(_06242_),
    .Y(_01712_),
    .A1(net734),
    .A2(net311));
 sg13g2_mux2_1 _24562_ (.A0(_06145_),
    .A1(\cpu.genblk1.mmu.r_vtop_i[24][7] ),
    .S(net311),
    .X(_01713_));
 sg13g2_mux2_1 _24563_ (.A0(net475),
    .A1(\cpu.genblk1.mmu.r_vtop_i[24][8] ),
    .S(_06234_),
    .X(_01714_));
 sg13g2_mux2_1 _24564_ (.A0(_06170_),
    .A1(\cpu.genblk1.mmu.r_vtop_i[24][9] ),
    .S(net391),
    .X(_01715_));
 sg13g2_nand3_1 _24565_ (.B(_06232_),
    .C(_06094_),
    .A(net978),
    .Y(_06243_));
 sg13g2_buf_1 _24566_ (.A(_06243_),
    .X(_06244_));
 sg13g2_buf_1 _24567_ (.A(net310),
    .X(_06245_));
 sg13g2_nand2_1 _24568_ (.Y(_06246_),
    .A(\cpu.genblk1.mmu.r_vtop_i[25][0] ),
    .B(net310));
 sg13g2_o21ai_1 _24569_ (.B1(_06246_),
    .Y(_01716_),
    .A1(net588),
    .A2(net249));
 sg13g2_mux2_1 _24570_ (.A0(net526),
    .A1(\cpu.genblk1.mmu.r_vtop_i[25][10] ),
    .S(net249),
    .X(_01717_));
 sg13g2_nand2_1 _24571_ (.Y(_06247_),
    .A(\cpu.genblk1.mmu.r_vtop_i[25][11] ),
    .B(_06244_));
 sg13g2_o21ai_1 _24572_ (.B1(_06247_),
    .Y(_01718_),
    .A1(net587),
    .A2(net249));
 sg13g2_buf_1 _24573_ (.A(net873),
    .X(_06248_));
 sg13g2_nand2_1 _24574_ (.Y(_06249_),
    .A(\cpu.genblk1.mmu.r_vtop_i[25][1] ),
    .B(net310));
 sg13g2_o21ai_1 _24575_ (.B1(_06249_),
    .Y(_01719_),
    .A1(net733),
    .A2(net249));
 sg13g2_buf_1 _24576_ (.A(net872),
    .X(_06250_));
 sg13g2_mux2_1 _24577_ (.A0(net732),
    .A1(\cpu.genblk1.mmu.r_vtop_i[25][2] ),
    .S(net249),
    .X(_01720_));
 sg13g2_buf_1 _24578_ (.A(net871),
    .X(_06251_));
 sg13g2_nand2_1 _24579_ (.Y(_06252_),
    .A(\cpu.genblk1.mmu.r_vtop_i[25][3] ),
    .B(net310));
 sg13g2_o21ai_1 _24580_ (.B1(_06252_),
    .Y(_01721_),
    .A1(net731),
    .A2(net249));
 sg13g2_buf_1 _24581_ (.A(net1037),
    .X(_06253_));
 sg13g2_nand2_1 _24582_ (.Y(_06254_),
    .A(\cpu.genblk1.mmu.r_vtop_i[25][4] ),
    .B(_06244_));
 sg13g2_o21ai_1 _24583_ (.B1(_06254_),
    .Y(_01722_),
    .A1(net847),
    .A2(_06245_));
 sg13g2_buf_1 _24584_ (.A(net869),
    .X(_06255_));
 sg13g2_nand2_1 _24585_ (.Y(_06256_),
    .A(\cpu.genblk1.mmu.r_vtop_i[25][5] ),
    .B(net310));
 sg13g2_o21ai_1 _24586_ (.B1(_06256_),
    .Y(_01723_),
    .A1(net730),
    .A2(_06245_));
 sg13g2_buf_1 _24587_ (.A(net889),
    .X(_06257_));
 sg13g2_nand2_1 _24588_ (.Y(_06258_),
    .A(\cpu.genblk1.mmu.r_vtop_i[25][6] ),
    .B(net310));
 sg13g2_o21ai_1 _24589_ (.B1(_06258_),
    .Y(_01724_),
    .A1(net729),
    .A2(net249));
 sg13g2_buf_1 _24590_ (.A(net999),
    .X(_06259_));
 sg13g2_mux2_1 _24591_ (.A0(net846),
    .A1(\cpu.genblk1.mmu.r_vtop_i[25][7] ),
    .S(net249),
    .X(_01725_));
 sg13g2_mux2_1 _24592_ (.A0(net475),
    .A1(\cpu.genblk1.mmu.r_vtop_i[25][8] ),
    .S(net310),
    .X(_01726_));
 sg13g2_mux2_1 _24593_ (.A0(net444),
    .A1(\cpu.genblk1.mmu.r_vtop_i[25][9] ),
    .S(net310),
    .X(_01727_));
 sg13g2_nand2_1 _24594_ (.Y(_06260_),
    .A(_05985_),
    .B(net477));
 sg13g2_buf_1 _24595_ (.A(_06260_),
    .X(_06261_));
 sg13g2_buf_1 _24596_ (.A(net390),
    .X(_06262_));
 sg13g2_nand2_1 _24597_ (.Y(_06263_),
    .A(\cpu.genblk1.mmu.r_vtop_i[26][0] ),
    .B(net390));
 sg13g2_o21ai_1 _24598_ (.B1(_06263_),
    .Y(_01728_),
    .A1(_06156_),
    .A2(net309));
 sg13g2_mux2_1 _24599_ (.A0(_06161_),
    .A1(\cpu.genblk1.mmu.r_vtop_i[26][10] ),
    .S(net309),
    .X(_01729_));
 sg13g2_nand2_1 _24600_ (.Y(_06264_),
    .A(\cpu.genblk1.mmu.r_vtop_i[26][11] ),
    .B(net390));
 sg13g2_o21ai_1 _24601_ (.B1(_06264_),
    .Y(_01730_),
    .A1(net587),
    .A2(net309));
 sg13g2_nand2_1 _24602_ (.Y(_06265_),
    .A(\cpu.genblk1.mmu.r_vtop_i[26][1] ),
    .B(net390));
 sg13g2_o21ai_1 _24603_ (.B1(_06265_),
    .Y(_01731_),
    .A1(net733),
    .A2(net309));
 sg13g2_mux2_1 _24604_ (.A0(net732),
    .A1(\cpu.genblk1.mmu.r_vtop_i[26][2] ),
    .S(net309),
    .X(_01732_));
 sg13g2_nand2_1 _24605_ (.Y(_06266_),
    .A(\cpu.genblk1.mmu.r_vtop_i[26][3] ),
    .B(net390));
 sg13g2_o21ai_1 _24606_ (.B1(_06266_),
    .Y(_01733_),
    .A1(net731),
    .A2(net309));
 sg13g2_nand2_1 _24607_ (.Y(_06267_),
    .A(\cpu.genblk1.mmu.r_vtop_i[26][4] ),
    .B(net390));
 sg13g2_o21ai_1 _24608_ (.B1(_06267_),
    .Y(_01734_),
    .A1(net847),
    .A2(_06262_));
 sg13g2_nand2_1 _24609_ (.Y(_06268_),
    .A(\cpu.genblk1.mmu.r_vtop_i[26][5] ),
    .B(net390));
 sg13g2_o21ai_1 _24610_ (.B1(_06268_),
    .Y(_01735_),
    .A1(net730),
    .A2(_06262_));
 sg13g2_nand2_1 _24611_ (.Y(_06269_),
    .A(\cpu.genblk1.mmu.r_vtop_i[26][6] ),
    .B(net390));
 sg13g2_o21ai_1 _24612_ (.B1(_06269_),
    .Y(_01736_),
    .A1(net729),
    .A2(net309));
 sg13g2_mux2_1 _24613_ (.A0(net846),
    .A1(\cpu.genblk1.mmu.r_vtop_i[26][7] ),
    .S(net309),
    .X(_01737_));
 sg13g2_mux2_1 _24614_ (.A0(_06169_),
    .A1(\cpu.genblk1.mmu.r_vtop_i[26][8] ),
    .S(_06261_),
    .X(_01738_));
 sg13g2_mux2_1 _24615_ (.A0(net444),
    .A1(\cpu.genblk1.mmu.r_vtop_i[26][9] ),
    .S(_06261_),
    .X(_01739_));
 sg13g2_buf_1 _24616_ (.A(net666),
    .X(_06270_));
 sg13g2_nand2_1 _24617_ (.Y(_06271_),
    .A(_05990_),
    .B(net477));
 sg13g2_buf_1 _24618_ (.A(_06271_),
    .X(_06272_));
 sg13g2_buf_1 _24619_ (.A(net389),
    .X(_06273_));
 sg13g2_nand2_1 _24620_ (.Y(_06274_),
    .A(\cpu.genblk1.mmu.r_vtop_i[27][0] ),
    .B(net389));
 sg13g2_o21ai_1 _24621_ (.B1(_06274_),
    .Y(_01740_),
    .A1(net586),
    .A2(net308));
 sg13g2_buf_1 _24622_ (.A(net605),
    .X(_06275_));
 sg13g2_mux2_1 _24623_ (.A0(net525),
    .A1(\cpu.genblk1.mmu.r_vtop_i[27][10] ),
    .S(net308),
    .X(_01741_));
 sg13g2_buf_1 _24624_ (.A(net699),
    .X(_06276_));
 sg13g2_nand2_1 _24625_ (.Y(_06277_),
    .A(\cpu.genblk1.mmu.r_vtop_i[27][11] ),
    .B(_06272_));
 sg13g2_o21ai_1 _24626_ (.B1(_06277_),
    .Y(_01742_),
    .A1(_06276_),
    .A2(net308));
 sg13g2_nand2_1 _24627_ (.Y(_06278_),
    .A(\cpu.genblk1.mmu.r_vtop_i[27][1] ),
    .B(net389));
 sg13g2_o21ai_1 _24628_ (.B1(_06278_),
    .Y(_01743_),
    .A1(net733),
    .A2(net308));
 sg13g2_mux2_1 _24629_ (.A0(net732),
    .A1(\cpu.genblk1.mmu.r_vtop_i[27][2] ),
    .S(net308),
    .X(_01744_));
 sg13g2_nand2_1 _24630_ (.Y(_06279_),
    .A(\cpu.genblk1.mmu.r_vtop_i[27][3] ),
    .B(net389));
 sg13g2_o21ai_1 _24631_ (.B1(_06279_),
    .Y(_01745_),
    .A1(net731),
    .A2(net308));
 sg13g2_nand2_1 _24632_ (.Y(_06280_),
    .A(\cpu.genblk1.mmu.r_vtop_i[27][4] ),
    .B(_06272_));
 sg13g2_o21ai_1 _24633_ (.B1(_06280_),
    .Y(_01746_),
    .A1(net847),
    .A2(_06273_));
 sg13g2_nand2_1 _24634_ (.Y(_06281_),
    .A(\cpu.genblk1.mmu.r_vtop_i[27][5] ),
    .B(net389));
 sg13g2_o21ai_1 _24635_ (.B1(_06281_),
    .Y(_01747_),
    .A1(net730),
    .A2(_06273_));
 sg13g2_nand2_1 _24636_ (.Y(_06282_),
    .A(\cpu.genblk1.mmu.r_vtop_i[27][6] ),
    .B(net389));
 sg13g2_o21ai_1 _24637_ (.B1(_06282_),
    .Y(_01748_),
    .A1(net729),
    .A2(net308));
 sg13g2_mux2_1 _24638_ (.A0(net846),
    .A1(\cpu.genblk1.mmu.r_vtop_i[27][7] ),
    .S(net308),
    .X(_01749_));
 sg13g2_buf_1 _24639_ (.A(net552),
    .X(_06283_));
 sg13g2_mux2_1 _24640_ (.A0(net474),
    .A1(\cpu.genblk1.mmu.r_vtop_i[27][8] ),
    .S(net389),
    .X(_01750_));
 sg13g2_buf_1 _24641_ (.A(net493),
    .X(_06284_));
 sg13g2_mux2_1 _24642_ (.A0(net443),
    .A1(\cpu.genblk1.mmu.r_vtop_i[27][9] ),
    .S(net389),
    .X(_01751_));
 sg13g2_nor2_1 _24643_ (.A(_05877_),
    .B(_05976_),
    .Y(_06285_));
 sg13g2_nand2_1 _24644_ (.Y(_06286_),
    .A(_06285_),
    .B(_06050_));
 sg13g2_buf_1 _24645_ (.A(_06286_),
    .X(_06287_));
 sg13g2_buf_1 _24646_ (.A(net307),
    .X(_06288_));
 sg13g2_nand2_1 _24647_ (.Y(_06289_),
    .A(\cpu.genblk1.mmu.r_vtop_i[28][0] ),
    .B(net307));
 sg13g2_o21ai_1 _24648_ (.B1(_06289_),
    .Y(_01752_),
    .A1(net586),
    .A2(net248));
 sg13g2_mux2_1 _24649_ (.A0(net525),
    .A1(\cpu.genblk1.mmu.r_vtop_i[28][10] ),
    .S(net248),
    .X(_01753_));
 sg13g2_nand2_1 _24650_ (.Y(_06290_),
    .A(\cpu.genblk1.mmu.r_vtop_i[28][11] ),
    .B(_06287_));
 sg13g2_o21ai_1 _24651_ (.B1(_06290_),
    .Y(_01754_),
    .A1(net585),
    .A2(_06288_));
 sg13g2_nand2_1 _24652_ (.Y(_06291_),
    .A(\cpu.genblk1.mmu.r_vtop_i[28][1] ),
    .B(net307));
 sg13g2_o21ai_1 _24653_ (.B1(_06291_),
    .Y(_01755_),
    .A1(net733),
    .A2(net248));
 sg13g2_mux2_1 _24654_ (.A0(net732),
    .A1(\cpu.genblk1.mmu.r_vtop_i[28][2] ),
    .S(net248),
    .X(_01756_));
 sg13g2_nand2_1 _24655_ (.Y(_06292_),
    .A(\cpu.genblk1.mmu.r_vtop_i[28][3] ),
    .B(net307));
 sg13g2_o21ai_1 _24656_ (.B1(_06292_),
    .Y(_01757_),
    .A1(net731),
    .A2(net248));
 sg13g2_nand2_1 _24657_ (.Y(_06293_),
    .A(\cpu.genblk1.mmu.r_vtop_i[28][4] ),
    .B(net307));
 sg13g2_o21ai_1 _24658_ (.B1(_06293_),
    .Y(_01758_),
    .A1(net847),
    .A2(_06288_));
 sg13g2_nand2_1 _24659_ (.Y(_06294_),
    .A(\cpu.genblk1.mmu.r_vtop_i[28][5] ),
    .B(net307));
 sg13g2_o21ai_1 _24660_ (.B1(_06294_),
    .Y(_01759_),
    .A1(net730),
    .A2(net248));
 sg13g2_nand2_1 _24661_ (.Y(_06295_),
    .A(\cpu.genblk1.mmu.r_vtop_i[28][6] ),
    .B(net307));
 sg13g2_o21ai_1 _24662_ (.B1(_06295_),
    .Y(_01760_),
    .A1(net729),
    .A2(net248));
 sg13g2_mux2_1 _24663_ (.A0(net846),
    .A1(\cpu.genblk1.mmu.r_vtop_i[28][7] ),
    .S(net248),
    .X(_01761_));
 sg13g2_mux2_1 _24664_ (.A0(net474),
    .A1(\cpu.genblk1.mmu.r_vtop_i[28][8] ),
    .S(_06287_),
    .X(_01762_));
 sg13g2_mux2_1 _24665_ (.A0(net443),
    .A1(\cpu.genblk1.mmu.r_vtop_i[28][9] ),
    .S(net307),
    .X(_01763_));
 sg13g2_nand2_1 _24666_ (.Y(_06296_),
    .A(_06285_),
    .B(_06094_));
 sg13g2_buf_1 _24667_ (.A(_06296_),
    .X(_06297_));
 sg13g2_buf_1 _24668_ (.A(net306),
    .X(_06298_));
 sg13g2_nand2_1 _24669_ (.Y(_06299_),
    .A(\cpu.genblk1.mmu.r_vtop_i[29][0] ),
    .B(net306));
 sg13g2_o21ai_1 _24670_ (.B1(_06299_),
    .Y(_01764_),
    .A1(net586),
    .A2(net247));
 sg13g2_mux2_1 _24671_ (.A0(net525),
    .A1(\cpu.genblk1.mmu.r_vtop_i[29][10] ),
    .S(net247),
    .X(_01765_));
 sg13g2_nand2_1 _24672_ (.Y(_06300_),
    .A(\cpu.genblk1.mmu.r_vtop_i[29][11] ),
    .B(_06297_));
 sg13g2_o21ai_1 _24673_ (.B1(_06300_),
    .Y(_01766_),
    .A1(net585),
    .A2(_06298_));
 sg13g2_nand2_1 _24674_ (.Y(_06301_),
    .A(\cpu.genblk1.mmu.r_vtop_i[29][1] ),
    .B(net306));
 sg13g2_o21ai_1 _24675_ (.B1(_06301_),
    .Y(_01767_),
    .A1(net733),
    .A2(net247));
 sg13g2_mux2_1 _24676_ (.A0(net732),
    .A1(\cpu.genblk1.mmu.r_vtop_i[29][2] ),
    .S(net247),
    .X(_01768_));
 sg13g2_nand2_1 _24677_ (.Y(_06302_),
    .A(\cpu.genblk1.mmu.r_vtop_i[29][3] ),
    .B(net306));
 sg13g2_o21ai_1 _24678_ (.B1(_06302_),
    .Y(_01769_),
    .A1(net731),
    .A2(net247));
 sg13g2_nand2_1 _24679_ (.Y(_06303_),
    .A(\cpu.genblk1.mmu.r_vtop_i[29][4] ),
    .B(net306));
 sg13g2_o21ai_1 _24680_ (.B1(_06303_),
    .Y(_01770_),
    .A1(net847),
    .A2(_06298_));
 sg13g2_nand2_1 _24681_ (.Y(_06304_),
    .A(\cpu.genblk1.mmu.r_vtop_i[29][5] ),
    .B(net306));
 sg13g2_o21ai_1 _24682_ (.B1(_06304_),
    .Y(_01771_),
    .A1(_06255_),
    .A2(net247));
 sg13g2_nand2_1 _24683_ (.Y(_06305_),
    .A(\cpu.genblk1.mmu.r_vtop_i[29][6] ),
    .B(net306));
 sg13g2_o21ai_1 _24684_ (.B1(_06305_),
    .Y(_01772_),
    .A1(net729),
    .A2(net247));
 sg13g2_mux2_1 _24685_ (.A0(net846),
    .A1(\cpu.genblk1.mmu.r_vtop_i[29][7] ),
    .S(net247),
    .X(_01773_));
 sg13g2_mux2_1 _24686_ (.A0(net474),
    .A1(\cpu.genblk1.mmu.r_vtop_i[29][8] ),
    .S(_06297_),
    .X(_01774_));
 sg13g2_mux2_1 _24687_ (.A0(net443),
    .A1(\cpu.genblk1.mmu.r_vtop_i[29][9] ),
    .S(net306),
    .X(_01775_));
 sg13g2_nand3_1 _24688_ (.B(_06046_),
    .C(net476),
    .A(_06105_),
    .Y(_06306_));
 sg13g2_buf_1 _24689_ (.A(_06306_),
    .X(_06307_));
 sg13g2_buf_1 _24690_ (.A(net388),
    .X(_06308_));
 sg13g2_nand2_1 _24691_ (.Y(_06309_),
    .A(\cpu.genblk1.mmu.r_vtop_i[2][0] ),
    .B(net388));
 sg13g2_o21ai_1 _24692_ (.B1(_06309_),
    .Y(_01776_),
    .A1(net586),
    .A2(net305));
 sg13g2_mux2_1 _24693_ (.A0(net525),
    .A1(\cpu.genblk1.mmu.r_vtop_i[2][10] ),
    .S(net305),
    .X(_01777_));
 sg13g2_nand2_1 _24694_ (.Y(_06310_),
    .A(\cpu.genblk1.mmu.r_vtop_i[2][11] ),
    .B(_06307_));
 sg13g2_o21ai_1 _24695_ (.B1(_06310_),
    .Y(_01778_),
    .A1(net585),
    .A2(net305));
 sg13g2_nand2_1 _24696_ (.Y(_06311_),
    .A(\cpu.genblk1.mmu.r_vtop_i[2][1] ),
    .B(net388));
 sg13g2_o21ai_1 _24697_ (.B1(_06311_),
    .Y(_01779_),
    .A1(net733),
    .A2(net305));
 sg13g2_mux2_1 _24698_ (.A0(_06250_),
    .A1(\cpu.genblk1.mmu.r_vtop_i[2][2] ),
    .S(net305),
    .X(_01780_));
 sg13g2_nand2_1 _24699_ (.Y(_06312_),
    .A(\cpu.genblk1.mmu.r_vtop_i[2][3] ),
    .B(net388));
 sg13g2_o21ai_1 _24700_ (.B1(_06312_),
    .Y(_01781_),
    .A1(net731),
    .A2(net305));
 sg13g2_nand2_1 _24701_ (.Y(_06313_),
    .A(\cpu.genblk1.mmu.r_vtop_i[2][4] ),
    .B(_06307_));
 sg13g2_o21ai_1 _24702_ (.B1(_06313_),
    .Y(_01782_),
    .A1(_06253_),
    .A2(_06308_));
 sg13g2_nand2_1 _24703_ (.Y(_06314_),
    .A(\cpu.genblk1.mmu.r_vtop_i[2][5] ),
    .B(net388));
 sg13g2_o21ai_1 _24704_ (.B1(_06314_),
    .Y(_01783_),
    .A1(net730),
    .A2(_06308_));
 sg13g2_nand2_1 _24705_ (.Y(_06315_),
    .A(\cpu.genblk1.mmu.r_vtop_i[2][6] ),
    .B(net388));
 sg13g2_o21ai_1 _24706_ (.B1(_06315_),
    .Y(_01784_),
    .A1(net729),
    .A2(net305));
 sg13g2_mux2_1 _24707_ (.A0(net846),
    .A1(\cpu.genblk1.mmu.r_vtop_i[2][7] ),
    .S(net305),
    .X(_01785_));
 sg13g2_mux2_1 _24708_ (.A0(net474),
    .A1(\cpu.genblk1.mmu.r_vtop_i[2][8] ),
    .S(net388),
    .X(_01786_));
 sg13g2_mux2_1 _24709_ (.A0(net443),
    .A1(\cpu.genblk1.mmu.r_vtop_i[2][9] ),
    .S(net388),
    .X(_01787_));
 sg13g2_nand3_1 _24710_ (.B(_06285_),
    .C(net476),
    .A(_06105_),
    .Y(_06316_));
 sg13g2_buf_1 _24711_ (.A(_06316_),
    .X(_06317_));
 sg13g2_buf_1 _24712_ (.A(net387),
    .X(_06318_));
 sg13g2_nand2_1 _24713_ (.Y(_06319_),
    .A(\cpu.genblk1.mmu.r_vtop_i[30][0] ),
    .B(net387));
 sg13g2_o21ai_1 _24714_ (.B1(_06319_),
    .Y(_01788_),
    .A1(net586),
    .A2(net304));
 sg13g2_mux2_1 _24715_ (.A0(net525),
    .A1(\cpu.genblk1.mmu.r_vtop_i[30][10] ),
    .S(net304),
    .X(_01789_));
 sg13g2_nand2_1 _24716_ (.Y(_06320_),
    .A(\cpu.genblk1.mmu.r_vtop_i[30][11] ),
    .B(_06317_));
 sg13g2_o21ai_1 _24717_ (.B1(_06320_),
    .Y(_01790_),
    .A1(net585),
    .A2(_06318_));
 sg13g2_nand2_1 _24718_ (.Y(_06321_),
    .A(\cpu.genblk1.mmu.r_vtop_i[30][1] ),
    .B(net387));
 sg13g2_o21ai_1 _24719_ (.B1(_06321_),
    .Y(_01791_),
    .A1(net733),
    .A2(net304));
 sg13g2_mux2_1 _24720_ (.A0(net732),
    .A1(\cpu.genblk1.mmu.r_vtop_i[30][2] ),
    .S(net304),
    .X(_01792_));
 sg13g2_nand2_1 _24721_ (.Y(_06322_),
    .A(\cpu.genblk1.mmu.r_vtop_i[30][3] ),
    .B(net387));
 sg13g2_o21ai_1 _24722_ (.B1(_06322_),
    .Y(_01793_),
    .A1(_06251_),
    .A2(net304));
 sg13g2_nand2_1 _24723_ (.Y(_06323_),
    .A(\cpu.genblk1.mmu.r_vtop_i[30][4] ),
    .B(net387));
 sg13g2_o21ai_1 _24724_ (.B1(_06323_),
    .Y(_01794_),
    .A1(net847),
    .A2(_06318_));
 sg13g2_nand2_1 _24725_ (.Y(_06324_),
    .A(\cpu.genblk1.mmu.r_vtop_i[30][5] ),
    .B(net387));
 sg13g2_o21ai_1 _24726_ (.B1(_06324_),
    .Y(_01795_),
    .A1(_06255_),
    .A2(net304));
 sg13g2_nand2_1 _24727_ (.Y(_06325_),
    .A(\cpu.genblk1.mmu.r_vtop_i[30][6] ),
    .B(net387));
 sg13g2_o21ai_1 _24728_ (.B1(_06325_),
    .Y(_01796_),
    .A1(net729),
    .A2(net304));
 sg13g2_mux2_1 _24729_ (.A0(_06259_),
    .A1(\cpu.genblk1.mmu.r_vtop_i[30][7] ),
    .S(net304),
    .X(_01797_));
 sg13g2_mux2_1 _24730_ (.A0(net474),
    .A1(\cpu.genblk1.mmu.r_vtop_i[30][8] ),
    .S(_06317_),
    .X(_01798_));
 sg13g2_mux2_1 _24731_ (.A0(net443),
    .A1(\cpu.genblk1.mmu.r_vtop_i[30][9] ),
    .S(net387),
    .X(_01799_));
 sg13g2_nand3_1 _24732_ (.B(_06285_),
    .C(net476),
    .A(_05844_),
    .Y(_06326_));
 sg13g2_buf_1 _24733_ (.A(_06326_),
    .X(_06327_));
 sg13g2_buf_1 _24734_ (.A(net386),
    .X(_06328_));
 sg13g2_nand2_1 _24735_ (.Y(_06329_),
    .A(\cpu.genblk1.mmu.r_vtop_i[31][0] ),
    .B(net386));
 sg13g2_o21ai_1 _24736_ (.B1(_06329_),
    .Y(_01800_),
    .A1(net586),
    .A2(net303));
 sg13g2_mux2_1 _24737_ (.A0(net525),
    .A1(\cpu.genblk1.mmu.r_vtop_i[31][10] ),
    .S(net303),
    .X(_01801_));
 sg13g2_nand2_1 _24738_ (.Y(_06330_),
    .A(\cpu.genblk1.mmu.r_vtop_i[31][11] ),
    .B(_06327_));
 sg13g2_o21ai_1 _24739_ (.B1(_06330_),
    .Y(_01802_),
    .A1(net585),
    .A2(net303));
 sg13g2_nand2_1 _24740_ (.Y(_06331_),
    .A(\cpu.genblk1.mmu.r_vtop_i[31][1] ),
    .B(net386));
 sg13g2_o21ai_1 _24741_ (.B1(_06331_),
    .Y(_01803_),
    .A1(net733),
    .A2(net303));
 sg13g2_mux2_1 _24742_ (.A0(net732),
    .A1(\cpu.genblk1.mmu.r_vtop_i[31][2] ),
    .S(net303),
    .X(_01804_));
 sg13g2_nand2_1 _24743_ (.Y(_06332_),
    .A(\cpu.genblk1.mmu.r_vtop_i[31][3] ),
    .B(net386));
 sg13g2_o21ai_1 _24744_ (.B1(_06332_),
    .Y(_01805_),
    .A1(_06251_),
    .A2(net303));
 sg13g2_nand2_1 _24745_ (.Y(_06333_),
    .A(\cpu.genblk1.mmu.r_vtop_i[31][4] ),
    .B(net386));
 sg13g2_o21ai_1 _24746_ (.B1(_06333_),
    .Y(_01806_),
    .A1(net847),
    .A2(_06328_));
 sg13g2_nand2_1 _24747_ (.Y(_06334_),
    .A(\cpu.genblk1.mmu.r_vtop_i[31][5] ),
    .B(net386));
 sg13g2_o21ai_1 _24748_ (.B1(_06334_),
    .Y(_01807_),
    .A1(net730),
    .A2(_06328_));
 sg13g2_nand2_1 _24749_ (.Y(_06335_),
    .A(\cpu.genblk1.mmu.r_vtop_i[31][6] ),
    .B(net386));
 sg13g2_o21ai_1 _24750_ (.B1(_06335_),
    .Y(_01808_),
    .A1(net729),
    .A2(net303));
 sg13g2_mux2_1 _24751_ (.A0(_06259_),
    .A1(\cpu.genblk1.mmu.r_vtop_i[31][7] ),
    .S(net303),
    .X(_01809_));
 sg13g2_mux2_1 _24752_ (.A0(net474),
    .A1(\cpu.genblk1.mmu.r_vtop_i[31][8] ),
    .S(_06327_),
    .X(_01810_));
 sg13g2_mux2_1 _24753_ (.A0(net443),
    .A1(\cpu.genblk1.mmu.r_vtop_i[31][9] ),
    .S(net386),
    .X(_01811_));
 sg13g2_nand3_1 _24754_ (.B(_06046_),
    .C(net476),
    .A(_05844_),
    .Y(_06336_));
 sg13g2_buf_1 _24755_ (.A(_06336_),
    .X(_06337_));
 sg13g2_buf_1 _24756_ (.A(net385),
    .X(_06338_));
 sg13g2_nand2_1 _24757_ (.Y(_06339_),
    .A(\cpu.genblk1.mmu.r_vtop_i[3][0] ),
    .B(net385));
 sg13g2_o21ai_1 _24758_ (.B1(_06339_),
    .Y(_01812_),
    .A1(net586),
    .A2(net302));
 sg13g2_mux2_1 _24759_ (.A0(net525),
    .A1(\cpu.genblk1.mmu.r_vtop_i[3][10] ),
    .S(net302),
    .X(_01813_));
 sg13g2_nand2_1 _24760_ (.Y(_06340_),
    .A(\cpu.genblk1.mmu.r_vtop_i[3][11] ),
    .B(_06337_));
 sg13g2_o21ai_1 _24761_ (.B1(_06340_),
    .Y(_01814_),
    .A1(_06276_),
    .A2(net302));
 sg13g2_nand2_1 _24762_ (.Y(_06341_),
    .A(\cpu.genblk1.mmu.r_vtop_i[3][1] ),
    .B(net385));
 sg13g2_o21ai_1 _24763_ (.B1(_06341_),
    .Y(_01815_),
    .A1(_06248_),
    .A2(net302));
 sg13g2_mux2_1 _24764_ (.A0(net732),
    .A1(\cpu.genblk1.mmu.r_vtop_i[3][2] ),
    .S(net302),
    .X(_01816_));
 sg13g2_nand2_1 _24765_ (.Y(_06342_),
    .A(\cpu.genblk1.mmu.r_vtop_i[3][3] ),
    .B(net385));
 sg13g2_o21ai_1 _24766_ (.B1(_06342_),
    .Y(_01817_),
    .A1(net731),
    .A2(net302));
 sg13g2_nand2_1 _24767_ (.Y(_06343_),
    .A(\cpu.genblk1.mmu.r_vtop_i[3][4] ),
    .B(_06337_));
 sg13g2_o21ai_1 _24768_ (.B1(_06343_),
    .Y(_01818_),
    .A1(net847),
    .A2(_06338_));
 sg13g2_nand2_1 _24769_ (.Y(_06344_),
    .A(\cpu.genblk1.mmu.r_vtop_i[3][5] ),
    .B(net385));
 sg13g2_o21ai_1 _24770_ (.B1(_06344_),
    .Y(_01819_),
    .A1(net730),
    .A2(_06338_));
 sg13g2_nand2_1 _24771_ (.Y(_06345_),
    .A(\cpu.genblk1.mmu.r_vtop_i[3][6] ),
    .B(net385));
 sg13g2_o21ai_1 _24772_ (.B1(_06345_),
    .Y(_01820_),
    .A1(_06257_),
    .A2(net302));
 sg13g2_mux2_1 _24773_ (.A0(net846),
    .A1(\cpu.genblk1.mmu.r_vtop_i[3][7] ),
    .S(net302),
    .X(_01821_));
 sg13g2_mux2_1 _24774_ (.A0(net474),
    .A1(\cpu.genblk1.mmu.r_vtop_i[3][8] ),
    .S(net385),
    .X(_01822_));
 sg13g2_mux2_1 _24775_ (.A0(_06284_),
    .A1(\cpu.genblk1.mmu.r_vtop_i[3][9] ),
    .S(net385),
    .X(_01823_));
 sg13g2_nand2b_1 _24776_ (.Y(_06346_),
    .B(_06050_),
    .A_N(_06019_));
 sg13g2_buf_1 _24777_ (.A(_06346_),
    .X(_06347_));
 sg13g2_buf_1 _24778_ (.A(net301),
    .X(_06348_));
 sg13g2_nand2_1 _24779_ (.Y(_06349_),
    .A(\cpu.genblk1.mmu.r_vtop_i[4][0] ),
    .B(net301));
 sg13g2_o21ai_1 _24780_ (.B1(_06349_),
    .Y(_01824_),
    .A1(net586),
    .A2(net246));
 sg13g2_mux2_1 _24781_ (.A0(net525),
    .A1(\cpu.genblk1.mmu.r_vtop_i[4][10] ),
    .S(net246),
    .X(_01825_));
 sg13g2_nand2_1 _24782_ (.Y(_06350_),
    .A(\cpu.genblk1.mmu.r_vtop_i[4][11] ),
    .B(net301));
 sg13g2_o21ai_1 _24783_ (.B1(_06350_),
    .Y(_01826_),
    .A1(net585),
    .A2(net246));
 sg13g2_nand2_1 _24784_ (.Y(_06351_),
    .A(\cpu.genblk1.mmu.r_vtop_i[4][1] ),
    .B(net301));
 sg13g2_o21ai_1 _24785_ (.B1(_06351_),
    .Y(_01827_),
    .A1(_06248_),
    .A2(net246));
 sg13g2_mux2_1 _24786_ (.A0(_06250_),
    .A1(\cpu.genblk1.mmu.r_vtop_i[4][2] ),
    .S(net246),
    .X(_01828_));
 sg13g2_nand2_1 _24787_ (.Y(_06352_),
    .A(\cpu.genblk1.mmu.r_vtop_i[4][3] ),
    .B(net301));
 sg13g2_o21ai_1 _24788_ (.B1(_06352_),
    .Y(_01829_),
    .A1(net731),
    .A2(net246));
 sg13g2_nand2_1 _24789_ (.Y(_06353_),
    .A(\cpu.genblk1.mmu.r_vtop_i[4][4] ),
    .B(net301));
 sg13g2_o21ai_1 _24790_ (.B1(_06353_),
    .Y(_01830_),
    .A1(_06253_),
    .A2(_06348_));
 sg13g2_nand2_1 _24791_ (.Y(_06354_),
    .A(\cpu.genblk1.mmu.r_vtop_i[4][5] ),
    .B(_06347_));
 sg13g2_o21ai_1 _24792_ (.B1(_06354_),
    .Y(_01831_),
    .A1(net730),
    .A2(_06348_));
 sg13g2_nand2_1 _24793_ (.Y(_06355_),
    .A(\cpu.genblk1.mmu.r_vtop_i[4][6] ),
    .B(net301));
 sg13g2_o21ai_1 _24794_ (.B1(_06355_),
    .Y(_01832_),
    .A1(_06257_),
    .A2(net246));
 sg13g2_mux2_1 _24795_ (.A0(net846),
    .A1(\cpu.genblk1.mmu.r_vtop_i[4][7] ),
    .S(net246),
    .X(_01833_));
 sg13g2_mux2_1 _24796_ (.A0(net474),
    .A1(\cpu.genblk1.mmu.r_vtop_i[4][8] ),
    .S(_06347_),
    .X(_01834_));
 sg13g2_mux2_1 _24797_ (.A0(net443),
    .A1(\cpu.genblk1.mmu.r_vtop_i[4][9] ),
    .S(net301),
    .X(_01835_));
 sg13g2_nand2_1 _24798_ (.Y(_06356_),
    .A(_06024_),
    .B(net477));
 sg13g2_buf_1 _24799_ (.A(_06356_),
    .X(_06357_));
 sg13g2_buf_1 _24800_ (.A(net384),
    .X(_06358_));
 sg13g2_nand2_1 _24801_ (.Y(_06359_),
    .A(\cpu.genblk1.mmu.r_vtop_i[5][0] ),
    .B(net384));
 sg13g2_o21ai_1 _24802_ (.B1(_06359_),
    .Y(_01836_),
    .A1(_06270_),
    .A2(net300));
 sg13g2_mux2_1 _24803_ (.A0(_06275_),
    .A1(\cpu.genblk1.mmu.r_vtop_i[5][10] ),
    .S(net300),
    .X(_01837_));
 sg13g2_nand2_1 _24804_ (.Y(_06360_),
    .A(\cpu.genblk1.mmu.r_vtop_i[5][11] ),
    .B(net384));
 sg13g2_o21ai_1 _24805_ (.B1(_06360_),
    .Y(_01838_),
    .A1(net585),
    .A2(net300));
 sg13g2_nand2_1 _24806_ (.Y(_06361_),
    .A(\cpu.genblk1.mmu.r_vtop_i[5][1] ),
    .B(net384));
 sg13g2_o21ai_1 _24807_ (.B1(_06361_),
    .Y(_01839_),
    .A1(net873),
    .A2(_06358_));
 sg13g2_mux2_1 _24808_ (.A0(net748),
    .A1(\cpu.genblk1.mmu.r_vtop_i[5][2] ),
    .S(net300),
    .X(_01840_));
 sg13g2_nand2_1 _24809_ (.Y(_06362_),
    .A(\cpu.genblk1.mmu.r_vtop_i[5][3] ),
    .B(net384));
 sg13g2_o21ai_1 _24810_ (.B1(_06362_),
    .Y(_01841_),
    .A1(net871),
    .A2(net300));
 sg13g2_nand2_1 _24811_ (.Y(_06363_),
    .A(\cpu.genblk1.mmu.r_vtop_i[5][4] ),
    .B(net384));
 sg13g2_o21ai_1 _24812_ (.B1(_06363_),
    .Y(_01842_),
    .A1(net1037),
    .A2(net300));
 sg13g2_nand2_1 _24813_ (.Y(_06364_),
    .A(\cpu.genblk1.mmu.r_vtop_i[5][5] ),
    .B(net384));
 sg13g2_o21ai_1 _24814_ (.B1(_06364_),
    .Y(_01843_),
    .A1(net869),
    .A2(_06358_));
 sg13g2_nand2_1 _24815_ (.Y(_06365_),
    .A(\cpu.genblk1.mmu.r_vtop_i[5][6] ),
    .B(net384));
 sg13g2_o21ai_1 _24816_ (.B1(_06365_),
    .Y(_01844_),
    .A1(net889),
    .A2(net300));
 sg13g2_mux2_1 _24817_ (.A0(net863),
    .A1(\cpu.genblk1.mmu.r_vtop_i[5][7] ),
    .S(net300),
    .X(_01845_));
 sg13g2_mux2_1 _24818_ (.A0(_06283_),
    .A1(\cpu.genblk1.mmu.r_vtop_i[5][8] ),
    .S(_06357_),
    .X(_01846_));
 sg13g2_mux2_1 _24819_ (.A0(net443),
    .A1(\cpu.genblk1.mmu.r_vtop_i[5][9] ),
    .S(_06357_),
    .X(_01847_));
 sg13g2_nand2_1 _24820_ (.Y(_06366_),
    .A(_06030_),
    .B(net477));
 sg13g2_buf_1 _24821_ (.A(_06366_),
    .X(_06367_));
 sg13g2_buf_1 _24822_ (.A(net383),
    .X(_06368_));
 sg13g2_nand2_1 _24823_ (.Y(_06369_),
    .A(\cpu.genblk1.mmu.r_vtop_i[6][0] ),
    .B(net383));
 sg13g2_o21ai_1 _24824_ (.B1(_06369_),
    .Y(_01848_),
    .A1(_06270_),
    .A2(net299));
 sg13g2_mux2_1 _24825_ (.A0(_06275_),
    .A1(\cpu.genblk1.mmu.r_vtop_i[6][10] ),
    .S(net299),
    .X(_01849_));
 sg13g2_nand2_1 _24826_ (.Y(_06370_),
    .A(\cpu.genblk1.mmu.r_vtop_i[6][11] ),
    .B(net383));
 sg13g2_o21ai_1 _24827_ (.B1(_06370_),
    .Y(_01850_),
    .A1(net585),
    .A2(net299));
 sg13g2_nand2_1 _24828_ (.Y(_06371_),
    .A(\cpu.genblk1.mmu.r_vtop_i[6][1] ),
    .B(net383));
 sg13g2_o21ai_1 _24829_ (.B1(_06371_),
    .Y(_01851_),
    .A1(net873),
    .A2(_06368_));
 sg13g2_mux2_1 _24830_ (.A0(net748),
    .A1(\cpu.genblk1.mmu.r_vtop_i[6][2] ),
    .S(net299),
    .X(_01852_));
 sg13g2_nand2_1 _24831_ (.Y(_06372_),
    .A(\cpu.genblk1.mmu.r_vtop_i[6][3] ),
    .B(net383));
 sg13g2_o21ai_1 _24832_ (.B1(_06372_),
    .Y(_01853_),
    .A1(net871),
    .A2(net299));
 sg13g2_nand2_1 _24833_ (.Y(_06373_),
    .A(\cpu.genblk1.mmu.r_vtop_i[6][4] ),
    .B(net383));
 sg13g2_o21ai_1 _24834_ (.B1(_06373_),
    .Y(_01854_),
    .A1(net1037),
    .A2(net299));
 sg13g2_nand2_1 _24835_ (.Y(_06374_),
    .A(\cpu.genblk1.mmu.r_vtop_i[6][5] ),
    .B(net383));
 sg13g2_o21ai_1 _24836_ (.B1(_06374_),
    .Y(_01855_),
    .A1(net869),
    .A2(_06368_));
 sg13g2_nand2_1 _24837_ (.Y(_06375_),
    .A(\cpu.genblk1.mmu.r_vtop_i[6][6] ),
    .B(net383));
 sg13g2_o21ai_1 _24838_ (.B1(_06375_),
    .Y(_01856_),
    .A1(net889),
    .A2(net299));
 sg13g2_mux2_1 _24839_ (.A0(net863),
    .A1(\cpu.genblk1.mmu.r_vtop_i[6][7] ),
    .S(net299),
    .X(_01857_));
 sg13g2_mux2_1 _24840_ (.A0(_06283_),
    .A1(\cpu.genblk1.mmu.r_vtop_i[6][8] ),
    .S(_06367_),
    .X(_01858_));
 sg13g2_mux2_1 _24841_ (.A0(_06284_),
    .A1(\cpu.genblk1.mmu.r_vtop_i[6][9] ),
    .S(_06367_),
    .X(_01859_));
 sg13g2_nand2_1 _24842_ (.Y(_06376_),
    .A(_06035_),
    .B(_06061_));
 sg13g2_buf_1 _24843_ (.A(_06376_),
    .X(_06377_));
 sg13g2_buf_1 _24844_ (.A(net298),
    .X(_06378_));
 sg13g2_nand2_1 _24845_ (.Y(_06379_),
    .A(\cpu.genblk1.mmu.r_vtop_i[7][0] ),
    .B(net298));
 sg13g2_o21ai_1 _24846_ (.B1(_06379_),
    .Y(_01860_),
    .A1(net666),
    .A2(net245));
 sg13g2_mux2_1 _24847_ (.A0(net551),
    .A1(\cpu.genblk1.mmu.r_vtop_i[7][10] ),
    .S(net245),
    .X(_01861_));
 sg13g2_nand2_1 _24848_ (.Y(_06380_),
    .A(\cpu.genblk1.mmu.r_vtop_i[7][11] ),
    .B(net298));
 sg13g2_o21ai_1 _24849_ (.B1(_06380_),
    .Y(_01862_),
    .A1(net699),
    .A2(net245));
 sg13g2_nand2_1 _24850_ (.Y(_06381_),
    .A(\cpu.genblk1.mmu.r_vtop_i[7][1] ),
    .B(net298));
 sg13g2_o21ai_1 _24851_ (.B1(_06381_),
    .Y(_01863_),
    .A1(net873),
    .A2(_06378_));
 sg13g2_mux2_1 _24852_ (.A0(net748),
    .A1(\cpu.genblk1.mmu.r_vtop_i[7][2] ),
    .S(net245),
    .X(_01864_));
 sg13g2_nand2_1 _24853_ (.Y(_06382_),
    .A(\cpu.genblk1.mmu.r_vtop_i[7][3] ),
    .B(net298));
 sg13g2_o21ai_1 _24854_ (.B1(_06382_),
    .Y(_01865_),
    .A1(net871),
    .A2(net245));
 sg13g2_nand2_1 _24855_ (.Y(_06383_),
    .A(\cpu.genblk1.mmu.r_vtop_i[7][4] ),
    .B(_06377_));
 sg13g2_o21ai_1 _24856_ (.B1(_06383_),
    .Y(_01866_),
    .A1(net1037),
    .A2(net245));
 sg13g2_nand2_1 _24857_ (.Y(_06384_),
    .A(\cpu.genblk1.mmu.r_vtop_i[7][5] ),
    .B(net298));
 sg13g2_o21ai_1 _24858_ (.B1(_06384_),
    .Y(_01867_),
    .A1(net869),
    .A2(_06378_));
 sg13g2_nand2_1 _24859_ (.Y(_06385_),
    .A(\cpu.genblk1.mmu.r_vtop_i[7][6] ),
    .B(net298));
 sg13g2_o21ai_1 _24860_ (.B1(_06385_),
    .Y(_01868_),
    .A1(net889),
    .A2(net245));
 sg13g2_mux2_1 _24861_ (.A0(net863),
    .A1(\cpu.genblk1.mmu.r_vtop_i[7][7] ),
    .S(net245),
    .X(_01869_));
 sg13g2_mux2_1 _24862_ (.A0(_03500_),
    .A1(\cpu.genblk1.mmu.r_vtop_i[7][8] ),
    .S(net298),
    .X(_01870_));
 sg13g2_mux2_1 _24863_ (.A0(net454),
    .A1(\cpu.genblk1.mmu.r_vtop_i[7][9] ),
    .S(_06377_),
    .X(_01871_));
 sg13g2_nor2_1 _24864_ (.A(net965),
    .B(net1044),
    .Y(_06386_));
 sg13g2_nand3_1 _24865_ (.B(_06128_),
    .C(_06116_),
    .A(_06386_),
    .Y(_06387_));
 sg13g2_buf_1 _24866_ (.A(_06387_),
    .X(_06388_));
 sg13g2_buf_1 _24867_ (.A(net382),
    .X(_06389_));
 sg13g2_nand2_1 _24868_ (.Y(_06390_),
    .A(\cpu.genblk1.mmu.r_vtop_i[8][0] ),
    .B(net382));
 sg13g2_o21ai_1 _24869_ (.B1(_06390_),
    .Y(_01872_),
    .A1(net666),
    .A2(net297));
 sg13g2_mux2_1 _24870_ (.A0(net551),
    .A1(\cpu.genblk1.mmu.r_vtop_i[8][10] ),
    .S(net297),
    .X(_01873_));
 sg13g2_nand2_1 _24871_ (.Y(_06391_),
    .A(\cpu.genblk1.mmu.r_vtop_i[8][11] ),
    .B(net382));
 sg13g2_o21ai_1 _24872_ (.B1(_06391_),
    .Y(_01874_),
    .A1(net699),
    .A2(net297));
 sg13g2_nand2_1 _24873_ (.Y(_06392_),
    .A(\cpu.genblk1.mmu.r_vtop_i[8][1] ),
    .B(net382));
 sg13g2_o21ai_1 _24874_ (.B1(_06392_),
    .Y(_01875_),
    .A1(net873),
    .A2(net297));
 sg13g2_mux2_1 _24875_ (.A0(net748),
    .A1(\cpu.genblk1.mmu.r_vtop_i[8][2] ),
    .S(net297),
    .X(_01876_));
 sg13g2_nand2_1 _24876_ (.Y(_06393_),
    .A(\cpu.genblk1.mmu.r_vtop_i[8][3] ),
    .B(net382));
 sg13g2_o21ai_1 _24877_ (.B1(_06393_),
    .Y(_01877_),
    .A1(net871),
    .A2(net297));
 sg13g2_nand2_1 _24878_ (.Y(_06394_),
    .A(\cpu.genblk1.mmu.r_vtop_i[8][4] ),
    .B(_06388_));
 sg13g2_o21ai_1 _24879_ (.B1(_06394_),
    .Y(_01878_),
    .A1(net1037),
    .A2(_06389_));
 sg13g2_nand2_1 _24880_ (.Y(_06395_),
    .A(\cpu.genblk1.mmu.r_vtop_i[8][5] ),
    .B(net382));
 sg13g2_o21ai_1 _24881_ (.B1(_06395_),
    .Y(_01879_),
    .A1(net869),
    .A2(_06389_));
 sg13g2_nand2_1 _24882_ (.Y(_06396_),
    .A(\cpu.genblk1.mmu.r_vtop_i[8][6] ),
    .B(net382));
 sg13g2_o21ai_1 _24883_ (.B1(_06396_),
    .Y(_01880_),
    .A1(net889),
    .A2(net297));
 sg13g2_mux2_1 _24884_ (.A0(net863),
    .A1(\cpu.genblk1.mmu.r_vtop_i[8][7] ),
    .S(net297),
    .X(_01881_));
 sg13g2_mux2_1 _24885_ (.A0(net494),
    .A1(\cpu.genblk1.mmu.r_vtop_i[8][8] ),
    .S(net382),
    .X(_01882_));
 sg13g2_mux2_1 _24886_ (.A0(net454),
    .A1(\cpu.genblk1.mmu.r_vtop_i[8][9] ),
    .S(_06388_),
    .X(_01883_));
 sg13g2_nand3_1 _24887_ (.B(_06386_),
    .C(_06094_),
    .A(net978),
    .Y(_06397_));
 sg13g2_buf_1 _24888_ (.A(_06397_),
    .X(_06398_));
 sg13g2_buf_1 _24889_ (.A(net296),
    .X(_06399_));
 sg13g2_nand2_1 _24890_ (.Y(_06400_),
    .A(\cpu.genblk1.mmu.r_vtop_i[9][0] ),
    .B(net296));
 sg13g2_o21ai_1 _24891_ (.B1(_06400_),
    .Y(_01884_),
    .A1(_03838_),
    .A2(net244));
 sg13g2_mux2_1 _24892_ (.A0(net551),
    .A1(\cpu.genblk1.mmu.r_vtop_i[9][10] ),
    .S(net244),
    .X(_01885_));
 sg13g2_nand2_1 _24893_ (.Y(_06401_),
    .A(\cpu.genblk1.mmu.r_vtop_i[9][11] ),
    .B(net296));
 sg13g2_o21ai_1 _24894_ (.B1(_06401_),
    .Y(_01886_),
    .A1(net699),
    .A2(net244));
 sg13g2_nand2_1 _24895_ (.Y(_06402_),
    .A(\cpu.genblk1.mmu.r_vtop_i[9][1] ),
    .B(net296));
 sg13g2_o21ai_1 _24896_ (.B1(_06402_),
    .Y(_01887_),
    .A1(net873),
    .A2(net244));
 sg13g2_mux2_1 _24897_ (.A0(net748),
    .A1(\cpu.genblk1.mmu.r_vtop_i[9][2] ),
    .S(net244),
    .X(_01888_));
 sg13g2_nand2_1 _24898_ (.Y(_06403_),
    .A(\cpu.genblk1.mmu.r_vtop_i[9][3] ),
    .B(net296));
 sg13g2_o21ai_1 _24899_ (.B1(_06403_),
    .Y(_01889_),
    .A1(net871),
    .A2(net244));
 sg13g2_nand2_1 _24900_ (.Y(_06404_),
    .A(\cpu.genblk1.mmu.r_vtop_i[9][4] ),
    .B(_06398_));
 sg13g2_o21ai_1 _24901_ (.B1(_06404_),
    .Y(_01890_),
    .A1(net1037),
    .A2(_06399_));
 sg13g2_nand2_1 _24902_ (.Y(_06405_),
    .A(\cpu.genblk1.mmu.r_vtop_i[9][5] ),
    .B(net296));
 sg13g2_o21ai_1 _24903_ (.B1(_06405_),
    .Y(_01891_),
    .A1(net869),
    .A2(_06399_));
 sg13g2_nand2_1 _24904_ (.Y(_06406_),
    .A(\cpu.genblk1.mmu.r_vtop_i[9][6] ),
    .B(net296));
 sg13g2_o21ai_1 _24905_ (.B1(_06406_),
    .Y(_01892_),
    .A1(net889),
    .A2(net244));
 sg13g2_mux2_1 _24906_ (.A0(net863),
    .A1(\cpu.genblk1.mmu.r_vtop_i[9][7] ),
    .S(net244),
    .X(_01893_));
 sg13g2_mux2_1 _24907_ (.A0(_03500_),
    .A1(\cpu.genblk1.mmu.r_vtop_i[9][8] ),
    .S(net296),
    .X(_01894_));
 sg13g2_mux2_1 _24908_ (.A0(net454),
    .A1(\cpu.genblk1.mmu.r_vtop_i[9][9] ),
    .S(_06398_),
    .X(_01895_));
 sg13g2_buf_1 _24909_ (.A(net491),
    .X(_06407_));
 sg13g2_mux2_1 _24910_ (.A0(\cpu.genblk1.mmu.r_writeable_d[0] ),
    .A1(net442),
    .S(_05886_),
    .X(_01896_));
 sg13g2_mux2_1 _24911_ (.A0(\cpu.genblk1.mmu.r_writeable_d[10] ),
    .A1(net442),
    .S(_05897_),
    .X(_01897_));
 sg13g2_mux2_1 _24912_ (.A0(\cpu.genblk1.mmu.r_writeable_d[11] ),
    .A1(net442),
    .S(_05902_),
    .X(_01898_));
 sg13g2_mux2_1 _24913_ (.A0(\cpu.genblk1.mmu.r_writeable_d[12] ),
    .A1(net442),
    .S(_05907_),
    .X(_01899_));
 sg13g2_mux2_1 _24914_ (.A0(\cpu.genblk1.mmu.r_writeable_d[13] ),
    .A1(net442),
    .S(_05913_),
    .X(_01900_));
 sg13g2_mux2_1 _24915_ (.A0(\cpu.genblk1.mmu.r_writeable_d[14] ),
    .A1(_06407_),
    .S(_05918_),
    .X(_01901_));
 sg13g2_mux2_1 _24916_ (.A0(\cpu.genblk1.mmu.r_writeable_d[15] ),
    .A1(_06407_),
    .S(_05925_),
    .X(_01902_));
 sg13g2_mux2_1 _24917_ (.A0(\cpu.genblk1.mmu.r_writeable_d[16] ),
    .A1(net442),
    .S(_05931_),
    .X(_01903_));
 sg13g2_mux2_1 _24918_ (.A0(\cpu.genblk1.mmu.r_writeable_d[17] ),
    .A1(net442),
    .S(_05936_),
    .X(_01904_));
 sg13g2_mux2_1 _24919_ (.A0(\cpu.genblk1.mmu.r_writeable_d[18] ),
    .A1(net442),
    .S(_05941_),
    .X(_01905_));
 sg13g2_buf_1 _24920_ (.A(net491),
    .X(_06408_));
 sg13g2_mux2_1 _24921_ (.A0(\cpu.genblk1.mmu.r_writeable_d[19] ),
    .A1(net441),
    .S(_05949_),
    .X(_01906_));
 sg13g2_mux2_1 _24922_ (.A0(\cpu.genblk1.mmu.r_writeable_d[1] ),
    .A1(net441),
    .S(_05954_),
    .X(_01907_));
 sg13g2_mux2_1 _24923_ (.A0(\cpu.genblk1.mmu.r_writeable_d[20] ),
    .A1(net441),
    .S(_05959_),
    .X(_01908_));
 sg13g2_mux2_1 _24924_ (.A0(\cpu.genblk1.mmu.r_writeable_d[21] ),
    .A1(net441),
    .S(_05962_),
    .X(_01909_));
 sg13g2_mux2_1 _24925_ (.A0(\cpu.genblk1.mmu.r_writeable_d[22] ),
    .A1(_06408_),
    .S(_05965_),
    .X(_01910_));
 sg13g2_mux2_1 _24926_ (.A0(\cpu.genblk1.mmu.r_writeable_d[23] ),
    .A1(net441),
    .S(_05969_),
    .X(_01911_));
 sg13g2_mux2_1 _24927_ (.A0(\cpu.genblk1.mmu.r_writeable_d[24] ),
    .A1(net441),
    .S(_05978_),
    .X(_01912_));
 sg13g2_mux2_1 _24928_ (.A0(\cpu.genblk1.mmu.r_writeable_d[25] ),
    .A1(net441),
    .S(_05981_),
    .X(_01913_));
 sg13g2_mux2_1 _24929_ (.A0(\cpu.genblk1.mmu.r_writeable_d[26] ),
    .A1(net441),
    .S(_05987_),
    .X(_01914_));
 sg13g2_mux2_1 _24930_ (.A0(\cpu.genblk1.mmu.r_writeable_d[27] ),
    .A1(_06408_),
    .S(_05992_),
    .X(_01915_));
 sg13g2_buf_1 _24931_ (.A(net491),
    .X(_06409_));
 sg13g2_mux2_1 _24932_ (.A0(\cpu.genblk1.mmu.r_writeable_d[28] ),
    .A1(net440),
    .S(_06000_),
    .X(_01916_));
 sg13g2_mux2_1 _24933_ (.A0(\cpu.genblk1.mmu.r_writeable_d[29] ),
    .A1(net440),
    .S(_06005_),
    .X(_01917_));
 sg13g2_mux2_1 _24934_ (.A0(\cpu.genblk1.mmu.r_writeable_d[2] ),
    .A1(_06409_),
    .S(_06008_),
    .X(_01918_));
 sg13g2_mux2_1 _24935_ (.A0(\cpu.genblk1.mmu.r_writeable_d[30] ),
    .A1(net440),
    .S(_06011_),
    .X(_01919_));
 sg13g2_mux2_1 _24936_ (.A0(\cpu.genblk1.mmu.r_writeable_d[31] ),
    .A1(net440),
    .S(_06014_),
    .X(_01920_));
 sg13g2_mux2_1 _24937_ (.A0(\cpu.genblk1.mmu.r_writeable_d[3] ),
    .A1(net440),
    .S(_06017_),
    .X(_01921_));
 sg13g2_mux2_1 _24938_ (.A0(\cpu.genblk1.mmu.r_writeable_d[4] ),
    .A1(net440),
    .S(_06021_),
    .X(_01922_));
 sg13g2_mux2_1 _24939_ (.A0(\cpu.genblk1.mmu.r_writeable_d[5] ),
    .A1(net440),
    .S(_06026_),
    .X(_01923_));
 sg13g2_mux2_1 _24940_ (.A0(\cpu.genblk1.mmu.r_writeable_d[6] ),
    .A1(_06409_),
    .S(_06032_),
    .X(_01924_));
 sg13g2_mux2_1 _24941_ (.A0(\cpu.genblk1.mmu.r_writeable_d[7] ),
    .A1(net440),
    .S(_06037_),
    .X(_01925_));
 sg13g2_mux2_1 _24942_ (.A0(\cpu.genblk1.mmu.r_writeable_d[8] ),
    .A1(_03509_),
    .S(_06040_),
    .X(_01926_));
 sg13g2_mux2_1 _24943_ (.A0(\cpu.genblk1.mmu.r_writeable_d[9] ),
    .A1(_03509_),
    .S(_06043_),
    .X(_01927_));
 sg13g2_inv_1 _24944_ (.Y(_06410_),
    .A(_00219_));
 sg13g2_nor4_1 _24945_ (.A(net1000),
    .B(_09223_),
    .C(_06410_),
    .D(_09246_),
    .Y(_06411_));
 sg13g2_buf_1 _24946_ (.A(_06411_),
    .X(_06412_));
 sg13g2_and2_1 _24947_ (.A(net928),
    .B(net112),
    .X(_06413_));
 sg13g2_buf_2 _24948_ (.A(_06413_),
    .X(_06414_));
 sg13g2_and2_1 _24949_ (.A(_05689_),
    .B(_06414_),
    .X(_06415_));
 sg13g2_buf_1 _24950_ (.A(_06415_),
    .X(_06416_));
 sg13g2_mux2_1 _24951_ (.A0(\cpu.gpio.genblk2[4].srcs_io[0] ),
    .A1(_10067_),
    .S(_06416_),
    .X(_01944_));
 sg13g2_mux2_1 _24952_ (.A0(\cpu.gpio.genblk2[5].srcs_io[0] ),
    .A1(net1058),
    .S(_06416_),
    .X(_01945_));
 sg13g2_mux2_1 _24953_ (.A0(\cpu.gpio.genblk2[6].srcs_io[0] ),
    .A1(net1057),
    .S(_06416_),
    .X(_01946_));
 sg13g2_mux2_1 _24954_ (.A0(\cpu.gpio.genblk2[7].srcs_io[0] ),
    .A1(net1023),
    .S(_06416_),
    .X(_01947_));
 sg13g2_buf_1 _24955_ (.A(net1128),
    .X(_06417_));
 sg13g2_nand3_1 _24956_ (.B(_10095_),
    .C(_06414_),
    .A(_04980_),
    .Y(_06418_));
 sg13g2_buf_2 _24957_ (.A(_06418_),
    .X(_06419_));
 sg13g2_mux2_1 _24958_ (.A0(net964),
    .A1(\cpu.gpio.genblk1[3].srcs_o[0] ),
    .S(_06419_),
    .X(_01948_));
 sg13g2_nand2_1 _24959_ (.Y(_06420_),
    .A(\cpu.gpio.genblk1[4].srcs_o[0] ),
    .B(_06419_));
 sg13g2_o21ai_1 _24960_ (.B1(_06420_),
    .Y(_01949_),
    .A1(net877),
    .A2(_06419_));
 sg13g2_nand2_1 _24961_ (.Y(_06421_),
    .A(\cpu.gpio.genblk1[5].srcs_o[0] ),
    .B(_06419_));
 sg13g2_o21ai_1 _24962_ (.B1(_06421_),
    .Y(_01950_),
    .A1(net876),
    .A2(_06419_));
 sg13g2_nand2_1 _24963_ (.Y(_06422_),
    .A(\cpu.gpio.genblk1[6].srcs_o[0] ),
    .B(_06419_));
 sg13g2_o21ai_1 _24964_ (.B1(_06422_),
    .Y(_01951_),
    .A1(net875),
    .A2(_06419_));
 sg13g2_mux2_1 _24965_ (.A0(net1056),
    .A1(\cpu.gpio.genblk1[7].srcs_o[0] ),
    .S(_06419_),
    .X(_01952_));
 sg13g2_nand2_1 _24966_ (.Y(_06423_),
    .A(_04924_),
    .B(_06414_));
 sg13g2_buf_1 _24967_ (.A(_06423_),
    .X(_06424_));
 sg13g2_mux2_1 _24968_ (.A0(net913),
    .A1(_04923_),
    .S(_06424_),
    .X(_01953_));
 sg13g2_buf_1 _24969_ (.A(\cpu.gpio.r_spi_miso_src[0][1] ),
    .X(_06425_));
 sg13g2_mux2_1 _24970_ (.A0(net853),
    .A1(_06425_),
    .S(net74),
    .X(_01954_));
 sg13g2_buf_1 _24971_ (.A(net1060),
    .X(_06426_));
 sg13g2_mux2_1 _24972_ (.A0(_06426_),
    .A1(\cpu.gpio.r_spi_miso_src[0][2] ),
    .S(net74),
    .X(_01955_));
 sg13g2_buf_1 _24973_ (.A(\cpu.gpio.r_spi_miso_src[0][3] ),
    .X(_06427_));
 sg13g2_mux2_1 _24974_ (.A0(net964),
    .A1(_06427_),
    .S(net74),
    .X(_01956_));
 sg13g2_nand2_1 _24975_ (.Y(_06428_),
    .A(_05550_),
    .B(net74));
 sg13g2_o21ai_1 _24976_ (.B1(_06428_),
    .Y(_01957_),
    .A1(_12761_),
    .A2(net74));
 sg13g2_nand2_1 _24977_ (.Y(_06429_),
    .A(\cpu.gpio.r_spi_miso_src[1][1] ),
    .B(net74));
 sg13g2_o21ai_1 _24978_ (.B1(_06429_),
    .Y(_01958_),
    .A1(_12766_),
    .A2(net74));
 sg13g2_nand2_1 _24979_ (.Y(_06430_),
    .A(\cpu.gpio.r_spi_miso_src[1][2] ),
    .B(_06423_));
 sg13g2_o21ai_1 _24980_ (.B1(_06430_),
    .Y(_01959_),
    .A1(_12769_),
    .A2(net74));
 sg13g2_buf_1 _24981_ (.A(\cpu.gpio.r_spi_miso_src[1][3] ),
    .X(_06431_));
 sg13g2_mux2_1 _24982_ (.A0(net1056),
    .A1(_06431_),
    .S(_06424_),
    .X(_01960_));
 sg13g2_nand3_1 _24983_ (.B(net486),
    .C(_06414_),
    .A(net622),
    .Y(_06432_));
 sg13g2_buf_1 _24984_ (.A(_06432_),
    .X(_06433_));
 sg13g2_buf_1 _24985_ (.A(_06433_),
    .X(_06434_));
 sg13g2_mux2_1 _24986_ (.A0(_10034_),
    .A1(_04915_),
    .S(net34),
    .X(_01961_));
 sg13g2_mux2_1 _24987_ (.A0(net853),
    .A1(_05354_),
    .S(net34),
    .X(_01962_));
 sg13g2_mux2_1 _24988_ (.A0(_06426_),
    .A1(_05421_),
    .S(_06434_),
    .X(_01963_));
 sg13g2_mux2_1 _24989_ (.A0(_06417_),
    .A1(_05493_),
    .S(net34),
    .X(_01964_));
 sg13g2_nand2_1 _24990_ (.Y(_06435_),
    .A(_05554_),
    .B(net34));
 sg13g2_o21ai_1 _24991_ (.B1(_06435_),
    .Y(_01965_),
    .A1(net877),
    .A2(net34));
 sg13g2_nand2_1 _24992_ (.Y(_06436_),
    .A(_05615_),
    .B(net34));
 sg13g2_o21ai_1 _24993_ (.B1(_06436_),
    .Y(_01966_),
    .A1(_12145_),
    .A2(net34));
 sg13g2_nand2_1 _24994_ (.Y(_06437_),
    .A(_05683_),
    .B(_06433_));
 sg13g2_o21ai_1 _24995_ (.B1(_06437_),
    .Y(_01967_),
    .A1(_12769_),
    .A2(net34));
 sg13g2_mux2_1 _24996_ (.A0(net1056),
    .A1(_05094_),
    .S(_06434_),
    .X(_01968_));
 sg13g2_and3_1 _24997_ (.X(_06438_),
    .A(net550),
    .B(net486),
    .C(_06414_));
 sg13g2_buf_4 _24998_ (.X(_06439_),
    .A(_06438_));
 sg13g2_mux2_1 _24999_ (.A0(_04916_),
    .A1(net911),
    .S(_06439_),
    .X(_01969_));
 sg13g2_buf_1 _25000_ (.A(\cpu.gpio.r_src_io[6][1] ),
    .X(_06440_));
 sg13g2_mux2_1 _25001_ (.A0(_06440_),
    .A1(net885),
    .S(_06439_),
    .X(_01970_));
 sg13g2_mux2_1 _25002_ (.A0(\cpu.gpio.r_src_io[6][2] ),
    .A1(net884),
    .S(_06439_),
    .X(_01971_));
 sg13g2_mux2_1 _25003_ (.A0(\cpu.gpio.r_src_io[6][3] ),
    .A1(net1024),
    .S(_06439_),
    .X(_01972_));
 sg13g2_mux2_1 _25004_ (.A0(_05555_),
    .A1(net1059),
    .S(_06439_),
    .X(_01973_));
 sg13g2_buf_1 _25005_ (.A(\cpu.gpio.r_src_io[7][1] ),
    .X(_06441_));
 sg13g2_mux2_1 _25006_ (.A0(_06441_),
    .A1(net1058),
    .S(_06439_),
    .X(_01974_));
 sg13g2_mux2_1 _25007_ (.A0(\cpu.gpio.r_src_io[7][2] ),
    .A1(net1057),
    .S(_06439_),
    .X(_01975_));
 sg13g2_mux2_1 _25008_ (.A0(\cpu.gpio.r_src_io[7][3] ),
    .A1(net1018),
    .S(_06439_),
    .X(_01976_));
 sg13g2_and3_1 _25009_ (.X(_06442_),
    .A(_02975_),
    .B(_04955_),
    .C(_06414_));
 sg13g2_buf_2 _25010_ (.A(_06442_),
    .X(_06443_));
 sg13g2_nand2_1 _25011_ (.Y(_06444_),
    .A(net1059),
    .B(_06443_));
 sg13g2_o21ai_1 _25012_ (.B1(_06444_),
    .Y(_01977_),
    .A1(_05561_),
    .A2(_06443_));
 sg13g2_buf_1 _25013_ (.A(\cpu.gpio.r_src_o[3][1] ),
    .X(_06445_));
 sg13g2_mux2_1 _25014_ (.A0(_06445_),
    .A1(net1058),
    .S(_06443_),
    .X(_01978_));
 sg13g2_mux2_1 _25015_ (.A0(\cpu.gpio.r_src_o[3][2] ),
    .A1(_10079_),
    .S(_06443_),
    .X(_01979_));
 sg13g2_mux2_1 _25016_ (.A0(\cpu.gpio.r_src_o[3][3] ),
    .A1(net1018),
    .S(_06443_),
    .X(_01980_));
 sg13g2_nand2_1 _25017_ (.Y(_06446_),
    .A(_04905_),
    .B(_06414_));
 sg13g2_buf_1 _25018_ (.A(_06446_),
    .X(_06447_));
 sg13g2_mux2_1 _25019_ (.A0(_10034_),
    .A1(_04901_),
    .S(net73),
    .X(_01981_));
 sg13g2_buf_1 _25020_ (.A(\cpu.gpio.r_src_o[4][1] ),
    .X(_06448_));
 sg13g2_mux2_1 _25021_ (.A0(_05807_),
    .A1(_06448_),
    .S(net73),
    .X(_01982_));
 sg13g2_mux2_1 _25022_ (.A0(net845),
    .A1(\cpu.gpio.r_src_o[4][2] ),
    .S(net73),
    .X(_01983_));
 sg13g2_mux2_1 _25023_ (.A0(_06417_),
    .A1(\cpu.gpio.r_src_o[4][3] ),
    .S(net73),
    .X(_01984_));
 sg13g2_nand2_1 _25024_ (.Y(_06449_),
    .A(_05564_),
    .B(net73));
 sg13g2_o21ai_1 _25025_ (.B1(_06449_),
    .Y(_01985_),
    .A1(_12137_),
    .A2(net73));
 sg13g2_buf_1 _25026_ (.A(\cpu.gpio.r_src_o[5][1] ),
    .X(_06450_));
 sg13g2_nand2_1 _25027_ (.Y(_06451_),
    .A(_06450_),
    .B(net73));
 sg13g2_o21ai_1 _25028_ (.B1(_06451_),
    .Y(_01986_),
    .A1(_12145_),
    .A2(net73));
 sg13g2_nand2_1 _25029_ (.Y(_06452_),
    .A(\cpu.gpio.r_src_o[5][2] ),
    .B(_06446_));
 sg13g2_o21ai_1 _25030_ (.B1(_06452_),
    .Y(_01987_),
    .A1(_12150_),
    .A2(_06447_));
 sg13g2_mux2_1 _25031_ (.A0(_10082_),
    .A1(\cpu.gpio.r_src_o[5][3] ),
    .S(_06447_),
    .X(_01988_));
 sg13g2_nand2_1 _25032_ (.Y(_06453_),
    .A(net408),
    .B(_06414_));
 sg13g2_buf_2 _25033_ (.A(_06453_),
    .X(_06454_));
 sg13g2_nand2_1 _25034_ (.Y(_06455_),
    .A(_05559_),
    .B(_06454_));
 sg13g2_o21ai_1 _25035_ (.B1(_06455_),
    .Y(_01993_),
    .A1(_12137_),
    .A2(_06454_));
 sg13g2_buf_1 _25036_ (.A(\cpu.gpio.r_src_o[7][1] ),
    .X(_06456_));
 sg13g2_nand2_1 _25037_ (.Y(_06457_),
    .A(_06456_),
    .B(_06454_));
 sg13g2_o21ai_1 _25038_ (.B1(_06457_),
    .Y(_01994_),
    .A1(net882),
    .A2(_06454_));
 sg13g2_nand2_1 _25039_ (.Y(_06458_),
    .A(\cpu.gpio.r_src_o[7][2] ),
    .B(_06454_));
 sg13g2_o21ai_1 _25040_ (.B1(_06458_),
    .Y(_01995_),
    .A1(_12150_),
    .A2(_06454_));
 sg13g2_mux2_1 _25041_ (.A0(_10082_),
    .A1(\cpu.gpio.r_src_o[7][3] ),
    .S(_06454_),
    .X(_01996_));
 sg13g2_buf_1 _25042_ (.A(net1004),
    .X(_06459_));
 sg13g2_and2_1 _25043_ (.A(_08536_),
    .B(_08734_),
    .X(_06460_));
 sg13g2_buf_4 _25044_ (.X(_06461_),
    .A(_06460_));
 sg13g2_buf_1 _25045_ (.A(_00237_),
    .X(_06462_));
 sg13g2_nor2_1 _25046_ (.A(\cpu.icache.r_offset[2] ),
    .B(_06462_),
    .Y(_06463_));
 sg13g2_buf_2 _25047_ (.A(_06463_),
    .X(_06464_));
 sg13g2_buf_1 _25048_ (.A(\cpu.icache.r_offset[1] ),
    .X(_06465_));
 sg13g2_buf_1 _25049_ (.A(\cpu.icache.r_offset[0] ),
    .X(_06466_));
 sg13g2_nor2b_1 _25050_ (.A(_06465_),
    .B_N(_06466_),
    .Y(_06467_));
 sg13g2_buf_1 _25051_ (.A(_06467_),
    .X(_06468_));
 sg13g2_and2_1 _25052_ (.A(_06464_),
    .B(_06468_),
    .X(_06469_));
 sg13g2_buf_2 _25053_ (.A(_06469_),
    .X(_06470_));
 sg13g2_nand2_2 _25054_ (.Y(_06471_),
    .A(_06461_),
    .B(_06470_));
 sg13g2_mux2_1 _25055_ (.A0(net844),
    .A1(\cpu.icache.r_data[0][0] ),
    .S(_06471_),
    .X(_02000_));
 sg13g2_buf_1 _25056_ (.A(net1003),
    .X(_06472_));
 sg13g2_inv_1 _25057_ (.Y(_06473_),
    .A(_00238_));
 sg13g2_nand2_1 _25058_ (.Y(_06474_),
    .A(_06465_),
    .B(_06466_));
 sg13g2_buf_2 _25059_ (.A(_06474_),
    .X(_06475_));
 sg13g2_nor3_2 _25060_ (.A(_06462_),
    .B(_06473_),
    .C(_06475_),
    .Y(_06476_));
 sg13g2_nand2_2 _25061_ (.Y(_06477_),
    .A(_06461_),
    .B(_06476_));
 sg13g2_mux2_1 _25062_ (.A0(net843),
    .A1(\cpu.icache.r_data[0][10] ),
    .S(_06477_),
    .X(_02001_));
 sg13g2_buf_1 _25063_ (.A(net1099),
    .X(_06478_));
 sg13g2_mux2_1 _25064_ (.A0(net963),
    .A1(\cpu.icache.r_data[0][11] ),
    .S(_06477_),
    .X(_02002_));
 sg13g2_nor2b_1 _25065_ (.A(_06466_),
    .B_N(_06465_),
    .Y(_06479_));
 sg13g2_buf_1 _25066_ (.A(_06479_),
    .X(_06480_));
 sg13g2_and2_1 _25067_ (.A(_06464_),
    .B(_06480_),
    .X(_06481_));
 sg13g2_buf_2 _25068_ (.A(_06481_),
    .X(_06482_));
 sg13g2_nand2_2 _25069_ (.Y(_06483_),
    .A(_06461_),
    .B(_06482_));
 sg13g2_mux2_1 _25070_ (.A0(_06459_),
    .A1(\cpu.icache.r_data[0][12] ),
    .S(_06483_),
    .X(_02003_));
 sg13g2_buf_1 _25071_ (.A(net1002),
    .X(_06484_));
 sg13g2_mux2_1 _25072_ (.A0(_06484_),
    .A1(\cpu.icache.r_data[0][13] ),
    .S(_06483_),
    .X(_02004_));
 sg13g2_mux2_1 _25073_ (.A0(net843),
    .A1(\cpu.icache.r_data[0][14] ),
    .S(_06483_),
    .X(_02005_));
 sg13g2_mux2_1 _25074_ (.A0(_06478_),
    .A1(\cpu.icache.r_data[0][15] ),
    .S(_06483_),
    .X(_02006_));
 sg13g2_nor2_1 _25075_ (.A(_06462_),
    .B(_00238_),
    .Y(_06485_));
 sg13g2_buf_2 _25076_ (.A(_06485_),
    .X(_06486_));
 sg13g2_and2_1 _25077_ (.A(_06468_),
    .B(_06486_),
    .X(_06487_));
 sg13g2_buf_2 _25078_ (.A(_06487_),
    .X(_06488_));
 sg13g2_nand2_2 _25079_ (.Y(_06489_),
    .A(_06461_),
    .B(_06488_));
 sg13g2_mux2_1 _25080_ (.A0(net844),
    .A1(\cpu.icache.r_data[0][16] ),
    .S(_06489_),
    .X(_02007_));
 sg13g2_mux2_1 _25081_ (.A0(net842),
    .A1(\cpu.icache.r_data[0][17] ),
    .S(_06489_),
    .X(_02008_));
 sg13g2_mux2_1 _25082_ (.A0(net843),
    .A1(\cpu.icache.r_data[0][18] ),
    .S(_06489_),
    .X(_02009_));
 sg13g2_mux2_1 _25083_ (.A0(net963),
    .A1(\cpu.icache.r_data[0][19] ),
    .S(_06489_),
    .X(_02010_));
 sg13g2_mux2_1 _25084_ (.A0(net842),
    .A1(\cpu.icache.r_data[0][1] ),
    .S(_06471_),
    .X(_02011_));
 sg13g2_nor2_2 _25085_ (.A(_06465_),
    .B(_06466_),
    .Y(_06490_));
 sg13g2_and2_1 _25086_ (.A(_06486_),
    .B(_06490_),
    .X(_06491_));
 sg13g2_buf_2 _25087_ (.A(_06491_),
    .X(_06492_));
 sg13g2_nand2_2 _25088_ (.Y(_06493_),
    .A(_06461_),
    .B(_06492_));
 sg13g2_mux2_1 _25089_ (.A0(_06459_),
    .A1(\cpu.icache.r_data[0][20] ),
    .S(_06493_),
    .X(_02012_));
 sg13g2_mux2_1 _25090_ (.A0(net842),
    .A1(\cpu.icache.r_data[0][21] ),
    .S(_06493_),
    .X(_02013_));
 sg13g2_mux2_1 _25091_ (.A0(_06472_),
    .A1(\cpu.icache.r_data[0][22] ),
    .S(_06493_),
    .X(_02014_));
 sg13g2_mux2_1 _25092_ (.A0(net963),
    .A1(\cpu.icache.r_data[0][23] ),
    .S(_06493_),
    .X(_02015_));
 sg13g2_inv_1 _25093_ (.Y(_06494_),
    .A(\cpu.i_wstrobe_d ));
 sg13g2_nor3_2 _25094_ (.A(_00238_),
    .B(_06494_),
    .C(_06475_),
    .Y(_06495_));
 sg13g2_nand2_1 _25095_ (.Y(_06496_),
    .A(_06461_),
    .B(_06495_));
 sg13g2_buf_1 _25096_ (.A(_06496_),
    .X(_06497_));
 sg13g2_buf_1 _25097_ (.A(net439),
    .X(_06498_));
 sg13g2_mux2_1 _25098_ (.A0(net844),
    .A1(\cpu.icache.r_data[0][24] ),
    .S(net381),
    .X(_02016_));
 sg13g2_mux2_1 _25099_ (.A0(net842),
    .A1(\cpu.icache.r_data[0][25] ),
    .S(net381),
    .X(_02017_));
 sg13g2_mux2_1 _25100_ (.A0(net843),
    .A1(\cpu.icache.r_data[0][26] ),
    .S(net381),
    .X(_02018_));
 sg13g2_mux2_1 _25101_ (.A0(net963),
    .A1(\cpu.icache.r_data[0][27] ),
    .S(net381),
    .X(_02019_));
 sg13g2_and2_1 _25102_ (.A(_06480_),
    .B(_06486_),
    .X(_06499_));
 sg13g2_buf_2 _25103_ (.A(_06499_),
    .X(_06500_));
 sg13g2_nand2_2 _25104_ (.Y(_06501_),
    .A(_06461_),
    .B(_06500_));
 sg13g2_mux2_1 _25105_ (.A0(net844),
    .A1(\cpu.icache.r_data[0][28] ),
    .S(_06501_),
    .X(_02020_));
 sg13g2_mux2_1 _25106_ (.A0(net842),
    .A1(\cpu.icache.r_data[0][29] ),
    .S(_06501_),
    .X(_02021_));
 sg13g2_mux2_1 _25107_ (.A0(net843),
    .A1(\cpu.icache.r_data[0][2] ),
    .S(_06471_),
    .X(_02022_));
 sg13g2_mux2_1 _25108_ (.A0(net843),
    .A1(\cpu.icache.r_data[0][30] ),
    .S(_06501_),
    .X(_02023_));
 sg13g2_mux2_1 _25109_ (.A0(net963),
    .A1(\cpu.icache.r_data[0][31] ),
    .S(_06501_),
    .X(_02024_));
 sg13g2_mux2_1 _25110_ (.A0(net963),
    .A1(\cpu.icache.r_data[0][3] ),
    .S(_06471_),
    .X(_02025_));
 sg13g2_and2_1 _25111_ (.A(_06464_),
    .B(_06490_),
    .X(_06502_));
 sg13g2_buf_2 _25112_ (.A(_06502_),
    .X(_06503_));
 sg13g2_nand2_2 _25113_ (.Y(_06504_),
    .A(_06461_),
    .B(_06503_));
 sg13g2_mux2_1 _25114_ (.A0(net844),
    .A1(\cpu.icache.r_data[0][4] ),
    .S(_06504_),
    .X(_02026_));
 sg13g2_mux2_1 _25115_ (.A0(_06484_),
    .A1(\cpu.icache.r_data[0][5] ),
    .S(_06504_),
    .X(_02027_));
 sg13g2_mux2_1 _25116_ (.A0(_06472_),
    .A1(\cpu.icache.r_data[0][6] ),
    .S(_06504_),
    .X(_02028_));
 sg13g2_mux2_1 _25117_ (.A0(_06478_),
    .A1(\cpu.icache.r_data[0][7] ),
    .S(_06504_),
    .X(_02029_));
 sg13g2_mux2_1 _25118_ (.A0(net844),
    .A1(\cpu.icache.r_data[0][8] ),
    .S(_06477_),
    .X(_02030_));
 sg13g2_mux2_1 _25119_ (.A0(net842),
    .A1(\cpu.icache.r_data[0][9] ),
    .S(_06477_),
    .X(_02031_));
 sg13g2_buf_1 _25120_ (.A(net1004),
    .X(_06505_));
 sg13g2_nand2b_1 _25121_ (.Y(_06506_),
    .B(net806),
    .A_N(_08502_));
 sg13g2_buf_4 _25122_ (.X(_06507_),
    .A(_06506_));
 sg13g2_nand2_2 _25123_ (.Y(_06508_),
    .A(_06464_),
    .B(_06468_));
 sg13g2_nor2_2 _25124_ (.A(_06507_),
    .B(_06508_),
    .Y(_06509_));
 sg13g2_mux2_1 _25125_ (.A0(\cpu.icache.r_data[1][0] ),
    .A1(net841),
    .S(_06509_),
    .X(_02032_));
 sg13g2_buf_1 _25126_ (.A(net1003),
    .X(_06510_));
 sg13g2_or3_1 _25127_ (.A(_06462_),
    .B(_06473_),
    .C(_06475_),
    .X(_06511_));
 sg13g2_buf_2 _25128_ (.A(_06511_),
    .X(_06512_));
 sg13g2_nor2_2 _25129_ (.A(_06507_),
    .B(_06512_),
    .Y(_06513_));
 sg13g2_mux2_1 _25130_ (.A0(\cpu.icache.r_data[1][10] ),
    .A1(net840),
    .S(_06513_),
    .X(_02033_));
 sg13g2_buf_1 _25131_ (.A(net1099),
    .X(_06514_));
 sg13g2_mux2_1 _25132_ (.A0(\cpu.icache.r_data[1][11] ),
    .A1(net962),
    .S(_06513_),
    .X(_02034_));
 sg13g2_buf_1 _25133_ (.A(net1004),
    .X(_06515_));
 sg13g2_nand2_2 _25134_ (.Y(_06516_),
    .A(_06464_),
    .B(_06480_));
 sg13g2_nor2_2 _25135_ (.A(_06507_),
    .B(_06516_),
    .Y(_06517_));
 sg13g2_mux2_1 _25136_ (.A0(\cpu.icache.r_data[1][12] ),
    .A1(net839),
    .S(_06517_),
    .X(_02035_));
 sg13g2_buf_1 _25137_ (.A(net1002),
    .X(_06518_));
 sg13g2_mux2_1 _25138_ (.A0(\cpu.icache.r_data[1][13] ),
    .A1(net838),
    .S(_06517_),
    .X(_02036_));
 sg13g2_buf_1 _25139_ (.A(net1003),
    .X(_06519_));
 sg13g2_mux2_1 _25140_ (.A0(\cpu.icache.r_data[1][14] ),
    .A1(net837),
    .S(_06517_),
    .X(_02037_));
 sg13g2_buf_1 _25141_ (.A(net1099),
    .X(_06520_));
 sg13g2_mux2_1 _25142_ (.A0(\cpu.icache.r_data[1][15] ),
    .A1(net961),
    .S(_06517_),
    .X(_02038_));
 sg13g2_nand2_2 _25143_ (.Y(_06521_),
    .A(_06468_),
    .B(_06486_));
 sg13g2_nor2_2 _25144_ (.A(_06507_),
    .B(_06521_),
    .Y(_06522_));
 sg13g2_mux2_1 _25145_ (.A0(\cpu.icache.r_data[1][16] ),
    .A1(net839),
    .S(_06522_),
    .X(_02039_));
 sg13g2_buf_1 _25146_ (.A(net1002),
    .X(_06523_));
 sg13g2_mux2_1 _25147_ (.A0(\cpu.icache.r_data[1][17] ),
    .A1(net836),
    .S(_06522_),
    .X(_02040_));
 sg13g2_mux2_1 _25148_ (.A0(\cpu.icache.r_data[1][18] ),
    .A1(net837),
    .S(_06522_),
    .X(_02041_));
 sg13g2_mux2_1 _25149_ (.A0(\cpu.icache.r_data[1][19] ),
    .A1(net961),
    .S(_06522_),
    .X(_02042_));
 sg13g2_mux2_1 _25150_ (.A0(\cpu.icache.r_data[1][1] ),
    .A1(net836),
    .S(_06509_),
    .X(_02043_));
 sg13g2_nand2_2 _25151_ (.Y(_06524_),
    .A(_06486_),
    .B(_06490_));
 sg13g2_nor2_2 _25152_ (.A(_06507_),
    .B(_06524_),
    .Y(_06525_));
 sg13g2_mux2_1 _25153_ (.A0(\cpu.icache.r_data[1][20] ),
    .A1(_06515_),
    .S(_06525_),
    .X(_02044_));
 sg13g2_mux2_1 _25154_ (.A0(\cpu.icache.r_data[1][21] ),
    .A1(net836),
    .S(_06525_),
    .X(_02045_));
 sg13g2_mux2_1 _25155_ (.A0(\cpu.icache.r_data[1][22] ),
    .A1(net837),
    .S(_06525_),
    .X(_02046_));
 sg13g2_mux2_1 _25156_ (.A0(\cpu.icache.r_data[1][23] ),
    .A1(net961),
    .S(_06525_),
    .X(_02047_));
 sg13g2_nand4_1 _25157_ (.B(_06466_),
    .C(_06473_),
    .A(_06465_),
    .Y(_06526_),
    .D(\cpu.i_wstrobe_d ));
 sg13g2_buf_1 _25158_ (.A(_06526_),
    .X(_06527_));
 sg13g2_nor2_1 _25159_ (.A(_06507_),
    .B(_06527_),
    .Y(_06528_));
 sg13g2_buf_2 _25160_ (.A(_06528_),
    .X(_06529_));
 sg13g2_mux2_1 _25161_ (.A0(\cpu.icache.r_data[1][24] ),
    .A1(_06515_),
    .S(_06529_),
    .X(_02048_));
 sg13g2_mux2_1 _25162_ (.A0(\cpu.icache.r_data[1][25] ),
    .A1(_06523_),
    .S(_06529_),
    .X(_02049_));
 sg13g2_mux2_1 _25163_ (.A0(\cpu.icache.r_data[1][26] ),
    .A1(_06519_),
    .S(_06529_),
    .X(_02050_));
 sg13g2_mux2_1 _25164_ (.A0(\cpu.icache.r_data[1][27] ),
    .A1(net961),
    .S(_06529_),
    .X(_02051_));
 sg13g2_nand2_2 _25165_ (.Y(_06530_),
    .A(_06480_),
    .B(_06486_));
 sg13g2_nor2_2 _25166_ (.A(_06507_),
    .B(_06530_),
    .Y(_06531_));
 sg13g2_mux2_1 _25167_ (.A0(\cpu.icache.r_data[1][28] ),
    .A1(net839),
    .S(_06531_),
    .X(_02052_));
 sg13g2_mux2_1 _25168_ (.A0(\cpu.icache.r_data[1][29] ),
    .A1(net836),
    .S(_06531_),
    .X(_02053_));
 sg13g2_mux2_1 _25169_ (.A0(\cpu.icache.r_data[1][2] ),
    .A1(net837),
    .S(_06509_),
    .X(_02054_));
 sg13g2_mux2_1 _25170_ (.A0(\cpu.icache.r_data[1][30] ),
    .A1(net837),
    .S(_06531_),
    .X(_02055_));
 sg13g2_mux2_1 _25171_ (.A0(\cpu.icache.r_data[1][31] ),
    .A1(net961),
    .S(_06531_),
    .X(_02056_));
 sg13g2_mux2_1 _25172_ (.A0(\cpu.icache.r_data[1][3] ),
    .A1(net961),
    .S(_06509_),
    .X(_02057_));
 sg13g2_nand2_2 _25173_ (.Y(_06532_),
    .A(_06464_),
    .B(_06490_));
 sg13g2_nor2_2 _25174_ (.A(_06507_),
    .B(_06532_),
    .Y(_06533_));
 sg13g2_mux2_1 _25175_ (.A0(\cpu.icache.r_data[1][4] ),
    .A1(net839),
    .S(_06533_),
    .X(_02058_));
 sg13g2_mux2_1 _25176_ (.A0(\cpu.icache.r_data[1][5] ),
    .A1(net836),
    .S(_06533_),
    .X(_02059_));
 sg13g2_mux2_1 _25177_ (.A0(\cpu.icache.r_data[1][6] ),
    .A1(net837),
    .S(_06533_),
    .X(_02060_));
 sg13g2_mux2_1 _25178_ (.A0(\cpu.icache.r_data[1][7] ),
    .A1(_06520_),
    .S(_06533_),
    .X(_02061_));
 sg13g2_mux2_1 _25179_ (.A0(\cpu.icache.r_data[1][8] ),
    .A1(net839),
    .S(_06513_),
    .X(_02062_));
 sg13g2_mux2_1 _25180_ (.A0(\cpu.icache.r_data[1][9] ),
    .A1(_06523_),
    .S(_06513_),
    .X(_02063_));
 sg13g2_nand2_1 _25181_ (.Y(_06534_),
    .A(_08950_),
    .B(_08501_));
 sg13g2_buf_4 _25182_ (.X(_06535_),
    .A(_06534_));
 sg13g2_nor2_2 _25183_ (.A(_06535_),
    .B(_06508_),
    .Y(_06536_));
 sg13g2_mux2_1 _25184_ (.A0(\cpu.icache.r_data[2][0] ),
    .A1(net839),
    .S(_06536_),
    .X(_02064_));
 sg13g2_nor2_2 _25185_ (.A(_06535_),
    .B(_06512_),
    .Y(_06537_));
 sg13g2_mux2_1 _25186_ (.A0(\cpu.icache.r_data[2][10] ),
    .A1(_06519_),
    .S(_06537_),
    .X(_02065_));
 sg13g2_mux2_1 _25187_ (.A0(\cpu.icache.r_data[2][11] ),
    .A1(_06520_),
    .S(_06537_),
    .X(_02066_));
 sg13g2_nor2_2 _25188_ (.A(_06535_),
    .B(_06516_),
    .Y(_06538_));
 sg13g2_mux2_1 _25189_ (.A0(\cpu.icache.r_data[2][12] ),
    .A1(net839),
    .S(_06538_),
    .X(_02067_));
 sg13g2_mux2_1 _25190_ (.A0(\cpu.icache.r_data[2][13] ),
    .A1(net836),
    .S(_06538_),
    .X(_02068_));
 sg13g2_mux2_1 _25191_ (.A0(\cpu.icache.r_data[2][14] ),
    .A1(net837),
    .S(_06538_),
    .X(_02069_));
 sg13g2_mux2_1 _25192_ (.A0(\cpu.icache.r_data[2][15] ),
    .A1(net961),
    .S(_06538_),
    .X(_02070_));
 sg13g2_nor2_2 _25193_ (.A(_06535_),
    .B(_06521_),
    .Y(_06539_));
 sg13g2_mux2_1 _25194_ (.A0(\cpu.icache.r_data[2][16] ),
    .A1(net839),
    .S(_06539_),
    .X(_02071_));
 sg13g2_mux2_1 _25195_ (.A0(\cpu.icache.r_data[2][17] ),
    .A1(net836),
    .S(_06539_),
    .X(_02072_));
 sg13g2_mux2_1 _25196_ (.A0(\cpu.icache.r_data[2][18] ),
    .A1(net837),
    .S(_06539_),
    .X(_02073_));
 sg13g2_mux2_1 _25197_ (.A0(\cpu.icache.r_data[2][19] ),
    .A1(net961),
    .S(_06539_),
    .X(_02074_));
 sg13g2_mux2_1 _25198_ (.A0(\cpu.icache.r_data[2][1] ),
    .A1(net836),
    .S(_06536_),
    .X(_02075_));
 sg13g2_buf_1 _25199_ (.A(_02836_),
    .X(_06540_));
 sg13g2_nor2_2 _25200_ (.A(_06535_),
    .B(_06524_),
    .Y(_06541_));
 sg13g2_mux2_1 _25201_ (.A0(\cpu.icache.r_data[2][20] ),
    .A1(net835),
    .S(_06541_),
    .X(_02076_));
 sg13g2_buf_1 _25202_ (.A(_02861_),
    .X(_06542_));
 sg13g2_mux2_1 _25203_ (.A0(\cpu.icache.r_data[2][21] ),
    .A1(net834),
    .S(_06541_),
    .X(_02077_));
 sg13g2_buf_1 _25204_ (.A(_02845_),
    .X(_06543_));
 sg13g2_mux2_1 _25205_ (.A0(\cpu.icache.r_data[2][22] ),
    .A1(net833),
    .S(_06541_),
    .X(_02078_));
 sg13g2_buf_1 _25206_ (.A(_02849_),
    .X(_06544_));
 sg13g2_mux2_1 _25207_ (.A0(\cpu.icache.r_data[2][23] ),
    .A1(net960),
    .S(_06541_),
    .X(_02079_));
 sg13g2_nor2_1 _25208_ (.A(_06535_),
    .B(_06527_),
    .Y(_06545_));
 sg13g2_buf_2 _25209_ (.A(_06545_),
    .X(_06546_));
 sg13g2_mux2_1 _25210_ (.A0(\cpu.icache.r_data[2][24] ),
    .A1(net835),
    .S(_06546_),
    .X(_02080_));
 sg13g2_mux2_1 _25211_ (.A0(\cpu.icache.r_data[2][25] ),
    .A1(net834),
    .S(_06546_),
    .X(_02081_));
 sg13g2_mux2_1 _25212_ (.A0(\cpu.icache.r_data[2][26] ),
    .A1(net833),
    .S(_06546_),
    .X(_02082_));
 sg13g2_mux2_1 _25213_ (.A0(\cpu.icache.r_data[2][27] ),
    .A1(net960),
    .S(_06546_),
    .X(_02083_));
 sg13g2_nor2_2 _25214_ (.A(_06535_),
    .B(_06530_),
    .Y(_06547_));
 sg13g2_mux2_1 _25215_ (.A0(\cpu.icache.r_data[2][28] ),
    .A1(net835),
    .S(_06547_),
    .X(_02084_));
 sg13g2_mux2_1 _25216_ (.A0(\cpu.icache.r_data[2][29] ),
    .A1(net834),
    .S(_06547_),
    .X(_02085_));
 sg13g2_mux2_1 _25217_ (.A0(\cpu.icache.r_data[2][2] ),
    .A1(net833),
    .S(_06536_),
    .X(_02086_));
 sg13g2_mux2_1 _25218_ (.A0(\cpu.icache.r_data[2][30] ),
    .A1(_06543_),
    .S(_06547_),
    .X(_02087_));
 sg13g2_mux2_1 _25219_ (.A0(\cpu.icache.r_data[2][31] ),
    .A1(net960),
    .S(_06547_),
    .X(_02088_));
 sg13g2_mux2_1 _25220_ (.A0(\cpu.icache.r_data[2][3] ),
    .A1(net960),
    .S(_06536_),
    .X(_02089_));
 sg13g2_nor2_2 _25221_ (.A(_06535_),
    .B(_06532_),
    .Y(_06548_));
 sg13g2_mux2_1 _25222_ (.A0(\cpu.icache.r_data[2][4] ),
    .A1(net835),
    .S(_06548_),
    .X(_02090_));
 sg13g2_mux2_1 _25223_ (.A0(\cpu.icache.r_data[2][5] ),
    .A1(net834),
    .S(_06548_),
    .X(_02091_));
 sg13g2_mux2_1 _25224_ (.A0(\cpu.icache.r_data[2][6] ),
    .A1(net833),
    .S(_06548_),
    .X(_02092_));
 sg13g2_mux2_1 _25225_ (.A0(\cpu.icache.r_data[2][7] ),
    .A1(net960),
    .S(_06548_),
    .X(_02093_));
 sg13g2_mux2_1 _25226_ (.A0(\cpu.icache.r_data[2][8] ),
    .A1(_06540_),
    .S(_06537_),
    .X(_02094_));
 sg13g2_mux2_1 _25227_ (.A0(\cpu.icache.r_data[2][9] ),
    .A1(net834),
    .S(_06537_),
    .X(_02095_));
 sg13g2_nand2_2 _25228_ (.Y(_06549_),
    .A(net518),
    .B(_06470_));
 sg13g2_mux2_1 _25229_ (.A0(net844),
    .A1(\cpu.icache.r_data[3][0] ),
    .S(_06549_),
    .X(_02096_));
 sg13g2_and2_1 _25230_ (.A(net518),
    .B(_06476_),
    .X(_06550_));
 sg13g2_buf_1 _25231_ (.A(_06550_),
    .X(_06551_));
 sg13g2_mux2_1 _25232_ (.A0(\cpu.icache.r_data[3][10] ),
    .A1(net833),
    .S(_06551_),
    .X(_02097_));
 sg13g2_mux2_1 _25233_ (.A0(\cpu.icache.r_data[3][11] ),
    .A1(net960),
    .S(_06551_),
    .X(_02098_));
 sg13g2_nand2_2 _25234_ (.Y(_06552_),
    .A(net518),
    .B(_06482_));
 sg13g2_mux2_1 _25235_ (.A0(net844),
    .A1(\cpu.icache.r_data[3][12] ),
    .S(_06552_),
    .X(_02099_));
 sg13g2_mux2_1 _25236_ (.A0(net842),
    .A1(\cpu.icache.r_data[3][13] ),
    .S(_06552_),
    .X(_02100_));
 sg13g2_mux2_1 _25237_ (.A0(net843),
    .A1(\cpu.icache.r_data[3][14] ),
    .S(_06552_),
    .X(_02101_));
 sg13g2_mux2_1 _25238_ (.A0(net963),
    .A1(\cpu.icache.r_data[3][15] ),
    .S(_06552_),
    .X(_02102_));
 sg13g2_buf_1 _25239_ (.A(_02836_),
    .X(_06553_));
 sg13g2_nand2_2 _25240_ (.Y(_06554_),
    .A(net518),
    .B(_06488_));
 sg13g2_mux2_1 _25241_ (.A0(net832),
    .A1(\cpu.icache.r_data[3][16] ),
    .S(_06554_),
    .X(_02103_));
 sg13g2_mux2_1 _25242_ (.A0(net842),
    .A1(\cpu.icache.r_data[3][17] ),
    .S(_06554_),
    .X(_02104_));
 sg13g2_mux2_1 _25243_ (.A0(net843),
    .A1(\cpu.icache.r_data[3][18] ),
    .S(_06554_),
    .X(_02105_));
 sg13g2_mux2_1 _25244_ (.A0(net963),
    .A1(\cpu.icache.r_data[3][19] ),
    .S(_06554_),
    .X(_02106_));
 sg13g2_buf_1 _25245_ (.A(_02861_),
    .X(_06555_));
 sg13g2_mux2_1 _25246_ (.A0(net831),
    .A1(\cpu.icache.r_data[3][1] ),
    .S(_06549_),
    .X(_02107_));
 sg13g2_nand2_2 _25247_ (.Y(_06556_),
    .A(_09031_),
    .B(_06492_));
 sg13g2_mux2_1 _25248_ (.A0(net832),
    .A1(\cpu.icache.r_data[3][20] ),
    .S(_06556_),
    .X(_02108_));
 sg13g2_mux2_1 _25249_ (.A0(_06555_),
    .A1(\cpu.icache.r_data[3][21] ),
    .S(_06556_),
    .X(_02109_));
 sg13g2_buf_1 _25250_ (.A(_02845_),
    .X(_06557_));
 sg13g2_mux2_1 _25251_ (.A0(net830),
    .A1(\cpu.icache.r_data[3][22] ),
    .S(_06556_),
    .X(_02110_));
 sg13g2_buf_1 _25252_ (.A(_02849_),
    .X(_06558_));
 sg13g2_mux2_1 _25253_ (.A0(net959),
    .A1(\cpu.icache.r_data[3][23] ),
    .S(_06556_),
    .X(_02111_));
 sg13g2_nand2_1 _25254_ (.Y(_06559_),
    .A(net518),
    .B(_06495_));
 sg13g2_buf_1 _25255_ (.A(_06559_),
    .X(_06560_));
 sg13g2_buf_1 _25256_ (.A(_06560_),
    .X(_06561_));
 sg13g2_mux2_1 _25257_ (.A0(_06553_),
    .A1(\cpu.icache.r_data[3][24] ),
    .S(net295),
    .X(_02112_));
 sg13g2_mux2_1 _25258_ (.A0(_06555_),
    .A1(\cpu.icache.r_data[3][25] ),
    .S(net295),
    .X(_02113_));
 sg13g2_mux2_1 _25259_ (.A0(_06557_),
    .A1(\cpu.icache.r_data[3][26] ),
    .S(net295),
    .X(_02114_));
 sg13g2_mux2_1 _25260_ (.A0(net959),
    .A1(\cpu.icache.r_data[3][27] ),
    .S(net295),
    .X(_02115_));
 sg13g2_nand2_2 _25261_ (.Y(_06562_),
    .A(net518),
    .B(_06500_));
 sg13g2_mux2_1 _25262_ (.A0(net832),
    .A1(\cpu.icache.r_data[3][28] ),
    .S(_06562_),
    .X(_02116_));
 sg13g2_mux2_1 _25263_ (.A0(net831),
    .A1(\cpu.icache.r_data[3][29] ),
    .S(_06562_),
    .X(_02117_));
 sg13g2_mux2_1 _25264_ (.A0(net830),
    .A1(\cpu.icache.r_data[3][2] ),
    .S(_06549_),
    .X(_02118_));
 sg13g2_mux2_1 _25265_ (.A0(net830),
    .A1(\cpu.icache.r_data[3][30] ),
    .S(_06562_),
    .X(_02119_));
 sg13g2_mux2_1 _25266_ (.A0(net959),
    .A1(\cpu.icache.r_data[3][31] ),
    .S(_06562_),
    .X(_02120_));
 sg13g2_mux2_1 _25267_ (.A0(net959),
    .A1(\cpu.icache.r_data[3][3] ),
    .S(_06549_),
    .X(_02121_));
 sg13g2_nand2_2 _25268_ (.Y(_06563_),
    .A(_09031_),
    .B(_06503_));
 sg13g2_mux2_1 _25269_ (.A0(_06553_),
    .A1(\cpu.icache.r_data[3][4] ),
    .S(_06563_),
    .X(_02122_));
 sg13g2_mux2_1 _25270_ (.A0(net831),
    .A1(\cpu.icache.r_data[3][5] ),
    .S(_06563_),
    .X(_02123_));
 sg13g2_mux2_1 _25271_ (.A0(net830),
    .A1(\cpu.icache.r_data[3][6] ),
    .S(_06563_),
    .X(_02124_));
 sg13g2_mux2_1 _25272_ (.A0(_06558_),
    .A1(\cpu.icache.r_data[3][7] ),
    .S(_06563_),
    .X(_02125_));
 sg13g2_mux2_1 _25273_ (.A0(\cpu.icache.r_data[3][8] ),
    .A1(_06540_),
    .S(_06551_),
    .X(_02126_));
 sg13g2_mux2_1 _25274_ (.A0(\cpu.icache.r_data[3][9] ),
    .A1(net834),
    .S(_06551_),
    .X(_02127_));
 sg13g2_nand2_2 _25275_ (.Y(_06564_),
    .A(net636),
    .B(_06470_));
 sg13g2_mux2_1 _25276_ (.A0(net832),
    .A1(\cpu.icache.r_data[4][0] ),
    .S(_06564_),
    .X(_02128_));
 sg13g2_and2_1 _25277_ (.A(net636),
    .B(_06476_),
    .X(_06565_));
 sg13g2_buf_1 _25278_ (.A(_06565_),
    .X(_06566_));
 sg13g2_mux2_1 _25279_ (.A0(\cpu.icache.r_data[4][10] ),
    .A1(net833),
    .S(_06566_),
    .X(_02129_));
 sg13g2_mux2_1 _25280_ (.A0(\cpu.icache.r_data[4][11] ),
    .A1(net960),
    .S(_06566_),
    .X(_02130_));
 sg13g2_nand2_2 _25281_ (.Y(_06567_),
    .A(net636),
    .B(_06482_));
 sg13g2_mux2_1 _25282_ (.A0(net832),
    .A1(\cpu.icache.r_data[4][12] ),
    .S(_06567_),
    .X(_02131_));
 sg13g2_mux2_1 _25283_ (.A0(net831),
    .A1(\cpu.icache.r_data[4][13] ),
    .S(_06567_),
    .X(_02132_));
 sg13g2_mux2_1 _25284_ (.A0(_06557_),
    .A1(\cpu.icache.r_data[4][14] ),
    .S(_06567_),
    .X(_02133_));
 sg13g2_mux2_1 _25285_ (.A0(_06558_),
    .A1(\cpu.icache.r_data[4][15] ),
    .S(_06567_),
    .X(_02134_));
 sg13g2_nand2_2 _25286_ (.Y(_06568_),
    .A(net636),
    .B(_06488_));
 sg13g2_mux2_1 _25287_ (.A0(net832),
    .A1(\cpu.icache.r_data[4][16] ),
    .S(_06568_),
    .X(_02135_));
 sg13g2_mux2_1 _25288_ (.A0(net831),
    .A1(\cpu.icache.r_data[4][17] ),
    .S(_06568_),
    .X(_02136_));
 sg13g2_mux2_1 _25289_ (.A0(net830),
    .A1(\cpu.icache.r_data[4][18] ),
    .S(_06568_),
    .X(_02137_));
 sg13g2_mux2_1 _25290_ (.A0(net959),
    .A1(\cpu.icache.r_data[4][19] ),
    .S(_06568_),
    .X(_02138_));
 sg13g2_mux2_1 _25291_ (.A0(net831),
    .A1(\cpu.icache.r_data[4][1] ),
    .S(_06564_),
    .X(_02139_));
 sg13g2_nand2_2 _25292_ (.Y(_06569_),
    .A(net636),
    .B(_06492_));
 sg13g2_mux2_1 _25293_ (.A0(net832),
    .A1(\cpu.icache.r_data[4][20] ),
    .S(_06569_),
    .X(_02140_));
 sg13g2_mux2_1 _25294_ (.A0(net831),
    .A1(\cpu.icache.r_data[4][21] ),
    .S(_06569_),
    .X(_02141_));
 sg13g2_mux2_1 _25295_ (.A0(net830),
    .A1(\cpu.icache.r_data[4][22] ),
    .S(_06569_),
    .X(_02142_));
 sg13g2_mux2_1 _25296_ (.A0(net959),
    .A1(\cpu.icache.r_data[4][23] ),
    .S(_06569_),
    .X(_02143_));
 sg13g2_and2_1 _25297_ (.A(_09035_),
    .B(_06495_),
    .X(_06570_));
 sg13g2_buf_2 _25298_ (.A(_06570_),
    .X(_06571_));
 sg13g2_mux2_1 _25299_ (.A0(\cpu.icache.r_data[4][24] ),
    .A1(net835),
    .S(_06571_),
    .X(_02144_));
 sg13g2_mux2_1 _25300_ (.A0(\cpu.icache.r_data[4][25] ),
    .A1(net834),
    .S(_06571_),
    .X(_02145_));
 sg13g2_mux2_1 _25301_ (.A0(\cpu.icache.r_data[4][26] ),
    .A1(_06543_),
    .S(_06571_),
    .X(_02146_));
 sg13g2_mux2_1 _25302_ (.A0(\cpu.icache.r_data[4][27] ),
    .A1(_06544_),
    .S(_06571_),
    .X(_02147_));
 sg13g2_nand2_2 _25303_ (.Y(_06572_),
    .A(net636),
    .B(_06500_));
 sg13g2_mux2_1 _25304_ (.A0(net832),
    .A1(\cpu.icache.r_data[4][28] ),
    .S(_06572_),
    .X(_02148_));
 sg13g2_mux2_1 _25305_ (.A0(net831),
    .A1(\cpu.icache.r_data[4][29] ),
    .S(_06572_),
    .X(_02149_));
 sg13g2_mux2_1 _25306_ (.A0(net830),
    .A1(\cpu.icache.r_data[4][2] ),
    .S(_06564_),
    .X(_02150_));
 sg13g2_mux2_1 _25307_ (.A0(net830),
    .A1(\cpu.icache.r_data[4][30] ),
    .S(_06572_),
    .X(_02151_));
 sg13g2_mux2_1 _25308_ (.A0(net959),
    .A1(\cpu.icache.r_data[4][31] ),
    .S(_06572_),
    .X(_02152_));
 sg13g2_mux2_1 _25309_ (.A0(net959),
    .A1(\cpu.icache.r_data[4][3] ),
    .S(_06564_),
    .X(_02153_));
 sg13g2_nand2_2 _25310_ (.Y(_06573_),
    .A(net636),
    .B(_06503_));
 sg13g2_mux2_1 _25311_ (.A0(net841),
    .A1(\cpu.icache.r_data[4][4] ),
    .S(_06573_),
    .X(_02154_));
 sg13g2_mux2_1 _25312_ (.A0(net838),
    .A1(\cpu.icache.r_data[4][5] ),
    .S(_06573_),
    .X(_02155_));
 sg13g2_mux2_1 _25313_ (.A0(net840),
    .A1(\cpu.icache.r_data[4][6] ),
    .S(_06573_),
    .X(_02156_));
 sg13g2_mux2_1 _25314_ (.A0(net962),
    .A1(\cpu.icache.r_data[4][7] ),
    .S(_06573_),
    .X(_02157_));
 sg13g2_mux2_1 _25315_ (.A0(\cpu.icache.r_data[4][8] ),
    .A1(net835),
    .S(_06566_),
    .X(_02158_));
 sg13g2_mux2_1 _25316_ (.A0(\cpu.icache.r_data[4][9] ),
    .A1(_06542_),
    .S(_06566_),
    .X(_02159_));
 sg13g2_nand2_1 _25317_ (.Y(_06574_),
    .A(net715),
    .B(net806));
 sg13g2_buf_4 _25318_ (.X(_06575_),
    .A(_06574_));
 sg13g2_nor2_2 _25319_ (.A(_06575_),
    .B(_06508_),
    .Y(_06576_));
 sg13g2_mux2_1 _25320_ (.A0(\cpu.icache.r_data[5][0] ),
    .A1(net835),
    .S(_06576_),
    .X(_02160_));
 sg13g2_nor2_2 _25321_ (.A(_06575_),
    .B(_06512_),
    .Y(_06577_));
 sg13g2_mux2_1 _25322_ (.A0(\cpu.icache.r_data[5][10] ),
    .A1(net833),
    .S(_06577_),
    .X(_02161_));
 sg13g2_mux2_1 _25323_ (.A0(\cpu.icache.r_data[5][11] ),
    .A1(_06544_),
    .S(_06577_),
    .X(_02162_));
 sg13g2_nor2_2 _25324_ (.A(_06575_),
    .B(_06516_),
    .Y(_06578_));
 sg13g2_mux2_1 _25325_ (.A0(\cpu.icache.r_data[5][12] ),
    .A1(net835),
    .S(_06578_),
    .X(_02163_));
 sg13g2_mux2_1 _25326_ (.A0(\cpu.icache.r_data[5][13] ),
    .A1(_06542_),
    .S(_06578_),
    .X(_02164_));
 sg13g2_mux2_1 _25327_ (.A0(\cpu.icache.r_data[5][14] ),
    .A1(net833),
    .S(_06578_),
    .X(_02165_));
 sg13g2_mux2_1 _25328_ (.A0(\cpu.icache.r_data[5][15] ),
    .A1(net960),
    .S(_06578_),
    .X(_02166_));
 sg13g2_buf_2 _25329_ (.A(net1110),
    .X(_06579_));
 sg13g2_nor2_2 _25330_ (.A(_06575_),
    .B(_06521_),
    .Y(_06580_));
 sg13g2_mux2_1 _25331_ (.A0(\cpu.icache.r_data[5][16] ),
    .A1(net958),
    .S(_06580_),
    .X(_02167_));
 sg13g2_mux2_1 _25332_ (.A0(\cpu.icache.r_data[5][17] ),
    .A1(net834),
    .S(_06580_),
    .X(_02168_));
 sg13g2_buf_2 _25333_ (.A(net1109),
    .X(_06581_));
 sg13g2_mux2_1 _25334_ (.A0(\cpu.icache.r_data[5][18] ),
    .A1(net957),
    .S(_06580_),
    .X(_02169_));
 sg13g2_buf_2 _25335_ (.A(net1108),
    .X(_06582_));
 sg13g2_mux2_1 _25336_ (.A0(\cpu.icache.r_data[5][19] ),
    .A1(net956),
    .S(_06580_),
    .X(_02170_));
 sg13g2_buf_2 _25337_ (.A(net1107),
    .X(_06583_));
 sg13g2_mux2_1 _25338_ (.A0(\cpu.icache.r_data[5][1] ),
    .A1(net955),
    .S(_06576_),
    .X(_02171_));
 sg13g2_nor2_2 _25339_ (.A(_06575_),
    .B(_06524_),
    .Y(_06584_));
 sg13g2_mux2_1 _25340_ (.A0(\cpu.icache.r_data[5][20] ),
    .A1(net958),
    .S(_06584_),
    .X(_02172_));
 sg13g2_mux2_1 _25341_ (.A0(\cpu.icache.r_data[5][21] ),
    .A1(net955),
    .S(_06584_),
    .X(_02173_));
 sg13g2_mux2_1 _25342_ (.A0(\cpu.icache.r_data[5][22] ),
    .A1(net957),
    .S(_06584_),
    .X(_02174_));
 sg13g2_mux2_1 _25343_ (.A0(\cpu.icache.r_data[5][23] ),
    .A1(net956),
    .S(_06584_),
    .X(_02175_));
 sg13g2_nor2_1 _25344_ (.A(_06575_),
    .B(_06527_),
    .Y(_06585_));
 sg13g2_buf_2 _25345_ (.A(_06585_),
    .X(_06586_));
 sg13g2_mux2_1 _25346_ (.A0(\cpu.icache.r_data[5][24] ),
    .A1(net958),
    .S(_06586_),
    .X(_02176_));
 sg13g2_mux2_1 _25347_ (.A0(\cpu.icache.r_data[5][25] ),
    .A1(net955),
    .S(_06586_),
    .X(_02177_));
 sg13g2_mux2_1 _25348_ (.A0(\cpu.icache.r_data[5][26] ),
    .A1(net957),
    .S(_06586_),
    .X(_02178_));
 sg13g2_mux2_1 _25349_ (.A0(\cpu.icache.r_data[5][27] ),
    .A1(net956),
    .S(_06586_),
    .X(_02179_));
 sg13g2_nor2_2 _25350_ (.A(_06575_),
    .B(_06530_),
    .Y(_06587_));
 sg13g2_mux2_1 _25351_ (.A0(\cpu.icache.r_data[5][28] ),
    .A1(net958),
    .S(_06587_),
    .X(_02180_));
 sg13g2_mux2_1 _25352_ (.A0(\cpu.icache.r_data[5][29] ),
    .A1(net955),
    .S(_06587_),
    .X(_02181_));
 sg13g2_mux2_1 _25353_ (.A0(\cpu.icache.r_data[5][2] ),
    .A1(_06581_),
    .S(_06576_),
    .X(_02182_));
 sg13g2_mux2_1 _25354_ (.A0(\cpu.icache.r_data[5][30] ),
    .A1(net957),
    .S(_06587_),
    .X(_02183_));
 sg13g2_mux2_1 _25355_ (.A0(\cpu.icache.r_data[5][31] ),
    .A1(net956),
    .S(_06587_),
    .X(_02184_));
 sg13g2_mux2_1 _25356_ (.A0(\cpu.icache.r_data[5][3] ),
    .A1(net956),
    .S(_06576_),
    .X(_02185_));
 sg13g2_nor2_2 _25357_ (.A(_06575_),
    .B(_06532_),
    .Y(_06588_));
 sg13g2_mux2_1 _25358_ (.A0(\cpu.icache.r_data[5][4] ),
    .A1(net958),
    .S(_06588_),
    .X(_02186_));
 sg13g2_mux2_1 _25359_ (.A0(\cpu.icache.r_data[5][5] ),
    .A1(net955),
    .S(_06588_),
    .X(_02187_));
 sg13g2_mux2_1 _25360_ (.A0(\cpu.icache.r_data[5][6] ),
    .A1(net957),
    .S(_06588_),
    .X(_02188_));
 sg13g2_mux2_1 _25361_ (.A0(\cpu.icache.r_data[5][7] ),
    .A1(_06582_),
    .S(_06588_),
    .X(_02189_));
 sg13g2_mux2_1 _25362_ (.A0(\cpu.icache.r_data[5][8] ),
    .A1(_06579_),
    .S(_06577_),
    .X(_02190_));
 sg13g2_mux2_1 _25363_ (.A0(\cpu.icache.r_data[5][9] ),
    .A1(_06583_),
    .S(_06577_),
    .X(_02191_));
 sg13g2_nand2_2 _25364_ (.Y(_06589_),
    .A(net635),
    .B(_06470_));
 sg13g2_mux2_1 _25365_ (.A0(net841),
    .A1(\cpu.icache.r_data[6][0] ),
    .S(_06589_),
    .X(_02192_));
 sg13g2_nand2_2 _25366_ (.Y(_06590_),
    .A(net635),
    .B(_06476_));
 sg13g2_mux2_1 _25367_ (.A0(_06510_),
    .A1(\cpu.icache.r_data[6][10] ),
    .S(_06590_),
    .X(_02193_));
 sg13g2_mux2_1 _25368_ (.A0(_06514_),
    .A1(\cpu.icache.r_data[6][11] ),
    .S(_06590_),
    .X(_02194_));
 sg13g2_nand2_2 _25369_ (.Y(_06591_),
    .A(net635),
    .B(_06482_));
 sg13g2_mux2_1 _25370_ (.A0(net841),
    .A1(\cpu.icache.r_data[6][12] ),
    .S(_06591_),
    .X(_02195_));
 sg13g2_mux2_1 _25371_ (.A0(net838),
    .A1(\cpu.icache.r_data[6][13] ),
    .S(_06591_),
    .X(_02196_));
 sg13g2_mux2_1 _25372_ (.A0(net840),
    .A1(\cpu.icache.r_data[6][14] ),
    .S(_06591_),
    .X(_02197_));
 sg13g2_mux2_1 _25373_ (.A0(net962),
    .A1(\cpu.icache.r_data[6][15] ),
    .S(_06591_),
    .X(_02198_));
 sg13g2_nand2_2 _25374_ (.Y(_06592_),
    .A(net635),
    .B(_06488_));
 sg13g2_mux2_1 _25375_ (.A0(net841),
    .A1(\cpu.icache.r_data[6][16] ),
    .S(_06592_),
    .X(_02199_));
 sg13g2_mux2_1 _25376_ (.A0(net838),
    .A1(\cpu.icache.r_data[6][17] ),
    .S(_06592_),
    .X(_02200_));
 sg13g2_mux2_1 _25377_ (.A0(net840),
    .A1(\cpu.icache.r_data[6][18] ),
    .S(_06592_),
    .X(_02201_));
 sg13g2_mux2_1 _25378_ (.A0(net962),
    .A1(\cpu.icache.r_data[6][19] ),
    .S(_06592_),
    .X(_02202_));
 sg13g2_mux2_1 _25379_ (.A0(net838),
    .A1(\cpu.icache.r_data[6][1] ),
    .S(_06589_),
    .X(_02203_));
 sg13g2_nand2_2 _25380_ (.Y(_06593_),
    .A(net635),
    .B(_06492_));
 sg13g2_mux2_1 _25381_ (.A0(net841),
    .A1(\cpu.icache.r_data[6][20] ),
    .S(_06593_),
    .X(_02204_));
 sg13g2_mux2_1 _25382_ (.A0(net838),
    .A1(\cpu.icache.r_data[6][21] ),
    .S(_06593_),
    .X(_02205_));
 sg13g2_mux2_1 _25383_ (.A0(net840),
    .A1(\cpu.icache.r_data[6][22] ),
    .S(_06593_),
    .X(_02206_));
 sg13g2_mux2_1 _25384_ (.A0(net962),
    .A1(\cpu.icache.r_data[6][23] ),
    .S(_06593_),
    .X(_02207_));
 sg13g2_nand2_1 _25385_ (.Y(_06594_),
    .A(_09037_),
    .B(_06495_));
 sg13g2_buf_2 _25386_ (.A(_06594_),
    .X(_06595_));
 sg13g2_mux2_1 _25387_ (.A0(_06505_),
    .A1(\cpu.icache.r_data[6][24] ),
    .S(_06595_),
    .X(_02208_));
 sg13g2_mux2_1 _25388_ (.A0(_06518_),
    .A1(\cpu.icache.r_data[6][25] ),
    .S(_06595_),
    .X(_02209_));
 sg13g2_mux2_1 _25389_ (.A0(_06510_),
    .A1(\cpu.icache.r_data[6][26] ),
    .S(_06595_),
    .X(_02210_));
 sg13g2_mux2_1 _25390_ (.A0(_06514_),
    .A1(\cpu.icache.r_data[6][27] ),
    .S(_06595_),
    .X(_02211_));
 sg13g2_nand2_2 _25391_ (.Y(_06596_),
    .A(net635),
    .B(_06500_));
 sg13g2_mux2_1 _25392_ (.A0(net841),
    .A1(\cpu.icache.r_data[6][28] ),
    .S(_06596_),
    .X(_02212_));
 sg13g2_mux2_1 _25393_ (.A0(net838),
    .A1(\cpu.icache.r_data[6][29] ),
    .S(_06596_),
    .X(_02213_));
 sg13g2_mux2_1 _25394_ (.A0(net840),
    .A1(\cpu.icache.r_data[6][2] ),
    .S(_06589_),
    .X(_02214_));
 sg13g2_mux2_1 _25395_ (.A0(net840),
    .A1(\cpu.icache.r_data[6][30] ),
    .S(_06596_),
    .X(_02215_));
 sg13g2_mux2_1 _25396_ (.A0(net962),
    .A1(\cpu.icache.r_data[6][31] ),
    .S(_06596_),
    .X(_02216_));
 sg13g2_mux2_1 _25397_ (.A0(net962),
    .A1(\cpu.icache.r_data[6][3] ),
    .S(_06589_),
    .X(_02217_));
 sg13g2_nand2_2 _25398_ (.Y(_06597_),
    .A(net635),
    .B(_06503_));
 sg13g2_mux2_1 _25399_ (.A0(net841),
    .A1(\cpu.icache.r_data[6][4] ),
    .S(_06597_),
    .X(_02218_));
 sg13g2_mux2_1 _25400_ (.A0(net838),
    .A1(\cpu.icache.r_data[6][5] ),
    .S(_06597_),
    .X(_02219_));
 sg13g2_mux2_1 _25401_ (.A0(net840),
    .A1(\cpu.icache.r_data[6][6] ),
    .S(_06597_),
    .X(_02220_));
 sg13g2_mux2_1 _25402_ (.A0(net962),
    .A1(\cpu.icache.r_data[6][7] ),
    .S(_06597_),
    .X(_02221_));
 sg13g2_mux2_1 _25403_ (.A0(_06505_),
    .A1(\cpu.icache.r_data[6][8] ),
    .S(_06590_),
    .X(_02222_));
 sg13g2_mux2_1 _25404_ (.A0(_06518_),
    .A1(\cpu.icache.r_data[6][9] ),
    .S(_06590_),
    .X(_02223_));
 sg13g2_nand2_1 _25405_ (.Y(_06598_),
    .A(net715),
    .B(net820));
 sg13g2_buf_4 _25406_ (.X(_06599_),
    .A(_06598_));
 sg13g2_nor2_2 _25407_ (.A(_06599_),
    .B(_06508_),
    .Y(_06600_));
 sg13g2_mux2_1 _25408_ (.A0(\cpu.icache.r_data[7][0] ),
    .A1(net958),
    .S(_06600_),
    .X(_02224_));
 sg13g2_nor2_2 _25409_ (.A(_06599_),
    .B(_06512_),
    .Y(_06601_));
 sg13g2_mux2_1 _25410_ (.A0(\cpu.icache.r_data[7][10] ),
    .A1(net957),
    .S(_06601_),
    .X(_02225_));
 sg13g2_mux2_1 _25411_ (.A0(\cpu.icache.r_data[7][11] ),
    .A1(net956),
    .S(_06601_),
    .X(_02226_));
 sg13g2_nor2_2 _25412_ (.A(_06599_),
    .B(_06516_),
    .Y(_06602_));
 sg13g2_mux2_1 _25413_ (.A0(\cpu.icache.r_data[7][12] ),
    .A1(_06579_),
    .S(_06602_),
    .X(_02227_));
 sg13g2_mux2_1 _25414_ (.A0(\cpu.icache.r_data[7][13] ),
    .A1(net955),
    .S(_06602_),
    .X(_02228_));
 sg13g2_mux2_1 _25415_ (.A0(\cpu.icache.r_data[7][14] ),
    .A1(net957),
    .S(_06602_),
    .X(_02229_));
 sg13g2_mux2_1 _25416_ (.A0(\cpu.icache.r_data[7][15] ),
    .A1(_06582_),
    .S(_06602_),
    .X(_02230_));
 sg13g2_nor2_2 _25417_ (.A(_06599_),
    .B(_06521_),
    .Y(_06603_));
 sg13g2_mux2_1 _25418_ (.A0(\cpu.icache.r_data[7][16] ),
    .A1(net958),
    .S(_06603_),
    .X(_02231_));
 sg13g2_mux2_1 _25419_ (.A0(\cpu.icache.r_data[7][17] ),
    .A1(net955),
    .S(_06603_),
    .X(_02232_));
 sg13g2_mux2_1 _25420_ (.A0(\cpu.icache.r_data[7][18] ),
    .A1(net957),
    .S(_06603_),
    .X(_02233_));
 sg13g2_mux2_1 _25421_ (.A0(\cpu.icache.r_data[7][19] ),
    .A1(net956),
    .S(_06603_),
    .X(_02234_));
 sg13g2_mux2_1 _25422_ (.A0(\cpu.icache.r_data[7][1] ),
    .A1(net955),
    .S(_06600_),
    .X(_02235_));
 sg13g2_nor2_2 _25423_ (.A(_06599_),
    .B(_06524_),
    .Y(_06604_));
 sg13g2_mux2_1 _25424_ (.A0(\cpu.icache.r_data[7][20] ),
    .A1(net958),
    .S(_06604_),
    .X(_02236_));
 sg13g2_mux2_1 _25425_ (.A0(\cpu.icache.r_data[7][21] ),
    .A1(_06583_),
    .S(_06604_),
    .X(_02237_));
 sg13g2_mux2_1 _25426_ (.A0(\cpu.icache.r_data[7][22] ),
    .A1(_06581_),
    .S(_06604_),
    .X(_02238_));
 sg13g2_mux2_1 _25427_ (.A0(\cpu.icache.r_data[7][23] ),
    .A1(net956),
    .S(_06604_),
    .X(_02239_));
 sg13g2_nor2_1 _25428_ (.A(_06599_),
    .B(_06527_),
    .Y(_06605_));
 sg13g2_buf_2 _25429_ (.A(_06605_),
    .X(_06606_));
 sg13g2_mux2_1 _25430_ (.A0(\cpu.icache.r_data[7][24] ),
    .A1(net1022),
    .S(_06606_),
    .X(_02240_));
 sg13g2_mux2_1 _25431_ (.A0(\cpu.icache.r_data[7][25] ),
    .A1(net1019),
    .S(_06606_),
    .X(_02241_));
 sg13g2_mux2_1 _25432_ (.A0(\cpu.icache.r_data[7][26] ),
    .A1(net1021),
    .S(_06606_),
    .X(_02242_));
 sg13g2_mux2_1 _25433_ (.A0(\cpu.icache.r_data[7][27] ),
    .A1(net1020),
    .S(_06606_),
    .X(_02243_));
 sg13g2_nor2_2 _25434_ (.A(_06599_),
    .B(_06530_),
    .Y(_06607_));
 sg13g2_mux2_1 _25435_ (.A0(\cpu.icache.r_data[7][28] ),
    .A1(net1022),
    .S(_06607_),
    .X(_02244_));
 sg13g2_mux2_1 _25436_ (.A0(\cpu.icache.r_data[7][29] ),
    .A1(net1019),
    .S(_06607_),
    .X(_02245_));
 sg13g2_mux2_1 _25437_ (.A0(\cpu.icache.r_data[7][2] ),
    .A1(net1021),
    .S(_06600_),
    .X(_02246_));
 sg13g2_mux2_1 _25438_ (.A0(\cpu.icache.r_data[7][30] ),
    .A1(_12218_),
    .S(_06607_),
    .X(_02247_));
 sg13g2_mux2_1 _25439_ (.A0(\cpu.icache.r_data[7][31] ),
    .A1(net1020),
    .S(_06607_),
    .X(_02248_));
 sg13g2_mux2_1 _25440_ (.A0(\cpu.icache.r_data[7][3] ),
    .A1(_12225_),
    .S(_06600_),
    .X(_02249_));
 sg13g2_nor2_2 _25441_ (.A(_06599_),
    .B(_06532_),
    .Y(_06608_));
 sg13g2_mux2_1 _25442_ (.A0(\cpu.icache.r_data[7][4] ),
    .A1(_12205_),
    .S(_06608_),
    .X(_02250_));
 sg13g2_mux2_1 _25443_ (.A0(\cpu.icache.r_data[7][5] ),
    .A1(_12236_),
    .S(_06608_),
    .X(_02251_));
 sg13g2_mux2_1 _25444_ (.A0(\cpu.icache.r_data[7][6] ),
    .A1(_12218_),
    .S(_06608_),
    .X(_02252_));
 sg13g2_mux2_1 _25445_ (.A0(\cpu.icache.r_data[7][7] ),
    .A1(_12225_),
    .S(_06608_),
    .X(_02253_));
 sg13g2_mux2_1 _25446_ (.A0(\cpu.icache.r_data[7][8] ),
    .A1(_12205_),
    .S(_06601_),
    .X(_02254_));
 sg13g2_mux2_1 _25447_ (.A0(\cpu.icache.r_data[7][9] ),
    .A1(_12236_),
    .S(_06601_),
    .X(_02255_));
 sg13g2_mux2_1 _25448_ (.A0(net989),
    .A1(\cpu.icache.r_tag[0][5] ),
    .S(net381),
    .X(_02259_));
 sg13g2_buf_1 _25449_ (.A(net439),
    .X(_06609_));
 sg13g2_buf_1 _25450_ (.A(_06496_),
    .X(_06610_));
 sg13g2_nand2_1 _25451_ (.Y(_06611_),
    .A(\cpu.icache.r_tag[0][15] ),
    .B(net438));
 sg13g2_o21ai_1 _25452_ (.B1(_06611_),
    .Y(_02260_),
    .A1(net428),
    .A2(net379));
 sg13g2_nand2_1 _25453_ (.Y(_06612_),
    .A(\cpu.icache.r_tag[0][16] ),
    .B(net438));
 sg13g2_o21ai_1 _25454_ (.B1(_06612_),
    .Y(_02261_),
    .A1(net465),
    .A2(net379));
 sg13g2_nand2_1 _25455_ (.Y(_06613_),
    .A(\cpu.icache.r_tag[0][17] ),
    .B(net438));
 sg13g2_o21ai_1 _25456_ (.B1(_06613_),
    .Y(_02262_),
    .A1(net370),
    .A2(net379));
 sg13g2_nand2_1 _25457_ (.Y(_06614_),
    .A(\cpu.icache.r_tag[0][18] ),
    .B(net438));
 sg13g2_o21ai_1 _25458_ (.B1(_06614_),
    .Y(_02263_),
    .A1(_08603_),
    .A2(net379));
 sg13g2_nand2_1 _25459_ (.Y(_06615_),
    .A(\cpu.icache.r_tag[0][19] ),
    .B(_06610_));
 sg13g2_o21ai_1 _25460_ (.B1(_06615_),
    .Y(_02264_),
    .A1(net427),
    .A2(_06609_));
 sg13g2_nand2_1 _25461_ (.Y(_06616_),
    .A(\cpu.icache.r_tag[0][20] ),
    .B(_06610_));
 sg13g2_o21ai_1 _25462_ (.B1(_06616_),
    .Y(_02265_),
    .A1(net425),
    .A2(net379));
 sg13g2_nand2_1 _25463_ (.Y(_06617_),
    .A(\cpu.icache.r_tag[0][21] ),
    .B(net439));
 sg13g2_o21ai_1 _25464_ (.B1(_06617_),
    .Y(_02266_),
    .A1(net464),
    .A2(net379));
 sg13g2_nand2_1 _25465_ (.Y(_06618_),
    .A(\cpu.icache.r_tag[0][22] ),
    .B(net439));
 sg13g2_o21ai_1 _25466_ (.B1(_06618_),
    .Y(_02267_),
    .A1(net424),
    .A2(net379));
 sg13g2_nand2_1 _25467_ (.Y(_06619_),
    .A(\cpu.icache.r_tag[0][23] ),
    .B(_06497_));
 sg13g2_o21ai_1 _25468_ (.B1(_06619_),
    .Y(_02268_),
    .A1(net519),
    .A2(net379));
 sg13g2_mux2_1 _25469_ (.A0(net988),
    .A1(\cpu.icache.r_tag[0][6] ),
    .S(net438),
    .X(_02269_));
 sg13g2_mux2_1 _25470_ (.A0(net987),
    .A1(\cpu.icache.r_tag[0][7] ),
    .S(net438),
    .X(_02270_));
 sg13g2_nand2_1 _25471_ (.Y(_06620_),
    .A(\cpu.icache.r_tag[0][8] ),
    .B(net439));
 sg13g2_o21ai_1 _25472_ (.B1(_06620_),
    .Y(_02271_),
    .A1(net1078),
    .A2(net381));
 sg13g2_mux2_1 _25473_ (.A0(net986),
    .A1(\cpu.icache.r_tag[0][9] ),
    .S(net438),
    .X(_02272_));
 sg13g2_mux2_1 _25474_ (.A0(net985),
    .A1(\cpu.icache.r_tag[0][10] ),
    .S(net438),
    .X(_02273_));
 sg13g2_nand2_1 _25475_ (.Y(_06621_),
    .A(\cpu.icache.r_tag[0][11] ),
    .B(net439));
 sg13g2_o21ai_1 _25476_ (.B1(_06621_),
    .Y(_02274_),
    .A1(net1077),
    .A2(net381));
 sg13g2_nand2_1 _25477_ (.Y(_06622_),
    .A(\cpu.icache.r_tag[0][12] ),
    .B(net439));
 sg13g2_o21ai_1 _25478_ (.B1(_06622_),
    .Y(_02275_),
    .A1(net430),
    .A2(net381));
 sg13g2_nand2_1 _25479_ (.Y(_06623_),
    .A(\cpu.icache.r_tag[0][13] ),
    .B(net439));
 sg13g2_o21ai_1 _25480_ (.B1(_06623_),
    .Y(_02276_),
    .A1(net431),
    .A2(_06498_));
 sg13g2_nand2_1 _25481_ (.Y(_06624_),
    .A(\cpu.icache.r_tag[0][14] ),
    .B(_06497_));
 sg13g2_o21ai_1 _25482_ (.B1(_06624_),
    .Y(_02277_),
    .A1(net426),
    .A2(_06498_));
 sg13g2_nor2b_1 _25483_ (.A(_06475_),
    .B_N(_06486_),
    .Y(_06625_));
 sg13g2_buf_1 _25484_ (.A(_06625_),
    .X(_06626_));
 sg13g2_nand2_1 _25485_ (.Y(_06627_),
    .A(_09010_),
    .B(_06626_));
 sg13g2_buf_1 _25486_ (.A(_06627_),
    .X(_06628_));
 sg13g2_buf_1 _25487_ (.A(_06628_),
    .X(_06629_));
 sg13g2_mux2_1 _25488_ (.A0(net989),
    .A1(\cpu.icache.r_tag[1][5] ),
    .S(_06629_),
    .X(_02278_));
 sg13g2_buf_1 _25489_ (.A(_06628_),
    .X(_06630_));
 sg13g2_nand2_1 _25490_ (.Y(_06631_),
    .A(\cpu.icache.r_tag[1][15] ),
    .B(net378));
 sg13g2_o21ai_1 _25491_ (.B1(_06631_),
    .Y(_02279_),
    .A1(net428),
    .A2(net377));
 sg13g2_buf_1 _25492_ (.A(_06628_),
    .X(_06632_));
 sg13g2_nand2_1 _25493_ (.Y(_06633_),
    .A(\cpu.icache.r_tag[1][16] ),
    .B(net376));
 sg13g2_o21ai_1 _25494_ (.B1(_06633_),
    .Y(_02280_),
    .A1(net465),
    .A2(net377));
 sg13g2_nand2_1 _25495_ (.Y(_06634_),
    .A(\cpu.icache.r_tag[1][17] ),
    .B(net376));
 sg13g2_o21ai_1 _25496_ (.B1(_06634_),
    .Y(_02281_),
    .A1(net370),
    .A2(net377));
 sg13g2_nand2_1 _25497_ (.Y(_06635_),
    .A(\cpu.icache.r_tag[1][18] ),
    .B(net376));
 sg13g2_o21ai_1 _25498_ (.B1(_06635_),
    .Y(_02282_),
    .A1(net429),
    .A2(net377));
 sg13g2_nand2_1 _25499_ (.Y(_06636_),
    .A(\cpu.icache.r_tag[1][19] ),
    .B(net376));
 sg13g2_o21ai_1 _25500_ (.B1(_06636_),
    .Y(_02283_),
    .A1(net427),
    .A2(net377));
 sg13g2_nand2_1 _25501_ (.Y(_06637_),
    .A(\cpu.icache.r_tag[1][20] ),
    .B(_06632_));
 sg13g2_o21ai_1 _25502_ (.B1(_06637_),
    .Y(_02284_),
    .A1(net425),
    .A2(_06630_));
 sg13g2_nand2_1 _25503_ (.Y(_06638_),
    .A(\cpu.icache.r_tag[1][21] ),
    .B(net376));
 sg13g2_o21ai_1 _25504_ (.B1(_06638_),
    .Y(_02285_),
    .A1(net464),
    .A2(net377));
 sg13g2_nand2_1 _25505_ (.Y(_06639_),
    .A(\cpu.icache.r_tag[1][22] ),
    .B(_06632_));
 sg13g2_o21ai_1 _25506_ (.B1(_06639_),
    .Y(_02286_),
    .A1(net424),
    .A2(_06630_));
 sg13g2_nand2_1 _25507_ (.Y(_06640_),
    .A(\cpu.icache.r_tag[1][23] ),
    .B(net376));
 sg13g2_o21ai_1 _25508_ (.B1(_06640_),
    .Y(_02287_),
    .A1(net519),
    .A2(net377));
 sg13g2_mux2_1 _25509_ (.A0(net988),
    .A1(\cpu.icache.r_tag[1][6] ),
    .S(net378),
    .X(_02288_));
 sg13g2_mux2_1 _25510_ (.A0(net987),
    .A1(\cpu.icache.r_tag[1][7] ),
    .S(net378),
    .X(_02289_));
 sg13g2_nand2_1 _25511_ (.Y(_06641_),
    .A(\cpu.icache.r_tag[1][8] ),
    .B(net376));
 sg13g2_o21ai_1 _25512_ (.B1(_06641_),
    .Y(_02290_),
    .A1(net1078),
    .A2(net377));
 sg13g2_mux2_1 _25513_ (.A0(net986),
    .A1(\cpu.icache.r_tag[1][9] ),
    .S(_06629_),
    .X(_02291_));
 sg13g2_mux2_1 _25514_ (.A0(net985),
    .A1(\cpu.icache.r_tag[1][10] ),
    .S(net378),
    .X(_02292_));
 sg13g2_nand2_1 _25515_ (.Y(_06642_),
    .A(\cpu.icache.r_tag[1][11] ),
    .B(net376));
 sg13g2_o21ai_1 _25516_ (.B1(_06642_),
    .Y(_02293_),
    .A1(net1077),
    .A2(net378));
 sg13g2_nand2_1 _25517_ (.Y(_06643_),
    .A(\cpu.icache.r_tag[1][12] ),
    .B(_06628_));
 sg13g2_o21ai_1 _25518_ (.B1(_06643_),
    .Y(_02294_),
    .A1(net430),
    .A2(net378));
 sg13g2_nand2_1 _25519_ (.Y(_06644_),
    .A(\cpu.icache.r_tag[1][13] ),
    .B(_06628_));
 sg13g2_o21ai_1 _25520_ (.B1(_06644_),
    .Y(_02295_),
    .A1(net431),
    .A2(net378));
 sg13g2_nand2_1 _25521_ (.Y(_06645_),
    .A(\cpu.icache.r_tag[1][14] ),
    .B(_06628_));
 sg13g2_o21ai_1 _25522_ (.B1(_06645_),
    .Y(_02296_),
    .A1(net426),
    .A2(net378));
 sg13g2_nand2_1 _25523_ (.Y(_06646_),
    .A(_08800_),
    .B(_06626_));
 sg13g2_buf_1 _25524_ (.A(_06646_),
    .X(_06647_));
 sg13g2_buf_1 _25525_ (.A(_06647_),
    .X(_06648_));
 sg13g2_mux2_1 _25526_ (.A0(net989),
    .A1(\cpu.icache.r_tag[2][5] ),
    .S(net375),
    .X(_02297_));
 sg13g2_buf_1 _25527_ (.A(_06647_),
    .X(_06649_));
 sg13g2_nand2_1 _25528_ (.Y(_06650_),
    .A(\cpu.icache.r_tag[2][15] ),
    .B(net375));
 sg13g2_o21ai_1 _25529_ (.B1(_06650_),
    .Y(_02298_),
    .A1(net428),
    .A2(net374));
 sg13g2_buf_1 _25530_ (.A(_06647_),
    .X(_06651_));
 sg13g2_nand2_1 _25531_ (.Y(_06652_),
    .A(\cpu.icache.r_tag[2][16] ),
    .B(net373));
 sg13g2_o21ai_1 _25532_ (.B1(_06652_),
    .Y(_02299_),
    .A1(net465),
    .A2(net374));
 sg13g2_nand2_1 _25533_ (.Y(_06653_),
    .A(\cpu.icache.r_tag[2][17] ),
    .B(net373));
 sg13g2_o21ai_1 _25534_ (.B1(_06653_),
    .Y(_02300_),
    .A1(net370),
    .A2(_06649_));
 sg13g2_nand2_1 _25535_ (.Y(_06654_),
    .A(\cpu.icache.r_tag[2][18] ),
    .B(net373));
 sg13g2_o21ai_1 _25536_ (.B1(_06654_),
    .Y(_02301_),
    .A1(net429),
    .A2(net374));
 sg13g2_nand2_1 _25537_ (.Y(_06655_),
    .A(\cpu.icache.r_tag[2][19] ),
    .B(net373));
 sg13g2_o21ai_1 _25538_ (.B1(_06655_),
    .Y(_02302_),
    .A1(net427),
    .A2(net374));
 sg13g2_nand2_1 _25539_ (.Y(_06656_),
    .A(\cpu.icache.r_tag[2][20] ),
    .B(net373));
 sg13g2_o21ai_1 _25540_ (.B1(_06656_),
    .Y(_02303_),
    .A1(net425),
    .A2(net374));
 sg13g2_nand2_1 _25541_ (.Y(_06657_),
    .A(\cpu.icache.r_tag[2][21] ),
    .B(net373));
 sg13g2_o21ai_1 _25542_ (.B1(_06657_),
    .Y(_02304_),
    .A1(net464),
    .A2(net374));
 sg13g2_nand2_1 _25543_ (.Y(_06658_),
    .A(\cpu.icache.r_tag[2][22] ),
    .B(_06651_));
 sg13g2_o21ai_1 _25544_ (.B1(_06658_),
    .Y(_02305_),
    .A1(net424),
    .A2(_06649_));
 sg13g2_nand2_1 _25545_ (.Y(_06659_),
    .A(\cpu.icache.r_tag[2][23] ),
    .B(net373));
 sg13g2_o21ai_1 _25546_ (.B1(_06659_),
    .Y(_02306_),
    .A1(net519),
    .A2(net374));
 sg13g2_mux2_1 _25547_ (.A0(net988),
    .A1(\cpu.icache.r_tag[2][6] ),
    .S(net375),
    .X(_02307_));
 sg13g2_mux2_1 _25548_ (.A0(net987),
    .A1(\cpu.icache.r_tag[2][7] ),
    .S(net375),
    .X(_02308_));
 sg13g2_nand2_1 _25549_ (.Y(_06660_),
    .A(\cpu.icache.r_tag[2][8] ),
    .B(net373));
 sg13g2_o21ai_1 _25550_ (.B1(_06660_),
    .Y(_02309_),
    .A1(net1078),
    .A2(net374));
 sg13g2_mux2_1 _25551_ (.A0(net986),
    .A1(\cpu.icache.r_tag[2][9] ),
    .S(net375),
    .X(_02310_));
 sg13g2_mux2_1 _25552_ (.A0(net985),
    .A1(\cpu.icache.r_tag[2][10] ),
    .S(net375),
    .X(_02311_));
 sg13g2_nand2_1 _25553_ (.Y(_06661_),
    .A(\cpu.icache.r_tag[2][11] ),
    .B(_06651_));
 sg13g2_o21ai_1 _25554_ (.B1(_06661_),
    .Y(_02312_),
    .A1(net1077),
    .A2(_06648_));
 sg13g2_nand2_1 _25555_ (.Y(_06662_),
    .A(\cpu.icache.r_tag[2][12] ),
    .B(_06647_));
 sg13g2_o21ai_1 _25556_ (.B1(_06662_),
    .Y(_02313_),
    .A1(net430),
    .A2(net375));
 sg13g2_nand2_1 _25557_ (.Y(_06663_),
    .A(\cpu.icache.r_tag[2][13] ),
    .B(_06647_));
 sg13g2_o21ai_1 _25558_ (.B1(_06663_),
    .Y(_02314_),
    .A1(net431),
    .A2(net375));
 sg13g2_nand2_1 _25559_ (.Y(_06664_),
    .A(\cpu.icache.r_tag[2][14] ),
    .B(_06647_));
 sg13g2_o21ai_1 _25560_ (.B1(_06664_),
    .Y(_02315_),
    .A1(net426),
    .A2(_06648_));
 sg13g2_mux2_1 _25561_ (.A0(net989),
    .A1(\cpu.icache.r_tag[3][5] ),
    .S(net295),
    .X(_02316_));
 sg13g2_buf_1 _25562_ (.A(net380),
    .X(_06665_));
 sg13g2_buf_1 _25563_ (.A(_06559_),
    .X(_06666_));
 sg13g2_nand2_1 _25564_ (.Y(_06667_),
    .A(\cpu.icache.r_tag[3][15] ),
    .B(net372));
 sg13g2_o21ai_1 _25565_ (.B1(_06667_),
    .Y(_02317_),
    .A1(net428),
    .A2(net294));
 sg13g2_nand2_1 _25566_ (.Y(_06668_),
    .A(\cpu.icache.r_tag[3][16] ),
    .B(net372));
 sg13g2_o21ai_1 _25567_ (.B1(_06668_),
    .Y(_02318_),
    .A1(net465),
    .A2(net294));
 sg13g2_nand2_1 _25568_ (.Y(_06669_),
    .A(\cpu.icache.r_tag[3][17] ),
    .B(_06666_));
 sg13g2_o21ai_1 _25569_ (.B1(_06669_),
    .Y(_02319_),
    .A1(net370),
    .A2(net294));
 sg13g2_nand2_1 _25570_ (.Y(_06670_),
    .A(\cpu.icache.r_tag[3][18] ),
    .B(net372));
 sg13g2_o21ai_1 _25571_ (.B1(_06670_),
    .Y(_02320_),
    .A1(net429),
    .A2(net294));
 sg13g2_nand2_1 _25572_ (.Y(_06671_),
    .A(\cpu.icache.r_tag[3][19] ),
    .B(_06666_));
 sg13g2_o21ai_1 _25573_ (.B1(_06671_),
    .Y(_02321_),
    .A1(net427),
    .A2(_06665_));
 sg13g2_nand2_1 _25574_ (.Y(_06672_),
    .A(\cpu.icache.r_tag[3][20] ),
    .B(net372));
 sg13g2_o21ai_1 _25575_ (.B1(_06672_),
    .Y(_02322_),
    .A1(net425),
    .A2(_06665_));
 sg13g2_nand2_1 _25576_ (.Y(_06673_),
    .A(\cpu.icache.r_tag[3][21] ),
    .B(net380));
 sg13g2_o21ai_1 _25577_ (.B1(_06673_),
    .Y(_02323_),
    .A1(net464),
    .A2(net294));
 sg13g2_nand2_1 _25578_ (.Y(_06674_),
    .A(\cpu.icache.r_tag[3][22] ),
    .B(_06560_));
 sg13g2_o21ai_1 _25579_ (.B1(_06674_),
    .Y(_02324_),
    .A1(net424),
    .A2(net294));
 sg13g2_nand2_1 _25580_ (.Y(_06675_),
    .A(\cpu.icache.r_tag[3][23] ),
    .B(net380));
 sg13g2_o21ai_1 _25581_ (.B1(_06675_),
    .Y(_02325_),
    .A1(net519),
    .A2(net294));
 sg13g2_mux2_1 _25582_ (.A0(net988),
    .A1(\cpu.icache.r_tag[3][6] ),
    .S(net372),
    .X(_02326_));
 sg13g2_mux2_1 _25583_ (.A0(net987),
    .A1(\cpu.icache.r_tag[3][7] ),
    .S(net372),
    .X(_02327_));
 sg13g2_nand2_1 _25584_ (.Y(_06676_),
    .A(\cpu.icache.r_tag[3][8] ),
    .B(net380));
 sg13g2_o21ai_1 _25585_ (.B1(_06676_),
    .Y(_02328_),
    .A1(net1078),
    .A2(_06561_));
 sg13g2_mux2_1 _25586_ (.A0(net986),
    .A1(\cpu.icache.r_tag[3][9] ),
    .S(net372),
    .X(_02329_));
 sg13g2_mux2_1 _25587_ (.A0(net985),
    .A1(\cpu.icache.r_tag[3][10] ),
    .S(net372),
    .X(_02330_));
 sg13g2_nand2_1 _25588_ (.Y(_06677_),
    .A(\cpu.icache.r_tag[3][11] ),
    .B(net380));
 sg13g2_o21ai_1 _25589_ (.B1(_06677_),
    .Y(_02331_),
    .A1(net1077),
    .A2(_06561_));
 sg13g2_nand2_1 _25590_ (.Y(_06678_),
    .A(\cpu.icache.r_tag[3][12] ),
    .B(net380));
 sg13g2_o21ai_1 _25591_ (.B1(_06678_),
    .Y(_02332_),
    .A1(net430),
    .A2(net295));
 sg13g2_nand2_1 _25592_ (.Y(_06679_),
    .A(\cpu.icache.r_tag[3][13] ),
    .B(net380));
 sg13g2_o21ai_1 _25593_ (.B1(_06679_),
    .Y(_02333_),
    .A1(_08497_),
    .A2(net295));
 sg13g2_nand2_1 _25594_ (.Y(_06680_),
    .A(\cpu.icache.r_tag[3][14] ),
    .B(net380));
 sg13g2_o21ai_1 _25595_ (.B1(_06680_),
    .Y(_02334_),
    .A1(net426),
    .A2(net295));
 sg13g2_nand2_1 _25596_ (.Y(_06681_),
    .A(_09035_),
    .B(_06626_));
 sg13g2_buf_1 _25597_ (.A(_06681_),
    .X(_06682_));
 sg13g2_buf_1 _25598_ (.A(_06682_),
    .X(_06683_));
 sg13g2_mux2_1 _25599_ (.A0(net989),
    .A1(\cpu.icache.r_tag[4][5] ),
    .S(net437),
    .X(_02335_));
 sg13g2_buf_1 _25600_ (.A(_06682_),
    .X(_06684_));
 sg13g2_nand2_1 _25601_ (.Y(_06685_),
    .A(\cpu.icache.r_tag[4][15] ),
    .B(net437));
 sg13g2_o21ai_1 _25602_ (.B1(_06685_),
    .Y(_02336_),
    .A1(net428),
    .A2(net436));
 sg13g2_buf_1 _25603_ (.A(_06682_),
    .X(_06686_));
 sg13g2_nand2_1 _25604_ (.Y(_06687_),
    .A(\cpu.icache.r_tag[4][16] ),
    .B(net435));
 sg13g2_o21ai_1 _25605_ (.B1(_06687_),
    .Y(_02337_),
    .A1(net465),
    .A2(net436));
 sg13g2_nand2_1 _25606_ (.Y(_06688_),
    .A(\cpu.icache.r_tag[4][17] ),
    .B(net435));
 sg13g2_o21ai_1 _25607_ (.B1(_06688_),
    .Y(_02338_),
    .A1(net370),
    .A2(net436));
 sg13g2_nand2_1 _25608_ (.Y(_06689_),
    .A(\cpu.icache.r_tag[4][18] ),
    .B(net435));
 sg13g2_o21ai_1 _25609_ (.B1(_06689_),
    .Y(_02339_),
    .A1(net429),
    .A2(net436));
 sg13g2_nand2_1 _25610_ (.Y(_06690_),
    .A(\cpu.icache.r_tag[4][19] ),
    .B(net435));
 sg13g2_o21ai_1 _25611_ (.B1(_06690_),
    .Y(_02340_),
    .A1(net427),
    .A2(net436));
 sg13g2_nand2_1 _25612_ (.Y(_06691_),
    .A(\cpu.icache.r_tag[4][20] ),
    .B(_06686_));
 sg13g2_o21ai_1 _25613_ (.B1(_06691_),
    .Y(_02341_),
    .A1(net425),
    .A2(_06684_));
 sg13g2_nand2_1 _25614_ (.Y(_06692_),
    .A(\cpu.icache.r_tag[4][21] ),
    .B(net435));
 sg13g2_o21ai_1 _25615_ (.B1(_06692_),
    .Y(_02342_),
    .A1(net464),
    .A2(net436));
 sg13g2_nand2_1 _25616_ (.Y(_06693_),
    .A(\cpu.icache.r_tag[4][22] ),
    .B(_06686_));
 sg13g2_o21ai_1 _25617_ (.B1(_06693_),
    .Y(_02343_),
    .A1(net424),
    .A2(_06684_));
 sg13g2_nand2_1 _25618_ (.Y(_06694_),
    .A(\cpu.icache.r_tag[4][23] ),
    .B(net435));
 sg13g2_o21ai_1 _25619_ (.B1(_06694_),
    .Y(_02344_),
    .A1(net519),
    .A2(net436));
 sg13g2_mux2_1 _25620_ (.A0(net988),
    .A1(\cpu.icache.r_tag[4][6] ),
    .S(net437),
    .X(_02345_));
 sg13g2_mux2_1 _25621_ (.A0(net987),
    .A1(\cpu.icache.r_tag[4][7] ),
    .S(_06683_),
    .X(_02346_));
 sg13g2_nand2_1 _25622_ (.Y(_06695_),
    .A(\cpu.icache.r_tag[4][8] ),
    .B(net435));
 sg13g2_o21ai_1 _25623_ (.B1(_06695_),
    .Y(_02347_),
    .A1(net1078),
    .A2(net436));
 sg13g2_mux2_1 _25624_ (.A0(net986),
    .A1(\cpu.icache.r_tag[4][9] ),
    .S(_06683_),
    .X(_02348_));
 sg13g2_mux2_1 _25625_ (.A0(net985),
    .A1(\cpu.icache.r_tag[4][10] ),
    .S(net437),
    .X(_02349_));
 sg13g2_nand2_1 _25626_ (.Y(_06696_),
    .A(\cpu.icache.r_tag[4][11] ),
    .B(net435));
 sg13g2_o21ai_1 _25627_ (.B1(_06696_),
    .Y(_02350_),
    .A1(net1077),
    .A2(net437));
 sg13g2_nand2_1 _25628_ (.Y(_06697_),
    .A(\cpu.icache.r_tag[4][12] ),
    .B(_06682_));
 sg13g2_o21ai_1 _25629_ (.B1(_06697_),
    .Y(_02351_),
    .A1(net430),
    .A2(net437));
 sg13g2_nand2_1 _25630_ (.Y(_06698_),
    .A(\cpu.icache.r_tag[4][13] ),
    .B(_06682_));
 sg13g2_o21ai_1 _25631_ (.B1(_06698_),
    .Y(_02352_),
    .A1(net431),
    .A2(net437));
 sg13g2_nand2_1 _25632_ (.Y(_06699_),
    .A(\cpu.icache.r_tag[4][14] ),
    .B(_06682_));
 sg13g2_o21ai_1 _25633_ (.B1(_06699_),
    .Y(_02353_),
    .A1(net426),
    .A2(net437));
 sg13g2_nand2_1 _25634_ (.Y(_06700_),
    .A(_08518_),
    .B(_06626_));
 sg13g2_buf_1 _25635_ (.A(_06700_),
    .X(_06701_));
 sg13g2_buf_1 _25636_ (.A(_06701_),
    .X(_06702_));
 sg13g2_mux2_1 _25637_ (.A0(net989),
    .A1(\cpu.icache.r_tag[5][5] ),
    .S(net473),
    .X(_02354_));
 sg13g2_buf_1 _25638_ (.A(_06701_),
    .X(_06703_));
 sg13g2_nand2_1 _25639_ (.Y(_06704_),
    .A(\cpu.icache.r_tag[5][15] ),
    .B(net473));
 sg13g2_o21ai_1 _25640_ (.B1(_06704_),
    .Y(_02355_),
    .A1(net428),
    .A2(net472));
 sg13g2_buf_1 _25641_ (.A(_06701_),
    .X(_06705_));
 sg13g2_nand2_1 _25642_ (.Y(_06706_),
    .A(\cpu.icache.r_tag[5][16] ),
    .B(net471));
 sg13g2_o21ai_1 _25643_ (.B1(_06706_),
    .Y(_02356_),
    .A1(net465),
    .A2(net472));
 sg13g2_nand2_1 _25644_ (.Y(_06707_),
    .A(\cpu.icache.r_tag[5][17] ),
    .B(net471));
 sg13g2_o21ai_1 _25645_ (.B1(_06707_),
    .Y(_02357_),
    .A1(net370),
    .A2(net472));
 sg13g2_nand2_1 _25646_ (.Y(_06708_),
    .A(\cpu.icache.r_tag[5][18] ),
    .B(net471));
 sg13g2_o21ai_1 _25647_ (.B1(_06708_),
    .Y(_02358_),
    .A1(net429),
    .A2(net472));
 sg13g2_nand2_1 _25648_ (.Y(_06709_),
    .A(\cpu.icache.r_tag[5][19] ),
    .B(net471));
 sg13g2_o21ai_1 _25649_ (.B1(_06709_),
    .Y(_02359_),
    .A1(net427),
    .A2(net472));
 sg13g2_nand2_1 _25650_ (.Y(_06710_),
    .A(\cpu.icache.r_tag[5][20] ),
    .B(_06705_));
 sg13g2_o21ai_1 _25651_ (.B1(_06710_),
    .Y(_02360_),
    .A1(net425),
    .A2(_06703_));
 sg13g2_nand2_1 _25652_ (.Y(_06711_),
    .A(\cpu.icache.r_tag[5][21] ),
    .B(net471));
 sg13g2_o21ai_1 _25653_ (.B1(_06711_),
    .Y(_02361_),
    .A1(net464),
    .A2(net472));
 sg13g2_nand2_1 _25654_ (.Y(_06712_),
    .A(\cpu.icache.r_tag[5][22] ),
    .B(net471));
 sg13g2_o21ai_1 _25655_ (.B1(_06712_),
    .Y(_02362_),
    .A1(net424),
    .A2(_06703_));
 sg13g2_nand2_1 _25656_ (.Y(_06713_),
    .A(\cpu.icache.r_tag[5][23] ),
    .B(net471));
 sg13g2_o21ai_1 _25657_ (.B1(_06713_),
    .Y(_02363_),
    .A1(net519),
    .A2(net472));
 sg13g2_mux2_1 _25658_ (.A0(net988),
    .A1(\cpu.icache.r_tag[5][6] ),
    .S(net473),
    .X(_02364_));
 sg13g2_mux2_1 _25659_ (.A0(net987),
    .A1(\cpu.icache.r_tag[5][7] ),
    .S(_06702_),
    .X(_02365_));
 sg13g2_nand2_1 _25660_ (.Y(_06714_),
    .A(\cpu.icache.r_tag[5][8] ),
    .B(net471));
 sg13g2_o21ai_1 _25661_ (.B1(_06714_),
    .Y(_02366_),
    .A1(net1078),
    .A2(net472));
 sg13g2_mux2_1 _25662_ (.A0(net986),
    .A1(\cpu.icache.r_tag[5][9] ),
    .S(_06702_),
    .X(_02367_));
 sg13g2_mux2_1 _25663_ (.A0(net985),
    .A1(\cpu.icache.r_tag[5][10] ),
    .S(net473),
    .X(_02368_));
 sg13g2_nand2_1 _25664_ (.Y(_06715_),
    .A(\cpu.icache.r_tag[5][11] ),
    .B(_06705_));
 sg13g2_o21ai_1 _25665_ (.B1(_06715_),
    .Y(_02369_),
    .A1(net1077),
    .A2(net473));
 sg13g2_nand2_1 _25666_ (.Y(_06716_),
    .A(\cpu.icache.r_tag[5][12] ),
    .B(_06701_));
 sg13g2_o21ai_1 _25667_ (.B1(_06716_),
    .Y(_02370_),
    .A1(net430),
    .A2(net473));
 sg13g2_nand2_1 _25668_ (.Y(_06717_),
    .A(\cpu.icache.r_tag[5][13] ),
    .B(_06701_));
 sg13g2_o21ai_1 _25669_ (.B1(_06717_),
    .Y(_02371_),
    .A1(net431),
    .A2(net473));
 sg13g2_nand2_1 _25670_ (.Y(_06718_),
    .A(\cpu.icache.r_tag[5][14] ),
    .B(_06701_));
 sg13g2_o21ai_1 _25671_ (.B1(_06718_),
    .Y(_02372_),
    .A1(net426),
    .A2(net473));
 sg13g2_nand2_1 _25672_ (.Y(_06719_),
    .A(_09037_),
    .B(_06626_));
 sg13g2_buf_1 _25673_ (.A(_06719_),
    .X(_06720_));
 sg13g2_buf_1 _25674_ (.A(_06720_),
    .X(_06721_));
 sg13g2_mux2_1 _25675_ (.A0(_04612_),
    .A1(\cpu.icache.r_tag[6][5] ),
    .S(net434),
    .X(_02373_));
 sg13g2_buf_1 _25676_ (.A(_06720_),
    .X(_06722_));
 sg13g2_nand2_1 _25677_ (.Y(_06723_),
    .A(\cpu.icache.r_tag[6][15] ),
    .B(net434));
 sg13g2_o21ai_1 _25678_ (.B1(_06723_),
    .Y(_02374_),
    .A1(net428),
    .A2(net433));
 sg13g2_buf_1 _25679_ (.A(_06720_),
    .X(_06724_));
 sg13g2_nand2_1 _25680_ (.Y(_06725_),
    .A(\cpu.icache.r_tag[6][16] ),
    .B(net432));
 sg13g2_o21ai_1 _25681_ (.B1(_06725_),
    .Y(_02375_),
    .A1(net465),
    .A2(net433));
 sg13g2_nand2_1 _25682_ (.Y(_06726_),
    .A(\cpu.icache.r_tag[6][17] ),
    .B(net432));
 sg13g2_o21ai_1 _25683_ (.B1(_06726_),
    .Y(_02376_),
    .A1(net370),
    .A2(_06722_));
 sg13g2_nand2_1 _25684_ (.Y(_06727_),
    .A(\cpu.icache.r_tag[6][18] ),
    .B(net432));
 sg13g2_o21ai_1 _25685_ (.B1(_06727_),
    .Y(_02377_),
    .A1(net429),
    .A2(net433));
 sg13g2_nand2_1 _25686_ (.Y(_06728_),
    .A(\cpu.icache.r_tag[6][19] ),
    .B(net432));
 sg13g2_o21ai_1 _25687_ (.B1(_06728_),
    .Y(_02378_),
    .A1(net427),
    .A2(net433));
 sg13g2_nand2_1 _25688_ (.Y(_06729_),
    .A(\cpu.icache.r_tag[6][20] ),
    .B(_06724_));
 sg13g2_o21ai_1 _25689_ (.B1(_06729_),
    .Y(_02379_),
    .A1(net425),
    .A2(_06722_));
 sg13g2_nand2_1 _25690_ (.Y(_06730_),
    .A(\cpu.icache.r_tag[6][21] ),
    .B(net432));
 sg13g2_o21ai_1 _25691_ (.B1(_06730_),
    .Y(_02380_),
    .A1(_08778_),
    .A2(net433));
 sg13g2_nand2_1 _25692_ (.Y(_06731_),
    .A(\cpu.icache.r_tag[6][22] ),
    .B(net432));
 sg13g2_o21ai_1 _25693_ (.B1(_06731_),
    .Y(_02381_),
    .A1(net424),
    .A2(net433));
 sg13g2_nand2_1 _25694_ (.Y(_06732_),
    .A(\cpu.icache.r_tag[6][23] ),
    .B(net432));
 sg13g2_o21ai_1 _25695_ (.B1(_06732_),
    .Y(_02382_),
    .A1(net519),
    .A2(net433));
 sg13g2_mux2_1 _25696_ (.A0(_04646_),
    .A1(\cpu.icache.r_tag[6][6] ),
    .S(net434),
    .X(_02383_));
 sg13g2_mux2_1 _25697_ (.A0(_04675_),
    .A1(\cpu.icache.r_tag[6][7] ),
    .S(_06721_),
    .X(_02384_));
 sg13g2_nand2_1 _25698_ (.Y(_06733_),
    .A(\cpu.icache.r_tag[6][8] ),
    .B(net432));
 sg13g2_o21ai_1 _25699_ (.B1(_06733_),
    .Y(_02385_),
    .A1(net1078),
    .A2(net433));
 sg13g2_mux2_1 _25700_ (.A0(_04741_),
    .A1(\cpu.icache.r_tag[6][9] ),
    .S(_06721_),
    .X(_02386_));
 sg13g2_mux2_1 _25701_ (.A0(_04774_),
    .A1(\cpu.icache.r_tag[6][10] ),
    .S(net434),
    .X(_02387_));
 sg13g2_nand2_1 _25702_ (.Y(_06734_),
    .A(\cpu.icache.r_tag[6][11] ),
    .B(_06724_));
 sg13g2_o21ai_1 _25703_ (.B1(_06734_),
    .Y(_02388_),
    .A1(_08731_),
    .A2(net434));
 sg13g2_nand2_1 _25704_ (.Y(_06735_),
    .A(\cpu.icache.r_tag[6][12] ),
    .B(_06720_));
 sg13g2_o21ai_1 _25705_ (.B1(_06735_),
    .Y(_02389_),
    .A1(net430),
    .A2(net434));
 sg13g2_nand2_1 _25706_ (.Y(_06736_),
    .A(\cpu.icache.r_tag[6][13] ),
    .B(_06720_));
 sg13g2_o21ai_1 _25707_ (.B1(_06736_),
    .Y(_02390_),
    .A1(net431),
    .A2(net434));
 sg13g2_nand2_1 _25708_ (.Y(_06737_),
    .A(\cpu.icache.r_tag[6][14] ),
    .B(_06720_));
 sg13g2_o21ai_1 _25709_ (.B1(_06737_),
    .Y(_02391_),
    .A1(net426),
    .A2(net434));
 sg13g2_nand2_1 _25710_ (.Y(_06738_),
    .A(_08639_),
    .B(_06626_));
 sg13g2_buf_1 _25711_ (.A(_06738_),
    .X(_06739_));
 sg13g2_buf_1 _25712_ (.A(_06739_),
    .X(_06740_));
 sg13g2_mux2_1 _25713_ (.A0(_04612_),
    .A1(\cpu.icache.r_tag[7][5] ),
    .S(net470),
    .X(_02392_));
 sg13g2_buf_1 _25714_ (.A(_06739_),
    .X(_06741_));
 sg13g2_nand2_1 _25715_ (.Y(_06742_),
    .A(\cpu.icache.r_tag[7][15] ),
    .B(net470));
 sg13g2_o21ai_1 _25716_ (.B1(_06742_),
    .Y(_02393_),
    .A1(_08663_),
    .A2(net469));
 sg13g2_buf_1 _25717_ (.A(_06739_),
    .X(_06743_));
 sg13g2_nand2_1 _25718_ (.Y(_06744_),
    .A(\cpu.icache.r_tag[7][16] ),
    .B(net468));
 sg13g2_o21ai_1 _25719_ (.B1(_06744_),
    .Y(_02394_),
    .A1(net465),
    .A2(net469));
 sg13g2_nand2_1 _25720_ (.Y(_06745_),
    .A(\cpu.icache.r_tag[7][17] ),
    .B(net468));
 sg13g2_o21ai_1 _25721_ (.B1(_06745_),
    .Y(_02395_),
    .A1(_09091_),
    .A2(net469));
 sg13g2_nand2_1 _25722_ (.Y(_06746_),
    .A(\cpu.icache.r_tag[7][18] ),
    .B(net468));
 sg13g2_o21ai_1 _25723_ (.B1(_06746_),
    .Y(_02396_),
    .A1(net429),
    .A2(net469));
 sg13g2_nand2_1 _25724_ (.Y(_06747_),
    .A(\cpu.icache.r_tag[7][19] ),
    .B(net468));
 sg13g2_o21ai_1 _25725_ (.B1(_06747_),
    .Y(_02397_),
    .A1(_08820_),
    .A2(_06741_));
 sg13g2_nand2_1 _25726_ (.Y(_06748_),
    .A(\cpu.icache.r_tag[7][20] ),
    .B(_06743_));
 sg13g2_o21ai_1 _25727_ (.B1(_06748_),
    .Y(_02398_),
    .A1(_08869_),
    .A2(_06741_));
 sg13g2_nand2_1 _25728_ (.Y(_06749_),
    .A(\cpu.icache.r_tag[7][21] ),
    .B(net468));
 sg13g2_o21ai_1 _25729_ (.B1(_06749_),
    .Y(_02399_),
    .A1(net464),
    .A2(net469));
 sg13g2_nand2_1 _25730_ (.Y(_06750_),
    .A(\cpu.icache.r_tag[7][22] ),
    .B(net468));
 sg13g2_o21ai_1 _25731_ (.B1(_06750_),
    .Y(_02400_),
    .A1(_08890_),
    .A2(net469));
 sg13g2_nand2_1 _25732_ (.Y(_06751_),
    .A(\cpu.icache.r_tag[7][23] ),
    .B(net468));
 sg13g2_o21ai_1 _25733_ (.B1(_06751_),
    .Y(_02401_),
    .A1(_08799_),
    .A2(net469));
 sg13g2_mux2_1 _25734_ (.A0(_04646_),
    .A1(\cpu.icache.r_tag[7][6] ),
    .S(net470),
    .X(_02402_));
 sg13g2_mux2_1 _25735_ (.A0(_04675_),
    .A1(\cpu.icache.r_tag[7][7] ),
    .S(_06740_),
    .X(_02403_));
 sg13g2_nand2_1 _25736_ (.Y(_06752_),
    .A(\cpu.icache.r_tag[7][8] ),
    .B(net468));
 sg13g2_o21ai_1 _25737_ (.B1(_06752_),
    .Y(_02404_),
    .A1(_08709_),
    .A2(net469));
 sg13g2_mux2_1 _25738_ (.A0(_04741_),
    .A1(\cpu.icache.r_tag[7][9] ),
    .S(_06740_),
    .X(_02405_));
 sg13g2_mux2_1 _25739_ (.A0(_04774_),
    .A1(\cpu.icache.r_tag[7][10] ),
    .S(net470),
    .X(_02406_));
 sg13g2_nand2_1 _25740_ (.Y(_06753_),
    .A(\cpu.icache.r_tag[7][11] ),
    .B(_06743_));
 sg13g2_o21ai_1 _25741_ (.B1(_06753_),
    .Y(_02407_),
    .A1(net1077),
    .A2(net470));
 sg13g2_nand2_1 _25742_ (.Y(_06754_),
    .A(\cpu.icache.r_tag[7][12] ),
    .B(_06739_));
 sg13g2_o21ai_1 _25743_ (.B1(_06754_),
    .Y(_02408_),
    .A1(_08565_),
    .A2(net470));
 sg13g2_nand2_1 _25744_ (.Y(_06755_),
    .A(\cpu.icache.r_tag[7][13] ),
    .B(_06739_));
 sg13g2_o21ai_1 _25745_ (.B1(_06755_),
    .Y(_02409_),
    .A1(net431),
    .A2(net470));
 sg13g2_nand2_1 _25746_ (.Y(_06756_),
    .A(\cpu.icache.r_tag[7][14] ),
    .B(_06739_));
 sg13g2_o21ai_1 _25747_ (.B1(_06756_),
    .Y(_02410_),
    .A1(_08848_),
    .A2(net470));
 sg13g2_buf_1 _25748_ (.A(_09953_),
    .X(_06757_));
 sg13g2_nand2_1 _25749_ (.Y(_06758_),
    .A(net103),
    .B(net405));
 sg13g2_buf_1 _25750_ (.A(_06758_),
    .X(_06759_));
 sg13g2_buf_1 _25751_ (.A(_06759_),
    .X(_06760_));
 sg13g2_mux2_1 _25752_ (.A0(net913),
    .A1(\cpu.intr.r_clock_cmp[0] ),
    .S(_06760_),
    .X(_02420_));
 sg13g2_buf_1 _25753_ (.A(_06759_),
    .X(_06761_));
 sg13g2_nand2_1 _25754_ (.Y(_06762_),
    .A(\cpu.intr.r_clock_cmp[10] ),
    .B(net71));
 sg13g2_o21ai_1 _25755_ (.B1(_06762_),
    .Y(_02421_),
    .A1(_12066_),
    .A2(net72));
 sg13g2_mux2_1 _25756_ (.A0(_10162_),
    .A1(\cpu.intr.r_clock_cmp[11] ),
    .S(net71),
    .X(_02422_));
 sg13g2_nand2_1 _25757_ (.Y(_06763_),
    .A(\cpu.intr.r_clock_cmp[12] ),
    .B(net71));
 sg13g2_o21ai_1 _25758_ (.B1(_06763_),
    .Y(_02423_),
    .A1(_12093_),
    .A2(net72));
 sg13g2_nand2_1 _25759_ (.Y(_06764_),
    .A(\cpu.intr.r_clock_cmp[13] ),
    .B(net71));
 sg13g2_o21ai_1 _25760_ (.B1(_06764_),
    .Y(_02424_),
    .A1(_12101_),
    .A2(net72));
 sg13g2_nand2_1 _25761_ (.Y(_06765_),
    .A(\cpu.intr.r_clock_cmp[14] ),
    .B(net71));
 sg13g2_o21ai_1 _25762_ (.B1(_06765_),
    .Y(_02425_),
    .A1(_12107_),
    .A2(net72));
 sg13g2_nand2_1 _25763_ (.Y(_06766_),
    .A(\cpu.intr.r_clock_cmp[15] ),
    .B(_06759_));
 sg13g2_o21ai_1 _25764_ (.B1(_06766_),
    .Y(_02426_),
    .A1(_12113_),
    .A2(_06760_));
 sg13g2_nand2_1 _25765_ (.Y(_06767_),
    .A(net103),
    .B(net407));
 sg13g2_buf_1 _25766_ (.A(_06767_),
    .X(_06768_));
 sg13g2_buf_1 _25767_ (.A(_06768_),
    .X(_06769_));
 sg13g2_mux2_1 _25768_ (.A0(net913),
    .A1(\cpu.intr.r_clock_cmp[16] ),
    .S(net70),
    .X(_02427_));
 sg13g2_buf_1 _25769_ (.A(_06768_),
    .X(_06770_));
 sg13g2_mux2_1 _25770_ (.A0(net853),
    .A1(\cpu.intr.r_clock_cmp[17] ),
    .S(net69),
    .X(_02428_));
 sg13g2_mux2_1 _25771_ (.A0(net845),
    .A1(\cpu.intr.r_clock_cmp[18] ),
    .S(_06770_),
    .X(_02429_));
 sg13g2_mux2_1 _25772_ (.A0(net964),
    .A1(\cpu.intr.r_clock_cmp[19] ),
    .S(net69),
    .X(_02430_));
 sg13g2_mux2_1 _25773_ (.A0(net853),
    .A1(\cpu.intr.r_clock_cmp[1] ),
    .S(_06761_),
    .X(_02431_));
 sg13g2_nand2_1 _25774_ (.Y(_06771_),
    .A(\cpu.intr.r_clock_cmp[20] ),
    .B(_06770_));
 sg13g2_o21ai_1 _25775_ (.B1(_06771_),
    .Y(_02432_),
    .A1(net883),
    .A2(_06769_));
 sg13g2_nand2_1 _25776_ (.Y(_06772_),
    .A(\cpu.intr.r_clock_cmp[21] ),
    .B(net69));
 sg13g2_o21ai_1 _25777_ (.B1(_06772_),
    .Y(_02433_),
    .A1(net882),
    .A2(net70));
 sg13g2_nand2_1 _25778_ (.Y(_06773_),
    .A(\cpu.intr.r_clock_cmp[22] ),
    .B(net69));
 sg13g2_o21ai_1 _25779_ (.B1(_06773_),
    .Y(_02434_),
    .A1(net881),
    .A2(_06769_));
 sg13g2_mux2_1 _25780_ (.A0(net1056),
    .A1(\cpu.intr.r_clock_cmp[23] ),
    .S(net69),
    .X(_02435_));
 sg13g2_mux2_1 _25781_ (.A0(_10146_),
    .A1(\cpu.intr.r_clock_cmp[24] ),
    .S(net69),
    .X(_02436_));
 sg13g2_nand2_1 _25782_ (.Y(_06774_),
    .A(\cpu.intr.r_clock_cmp[25] ),
    .B(net69));
 sg13g2_o21ai_1 _25783_ (.B1(_06774_),
    .Y(_02437_),
    .A1(_12170_),
    .A2(net70));
 sg13g2_nand2_1 _25784_ (.Y(_06775_),
    .A(\cpu.intr.r_clock_cmp[26] ),
    .B(_06768_));
 sg13g2_o21ai_1 _25785_ (.B1(_06775_),
    .Y(_02438_),
    .A1(_12066_),
    .A2(net70));
 sg13g2_mux2_1 _25786_ (.A0(_10162_),
    .A1(\cpu.intr.r_clock_cmp[27] ),
    .S(net69),
    .X(_02439_));
 sg13g2_nand2_1 _25787_ (.Y(_06776_),
    .A(\cpu.intr.r_clock_cmp[28] ),
    .B(_06768_));
 sg13g2_o21ai_1 _25788_ (.B1(_06776_),
    .Y(_02440_),
    .A1(_12093_),
    .A2(net70));
 sg13g2_nand2_1 _25789_ (.Y(_06777_),
    .A(\cpu.intr.r_clock_cmp[29] ),
    .B(_06768_));
 sg13g2_o21ai_1 _25790_ (.B1(_06777_),
    .Y(_02441_),
    .A1(_12101_),
    .A2(net70));
 sg13g2_mux2_1 _25791_ (.A0(net845),
    .A1(\cpu.intr.r_clock_cmp[2] ),
    .S(net71),
    .X(_02442_));
 sg13g2_nand2_1 _25792_ (.Y(_06778_),
    .A(\cpu.intr.r_clock_cmp[30] ),
    .B(_06768_));
 sg13g2_o21ai_1 _25793_ (.B1(_06778_),
    .Y(_02443_),
    .A1(_12107_),
    .A2(net70));
 sg13g2_nand2_1 _25794_ (.Y(_06779_),
    .A(\cpu.intr.r_clock_cmp[31] ),
    .B(_06768_));
 sg13g2_o21ai_1 _25795_ (.B1(_06779_),
    .Y(_02444_),
    .A1(_12113_),
    .A2(net70));
 sg13g2_mux2_1 _25796_ (.A0(net964),
    .A1(\cpu.intr.r_clock_cmp[3] ),
    .S(_06761_),
    .X(_02445_));
 sg13g2_nand2_1 _25797_ (.Y(_06780_),
    .A(\cpu.intr.r_clock_cmp[4] ),
    .B(_06759_));
 sg13g2_o21ai_1 _25798_ (.B1(_06780_),
    .Y(_02446_),
    .A1(net883),
    .A2(net72));
 sg13g2_nand2_1 _25799_ (.Y(_06781_),
    .A(\cpu.intr.r_clock_cmp[5] ),
    .B(_06759_));
 sg13g2_o21ai_1 _25800_ (.B1(_06781_),
    .Y(_02447_),
    .A1(net882),
    .A2(net72));
 sg13g2_nand2_1 _25801_ (.Y(_06782_),
    .A(\cpu.intr.r_clock_cmp[6] ),
    .B(_06759_));
 sg13g2_o21ai_1 _25802_ (.B1(_06782_),
    .Y(_02448_),
    .A1(net881),
    .A2(net72));
 sg13g2_mux2_1 _25803_ (.A0(net1056),
    .A1(\cpu.intr.r_clock_cmp[7] ),
    .S(net71),
    .X(_02449_));
 sg13g2_mux2_1 _25804_ (.A0(_10146_),
    .A1(\cpu.intr.r_clock_cmp[8] ),
    .S(net71),
    .X(_02450_));
 sg13g2_nand2_1 _25805_ (.Y(_06783_),
    .A(\cpu.intr.r_clock_cmp[9] ),
    .B(_06759_));
 sg13g2_o21ai_1 _25806_ (.B1(_06783_),
    .Y(_02451_),
    .A1(_12170_),
    .A2(net72));
 sg13g2_nand2_1 _25807_ (.Y(_06784_),
    .A(net103),
    .B(net449));
 sg13g2_buf_1 _25808_ (.A(_06784_),
    .X(_06785_));
 sg13g2_buf_1 _25809_ (.A(_06785_),
    .X(_06786_));
 sg13g2_mux2_1 _25810_ (.A0(net913),
    .A1(\cpu.intr.r_timer_reload[0] ),
    .S(net68),
    .X(_02475_));
 sg13g2_buf_1 _25811_ (.A(_06785_),
    .X(_06787_));
 sg13g2_nand2_1 _25812_ (.Y(_06788_),
    .A(\cpu.intr.r_timer_reload[10] ),
    .B(net67));
 sg13g2_o21ai_1 _25813_ (.B1(_06788_),
    .Y(_02476_),
    .A1(_12066_),
    .A2(net68));
 sg13g2_mux2_1 _25814_ (.A0(_10162_),
    .A1(\cpu.intr.r_timer_reload[11] ),
    .S(net67),
    .X(_02477_));
 sg13g2_nand2_1 _25815_ (.Y(_06789_),
    .A(\cpu.intr.r_timer_reload[12] ),
    .B(net67));
 sg13g2_o21ai_1 _25816_ (.B1(_06789_),
    .Y(_02478_),
    .A1(_12093_),
    .A2(net68));
 sg13g2_nand2_1 _25817_ (.Y(_06790_),
    .A(\cpu.intr.r_timer_reload[13] ),
    .B(net67));
 sg13g2_o21ai_1 _25818_ (.B1(_06790_),
    .Y(_02479_),
    .A1(_12101_),
    .A2(net68));
 sg13g2_nand2_1 _25819_ (.Y(_06791_),
    .A(\cpu.intr.r_timer_reload[14] ),
    .B(net67));
 sg13g2_o21ai_1 _25820_ (.B1(_06791_),
    .Y(_02480_),
    .A1(_12107_),
    .A2(net68));
 sg13g2_nand2_1 _25821_ (.Y(_06792_),
    .A(\cpu.intr.r_timer_reload[15] ),
    .B(_06785_));
 sg13g2_o21ai_1 _25822_ (.B1(_06792_),
    .Y(_02481_),
    .A1(_12113_),
    .A2(_06786_));
 sg13g2_mux2_1 _25823_ (.A0(\cpu.intr.r_timer_reload[16] ),
    .A1(net911),
    .S(_10046_),
    .X(_02482_));
 sg13g2_inv_1 _25824_ (.Y(_06793_),
    .A(\cpu.intr.r_timer_reload[17] ));
 sg13g2_o21ai_1 _25825_ (.B1(_10052_),
    .Y(_02483_),
    .A1(_06793_),
    .A2(net110));
 sg13g2_inv_1 _25826_ (.Y(_06794_),
    .A(\cpu.intr.r_timer_reload[18] ));
 sg13g2_o21ai_1 _25827_ (.B1(_10057_),
    .Y(_02484_),
    .A1(_06794_),
    .A2(net110));
 sg13g2_inv_1 _25828_ (.Y(_06795_),
    .A(\cpu.intr.r_timer_reload[19] ));
 sg13g2_o21ai_1 _25829_ (.B1(_10061_),
    .Y(_02485_),
    .A1(_06795_),
    .A2(_10047_));
 sg13g2_mux2_1 _25830_ (.A0(net853),
    .A1(\cpu.intr.r_timer_reload[1] ),
    .S(net67),
    .X(_02486_));
 sg13g2_o21ai_1 _25831_ (.B1(_10068_),
    .Y(_02487_),
    .A1(_10062_),
    .A2(net110));
 sg13g2_inv_1 _25832_ (.Y(_06796_),
    .A(\cpu.intr.r_timer_reload[21] ));
 sg13g2_o21ai_1 _25833_ (.B1(_10074_),
    .Y(_02488_),
    .A1(_06796_),
    .A2(net110));
 sg13g2_inv_1 _25834_ (.Y(_06797_),
    .A(\cpu.intr.r_timer_reload[22] ));
 sg13g2_o21ai_1 _25835_ (.B1(_10080_),
    .Y(_02489_),
    .A1(_06797_),
    .A2(net110));
 sg13g2_mux2_1 _25836_ (.A0(\cpu.intr.r_timer_reload[23] ),
    .A1(net1018),
    .S(net125),
    .X(_02490_));
 sg13g2_mux2_1 _25837_ (.A0(net845),
    .A1(\cpu.intr.r_timer_reload[2] ),
    .S(net67),
    .X(_02491_));
 sg13g2_mux2_1 _25838_ (.A0(net964),
    .A1(\cpu.intr.r_timer_reload[3] ),
    .S(_06787_),
    .X(_02492_));
 sg13g2_nand2_1 _25839_ (.Y(_06798_),
    .A(\cpu.intr.r_timer_reload[4] ),
    .B(_06785_));
 sg13g2_o21ai_1 _25840_ (.B1(_06798_),
    .Y(_02493_),
    .A1(net883),
    .A2(net68));
 sg13g2_nand2_1 _25841_ (.Y(_06799_),
    .A(\cpu.intr.r_timer_reload[5] ),
    .B(_06785_));
 sg13g2_o21ai_1 _25842_ (.B1(_06799_),
    .Y(_02494_),
    .A1(net882),
    .A2(_06786_));
 sg13g2_nand2_1 _25843_ (.Y(_06800_),
    .A(\cpu.intr.r_timer_reload[6] ),
    .B(_06785_));
 sg13g2_o21ai_1 _25844_ (.B1(_06800_),
    .Y(_02495_),
    .A1(net881),
    .A2(net68));
 sg13g2_mux2_1 _25845_ (.A0(net1056),
    .A1(\cpu.intr.r_timer_reload[7] ),
    .S(_06787_),
    .X(_02496_));
 sg13g2_mux2_1 _25846_ (.A0(_10146_),
    .A1(\cpu.intr.r_timer_reload[8] ),
    .S(net67),
    .X(_02497_));
 sg13g2_nand2_1 _25847_ (.Y(_06801_),
    .A(\cpu.intr.r_timer_reload[9] ),
    .B(_06785_));
 sg13g2_o21ai_1 _25848_ (.B1(_06801_),
    .Y(_02498_),
    .A1(_12170_),
    .A2(net68));
 sg13g2_inv_1 _25849_ (.Y(_06802_),
    .A(_09830_));
 sg13g2_a21oi_1 _25850_ (.A1(_09824_),
    .A2(_09869_),
    .Y(_06803_),
    .B1(_09360_));
 sg13g2_nor4_2 _25851_ (.A(_11916_),
    .B(_11938_),
    .C(_09886_),
    .Y(_06804_),
    .D(_11914_));
 sg13g2_nor3_1 _25852_ (.A(_11942_),
    .B(_11918_),
    .C(_11939_),
    .Y(_06805_));
 sg13g2_nand2_1 _25853_ (.Y(_06806_),
    .A(_06804_),
    .B(_06805_));
 sg13g2_nor4_1 _25854_ (.A(_09839_),
    .B(_09827_),
    .C(_06803_),
    .D(_06806_),
    .Y(_06807_));
 sg13g2_buf_1 _25855_ (.A(_06807_),
    .X(_06808_));
 sg13g2_and2_1 _25856_ (.A(\cpu.qspi.r_read_delay[1][0] ),
    .B(net81),
    .X(_06809_));
 sg13g2_a221oi_1 _25857_ (.B2(\cpu.qspi.r_read_delay[0][0] ),
    .C1(_06809_),
    .B1(_09866_),
    .A1(\cpu.qspi.r_read_delay[2][0] ),
    .Y(_06810_),
    .A2(net224));
 sg13g2_or4_1 _25858_ (.A(_09838_),
    .B(_09854_),
    .C(net1064),
    .D(_09841_),
    .X(_06811_));
 sg13g2_buf_1 _25859_ (.A(_06811_),
    .X(_06812_));
 sg13g2_a221oi_1 _25860_ (.B2(_06812_),
    .C1(_09846_),
    .B1(_00173_),
    .A1(_09873_),
    .Y(_06813_),
    .A2(_06802_));
 sg13g2_o21ai_1 _25861_ (.B1(_06813_),
    .Y(_06814_),
    .A1(_09889_),
    .A2(_06810_));
 sg13g2_nand2_1 _25862_ (.Y(_06815_),
    .A(_06808_),
    .B(_06814_));
 sg13g2_o21ai_1 _25863_ (.B1(_06815_),
    .Y(_02499_),
    .A1(_06802_),
    .A2(net27));
 sg13g2_inv_1 _25864_ (.Y(_06816_),
    .A(_09831_));
 sg13g2_and2_1 _25865_ (.A(\cpu.qspi.r_read_delay[1][1] ),
    .B(net81),
    .X(_06817_));
 sg13g2_a221oi_1 _25866_ (.B2(\cpu.qspi.r_read_delay[0][1] ),
    .C1(_06817_),
    .B1(_09866_),
    .A1(\cpu.qspi.r_read_delay[2][1] ),
    .Y(_06818_),
    .A2(net224));
 sg13g2_nor2_1 _25867_ (.A(_09873_),
    .B(_06812_),
    .Y(_06819_));
 sg13g2_xor2_1 _25868_ (.B(_09831_),
    .A(_09830_),
    .X(_06820_));
 sg13g2_nor2_1 _25869_ (.A(_06819_),
    .B(_06820_),
    .Y(_06821_));
 sg13g2_a21oi_1 _25870_ (.A1(_09889_),
    .A2(_06819_),
    .Y(_06822_),
    .B1(_06821_));
 sg13g2_o21ai_1 _25871_ (.B1(_06822_),
    .Y(_06823_),
    .A1(_09889_),
    .A2(_06818_));
 sg13g2_o21ai_1 _25872_ (.B1(net27),
    .Y(_06824_),
    .A1(_09846_),
    .A2(_06823_));
 sg13g2_o21ai_1 _25873_ (.B1(_06824_),
    .Y(_02500_),
    .A1(_06816_),
    .A2(_06808_));
 sg13g2_nor2_1 _25874_ (.A(_09830_),
    .B(_09831_),
    .Y(_06825_));
 sg13g2_xor2_1 _25875_ (.B(_06825_),
    .A(_00174_),
    .X(_06826_));
 sg13g2_nor4_2 _25876_ (.A(_09838_),
    .B(_09854_),
    .C(net1064),
    .Y(_06827_),
    .D(_09841_));
 sg13g2_o21ai_1 _25877_ (.B1(_09890_),
    .Y(_06828_),
    .A1(_09873_),
    .A2(_06827_));
 sg13g2_a22oi_1 _25878_ (.Y(_06829_),
    .B1(_06826_),
    .B2(_06828_),
    .A2(_06819_),
    .A1(_09888_));
 sg13g2_a22oi_1 _25879_ (.Y(_06830_),
    .B1(net81),
    .B2(\cpu.qspi.r_read_delay[1][2] ),
    .A2(net224),
    .A1(\cpu.qspi.r_read_delay[2][2] ));
 sg13g2_nand2_1 _25880_ (.Y(_06831_),
    .A(\cpu.qspi.r_read_delay[0][2] ),
    .B(_09866_));
 sg13g2_a21oi_1 _25881_ (.A1(_06830_),
    .A2(_06831_),
    .Y(_06832_),
    .B1(_09889_));
 sg13g2_nor3_1 _25882_ (.A(_09846_),
    .B(_06829_),
    .C(_06832_),
    .Y(_06833_));
 sg13g2_nor2_1 _25883_ (.A(_09832_),
    .B(net27),
    .Y(_06834_));
 sg13g2_a21oi_1 _25884_ (.A1(net27),
    .A2(_06833_),
    .Y(_02501_),
    .B1(_06834_));
 sg13g2_a21oi_1 _25885_ (.A1(_09890_),
    .A2(_06827_),
    .Y(_06835_),
    .B1(_09833_));
 sg13g2_nand2b_1 _25886_ (.Y(_06836_),
    .B(net27),
    .A_N(_06835_));
 sg13g2_nand2_1 _25887_ (.Y(_06837_),
    .A(_09890_),
    .B(_06827_));
 sg13g2_inv_1 _25888_ (.Y(_06838_),
    .A(\cpu.qspi.r_read_delay[0][3] ));
 sg13g2_or2_1 _25889_ (.X(_06839_),
    .B(_09863_),
    .A(net224));
 sg13g2_a22oi_1 _25890_ (.Y(_06840_),
    .B1(net81),
    .B2(\cpu.qspi.r_read_delay[1][3] ),
    .A2(net224),
    .A1(\cpu.qspi.r_read_delay[2][3] ));
 sg13g2_o21ai_1 _25891_ (.B1(_06840_),
    .Y(_06841_),
    .A1(_06838_),
    .A2(_06839_));
 sg13g2_a22oi_1 _25892_ (.Y(_06842_),
    .B1(_06841_),
    .B2(_09888_),
    .A2(_06837_),
    .A1(_09835_));
 sg13g2_nor2b_1 _25893_ (.A(_06842_),
    .B_N(net27),
    .Y(_06843_));
 sg13g2_a21o_1 _25894_ (.A2(_06836_),
    .A1(\cpu.qspi.r_count[3] ),
    .B1(_06843_),
    .X(_02502_));
 sg13g2_and2_1 _25895_ (.A(_09835_),
    .B(_06812_),
    .X(_06844_));
 sg13g2_nor3_1 _25896_ (.A(_09829_),
    .B(_09835_),
    .C(_06819_),
    .Y(_06845_));
 sg13g2_a21oi_1 _25897_ (.A1(_09829_),
    .A2(_06844_),
    .Y(_06846_),
    .B1(_06845_));
 sg13g2_nor2_1 _25898_ (.A(\cpu.qspi.r_count[4] ),
    .B(net27),
    .Y(_06847_));
 sg13g2_a21oi_1 _25899_ (.A1(net27),
    .A2(_06846_),
    .Y(_02503_),
    .B1(_06847_));
 sg13g2_nor2_1 _25900_ (.A(_09220_),
    .B(_09246_),
    .Y(_06848_));
 sg13g2_and2_1 _25901_ (.A(_09949_),
    .B(_06848_),
    .X(_06849_));
 sg13g2_buf_1 _25902_ (.A(_06849_),
    .X(_06850_));
 sg13g2_and2_1 _25903_ (.A(_09235_),
    .B(_06850_),
    .X(_06851_));
 sg13g2_buf_1 _25904_ (.A(_06851_),
    .X(_06852_));
 sg13g2_nand2_1 _25905_ (.Y(_06853_),
    .A(net874),
    .B(_06852_));
 sg13g2_nand2_1 _25906_ (.Y(_06854_),
    .A(_09235_),
    .B(_06850_));
 sg13g2_buf_1 _25907_ (.A(_06854_),
    .X(_06855_));
 sg13g2_nand2_1 _25908_ (.Y(_06856_),
    .A(\cpu.qspi.r_read_delay[0][0] ),
    .B(_06855_));
 sg13g2_a21oi_1 _25909_ (.A1(_06853_),
    .A2(_06856_),
    .Y(_02514_),
    .B1(net687));
 sg13g2_nand2_1 _25910_ (.Y(_06857_),
    .A(net1055),
    .B(_06852_));
 sg13g2_nand2_1 _25911_ (.Y(_06858_),
    .A(\cpu.qspi.r_read_delay[0][1] ),
    .B(_06855_));
 sg13g2_a21oi_1 _25912_ (.A1(_06857_),
    .A2(_06858_),
    .Y(_02515_),
    .B1(net687));
 sg13g2_nand2_1 _25913_ (.Y(_06859_),
    .A(net910),
    .B(_06852_));
 sg13g2_nand2_1 _25914_ (.Y(_06860_),
    .A(\cpu.qspi.r_read_delay[0][2] ),
    .B(_06855_));
 sg13g2_nand3_1 _25915_ (.B(_06859_),
    .C(_06860_),
    .A(net634),
    .Y(_02516_));
 sg13g2_buf_1 _25916_ (.A(net1128),
    .X(_06861_));
 sg13g2_nand2_1 _25917_ (.Y(_06862_),
    .A(net954),
    .B(_06852_));
 sg13g2_nand2_1 _25918_ (.Y(_06863_),
    .A(\cpu.qspi.r_read_delay[0][3] ),
    .B(_06855_));
 sg13g2_a21oi_1 _25919_ (.A1(_06862_),
    .A2(_06863_),
    .Y(_02517_),
    .B1(net687));
 sg13g2_nand2_1 _25920_ (.Y(_06864_),
    .A(_12124_),
    .B(net540));
 sg13g2_nand2_1 _25921_ (.Y(_06865_),
    .A(_09949_),
    .B(_06848_));
 sg13g2_nor2_1 _25922_ (.A(_06864_),
    .B(_06865_),
    .Y(_06866_));
 sg13g2_nand2_1 _25923_ (.Y(_06867_),
    .A(_02704_),
    .B(_06866_));
 sg13g2_nand2_1 _25924_ (.Y(_06868_),
    .A(_10112_),
    .B(_06850_));
 sg13g2_buf_1 _25925_ (.A(_06868_),
    .X(_06869_));
 sg13g2_nand2_1 _25926_ (.Y(_06870_),
    .A(\cpu.qspi.r_read_delay[1][0] ),
    .B(_06869_));
 sg13g2_a21oi_1 _25927_ (.A1(_06867_),
    .A2(_06870_),
    .Y(_02518_),
    .B1(net687));
 sg13g2_nand2_1 _25928_ (.Y(_06871_),
    .A(_10101_),
    .B(_06866_));
 sg13g2_nand2_1 _25929_ (.Y(_06872_),
    .A(\cpu.qspi.r_read_delay[1][1] ),
    .B(_06869_));
 sg13g2_a21oi_1 _25930_ (.A1(_06871_),
    .A2(_06872_),
    .Y(_02519_),
    .B1(net687));
 sg13g2_nand2_1 _25931_ (.Y(_06873_),
    .A(net910),
    .B(_06866_));
 sg13g2_nand2_1 _25932_ (.Y(_06874_),
    .A(\cpu.qspi.r_read_delay[1][2] ),
    .B(_06869_));
 sg13g2_nand3_1 _25933_ (.B(_06873_),
    .C(_06874_),
    .A(net634),
    .Y(_02520_));
 sg13g2_nand2_1 _25934_ (.Y(_06875_),
    .A(net954),
    .B(_06866_));
 sg13g2_nand2_1 _25935_ (.Y(_06876_),
    .A(\cpu.qspi.r_read_delay[1][3] ),
    .B(_06869_));
 sg13g2_a21oi_1 _25936_ (.A1(_06875_),
    .A2(_06876_),
    .Y(_02521_),
    .B1(net687));
 sg13g2_nor2_1 _25937_ (.A(_04886_),
    .B(_06865_),
    .Y(_06877_));
 sg13g2_buf_1 _25938_ (.A(_06877_),
    .X(_06878_));
 sg13g2_nand2_1 _25939_ (.Y(_06879_),
    .A(net874),
    .B(_06878_));
 sg13g2_nand2_1 _25940_ (.Y(_06880_),
    .A(_04895_),
    .B(_06850_));
 sg13g2_buf_1 _25941_ (.A(_06880_),
    .X(_06881_));
 sg13g2_nand2_1 _25942_ (.Y(_06882_),
    .A(\cpu.qspi.r_read_delay[2][0] ),
    .B(_06881_));
 sg13g2_a21oi_1 _25943_ (.A1(_06879_),
    .A2(_06882_),
    .Y(_02522_),
    .B1(net687));
 sg13g2_nand2_1 _25944_ (.Y(_06883_),
    .A(net1055),
    .B(_06878_));
 sg13g2_nand2_1 _25945_ (.Y(_06884_),
    .A(\cpu.qspi.r_read_delay[2][1] ),
    .B(_06881_));
 sg13g2_buf_2 _25946_ (.A(_09330_),
    .X(_06885_));
 sg13g2_a21oi_1 _25947_ (.A1(_06883_),
    .A2(_06884_),
    .Y(_02523_),
    .B1(net656));
 sg13g2_nand2_1 _25948_ (.Y(_06886_),
    .A(_10107_),
    .B(_06878_));
 sg13g2_nand2_1 _25949_ (.Y(_06887_),
    .A(\cpu.qspi.r_read_delay[2][2] ),
    .B(_06881_));
 sg13g2_nand3_1 _25950_ (.B(_06886_),
    .C(_06887_),
    .A(net634),
    .Y(_02524_));
 sg13g2_nand2_1 _25951_ (.Y(_06888_),
    .A(net954),
    .B(_06878_));
 sg13g2_nand2_1 _25952_ (.Y(_06889_),
    .A(\cpu.qspi.r_read_delay[2][3] ),
    .B(_06881_));
 sg13g2_a21oi_1 _25953_ (.A1(_06888_),
    .A2(_06889_),
    .Y(_02525_),
    .B1(net656));
 sg13g2_a22oi_1 _25954_ (.Y(_06890_),
    .B1(net81),
    .B2(\cpu.qspi.r_mask[1] ),
    .A2(net224),
    .A1(\cpu.qspi.r_mask[2] ));
 sg13g2_nand2_1 _25955_ (.Y(_06891_),
    .A(\cpu.qspi.r_mask[0] ),
    .B(_09866_));
 sg13g2_nand3_1 _25956_ (.B(_06890_),
    .C(_06891_),
    .A(_11916_),
    .Y(_06892_));
 sg13g2_nor2_1 _25957_ (.A(_09873_),
    .B(_09825_),
    .Y(_06893_));
 sg13g2_nor3_2 _25958_ (.A(_09838_),
    .B(_09839_),
    .C(_09827_),
    .Y(_06894_));
 sg13g2_nand4_1 _25959_ (.B(_06892_),
    .C(_06893_),
    .A(_09889_),
    .Y(_06895_),
    .D(_06894_));
 sg13g2_buf_2 _25960_ (.A(_06895_),
    .X(_06896_));
 sg13g2_buf_1 _25961_ (.A(_08346_),
    .X(_06897_));
 sg13g2_buf_1 _25962_ (.A(net829),
    .X(_06898_));
 sg13g2_buf_1 _25963_ (.A(net829),
    .X(_06899_));
 sg13g2_buf_1 _25964_ (.A(_09819_),
    .X(_06900_));
 sg13g2_mux2_1 _25965_ (.A0(_09800_),
    .A1(net418),
    .S(net96),
    .X(_06901_));
 sg13g2_nand2_1 _25966_ (.Y(_06902_),
    .A(_06899_),
    .B(_06901_));
 sg13g2_o21ai_1 _25967_ (.B1(_06902_),
    .Y(_06903_),
    .A1(net728),
    .A2(_08758_));
 sg13g2_buf_1 _25968_ (.A(_09819_),
    .X(_06904_));
 sg13g2_and2_1 _25969_ (.A(_09397_),
    .B(net95),
    .X(_06905_));
 sg13g2_nor2_1 _25970_ (.A(_09434_),
    .B(net95),
    .Y(_06906_));
 sg13g2_o21ai_1 _25971_ (.B1(net727),
    .Y(_06907_),
    .A1(_06905_),
    .A2(_06906_));
 sg13g2_o21ai_1 _25972_ (.B1(_06907_),
    .Y(_06908_),
    .A1(net728),
    .A2(_08565_));
 sg13g2_nor2_1 _25973_ (.A(_09627_),
    .B(_09819_),
    .Y(_06909_));
 sg13g2_a21oi_1 _25974_ (.A1(_00219_),
    .A2(net96),
    .Y(_06910_),
    .B1(_06909_));
 sg13g2_nand2_1 _25975_ (.Y(_06911_),
    .A(net829),
    .B(_06910_));
 sg13g2_o21ai_1 _25976_ (.B1(_06911_),
    .Y(_06912_),
    .A1(net727),
    .A2(_10487_));
 sg13g2_nand2b_1 _25977_ (.Y(_06913_),
    .B(_09886_),
    .A_N(net111));
 sg13g2_mux2_1 _25978_ (.A0(_05226_),
    .A1(_04873_),
    .S(_12026_),
    .X(_06914_));
 sg13g2_nand2_1 _25979_ (.Y(_06915_),
    .A(_12026_),
    .B(_04866_));
 sg13g2_o21ai_1 _25980_ (.B1(_06915_),
    .Y(_06916_),
    .A1(_12027_),
    .A2(_05219_));
 sg13g2_a22oi_1 _25981_ (.Y(_06917_),
    .B1(_06916_),
    .B2(net1027),
    .A2(_06914_),
    .A1(net1001));
 sg13g2_inv_1 _25982_ (.Y(_06918_),
    .A(_12030_));
 sg13g2_nand2_1 _25983_ (.Y(_06919_),
    .A(_12047_),
    .B(_04843_));
 sg13g2_o21ai_1 _25984_ (.B1(_06919_),
    .Y(_06920_),
    .A1(_06918_),
    .A2(_04851_));
 sg13g2_nor2b_1 _25985_ (.A(net1028),
    .B_N(_12047_),
    .Y(_06921_));
 sg13g2_a221oi_1 _25986_ (.B2(_05582_),
    .C1(_12025_),
    .B1(_06921_),
    .A1(_12027_),
    .Y(_06922_),
    .A2(_06920_));
 sg13g2_a21oi_1 _25987_ (.A1(_12025_),
    .A2(_06917_),
    .Y(_06923_),
    .B1(_06922_));
 sg13g2_nor2b_1 _25988_ (.A(_12139_),
    .B_N(_12030_),
    .Y(_06924_));
 sg13g2_nor2_1 _25989_ (.A(_12047_),
    .B(_06924_),
    .Y(_06925_));
 sg13g2_buf_1 _25990_ (.A(_06925_),
    .X(_06926_));
 sg13g2_and2_1 _25991_ (.A(_05590_),
    .B(_06926_),
    .X(_06927_));
 sg13g2_o21ai_1 _25992_ (.B1(_09841_),
    .Y(_06928_),
    .A1(_06923_),
    .A2(_06927_));
 sg13g2_nand2_1 _25993_ (.Y(_06929_),
    .A(_11912_),
    .B(_09848_));
 sg13g2_nand3b_1 _25994_ (.B(_11919_),
    .C(_06805_),
    .Y(_06930_),
    .A_N(_09854_));
 sg13g2_buf_1 _25995_ (.A(_06930_),
    .X(_06931_));
 sg13g2_nor2b_1 _25996_ (.A(_09849_),
    .B_N(_06804_),
    .Y(_06932_));
 sg13g2_inv_1 _25997_ (.Y(_06933_),
    .A(_06932_));
 sg13g2_nor3_2 _25998_ (.A(_06929_),
    .B(_06931_),
    .C(_06933_),
    .Y(_06934_));
 sg13g2_nor2_1 _25999_ (.A(_11916_),
    .B(_06934_),
    .Y(_06935_));
 sg13g2_buf_1 _26000_ (.A(\cpu.qspi.r_state[0] ),
    .X(_06936_));
 sg13g2_buf_1 _26001_ (.A(_08345_),
    .X(_06937_));
 sg13g2_nand2_1 _26002_ (.Y(_06938_),
    .A(net1141),
    .B(_08345_));
 sg13g2_o21ai_1 _26003_ (.B1(_06938_),
    .Y(_06939_),
    .A1(net953),
    .A2(_09810_));
 sg13g2_a22oi_1 _26004_ (.Y(_06940_),
    .B1(_06939_),
    .B2(_11939_),
    .A2(_06936_),
    .A1(_09875_));
 sg13g2_nand4_1 _26005_ (.B(_06928_),
    .C(_06935_),
    .A(_06913_),
    .Y(_06941_),
    .D(_06940_));
 sg13g2_a21o_1 _26006_ (.A2(_06912_),
    .A1(_11938_),
    .B1(_06941_),
    .X(_06942_));
 sg13g2_a221oi_1 _26007_ (.B2(_11918_),
    .C1(_06942_),
    .B1(_06908_),
    .A1(_11942_),
    .Y(_06943_),
    .A2(_06903_));
 sg13g2_nand2_1 _26008_ (.Y(_06944_),
    .A(_09849_),
    .B(_09828_));
 sg13g2_nand3_1 _26009_ (.B(_09831_),
    .C(_06944_),
    .A(_06802_),
    .Y(_06945_));
 sg13g2_o21ai_1 _26010_ (.B1(_06945_),
    .Y(_06946_),
    .A1(_06802_),
    .A2(_06944_));
 sg13g2_nor2_1 _26011_ (.A(_09832_),
    .B(_06946_),
    .Y(_06947_));
 sg13g2_nand3b_1 _26012_ (.B(_00173_),
    .C(_06944_),
    .Y(_06948_),
    .A_N(_09831_));
 sg13g2_nor2b_1 _26013_ (.A(net1064),
    .B_N(_09845_),
    .Y(_06949_));
 sg13g2_o21ai_1 _26014_ (.B1(_09832_),
    .Y(_06950_),
    .A1(_06948_),
    .A2(_06949_));
 sg13g2_nor3_1 _26015_ (.A(_09850_),
    .B(_09830_),
    .C(_06950_),
    .Y(_06951_));
 sg13g2_nor2_1 _26016_ (.A(_06947_),
    .B(_06951_),
    .Y(_06952_));
 sg13g2_o21ai_1 _26017_ (.B1(_06947_),
    .Y(_06953_),
    .A1(_09850_),
    .A2(_09831_));
 sg13g2_o21ai_1 _26018_ (.B1(_06953_),
    .Y(_06954_),
    .A1(_09831_),
    .A2(_06950_));
 sg13g2_inv_1 _26019_ (.Y(_06955_),
    .A(_06954_));
 sg13g2_o21ai_1 _26020_ (.B1(_06955_),
    .Y(_06956_),
    .A1(net111),
    .A2(_06952_));
 sg13g2_o21ai_1 _26021_ (.B1(_06956_),
    .Y(_06957_),
    .A1(_09854_),
    .A2(net1064));
 sg13g2_xnor2_1 _26022_ (.Y(_06958_),
    .A(net111),
    .B(_09869_));
 sg13g2_a221oi_1 _26023_ (.B2(_06934_),
    .C1(_06896_),
    .B1(_06958_),
    .A1(_06943_),
    .Y(_06959_),
    .A2(_06957_));
 sg13g2_a21o_1 _26024_ (.A2(_06896_),
    .A1(net11),
    .B1(_06959_),
    .X(_02530_));
 sg13g2_mux2_1 _26025_ (.A0(_09470_),
    .A1(_09451_),
    .S(net95),
    .X(_06960_));
 sg13g2_nand2_1 _26026_ (.Y(_06961_),
    .A(net728),
    .B(_06960_));
 sg13g2_o21ai_1 _26027_ (.B1(_06961_),
    .Y(_06962_),
    .A1(net728),
    .A2(_08497_));
 sg13g2_inv_1 _26028_ (.Y(_06963_),
    .A(_05653_));
 sg13g2_a22oi_1 _26029_ (.Y(_06964_),
    .B1(_05250_),
    .B2(net1001),
    .A2(_05257_),
    .A1(net1027));
 sg13g2_a22oi_1 _26030_ (.Y(_06965_),
    .B1(_05329_),
    .B2(net1001),
    .A2(_05322_),
    .A1(net1027));
 sg13g2_a22oi_1 _26031_ (.Y(_06966_),
    .B1(_05347_),
    .B2(net1001),
    .A2(_05339_),
    .A1(net1027));
 sg13g2_mux4_1 _26032_ (.S0(net1029),
    .A0(_06963_),
    .A1(_06964_),
    .A2(_06965_),
    .A3(_06966_),
    .S1(net1028),
    .X(_06967_));
 sg13g2_nand2b_1 _26033_ (.Y(_06968_),
    .B(_06926_),
    .A_N(_05662_));
 sg13g2_o21ai_1 _26034_ (.B1(_06968_),
    .Y(_06969_),
    .A1(_06926_),
    .A2(_06967_));
 sg13g2_a21oi_1 _26035_ (.A1(_09841_),
    .A2(_06969_),
    .Y(_06970_),
    .B1(_11916_));
 sg13g2_nand2_1 _26036_ (.Y(_06971_),
    .A(_06913_),
    .B(_06970_));
 sg13g2_a21oi_1 _26037_ (.A1(_11918_),
    .A2(_06962_),
    .Y(_06972_),
    .B1(_06971_));
 sg13g2_mux2_1 _26038_ (.A0(_09602_),
    .A1(_00221_),
    .S(net95),
    .X(_06973_));
 sg13g2_nand2_1 _26039_ (.Y(_06974_),
    .A(net953),
    .B(_10548_));
 sg13g2_o21ai_1 _26040_ (.B1(_06974_),
    .Y(_06975_),
    .A1(net953),
    .A2(_06973_));
 sg13g2_mux2_1 _26041_ (.A0(_09732_),
    .A1(net420),
    .S(net95),
    .X(_06976_));
 sg13g2_nand2_1 _26042_ (.Y(_06977_),
    .A(_06899_),
    .B(_06976_));
 sg13g2_o21ai_1 _26043_ (.B1(_06977_),
    .Y(_06978_),
    .A1(net728),
    .A2(_09091_));
 sg13g2_nand2_1 _26044_ (.Y(_06979_),
    .A(net953),
    .B(_10740_));
 sg13g2_nor2_1 _26045_ (.A(_09616_),
    .B(net95),
    .Y(_06980_));
 sg13g2_a21oi_1 _26046_ (.A1(_04980_),
    .A2(net95),
    .Y(_06981_),
    .B1(_06980_));
 sg13g2_nand2_1 _26047_ (.Y(_06982_),
    .A(net728),
    .B(_06981_));
 sg13g2_a21oi_1 _26048_ (.A1(_06979_),
    .A2(_06982_),
    .Y(_06983_),
    .B1(_11940_));
 sg13g2_a221oi_1 _26049_ (.B2(_11942_),
    .C1(_06983_),
    .B1(_06978_),
    .A1(_11938_),
    .Y(_06984_),
    .A2(_06975_));
 sg13g2_nand2b_1 _26050_ (.Y(_06985_),
    .B(_06934_),
    .A_N(_09869_));
 sg13g2_nand3_1 _26051_ (.B(_06984_),
    .C(_06985_),
    .A(_06972_),
    .Y(_06986_));
 sg13g2_mux2_1 _26052_ (.A0(_06986_),
    .A1(net12),
    .S(_06896_),
    .X(_02531_));
 sg13g2_mux2_1 _26053_ (.A0(_09584_),
    .A1(_09571_),
    .S(_06904_),
    .X(_06987_));
 sg13g2_nand2_1 _26054_ (.Y(_06988_),
    .A(net728),
    .B(_06987_));
 sg13g2_o21ai_1 _26055_ (.B1(_06988_),
    .Y(_06989_),
    .A1(net728),
    .A2(_10679_));
 sg13g2_mux2_1 _26056_ (.A0(_09557_),
    .A1(net366),
    .S(_09819_),
    .X(_06990_));
 sg13g2_nand2_1 _26057_ (.Y(_06991_),
    .A(net829),
    .B(_06990_));
 sg13g2_o21ai_1 _26058_ (.B1(_06991_),
    .Y(_06992_),
    .A1(net727),
    .A2(_08603_));
 sg13g2_mux2_1 _26059_ (.A0(_09664_),
    .A1(_09658_),
    .S(net96),
    .X(_06993_));
 sg13g2_nand2_1 _26060_ (.Y(_06994_),
    .A(net829),
    .B(_06993_));
 sg13g2_o21ai_1 _26061_ (.B1(_06994_),
    .Y(_06995_),
    .A1(net727),
    .A2(_08848_));
 sg13g2_a22oi_1 _26062_ (.Y(_06996_),
    .B1(_06995_),
    .B2(_11918_),
    .A2(_06992_),
    .A1(_11942_));
 sg13g2_mux2_1 _26063_ (.A0(_09569_),
    .A1(_00223_),
    .S(_06900_),
    .X(_06997_));
 sg13g2_nand2_1 _26064_ (.Y(_06998_),
    .A(net953),
    .B(_10389_));
 sg13g2_o21ai_1 _26065_ (.B1(_06998_),
    .Y(_06999_),
    .A1(_06937_),
    .A2(_06997_));
 sg13g2_nand2_1 _26066_ (.Y(_07000_),
    .A(_12118_),
    .B(_05404_));
 sg13g2_o21ai_1 _26067_ (.B1(_07000_),
    .Y(_07001_),
    .A1(_12087_),
    .A2(_05277_));
 sg13g2_and2_1 _26068_ (.A(_12031_),
    .B(_02941_),
    .X(_07002_));
 sg13g2_inv_1 _26069_ (.Y(_07003_),
    .A(_05145_));
 sg13g2_a221oi_1 _26070_ (.B2(_07003_),
    .C1(_06926_),
    .B1(_07002_),
    .A1(_02939_),
    .Y(_07004_),
    .A2(_07001_));
 sg13g2_nand2_1 _26071_ (.Y(_07005_),
    .A(net1001),
    .B(_05728_));
 sg13g2_nand3_1 _26072_ (.B(net1027),
    .C(_05284_),
    .A(net1029),
    .Y(_07006_));
 sg13g2_o21ai_1 _26073_ (.B1(_07006_),
    .Y(_07007_),
    .A1(net1029),
    .A2(_07005_));
 sg13g2_nand3_1 _26074_ (.B(net1001),
    .C(_05138_),
    .A(net1029),
    .Y(_07008_));
 sg13g2_nor2b_1 _26075_ (.A(_12024_),
    .B_N(_12030_),
    .Y(_07009_));
 sg13g2_nand2b_1 _26076_ (.Y(_07010_),
    .B(_07009_),
    .A_N(_05411_));
 sg13g2_nand3_1 _26077_ (.B(_07008_),
    .C(_07010_),
    .A(net1028),
    .Y(_07011_));
 sg13g2_o21ai_1 _26078_ (.B1(_07011_),
    .Y(_07012_),
    .A1(net1028),
    .A2(_07007_));
 sg13g2_nand2_1 _26079_ (.Y(_07013_),
    .A(_07004_),
    .B(_07012_));
 sg13g2_a21oi_1 _26080_ (.A1(_05721_),
    .A2(_06926_),
    .Y(_07014_),
    .B1(_11919_));
 sg13g2_mux2_1 _26081_ (.A0(_08950_),
    .A1(net540),
    .S(net829),
    .X(_07015_));
 sg13g2_o21ai_1 _26082_ (.B1(_06935_),
    .Y(_07016_),
    .A1(_00175_),
    .A2(_07015_));
 sg13g2_a221oi_1 _26083_ (.B2(_07014_),
    .C1(_07016_),
    .B1(_07013_),
    .A1(_11938_),
    .Y(_07017_),
    .A2(_06999_));
 sg13g2_nand2_1 _26084_ (.Y(_07018_),
    .A(_06996_),
    .B(_07017_));
 sg13g2_a21oi_1 _26085_ (.A1(_11939_),
    .A2(_06989_),
    .Y(_07019_),
    .B1(_07018_));
 sg13g2_nor2_1 _26086_ (.A(net111),
    .B(_09869_),
    .Y(_07020_));
 sg13g2_nor4_1 _26087_ (.A(_06929_),
    .B(_06931_),
    .C(_06933_),
    .D(_07020_),
    .Y(_07021_));
 sg13g2_nor3_1 _26088_ (.A(_06896_),
    .B(_07019_),
    .C(_07021_),
    .Y(_07022_));
 sg13g2_a21o_1 _26089_ (.A2(_06896_),
    .A1(net13),
    .B1(_07022_),
    .X(_02532_));
 sg13g2_mux2_1 _26090_ (.A0(_09593_),
    .A1(_00225_),
    .S(_06904_),
    .X(_07023_));
 sg13g2_nand2_1 _26091_ (.Y(_07024_),
    .A(net953),
    .B(_10385_));
 sg13g2_o21ai_1 _26092_ (.B1(_07024_),
    .Y(_07025_),
    .A1(_06937_),
    .A2(_07023_));
 sg13g2_nand2_1 _26093_ (.Y(_07026_),
    .A(net363),
    .B(net96));
 sg13g2_o21ai_1 _26094_ (.B1(_07026_),
    .Y(_07027_),
    .A1(_09755_),
    .A2(net96));
 sg13g2_a21oi_1 _26095_ (.A1(_06897_),
    .A2(_07027_),
    .Y(_07028_),
    .B1(_09858_));
 sg13g2_nand2_1 _26096_ (.Y(_07029_),
    .A(_09856_),
    .B(_11914_));
 sg13g2_nor3_1 _26097_ (.A(_09855_),
    .B(_07028_),
    .C(_07029_),
    .Y(_07030_));
 sg13g2_a21oi_1 _26098_ (.A1(_11938_),
    .A2(_07025_),
    .Y(_07031_),
    .B1(_07030_));
 sg13g2_and2_1 _26099_ (.A(net367),
    .B(net96),
    .X(_07032_));
 sg13g2_nor2_1 _26100_ (.A(_09530_),
    .B(net95),
    .Y(_07033_));
 sg13g2_o21ai_1 _26101_ (.B1(net829),
    .Y(_07034_),
    .A1(_07032_),
    .A2(_07033_));
 sg13g2_o21ai_1 _26102_ (.B1(_07034_),
    .Y(_07035_),
    .A1(net727),
    .A2(_08820_));
 sg13g2_nand2b_1 _26103_ (.Y(_07036_),
    .B(net1027),
    .A_N(net1028));
 sg13g2_nand3_1 _26104_ (.B(net1001),
    .C(_05182_),
    .A(net1028),
    .Y(_07037_));
 sg13g2_o21ai_1 _26105_ (.B1(_07037_),
    .Y(_07038_),
    .A1(_05073_),
    .A2(_07036_));
 sg13g2_mux2_1 _26106_ (.A0(_05054_),
    .A1(_05304_),
    .S(net1029),
    .X(_07039_));
 sg13g2_nand2_1 _26107_ (.Y(_07040_),
    .A(net1028),
    .B(net1027));
 sg13g2_mux2_1 _26108_ (.A0(_05480_),
    .A1(_05191_),
    .S(net1029),
    .X(_07041_));
 sg13g2_and2_1 _26109_ (.A(_12047_),
    .B(_12118_),
    .X(_07042_));
 sg13g2_a22oi_1 _26110_ (.Y(_07043_),
    .B1(_07042_),
    .B2(_05473_),
    .A2(_06926_),
    .A1(_05046_));
 sg13g2_o21ai_1 _26111_ (.B1(_07043_),
    .Y(_07044_),
    .A1(_07040_),
    .A2(_07041_));
 sg13g2_a221oi_1 _26112_ (.B2(_06921_),
    .C1(_07044_),
    .B1(_07039_),
    .A1(net1029),
    .Y(_07045_),
    .A2(_07038_));
 sg13g2_nand2_1 _26113_ (.Y(_07046_),
    .A(_08826_),
    .B(net953));
 sg13g2_nand2_1 _26114_ (.Y(_07047_),
    .A(net829),
    .B(net463));
 sg13g2_a21oi_1 _26115_ (.A1(_07046_),
    .A2(_07047_),
    .Y(_07048_),
    .B1(_00175_));
 sg13g2_nor4_1 _26116_ (.A(_11916_),
    .B(_09886_),
    .C(_06934_),
    .D(_07048_),
    .Y(_07049_));
 sg13g2_o21ai_1 _26117_ (.B1(_07049_),
    .Y(_07050_),
    .A1(_11919_),
    .A2(_07045_));
 sg13g2_a21oi_1 _26118_ (.A1(_11942_),
    .A2(_07035_),
    .Y(_07051_),
    .B1(_07050_));
 sg13g2_nor2_1 _26119_ (.A(_09638_),
    .B(_06900_),
    .Y(_07052_));
 sg13g2_a21oi_1 _26120_ (.A1(_00217_),
    .A2(net96),
    .Y(_07053_),
    .B1(_07052_));
 sg13g2_nand2_1 _26121_ (.Y(_07054_),
    .A(_06897_),
    .B(_07053_));
 sg13g2_o21ai_1 _26122_ (.B1(_07054_),
    .Y(_07055_),
    .A1(net727),
    .A2(_10733_));
 sg13g2_mux2_1 _26123_ (.A0(_09777_),
    .A1(net419),
    .S(net96),
    .X(_07056_));
 sg13g2_nand2_1 _26124_ (.Y(_07057_),
    .A(net727),
    .B(_07056_));
 sg13g2_o21ai_1 _26125_ (.B1(_07057_),
    .Y(_07058_),
    .A1(net727),
    .A2(_08663_));
 sg13g2_a22oi_1 _26126_ (.Y(_07059_),
    .B1(_07058_),
    .B2(_11918_),
    .A2(_07055_),
    .A1(_11939_));
 sg13g2_and3_1 _26127_ (.X(_07060_),
    .A(_07031_),
    .B(_07051_),
    .C(_07059_));
 sg13g2_nor3_1 _26128_ (.A(_06896_),
    .B(_07021_),
    .C(_07060_),
    .Y(_07061_));
 sg13g2_a21o_1 _26129_ (.A2(_06896_),
    .A1(net14),
    .B1(_07061_),
    .X(_02533_));
 sg13g2_nand2_1 _26130_ (.Y(_07062_),
    .A(_09248_),
    .B(net404));
 sg13g2_buf_1 _26131_ (.A(_07062_),
    .X(_07063_));
 sg13g2_mux2_1 _26132_ (.A0(net913),
    .A1(\cpu.spi.r_clk_count[0][0] ),
    .S(net94),
    .X(_02538_));
 sg13g2_mux2_1 _26133_ (.A0(net853),
    .A1(\cpu.spi.r_clk_count[0][1] ),
    .S(net94),
    .X(_02539_));
 sg13g2_mux2_1 _26134_ (.A0(net845),
    .A1(\cpu.spi.r_clk_count[0][2] ),
    .S(_07063_),
    .X(_02540_));
 sg13g2_mux2_1 _26135_ (.A0(net964),
    .A1(\cpu.spi.r_clk_count[0][3] ),
    .S(net94),
    .X(_02541_));
 sg13g2_nand2_1 _26136_ (.Y(_07064_),
    .A(\cpu.spi.r_clk_count[0][4] ),
    .B(net94));
 sg13g2_o21ai_1 _26137_ (.B1(_07064_),
    .Y(_02542_),
    .A1(net883),
    .A2(net94));
 sg13g2_nand2_1 _26138_ (.Y(_07065_),
    .A(\cpu.spi.r_clk_count[0][5] ),
    .B(net94));
 sg13g2_o21ai_1 _26139_ (.B1(_07065_),
    .Y(_02543_),
    .A1(net882),
    .A2(net94));
 sg13g2_nand2_1 _26140_ (.Y(_07066_),
    .A(\cpu.spi.r_clk_count[0][6] ),
    .B(_07062_));
 sg13g2_o21ai_1 _26141_ (.B1(_07066_),
    .Y(_02544_),
    .A1(net881),
    .A2(net94));
 sg13g2_mux2_1 _26142_ (.A0(net1023),
    .A1(\cpu.spi.r_clk_count[0][7] ),
    .S(_07063_),
    .X(_02545_));
 sg13g2_nand4_1 _26143_ (.B(net550),
    .C(_09248_),
    .A(net1043),
    .Y(_07067_),
    .D(net499));
 sg13g2_buf_1 _26144_ (.A(_07067_),
    .X(_07068_));
 sg13g2_buf_1 _26145_ (.A(_07068_),
    .X(_07069_));
 sg13g2_mux2_1 _26146_ (.A0(net913),
    .A1(\cpu.spi.r_clk_count[1][0] ),
    .S(net84),
    .X(_02546_));
 sg13g2_mux2_1 _26147_ (.A0(net853),
    .A1(\cpu.spi.r_clk_count[1][1] ),
    .S(net84),
    .X(_02547_));
 sg13g2_mux2_1 _26148_ (.A0(net845),
    .A1(\cpu.spi.r_clk_count[1][2] ),
    .S(net84),
    .X(_02548_));
 sg13g2_mux2_1 _26149_ (.A0(net964),
    .A1(\cpu.spi.r_clk_count[1][3] ),
    .S(net84),
    .X(_02549_));
 sg13g2_nand2_1 _26150_ (.Y(_07070_),
    .A(\cpu.spi.r_clk_count[1][4] ),
    .B(net84));
 sg13g2_o21ai_1 _26151_ (.B1(_07070_),
    .Y(_02550_),
    .A1(net883),
    .A2(net84));
 sg13g2_nand2_1 _26152_ (.Y(_07071_),
    .A(\cpu.spi.r_clk_count[1][5] ),
    .B(net84));
 sg13g2_o21ai_1 _26153_ (.B1(_07071_),
    .Y(_02551_),
    .A1(net882),
    .A2(net84));
 sg13g2_nand2_1 _26154_ (.Y(_07072_),
    .A(\cpu.spi.r_clk_count[1][6] ),
    .B(_07068_));
 sg13g2_o21ai_1 _26155_ (.B1(_07072_),
    .Y(_02552_),
    .A1(net881),
    .A2(_07069_));
 sg13g2_mux2_1 _26156_ (.A0(net1023),
    .A1(\cpu.spi.r_clk_count[1][7] ),
    .S(_07069_),
    .X(_02553_));
 sg13g2_nand2_1 _26157_ (.Y(_07073_),
    .A(net888),
    .B(_04968_));
 sg13g2_nor4_1 _26158_ (.A(net622),
    .B(net926),
    .C(_09300_),
    .D(_07073_),
    .Y(_07074_));
 sg13g2_buf_4 _26159_ (.X(_07075_),
    .A(_07074_));
 sg13g2_mux2_1 _26160_ (.A0(_04983_),
    .A1(net911),
    .S(_07075_),
    .X(_02554_));
 sg13g2_mux2_1 _26161_ (.A0(_05372_),
    .A1(net885),
    .S(_07075_),
    .X(_02555_));
 sg13g2_mux2_1 _26162_ (.A0(_05445_),
    .A1(net884),
    .S(_07075_),
    .X(_02556_));
 sg13g2_mux2_1 _26163_ (.A0(_05487_),
    .A1(net1024),
    .S(_07075_),
    .X(_02557_));
 sg13g2_mux2_1 _26164_ (.A0(_05530_),
    .A1(net1059),
    .S(_07075_),
    .X(_02558_));
 sg13g2_mux2_1 _26165_ (.A0(_05626_),
    .A1(net1058),
    .S(_07075_),
    .X(_02559_));
 sg13g2_mux2_1 _26166_ (.A0(_05696_),
    .A1(net1057),
    .S(_07075_),
    .X(_02560_));
 sg13g2_mux2_1 _26167_ (.A0(_05114_),
    .A1(net1018),
    .S(_07075_),
    .X(_02561_));
 sg13g2_inv_1 _26168_ (.Y(_07076_),
    .A(_09325_));
 sg13g2_buf_2 _26169_ (.A(_00210_),
    .X(_07077_));
 sg13g2_nor4_2 _26170_ (.A(\cpu.spi.r_state[5] ),
    .B(net1135),
    .C(_09321_),
    .Y(_07078_),
    .D(_11945_));
 sg13g2_nand3_1 _26171_ (.B(_07077_),
    .C(_07078_),
    .A(_07076_),
    .Y(_07079_));
 sg13g2_inv_1 _26172_ (.Y(_07080_),
    .A(_07077_));
 sg13g2_nand3_1 _26173_ (.B(_09302_),
    .C(_09308_),
    .A(_07080_),
    .Y(_07081_));
 sg13g2_o21ai_1 _26174_ (.B1(_09320_),
    .Y(_07082_),
    .A1(_09237_),
    .A2(net517));
 sg13g2_nand4_1 _26175_ (.B(_07079_),
    .C(_07081_),
    .A(_09359_),
    .Y(_07083_),
    .D(_07082_));
 sg13g2_buf_2 _26176_ (.A(_07083_),
    .X(_07084_));
 sg13g2_buf_1 _26177_ (.A(_07084_),
    .X(_07085_));
 sg13g2_buf_1 _26178_ (.A(net563),
    .X(_07086_));
 sg13g2_nand2b_1 _26179_ (.Y(_07087_),
    .B(net467),
    .A_N(\cpu.spi.r_clk_count[0][0] ));
 sg13g2_o21ai_1 _26180_ (.B1(_07087_),
    .Y(_07088_),
    .A1(net490),
    .A2(_04983_));
 sg13g2_mux2_1 _26181_ (.A0(\cpu.spi.r_clk_count[0][0] ),
    .A1(\cpu.spi.r_clk_count[1][0] ),
    .S(net563),
    .X(_07089_));
 sg13g2_nor2_1 _26182_ (.A(net749),
    .B(_07089_),
    .Y(_07090_));
 sg13g2_a21oi_1 _26183_ (.A1(net749),
    .A2(_07088_),
    .Y(_07091_),
    .B1(_07090_));
 sg13g2_nand2_1 _26184_ (.Y(_07092_),
    .A(_07077_),
    .B(_07078_));
 sg13g2_buf_1 _26185_ (.A(_07092_),
    .X(_07093_));
 sg13g2_buf_1 _26186_ (.A(_07093_),
    .X(_07094_));
 sg13g2_buf_1 _26187_ (.A(net1115),
    .X(_07095_));
 sg13g2_mux2_1 _26188_ (.A0(_00298_),
    .A1(_00297_),
    .S(net952),
    .X(_07096_));
 sg13g2_buf_1 _26189_ (.A(_11951_),
    .X(_07097_));
 sg13g2_nor2_1 _26190_ (.A(net1032),
    .B(_04983_),
    .Y(_07098_));
 sg13g2_a21oi_1 _26191_ (.A1(_07095_),
    .A2(_00298_),
    .Y(_07099_),
    .B1(_07098_));
 sg13g2_nand2_1 _26192_ (.Y(_07100_),
    .A(_07097_),
    .B(_07099_));
 sg13g2_o21ai_1 _26193_ (.B1(_07100_),
    .Y(_07101_),
    .A1(net1033),
    .A2(_07096_));
 sg13g2_nand2_1 _26194_ (.Y(_07102_),
    .A(net100),
    .B(_07101_));
 sg13g2_o21ai_1 _26195_ (.B1(_07102_),
    .Y(_07103_),
    .A1(_09279_),
    .A2(_09303_));
 sg13g2_buf_1 _26196_ (.A(_07078_),
    .X(_07104_));
 sg13g2_nor2_1 _26197_ (.A(net422),
    .B(_07101_),
    .Y(_07105_));
 sg13g2_nor3_1 _26198_ (.A(_09279_),
    .B(_07104_),
    .C(_07105_),
    .Y(_07106_));
 sg13g2_a21oi_1 _26199_ (.A1(_09289_),
    .A2(_07103_),
    .Y(_07107_),
    .B1(_07106_));
 sg13g2_nand2_1 _26200_ (.Y(_07108_),
    .A(net524),
    .B(_07107_));
 sg13g2_o21ai_1 _26201_ (.B1(_07108_),
    .Y(_07109_),
    .A1(_07091_),
    .A2(net524));
 sg13g2_nand2_1 _26202_ (.Y(_07110_),
    .A(_09279_),
    .B(net30));
 sg13g2_o21ai_1 _26203_ (.B1(_07110_),
    .Y(_02562_),
    .A1(net30),
    .A2(_07109_));
 sg13g2_nand2b_1 _26204_ (.Y(_07111_),
    .B(net490),
    .A_N(\cpu.spi.r_clk_count[0][1] ));
 sg13g2_o21ai_1 _26205_ (.B1(_07111_),
    .Y(_07112_),
    .A1(net490),
    .A2(_05372_));
 sg13g2_mux2_1 _26206_ (.A0(\cpu.spi.r_clk_count[0][1] ),
    .A1(\cpu.spi.r_clk_count[1][1] ),
    .S(_07086_),
    .X(_07113_));
 sg13g2_nor2_1 _26207_ (.A(net749),
    .B(_07113_),
    .Y(_07114_));
 sg13g2_a21oi_1 _26208_ (.A1(net745),
    .A2(_07112_),
    .Y(_07115_),
    .B1(_07114_));
 sg13g2_xor2_1 _26209_ (.B(\cpu.spi.r_count[1] ),
    .A(_09279_),
    .X(_07116_));
 sg13g2_nand2_1 _26210_ (.Y(_07117_),
    .A(net1032),
    .B(_00302_));
 sg13g2_o21ai_1 _26211_ (.B1(_07117_),
    .Y(_07118_),
    .A1(net1031),
    .A2(_05370_));
 sg13g2_nor2_1 _26212_ (.A(net1032),
    .B(_05372_),
    .Y(_07119_));
 sg13g2_a21oi_1 _26213_ (.A1(_07095_),
    .A2(_00091_),
    .Y(_07120_),
    .B1(_07119_));
 sg13g2_nand2_1 _26214_ (.Y(_07121_),
    .A(net951),
    .B(_07120_));
 sg13g2_o21ai_1 _26215_ (.B1(_07121_),
    .Y(_07122_),
    .A1(net1033),
    .A2(_07118_));
 sg13g2_nand2_1 _26216_ (.Y(_07123_),
    .A(net100),
    .B(_07122_));
 sg13g2_o21ai_1 _26217_ (.B1(_07123_),
    .Y(_07124_),
    .A1(net91),
    .A2(_07116_));
 sg13g2_nor2_1 _26218_ (.A(net462),
    .B(_07122_),
    .Y(_07125_));
 sg13g2_nor3_1 _26219_ (.A(_07104_),
    .B(_07125_),
    .C(_07116_),
    .Y(_07126_));
 sg13g2_a21oi_1 _26220_ (.A1(net1070),
    .A2(_07124_),
    .Y(_07127_),
    .B1(_07126_));
 sg13g2_nand2_1 _26221_ (.Y(_07128_),
    .A(_07094_),
    .B(_07127_));
 sg13g2_o21ai_1 _26222_ (.B1(_07128_),
    .Y(_07129_),
    .A1(_07094_),
    .A2(_07115_));
 sg13g2_nand2_1 _26223_ (.Y(_07130_),
    .A(\cpu.spi.r_count[1] ),
    .B(_07085_));
 sg13g2_o21ai_1 _26224_ (.B1(_07130_),
    .Y(_02563_),
    .A1(net30),
    .A2(_07129_));
 sg13g2_nand2b_1 _26225_ (.Y(_07131_),
    .B(_03512_),
    .A_N(\cpu.spi.r_clk_count[0][2] ));
 sg13g2_o21ai_1 _26226_ (.B1(_07131_),
    .Y(_07132_),
    .A1(_03512_),
    .A2(_05445_));
 sg13g2_mux2_1 _26227_ (.A0(\cpu.spi.r_clk_count[0][2] ),
    .A1(\cpu.spi.r_clk_count[1][2] ),
    .S(net467),
    .X(_07133_));
 sg13g2_nor2_1 _26228_ (.A(net749),
    .B(_07133_),
    .Y(_07134_));
 sg13g2_a21oi_1 _26229_ (.A1(net745),
    .A2(_07132_),
    .Y(_07135_),
    .B1(_07134_));
 sg13g2_xnor2_1 _26230_ (.Y(_07136_),
    .A(\cpu.spi.r_count[2] ),
    .B(_09280_));
 sg13g2_nand2_1 _26231_ (.Y(_07137_),
    .A(net1032),
    .B(_00100_));
 sg13g2_o21ai_1 _26232_ (.B1(_07137_),
    .Y(_07138_),
    .A1(net1031),
    .A2(_05444_));
 sg13g2_nor2_1 _26233_ (.A(net1115),
    .B(_05445_),
    .Y(_07139_));
 sg13g2_a21oi_1 _26234_ (.A1(net952),
    .A2(_00101_),
    .Y(_07140_),
    .B1(_07139_));
 sg13g2_nand2_1 _26235_ (.Y(_07141_),
    .A(_07097_),
    .B(_07140_));
 sg13g2_o21ai_1 _26236_ (.B1(_07141_),
    .Y(_07142_),
    .A1(net1033),
    .A2(_07138_));
 sg13g2_nand2_1 _26237_ (.Y(_07143_),
    .A(net100),
    .B(_07142_));
 sg13g2_o21ai_1 _26238_ (.B1(_07143_),
    .Y(_07144_),
    .A1(net91),
    .A2(_07136_));
 sg13g2_nor2_1 _26239_ (.A(net462),
    .B(_07142_),
    .Y(_07145_));
 sg13g2_nor3_1 _26240_ (.A(net655),
    .B(_07145_),
    .C(_07136_),
    .Y(_07146_));
 sg13g2_a21oi_1 _26241_ (.A1(net1070),
    .A2(_07144_),
    .Y(_07147_),
    .B1(_07146_));
 sg13g2_nand2_1 _26242_ (.Y(_07148_),
    .A(net524),
    .B(_07147_));
 sg13g2_o21ai_1 _26243_ (.B1(_07148_),
    .Y(_07149_),
    .A1(net524),
    .A2(_07135_));
 sg13g2_nand2_1 _26244_ (.Y(_07150_),
    .A(\cpu.spi.r_count[2] ),
    .B(_07084_));
 sg13g2_o21ai_1 _26245_ (.B1(_07150_),
    .Y(_02564_),
    .A1(_07085_),
    .A2(_07149_));
 sg13g2_nand2b_1 _26246_ (.Y(_07151_),
    .B(net467),
    .A_N(\cpu.spi.r_clk_count[0][3] ));
 sg13g2_o21ai_1 _26247_ (.B1(_07151_),
    .Y(_07152_),
    .A1(net490),
    .A2(_05487_));
 sg13g2_mux2_1 _26248_ (.A0(\cpu.spi.r_clk_count[0][3] ),
    .A1(\cpu.spi.r_clk_count[1][3] ),
    .S(net467),
    .X(_07153_));
 sg13g2_nor2_1 _26249_ (.A(net749),
    .B(_07153_),
    .Y(_07154_));
 sg13g2_a21oi_1 _26250_ (.A1(net745),
    .A2(_07152_),
    .Y(_07155_),
    .B1(_07154_));
 sg13g2_xor2_1 _26251_ (.B(_09281_),
    .A(_09278_),
    .X(_07156_));
 sg13g2_mux2_1 _26252_ (.A0(_00111_),
    .A1(_00110_),
    .S(net952),
    .X(_07157_));
 sg13g2_nor2_1 _26253_ (.A(net1032),
    .B(_05487_),
    .Y(_07158_));
 sg13g2_a21oi_1 _26254_ (.A1(net952),
    .A2(_00111_),
    .Y(_07159_),
    .B1(_07158_));
 sg13g2_nand2_1 _26255_ (.Y(_07160_),
    .A(net951),
    .B(_07159_));
 sg13g2_o21ai_1 _26256_ (.B1(_07160_),
    .Y(_07161_),
    .A1(net1033),
    .A2(_07157_));
 sg13g2_nand2_1 _26257_ (.Y(_07162_),
    .A(net100),
    .B(_07161_));
 sg13g2_o21ai_1 _26258_ (.B1(_07162_),
    .Y(_07163_),
    .A1(net91),
    .A2(_07156_));
 sg13g2_nor2_1 _26259_ (.A(net462),
    .B(_07161_),
    .Y(_07164_));
 sg13g2_nor3_1 _26260_ (.A(net655),
    .B(_07156_),
    .C(_07164_),
    .Y(_07165_));
 sg13g2_a21oi_1 _26261_ (.A1(net1070),
    .A2(_07163_),
    .Y(_07166_),
    .B1(_07165_));
 sg13g2_nand2_1 _26262_ (.Y(_07167_),
    .A(_07093_),
    .B(_07166_));
 sg13g2_o21ai_1 _26263_ (.B1(_07167_),
    .Y(_07168_),
    .A1(net524),
    .A2(_07155_));
 sg13g2_nand2_1 _26264_ (.Y(_07169_),
    .A(_09278_),
    .B(_07084_));
 sg13g2_o21ai_1 _26265_ (.B1(_07169_),
    .Y(_02565_),
    .A1(net30),
    .A2(_07168_));
 sg13g2_nand2b_1 _26266_ (.Y(_07170_),
    .B(net467),
    .A_N(\cpu.spi.r_clk_count[0][4] ));
 sg13g2_o21ai_1 _26267_ (.B1(_07170_),
    .Y(_07171_),
    .A1(net490),
    .A2(_05530_));
 sg13g2_mux2_1 _26268_ (.A0(\cpu.spi.r_clk_count[0][4] ),
    .A1(\cpu.spi.r_clk_count[1][4] ),
    .S(net467),
    .X(_07172_));
 sg13g2_nor2_1 _26269_ (.A(net749),
    .B(_07172_),
    .Y(_07173_));
 sg13g2_a21oi_1 _26270_ (.A1(net745),
    .A2(_07171_),
    .Y(_07174_),
    .B1(_07173_));
 sg13g2_nor2_1 _26271_ (.A(_09278_),
    .B(_09281_),
    .Y(_07175_));
 sg13g2_xnor2_1 _26272_ (.Y(_07176_),
    .A(\cpu.spi.r_count[4] ),
    .B(_07175_));
 sg13g2_mux2_1 _26273_ (.A0(_00121_),
    .A1(_00120_),
    .S(net952),
    .X(_07177_));
 sg13g2_nor2_1 _26274_ (.A(net1032),
    .B(_05530_),
    .Y(_07178_));
 sg13g2_a21oi_1 _26275_ (.A1(net952),
    .A2(_00121_),
    .Y(_07179_),
    .B1(_07178_));
 sg13g2_nand2_1 _26276_ (.Y(_07180_),
    .A(net951),
    .B(_07179_));
 sg13g2_o21ai_1 _26277_ (.B1(_07180_),
    .Y(_07181_),
    .A1(net1033),
    .A2(_07177_));
 sg13g2_nand2_1 _26278_ (.Y(_07182_),
    .A(net100),
    .B(_07181_));
 sg13g2_o21ai_1 _26279_ (.B1(_07182_),
    .Y(_07183_),
    .A1(net91),
    .A2(_07176_));
 sg13g2_nor2_1 _26280_ (.A(net462),
    .B(_07181_),
    .Y(_07184_));
 sg13g2_nor3_1 _26281_ (.A(net655),
    .B(_07176_),
    .C(_07184_),
    .Y(_07185_));
 sg13g2_a21oi_1 _26282_ (.A1(net1070),
    .A2(_07183_),
    .Y(_07186_),
    .B1(_07185_));
 sg13g2_nand2_1 _26283_ (.Y(_07187_),
    .A(_07093_),
    .B(_07186_));
 sg13g2_o21ai_1 _26284_ (.B1(_07187_),
    .Y(_07188_),
    .A1(net524),
    .A2(_07174_));
 sg13g2_nand2_1 _26285_ (.Y(_07189_),
    .A(\cpu.spi.r_count[4] ),
    .B(_07084_));
 sg13g2_o21ai_1 _26286_ (.B1(_07189_),
    .Y(_02566_),
    .A1(net30),
    .A2(_07188_));
 sg13g2_nand2b_1 _26287_ (.Y(_07190_),
    .B(net467),
    .A_N(\cpu.spi.r_clk_count[0][5] ));
 sg13g2_o21ai_1 _26288_ (.B1(_07190_),
    .Y(_07191_),
    .A1(net490),
    .A2(_05626_));
 sg13g2_mux2_1 _26289_ (.A0(\cpu.spi.r_clk_count[0][5] ),
    .A1(\cpu.spi.r_clk_count[1][5] ),
    .S(net467),
    .X(_07192_));
 sg13g2_nor2_1 _26290_ (.A(net749),
    .B(_07192_),
    .Y(_07193_));
 sg13g2_a21oi_1 _26291_ (.A1(net745),
    .A2(_07191_),
    .Y(_07194_),
    .B1(_07193_));
 sg13g2_xnor2_1 _26292_ (.Y(_07195_),
    .A(\cpu.spi.r_count[5] ),
    .B(_09282_));
 sg13g2_mux2_1 _26293_ (.A0(_00127_),
    .A1(_00126_),
    .S(net1032),
    .X(_07196_));
 sg13g2_nor2_1 _26294_ (.A(net1115),
    .B(_05626_),
    .Y(_07197_));
 sg13g2_a21oi_1 _26295_ (.A1(net952),
    .A2(_00127_),
    .Y(_07198_),
    .B1(_07197_));
 sg13g2_nand2_1 _26296_ (.Y(_07199_),
    .A(net951),
    .B(_07198_));
 sg13g2_o21ai_1 _26297_ (.B1(_07199_),
    .Y(_07200_),
    .A1(net951),
    .A2(_07196_));
 sg13g2_nand2_1 _26298_ (.Y(_07201_),
    .A(net100),
    .B(_07200_));
 sg13g2_o21ai_1 _26299_ (.B1(_07201_),
    .Y(_07202_),
    .A1(net91),
    .A2(_07195_));
 sg13g2_nor2_1 _26300_ (.A(net462),
    .B(_07200_),
    .Y(_07203_));
 sg13g2_nor3_1 _26301_ (.A(net655),
    .B(_07203_),
    .C(_07195_),
    .Y(_07204_));
 sg13g2_a21oi_1 _26302_ (.A1(net1070),
    .A2(_07202_),
    .Y(_07205_),
    .B1(_07204_));
 sg13g2_nand2_1 _26303_ (.Y(_07206_),
    .A(_07093_),
    .B(_07205_));
 sg13g2_o21ai_1 _26304_ (.B1(_07206_),
    .Y(_07207_),
    .A1(net524),
    .A2(_07194_));
 sg13g2_nand2_1 _26305_ (.Y(_07208_),
    .A(\cpu.spi.r_count[5] ),
    .B(_07084_));
 sg13g2_o21ai_1 _26306_ (.B1(_07208_),
    .Y(_02567_),
    .A1(net30),
    .A2(_07207_));
 sg13g2_nand2b_1 _26307_ (.Y(_07209_),
    .B(_07086_),
    .A_N(\cpu.spi.r_clk_count[0][6] ));
 sg13g2_o21ai_1 _26308_ (.B1(_07209_),
    .Y(_07210_),
    .A1(net490),
    .A2(_05696_));
 sg13g2_mux2_1 _26309_ (.A0(\cpu.spi.r_clk_count[0][6] ),
    .A1(\cpu.spi.r_clk_count[1][6] ),
    .S(net563),
    .X(_07211_));
 sg13g2_nor2_1 _26310_ (.A(net749),
    .B(_07211_),
    .Y(_07212_));
 sg13g2_a21oi_1 _26311_ (.A1(net745),
    .A2(_07210_),
    .Y(_07213_),
    .B1(_07212_));
 sg13g2_xnor2_1 _26312_ (.Y(_07214_),
    .A(\cpu.spi.r_count[6] ),
    .B(_09283_));
 sg13g2_mux2_1 _26313_ (.A0(_00138_),
    .A1(_00137_),
    .S(net1032),
    .X(_07215_));
 sg13g2_nor2_1 _26314_ (.A(net1115),
    .B(_05696_),
    .Y(_07216_));
 sg13g2_a21oi_1 _26315_ (.A1(net952),
    .A2(_00138_),
    .Y(_07217_),
    .B1(_07216_));
 sg13g2_nand2_1 _26316_ (.Y(_07218_),
    .A(net951),
    .B(_07217_));
 sg13g2_o21ai_1 _26317_ (.B1(_07218_),
    .Y(_07219_),
    .A1(net951),
    .A2(_07215_));
 sg13g2_nand2_1 _26318_ (.Y(_07220_),
    .A(net100),
    .B(_07219_));
 sg13g2_o21ai_1 _26319_ (.B1(_07220_),
    .Y(_07221_),
    .A1(net91),
    .A2(_07214_));
 sg13g2_nor2_1 _26320_ (.A(net462),
    .B(_07219_),
    .Y(_07222_));
 sg13g2_nor3_1 _26321_ (.A(net655),
    .B(_07222_),
    .C(_07214_),
    .Y(_07223_));
 sg13g2_a21oi_1 _26322_ (.A1(net1070),
    .A2(_07221_),
    .Y(_07224_),
    .B1(_07223_));
 sg13g2_nand2_1 _26323_ (.Y(_07225_),
    .A(_07093_),
    .B(_07224_));
 sg13g2_o21ai_1 _26324_ (.B1(_07225_),
    .Y(_07226_),
    .A1(net524),
    .A2(_07213_));
 sg13g2_nand2_1 _26325_ (.Y(_07227_),
    .A(\cpu.spi.r_count[6] ),
    .B(_07084_));
 sg13g2_o21ai_1 _26326_ (.B1(_07227_),
    .Y(_02568_),
    .A1(net30),
    .A2(_07226_));
 sg13g2_nor2_1 _26327_ (.A(net1031),
    .B(_05114_),
    .Y(_07228_));
 sg13g2_a21oi_1 _26328_ (.A1(net1031),
    .A2(_00149_),
    .Y(_07229_),
    .B1(_07228_));
 sg13g2_mux2_1 _26329_ (.A0(_00149_),
    .A1(_00148_),
    .S(net1031),
    .X(_07230_));
 sg13g2_nor2_1 _26330_ (.A(net1033),
    .B(_07230_),
    .Y(_07231_));
 sg13g2_a21oi_1 _26331_ (.A1(net1033),
    .A2(_07229_),
    .Y(_07232_),
    .B1(_07231_));
 sg13g2_nor2b_1 _26332_ (.A(_09284_),
    .B_N(_09277_),
    .Y(_07233_));
 sg13g2_o21ai_1 _26333_ (.B1(_09249_),
    .Y(_07234_),
    .A1(net517),
    .A2(_07233_));
 sg13g2_o21ai_1 _26334_ (.B1(_07234_),
    .Y(_07235_),
    .A1(_09249_),
    .A2(_07232_));
 sg13g2_buf_1 _26335_ (.A(_09319_),
    .X(_07236_));
 sg13g2_a21oi_1 _26336_ (.A1(_07077_),
    .A2(net655),
    .Y(_07237_),
    .B1(_07236_));
 sg13g2_and2_1 _26337_ (.A(net563),
    .B(\cpu.spi.r_clk_count[1][7] ),
    .X(_07238_));
 sg13g2_a21oi_1 _26338_ (.A1(net783),
    .A2(\cpu.spi.r_clk_count[0][7] ),
    .Y(_07239_),
    .B1(_07238_));
 sg13g2_mux2_1 _26339_ (.A0(_05114_),
    .A1(\cpu.spi.r_clk_count[0][7] ),
    .S(net563),
    .X(_07240_));
 sg13g2_nand2_1 _26340_ (.Y(_07241_),
    .A(net888),
    .B(_07240_));
 sg13g2_o21ai_1 _26341_ (.B1(_07241_),
    .Y(_07242_),
    .A1(net888),
    .A2(_07239_));
 sg13g2_nand2_1 _26342_ (.Y(_07243_),
    .A(_07077_),
    .B(_07242_));
 sg13g2_nor2_1 _26343_ (.A(net422),
    .B(_07232_),
    .Y(_07244_));
 sg13g2_nor3_1 _26344_ (.A(net655),
    .B(_07233_),
    .C(_07244_),
    .Y(_07245_));
 sg13g2_a21oi_1 _26345_ (.A1(net655),
    .A2(_07243_),
    .Y(_07246_),
    .B1(_07245_));
 sg13g2_a21oi_1 _26346_ (.A1(_07235_),
    .A2(_07237_),
    .Y(_07247_),
    .B1(_07246_));
 sg13g2_nand2_1 _26347_ (.Y(_07248_),
    .A(_09277_),
    .B(_07084_));
 sg13g2_o21ai_1 _26348_ (.B1(_07248_),
    .Y(_02569_),
    .A1(net30),
    .A2(_07247_));
 sg13g2_inv_1 _26349_ (.Y(_07249_),
    .A(\cpu.gpio.r_spi_miso_src[1][1] ));
 sg13g2_mux4_1 _26350_ (.S0(_05550_),
    .A0(_09180_),
    .A1(_09182_),
    .A2(_09177_),
    .A3(_09193_),
    .S1(\cpu.gpio.r_spi_miso_src[1][2] ),
    .X(_07250_));
 sg13g2_nand2_1 _26351_ (.Y(_07251_),
    .A(_09195_),
    .B(_05550_));
 sg13g2_nand2b_1 _26352_ (.Y(_07252_),
    .B(_09200_),
    .A_N(_05550_));
 sg13g2_nand3_1 _26353_ (.B(_07251_),
    .C(_07252_),
    .A(_06431_),
    .Y(_07253_));
 sg13g2_o21ai_1 _26354_ (.B1(_07253_),
    .Y(_07254_),
    .A1(_06431_),
    .A2(_07250_));
 sg13g2_nand2b_1 _26355_ (.Y(_07255_),
    .B(_05550_),
    .A_N(_09191_));
 sg13g2_o21ai_1 _26356_ (.B1(_07255_),
    .Y(_07256_),
    .A1(_09188_),
    .A2(_05550_));
 sg13g2_a21o_1 _26357_ (.A2(_07256_),
    .A1(\cpu.gpio.r_spi_miso_src[1][1] ),
    .B1(_00143_),
    .X(_07257_));
 sg13g2_mux4_1 _26358_ (.S0(_05550_),
    .A0(_09190_),
    .A1(_09198_),
    .A2(_09175_),
    .A3(_09186_),
    .S1(\cpu.gpio.r_spi_miso_src[1][2] ),
    .X(_07258_));
 sg13g2_nor3_1 _26359_ (.A(_07249_),
    .B(_06431_),
    .C(_07258_),
    .Y(_07259_));
 sg13g2_a221oi_1 _26360_ (.B2(_06431_),
    .C1(_07259_),
    .B1(_07257_),
    .A1(_07249_),
    .Y(_07260_),
    .A2(_07254_));
 sg13g2_mux4_1 _26361_ (.S0(_04923_),
    .A0(_09190_),
    .A1(_09198_),
    .A2(_09175_),
    .A3(_09186_),
    .S1(\cpu.gpio.r_spi_miso_src[0][2] ),
    .X(_07261_));
 sg13g2_nand2_1 _26362_ (.Y(_07262_),
    .A(_09191_),
    .B(_04923_));
 sg13g2_nand2b_1 _26363_ (.Y(_07263_),
    .B(_09188_),
    .A_N(_04923_));
 sg13g2_nand3_1 _26364_ (.B(_07262_),
    .C(_07263_),
    .A(_06427_),
    .Y(_07264_));
 sg13g2_o21ai_1 _26365_ (.B1(_07264_),
    .Y(_07265_),
    .A1(_06427_),
    .A2(_07261_));
 sg13g2_mux2_1 _26366_ (.A0(_09200_),
    .A1(_09195_),
    .S(_04923_),
    .X(_07266_));
 sg13g2_o21ai_1 _26367_ (.B1(_05425_),
    .Y(_07267_),
    .A1(_06425_),
    .A2(_07266_));
 sg13g2_mux4_1 _26368_ (.S0(_04923_),
    .A0(_09180_),
    .A1(_09182_),
    .A2(_09177_),
    .A3(_09193_),
    .S1(\cpu.gpio.r_spi_miso_src[0][2] ),
    .X(_07268_));
 sg13g2_nor3_1 _26369_ (.A(_06425_),
    .B(_06427_),
    .C(_07268_),
    .Y(_07269_));
 sg13g2_a221oi_1 _26370_ (.B2(_06427_),
    .C1(_07269_),
    .B1(_07267_),
    .A1(_06425_),
    .Y(_07270_),
    .A2(_07265_));
 sg13g2_mux2_1 _26371_ (.A0(_07260_),
    .A1(_07270_),
    .S(_11961_),
    .X(_07271_));
 sg13g2_nor2_1 _26372_ (.A(net1134),
    .B(net672),
    .Y(_07272_));
 sg13g2_nor2b_1 _26373_ (.A(_09252_),
    .B_N(net1134),
    .Y(_07273_));
 sg13g2_a22oi_1 _26374_ (.Y(_07274_),
    .B1(_07273_),
    .B2(net672),
    .A2(_07272_),
    .A1(_09252_));
 sg13g2_nor3_1 _26375_ (.A(net923),
    .B(net422),
    .C(_07274_),
    .Y(_07275_));
 sg13g2_buf_4 _26376_ (.X(_07276_),
    .A(_07275_));
 sg13g2_mux2_1 _26377_ (.A0(_09267_),
    .A1(_07271_),
    .S(_07276_),
    .X(_02573_));
 sg13g2_mux2_1 _26378_ (.A0(_09266_),
    .A1(_09267_),
    .S(_07276_),
    .X(_02574_));
 sg13g2_mux2_1 _26379_ (.A0(_09270_),
    .A1(_09266_),
    .S(_07276_),
    .X(_02575_));
 sg13g2_mux2_1 _26380_ (.A0(_09264_),
    .A1(_09270_),
    .S(_07276_),
    .X(_02576_));
 sg13g2_mux2_1 _26381_ (.A0(_09272_),
    .A1(_09264_),
    .S(_07276_),
    .X(_02577_));
 sg13g2_mux2_1 _26382_ (.A0(_09271_),
    .A1(_09272_),
    .S(_07276_),
    .X(_02578_));
 sg13g2_mux2_1 _26383_ (.A0(_09265_),
    .A1(_09271_),
    .S(_07276_),
    .X(_02579_));
 sg13g2_mux2_1 _26384_ (.A0(\cpu.spi.r_in[7] ),
    .A1(_09265_),
    .S(_07276_),
    .X(_02580_));
 sg13g2_nand3_1 _26385_ (.B(_09248_),
    .C(_04885_),
    .A(_04967_),
    .Y(_07277_));
 sg13g2_nor3_2 _26386_ (.A(net491),
    .B(net452),
    .C(_07277_),
    .Y(_07278_));
 sg13g2_mux2_1 _26387_ (.A0(\cpu.spi.r_mode[0][0] ),
    .A1(_10099_),
    .S(_07278_),
    .X(_02582_));
 sg13g2_mux2_1 _26388_ (.A0(_11965_),
    .A1(net885),
    .S(_07278_),
    .X(_02583_));
 sg13g2_nor3_2 _26389_ (.A(net491),
    .B(net666),
    .C(_07277_),
    .Y(_07279_));
 sg13g2_mux2_1 _26390_ (.A0(\cpu.spi.r_mode[1][0] ),
    .A1(net911),
    .S(_07279_),
    .X(_02584_));
 sg13g2_mux2_1 _26391_ (.A0(_11966_),
    .A1(net885),
    .S(_07279_),
    .X(_02585_));
 sg13g2_nor4_2 _26392_ (.A(net550),
    .B(_09226_),
    .C(_09300_),
    .Y(_07280_),
    .D(_07073_));
 sg13g2_mux2_1 _26393_ (.A0(_12003_),
    .A1(net911),
    .S(_07280_),
    .X(_02586_));
 sg13g2_mux2_1 _26394_ (.A0(_11970_),
    .A1(net885),
    .S(_07280_),
    .X(_02587_));
 sg13g2_a21o_1 _26395_ (.A2(_11969_),
    .A1(_12003_),
    .B1(_12006_),
    .X(_07281_));
 sg13g2_buf_2 _26396_ (.A(_07281_),
    .X(_07282_));
 sg13g2_a21o_1 _26397_ (.A2(_07282_),
    .A1(_00208_),
    .B1(_07077_),
    .X(_07283_));
 sg13g2_a21oi_1 _26398_ (.A1(net828),
    .A2(_10032_),
    .Y(_07284_),
    .B1(net887));
 sg13g2_o21ai_1 _26399_ (.B1(_07284_),
    .Y(_07285_),
    .A1(net828),
    .A2(_07283_));
 sg13g2_nor2_1 _26400_ (.A(_09238_),
    .B(net887),
    .Y(_07286_));
 sg13g2_buf_2 _26401_ (.A(_07286_),
    .X(_07287_));
 sg13g2_a22oi_1 _26402_ (.Y(_07288_),
    .B1(_07287_),
    .B2(_07076_),
    .A2(_12010_),
    .A1(_09305_));
 sg13g2_nand2_1 _26403_ (.Y(_07289_),
    .A(_09357_),
    .B(_07288_));
 sg13g2_nor2_1 _26404_ (.A(_12015_),
    .B(_07289_),
    .Y(_07290_));
 sg13g2_buf_4 _26405_ (.X(_07291_),
    .A(_07290_));
 sg13g2_mux2_1 _26406_ (.A0(\cpu.spi.r_out[0] ),
    .A1(_07285_),
    .S(_07291_),
    .X(_02588_));
 sg13g2_mux2_1 _26407_ (.A0(_00208_),
    .A1(_00168_),
    .S(_07282_),
    .X(_07292_));
 sg13g2_a22oi_1 _26408_ (.Y(_07293_),
    .B1(_07287_),
    .B2(_10050_),
    .A2(net887),
    .A1(\cpu.spi.r_out[0] ));
 sg13g2_o21ai_1 _26409_ (.B1(_07293_),
    .Y(_07294_),
    .A1(net828),
    .A2(_07292_));
 sg13g2_mux2_1 _26410_ (.A0(\cpu.spi.r_out[1] ),
    .A1(_07294_),
    .S(_07291_),
    .X(_02589_));
 sg13g2_mux2_1 _26411_ (.A0(_00168_),
    .A1(_00169_),
    .S(_07282_),
    .X(_07295_));
 sg13g2_a22oi_1 _26412_ (.Y(_07296_),
    .B1(_07287_),
    .B2(net1060),
    .A2(net887),
    .A1(\cpu.spi.r_out[1] ));
 sg13g2_o21ai_1 _26413_ (.B1(_07296_),
    .Y(_07297_),
    .A1(_07236_),
    .A2(_07295_));
 sg13g2_mux2_1 _26414_ (.A0(\cpu.spi.r_out[2] ),
    .A1(_07297_),
    .S(_07291_),
    .X(_02590_));
 sg13g2_mux2_1 _26415_ (.A0(_00169_),
    .A1(_00271_),
    .S(_07282_),
    .X(_07298_));
 sg13g2_a22oi_1 _26416_ (.Y(_07299_),
    .B1(_07287_),
    .B2(net1128),
    .A2(_11994_),
    .A1(\cpu.spi.r_out[2] ));
 sg13g2_o21ai_1 _26417_ (.B1(_07299_),
    .Y(_07300_),
    .A1(net828),
    .A2(_07298_));
 sg13g2_mux2_1 _26418_ (.A0(\cpu.spi.r_out[3] ),
    .A1(_07300_),
    .S(_07291_),
    .X(_02591_));
 sg13g2_mux2_1 _26419_ (.A0(_00271_),
    .A1(_00170_),
    .S(_07282_),
    .X(_07301_));
 sg13g2_a22oi_1 _26420_ (.Y(_07302_),
    .B1(_07287_),
    .B2(_10066_),
    .A2(net887),
    .A1(\cpu.spi.r_out[3] ));
 sg13g2_o21ai_1 _26421_ (.B1(_07302_),
    .Y(_07303_),
    .A1(net828),
    .A2(_07301_));
 sg13g2_mux2_1 _26422_ (.A0(\cpu.spi.r_out[4] ),
    .A1(_07303_),
    .S(_07291_),
    .X(_02592_));
 sg13g2_mux2_1 _26423_ (.A0(_00170_),
    .A1(_00171_),
    .S(_07282_),
    .X(_07304_));
 sg13g2_a22oi_1 _26424_ (.Y(_07305_),
    .B1(_07287_),
    .B2(_10072_),
    .A2(_11994_),
    .A1(\cpu.spi.r_out[4] ));
 sg13g2_o21ai_1 _26425_ (.B1(_07305_),
    .Y(_07306_),
    .A1(net828),
    .A2(_07304_));
 sg13g2_mux2_1 _26426_ (.A0(\cpu.spi.r_out[5] ),
    .A1(_07306_),
    .S(_07291_),
    .X(_02593_));
 sg13g2_inv_1 _26427_ (.Y(_07307_),
    .A(_00172_));
 sg13g2_nand2_1 _26428_ (.Y(_07308_),
    .A(_00171_),
    .B(net672));
 sg13g2_o21ai_1 _26429_ (.B1(_07308_),
    .Y(_07309_),
    .A1(_07307_),
    .A2(net672));
 sg13g2_a22oi_1 _26430_ (.Y(_07310_),
    .B1(_07287_),
    .B2(_10078_),
    .A2(net887),
    .A1(\cpu.spi.r_out[5] ));
 sg13g2_o21ai_1 _26431_ (.B1(_07310_),
    .Y(_07311_),
    .A1(net828),
    .A2(_07309_));
 sg13g2_mux2_1 _26432_ (.A0(\cpu.spi.r_out[6] ),
    .A1(_07311_),
    .S(_07291_),
    .X(_02594_));
 sg13g2_buf_1 _26433_ (.A(_00265_),
    .X(_07312_));
 sg13g2_nor2_1 _26434_ (.A(_07312_),
    .B(net672),
    .Y(_07313_));
 sg13g2_a21oi_1 _26435_ (.A1(_07307_),
    .A2(_12008_),
    .Y(_07314_),
    .B1(_07313_));
 sg13g2_a22oi_1 _26436_ (.Y(_07315_),
    .B1(_07287_),
    .B2(_10081_),
    .A2(net887),
    .A1(\cpu.spi.r_out[6] ));
 sg13g2_o21ai_1 _26437_ (.B1(_07315_),
    .Y(_07316_),
    .A1(net828),
    .A2(_07314_));
 sg13g2_mux2_1 _26438_ (.A0(\cpu.spi.r_out[7] ),
    .A1(_07316_),
    .S(_07291_),
    .X(_02595_));
 sg13g2_nand3_1 _26439_ (.B(net928),
    .C(_09324_),
    .A(_09325_),
    .Y(_07317_));
 sg13g2_buf_1 _26440_ (.A(_07317_),
    .X(_07318_));
 sg13g2_nand2_1 _26441_ (.Y(_07319_),
    .A(net1031),
    .B(_07318_));
 sg13g2_o21ai_1 _26442_ (.B1(_07319_),
    .Y(_02598_),
    .A1(net666),
    .A2(_07318_));
 sg13g2_nand2_1 _26443_ (.Y(_07320_),
    .A(_11952_),
    .B(_07318_));
 sg13g2_o21ai_1 _26444_ (.B1(_07320_),
    .Y(_02599_),
    .A1(_02954_),
    .A2(_07318_));
 sg13g2_mux2_1 _26445_ (.A0(\cpu.spi.r_src[0] ),
    .A1(net884),
    .S(_07278_),
    .X(_02600_));
 sg13g2_mux2_1 _26446_ (.A0(\cpu.spi.r_src[1] ),
    .A1(net884),
    .S(_07279_),
    .X(_02601_));
 sg13g2_mux2_1 _26447_ (.A0(_11953_),
    .A1(net884),
    .S(_07280_),
    .X(_02602_));
 sg13g2_nand2_1 _26448_ (.Y(_07321_),
    .A(_09248_),
    .B(_05116_));
 sg13g2_buf_1 _26449_ (.A(_07321_),
    .X(_07322_));
 sg13g2_mux2_1 _26450_ (.A0(net911),
    .A1(\cpu.spi.r_timeout[0] ),
    .S(net93),
    .X(_02603_));
 sg13g2_mux2_1 _26451_ (.A0(net853),
    .A1(\cpu.spi.r_timeout[1] ),
    .S(_07322_),
    .X(_02604_));
 sg13g2_mux2_1 _26452_ (.A0(net845),
    .A1(\cpu.spi.r_timeout[2] ),
    .S(_07322_),
    .X(_02605_));
 sg13g2_mux2_1 _26453_ (.A0(net964),
    .A1(\cpu.spi.r_timeout[3] ),
    .S(net93),
    .X(_02606_));
 sg13g2_nand2_1 _26454_ (.Y(_07323_),
    .A(\cpu.spi.r_timeout[4] ),
    .B(net93));
 sg13g2_o21ai_1 _26455_ (.B1(_07323_),
    .Y(_02607_),
    .A1(net883),
    .A2(net93));
 sg13g2_nand2_1 _26456_ (.Y(_07324_),
    .A(\cpu.spi.r_timeout[5] ),
    .B(net93));
 sg13g2_o21ai_1 _26457_ (.B1(_07324_),
    .Y(_02608_),
    .A1(net882),
    .A2(net93));
 sg13g2_nand2_1 _26458_ (.Y(_07325_),
    .A(\cpu.spi.r_timeout[6] ),
    .B(_07321_));
 sg13g2_o21ai_1 _26459_ (.B1(_07325_),
    .Y(_02609_),
    .A1(net881),
    .A2(net93));
 sg13g2_mux2_1 _26460_ (.A0(net1023),
    .A1(\cpu.spi.r_timeout[7] ),
    .S(net93),
    .X(_02610_));
 sg13g2_inv_1 _26461_ (.Y(_07326_),
    .A(\cpu.spi.r_timeout_count[0] ));
 sg13g2_nor4_1 _26462_ (.A(_00211_),
    .B(_09255_),
    .C(_09276_),
    .D(net462),
    .Y(_07327_));
 sg13g2_o21ai_1 _26463_ (.B1(_09251_),
    .Y(_07328_),
    .A1(_09276_),
    .A2(_09307_));
 sg13g2_o21ai_1 _26464_ (.B1(_07328_),
    .Y(_07329_),
    .A1(_09251_),
    .A2(net1137));
 sg13g2_nor4_1 _26465_ (.A(_09316_),
    .B(_09320_),
    .C(_07327_),
    .D(_07329_),
    .Y(_07330_));
 sg13g2_buf_2 _26466_ (.A(_07330_),
    .X(_07331_));
 sg13g2_buf_1 _26467_ (.A(_07331_),
    .X(_07332_));
 sg13g2_mux2_1 _26468_ (.A0(_00268_),
    .A1(\cpu.spi.r_timeout[0] ),
    .S(net886),
    .X(_07333_));
 sg13g2_nand2_1 _26469_ (.Y(_07334_),
    .A(net33),
    .B(_07333_));
 sg13g2_o21ai_1 _26470_ (.B1(_07334_),
    .Y(_02611_),
    .A1(_07326_),
    .A2(net33));
 sg13g2_o21ai_1 _26471_ (.B1(net33),
    .Y(_07335_),
    .A1(_07326_),
    .A2(net925));
 sg13g2_nor2_1 _26472_ (.A(\cpu.spi.r_timeout_count[0] ),
    .B(\cpu.spi.r_timeout_count[1] ),
    .Y(_07336_));
 sg13g2_mux2_1 _26473_ (.A0(\cpu.spi.r_timeout[1] ),
    .A1(_07336_),
    .S(_09319_),
    .X(_07337_));
 sg13g2_a22oi_1 _26474_ (.Y(_07338_),
    .B1(_07337_),
    .B2(net33),
    .A2(_07335_),
    .A1(\cpu.spi.r_timeout_count[1] ));
 sg13g2_inv_1 _26475_ (.Y(_02612_),
    .A(_07338_));
 sg13g2_o21ai_1 _26476_ (.B1(_07331_),
    .Y(_07339_),
    .A1(net925),
    .A2(_07336_));
 sg13g2_mux2_1 _26477_ (.A0(\cpu.spi.r_timeout[2] ),
    .A1(_09256_),
    .S(_09319_),
    .X(_07340_));
 sg13g2_a22oi_1 _26478_ (.Y(_07341_),
    .B1(_07340_),
    .B2(net33),
    .A2(_07339_),
    .A1(\cpu.spi.r_timeout_count[2] ));
 sg13g2_inv_1 _26479_ (.Y(_02613_),
    .A(_07341_));
 sg13g2_o21ai_1 _26480_ (.B1(_07331_),
    .Y(_07342_),
    .A1(net925),
    .A2(_09256_));
 sg13g2_nand2b_1 _26481_ (.Y(_07343_),
    .B(_09256_),
    .A_N(\cpu.spi.r_timeout_count[3] ));
 sg13g2_nand2_1 _26482_ (.Y(_07344_),
    .A(net886),
    .B(\cpu.spi.r_timeout[3] ));
 sg13g2_o21ai_1 _26483_ (.B1(_07344_),
    .Y(_07345_),
    .A1(net925),
    .A2(_07343_));
 sg13g2_a22oi_1 _26484_ (.Y(_07346_),
    .B1(_07345_),
    .B2(net33),
    .A2(_07342_),
    .A1(\cpu.spi.r_timeout_count[3] ));
 sg13g2_inv_1 _26485_ (.Y(_02614_),
    .A(_07346_));
 sg13g2_o21ai_1 _26486_ (.B1(_07331_),
    .Y(_07347_),
    .A1(net925),
    .A2(_09257_));
 sg13g2_nand2_1 _26487_ (.Y(_07348_),
    .A(net886),
    .B(\cpu.spi.r_timeout[4] ));
 sg13g2_o21ai_1 _26488_ (.B1(_07348_),
    .Y(_07349_),
    .A1(net925),
    .A2(_09258_));
 sg13g2_a22oi_1 _26489_ (.Y(_07350_),
    .B1(_07349_),
    .B2(net33),
    .A2(_07347_),
    .A1(\cpu.spi.r_timeout_count[4] ));
 sg13g2_inv_1 _26490_ (.Y(_02615_),
    .A(_07350_));
 sg13g2_nor2_1 _26491_ (.A(\cpu.spi.r_timeout_count[4] ),
    .B(_07343_),
    .Y(_07351_));
 sg13g2_o21ai_1 _26492_ (.B1(_07331_),
    .Y(_07352_),
    .A1(net886),
    .A2(_07351_));
 sg13g2_mux2_1 _26493_ (.A0(\cpu.spi.r_timeout[5] ),
    .A1(_09259_),
    .S(_09319_),
    .X(_07353_));
 sg13g2_a22oi_1 _26494_ (.Y(_07354_),
    .B1(_07353_),
    .B2(net33),
    .A2(_07352_),
    .A1(\cpu.spi.r_timeout_count[5] ));
 sg13g2_inv_1 _26495_ (.Y(_02616_),
    .A(_07354_));
 sg13g2_o21ai_1 _26496_ (.B1(_07331_),
    .Y(_07355_),
    .A1(net886),
    .A2(_09259_));
 sg13g2_nand2_1 _26497_ (.Y(_07356_),
    .A(net886),
    .B(\cpu.spi.r_timeout[6] ));
 sg13g2_o21ai_1 _26498_ (.B1(_07356_),
    .Y(_07357_),
    .A1(net925),
    .A2(_09261_));
 sg13g2_a22oi_1 _26499_ (.Y(_07358_),
    .B1(_07357_),
    .B2(_07332_),
    .A2(_07355_),
    .A1(\cpu.spi.r_timeout_count[6] ));
 sg13g2_inv_1 _26500_ (.Y(_02617_),
    .A(_07358_));
 sg13g2_inv_1 _26501_ (.Y(_07359_),
    .A(_09261_));
 sg13g2_o21ai_1 _26502_ (.B1(_07331_),
    .Y(_07360_),
    .A1(net886),
    .A2(_07359_));
 sg13g2_nor3_1 _26503_ (.A(\cpu.spi.r_timeout_count[7] ),
    .B(net886),
    .C(_09261_),
    .Y(_07361_));
 sg13g2_a21o_1 _26504_ (.A2(\cpu.spi.r_timeout[7] ),
    .A1(net925),
    .B1(_07361_),
    .X(_07362_));
 sg13g2_a22oi_1 _26505_ (.Y(_07363_),
    .B1(_07362_),
    .B2(_07332_),
    .A2(_07360_),
    .A1(\cpu.spi.r_timeout_count[7] ));
 sg13g2_inv_1 _26506_ (.Y(_02618_),
    .A(_07363_));
 sg13g2_buf_1 _26507_ (.A(\cpu.uart.r_rcnt[0] ),
    .X(_07364_));
 sg13g2_nand2b_1 _26508_ (.Y(_07365_),
    .B(_09939_),
    .A_N(_09900_));
 sg13g2_buf_1 _26509_ (.A(_07365_),
    .X(_07366_));
 sg13g2_or3_1 _26510_ (.A(_07364_),
    .B(\cpu.uart.r_rcnt[1] ),
    .C(_07366_),
    .X(_07367_));
 sg13g2_buf_1 _26511_ (.A(_07367_),
    .X(_07368_));
 sg13g2_nor2_1 _26512_ (.A(net923),
    .B(_07368_),
    .Y(_07369_));
 sg13g2_buf_1 _26513_ (.A(\cpu.uart.r_rstate[3] ),
    .X(_07370_));
 sg13g2_buf_1 _26514_ (.A(_07370_),
    .X(_07371_));
 sg13g2_buf_1 _26515_ (.A(\cpu.uart.r_rstate[1] ),
    .X(_07372_));
 sg13g2_buf_1 _26516_ (.A(\cpu.uart.r_rstate[2] ),
    .X(_07373_));
 sg13g2_buf_1 _26517_ (.A(_07373_),
    .X(_07374_));
 sg13g2_nor2_2 _26518_ (.A(net1097),
    .B(net949),
    .Y(_07375_));
 sg13g2_buf_2 _26519_ (.A(\cpu.uart.r_rstate[0] ),
    .X(_07376_));
 sg13g2_inv_1 _26520_ (.Y(_07377_),
    .A(_07376_));
 sg13g2_nand3_1 _26521_ (.B(net950),
    .C(_07375_),
    .A(_07377_),
    .Y(_07378_));
 sg13g2_o21ai_1 _26522_ (.B1(_07378_),
    .Y(_07379_),
    .A1(net950),
    .A2(_07375_));
 sg13g2_and2_1 _26523_ (.A(_07369_),
    .B(_07379_),
    .X(_07380_));
 sg13g2_buf_2 _26524_ (.A(_07380_),
    .X(_07381_));
 sg13g2_mux2_1 _26525_ (.A0(\cpu.uart.r_ib[0] ),
    .A1(\cpu.uart.r_ib[1] ),
    .S(_07381_),
    .X(_02631_));
 sg13g2_mux2_1 _26526_ (.A0(\cpu.uart.r_ib[1] ),
    .A1(\cpu.uart.r_ib[2] ),
    .S(_07381_),
    .X(_02632_));
 sg13g2_mux2_1 _26527_ (.A0(\cpu.uart.r_ib[2] ),
    .A1(\cpu.uart.r_ib[3] ),
    .S(_07381_),
    .X(_02633_));
 sg13g2_mux2_1 _26528_ (.A0(\cpu.uart.r_ib[3] ),
    .A1(\cpu.uart.r_ib[4] ),
    .S(_07381_),
    .X(_02634_));
 sg13g2_mux2_1 _26529_ (.A0(\cpu.uart.r_ib[4] ),
    .A1(\cpu.uart.r_ib[5] ),
    .S(_07381_),
    .X(_02635_));
 sg13g2_mux2_1 _26530_ (.A0(\cpu.uart.r_ib[5] ),
    .A1(\cpu.uart.r_ib[6] ),
    .S(_07381_),
    .X(_02636_));
 sg13g2_xor2_1 _26531_ (.B(\cpu.uart.r_r ),
    .A(\cpu.uart.r_r_invert ),
    .X(_07382_));
 sg13g2_mux2_1 _26532_ (.A0(\cpu.uart.r_ib[6] ),
    .A1(_07382_),
    .S(_07381_),
    .X(_02637_));
 sg13g2_and4_1 _26533_ (.A(_07376_),
    .B(net950),
    .C(_07369_),
    .D(_07375_),
    .X(_07383_));
 sg13g2_buf_1 _26534_ (.A(_07383_),
    .X(_07384_));
 sg13g2_mux2_1 _26535_ (.A0(\cpu.uart.r_in[0] ),
    .A1(\cpu.uart.r_ib[0] ),
    .S(net129),
    .X(_02638_));
 sg13g2_mux2_1 _26536_ (.A0(\cpu.uart.r_in[1] ),
    .A1(\cpu.uart.r_ib[1] ),
    .S(net129),
    .X(_02639_));
 sg13g2_mux2_1 _26537_ (.A0(\cpu.uart.r_in[2] ),
    .A1(\cpu.uart.r_ib[2] ),
    .S(net129),
    .X(_02640_));
 sg13g2_mux2_1 _26538_ (.A0(\cpu.uart.r_in[3] ),
    .A1(\cpu.uart.r_ib[3] ),
    .S(net129),
    .X(_02641_));
 sg13g2_mux2_1 _26539_ (.A0(\cpu.uart.r_in[4] ),
    .A1(\cpu.uart.r_ib[4] ),
    .S(net129),
    .X(_02642_));
 sg13g2_mux2_1 _26540_ (.A0(\cpu.uart.r_in[5] ),
    .A1(\cpu.uart.r_ib[5] ),
    .S(net129),
    .X(_02643_));
 sg13g2_mux2_1 _26541_ (.A0(\cpu.uart.r_in[6] ),
    .A1(\cpu.uart.r_ib[6] ),
    .S(net129),
    .X(_02644_));
 sg13g2_mux2_1 _26542_ (.A0(\cpu.uart.r_in[7] ),
    .A1(_07382_),
    .S(_07384_),
    .X(_02645_));
 sg13g2_buf_2 _26543_ (.A(\cpu.uart.r_xstate[2] ),
    .X(_07385_));
 sg13g2_nor2_1 _26544_ (.A(net1139),
    .B(net1138),
    .Y(_07386_));
 sg13g2_and3_1 _26545_ (.X(_07387_),
    .A(net1030),
    .B(_07386_),
    .C(_06848_));
 sg13g2_buf_2 _26546_ (.A(_07387_),
    .X(_07388_));
 sg13g2_nand2_2 _26547_ (.Y(_07389_),
    .A(_04955_),
    .B(_07388_));
 sg13g2_buf_1 _26548_ (.A(\cpu.uart.r_xstate[1] ),
    .X(_07390_));
 sg13g2_inv_1 _26549_ (.Y(_07391_),
    .A(_07390_));
 sg13g2_buf_1 _26550_ (.A(_07391_),
    .X(_07392_));
 sg13g2_buf_1 _26551_ (.A(\cpu.uart.r_xstate[0] ),
    .X(_07393_));
 sg13g2_inv_1 _26552_ (.Y(_07394_),
    .A(_07393_));
 sg13g2_buf_2 _26553_ (.A(\cpu.uart.r_xstate[3] ),
    .X(_07395_));
 sg13g2_inv_2 _26554_ (.Y(_07396_),
    .A(_07395_));
 sg13g2_nor3_1 _26555_ (.A(net827),
    .B(_07394_),
    .C(_07396_),
    .Y(_07397_));
 sg13g2_nor2_1 _26556_ (.A(net1096),
    .B(_07389_),
    .Y(_07398_));
 sg13g2_nor3_1 _26557_ (.A(_07390_),
    .B(_07395_),
    .C(_07398_),
    .Y(_07399_));
 sg13g2_a21oi_1 _26558_ (.A1(_07389_),
    .A2(_07397_),
    .Y(_07400_),
    .B1(_07399_));
 sg13g2_buf_1 _26559_ (.A(\cpu.uart.r_xcnt[0] ),
    .X(_07401_));
 sg13g2_nor2_1 _26560_ (.A(_07401_),
    .B(\cpu.uart.r_xcnt[1] ),
    .Y(_07402_));
 sg13g2_nand2_1 _26561_ (.Y(_07403_),
    .A(_09911_),
    .B(_07402_));
 sg13g2_a21oi_1 _26562_ (.A1(_07395_),
    .A2(_07403_),
    .Y(_07404_),
    .B1(_07390_));
 sg13g2_inv_1 _26563_ (.Y(_07405_),
    .A(_07385_));
 sg13g2_o21ai_1 _26564_ (.B1(_07405_),
    .Y(_07406_),
    .A1(_07397_),
    .A2(_07404_));
 sg13g2_and2_1 _26565_ (.A(_09911_),
    .B(_07402_),
    .X(_07407_));
 sg13g2_buf_1 _26566_ (.A(_07407_),
    .X(_07408_));
 sg13g2_nand2_1 _26567_ (.Y(_07409_),
    .A(_07396_),
    .B(_07408_));
 sg13g2_a21oi_1 _26568_ (.A1(_07406_),
    .A2(_07409_),
    .Y(_07410_),
    .B1(_09316_));
 sg13g2_o21ai_1 _26569_ (.B1(_07410_),
    .Y(_07411_),
    .A1(_07385_),
    .A2(_07400_));
 sg13g2_buf_2 _26570_ (.A(_07411_),
    .X(_07412_));
 sg13g2_buf_1 _26571_ (.A(_07412_),
    .X(_07413_));
 sg13g2_nor2_1 _26572_ (.A(_07385_),
    .B(_07395_),
    .Y(_07414_));
 sg13g2_a21oi_1 _26573_ (.A1(net827),
    .A2(_07405_),
    .Y(_07415_),
    .B1(_07396_));
 sg13g2_a21oi_1 _26574_ (.A1(net827),
    .A2(_07414_),
    .Y(_07416_),
    .B1(_07415_));
 sg13g2_buf_2 _26575_ (.A(_07416_),
    .X(_07417_));
 sg13g2_buf_1 _26576_ (.A(_07417_),
    .X(_07418_));
 sg13g2_nor2b_1 _26577_ (.A(_07417_),
    .B_N(_10032_),
    .Y(_07419_));
 sg13g2_a21oi_1 _26578_ (.A1(\cpu.uart.r_out[1] ),
    .A2(net523),
    .Y(_07420_),
    .B1(_07419_));
 sg13g2_nand2_1 _26579_ (.Y(_07421_),
    .A(\cpu.uart.r_out[0] ),
    .B(net29));
 sg13g2_o21ai_1 _26580_ (.B1(_07421_),
    .Y(_02646_),
    .A1(net29),
    .A2(_07420_));
 sg13g2_nor2b_1 _26581_ (.A(_07417_),
    .B_N(_10050_),
    .Y(_07422_));
 sg13g2_a21oi_1 _26582_ (.A1(\cpu.uart.r_out[2] ),
    .A2(net523),
    .Y(_07423_),
    .B1(_07422_));
 sg13g2_nand2_1 _26583_ (.Y(_07424_),
    .A(\cpu.uart.r_out[1] ),
    .B(net29));
 sg13g2_o21ai_1 _26584_ (.B1(_07424_),
    .Y(_02647_),
    .A1(net29),
    .A2(_07423_));
 sg13g2_nor2b_1 _26585_ (.A(_07417_),
    .B_N(_10055_),
    .Y(_07425_));
 sg13g2_a21oi_1 _26586_ (.A1(\cpu.uart.r_out[3] ),
    .A2(net523),
    .Y(_07426_),
    .B1(_07425_));
 sg13g2_nand2_1 _26587_ (.Y(_07427_),
    .A(\cpu.uart.r_out[2] ),
    .B(_07412_));
 sg13g2_o21ai_1 _26588_ (.B1(_07427_),
    .Y(_02648_),
    .A1(net29),
    .A2(_07426_));
 sg13g2_nor2b_1 _26589_ (.A(_07417_),
    .B_N(_10060_),
    .Y(_07428_));
 sg13g2_a21oi_1 _26590_ (.A1(\cpu.uart.r_out[4] ),
    .A2(net523),
    .Y(_07429_),
    .B1(_07428_));
 sg13g2_nand2_1 _26591_ (.Y(_07430_),
    .A(\cpu.uart.r_out[3] ),
    .B(_07412_));
 sg13g2_o21ai_1 _26592_ (.B1(_07430_),
    .Y(_02649_),
    .A1(net29),
    .A2(_07429_));
 sg13g2_nor2_1 _26593_ (.A(_12136_),
    .B(_07418_),
    .Y(_07431_));
 sg13g2_a21oi_1 _26594_ (.A1(\cpu.uart.r_out[5] ),
    .A2(_07418_),
    .Y(_07432_),
    .B1(_07431_));
 sg13g2_nand2_1 _26595_ (.Y(_07433_),
    .A(\cpu.uart.r_out[4] ),
    .B(_07412_));
 sg13g2_o21ai_1 _26596_ (.B1(_07433_),
    .Y(_02650_),
    .A1(_07413_),
    .A2(_07432_));
 sg13g2_nor2_1 _26597_ (.A(_12144_),
    .B(net523),
    .Y(_07434_));
 sg13g2_a21oi_1 _26598_ (.A1(\cpu.uart.r_out[6] ),
    .A2(net523),
    .Y(_07435_),
    .B1(_07434_));
 sg13g2_nand2_1 _26599_ (.Y(_07436_),
    .A(\cpu.uart.r_out[5] ),
    .B(_07412_));
 sg13g2_o21ai_1 _26600_ (.B1(_07436_),
    .Y(_02651_),
    .A1(_07413_),
    .A2(_07435_));
 sg13g2_nor2_1 _26601_ (.A(_12149_),
    .B(_07417_),
    .Y(_07437_));
 sg13g2_a21oi_1 _26602_ (.A1(\cpu.uart.r_out[7] ),
    .A2(net523),
    .Y(_07438_),
    .B1(_07437_));
 sg13g2_nand2_1 _26603_ (.Y(_07439_),
    .A(\cpu.uart.r_out[6] ),
    .B(_07412_));
 sg13g2_o21ai_1 _26604_ (.B1(_07439_),
    .Y(_02652_),
    .A1(net29),
    .A2(_07438_));
 sg13g2_nor3_1 _26605_ (.A(_07312_),
    .B(_07412_),
    .C(net523),
    .Y(_07440_));
 sg13g2_a21o_1 _26606_ (.A2(net29),
    .A1(\cpu.uart.r_out[7] ),
    .B1(_07440_),
    .X(_02653_));
 sg13g2_nor3_1 _26607_ (.A(net1097),
    .B(_07373_),
    .C(net1098),
    .Y(_07441_));
 sg13g2_a22oi_1 _26608_ (.Y(_07442_),
    .B1(_07366_),
    .B2(_07441_),
    .A2(net1098),
    .A1(net1097));
 sg13g2_nor4_1 _26609_ (.A(_07376_),
    .B(\cpu.uart.r_rstate[1] ),
    .C(_07373_),
    .D(net1098),
    .Y(_07443_));
 sg13g2_a21o_1 _26610_ (.A2(_07366_),
    .A1(net1097),
    .B1(_07373_),
    .X(_07444_));
 sg13g2_a22oi_1 _26611_ (.Y(_07445_),
    .B1(_07444_),
    .B2(net1098),
    .A2(_07443_),
    .A1(_07382_));
 sg13g2_o21ai_1 _26612_ (.B1(_07445_),
    .Y(_07446_),
    .A1(_07377_),
    .A2(_07442_));
 sg13g2_nor2_1 _26613_ (.A(_07377_),
    .B(_07372_),
    .Y(_07447_));
 sg13g2_nor2b_1 _26614_ (.A(net1098),
    .B_N(_07382_),
    .Y(_07448_));
 sg13g2_nand2_1 _26615_ (.Y(_07449_),
    .A(net1097),
    .B(net1098));
 sg13g2_nor2_1 _26616_ (.A(_07376_),
    .B(_07449_),
    .Y(_07450_));
 sg13g2_a21oi_1 _26617_ (.A1(_07447_),
    .A2(_07448_),
    .Y(_07451_),
    .B1(_07450_));
 sg13g2_nor3_1 _26618_ (.A(net949),
    .B(_07368_),
    .C(_07451_),
    .Y(_07452_));
 sg13g2_xor2_1 _26619_ (.B(_07375_),
    .A(net950),
    .X(_07453_));
 sg13g2_o21ai_1 _26620_ (.B1(net928),
    .Y(_07454_),
    .A1(_09911_),
    .A2(_07453_));
 sg13g2_nor3_2 _26621_ (.A(_07446_),
    .B(_07452_),
    .C(_07454_),
    .Y(_07455_));
 sg13g2_and2_1 _26622_ (.A(_07376_),
    .B(net1097),
    .X(_07456_));
 sg13g2_buf_1 _26623_ (.A(_07456_),
    .X(_07457_));
 sg13g2_o21ai_1 _26624_ (.B1(_07371_),
    .Y(_07458_),
    .A1(net949),
    .A2(_07457_));
 sg13g2_nor2b_1 _26625_ (.A(_07443_),
    .B_N(_07458_),
    .Y(_07459_));
 sg13g2_nand3_1 _26626_ (.B(_07455_),
    .C(_07459_),
    .A(_07364_),
    .Y(_07460_));
 sg13g2_o21ai_1 _26627_ (.B1(_07460_),
    .Y(_07461_),
    .A1(_07364_),
    .A2(_07455_));
 sg13g2_inv_1 _26628_ (.Y(_02656_),
    .A(_07461_));
 sg13g2_nand3b_1 _26629_ (.B(_07455_),
    .C(_07459_),
    .Y(_07462_),
    .A_N(_07364_));
 sg13g2_nand2_1 _26630_ (.Y(_07463_),
    .A(_07364_),
    .B(_07459_));
 sg13g2_nand2_1 _26631_ (.Y(_07464_),
    .A(_07455_),
    .B(_07463_));
 sg13g2_nand2_1 _26632_ (.Y(_07465_),
    .A(\cpu.uart.r_rcnt[1] ),
    .B(_07464_));
 sg13g2_o21ai_1 _26633_ (.B1(_07465_),
    .Y(_02657_),
    .A1(\cpu.uart.r_rcnt[1] ),
    .A2(_07462_));
 sg13g2_nand2_1 _26634_ (.Y(_07466_),
    .A(\cpu.uart.r_out[0] ),
    .B(_07417_));
 sg13g2_xnor2_1 _26635_ (.Y(_07467_),
    .A(\cpu.uart.r_x_invert ),
    .B(_07466_));
 sg13g2_nand2_1 _26636_ (.Y(_07468_),
    .A(_07405_),
    .B(_07396_));
 sg13g2_nand2_1 _26637_ (.Y(_07469_),
    .A(_07385_),
    .B(_07395_));
 sg13g2_buf_1 _26638_ (.A(_07469_),
    .X(_07470_));
 sg13g2_a21oi_1 _26639_ (.A1(_07468_),
    .A2(_07470_),
    .Y(_07471_),
    .B1(_07393_));
 sg13g2_nand2_1 _26640_ (.Y(_07472_),
    .A(net827),
    .B(_07471_));
 sg13g2_nor2_1 _26641_ (.A(_07385_),
    .B(_07396_),
    .Y(_07473_));
 sg13g2_nand2_1 _26642_ (.Y(_07474_),
    .A(_07390_),
    .B(_07473_));
 sg13g2_nand3_1 _26643_ (.B(_07472_),
    .C(_07474_),
    .A(net803),
    .Y(_07475_));
 sg13g2_mux2_1 _26644_ (.A0(_07467_),
    .A1(_00264_),
    .S(_07475_),
    .X(_07476_));
 sg13g2_buf_1 _26645_ (.A(\cpu.gpio.genblk1[3].srcs_o[1] ),
    .X(_07477_));
 sg13g2_nor2_2 _26646_ (.A(net827),
    .B(_07394_),
    .Y(_07478_));
 sg13g2_nand2_2 _26647_ (.Y(_07479_),
    .A(_07478_),
    .B(_07473_));
 sg13g2_nor2_2 _26648_ (.A(_07389_),
    .B(_07479_),
    .Y(_07480_));
 sg13g2_inv_1 _26649_ (.Y(_07481_),
    .A(_07480_));
 sg13g2_nor2_1 _26650_ (.A(_07366_),
    .B(_07468_),
    .Y(_07482_));
 sg13g2_nor2_1 _26651_ (.A(_07471_),
    .B(_07482_),
    .Y(_07483_));
 sg13g2_nand2b_1 _26652_ (.Y(_07484_),
    .B(_07403_),
    .A_N(_07397_));
 sg13g2_a22oi_1 _26653_ (.Y(_07485_),
    .B1(_07484_),
    .B2(_07405_),
    .A2(_07408_),
    .A1(_07396_));
 sg13g2_o21ai_1 _26654_ (.B1(_07485_),
    .Y(_07486_),
    .A1(_07390_),
    .A2(_07483_));
 sg13g2_a21oi_1 _26655_ (.A1(_07481_),
    .A2(_07486_),
    .Y(_07487_),
    .B1(net923));
 sg13g2_mux2_1 _26656_ (.A0(_07476_),
    .A1(_07477_),
    .S(_07487_),
    .X(_02662_));
 sg13g2_a21oi_1 _26657_ (.A1(net1096),
    .A2(_07402_),
    .Y(_07488_),
    .B1(_07385_));
 sg13g2_o21ai_1 _26658_ (.B1(_07385_),
    .Y(_07489_),
    .A1(net1096),
    .A2(_07402_));
 sg13g2_o21ai_1 _26659_ (.B1(_07489_),
    .Y(_07490_),
    .A1(net827),
    .A2(_07488_));
 sg13g2_nand2_1 _26660_ (.Y(_07491_),
    .A(_07395_),
    .B(_07490_));
 sg13g2_nor2_1 _26661_ (.A(_07390_),
    .B(net1096),
    .Y(_07492_));
 sg13g2_nand2_1 _26662_ (.Y(_07493_),
    .A(_07414_),
    .B(_07492_));
 sg13g2_nand4_1 _26663_ (.B(_09911_),
    .C(_07491_),
    .A(net928),
    .Y(_07494_),
    .D(_07493_));
 sg13g2_nor2_1 _26664_ (.A(_07480_),
    .B(_07494_),
    .Y(_07495_));
 sg13g2_nor2_1 _26665_ (.A(_07470_),
    .B(_07492_),
    .Y(_07496_));
 sg13g2_a21oi_1 _26666_ (.A1(net827),
    .A2(_07414_),
    .Y(_07497_),
    .B1(_07496_));
 sg13g2_nand2_1 _26667_ (.Y(_07498_),
    .A(_07495_),
    .B(_07497_));
 sg13g2_nor3_1 _26668_ (.A(_07401_),
    .B(_07480_),
    .C(_07494_),
    .Y(_07499_));
 sg13g2_a21oi_1 _26669_ (.A1(_07401_),
    .A2(_07498_),
    .Y(_07500_),
    .B1(_07499_));
 sg13g2_inv_1 _26670_ (.Y(_02665_),
    .A(_07500_));
 sg13g2_nand2_1 _26671_ (.Y(_07501_),
    .A(_07401_),
    .B(_07497_));
 sg13g2_nand2_1 _26672_ (.Y(_07502_),
    .A(_07495_),
    .B(_07501_));
 sg13g2_o21ai_1 _26673_ (.B1(\cpu.uart.r_xcnt[1] ),
    .Y(_07503_),
    .A1(_07401_),
    .A2(_07498_));
 sg13g2_o21ai_1 _26674_ (.B1(_07503_),
    .Y(_02666_),
    .A1(\cpu.uart.r_xcnt[1] ),
    .A2(_07502_));
 sg13g2_nor3_1 _26675_ (.A(_09246_),
    .B(net684),
    .C(_09951_),
    .Y(_07504_));
 sg13g2_buf_1 _26676_ (.A(_07504_),
    .X(_07505_));
 sg13g2_buf_1 _26677_ (.A(_07505_),
    .X(_07506_));
 sg13g2_nand3_1 _26678_ (.B(_10179_),
    .C(_10184_),
    .A(_10173_),
    .Y(_07507_));
 sg13g2_nor3_2 _26679_ (.A(_10148_),
    .B(_10175_),
    .C(_07507_),
    .Y(_07508_));
 sg13g2_nand2_1 _26680_ (.Y(_07509_),
    .A(_09953_),
    .B(_10095_));
 sg13g2_buf_1 _26681_ (.A(_07509_),
    .X(_07510_));
 sg13g2_o21ai_1 _26682_ (.B1(net92),
    .Y(_07511_),
    .A1(net102),
    .A2(_07508_));
 sg13g2_nand2_1 _26683_ (.Y(_07512_),
    .A(_04945_),
    .B(_07511_));
 sg13g2_buf_1 _26684_ (.A(_10118_),
    .X(_07513_));
 sg13g2_nor2b_1 _26685_ (.A(_04945_),
    .B_N(_07508_),
    .Y(_07514_));
 sg13g2_a22oi_1 _26686_ (.Y(_07515_),
    .B1(_07514_),
    .B2(net90),
    .A2(net83),
    .A1(net1062));
 sg13g2_nand2_1 _26687_ (.Y(_02452_),
    .A(_07512_),
    .B(_07515_));
 sg13g2_a21o_1 _26688_ (.A2(_07508_),
    .A1(_04945_),
    .B1(_07505_),
    .X(_07516_));
 sg13g2_a21oi_1 _26689_ (.A1(net92),
    .A2(_07516_),
    .Y(_07517_),
    .B1(_05384_));
 sg13g2_nand2_1 _26690_ (.Y(_07518_),
    .A(net103),
    .B(net362));
 sg13g2_buf_1 _26691_ (.A(_07518_),
    .X(_07519_));
 sg13g2_nor2_1 _26692_ (.A(net1061),
    .B(_07519_),
    .Y(_07520_));
 sg13g2_nand3_1 _26693_ (.B(_05384_),
    .C(_07508_),
    .A(_04945_),
    .Y(_07521_));
 sg13g2_nor2_1 _26694_ (.A(_07505_),
    .B(_07521_),
    .Y(_07522_));
 sg13g2_nor3_1 _26695_ (.A(_07517_),
    .B(_07520_),
    .C(_07522_),
    .Y(_02453_));
 sg13g2_a21oi_1 _26696_ (.A1(_10089_),
    .A2(_07521_),
    .Y(_07523_),
    .B1(_10097_));
 sg13g2_nor2_1 _26697_ (.A(_05433_),
    .B(_07522_),
    .Y(_07524_));
 sg13g2_a21oi_1 _26698_ (.A1(_05433_),
    .A2(_07523_),
    .Y(_07525_),
    .B1(_07524_));
 sg13g2_a21o_1 _26699_ (.A2(net83),
    .A1(net845),
    .B1(_07525_),
    .X(_02454_));
 sg13g2_inv_1 _26700_ (.Y(_07526_),
    .A(_05506_));
 sg13g2_nand3_1 _26701_ (.B(_05384_),
    .C(_05433_),
    .A(_04945_),
    .Y(_07527_));
 sg13g2_nor2_1 _26702_ (.A(_07507_),
    .B(_07527_),
    .Y(_07528_));
 sg13g2_and2_1 _26703_ (.A(_10176_),
    .B(_07528_),
    .X(_07529_));
 sg13g2_buf_1 _26704_ (.A(_07529_),
    .X(_07530_));
 sg13g2_o21ai_1 _26705_ (.B1(net92),
    .Y(_07531_),
    .A1(net102),
    .A2(_07530_));
 sg13g2_nand3_1 _26706_ (.B(net90),
    .C(_07530_),
    .A(_05506_),
    .Y(_07532_));
 sg13g2_o21ai_1 _26707_ (.B1(_07532_),
    .Y(_07533_),
    .A1(net954),
    .A2(_07519_));
 sg13g2_a21oi_1 _26708_ (.A1(_07526_),
    .A2(_07531_),
    .Y(_02455_),
    .B1(_07533_));
 sg13g2_and3_1 _26709_ (.X(_07534_),
    .A(_05506_),
    .B(_10180_),
    .C(_07528_));
 sg13g2_buf_1 _26710_ (.A(_07534_),
    .X(_07535_));
 sg13g2_o21ai_1 _26711_ (.B1(net92),
    .Y(_07536_),
    .A1(net102),
    .A2(_07535_));
 sg13g2_nor2b_1 _26712_ (.A(_05541_),
    .B_N(_07535_),
    .Y(_07537_));
 sg13g2_a22oi_1 _26713_ (.Y(_07538_),
    .B1(_07537_),
    .B2(net90),
    .A2(_07536_),
    .A1(_05541_));
 sg13g2_o21ai_1 _26714_ (.B1(_07538_),
    .Y(_02456_),
    .A1(net883),
    .A2(_07519_));
 sg13g2_buf_1 _26715_ (.A(_10089_),
    .X(_07539_));
 sg13g2_nand3_1 _26716_ (.B(_05541_),
    .C(_07530_),
    .A(_05506_),
    .Y(_07540_));
 sg13g2_buf_1 _26717_ (.A(_07540_),
    .X(_07541_));
 sg13g2_a21oi_1 _26718_ (.A1(_07539_),
    .A2(_07541_),
    .Y(_07542_),
    .B1(net88));
 sg13g2_nand2b_1 _26719_ (.Y(_07543_),
    .B(_07542_),
    .A_N(_05634_));
 sg13g2_o21ai_1 _26720_ (.B1(_05634_),
    .Y(_07544_),
    .A1(net102),
    .A2(_07541_));
 sg13g2_a22oi_1 _26721_ (.Y(_02457_),
    .B1(_07543_),
    .B2(_07544_),
    .A2(_07513_),
    .A1(net876));
 sg13g2_and3_1 _26722_ (.X(_07545_),
    .A(_05541_),
    .B(_05634_),
    .C(_07535_));
 sg13g2_o21ai_1 _26723_ (.B1(_07510_),
    .Y(_07546_),
    .A1(_07505_),
    .A2(_07545_));
 sg13g2_nor2b_1 _26724_ (.A(_05702_),
    .B_N(_07545_),
    .Y(_07547_));
 sg13g2_a22oi_1 _26725_ (.Y(_07548_),
    .B1(_07547_),
    .B2(_10090_),
    .A2(_07546_),
    .A1(_05702_));
 sg13g2_o21ai_1 _26726_ (.B1(_07548_),
    .Y(_02458_),
    .A1(net881),
    .A2(_07519_));
 sg13g2_nand2_1 _26727_ (.Y(_07549_),
    .A(_05634_),
    .B(_05702_));
 sg13g2_nor2_1 _26728_ (.A(_07541_),
    .B(_07549_),
    .Y(_07550_));
 sg13g2_o21ai_1 _26729_ (.B1(net92),
    .Y(_07551_),
    .A1(_07506_),
    .A2(_07550_));
 sg13g2_nor4_1 _26730_ (.A(_05110_),
    .B(_07506_),
    .C(_07541_),
    .D(_07549_),
    .Y(_07552_));
 sg13g2_a221oi_1 _26731_ (.B2(_05110_),
    .C1(_07552_),
    .B1(_07551_),
    .A1(net1053),
    .Y(_07553_),
    .A2(_07513_));
 sg13g2_inv_1 _26732_ (.Y(_02459_),
    .A(_07553_));
 sg13g2_nand2_1 _26733_ (.Y(_07554_),
    .A(_05541_),
    .B(_07535_));
 sg13g2_nand3_1 _26734_ (.B(_05702_),
    .C(_05110_),
    .A(_05634_),
    .Y(_07555_));
 sg13g2_o21ai_1 _26735_ (.B1(_07539_),
    .Y(_07556_),
    .A1(_07554_),
    .A2(_07555_));
 sg13g2_a21oi_1 _26736_ (.A1(net92),
    .A2(_07556_),
    .Y(_07557_),
    .B1(_05752_));
 sg13g2_inv_1 _26737_ (.Y(_07558_),
    .A(_05752_));
 sg13g2_nor2_1 _26738_ (.A(_07558_),
    .B(_07555_),
    .Y(_07559_));
 sg13g2_nor2b_1 _26739_ (.A(_07554_),
    .B_N(_07559_),
    .Y(_07560_));
 sg13g2_nand2_1 _26740_ (.Y(_07561_),
    .A(net82),
    .B(_07560_));
 sg13g2_o21ai_1 _26741_ (.B1(_07561_),
    .Y(_07562_),
    .A1(_10146_),
    .A2(_07519_));
 sg13g2_nor2_1 _26742_ (.A(_07557_),
    .B(_07562_),
    .Y(_02460_));
 sg13g2_o21ai_1 _26743_ (.B1(net92),
    .Y(_07563_),
    .A1(_07505_),
    .A2(_07560_));
 sg13g2_nor2_1 _26744_ (.A(_05767_),
    .B(_07563_),
    .Y(_07564_));
 sg13g2_a21oi_1 _26745_ (.A1(_05767_),
    .A2(_07561_),
    .Y(_07565_),
    .B1(_07564_));
 sg13g2_a21oi_1 _26746_ (.A1(_12170_),
    .A2(net83),
    .Y(_02461_),
    .B1(_07565_));
 sg13g2_nand2_1 _26747_ (.Y(_07566_),
    .A(_05767_),
    .B(_07560_));
 sg13g2_a21oi_1 _26748_ (.A1(net82),
    .A2(_07566_),
    .Y(_07567_),
    .B1(net88));
 sg13g2_nand2b_1 _26749_ (.Y(_07568_),
    .B(_07567_),
    .A_N(_05152_));
 sg13g2_o21ai_1 _26750_ (.B1(_05152_),
    .Y(_07569_),
    .A1(net102),
    .A2(_07566_));
 sg13g2_a22oi_1 _26751_ (.Y(_02462_),
    .B1(_07568_),
    .B2(_07569_),
    .A2(net83),
    .A1(_12066_));
 sg13g2_inv_1 _26752_ (.Y(_07570_),
    .A(_05196_));
 sg13g2_nand3_1 _26753_ (.B(_05152_),
    .C(_07559_),
    .A(_05767_),
    .Y(_07571_));
 sg13g2_nor2_1 _26754_ (.A(_07541_),
    .B(_07571_),
    .Y(_07572_));
 sg13g2_o21ai_1 _26755_ (.B1(net92),
    .Y(_07573_),
    .A1(net102),
    .A2(_07572_));
 sg13g2_nand3_1 _26756_ (.B(net90),
    .C(_07572_),
    .A(_05196_),
    .Y(_07574_));
 sg13g2_o21ai_1 _26757_ (.B1(_07574_),
    .Y(_07575_),
    .A1(_10162_),
    .A2(_07519_));
 sg13g2_a21oi_1 _26758_ (.A1(_07570_),
    .A2(_07573_),
    .Y(_02463_),
    .B1(_07575_));
 sg13g2_nand4_1 _26759_ (.B(_05152_),
    .C(_05196_),
    .A(_05767_),
    .Y(_07576_),
    .D(_07560_));
 sg13g2_a21oi_1 _26760_ (.A1(net82),
    .A2(_07576_),
    .Y(_07577_),
    .B1(_10097_));
 sg13g2_inv_1 _26761_ (.Y(_07578_),
    .A(_07576_));
 sg13g2_nand3_1 _26762_ (.B(net82),
    .C(_07578_),
    .A(_05208_),
    .Y(_07579_));
 sg13g2_o21ai_1 _26763_ (.B1(_07579_),
    .Y(_07580_),
    .A1(_05208_),
    .A2(_07577_));
 sg13g2_a21oi_1 _26764_ (.A1(_12093_),
    .A2(net83),
    .Y(_02464_),
    .B1(_07580_));
 sg13g2_nand3_1 _26765_ (.B(_05208_),
    .C(_07572_),
    .A(_05196_),
    .Y(_07581_));
 sg13g2_a21oi_1 _26766_ (.A1(net82),
    .A2(_07581_),
    .Y(_07582_),
    .B1(_10097_));
 sg13g2_inv_1 _26767_ (.Y(_07583_),
    .A(_07581_));
 sg13g2_nand3_1 _26768_ (.B(net82),
    .C(_07583_),
    .A(_05239_),
    .Y(_07584_));
 sg13g2_o21ai_1 _26769_ (.B1(_07584_),
    .Y(_07585_),
    .A1(_05239_),
    .A2(_07582_));
 sg13g2_a21oi_1 _26770_ (.A1(_12101_),
    .A2(net83),
    .Y(_02465_),
    .B1(_07585_));
 sg13g2_nand3_1 _26771_ (.B(_05239_),
    .C(_07578_),
    .A(_05208_),
    .Y(_07586_));
 sg13g2_a21oi_1 _26772_ (.A1(net82),
    .A2(_07586_),
    .Y(_07587_),
    .B1(net88));
 sg13g2_nand2b_1 _26773_ (.Y(_07588_),
    .B(_07587_),
    .A_N(_05268_));
 sg13g2_o21ai_1 _26774_ (.B1(_05268_),
    .Y(_07589_),
    .A1(net102),
    .A2(_07586_));
 sg13g2_a22oi_1 _26775_ (.Y(_02466_),
    .B1(_07588_),
    .B2(_07589_),
    .A2(net83),
    .A1(_12107_));
 sg13g2_nand3_1 _26776_ (.B(_05268_),
    .C(_07583_),
    .A(_05239_),
    .Y(_07590_));
 sg13g2_a21oi_1 _26777_ (.A1(net82),
    .A2(_07590_),
    .Y(_07591_),
    .B1(net88));
 sg13g2_nand2b_1 _26778_ (.Y(_07592_),
    .B(_07591_),
    .A_N(_05301_));
 sg13g2_o21ai_1 _26779_ (.B1(_05301_),
    .Y(_07593_),
    .A1(net102),
    .A2(_07590_));
 sg13g2_a22oi_1 _26780_ (.Y(_02467_),
    .B1(_07592_),
    .B2(_07593_),
    .A2(net83),
    .A1(_12113_));
 sg13g2_nor2_1 _26781_ (.A(\cpu.r_clk_invert ),
    .B(net800),
    .Y(_07594_));
 sg13g2_a21oi_1 _26782_ (.A1(_09186_),
    .A2(_09876_),
    .Y(_02534_),
    .B1(_07594_));
 sg13g2_inv_1 _26783_ (.Y(_07595_),
    .A(\cpu.dcache.r_valid[0] ));
 sg13g2_nand4_1 _26784_ (.B(_02934_),
    .C(_02939_),
    .A(_09361_),
    .Y(_07596_),
    .D(_02941_));
 sg13g2_buf_2 _26785_ (.A(_07596_),
    .X(_07597_));
 sg13g2_inv_1 _26786_ (.Y(_07598_),
    .A(_07597_));
 sg13g2_nand2b_1 _26787_ (.Y(_07599_),
    .B(_09157_),
    .A_N(\cpu.d_flush_all ));
 sg13g2_buf_2 _26788_ (.A(_07599_),
    .X(_07600_));
 sg13g2_a221oi_1 _26789_ (.B2(_12045_),
    .C1(_07600_),
    .B1(_07598_),
    .A1(_07595_),
    .Y(_00729_),
    .A2(net555));
 sg13g2_nor2_1 _26790_ (.A(\cpu.dcache.r_valid[1] ),
    .B(net496),
    .Y(_07601_));
 sg13g2_nor2_1 _26791_ (.A(_12207_),
    .B(_07597_),
    .Y(_07602_));
 sg13g2_nor3_1 _26792_ (.A(_07600_),
    .B(_07601_),
    .C(_07602_),
    .Y(_00730_));
 sg13g2_nor2_1 _26793_ (.A(\cpu.dcache.r_valid[2] ),
    .B(net501),
    .Y(_07603_));
 sg13g2_nor2_1 _26794_ (.A(net669),
    .B(_07597_),
    .Y(_07604_));
 sg13g2_nor3_1 _26795_ (.A(_07600_),
    .B(_07603_),
    .C(_07604_),
    .Y(_00731_));
 sg13g2_nor2_1 _26796_ (.A(\cpu.dcache.r_valid[3] ),
    .B(net273),
    .Y(_07605_));
 sg13g2_nor2_1 _26797_ (.A(_12477_),
    .B(_07597_),
    .Y(_07606_));
 sg13g2_nor3_1 _26798_ (.A(_07600_),
    .B(_07605_),
    .C(_07606_),
    .Y(_00732_));
 sg13g2_inv_1 _26799_ (.Y(_07607_),
    .A(\cpu.dcache.r_valid[4] ));
 sg13g2_a221oi_1 _26800_ (.B2(_10087_),
    .C1(_07600_),
    .B1(_07598_),
    .A1(_07607_),
    .Y(_00733_),
    .A2(net414));
 sg13g2_nor2_1 _26801_ (.A(\cpu.dcache.r_valid[5] ),
    .B(net356),
    .Y(_07608_));
 sg13g2_nor2_1 _26802_ (.A(net500),
    .B(_07597_),
    .Y(_07609_));
 sg13g2_nor3_1 _26803_ (.A(_07600_),
    .B(_07608_),
    .C(_07609_),
    .Y(_00734_));
 sg13g2_nor2_1 _26804_ (.A(\cpu.dcache.r_valid[6] ),
    .B(net354),
    .Y(_07610_));
 sg13g2_nor2_1 _26805_ (.A(net498),
    .B(_07597_),
    .Y(_07611_));
 sg13g2_nor3_1 _26806_ (.A(_07600_),
    .B(_07610_),
    .C(_07611_),
    .Y(_00735_));
 sg13g2_nor2_1 _26807_ (.A(\cpu.dcache.r_valid[7] ),
    .B(net411),
    .Y(_07612_));
 sg13g2_nor2_1 _26808_ (.A(_10044_),
    .B(_07597_),
    .Y(_07613_));
 sg13g2_nor3_1 _26809_ (.A(_07600_),
    .B(_07612_),
    .C(_07613_),
    .Y(_00736_));
 sg13g2_nor3_1 _26810_ (.A(net1125),
    .B(net1124),
    .C(_10194_),
    .Y(_07614_));
 sg13g2_nand2_1 _26811_ (.Y(_07615_),
    .A(_04788_),
    .B(_07614_));
 sg13g2_buf_1 _26812_ (.A(_07615_),
    .X(_07616_));
 sg13g2_nand2_1 _26813_ (.Y(_07617_),
    .A(_08347_),
    .B(net522));
 sg13g2_o21ai_1 _26814_ (.B1(_07617_),
    .Y(_07618_),
    .A1(_03838_),
    .A2(net522));
 sg13g2_inv_1 _26815_ (.Y(_07619_),
    .A(_07618_));
 sg13g2_nor3_1 _26816_ (.A(net270),
    .B(_09318_),
    .C(_07619_),
    .Y(_00784_));
 sg13g2_and4_1 _26817_ (.A(net994),
    .B(_10651_),
    .C(\cpu.dec.do_flush_all ),
    .D(_03950_),
    .X(_00917_));
 sg13g2_and4_1 _26818_ (.A(net994),
    .B(_10645_),
    .C(\cpu.dec.do_flush_all ),
    .D(net665),
    .X(_00935_));
 sg13g2_nand4_1 _26819_ (.B(_04096_),
    .C(net665),
    .A(net994),
    .Y(_07620_),
    .D(_10932_));
 sg13g2_mux2_1 _26820_ (.A0(_10625_),
    .A1(_09160_),
    .S(_07620_),
    .X(_07621_));
 sg13g2_nand2_1 _26821_ (.Y(_07622_),
    .A(net522),
    .B(_07621_));
 sg13g2_o21ai_1 _26822_ (.B1(_07622_),
    .Y(_07623_),
    .A1(_11056_),
    .A2(_07616_));
 sg13g2_nand3_1 _26823_ (.B(_11466_),
    .C(_07623_),
    .A(_09158_),
    .Y(_07624_));
 sg13g2_a21oi_1 _26824_ (.A1(net665),
    .A2(net153),
    .Y(_00936_),
    .B1(_07624_));
 sg13g2_nor3_1 _26825_ (.A(_00294_),
    .B(_09244_),
    .C(_11475_),
    .Y(_07625_));
 sg13g2_o21ai_1 _26826_ (.B1(_07625_),
    .Y(_07626_),
    .A1(_00282_),
    .A2(_05035_));
 sg13g2_a221oi_1 _26827_ (.B2(net928),
    .C1(_11490_),
    .B1(_12156_),
    .A1(_09361_),
    .Y(_07627_),
    .A2(_09813_));
 sg13g2_or2_1 _26828_ (.X(_07628_),
    .B(_07627_),
    .A(_08343_));
 sg13g2_and2_1 _26829_ (.A(net803),
    .B(_07628_),
    .X(_07629_));
 sg13g2_inv_1 _26830_ (.Y(_07630_),
    .A(_07629_));
 sg13g2_a21oi_1 _26831_ (.A1(_09243_),
    .A2(_07626_),
    .Y(_01055_),
    .B1(_07630_));
 sg13g2_nor3_1 _26832_ (.A(_09213_),
    .B(_05012_),
    .C(_05034_),
    .Y(_07631_));
 sg13g2_nand2b_1 _26833_ (.Y(_07632_),
    .B(_07625_),
    .A_N(_07631_));
 sg13g2_a21oi_1 _26834_ (.A1(_09242_),
    .A2(_07632_),
    .Y(_01056_),
    .B1(_07630_));
 sg13g2_inv_1 _26835_ (.Y(_07633_),
    .A(\cpu.icache.r_valid[0] ));
 sg13g2_nand2b_1 _26836_ (.Y(_07634_),
    .B(net803),
    .A_N(\cpu.ex.i_flush_all ));
 sg13g2_buf_2 _26837_ (.A(_07634_),
    .X(_07635_));
 sg13g2_a21oi_1 _26838_ (.A1(_07633_),
    .A2(_06609_),
    .Y(_02411_),
    .B1(_07635_));
 sg13g2_nor2_1 _26839_ (.A(\cpu.icache.r_valid[1] ),
    .B(_06529_),
    .Y(_07636_));
 sg13g2_nor2_1 _26840_ (.A(_07635_),
    .B(_07636_),
    .Y(_02412_));
 sg13g2_nor2_1 _26841_ (.A(\cpu.icache.r_valid[2] ),
    .B(_06546_),
    .Y(_07637_));
 sg13g2_nor2_1 _26842_ (.A(_07635_),
    .B(_07637_),
    .Y(_02413_));
 sg13g2_inv_1 _26843_ (.Y(_07638_),
    .A(\cpu.icache.r_valid[3] ));
 sg13g2_a21oi_1 _26844_ (.A1(_07638_),
    .A2(net294),
    .Y(_02414_),
    .B1(_07635_));
 sg13g2_nor2_1 _26845_ (.A(\cpu.icache.r_valid[4] ),
    .B(_06571_),
    .Y(_07639_));
 sg13g2_nor2_1 _26846_ (.A(_07635_),
    .B(_07639_),
    .Y(_02415_));
 sg13g2_nor2_1 _26847_ (.A(\cpu.icache.r_valid[5] ),
    .B(_06586_),
    .Y(_07640_));
 sg13g2_nor2_1 _26848_ (.A(_07635_),
    .B(_07640_),
    .Y(_02416_));
 sg13g2_inv_1 _26849_ (.Y(_07641_),
    .A(\cpu.icache.r_valid[6] ));
 sg13g2_a21oi_1 _26850_ (.A1(_07641_),
    .A2(_06595_),
    .Y(_02417_),
    .B1(_07635_));
 sg13g2_nor2_1 _26851_ (.A(\cpu.icache.r_valid[7] ),
    .B(_06606_),
    .Y(_07642_));
 sg13g2_nor2_1 _26852_ (.A(_07635_),
    .B(_07642_),
    .Y(_02418_));
 sg13g2_nand3_1 _26853_ (.B(net103),
    .C(net445),
    .A(net1128),
    .Y(_07643_));
 sg13g2_and2_1 _26854_ (.A(net103),
    .B(net406),
    .X(_07644_));
 sg13g2_buf_1 _26855_ (.A(_07644_),
    .X(_07645_));
 sg13g2_a22oi_1 _26856_ (.Y(_07646_),
    .B1(_07645_),
    .B2(net954),
    .A2(_07643_),
    .A1(_09163_));
 sg13g2_nor2_1 _26857_ (.A(net705),
    .B(_07646_),
    .Y(_00305_));
 sg13g2_nor2_1 _26858_ (.A(_02934_),
    .B(_12029_),
    .Y(_07647_));
 sg13g2_nor2b_1 _26859_ (.A(_07647_),
    .B_N(_00303_),
    .Y(_00574_));
 sg13g2_a21oi_1 _26860_ (.A1(_12028_),
    .A2(_12087_),
    .Y(_00575_),
    .B1(_07647_));
 sg13g2_xnor2_1 _26861_ (.Y(_07648_),
    .A(_12031_),
    .B(_12046_));
 sg13g2_nor2_1 _26862_ (.A(_07647_),
    .B(_07648_),
    .Y(_00576_));
 sg13g2_nor2_1 _26863_ (.A(_09241_),
    .B(net522),
    .Y(_07649_));
 sg13g2_a21oi_1 _26864_ (.A1(net1083),
    .A2(net522),
    .Y(_07650_),
    .B1(_07649_));
 sg13g2_nor2_1 _26865_ (.A(_09323_),
    .B(_07650_),
    .Y(_00785_));
 sg13g2_nand2_1 _26866_ (.Y(_07651_),
    .A(_08454_),
    .B(net665));
 sg13g2_o21ai_1 _26867_ (.B1(_11466_),
    .Y(_07652_),
    .A1(_04100_),
    .A2(_07651_));
 sg13g2_buf_1 _26868_ (.A(_07652_),
    .X(_07653_));
 sg13g2_nand2_1 _26869_ (.Y(_07654_),
    .A(net994),
    .B(_07653_));
 sg13g2_nor2_1 _26870_ (.A(_10657_),
    .B(_09336_),
    .Y(_07655_));
 sg13g2_nand3_1 _26871_ (.B(_10932_),
    .C(_07655_),
    .A(_04096_),
    .Y(_07656_));
 sg13g2_a21oi_1 _26872_ (.A1(net994),
    .A2(_07656_),
    .Y(_07657_),
    .B1(_09316_));
 sg13g2_nor2_1 _26873_ (.A(_03820_),
    .B(_07657_),
    .Y(_07658_));
 sg13g2_nor2_1 _26874_ (.A(_10657_),
    .B(_07658_),
    .Y(_07659_));
 sg13g2_a21oi_1 _26875_ (.A1(_11056_),
    .A2(_07658_),
    .Y(_07660_),
    .B1(_07659_));
 sg13g2_nand2b_1 _26876_ (.Y(_07661_),
    .B(_07660_),
    .A_N(_07653_));
 sg13g2_nand3_1 _26877_ (.B(_07654_),
    .C(_07661_),
    .A(_09159_),
    .Y(_00786_));
 sg13g2_nand2_1 _26878_ (.Y(_07662_),
    .A(_10723_),
    .B(net522));
 sg13g2_o21ai_1 _26879_ (.B1(_07662_),
    .Y(_07663_),
    .A1(_02962_),
    .A2(net522));
 sg13g2_and2_1 _26880_ (.A(_11913_),
    .B(_07663_),
    .X(_00787_));
 sg13g2_nor3_1 _26881_ (.A(\cpu.ex.r_branch_stall ),
    .B(_11465_),
    .C(_03448_),
    .Y(_07664_));
 sg13g2_nand3_1 _26882_ (.B(net665),
    .C(_07664_),
    .A(_08343_),
    .Y(_07665_));
 sg13g2_nand3_1 _26883_ (.B(_07628_),
    .C(_07665_),
    .A(_11459_),
    .Y(_07666_));
 sg13g2_nand3_1 _26884_ (.B(_11470_),
    .C(_07666_),
    .A(net1143),
    .Y(_07667_));
 sg13g2_and3_1 _26885_ (.X(_07668_),
    .A(_06898_),
    .B(net36),
    .C(_07667_));
 sg13g2_nor2_1 _26886_ (.A(_06898_),
    .B(net166),
    .Y(_07669_));
 sg13g2_o21ai_1 _26887_ (.B1(_05863_),
    .Y(_00933_),
    .A1(_07668_),
    .A2(_07669_));
 sg13g2_nand2_1 _26888_ (.Y(_07670_),
    .A(_09361_),
    .B(_09336_));
 sg13g2_nand3_1 _26889_ (.B(\cpu.dec.do_flush_write ),
    .C(_11474_),
    .A(net994),
    .Y(_07671_));
 sg13g2_a21oi_1 _26890_ (.A1(_07670_),
    .A2(_07671_),
    .Y(_00934_),
    .B1(net656));
 sg13g2_nand2_1 _26891_ (.Y(_07672_),
    .A(\cpu.dec.io ),
    .B(_11474_));
 sg13g2_nand2_1 _26892_ (.Y(_07673_),
    .A(_04834_),
    .B(_09336_));
 sg13g2_a21oi_1 _26893_ (.A1(_07672_),
    .A2(_07673_),
    .Y(_00937_),
    .B1(net656));
 sg13g2_nor2b_1 _26894_ (.A(_09160_),
    .B_N(_07653_),
    .Y(_07674_));
 sg13g2_nand2_1 _26895_ (.Y(_07675_),
    .A(_10625_),
    .B(_07616_));
 sg13g2_o21ai_1 _26896_ (.B1(_07675_),
    .Y(_07676_),
    .A1(net622),
    .A2(net522));
 sg13g2_nor2_1 _26897_ (.A(_07653_),
    .B(_07676_),
    .Y(_07677_));
 sg13g2_nor3_1 _26898_ (.A(net800),
    .B(_07674_),
    .C(_07677_),
    .Y(_00984_));
 sg13g2_buf_1 _26899_ (.A(_09852_),
    .X(_07678_));
 sg13g2_a22oi_1 _26900_ (.Y(_07679_),
    .B1(_11492_),
    .B2(_09214_),
    .A2(_11474_),
    .A1(_11465_));
 sg13g2_nor2_1 _26901_ (.A(_07678_),
    .B(_07679_),
    .Y(_00985_));
 sg13g2_nor2_2 _26902_ (.A(net993),
    .B(_05829_),
    .Y(_07680_));
 sg13g2_mux2_1 _26903_ (.A0(_10604_),
    .A1(_09298_),
    .S(_07680_),
    .X(_07681_));
 sg13g2_nand2b_1 _26904_ (.Y(_07682_),
    .B(_07681_),
    .A_N(net270));
 sg13g2_a21oi_1 _26905_ (.A1(_11466_),
    .A2(_07682_),
    .Y(_01061_),
    .B1(net656));
 sg13g2_mux2_1 _26906_ (.A0(net965),
    .A1(_12475_),
    .S(_07680_),
    .X(_07683_));
 sg13g2_nand2_1 _26907_ (.Y(_07684_),
    .A(_09363_),
    .B(_04573_));
 sg13g2_o21ai_1 _26908_ (.B1(_07684_),
    .Y(_07685_),
    .A1(net270),
    .A2(_07683_));
 sg13g2_nor2_1 _26909_ (.A(_07678_),
    .B(_07685_),
    .Y(_01062_));
 sg13g2_mux2_1 _26910_ (.A0(\cpu.ex.mmu_read[1] ),
    .A1(_03507_),
    .S(_07680_),
    .X(_07686_));
 sg13g2_nand2_1 _26911_ (.Y(_07687_),
    .A(_08388_),
    .B(_07686_));
 sg13g2_a21oi_1 _26912_ (.A1(_04462_),
    .A2(_07687_),
    .Y(_01063_),
    .B1(net656));
 sg13g2_nor4_2 _26913_ (.A(_10558_),
    .B(_05865_),
    .C(_05831_),
    .Y(_07688_),
    .D(_05929_));
 sg13g2_nor2b_1 _26914_ (.A(_00241_),
    .B_N(_05828_),
    .Y(_07689_));
 sg13g2_o21ai_1 _26915_ (.B1(_07689_),
    .Y(_07690_),
    .A1(_11056_),
    .A2(_00239_));
 sg13g2_a21oi_1 _26916_ (.A1(net660),
    .A2(_07690_),
    .Y(_07691_),
    .B1(net371));
 sg13g2_nand2_1 _26917_ (.Y(_07692_),
    .A(net660),
    .B(_07691_));
 sg13g2_buf_1 _26918_ (.A(_07692_),
    .X(_07693_));
 sg13g2_buf_1 _26919_ (.A(_07693_),
    .X(_07694_));
 sg13g2_a21oi_1 _26920_ (.A1(_03328_),
    .A2(_10651_),
    .Y(_07695_),
    .B1(net660));
 sg13g2_nor2b_1 _26921_ (.A(_07695_),
    .B_N(_07691_),
    .Y(_07696_));
 sg13g2_buf_2 _26922_ (.A(_07696_),
    .X(_07697_));
 sg13g2_o21ai_1 _26923_ (.B1(_07697_),
    .Y(_07698_),
    .A1(_07688_),
    .A2(_07694_));
 sg13g2_nor2_1 _26924_ (.A(_10042_),
    .B(_07693_),
    .Y(_07699_));
 sg13g2_buf_2 _26925_ (.A(_07699_),
    .X(_07700_));
 sg13g2_buf_1 _26926_ (.A(_07700_),
    .X(_07701_));
 sg13g2_a22oi_1 _26927_ (.Y(_07702_),
    .B1(_07701_),
    .B2(_07688_),
    .A2(_07698_),
    .A1(\cpu.genblk1.mmu.r_valid_d[0] ));
 sg13g2_nor2_1 _26928_ (.A(net654),
    .B(_07702_),
    .Y(_01064_));
 sg13g2_o21ai_1 _26929_ (.B1(_07697_),
    .Y(_07703_),
    .A1(_05895_),
    .A2(_07694_));
 sg13g2_nor3_1 _26930_ (.A(net852),
    .B(net983),
    .C(net659),
    .Y(_07704_));
 sg13g2_buf_2 _26931_ (.A(_07704_),
    .X(_07705_));
 sg13g2_and2_1 _26932_ (.A(net660),
    .B(_07691_),
    .X(_07706_));
 sg13g2_buf_1 _26933_ (.A(_07706_),
    .X(_07707_));
 sg13g2_nor4_1 _26934_ (.A(net979),
    .B(_10474_),
    .C(net977),
    .D(_05831_),
    .Y(_07708_));
 sg13g2_nor2_1 _26935_ (.A(net979),
    .B(_10474_),
    .Y(_07709_));
 sg13g2_a21oi_1 _26936_ (.A1(_05830_),
    .A2(_07709_),
    .Y(_07710_),
    .B1(net1044));
 sg13g2_a21oi_1 _26937_ (.A1(net980),
    .A2(_07708_),
    .Y(_07711_),
    .B1(_07710_));
 sg13g2_nand2b_1 _26938_ (.Y(_07712_),
    .B(_07708_),
    .A_N(_05938_));
 sg13g2_o21ai_1 _26939_ (.B1(_07712_),
    .Y(_07713_),
    .A1(net965),
    .A2(_07711_));
 sg13g2_buf_1 _26940_ (.A(_07713_),
    .X(_07714_));
 sg13g2_and2_1 _26941_ (.A(_07707_),
    .B(_07714_),
    .X(_07715_));
 sg13g2_buf_1 _26942_ (.A(_07715_),
    .X(_07716_));
 sg13g2_a22oi_1 _26943_ (.Y(_07717_),
    .B1(_07705_),
    .B2(_07716_),
    .A2(_07703_),
    .A1(\cpu.genblk1.mmu.r_valid_d[10] ));
 sg13g2_nor2_1 _26944_ (.A(net654),
    .B(_07717_),
    .Y(_01065_));
 sg13g2_buf_1 _26945_ (.A(_07693_),
    .X(_07718_));
 sg13g2_buf_1 _26946_ (.A(_07697_),
    .X(_07719_));
 sg13g2_o21ai_1 _26947_ (.B1(_07719_),
    .Y(_07720_),
    .A1(_05900_),
    .A2(_07718_));
 sg13g2_a22oi_1 _26948_ (.Y(_07721_),
    .B1(_07720_),
    .B2(\cpu.genblk1.mmu.r_valid_d[11] ),
    .A2(_07700_),
    .A1(_05900_));
 sg13g2_nor2_1 _26949_ (.A(net654),
    .B(_07721_),
    .Y(_01066_));
 sg13g2_nand2_1 _26950_ (.Y(_07722_),
    .A(net978),
    .B(_05844_));
 sg13g2_nand3_1 _26951_ (.B(_05842_),
    .C(net976),
    .A(_05840_),
    .Y(_07723_));
 sg13g2_a21oi_2 _26952_ (.B1(_05831_),
    .Y(_07724_),
    .A2(_07723_),
    .A1(_07722_));
 sg13g2_nand2_1 _26953_ (.Y(_07725_),
    .A(_07714_),
    .B(_07724_));
 sg13g2_inv_1 _26954_ (.Y(_07726_),
    .A(_07725_));
 sg13g2_o21ai_1 _26955_ (.B1(_07697_),
    .Y(_07727_),
    .A1(net183),
    .A2(_07726_));
 sg13g2_nand2b_1 _26956_ (.Y(_07728_),
    .B(net852),
    .A_N(net983));
 sg13g2_nor3_1 _26957_ (.A(net980),
    .B(net979),
    .C(_07728_),
    .Y(_07729_));
 sg13g2_buf_2 _26958_ (.A(_07729_),
    .X(_07730_));
 sg13g2_a22oi_1 _26959_ (.Y(_07731_),
    .B1(_07730_),
    .B2(_07716_),
    .A2(_07727_),
    .A1(\cpu.genblk1.mmu.r_valid_d[12] ));
 sg13g2_nor2_1 _26960_ (.A(net654),
    .B(_07731_),
    .Y(_01067_));
 sg13g2_nor2_1 _26961_ (.A(_05852_),
    .B(_05909_),
    .Y(_07732_));
 sg13g2_and2_1 _26962_ (.A(_07714_),
    .B(_07732_),
    .X(_07733_));
 sg13g2_buf_1 _26963_ (.A(_07733_),
    .X(_07734_));
 sg13g2_o21ai_1 _26964_ (.B1(net181),
    .Y(_07735_),
    .A1(net182),
    .A2(_07734_));
 sg13g2_a22oi_1 _26965_ (.Y(_07736_),
    .B1(_07735_),
    .B2(\cpu.genblk1.mmu.r_valid_d[13] ),
    .A2(_07734_),
    .A1(net128));
 sg13g2_nor2_1 _26966_ (.A(net654),
    .B(_07736_),
    .Y(_01068_));
 sg13g2_and2_1 _26967_ (.A(_06028_),
    .B(_07714_),
    .X(_07737_));
 sg13g2_o21ai_1 _26968_ (.B1(_07697_),
    .Y(_07738_),
    .A1(net183),
    .A2(_07737_));
 sg13g2_nor2_1 _26969_ (.A(net659),
    .B(_07728_),
    .Y(_07739_));
 sg13g2_buf_2 _26970_ (.A(_07739_),
    .X(_07740_));
 sg13g2_a22oi_1 _26971_ (.Y(_07741_),
    .B1(_07740_),
    .B2(_07716_),
    .A2(_07738_),
    .A1(\cpu.genblk1.mmu.r_valid_d[14] ));
 sg13g2_nor2_1 _26972_ (.A(net654),
    .B(_07741_),
    .Y(_01069_));
 sg13g2_nor2_2 _26973_ (.A(_05868_),
    .B(_05894_),
    .Y(_07742_));
 sg13g2_o21ai_1 _26974_ (.B1(net181),
    .Y(_07743_),
    .A1(net182),
    .A2(_07742_));
 sg13g2_a22oi_1 _26975_ (.Y(_07744_),
    .B1(_07743_),
    .B2(\cpu.genblk1.mmu.r_valid_d[15] ),
    .A2(_07742_),
    .A1(_07701_));
 sg13g2_nor2_1 _26976_ (.A(net654),
    .B(_07744_),
    .Y(_01070_));
 sg13g2_nor4_1 _26977_ (.A(net979),
    .B(net852),
    .C(net977),
    .D(_05938_),
    .Y(_07745_));
 sg13g2_o21ai_1 _26978_ (.B1(_05830_),
    .Y(_07746_),
    .A1(_07742_),
    .A2(_07745_));
 sg13g2_inv_1 _26979_ (.Y(_07747_),
    .A(_07746_));
 sg13g2_a21oi_1 _26980_ (.A1(_03328_),
    .A2(_10583_),
    .Y(_07748_),
    .B1(_05827_));
 sg13g2_nor2b_1 _26981_ (.A(_07748_),
    .B_N(_07691_),
    .Y(_07749_));
 sg13g2_buf_2 _26982_ (.A(_07749_),
    .X(_07750_));
 sg13g2_o21ai_1 _26983_ (.B1(_07750_),
    .Y(_07751_),
    .A1(_07693_),
    .A2(_07747_));
 sg13g2_a21oi_1 _26984_ (.A1(_05830_),
    .A2(_05879_),
    .Y(_07752_),
    .B1(_04852_));
 sg13g2_and2_1 _26985_ (.A(_06128_),
    .B(_07752_),
    .X(_07753_));
 sg13g2_buf_2 _26986_ (.A(_07753_),
    .X(_07754_));
 sg13g2_a22oi_1 _26987_ (.Y(_07755_),
    .B1(_07754_),
    .B2(_07716_),
    .A2(_07751_),
    .A1(\cpu.genblk1.mmu.r_valid_d[16] ));
 sg13g2_nor2_1 _26988_ (.A(net654),
    .B(_07755_),
    .Y(_01071_));
 sg13g2_buf_1 _26989_ (.A(_09852_),
    .X(_07756_));
 sg13g2_nor2_1 _26990_ (.A(net852),
    .B(_05909_),
    .Y(_07757_));
 sg13g2_nand2_1 _26991_ (.Y(_07758_),
    .A(net980),
    .B(_05831_));
 sg13g2_a21oi_1 _26992_ (.A1(_07709_),
    .A2(_07758_),
    .Y(_07759_),
    .B1(net977));
 sg13g2_nor4_1 _26993_ (.A(_10558_),
    .B(net980),
    .C(net977),
    .D(_05830_),
    .Y(_07760_));
 sg13g2_a21oi_1 _26994_ (.A1(_05830_),
    .A2(_06232_),
    .Y(_07761_),
    .B1(_07760_));
 sg13g2_nor2b_1 _26995_ (.A(_07761_),
    .B_N(_07709_),
    .Y(_07762_));
 sg13g2_a21o_1 _26996_ (.A2(_07759_),
    .A1(net965),
    .B1(_07762_),
    .X(_07763_));
 sg13g2_buf_1 _26997_ (.A(_07763_),
    .X(_07764_));
 sg13g2_and2_1 _26998_ (.A(_07757_),
    .B(_07764_),
    .X(_07765_));
 sg13g2_buf_1 _26999_ (.A(_07765_),
    .X(_07766_));
 sg13g2_buf_1 _27000_ (.A(_07750_),
    .X(_07767_));
 sg13g2_o21ai_1 _27001_ (.B1(net180),
    .Y(_07768_),
    .A1(net182),
    .A2(_07766_));
 sg13g2_a22oi_1 _27002_ (.Y(_07769_),
    .B1(_07768_),
    .B2(\cpu.genblk1.mmu.r_valid_d[17] ),
    .A2(_07766_),
    .A1(net128));
 sg13g2_nor2_1 _27003_ (.A(net653),
    .B(_07769_),
    .Y(_01072_));
 sg13g2_o21ai_1 _27004_ (.B1(_07750_),
    .Y(_07770_),
    .A1(_05939_),
    .A2(net183));
 sg13g2_and2_1 _27005_ (.A(net202),
    .B(_07764_),
    .X(_07771_));
 sg13g2_buf_1 _27006_ (.A(_07771_),
    .X(_07772_));
 sg13g2_a22oi_1 _27007_ (.Y(_07773_),
    .B1(_07772_),
    .B2(_07705_),
    .A2(_07770_),
    .A1(\cpu.genblk1.mmu.r_valid_d[18] ));
 sg13g2_nor2_1 _27008_ (.A(net653),
    .B(_07773_),
    .Y(_01073_));
 sg13g2_o21ai_1 _27009_ (.B1(net180),
    .Y(_07774_),
    .A1(_05947_),
    .A2(net182));
 sg13g2_a22oi_1 _27010_ (.Y(_07775_),
    .B1(_07774_),
    .B2(\cpu.genblk1.mmu.r_valid_d[19] ),
    .A2(_07700_),
    .A1(_05947_));
 sg13g2_nor2_1 _27011_ (.A(net653),
    .B(_07775_),
    .Y(_01074_));
 sg13g2_nand2b_1 _27012_ (.Y(_07776_),
    .B(_07759_),
    .A_N(net965));
 sg13g2_nor2_1 _27013_ (.A(_05831_),
    .B(_05894_),
    .Y(_07777_));
 sg13g2_nor3_1 _27014_ (.A(net977),
    .B(_05830_),
    .C(_05938_),
    .Y(_07778_));
 sg13g2_o21ai_1 _27015_ (.B1(_07709_),
    .Y(_07779_),
    .A1(_07777_),
    .A2(_07778_));
 sg13g2_nand2_1 _27016_ (.Y(_07780_),
    .A(_07776_),
    .B(_07779_));
 sg13g2_buf_1 _27017_ (.A(_07780_),
    .X(_07781_));
 sg13g2_and2_1 _27018_ (.A(_07757_),
    .B(_07781_),
    .X(_07782_));
 sg13g2_buf_1 _27019_ (.A(_07782_),
    .X(_07783_));
 sg13g2_buf_1 _27020_ (.A(_07693_),
    .X(_07784_));
 sg13g2_o21ai_1 _27021_ (.B1(net181),
    .Y(_07785_),
    .A1(net179),
    .A2(_07783_));
 sg13g2_a22oi_1 _27022_ (.Y(_07786_),
    .B1(_07785_),
    .B2(\cpu.genblk1.mmu.r_valid_d[1] ),
    .A2(_07783_),
    .A1(net128));
 sg13g2_nor2_1 _27023_ (.A(_07756_),
    .B(_07786_),
    .Y(_01075_));
 sg13g2_and2_1 _27024_ (.A(_07724_),
    .B(_07764_),
    .X(_07787_));
 sg13g2_o21ai_1 _27025_ (.B1(net180),
    .Y(_07788_),
    .A1(net179),
    .A2(_07787_));
 sg13g2_a22oi_1 _27026_ (.Y(_07789_),
    .B1(_07788_),
    .B2(\cpu.genblk1.mmu.r_valid_d[20] ),
    .A2(_07772_),
    .A1(_07730_));
 sg13g2_nor2_1 _27027_ (.A(net653),
    .B(_07789_),
    .Y(_01076_));
 sg13g2_and2_1 _27028_ (.A(_07732_),
    .B(_07764_),
    .X(_07790_));
 sg13g2_buf_1 _27029_ (.A(_07790_),
    .X(_07791_));
 sg13g2_o21ai_1 _27030_ (.B1(net180),
    .Y(_07792_),
    .A1(net179),
    .A2(_07791_));
 sg13g2_a22oi_1 _27031_ (.Y(_07793_),
    .B1(_07792_),
    .B2(\cpu.genblk1.mmu.r_valid_d[21] ),
    .A2(_07791_),
    .A1(net128));
 sg13g2_nor2_1 _27032_ (.A(net653),
    .B(_07793_),
    .Y(_01077_));
 sg13g2_nand2_1 _27033_ (.Y(_07794_),
    .A(_06028_),
    .B(_07764_));
 sg13g2_inv_1 _27034_ (.Y(_07795_),
    .A(_07794_));
 sg13g2_o21ai_1 _27035_ (.B1(net180),
    .Y(_07796_),
    .A1(net179),
    .A2(_07795_));
 sg13g2_a22oi_1 _27036_ (.Y(_07797_),
    .B1(_07796_),
    .B2(\cpu.genblk1.mmu.r_valid_d[22] ),
    .A2(_07772_),
    .A1(_07740_));
 sg13g2_nor2_1 _27037_ (.A(net653),
    .B(_07797_),
    .Y(_01078_));
 sg13g2_nor2_2 _27038_ (.A(_05868_),
    .B(_05928_),
    .Y(_07798_));
 sg13g2_o21ai_1 _27039_ (.B1(net180),
    .Y(_07799_),
    .A1(net179),
    .A2(_07798_));
 sg13g2_a22oi_1 _27040_ (.Y(_07800_),
    .B1(_07799_),
    .B2(\cpu.genblk1.mmu.r_valid_d[23] ),
    .A2(_07798_),
    .A1(net128));
 sg13g2_nor2_1 _27041_ (.A(net653),
    .B(_07800_),
    .Y(_01079_));
 sg13g2_a21oi_1 _27042_ (.A1(net977),
    .A2(_06128_),
    .Y(_07801_),
    .B1(_05869_));
 sg13g2_nand3b_1 _27043_ (.B(_05830_),
    .C(net965),
    .Y(_07802_),
    .A_N(_07801_));
 sg13g2_inv_1 _27044_ (.Y(_07803_),
    .A(_07802_));
 sg13g2_o21ai_1 _27045_ (.B1(net180),
    .Y(_07804_),
    .A1(net179),
    .A2(_07803_));
 sg13g2_a22oi_1 _27046_ (.Y(_07805_),
    .B1(_07804_),
    .B2(\cpu.genblk1.mmu.r_valid_d[24] ),
    .A2(_07772_),
    .A1(_07754_));
 sg13g2_nor2_1 _27047_ (.A(net653),
    .B(_07805_),
    .Y(_01080_));
 sg13g2_nand2b_1 _27048_ (.Y(_07806_),
    .B(_06127_),
    .A_N(_07711_));
 sg13g2_nand2b_1 _27049_ (.Y(_07807_),
    .B(_07806_),
    .A_N(_07688_));
 sg13g2_buf_1 _27050_ (.A(_07807_),
    .X(_07808_));
 sg13g2_and2_1 _27051_ (.A(_07757_),
    .B(net466),
    .X(_07809_));
 sg13g2_buf_1 _27052_ (.A(_07809_),
    .X(_07810_));
 sg13g2_o21ai_1 _27053_ (.B1(_07767_),
    .Y(_07811_),
    .A1(net179),
    .A2(_07810_));
 sg13g2_a22oi_1 _27054_ (.Y(_07812_),
    .B1(_07811_),
    .B2(\cpu.genblk1.mmu.r_valid_d[25] ),
    .A2(_07810_),
    .A1(net128));
 sg13g2_nor2_1 _27055_ (.A(_07756_),
    .B(_07812_),
    .Y(_01081_));
 sg13g2_o21ai_1 _27056_ (.B1(_07750_),
    .Y(_07813_),
    .A1(_05985_),
    .A2(net182));
 sg13g2_nand2_1 _27057_ (.Y(_07814_),
    .A(\cpu.genblk1.mmu.r_valid_d[26] ),
    .B(_07813_));
 sg13g2_nand3_1 _27058_ (.B(_07705_),
    .C(net466),
    .A(net202),
    .Y(_07815_));
 sg13g2_a21oi_1 _27059_ (.A1(_07814_),
    .A2(_07815_),
    .Y(_01082_),
    .B1(net656));
 sg13g2_buf_1 _27060_ (.A(_09852_),
    .X(_07816_));
 sg13g2_o21ai_1 _27061_ (.B1(net180),
    .Y(_07817_),
    .A1(_05990_),
    .A2(net182));
 sg13g2_a22oi_1 _27062_ (.Y(_07818_),
    .B1(_07817_),
    .B2(\cpu.genblk1.mmu.r_valid_d[27] ),
    .A2(_07700_),
    .A1(_05990_));
 sg13g2_nor2_1 _27063_ (.A(net652),
    .B(_07818_),
    .Y(_01083_));
 sg13g2_and2_1 _27064_ (.A(_07724_),
    .B(net466),
    .X(_07819_));
 sg13g2_o21ai_1 _27065_ (.B1(_07750_),
    .Y(_07820_),
    .A1(net183),
    .A2(_07819_));
 sg13g2_nand2_1 _27066_ (.Y(_07821_),
    .A(\cpu.genblk1.mmu.r_valid_d[28] ),
    .B(_07820_));
 sg13g2_nand3_1 _27067_ (.B(_07730_),
    .C(net466),
    .A(net202),
    .Y(_07822_));
 sg13g2_a21oi_1 _27068_ (.A1(_07821_),
    .A2(_07822_),
    .Y(_01084_),
    .B1(net656));
 sg13g2_and2_1 _27069_ (.A(_07732_),
    .B(net466),
    .X(_07823_));
 sg13g2_buf_1 _27070_ (.A(_07823_),
    .X(_07824_));
 sg13g2_o21ai_1 _27071_ (.B1(_07767_),
    .Y(_07825_),
    .A1(net179),
    .A2(_07824_));
 sg13g2_a22oi_1 _27072_ (.Y(_07826_),
    .B1(_07825_),
    .B2(\cpu.genblk1.mmu.r_valid_d[29] ),
    .A2(_07824_),
    .A1(net128));
 sg13g2_nor2_1 _27073_ (.A(net652),
    .B(_07826_),
    .Y(_01085_));
 sg13g2_inv_1 _27074_ (.Y(_07827_),
    .A(_07781_));
 sg13g2_nor3_1 _27075_ (.A(net852),
    .B(net659),
    .C(_07827_),
    .Y(_07828_));
 sg13g2_o21ai_1 _27076_ (.B1(_07697_),
    .Y(_07829_),
    .A1(_07693_),
    .A2(_07828_));
 sg13g2_nor2b_1 _27077_ (.A(_04852_),
    .B_N(_07828_),
    .Y(_07830_));
 sg13g2_a22oi_1 _27078_ (.Y(_07831_),
    .B1(_07830_),
    .B2(net202),
    .A2(_07829_),
    .A1(\cpu.genblk1.mmu.r_valid_d[2] ));
 sg13g2_nor2_1 _27079_ (.A(_07816_),
    .B(_07831_),
    .Y(_01086_));
 sg13g2_and2_1 _27080_ (.A(_06028_),
    .B(net466),
    .X(_07832_));
 sg13g2_o21ai_1 _27081_ (.B1(_07750_),
    .Y(_07833_),
    .A1(net183),
    .A2(_07832_));
 sg13g2_nand2_1 _27082_ (.Y(_07834_),
    .A(\cpu.genblk1.mmu.r_valid_d[30] ),
    .B(_07833_));
 sg13g2_nand3_1 _27083_ (.B(_07740_),
    .C(_07808_),
    .A(net202),
    .Y(_07835_));
 sg13g2_a21oi_1 _27084_ (.A1(_07834_),
    .A2(_07835_),
    .Y(_01087_),
    .B1(_06885_));
 sg13g2_nor2b_2 _27085_ (.A(_05868_),
    .B_N(net466),
    .Y(_07836_));
 sg13g2_o21ai_1 _27086_ (.B1(_07750_),
    .Y(_07837_),
    .A1(_07784_),
    .A2(_07836_));
 sg13g2_a22oi_1 _27087_ (.Y(_07838_),
    .B1(_07837_),
    .B2(\cpu.genblk1.mmu.r_valid_d[31] ),
    .A2(_07836_),
    .A1(net128));
 sg13g2_nor2_1 _27088_ (.A(net652),
    .B(_07838_),
    .Y(_01088_));
 sg13g2_nor2_2 _27089_ (.A(_07722_),
    .B(_07827_),
    .Y(_07839_));
 sg13g2_o21ai_1 _27090_ (.B1(net181),
    .Y(_07840_),
    .A1(_07784_),
    .A2(_07839_));
 sg13g2_a22oi_1 _27091_ (.Y(_07841_),
    .B1(_07840_),
    .B2(\cpu.genblk1.mmu.r_valid_d[3] ),
    .A2(_07839_),
    .A1(_07700_));
 sg13g2_nor2_1 _27092_ (.A(net652),
    .B(_07841_),
    .Y(_01089_));
 sg13g2_nand3_1 _27093_ (.B(_07730_),
    .C(_07781_),
    .A(net202),
    .Y(_07842_));
 sg13g2_and2_1 _27094_ (.A(_07724_),
    .B(_07781_),
    .X(_07843_));
 sg13g2_o21ai_1 _27095_ (.B1(_07697_),
    .Y(_07844_),
    .A1(net183),
    .A2(_07843_));
 sg13g2_nand2_1 _27096_ (.Y(_07845_),
    .A(\cpu.genblk1.mmu.r_valid_d[4] ),
    .B(_07844_));
 sg13g2_a21oi_1 _27097_ (.A1(_07842_),
    .A2(_07845_),
    .Y(_01090_),
    .B1(_06885_));
 sg13g2_o21ai_1 _27098_ (.B1(net181),
    .Y(_07846_),
    .A1(_06024_),
    .A2(net182));
 sg13g2_a22oi_1 _27099_ (.Y(_07847_),
    .B1(_07846_),
    .B2(\cpu.genblk1.mmu.r_valid_d[5] ),
    .A2(_07700_),
    .A1(_06024_));
 sg13g2_nor2_1 _27100_ (.A(net652),
    .B(_07847_),
    .Y(_01091_));
 sg13g2_o21ai_1 _27101_ (.B1(net181),
    .Y(_07848_),
    .A1(_06030_),
    .A2(net182));
 sg13g2_nand2_1 _27102_ (.Y(_07849_),
    .A(\cpu.genblk1.mmu.r_valid_d[6] ),
    .B(_07848_));
 sg13g2_nand3_1 _27103_ (.B(_07740_),
    .C(_07781_),
    .A(net202),
    .Y(_07850_));
 sg13g2_buf_1 _27104_ (.A(_09330_),
    .X(_07851_));
 sg13g2_a21oi_1 _27105_ (.A1(_07849_),
    .A2(_07850_),
    .Y(_01092_),
    .B1(_07851_));
 sg13g2_o21ai_1 _27106_ (.B1(_07719_),
    .Y(_07852_),
    .A1(_06035_),
    .A2(_07718_));
 sg13g2_a22oi_1 _27107_ (.Y(_07853_),
    .B1(_07852_),
    .B2(\cpu.genblk1.mmu.r_valid_d[7] ),
    .A2(_07700_),
    .A1(_06035_));
 sg13g2_nor2_1 _27108_ (.A(net652),
    .B(_07853_),
    .Y(_01093_));
 sg13g2_nor3_1 _27109_ (.A(_06127_),
    .B(_05831_),
    .C(_07801_),
    .Y(_07854_));
 sg13g2_o21ai_1 _27110_ (.B1(net181),
    .Y(_07855_),
    .A1(net183),
    .A2(_07854_));
 sg13g2_nand2_1 _27111_ (.Y(_07856_),
    .A(\cpu.genblk1.mmu.r_valid_d[8] ),
    .B(_07855_));
 sg13g2_nand3_1 _27112_ (.B(_07754_),
    .C(_07781_),
    .A(net202),
    .Y(_07857_));
 sg13g2_a21oi_1 _27113_ (.A1(_07856_),
    .A2(_07857_),
    .Y(_01094_),
    .B1(_07851_));
 sg13g2_and2_1 _27114_ (.A(_07714_),
    .B(_07757_),
    .X(_07858_));
 sg13g2_buf_1 _27115_ (.A(_07858_),
    .X(_07859_));
 sg13g2_o21ai_1 _27116_ (.B1(net181),
    .Y(_07860_),
    .A1(net183),
    .A2(_07859_));
 sg13g2_a22oi_1 _27117_ (.Y(_07861_),
    .B1(_07860_),
    .B2(\cpu.genblk1.mmu.r_valid_d[9] ),
    .A2(_07859_),
    .A1(_07700_));
 sg13g2_nor2_1 _27118_ (.A(net652),
    .B(_07861_),
    .Y(_01095_));
 sg13g2_inv_1 _27119_ (.Y(_07862_),
    .A(_00239_));
 sg13g2_o21ai_1 _27120_ (.B1(_07689_),
    .Y(_07863_),
    .A1(_11056_),
    .A2(_07862_));
 sg13g2_a21oi_1 _27121_ (.A1(_05826_),
    .A2(_07863_),
    .Y(_07864_),
    .B1(net371));
 sg13g2_nand2_1 _27122_ (.Y(_07865_),
    .A(net660),
    .B(_07864_));
 sg13g2_buf_1 _27123_ (.A(_07865_),
    .X(_07866_));
 sg13g2_nand3b_1 _27124_ (.B(_05824_),
    .C(_03328_),
    .Y(_07867_),
    .A_N(_10645_));
 sg13g2_and2_1 _27125_ (.A(_07864_),
    .B(_07867_),
    .X(_07868_));
 sg13g2_buf_2 _27126_ (.A(_07868_),
    .X(_07869_));
 sg13g2_o21ai_1 _27127_ (.B1(_07869_),
    .Y(_07870_),
    .A1(_07688_),
    .A2(_07866_));
 sg13g2_nor2_1 _27128_ (.A(_10042_),
    .B(_07866_),
    .Y(_07871_));
 sg13g2_buf_2 _27129_ (.A(_07871_),
    .X(_07872_));
 sg13g2_buf_1 _27130_ (.A(_07872_),
    .X(_07873_));
 sg13g2_a22oi_1 _27131_ (.Y(_07874_),
    .B1(net127),
    .B2(_07688_),
    .A2(_07870_),
    .A1(\cpu.genblk1.mmu.r_valid_i[0] ));
 sg13g2_nor2_1 _27132_ (.A(net652),
    .B(_07874_),
    .Y(_01096_));
 sg13g2_and2_1 _27133_ (.A(net660),
    .B(_07864_),
    .X(_07875_));
 sg13g2_buf_1 _27134_ (.A(_07875_),
    .X(_07876_));
 sg13g2_and2_1 _27135_ (.A(_07714_),
    .B(_07876_),
    .X(_07877_));
 sg13g2_buf_1 _27136_ (.A(_07877_),
    .X(_07878_));
 sg13g2_buf_1 _27137_ (.A(_07866_),
    .X(_07879_));
 sg13g2_buf_1 _27138_ (.A(_07869_),
    .X(_07880_));
 sg13g2_o21ai_1 _27139_ (.B1(net177),
    .Y(_07881_),
    .A1(_05895_),
    .A2(net178));
 sg13g2_a22oi_1 _27140_ (.Y(_07882_),
    .B1(_07881_),
    .B2(\cpu.genblk1.mmu.r_valid_i[10] ),
    .A2(_07878_),
    .A1(_07705_));
 sg13g2_nor2_1 _27141_ (.A(_07816_),
    .B(_07882_),
    .Y(_01097_));
 sg13g2_buf_1 _27142_ (.A(_09852_),
    .X(_07883_));
 sg13g2_o21ai_1 _27143_ (.B1(net177),
    .Y(_07884_),
    .A1(_05900_),
    .A2(_07879_));
 sg13g2_a22oi_1 _27144_ (.Y(_07885_),
    .B1(_07884_),
    .B2(\cpu.genblk1.mmu.r_valid_i[11] ),
    .A2(_07873_),
    .A1(_05900_));
 sg13g2_nor2_1 _27145_ (.A(net650),
    .B(_07885_),
    .Y(_01098_));
 sg13g2_o21ai_1 _27146_ (.B1(net177),
    .Y(_07886_),
    .A1(_07726_),
    .A2(net178));
 sg13g2_a22oi_1 _27147_ (.Y(_07887_),
    .B1(_07886_),
    .B2(\cpu.genblk1.mmu.r_valid_i[12] ),
    .A2(_07878_),
    .A1(_07730_));
 sg13g2_nor2_1 _27148_ (.A(net650),
    .B(_07887_),
    .Y(_01099_));
 sg13g2_o21ai_1 _27149_ (.B1(net177),
    .Y(_07888_),
    .A1(_07734_),
    .A2(_07879_));
 sg13g2_a22oi_1 _27150_ (.Y(_07889_),
    .B1(_07888_),
    .B2(\cpu.genblk1.mmu.r_valid_i[13] ),
    .A2(net127),
    .A1(_07734_));
 sg13g2_nor2_1 _27151_ (.A(_07883_),
    .B(_07889_),
    .Y(_01100_));
 sg13g2_o21ai_1 _27152_ (.B1(net177),
    .Y(_07890_),
    .A1(_07737_),
    .A2(net178));
 sg13g2_a22oi_1 _27153_ (.Y(_07891_),
    .B1(_07890_),
    .B2(\cpu.genblk1.mmu.r_valid_i[14] ),
    .A2(_07878_),
    .A1(_07740_));
 sg13g2_nor2_1 _27154_ (.A(net650),
    .B(_07891_),
    .Y(_01101_));
 sg13g2_o21ai_1 _27155_ (.B1(net177),
    .Y(_07892_),
    .A1(_07742_),
    .A2(net178));
 sg13g2_a22oi_1 _27156_ (.Y(_07893_),
    .B1(_07892_),
    .B2(\cpu.genblk1.mmu.r_valid_i[15] ),
    .A2(_07873_),
    .A1(_07742_));
 sg13g2_nor2_1 _27157_ (.A(_07883_),
    .B(_07893_),
    .Y(_01102_));
 sg13g2_a21oi_1 _27158_ (.A1(_03328_),
    .A2(_10613_),
    .Y(_07894_),
    .B1(_05827_));
 sg13g2_nor2b_1 _27159_ (.A(_07894_),
    .B_N(_07864_),
    .Y(_07895_));
 sg13g2_buf_2 _27160_ (.A(_07895_),
    .X(_07896_));
 sg13g2_buf_1 _27161_ (.A(_07896_),
    .X(_07897_));
 sg13g2_o21ai_1 _27162_ (.B1(_07897_),
    .Y(_07898_),
    .A1(_07747_),
    .A2(net178));
 sg13g2_a22oi_1 _27163_ (.Y(_07899_),
    .B1(_07898_),
    .B2(\cpu.genblk1.mmu.r_valid_i[16] ),
    .A2(_07878_),
    .A1(_07754_));
 sg13g2_nor2_1 _27164_ (.A(net650),
    .B(_07899_),
    .Y(_01103_));
 sg13g2_o21ai_1 _27165_ (.B1(net176),
    .Y(_07900_),
    .A1(_07766_),
    .A2(net178));
 sg13g2_a22oi_1 _27166_ (.Y(_07901_),
    .B1(_07900_),
    .B2(\cpu.genblk1.mmu.r_valid_i[17] ),
    .A2(net127),
    .A1(_07766_));
 sg13g2_nor2_1 _27167_ (.A(net650),
    .B(_07901_),
    .Y(_01104_));
 sg13g2_and2_1 _27168_ (.A(_07764_),
    .B(_07876_),
    .X(_07902_));
 sg13g2_buf_1 _27169_ (.A(_07902_),
    .X(_07903_));
 sg13g2_o21ai_1 _27170_ (.B1(net176),
    .Y(_07904_),
    .A1(_05939_),
    .A2(net178));
 sg13g2_a22oi_1 _27171_ (.Y(_07905_),
    .B1(_07904_),
    .B2(\cpu.genblk1.mmu.r_valid_i[18] ),
    .A2(_07903_),
    .A1(_07705_));
 sg13g2_nor2_1 _27172_ (.A(net650),
    .B(_07905_),
    .Y(_01105_));
 sg13g2_o21ai_1 _27173_ (.B1(net176),
    .Y(_07906_),
    .A1(_05947_),
    .A2(net178));
 sg13g2_a22oi_1 _27174_ (.Y(_07907_),
    .B1(_07906_),
    .B2(\cpu.genblk1.mmu.r_valid_i[19] ),
    .A2(net127),
    .A1(_05947_));
 sg13g2_nor2_1 _27175_ (.A(net650),
    .B(_07907_),
    .Y(_01106_));
 sg13g2_buf_1 _27176_ (.A(_07866_),
    .X(_07908_));
 sg13g2_o21ai_1 _27177_ (.B1(net177),
    .Y(_07909_),
    .A1(_07783_),
    .A2(_07908_));
 sg13g2_a22oi_1 _27178_ (.Y(_07910_),
    .B1(_07909_),
    .B2(\cpu.genblk1.mmu.r_valid_i[1] ),
    .A2(net127),
    .A1(_07783_));
 sg13g2_nor2_1 _27179_ (.A(net650),
    .B(_07910_),
    .Y(_01107_));
 sg13g2_buf_1 _27180_ (.A(_09852_),
    .X(_07911_));
 sg13g2_o21ai_1 _27181_ (.B1(net176),
    .Y(_07912_),
    .A1(_07787_),
    .A2(net175));
 sg13g2_a22oi_1 _27182_ (.Y(_07913_),
    .B1(_07912_),
    .B2(\cpu.genblk1.mmu.r_valid_i[20] ),
    .A2(_07903_),
    .A1(_07730_));
 sg13g2_nor2_1 _27183_ (.A(net649),
    .B(_07913_),
    .Y(_01108_));
 sg13g2_o21ai_1 _27184_ (.B1(net176),
    .Y(_07914_),
    .A1(_07791_),
    .A2(net175));
 sg13g2_a22oi_1 _27185_ (.Y(_07915_),
    .B1(_07914_),
    .B2(\cpu.genblk1.mmu.r_valid_i[21] ),
    .A2(net127),
    .A1(_07791_));
 sg13g2_nor2_1 _27186_ (.A(net649),
    .B(_07915_),
    .Y(_01109_));
 sg13g2_o21ai_1 _27187_ (.B1(net176),
    .Y(_07916_),
    .A1(_07795_),
    .A2(net175));
 sg13g2_a22oi_1 _27188_ (.Y(_07917_),
    .B1(_07916_),
    .B2(\cpu.genblk1.mmu.r_valid_i[22] ),
    .A2(_07903_),
    .A1(_07740_));
 sg13g2_nor2_1 _27189_ (.A(net649),
    .B(_07917_),
    .Y(_01110_));
 sg13g2_o21ai_1 _27190_ (.B1(net176),
    .Y(_07918_),
    .A1(_07798_),
    .A2(net175));
 sg13g2_a22oi_1 _27191_ (.Y(_07919_),
    .B1(_07918_),
    .B2(\cpu.genblk1.mmu.r_valid_i[23] ),
    .A2(net127),
    .A1(_07798_));
 sg13g2_nor2_1 _27192_ (.A(net649),
    .B(_07919_),
    .Y(_01111_));
 sg13g2_o21ai_1 _27193_ (.B1(net176),
    .Y(_07920_),
    .A1(_07803_),
    .A2(net175));
 sg13g2_a22oi_1 _27194_ (.Y(_07921_),
    .B1(_07920_),
    .B2(\cpu.genblk1.mmu.r_valid_i[24] ),
    .A2(_07903_),
    .A1(_07754_));
 sg13g2_nor2_1 _27195_ (.A(_07911_),
    .B(_07921_),
    .Y(_01112_));
 sg13g2_o21ai_1 _27196_ (.B1(_07897_),
    .Y(_07922_),
    .A1(_07810_),
    .A2(net175));
 sg13g2_a22oi_1 _27197_ (.Y(_07923_),
    .B1(_07922_),
    .B2(\cpu.genblk1.mmu.r_valid_i[25] ),
    .A2(net127),
    .A1(_07810_));
 sg13g2_nor2_1 _27198_ (.A(net649),
    .B(_07923_),
    .Y(_01113_));
 sg13g2_and2_1 _27199_ (.A(net466),
    .B(_07876_),
    .X(_07924_));
 sg13g2_buf_1 _27200_ (.A(_07924_),
    .X(_07925_));
 sg13g2_o21ai_1 _27201_ (.B1(_07896_),
    .Y(_07926_),
    .A1(_05985_),
    .A2(net175));
 sg13g2_a22oi_1 _27202_ (.Y(_07927_),
    .B1(_07926_),
    .B2(\cpu.genblk1.mmu.r_valid_i[26] ),
    .A2(_07925_),
    .A1(_07705_));
 sg13g2_nor2_1 _27203_ (.A(_07911_),
    .B(_07927_),
    .Y(_01114_));
 sg13g2_o21ai_1 _27204_ (.B1(_07896_),
    .Y(_07928_),
    .A1(_05990_),
    .A2(net175));
 sg13g2_a22oi_1 _27205_ (.Y(_07929_),
    .B1(_07928_),
    .B2(\cpu.genblk1.mmu.r_valid_i[27] ),
    .A2(_07872_),
    .A1(_05990_));
 sg13g2_nor2_1 _27206_ (.A(net649),
    .B(_07929_),
    .Y(_01115_));
 sg13g2_o21ai_1 _27207_ (.B1(_07896_),
    .Y(_07930_),
    .A1(_07819_),
    .A2(_07908_));
 sg13g2_a22oi_1 _27208_ (.Y(_07931_),
    .B1(_07930_),
    .B2(\cpu.genblk1.mmu.r_valid_i[28] ),
    .A2(_07925_),
    .A1(_07730_));
 sg13g2_nor2_1 _27209_ (.A(net649),
    .B(_07931_),
    .Y(_01116_));
 sg13g2_buf_1 _27210_ (.A(_07866_),
    .X(_07932_));
 sg13g2_o21ai_1 _27211_ (.B1(_07896_),
    .Y(_07933_),
    .A1(_07824_),
    .A2(net174));
 sg13g2_a22oi_1 _27212_ (.Y(_07934_),
    .B1(_07933_),
    .B2(\cpu.genblk1.mmu.r_valid_i[29] ),
    .A2(_07872_),
    .A1(_07824_));
 sg13g2_nor2_1 _27213_ (.A(net649),
    .B(_07934_),
    .Y(_01117_));
 sg13g2_buf_1 _27214_ (.A(_09852_),
    .X(_07935_));
 sg13g2_o21ai_1 _27215_ (.B1(_07880_),
    .Y(_07936_),
    .A1(_07828_),
    .A2(_07932_));
 sg13g2_a22oi_1 _27216_ (.Y(_07937_),
    .B1(_07936_),
    .B2(\cpu.genblk1.mmu.r_valid_i[2] ),
    .A2(_07876_),
    .A1(_07830_));
 sg13g2_nor2_1 _27217_ (.A(net648),
    .B(_07937_),
    .Y(_01118_));
 sg13g2_o21ai_1 _27218_ (.B1(_07896_),
    .Y(_07938_),
    .A1(_07832_),
    .A2(net174));
 sg13g2_a22oi_1 _27219_ (.Y(_07939_),
    .B1(_07938_),
    .B2(\cpu.genblk1.mmu.r_valid_i[30] ),
    .A2(_07925_),
    .A1(_07740_));
 sg13g2_nor2_1 _27220_ (.A(net648),
    .B(_07939_),
    .Y(_01119_));
 sg13g2_o21ai_1 _27221_ (.B1(_07896_),
    .Y(_07940_),
    .A1(_07836_),
    .A2(net174));
 sg13g2_a22oi_1 _27222_ (.Y(_07941_),
    .B1(_07940_),
    .B2(\cpu.genblk1.mmu.r_valid_i[31] ),
    .A2(_07872_),
    .A1(_07836_));
 sg13g2_nor2_1 _27223_ (.A(net648),
    .B(_07941_),
    .Y(_01120_));
 sg13g2_o21ai_1 _27224_ (.B1(net177),
    .Y(_07942_),
    .A1(_07839_),
    .A2(net174));
 sg13g2_a22oi_1 _27225_ (.Y(_07943_),
    .B1(_07942_),
    .B2(\cpu.genblk1.mmu.r_valid_i[3] ),
    .A2(_07872_),
    .A1(_07839_));
 sg13g2_nor2_1 _27226_ (.A(_07935_),
    .B(_07943_),
    .Y(_01121_));
 sg13g2_nor2_1 _27227_ (.A(_07827_),
    .B(_07866_),
    .Y(_07944_));
 sg13g2_o21ai_1 _27228_ (.B1(_07880_),
    .Y(_07945_),
    .A1(_07843_),
    .A2(net174));
 sg13g2_a22oi_1 _27229_ (.Y(_07946_),
    .B1(_07945_),
    .B2(\cpu.genblk1.mmu.r_valid_i[4] ),
    .A2(_07944_),
    .A1(_07730_));
 sg13g2_nor2_1 _27230_ (.A(_07935_),
    .B(_07946_),
    .Y(_01122_));
 sg13g2_o21ai_1 _27231_ (.B1(_07869_),
    .Y(_07947_),
    .A1(_06024_),
    .A2(net174));
 sg13g2_a22oi_1 _27232_ (.Y(_07948_),
    .B1(_07947_),
    .B2(\cpu.genblk1.mmu.r_valid_i[5] ),
    .A2(_07872_),
    .A1(_06024_));
 sg13g2_nor2_1 _27233_ (.A(net648),
    .B(_07948_),
    .Y(_01123_));
 sg13g2_o21ai_1 _27234_ (.B1(_07869_),
    .Y(_07949_),
    .A1(_06030_),
    .A2(_07932_));
 sg13g2_a22oi_1 _27235_ (.Y(_07950_),
    .B1(_07949_),
    .B2(\cpu.genblk1.mmu.r_valid_i[6] ),
    .A2(_07944_),
    .A1(_07740_));
 sg13g2_nor2_1 _27236_ (.A(net648),
    .B(_07950_),
    .Y(_01124_));
 sg13g2_o21ai_1 _27237_ (.B1(_07869_),
    .Y(_07951_),
    .A1(_06035_),
    .A2(net174));
 sg13g2_a22oi_1 _27238_ (.Y(_07952_),
    .B1(_07951_),
    .B2(\cpu.genblk1.mmu.r_valid_i[7] ),
    .A2(_07872_),
    .A1(_06035_));
 sg13g2_nor2_1 _27239_ (.A(net648),
    .B(_07952_),
    .Y(_01125_));
 sg13g2_o21ai_1 _27240_ (.B1(_07869_),
    .Y(_07953_),
    .A1(_07854_),
    .A2(net174));
 sg13g2_a22oi_1 _27241_ (.Y(_07954_),
    .B1(_07953_),
    .B2(\cpu.genblk1.mmu.r_valid_i[8] ),
    .A2(_07944_),
    .A1(_07754_));
 sg13g2_nor2_1 _27242_ (.A(net648),
    .B(_07954_),
    .Y(_01126_));
 sg13g2_o21ai_1 _27243_ (.B1(_07869_),
    .Y(_07955_),
    .A1(_07859_),
    .A2(_07866_));
 sg13g2_a22oi_1 _27244_ (.Y(_07956_),
    .B1(_07955_),
    .B2(\cpu.genblk1.mmu.r_valid_i[9] ),
    .A2(_07872_),
    .A1(_07859_));
 sg13g2_nor2_1 _27245_ (.A(net648),
    .B(_07956_),
    .Y(_01127_));
 sg13g2_and2_1 _27246_ (.A(net348),
    .B(net112),
    .X(_07957_));
 sg13g2_buf_2 _27247_ (.A(_07957_),
    .X(_07958_));
 sg13g2_nand2_1 _27248_ (.Y(_07959_),
    .A(_02704_),
    .B(_07958_));
 sg13g2_nand2_1 _27249_ (.Y(_07960_),
    .A(_04921_),
    .B(net112));
 sg13g2_buf_2 _27250_ (.A(_07960_),
    .X(_07961_));
 sg13g2_nand2_1 _27251_ (.Y(_07962_),
    .A(_09179_),
    .B(_07961_));
 sg13g2_a21oi_1 _27252_ (.A1(_07959_),
    .A2(_07962_),
    .Y(_01928_),
    .B1(net651));
 sg13g2_nand2_1 _27253_ (.Y(_07963_),
    .A(_10101_),
    .B(_07958_));
 sg13g2_nand2_1 _27254_ (.Y(_07964_),
    .A(_09181_),
    .B(_07961_));
 sg13g2_a21oi_1 _27255_ (.A1(_07963_),
    .A2(_07964_),
    .Y(_01929_),
    .B1(net651));
 sg13g2_nand2_1 _27256_ (.Y(_07965_),
    .A(net910),
    .B(_07958_));
 sg13g2_nand2_1 _27257_ (.Y(_07966_),
    .A(\cpu.gpio.r_enable_in[2] ),
    .B(_07961_));
 sg13g2_a21oi_1 _27258_ (.A1(_07965_),
    .A2(_07966_),
    .Y(_01930_),
    .B1(net651));
 sg13g2_nand2_1 _27259_ (.Y(_07967_),
    .A(_06861_),
    .B(_07958_));
 sg13g2_nand2_1 _27260_ (.Y(_07968_),
    .A(_09197_),
    .B(_07961_));
 sg13g2_a21oi_1 _27261_ (.A1(_07967_),
    .A2(_07968_),
    .Y(_01931_),
    .B1(net651));
 sg13g2_nand2_1 _27262_ (.Y(_07969_),
    .A(_10067_),
    .B(_07958_));
 sg13g2_nand2_1 _27263_ (.Y(_07970_),
    .A(\cpu.gpio.r_enable_in[4] ),
    .B(_07961_));
 sg13g2_a21oi_1 _27264_ (.A1(_07969_),
    .A2(_07970_),
    .Y(_01932_),
    .B1(net651));
 sg13g2_nand2_1 _27265_ (.Y(_07971_),
    .A(_10073_),
    .B(_07958_));
 sg13g2_nand2_1 _27266_ (.Y(_07972_),
    .A(\cpu.gpio.r_enable_in[5] ),
    .B(_07961_));
 sg13g2_a21oi_1 _27267_ (.A1(_07971_),
    .A2(_07972_),
    .Y(_01933_),
    .B1(net651));
 sg13g2_nand2_1 _27268_ (.Y(_07973_),
    .A(_10079_),
    .B(_07958_));
 sg13g2_nand2_1 _27269_ (.Y(_07974_),
    .A(\cpu.gpio.r_enable_in[6] ),
    .B(_07961_));
 sg13g2_a21oi_1 _27270_ (.A1(_07973_),
    .A2(_07974_),
    .Y(_01934_),
    .B1(net651));
 sg13g2_nand2_1 _27271_ (.Y(_07975_),
    .A(net1053),
    .B(_07958_));
 sg13g2_nand2_1 _27272_ (.Y(_07976_),
    .A(_09185_),
    .B(_07961_));
 sg13g2_a21oi_1 _27273_ (.A1(_07975_),
    .A2(_07976_),
    .Y(_01935_),
    .B1(net651));
 sg13g2_buf_1 _27274_ (.A(net112),
    .X(_07977_));
 sg13g2_nand3_1 _27275_ (.B(net404),
    .C(net101),
    .A(net1059),
    .Y(_07978_));
 sg13g2_nand2_1 _27276_ (.Y(_07979_),
    .A(net404),
    .B(net112));
 sg13g2_nand2_1 _27277_ (.Y(_07980_),
    .A(_09199_),
    .B(_07979_));
 sg13g2_buf_1 _27278_ (.A(_09330_),
    .X(_07981_));
 sg13g2_a21oi_1 _27279_ (.A1(_07978_),
    .A2(_07980_),
    .Y(_01936_),
    .B1(net647));
 sg13g2_nand3_1 _27280_ (.B(net404),
    .C(_07977_),
    .A(net1058),
    .Y(_07982_));
 sg13g2_nand2_1 _27281_ (.Y(_07983_),
    .A(_09194_),
    .B(_07979_));
 sg13g2_a21oi_1 _27282_ (.A1(_07982_),
    .A2(_07983_),
    .Y(_01937_),
    .B1(_07981_));
 sg13g2_nand3_1 _27283_ (.B(_05371_),
    .C(_07977_),
    .A(net1057),
    .Y(_07984_));
 sg13g2_nand2_1 _27284_ (.Y(_07985_),
    .A(_09187_),
    .B(_07979_));
 sg13g2_a21oi_1 _27285_ (.A1(_07984_),
    .A2(_07985_),
    .Y(_01938_),
    .B1(_07981_));
 sg13g2_nand3_1 _27286_ (.B(_05371_),
    .C(net101),
    .A(_10140_),
    .Y(_07986_));
 sg13g2_nand2_1 _27287_ (.Y(_07987_),
    .A(\cpu.gpio.r_enable_io[7] ),
    .B(_07979_));
 sg13g2_a21oi_1 _27288_ (.A1(_07986_),
    .A2(_07987_),
    .Y(_01939_),
    .B1(net647));
 sg13g2_nand3_1 _27289_ (.B(_05153_),
    .C(net112),
    .A(net982),
    .Y(_07988_));
 sg13g2_buf_2 _27290_ (.A(_07988_),
    .X(_07989_));
 sg13g2_mux2_1 _27291_ (.A0(_10066_),
    .A1(net7),
    .S(_07989_),
    .X(_07990_));
 sg13g2_and2_1 _27292_ (.A(net614),
    .B(_07990_),
    .X(_01940_));
 sg13g2_nand2_1 _27293_ (.Y(_07991_),
    .A(net8),
    .B(_07989_));
 sg13g2_o21ai_1 _27294_ (.B1(_07991_),
    .Y(_07992_),
    .A1(_12144_),
    .A2(_07989_));
 sg13g2_and2_1 _27295_ (.A(net614),
    .B(_07992_),
    .X(_01941_));
 sg13g2_mux2_1 _27296_ (.A0(_10078_),
    .A1(net9),
    .S(_07989_),
    .X(_07993_));
 sg13g2_and2_1 _27297_ (.A(net614),
    .B(_07993_),
    .X(_01942_));
 sg13g2_mux2_1 _27298_ (.A0(_10081_),
    .A1(net10),
    .S(_07989_),
    .X(_07994_));
 sg13g2_and2_1 _27299_ (.A(net614),
    .B(_07994_),
    .X(_01943_));
 sg13g2_nand3_1 _27300_ (.B(net408),
    .C(net101),
    .A(net1062),
    .Y(_07995_));
 sg13g2_nand2_1 _27301_ (.Y(_07996_),
    .A(_04909_),
    .B(net112));
 sg13g2_nand2_1 _27302_ (.Y(_07997_),
    .A(_04910_),
    .B(_07996_));
 sg13g2_nand3_1 _27303_ (.B(_07995_),
    .C(_07997_),
    .A(net634),
    .Y(_01989_));
 sg13g2_nand3_1 _27304_ (.B(net408),
    .C(net101),
    .A(_10051_),
    .Y(_07998_));
 sg13g2_buf_1 _27305_ (.A(\cpu.gpio.r_src_o[6][1] ),
    .X(_07999_));
 sg13g2_nand2_1 _27306_ (.Y(_08000_),
    .A(_07999_),
    .B(_07996_));
 sg13g2_a21oi_1 _27307_ (.A1(_07998_),
    .A2(_08000_),
    .Y(_01990_),
    .B1(net647));
 sg13g2_nand3_1 _27308_ (.B(net408),
    .C(net101),
    .A(_10056_),
    .Y(_08001_));
 sg13g2_nand2_1 _27309_ (.Y(_08002_),
    .A(\cpu.gpio.r_src_o[6][2] ),
    .B(_07996_));
 sg13g2_a21oi_1 _27310_ (.A1(_08001_),
    .A2(_08002_),
    .Y(_01991_),
    .B1(net647));
 sg13g2_nand3_1 _27311_ (.B(net408),
    .C(net101),
    .A(_06861_),
    .Y(_08003_));
 sg13g2_nand2_1 _27312_ (.Y(_08004_),
    .A(\cpu.gpio.r_src_o[6][3] ),
    .B(_07996_));
 sg13g2_a21oi_1 _27313_ (.A1(_08003_),
    .A2(_08004_),
    .Y(_01992_),
    .B1(net647));
 sg13g2_nand3_1 _27314_ (.B(net450),
    .C(net101),
    .A(net1062),
    .Y(_08005_));
 sg13g2_nand2_1 _27315_ (.Y(_08006_),
    .A(net450),
    .B(net112));
 sg13g2_nand2_1 _27316_ (.Y(_08007_),
    .A(_04927_),
    .B(_08006_));
 sg13g2_a21oi_1 _27317_ (.A1(_08005_),
    .A2(_08007_),
    .Y(_01997_),
    .B1(net647));
 sg13g2_nand3_1 _27318_ (.B(_04926_),
    .C(net101),
    .A(_10051_),
    .Y(_08008_));
 sg13g2_nand2_1 _27319_ (.Y(_08009_),
    .A(\cpu.gpio.r_uart_rx_src[1] ),
    .B(_08006_));
 sg13g2_a21oi_1 _27320_ (.A1(_08008_),
    .A2(_08009_),
    .Y(_01998_),
    .B1(net647));
 sg13g2_nand3_1 _27321_ (.B(_04926_),
    .C(_06412_),
    .A(net1060),
    .Y(_08010_));
 sg13g2_nand2_1 _27322_ (.Y(_08011_),
    .A(\cpu.gpio.r_uart_rx_src[2] ),
    .B(_08006_));
 sg13g2_a21oi_1 _27323_ (.A1(_08010_),
    .A2(_08011_),
    .Y(_01999_),
    .B1(net647));
 sg13g2_and2_1 _27324_ (.A(\cpu.i_wstrobe_d ),
    .B(_00304_),
    .X(_02256_));
 sg13g2_nor2_1 _27325_ (.A(_06468_),
    .B(_06480_),
    .Y(_08012_));
 sg13g2_nor2_1 _27326_ (.A(_06494_),
    .B(_08012_),
    .Y(_02257_));
 sg13g2_xor2_1 _27327_ (.B(_06475_),
    .A(\cpu.icache.r_offset[2] ),
    .X(_08013_));
 sg13g2_nor2_1 _27328_ (.A(_06494_),
    .B(_08013_),
    .Y(_02258_));
 sg13g2_xnor2_1 _27329_ (.Y(_08014_),
    .A(\cpu.intr.r_clock_cmp[31] ),
    .B(_05301_));
 sg13g2_xnor2_1 _27330_ (.Y(_08015_),
    .A(\cpu.intr.r_clock_cmp[1] ),
    .B(_10103_));
 sg13g2_xnor2_1 _27331_ (.Y(_08016_),
    .A(\cpu.intr.r_clock_cmp[21] ),
    .B(_05634_));
 sg13g2_xnor2_1 _27332_ (.Y(_08017_),
    .A(\cpu.intr.r_clock_cmp[14] ),
    .B(_10179_));
 sg13g2_nand4_1 _27333_ (.B(_08015_),
    .C(_08016_),
    .A(_08014_),
    .Y(_08018_),
    .D(_08017_));
 sg13g2_xnor2_1 _27334_ (.Y(_08019_),
    .A(\cpu.intr.r_clock_cmp[16] ),
    .B(_04945_));
 sg13g2_xnor2_1 _27335_ (.Y(_08020_),
    .A(\cpu.intr.r_clock_cmp[15] ),
    .B(_10184_));
 sg13g2_xnor2_1 _27336_ (.Y(_08021_),
    .A(\cpu.intr.r_clock_cmp[25] ),
    .B(_05767_));
 sg13g2_xnor2_1 _27337_ (.Y(_08022_),
    .A(\cpu.intr.r_clock_cmp[4] ),
    .B(_10127_));
 sg13g2_nand4_1 _27338_ (.B(_08020_),
    .C(_08021_),
    .A(_08019_),
    .Y(_08023_),
    .D(_08022_));
 sg13g2_xnor2_1 _27339_ (.Y(_08024_),
    .A(\cpu.intr.r_clock_cmp[3] ),
    .B(_10122_));
 sg13g2_xnor2_1 _27340_ (.Y(_08025_),
    .A(\cpu.intr.r_clock_cmp[23] ),
    .B(_05110_));
 sg13g2_xnor2_1 _27341_ (.Y(_08026_),
    .A(\cpu.intr.r_clock_cmp[11] ),
    .B(_10163_));
 sg13g2_xnor2_1 _27342_ (.Y(_08027_),
    .A(\cpu.intr.r_clock_cmp[27] ),
    .B(_05196_));
 sg13g2_nand4_1 _27343_ (.B(_08025_),
    .C(_08026_),
    .A(_08024_),
    .Y(_08028_),
    .D(_08027_));
 sg13g2_xnor2_1 _27344_ (.Y(_08029_),
    .A(\cpu.intr.r_clock_cmp[28] ),
    .B(_05208_));
 sg13g2_xnor2_1 _27345_ (.Y(_08030_),
    .A(\cpu.intr.r_clock_cmp[10] ),
    .B(_10158_));
 sg13g2_xnor2_1 _27346_ (.Y(_08031_),
    .A(\cpu.intr.r_clock_cmp[17] ),
    .B(_05384_));
 sg13g2_xnor2_1 _27347_ (.Y(_08032_),
    .A(\cpu.intr.r_clock_cmp[12] ),
    .B(_10169_));
 sg13g2_nand4_1 _27348_ (.B(_08030_),
    .C(_08031_),
    .A(_08029_),
    .Y(_08033_),
    .D(_08032_));
 sg13g2_nor4_1 _27349_ (.A(_08018_),
    .B(_08023_),
    .C(_08028_),
    .D(_08033_),
    .Y(_08034_));
 sg13g2_xnor2_1 _27350_ (.Y(_08035_),
    .A(\cpu.intr.r_clock_cmp[19] ),
    .B(_05506_));
 sg13g2_xnor2_1 _27351_ (.Y(_08036_),
    .A(\cpu.intr.r_clock_cmp[20] ),
    .B(_05541_));
 sg13g2_xnor2_1 _27352_ (.Y(_08037_),
    .A(\cpu.intr.r_clock_cmp[13] ),
    .B(_10173_));
 sg13g2_xnor2_1 _27353_ (.Y(_08038_),
    .A(\cpu.intr.r_clock_cmp[6] ),
    .B(_10136_));
 sg13g2_nand4_1 _27354_ (.B(_08036_),
    .C(_08037_),
    .A(_08035_),
    .Y(_08039_),
    .D(_08038_));
 sg13g2_xnor2_1 _27355_ (.Y(_08040_),
    .A(\cpu.intr.r_clock_cmp[8] ),
    .B(_10147_));
 sg13g2_xnor2_1 _27356_ (.Y(_08041_),
    .A(\cpu.intr.r_clock_cmp[7] ),
    .B(_10141_));
 sg13g2_xnor2_1 _27357_ (.Y(_08042_),
    .A(\cpu.intr.r_clock_cmp[22] ),
    .B(_05702_));
 sg13g2_xnor2_1 _27358_ (.Y(_08043_),
    .A(\cpu.intr.r_clock_cmp[30] ),
    .B(_05268_));
 sg13g2_nand4_1 _27359_ (.B(_08041_),
    .C(_08042_),
    .A(_08040_),
    .Y(_08044_),
    .D(_08043_));
 sg13g2_xnor2_1 _27360_ (.Y(_08045_),
    .A(\cpu.intr.r_clock_cmp[29] ),
    .B(_05239_));
 sg13g2_xnor2_1 _27361_ (.Y(_08046_),
    .A(\cpu.intr.r_clock_cmp[24] ),
    .B(_05752_));
 sg13g2_xnor2_1 _27362_ (.Y(_08047_),
    .A(\cpu.intr.r_clock_cmp[5] ),
    .B(_10132_));
 sg13g2_xnor2_1 _27363_ (.Y(_08048_),
    .A(\cpu.intr.r_clock_cmp[9] ),
    .B(_10153_));
 sg13g2_nand4_1 _27364_ (.B(_08046_),
    .C(_08047_),
    .A(_08045_),
    .Y(_08049_),
    .D(_08048_));
 sg13g2_xnor2_1 _27365_ (.Y(_08050_),
    .A(\cpu.intr.r_clock_cmp[2] ),
    .B(_10108_));
 sg13g2_xnor2_1 _27366_ (.Y(_08051_),
    .A(\cpu.intr.r_clock_cmp[0] ),
    .B(_10102_));
 sg13g2_xnor2_1 _27367_ (.Y(_08052_),
    .A(\cpu.intr.r_clock_cmp[26] ),
    .B(_05152_));
 sg13g2_xnor2_1 _27368_ (.Y(_08053_),
    .A(\cpu.intr.r_clock_cmp[18] ),
    .B(_05433_));
 sg13g2_nand4_1 _27369_ (.B(_08051_),
    .C(_08052_),
    .A(_08050_),
    .Y(_08054_),
    .D(_08053_));
 sg13g2_nor4_1 _27370_ (.A(_08039_),
    .B(_08044_),
    .C(_08049_),
    .D(_08054_),
    .Y(_08055_));
 sg13g2_a22oi_1 _27371_ (.Y(_08056_),
    .B1(_08034_),
    .B2(_08055_),
    .A2(_07645_),
    .A1(net1061));
 sg13g2_nand3_1 _27372_ (.B(net103),
    .C(net445),
    .A(net1061),
    .Y(_08057_));
 sg13g2_nand2_1 _27373_ (.Y(_08058_),
    .A(\cpu.intr.r_clock ),
    .B(_08057_));
 sg13g2_buf_1 _27374_ (.A(_09330_),
    .X(_08059_));
 sg13g2_a21oi_1 _27375_ (.A1(_08056_),
    .A2(_08058_),
    .Y(_02419_),
    .B1(net646));
 sg13g2_and2_1 _27376_ (.A(net103),
    .B(net448),
    .X(_08060_));
 sg13g2_buf_1 _27377_ (.A(_08060_),
    .X(_08061_));
 sg13g2_nand2_1 _27378_ (.Y(_08062_),
    .A(net874),
    .B(_08061_));
 sg13g2_nand2_1 _27379_ (.Y(_08063_),
    .A(_06757_),
    .B(net448));
 sg13g2_buf_1 _27380_ (.A(_08063_),
    .X(_08064_));
 sg13g2_nand2_1 _27381_ (.Y(_08065_),
    .A(_09167_),
    .B(_08064_));
 sg13g2_a21oi_1 _27382_ (.A1(_08062_),
    .A2(_08065_),
    .Y(_02468_),
    .B1(_08059_));
 sg13g2_nand2_1 _27383_ (.Y(_08066_),
    .A(net1055),
    .B(_08061_));
 sg13g2_nand2_1 _27384_ (.Y(_08067_),
    .A(_09169_),
    .B(_08064_));
 sg13g2_a21oi_1 _27385_ (.A1(_08066_),
    .A2(_08067_),
    .Y(_02469_),
    .B1(_08059_));
 sg13g2_nand2_1 _27386_ (.Y(_08068_),
    .A(net910),
    .B(_08061_));
 sg13g2_nand2_1 _27387_ (.Y(_08069_),
    .A(_09162_),
    .B(_08064_));
 sg13g2_a21oi_1 _27388_ (.A1(_08068_),
    .A2(_08069_),
    .Y(_02470_),
    .B1(net646));
 sg13g2_nand2_1 _27389_ (.Y(_08070_),
    .A(net954),
    .B(_08061_));
 sg13g2_nand2_1 _27390_ (.Y(_08071_),
    .A(\cpu.intr.r_enable[3] ),
    .B(_08064_));
 sg13g2_a21oi_1 _27391_ (.A1(_08070_),
    .A2(_08071_),
    .Y(_02471_),
    .B1(net646));
 sg13g2_nand2_1 _27392_ (.Y(_08072_),
    .A(net1059),
    .B(_08061_));
 sg13g2_nand2_1 _27393_ (.Y(_08073_),
    .A(_09203_),
    .B(_08064_));
 sg13g2_a21oi_1 _27394_ (.A1(_08072_),
    .A2(_08073_),
    .Y(_02472_),
    .B1(net646));
 sg13g2_nand2_1 _27395_ (.Y(_08074_),
    .A(net1058),
    .B(_08061_));
 sg13g2_nand2_1 _27396_ (.Y(_08075_),
    .A(\cpu.intr.r_enable[5] ),
    .B(_08064_));
 sg13g2_a21oi_1 _27397_ (.A1(_08074_),
    .A2(_08075_),
    .Y(_02473_),
    .B1(net646));
 sg13g2_nand3_1 _27398_ (.B(_06757_),
    .C(net445),
    .A(net1060),
    .Y(_08076_));
 sg13g2_inv_1 _27399_ (.Y(_08077_),
    .A(_09990_));
 sg13g2_a221oi_1 _27400_ (.B2(_09161_),
    .C1(_08077_),
    .B1(_08076_),
    .A1(net1060),
    .Y(_08078_),
    .A2(_07645_));
 sg13g2_nor2_1 _27401_ (.A(net704),
    .B(_08078_),
    .Y(_02474_));
 sg13g2_nor3_2 _27402_ (.A(_09888_),
    .B(_09846_),
    .C(_06931_),
    .Y(_08079_));
 sg13g2_nand4_1 _27403_ (.B(_06893_),
    .C(_06932_),
    .A(_09872_),
    .Y(_08080_),
    .D(_08079_));
 sg13g2_buf_1 _27404_ (.A(_08080_),
    .X(_08081_));
 sg13g2_a21o_1 _27405_ (.A2(_06839_),
    .A1(_09848_),
    .B1(_08081_),
    .X(_08082_));
 sg13g2_o21ai_1 _27406_ (.B1(net803),
    .Y(_08083_),
    .A1(_06894_),
    .A2(_08081_));
 sg13g2_a21o_1 _27407_ (.A2(_08082_),
    .A1(net19),
    .B1(_08083_),
    .X(_02504_));
 sg13g2_nand3b_1 _27408_ (.B(_06936_),
    .C(_09828_),
    .Y(_08084_),
    .A_N(_09848_));
 sg13g2_a21o_1 _27409_ (.A2(_08084_),
    .A1(_06894_),
    .B1(_08081_),
    .X(_08085_));
 sg13g2_nand2_1 _27410_ (.Y(_08086_),
    .A(_09848_),
    .B(_06894_));
 sg13g2_nor2_1 _27411_ (.A(net81),
    .B(_08086_),
    .Y(_08087_));
 sg13g2_o21ai_1 _27412_ (.B1(net20),
    .Y(_08088_),
    .A1(_08081_),
    .A2(_08087_));
 sg13g2_nand3_1 _27413_ (.B(_08085_),
    .C(_08088_),
    .A(net634),
    .Y(_02505_));
 sg13g2_nor2b_1 _27414_ (.A(_09865_),
    .B_N(_09848_),
    .Y(_08089_));
 sg13g2_buf_1 _27415_ (.A(\cpu.gpio.genblk1[3].srcs_o[11] ),
    .X(_08090_));
 sg13g2_o21ai_1 _27416_ (.B1(_08090_),
    .Y(_08091_),
    .A1(_08081_),
    .A2(_08089_));
 sg13g2_nand2b_1 _27417_ (.Y(_02506_),
    .B(_08091_),
    .A_N(_08083_));
 sg13g2_nor4_1 _27418_ (.A(\cpu.qspi.r_state[17] ),
    .B(_09838_),
    .C(net1064),
    .D(_06936_),
    .Y(_08092_));
 sg13g2_nand2_1 _27419_ (.Y(_08093_),
    .A(_06804_),
    .B(_08092_));
 sg13g2_nor3_1 _27420_ (.A(_09839_),
    .B(_09873_),
    .C(_08093_),
    .Y(_08094_));
 sg13g2_a21oi_1 _27421_ (.A1(_08079_),
    .A2(_08094_),
    .Y(_08095_),
    .B1(_09828_));
 sg13g2_nor2_1 _27422_ (.A(net704),
    .B(_08095_),
    .Y(_02507_));
 sg13g2_nand2_1 _27423_ (.Y(_08096_),
    .A(net1053),
    .B(_06852_));
 sg13g2_nand2_1 _27424_ (.Y(_08097_),
    .A(\cpu.qspi.r_mask[0] ),
    .B(_06855_));
 sg13g2_a21oi_1 _27425_ (.A1(_08096_),
    .A2(_08097_),
    .Y(_02508_),
    .B1(net646));
 sg13g2_nor3_1 _27426_ (.A(net983),
    .B(_04950_),
    .C(_06865_),
    .Y(_08098_));
 sg13g2_inv_1 _27427_ (.Y(_08099_),
    .A(_07312_));
 sg13g2_a22oi_1 _27428_ (.Y(_08100_),
    .B1(_08098_),
    .B2(_08099_),
    .A2(_06869_),
    .A1(\cpu.qspi.r_mask[1] ));
 sg13g2_nand2_1 _27429_ (.Y(_02509_),
    .A(net591),
    .B(_08100_));
 sg13g2_nor2_1 _27430_ (.A(_07312_),
    .B(_06881_),
    .Y(_08101_));
 sg13g2_a21oi_1 _27431_ (.A1(\cpu.qspi.r_mask[2] ),
    .A2(_06881_),
    .Y(_08102_),
    .B1(_08101_));
 sg13g2_nor2_1 _27432_ (.A(_09331_),
    .B(_08102_),
    .Y(_02510_));
 sg13g2_nand2_1 _27433_ (.Y(_08103_),
    .A(\cpu.qspi.r_quad[0] ),
    .B(_06855_));
 sg13g2_nand2_1 _27434_ (.Y(_08104_),
    .A(net1057),
    .B(_06852_));
 sg13g2_nand3_1 _27435_ (.B(_08103_),
    .C(_08104_),
    .A(net634),
    .Y(_02511_));
 sg13g2_a22oi_1 _27436_ (.Y(_08105_),
    .B1(_08098_),
    .B2(_07307_),
    .A2(_06869_),
    .A1(\cpu.qspi.r_quad[1] ));
 sg13g2_nor2_1 _27437_ (.A(_09331_),
    .B(_08105_),
    .Y(_02512_));
 sg13g2_nand2_1 _27438_ (.Y(_08106_),
    .A(_00172_),
    .B(_06878_));
 sg13g2_o21ai_1 _27439_ (.B1(_08106_),
    .Y(_08107_),
    .A1(\cpu.qspi.r_quad[2] ),
    .A2(_06878_));
 sg13g2_nand2_1 _27440_ (.Y(_02513_),
    .A(net591),
    .B(_08107_));
 sg13g2_nand3_1 _27441_ (.B(net558),
    .C(_06850_),
    .A(net550),
    .Y(_08108_));
 sg13g2_mux2_1 _27442_ (.A0(net1062),
    .A1(_09856_),
    .S(_08108_),
    .X(_08109_));
 sg13g2_nand2b_1 _27443_ (.Y(_02526_),
    .B(net591),
    .A_N(_08109_));
 sg13g2_mux2_1 _27444_ (.A0(net1061),
    .A1(_09855_),
    .S(_08108_),
    .X(_08110_));
 sg13g2_nand2b_1 _27445_ (.Y(_02527_),
    .B(net591),
    .A_N(_08110_));
 sg13g2_a21o_1 _27446_ (.A2(_06891_),
    .A1(_06890_),
    .B1(_11917_),
    .X(_08111_));
 sg13g2_nor4_1 _27447_ (.A(_11938_),
    .B(_09838_),
    .C(net1064),
    .D(_09886_),
    .Y(_08112_));
 sg13g2_nand4_1 _27448_ (.B(_08079_),
    .C(_08111_),
    .A(_09826_),
    .Y(_08113_),
    .D(_08112_));
 sg13g2_buf_1 _27449_ (.A(_08113_),
    .X(_08114_));
 sg13g2_nor2b_1 _27450_ (.A(net3),
    .B_N(_08114_),
    .Y(_08115_));
 sg13g2_nor4_1 _27451_ (.A(_11916_),
    .B(_09839_),
    .C(_09827_),
    .D(_09873_),
    .Y(_08116_));
 sg13g2_nor4_1 _27452_ (.A(_11914_),
    .B(_06936_),
    .C(_08114_),
    .D(_08116_),
    .Y(_08117_));
 sg13g2_nor3_1 _27453_ (.A(net800),
    .B(_08115_),
    .C(_08117_),
    .Y(_02528_));
 sg13g2_nor2b_1 _27454_ (.A(net6),
    .B_N(_08114_),
    .Y(_08118_));
 sg13g2_nand2b_1 _27455_ (.Y(_08119_),
    .B(_08116_),
    .A_N(_06936_));
 sg13g2_o21ai_1 _27456_ (.B1(_11915_),
    .Y(_08120_),
    .A1(_09869_),
    .A2(_08119_));
 sg13g2_nor2_1 _27457_ (.A(_08114_),
    .B(_08120_),
    .Y(_08121_));
 sg13g2_nor3_1 _27458_ (.A(net800),
    .B(_08118_),
    .C(_08121_),
    .Y(_02529_));
 sg13g2_nor3_1 _27459_ (.A(_09251_),
    .B(net1137),
    .C(_09325_),
    .Y(_08122_));
 sg13g2_a221oi_1 _27460_ (.B2(net1071),
    .C1(_08122_),
    .B1(_09309_),
    .A1(_09289_),
    .Y(_08123_),
    .A2(_09249_));
 sg13g2_buf_1 _27461_ (.A(_08123_),
    .X(_08124_));
 sg13g2_nand3_1 _27462_ (.B(net1071),
    .C(_08124_),
    .A(_09253_),
    .Y(_08125_));
 sg13g2_o21ai_1 _27463_ (.B1(_08125_),
    .Y(_08126_),
    .A1(_09253_),
    .A2(_08124_));
 sg13g2_nand2_1 _27464_ (.Y(_02535_),
    .A(net591),
    .B(_08126_));
 sg13g2_nand2_1 _27465_ (.Y(_08127_),
    .A(_09253_),
    .B(_11949_));
 sg13g2_a21oi_1 _27466_ (.A1(_08124_),
    .A2(_08127_),
    .Y(_08128_),
    .B1(_09254_));
 sg13g2_inv_1 _27467_ (.Y(_08129_),
    .A(_09253_));
 sg13g2_and4_1 _27468_ (.A(_08129_),
    .B(_09254_),
    .C(_11949_),
    .D(_08124_),
    .X(_08130_));
 sg13g2_o21ai_1 _27469_ (.B1(net591),
    .Y(_02536_),
    .A1(_08128_),
    .A2(_08130_));
 sg13g2_nor2_1 _27470_ (.A(_09253_),
    .B(_09254_),
    .Y(_08131_));
 sg13g2_or2_1 _27471_ (.X(_08132_),
    .B(_08131_),
    .A(_00211_));
 sg13g2_a21oi_1 _27472_ (.A1(_08124_),
    .A2(_08132_),
    .Y(_08133_),
    .B1(\cpu.spi.r_bits[2] ));
 sg13g2_and4_1 _27473_ (.A(\cpu.spi.r_bits[2] ),
    .B(_11949_),
    .C(_08131_),
    .D(_08124_),
    .X(_08134_));
 sg13g2_o21ai_1 _27474_ (.B1(net591),
    .Y(_02537_),
    .A1(_08133_),
    .A2(_08134_));
 sg13g2_o21ai_1 _27475_ (.B1(net517),
    .Y(_08135_),
    .A1(net1137),
    .A2(_09321_));
 sg13g2_nand2_1 _27476_ (.Y(_08136_),
    .A(_09237_),
    .B(_09249_));
 sg13g2_nor4_1 _27477_ (.A(net1137),
    .B(net1135),
    .C(_09321_),
    .D(net517),
    .Y(_08137_));
 sg13g2_a21oi_1 _27478_ (.A1(net951),
    .A2(net1031),
    .Y(_08138_),
    .B1(_09308_));
 sg13g2_nor3_1 _27479_ (.A(_00262_),
    .B(_08137_),
    .C(_08138_),
    .Y(_08139_));
 sg13g2_a221oi_1 _27480_ (.B2(_07080_),
    .C1(_08139_),
    .B1(_08136_),
    .A1(_00262_),
    .Y(_08140_),
    .A2(_08135_));
 sg13g2_buf_1 _27481_ (.A(_08140_),
    .X(_08141_));
 sg13g2_o21ai_1 _27482_ (.B1(_08141_),
    .Y(_08142_),
    .A1(_12000_),
    .A2(_09321_));
 sg13g2_nand2_1 _27483_ (.Y(_08143_),
    .A(net803),
    .B(_08142_));
 sg13g2_nand2b_1 _27484_ (.Y(_08144_),
    .B(_08141_),
    .A_N(_11967_));
 sg13g2_buf_1 _27485_ (.A(\cpu.gpio.genblk1[3].srcs_o[6] ),
    .X(_08145_));
 sg13g2_o21ai_1 _27486_ (.B1(net1093),
    .Y(_08146_),
    .A1(_11952_),
    .A2(_08144_));
 sg13g2_nand2b_1 _27487_ (.Y(_02570_),
    .B(_08146_),
    .A_N(_08143_));
 sg13g2_buf_1 _27488_ (.A(\cpu.gpio.genblk1[3].srcs_o[7] ),
    .X(_08147_));
 sg13g2_nand3_1 _27489_ (.B(_11967_),
    .C(_08141_),
    .A(_11964_),
    .Y(_08148_));
 sg13g2_a21o_1 _27490_ (.A2(_08148_),
    .A1(net1092),
    .B1(_08143_),
    .X(_02571_));
 sg13g2_buf_1 _27491_ (.A(\cpu.gpio.genblk1[3].srcs_o[8] ),
    .X(_08149_));
 sg13g2_o21ai_1 _27492_ (.B1(net1091),
    .Y(_08150_),
    .A1(_11964_),
    .A2(_08144_));
 sg13g2_nand2b_1 _27493_ (.Y(_02572_),
    .B(_08150_),
    .A_N(_08143_));
 sg13g2_or3_1 _27494_ (.A(_07077_),
    .B(_09237_),
    .C(_09302_),
    .X(_08151_));
 sg13g2_nand2_1 _27495_ (.Y(_08152_),
    .A(_09276_),
    .B(net517));
 sg13g2_a21oi_1 _27496_ (.A1(net1071),
    .A2(_08152_),
    .Y(_08153_),
    .B1(_08122_));
 sg13g2_nand3_1 _27497_ (.B(_08151_),
    .C(_08153_),
    .A(_09357_),
    .Y(_08154_));
 sg13g2_nand2_1 _27498_ (.Y(_08155_),
    .A(_09170_),
    .B(_08154_));
 sg13g2_o21ai_1 _27499_ (.B1(_08155_),
    .Y(_08156_),
    .A1(_09304_),
    .A2(_08154_));
 sg13g2_and2_1 _27500_ (.A(net614),
    .B(_08156_),
    .X(_02581_));
 sg13g2_inv_1 _27501_ (.Y(_08157_),
    .A(\cpu.spi.r_ready ));
 sg13g2_nor4_1 _27502_ (.A(_09251_),
    .B(net1137),
    .C(_09321_),
    .D(_09325_),
    .Y(_08158_));
 sg13g2_a21oi_1 _27503_ (.A1(net1071),
    .A2(_08152_),
    .Y(_08159_),
    .B1(_08158_));
 sg13g2_and3_1 _27504_ (.X(_08160_),
    .A(_09357_),
    .B(_08151_),
    .C(_08159_));
 sg13g2_nor2_1 _27505_ (.A(_09321_),
    .B(_09320_),
    .Y(_08161_));
 sg13g2_a22oi_1 _27506_ (.Y(_08162_),
    .B1(_08160_),
    .B2(_08161_),
    .A2(net422),
    .A1(_08157_));
 sg13g2_nor2_1 _27507_ (.A(net1071),
    .B(_08162_),
    .Y(_08163_));
 sg13g2_nor2_1 _27508_ (.A(\cpu.spi.r_ready ),
    .B(_08160_),
    .Y(_08164_));
 sg13g2_o21ai_1 _27509_ (.B1(net591),
    .Y(_02596_),
    .A1(_08163_),
    .A2(_08164_));
 sg13g2_nand2_1 _27510_ (.Y(_08165_),
    .A(_09250_),
    .B(_08153_));
 sg13g2_nand2_1 _27511_ (.Y(_08166_),
    .A(\cpu.spi.r_searching ),
    .B(_08165_));
 sg13g2_nand4_1 _27512_ (.B(_09236_),
    .C(_09250_),
    .A(_07080_),
    .Y(_08167_),
    .D(_08153_));
 sg13g2_a21oi_1 _27513_ (.A1(_08166_),
    .A2(_08167_),
    .Y(_02597_),
    .B1(net646));
 sg13g2_and2_1 _27514_ (.A(_04962_),
    .B(_07388_),
    .X(_08168_));
 sg13g2_buf_2 _27515_ (.A(_08168_),
    .X(_08169_));
 sg13g2_nand2_1 _27516_ (.Y(_08170_),
    .A(net874),
    .B(_08169_));
 sg13g2_nand2_1 _27517_ (.Y(_08171_),
    .A(_04962_),
    .B(_07388_));
 sg13g2_buf_2 _27518_ (.A(_08171_),
    .X(_08172_));
 sg13g2_nand2_1 _27519_ (.Y(_08173_),
    .A(\cpu.uart.r_div_value[0] ),
    .B(_08172_));
 sg13g2_nand3_1 _27520_ (.B(_08170_),
    .C(_08173_),
    .A(net634),
    .Y(_02619_));
 sg13g2_and2_1 _27521_ (.A(net445),
    .B(_07388_),
    .X(_08174_));
 sg13g2_buf_2 _27522_ (.A(_08174_),
    .X(_08175_));
 sg13g2_nand2_1 _27523_ (.Y(_08176_),
    .A(net910),
    .B(_08175_));
 sg13g2_nand2b_1 _27524_ (.Y(_08177_),
    .B(_09933_),
    .A_N(_08175_));
 sg13g2_a21oi_1 _27525_ (.A1(_08176_),
    .A2(_08177_),
    .Y(_02620_),
    .B1(net646));
 sg13g2_nand2_1 _27526_ (.Y(_08178_),
    .A(net954),
    .B(_08175_));
 sg13g2_nand2b_1 _27527_ (.Y(_08179_),
    .B(\cpu.uart.r_div_value[11] ),
    .A_N(_08175_));
 sg13g2_buf_1 _27528_ (.A(_09330_),
    .X(_08180_));
 sg13g2_a21oi_1 _27529_ (.A1(_08178_),
    .A2(_08179_),
    .Y(_02621_),
    .B1(net645));
 sg13g2_nand2_1 _27530_ (.Y(_08181_),
    .A(net1055),
    .B(_08169_));
 sg13g2_nand2_1 _27531_ (.Y(_08182_),
    .A(\cpu.uart.r_div_value[1] ),
    .B(_08172_));
 sg13g2_a21oi_1 _27532_ (.A1(_08181_),
    .A2(_08182_),
    .Y(_02622_),
    .B1(net645));
 sg13g2_nand2_1 _27533_ (.Y(_08183_),
    .A(net910),
    .B(_08169_));
 sg13g2_nand2_1 _27534_ (.Y(_08184_),
    .A(\cpu.uart.r_div_value[2] ),
    .B(_08172_));
 sg13g2_a21oi_1 _27535_ (.A1(_08183_),
    .A2(_08184_),
    .Y(_02623_),
    .B1(_08180_));
 sg13g2_nand2_1 _27536_ (.Y(_08185_),
    .A(net954),
    .B(_08169_));
 sg13g2_nand2_1 _27537_ (.Y(_08186_),
    .A(\cpu.uart.r_div_value[3] ),
    .B(_08172_));
 sg13g2_a21oi_1 _27538_ (.A1(_08185_),
    .A2(_08186_),
    .Y(_02624_),
    .B1(net645));
 sg13g2_nand2_1 _27539_ (.Y(_08187_),
    .A(net1059),
    .B(_08169_));
 sg13g2_nand2_1 _27540_ (.Y(_08188_),
    .A(\cpu.uart.r_div_value[4] ),
    .B(_08172_));
 sg13g2_a21oi_1 _27541_ (.A1(_08187_),
    .A2(_08188_),
    .Y(_02625_),
    .B1(net645));
 sg13g2_nand2_1 _27542_ (.Y(_08189_),
    .A(_10073_),
    .B(_08169_));
 sg13g2_nand2_1 _27543_ (.Y(_08190_),
    .A(\cpu.uart.r_div_value[5] ),
    .B(_08172_));
 sg13g2_a21oi_1 _27544_ (.A1(_08189_),
    .A2(_08190_),
    .Y(_02626_),
    .B1(net645));
 sg13g2_nand2_1 _27545_ (.Y(_08191_),
    .A(net1057),
    .B(_08169_));
 sg13g2_nand2_1 _27546_ (.Y(_08192_),
    .A(\cpu.uart.r_div_value[6] ),
    .B(_08172_));
 sg13g2_a21oi_1 _27547_ (.A1(_08191_),
    .A2(_08192_),
    .Y(_02627_),
    .B1(net645));
 sg13g2_nand2_1 _27548_ (.Y(_08193_),
    .A(_10140_),
    .B(_08169_));
 sg13g2_nand2_1 _27549_ (.Y(_08194_),
    .A(\cpu.uart.r_div_value[7] ),
    .B(_08172_));
 sg13g2_a21oi_1 _27550_ (.A1(_08193_),
    .A2(_08194_),
    .Y(_02628_),
    .B1(_08180_));
 sg13g2_nand2_1 _27551_ (.Y(_08195_),
    .A(net1062),
    .B(_08175_));
 sg13g2_nand2b_1 _27552_ (.Y(_08196_),
    .B(\cpu.uart.r_div_value[8] ),
    .A_N(_08175_));
 sg13g2_a21oi_1 _27553_ (.A1(_08195_),
    .A2(_08196_),
    .Y(_02629_),
    .B1(net645));
 sg13g2_nand2_1 _27554_ (.Y(_08197_),
    .A(net1055),
    .B(_08175_));
 sg13g2_nand2b_1 _27555_ (.Y(_08198_),
    .B(\cpu.uart.r_div_value[9] ),
    .A_N(_08175_));
 sg13g2_a21oi_1 _27556_ (.A1(_08197_),
    .A2(_08198_),
    .Y(_02630_),
    .B1(net645));
 sg13g2_nand3_1 _27557_ (.B(_04946_),
    .C(_07388_),
    .A(_10050_),
    .Y(_08199_));
 sg13g2_nor2_1 _27558_ (.A(net1000),
    .B(net463),
    .Y(_08200_));
 sg13g2_nand3_1 _27559_ (.B(_07386_),
    .C(_08200_),
    .A(_08455_),
    .Y(_08201_));
 sg13g2_or4_1 _27560_ (.A(net550),
    .B(_09212_),
    .C(_07073_),
    .D(_08201_),
    .X(_08202_));
 sg13g2_nand4_1 _27561_ (.B(net708),
    .C(_08199_),
    .A(_09166_),
    .Y(_08203_),
    .D(_08202_));
 sg13g2_nand2b_1 _27562_ (.Y(_02654_),
    .B(_08203_),
    .A_N(net129));
 sg13g2_and2_1 _27563_ (.A(net487),
    .B(_07388_),
    .X(_08204_));
 sg13g2_buf_1 _27564_ (.A(_08204_),
    .X(_08205_));
 sg13g2_nand2_1 _27565_ (.Y(_08206_),
    .A(net1055),
    .B(_08205_));
 sg13g2_nand2b_1 _27566_ (.Y(_08207_),
    .B(\cpu.uart.r_r_invert ),
    .A_N(_08205_));
 sg13g2_a21oi_1 _27567_ (.A1(_08206_),
    .A2(_08207_),
    .Y(_02655_),
    .B1(net782));
 sg13g2_a21oi_1 _27568_ (.A1(_07376_),
    .A2(_09911_),
    .Y(_08208_),
    .B1(net1098));
 sg13g2_a21oi_1 _27569_ (.A1(_07377_),
    .A2(_09911_),
    .Y(_08209_),
    .B1(_07449_));
 sg13g2_a221oi_1 _27570_ (.B2(_08208_),
    .C1(_08209_),
    .B1(_07375_),
    .A1(net949),
    .Y(_08210_),
    .A2(net1098));
 sg13g2_a21oi_1 _27571_ (.A1(_07368_),
    .A2(_08210_),
    .Y(_08211_),
    .B1(_07446_));
 sg13g2_buf_2 _27572_ (.A(_08211_),
    .X(_08212_));
 sg13g2_o21ai_1 _27573_ (.B1(_08212_),
    .Y(_08213_),
    .A1(net949),
    .A2(_07449_));
 sg13g2_xnor2_1 _27574_ (.Y(_08214_),
    .A(_07377_),
    .B(_08213_));
 sg13g2_nor2_1 _27575_ (.A(net704),
    .B(_08214_),
    .Y(_02658_));
 sg13g2_o21ai_1 _27576_ (.B1(_08212_),
    .Y(_08215_),
    .A1(_07376_),
    .A2(net950));
 sg13g2_nand2_1 _27577_ (.Y(_08216_),
    .A(_07372_),
    .B(_08215_));
 sg13g2_nand2b_1 _27578_ (.Y(_08217_),
    .B(_07374_),
    .A_N(_07371_));
 sg13g2_o21ai_1 _27579_ (.B1(_08217_),
    .Y(_08218_),
    .A1(_07374_),
    .A2(_07448_));
 sg13g2_nand3_1 _27580_ (.B(_08212_),
    .C(_08218_),
    .A(_07447_),
    .Y(_08219_));
 sg13g2_a21oi_1 _27581_ (.A1(_08216_),
    .A2(_08219_),
    .Y(_02659_),
    .B1(net782));
 sg13g2_nand2_1 _27582_ (.Y(_08220_),
    .A(_07376_),
    .B(net1097));
 sg13g2_nor3_1 _27583_ (.A(net949),
    .B(net950),
    .C(_08220_),
    .Y(_08221_));
 sg13g2_o21ai_1 _27584_ (.B1(_08212_),
    .Y(_08222_),
    .A1(net950),
    .A2(_07457_));
 sg13g2_a22oi_1 _27585_ (.Y(_08223_),
    .B1(_08222_),
    .B2(net949),
    .A2(_08221_),
    .A1(_08212_));
 sg13g2_nor2_1 _27586_ (.A(net704),
    .B(_08223_),
    .Y(_02660_));
 sg13g2_a21oi_1 _27587_ (.A1(_07457_),
    .A2(_08212_),
    .Y(_08224_),
    .B1(net950));
 sg13g2_nor2b_1 _27588_ (.A(net949),
    .B_N(net1097),
    .Y(_08225_));
 sg13g2_a21oi_1 _27589_ (.A1(_08212_),
    .A2(_08225_),
    .Y(_08226_),
    .B1(_09852_));
 sg13g2_nor2b_1 _27590_ (.A(_08224_),
    .B_N(_08226_),
    .Y(_02661_));
 sg13g2_nor2b_1 _27591_ (.A(_07474_),
    .B_N(_07479_),
    .Y(_08227_));
 sg13g2_o21ai_1 _27592_ (.B1(_06864_),
    .Y(_08228_),
    .A1(_00208_),
    .A2(_04886_));
 sg13g2_nand4_1 _27593_ (.B(_07414_),
    .C(_07492_),
    .A(_09581_),
    .Y(_08229_),
    .D(_08228_));
 sg13g2_a221oi_1 _27594_ (.B2(_10032_),
    .C1(_07479_),
    .B1(_04946_),
    .A1(_09581_),
    .Y(_08230_),
    .A2(_10112_));
 sg13g2_a21oi_1 _27595_ (.A1(_07474_),
    .A2(_08229_),
    .Y(_08231_),
    .B1(_08230_));
 sg13g2_a21o_1 _27596_ (.A2(_08231_),
    .A1(_07408_),
    .B1(_09165_),
    .X(_08232_));
 sg13g2_nand2_1 _27597_ (.Y(_08233_),
    .A(_07388_),
    .B(_08231_));
 sg13g2_a22oi_1 _27598_ (.Y(_08234_),
    .B1(_08233_),
    .B2(_09165_),
    .A2(_08232_),
    .A1(_08227_));
 sg13g2_nor2_1 _27599_ (.A(net704),
    .B(_08234_),
    .Y(_02663_));
 sg13g2_nand2_1 _27600_ (.Y(_08235_),
    .A(net1062),
    .B(_08205_));
 sg13g2_nand2b_1 _27601_ (.Y(_08236_),
    .B(\cpu.uart.r_x_invert ),
    .A_N(_08205_));
 sg13g2_a21oi_1 _27602_ (.A1(_08235_),
    .A2(_08236_),
    .Y(_02664_),
    .B1(net782));
 sg13g2_a21oi_1 _27603_ (.A1(_07403_),
    .A2(_07468_),
    .Y(_08237_),
    .B1(net1096));
 sg13g2_o21ai_1 _27604_ (.B1(net827),
    .Y(_08238_),
    .A1(_07482_),
    .A2(_08237_));
 sg13g2_o21ai_1 _27605_ (.B1(_07493_),
    .Y(_08239_),
    .A1(_07408_),
    .A2(_07479_));
 sg13g2_a22oi_1 _27606_ (.Y(_08240_),
    .B1(_08239_),
    .B2(_07389_),
    .A2(_08238_),
    .A1(_07485_));
 sg13g2_buf_2 _27607_ (.A(_08240_),
    .X(_08241_));
 sg13g2_nand2_1 _27608_ (.Y(_08242_),
    .A(_07408_),
    .B(_07480_));
 sg13g2_nand4_1 _27609_ (.B(_07470_),
    .C(_08241_),
    .A(net1096),
    .Y(_08243_),
    .D(_08242_));
 sg13g2_o21ai_1 _27610_ (.B1(_08243_),
    .Y(_08244_),
    .A1(net1096),
    .A2(_08241_));
 sg13g2_nor2_1 _27611_ (.A(net704),
    .B(_08244_),
    .Y(_02667_));
 sg13g2_nand2_1 _27612_ (.Y(_08245_),
    .A(_07394_),
    .B(_07470_));
 sg13g2_a21o_1 _27613_ (.A2(_08245_),
    .A1(_08241_),
    .B1(_07392_),
    .X(_08246_));
 sg13g2_nand4_1 _27614_ (.B(net1096),
    .C(_07470_),
    .A(_07392_),
    .Y(_08247_),
    .D(_08241_));
 sg13g2_a21oi_1 _27615_ (.A1(_08246_),
    .A2(_08247_),
    .Y(_02668_),
    .B1(net782));
 sg13g2_o21ai_1 _27616_ (.B1(_08241_),
    .Y(_08248_),
    .A1(_07395_),
    .A2(_07478_));
 sg13g2_nand2_1 _27617_ (.Y(_08249_),
    .A(_07385_),
    .B(_08248_));
 sg13g2_nand2_1 _27618_ (.Y(_08250_),
    .A(_07403_),
    .B(_07480_));
 sg13g2_o21ai_1 _27619_ (.B1(_08250_),
    .Y(_08251_),
    .A1(_07394_),
    .A2(_07395_));
 sg13g2_nand4_1 _27620_ (.B(_07405_),
    .C(_08241_),
    .A(_07390_),
    .Y(_08252_),
    .D(_08251_));
 sg13g2_a21oi_1 _27621_ (.A1(_08249_),
    .A2(_08252_),
    .Y(_02669_),
    .B1(net782));
 sg13g2_nand3_1 _27622_ (.B(_07478_),
    .C(_08250_),
    .A(_07405_),
    .Y(_08253_));
 sg13g2_nand2_1 _27623_ (.Y(_08254_),
    .A(_07470_),
    .B(_08253_));
 sg13g2_nand2_1 _27624_ (.Y(_08255_),
    .A(_07478_),
    .B(_08241_));
 sg13g2_a221oi_1 _27625_ (.B2(_07396_),
    .C1(net782),
    .B1(_08255_),
    .A1(_08241_),
    .Y(_02670_),
    .A2(_08254_));
 sg13g2_nand2b_1 _27626_ (.Y(\cpu.ex.genblk3.c_supmode ),
    .B(_07657_),
    .A_N(_07653_));
 sg13g2_nor3_1 _27627_ (.A(_09888_),
    .B(_09827_),
    .C(_06931_),
    .Y(_08256_));
 sg13g2_and3_1 _27628_ (.X(_08257_),
    .A(net111),
    .B(_08094_),
    .C(_08256_));
 sg13g2_a21oi_1 _27629_ (.A1(_09841_),
    .A2(net624),
    .Y(_08258_),
    .B1(_08257_));
 sg13g2_inv_1 _27630_ (.Y(\cpu.qspi.c_rstrobe_d ),
    .A(_08258_));
 sg13g2_nor4_1 _27631_ (.A(_09839_),
    .B(_09827_),
    .C(net624),
    .D(_08093_),
    .Y(_08259_));
 sg13g2_a22oi_1 _27632_ (.Y(_08260_),
    .B1(_08079_),
    .B2(_08259_),
    .A2(net624),
    .A1(_09838_));
 sg13g2_nor2_1 _27633_ (.A(net953),
    .B(_08260_),
    .Y(\cpu.qspi.c_wstrobe_d ));
 sg13g2_nor2_1 _27634_ (.A(_00179_),
    .B(_08260_),
    .Y(\cpu.qspi.c_wstrobe_i ));
 sg13g2_mux4_1 _27635_ (.S0(_04927_),
    .A0(_09180_),
    .A1(_09182_),
    .A2(_09190_),
    .A3(_09198_),
    .S1(\cpu.gpio.r_uart_rx_src[1] ),
    .X(_08261_));
 sg13g2_mux4_1 _27636_ (.S0(_04927_),
    .A0(_09177_),
    .A1(_09193_),
    .A2(_09175_),
    .A3(_09186_),
    .S1(\cpu.gpio.r_uart_rx_src[1] ),
    .X(_08262_));
 sg13g2_mux2_1 _27637_ (.A0(_08261_),
    .A1(_08262_),
    .S(\cpu.gpio.r_uart_rx_src[2] ),
    .X(\cpu.gpio.uart_rx ));
 sg13g2_mux4_1 _27638_ (.S0(_04915_),
    .A0(_11997_),
    .A1(net1114),
    .A2(_08145_),
    .A3(net1092),
    .S1(_05354_),
    .X(_08263_));
 sg13g2_mux4_1 _27639_ (.S0(_04915_),
    .A0(\cpu.gpio.genblk2[4].srcs_io[0] ),
    .A1(_07477_),
    .A2(net1111),
    .A3(net1112),
    .S1(_05354_),
    .X(_08264_));
 sg13g2_nor2b_1 _27640_ (.A(_05421_),
    .B_N(_08264_),
    .Y(_08265_));
 sg13g2_a21oi_1 _27641_ (.A1(_05421_),
    .A2(_08263_),
    .Y(_08266_),
    .B1(_08265_));
 sg13g2_nand2b_1 _27642_ (.Y(_08267_),
    .B(net1091),
    .A_N(_04915_));
 sg13g2_nand3_1 _27643_ (.B(_05354_),
    .C(net1094),
    .A(_04915_),
    .Y(_08268_));
 sg13g2_o21ai_1 _27644_ (.B1(_08268_),
    .Y(_08269_),
    .A1(_05354_),
    .A2(_08267_));
 sg13g2_nand3_1 _27645_ (.B(_00177_),
    .C(_08269_),
    .A(_05493_),
    .Y(_08270_));
 sg13g2_o21ai_1 _27646_ (.B1(_08270_),
    .Y(net15),
    .A1(_05493_),
    .A2(_08266_));
 sg13g2_mux4_1 _27647_ (.S0(_05554_),
    .A0(net1113),
    .A1(net1114),
    .A2(_08145_),
    .A3(_08147_),
    .S1(_05615_),
    .X(_08271_));
 sg13g2_mux4_1 _27648_ (.S0(_05554_),
    .A0(\cpu.gpio.genblk2[5].srcs_io[0] ),
    .A1(net1095),
    .A2(_12018_),
    .A3(_11999_),
    .S1(_05615_),
    .X(_08272_));
 sg13g2_nor2b_1 _27649_ (.A(_05683_),
    .B_N(_08272_),
    .Y(_08273_));
 sg13g2_a21oi_1 _27650_ (.A1(_05683_),
    .A2(_08271_),
    .Y(_08274_),
    .B1(_08273_));
 sg13g2_nand2b_1 _27651_ (.Y(_08275_),
    .B(_08149_),
    .A_N(_05554_));
 sg13g2_nand3_1 _27652_ (.B(_05615_),
    .C(net1094),
    .A(_05554_),
    .Y(_08276_));
 sg13g2_o21ai_1 _27653_ (.B1(_08276_),
    .Y(_08277_),
    .A1(_05615_),
    .A2(_08275_));
 sg13g2_nand3_1 _27654_ (.B(_00176_),
    .C(_08277_),
    .A(_05094_),
    .Y(_08278_));
 sg13g2_o21ai_1 _27655_ (.B1(_08278_),
    .Y(net16),
    .A1(_05094_),
    .A2(_08274_));
 sg13g2_mux4_1 _27656_ (.S0(_04916_),
    .A0(net1113),
    .A1(net1114),
    .A2(net1093),
    .A3(net1092),
    .S1(_06440_),
    .X(_08279_));
 sg13g2_mux4_1 _27657_ (.S0(_04916_),
    .A0(\cpu.gpio.genblk2[6].srcs_io[0] ),
    .A1(net1095),
    .A2(net1111),
    .A3(net1112),
    .S1(_06440_),
    .X(_08280_));
 sg13g2_nor2b_1 _27658_ (.A(\cpu.gpio.r_src_io[6][2] ),
    .B_N(_08280_),
    .Y(_08281_));
 sg13g2_a21oi_1 _27659_ (.A1(\cpu.gpio.r_src_io[6][2] ),
    .A2(_08279_),
    .Y(_08282_),
    .B1(_08281_));
 sg13g2_nand2b_1 _27660_ (.Y(_08283_),
    .B(net1091),
    .A_N(_04916_));
 sg13g2_nand3_1 _27661_ (.B(net1094),
    .C(_06440_),
    .A(_04916_),
    .Y(_08284_));
 sg13g2_o21ai_1 _27662_ (.B1(_08284_),
    .Y(_08285_),
    .A1(_06440_),
    .A2(_08283_));
 sg13g2_nand3_1 _27663_ (.B(\cpu.gpio.r_src_io[6][3] ),
    .C(_08285_),
    .A(_00102_),
    .Y(_08286_));
 sg13g2_o21ai_1 _27664_ (.B1(_08286_),
    .Y(net17),
    .A1(\cpu.gpio.r_src_io[6][3] ),
    .A2(_08282_));
 sg13g2_mux4_1 _27665_ (.S0(_05555_),
    .A0(_11997_),
    .A1(_11990_),
    .A2(net1093),
    .A3(net1092),
    .S1(_06441_),
    .X(_08287_));
 sg13g2_mux4_1 _27666_ (.S0(_05555_),
    .A0(\cpu.gpio.genblk2[7].srcs_io[0] ),
    .A1(net1095),
    .A2(net1111),
    .A3(net1112),
    .S1(_06441_),
    .X(_08288_));
 sg13g2_nor2b_1 _27667_ (.A(\cpu.gpio.r_src_io[7][2] ),
    .B_N(_08288_),
    .Y(_08289_));
 sg13g2_a21oi_1 _27668_ (.A1(\cpu.gpio.r_src_io[7][2] ),
    .A2(_08287_),
    .Y(_08290_),
    .B1(_08289_));
 sg13g2_nand2b_1 _27669_ (.Y(_08291_),
    .B(net1091),
    .A_N(_05555_));
 sg13g2_nand3_1 _27670_ (.B(net1094),
    .C(_06441_),
    .A(_05555_),
    .Y(_08292_));
 sg13g2_o21ai_1 _27671_ (.B1(_08292_),
    .Y(_08293_),
    .A1(_06441_),
    .A2(_08291_));
 sg13g2_nand3_1 _27672_ (.B(\cpu.gpio.r_src_io[7][3] ),
    .C(_08293_),
    .A(_00139_),
    .Y(_08294_));
 sg13g2_o21ai_1 _27673_ (.B1(_08294_),
    .Y(net18),
    .A1(\cpu.gpio.r_src_io[7][3] ),
    .A2(_08290_));
 sg13g2_xor2_1 _27674_ (.B(clknet_leaf_79_clk),
    .A(\cpu.r_clk_invert ),
    .X(net21));
 sg13g2_mux4_1 _27675_ (.S0(_05560_),
    .A0(net1113),
    .A1(net1114),
    .A2(net1093),
    .A3(net1092),
    .S1(_06445_),
    .X(_08295_));
 sg13g2_mux4_1 _27676_ (.S0(_05560_),
    .A0(\cpu.gpio.genblk1[3].srcs_o[0] ),
    .A1(net1095),
    .A2(net1111),
    .A3(net1112),
    .S1(_06445_),
    .X(_08296_));
 sg13g2_nor2b_1 _27677_ (.A(\cpu.gpio.r_src_o[3][2] ),
    .B_N(_08296_),
    .Y(_08297_));
 sg13g2_a21oi_1 _27678_ (.A1(\cpu.gpio.r_src_o[3][2] ),
    .A2(_08295_),
    .Y(_08298_),
    .B1(_08297_));
 sg13g2_nand2_1 _27679_ (.Y(_08299_),
    .A(net1091),
    .B(_05561_));
 sg13g2_nand3_1 _27680_ (.B(net1094),
    .C(_06445_),
    .A(_05560_),
    .Y(_08300_));
 sg13g2_o21ai_1 _27681_ (.B1(_08300_),
    .Y(_08301_),
    .A1(_06445_),
    .A2(_08299_));
 sg13g2_nand3_1 _27682_ (.B(\cpu.gpio.r_src_o[3][3] ),
    .C(_08301_),
    .A(_00142_),
    .Y(_08302_));
 sg13g2_o21ai_1 _27683_ (.B1(_08302_),
    .Y(net22),
    .A1(\cpu.gpio.r_src_o[3][3] ),
    .A2(_08298_));
 sg13g2_mux4_1 _27684_ (.S0(_04901_),
    .A0(net1113),
    .A1(_11990_),
    .A2(net1093),
    .A3(net1092),
    .S1(_06448_),
    .X(_08303_));
 sg13g2_mux4_1 _27685_ (.S0(_04901_),
    .A0(\cpu.gpio.genblk1[4].srcs_o[0] ),
    .A1(net1095),
    .A2(net1111),
    .A3(net1112),
    .S1(_06448_),
    .X(_08304_));
 sg13g2_nor2b_1 _27686_ (.A(\cpu.gpio.r_src_o[4][2] ),
    .B_N(_08304_),
    .Y(_08305_));
 sg13g2_a21oi_1 _27687_ (.A1(\cpu.gpio.r_src_o[4][2] ),
    .A2(_08303_),
    .Y(_08306_),
    .B1(_08305_));
 sg13g2_nand2b_1 _27688_ (.Y(_08307_),
    .B(_08149_),
    .A_N(_04901_));
 sg13g2_nand3_1 _27689_ (.B(net1094),
    .C(_06448_),
    .A(_04901_),
    .Y(_08308_));
 sg13g2_o21ai_1 _27690_ (.B1(_08308_),
    .Y(_08309_),
    .A1(_06448_),
    .A2(_08307_));
 sg13g2_nand3_1 _27691_ (.B(\cpu.gpio.r_src_o[4][3] ),
    .C(_08309_),
    .A(_00104_),
    .Y(_08310_));
 sg13g2_o21ai_1 _27692_ (.B1(_08310_),
    .Y(net23),
    .A1(\cpu.gpio.r_src_o[4][3] ),
    .A2(_08306_));
 sg13g2_mux4_1 _27693_ (.S0(_05564_),
    .A0(net1113),
    .A1(net1114),
    .A2(net1093),
    .A3(_08147_),
    .S1(_06450_),
    .X(_08311_));
 sg13g2_mux4_1 _27694_ (.S0(_05564_),
    .A0(\cpu.gpio.genblk1[5].srcs_o[0] ),
    .A1(net1095),
    .A2(net1111),
    .A3(net1112),
    .S1(_06450_),
    .X(_08312_));
 sg13g2_nor2b_1 _27695_ (.A(\cpu.gpio.r_src_o[5][2] ),
    .B_N(_08312_),
    .Y(_08313_));
 sg13g2_a21oi_1 _27696_ (.A1(\cpu.gpio.r_src_o[5][2] ),
    .A2(_08311_),
    .Y(_08314_),
    .B1(_08313_));
 sg13g2_nand2b_1 _27697_ (.Y(_08315_),
    .B(net1091),
    .A_N(_05564_));
 sg13g2_nand3_1 _27698_ (.B(net1094),
    .C(_06450_),
    .A(_05564_),
    .Y(_08316_));
 sg13g2_o21ai_1 _27699_ (.B1(_08316_),
    .Y(_08317_),
    .A1(_06450_),
    .A2(_08315_));
 sg13g2_nand3_1 _27700_ (.B(\cpu.gpio.r_src_o[5][3] ),
    .C(_08317_),
    .A(_00141_),
    .Y(_08318_));
 sg13g2_o21ai_1 _27701_ (.B1(_08318_),
    .Y(net24),
    .A1(\cpu.gpio.r_src_o[5][3] ),
    .A2(_08314_));
 sg13g2_mux4_1 _27702_ (.S0(_04910_),
    .A0(net1113),
    .A1(net1114),
    .A2(net1093),
    .A3(net1092),
    .S1(_07999_),
    .X(_08319_));
 sg13g2_mux4_1 _27703_ (.S0(_04910_),
    .A0(\cpu.gpio.genblk1[6].srcs_o[0] ),
    .A1(net1095),
    .A2(_12018_),
    .A3(_11999_),
    .S1(_07999_),
    .X(_08320_));
 sg13g2_nor2b_1 _27704_ (.A(\cpu.gpio.r_src_o[6][2] ),
    .B_N(_08320_),
    .Y(_08321_));
 sg13g2_a21oi_1 _27705_ (.A1(\cpu.gpio.r_src_o[6][2] ),
    .A2(_08319_),
    .Y(_08322_),
    .B1(_08321_));
 sg13g2_nand2b_1 _27706_ (.Y(_08323_),
    .B(net1091),
    .A_N(_04910_));
 sg13g2_nand3_1 _27707_ (.B(net1094),
    .C(_07999_),
    .A(_04910_),
    .Y(_08324_));
 sg13g2_o21ai_1 _27708_ (.B1(_08324_),
    .Y(_08325_),
    .A1(_07999_),
    .A2(_08323_));
 sg13g2_nand3_1 _27709_ (.B(\cpu.gpio.r_src_o[6][3] ),
    .C(_08325_),
    .A(_00103_),
    .Y(_08326_));
 sg13g2_o21ai_1 _27710_ (.B1(_08326_),
    .Y(net25),
    .A1(\cpu.gpio.r_src_o[6][3] ),
    .A2(_08322_));
 sg13g2_mux4_1 _27711_ (.S0(_05559_),
    .A0(net1113),
    .A1(net1114),
    .A2(net1093),
    .A3(net1092),
    .S1(_06456_),
    .X(_08327_));
 sg13g2_mux4_1 _27712_ (.S0(_05559_),
    .A0(\cpu.gpio.genblk1[7].srcs_o[0] ),
    .A1(net1095),
    .A2(net1111),
    .A3(net1112),
    .S1(_06456_),
    .X(_08328_));
 sg13g2_nor2b_1 _27713_ (.A(\cpu.gpio.r_src_o[7][2] ),
    .B_N(_08328_),
    .Y(_08329_));
 sg13g2_a21oi_1 _27714_ (.A1(\cpu.gpio.r_src_o[7][2] ),
    .A2(_08327_),
    .Y(_08330_),
    .B1(_08329_));
 sg13g2_nand2b_1 _27715_ (.Y(_08331_),
    .B(net1091),
    .A_N(_05559_));
 sg13g2_nand3_1 _27716_ (.B(_08090_),
    .C(_06456_),
    .A(_05559_),
    .Y(_08332_));
 sg13g2_o21ai_1 _27717_ (.B1(_08332_),
    .Y(_08333_),
    .A1(_06456_),
    .A2(_08331_));
 sg13g2_nand3_1 _27718_ (.B(\cpu.gpio.r_src_o[7][3] ),
    .C(_08333_),
    .A(_00140_),
    .Y(_08334_));
 sg13g2_o21ai_1 _27719_ (.B1(_08334_),
    .Y(net26),
    .A1(\cpu.gpio.r_src_o[7][3] ),
    .A2(_08330_));
 sg13g2_dfrbp_1 _27720_ (.CLK(clknet_leaf_16_clk),
    .RESET_B(net1150),
    .D(_00305_),
    .Q_N(_14973_),
    .Q(\cpu.intr.r_swi ));
 sg13g2_dfrbp_1 _27721_ (.CLK(clknet_leaf_59_clk),
    .RESET_B(net1151),
    .D(_00306_),
    .Q_N(_14972_),
    .Q(\cpu.gpio.genblk1[3].srcs_o[5] ));
 sg13g2_dfrbp_1 _27722_ (.CLK(clknet_leaf_59_clk),
    .RESET_B(net1152),
    .D(_00307_),
    .Q_N(_14971_),
    .Q(\cpu.gpio.genblk1[3].srcs_o[4] ));
 sg13g2_dfrbp_1 _27723_ (.CLK(clknet_leaf_64_clk),
    .RESET_B(net1153),
    .D(_00308_),
    .Q_N(_14970_),
    .Q(\cpu.gpio.genblk1[3].srcs_o[3] ));
 sg13g2_dfrbp_1 _27724_ (.CLK(clknet_leaf_64_clk),
    .RESET_B(net1154),
    .D(_00309_),
    .Q_N(_14969_),
    .Q(\cpu.gpio.genblk1[3].srcs_o[2] ));
 sg13g2_buf_8 clkbuf_leaf_0_clk (.A(clknet_6_0__leaf_clk),
    .X(clknet_leaf_0_clk));
 sg13g2_buf_1 _27726_ (.A(net6),
    .X(net4));
 sg13g2_buf_1 _27727_ (.A(net6),
    .X(net5));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[0][0]$_DFFE_PP_  (.CLK(clknet_leaf_66_clk),
    .RESET_B(net1155),
    .D(_00310_),
    .Q_N(_14968_),
    .Q(\cpu.dcache.r_data[0][0] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[0][10]$_DFFE_PP_  (.CLK(clknet_leaf_46_clk),
    .RESET_B(net1156),
    .D(_00311_),
    .Q_N(_00099_),
    .Q(\cpu.dcache.r_data[0][10] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[0][11]$_DFFE_PP_  (.CLK(clknet_leaf_46_clk),
    .RESET_B(net1157),
    .D(_00312_),
    .Q_N(_00109_),
    .Q(\cpu.dcache.r_data[0][11] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[0][12]$_DFFE_PP_  (.CLK(clknet_leaf_34_clk),
    .RESET_B(net1158),
    .D(_00313_),
    .Q_N(_00119_),
    .Q(\cpu.dcache.r_data[0][12] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[0][13]$_DFFE_PP_  (.CLK(clknet_leaf_34_clk),
    .RESET_B(net1159),
    .D(_00314_),
    .Q_N(_00125_),
    .Q(\cpu.dcache.r_data[0][13] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[0][14]$_DFFE_PP_  (.CLK(clknet_leaf_35_clk),
    .RESET_B(net1160),
    .D(_00315_),
    .Q_N(_00136_),
    .Q(\cpu.dcache.r_data[0][14] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[0][15]$_DFFE_PP_  (.CLK(clknet_leaf_34_clk),
    .RESET_B(net1161),
    .D(_00316_),
    .Q_N(_00147_),
    .Q(\cpu.dcache.r_data[0][15] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[0][16]$_DFFE_PP_  (.CLK(clknet_leaf_66_clk),
    .RESET_B(net1162),
    .D(_00317_),
    .Q_N(_14967_),
    .Q(\cpu.dcache.r_data[0][16] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[0][17]$_DFFE_PP_  (.CLK(clknet_leaf_52_clk),
    .RESET_B(net1163),
    .D(_00318_),
    .Q_N(_00299_),
    .Q(\cpu.dcache.r_data[0][17] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[0][18]$_DFFE_PP_  (.CLK(clknet_leaf_52_clk),
    .RESET_B(net1164),
    .D(_00319_),
    .Q_N(_00097_),
    .Q(\cpu.dcache.r_data[0][18] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[0][19]$_DFFE_PP_  (.CLK(clknet_leaf_52_clk),
    .RESET_B(net1165),
    .D(_00320_),
    .Q_N(_00107_),
    .Q(\cpu.dcache.r_data[0][19] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[0][1]$_DFFE_PP_  (.CLK(clknet_leaf_52_clk),
    .RESET_B(net1166),
    .D(_00321_),
    .Q_N(_14966_),
    .Q(\cpu.dcache.r_data[0][1] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[0][20]$_DFFE_PP_  (.CLK(clknet_leaf_54_clk),
    .RESET_B(net1167),
    .D(_00322_),
    .Q_N(_00117_),
    .Q(\cpu.dcache.r_data[0][20] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[0][21]$_DFFE_PP_  (.CLK(clknet_leaf_54_clk),
    .RESET_B(net1168),
    .D(_00323_),
    .Q_N(_00123_),
    .Q(\cpu.dcache.r_data[0][21] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[0][22]$_DFFE_PP_  (.CLK(clknet_leaf_54_clk),
    .RESET_B(net1169),
    .D(_00324_),
    .Q_N(_00134_),
    .Q(\cpu.dcache.r_data[0][22] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[0][23]$_DFFE_PP_  (.CLK(clknet_leaf_53_clk),
    .RESET_B(net1170),
    .D(_00325_),
    .Q_N(_00145_),
    .Q(\cpu.dcache.r_data[0][23] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[0][24]$_DFFE_PP_  (.CLK(clknet_leaf_47_clk),
    .RESET_B(net1171),
    .D(_00326_),
    .Q_N(_00295_),
    .Q(\cpu.dcache.r_data[0][24] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[0][25]$_DFFE_PP_  (.CLK(clknet_leaf_46_clk),
    .RESET_B(net1172),
    .D(_00327_),
    .Q_N(_00300_),
    .Q(\cpu.dcache.r_data[0][25] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[0][26]$_DFFE_PP_  (.CLK(clknet_leaf_47_clk),
    .RESET_B(net1173),
    .D(_00328_),
    .Q_N(_00098_),
    .Q(\cpu.dcache.r_data[0][26] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[0][27]$_DFFE_PP_  (.CLK(clknet_leaf_47_clk),
    .RESET_B(net1174),
    .D(_00329_),
    .Q_N(_00108_),
    .Q(\cpu.dcache.r_data[0][27] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[0][28]$_DFFE_PP_  (.CLK(clknet_leaf_23_clk),
    .RESET_B(net1175),
    .D(_00330_),
    .Q_N(_00118_),
    .Q(\cpu.dcache.r_data[0][28] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[0][29]$_DFFE_PP_  (.CLK(clknet_leaf_23_clk),
    .RESET_B(net1176),
    .D(_00331_),
    .Q_N(_00124_),
    .Q(\cpu.dcache.r_data[0][29] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[0][2]$_DFFE_PP_  (.CLK(clknet_leaf_52_clk),
    .RESET_B(net1177),
    .D(_00332_),
    .Q_N(_14965_),
    .Q(\cpu.dcache.r_data[0][2] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[0][30]$_DFFE_PP_  (.CLK(clknet_leaf_46_clk),
    .RESET_B(net1178),
    .D(_00333_),
    .Q_N(_00135_),
    .Q(\cpu.dcache.r_data[0][30] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[0][31]$_DFFE_PP_  (.CLK(clknet_leaf_33_clk),
    .RESET_B(net1179),
    .D(_00334_),
    .Q_N(_00146_),
    .Q(\cpu.dcache.r_data[0][31] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[0][3]$_DFFE_PP_  (.CLK(clknet_leaf_66_clk),
    .RESET_B(net1180),
    .D(_00335_),
    .Q_N(_14964_),
    .Q(\cpu.dcache.r_data[0][3] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[0][4]$_DFFE_PP_  (.CLK(clknet_leaf_53_clk),
    .RESET_B(net1181),
    .D(_00336_),
    .Q_N(_00116_),
    .Q(\cpu.dcache.r_data[0][4] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[0][5]$_DFFE_PP_  (.CLK(clknet_leaf_53_clk),
    .RESET_B(net1182),
    .D(_00337_),
    .Q_N(_00122_),
    .Q(\cpu.dcache.r_data[0][5] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[0][6]$_DFFE_PP_  (.CLK(clknet_leaf_53_clk),
    .RESET_B(net1183),
    .D(_00338_),
    .Q_N(_00133_),
    .Q(\cpu.dcache.r_data[0][6] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[0][7]$_DFFE_PP_  (.CLK(clknet_leaf_53_clk),
    .RESET_B(net1184),
    .D(_00339_),
    .Q_N(_00144_),
    .Q(\cpu.dcache.r_data[0][7] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[0][8]$_DFFE_PP_  (.CLK(clknet_leaf_46_clk),
    .RESET_B(net1185),
    .D(_00340_),
    .Q_N(_00296_),
    .Q(\cpu.dcache.r_data[0][8] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[0][9]$_DFFE_PP_  (.CLK(clknet_leaf_46_clk),
    .RESET_B(net1186),
    .D(_00341_),
    .Q_N(_00301_),
    .Q(\cpu.dcache.r_data[0][9] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[1][0]$_DFFE_PP_  (.CLK(clknet_leaf_24_clk),
    .RESET_B(net1187),
    .D(_00342_),
    .Q_N(_14963_),
    .Q(\cpu.dcache.r_data[1][0] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[1][10]$_DFFE_PP_  (.CLK(clknet_leaf_29_clk),
    .RESET_B(net1188),
    .D(_00343_),
    .Q_N(_14962_),
    .Q(\cpu.dcache.r_data[1][10] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[1][11]$_DFFE_PP_  (.CLK(clknet_leaf_27_clk),
    .RESET_B(net1189),
    .D(_00344_),
    .Q_N(_14961_),
    .Q(\cpu.dcache.r_data[1][11] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[1][12]$_DFFE_PP_  (.CLK(clknet_leaf_32_clk),
    .RESET_B(net1190),
    .D(_00345_),
    .Q_N(_14960_),
    .Q(\cpu.dcache.r_data[1][12] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[1][13]$_DFFE_PP_  (.CLK(clknet_leaf_29_clk),
    .RESET_B(net1191),
    .D(_00346_),
    .Q_N(_14959_),
    .Q(\cpu.dcache.r_data[1][13] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[1][14]$_DFFE_PP_  (.CLK(clknet_leaf_29_clk),
    .RESET_B(net1192),
    .D(_00347_),
    .Q_N(_14958_),
    .Q(\cpu.dcache.r_data[1][14] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[1][15]$_DFFE_PP_  (.CLK(clknet_leaf_29_clk),
    .RESET_B(net1193),
    .D(_00348_),
    .Q_N(_14957_),
    .Q(\cpu.dcache.r_data[1][15] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[1][16]$_DFFE_PP_  (.CLK(clknet_leaf_23_clk),
    .RESET_B(net1194),
    .D(_00349_),
    .Q_N(_14956_),
    .Q(\cpu.dcache.r_data[1][16] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[1][17]$_DFFE_PP_  (.CLK(clknet_leaf_23_clk),
    .RESET_B(net1195),
    .D(_00350_),
    .Q_N(_14955_),
    .Q(\cpu.dcache.r_data[1][17] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[1][18]$_DFFE_PP_  (.CLK(clknet_leaf_54_clk),
    .RESET_B(net1196),
    .D(_00351_),
    .Q_N(_14954_),
    .Q(\cpu.dcache.r_data[1][18] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[1][19]$_DFFE_PP_  (.CLK(clknet_leaf_54_clk),
    .RESET_B(net1197),
    .D(_00352_),
    .Q_N(_14953_),
    .Q(\cpu.dcache.r_data[1][19] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[1][1]$_DFFE_PP_  (.CLK(clknet_leaf_25_clk),
    .RESET_B(net1198),
    .D(_00353_),
    .Q_N(_14952_),
    .Q(\cpu.dcache.r_data[1][1] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[1][20]$_DFFE_PP_  (.CLK(clknet_leaf_54_clk),
    .RESET_B(net1199),
    .D(_00354_),
    .Q_N(_14951_),
    .Q(\cpu.dcache.r_data[1][20] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[1][21]$_DFFE_PP_  (.CLK(clknet_leaf_22_clk),
    .RESET_B(net1200),
    .D(_00355_),
    .Q_N(_14950_),
    .Q(\cpu.dcache.r_data[1][21] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[1][22]$_DFFE_PP_  (.CLK(clknet_leaf_23_clk),
    .RESET_B(net1201),
    .D(_00356_),
    .Q_N(_14949_),
    .Q(\cpu.dcache.r_data[1][22] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[1][23]$_DFFE_PP_  (.CLK(clknet_leaf_54_clk),
    .RESET_B(net1202),
    .D(_00357_),
    .Q_N(_14948_),
    .Q(\cpu.dcache.r_data[1][23] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[1][24]$_DFFE_PP_  (.CLK(clknet_leaf_24_clk),
    .RESET_B(net1203),
    .D(_00358_),
    .Q_N(_14947_),
    .Q(\cpu.dcache.r_data[1][24] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[1][25]$_DFFE_PP_  (.CLK(clknet_leaf_24_clk),
    .RESET_B(net1204),
    .D(_00359_),
    .Q_N(_14946_),
    .Q(\cpu.dcache.r_data[1][25] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[1][26]$_DFFE_PP_  (.CLK(clknet_leaf_33_clk),
    .RESET_B(net1205),
    .D(_00360_),
    .Q_N(_14945_),
    .Q(\cpu.dcache.r_data[1][26] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[1][27]$_DFFE_PP_  (.CLK(clknet_leaf_33_clk),
    .RESET_B(net1206),
    .D(_00361_),
    .Q_N(_14944_),
    .Q(\cpu.dcache.r_data[1][27] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[1][28]$_DFFE_PP_  (.CLK(clknet_leaf_24_clk),
    .RESET_B(net1207),
    .D(_00362_),
    .Q_N(_14943_),
    .Q(\cpu.dcache.r_data[1][28] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[1][29]$_DFFE_PP_  (.CLK(clknet_leaf_33_clk),
    .RESET_B(net1208),
    .D(_00363_),
    .Q_N(_14942_),
    .Q(\cpu.dcache.r_data[1][29] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[1][2]$_DFFE_PP_  (.CLK(clknet_leaf_25_clk),
    .RESET_B(net1209),
    .D(_00364_),
    .Q_N(_14941_),
    .Q(\cpu.dcache.r_data[1][2] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[1][30]$_DFFE_PP_  (.CLK(clknet_leaf_32_clk),
    .RESET_B(net1210),
    .D(_00365_),
    .Q_N(_14940_),
    .Q(\cpu.dcache.r_data[1][30] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[1][31]$_DFFE_PP_  (.CLK(clknet_leaf_24_clk),
    .RESET_B(net1211),
    .D(_00366_),
    .Q_N(_14939_),
    .Q(\cpu.dcache.r_data[1][31] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[1][3]$_DFFE_PP_  (.CLK(clknet_leaf_25_clk),
    .RESET_B(net1212),
    .D(_00367_),
    .Q_N(_14938_),
    .Q(\cpu.dcache.r_data[1][3] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[1][4]$_DFFE_PP_  (.CLK(clknet_leaf_25_clk),
    .RESET_B(net1213),
    .D(_00368_),
    .Q_N(_14937_),
    .Q(\cpu.dcache.r_data[1][4] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[1][5]$_DFFE_PP_  (.CLK(clknet_leaf_21_clk),
    .RESET_B(net1214),
    .D(_00369_),
    .Q_N(_14936_),
    .Q(\cpu.dcache.r_data[1][5] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[1][6]$_DFFE_PP_  (.CLK(clknet_leaf_23_clk),
    .RESET_B(net1215),
    .D(_00370_),
    .Q_N(_14935_),
    .Q(\cpu.dcache.r_data[1][6] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[1][7]$_DFFE_PP_  (.CLK(clknet_leaf_25_clk),
    .RESET_B(net1216),
    .D(_00371_),
    .Q_N(_14934_),
    .Q(\cpu.dcache.r_data[1][7] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[1][8]$_DFFE_PP_  (.CLK(clknet_leaf_32_clk),
    .RESET_B(net1217),
    .D(_00372_),
    .Q_N(_14933_),
    .Q(\cpu.dcache.r_data[1][8] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[1][9]$_DFFE_PP_  (.CLK(clknet_leaf_27_clk),
    .RESET_B(net1218),
    .D(_00373_),
    .Q_N(_14932_),
    .Q(\cpu.dcache.r_data[1][9] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[2][0]$_DFFE_PP_  (.CLK(clknet_leaf_27_clk),
    .RESET_B(net1219),
    .D(_00374_),
    .Q_N(_14931_),
    .Q(\cpu.dcache.r_data[2][0] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[2][10]$_DFFE_PP_  (.CLK(clknet_leaf_30_clk),
    .RESET_B(net1220),
    .D(_00375_),
    .Q_N(_14930_),
    .Q(\cpu.dcache.r_data[2][10] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[2][11]$_DFFE_PP_  (.CLK(clknet_leaf_29_clk),
    .RESET_B(net1221),
    .D(_00376_),
    .Q_N(_14929_),
    .Q(\cpu.dcache.r_data[2][11] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[2][12]$_DFFE_PP_  (.CLK(clknet_leaf_29_clk),
    .RESET_B(net1222),
    .D(_00377_),
    .Q_N(_14928_),
    .Q(\cpu.dcache.r_data[2][12] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[2][13]$_DFFE_PP_  (.CLK(clknet_leaf_30_clk),
    .RESET_B(net1223),
    .D(_00378_),
    .Q_N(_14927_),
    .Q(\cpu.dcache.r_data[2][13] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[2][14]$_DFFE_PP_  (.CLK(clknet_leaf_30_clk),
    .RESET_B(net1224),
    .D(_00379_),
    .Q_N(_14926_),
    .Q(\cpu.dcache.r_data[2][14] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[2][15]$_DFFE_PP_  (.CLK(clknet_leaf_29_clk),
    .RESET_B(net1225),
    .D(_00380_),
    .Q_N(_14925_),
    .Q(\cpu.dcache.r_data[2][15] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[2][16]$_DFFE_PP_  (.CLK(clknet_leaf_24_clk),
    .RESET_B(net1226),
    .D(_00381_),
    .Q_N(_14924_),
    .Q(\cpu.dcache.r_data[2][16] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[2][17]$_DFFE_PP_  (.CLK(clknet_leaf_24_clk),
    .RESET_B(net1227),
    .D(_00382_),
    .Q_N(_14923_),
    .Q(\cpu.dcache.r_data[2][17] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[2][18]$_DFFE_PP_  (.CLK(clknet_leaf_23_clk),
    .RESET_B(net1228),
    .D(_00383_),
    .Q_N(_14922_),
    .Q(\cpu.dcache.r_data[2][18] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[2][19]$_DFFE_PP_  (.CLK(clknet_leaf_24_clk),
    .RESET_B(net1229),
    .D(_00384_),
    .Q_N(_14921_),
    .Q(\cpu.dcache.r_data[2][19] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[2][1]$_DFFE_PP_  (.CLK(clknet_leaf_27_clk),
    .RESET_B(net1230),
    .D(_00385_),
    .Q_N(_14920_),
    .Q(\cpu.dcache.r_data[2][1] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[2][20]$_DFFE_PP_  (.CLK(clknet_leaf_22_clk),
    .RESET_B(net1231),
    .D(_00386_),
    .Q_N(_14919_),
    .Q(\cpu.dcache.r_data[2][20] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[2][21]$_DFFE_PP_  (.CLK(clknet_leaf_22_clk),
    .RESET_B(net1232),
    .D(_00387_),
    .Q_N(_14918_),
    .Q(\cpu.dcache.r_data[2][21] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[2][22]$_DFFE_PP_  (.CLK(clknet_leaf_23_clk),
    .RESET_B(net1233),
    .D(_00388_),
    .Q_N(_14917_),
    .Q(\cpu.dcache.r_data[2][22] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[2][23]$_DFFE_PP_  (.CLK(clknet_leaf_22_clk),
    .RESET_B(net1234),
    .D(_00389_),
    .Q_N(_14916_),
    .Q(\cpu.dcache.r_data[2][23] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[2][24]$_DFFE_PP_  (.CLK(clknet_leaf_34_clk),
    .RESET_B(net1235),
    .D(_00390_),
    .Q_N(_14915_),
    .Q(\cpu.dcache.r_data[2][24] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[2][25]$_DFFE_PP_  (.CLK(clknet_leaf_34_clk),
    .RESET_B(net1236),
    .D(_00391_),
    .Q_N(_14914_),
    .Q(\cpu.dcache.r_data[2][25] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[2][26]$_DFFE_PP_  (.CLK(clknet_leaf_34_clk),
    .RESET_B(net1237),
    .D(_00392_),
    .Q_N(_14913_),
    .Q(\cpu.dcache.r_data[2][26] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[2][27]$_DFFE_PP_  (.CLK(clknet_leaf_34_clk),
    .RESET_B(net1238),
    .D(_00393_),
    .Q_N(_14912_),
    .Q(\cpu.dcache.r_data[2][27] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[2][28]$_DFFE_PP_  (.CLK(clknet_leaf_32_clk),
    .RESET_B(net1239),
    .D(_00394_),
    .Q_N(_14911_),
    .Q(\cpu.dcache.r_data[2][28] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[2][29]$_DFFE_PP_  (.CLK(clknet_leaf_31_clk),
    .RESET_B(net1240),
    .D(_00395_),
    .Q_N(_14910_),
    .Q(\cpu.dcache.r_data[2][29] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[2][2]$_DFFE_PP_  (.CLK(clknet_leaf_27_clk),
    .RESET_B(net1241),
    .D(_00396_),
    .Q_N(_14909_),
    .Q(\cpu.dcache.r_data[2][2] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[2][30]$_DFFE_PP_  (.CLK(clknet_leaf_32_clk),
    .RESET_B(net1242),
    .D(_00397_),
    .Q_N(_14908_),
    .Q(\cpu.dcache.r_data[2][30] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[2][31]$_DFFE_PP_  (.CLK(clknet_leaf_32_clk),
    .RESET_B(net1243),
    .D(_00398_),
    .Q_N(_14907_),
    .Q(\cpu.dcache.r_data[2][31] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[2][3]$_DFFE_PP_  (.CLK(clknet_leaf_27_clk),
    .RESET_B(net1244),
    .D(_00399_),
    .Q_N(_14906_),
    .Q(\cpu.dcache.r_data[2][3] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[2][4]$_DFFE_PP_  (.CLK(clknet_leaf_11_clk),
    .RESET_B(net1245),
    .D(_00400_),
    .Q_N(_14905_),
    .Q(\cpu.dcache.r_data[2][4] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[2][5]$_DFFE_PP_  (.CLK(clknet_leaf_26_clk),
    .RESET_B(net1246),
    .D(_00401_),
    .Q_N(_14904_),
    .Q(\cpu.dcache.r_data[2][5] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[2][6]$_DFFE_PP_  (.CLK(clknet_leaf_26_clk),
    .RESET_B(net1247),
    .D(_00402_),
    .Q_N(_14903_),
    .Q(\cpu.dcache.r_data[2][6] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[2][7]$_DFFE_PP_  (.CLK(clknet_leaf_27_clk),
    .RESET_B(net1248),
    .D(_00403_),
    .Q_N(_14902_),
    .Q(\cpu.dcache.r_data[2][7] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[2][8]$_DFFE_PP_  (.CLK(clknet_leaf_32_clk),
    .RESET_B(net1249),
    .D(_00404_),
    .Q_N(_14901_),
    .Q(\cpu.dcache.r_data[2][8] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[2][9]$_DFFE_PP_  (.CLK(clknet_leaf_30_clk),
    .RESET_B(net1250),
    .D(_00405_),
    .Q_N(_14900_),
    .Q(\cpu.dcache.r_data[2][9] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[3][0]$_DFFE_PP_  (.CLK(clknet_leaf_28_clk),
    .RESET_B(net1251),
    .D(_00406_),
    .Q_N(_14899_),
    .Q(\cpu.dcache.r_data[3][0] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[3][10]$_DFFE_PP_  (.CLK(clknet_leaf_274_clk),
    .RESET_B(net1252),
    .D(_00407_),
    .Q_N(_14898_),
    .Q(\cpu.dcache.r_data[3][10] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[3][11]$_DFFE_PP_  (.CLK(clknet_leaf_274_clk),
    .RESET_B(net1253),
    .D(_00408_),
    .Q_N(_14897_),
    .Q(\cpu.dcache.r_data[3][11] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[3][12]$_DFFE_PP_  (.CLK(clknet_leaf_274_clk),
    .RESET_B(net1254),
    .D(_00409_),
    .Q_N(_14896_),
    .Q(\cpu.dcache.r_data[3][12] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[3][13]$_DFFE_PP_  (.CLK(clknet_leaf_274_clk),
    .RESET_B(net1255),
    .D(_00410_),
    .Q_N(_14895_),
    .Q(\cpu.dcache.r_data[3][13] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[3][14]$_DFFE_PP_  (.CLK(clknet_leaf_274_clk),
    .RESET_B(net1256),
    .D(_00411_),
    .Q_N(_14894_),
    .Q(\cpu.dcache.r_data[3][14] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[3][15]$_DFFE_PP_  (.CLK(clknet_leaf_274_clk),
    .RESET_B(net1257),
    .D(_00412_),
    .Q_N(_14893_),
    .Q(\cpu.dcache.r_data[3][15] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[3][16]$_DFFE_PP_  (.CLK(clknet_leaf_10_clk),
    .RESET_B(net1258),
    .D(_00413_),
    .Q_N(_14892_),
    .Q(\cpu.dcache.r_data[3][16] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[3][17]$_DFFE_PP_  (.CLK(clknet_leaf_26_clk),
    .RESET_B(net1259),
    .D(_00414_),
    .Q_N(_14891_),
    .Q(\cpu.dcache.r_data[3][17] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[3][18]$_DFFE_PP_  (.CLK(clknet_leaf_9_clk),
    .RESET_B(net1260),
    .D(_00415_),
    .Q_N(_14890_),
    .Q(\cpu.dcache.r_data[3][18] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[3][19]$_DFFE_PP_  (.CLK(clknet_leaf_26_clk),
    .RESET_B(net1261),
    .D(_00416_),
    .Q_N(_14889_),
    .Q(\cpu.dcache.r_data[3][19] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[3][1]$_DFFE_PP_  (.CLK(clknet_leaf_9_clk),
    .RESET_B(net1262),
    .D(_00417_),
    .Q_N(_14888_),
    .Q(\cpu.dcache.r_data[3][1] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[3][20]$_DFFE_PP_  (.CLK(clknet_leaf_55_clk),
    .RESET_B(net1263),
    .D(_00418_),
    .Q_N(_14887_),
    .Q(\cpu.dcache.r_data[3][20] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[3][21]$_DFFE_PP_  (.CLK(clknet_leaf_25_clk),
    .RESET_B(net1264),
    .D(_00419_),
    .Q_N(_14886_),
    .Q(\cpu.dcache.r_data[3][21] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[3][22]$_DFFE_PP_  (.CLK(clknet_leaf_11_clk),
    .RESET_B(net1265),
    .D(_00420_),
    .Q_N(_14885_),
    .Q(\cpu.dcache.r_data[3][22] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[3][23]$_DFFE_PP_  (.CLK(clknet_leaf_54_clk),
    .RESET_B(net1266),
    .D(_00421_),
    .Q_N(_14884_),
    .Q(\cpu.dcache.r_data[3][23] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[3][24]$_DFFE_PP_  (.CLK(clknet_leaf_29_clk),
    .RESET_B(net1267),
    .D(_00422_),
    .Q_N(_14883_),
    .Q(\cpu.dcache.r_data[3][24] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[3][25]$_DFFE_PP_  (.CLK(clknet_leaf_273_clk),
    .RESET_B(net1268),
    .D(_00423_),
    .Q_N(_14882_),
    .Q(\cpu.dcache.r_data[3][25] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[3][26]$_DFFE_PP_  (.CLK(clknet_leaf_300_clk),
    .RESET_B(net1269),
    .D(_00424_),
    .Q_N(_14881_),
    .Q(\cpu.dcache.r_data[3][26] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[3][27]$_DFFE_PP_  (.CLK(clknet_leaf_299_clk),
    .RESET_B(net1270),
    .D(_00425_),
    .Q_N(_14880_),
    .Q(\cpu.dcache.r_data[3][27] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[3][28]$_DFFE_PP_  (.CLK(clknet_leaf_300_clk),
    .RESET_B(net1271),
    .D(_00426_),
    .Q_N(_14879_),
    .Q(\cpu.dcache.r_data[3][28] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[3][29]$_DFFE_PP_  (.CLK(clknet_leaf_300_clk),
    .RESET_B(net1272),
    .D(_00427_),
    .Q_N(_14878_),
    .Q(\cpu.dcache.r_data[3][29] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[3][2]$_DFFE_PP_  (.CLK(clknet_leaf_9_clk),
    .RESET_B(net1273),
    .D(_00428_),
    .Q_N(_14877_),
    .Q(\cpu.dcache.r_data[3][2] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[3][30]$_DFFE_PP_  (.CLK(clknet_leaf_300_clk),
    .RESET_B(net1274),
    .D(_00429_),
    .Q_N(_14876_),
    .Q(\cpu.dcache.r_data[3][30] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[3][31]$_DFFE_PP_  (.CLK(clknet_leaf_274_clk),
    .RESET_B(net1275),
    .D(_00430_),
    .Q_N(_14875_),
    .Q(\cpu.dcache.r_data[3][31] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[3][3]$_DFFE_PP_  (.CLK(clknet_leaf_10_clk),
    .RESET_B(net1276),
    .D(_00431_),
    .Q_N(_14874_),
    .Q(\cpu.dcache.r_data[3][3] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[3][4]$_DFFE_PP_  (.CLK(clknet_leaf_10_clk),
    .RESET_B(net1277),
    .D(_00432_),
    .Q_N(_14873_),
    .Q(\cpu.dcache.r_data[3][4] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[3][5]$_DFFE_PP_  (.CLK(clknet_leaf_8_clk),
    .RESET_B(net1278),
    .D(_00433_),
    .Q_N(_14872_),
    .Q(\cpu.dcache.r_data[3][5] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[3][6]$_DFFE_PP_  (.CLK(clknet_leaf_9_clk),
    .RESET_B(net1279),
    .D(_00434_),
    .Q_N(_14871_),
    .Q(\cpu.dcache.r_data[3][6] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[3][7]$_DFFE_PP_  (.CLK(clknet_leaf_10_clk),
    .RESET_B(net1280),
    .D(_00435_),
    .Q_N(_14870_),
    .Q(\cpu.dcache.r_data[3][7] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[3][8]$_DFFE_PP_  (.CLK(clknet_leaf_274_clk),
    .RESET_B(net1281),
    .D(_00436_),
    .Q_N(_14869_),
    .Q(\cpu.dcache.r_data[3][8] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[3][9]$_DFFE_PP_  (.CLK(clknet_leaf_275_clk),
    .RESET_B(net1282),
    .D(_00437_),
    .Q_N(_14868_),
    .Q(\cpu.dcache.r_data[3][9] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[4][0]$_DFFE_PP_  (.CLK(clknet_leaf_306_clk),
    .RESET_B(net1283),
    .D(_00438_),
    .Q_N(_14867_),
    .Q(\cpu.dcache.r_data[4][0] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[4][10]$_DFFE_PP_  (.CLK(clknet_leaf_296_clk),
    .RESET_B(net1284),
    .D(_00439_),
    .Q_N(_14866_),
    .Q(\cpu.dcache.r_data[4][10] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[4][11]$_DFFE_PP_  (.CLK(clknet_leaf_295_clk),
    .RESET_B(net1285),
    .D(_00440_),
    .Q_N(_14865_),
    .Q(\cpu.dcache.r_data[4][11] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[4][12]$_DFFE_PP_  (.CLK(clknet_leaf_294_clk),
    .RESET_B(net1286),
    .D(_00441_),
    .Q_N(_14864_),
    .Q(\cpu.dcache.r_data[4][12] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[4][13]$_DFFE_PP_  (.CLK(clknet_leaf_294_clk),
    .RESET_B(net1287),
    .D(_00442_),
    .Q_N(_14863_),
    .Q(\cpu.dcache.r_data[4][13] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[4][14]$_DFFE_PP_  (.CLK(clknet_leaf_296_clk),
    .RESET_B(net1288),
    .D(_00443_),
    .Q_N(_14862_),
    .Q(\cpu.dcache.r_data[4][14] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[4][15]$_DFFE_PP_  (.CLK(clknet_leaf_297_clk),
    .RESET_B(net1289),
    .D(_00444_),
    .Q_N(_14861_),
    .Q(\cpu.dcache.r_data[4][15] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[4][16]$_DFFE_PP_  (.CLK(clknet_leaf_307_clk),
    .RESET_B(net1290),
    .D(_00445_),
    .Q_N(_14860_),
    .Q(\cpu.dcache.r_data[4][16] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[4][17]$_DFFE_PP_  (.CLK(clknet_leaf_307_clk),
    .RESET_B(net1291),
    .D(_00446_),
    .Q_N(_14859_),
    .Q(\cpu.dcache.r_data[4][17] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[4][18]$_DFFE_PP_  (.CLK(clknet_leaf_304_clk),
    .RESET_B(net1292),
    .D(_00447_),
    .Q_N(_14858_),
    .Q(\cpu.dcache.r_data[4][18] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[4][19]$_DFFE_PP_  (.CLK(clknet_leaf_304_clk),
    .RESET_B(net1293),
    .D(_00448_),
    .Q_N(_14857_),
    .Q(\cpu.dcache.r_data[4][19] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[4][1]$_DFFE_PP_  (.CLK(clknet_leaf_305_clk),
    .RESET_B(net1294),
    .D(_00449_),
    .Q_N(_14856_),
    .Q(\cpu.dcache.r_data[4][1] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[4][20]$_DFFE_PP_  (.CLK(clknet_leaf_11_clk),
    .RESET_B(net1295),
    .D(_00450_),
    .Q_N(_14855_),
    .Q(\cpu.dcache.r_data[4][20] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[4][21]$_DFFE_PP_  (.CLK(clknet_leaf_22_clk),
    .RESET_B(net1296),
    .D(_00451_),
    .Q_N(_14854_),
    .Q(\cpu.dcache.r_data[4][21] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[4][22]$_DFFE_PP_  (.CLK(clknet_leaf_21_clk),
    .RESET_B(net1297),
    .D(_00452_),
    .Q_N(_14853_),
    .Q(\cpu.dcache.r_data[4][22] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[4][23]$_DFFE_PP_  (.CLK(clknet_leaf_25_clk),
    .RESET_B(net1298),
    .D(_00453_),
    .Q_N(_14852_),
    .Q(\cpu.dcache.r_data[4][23] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[4][24]$_DFFE_PP_  (.CLK(clknet_leaf_33_clk),
    .RESET_B(net1299),
    .D(_00454_),
    .Q_N(_14851_),
    .Q(\cpu.dcache.r_data[4][24] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[4][25]$_DFFE_PP_  (.CLK(clknet_leaf_33_clk),
    .RESET_B(net1300),
    .D(_00455_),
    .Q_N(_14850_),
    .Q(\cpu.dcache.r_data[4][25] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[4][26]$_DFFE_PP_  (.CLK(clknet_leaf_33_clk),
    .RESET_B(net1301),
    .D(_00456_),
    .Q_N(_14849_),
    .Q(\cpu.dcache.r_data[4][26] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[4][27]$_DFFE_PP_  (.CLK(clknet_leaf_33_clk),
    .RESET_B(net1302),
    .D(_00457_),
    .Q_N(_14848_),
    .Q(\cpu.dcache.r_data[4][27] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[4][28]$_DFFE_PP_  (.CLK(clknet_leaf_28_clk),
    .RESET_B(net1303),
    .D(_00458_),
    .Q_N(_14847_),
    .Q(\cpu.dcache.r_data[4][28] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[4][29]$_DFFE_PP_  (.CLK(clknet_leaf_300_clk),
    .RESET_B(net1304),
    .D(_00459_),
    .Q_N(_14846_),
    .Q(\cpu.dcache.r_data[4][29] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[4][2]$_DFFE_PP_  (.CLK(clknet_leaf_302_clk),
    .RESET_B(net1305),
    .D(_00460_),
    .Q_N(_14845_),
    .Q(\cpu.dcache.r_data[4][2] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[4][30]$_DFFE_PP_  (.CLK(clknet_leaf_28_clk),
    .RESET_B(net1306),
    .D(_00461_),
    .Q_N(_14844_),
    .Q(\cpu.dcache.r_data[4][30] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[4][31]$_DFFE_PP_  (.CLK(clknet_leaf_28_clk),
    .RESET_B(net1307),
    .D(_00462_),
    .Q_N(_14843_),
    .Q(\cpu.dcache.r_data[4][31] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[4][3]$_DFFE_PP_  (.CLK(clknet_leaf_304_clk),
    .RESET_B(net1308),
    .D(_00463_),
    .Q_N(_14842_),
    .Q(\cpu.dcache.r_data[4][3] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[4][4]$_DFFE_PP_  (.CLK(clknet_leaf_10_clk),
    .RESET_B(net1309),
    .D(_00464_),
    .Q_N(_14841_),
    .Q(\cpu.dcache.r_data[4][4] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[4][5]$_DFFE_PP_  (.CLK(clknet_leaf_10_clk),
    .RESET_B(net1310),
    .D(_00465_),
    .Q_N(_14840_),
    .Q(\cpu.dcache.r_data[4][5] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[4][6]$_DFFE_PP_  (.CLK(clknet_leaf_8_clk),
    .RESET_B(net1311),
    .D(_00466_),
    .Q_N(_14839_),
    .Q(\cpu.dcache.r_data[4][6] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[4][7]$_DFFE_PP_  (.CLK(clknet_leaf_11_clk),
    .RESET_B(net1312),
    .D(_00467_),
    .Q_N(_14838_),
    .Q(\cpu.dcache.r_data[4][7] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[4][8]$_DFFE_PP_  (.CLK(clknet_leaf_296_clk),
    .RESET_B(net1313),
    .D(_00468_),
    .Q_N(_14837_),
    .Q(\cpu.dcache.r_data[4][8] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[4][9]$_DFFE_PP_  (.CLK(clknet_leaf_297_clk),
    .RESET_B(net1314),
    .D(_00469_),
    .Q_N(_14836_),
    .Q(\cpu.dcache.r_data[4][9] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[5][0]$_DFFE_PP_  (.CLK(clknet_leaf_307_clk),
    .RESET_B(net1315),
    .D(_00470_),
    .Q_N(_14835_),
    .Q(\cpu.dcache.r_data[5][0] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[5][10]$_DFFE_PP_  (.CLK(clknet_leaf_304_clk),
    .RESET_B(net1316),
    .D(_00471_),
    .Q_N(_14834_),
    .Q(\cpu.dcache.r_data[5][10] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[5][11]$_DFFE_PP_  (.CLK(clknet_leaf_304_clk),
    .RESET_B(net1317),
    .D(_00472_),
    .Q_N(_14833_),
    .Q(\cpu.dcache.r_data[5][11] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[5][12]$_DFFE_PP_  (.CLK(clknet_leaf_305_clk),
    .RESET_B(net1318),
    .D(_00473_),
    .Q_N(_14832_),
    .Q(\cpu.dcache.r_data[5][12] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[5][13]$_DFFE_PP_  (.CLK(clknet_leaf_306_clk),
    .RESET_B(net1319),
    .D(_00474_),
    .Q_N(_14831_),
    .Q(\cpu.dcache.r_data[5][13] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[5][14]$_DFFE_PP_  (.CLK(clknet_leaf_305_clk),
    .RESET_B(net1320),
    .D(_00475_),
    .Q_N(_14830_),
    .Q(\cpu.dcache.r_data[5][14] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[5][15]$_DFFE_PP_  (.CLK(clknet_leaf_305_clk),
    .RESET_B(net1321),
    .D(_00476_),
    .Q_N(_14829_),
    .Q(\cpu.dcache.r_data[5][15] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[5][16]$_DFFE_PP_  (.CLK(clknet_leaf_9_clk),
    .RESET_B(net1322),
    .D(_00477_),
    .Q_N(_14828_),
    .Q(\cpu.dcache.r_data[5][16] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[5][17]$_DFFE_PP_  (.CLK(clknet_leaf_303_clk),
    .RESET_B(net1323),
    .D(_00478_),
    .Q_N(_14827_),
    .Q(\cpu.dcache.r_data[5][17] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[5][18]$_DFFE_PP_  (.CLK(clknet_leaf_303_clk),
    .RESET_B(net1324),
    .D(_00479_),
    .Q_N(_14826_),
    .Q(\cpu.dcache.r_data[5][18] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[5][19]$_DFFE_PP_  (.CLK(clknet_leaf_303_clk),
    .RESET_B(net1325),
    .D(_00480_),
    .Q_N(_14825_),
    .Q(\cpu.dcache.r_data[5][19] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[5][1]$_DFFE_PP_  (.CLK(clknet_leaf_307_clk),
    .RESET_B(net1326),
    .D(_00481_),
    .Q_N(_14824_),
    .Q(\cpu.dcache.r_data[5][1] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[5][20]$_DFFE_PP_  (.CLK(clknet_leaf_22_clk),
    .RESET_B(net1327),
    .D(_00482_),
    .Q_N(_14823_),
    .Q(\cpu.dcache.r_data[5][20] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[5][21]$_DFFE_PP_  (.CLK(clknet_leaf_21_clk),
    .RESET_B(net1328),
    .D(_00483_),
    .Q_N(_14822_),
    .Q(\cpu.dcache.r_data[5][21] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[5][22]$_DFFE_PP_  (.CLK(clknet_leaf_22_clk),
    .RESET_B(net1329),
    .D(_00484_),
    .Q_N(_14821_),
    .Q(\cpu.dcache.r_data[5][22] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[5][23]$_DFFE_PP_  (.CLK(clknet_leaf_21_clk),
    .RESET_B(net1330),
    .D(_00485_),
    .Q_N(_14820_),
    .Q(\cpu.dcache.r_data[5][23] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[5][24]$_DFFE_PP_  (.CLK(clknet_leaf_301_clk),
    .RESET_B(net1331),
    .D(_00486_),
    .Q_N(_14819_),
    .Q(\cpu.dcache.r_data[5][24] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[5][25]$_DFFE_PP_  (.CLK(clknet_leaf_27_clk),
    .RESET_B(net1332),
    .D(_00487_),
    .Q_N(_14818_),
    .Q(\cpu.dcache.r_data[5][25] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[5][26]$_DFFE_PP_  (.CLK(clknet_leaf_9_clk),
    .RESET_B(net1333),
    .D(_00488_),
    .Q_N(_14817_),
    .Q(\cpu.dcache.r_data[5][26] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[5][27]$_DFFE_PP_  (.CLK(clknet_leaf_28_clk),
    .RESET_B(net1334),
    .D(_00489_),
    .Q_N(_14816_),
    .Q(\cpu.dcache.r_data[5][27] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[5][28]$_DFFE_PP_  (.CLK(clknet_leaf_301_clk),
    .RESET_B(net1335),
    .D(_00490_),
    .Q_N(_14815_),
    .Q(\cpu.dcache.r_data[5][28] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[5][29]$_DFFE_PP_  (.CLK(clknet_leaf_301_clk),
    .RESET_B(net1336),
    .D(_00491_),
    .Q_N(_14814_),
    .Q(\cpu.dcache.r_data[5][29] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[5][2]$_DFFE_PP_  (.CLK(clknet_leaf_308_clk),
    .RESET_B(net1337),
    .D(_00492_),
    .Q_N(_14813_),
    .Q(\cpu.dcache.r_data[5][2] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[5][30]$_DFFE_PP_  (.CLK(clknet_leaf_301_clk),
    .RESET_B(net1338),
    .D(_00493_),
    .Q_N(_14812_),
    .Q(\cpu.dcache.r_data[5][30] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[5][31]$_DFFE_PP_  (.CLK(clknet_leaf_301_clk),
    .RESET_B(net1339),
    .D(_00494_),
    .Q_N(_14811_),
    .Q(\cpu.dcache.r_data[5][31] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[5][3]$_DFFE_PP_  (.CLK(clknet_leaf_308_clk),
    .RESET_B(net1340),
    .D(_00495_),
    .Q_N(_14810_),
    .Q(\cpu.dcache.r_data[5][3] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[5][4]$_DFFE_PP_  (.CLK(clknet_leaf_9_clk),
    .RESET_B(net1341),
    .D(_00496_),
    .Q_N(_14809_),
    .Q(\cpu.dcache.r_data[5][4] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[5][5]$_DFFE_PP_  (.CLK(clknet_leaf_7_clk),
    .RESET_B(net1342),
    .D(_00497_),
    .Q_N(_14808_),
    .Q(\cpu.dcache.r_data[5][5] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[5][6]$_DFFE_PP_  (.CLK(clknet_leaf_8_clk),
    .RESET_B(net1343),
    .D(_00498_),
    .Q_N(_14807_),
    .Q(\cpu.dcache.r_data[5][6] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[5][7]$_DFFE_PP_  (.CLK(clknet_leaf_7_clk),
    .RESET_B(net1344),
    .D(_00499_),
    .Q_N(_14806_),
    .Q(\cpu.dcache.r_data[5][7] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[5][8]$_DFFE_PP_  (.CLK(clknet_leaf_306_clk),
    .RESET_B(net1345),
    .D(_00500_),
    .Q_N(_14805_),
    .Q(\cpu.dcache.r_data[5][8] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[5][9]$_DFFE_PP_  (.CLK(clknet_leaf_306_clk),
    .RESET_B(net1346),
    .D(_00501_),
    .Q_N(_14804_),
    .Q(\cpu.dcache.r_data[5][9] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[6][0]$_DFFE_PP_  (.CLK(clknet_leaf_306_clk),
    .RESET_B(net1347),
    .D(_00502_),
    .Q_N(_14803_),
    .Q(\cpu.dcache.r_data[6][0] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[6][10]$_DFFE_PP_  (.CLK(clknet_leaf_296_clk),
    .RESET_B(net1348),
    .D(_00503_),
    .Q_N(_14802_),
    .Q(\cpu.dcache.r_data[6][10] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[6][11]$_DFFE_PP_  (.CLK(clknet_leaf_296_clk),
    .RESET_B(net1349),
    .D(_00504_),
    .Q_N(_14801_),
    .Q(\cpu.dcache.r_data[6][11] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[6][12]$_DFFE_PP_  (.CLK(clknet_leaf_295_clk),
    .RESET_B(net1350),
    .D(_00505_),
    .Q_N(_14800_),
    .Q(\cpu.dcache.r_data[6][12] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[6][13]$_DFFE_PP_  (.CLK(clknet_leaf_295_clk),
    .RESET_B(net1351),
    .D(_00506_),
    .Q_N(_14799_),
    .Q(\cpu.dcache.r_data[6][13] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[6][14]$_DFFE_PP_  (.CLK(clknet_leaf_296_clk),
    .RESET_B(net1352),
    .D(_00507_),
    .Q_N(_14798_),
    .Q(\cpu.dcache.r_data[6][14] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[6][15]$_DFFE_PP_  (.CLK(clknet_leaf_296_clk),
    .RESET_B(net1353),
    .D(_00508_),
    .Q_N(_14797_),
    .Q(\cpu.dcache.r_data[6][15] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[6][16]$_DFFE_PP_  (.CLK(clknet_leaf_307_clk),
    .RESET_B(net1354),
    .D(_00509_),
    .Q_N(_14796_),
    .Q(\cpu.dcache.r_data[6][16] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[6][17]$_DFFE_PP_  (.CLK(clknet_leaf_306_clk),
    .RESET_B(net1355),
    .D(_00510_),
    .Q_N(_14795_),
    .Q(\cpu.dcache.r_data[6][17] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[6][18]$_DFFE_PP_  (.CLK(clknet_leaf_304_clk),
    .RESET_B(net1356),
    .D(_00511_),
    .Q_N(_14794_),
    .Q(\cpu.dcache.r_data[6][18] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[6][19]$_DFFE_PP_  (.CLK(clknet_leaf_304_clk),
    .RESET_B(net1357),
    .D(_00512_),
    .Q_N(_14793_),
    .Q(\cpu.dcache.r_data[6][19] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[6][1]$_DFFE_PP_  (.CLK(clknet_leaf_306_clk),
    .RESET_B(net1358),
    .D(_00513_),
    .Q_N(_14792_),
    .Q(\cpu.dcache.r_data[6][1] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[6][20]$_DFFE_PP_  (.CLK(clknet_leaf_12_clk),
    .RESET_B(net1359),
    .D(_00514_),
    .Q_N(_14791_),
    .Q(\cpu.dcache.r_data[6][20] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[6][21]$_DFFE_PP_  (.CLK(clknet_leaf_26_clk),
    .RESET_B(net1360),
    .D(_00515_),
    .Q_N(_14790_),
    .Q(\cpu.dcache.r_data[6][21] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[6][22]$_DFFE_PP_  (.CLK(clknet_leaf_21_clk),
    .RESET_B(net1361),
    .D(_00516_),
    .Q_N(_14789_),
    .Q(\cpu.dcache.r_data[6][22] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[6][23]$_DFFE_PP_  (.CLK(clknet_leaf_25_clk),
    .RESET_B(net1362),
    .D(_00517_),
    .Q_N(_14788_),
    .Q(\cpu.dcache.r_data[6][23] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[6][24]$_DFFE_PP_  (.CLK(clknet_leaf_301_clk),
    .RESET_B(net1363),
    .D(_00518_),
    .Q_N(_14787_),
    .Q(\cpu.dcache.r_data[6][24] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[6][25]$_DFFE_PP_  (.CLK(clknet_leaf_28_clk),
    .RESET_B(net1364),
    .D(_00519_),
    .Q_N(_14786_),
    .Q(\cpu.dcache.r_data[6][25] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[6][26]$_DFFE_PP_  (.CLK(clknet_leaf_301_clk),
    .RESET_B(net1365),
    .D(_00520_),
    .Q_N(_14785_),
    .Q(\cpu.dcache.r_data[6][26] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[6][27]$_DFFE_PP_  (.CLK(clknet_leaf_300_clk),
    .RESET_B(net1366),
    .D(_00521_),
    .Q_N(_14784_),
    .Q(\cpu.dcache.r_data[6][27] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[6][28]$_DFFE_PP_  (.CLK(clknet_leaf_300_clk),
    .RESET_B(net1367),
    .D(_00522_),
    .Q_N(_14783_),
    .Q(\cpu.dcache.r_data[6][28] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[6][29]$_DFFE_PP_  (.CLK(clknet_leaf_299_clk),
    .RESET_B(net1368),
    .D(_00523_),
    .Q_N(_14782_),
    .Q(\cpu.dcache.r_data[6][29] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[6][2]$_DFFE_PP_  (.CLK(clknet_leaf_302_clk),
    .RESET_B(net1369),
    .D(_00524_),
    .Q_N(_14781_),
    .Q(\cpu.dcache.r_data[6][2] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[6][30]$_DFFE_PP_  (.CLK(clknet_leaf_299_clk),
    .RESET_B(net1370),
    .D(_00525_),
    .Q_N(_14780_),
    .Q(\cpu.dcache.r_data[6][30] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[6][31]$_DFFE_PP_  (.CLK(clknet_leaf_300_clk),
    .RESET_B(net1371),
    .D(_00526_),
    .Q_N(_14779_),
    .Q(\cpu.dcache.r_data[6][31] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[6][3]$_DFFE_PP_  (.CLK(clknet_leaf_301_clk),
    .RESET_B(net1372),
    .D(_00527_),
    .Q_N(_14778_),
    .Q(\cpu.dcache.r_data[6][3] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[6][4]$_DFFE_PP_  (.CLK(clknet_leaf_8_clk),
    .RESET_B(net1373),
    .D(_00528_),
    .Q_N(_14777_),
    .Q(\cpu.dcache.r_data[6][4] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[6][5]$_DFFE_PP_  (.CLK(clknet_leaf_7_clk),
    .RESET_B(net1374),
    .D(_00529_),
    .Q_N(_14776_),
    .Q(\cpu.dcache.r_data[6][5] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[6][6]$_DFFE_PP_  (.CLK(clknet_leaf_8_clk),
    .RESET_B(net1375),
    .D(_00530_),
    .Q_N(_14775_),
    .Q(\cpu.dcache.r_data[6][6] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[6][7]$_DFFE_PP_  (.CLK(clknet_leaf_7_clk),
    .RESET_B(net1376),
    .D(_00531_),
    .Q_N(_14774_),
    .Q(\cpu.dcache.r_data[6][7] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[6][8]$_DFFE_PP_  (.CLK(clknet_leaf_295_clk),
    .RESET_B(net1377),
    .D(_00532_),
    .Q_N(_14773_),
    .Q(\cpu.dcache.r_data[6][8] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[6][9]$_DFFE_PP_  (.CLK(clknet_leaf_295_clk),
    .RESET_B(net1378),
    .D(_00533_),
    .Q_N(_14772_),
    .Q(\cpu.dcache.r_data[6][9] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[7][0]$_DFFE_PP_  (.CLK(clknet_leaf_302_clk),
    .RESET_B(net1379),
    .D(_00534_),
    .Q_N(_14771_),
    .Q(\cpu.dcache.r_data[7][0] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[7][10]$_DFFE_PP_  (.CLK(clknet_leaf_305_clk),
    .RESET_B(net1380),
    .D(_00535_),
    .Q_N(_14770_),
    .Q(\cpu.dcache.r_data[7][10] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[7][11]$_DFFE_PP_  (.CLK(clknet_leaf_295_clk),
    .RESET_B(net1381),
    .D(_00536_),
    .Q_N(_14769_),
    .Q(\cpu.dcache.r_data[7][11] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[7][12]$_DFFE_PP_  (.CLK(clknet_leaf_295_clk),
    .RESET_B(net1382),
    .D(_00537_),
    .Q_N(_14768_),
    .Q(\cpu.dcache.r_data[7][12] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[7][13]$_DFFE_PP_  (.CLK(clknet_leaf_306_clk),
    .RESET_B(net1383),
    .D(_00538_),
    .Q_N(_14767_),
    .Q(\cpu.dcache.r_data[7][13] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[7][14]$_DFFE_PP_  (.CLK(clknet_leaf_305_clk),
    .RESET_B(net1384),
    .D(_00539_),
    .Q_N(_14766_),
    .Q(\cpu.dcache.r_data[7][14] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[7][15]$_DFFE_PP_  (.CLK(clknet_leaf_296_clk),
    .RESET_B(net1385),
    .D(_00540_),
    .Q_N(_14765_),
    .Q(\cpu.dcache.r_data[7][15] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[7][16]$_DFFE_PP_  (.CLK(clknet_leaf_307_clk),
    .RESET_B(net1386),
    .D(_00541_),
    .Q_N(_14764_),
    .Q(\cpu.dcache.r_data[7][16] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[7][17]$_DFFE_PP_  (.CLK(clknet_leaf_305_clk),
    .RESET_B(net1387),
    .D(_00542_),
    .Q_N(_14763_),
    .Q(\cpu.dcache.r_data[7][17] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[7][18]$_DFFE_PP_  (.CLK(clknet_leaf_308_clk),
    .RESET_B(net1388),
    .D(_00543_),
    .Q_N(_14762_),
    .Q(\cpu.dcache.r_data[7][18] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[7][19]$_DFFE_PP_  (.CLK(clknet_leaf_304_clk),
    .RESET_B(net1389),
    .D(_00544_),
    .Q_N(_14761_),
    .Q(\cpu.dcache.r_data[7][19] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[7][1]$_DFFE_PP_  (.CLK(clknet_leaf_303_clk),
    .RESET_B(net1390),
    .D(_00545_),
    .Q_N(_14760_),
    .Q(\cpu.dcache.r_data[7][1] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[7][20]$_DFFE_PP_  (.CLK(clknet_leaf_11_clk),
    .RESET_B(net1391),
    .D(_00546_),
    .Q_N(_14759_),
    .Q(\cpu.dcache.r_data[7][20] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[7][21]$_DFFE_PP_  (.CLK(clknet_leaf_11_clk),
    .RESET_B(net1392),
    .D(_00547_),
    .Q_N(_14758_),
    .Q(\cpu.dcache.r_data[7][21] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[7][22]$_DFFE_PP_  (.CLK(clknet_leaf_26_clk),
    .RESET_B(net1393),
    .D(_00548_),
    .Q_N(_14757_),
    .Q(\cpu.dcache.r_data[7][22] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[7][23]$_DFFE_PP_  (.CLK(clknet_leaf_26_clk),
    .RESET_B(net1394),
    .D(_00549_),
    .Q_N(_14756_),
    .Q(\cpu.dcache.r_data[7][23] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[7][24]$_DFFE_PP_  (.CLK(clknet_leaf_302_clk),
    .RESET_B(net1395),
    .D(_00550_),
    .Q_N(_14755_),
    .Q(\cpu.dcache.r_data[7][24] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[7][25]$_DFFE_PP_  (.CLK(clknet_leaf_28_clk),
    .RESET_B(net1396),
    .D(_00551_),
    .Q_N(_14754_),
    .Q(\cpu.dcache.r_data[7][25] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[7][26]$_DFFE_PP_  (.CLK(clknet_leaf_9_clk),
    .RESET_B(net1397),
    .D(_00552_),
    .Q_N(_14753_),
    .Q(\cpu.dcache.r_data[7][26] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[7][27]$_DFFE_PP_  (.CLK(clknet_leaf_28_clk),
    .RESET_B(net1398),
    .D(_00553_),
    .Q_N(_14752_),
    .Q(\cpu.dcache.r_data[7][27] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[7][28]$_DFFE_PP_  (.CLK(clknet_leaf_302_clk),
    .RESET_B(net1399),
    .D(_00554_),
    .Q_N(_14751_),
    .Q(\cpu.dcache.r_data[7][28] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[7][29]$_DFFE_PP_  (.CLK(clknet_leaf_302_clk),
    .RESET_B(net1400),
    .D(_00555_),
    .Q_N(_14750_),
    .Q(\cpu.dcache.r_data[7][29] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[7][2]$_DFFE_PP_  (.CLK(clknet_leaf_303_clk),
    .RESET_B(net1401),
    .D(_00556_),
    .Q_N(_14749_),
    .Q(\cpu.dcache.r_data[7][2] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[7][30]$_DFFE_PP_  (.CLK(clknet_leaf_302_clk),
    .RESET_B(net1402),
    .D(_00557_),
    .Q_N(_14748_),
    .Q(\cpu.dcache.r_data[7][30] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[7][31]$_DFFE_PP_  (.CLK(clknet_leaf_302_clk),
    .RESET_B(net1403),
    .D(_00558_),
    .Q_N(_14747_),
    .Q(\cpu.dcache.r_data[7][31] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[7][3]$_DFFE_PP_  (.CLK(clknet_leaf_303_clk),
    .RESET_B(net1404),
    .D(_00559_),
    .Q_N(_14746_),
    .Q(\cpu.dcache.r_data[7][3] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[7][4]$_DFFE_PP_  (.CLK(clknet_leaf_11_clk),
    .RESET_B(net1405),
    .D(_00560_),
    .Q_N(_14745_),
    .Q(\cpu.dcache.r_data[7][4] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[7][5]$_DFFE_PP_  (.CLK(clknet_leaf_8_clk),
    .RESET_B(net1406),
    .D(_00561_),
    .Q_N(_14744_),
    .Q(\cpu.dcache.r_data[7][5] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[7][6]$_DFFE_PP_  (.CLK(clknet_leaf_8_clk),
    .RESET_B(net1407),
    .D(_00562_),
    .Q_N(_14743_),
    .Q(\cpu.dcache.r_data[7][6] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[7][7]$_DFFE_PP_  (.CLK(clknet_leaf_10_clk),
    .RESET_B(net1408),
    .D(_00563_),
    .Q_N(_14742_),
    .Q(\cpu.dcache.r_data[7][7] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[7][8]$_DFFE_PP_  (.CLK(clknet_leaf_305_clk),
    .RESET_B(net1409),
    .D(_00564_),
    .Q_N(_14741_),
    .Q(\cpu.dcache.r_data[7][8] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[7][9]$_DFFE_PP_  (.CLK(clknet_leaf_295_clk),
    .RESET_B(net1410),
    .D(_00565_),
    .Q_N(_14740_),
    .Q(\cpu.dcache.r_data[7][9] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_dirty[0]$_SDFFCE_PP1P_  (.CLK(clknet_leaf_50_clk),
    .RESET_B(net1411),
    .D(_00566_),
    .Q_N(_14739_),
    .Q(\cpu.dcache.r_dirty[0] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_dirty[1]$_SDFFCE_PP1P_  (.CLK(clknet_leaf_50_clk),
    .RESET_B(net1412),
    .D(_00567_),
    .Q_N(_14738_),
    .Q(\cpu.dcache.r_dirty[1] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_dirty[2]$_SDFFCE_PP1P_  (.CLK(clknet_leaf_47_clk),
    .RESET_B(net1413),
    .D(_00568_),
    .Q_N(_14737_),
    .Q(\cpu.dcache.r_dirty[2] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_dirty[3]$_SDFFCE_PP1P_  (.CLK(clknet_leaf_49_clk),
    .RESET_B(net1414),
    .D(_00569_),
    .Q_N(_14736_),
    .Q(\cpu.dcache.r_dirty[3] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_dirty[4]$_SDFFCE_PP1P_  (.CLK(clknet_leaf_51_clk),
    .RESET_B(net1415),
    .D(_00570_),
    .Q_N(_14735_),
    .Q(\cpu.dcache.r_dirty[4] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_dirty[5]$_SDFFCE_PP1P_  (.CLK(clknet_leaf_51_clk),
    .RESET_B(net1416),
    .D(_00571_),
    .Q_N(_14734_),
    .Q(\cpu.dcache.r_dirty[5] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_dirty[6]$_SDFFCE_PP1P_  (.CLK(clknet_leaf_50_clk),
    .RESET_B(net1417),
    .D(_00572_),
    .Q_N(_14733_),
    .Q(\cpu.dcache.r_dirty[6] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_dirty[7]$_SDFFCE_PP1P_  (.CLK(clknet_leaf_51_clk),
    .RESET_B(net1418),
    .D(_00573_),
    .Q_N(_14732_),
    .Q(\cpu.dcache.r_dirty[7] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_offset[0]$_SDFF_PN0_  (.CLK(clknet_leaf_52_clk),
    .RESET_B(net1419),
    .D(_00574_),
    .Q_N(_00303_),
    .Q(\cpu.dcache.r_offset[0] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_offset[1]$_SDFF_PN0_  (.CLK(clknet_leaf_52_clk),
    .RESET_B(net1420),
    .D(_00575_),
    .Q_N(_14731_),
    .Q(\cpu.dcache.r_offset[1] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_offset[2]$_SDFF_PN0_  (.CLK(clknet_leaf_52_clk),
    .RESET_B(net1421),
    .D(_00576_),
    .Q_N(_00260_),
    .Q(\cpu.dcache.r_offset[2] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[0][0]$_DFFE_PP_  (.CLK(clknet_leaf_106_clk),
    .RESET_B(net1422),
    .D(_00577_),
    .Q_N(_00214_),
    .Q(\cpu.dcache.r_tag[0][5] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[0][10]$_DFFE_PP_  (.CLK(clknet_leaf_108_clk),
    .RESET_B(net1423),
    .D(_00578_),
    .Q_N(_00230_),
    .Q(\cpu.dcache.r_tag[0][15] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[0][11]$_DFFE_PP_  (.CLK(clknet_leaf_89_clk),
    .RESET_B(net1424),
    .D(_00579_),
    .Q_N(_00231_),
    .Q(\cpu.dcache.r_tag[0][16] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[0][12]$_DFFE_PP_  (.CLK(clknet_leaf_107_clk),
    .RESET_B(net1425),
    .D(_00580_),
    .Q_N(_00232_),
    .Q(\cpu.dcache.r_tag[0][17] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[0][13]$_DFFE_PP_  (.CLK(clknet_leaf_88_clk),
    .RESET_B(net1426),
    .D(_00581_),
    .Q_N(_00233_),
    .Q(\cpu.dcache.r_tag[0][18] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[0][14]$_DFFE_PP_  (.CLK(clknet_leaf_88_clk),
    .RESET_B(net1427),
    .D(_00582_),
    .Q_N(_00234_),
    .Q(\cpu.dcache.r_tag[0][19] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[0][15]$_DFFE_PP_  (.CLK(clknet_leaf_88_clk),
    .RESET_B(net1428),
    .D(_00583_),
    .Q_N(_14730_),
    .Q(\cpu.dcache.r_tag[0][20] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[0][16]$_DFFE_PP_  (.CLK(clknet_leaf_107_clk),
    .RESET_B(net1429),
    .D(_00584_),
    .Q_N(_14729_),
    .Q(\cpu.dcache.r_tag[0][21] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[0][17]$_DFFE_PP_  (.CLK(clknet_leaf_88_clk),
    .RESET_B(net1430),
    .D(_00585_),
    .Q_N(_14728_),
    .Q(\cpu.dcache.r_tag[0][22] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[0][18]$_DFFE_PP_  (.CLK(clknet_leaf_107_clk),
    .RESET_B(net1431),
    .D(_00586_),
    .Q_N(_00235_),
    .Q(\cpu.dcache.r_tag[0][23] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[0][1]$_DFFE_PP_  (.CLK(clknet_leaf_108_clk),
    .RESET_B(net1432),
    .D(_00587_),
    .Q_N(_00216_),
    .Q(\cpu.dcache.r_tag[0][6] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[0][2]$_DFFE_PP_  (.CLK(clknet_leaf_106_clk),
    .RESET_B(net1433),
    .D(_00588_),
    .Q_N(_00218_),
    .Q(\cpu.dcache.r_tag[0][7] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[0][3]$_DFFE_PP_  (.CLK(clknet_leaf_106_clk),
    .RESET_B(net1434),
    .D(_00589_),
    .Q_N(_00220_),
    .Q(\cpu.dcache.r_tag[0][8] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[0][4]$_DFFE_PP_  (.CLK(clknet_leaf_107_clk),
    .RESET_B(net1435),
    .D(_00590_),
    .Q_N(_00222_),
    .Q(\cpu.dcache.r_tag[0][9] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[0][5]$_DFFE_PP_  (.CLK(clknet_leaf_109_clk),
    .RESET_B(net1436),
    .D(_00591_),
    .Q_N(_00224_),
    .Q(\cpu.dcache.r_tag[0][10] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[0][6]$_DFFE_PP_  (.CLK(clknet_leaf_108_clk),
    .RESET_B(net1437),
    .D(_00592_),
    .Q_N(_00226_),
    .Q(\cpu.dcache.r_tag[0][11] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[0][7]$_DFFE_PP_  (.CLK(clknet_leaf_107_clk),
    .RESET_B(net1438),
    .D(_00593_),
    .Q_N(_00227_),
    .Q(\cpu.dcache.r_tag[0][12] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[0][8]$_DFFE_PP_  (.CLK(clknet_leaf_87_clk),
    .RESET_B(net1439),
    .D(_00594_),
    .Q_N(_00228_),
    .Q(\cpu.dcache.r_tag[0][13] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[0][9]$_DFFE_PP_  (.CLK(clknet_leaf_108_clk),
    .RESET_B(net1440),
    .D(_00595_),
    .Q_N(_00229_),
    .Q(\cpu.dcache.r_tag[0][14] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[1][0]$_DFFE_PP_  (.CLK(clknet_leaf_94_clk),
    .RESET_B(net1441),
    .D(_00596_),
    .Q_N(_14727_),
    .Q(\cpu.dcache.r_tag[1][5] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[1][10]$_DFFE_PP_  (.CLK(clknet_leaf_108_clk),
    .RESET_B(net1442),
    .D(_00597_),
    .Q_N(_14726_),
    .Q(\cpu.dcache.r_tag[1][15] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[1][11]$_DFFE_PP_  (.CLK(clknet_leaf_90_clk),
    .RESET_B(net1443),
    .D(_00598_),
    .Q_N(_14725_),
    .Q(\cpu.dcache.r_tag[1][16] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[1][12]$_DFFE_PP_  (.CLK(clknet_leaf_89_clk),
    .RESET_B(net1444),
    .D(_00599_),
    .Q_N(_14724_),
    .Q(\cpu.dcache.r_tag[1][17] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[1][13]$_DFFE_PP_  (.CLK(clknet_leaf_91_clk),
    .RESET_B(net1445),
    .D(_00600_),
    .Q_N(_14723_),
    .Q(\cpu.dcache.r_tag[1][18] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[1][14]$_DFFE_PP_  (.CLK(clknet_leaf_88_clk),
    .RESET_B(net1446),
    .D(_00601_),
    .Q_N(_14722_),
    .Q(\cpu.dcache.r_tag[1][19] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[1][15]$_DFFE_PP_  (.CLK(clknet_leaf_93_clk),
    .RESET_B(net1447),
    .D(_00602_),
    .Q_N(_14721_),
    .Q(\cpu.dcache.r_tag[1][20] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[1][16]$_DFFE_PP_  (.CLK(clknet_leaf_87_clk),
    .RESET_B(net1448),
    .D(_00603_),
    .Q_N(_14720_),
    .Q(\cpu.dcache.r_tag[1][21] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[1][17]$_DFFE_PP_  (.CLK(clknet_leaf_92_clk),
    .RESET_B(net1449),
    .D(_00604_),
    .Q_N(_14719_),
    .Q(\cpu.dcache.r_tag[1][22] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[1][18]$_DFFE_PP_  (.CLK(clknet_leaf_89_clk),
    .RESET_B(net1450),
    .D(_00605_),
    .Q_N(_14718_),
    .Q(\cpu.dcache.r_tag[1][23] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[1][1]$_DFFE_PP_  (.CLK(clknet_leaf_48_clk),
    .RESET_B(net1451),
    .D(_00606_),
    .Q_N(_14717_),
    .Q(\cpu.dcache.r_tag[1][6] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[1][2]$_DFFE_PP_  (.CLK(clknet_leaf_95_clk),
    .RESET_B(net1452),
    .D(_00607_),
    .Q_N(_14716_),
    .Q(\cpu.dcache.r_tag[1][7] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[1][3]$_DFFE_PP_  (.CLK(clknet_leaf_94_clk),
    .RESET_B(net1453),
    .D(_00608_),
    .Q_N(_14715_),
    .Q(\cpu.dcache.r_tag[1][8] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[1][4]$_DFFE_PP_  (.CLK(clknet_leaf_106_clk),
    .RESET_B(net1454),
    .D(_00609_),
    .Q_N(_14714_),
    .Q(\cpu.dcache.r_tag[1][9] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[1][5]$_DFFE_PP_  (.CLK(clknet_leaf_109_clk),
    .RESET_B(net1455),
    .D(_00610_),
    .Q_N(_14713_),
    .Q(\cpu.dcache.r_tag[1][10] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[1][6]$_DFFE_PP_  (.CLK(clknet_leaf_48_clk),
    .RESET_B(net1456),
    .D(_00611_),
    .Q_N(_14712_),
    .Q(\cpu.dcache.r_tag[1][11] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[1][7]$_DFFE_PP_  (.CLK(clknet_leaf_86_clk),
    .RESET_B(net1457),
    .D(_00612_),
    .Q_N(_14711_),
    .Q(\cpu.dcache.r_tag[1][12] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[1][8]$_DFFE_PP_  (.CLK(clknet_leaf_91_clk),
    .RESET_B(net1458),
    .D(_00613_),
    .Q_N(_14710_),
    .Q(\cpu.dcache.r_tag[1][13] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[1][9]$_DFFE_PP_  (.CLK(clknet_leaf_108_clk),
    .RESET_B(net1459),
    .D(_00614_),
    .Q_N(_14709_),
    .Q(\cpu.dcache.r_tag[1][14] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[2][0]$_DFFE_PP_  (.CLK(clknet_leaf_106_clk),
    .RESET_B(net1460),
    .D(_00615_),
    .Q_N(_14708_),
    .Q(\cpu.dcache.r_tag[2][5] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[2][10]$_DFFE_PP_  (.CLK(clknet_leaf_107_clk),
    .RESET_B(net1461),
    .D(_00616_),
    .Q_N(_14707_),
    .Q(\cpu.dcache.r_tag[2][15] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[2][11]$_DFFE_PP_  (.CLK(clknet_leaf_90_clk),
    .RESET_B(net1462),
    .D(_00617_),
    .Q_N(_14706_),
    .Q(\cpu.dcache.r_tag[2][16] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[2][12]$_DFFE_PP_  (.CLK(clknet_leaf_106_clk),
    .RESET_B(net1463),
    .D(_00618_),
    .Q_N(_14705_),
    .Q(\cpu.dcache.r_tag[2][17] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[2][13]$_DFFE_PP_  (.CLK(clknet_leaf_92_clk),
    .RESET_B(net1464),
    .D(_00619_),
    .Q_N(_14704_),
    .Q(\cpu.dcache.r_tag[2][18] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[2][14]$_DFFE_PP_  (.CLK(clknet_leaf_88_clk),
    .RESET_B(net1465),
    .D(_00620_),
    .Q_N(_14703_),
    .Q(\cpu.dcache.r_tag[2][19] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[2][15]$_DFFE_PP_  (.CLK(clknet_leaf_91_clk),
    .RESET_B(net1466),
    .D(_00621_),
    .Q_N(_14702_),
    .Q(\cpu.dcache.r_tag[2][20] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[2][16]$_DFFE_PP_  (.CLK(clknet_leaf_87_clk),
    .RESET_B(net1467),
    .D(_00622_),
    .Q_N(_14701_),
    .Q(\cpu.dcache.r_tag[2][21] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[2][17]$_DFFE_PP_  (.CLK(clknet_leaf_91_clk),
    .RESET_B(net1468),
    .D(_00623_),
    .Q_N(_14700_),
    .Q(\cpu.dcache.r_tag[2][22] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[2][18]$_DFFE_PP_  (.CLK(clknet_leaf_89_clk),
    .RESET_B(net1469),
    .D(_00624_),
    .Q_N(_14699_),
    .Q(\cpu.dcache.r_tag[2][23] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[2][1]$_DFFE_PP_  (.CLK(clknet_leaf_45_clk),
    .RESET_B(net1470),
    .D(_00625_),
    .Q_N(_14698_),
    .Q(\cpu.dcache.r_tag[2][6] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[2][2]$_DFFE_PP_  (.CLK(clknet_leaf_104_clk),
    .RESET_B(net1471),
    .D(_00626_),
    .Q_N(_14697_),
    .Q(\cpu.dcache.r_tag[2][7] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[2][3]$_DFFE_PP_  (.CLK(clknet_leaf_104_clk),
    .RESET_B(net1472),
    .D(_00627_),
    .Q_N(_14696_),
    .Q(\cpu.dcache.r_tag[2][8] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[2][4]$_DFFE_PP_  (.CLK(clknet_leaf_95_clk),
    .RESET_B(net1473),
    .D(_00628_),
    .Q_N(_14695_),
    .Q(\cpu.dcache.r_tag[2][9] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[2][5]$_DFFE_PP_  (.CLK(clknet_leaf_48_clk),
    .RESET_B(net1474),
    .D(_00629_),
    .Q_N(_14694_),
    .Q(\cpu.dcache.r_tag[2][10] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[2][6]$_DFFE_PP_  (.CLK(clknet_leaf_44_clk),
    .RESET_B(net1475),
    .D(_00630_),
    .Q_N(_14693_),
    .Q(\cpu.dcache.r_tag[2][11] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[2][7]$_DFFE_PP_  (.CLK(clknet_leaf_86_clk),
    .RESET_B(net1476),
    .D(_00631_),
    .Q_N(_14692_),
    .Q(\cpu.dcache.r_tag[2][12] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[2][8]$_DFFE_PP_  (.CLK(clknet_leaf_82_clk),
    .RESET_B(net1477),
    .D(_00632_),
    .Q_N(_14691_),
    .Q(\cpu.dcache.r_tag[2][13] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[2][9]$_DFFE_PP_  (.CLK(clknet_leaf_47_clk),
    .RESET_B(net1478),
    .D(_00633_),
    .Q_N(_14690_),
    .Q(\cpu.dcache.r_tag[2][14] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[3][0]$_DFFE_PP_  (.CLK(clknet_leaf_94_clk),
    .RESET_B(net1479),
    .D(_00634_),
    .Q_N(_14689_),
    .Q(\cpu.dcache.r_tag[3][5] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[3][10]$_DFFE_PP_  (.CLK(clknet_leaf_108_clk),
    .RESET_B(net1480),
    .D(_00635_),
    .Q_N(_14688_),
    .Q(\cpu.dcache.r_tag[3][15] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[3][11]$_DFFE_PP_  (.CLK(clknet_leaf_90_clk),
    .RESET_B(net1481),
    .D(_00636_),
    .Q_N(_14687_),
    .Q(\cpu.dcache.r_tag[3][16] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[3][12]$_DFFE_PP_  (.CLK(clknet_leaf_89_clk),
    .RESET_B(net1482),
    .D(_00637_),
    .Q_N(_14686_),
    .Q(\cpu.dcache.r_tag[3][17] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[3][13]$_DFFE_PP_  (.CLK(clknet_leaf_91_clk),
    .RESET_B(net1483),
    .D(_00638_),
    .Q_N(_14685_),
    .Q(\cpu.dcache.r_tag[3][18] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[3][14]$_DFFE_PP_  (.CLK(clknet_leaf_87_clk),
    .RESET_B(net1484),
    .D(_00639_),
    .Q_N(_14684_),
    .Q(\cpu.dcache.r_tag[3][19] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[3][15]$_DFFE_PP_  (.CLK(clknet_leaf_92_clk),
    .RESET_B(net1485),
    .D(_00640_),
    .Q_N(_14683_),
    .Q(\cpu.dcache.r_tag[3][20] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[3][16]$_DFFE_PP_  (.CLK(clknet_leaf_107_clk),
    .RESET_B(net1486),
    .D(_00641_),
    .Q_N(_14682_),
    .Q(\cpu.dcache.r_tag[3][21] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[3][17]$_DFFE_PP_  (.CLK(clknet_leaf_92_clk),
    .RESET_B(net1487),
    .D(_00642_),
    .Q_N(_14681_),
    .Q(\cpu.dcache.r_tag[3][22] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[3][18]$_DFFE_PP_  (.CLK(clknet_leaf_90_clk),
    .RESET_B(net1488),
    .D(_00643_),
    .Q_N(_14680_),
    .Q(\cpu.dcache.r_tag[3][23] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[3][1]$_DFFE_PP_  (.CLK(clknet_leaf_49_clk),
    .RESET_B(net1489),
    .D(_00644_),
    .Q_N(_14679_),
    .Q(\cpu.dcache.r_tag[3][6] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[3][2]$_DFFE_PP_  (.CLK(clknet_leaf_97_clk),
    .RESET_B(net1490),
    .D(_00645_),
    .Q_N(_14678_),
    .Q(\cpu.dcache.r_tag[3][7] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[3][3]$_DFFE_PP_  (.CLK(clknet_leaf_97_clk),
    .RESET_B(net1491),
    .D(_00646_),
    .Q_N(_14677_),
    .Q(\cpu.dcache.r_tag[3][8] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[3][4]$_DFFE_PP_  (.CLK(clknet_leaf_97_clk),
    .RESET_B(net1492),
    .D(_00647_),
    .Q_N(_14676_),
    .Q(\cpu.dcache.r_tag[3][9] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[3][5]$_DFFE_PP_  (.CLK(clknet_leaf_109_clk),
    .RESET_B(net1493),
    .D(_00648_),
    .Q_N(_14675_),
    .Q(\cpu.dcache.r_tag[3][10] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[3][6]$_DFFE_PP_  (.CLK(clknet_leaf_109_clk),
    .RESET_B(net1494),
    .D(_00649_),
    .Q_N(_14674_),
    .Q(\cpu.dcache.r_tag[3][11] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[3][7]$_DFFE_PP_  (.CLK(clknet_leaf_86_clk),
    .RESET_B(net1495),
    .D(_00650_),
    .Q_N(_14673_),
    .Q(\cpu.dcache.r_tag[3][12] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[3][8]$_DFFE_PP_  (.CLK(clknet_leaf_82_clk),
    .RESET_B(net1496),
    .D(_00651_),
    .Q_N(_14672_),
    .Q(\cpu.dcache.r_tag[3][13] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[3][9]$_DFFE_PP_  (.CLK(clknet_leaf_49_clk),
    .RESET_B(net1497),
    .D(_00652_),
    .Q_N(_14671_),
    .Q(\cpu.dcache.r_tag[3][14] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[4][0]$_DFFE_PP_  (.CLK(clknet_leaf_95_clk),
    .RESET_B(net1498),
    .D(_00653_),
    .Q_N(_14670_),
    .Q(\cpu.dcache.r_tag[4][5] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[4][10]$_DFFE_PP_  (.CLK(clknet_leaf_49_clk),
    .RESET_B(net1499),
    .D(_00654_),
    .Q_N(_14669_),
    .Q(\cpu.dcache.r_tag[4][15] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[4][11]$_DFFE_PP_  (.CLK(clknet_leaf_89_clk),
    .RESET_B(net1500),
    .D(_00655_),
    .Q_N(_14668_),
    .Q(\cpu.dcache.r_tag[4][16] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[4][12]$_DFFE_PP_  (.CLK(clknet_leaf_89_clk),
    .RESET_B(net1501),
    .D(_00656_),
    .Q_N(_14667_),
    .Q(\cpu.dcache.r_tag[4][17] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[4][13]$_DFFE_PP_  (.CLK(clknet_leaf_91_clk),
    .RESET_B(net1502),
    .D(_00657_),
    .Q_N(_14666_),
    .Q(\cpu.dcache.r_tag[4][18] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[4][14]$_DFFE_PP_  (.CLK(clknet_leaf_93_clk),
    .RESET_B(net1503),
    .D(_00658_),
    .Q_N(_14665_),
    .Q(\cpu.dcache.r_tag[4][19] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[4][15]$_DFFE_PP_  (.CLK(clknet_leaf_90_clk),
    .RESET_B(net1504),
    .D(_00659_),
    .Q_N(_14664_),
    .Q(\cpu.dcache.r_tag[4][20] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[4][16]$_DFFE_PP_  (.CLK(clknet_leaf_87_clk),
    .RESET_B(net1505),
    .D(_00660_),
    .Q_N(_14663_),
    .Q(\cpu.dcache.r_tag[4][21] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[4][17]$_DFFE_PP_  (.CLK(clknet_leaf_81_clk),
    .RESET_B(net1506),
    .D(_00661_),
    .Q_N(_14662_),
    .Q(\cpu.dcache.r_tag[4][22] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[4][18]$_DFFE_PP_  (.CLK(clknet_leaf_94_clk),
    .RESET_B(net1507),
    .D(_00662_),
    .Q_N(_14661_),
    .Q(\cpu.dcache.r_tag[4][23] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[4][1]$_DFFE_PP_  (.CLK(clknet_leaf_109_clk),
    .RESET_B(net1508),
    .D(_00663_),
    .Q_N(_14660_),
    .Q(\cpu.dcache.r_tag[4][6] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[4][2]$_DFFE_PP_  (.CLK(clknet_leaf_106_clk),
    .RESET_B(net1509),
    .D(_00664_),
    .Q_N(_14659_),
    .Q(\cpu.dcache.r_tag[4][7] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[4][3]$_DFFE_PP_  (.CLK(clknet_leaf_102_clk),
    .RESET_B(net1510),
    .D(_00665_),
    .Q_N(_14658_),
    .Q(\cpu.dcache.r_tag[4][8] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[4][4]$_DFFE_PP_  (.CLK(clknet_leaf_106_clk),
    .RESET_B(net1511),
    .D(_00666_),
    .Q_N(_14657_),
    .Q(\cpu.dcache.r_tag[4][9] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[4][5]$_DFFE_PP_  (.CLK(clknet_leaf_109_clk),
    .RESET_B(net1512),
    .D(_00667_),
    .Q_N(_14656_),
    .Q(\cpu.dcache.r_tag[4][10] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[4][6]$_DFFE_PP_  (.CLK(clknet_leaf_49_clk),
    .RESET_B(net1513),
    .D(_00668_),
    .Q_N(_14655_),
    .Q(\cpu.dcache.r_tag[4][11] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[4][7]$_DFFE_PP_  (.CLK(clknet_leaf_87_clk),
    .RESET_B(net1514),
    .D(_00669_),
    .Q_N(_14654_),
    .Q(\cpu.dcache.r_tag[4][12] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[4][8]$_DFFE_PP_  (.CLK(clknet_leaf_81_clk),
    .RESET_B(net1515),
    .D(_00670_),
    .Q_N(_14653_),
    .Q(\cpu.dcache.r_tag[4][13] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[4][9]$_DFFE_PP_  (.CLK(clknet_leaf_50_clk),
    .RESET_B(net1516),
    .D(_00671_),
    .Q_N(_14652_),
    .Q(\cpu.dcache.r_tag[4][14] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[5][0]$_DFFE_PP_  (.CLK(clknet_leaf_94_clk),
    .RESET_B(net1517),
    .D(_00672_),
    .Q_N(_14651_),
    .Q(\cpu.dcache.r_tag[5][5] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[5][10]$_DFFE_PP_  (.CLK(clknet_leaf_44_clk),
    .RESET_B(net1518),
    .D(_00673_),
    .Q_N(_14650_),
    .Q(\cpu.dcache.r_tag[5][15] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[5][11]$_DFFE_PP_  (.CLK(clknet_leaf_94_clk),
    .RESET_B(net1519),
    .D(_00674_),
    .Q_N(_14649_),
    .Q(\cpu.dcache.r_tag[5][16] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[5][12]$_DFFE_PP_  (.CLK(clknet_leaf_90_clk),
    .RESET_B(net1520),
    .D(_00675_),
    .Q_N(_14648_),
    .Q(\cpu.dcache.r_tag[5][17] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[5][13]$_DFFE_PP_  (.CLK(clknet_leaf_92_clk),
    .RESET_B(net1521),
    .D(_00676_),
    .Q_N(_14647_),
    .Q(\cpu.dcache.r_tag[5][18] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[5][14]$_DFFE_PP_  (.CLK(clknet_leaf_88_clk),
    .RESET_B(net1522),
    .D(_00677_),
    .Q_N(_14646_),
    .Q(\cpu.dcache.r_tag[5][19] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[5][15]$_DFFE_PP_  (.CLK(clknet_leaf_93_clk),
    .RESET_B(net1523),
    .D(_00678_),
    .Q_N(_14645_),
    .Q(\cpu.dcache.r_tag[5][20] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[5][16]$_DFFE_PP_  (.CLK(clknet_leaf_107_clk),
    .RESET_B(net1524),
    .D(_00679_),
    .Q_N(_14644_),
    .Q(\cpu.dcache.r_tag[5][21] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[5][17]$_DFFE_PP_  (.CLK(clknet_leaf_81_clk),
    .RESET_B(net1525),
    .D(_00680_),
    .Q_N(_14643_),
    .Q(\cpu.dcache.r_tag[5][22] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[5][18]$_DFFE_PP_  (.CLK(clknet_leaf_93_clk),
    .RESET_B(net1526),
    .D(_00681_),
    .Q_N(_14642_),
    .Q(\cpu.dcache.r_tag[5][23] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[5][1]$_DFFE_PP_  (.CLK(clknet_leaf_48_clk),
    .RESET_B(net1527),
    .D(_00682_),
    .Q_N(_14641_),
    .Q(\cpu.dcache.r_tag[5][6] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[5][2]$_DFFE_PP_  (.CLK(clknet_leaf_97_clk),
    .RESET_B(net1528),
    .D(_00683_),
    .Q_N(_14640_),
    .Q(\cpu.dcache.r_tag[5][7] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[5][3]$_DFFE_PP_  (.CLK(clknet_leaf_94_clk),
    .RESET_B(net1529),
    .D(_00684_),
    .Q_N(_14639_),
    .Q(\cpu.dcache.r_tag[5][8] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[5][4]$_DFFE_PP_  (.CLK(clknet_leaf_89_clk),
    .RESET_B(net1530),
    .D(_00685_),
    .Q_N(_14638_),
    .Q(\cpu.dcache.r_tag[5][9] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[5][5]$_DFFE_PP_  (.CLK(clknet_leaf_109_clk),
    .RESET_B(net1531),
    .D(_00686_),
    .Q_N(_14637_),
    .Q(\cpu.dcache.r_tag[5][10] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[5][6]$_DFFE_PP_  (.CLK(clknet_leaf_44_clk),
    .RESET_B(net1532),
    .D(_00687_),
    .Q_N(_14636_),
    .Q(\cpu.dcache.r_tag[5][11] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[5][7]$_DFFE_PP_  (.CLK(clknet_leaf_85_clk),
    .RESET_B(net1533),
    .D(_00688_),
    .Q_N(_14635_),
    .Q(\cpu.dcache.r_tag[5][12] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[5][8]$_DFFE_PP_  (.CLK(clknet_leaf_87_clk),
    .RESET_B(net1534),
    .D(_00689_),
    .Q_N(_14634_),
    .Q(\cpu.dcache.r_tag[5][13] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[5][9]$_DFFE_PP_  (.CLK(clknet_leaf_47_clk),
    .RESET_B(net1535),
    .D(_00690_),
    .Q_N(_14633_),
    .Q(\cpu.dcache.r_tag[5][14] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[6][0]$_DFFE_PP_  (.CLK(clknet_leaf_95_clk),
    .RESET_B(net1536),
    .D(_00691_),
    .Q_N(_14632_),
    .Q(\cpu.dcache.r_tag[6][5] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[6][10]$_DFFE_PP_  (.CLK(clknet_leaf_108_clk),
    .RESET_B(net1537),
    .D(_00692_),
    .Q_N(_14631_),
    .Q(\cpu.dcache.r_tag[6][15] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[6][11]$_DFFE_PP_  (.CLK(clknet_leaf_93_clk),
    .RESET_B(net1538),
    .D(_00693_),
    .Q_N(_14630_),
    .Q(\cpu.dcache.r_tag[6][16] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[6][12]$_DFFE_PP_  (.CLK(clknet_leaf_90_clk),
    .RESET_B(net1539),
    .D(_00694_),
    .Q_N(_14629_),
    .Q(\cpu.dcache.r_tag[6][17] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[6][13]$_DFFE_PP_  (.CLK(clknet_leaf_92_clk),
    .RESET_B(net1540),
    .D(_00695_),
    .Q_N(_14628_),
    .Q(\cpu.dcache.r_tag[6][18] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[6][14]$_DFFE_PP_  (.CLK(clknet_leaf_93_clk),
    .RESET_B(net1541),
    .D(_00696_),
    .Q_N(_14627_),
    .Q(\cpu.dcache.r_tag[6][19] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[6][15]$_DFFE_PP_  (.CLK(clknet_leaf_91_clk),
    .RESET_B(net1542),
    .D(_00697_),
    .Q_N(_14626_),
    .Q(\cpu.dcache.r_tag[6][20] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[6][16]$_DFFE_PP_  (.CLK(clknet_leaf_49_clk),
    .RESET_B(net1543),
    .D(_00698_),
    .Q_N(_14625_),
    .Q(\cpu.dcache.r_tag[6][21] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[6][17]$_DFFE_PP_  (.CLK(clknet_leaf_92_clk),
    .RESET_B(net1544),
    .D(_00699_),
    .Q_N(_14624_),
    .Q(\cpu.dcache.r_tag[6][22] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[6][18]$_DFFE_PP_  (.CLK(clknet_leaf_95_clk),
    .RESET_B(net1545),
    .D(_00700_),
    .Q_N(_14623_),
    .Q(\cpu.dcache.r_tag[6][23] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[6][1]$_DFFE_PP_  (.CLK(clknet_leaf_49_clk),
    .RESET_B(net1546),
    .D(_00701_),
    .Q_N(_14622_),
    .Q(\cpu.dcache.r_tag[6][6] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[6][2]$_DFFE_PP_  (.CLK(clknet_leaf_105_clk),
    .RESET_B(net1547),
    .D(_00702_),
    .Q_N(_14621_),
    .Q(\cpu.dcache.r_tag[6][7] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[6][3]$_DFFE_PP_  (.CLK(clknet_leaf_96_clk),
    .RESET_B(net1548),
    .D(_00703_),
    .Q_N(_14620_),
    .Q(\cpu.dcache.r_tag[6][8] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[6][4]$_DFFE_PP_  (.CLK(clknet_leaf_95_clk),
    .RESET_B(net1549),
    .D(_00704_),
    .Q_N(_14619_),
    .Q(\cpu.dcache.r_tag[6][9] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[6][5]$_DFFE_PP_  (.CLK(clknet_leaf_48_clk),
    .RESET_B(net1550),
    .D(_00705_),
    .Q_N(_14618_),
    .Q(\cpu.dcache.r_tag[6][10] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[6][6]$_DFFE_PP_  (.CLK(clknet_leaf_48_clk),
    .RESET_B(net1551),
    .D(_00706_),
    .Q_N(_14617_),
    .Q(\cpu.dcache.r_tag[6][11] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[6][7]$_DFFE_PP_  (.CLK(clknet_leaf_87_clk),
    .RESET_B(net1552),
    .D(_00707_),
    .Q_N(_14616_),
    .Q(\cpu.dcache.r_tag[6][12] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[6][8]$_DFFE_PP_  (.CLK(clknet_leaf_81_clk),
    .RESET_B(net1553),
    .D(_00708_),
    .Q_N(_14615_),
    .Q(\cpu.dcache.r_tag[6][13] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[6][9]$_DFFE_PP_  (.CLK(clknet_leaf_49_clk),
    .RESET_B(net1554),
    .D(_00709_),
    .Q_N(_14614_),
    .Q(\cpu.dcache.r_tag[6][14] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[7][0]$_DFFE_PP_  (.CLK(clknet_leaf_95_clk),
    .RESET_B(net1555),
    .D(_00710_),
    .Q_N(_14613_),
    .Q(\cpu.dcache.r_tag[7][5] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[7][10]$_DFFE_PP_  (.CLK(clknet_leaf_48_clk),
    .RESET_B(net1556),
    .D(_00711_),
    .Q_N(_14612_),
    .Q(\cpu.dcache.r_tag[7][15] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[7][11]$_DFFE_PP_  (.CLK(clknet_leaf_94_clk),
    .RESET_B(net1557),
    .D(_00712_),
    .Q_N(_14611_),
    .Q(\cpu.dcache.r_tag[7][16] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[7][12]$_DFFE_PP_  (.CLK(clknet_leaf_95_clk),
    .RESET_B(net1558),
    .D(_00713_),
    .Q_N(_14610_),
    .Q(\cpu.dcache.r_tag[7][17] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[7][13]$_DFFE_PP_  (.CLK(clknet_leaf_93_clk),
    .RESET_B(net1559),
    .D(_00714_),
    .Q_N(_14609_),
    .Q(\cpu.dcache.r_tag[7][18] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[7][14]$_DFFE_PP_  (.CLK(clknet_leaf_90_clk),
    .RESET_B(net1560),
    .D(_00715_),
    .Q_N(_14608_),
    .Q(\cpu.dcache.r_tag[7][19] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[7][15]$_DFFE_PP_  (.CLK(clknet_leaf_88_clk),
    .RESET_B(net1561),
    .D(_00716_),
    .Q_N(_14607_),
    .Q(\cpu.dcache.r_tag[7][20] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[7][16]$_DFFE_PP_  (.CLK(clknet_leaf_47_clk),
    .RESET_B(net1562),
    .D(_00717_),
    .Q_N(_14606_),
    .Q(\cpu.dcache.r_tag[7][21] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[7][17]$_DFFE_PP_  (.CLK(clknet_leaf_92_clk),
    .RESET_B(net1563),
    .D(_00718_),
    .Q_N(_14605_),
    .Q(\cpu.dcache.r_tag[7][22] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[7][18]$_DFFE_PP_  (.CLK(clknet_leaf_93_clk),
    .RESET_B(net1564),
    .D(_00719_),
    .Q_N(_14604_),
    .Q(\cpu.dcache.r_tag[7][23] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[7][1]$_DFFE_PP_  (.CLK(clknet_leaf_96_clk),
    .RESET_B(net1565),
    .D(_00720_),
    .Q_N(_14603_),
    .Q(\cpu.dcache.r_tag[7][6] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[7][2]$_DFFE_PP_  (.CLK(clknet_leaf_105_clk),
    .RESET_B(net1566),
    .D(_00721_),
    .Q_N(_14602_),
    .Q(\cpu.dcache.r_tag[7][7] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[7][3]$_DFFE_PP_  (.CLK(clknet_leaf_96_clk),
    .RESET_B(net1567),
    .D(_00722_),
    .Q_N(_14601_),
    .Q(\cpu.dcache.r_tag[7][8] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[7][4]$_DFFE_PP_  (.CLK(clknet_leaf_96_clk),
    .RESET_B(net1568),
    .D(_00723_),
    .Q_N(_14600_),
    .Q(\cpu.dcache.r_tag[7][9] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[7][5]$_DFFE_PP_  (.CLK(clknet_leaf_110_clk),
    .RESET_B(net1569),
    .D(_00724_),
    .Q_N(_14599_),
    .Q(\cpu.dcache.r_tag[7][10] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[7][6]$_DFFE_PP_  (.CLK(clknet_leaf_111_clk),
    .RESET_B(net1570),
    .D(_00725_),
    .Q_N(_14598_),
    .Q(\cpu.dcache.r_tag[7][11] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[7][7]$_DFFE_PP_  (.CLK(clknet_leaf_86_clk),
    .RESET_B(net1571),
    .D(_00726_),
    .Q_N(_14597_),
    .Q(\cpu.dcache.r_tag[7][12] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[7][8]$_DFFE_PP_  (.CLK(clknet_leaf_91_clk),
    .RESET_B(net1572),
    .D(_00727_),
    .Q_N(_14596_),
    .Q(\cpu.dcache.r_tag[7][13] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[7][9]$_DFFE_PP_  (.CLK(clknet_leaf_47_clk),
    .RESET_B(net1573),
    .D(_00728_),
    .Q_N(_14595_),
    .Q(\cpu.dcache.r_tag[7][14] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_valid[0]$_SDFFE_PP0P_  (.CLK(clknet_leaf_50_clk),
    .RESET_B(net1574),
    .D(_00729_),
    .Q_N(_14594_),
    .Q(\cpu.dcache.r_valid[0] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_valid[1]$_SDFFE_PP0P_  (.CLK(clknet_leaf_51_clk),
    .RESET_B(net1575),
    .D(_00730_),
    .Q_N(_14593_),
    .Q(\cpu.dcache.r_valid[1] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_valid[2]$_SDFFE_PP0P_  (.CLK(clknet_leaf_50_clk),
    .RESET_B(net1576),
    .D(_00731_),
    .Q_N(_14592_),
    .Q(\cpu.dcache.r_valid[2] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_valid[3]$_SDFFE_PP0P_  (.CLK(clknet_leaf_50_clk),
    .RESET_B(net1577),
    .D(_00732_),
    .Q_N(_14591_),
    .Q(\cpu.dcache.r_valid[3] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_valid[4]$_SDFFE_PP0P_  (.CLK(clknet_leaf_50_clk),
    .RESET_B(net1578),
    .D(_00733_),
    .Q_N(_14590_),
    .Q(\cpu.dcache.r_valid[4] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_valid[5]$_SDFFE_PP0P_  (.CLK(clknet_leaf_51_clk),
    .RESET_B(net1579),
    .D(_00734_),
    .Q_N(_14589_),
    .Q(\cpu.dcache.r_valid[5] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_valid[6]$_SDFFE_PP0P_  (.CLK(clknet_leaf_51_clk),
    .RESET_B(net1580),
    .D(_00735_),
    .Q_N(_14588_),
    .Q(\cpu.dcache.r_valid[6] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_valid[7]$_SDFFE_PP0P_  (.CLK(clknet_leaf_51_clk),
    .RESET_B(net1581),
    .D(_00736_),
    .Q_N(_14587_),
    .Q(\cpu.dcache.r_valid[7] ));
 sg13g2_dfrbp_1 \cpu.dec.r_br$_DFFE_PP_  (.CLK(clknet_leaf_175_clk),
    .RESET_B(net1582),
    .D(_00737_),
    .Q_N(_14586_),
    .Q(\cpu.br ));
 sg13g2_dfrbp_1 \cpu.dec.r_cond[0]$_DFFE_PP_  (.CLK(clknet_leaf_176_clk),
    .RESET_B(net1583),
    .D(_00738_),
    .Q_N(_00282_),
    .Q(\cpu.cond[0] ));
 sg13g2_dfrbp_1 \cpu.dec.r_cond[1]$_DFFE_PP_  (.CLK(clknet_leaf_180_clk),
    .RESET_B(net1584),
    .D(_00739_),
    .Q_N(_14585_),
    .Q(\cpu.cond[1] ));
 sg13g2_dfrbp_1 \cpu.dec.r_cond[2]$_DFFE_PP_  (.CLK(clknet_leaf_179_clk),
    .RESET_B(net1585),
    .D(_00740_),
    .Q_N(_00257_),
    .Q(\cpu.cond[2] ));
 sg13g2_dfrbp_1 \cpu.dec.r_div$_DFFE_PP_  (.CLK(clknet_leaf_174_clk),
    .RESET_B(net1586),
    .D(_00741_),
    .Q_N(_14584_),
    .Q(\cpu.dec.div ));
 sg13g2_dfrbp_1 \cpu.dec.r_flush_all$_DFFE_PP_  (.CLK(clknet_leaf_179_clk),
    .RESET_B(net1587),
    .D(_00742_),
    .Q_N(_14583_),
    .Q(\cpu.dec.do_flush_all ));
 sg13g2_dfrbp_1 \cpu.dec.r_flush_write$_DFFE_PP_  (.CLK(clknet_leaf_179_clk),
    .RESET_B(net1588),
    .D(_00743_),
    .Q_N(_14582_),
    .Q(\cpu.dec.do_flush_write ));
 sg13g2_dfrbp_1 \cpu.dec.r_imm[0]$_DFFE_PP_  (.CLK(clknet_leaf_255_clk),
    .RESET_B(net1589),
    .D(_00744_),
    .Q_N(_14581_),
    .Q(\cpu.dec.imm[0] ));
 sg13g2_dfrbp_1 \cpu.dec.r_imm[10]$_DFFE_PP_  (.CLK(clknet_leaf_181_clk),
    .RESET_B(net1590),
    .D(_00745_),
    .Q_N(_14580_),
    .Q(\cpu.dec.imm[10] ));
 sg13g2_dfrbp_1 \cpu.dec.r_imm[11]$_DFFE_PP_  (.CLK(clknet_leaf_174_clk),
    .RESET_B(net1591),
    .D(_00746_),
    .Q_N(_14579_),
    .Q(\cpu.dec.imm[11] ));
 sg13g2_dfrbp_1 \cpu.dec.r_imm[12]$_DFFE_PP_  (.CLK(clknet_leaf_174_clk),
    .RESET_B(net1592),
    .D(_00747_),
    .Q_N(_14578_),
    .Q(\cpu.dec.imm[12] ));
 sg13g2_dfrbp_1 \cpu.dec.r_imm[13]$_DFFE_PP_  (.CLK(clknet_leaf_174_clk),
    .RESET_B(net1593),
    .D(_00748_),
    .Q_N(_14577_),
    .Q(\cpu.dec.imm[13] ));
 sg13g2_dfrbp_1 \cpu.dec.r_imm[14]$_DFFE_PP_  (.CLK(clknet_leaf_175_clk),
    .RESET_B(net1594),
    .D(_00749_),
    .Q_N(_14576_),
    .Q(\cpu.dec.imm[14] ));
 sg13g2_dfrbp_1 \cpu.dec.r_imm[15]$_DFFE_PP_  (.CLK(clknet_leaf_175_clk),
    .RESET_B(net1595),
    .D(_00750_),
    .Q_N(_14575_),
    .Q(\cpu.dec.imm[15] ));
 sg13g2_dfrbp_1 \cpu.dec.r_imm[1]$_DFFE_PP_  (.CLK(clknet_leaf_260_clk),
    .RESET_B(net1596),
    .D(_00751_),
    .Q_N(_14574_),
    .Q(\cpu.dec.imm[1] ));
 sg13g2_dfrbp_1 \cpu.dec.r_imm[2]$_DFFE_PP_  (.CLK(clknet_leaf_180_clk),
    .RESET_B(net1597),
    .D(_00752_),
    .Q_N(_14573_),
    .Q(\cpu.dec.imm[2] ));
 sg13g2_dfrbp_1 \cpu.dec.r_imm[3]$_DFFE_PP_  (.CLK(clknet_leaf_255_clk),
    .RESET_B(net1598),
    .D(_00753_),
    .Q_N(_14572_),
    .Q(\cpu.dec.imm[3] ));
 sg13g2_dfrbp_1 \cpu.dec.r_imm[4]$_DFFE_PP_  (.CLK(clknet_leaf_179_clk),
    .RESET_B(net1599),
    .D(_00754_),
    .Q_N(_14571_),
    .Q(\cpu.dec.imm[4] ));
 sg13g2_dfrbp_1 \cpu.dec.r_imm[5]$_DFFE_PP_  (.CLK(clknet_leaf_180_clk),
    .RESET_B(net1600),
    .D(_00755_),
    .Q_N(_14570_),
    .Q(\cpu.dec.imm[5] ));
 sg13g2_dfrbp_1 \cpu.dec.r_imm[6]$_DFFE_PP_  (.CLK(clknet_leaf_255_clk),
    .RESET_B(net1601),
    .D(_00756_),
    .Q_N(_14569_),
    .Q(\cpu.dec.imm[6] ));
 sg13g2_dfrbp_1 \cpu.dec.r_imm[7]$_DFFE_PP_  (.CLK(clknet_leaf_178_clk),
    .RESET_B(net1602),
    .D(_00757_),
    .Q_N(_14568_),
    .Q(\cpu.dec.imm[7] ));
 sg13g2_dfrbp_1 \cpu.dec.r_imm[8]$_DFFE_PP_  (.CLK(clknet_leaf_174_clk),
    .RESET_B(net1603),
    .D(_00758_),
    .Q_N(_14567_),
    .Q(\cpu.dec.imm[8] ));
 sg13g2_dfrbp_1 \cpu.dec.r_imm[9]$_DFFE_PP_  (.CLK(clknet_leaf_174_clk),
    .RESET_B(net1604),
    .D(_00759_),
    .Q_N(_14566_),
    .Q(\cpu.dec.imm[9] ));
 sg13g2_dfrbp_1 \cpu.dec.r_inv_mmu$_DFFE_PP_  (.CLK(clknet_leaf_260_clk),
    .RESET_B(net1605),
    .D(_00760_),
    .Q_N(_14565_),
    .Q(\cpu.dec.do_inv_mmu ));
 sg13g2_dfrbp_1 \cpu.dec.r_io$_DFFE_PP_  (.CLK(clknet_leaf_180_clk),
    .RESET_B(net1606),
    .D(_00761_),
    .Q_N(_14564_),
    .Q(\cpu.dec.io ));
 sg13g2_dfrbp_1 \cpu.dec.r_jmp$_SDFFCE_PP0P_  (.CLK(clknet_leaf_179_clk),
    .RESET_B(net1607),
    .D(_00762_),
    .Q_N(_00242_),
    .Q(\cpu.dec.jmp ));
 sg13g2_dfrbp_1 \cpu.dec.r_load$_DFFE_PP_  (.CLK(clknet_leaf_260_clk),
    .RESET_B(net1608),
    .D(_00763_),
    .Q_N(_14563_),
    .Q(\cpu.dec.load ));
 sg13g2_dfrbp_1 \cpu.dec.r_mult$_DFFE_PP_  (.CLK(clknet_leaf_179_clk),
    .RESET_B(net1609),
    .D(_00764_),
    .Q_N(_14562_),
    .Q(\cpu.dec.mult ));
 sg13g2_dfrbp_1 \cpu.dec.r_needs_rs2$_DFFE_PP_  (.CLK(clknet_leaf_175_clk),
    .RESET_B(net1610),
    .D(_00765_),
    .Q_N(_14974_),
    .Q(\cpu.dec.needs_rs2 ));
 sg13g2_dfrbp_1 \cpu.dec.r_op[10]$_DFF_P_  (.CLK(clknet_leaf_182_clk),
    .RESET_B(net1611),
    .D(_00011_),
    .Q_N(_14975_),
    .Q(\cpu.dec.r_op[10] ));
 sg13g2_dfrbp_1 \cpu.dec.r_op[1]$_DFF_P_  (.CLK(clknet_leaf_181_clk),
    .RESET_B(net1612),
    .D(_00012_),
    .Q_N(_14976_),
    .Q(\cpu.dec.r_op[1] ));
 sg13g2_dfrbp_1 \cpu.dec.r_op[2]$_DFF_P_  (.CLK(clknet_leaf_181_clk),
    .RESET_B(net1613),
    .D(_00013_),
    .Q_N(_14977_),
    .Q(\cpu.dec.r_op[2] ));
 sg13g2_dfrbp_1 \cpu.dec.r_op[3]$_DFF_P_  (.CLK(clknet_leaf_174_clk),
    .RESET_B(net1614),
    .D(_00014_),
    .Q_N(_14978_),
    .Q(\cpu.dec.r_op[3] ));
 sg13g2_dfrbp_1 \cpu.dec.r_op[4]$_DFF_P_  (.CLK(clknet_leaf_181_clk),
    .RESET_B(net1615),
    .D(_00015_),
    .Q_N(_14979_),
    .Q(\cpu.dec.r_op[4] ));
 sg13g2_dfrbp_1 \cpu.dec.r_op[5]$_DFF_P_  (.CLK(clknet_leaf_182_clk),
    .RESET_B(net1616),
    .D(_00016_),
    .Q_N(_14980_),
    .Q(\cpu.dec.r_op[5] ));
 sg13g2_dfrbp_1 \cpu.dec.r_op[6]$_DFF_P_  (.CLK(clknet_leaf_181_clk),
    .RESET_B(net1617),
    .D(_00017_),
    .Q_N(_14981_),
    .Q(\cpu.dec.r_op[6] ));
 sg13g2_dfrbp_1 \cpu.dec.r_op[7]$_DFF_P_  (.CLK(clknet_leaf_182_clk),
    .RESET_B(net1618),
    .D(_00018_),
    .Q_N(_14982_),
    .Q(\cpu.dec.r_op[7] ));
 sg13g2_dfrbp_1 \cpu.dec.r_op[8]$_DFF_P_  (.CLK(clknet_leaf_181_clk),
    .RESET_B(net1619),
    .D(_00019_),
    .Q_N(_14983_),
    .Q(\cpu.dec.r_op[8] ));
 sg13g2_dfrbp_1 \cpu.dec.r_op[9]$_DFF_P_  (.CLK(clknet_leaf_181_clk),
    .RESET_B(net1620),
    .D(_00020_),
    .Q_N(_14561_),
    .Q(\cpu.dec.r_op[9] ));
 sg13g2_dfrbp_1 \cpu.dec.r_rd[0]$_DFFE_PP_  (.CLK(clknet_leaf_180_clk),
    .RESET_B(net1621),
    .D(_00766_),
    .Q_N(_14560_),
    .Q(\cpu.dec.r_rd[0] ));
 sg13g2_dfrbp_1 \cpu.dec.r_rd[1]$_DFFE_PP_  (.CLK(clknet_leaf_179_clk),
    .RESET_B(net1622),
    .D(_00767_),
    .Q_N(_14559_),
    .Q(\cpu.dec.r_rd[1] ));
 sg13g2_dfrbp_1 \cpu.dec.r_rd[2]$_DFFE_PP_  (.CLK(clknet_leaf_178_clk),
    .RESET_B(net1623),
    .D(_00768_),
    .Q_N(_14558_),
    .Q(\cpu.dec.r_rd[2] ));
 sg13g2_dfrbp_1 \cpu.dec.r_rd[3]$_DFFE_PP_  (.CLK(clknet_leaf_255_clk),
    .RESET_B(net1624),
    .D(_00769_),
    .Q_N(_14984_),
    .Q(\cpu.dec.r_rd[3] ));
 sg13g2_dfrbp_1 \cpu.dec.r_ready$_DFF_P_  (.CLK(clknet_leaf_177_clk),
    .RESET_B(net1625),
    .D(_00052_),
    .Q_N(_14557_),
    .Q(\cpu.dec.iready ));
 sg13g2_dfrbp_1 \cpu.dec.r_rs1[0]$_DFFE_PP_  (.CLK(clknet_leaf_177_clk),
    .RESET_B(net1626),
    .D(_00770_),
    .Q_N(_14556_),
    .Q(\cpu.dec.r_rs1[0] ));
 sg13g2_dfrbp_1 \cpu.dec.r_rs1[1]$_DFFE_PP_  (.CLK(clknet_leaf_178_clk),
    .RESET_B(net1627),
    .D(_00771_),
    .Q_N(_14555_),
    .Q(\cpu.dec.r_rs1[1] ));
 sg13g2_dfrbp_1 \cpu.dec.r_rs1[2]$_DFFE_PP_  (.CLK(clknet_leaf_177_clk),
    .RESET_B(net1628),
    .D(_00772_),
    .Q_N(_14554_),
    .Q(\cpu.dec.r_rs1[2] ));
 sg13g2_dfrbp_1 \cpu.dec.r_rs1[3]$_DFFE_PP_  (.CLK(clknet_leaf_178_clk),
    .RESET_B(net1629),
    .D(_00773_),
    .Q_N(_14553_),
    .Q(\cpu.dec.r_rs1[3] ));
 sg13g2_dfrbp_1 \cpu.dec.r_rs2[0]$_DFFE_PP_  (.CLK(clknet_leaf_177_clk),
    .RESET_B(net1630),
    .D(_00774_),
    .Q_N(_14552_),
    .Q(\cpu.dec.r_rs2[0] ));
 sg13g2_dfrbp_1 \cpu.dec.r_rs2[1]$_DFFE_PP_  (.CLK(clknet_leaf_116_clk),
    .RESET_B(net1631),
    .D(_00775_),
    .Q_N(_14551_),
    .Q(\cpu.dec.r_rs2[1] ));
 sg13g2_dfrbp_1 \cpu.dec.r_rs2[2]$_DFFE_PP_  (.CLK(clknet_leaf_177_clk),
    .RESET_B(net1632),
    .D(_00776_),
    .Q_N(_14550_),
    .Q(\cpu.dec.r_rs2[2] ));
 sg13g2_dfrbp_1 \cpu.dec.r_rs2[3]$_DFFE_PP_  (.CLK(clknet_leaf_262_clk),
    .RESET_B(net1633),
    .D(_00777_),
    .Q_N(_14549_),
    .Q(\cpu.dec.r_rs2[3] ));
 sg13g2_dfrbp_1 \cpu.dec.r_rs2_pc$_DFFE_PP_  (.CLK(clknet_leaf_175_clk),
    .RESET_B(net1634),
    .D(_00778_),
    .Q_N(_14548_),
    .Q(\cpu.dec.r_rs2_pc ));
 sg13g2_dfrbp_1 \cpu.dec.r_set_cc$_SDFFCE_PP0P_  (.CLK(clknet_leaf_179_clk),
    .RESET_B(net1635),
    .D(_00779_),
    .Q_N(_14547_),
    .Q(\cpu.dec.r_set_cc ));
 sg13g2_dfrbp_1 \cpu.dec.r_store$_DFFE_PP_  (.CLK(clknet_leaf_178_clk),
    .RESET_B(net1636),
    .D(_00780_),
    .Q_N(_00294_),
    .Q(\cpu.dec.r_store ));
 sg13g2_dfrbp_1 \cpu.dec.r_swapsp$_DFFE_PP_  (.CLK(clknet_leaf_180_clk),
    .RESET_B(net1637),
    .D(_00781_),
    .Q_N(_14546_),
    .Q(\cpu.dec.r_swapsp ));
 sg13g2_dfrbp_1 \cpu.dec.r_sys_call$_DFFE_PP_  (.CLK(clknet_leaf_174_clk),
    .RESET_B(net1638),
    .D(_00782_),
    .Q_N(_00258_),
    .Q(\cpu.dec.r_sys_call ));
 sg13g2_dfrbp_1 \cpu.dec.r_trap$_DFFE_PP_  (.CLK(clknet_leaf_180_clk),
    .RESET_B(net1639),
    .D(_00783_),
    .Q_N(_14545_),
    .Q(\cpu.dec.r_trap ));
 sg13g2_dfrbp_1 \cpu.ex.genblk3.r_mmu_d_proxy$_SDFFE_PP0P_  (.CLK(clknet_leaf_178_clk),
    .RESET_B(net1640),
    .D(_00784_),
    .Q_N(_14544_),
    .Q(\cpu.ex.genblk3.r_mmu_d_proxy ));
 sg13g2_dfrbp_1 \cpu.ex.genblk3.r_mmu_enable$_SDFFE_PN0P_  (.CLK(clknet_leaf_182_clk),
    .RESET_B(net1641),
    .D(_00785_),
    .Q_N(_00182_),
    .Q(\cpu.ex.genblk3.r_mmu_enable ));
 sg13g2_dfrbp_1 \cpu.ex.genblk3.r_prev_supmode$_SDFFE_PN1P_  (.CLK(clknet_leaf_116_clk),
    .RESET_B(net1642),
    .D(_00786_),
    .Q_N(_14985_),
    .Q(\cpu.ex.genblk3.r_prev_supmode ));
 sg13g2_dfrbp_1 \cpu.ex.genblk3.r_supmode$_DFF_P_  (.CLK(clknet_leaf_178_clk),
    .RESET_B(net1643),
    .D(\cpu.ex.genblk3.c_supmode ),
    .Q_N(_00183_),
    .Q(\cpu.dec.supmode ));
 sg13g2_dfrbp_1 \cpu.ex.genblk3.r_user_io$_SDFFE_PN0P_  (.CLK(clknet_leaf_43_clk),
    .RESET_B(net1644),
    .D(_00787_),
    .Q_N(_14543_),
    .Q(\cpu.dec.user_io ));
 sg13g2_dfrbp_1 \cpu.ex.r_10[0]$_DFFE_PP_  (.CLK(clknet_leaf_122_clk),
    .RESET_B(net1645),
    .D(_00788_),
    .Q_N(_14542_),
    .Q(\cpu.ex.r_10[0] ));
 sg13g2_dfrbp_1 \cpu.ex.r_10[10]$_DFFE_PP_  (.CLK(clknet_leaf_112_clk),
    .RESET_B(net1646),
    .D(_00789_),
    .Q_N(_14541_),
    .Q(\cpu.ex.r_10[10] ));
 sg13g2_dfrbp_1 \cpu.ex.r_10[11]$_DFFE_PP_  (.CLK(clknet_leaf_105_clk),
    .RESET_B(net1647),
    .D(_00790_),
    .Q_N(_14540_),
    .Q(\cpu.ex.r_10[11] ));
 sg13g2_dfrbp_1 \cpu.ex.r_10[12]$_DFFE_PP_  (.CLK(clknet_leaf_42_clk),
    .RESET_B(net1648),
    .D(_00791_),
    .Q_N(_14539_),
    .Q(\cpu.ex.r_10[12] ));
 sg13g2_dfrbp_1 \cpu.ex.r_10[13]$_DFFE_PP_  (.CLK(clknet_leaf_263_clk),
    .RESET_B(net1649),
    .D(_00792_),
    .Q_N(_14538_),
    .Q(\cpu.ex.r_10[13] ));
 sg13g2_dfrbp_1 \cpu.ex.r_10[14]$_DFFE_PP_  (.CLK(clknet_leaf_110_clk),
    .RESET_B(net1650),
    .D(_00793_),
    .Q_N(_14537_),
    .Q(\cpu.ex.r_10[14] ));
 sg13g2_dfrbp_1 \cpu.ex.r_10[15]$_DFFE_PP_  (.CLK(clknet_leaf_40_clk),
    .RESET_B(net1651),
    .D(_00794_),
    .Q_N(_14536_),
    .Q(\cpu.ex.r_10[15] ));
 sg13g2_dfrbp_1 \cpu.ex.r_10[1]$_DFFE_PP_  (.CLK(clknet_leaf_113_clk),
    .RESET_B(net1652),
    .D(_00795_),
    .Q_N(_14535_),
    .Q(\cpu.ex.r_10[1] ));
 sg13g2_dfrbp_1 \cpu.ex.r_10[2]$_DFFE_PP_  (.CLK(clknet_leaf_262_clk),
    .RESET_B(net1653),
    .D(_00796_),
    .Q_N(_14534_),
    .Q(\cpu.ex.r_10[2] ));
 sg13g2_dfrbp_1 \cpu.ex.r_10[3]$_DFFE_PP_  (.CLK(clknet_leaf_104_clk),
    .RESET_B(net1654),
    .D(_00797_),
    .Q_N(_14533_),
    .Q(\cpu.ex.r_10[3] ));
 sg13g2_dfrbp_1 \cpu.ex.r_10[4]$_DFFE_PP_  (.CLK(clknet_leaf_103_clk),
    .RESET_B(net1655),
    .D(_00798_),
    .Q_N(_14532_),
    .Q(\cpu.ex.r_10[4] ));
 sg13g2_dfrbp_1 \cpu.ex.r_10[5]$_DFFE_PP_  (.CLK(clknet_leaf_97_clk),
    .RESET_B(net1656),
    .D(_00799_),
    .Q_N(_14531_),
    .Q(\cpu.ex.r_10[5] ));
 sg13g2_dfrbp_1 \cpu.ex.r_10[6]$_DFFE_PP_  (.CLK(clknet_leaf_124_clk),
    .RESET_B(net1657),
    .D(_00800_),
    .Q_N(_14530_),
    .Q(\cpu.ex.r_10[6] ));
 sg13g2_dfrbp_1 \cpu.ex.r_10[7]$_DFFE_PP_  (.CLK(clknet_leaf_96_clk),
    .RESET_B(net1658),
    .D(_00801_),
    .Q_N(_14529_),
    .Q(\cpu.ex.r_10[7] ));
 sg13g2_dfrbp_1 \cpu.ex.r_10[8]$_DFFE_PP_  (.CLK(clknet_leaf_97_clk),
    .RESET_B(net1659),
    .D(_00802_),
    .Q_N(_14528_),
    .Q(\cpu.ex.r_10[8] ));
 sg13g2_dfrbp_1 \cpu.ex.r_10[9]$_DFFE_PP_  (.CLK(clknet_leaf_101_clk),
    .RESET_B(net1660),
    .D(_00803_),
    .Q_N(_14527_),
    .Q(\cpu.ex.r_10[9] ));
 sg13g2_dfrbp_1 \cpu.ex.r_11[0]$_DFFE_PP_  (.CLK(clknet_leaf_123_clk),
    .RESET_B(net1661),
    .D(_00804_),
    .Q_N(_14526_),
    .Q(\cpu.ex.r_11[0] ));
 sg13g2_dfrbp_1 \cpu.ex.r_11[10]$_DFFE_PP_  (.CLK(clknet_leaf_110_clk),
    .RESET_B(net1662),
    .D(_00805_),
    .Q_N(_14525_),
    .Q(\cpu.ex.r_11[10] ));
 sg13g2_dfrbp_1 \cpu.ex.r_11[11]$_DFFE_PP_  (.CLK(clknet_leaf_104_clk),
    .RESET_B(net1663),
    .D(_00806_),
    .Q_N(_14524_),
    .Q(\cpu.ex.r_11[11] ));
 sg13g2_dfrbp_1 \cpu.ex.r_11[12]$_DFFE_PP_  (.CLK(clknet_leaf_115_clk),
    .RESET_B(net1664),
    .D(_00807_),
    .Q_N(_14523_),
    .Q(\cpu.ex.r_11[12] ));
 sg13g2_dfrbp_1 \cpu.ex.r_11[13]$_DFFE_PP_  (.CLK(clknet_leaf_263_clk),
    .RESET_B(net1665),
    .D(_00808_),
    .Q_N(_14522_),
    .Q(\cpu.ex.r_11[13] ));
 sg13g2_dfrbp_1 \cpu.ex.r_11[14]$_DFFE_PP_  (.CLK(clknet_leaf_113_clk),
    .RESET_B(net1666),
    .D(_00809_),
    .Q_N(_14521_),
    .Q(\cpu.ex.r_11[14] ));
 sg13g2_dfrbp_1 \cpu.ex.r_11[15]$_DFFE_PP_  (.CLK(clknet_leaf_40_clk),
    .RESET_B(net1667),
    .D(_00810_),
    .Q_N(_14520_),
    .Q(\cpu.ex.r_11[15] ));
 sg13g2_dfrbp_1 \cpu.ex.r_11[1]$_DFFE_PP_  (.CLK(clknet_leaf_114_clk),
    .RESET_B(net1668),
    .D(_00811_),
    .Q_N(_14519_),
    .Q(\cpu.ex.r_11[1] ));
 sg13g2_dfrbp_1 \cpu.ex.r_11[2]$_DFFE_PP_  (.CLK(clknet_leaf_262_clk),
    .RESET_B(net1669),
    .D(_00812_),
    .Q_N(_14518_),
    .Q(\cpu.ex.r_11[2] ));
 sg13g2_dfrbp_1 \cpu.ex.r_11[3]$_DFFE_PP_  (.CLK(clknet_leaf_104_clk),
    .RESET_B(net1670),
    .D(_00813_),
    .Q_N(_14517_),
    .Q(\cpu.ex.r_11[3] ));
 sg13g2_dfrbp_1 \cpu.ex.r_11[4]$_DFFE_PP_  (.CLK(clknet_leaf_99_clk),
    .RESET_B(net1671),
    .D(_00814_),
    .Q_N(_14516_),
    .Q(\cpu.ex.r_11[4] ));
 sg13g2_dfrbp_1 \cpu.ex.r_11[5]$_DFFE_PP_  (.CLK(clknet_leaf_99_clk),
    .RESET_B(net1672),
    .D(_00815_),
    .Q_N(_14515_),
    .Q(\cpu.ex.r_11[5] ));
 sg13g2_dfrbp_1 \cpu.ex.r_11[6]$_DFFE_PP_  (.CLK(clknet_leaf_99_clk),
    .RESET_B(net1673),
    .D(_00816_),
    .Q_N(_14514_),
    .Q(\cpu.ex.r_11[6] ));
 sg13g2_dfrbp_1 \cpu.ex.r_11[7]$_DFFE_PP_  (.CLK(clknet_leaf_97_clk),
    .RESET_B(net1674),
    .D(_00817_),
    .Q_N(_14513_),
    .Q(\cpu.ex.r_11[7] ));
 sg13g2_dfrbp_1 \cpu.ex.r_11[8]$_DFFE_PP_  (.CLK(clknet_leaf_97_clk),
    .RESET_B(net1675),
    .D(_00818_),
    .Q_N(_14512_),
    .Q(\cpu.ex.r_11[8] ));
 sg13g2_dfrbp_1 \cpu.ex.r_11[9]$_DFFE_PP_  (.CLK(clknet_leaf_124_clk),
    .RESET_B(net1676),
    .D(_00819_),
    .Q_N(_14511_),
    .Q(\cpu.ex.r_11[9] ));
 sg13g2_dfrbp_1 \cpu.ex.r_12[0]$_DFFE_PP_  (.CLK(clknet_leaf_122_clk),
    .RESET_B(net1677),
    .D(_00820_),
    .Q_N(_14510_),
    .Q(\cpu.ex.r_12[0] ));
 sg13g2_dfrbp_1 \cpu.ex.r_12[10]$_DFFE_PP_  (.CLK(clknet_leaf_111_clk),
    .RESET_B(net1678),
    .D(_00821_),
    .Q_N(_14509_),
    .Q(\cpu.ex.r_12[10] ));
 sg13g2_dfrbp_1 \cpu.ex.r_12[11]$_DFFE_PP_  (.CLK(clknet_leaf_111_clk),
    .RESET_B(net1679),
    .D(_00822_),
    .Q_N(_14508_),
    .Q(\cpu.ex.r_12[11] ));
 sg13g2_dfrbp_1 \cpu.ex.r_12[12]$_DFFE_PP_  (.CLK(clknet_leaf_41_clk),
    .RESET_B(net1680),
    .D(_00823_),
    .Q_N(_14507_),
    .Q(\cpu.ex.r_12[12] ));
 sg13g2_dfrbp_1 \cpu.ex.r_12[13]$_DFFE_PP_  (.CLK(clknet_leaf_41_clk),
    .RESET_B(net1681),
    .D(_00824_),
    .Q_N(_14506_),
    .Q(\cpu.ex.r_12[13] ));
 sg13g2_dfrbp_1 \cpu.ex.r_12[14]$_DFFE_PP_  (.CLK(clknet_leaf_110_clk),
    .RESET_B(net1682),
    .D(_00825_),
    .Q_N(_14505_),
    .Q(\cpu.ex.r_12[14] ));
 sg13g2_dfrbp_1 \cpu.ex.r_12[15]$_DFFE_PP_  (.CLK(clknet_leaf_41_clk),
    .RESET_B(net1683),
    .D(_00826_),
    .Q_N(_14504_),
    .Q(\cpu.ex.r_12[15] ));
 sg13g2_dfrbp_1 \cpu.ex.r_12[1]$_DFFE_PP_  (.CLK(clknet_leaf_44_clk),
    .RESET_B(net1684),
    .D(_00827_),
    .Q_N(_14503_),
    .Q(\cpu.ex.r_12[1] ));
 sg13g2_dfrbp_1 \cpu.ex.r_12[2]$_DFFE_PP_  (.CLK(clknet_leaf_177_clk),
    .RESET_B(net1685),
    .D(_00828_),
    .Q_N(_14502_),
    .Q(\cpu.ex.r_12[2] ));
 sg13g2_dfrbp_1 \cpu.ex.r_12[3]$_DFFE_PP_  (.CLK(clknet_leaf_105_clk),
    .RESET_B(net1686),
    .D(_00829_),
    .Q_N(_14501_),
    .Q(\cpu.ex.r_12[3] ));
 sg13g2_dfrbp_1 \cpu.ex.r_12[4]$_DFFE_PP_  (.CLK(clknet_leaf_126_clk),
    .RESET_B(net1687),
    .D(_00830_),
    .Q_N(_14500_),
    .Q(\cpu.ex.r_12[4] ));
 sg13g2_dfrbp_1 \cpu.ex.r_12[5]$_DFFE_PP_  (.CLK(clknet_leaf_99_clk),
    .RESET_B(net1688),
    .D(_00831_),
    .Q_N(_14499_),
    .Q(\cpu.ex.r_12[5] ));
 sg13g2_dfrbp_1 \cpu.ex.r_12[6]$_DFFE_PP_  (.CLK(clknet_leaf_125_clk),
    .RESET_B(net1689),
    .D(_00832_),
    .Q_N(_14498_),
    .Q(\cpu.ex.r_12[6] ));
 sg13g2_dfrbp_1 \cpu.ex.r_12[7]$_DFFE_PP_  (.CLK(clknet_leaf_96_clk),
    .RESET_B(net1690),
    .D(_00833_),
    .Q_N(_14497_),
    .Q(\cpu.ex.r_12[7] ));
 sg13g2_dfrbp_1 \cpu.ex.r_12[8]$_DFFE_PP_  (.CLK(clknet_leaf_98_clk),
    .RESET_B(net1691),
    .D(_00834_),
    .Q_N(_14496_),
    .Q(\cpu.ex.r_12[8] ));
 sg13g2_dfrbp_1 \cpu.ex.r_12[9]$_DFFE_PP_  (.CLK(clknet_leaf_124_clk),
    .RESET_B(net1692),
    .D(_00835_),
    .Q_N(_14495_),
    .Q(\cpu.ex.r_12[9] ));
 sg13g2_dfrbp_1 \cpu.ex.r_13[0]$_DFFE_PP_  (.CLK(clknet_leaf_122_clk),
    .RESET_B(net1693),
    .D(_00836_),
    .Q_N(_14494_),
    .Q(\cpu.ex.r_13[0] ));
 sg13g2_dfrbp_1 \cpu.ex.r_13[10]$_DFFE_PP_  (.CLK(clknet_leaf_110_clk),
    .RESET_B(net1694),
    .D(_00837_),
    .Q_N(_14493_),
    .Q(\cpu.ex.r_13[10] ));
 sg13g2_dfrbp_1 \cpu.ex.r_13[11]$_DFFE_PP_  (.CLK(clknet_leaf_112_clk),
    .RESET_B(net1695),
    .D(_00838_),
    .Q_N(_14492_),
    .Q(\cpu.ex.r_13[11] ));
 sg13g2_dfrbp_1 \cpu.ex.r_13[12]$_DFFE_PP_  (.CLK(clknet_leaf_115_clk),
    .RESET_B(net1696),
    .D(_00839_),
    .Q_N(_14491_),
    .Q(\cpu.ex.r_13[12] ));
 sg13g2_dfrbp_1 \cpu.ex.r_13[13]$_DFFE_PP_  (.CLK(clknet_leaf_41_clk),
    .RESET_B(net1697),
    .D(_00840_),
    .Q_N(_14490_),
    .Q(\cpu.ex.r_13[13] ));
 sg13g2_dfrbp_1 \cpu.ex.r_13[14]$_DFFE_PP_  (.CLK(clknet_leaf_111_clk),
    .RESET_B(net1698),
    .D(_00841_),
    .Q_N(_14489_),
    .Q(\cpu.ex.r_13[14] ));
 sg13g2_dfrbp_1 \cpu.ex.r_13[15]$_DFFE_PP_  (.CLK(clknet_leaf_40_clk),
    .RESET_B(net1699),
    .D(_00842_),
    .Q_N(_14488_),
    .Q(\cpu.ex.r_13[15] ));
 sg13g2_dfrbp_1 \cpu.ex.r_13[1]$_DFFE_PP_  (.CLK(clknet_leaf_114_clk),
    .RESET_B(net1700),
    .D(_00843_),
    .Q_N(_14487_),
    .Q(\cpu.ex.r_13[1] ));
 sg13g2_dfrbp_1 \cpu.ex.r_13[2]$_DFFE_PP_  (.CLK(clknet_leaf_262_clk),
    .RESET_B(net1701),
    .D(_00844_),
    .Q_N(_14486_),
    .Q(\cpu.ex.r_13[2] ));
 sg13g2_dfrbp_1 \cpu.ex.r_13[3]$_DFFE_PP_  (.CLK(clknet_leaf_102_clk),
    .RESET_B(net1702),
    .D(_00845_),
    .Q_N(_14485_),
    .Q(\cpu.ex.r_13[3] ));
 sg13g2_dfrbp_1 \cpu.ex.r_13[4]$_DFFE_PP_  (.CLK(clknet_leaf_100_clk),
    .RESET_B(net1703),
    .D(_00846_),
    .Q_N(_14484_),
    .Q(\cpu.ex.r_13[4] ));
 sg13g2_dfrbp_1 \cpu.ex.r_13[5]$_DFFE_PP_  (.CLK(clknet_leaf_99_clk),
    .RESET_B(net1704),
    .D(_00847_),
    .Q_N(_14483_),
    .Q(\cpu.ex.r_13[5] ));
 sg13g2_dfrbp_1 \cpu.ex.r_13[6]$_DFFE_PP_  (.CLK(clknet_leaf_125_clk),
    .RESET_B(net1705),
    .D(_00848_),
    .Q_N(_14482_),
    .Q(\cpu.ex.r_13[6] ));
 sg13g2_dfrbp_1 \cpu.ex.r_13[7]$_DFFE_PP_  (.CLK(clknet_leaf_96_clk),
    .RESET_B(net1706),
    .D(_00849_),
    .Q_N(_14481_),
    .Q(\cpu.ex.r_13[7] ));
 sg13g2_dfrbp_1 \cpu.ex.r_13[8]$_DFFE_PP_  (.CLK(clknet_leaf_98_clk),
    .RESET_B(net1707),
    .D(_00850_),
    .Q_N(_14480_),
    .Q(\cpu.ex.r_13[8] ));
 sg13g2_dfrbp_1 \cpu.ex.r_13[9]$_DFFE_PP_  (.CLK(clknet_leaf_100_clk),
    .RESET_B(net1708),
    .D(_00851_),
    .Q_N(_14479_),
    .Q(\cpu.ex.r_13[9] ));
 sg13g2_dfrbp_1 \cpu.ex.r_14[0]$_DFFE_PP_  (.CLK(clknet_leaf_122_clk),
    .RESET_B(net1709),
    .D(_00852_),
    .Q_N(_14478_),
    .Q(\cpu.ex.r_14[0] ));
 sg13g2_dfrbp_1 \cpu.ex.r_14[10]$_DFFE_PP_  (.CLK(clknet_leaf_111_clk),
    .RESET_B(net1710),
    .D(_00853_),
    .Q_N(_14477_),
    .Q(\cpu.ex.r_14[10] ));
 sg13g2_dfrbp_1 \cpu.ex.r_14[11]$_DFFE_PP_  (.CLK(clknet_leaf_112_clk),
    .RESET_B(net1711),
    .D(_00854_),
    .Q_N(_14476_),
    .Q(\cpu.ex.r_14[11] ));
 sg13g2_dfrbp_1 \cpu.ex.r_14[12]$_DFFE_PP_  (.CLK(clknet_leaf_41_clk),
    .RESET_B(net1712),
    .D(_00855_),
    .Q_N(_14475_),
    .Q(\cpu.ex.r_14[12] ));
 sg13g2_dfrbp_1 \cpu.ex.r_14[13]$_DFFE_PP_  (.CLK(clknet_leaf_41_clk),
    .RESET_B(net1713),
    .D(_00856_),
    .Q_N(_14474_),
    .Q(\cpu.ex.r_14[13] ));
 sg13g2_dfrbp_1 \cpu.ex.r_14[14]$_DFFE_PP_  (.CLK(clknet_leaf_112_clk),
    .RESET_B(net1714),
    .D(_00857_),
    .Q_N(_14473_),
    .Q(\cpu.ex.r_14[14] ));
 sg13g2_dfrbp_1 \cpu.ex.r_14[15]$_DFFE_PP_  (.CLK(clknet_leaf_40_clk),
    .RESET_B(net1715),
    .D(_00858_),
    .Q_N(_14472_),
    .Q(\cpu.ex.r_14[15] ));
 sg13g2_dfrbp_1 \cpu.ex.r_14[1]$_DFFE_PP_  (.CLK(clknet_leaf_114_clk),
    .RESET_B(net1716),
    .D(_00859_),
    .Q_N(_14471_),
    .Q(\cpu.ex.r_14[1] ));
 sg13g2_dfrbp_1 \cpu.ex.r_14[2]$_DFFE_PP_  (.CLK(clknet_leaf_262_clk),
    .RESET_B(net1717),
    .D(_00860_),
    .Q_N(_14470_),
    .Q(\cpu.ex.r_14[2] ));
 sg13g2_dfrbp_1 \cpu.ex.r_14[3]$_DFFE_PP_  (.CLK(clknet_leaf_105_clk),
    .RESET_B(net1718),
    .D(_00861_),
    .Q_N(_14469_),
    .Q(\cpu.ex.r_14[3] ));
 sg13g2_dfrbp_1 \cpu.ex.r_14[4]$_DFFE_PP_  (.CLK(clknet_leaf_98_clk),
    .RESET_B(net1719),
    .D(_00862_),
    .Q_N(_14468_),
    .Q(\cpu.ex.r_14[4] ));
 sg13g2_dfrbp_1 \cpu.ex.r_14[5]$_DFFE_PP_  (.CLK(clknet_leaf_99_clk),
    .RESET_B(net1720),
    .D(_00863_),
    .Q_N(_14467_),
    .Q(\cpu.ex.r_14[5] ));
 sg13g2_dfrbp_1 \cpu.ex.r_14[6]$_DFFE_PP_  (.CLK(clknet_leaf_125_clk),
    .RESET_B(net1721),
    .D(_00864_),
    .Q_N(_14466_),
    .Q(\cpu.ex.r_14[6] ));
 sg13g2_dfrbp_1 \cpu.ex.r_14[7]$_DFFE_PP_  (.CLK(clknet_leaf_96_clk),
    .RESET_B(net1722),
    .D(_00865_),
    .Q_N(_14465_),
    .Q(\cpu.ex.r_14[7] ));
 sg13g2_dfrbp_1 \cpu.ex.r_14[8]$_DFFE_PP_  (.CLK(clknet_leaf_98_clk),
    .RESET_B(net1723),
    .D(_00866_),
    .Q_N(_14464_),
    .Q(\cpu.ex.r_14[8] ));
 sg13g2_dfrbp_1 \cpu.ex.r_14[9]$_DFFE_PP_  (.CLK(clknet_leaf_126_clk),
    .RESET_B(net1724),
    .D(_00867_),
    .Q_N(_14463_),
    .Q(\cpu.ex.r_14[9] ));
 sg13g2_dfrbp_1 \cpu.ex.r_15[0]$_DFFE_PP_  (.CLK(clknet_leaf_122_clk),
    .RESET_B(net1725),
    .D(_00868_),
    .Q_N(_14462_),
    .Q(\cpu.ex.r_15[0] ));
 sg13g2_dfrbp_1 \cpu.ex.r_15[10]$_DFFE_PP_  (.CLK(clknet_leaf_113_clk),
    .RESET_B(net1726),
    .D(_00869_),
    .Q_N(_00252_),
    .Q(\cpu.ex.r_15[10] ));
 sg13g2_dfrbp_1 \cpu.ex.r_15[11]$_DFFE_PP_  (.CLK(clknet_leaf_112_clk),
    .RESET_B(net1727),
    .D(_00870_),
    .Q_N(_00253_),
    .Q(\cpu.ex.r_15[11] ));
 sg13g2_dfrbp_1 \cpu.ex.r_15[12]$_DFFE_PP_  (.CLK(clknet_leaf_43_clk),
    .RESET_B(net1728),
    .D(_00871_),
    .Q_N(_00254_),
    .Q(\cpu.ex.r_15[12] ));
 sg13g2_dfrbp_1 \cpu.ex.r_15[13]$_DFFE_PP_  (.CLK(clknet_leaf_263_clk),
    .RESET_B(net1729),
    .D(_00872_),
    .Q_N(_00255_),
    .Q(\cpu.ex.r_15[13] ));
 sg13g2_dfrbp_1 \cpu.ex.r_15[14]$_DFFE_PP_  (.CLK(clknet_leaf_110_clk),
    .RESET_B(net1730),
    .D(_00873_),
    .Q_N(_00256_),
    .Q(\cpu.ex.r_15[14] ));
 sg13g2_dfrbp_1 \cpu.ex.r_15[15]$_DFFE_PP_  (.CLK(clknet_leaf_263_clk),
    .RESET_B(net1731),
    .D(_00874_),
    .Q_N(_14461_),
    .Q(\cpu.ex.r_15[15] ));
 sg13g2_dfrbp_1 \cpu.ex.r_15[1]$_DFFE_PP_  (.CLK(clknet_leaf_114_clk),
    .RESET_B(net1732),
    .D(_00875_),
    .Q_N(_00243_),
    .Q(\cpu.ex.r_15[1] ));
 sg13g2_dfrbp_1 \cpu.ex.r_15[2]$_DFFE_PP_  (.CLK(clknet_leaf_262_clk),
    .RESET_B(net1733),
    .D(_00876_),
    .Q_N(_00244_),
    .Q(\cpu.ex.r_15[2] ));
 sg13g2_dfrbp_1 \cpu.ex.r_15[3]$_DFFE_PP_  (.CLK(clknet_leaf_103_clk),
    .RESET_B(net1734),
    .D(_00877_),
    .Q_N(_00245_),
    .Q(\cpu.ex.r_15[3] ));
 sg13g2_dfrbp_1 \cpu.ex.r_15[4]$_DFFE_PP_  (.CLK(clknet_leaf_100_clk),
    .RESET_B(net1735),
    .D(_00878_),
    .Q_N(_00246_),
    .Q(\cpu.ex.r_15[4] ));
 sg13g2_dfrbp_1 \cpu.ex.r_15[5]$_DFFE_PP_  (.CLK(clknet_leaf_100_clk),
    .RESET_B(net1736),
    .D(_00879_),
    .Q_N(_00247_),
    .Q(\cpu.ex.r_15[5] ));
 sg13g2_dfrbp_1 \cpu.ex.r_15[6]$_DFFE_PP_  (.CLK(clknet_leaf_125_clk),
    .RESET_B(net1737),
    .D(_00880_),
    .Q_N(_00248_),
    .Q(\cpu.ex.r_15[6] ));
 sg13g2_dfrbp_1 \cpu.ex.r_15[7]$_DFFE_PP_  (.CLK(clknet_leaf_99_clk),
    .RESET_B(net1738),
    .D(_00881_),
    .Q_N(_00249_),
    .Q(\cpu.ex.r_15[7] ));
 sg13g2_dfrbp_1 \cpu.ex.r_15[8]$_DFFE_PP_  (.CLK(clknet_leaf_100_clk),
    .RESET_B(net1739),
    .D(_00882_),
    .Q_N(_00250_),
    .Q(\cpu.ex.r_15[8] ));
 sg13g2_dfrbp_1 \cpu.ex.r_15[9]$_DFFE_PP_  (.CLK(clknet_leaf_126_clk),
    .RESET_B(net1740),
    .D(_00883_),
    .Q_N(_00251_),
    .Q(\cpu.ex.r_15[9] ));
 sg13g2_dfrbp_1 \cpu.ex.r_8[0]$_DFFE_PP_  (.CLK(clknet_leaf_124_clk),
    .RESET_B(net1741),
    .D(_00884_),
    .Q_N(_14460_),
    .Q(\cpu.ex.r_8[0] ));
 sg13g2_dfrbp_1 \cpu.ex.r_8[10]$_DFFE_PP_  (.CLK(clknet_leaf_115_clk),
    .RESET_B(net1742),
    .D(_00885_),
    .Q_N(_14459_),
    .Q(\cpu.ex.r_8[10] ));
 sg13g2_dfrbp_1 \cpu.ex.r_8[11]$_DFFE_PP_  (.CLK(clknet_leaf_104_clk),
    .RESET_B(net1743),
    .D(_00886_),
    .Q_N(_14458_),
    .Q(\cpu.ex.r_8[11] ));
 sg13g2_dfrbp_1 \cpu.ex.r_8[12]$_DFFE_PP_  (.CLK(clknet_leaf_43_clk),
    .RESET_B(net1744),
    .D(_00887_),
    .Q_N(_14457_),
    .Q(\cpu.ex.r_8[12] ));
 sg13g2_dfrbp_1 \cpu.ex.r_8[13]$_DFFE_PP_  (.CLK(clknet_leaf_263_clk),
    .RESET_B(net1745),
    .D(_00888_),
    .Q_N(_14456_),
    .Q(\cpu.ex.r_8[13] ));
 sg13g2_dfrbp_1 \cpu.ex.r_8[14]$_DFFE_PP_  (.CLK(clknet_leaf_113_clk),
    .RESET_B(net1746),
    .D(_00889_),
    .Q_N(_14455_),
    .Q(\cpu.ex.r_8[14] ));
 sg13g2_dfrbp_1 \cpu.ex.r_8[15]$_DFFE_PP_  (.CLK(clknet_leaf_40_clk),
    .RESET_B(net1747),
    .D(_00890_),
    .Q_N(_14454_),
    .Q(\cpu.ex.r_8[15] ));
 sg13g2_dfrbp_1 \cpu.ex.r_8[1]$_DFFE_PP_  (.CLK(clknet_leaf_43_clk),
    .RESET_B(net1748),
    .D(_00891_),
    .Q_N(_14453_),
    .Q(\cpu.ex.r_8[1] ));
 sg13g2_dfrbp_1 \cpu.ex.r_8[2]$_DFFE_PP_  (.CLK(clknet_leaf_262_clk),
    .RESET_B(net1749),
    .D(_00892_),
    .Q_N(_14452_),
    .Q(\cpu.ex.r_8[2] ));
 sg13g2_dfrbp_1 \cpu.ex.r_8[3]$_DFFE_PP_  (.CLK(clknet_leaf_102_clk),
    .RESET_B(net1750),
    .D(_00893_),
    .Q_N(_14451_),
    .Q(\cpu.ex.r_8[3] ));
 sg13g2_dfrbp_1 \cpu.ex.r_8[4]$_DFFE_PP_  (.CLK(clknet_leaf_124_clk),
    .RESET_B(net1751),
    .D(_00894_),
    .Q_N(_14450_),
    .Q(\cpu.ex.r_8[4] ));
 sg13g2_dfrbp_1 \cpu.ex.r_8[5]$_DFFE_PP_  (.CLK(clknet_leaf_98_clk),
    .RESET_B(net1752),
    .D(_00895_),
    .Q_N(_14449_),
    .Q(\cpu.ex.r_8[5] ));
 sg13g2_dfrbp_1 \cpu.ex.r_8[6]$_DFFE_PP_  (.CLK(clknet_leaf_98_clk),
    .RESET_B(net1753),
    .D(_00896_),
    .Q_N(_14448_),
    .Q(\cpu.ex.r_8[6] ));
 sg13g2_dfrbp_1 \cpu.ex.r_8[7]$_DFFE_PP_  (.CLK(clknet_leaf_100_clk),
    .RESET_B(net1754),
    .D(_00897_),
    .Q_N(_14447_),
    .Q(\cpu.ex.r_8[7] ));
 sg13g2_dfrbp_1 \cpu.ex.r_8[8]$_DFFE_PP_  (.CLK(clknet_leaf_101_clk),
    .RESET_B(net1755),
    .D(_00898_),
    .Q_N(_14446_),
    .Q(\cpu.ex.r_8[8] ));
 sg13g2_dfrbp_1 \cpu.ex.r_8[9]$_DFFE_PP_  (.CLK(clknet_leaf_124_clk),
    .RESET_B(net1756),
    .D(_00899_),
    .Q_N(_14445_),
    .Q(\cpu.ex.r_8[9] ));
 sg13g2_dfrbp_1 \cpu.ex.r_9[0]$_DFFE_PP_  (.CLK(clknet_leaf_124_clk),
    .RESET_B(net1757),
    .D(_00900_),
    .Q_N(_14444_),
    .Q(\cpu.ex.r_9[0] ));
 sg13g2_dfrbp_1 \cpu.ex.r_9[10]$_DFFE_PP_  (.CLK(clknet_leaf_115_clk),
    .RESET_B(net1758),
    .D(_00901_),
    .Q_N(_14443_),
    .Q(\cpu.ex.r_9[10] ));
 sg13g2_dfrbp_1 \cpu.ex.r_9[11]$_DFFE_PP_  (.CLK(clknet_leaf_103_clk),
    .RESET_B(net1759),
    .D(_00902_),
    .Q_N(_14442_),
    .Q(\cpu.ex.r_9[11] ));
 sg13g2_dfrbp_1 \cpu.ex.r_9[12]$_DFFE_PP_  (.CLK(clknet_leaf_264_clk),
    .RESET_B(net1760),
    .D(_00903_),
    .Q_N(_14441_),
    .Q(\cpu.ex.r_9[12] ));
 sg13g2_dfrbp_1 \cpu.ex.r_9[13]$_DFFE_PP_  (.CLK(clknet_leaf_264_clk),
    .RESET_B(net1761),
    .D(_00904_),
    .Q_N(_14440_),
    .Q(\cpu.ex.r_9[13] ));
 sg13g2_dfrbp_1 \cpu.ex.r_9[14]$_DFFE_PP_  (.CLK(clknet_leaf_113_clk),
    .RESET_B(net1762),
    .D(_00905_),
    .Q_N(_14439_),
    .Q(\cpu.ex.r_9[14] ));
 sg13g2_dfrbp_1 \cpu.ex.r_9[15]$_DFFE_PP_  (.CLK(clknet_leaf_263_clk),
    .RESET_B(net1763),
    .D(_00906_),
    .Q_N(_14438_),
    .Q(\cpu.ex.r_9[15] ));
 sg13g2_dfrbp_1 \cpu.ex.r_9[1]$_DFFE_PP_  (.CLK(clknet_leaf_115_clk),
    .RESET_B(net1764),
    .D(_00907_),
    .Q_N(_14437_),
    .Q(\cpu.ex.r_9[1] ));
 sg13g2_dfrbp_1 \cpu.ex.r_9[2]$_DFFE_PP_  (.CLK(clknet_leaf_261_clk),
    .RESET_B(net1765),
    .D(_00908_),
    .Q_N(_14436_),
    .Q(\cpu.ex.r_9[2] ));
 sg13g2_dfrbp_1 \cpu.ex.r_9[3]$_DFFE_PP_  (.CLK(clknet_leaf_104_clk),
    .RESET_B(net1766),
    .D(_00909_),
    .Q_N(_14435_),
    .Q(\cpu.ex.r_9[3] ));
 sg13g2_dfrbp_1 \cpu.ex.r_9[4]$_DFFE_PP_  (.CLK(clknet_leaf_124_clk),
    .RESET_B(net1767),
    .D(_00910_),
    .Q_N(_14434_),
    .Q(\cpu.ex.r_9[4] ));
 sg13g2_dfrbp_1 \cpu.ex.r_9[5]$_DFFE_PP_  (.CLK(clknet_leaf_100_clk),
    .RESET_B(net1768),
    .D(_00911_),
    .Q_N(_14433_),
    .Q(\cpu.ex.r_9[5] ));
 sg13g2_dfrbp_1 \cpu.ex.r_9[6]$_DFFE_PP_  (.CLK(clknet_leaf_98_clk),
    .RESET_B(net1769),
    .D(_00912_),
    .Q_N(_14432_),
    .Q(\cpu.ex.r_9[6] ));
 sg13g2_dfrbp_1 \cpu.ex.r_9[7]$_DFFE_PP_  (.CLK(clknet_leaf_101_clk),
    .RESET_B(net1770),
    .D(_00913_),
    .Q_N(_14431_),
    .Q(\cpu.ex.r_9[7] ));
 sg13g2_dfrbp_1 \cpu.ex.r_9[8]$_DFFE_PP_  (.CLK(clknet_leaf_101_clk),
    .RESET_B(net1771),
    .D(_00914_),
    .Q_N(_14430_),
    .Q(\cpu.ex.r_9[8] ));
 sg13g2_dfrbp_1 \cpu.ex.r_9[9]$_DFFE_PP_  (.CLK(clknet_leaf_123_clk),
    .RESET_B(net1772),
    .D(_00915_),
    .Q_N(_14986_),
    .Q(\cpu.ex.r_9[9] ));
 sg13g2_dfrbp_1 \cpu.ex.r_branch_stall$_DFF_P_  (.CLK(clknet_leaf_117_clk),
    .RESET_B(net1773),
    .D(_00053_),
    .Q_N(_14429_),
    .Q(\cpu.ex.r_branch_stall ));
 sg13g2_dfrbp_1 \cpu.ex.r_cc$_DFFE_PP_  (.CLK(clknet_leaf_128_clk),
    .RESET_B(net1774),
    .D(_00916_),
    .Q_N(_14428_),
    .Q(\cpu.ex.r_cc ));
 sg13g2_dfrbp_1 \cpu.ex.r_d_flush_all$_SDFF_PP0_  (.CLK(clknet_leaf_178_clk),
    .RESET_B(net1775),
    .D(_00917_),
    .Q_N(_14987_),
    .Q(\cpu.d_flush_all ));
 sg13g2_dfrbp_1 \cpu.ex.r_div_running$_DFF_P_  (.CLK(clknet_leaf_118_clk),
    .RESET_B(net1776),
    .D(\cpu.ex.c_div_running ),
    .Q_N(_14427_),
    .Q(\cpu.ex.r_div_running ));
 sg13g2_dfrbp_1 \cpu.ex.r_epc[0]$_DFFE_PP_  (.CLK(clknet_leaf_114_clk),
    .RESET_B(net1777),
    .D(_00918_),
    .Q_N(_14426_),
    .Q(\cpu.ex.r_epc[1] ));
 sg13g2_dfrbp_1 \cpu.ex.r_epc[10]$_DFFE_PP_  (.CLK(clknet_leaf_112_clk),
    .RESET_B(net1778),
    .D(_00919_),
    .Q_N(_14425_),
    .Q(\cpu.ex.r_epc[11] ));
 sg13g2_dfrbp_1 \cpu.ex.r_epc[11]$_DFFE_PP_  (.CLK(clknet_leaf_263_clk),
    .RESET_B(net1779),
    .D(_00920_),
    .Q_N(_14424_),
    .Q(\cpu.ex.r_epc[12] ));
 sg13g2_dfrbp_1 \cpu.ex.r_epc[12]$_DFFE_PP_  (.CLK(clknet_leaf_264_clk),
    .RESET_B(net1780),
    .D(_00921_),
    .Q_N(_14423_),
    .Q(\cpu.ex.r_epc[13] ));
 sg13g2_dfrbp_1 \cpu.ex.r_epc[13]$_DFFE_PP_  (.CLK(clknet_leaf_112_clk),
    .RESET_B(net1781),
    .D(_00922_),
    .Q_N(_14422_),
    .Q(\cpu.ex.r_epc[14] ));
 sg13g2_dfrbp_1 \cpu.ex.r_epc[14]$_DFFE_PP_  (.CLK(clknet_leaf_40_clk),
    .RESET_B(net1782),
    .D(_00923_),
    .Q_N(_14421_),
    .Q(\cpu.ex.r_epc[15] ));
 sg13g2_dfrbp_1 \cpu.ex.r_epc[1]$_DFFE_PP_  (.CLK(clknet_leaf_261_clk),
    .RESET_B(net1783),
    .D(_00924_),
    .Q_N(_14420_),
    .Q(\cpu.ex.r_epc[2] ));
 sg13g2_dfrbp_1 \cpu.ex.r_epc[2]$_DFFE_PP_  (.CLK(clknet_leaf_105_clk),
    .RESET_B(net1784),
    .D(_00925_),
    .Q_N(_14419_),
    .Q(\cpu.ex.r_epc[3] ));
 sg13g2_dfrbp_1 \cpu.ex.r_epc[3]$_DFFE_PP_  (.CLK(clknet_leaf_100_clk),
    .RESET_B(net1785),
    .D(_00926_),
    .Q_N(_14418_),
    .Q(\cpu.ex.r_epc[4] ));
 sg13g2_dfrbp_1 \cpu.ex.r_epc[4]$_DFFE_PP_  (.CLK(clknet_leaf_101_clk),
    .RESET_B(net1786),
    .D(_00927_),
    .Q_N(_14417_),
    .Q(\cpu.ex.r_epc[5] ));
 sg13g2_dfrbp_1 \cpu.ex.r_epc[5]$_DFFE_PP_  (.CLK(clknet_leaf_101_clk),
    .RESET_B(net1787),
    .D(_00928_),
    .Q_N(_14416_),
    .Q(\cpu.ex.r_epc[6] ));
 sg13g2_dfrbp_1 \cpu.ex.r_epc[6]$_DFFE_PP_  (.CLK(clknet_leaf_101_clk),
    .RESET_B(net1788),
    .D(_00929_),
    .Q_N(_14415_),
    .Q(\cpu.ex.r_epc[7] ));
 sg13g2_dfrbp_1 \cpu.ex.r_epc[7]$_DFFE_PP_  (.CLK(clknet_leaf_101_clk),
    .RESET_B(net1789),
    .D(_00930_),
    .Q_N(_14414_),
    .Q(\cpu.ex.r_epc[8] ));
 sg13g2_dfrbp_1 \cpu.ex.r_epc[8]$_DFFE_PP_  (.CLK(clknet_leaf_123_clk),
    .RESET_B(net1790),
    .D(_00931_),
    .Q_N(_14413_),
    .Q(\cpu.ex.r_epc[9] ));
 sg13g2_dfrbp_1 \cpu.ex.r_epc[9]$_DFFE_PP_  (.CLK(clknet_leaf_113_clk),
    .RESET_B(net1791),
    .D(_00932_),
    .Q_N(_14412_),
    .Q(\cpu.ex.r_epc[10] ));
 sg13g2_dfrbp_1 \cpu.ex.r_fetch$_SDFF_PN1_  (.CLK(clknet_leaf_176_clk),
    .RESET_B(net1792),
    .D(_00933_),
    .Q_N(_00179_),
    .Q(\cpu.ex.ifetch ));
 sg13g2_dfrbp_1 \cpu.ex.r_flush_write$_SDFFE_PN0P_  (.CLK(clknet_leaf_176_clk),
    .RESET_B(net1793),
    .D(_00934_),
    .Q_N(_14411_),
    .Q(\cpu.dcache.flush_write ));
 sg13g2_dfrbp_1 \cpu.ex.r_i_flush_all$_SDFF_PP0_  (.CLK(clknet_leaf_177_clk),
    .RESET_B(net1794),
    .D(_00935_),
    .Q_N(_14410_),
    .Q(\cpu.ex.i_flush_all ));
 sg13g2_dfrbp_1 \cpu.ex.r_ie$_SDFFE_PP0P_  (.CLK(clknet_leaf_116_clk),
    .RESET_B(net1795),
    .D(_00936_),
    .Q_N(_14409_),
    .Q(\cpu.ex.r_ie ));
 sg13g2_dfrbp_1 \cpu.ex.r_io_access$_SDFFE_PN0P_  (.CLK(clknet_leaf_116_clk),
    .RESET_B(net1796),
    .D(_00937_),
    .Q_N(_00187_),
    .Q(\cpu.ex.io_access ));
 sg13g2_dfrbp_1 \cpu.ex.r_lr[0]$_DFFE_PP_  (.CLK(clknet_leaf_42_clk),
    .RESET_B(net1797),
    .D(_00938_),
    .Q_N(_14408_),
    .Q(\cpu.ex.r_lr[1] ));
 sg13g2_dfrbp_1 \cpu.ex.r_lr[10]$_DFFE_PP_  (.CLK(clknet_leaf_111_clk),
    .RESET_B(net1798),
    .D(_00939_),
    .Q_N(_14407_),
    .Q(\cpu.ex.r_lr[11] ));
 sg13g2_dfrbp_1 \cpu.ex.r_lr[11]$_DFFE_PP_  (.CLK(clknet_leaf_264_clk),
    .RESET_B(net1799),
    .D(_00940_),
    .Q_N(_14406_),
    .Q(\cpu.ex.r_lr[12] ));
 sg13g2_dfrbp_1 \cpu.ex.r_lr[12]$_DFFE_PP_  (.CLK(clknet_leaf_267_clk),
    .RESET_B(net1800),
    .D(_00941_),
    .Q_N(_14405_),
    .Q(\cpu.ex.r_lr[13] ));
 sg13g2_dfrbp_1 \cpu.ex.r_lr[13]$_DFFE_PP_  (.CLK(clknet_leaf_44_clk),
    .RESET_B(net1801),
    .D(_00942_),
    .Q_N(_14404_),
    .Q(\cpu.ex.r_lr[14] ));
 sg13g2_dfrbp_1 \cpu.ex.r_lr[14]$_DFFE_PP_  (.CLK(clknet_leaf_42_clk),
    .RESET_B(net1802),
    .D(_00943_),
    .Q_N(_14403_),
    .Q(\cpu.ex.r_lr[15] ));
 sg13g2_dfrbp_1 \cpu.ex.r_lr[1]$_DFFE_PP_  (.CLK(clknet_leaf_114_clk),
    .RESET_B(net1803),
    .D(_00944_),
    .Q_N(_14402_),
    .Q(\cpu.ex.r_lr[2] ));
 sg13g2_dfrbp_1 \cpu.ex.r_lr[2]$_DFFE_PP_  (.CLK(clknet_leaf_104_clk),
    .RESET_B(net1804),
    .D(_00945_),
    .Q_N(_14401_),
    .Q(\cpu.ex.r_lr[3] ));
 sg13g2_dfrbp_1 \cpu.ex.r_lr[3]$_DFFE_PP_  (.CLK(clknet_leaf_43_clk),
    .RESET_B(net1805),
    .D(_00946_),
    .Q_N(_14400_),
    .Q(\cpu.ex.r_lr[4] ));
 sg13g2_dfrbp_1 \cpu.ex.r_lr[4]$_DFFE_PP_  (.CLK(clknet_leaf_102_clk),
    .RESET_B(net1806),
    .D(_00947_),
    .Q_N(_14399_),
    .Q(\cpu.ex.r_lr[5] ));
 sg13g2_dfrbp_1 \cpu.ex.r_lr[5]$_DFFE_PP_  (.CLK(clknet_leaf_111_clk),
    .RESET_B(net1807),
    .D(_00948_),
    .Q_N(_14398_),
    .Q(\cpu.ex.r_lr[6] ));
 sg13g2_dfrbp_1 \cpu.ex.r_lr[6]$_DFFE_PP_  (.CLK(clknet_leaf_102_clk),
    .RESET_B(net1808),
    .D(_00949_),
    .Q_N(_14397_),
    .Q(\cpu.ex.r_lr[7] ));
 sg13g2_dfrbp_1 \cpu.ex.r_lr[7]$_DFFE_PP_  (.CLK(clknet_leaf_105_clk),
    .RESET_B(net1809),
    .D(_00950_),
    .Q_N(_14396_),
    .Q(\cpu.ex.r_lr[8] ));
 sg13g2_dfrbp_1 \cpu.ex.r_lr[8]$_DFFE_PP_  (.CLK(clknet_leaf_102_clk),
    .RESET_B(net1810),
    .D(_00951_),
    .Q_N(_14395_),
    .Q(\cpu.ex.r_lr[9] ));
 sg13g2_dfrbp_1 \cpu.ex.r_lr[9]$_DFFE_PP_  (.CLK(clknet_leaf_111_clk),
    .RESET_B(net1811),
    .D(_00952_),
    .Q_N(_14988_),
    .Q(\cpu.ex.r_lr[10] ));
 sg13g2_dfrbp_1 \cpu.ex.r_mult[0]$_DFF_P_  (.CLK(clknet_leaf_121_clk),
    .RESET_B(net1812),
    .D(\cpu.ex.c_mult[0] ),
    .Q_N(_14989_),
    .Q(\cpu.ex.r_mult[0] ));
 sg13g2_dfrbp_1 \cpu.ex.r_mult[10]$_DFF_P_  (.CLK(clknet_leaf_127_clk),
    .RESET_B(net1813),
    .D(\cpu.ex.c_mult[10] ),
    .Q_N(_14990_),
    .Q(\cpu.ex.r_mult[10] ));
 sg13g2_dfrbp_1 \cpu.ex.r_mult[11]$_DFF_P_  (.CLK(clknet_leaf_127_clk),
    .RESET_B(net1814),
    .D(\cpu.ex.c_mult[11] ),
    .Q_N(_14991_),
    .Q(\cpu.ex.r_mult[11] ));
 sg13g2_dfrbp_1 \cpu.ex.r_mult[12]$_DFF_P_  (.CLK(clknet_leaf_127_clk),
    .RESET_B(net1815),
    .D(\cpu.ex.c_mult[12] ),
    .Q_N(_14992_),
    .Q(\cpu.ex.r_mult[12] ));
 sg13g2_dfrbp_1 \cpu.ex.r_mult[13]$_DFF_P_  (.CLK(clknet_leaf_126_clk),
    .RESET_B(net1816),
    .D(\cpu.ex.c_mult[13] ),
    .Q_N(_14993_),
    .Q(\cpu.ex.r_mult[13] ));
 sg13g2_dfrbp_1 \cpu.ex.r_mult[14]$_DFF_P_  (.CLK(clknet_leaf_126_clk),
    .RESET_B(net1817),
    .D(\cpu.ex.c_mult[14] ),
    .Q_N(_00155_),
    .Q(\cpu.ex.r_mult[14] ));
 sg13g2_dfrbp_1 \cpu.ex.r_mult[15]$_DFF_P_  (.CLK(clknet_leaf_127_clk),
    .RESET_B(net1818),
    .D(\cpu.ex.c_mult[15] ),
    .Q_N(_14394_),
    .Q(\cpu.ex.r_mult[15] ));
 sg13g2_dfrbp_1 \cpu.ex.r_mult[16]$_DFFE_PP_  (.CLK(clknet_leaf_123_clk),
    .RESET_B(net1819),
    .D(_00953_),
    .Q_N(_00293_),
    .Q(\cpu.ex.r_mult[16] ));
 sg13g2_dfrbp_1 \cpu.ex.r_mult[17]$_DFFE_PP_  (.CLK(clknet_leaf_121_clk),
    .RESET_B(net1820),
    .D(_00954_),
    .Q_N(_00292_),
    .Q(\cpu.ex.r_mult[17] ));
 sg13g2_dfrbp_1 \cpu.ex.r_mult[18]$_DFFE_PP_  (.CLK(clknet_leaf_121_clk),
    .RESET_B(net1821),
    .D(_00955_),
    .Q_N(_00291_),
    .Q(\cpu.ex.r_mult[18] ));
 sg13g2_dfrbp_1 \cpu.ex.r_mult[19]$_DFFE_PP_  (.CLK(clknet_leaf_121_clk),
    .RESET_B(net1822),
    .D(_00956_),
    .Q_N(_00290_),
    .Q(\cpu.ex.r_mult[19] ));
 sg13g2_dfrbp_1 \cpu.ex.r_mult[1]$_DFF_P_  (.CLK(clknet_leaf_120_clk),
    .RESET_B(net1823),
    .D(\cpu.ex.c_mult[1] ),
    .Q_N(_14393_),
    .Q(\cpu.ex.r_mult[1] ));
 sg13g2_dfrbp_1 \cpu.ex.r_mult[20]$_DFFE_PP_  (.CLK(clknet_leaf_121_clk),
    .RESET_B(net1824),
    .D(_00957_),
    .Q_N(_00289_),
    .Q(\cpu.ex.r_mult[20] ));
 sg13g2_dfrbp_1 \cpu.ex.r_mult[21]$_DFFE_PP_  (.CLK(clknet_leaf_123_clk),
    .RESET_B(net1825),
    .D(_00958_),
    .Q_N(_00288_),
    .Q(\cpu.ex.r_mult[21] ));
 sg13g2_dfrbp_1 \cpu.ex.r_mult[22]$_DFFE_PP_  (.CLK(clknet_leaf_122_clk),
    .RESET_B(net1826),
    .D(_00959_),
    .Q_N(_14392_),
    .Q(\cpu.ex.r_mult[22] ));
 sg13g2_dfrbp_1 \cpu.ex.r_mult[23]$_DFFE_PP_  (.CLK(clknet_leaf_123_clk),
    .RESET_B(net1827),
    .D(_00960_),
    .Q_N(_00287_),
    .Q(\cpu.ex.r_mult[23] ));
 sg13g2_dfrbp_1 \cpu.ex.r_mult[24]$_DFFE_PP_  (.CLK(clknet_leaf_122_clk),
    .RESET_B(net1828),
    .D(_00961_),
    .Q_N(_00286_),
    .Q(\cpu.ex.r_mult[24] ));
 sg13g2_dfrbp_1 \cpu.ex.r_mult[25]$_DFFE_PP_  (.CLK(clknet_leaf_123_clk),
    .RESET_B(net1829),
    .D(_00962_),
    .Q_N(_00285_),
    .Q(\cpu.ex.r_mult[25] ));
 sg13g2_dfrbp_1 \cpu.ex.r_mult[26]$_DFFE_PP_  (.CLK(clknet_leaf_123_clk),
    .RESET_B(net1830),
    .D(_00963_),
    .Q_N(_14391_),
    .Q(\cpu.ex.r_mult[26] ));
 sg13g2_dfrbp_1 \cpu.ex.r_mult[27]$_DFFE_PP_  (.CLK(clknet_leaf_126_clk),
    .RESET_B(net1831),
    .D(_00964_),
    .Q_N(_00284_),
    .Q(\cpu.ex.r_mult[27] ));
 sg13g2_dfrbp_1 \cpu.ex.r_mult[28]$_DFFE_PP_  (.CLK(clknet_leaf_125_clk),
    .RESET_B(net1832),
    .D(_00965_),
    .Q_N(_14390_),
    .Q(\cpu.ex.r_mult[28] ));
 sg13g2_dfrbp_1 \cpu.ex.r_mult[29]$_DFFE_PP_  (.CLK(clknet_leaf_125_clk),
    .RESET_B(net1833),
    .D(_00966_),
    .Q_N(_14994_),
    .Q(\cpu.ex.r_mult[29] ));
 sg13g2_dfrbp_1 \cpu.ex.r_mult[2]$_DFF_P_  (.CLK(clknet_leaf_120_clk),
    .RESET_B(net1834),
    .D(\cpu.ex.c_mult[2] ),
    .Q_N(_14389_),
    .Q(\cpu.ex.r_mult[2] ));
 sg13g2_dfrbp_1 \cpu.ex.r_mult[30]$_DFFE_PP_  (.CLK(clknet_leaf_126_clk),
    .RESET_B(net1835),
    .D(_00967_),
    .Q_N(_00283_),
    .Q(\cpu.ex.r_mult[30] ));
 sg13g2_dfrbp_1 \cpu.ex.r_mult[31]$_DFFE_PP_  (.CLK(clknet_leaf_126_clk),
    .RESET_B(net1836),
    .D(_00968_),
    .Q_N(_14995_),
    .Q(\cpu.ex.r_mult[31] ));
 sg13g2_dfrbp_1 \cpu.ex.r_mult[3]$_DFF_P_  (.CLK(clknet_leaf_129_clk),
    .RESET_B(net1837),
    .D(\cpu.ex.c_mult[3] ),
    .Q_N(_14996_),
    .Q(\cpu.ex.r_mult[3] ));
 sg13g2_dfrbp_1 \cpu.ex.r_mult[4]$_DFF_P_  (.CLK(clknet_leaf_127_clk),
    .RESET_B(net1838),
    .D(\cpu.ex.c_mult[4] ),
    .Q_N(_14997_),
    .Q(\cpu.ex.r_mult[4] ));
 sg13g2_dfrbp_1 \cpu.ex.r_mult[5]$_DFF_P_  (.CLK(clknet_leaf_128_clk),
    .RESET_B(net1839),
    .D(\cpu.ex.c_mult[5] ),
    .Q_N(_14998_),
    .Q(\cpu.ex.r_mult[5] ));
 sg13g2_dfrbp_1 \cpu.ex.r_mult[6]$_DFF_P_  (.CLK(clknet_leaf_128_clk),
    .RESET_B(net1840),
    .D(\cpu.ex.c_mult[6] ),
    .Q_N(_14999_),
    .Q(\cpu.ex.r_mult[6] ));
 sg13g2_dfrbp_1 \cpu.ex.r_mult[7]$_DFF_P_  (.CLK(clknet_leaf_128_clk),
    .RESET_B(net1841),
    .D(\cpu.ex.c_mult[7] ),
    .Q_N(_15000_),
    .Q(\cpu.ex.r_mult[7] ));
 sg13g2_dfrbp_1 \cpu.ex.r_mult[8]$_DFF_P_  (.CLK(clknet_leaf_128_clk),
    .RESET_B(net1842),
    .D(\cpu.ex.c_mult[8] ),
    .Q_N(_15001_),
    .Q(\cpu.ex.r_mult[8] ));
 sg13g2_dfrbp_1 \cpu.ex.r_mult[9]$_DFF_P_  (.CLK(clknet_leaf_127_clk),
    .RESET_B(net1843),
    .D(\cpu.ex.c_mult[9] ),
    .Q_N(_15002_),
    .Q(\cpu.ex.r_mult[9] ));
 sg13g2_dfrbp_1 \cpu.ex.r_mult_off[0]$_DFF_P_  (.CLK(clknet_leaf_119_clk),
    .RESET_B(net1844),
    .D(\cpu.ex.c_mult_off[0] ),
    .Q_N(_15003_),
    .Q(\cpu.ex.r_mult_off[0] ));
 sg13g2_dfrbp_1 \cpu.ex.r_mult_off[1]$_DFF_P_  (.CLK(clknet_leaf_119_clk),
    .RESET_B(net1845),
    .D(\cpu.ex.c_mult_off[1] ),
    .Q_N(_15004_),
    .Q(\cpu.ex.r_mult_off[1] ));
 sg13g2_dfrbp_1 \cpu.ex.r_mult_off[2]$_DFF_P_  (.CLK(clknet_leaf_121_clk),
    .RESET_B(net1846),
    .D(\cpu.ex.c_mult_off[2] ),
    .Q_N(_15005_),
    .Q(\cpu.ex.r_mult_off[2] ));
 sg13g2_dfrbp_1 \cpu.ex.r_mult_off[3]$_DFF_P_  (.CLK(clknet_leaf_119_clk),
    .RESET_B(net1847),
    .D(\cpu.ex.c_mult_off[3] ),
    .Q_N(_15006_),
    .Q(\cpu.ex.r_mult_off[3] ));
 sg13g2_dfrbp_1 \cpu.ex.r_mult_running$_DFF_P_  (.CLK(clknet_leaf_121_clk),
    .RESET_B(net1848),
    .D(\cpu.ex.c_mult_running ),
    .Q_N(_00189_),
    .Q(\cpu.ex.r_mult_running ));
 sg13g2_dfrbp_1 \cpu.ex.r_pc[0]$_DFFE_PP_  (.CLK(clknet_leaf_175_clk),
    .RESET_B(net1849),
    .D(_00969_),
    .Q_N(_00190_),
    .Q(\cpu.ex.pc[1] ));
 sg13g2_dfrbp_1 \cpu.ex.r_pc[10]$_DFFE_PP_  (.CLK(clknet_leaf_120_clk),
    .RESET_B(net1850),
    .D(_00970_),
    .Q_N(_00274_),
    .Q(\cpu.ex.pc[11] ));
 sg13g2_dfrbp_1 \cpu.ex.r_pc[11]$_DFFE_PP_  (.CLK(clknet_leaf_175_clk),
    .RESET_B(net1851),
    .D(_00971_),
    .Q_N(_00273_),
    .Q(\cpu.ex.pc[12] ));
 sg13g2_dfrbp_1 \cpu.ex.r_pc[12]$_DFFE_PP_  (.CLK(clknet_leaf_120_clk),
    .RESET_B(net1852),
    .D(_00972_),
    .Q_N(_00186_),
    .Q(\cpu.ex.pc[13] ));
 sg13g2_dfrbp_1 \cpu.ex.r_pc[13]$_DFFE_PP_  (.CLK(clknet_leaf_120_clk),
    .RESET_B(net1853),
    .D(_00973_),
    .Q_N(_00185_),
    .Q(\cpu.ex.pc[14] ));
 sg13g2_dfrbp_1 \cpu.ex.r_pc[14]$_DFFE_PP_  (.CLK(clknet_leaf_119_clk),
    .RESET_B(net1854),
    .D(_00974_),
    .Q_N(_00184_),
    .Q(\cpu.ex.pc[15] ));
 sg13g2_dfrbp_1 \cpu.ex.r_pc[1]$_DFFE_PP_  (.CLK(clknet_leaf_175_clk),
    .RESET_B(net1855),
    .D(_00975_),
    .Q_N(_00281_),
    .Q(\cpu.ex.pc[2] ));
 sg13g2_dfrbp_1 \cpu.ex.r_pc[2]$_DFFE_PP_  (.CLK(clknet_leaf_173_clk),
    .RESET_B(net1856),
    .D(_00976_),
    .Q_N(_00181_),
    .Q(\cpu.ex.pc[3] ));
 sg13g2_dfrbp_1 \cpu.ex.r_pc[3]$_DFFE_PP_  (.CLK(clknet_leaf_171_clk),
    .RESET_B(net1857),
    .D(_00977_),
    .Q_N(_00180_),
    .Q(\cpu.ex.pc[4] ));
 sg13g2_dfrbp_1 \cpu.ex.r_pc[4]$_DFFE_PP_  (.CLK(clknet_leaf_173_clk),
    .RESET_B(net1858),
    .D(_00978_),
    .Q_N(_00280_),
    .Q(\cpu.ex.pc[5] ));
 sg13g2_dfrbp_1 \cpu.ex.r_pc[5]$_DFFE_PP_  (.CLK(clknet_leaf_119_clk),
    .RESET_B(net1859),
    .D(_00979_),
    .Q_N(_00279_),
    .Q(\cpu.ex.pc[6] ));
 sg13g2_dfrbp_1 \cpu.ex.r_pc[6]$_DFFE_PP_  (.CLK(clknet_leaf_119_clk),
    .RESET_B(net1860),
    .D(_00980_),
    .Q_N(_00278_),
    .Q(\cpu.ex.pc[7] ));
 sg13g2_dfrbp_1 \cpu.ex.r_pc[7]$_DFFE_PP_  (.CLK(clknet_leaf_120_clk),
    .RESET_B(net1861),
    .D(_00981_),
    .Q_N(_00277_),
    .Q(\cpu.ex.pc[8] ));
 sg13g2_dfrbp_1 \cpu.ex.r_pc[8]$_DFFE_PP_  (.CLK(clknet_leaf_120_clk),
    .RESET_B(net1862),
    .D(_00982_),
    .Q_N(_00276_),
    .Q(\cpu.ex.pc[9] ));
 sg13g2_dfrbp_1 \cpu.ex.r_pc[9]$_DFFE_PP_  (.CLK(clknet_leaf_120_clk),
    .RESET_B(net1863),
    .D(_00983_),
    .Q_N(_00275_),
    .Q(\cpu.ex.pc[10] ));
 sg13g2_dfrbp_1 \cpu.ex.r_prev_ie$_SDFFE_PN0P_  (.CLK(clknet_leaf_177_clk),
    .RESET_B(net1864),
    .D(_00984_),
    .Q_N(_14388_),
    .Q(\cpu.ex.r_prev_ie ));
 sg13g2_dfrbp_1 \cpu.ex.r_read_stall$_SDFFE_PN0P_  (.CLK(clknet_leaf_176_clk),
    .RESET_B(net1865),
    .D(_00985_),
    .Q_N(_00188_),
    .Q(\cpu.ex.r_read_stall ));
 sg13g2_dfrbp_1 \cpu.ex.r_set_cc$_DFFE_PP_  (.CLK(clknet_leaf_176_clk),
    .RESET_B(net1866),
    .D(_00986_),
    .Q_N(_14387_),
    .Q(\cpu.ex.r_set_cc ));
 sg13g2_dfrbp_1 \cpu.ex.r_sp[0]$_DFFE_PP_  (.CLK(clknet_leaf_114_clk),
    .RESET_B(net1867),
    .D(_00987_),
    .Q_N(_14386_),
    .Q(\cpu.ex.r_sp[1] ));
 sg13g2_dfrbp_1 \cpu.ex.r_sp[10]$_DFFE_PP_  (.CLK(clknet_leaf_260_clk),
    .RESET_B(net1868),
    .D(_00988_),
    .Q_N(_14385_),
    .Q(\cpu.ex.r_sp[11] ));
 sg13g2_dfrbp_1 \cpu.ex.r_sp[11]$_DFFE_PP_  (.CLK(clknet_leaf_263_clk),
    .RESET_B(net1869),
    .D(_00989_),
    .Q_N(_14384_),
    .Q(\cpu.ex.r_sp[12] ));
 sg13g2_dfrbp_1 \cpu.ex.r_sp[12]$_DFFE_PP_  (.CLK(clknet_leaf_261_clk),
    .RESET_B(net1870),
    .D(_00990_),
    .Q_N(_14383_),
    .Q(\cpu.ex.r_sp[13] ));
 sg13g2_dfrbp_1 \cpu.ex.r_sp[13]$_DFFE_PP_  (.CLK(clknet_leaf_260_clk),
    .RESET_B(net1871),
    .D(_00991_),
    .Q_N(_14382_),
    .Q(\cpu.ex.r_sp[14] ));
 sg13g2_dfrbp_1 \cpu.ex.r_sp[14]$_DFFE_PP_  (.CLK(clknet_leaf_40_clk),
    .RESET_B(net1872),
    .D(_00992_),
    .Q_N(_14381_),
    .Q(\cpu.ex.r_sp[15] ));
 sg13g2_dfrbp_1 \cpu.ex.r_sp[1]$_DFFE_PP_  (.CLK(clknet_leaf_261_clk),
    .RESET_B(net1873),
    .D(_00993_),
    .Q_N(_14380_),
    .Q(\cpu.ex.r_sp[2] ));
 sg13g2_dfrbp_1 \cpu.ex.r_sp[2]$_DFFE_PP_  (.CLK(clknet_leaf_105_clk),
    .RESET_B(net1874),
    .D(_00994_),
    .Q_N(_14379_),
    .Q(\cpu.ex.r_sp[3] ));
 sg13g2_dfrbp_1 \cpu.ex.r_sp[3]$_DFFE_PP_  (.CLK(clknet_leaf_102_clk),
    .RESET_B(net1875),
    .D(_00995_),
    .Q_N(_14378_),
    .Q(\cpu.ex.r_sp[4] ));
 sg13g2_dfrbp_1 \cpu.ex.r_sp[4]$_DFFE_PP_  (.CLK(clknet_leaf_102_clk),
    .RESET_B(net1876),
    .D(_00996_),
    .Q_N(_14377_),
    .Q(\cpu.ex.r_sp[5] ));
 sg13g2_dfrbp_1 \cpu.ex.r_sp[5]$_DFFE_PP_  (.CLK(clknet_leaf_125_clk),
    .RESET_B(net1877),
    .D(_00997_),
    .Q_N(_14376_),
    .Q(\cpu.ex.r_sp[6] ));
 sg13g2_dfrbp_1 \cpu.ex.r_sp[6]$_DFFE_PP_  (.CLK(clknet_leaf_98_clk),
    .RESET_B(net1878),
    .D(_00998_),
    .Q_N(_14375_),
    .Q(\cpu.ex.r_sp[7] ));
 sg13g2_dfrbp_1 \cpu.ex.r_sp[7]$_DFFE_PP_  (.CLK(clknet_leaf_99_clk),
    .RESET_B(net1879),
    .D(_00999_),
    .Q_N(_14374_),
    .Q(\cpu.ex.r_sp[8] ));
 sg13g2_dfrbp_1 \cpu.ex.r_sp[8]$_DFFE_PP_  (.CLK(clknet_leaf_125_clk),
    .RESET_B(net1880),
    .D(_01000_),
    .Q_N(_14373_),
    .Q(\cpu.ex.r_sp[9] ));
 sg13g2_dfrbp_1 \cpu.ex.r_sp[9]$_DFFE_PP_  (.CLK(clknet_leaf_117_clk),
    .RESET_B(net1881),
    .D(_01001_),
    .Q_N(_14372_),
    .Q(\cpu.ex.r_sp[10] ));
 sg13g2_dfrbp_1 \cpu.ex.r_stmp[0]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_117_clk),
    .RESET_B(net1882),
    .D(_01002_),
    .Q_N(_14371_),
    .Q(\cpu.ex.r_stmp[0] ));
 sg13g2_dfrbp_1 \cpu.ex.r_stmp[10]$_DFFE_PP_  (.CLK(clknet_leaf_113_clk),
    .RESET_B(net1883),
    .D(_01003_),
    .Q_N(_14370_),
    .Q(\cpu.ex.r_stmp[10] ));
 sg13g2_dfrbp_1 \cpu.ex.r_stmp[11]$_DFFE_PP_  (.CLK(clknet_leaf_113_clk),
    .RESET_B(net1884),
    .D(_01004_),
    .Q_N(_14369_),
    .Q(\cpu.ex.r_stmp[11] ));
 sg13g2_dfrbp_1 \cpu.ex.r_stmp[12]$_DFFE_PP_  (.CLK(clknet_leaf_41_clk),
    .RESET_B(net1885),
    .D(_01005_),
    .Q_N(_14368_),
    .Q(\cpu.ex.r_stmp[12] ));
 sg13g2_dfrbp_1 \cpu.ex.r_stmp[13]$_DFFE_PP_  (.CLK(clknet_leaf_116_clk),
    .RESET_B(net1886),
    .D(_01006_),
    .Q_N(_14367_),
    .Q(\cpu.ex.r_stmp[13] ));
 sg13g2_dfrbp_1 \cpu.ex.r_stmp[14]$_DFFE_PP_  (.CLK(clknet_leaf_118_clk),
    .RESET_B(net1887),
    .D(_01007_),
    .Q_N(_14366_),
    .Q(\cpu.ex.r_stmp[14] ));
 sg13g2_dfrbp_1 \cpu.ex.r_stmp[15]$_DFFE_PP_  (.CLK(clknet_leaf_41_clk),
    .RESET_B(net1888),
    .D(_01008_),
    .Q_N(_14365_),
    .Q(\cpu.ex.r_stmp[15] ));
 sg13g2_dfrbp_1 \cpu.ex.r_stmp[1]$_DFFE_PP_  (.CLK(clknet_leaf_114_clk),
    .RESET_B(net1889),
    .D(_01009_),
    .Q_N(_14364_),
    .Q(\cpu.ex.r_stmp[1] ));
 sg13g2_dfrbp_1 \cpu.ex.r_stmp[2]$_DFFE_PP_  (.CLK(clknet_leaf_43_clk),
    .RESET_B(net1890),
    .D(_01010_),
    .Q_N(_14363_),
    .Q(\cpu.ex.r_stmp[2] ));
 sg13g2_dfrbp_1 \cpu.ex.r_stmp[3]$_DFFE_PP_  (.CLK(clknet_leaf_103_clk),
    .RESET_B(net1891),
    .D(_01011_),
    .Q_N(_14362_),
    .Q(\cpu.ex.r_stmp[3] ));
 sg13g2_dfrbp_1 \cpu.ex.r_stmp[4]$_DFFE_PP_  (.CLK(clknet_leaf_103_clk),
    .RESET_B(net1892),
    .D(_01012_),
    .Q_N(_14361_),
    .Q(\cpu.ex.r_stmp[4] ));
 sg13g2_dfrbp_1 \cpu.ex.r_stmp[5]$_DFFE_PP_  (.CLK(clknet_leaf_103_clk),
    .RESET_B(net1893),
    .D(_01013_),
    .Q_N(_14360_),
    .Q(\cpu.ex.r_stmp[5] ));
 sg13g2_dfrbp_1 \cpu.ex.r_stmp[6]$_DFFE_PP_  (.CLK(clknet_leaf_121_clk),
    .RESET_B(net1894),
    .D(_01014_),
    .Q_N(_14359_),
    .Q(\cpu.ex.r_stmp[6] ));
 sg13g2_dfrbp_1 \cpu.ex.r_stmp[7]$_DFFE_PP_  (.CLK(clknet_leaf_103_clk),
    .RESET_B(net1895),
    .D(_01015_),
    .Q_N(_14358_),
    .Q(\cpu.ex.r_stmp[7] ));
 sg13g2_dfrbp_1 \cpu.ex.r_stmp[8]$_DFFE_PP_  (.CLK(clknet_leaf_103_clk),
    .RESET_B(net1896),
    .D(_01016_),
    .Q_N(_14357_),
    .Q(\cpu.ex.r_stmp[8] ));
 sg13g2_dfrbp_1 \cpu.ex.r_stmp[9]$_DFFE_PP_  (.CLK(clknet_leaf_122_clk),
    .RESET_B(net1897),
    .D(_01017_),
    .Q_N(_14356_),
    .Q(\cpu.ex.r_stmp[9] ));
 sg13g2_dfrbp_1 \cpu.ex.r_wb[0]$_DFFE_PP_  (.CLK(clknet_leaf_116_clk),
    .RESET_B(net1898),
    .D(_01018_),
    .Q_N(_00241_),
    .Q(\cpu.ex.mmu_reg_data[0] ));
 sg13g2_dfrbp_1 \cpu.ex.r_wb[10]$_DFFE_PP_  (.CLK(clknet_leaf_118_clk),
    .RESET_B(net1899),
    .D(_01019_),
    .Q_N(_00223_),
    .Q(\cpu.addr[10] ));
 sg13g2_dfrbp_1 \cpu.ex.r_wb[11]$_DFFE_PP_  (.CLK(clknet_leaf_118_clk),
    .RESET_B(net1900),
    .D(_01020_),
    .Q_N(_00225_),
    .Q(\cpu.addr[11] ));
 sg13g2_dfrbp_1 \cpu.ex.r_wb[12]$_DFFE_PP_  (.CLK(clknet_leaf_180_clk),
    .RESET_B(net1901),
    .D(_01021_),
    .Q_N(_14355_),
    .Q(\cpu.addr[12] ));
 sg13g2_dfrbp_1 \cpu.ex.r_wb[13]$_DFFE_PP_  (.CLK(clknet_leaf_176_clk),
    .RESET_B(net1902),
    .D(_01022_),
    .Q_N(_14354_),
    .Q(\cpu.addr[13] ));
 sg13g2_dfrbp_1 \cpu.ex.r_wb[14]$_DFFE_PP_  (.CLK(clknet_leaf_119_clk),
    .RESET_B(net1903),
    .D(_01023_),
    .Q_N(_14353_),
    .Q(\cpu.addr[14] ));
 sg13g2_dfrbp_1 \cpu.ex.r_wb[15]$_DFFE_PP_  (.CLK(clknet_leaf_176_clk),
    .RESET_B(net1904),
    .D(_01024_),
    .Q_N(_14352_),
    .Q(\cpu.addr[15] ));
 sg13g2_dfrbp_1 \cpu.ex.r_wb[1]$_DFFE_PP_  (.CLK(clknet_leaf_48_clk),
    .RESET_B(net1905),
    .D(_01025_),
    .Q_N(_00259_),
    .Q(\cpu.addr[1] ));
 sg13g2_dfrbp_1 \cpu.ex.r_wb[2]$_DFFE_PP_  (.CLK(clknet_leaf_44_clk),
    .RESET_B(net1906),
    .D(_01026_),
    .Q_N(_14351_),
    .Q(\cpu.addr[2] ));
 sg13g2_dfrbp_1 \cpu.ex.r_wb[3]$_DFFE_PP_  (.CLK(clknet_leaf_44_clk),
    .RESET_B(net1907),
    .D(_01027_),
    .Q_N(_00207_),
    .Q(\cpu.addr[3] ));
 sg13g2_dfrbp_1 \cpu.ex.r_wb[4]$_DFFE_PP_  (.CLK(clknet_leaf_110_clk),
    .RESET_B(net1908),
    .D(_01028_),
    .Q_N(_00212_),
    .Q(\cpu.addr[4] ));
 sg13g2_dfrbp_1 \cpu.ex.r_wb[5]$_DFFE_PP_  (.CLK(clknet_leaf_109_clk),
    .RESET_B(net1909),
    .D(_01029_),
    .Q_N(_00213_),
    .Q(\cpu.addr[5] ));
 sg13g2_dfrbp_1 \cpu.ex.r_wb[6]$_DFFE_PP_  (.CLK(clknet_leaf_110_clk),
    .RESET_B(net1910),
    .D(_01030_),
    .Q_N(_00215_),
    .Q(\cpu.addr[6] ));
 sg13g2_dfrbp_1 \cpu.ex.r_wb[7]$_DFFE_PP_  (.CLK(clknet_leaf_118_clk),
    .RESET_B(net1911),
    .D(_01031_),
    .Q_N(_00217_),
    .Q(\cpu.addr[7] ));
 sg13g2_dfrbp_1 \cpu.ex.r_wb[8]$_DFFE_PP_  (.CLK(clknet_leaf_112_clk),
    .RESET_B(net1912),
    .D(_01032_),
    .Q_N(_00219_),
    .Q(\cpu.addr[8] ));
 sg13g2_dfrbp_1 \cpu.ex.r_wb[9]$_DFFE_PP_  (.CLK(clknet_leaf_118_clk),
    .RESET_B(net1913),
    .D(_01033_),
    .Q_N(_00221_),
    .Q(\cpu.addr[9] ));
 sg13g2_dfrbp_1 \cpu.ex.r_wb_addr[0]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_118_clk),
    .RESET_B(net1914),
    .D(_01034_),
    .Q_N(_14350_),
    .Q(\cpu.ex.r_wb_addr[0] ));
 sg13g2_dfrbp_1 \cpu.ex.r_wb_addr[1]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_117_clk),
    .RESET_B(net1915),
    .D(_01035_),
    .Q_N(_14349_),
    .Q(\cpu.ex.r_wb_addr[1] ));
 sg13g2_dfrbp_1 \cpu.ex.r_wb_addr[2]$_SDFFCE_PP0P_  (.CLK(clknet_leaf_117_clk),
    .RESET_B(net1916),
    .D(_01036_),
    .Q_N(_14348_),
    .Q(\cpu.ex.r_wb_addr[2] ));
 sg13g2_dfrbp_1 \cpu.ex.r_wb_addr[3]$_SDFFCE_PP0P_  (.CLK(clknet_leaf_118_clk),
    .RESET_B(net1917),
    .D(_01037_),
    .Q_N(_14347_),
    .Q(\cpu.ex.r_wb_addr[3] ));
 sg13g2_dfrbp_1 \cpu.ex.r_wb_swapsp$_DFFE_PP_  (.CLK(clknet_leaf_117_clk),
    .RESET_B(net1918),
    .D(_01038_),
    .Q_N(_15007_),
    .Q(\cpu.ex.r_wb_swapsp ));
 sg13g2_dfrbp_1 \cpu.ex.r_wb_valid$_DFF_P_  (.CLK(clknet_leaf_119_clk),
    .RESET_B(net1919),
    .D(_00054_),
    .Q_N(_00240_),
    .Q(\cpu.ex.r_wb_valid ));
 sg13g2_dfrbp_1 \cpu.ex.r_wdata[0]$_DFFE_PP_  (.CLK(clknet_leaf_53_clk),
    .RESET_B(net1920),
    .D(_01039_),
    .Q_N(_00208_),
    .Q(\cpu.dcache.wdata[0] ));
 sg13g2_dfrbp_1 \cpu.ex.r_wdata[10]$_DFFE_PP_  (.CLK(clknet_leaf_43_clk),
    .RESET_B(net1921),
    .D(_01040_),
    .Q_N(_14346_),
    .Q(\cpu.dcache.wdata[10] ));
 sg13g2_dfrbp_1 \cpu.ex.r_wdata[11]$_DFFE_PP_  (.CLK(clknet_leaf_45_clk),
    .RESET_B(net1922),
    .D(_01041_),
    .Q_N(_14345_),
    .Q(\cpu.dcache.wdata[11] ));
 sg13g2_dfrbp_1 \cpu.ex.r_wdata[12]$_DFFE_PP_  (.CLK(clknet_leaf_45_clk),
    .RESET_B(net1923),
    .D(_01042_),
    .Q_N(_14344_),
    .Q(\cpu.dcache.wdata[12] ));
 sg13g2_dfrbp_1 \cpu.ex.r_wdata[13]$_DFFE_PP_  (.CLK(clknet_leaf_308_clk),
    .RESET_B(net1924),
    .D(_01043_),
    .Q_N(_14343_),
    .Q(\cpu.dcache.wdata[13] ));
 sg13g2_dfrbp_1 \cpu.ex.r_wdata[14]$_DFFE_PP_  (.CLK(clknet_leaf_303_clk),
    .RESET_B(net1925),
    .D(_01044_),
    .Q_N(_14342_),
    .Q(\cpu.dcache.wdata[14] ));
 sg13g2_dfrbp_1 \cpu.ex.r_wdata[15]$_DFFE_PP_  (.CLK(clknet_leaf_44_clk),
    .RESET_B(net1926),
    .D(_01045_),
    .Q_N(_14341_),
    .Q(\cpu.dcache.wdata[15] ));
 sg13g2_dfrbp_1 \cpu.ex.r_wdata[1]$_DFFE_PP_  (.CLK(clknet_leaf_56_clk),
    .RESET_B(net1927),
    .D(_01046_),
    .Q_N(_00168_),
    .Q(\cpu.dcache.wdata[1] ));
 sg13g2_dfrbp_1 \cpu.ex.r_wdata[2]$_DFFE_PP_  (.CLK(clknet_leaf_55_clk),
    .RESET_B(net1928),
    .D(_01047_),
    .Q_N(_00169_),
    .Q(\cpu.dcache.wdata[2] ));
 sg13g2_dfrbp_1 \cpu.ex.r_wdata[3]$_DFFE_PP_  (.CLK(clknet_leaf_55_clk),
    .RESET_B(net1929),
    .D(_01048_),
    .Q_N(_00271_),
    .Q(\cpu.dcache.wdata[3] ));
 sg13g2_dfrbp_1 \cpu.ex.r_wdata[4]$_DFFE_PP_  (.CLK(clknet_leaf_53_clk),
    .RESET_B(net1930),
    .D(_01049_),
    .Q_N(_00170_),
    .Q(\cpu.dcache.wdata[4] ));
 sg13g2_dfrbp_1 \cpu.ex.r_wdata[5]$_DFFE_PP_  (.CLK(clknet_leaf_55_clk),
    .RESET_B(net1931),
    .D(_01050_),
    .Q_N(_00171_),
    .Q(\cpu.dcache.wdata[5] ));
 sg13g2_dfrbp_1 \cpu.ex.r_wdata[6]$_DFFE_PP_  (.CLK(clknet_leaf_65_clk),
    .RESET_B(net1932),
    .D(_01051_),
    .Q_N(_00172_),
    .Q(\cpu.dcache.wdata[6] ));
 sg13g2_dfrbp_1 \cpu.ex.r_wdata[7]$_DFFE_PP_  (.CLK(clknet_leaf_65_clk),
    .RESET_B(net1933),
    .D(_01052_),
    .Q_N(_00265_),
    .Q(\cpu.dcache.wdata[7] ));
 sg13g2_dfrbp_1 \cpu.ex.r_wdata[8]$_DFFE_PP_  (.CLK(clknet_leaf_45_clk),
    .RESET_B(net1934),
    .D(_01053_),
    .Q_N(_14340_),
    .Q(\cpu.dcache.wdata[8] ));
 sg13g2_dfrbp_1 \cpu.ex.r_wdata[9]$_DFFE_PP_  (.CLK(clknet_leaf_43_clk),
    .RESET_B(net1935),
    .D(_01054_),
    .Q_N(_14339_),
    .Q(\cpu.dcache.wdata[9] ));
 sg13g2_dfrbp_1 \cpu.ex.r_wmask[0]$_SDFFE_PP0P_  (.CLK(clknet_leaf_46_clk),
    .RESET_B(net1936),
    .D(_01055_),
    .Q_N(_14338_),
    .Q(\cpu.ex.r_wmask[0] ));
 sg13g2_dfrbp_1 \cpu.ex.r_wmask[1]$_SDFFE_PP0P_  (.CLK(clknet_leaf_46_clk),
    .RESET_B(net1937),
    .D(_01056_),
    .Q_N(_14337_),
    .Q(\cpu.ex.r_wmask[1] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_fault_address[0]$_DFFE_PP_  (.CLK(clknet_leaf_259_clk),
    .RESET_B(net1938),
    .D(_01057_),
    .Q_N(_00272_),
    .Q(\cpu.ex.mmu_read[12] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_fault_address[1]$_DFFE_PP_  (.CLK(clknet_leaf_261_clk),
    .RESET_B(net1939),
    .D(_01058_),
    .Q_N(_14336_),
    .Q(\cpu.ex.mmu_read[13] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_fault_address[2]$_DFFE_PP_  (.CLK(clknet_leaf_256_clk),
    .RESET_B(net1940),
    .D(_01059_),
    .Q_N(_00178_),
    .Q(\cpu.ex.mmu_read[14] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_fault_address[3]$_DFFE_PP_  (.CLK(clknet_leaf_260_clk),
    .RESET_B(net1941),
    .D(_01060_),
    .Q_N(_14335_),
    .Q(\cpu.ex.mmu_read[15] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_fault_ins$_SDFFE_PN0P_  (.CLK(clknet_leaf_260_clk),
    .RESET_B(net1942),
    .D(_01061_),
    .Q_N(_00239_),
    .Q(\cpu.ex.mmu_read[3] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_fault_sup$_SDFFE_PN0P_  (.CLK(clknet_leaf_260_clk),
    .RESET_B(net1943),
    .D(_01062_),
    .Q_N(_14334_),
    .Q(\cpu.ex.mmu_read[2] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_fault_type$_SDFFE_PN0P_  (.CLK(clknet_leaf_176_clk),
    .RESET_B(net1944),
    .D(_01063_),
    .Q_N(_14333_),
    .Q(\cpu.ex.mmu_read[1] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_valid_d[0]$_SDFFE_PN0P_  (.CLK(clknet_leaf_252_clk),
    .RESET_B(net1945),
    .D(_01064_),
    .Q_N(_14332_),
    .Q(\cpu.genblk1.mmu.r_valid_d[0] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_valid_d[10]$_SDFFE_PN0P_  (.CLK(clknet_leaf_250_clk),
    .RESET_B(net1946),
    .D(_01065_),
    .Q_N(_14331_),
    .Q(\cpu.genblk1.mmu.r_valid_d[10] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_valid_d[11]$_SDFFE_PN0P_  (.CLK(clknet_leaf_252_clk),
    .RESET_B(net1947),
    .D(_01066_),
    .Q_N(_14330_),
    .Q(\cpu.genblk1.mmu.r_valid_d[11] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_valid_d[12]$_SDFFE_PN0P_  (.CLK(clknet_leaf_250_clk),
    .RESET_B(net1948),
    .D(_01067_),
    .Q_N(_14329_),
    .Q(\cpu.genblk1.mmu.r_valid_d[12] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_valid_d[13]$_SDFFE_PN0P_  (.CLK(clknet_leaf_251_clk),
    .RESET_B(net1949),
    .D(_01068_),
    .Q_N(_14328_),
    .Q(\cpu.genblk1.mmu.r_valid_d[13] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_valid_d[14]$_SDFFE_PN0P_  (.CLK(clknet_leaf_250_clk),
    .RESET_B(net1950),
    .D(_01069_),
    .Q_N(_14327_),
    .Q(\cpu.genblk1.mmu.r_valid_d[14] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_valid_d[15]$_SDFFE_PN0P_  (.CLK(clknet_leaf_252_clk),
    .RESET_B(net1951),
    .D(_01070_),
    .Q_N(_14326_),
    .Q(\cpu.genblk1.mmu.r_valid_d[15] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_valid_d[16]$_SDFFE_PN0P_  (.CLK(clknet_leaf_250_clk),
    .RESET_B(net1952),
    .D(_01071_),
    .Q_N(_14325_),
    .Q(\cpu.genblk1.mmu.r_valid_d[16] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_valid_d[17]$_SDFFE_PN0P_  (.CLK(clknet_leaf_240_clk),
    .RESET_B(net1953),
    .D(_01072_),
    .Q_N(_14324_),
    .Q(\cpu.genblk1.mmu.r_valid_d[17] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_valid_d[18]$_SDFFE_PN0P_  (.CLK(clknet_leaf_241_clk),
    .RESET_B(net1954),
    .D(_01073_),
    .Q_N(_14323_),
    .Q(\cpu.genblk1.mmu.r_valid_d[18] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_valid_d[19]$_SDFFE_PN0P_  (.CLK(clknet_leaf_240_clk),
    .RESET_B(net1955),
    .D(_01074_),
    .Q_N(_14322_),
    .Q(\cpu.genblk1.mmu.r_valid_d[19] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_valid_d[1]$_SDFFE_PN0P_  (.CLK(clknet_leaf_251_clk),
    .RESET_B(net1956),
    .D(_01075_),
    .Q_N(_14321_),
    .Q(\cpu.genblk1.mmu.r_valid_d[1] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_valid_d[20]$_SDFFE_PN0P_  (.CLK(clknet_leaf_241_clk),
    .RESET_B(net1957),
    .D(_01076_),
    .Q_N(_14320_),
    .Q(\cpu.genblk1.mmu.r_valid_d[20] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_valid_d[21]$_SDFFE_PN0P_  (.CLK(clknet_leaf_239_clk),
    .RESET_B(net1958),
    .D(_01077_),
    .Q_N(_14319_),
    .Q(\cpu.genblk1.mmu.r_valid_d[21] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_valid_d[22]$_SDFFE_PN0P_  (.CLK(clknet_leaf_241_clk),
    .RESET_B(net1959),
    .D(_01078_),
    .Q_N(_14318_),
    .Q(\cpu.genblk1.mmu.r_valid_d[22] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_valid_d[23]$_SDFFE_PN0P_  (.CLK(clknet_leaf_241_clk),
    .RESET_B(net1960),
    .D(_01079_),
    .Q_N(_14317_),
    .Q(\cpu.genblk1.mmu.r_valid_d[23] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_valid_d[24]$_SDFFE_PN0P_  (.CLK(clknet_leaf_242_clk),
    .RESET_B(net1961),
    .D(_01080_),
    .Q_N(_14316_),
    .Q(\cpu.genblk1.mmu.r_valid_d[24] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_valid_d[25]$_SDFFE_PN0P_  (.CLK(clknet_leaf_239_clk),
    .RESET_B(net1962),
    .D(_01081_),
    .Q_N(_14315_),
    .Q(\cpu.genblk1.mmu.r_valid_d[25] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_valid_d[26]$_SDFFE_PN0P_  (.CLK(clknet_leaf_247_clk),
    .RESET_B(net1963),
    .D(_01082_),
    .Q_N(_14314_),
    .Q(\cpu.genblk1.mmu.r_valid_d[26] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_valid_d[27]$_SDFFE_PN0P_  (.CLK(clknet_leaf_240_clk),
    .RESET_B(net1964),
    .D(_01083_),
    .Q_N(_14313_),
    .Q(\cpu.genblk1.mmu.r_valid_d[27] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_valid_d[28]$_SDFFE_PN0P_  (.CLK(clknet_leaf_240_clk),
    .RESET_B(net1965),
    .D(_01084_),
    .Q_N(_14312_),
    .Q(\cpu.genblk1.mmu.r_valid_d[28] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_valid_d[29]$_SDFFE_PN0P_  (.CLK(clknet_leaf_240_clk),
    .RESET_B(net1966),
    .D(_01085_),
    .Q_N(_14311_),
    .Q(\cpu.genblk1.mmu.r_valid_d[29] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_valid_d[2]$_SDFFE_PN0P_  (.CLK(clknet_leaf_256_clk),
    .RESET_B(net1967),
    .D(_01086_),
    .Q_N(_14310_),
    .Q(\cpu.genblk1.mmu.r_valid_d[2] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_valid_d[30]$_SDFFE_PN0P_  (.CLK(clknet_leaf_251_clk),
    .RESET_B(net1968),
    .D(_01087_),
    .Q_N(_14309_),
    .Q(\cpu.genblk1.mmu.r_valid_d[30] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_valid_d[31]$_SDFFE_PN0P_  (.CLK(clknet_leaf_240_clk),
    .RESET_B(net1969),
    .D(_01088_),
    .Q_N(_14308_),
    .Q(\cpu.genblk1.mmu.r_valid_d[31] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_valid_d[3]$_SDFFE_PN0P_  (.CLK(clknet_leaf_251_clk),
    .RESET_B(net1970),
    .D(_01089_),
    .Q_N(_14307_),
    .Q(\cpu.genblk1.mmu.r_valid_d[3] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_valid_d[4]$_SDFFE_PN0P_  (.CLK(clknet_leaf_256_clk),
    .RESET_B(net1971),
    .D(_01090_),
    .Q_N(_14306_),
    .Q(\cpu.genblk1.mmu.r_valid_d[4] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_valid_d[5]$_SDFFE_PN0P_  (.CLK(clknet_leaf_255_clk),
    .RESET_B(net1972),
    .D(_01091_),
    .Q_N(_14305_),
    .Q(\cpu.genblk1.mmu.r_valid_d[5] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_valid_d[6]$_SDFFE_PN0P_  (.CLK(clknet_leaf_256_clk),
    .RESET_B(net1973),
    .D(_01092_),
    .Q_N(_14304_),
    .Q(\cpu.genblk1.mmu.r_valid_d[6] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_valid_d[7]$_SDFFE_PN0P_  (.CLK(clknet_leaf_255_clk),
    .RESET_B(net1974),
    .D(_01093_),
    .Q_N(_14303_),
    .Q(\cpu.genblk1.mmu.r_valid_d[7] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_valid_d[8]$_SDFFE_PN0P_  (.CLK(clknet_leaf_256_clk),
    .RESET_B(net1975),
    .D(_01094_),
    .Q_N(_14302_),
    .Q(\cpu.genblk1.mmu.r_valid_d[8] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_valid_d[9]$_SDFFE_PN0P_  (.CLK(clknet_leaf_252_clk),
    .RESET_B(net1976),
    .D(_01095_),
    .Q_N(_14301_),
    .Q(\cpu.genblk1.mmu.r_valid_d[9] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_valid_i[0]$_SDFFE_PN0P_  (.CLK(clknet_leaf_256_clk),
    .RESET_B(net1977),
    .D(_01096_),
    .Q_N(_14300_),
    .Q(\cpu.genblk1.mmu.r_valid_i[0] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_valid_i[10]$_SDFFE_PN0P_  (.CLK(clknet_leaf_250_clk),
    .RESET_B(net1978),
    .D(_01097_),
    .Q_N(_14299_),
    .Q(\cpu.genblk1.mmu.r_valid_i[10] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_valid_i[11]$_SDFFE_PN0P_  (.CLK(clknet_leaf_247_clk),
    .RESET_B(net1979),
    .D(_01098_),
    .Q_N(_14298_),
    .Q(\cpu.genblk1.mmu.r_valid_i[11] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_valid_i[12]$_SDFFE_PN0P_  (.CLK(clknet_leaf_251_clk),
    .RESET_B(net1980),
    .D(_01099_),
    .Q_N(_14297_),
    .Q(\cpu.genblk1.mmu.r_valid_i[12] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_valid_i[13]$_SDFFE_PN0P_  (.CLK(clknet_leaf_247_clk),
    .RESET_B(net1981),
    .D(_01100_),
    .Q_N(_14296_),
    .Q(\cpu.genblk1.mmu.r_valid_i[13] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_valid_i[14]$_SDFFE_PN0P_  (.CLK(clknet_leaf_251_clk),
    .RESET_B(net1982),
    .D(_01101_),
    .Q_N(_14295_),
    .Q(\cpu.genblk1.mmu.r_valid_i[14] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_valid_i[15]$_SDFFE_PN0P_  (.CLK(clknet_leaf_247_clk),
    .RESET_B(net1983),
    .D(_01102_),
    .Q_N(_14294_),
    .Q(\cpu.genblk1.mmu.r_valid_i[15] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_valid_i[16]$_SDFFE_PN0P_  (.CLK(clknet_leaf_246_clk),
    .RESET_B(net1984),
    .D(_01103_),
    .Q_N(_14293_),
    .Q(\cpu.genblk1.mmu.r_valid_i[16] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_valid_i[17]$_SDFFE_PN0P_  (.CLK(clknet_leaf_241_clk),
    .RESET_B(net1985),
    .D(_01104_),
    .Q_N(_14292_),
    .Q(\cpu.genblk1.mmu.r_valid_i[17] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_valid_i[18]$_SDFFE_PN0P_  (.CLK(clknet_leaf_241_clk),
    .RESET_B(net1986),
    .D(_01105_),
    .Q_N(_14291_),
    .Q(\cpu.genblk1.mmu.r_valid_i[18] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_valid_i[19]$_SDFFE_PN0P_  (.CLK(clknet_leaf_246_clk),
    .RESET_B(net1987),
    .D(_01106_),
    .Q_N(_14290_),
    .Q(\cpu.genblk1.mmu.r_valid_i[19] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_valid_i[1]$_SDFFE_PN0P_  (.CLK(clknet_leaf_247_clk),
    .RESET_B(net1988),
    .D(_01107_),
    .Q_N(_14289_),
    .Q(\cpu.genblk1.mmu.r_valid_i[1] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_valid_i[20]$_SDFFE_PN0P_  (.CLK(clknet_leaf_243_clk),
    .RESET_B(net1989),
    .D(_01108_),
    .Q_N(_14288_),
    .Q(\cpu.genblk1.mmu.r_valid_i[20] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_valid_i[21]$_SDFFE_PN0P_  (.CLK(clknet_leaf_242_clk),
    .RESET_B(net1990),
    .D(_01109_),
    .Q_N(_14287_),
    .Q(\cpu.genblk1.mmu.r_valid_i[21] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_valid_i[22]$_SDFFE_PN0P_  (.CLK(clknet_leaf_242_clk),
    .RESET_B(net1991),
    .D(_01110_),
    .Q_N(_14286_),
    .Q(\cpu.genblk1.mmu.r_valid_i[22] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_valid_i[23]$_SDFFE_PN0P_  (.CLK(clknet_leaf_242_clk),
    .RESET_B(net1992),
    .D(_01111_),
    .Q_N(_14285_),
    .Q(\cpu.genblk1.mmu.r_valid_i[23] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_valid_i[24]$_SDFFE_PN0P_  (.CLK(clknet_leaf_242_clk),
    .RESET_B(net1993),
    .D(_01112_),
    .Q_N(_14284_),
    .Q(\cpu.genblk1.mmu.r_valid_i[24] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_valid_i[25]$_SDFFE_PN0P_  (.CLK(clknet_leaf_242_clk),
    .RESET_B(net1994),
    .D(_01113_),
    .Q_N(_14283_),
    .Q(\cpu.genblk1.mmu.r_valid_i[25] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_valid_i[26]$_SDFFE_PN0P_  (.CLK(clknet_leaf_247_clk),
    .RESET_B(net1995),
    .D(_01114_),
    .Q_N(_14282_),
    .Q(\cpu.genblk1.mmu.r_valid_i[26] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_valid_i[27]$_SDFFE_PN0P_  (.CLK(clknet_leaf_242_clk),
    .RESET_B(net1996),
    .D(_01115_),
    .Q_N(_14281_),
    .Q(\cpu.genblk1.mmu.r_valid_i[27] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_valid_i[28]$_SDFFE_PN0P_  (.CLK(clknet_leaf_247_clk),
    .RESET_B(net1997),
    .D(_01116_),
    .Q_N(_14280_),
    .Q(\cpu.genblk1.mmu.r_valid_i[28] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_valid_i[29]$_SDFFE_PN0P_  (.CLK(clknet_leaf_242_clk),
    .RESET_B(net1998),
    .D(_01117_),
    .Q_N(_14279_),
    .Q(\cpu.genblk1.mmu.r_valid_i[29] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_valid_i[2]$_SDFFE_PN0P_  (.CLK(clknet_leaf_256_clk),
    .RESET_B(net1999),
    .D(_01118_),
    .Q_N(_14278_),
    .Q(\cpu.genblk1.mmu.r_valid_i[2] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_valid_i[30]$_SDFFE_PN0P_  (.CLK(clknet_leaf_241_clk),
    .RESET_B(net2000),
    .D(_01119_),
    .Q_N(_14277_),
    .Q(\cpu.genblk1.mmu.r_valid_i[30] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_valid_i[31]$_SDFFE_PN0P_  (.CLK(clknet_leaf_241_clk),
    .RESET_B(net2001),
    .D(_01120_),
    .Q_N(_14276_),
    .Q(\cpu.genblk1.mmu.r_valid_i[31] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_valid_i[3]$_SDFFE_PN0P_  (.CLK(clknet_leaf_250_clk),
    .RESET_B(net2002),
    .D(_01121_),
    .Q_N(_14275_),
    .Q(\cpu.genblk1.mmu.r_valid_i[3] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_valid_i[4]$_SDFFE_PN0P_  (.CLK(clknet_leaf_256_clk),
    .RESET_B(net2003),
    .D(_01122_),
    .Q_N(_14274_),
    .Q(\cpu.genblk1.mmu.r_valid_i[4] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_valid_i[5]$_SDFFE_PN0P_  (.CLK(clknet_leaf_250_clk),
    .RESET_B(net2004),
    .D(_01123_),
    .Q_N(_14273_),
    .Q(\cpu.genblk1.mmu.r_valid_i[5] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_valid_i[6]$_SDFFE_PN0P_  (.CLK(clknet_leaf_255_clk),
    .RESET_B(net2005),
    .D(_01124_),
    .Q_N(_14272_),
    .Q(\cpu.genblk1.mmu.r_valid_i[6] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_valid_i[7]$_SDFFE_PN0P_  (.CLK(clknet_leaf_250_clk),
    .RESET_B(net2006),
    .D(_01125_),
    .Q_N(_14271_),
    .Q(\cpu.genblk1.mmu.r_valid_i[7] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_valid_i[8]$_SDFFE_PN0P_  (.CLK(clknet_leaf_257_clk),
    .RESET_B(net2007),
    .D(_01126_),
    .Q_N(_14270_),
    .Q(\cpu.genblk1.mmu.r_valid_i[8] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_valid_i[9]$_SDFFE_PN0P_  (.CLK(clknet_leaf_251_clk),
    .RESET_B(net2008),
    .D(_01127_),
    .Q_N(_14269_),
    .Q(\cpu.genblk1.mmu.r_valid_i[9] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[0][0]$_DFFE_PP_  (.CLK(clknet_leaf_130_clk),
    .RESET_B(net2009),
    .D(_01128_),
    .Q_N(_14268_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[0][0] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[0][10]$_DFFE_PP_  (.CLK(clknet_leaf_185_clk),
    .RESET_B(net2010),
    .D(_01129_),
    .Q_N(_14267_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[0][10] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[0][11]$_DFFE_PP_  (.CLK(clknet_leaf_171_clk),
    .RESET_B(net2011),
    .D(_01130_),
    .Q_N(_14266_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[0][11] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[0][1]$_DFFE_PP_  (.CLK(clknet_leaf_130_clk),
    .RESET_B(net2012),
    .D(_01131_),
    .Q_N(_14265_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[0][1] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[0][2]$_DFFE_PP_  (.CLK(clknet_leaf_169_clk),
    .RESET_B(net2013),
    .D(_01132_),
    .Q_N(_14264_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[0][2] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[0][3]$_DFFE_PP_  (.CLK(clknet_leaf_169_clk),
    .RESET_B(net2014),
    .D(_01133_),
    .Q_N(_14263_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[0][3] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[0][4]$_DFFE_PP_  (.CLK(clknet_leaf_150_clk),
    .RESET_B(net2015),
    .D(_01134_),
    .Q_N(_14262_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[0][4] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[0][5]$_DFFE_PP_  (.CLK(clknet_leaf_130_clk),
    .RESET_B(net2016),
    .D(_01135_),
    .Q_N(_14261_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[0][5] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[0][6]$_DFFE_PP_  (.CLK(clknet_leaf_229_clk),
    .RESET_B(net2017),
    .D(_01136_),
    .Q_N(_14260_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[0][6] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[0][7]$_DFFE_PP_  (.CLK(clknet_leaf_230_clk),
    .RESET_B(net2018),
    .D(_01137_),
    .Q_N(_14259_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[0][7] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[0][8]$_DFFE_PP_  (.CLK(clknet_leaf_232_clk),
    .RESET_B(net2019),
    .D(_01138_),
    .Q_N(_14258_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[0][8] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[0][9]$_DFFE_PP_  (.CLK(clknet_leaf_232_clk),
    .RESET_B(net2020),
    .D(_01139_),
    .Q_N(_14257_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[0][9] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[10][0]$_DFFE_PP_  (.CLK(clknet_leaf_136_clk),
    .RESET_B(net2021),
    .D(_01140_),
    .Q_N(_14256_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[10][0] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[10][10]$_DFFE_PP_  (.CLK(clknet_leaf_184_clk),
    .RESET_B(net2022),
    .D(_01141_),
    .Q_N(_14255_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[10][10] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[10][11]$_DFFE_PP_  (.CLK(clknet_leaf_152_clk),
    .RESET_B(net2023),
    .D(_01142_),
    .Q_N(_14254_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[10][11] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[10][1]$_DFFE_PP_  (.CLK(clknet_leaf_133_clk),
    .RESET_B(net2024),
    .D(_01143_),
    .Q_N(_14253_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[10][1] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[10][2]$_DFFE_PP_  (.CLK(clknet_leaf_127_clk),
    .RESET_B(net2025),
    .D(_01144_),
    .Q_N(_14252_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[10][2] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[10][3]$_DFFE_PP_  (.CLK(clknet_leaf_129_clk),
    .RESET_B(net2026),
    .D(_01145_),
    .Q_N(_14251_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[10][3] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[10][4]$_DFFE_PP_  (.CLK(clknet_leaf_134_clk),
    .RESET_B(net2027),
    .D(_01146_),
    .Q_N(_14250_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[10][4] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[10][5]$_DFFE_PP_  (.CLK(clknet_leaf_133_clk),
    .RESET_B(net2028),
    .D(_01147_),
    .Q_N(_14249_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[10][5] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[10][6]$_DFFE_PP_  (.CLK(clknet_leaf_231_clk),
    .RESET_B(net2029),
    .D(_01148_),
    .Q_N(_14248_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[10][6] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[10][7]$_DFFE_PP_  (.CLK(clknet_leaf_231_clk),
    .RESET_B(net2030),
    .D(_01149_),
    .Q_N(_14247_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[10][7] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[10][8]$_DFFE_PP_  (.CLK(clknet_leaf_253_clk),
    .RESET_B(net2031),
    .D(_01150_),
    .Q_N(_14246_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[10][8] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[10][9]$_DFFE_PP_  (.CLK(clknet_leaf_254_clk),
    .RESET_B(net2032),
    .D(_01151_),
    .Q_N(_14245_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[10][9] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[11][0]$_DFFE_PP_  (.CLK(clknet_leaf_136_clk),
    .RESET_B(net2033),
    .D(_01152_),
    .Q_N(_14244_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[11][0] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[11][10]$_DFFE_PP_  (.CLK(clknet_leaf_184_clk),
    .RESET_B(net2034),
    .D(_01153_),
    .Q_N(_14243_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[11][10] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[11][11]$_DFFE_PP_  (.CLK(clknet_leaf_152_clk),
    .RESET_B(net2035),
    .D(_01154_),
    .Q_N(_14242_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[11][11] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[11][1]$_DFFE_PP_  (.CLK(clknet_leaf_135_clk),
    .RESET_B(net2036),
    .D(_01155_),
    .Q_N(_14241_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[11][1] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[11][2]$_DFFE_PP_  (.CLK(clknet_leaf_134_clk),
    .RESET_B(net2037),
    .D(_01156_),
    .Q_N(_14240_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[11][2] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[11][3]$_DFFE_PP_  (.CLK(clknet_leaf_130_clk),
    .RESET_B(net2038),
    .D(_01157_),
    .Q_N(_14239_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[11][3] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[11][4]$_DFFE_PP_  (.CLK(clknet_leaf_135_clk),
    .RESET_B(net2039),
    .D(_01158_),
    .Q_N(_14238_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[11][4] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[11][5]$_DFFE_PP_  (.CLK(clknet_leaf_133_clk),
    .RESET_B(net2040),
    .D(_01159_),
    .Q_N(_14237_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[11][5] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[11][6]$_DFFE_PP_  (.CLK(clknet_leaf_211_clk),
    .RESET_B(net2041),
    .D(_01160_),
    .Q_N(_14236_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[11][6] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[11][7]$_DFFE_PP_  (.CLK(clknet_leaf_231_clk),
    .RESET_B(net2042),
    .D(_01161_),
    .Q_N(_14235_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[11][7] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[11][8]$_DFFE_PP_  (.CLK(clknet_leaf_253_clk),
    .RESET_B(net2043),
    .D(_01162_),
    .Q_N(_14234_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[11][8] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[11][9]$_DFFE_PP_  (.CLK(clknet_leaf_254_clk),
    .RESET_B(net2044),
    .D(_01163_),
    .Q_N(_14233_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[11][9] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[12][0]$_DFFE_PP_  (.CLK(clknet_leaf_131_clk),
    .RESET_B(net2045),
    .D(_01164_),
    .Q_N(_14232_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[12][0] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[12][10]$_DFFE_PP_  (.CLK(clknet_leaf_184_clk),
    .RESET_B(net2046),
    .D(_01165_),
    .Q_N(_14231_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[12][10] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[12][11]$_DFFE_PP_  (.CLK(clknet_leaf_153_clk),
    .RESET_B(net2047),
    .D(_01166_),
    .Q_N(_14230_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[12][11] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[12][1]$_DFFE_PP_  (.CLK(clknet_leaf_132_clk),
    .RESET_B(net2048),
    .D(_01167_),
    .Q_N(_14229_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[12][1] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[12][2]$_DFFE_PP_  (.CLK(clknet_leaf_129_clk),
    .RESET_B(net2049),
    .D(_01168_),
    .Q_N(_14228_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[12][2] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[12][3]$_DFFE_PP_  (.CLK(clknet_leaf_169_clk),
    .RESET_B(net2050),
    .D(_01169_),
    .Q_N(_14227_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[12][3] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[12][4]$_DFFE_PP_  (.CLK(clknet_leaf_152_clk),
    .RESET_B(net2051),
    .D(_01170_),
    .Q_N(_14226_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[12][4] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[12][5]$_DFFE_PP_  (.CLK(clknet_leaf_132_clk),
    .RESET_B(net2052),
    .D(_01171_),
    .Q_N(_14225_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[12][5] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[12][6]$_DFFE_PP_  (.CLK(clknet_leaf_211_clk),
    .RESET_B(net2053),
    .D(_01172_),
    .Q_N(_14224_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[12][6] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[12][7]$_DFFE_PP_  (.CLK(clknet_leaf_210_clk),
    .RESET_B(net2054),
    .D(_01173_),
    .Q_N(_14223_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[12][7] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[12][8]$_DFFE_PP_  (.CLK(clknet_leaf_254_clk),
    .RESET_B(net2055),
    .D(_01174_),
    .Q_N(_14222_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[12][8] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[12][9]$_DFFE_PP_  (.CLK(clknet_leaf_185_clk),
    .RESET_B(net2056),
    .D(_01175_),
    .Q_N(_14221_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[12][9] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[13][0]$_DFFE_PP_  (.CLK(clknet_leaf_131_clk),
    .RESET_B(net2057),
    .D(_01176_),
    .Q_N(_14220_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[13][0] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[13][10]$_DFFE_PP_  (.CLK(clknet_leaf_183_clk),
    .RESET_B(net2058),
    .D(_01177_),
    .Q_N(_14219_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[13][10] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[13][11]$_DFFE_PP_  (.CLK(clknet_leaf_153_clk),
    .RESET_B(net2059),
    .D(_01178_),
    .Q_N(_14218_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[13][11] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[13][1]$_DFFE_PP_  (.CLK(clknet_leaf_132_clk),
    .RESET_B(net2060),
    .D(_01179_),
    .Q_N(_14217_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[13][1] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[13][2]$_DFFE_PP_  (.CLK(clknet_leaf_151_clk),
    .RESET_B(net2061),
    .D(_01180_),
    .Q_N(_14216_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[13][2] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[13][3]$_DFFE_PP_  (.CLK(clknet_leaf_169_clk),
    .RESET_B(net2062),
    .D(_01181_),
    .Q_N(_14215_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[13][3] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[13][4]$_DFFE_PP_  (.CLK(clknet_leaf_150_clk),
    .RESET_B(net2063),
    .D(_01182_),
    .Q_N(_14214_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[13][4] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[13][5]$_DFFE_PP_  (.CLK(clknet_leaf_132_clk),
    .RESET_B(net2064),
    .D(_01183_),
    .Q_N(_14213_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[13][5] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[13][6]$_DFFE_PP_  (.CLK(clknet_leaf_211_clk),
    .RESET_B(net2065),
    .D(_01184_),
    .Q_N(_14212_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[13][6] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[13][7]$_DFFE_PP_  (.CLK(clknet_leaf_210_clk),
    .RESET_B(net2066),
    .D(_01185_),
    .Q_N(_14211_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[13][7] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[13][8]$_DFFE_PP_  (.CLK(clknet_leaf_183_clk),
    .RESET_B(net2067),
    .D(_01186_),
    .Q_N(_14210_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[13][8] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[13][9]$_DFFE_PP_  (.CLK(clknet_leaf_185_clk),
    .RESET_B(net2068),
    .D(_01187_),
    .Q_N(_14209_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[13][9] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[14][0]$_DFFE_PP_  (.CLK(clknet_leaf_131_clk),
    .RESET_B(net2069),
    .D(_01188_),
    .Q_N(_14208_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[14][0] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[14][10]$_DFFE_PP_  (.CLK(clknet_leaf_183_clk),
    .RESET_B(net2070),
    .D(_01189_),
    .Q_N(_14207_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[14][10] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[14][11]$_DFFE_PP_  (.CLK(clknet_leaf_151_clk),
    .RESET_B(net2071),
    .D(_01190_),
    .Q_N(_14206_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[14][11] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[14][1]$_DFFE_PP_  (.CLK(clknet_leaf_132_clk),
    .RESET_B(net2072),
    .D(_01191_),
    .Q_N(_14205_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[14][1] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[14][2]$_DFFE_PP_  (.CLK(clknet_leaf_151_clk),
    .RESET_B(net2073),
    .D(_01192_),
    .Q_N(_14204_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[14][2] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[14][3]$_DFFE_PP_  (.CLK(clknet_leaf_169_clk),
    .RESET_B(net2074),
    .D(_01193_),
    .Q_N(_14203_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[14][3] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[14][4]$_DFFE_PP_  (.CLK(clknet_leaf_151_clk),
    .RESET_B(net2075),
    .D(_01194_),
    .Q_N(_14202_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[14][4] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[14][5]$_DFFE_PP_  (.CLK(clknet_leaf_132_clk),
    .RESET_B(net2076),
    .D(_01195_),
    .Q_N(_14201_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[14][5] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[14][6]$_DFFE_PP_  (.CLK(clknet_leaf_211_clk),
    .RESET_B(net2077),
    .D(_01196_),
    .Q_N(_14200_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[14][6] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[14][7]$_DFFE_PP_  (.CLK(clknet_leaf_231_clk),
    .RESET_B(net2078),
    .D(_01197_),
    .Q_N(_14199_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[14][7] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[14][8]$_DFFE_PP_  (.CLK(clknet_leaf_185_clk),
    .RESET_B(net2079),
    .D(_01198_),
    .Q_N(_14198_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[14][8] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[14][9]$_DFFE_PP_  (.CLK(clknet_leaf_185_clk),
    .RESET_B(net2080),
    .D(_01199_),
    .Q_N(_14197_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[14][9] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[15][0]$_DFFE_PP_  (.CLK(clknet_leaf_131_clk),
    .RESET_B(net2081),
    .D(_01200_),
    .Q_N(_14196_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[15][0] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[15][10]$_DFFE_PP_  (.CLK(clknet_leaf_184_clk),
    .RESET_B(net2082),
    .D(_01201_),
    .Q_N(_14195_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[15][10] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[15][11]$_DFFE_PP_  (.CLK(clknet_leaf_153_clk),
    .RESET_B(net2083),
    .D(_01202_),
    .Q_N(_14194_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[15][11] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[15][1]$_DFFE_PP_  (.CLK(clknet_leaf_132_clk),
    .RESET_B(net2084),
    .D(_01203_),
    .Q_N(_14193_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[15][1] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[15][2]$_DFFE_PP_  (.CLK(clknet_leaf_129_clk),
    .RESET_B(net2085),
    .D(_01204_),
    .Q_N(_14192_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[15][2] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[15][3]$_DFFE_PP_  (.CLK(clknet_leaf_169_clk),
    .RESET_B(net2086),
    .D(_01205_),
    .Q_N(_14191_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[15][3] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[15][4]$_DFFE_PP_  (.CLK(clknet_leaf_151_clk),
    .RESET_B(net2087),
    .D(_01206_),
    .Q_N(_14190_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[15][4] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[15][5]$_DFFE_PP_  (.CLK(clknet_leaf_132_clk),
    .RESET_B(net2088),
    .D(_01207_),
    .Q_N(_14189_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[15][5] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[15][6]$_DFFE_PP_  (.CLK(clknet_leaf_211_clk),
    .RESET_B(net2089),
    .D(_01208_),
    .Q_N(_14188_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[15][6] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[15][7]$_DFFE_PP_  (.CLK(clknet_leaf_230_clk),
    .RESET_B(net2090),
    .D(_01209_),
    .Q_N(_14187_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[15][7] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[15][8]$_DFFE_PP_  (.CLK(clknet_leaf_254_clk),
    .RESET_B(net2091),
    .D(_01210_),
    .Q_N(_14186_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[15][8] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[15][9]$_DFFE_PP_  (.CLK(clknet_leaf_184_clk),
    .RESET_B(net2092),
    .D(_01211_),
    .Q_N(_14185_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[15][9] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[16][0]$_DFFE_PP_  (.CLK(clknet_leaf_167_clk),
    .RESET_B(net2093),
    .D(_01212_),
    .Q_N(_14184_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[16][0] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[16][10]$_DFFE_PP_  (.CLK(clknet_leaf_186_clk),
    .RESET_B(net2094),
    .D(_01213_),
    .Q_N(_14183_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[16][10] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[16][11]$_DFFE_PP_  (.CLK(clknet_leaf_166_clk),
    .RESET_B(net2095),
    .D(_01214_),
    .Q_N(_14182_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[16][11] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[16][1]$_DFFE_PP_  (.CLK(clknet_leaf_223_clk),
    .RESET_B(net2096),
    .D(_01215_),
    .Q_N(_14181_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[16][1] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[16][2]$_DFFE_PP_  (.CLK(clknet_leaf_169_clk),
    .RESET_B(net2097),
    .D(_01216_),
    .Q_N(_14180_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[16][2] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[16][3]$_DFFE_PP_  (.CLK(clknet_leaf_170_clk),
    .RESET_B(net2098),
    .D(_01217_),
    .Q_N(_14179_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[16][3] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[16][4]$_DFFE_PP_  (.CLK(clknet_leaf_193_clk),
    .RESET_B(net2099),
    .D(_01218_),
    .Q_N(_14178_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[16][4] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[16][5]$_DFFE_PP_  (.CLK(clknet_leaf_168_clk),
    .RESET_B(net2100),
    .D(_01219_),
    .Q_N(_14177_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[16][5] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[16][6]$_DFFE_PP_  (.CLK(clknet_leaf_227_clk),
    .RESET_B(net2101),
    .D(_01220_),
    .Q_N(_14176_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[16][6] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[16][7]$_DFFE_PP_  (.CLK(clknet_leaf_230_clk),
    .RESET_B(net2102),
    .D(_01221_),
    .Q_N(_14175_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[16][7] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[16][8]$_DFFE_PP_  (.CLK(clknet_leaf_235_clk),
    .RESET_B(net2103),
    .D(_01222_),
    .Q_N(_14174_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[16][8] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[16][9]$_DFFE_PP_  (.CLK(clknet_leaf_227_clk),
    .RESET_B(net2104),
    .D(_01223_),
    .Q_N(_14173_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[16][9] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[17][0]$_DFFE_PP_  (.CLK(clknet_leaf_168_clk),
    .RESET_B(net2105),
    .D(_01224_),
    .Q_N(_14172_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[17][0] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[17][10]$_DFFE_PP_  (.CLK(clknet_leaf_186_clk),
    .RESET_B(net2106),
    .D(_01225_),
    .Q_N(_14171_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[17][10] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[17][11]$_DFFE_PP_  (.CLK(clknet_leaf_166_clk),
    .RESET_B(net2107),
    .D(_01226_),
    .Q_N(_14170_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[17][11] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[17][1]$_DFFE_PP_  (.CLK(clknet_leaf_222_clk),
    .RESET_B(net2108),
    .D(_01227_),
    .Q_N(_14169_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[17][1] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[17][2]$_DFFE_PP_  (.CLK(clknet_leaf_169_clk),
    .RESET_B(net2109),
    .D(_01228_),
    .Q_N(_14168_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[17][2] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[17][3]$_DFFE_PP_  (.CLK(clknet_leaf_170_clk),
    .RESET_B(net2110),
    .D(_01229_),
    .Q_N(_14167_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[17][3] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[17][4]$_DFFE_PP_  (.CLK(clknet_leaf_193_clk),
    .RESET_B(net2111),
    .D(_01230_),
    .Q_N(_14166_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[17][4] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[17][5]$_DFFE_PP_  (.CLK(clknet_leaf_168_clk),
    .RESET_B(net2112),
    .D(_01231_),
    .Q_N(_14165_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[17][5] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[17][6]$_DFFE_PP_  (.CLK(clknet_leaf_226_clk),
    .RESET_B(net2113),
    .D(_01232_),
    .Q_N(_14164_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[17][6] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[17][7]$_DFFE_PP_  (.CLK(clknet_leaf_230_clk),
    .RESET_B(net2114),
    .D(_01233_),
    .Q_N(_14163_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[17][7] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[17][8]$_DFFE_PP_  (.CLK(clknet_leaf_236_clk),
    .RESET_B(net2115),
    .D(_01234_),
    .Q_N(_14162_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[17][8] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[17][9]$_DFFE_PP_  (.CLK(clknet_leaf_226_clk),
    .RESET_B(net2116),
    .D(_01235_),
    .Q_N(_14161_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[17][9] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[18][0]$_DFFE_PP_  (.CLK(clknet_leaf_167_clk),
    .RESET_B(net2117),
    .D(_01236_),
    .Q_N(_14160_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[18][0] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[18][10]$_DFFE_PP_  (.CLK(clknet_leaf_186_clk),
    .RESET_B(net2118),
    .D(_01237_),
    .Q_N(_14159_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[18][10] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[18][11]$_DFFE_PP_  (.CLK(clknet_leaf_166_clk),
    .RESET_B(net2119),
    .D(_01238_),
    .Q_N(_14158_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[18][11] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[18][1]$_DFFE_PP_  (.CLK(clknet_leaf_223_clk),
    .RESET_B(net2120),
    .D(_01239_),
    .Q_N(_14157_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[18][1] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[18][2]$_DFFE_PP_  (.CLK(clknet_leaf_168_clk),
    .RESET_B(net2121),
    .D(_01240_),
    .Q_N(_14156_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[18][2] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[18][3]$_DFFE_PP_  (.CLK(clknet_leaf_168_clk),
    .RESET_B(net2122),
    .D(_01241_),
    .Q_N(_14155_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[18][3] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[18][4]$_DFFE_PP_  (.CLK(clknet_leaf_194_clk),
    .RESET_B(net2123),
    .D(_01242_),
    .Q_N(_14154_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[18][4] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[18][5]$_DFFE_PP_  (.CLK(clknet_leaf_192_clk),
    .RESET_B(net2124),
    .D(_01243_),
    .Q_N(_14153_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[18][5] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[18][6]$_DFFE_PP_  (.CLK(clknet_leaf_227_clk),
    .RESET_B(net2125),
    .D(_01244_),
    .Q_N(_14152_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[18][6] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[18][7]$_DFFE_PP_  (.CLK(clknet_leaf_229_clk),
    .RESET_B(net2126),
    .D(_01245_),
    .Q_N(_14151_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[18][7] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[18][8]$_DFFE_PP_  (.CLK(clknet_leaf_236_clk),
    .RESET_B(net2127),
    .D(_01246_),
    .Q_N(_14150_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[18][8] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[18][9]$_DFFE_PP_  (.CLK(clknet_leaf_227_clk),
    .RESET_B(net2128),
    .D(_01247_),
    .Q_N(_14149_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[18][9] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[19][0]$_DFFE_PP_  (.CLK(clknet_leaf_167_clk),
    .RESET_B(net2129),
    .D(_01248_),
    .Q_N(_14148_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[19][0] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[19][10]$_DFFE_PP_  (.CLK(clknet_leaf_210_clk),
    .RESET_B(net2130),
    .D(_01249_),
    .Q_N(_14147_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[19][10] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[19][11]$_DFFE_PP_  (.CLK(clknet_leaf_170_clk),
    .RESET_B(net2131),
    .D(_01250_),
    .Q_N(_14146_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[19][11] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[19][1]$_DFFE_PP_  (.CLK(clknet_leaf_222_clk),
    .RESET_B(net2132),
    .D(_01251_),
    .Q_N(_14145_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[19][1] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[19][2]$_DFFE_PP_  (.CLK(clknet_leaf_168_clk),
    .RESET_B(net2133),
    .D(_01252_),
    .Q_N(_14144_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[19][2] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[19][3]$_DFFE_PP_  (.CLK(clknet_leaf_170_clk),
    .RESET_B(net2134),
    .D(_01253_),
    .Q_N(_14143_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[19][3] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[19][4]$_DFFE_PP_  (.CLK(clknet_leaf_193_clk),
    .RESET_B(net2135),
    .D(_01254_),
    .Q_N(_14142_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[19][4] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[19][5]$_DFFE_PP_  (.CLK(clknet_leaf_192_clk),
    .RESET_B(net2136),
    .D(_01255_),
    .Q_N(_14141_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[19][5] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[19][6]$_DFFE_PP_  (.CLK(clknet_leaf_227_clk),
    .RESET_B(net2137),
    .D(_01256_),
    .Q_N(_14140_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[19][6] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[19][7]$_DFFE_PP_  (.CLK(clknet_leaf_227_clk),
    .RESET_B(net2138),
    .D(_01257_),
    .Q_N(_14139_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[19][7] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[19][8]$_DFFE_PP_  (.CLK(clknet_leaf_236_clk),
    .RESET_B(net2139),
    .D(_01258_),
    .Q_N(_14138_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[19][8] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[19][9]$_DFFE_PP_  (.CLK(clknet_leaf_226_clk),
    .RESET_B(net2140),
    .D(_01259_),
    .Q_N(_14137_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[19][9] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[1][0]$_DFFE_PP_  (.CLK(clknet_leaf_171_clk),
    .RESET_B(net2141),
    .D(_01260_),
    .Q_N(_14136_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[1][0] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[1][10]$_DFFE_PP_  (.CLK(clknet_leaf_186_clk),
    .RESET_B(net2142),
    .D(_01261_),
    .Q_N(_14135_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[1][10] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[1][11]$_DFFE_PP_  (.CLK(clknet_leaf_170_clk),
    .RESET_B(net2143),
    .D(_01262_),
    .Q_N(_14134_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[1][11] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[1][1]$_DFFE_PP_  (.CLK(clknet_leaf_131_clk),
    .RESET_B(net2144),
    .D(_01263_),
    .Q_N(_14133_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[1][1] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[1][2]$_DFFE_PP_  (.CLK(clknet_leaf_192_clk),
    .RESET_B(net2145),
    .D(_01264_),
    .Q_N(_14132_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[1][2] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[1][3]$_DFFE_PP_  (.CLK(clknet_leaf_171_clk),
    .RESET_B(net2146),
    .D(_01265_),
    .Q_N(_14131_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[1][3] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[1][4]$_DFFE_PP_  (.CLK(clknet_leaf_172_clk),
    .RESET_B(net2147),
    .D(_01266_),
    .Q_N(_14130_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[1][4] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[1][5]$_DFFE_PP_  (.CLK(clknet_leaf_129_clk),
    .RESET_B(net2148),
    .D(_01267_),
    .Q_N(_14129_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[1][5] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[1][6]$_DFFE_PP_  (.CLK(clknet_leaf_229_clk),
    .RESET_B(net2149),
    .D(_01268_),
    .Q_N(_14128_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[1][6] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[1][7]$_DFFE_PP_  (.CLK(clknet_leaf_230_clk),
    .RESET_B(net2150),
    .D(_01269_),
    .Q_N(_14127_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[1][7] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[1][8]$_DFFE_PP_  (.CLK(clknet_leaf_233_clk),
    .RESET_B(net2151),
    .D(_01270_),
    .Q_N(_14126_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[1][8] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[1][9]$_DFFE_PP_  (.CLK(clknet_leaf_233_clk),
    .RESET_B(net2152),
    .D(_01271_),
    .Q_N(_14125_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[1][9] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[20][0]$_DFFE_PP_  (.CLK(clknet_leaf_212_clk),
    .RESET_B(net2153),
    .D(_01272_),
    .Q_N(_14124_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[20][0] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[20][10]$_DFFE_PP_  (.CLK(clknet_leaf_213_clk),
    .RESET_B(net2154),
    .D(_01273_),
    .Q_N(_14123_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[20][10] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[20][11]$_DFFE_PP_  (.CLK(clknet_leaf_193_clk),
    .RESET_B(net2155),
    .D(_01274_),
    .Q_N(_14122_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[20][11] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[20][1]$_DFFE_PP_  (.CLK(clknet_leaf_222_clk),
    .RESET_B(net2156),
    .D(_01275_),
    .Q_N(_14121_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[20][1] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[20][2]$_DFFE_PP_  (.CLK(clknet_leaf_187_clk),
    .RESET_B(net2157),
    .D(_01276_),
    .Q_N(_14120_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[20][2] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[20][3]$_DFFE_PP_  (.CLK(clknet_leaf_192_clk),
    .RESET_B(net2158),
    .D(_01277_),
    .Q_N(_14119_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[20][3] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[20][4]$_DFFE_PP_  (.CLK(clknet_leaf_193_clk),
    .RESET_B(net2159),
    .D(_01278_),
    .Q_N(_14118_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[20][4] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[20][5]$_DFFE_PP_  (.CLK(clknet_leaf_192_clk),
    .RESET_B(net2160),
    .D(_01279_),
    .Q_N(_14117_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[20][5] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[20][6]$_DFFE_PP_  (.CLK(clknet_leaf_225_clk),
    .RESET_B(net2161),
    .D(_01280_),
    .Q_N(_14116_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[20][6] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[20][7]$_DFFE_PP_  (.CLK(clknet_leaf_224_clk),
    .RESET_B(net2162),
    .D(_01281_),
    .Q_N(_14115_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[20][7] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[20][8]$_DFFE_PP_  (.CLK(clknet_leaf_238_clk),
    .RESET_B(net2163),
    .D(_01282_),
    .Q_N(_14114_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[20][8] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[20][9]$_DFFE_PP_  (.CLK(clknet_leaf_237_clk),
    .RESET_B(net2164),
    .D(_01283_),
    .Q_N(_14113_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[20][9] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[21][0]$_DFFE_PP_  (.CLK(clknet_leaf_212_clk),
    .RESET_B(net2165),
    .D(_01284_),
    .Q_N(_14112_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[21][0] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[21][10]$_DFFE_PP_  (.CLK(clknet_leaf_211_clk),
    .RESET_B(net2166),
    .D(_01285_),
    .Q_N(_14111_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[21][10] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[21][11]$_DFFE_PP_  (.CLK(clknet_leaf_194_clk),
    .RESET_B(net2167),
    .D(_01286_),
    .Q_N(_14110_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[21][11] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[21][1]$_DFFE_PP_  (.CLK(clknet_leaf_228_clk),
    .RESET_B(net2168),
    .D(_01287_),
    .Q_N(_14109_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[21][1] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[21][2]$_DFFE_PP_  (.CLK(clknet_leaf_186_clk),
    .RESET_B(net2169),
    .D(_01288_),
    .Q_N(_14108_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[21][2] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[21][3]$_DFFE_PP_  (.CLK(clknet_leaf_192_clk),
    .RESET_B(net2170),
    .D(_01289_),
    .Q_N(_14107_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[21][3] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[21][4]$_DFFE_PP_  (.CLK(clknet_leaf_193_clk),
    .RESET_B(net2171),
    .D(_01290_),
    .Q_N(_14106_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[21][4] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[21][5]$_DFFE_PP_  (.CLK(clknet_leaf_191_clk),
    .RESET_B(net2172),
    .D(_01291_),
    .Q_N(_14105_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[21][5] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[21][6]$_DFFE_PP_  (.CLK(clknet_leaf_224_clk),
    .RESET_B(net2173),
    .D(_01292_),
    .Q_N(_14104_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[21][6] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[21][7]$_DFFE_PP_  (.CLK(clknet_leaf_225_clk),
    .RESET_B(net2174),
    .D(_01293_),
    .Q_N(_14103_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[21][7] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[21][8]$_DFFE_PP_  (.CLK(clknet_leaf_238_clk),
    .RESET_B(net2175),
    .D(_01294_),
    .Q_N(_14102_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[21][8] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[21][9]$_DFFE_PP_  (.CLK(clknet_leaf_237_clk),
    .RESET_B(net2176),
    .D(_01295_),
    .Q_N(_14101_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[21][9] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[22][0]$_DFFE_PP_  (.CLK(clknet_leaf_213_clk),
    .RESET_B(net2177),
    .D(_01296_),
    .Q_N(_14100_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[22][0] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[22][10]$_DFFE_PP_  (.CLK(clknet_leaf_213_clk),
    .RESET_B(net2178),
    .D(_01297_),
    .Q_N(_14099_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[22][10] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[22][11]$_DFFE_PP_  (.CLK(clknet_leaf_193_clk),
    .RESET_B(net2179),
    .D(_01298_),
    .Q_N(_14098_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[22][11] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[22][1]$_DFFE_PP_  (.CLK(clknet_leaf_222_clk),
    .RESET_B(net2180),
    .D(_01299_),
    .Q_N(_14097_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[22][1] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[22][2]$_DFFE_PP_  (.CLK(clknet_leaf_187_clk),
    .RESET_B(net2181),
    .D(_01300_),
    .Q_N(_14096_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[22][2] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[22][3]$_DFFE_PP_  (.CLK(clknet_leaf_168_clk),
    .RESET_B(net2182),
    .D(_01301_),
    .Q_N(_14095_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[22][3] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[22][4]$_DFFE_PP_  (.CLK(clknet_leaf_167_clk),
    .RESET_B(net2183),
    .D(_01302_),
    .Q_N(_14094_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[22][4] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[22][5]$_DFFE_PP_  (.CLK(clknet_leaf_191_clk),
    .RESET_B(net2184),
    .D(_01303_),
    .Q_N(_14093_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[22][5] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[22][6]$_DFFE_PP_  (.CLK(clknet_leaf_225_clk),
    .RESET_B(net2185),
    .D(_01304_),
    .Q_N(_14092_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[22][6] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[22][7]$_DFFE_PP_  (.CLK(clknet_leaf_224_clk),
    .RESET_B(net2186),
    .D(_01305_),
    .Q_N(_14091_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[22][7] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[22][8]$_DFFE_PP_  (.CLK(clknet_leaf_237_clk),
    .RESET_B(net2187),
    .D(_01306_),
    .Q_N(_14090_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[22][8] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[22][9]$_DFFE_PP_  (.CLK(clknet_leaf_225_clk),
    .RESET_B(net2188),
    .D(_01307_),
    .Q_N(_14089_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[22][9] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[23][0]$_DFFE_PP_  (.CLK(clknet_leaf_212_clk),
    .RESET_B(net2189),
    .D(_01308_),
    .Q_N(_14088_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[23][0] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[23][10]$_DFFE_PP_  (.CLK(clknet_leaf_213_clk),
    .RESET_B(net2190),
    .D(_01309_),
    .Q_N(_14087_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[23][10] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[23][11]$_DFFE_PP_  (.CLK(clknet_leaf_194_clk),
    .RESET_B(net2191),
    .D(_01310_),
    .Q_N(_14086_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[23][11] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[23][1]$_DFFE_PP_  (.CLK(clknet_leaf_223_clk),
    .RESET_B(net2192),
    .D(_01311_),
    .Q_N(_14085_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[23][1] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[23][2]$_DFFE_PP_  (.CLK(clknet_leaf_187_clk),
    .RESET_B(net2193),
    .D(_01312_),
    .Q_N(_14084_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[23][2] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[23][3]$_DFFE_PP_  (.CLK(clknet_leaf_168_clk),
    .RESET_B(net2194),
    .D(_01313_),
    .Q_N(_14083_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[23][3] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[23][4]$_DFFE_PP_  (.CLK(clknet_leaf_193_clk),
    .RESET_B(net2195),
    .D(_01314_),
    .Q_N(_14082_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[23][4] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[23][5]$_DFFE_PP_  (.CLK(clknet_leaf_191_clk),
    .RESET_B(net2196),
    .D(_01315_),
    .Q_N(_14081_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[23][5] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[23][6]$_DFFE_PP_  (.CLK(clknet_leaf_224_clk),
    .RESET_B(net2197),
    .D(_01316_),
    .Q_N(_14080_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[23][6] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[23][7]$_DFFE_PP_  (.CLK(clknet_leaf_225_clk),
    .RESET_B(net2198),
    .D(_01317_),
    .Q_N(_14079_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[23][7] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[23][8]$_DFFE_PP_  (.CLK(clknet_leaf_237_clk),
    .RESET_B(net2199),
    .D(_01318_),
    .Q_N(_14078_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[23][8] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[23][9]$_DFFE_PP_  (.CLK(clknet_leaf_225_clk),
    .RESET_B(net2200),
    .D(_01319_),
    .Q_N(_14077_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[23][9] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[24][0]$_DFFE_PP_  (.CLK(clknet_leaf_189_clk),
    .RESET_B(net2201),
    .D(_01320_),
    .Q_N(_14076_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[24][0] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[24][10]$_DFFE_PP_  (.CLK(clknet_leaf_186_clk),
    .RESET_B(net2202),
    .D(_01321_),
    .Q_N(_14075_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[24][10] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[24][11]$_DFFE_PP_  (.CLK(clknet_leaf_189_clk),
    .RESET_B(net2203),
    .D(_01322_),
    .Q_N(_14074_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[24][11] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[24][1]$_DFFE_PP_  (.CLK(clknet_leaf_223_clk),
    .RESET_B(net2204),
    .D(_01323_),
    .Q_N(_14073_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[24][1] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[24][2]$_DFFE_PP_  (.CLK(clknet_leaf_184_clk),
    .RESET_B(net2205),
    .D(_01324_),
    .Q_N(_14072_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[24][2] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[24][3]$_DFFE_PP_  (.CLK(clknet_leaf_190_clk),
    .RESET_B(net2206),
    .D(_01325_),
    .Q_N(_14071_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[24][3] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[24][4]$_DFFE_PP_  (.CLK(clknet_leaf_190_clk),
    .RESET_B(net2207),
    .D(_01326_),
    .Q_N(_14070_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[24][4] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[24][5]$_DFFE_PP_  (.CLK(clknet_leaf_187_clk),
    .RESET_B(net2208),
    .D(_01327_),
    .Q_N(_14069_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[24][5] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[24][6]$_DFFE_PP_  (.CLK(clknet_leaf_224_clk),
    .RESET_B(net2209),
    .D(_01328_),
    .Q_N(_14068_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[24][6] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[24][7]$_DFFE_PP_  (.CLK(clknet_leaf_225_clk),
    .RESET_B(net2210),
    .D(_01329_),
    .Q_N(_14067_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[24][7] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[24][8]$_DFFE_PP_  (.CLK(clknet_leaf_238_clk),
    .RESET_B(net2211),
    .D(_01330_),
    .Q_N(_14066_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[24][8] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[24][9]$_DFFE_PP_  (.CLK(clknet_leaf_237_clk),
    .RESET_B(net2212),
    .D(_01331_),
    .Q_N(_14065_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[24][9] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[25][0]$_DFFE_PP_  (.CLK(clknet_leaf_208_clk),
    .RESET_B(net2213),
    .D(_01332_),
    .Q_N(_14064_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[25][0] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[25][10]$_DFFE_PP_  (.CLK(clknet_leaf_210_clk),
    .RESET_B(net2214),
    .D(_01333_),
    .Q_N(_14063_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[25][10] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[25][11]$_DFFE_PP_  (.CLK(clknet_leaf_189_clk),
    .RESET_B(net2215),
    .D(_01334_),
    .Q_N(_14062_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[25][11] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[25][1]$_DFFE_PP_  (.CLK(clknet_leaf_223_clk),
    .RESET_B(net2216),
    .D(_01335_),
    .Q_N(_14061_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[25][1] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[25][2]$_DFFE_PP_  (.CLK(clknet_leaf_190_clk),
    .RESET_B(net2217),
    .D(_01336_),
    .Q_N(_14060_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[25][2] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[25][3]$_DFFE_PP_  (.CLK(clknet_leaf_187_clk),
    .RESET_B(net2218),
    .D(_01337_),
    .Q_N(_14059_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[25][3] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[25][4]$_DFFE_PP_  (.CLK(clknet_leaf_190_clk),
    .RESET_B(net2219),
    .D(_01338_),
    .Q_N(_14058_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[25][4] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[25][5]$_DFFE_PP_  (.CLK(clknet_leaf_187_clk),
    .RESET_B(net2220),
    .D(_01339_),
    .Q_N(_14057_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[25][5] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[25][6]$_DFFE_PP_  (.CLK(clknet_leaf_224_clk),
    .RESET_B(net2221),
    .D(_01340_),
    .Q_N(_14056_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[25][6] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[25][7]$_DFFE_PP_  (.CLK(clknet_leaf_225_clk),
    .RESET_B(net2222),
    .D(_01341_),
    .Q_N(_14055_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[25][7] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[25][8]$_DFFE_PP_  (.CLK(clknet_leaf_238_clk),
    .RESET_B(net2223),
    .D(_01342_),
    .Q_N(_14054_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[25][8] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[25][9]$_DFFE_PP_  (.CLK(clknet_leaf_237_clk),
    .RESET_B(net2224),
    .D(_01343_),
    .Q_N(_14053_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[25][9] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[26][0]$_DFFE_PP_  (.CLK(clknet_leaf_208_clk),
    .RESET_B(net2225),
    .D(_01344_),
    .Q_N(_14052_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[26][0] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[26][10]$_DFFE_PP_  (.CLK(clknet_leaf_210_clk),
    .RESET_B(net2226),
    .D(_01345_),
    .Q_N(_14051_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[26][10] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[26][11]$_DFFE_PP_  (.CLK(clknet_leaf_195_clk),
    .RESET_B(net2227),
    .D(_01346_),
    .Q_N(_14050_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[26][11] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[26][1]$_DFFE_PP_  (.CLK(clknet_leaf_223_clk),
    .RESET_B(net2228),
    .D(_01347_),
    .Q_N(_14049_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[26][1] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[26][2]$_DFFE_PP_  (.CLK(clknet_leaf_190_clk),
    .RESET_B(net2229),
    .D(_01348_),
    .Q_N(_14048_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[26][2] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[26][3]$_DFFE_PP_  (.CLK(clknet_leaf_191_clk),
    .RESET_B(net2230),
    .D(_01349_),
    .Q_N(_14047_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[26][3] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[26][4]$_DFFE_PP_  (.CLK(clknet_leaf_188_clk),
    .RESET_B(net2231),
    .D(_01350_),
    .Q_N(_14046_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[26][4] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[26][5]$_DFFE_PP_  (.CLK(clknet_leaf_187_clk),
    .RESET_B(net2232),
    .D(_01351_),
    .Q_N(_14045_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[26][5] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[26][6]$_DFFE_PP_  (.CLK(clknet_leaf_224_clk),
    .RESET_B(net2233),
    .D(_01352_),
    .Q_N(_14044_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[26][6] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[26][7]$_DFFE_PP_  (.CLK(clknet_leaf_226_clk),
    .RESET_B(net2234),
    .D(_01353_),
    .Q_N(_14043_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[26][7] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[26][8]$_DFFE_PP_  (.CLK(clknet_leaf_238_clk),
    .RESET_B(net2235),
    .D(_01354_),
    .Q_N(_14042_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[26][8] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[26][9]$_DFFE_PP_  (.CLK(clknet_leaf_236_clk),
    .RESET_B(net2236),
    .D(_01355_),
    .Q_N(_14041_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[26][9] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[27][0]$_DFFE_PP_  (.CLK(clknet_leaf_209_clk),
    .RESET_B(net2237),
    .D(_01356_),
    .Q_N(_14040_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[27][0] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[27][10]$_DFFE_PP_  (.CLK(clknet_leaf_210_clk),
    .RESET_B(net2238),
    .D(_01357_),
    .Q_N(_14039_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[27][10] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[27][11]$_DFFE_PP_  (.CLK(clknet_leaf_195_clk),
    .RESET_B(net2239),
    .D(_01358_),
    .Q_N(_14038_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[27][11] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[27][1]$_DFFE_PP_  (.CLK(clknet_leaf_223_clk),
    .RESET_B(net2240),
    .D(_01359_),
    .Q_N(_14037_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[27][1] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[27][2]$_DFFE_PP_  (.CLK(clknet_leaf_191_clk),
    .RESET_B(net2241),
    .D(_01360_),
    .Q_N(_14036_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[27][2] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[27][3]$_DFFE_PP_  (.CLK(clknet_leaf_191_clk),
    .RESET_B(net2242),
    .D(_01361_),
    .Q_N(_14035_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[27][3] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[27][4]$_DFFE_PP_  (.CLK(clknet_leaf_190_clk),
    .RESET_B(net2243),
    .D(_01362_),
    .Q_N(_14034_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[27][4] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[27][5]$_DFFE_PP_  (.CLK(clknet_leaf_187_clk),
    .RESET_B(net2244),
    .D(_01363_),
    .Q_N(_14033_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[27][5] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[27][6]$_DFFE_PP_  (.CLK(clknet_leaf_224_clk),
    .RESET_B(net2245),
    .D(_01364_),
    .Q_N(_14032_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[27][6] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[27][7]$_DFFE_PP_  (.CLK(clknet_leaf_226_clk),
    .RESET_B(net2246),
    .D(_01365_),
    .Q_N(_14031_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[27][7] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[27][8]$_DFFE_PP_  (.CLK(clknet_leaf_236_clk),
    .RESET_B(net2247),
    .D(_01366_),
    .Q_N(_14030_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[27][8] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[27][9]$_DFFE_PP_  (.CLK(clknet_leaf_236_clk),
    .RESET_B(net2248),
    .D(_01367_),
    .Q_N(_14029_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[27][9] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[28][0]$_DFFE_PP_  (.CLK(clknet_leaf_212_clk),
    .RESET_B(net2249),
    .D(_01368_),
    .Q_N(_14028_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[28][0] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[28][10]$_DFFE_PP_  (.CLK(clknet_leaf_209_clk),
    .RESET_B(net2250),
    .D(_01369_),
    .Q_N(_14027_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[28][10] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[28][11]$_DFFE_PP_  (.CLK(clknet_leaf_190_clk),
    .RESET_B(net2251),
    .D(_01370_),
    .Q_N(_14026_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[28][11] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[28][1]$_DFFE_PP_  (.CLK(clknet_leaf_228_clk),
    .RESET_B(net2252),
    .D(_01371_),
    .Q_N(_14025_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[28][1] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[28][2]$_DFFE_PP_  (.CLK(clknet_leaf_183_clk),
    .RESET_B(net2253),
    .D(_01372_),
    .Q_N(_14024_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[28][2] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[28][3]$_DFFE_PP_  (.CLK(clknet_leaf_188_clk),
    .RESET_B(net2254),
    .D(_01373_),
    .Q_N(_14023_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[28][3] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[28][4]$_DFFE_PP_  (.CLK(clknet_leaf_188_clk),
    .RESET_B(net2255),
    .D(_01374_),
    .Q_N(_14022_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[28][4] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[28][5]$_DFFE_PP_  (.CLK(clknet_leaf_191_clk),
    .RESET_B(net2256),
    .D(_01375_),
    .Q_N(_14021_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[28][5] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[28][6]$_DFFE_PP_  (.CLK(clknet_leaf_227_clk),
    .RESET_B(net2257),
    .D(_01376_),
    .Q_N(_14020_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[28][6] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[28][7]$_DFFE_PP_  (.CLK(clknet_leaf_226_clk),
    .RESET_B(net2258),
    .D(_01377_),
    .Q_N(_14019_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[28][7] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[28][8]$_DFFE_PP_  (.CLK(clknet_leaf_235_clk),
    .RESET_B(net2259),
    .D(_01378_),
    .Q_N(_14018_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[28][8] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[28][9]$_DFFE_PP_  (.CLK(clknet_leaf_237_clk),
    .RESET_B(net2260),
    .D(_01379_),
    .Q_N(_14017_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[28][9] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[29][0]$_DFFE_PP_  (.CLK(clknet_leaf_208_clk),
    .RESET_B(net2261),
    .D(_01380_),
    .Q_N(_14016_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[29][0] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[29][10]$_DFFE_PP_  (.CLK(clknet_leaf_210_clk),
    .RESET_B(net2262),
    .D(_01381_),
    .Q_N(_14015_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[29][10] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[29][11]$_DFFE_PP_  (.CLK(clknet_leaf_189_clk),
    .RESET_B(net2263),
    .D(_01382_),
    .Q_N(_14014_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[29][11] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[29][1]$_DFFE_PP_  (.CLK(clknet_leaf_228_clk),
    .RESET_B(net2264),
    .D(_01383_),
    .Q_N(_14013_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[29][1] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[29][2]$_DFFE_PP_  (.CLK(clknet_leaf_183_clk),
    .RESET_B(net2265),
    .D(_01384_),
    .Q_N(_14012_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[29][2] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[29][3]$_DFFE_PP_  (.CLK(clknet_leaf_188_clk),
    .RESET_B(net2266),
    .D(_01385_),
    .Q_N(_14011_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[29][3] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[29][4]$_DFFE_PP_  (.CLK(clknet_leaf_188_clk),
    .RESET_B(net2267),
    .D(_01386_),
    .Q_N(_14010_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[29][4] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[29][5]$_DFFE_PP_  (.CLK(clknet_leaf_191_clk),
    .RESET_B(net2268),
    .D(_01387_),
    .Q_N(_14009_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[29][5] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[29][6]$_DFFE_PP_  (.CLK(clknet_leaf_228_clk),
    .RESET_B(net2269),
    .D(_01388_),
    .Q_N(_14008_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[29][6] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[29][7]$_DFFE_PP_  (.CLK(clknet_leaf_226_clk),
    .RESET_B(net2270),
    .D(_01389_),
    .Q_N(_14007_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[29][7] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[29][8]$_DFFE_PP_  (.CLK(clknet_leaf_235_clk),
    .RESET_B(net2271),
    .D(_01390_),
    .Q_N(_14006_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[29][8] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[29][9]$_DFFE_PP_  (.CLK(clknet_leaf_237_clk),
    .RESET_B(net2272),
    .D(_01391_),
    .Q_N(_14005_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[29][9] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[2][0]$_DFFE_PP_  (.CLK(clknet_leaf_149_clk),
    .RESET_B(net2273),
    .D(_01392_),
    .Q_N(_14004_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[2][0] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[2][10]$_DFFE_PP_  (.CLK(clknet_leaf_186_clk),
    .RESET_B(net2274),
    .D(_01393_),
    .Q_N(_14003_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[2][10] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[2][11]$_DFFE_PP_  (.CLK(clknet_leaf_170_clk),
    .RESET_B(net2275),
    .D(_01394_),
    .Q_N(_14002_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[2][11] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[2][1]$_DFFE_PP_  (.CLK(clknet_leaf_130_clk),
    .RESET_B(net2276),
    .D(_01395_),
    .Q_N(_14001_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[2][1] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[2][2]$_DFFE_PP_  (.CLK(clknet_leaf_181_clk),
    .RESET_B(net2277),
    .D(_01396_),
    .Q_N(_14000_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[2][2] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[2][3]$_DFFE_PP_  (.CLK(clknet_leaf_172_clk),
    .RESET_B(net2278),
    .D(_01397_),
    .Q_N(_13999_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[2][3] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[2][4]$_DFFE_PP_  (.CLK(clknet_leaf_171_clk),
    .RESET_B(net2279),
    .D(_01398_),
    .Q_N(_13998_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[2][4] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[2][5]$_DFFE_PP_  (.CLK(clknet_leaf_129_clk),
    .RESET_B(net2280),
    .D(_01399_),
    .Q_N(_13997_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[2][5] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[2][6]$_DFFE_PP_  (.CLK(clknet_leaf_229_clk),
    .RESET_B(net2281),
    .D(_01400_),
    .Q_N(_13996_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[2][6] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[2][7]$_DFFE_PP_  (.CLK(clknet_leaf_230_clk),
    .RESET_B(net2282),
    .D(_01401_),
    .Q_N(_13995_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[2][7] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[2][8]$_DFFE_PP_  (.CLK(clknet_leaf_233_clk),
    .RESET_B(net2283),
    .D(_01402_),
    .Q_N(_13994_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[2][8] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[2][9]$_DFFE_PP_  (.CLK(clknet_leaf_233_clk),
    .RESET_B(net2284),
    .D(_01403_),
    .Q_N(_13993_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[2][9] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[30][0]$_DFFE_PP_  (.CLK(clknet_leaf_210_clk),
    .RESET_B(net2285),
    .D(_01404_),
    .Q_N(_13992_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[30][0] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[30][10]$_DFFE_PP_  (.CLK(clknet_leaf_209_clk),
    .RESET_B(net2286),
    .D(_01405_),
    .Q_N(_13991_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[30][10] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[30][11]$_DFFE_PP_  (.CLK(clknet_leaf_189_clk),
    .RESET_B(net2287),
    .D(_01406_),
    .Q_N(_13990_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[30][11] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[30][1]$_DFFE_PP_  (.CLK(clknet_leaf_229_clk),
    .RESET_B(net2288),
    .D(_01407_),
    .Q_N(_13989_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[30][1] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[30][2]$_DFFE_PP_  (.CLK(clknet_leaf_183_clk),
    .RESET_B(net2289),
    .D(_01408_),
    .Q_N(_13988_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[30][2] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[30][3]$_DFFE_PP_  (.CLK(clknet_leaf_188_clk),
    .RESET_B(net2290),
    .D(_01409_),
    .Q_N(_13987_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[30][3] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[30][4]$_DFFE_PP_  (.CLK(clknet_leaf_208_clk),
    .RESET_B(net2291),
    .D(_01410_),
    .Q_N(_13986_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[30][4] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[30][5]$_DFFE_PP_  (.CLK(clknet_leaf_190_clk),
    .RESET_B(net2292),
    .D(_01411_),
    .Q_N(_13985_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[30][5] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[30][6]$_DFFE_PP_  (.CLK(clknet_leaf_228_clk),
    .RESET_B(net2293),
    .D(_01412_),
    .Q_N(_13984_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[30][6] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[30][7]$_DFFE_PP_  (.CLK(clknet_leaf_227_clk),
    .RESET_B(net2294),
    .D(_01413_),
    .Q_N(_13983_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[30][7] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[30][8]$_DFFE_PP_  (.CLK(clknet_leaf_235_clk),
    .RESET_B(net2295),
    .D(_01414_),
    .Q_N(_13982_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[30][8] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[30][9]$_DFFE_PP_  (.CLK(clknet_leaf_236_clk),
    .RESET_B(net2296),
    .D(_01415_),
    .Q_N(_13981_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[30][9] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[31][0]$_DFFE_PP_  (.CLK(clknet_leaf_209_clk),
    .RESET_B(net2297),
    .D(_01416_),
    .Q_N(_13980_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[31][0] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[31][10]$_DFFE_PP_  (.CLK(clknet_leaf_209_clk),
    .RESET_B(net2298),
    .D(_01417_),
    .Q_N(_13979_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[31][10] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[31][11]$_DFFE_PP_  (.CLK(clknet_leaf_194_clk),
    .RESET_B(net2299),
    .D(_01418_),
    .Q_N(_13978_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[31][11] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[31][1]$_DFFE_PP_  (.CLK(clknet_leaf_228_clk),
    .RESET_B(net2300),
    .D(_01419_),
    .Q_N(_13977_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[31][1] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[31][2]$_DFFE_PP_  (.CLK(clknet_leaf_183_clk),
    .RESET_B(net2301),
    .D(_01420_),
    .Q_N(_13976_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[31][2] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[31][3]$_DFFE_PP_  (.CLK(clknet_leaf_188_clk),
    .RESET_B(net2302),
    .D(_01421_),
    .Q_N(_13975_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[31][3] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[31][4]$_DFFE_PP_  (.CLK(clknet_leaf_188_clk),
    .RESET_B(net2303),
    .D(_01422_),
    .Q_N(_13974_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[31][4] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[31][5]$_DFFE_PP_  (.CLK(clknet_leaf_192_clk),
    .RESET_B(net2304),
    .D(_01423_),
    .Q_N(_13973_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[31][5] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[31][6]$_DFFE_PP_  (.CLK(clknet_leaf_223_clk),
    .RESET_B(net2305),
    .D(_01424_),
    .Q_N(_13972_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[31][6] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[31][7]$_DFFE_PP_  (.CLK(clknet_leaf_226_clk),
    .RESET_B(net2306),
    .D(_01425_),
    .Q_N(_13971_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[31][7] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[31][8]$_DFFE_PP_  (.CLK(clknet_leaf_235_clk),
    .RESET_B(net2307),
    .D(_01426_),
    .Q_N(_13970_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[31][8] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[31][9]$_DFFE_PP_  (.CLK(clknet_leaf_236_clk),
    .RESET_B(net2308),
    .D(_01427_),
    .Q_N(_13969_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[31][9] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[3][0]$_DFFE_PP_  (.CLK(clknet_leaf_150_clk),
    .RESET_B(net2309),
    .D(_01428_),
    .Q_N(_13968_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[3][0] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[3][10]$_DFFE_PP_  (.CLK(clknet_leaf_186_clk),
    .RESET_B(net2310),
    .D(_01429_),
    .Q_N(_13967_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[3][10] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[3][11]$_DFFE_PP_  (.CLK(clknet_leaf_171_clk),
    .RESET_B(net2311),
    .D(_01430_),
    .Q_N(_13966_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[3][11] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[3][1]$_DFFE_PP_  (.CLK(clknet_leaf_130_clk),
    .RESET_B(net2312),
    .D(_01431_),
    .Q_N(_13965_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[3][1] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[3][2]$_DFFE_PP_  (.CLK(clknet_leaf_192_clk),
    .RESET_B(net2313),
    .D(_01432_),
    .Q_N(_13964_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[3][2] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[3][3]$_DFFE_PP_  (.CLK(clknet_leaf_171_clk),
    .RESET_B(net2314),
    .D(_01433_),
    .Q_N(_13963_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[3][3] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[3][4]$_DFFE_PP_  (.CLK(clknet_leaf_150_clk),
    .RESET_B(net2315),
    .D(_01434_),
    .Q_N(_13962_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[3][4] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[3][5]$_DFFE_PP_  (.CLK(clknet_leaf_129_clk),
    .RESET_B(net2316),
    .D(_01435_),
    .Q_N(_13961_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[3][5] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[3][6]$_DFFE_PP_  (.CLK(clknet_leaf_229_clk),
    .RESET_B(net2317),
    .D(_01436_),
    .Q_N(_13960_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[3][6] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[3][7]$_DFFE_PP_  (.CLK(clknet_leaf_230_clk),
    .RESET_B(net2318),
    .D(_01437_),
    .Q_N(_13959_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[3][7] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[3][8]$_DFFE_PP_  (.CLK(clknet_leaf_232_clk),
    .RESET_B(net2319),
    .D(_01438_),
    .Q_N(_13958_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[3][8] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[3][9]$_DFFE_PP_  (.CLK(clknet_leaf_233_clk),
    .RESET_B(net2320),
    .D(_01439_),
    .Q_N(_13957_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[3][9] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[4][0]$_DFFE_PP_  (.CLK(clknet_leaf_135_clk),
    .RESET_B(net2321),
    .D(_01440_),
    .Q_N(_13956_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[4][0] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[4][10]$_DFFE_PP_  (.CLK(clknet_leaf_185_clk),
    .RESET_B(net2322),
    .D(_01441_),
    .Q_N(_13955_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[4][10] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[4][11]$_DFFE_PP_  (.CLK(clknet_leaf_149_clk),
    .RESET_B(net2323),
    .D(_01442_),
    .Q_N(_13954_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[4][11] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[4][1]$_DFFE_PP_  (.CLK(clknet_leaf_134_clk),
    .RESET_B(net2324),
    .D(_01443_),
    .Q_N(_13953_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[4][1] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[4][2]$_DFFE_PP_  (.CLK(clknet_leaf_182_clk),
    .RESET_B(net2325),
    .D(_01444_),
    .Q_N(_13952_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[4][2] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[4][3]$_DFFE_PP_  (.CLK(clknet_leaf_172_clk),
    .RESET_B(net2326),
    .D(_01445_),
    .Q_N(_13951_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[4][3] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[4][4]$_DFFE_PP_  (.CLK(clknet_leaf_151_clk),
    .RESET_B(net2327),
    .D(_01446_),
    .Q_N(_13950_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[4][4] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[4][5]$_DFFE_PP_  (.CLK(clknet_leaf_134_clk),
    .RESET_B(net2328),
    .D(_01447_),
    .Q_N(_13949_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[4][5] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[4][6]$_DFFE_PP_  (.CLK(clknet_leaf_211_clk),
    .RESET_B(net2329),
    .D(_01448_),
    .Q_N(_13948_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[4][6] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[4][7]$_DFFE_PP_  (.CLK(clknet_leaf_233_clk),
    .RESET_B(net2330),
    .D(_01449_),
    .Q_N(_13947_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[4][7] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[4][8]$_DFFE_PP_  (.CLK(clknet_leaf_233_clk),
    .RESET_B(net2331),
    .D(_01450_),
    .Q_N(_13946_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[4][8] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[4][9]$_DFFE_PP_  (.CLK(clknet_leaf_233_clk),
    .RESET_B(net2332),
    .D(_01451_),
    .Q_N(_13945_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[4][9] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[5][0]$_DFFE_PP_  (.CLK(clknet_leaf_135_clk),
    .RESET_B(net2333),
    .D(_01452_),
    .Q_N(_13944_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[5][0] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[5][10]$_DFFE_PP_  (.CLK(clknet_leaf_185_clk),
    .RESET_B(net2334),
    .D(_01453_),
    .Q_N(_13943_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[5][10] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[5][11]$_DFFE_PP_  (.CLK(clknet_leaf_149_clk),
    .RESET_B(net2335),
    .D(_01454_),
    .Q_N(_13942_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[5][11] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[5][1]$_DFFE_PP_  (.CLK(clknet_leaf_134_clk),
    .RESET_B(net2336),
    .D(_01455_),
    .Q_N(_13941_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[5][1] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[5][2]$_DFFE_PP_  (.CLK(clknet_leaf_182_clk),
    .RESET_B(net2337),
    .D(_01456_),
    .Q_N(_13940_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[5][2] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[5][3]$_DFFE_PP_  (.CLK(clknet_leaf_172_clk),
    .RESET_B(net2338),
    .D(_01457_),
    .Q_N(_13939_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[5][3] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[5][4]$_DFFE_PP_  (.CLK(clknet_leaf_151_clk),
    .RESET_B(net2339),
    .D(_01458_),
    .Q_N(_13938_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[5][4] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[5][5]$_DFFE_PP_  (.CLK(clknet_leaf_133_clk),
    .RESET_B(net2340),
    .D(_01459_),
    .Q_N(_13937_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[5][5] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[5][6]$_DFFE_PP_  (.CLK(clknet_leaf_229_clk),
    .RESET_B(net2341),
    .D(_01460_),
    .Q_N(_13936_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[5][6] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[5][7]$_DFFE_PP_  (.CLK(clknet_leaf_231_clk),
    .RESET_B(net2342),
    .D(_01461_),
    .Q_N(_13935_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[5][7] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[5][8]$_DFFE_PP_  (.CLK(clknet_leaf_234_clk),
    .RESET_B(net2343),
    .D(_01462_),
    .Q_N(_13934_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[5][8] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[5][9]$_DFFE_PP_  (.CLK(clknet_leaf_232_clk),
    .RESET_B(net2344),
    .D(_01463_),
    .Q_N(_13933_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[5][9] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[6][0]$_DFFE_PP_  (.CLK(clknet_leaf_136_clk),
    .RESET_B(net2345),
    .D(_01464_),
    .Q_N(_13932_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[6][0] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[6][10]$_DFFE_PP_  (.CLK(clknet_leaf_185_clk),
    .RESET_B(net2346),
    .D(_01465_),
    .Q_N(_13931_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[6][10] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[6][11]$_DFFE_PP_  (.CLK(clknet_leaf_130_clk),
    .RESET_B(net2347),
    .D(_01466_),
    .Q_N(_13930_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[6][11] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[6][1]$_DFFE_PP_  (.CLK(clknet_leaf_134_clk),
    .RESET_B(net2348),
    .D(_01467_),
    .Q_N(_13929_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[6][1] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[6][2]$_DFFE_PP_  (.CLK(clknet_leaf_182_clk),
    .RESET_B(net2349),
    .D(_01468_),
    .Q_N(_13928_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[6][2] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[6][3]$_DFFE_PP_  (.CLK(clknet_leaf_172_clk),
    .RESET_B(net2350),
    .D(_01469_),
    .Q_N(_13927_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[6][3] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[6][4]$_DFFE_PP_  (.CLK(clknet_leaf_151_clk),
    .RESET_B(net2351),
    .D(_01470_),
    .Q_N(_13926_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[6][4] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[6][5]$_DFFE_PP_  (.CLK(clknet_leaf_133_clk),
    .RESET_B(net2352),
    .D(_01471_),
    .Q_N(_13925_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[6][5] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[6][6]$_DFFE_PP_  (.CLK(clknet_leaf_213_clk),
    .RESET_B(net2353),
    .D(_01472_),
    .Q_N(_13924_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[6][6] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[6][7]$_DFFE_PP_  (.CLK(clknet_leaf_231_clk),
    .RESET_B(net2354),
    .D(_01473_),
    .Q_N(_13923_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[6][7] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[6][8]$_DFFE_PP_  (.CLK(clknet_leaf_253_clk),
    .RESET_B(net2355),
    .D(_01474_),
    .Q_N(_13922_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[6][8] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[6][9]$_DFFE_PP_  (.CLK(clknet_leaf_232_clk),
    .RESET_B(net2356),
    .D(_01475_),
    .Q_N(_13921_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[6][9] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[7][0]$_DFFE_PP_  (.CLK(clknet_leaf_136_clk),
    .RESET_B(net2357),
    .D(_01476_),
    .Q_N(_13920_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[7][0] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[7][10]$_DFFE_PP_  (.CLK(clknet_leaf_184_clk),
    .RESET_B(net2358),
    .D(_01477_),
    .Q_N(_13919_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[7][10] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[7][11]$_DFFE_PP_  (.CLK(clknet_leaf_149_clk),
    .RESET_B(net2359),
    .D(_01478_),
    .Q_N(_13918_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[7][11] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[7][1]$_DFFE_PP_  (.CLK(clknet_leaf_133_clk),
    .RESET_B(net2360),
    .D(_01479_),
    .Q_N(_13917_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[7][1] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[7][2]$_DFFE_PP_  (.CLK(clknet_leaf_182_clk),
    .RESET_B(net2361),
    .D(_01480_),
    .Q_N(_13916_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[7][2] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[7][3]$_DFFE_PP_  (.CLK(clknet_leaf_172_clk),
    .RESET_B(net2362),
    .D(_01481_),
    .Q_N(_13915_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[7][3] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[7][4]$_DFFE_PP_  (.CLK(clknet_leaf_150_clk),
    .RESET_B(net2363),
    .D(_01482_),
    .Q_N(_13914_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[7][4] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[7][5]$_DFFE_PP_  (.CLK(clknet_leaf_133_clk),
    .RESET_B(net2364),
    .D(_01483_),
    .Q_N(_13913_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[7][5] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[7][6]$_DFFE_PP_  (.CLK(clknet_leaf_229_clk),
    .RESET_B(net2365),
    .D(_01484_),
    .Q_N(_13912_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[7][6] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[7][7]$_DFFE_PP_  (.CLK(clknet_leaf_232_clk),
    .RESET_B(net2366),
    .D(_01485_),
    .Q_N(_13911_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[7][7] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[7][8]$_DFFE_PP_  (.CLK(clknet_leaf_232_clk),
    .RESET_B(net2367),
    .D(_01486_),
    .Q_N(_13910_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[7][8] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[7][9]$_DFFE_PP_  (.CLK(clknet_leaf_232_clk),
    .RESET_B(net2368),
    .D(_01487_),
    .Q_N(_13909_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[7][9] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[8][0]$_DFFE_PP_  (.CLK(clknet_leaf_135_clk),
    .RESET_B(net2369),
    .D(_01488_),
    .Q_N(_13908_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[8][0] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[8][10]$_DFFE_PP_  (.CLK(clknet_leaf_183_clk),
    .RESET_B(net2370),
    .D(_01489_),
    .Q_N(_13907_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[8][10] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[8][11]$_DFFE_PP_  (.CLK(clknet_leaf_150_clk),
    .RESET_B(net2371),
    .D(_01490_),
    .Q_N(_13906_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[8][11] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[8][1]$_DFFE_PP_  (.CLK(clknet_leaf_134_clk),
    .RESET_B(net2372),
    .D(_01491_),
    .Q_N(_13905_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[8][1] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[8][2]$_DFFE_PP_  (.CLK(clknet_leaf_127_clk),
    .RESET_B(net2373),
    .D(_01492_),
    .Q_N(_13904_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[8][2] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[8][3]$_DFFE_PP_  (.CLK(clknet_leaf_129_clk),
    .RESET_B(net2374),
    .D(_01493_),
    .Q_N(_13903_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[8][3] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[8][4]$_DFFE_PP_  (.CLK(clknet_leaf_134_clk),
    .RESET_B(net2375),
    .D(_01494_),
    .Q_N(_13902_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[8][4] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[8][5]$_DFFE_PP_  (.CLK(clknet_leaf_128_clk),
    .RESET_B(net2376),
    .D(_01495_),
    .Q_N(_13901_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[8][5] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[8][6]$_DFFE_PP_  (.CLK(clknet_leaf_230_clk),
    .RESET_B(net2377),
    .D(_01496_),
    .Q_N(_13900_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[8][6] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[8][7]$_DFFE_PP_  (.CLK(clknet_leaf_231_clk),
    .RESET_B(net2378),
    .D(_01497_),
    .Q_N(_13899_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[8][7] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[8][8]$_DFFE_PP_  (.CLK(clknet_leaf_253_clk),
    .RESET_B(net2379),
    .D(_01498_),
    .Q_N(_13898_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[8][8] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[8][9]$_DFFE_PP_  (.CLK(clknet_leaf_254_clk),
    .RESET_B(net2380),
    .D(_01499_),
    .Q_N(_13897_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[8][9] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[9][0]$_DFFE_PP_  (.CLK(clknet_leaf_131_clk),
    .RESET_B(net2381),
    .D(_01500_),
    .Q_N(_13896_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[9][0] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[9][10]$_DFFE_PP_  (.CLK(clknet_leaf_184_clk),
    .RESET_B(net2382),
    .D(_01501_),
    .Q_N(_13895_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[9][10] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[9][11]$_DFFE_PP_  (.CLK(clknet_leaf_152_clk),
    .RESET_B(net2383),
    .D(_01502_),
    .Q_N(_13894_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[9][11] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[9][1]$_DFFE_PP_  (.CLK(clknet_leaf_133_clk),
    .RESET_B(net2384),
    .D(_01503_),
    .Q_N(_13893_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[9][1] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[9][2]$_DFFE_PP_  (.CLK(clknet_leaf_128_clk),
    .RESET_B(net2385),
    .D(_01504_),
    .Q_N(_13892_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[9][2] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[9][3]$_DFFE_PP_  (.CLK(clknet_leaf_130_clk),
    .RESET_B(net2386),
    .D(_01505_),
    .Q_N(_13891_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[9][3] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[9][4]$_DFFE_PP_  (.CLK(clknet_leaf_135_clk),
    .RESET_B(net2387),
    .D(_01506_),
    .Q_N(_13890_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[9][4] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[9][5]$_DFFE_PP_  (.CLK(clknet_leaf_128_clk),
    .RESET_B(net2388),
    .D(_01507_),
    .Q_N(_13889_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[9][5] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[9][6]$_DFFE_PP_  (.CLK(clknet_leaf_211_clk),
    .RESET_B(net2389),
    .D(_01508_),
    .Q_N(_13888_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[9][6] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[9][7]$_DFFE_PP_  (.CLK(clknet_leaf_231_clk),
    .RESET_B(net2390),
    .D(_01509_),
    .Q_N(_13887_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[9][7] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[9][8]$_DFFE_PP_  (.CLK(clknet_leaf_253_clk),
    .RESET_B(net2391),
    .D(_01510_),
    .Q_N(_13886_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[9][8] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[9][9]$_DFFE_PP_  (.CLK(clknet_leaf_253_clk),
    .RESET_B(net2392),
    .D(_01511_),
    .Q_N(_13885_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[9][9] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[0][0]$_DFFE_PP_  (.CLK(clknet_leaf_279_clk),
    .RESET_B(net2393),
    .D(_01512_),
    .Q_N(_13884_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[0][0] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[0][10]$_DFFE_PP_  (.CLK(clknet_leaf_275_clk),
    .RESET_B(net2394),
    .D(_01513_),
    .Q_N(_13883_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[0][10] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[0][11]$_DFFE_PP_  (.CLK(clknet_leaf_281_clk),
    .RESET_B(net2395),
    .D(_01514_),
    .Q_N(_13882_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[0][11] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[0][1]$_DFFE_PP_  (.CLK(clknet_leaf_271_clk),
    .RESET_B(net2396),
    .D(_01515_),
    .Q_N(_13881_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[0][1] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[0][2]$_DFFE_PP_  (.CLK(clknet_leaf_35_clk),
    .RESET_B(net2397),
    .D(_01516_),
    .Q_N(_13880_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[0][2] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[0][3]$_DFFE_PP_  (.CLK(clknet_leaf_279_clk),
    .RESET_B(net2398),
    .D(_01517_),
    .Q_N(_13879_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[0][3] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[0][4]$_DFFE_PP_  (.CLK(clknet_leaf_268_clk),
    .RESET_B(net2399),
    .D(_01518_),
    .Q_N(_13878_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[0][4] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[0][5]$_DFFE_PP_  (.CLK(clknet_leaf_269_clk),
    .RESET_B(net2400),
    .D(_01519_),
    .Q_N(_13877_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[0][5] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[0][6]$_DFFE_PP_  (.CLK(clknet_leaf_271_clk),
    .RESET_B(net2401),
    .D(_01520_),
    .Q_N(_13876_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[0][6] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[0][7]$_DFFE_PP_  (.CLK(clknet_leaf_32_clk),
    .RESET_B(net2402),
    .D(_01521_),
    .Q_N(_13875_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[0][7] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[0][8]$_DFFE_PP_  (.CLK(clknet_leaf_257_clk),
    .RESET_B(net2403),
    .D(_01522_),
    .Q_N(_13874_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[0][8] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[0][9]$_DFFE_PP_  (.CLK(clknet_leaf_249_clk),
    .RESET_B(net2404),
    .D(_01523_),
    .Q_N(_13873_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[0][9] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[10][0]$_DFFE_PP_  (.CLK(clknet_leaf_266_clk),
    .RESET_B(net2405),
    .D(_01524_),
    .Q_N(_13872_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[10][0] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[10][10]$_DFFE_PP_  (.CLK(clknet_leaf_30_clk),
    .RESET_B(net2406),
    .D(_01525_),
    .Q_N(_13871_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[10][10] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[10][11]$_DFFE_PP_  (.CLK(clknet_leaf_267_clk),
    .RESET_B(net2407),
    .D(_01526_),
    .Q_N(_13870_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[10][11] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[10][1]$_DFFE_PP_  (.CLK(clknet_leaf_266_clk),
    .RESET_B(net2408),
    .D(_01527_),
    .Q_N(_13869_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[10][1] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[10][2]$_DFFE_PP_  (.CLK(clknet_leaf_34_clk),
    .RESET_B(net2409),
    .D(_01528_),
    .Q_N(_13868_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[10][2] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[10][3]$_DFFE_PP_  (.CLK(clknet_leaf_271_clk),
    .RESET_B(net2410),
    .D(_01529_),
    .Q_N(_13867_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[10][3] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[10][4]$_DFFE_PP_  (.CLK(clknet_leaf_264_clk),
    .RESET_B(net2411),
    .D(_01530_),
    .Q_N(_13866_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[10][4] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[10][5]$_DFFE_PP_  (.CLK(clknet_leaf_266_clk),
    .RESET_B(net2412),
    .D(_01531_),
    .Q_N(_13865_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[10][5] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[10][6]$_DFFE_PP_  (.CLK(clknet_leaf_37_clk),
    .RESET_B(net2413),
    .D(_01532_),
    .Q_N(_13864_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[10][6] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[10][7]$_DFFE_PP_  (.CLK(clknet_leaf_36_clk),
    .RESET_B(net2414),
    .D(_01533_),
    .Q_N(_13863_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[10][7] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[10][8]$_DFFE_PP_  (.CLK(clknet_leaf_259_clk),
    .RESET_B(net2415),
    .D(_01534_),
    .Q_N(_13862_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[10][8] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[10][9]$_DFFE_PP_  (.CLK(clknet_leaf_257_clk),
    .RESET_B(net2416),
    .D(_01535_),
    .Q_N(_13861_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[10][9] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[11][0]$_DFFE_PP_  (.CLK(clknet_leaf_266_clk),
    .RESET_B(net2417),
    .D(_01536_),
    .Q_N(_13860_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[11][0] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[11][10]$_DFFE_PP_  (.CLK(clknet_leaf_30_clk),
    .RESET_B(net2418),
    .D(_01537_),
    .Q_N(_13859_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[11][10] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[11][11]$_DFFE_PP_  (.CLK(clknet_leaf_267_clk),
    .RESET_B(net2419),
    .D(_01538_),
    .Q_N(_13858_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[11][11] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[11][1]$_DFFE_PP_  (.CLK(clknet_leaf_266_clk),
    .RESET_B(net2420),
    .D(_01539_),
    .Q_N(_13857_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[11][1] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[11][2]$_DFFE_PP_  (.CLK(clknet_leaf_36_clk),
    .RESET_B(net2421),
    .D(_01540_),
    .Q_N(_13856_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[11][2] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[11][3]$_DFFE_PP_  (.CLK(clknet_leaf_37_clk),
    .RESET_B(net2422),
    .D(_01541_),
    .Q_N(_13855_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[11][3] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[11][4]$_DFFE_PP_  (.CLK(clknet_leaf_264_clk),
    .RESET_B(net2423),
    .D(_01542_),
    .Q_N(_13854_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[11][4] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[11][5]$_DFFE_PP_  (.CLK(clknet_leaf_265_clk),
    .RESET_B(net2424),
    .D(_01543_),
    .Q_N(_13853_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[11][5] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[11][6]$_DFFE_PP_  (.CLK(clknet_leaf_38_clk),
    .RESET_B(net2425),
    .D(_01544_),
    .Q_N(_13852_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[11][6] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[11][7]$_DFFE_PP_  (.CLK(clknet_leaf_37_clk),
    .RESET_B(net2426),
    .D(_01545_),
    .Q_N(_13851_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[11][7] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[11][8]$_DFFE_PP_  (.CLK(clknet_leaf_259_clk),
    .RESET_B(net2427),
    .D(_01546_),
    .Q_N(_13850_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[11][8] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[11][9]$_DFFE_PP_  (.CLK(clknet_leaf_258_clk),
    .RESET_B(net2428),
    .D(_01547_),
    .Q_N(_13849_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[11][9] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[12][0]$_DFFE_PP_  (.CLK(clknet_leaf_39_clk),
    .RESET_B(net2429),
    .D(_01548_),
    .Q_N(_13848_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[12][0] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[12][10]$_DFFE_PP_  (.CLK(clknet_leaf_35_clk),
    .RESET_B(net2430),
    .D(_01549_),
    .Q_N(_13847_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[12][10] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[12][11]$_DFFE_PP_  (.CLK(clknet_leaf_40_clk),
    .RESET_B(net2431),
    .D(_01550_),
    .Q_N(_13846_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[12][11] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[12][1]$_DFFE_PP_  (.CLK(clknet_leaf_38_clk),
    .RESET_B(net2432),
    .D(_01551_),
    .Q_N(_13845_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[12][1] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[12][2]$_DFFE_PP_  (.CLK(clknet_leaf_45_clk),
    .RESET_B(net2433),
    .D(_01552_),
    .Q_N(_13844_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[12][2] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[12][3]$_DFFE_PP_  (.CLK(clknet_leaf_36_clk),
    .RESET_B(net2434),
    .D(_01553_),
    .Q_N(_13843_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[12][3] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[12][4]$_DFFE_PP_  (.CLK(clknet_leaf_38_clk),
    .RESET_B(net2435),
    .D(_01554_),
    .Q_N(_13842_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[12][4] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[12][5]$_DFFE_PP_  (.CLK(clknet_leaf_45_clk),
    .RESET_B(net2436),
    .D(_01555_),
    .Q_N(_13841_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[12][5] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[12][6]$_DFFE_PP_  (.CLK(clknet_leaf_39_clk),
    .RESET_B(net2437),
    .D(_01556_),
    .Q_N(_13840_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[12][6] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[12][7]$_DFFE_PP_  (.CLK(clknet_leaf_45_clk),
    .RESET_B(net2438),
    .D(_01557_),
    .Q_N(_13839_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[12][7] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[12][8]$_DFFE_PP_  (.CLK(clknet_leaf_261_clk),
    .RESET_B(net2439),
    .D(_01558_),
    .Q_N(_13838_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[12][8] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[12][9]$_DFFE_PP_  (.CLK(clknet_leaf_258_clk),
    .RESET_B(net2440),
    .D(_01559_),
    .Q_N(_13837_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[12][9] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[13][0]$_DFFE_PP_  (.CLK(clknet_leaf_42_clk),
    .RESET_B(net2441),
    .D(_01560_),
    .Q_N(_13836_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[13][0] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[13][10]$_DFFE_PP_  (.CLK(clknet_leaf_36_clk),
    .RESET_B(net2442),
    .D(_01561_),
    .Q_N(_13835_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[13][10] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[13][11]$_DFFE_PP_  (.CLK(clknet_leaf_39_clk),
    .RESET_B(net2443),
    .D(_01562_),
    .Q_N(_13834_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[13][11] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[13][1]$_DFFE_PP_  (.CLK(clknet_leaf_38_clk),
    .RESET_B(net2444),
    .D(_01563_),
    .Q_N(_13833_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[13][1] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[13][2]$_DFFE_PP_  (.CLK(clknet_leaf_42_clk),
    .RESET_B(net2445),
    .D(_01564_),
    .Q_N(_13832_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[13][2] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[13][3]$_DFFE_PP_  (.CLK(clknet_leaf_36_clk),
    .RESET_B(net2446),
    .D(_01565_),
    .Q_N(_13831_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[13][3] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[13][4]$_DFFE_PP_  (.CLK(clknet_leaf_38_clk),
    .RESET_B(net2447),
    .D(_01566_),
    .Q_N(_13830_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[13][4] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[13][5]$_DFFE_PP_  (.CLK(clknet_leaf_35_clk),
    .RESET_B(net2448),
    .D(_01567_),
    .Q_N(_13829_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[13][5] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[13][6]$_DFFE_PP_  (.CLK(clknet_leaf_42_clk),
    .RESET_B(net2449),
    .D(_01568_),
    .Q_N(_13828_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[13][6] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[13][7]$_DFFE_PP_  (.CLK(clknet_leaf_45_clk),
    .RESET_B(net2450),
    .D(_01569_),
    .Q_N(_13827_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[13][7] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[13][8]$_DFFE_PP_  (.CLK(clknet_leaf_261_clk),
    .RESET_B(net2451),
    .D(_01570_),
    .Q_N(_13826_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[13][8] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[13][9]$_DFFE_PP_  (.CLK(clknet_leaf_258_clk),
    .RESET_B(net2452),
    .D(_01571_),
    .Q_N(_13825_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[13][9] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[14][0]$_DFFE_PP_  (.CLK(clknet_leaf_39_clk),
    .RESET_B(net2453),
    .D(_01572_),
    .Q_N(_13824_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[14][0] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[14][10]$_DFFE_PP_  (.CLK(clknet_leaf_35_clk),
    .RESET_B(net2454),
    .D(_01573_),
    .Q_N(_13823_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[14][10] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[14][11]$_DFFE_PP_  (.CLK(clknet_leaf_39_clk),
    .RESET_B(net2455),
    .D(_01574_),
    .Q_N(_13822_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[14][11] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[14][1]$_DFFE_PP_  (.CLK(clknet_leaf_38_clk),
    .RESET_B(net2456),
    .D(_01575_),
    .Q_N(_13821_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[14][1] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[14][2]$_DFFE_PP_  (.CLK(clknet_leaf_42_clk),
    .RESET_B(net2457),
    .D(_01576_),
    .Q_N(_13820_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[14][2] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[14][3]$_DFFE_PP_  (.CLK(clknet_leaf_37_clk),
    .RESET_B(net2458),
    .D(_01577_),
    .Q_N(_13819_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[14][3] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[14][4]$_DFFE_PP_  (.CLK(clknet_leaf_265_clk),
    .RESET_B(net2459),
    .D(_01578_),
    .Q_N(_13818_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[14][4] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[14][5]$_DFFE_PP_  (.CLK(clknet_leaf_36_clk),
    .RESET_B(net2460),
    .D(_01579_),
    .Q_N(_13817_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[14][5] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[14][6]$_DFFE_PP_  (.CLK(clknet_leaf_38_clk),
    .RESET_B(net2461),
    .D(_01580_),
    .Q_N(_13816_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[14][6] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[14][7]$_DFFE_PP_  (.CLK(clknet_leaf_35_clk),
    .RESET_B(net2462),
    .D(_01581_),
    .Q_N(_13815_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[14][7] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[14][8]$_DFFE_PP_  (.CLK(clknet_leaf_261_clk),
    .RESET_B(net2463),
    .D(_01582_),
    .Q_N(_13814_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[14][8] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[14][9]$_DFFE_PP_  (.CLK(clknet_leaf_259_clk),
    .RESET_B(net2464),
    .D(_01583_),
    .Q_N(_13813_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[14][9] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[15][0]$_DFFE_PP_  (.CLK(clknet_leaf_39_clk),
    .RESET_B(net2465),
    .D(_01584_),
    .Q_N(_13812_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[15][0] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[15][10]$_DFFE_PP_  (.CLK(clknet_leaf_36_clk),
    .RESET_B(net2466),
    .D(_01585_),
    .Q_N(_13811_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[15][10] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[15][11]$_DFFE_PP_  (.CLK(clknet_leaf_39_clk),
    .RESET_B(net2467),
    .D(_01586_),
    .Q_N(_13810_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[15][11] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[15][1]$_DFFE_PP_  (.CLK(clknet_leaf_38_clk),
    .RESET_B(net2468),
    .D(_01587_),
    .Q_N(_13809_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[15][1] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[15][2]$_DFFE_PP_  (.CLK(clknet_leaf_42_clk),
    .RESET_B(net2469),
    .D(_01588_),
    .Q_N(_13808_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[15][2] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[15][3]$_DFFE_PP_  (.CLK(clknet_leaf_37_clk),
    .RESET_B(net2470),
    .D(_01589_),
    .Q_N(_13807_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[15][3] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[15][4]$_DFFE_PP_  (.CLK(clknet_leaf_265_clk),
    .RESET_B(net2471),
    .D(_01590_),
    .Q_N(_13806_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[15][4] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[15][5]$_DFFE_PP_  (.CLK(clknet_leaf_35_clk),
    .RESET_B(net2472),
    .D(_01591_),
    .Q_N(_13805_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[15][5] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[15][6]$_DFFE_PP_  (.CLK(clknet_leaf_39_clk),
    .RESET_B(net2473),
    .D(_01592_),
    .Q_N(_13804_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[15][6] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[15][7]$_DFFE_PP_  (.CLK(clknet_leaf_35_clk),
    .RESET_B(net2474),
    .D(_01593_),
    .Q_N(_13803_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[15][7] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[15][8]$_DFFE_PP_  (.CLK(clknet_leaf_262_clk),
    .RESET_B(net2475),
    .D(_01594_),
    .Q_N(_13802_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[15][8] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[15][9]$_DFFE_PP_  (.CLK(clknet_leaf_258_clk),
    .RESET_B(net2476),
    .D(_01595_),
    .Q_N(_13801_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[15][9] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[16][0]$_DFFE_PP_  (.CLK(clknet_leaf_285_clk),
    .RESET_B(net2477),
    .D(_01596_),
    .Q_N(_13800_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[16][0] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[16][10]$_DFFE_PP_  (.CLK(clknet_leaf_292_clk),
    .RESET_B(net2478),
    .D(_01597_),
    .Q_N(_13799_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[16][10] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[16][11]$_DFFE_PP_  (.CLK(clknet_leaf_286_clk),
    .RESET_B(net2479),
    .D(_01598_),
    .Q_N(_13798_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[16][11] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[16][1]$_DFFE_PP_  (.CLK(clknet_leaf_291_clk),
    .RESET_B(net2480),
    .D(_01599_),
    .Q_N(_13797_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[16][1] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[16][2]$_DFFE_PP_  (.CLK(clknet_leaf_297_clk),
    .RESET_B(net2481),
    .D(_01600_),
    .Q_N(_13796_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[16][2] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[16][3]$_DFFE_PP_  (.CLK(clknet_leaf_291_clk),
    .RESET_B(net2482),
    .D(_01601_),
    .Q_N(_13795_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[16][3] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[16][4]$_DFFE_PP_  (.CLK(clknet_leaf_286_clk),
    .RESET_B(net2483),
    .D(_01602_),
    .Q_N(_13794_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[16][4] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[16][5]$_DFFE_PP_  (.CLK(clknet_leaf_285_clk),
    .RESET_B(net2484),
    .D(_01603_),
    .Q_N(_13793_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[16][5] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[16][6]$_DFFE_PP_  (.CLK(clknet_leaf_291_clk),
    .RESET_B(net2485),
    .D(_01604_),
    .Q_N(_13792_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[16][6] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[16][7]$_DFFE_PP_  (.CLK(clknet_leaf_292_clk),
    .RESET_B(net2486),
    .D(_01605_),
    .Q_N(_13791_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[16][7] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[16][8]$_DFFE_PP_  (.CLK(clknet_leaf_245_clk),
    .RESET_B(net2487),
    .D(_01606_),
    .Q_N(_13790_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[16][8] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[16][9]$_DFFE_PP_  (.CLK(clknet_leaf_244_clk),
    .RESET_B(net2488),
    .D(_01607_),
    .Q_N(_13789_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[16][9] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[17][0]$_DFFE_PP_  (.CLK(clknet_leaf_290_clk),
    .RESET_B(net2489),
    .D(_01608_),
    .Q_N(_13788_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[17][0] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[17][10]$_DFFE_PP_  (.CLK(clknet_leaf_292_clk),
    .RESET_B(net2490),
    .D(_01609_),
    .Q_N(_13787_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[17][10] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[17][11]$_DFFE_PP_  (.CLK(clknet_leaf_286_clk),
    .RESET_B(net2491),
    .D(_01610_),
    .Q_N(_13786_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[17][11] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[17][1]$_DFFE_PP_  (.CLK(clknet_leaf_290_clk),
    .RESET_B(net2492),
    .D(_01611_),
    .Q_N(_13785_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[17][1] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[17][2]$_DFFE_PP_  (.CLK(clknet_leaf_297_clk),
    .RESET_B(net2493),
    .D(_01612_),
    .Q_N(_13784_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[17][2] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[17][3]$_DFFE_PP_  (.CLK(clknet_leaf_291_clk),
    .RESET_B(net2494),
    .D(_01613_),
    .Q_N(_13783_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[17][3] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[17][4]$_DFFE_PP_  (.CLK(clknet_leaf_286_clk),
    .RESET_B(net2495),
    .D(_01614_),
    .Q_N(_13782_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[17][4] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[17][5]$_DFFE_PP_  (.CLK(clknet_leaf_287_clk),
    .RESET_B(net2496),
    .D(_01615_),
    .Q_N(_13781_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[17][5] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[17][6]$_DFFE_PP_  (.CLK(clknet_leaf_291_clk),
    .RESET_B(net2497),
    .D(_01616_),
    .Q_N(_13780_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[17][6] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[17][7]$_DFFE_PP_  (.CLK(clknet_leaf_292_clk),
    .RESET_B(net2498),
    .D(_01617_),
    .Q_N(_13779_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[17][7] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[17][8]$_DFFE_PP_  (.CLK(clknet_leaf_244_clk),
    .RESET_B(net2499),
    .D(_01618_),
    .Q_N(_13778_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[17][8] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[17][9]$_DFFE_PP_  (.CLK(clknet_leaf_244_clk),
    .RESET_B(net2500),
    .D(_01619_),
    .Q_N(_13777_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[17][9] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[18][0]$_DFFE_PP_  (.CLK(clknet_leaf_285_clk),
    .RESET_B(net2501),
    .D(_01620_),
    .Q_N(_13776_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[18][0] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[18][10]$_DFFE_PP_  (.CLK(clknet_leaf_292_clk),
    .RESET_B(net2502),
    .D(_01621_),
    .Q_N(_13775_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[18][10] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[18][11]$_DFFE_PP_  (.CLK(clknet_leaf_286_clk),
    .RESET_B(net2503),
    .D(_01622_),
    .Q_N(_13774_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[18][11] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[18][1]$_DFFE_PP_  (.CLK(clknet_leaf_290_clk),
    .RESET_B(net2504),
    .D(_01623_),
    .Q_N(_13773_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[18][1] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[18][2]$_DFFE_PP_  (.CLK(clknet_leaf_297_clk),
    .RESET_B(net2505),
    .D(_01624_),
    .Q_N(_13772_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[18][2] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[18][3]$_DFFE_PP_  (.CLK(clknet_leaf_291_clk),
    .RESET_B(net2506),
    .D(_01625_),
    .Q_N(_13771_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[18][3] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[18][4]$_DFFE_PP_  (.CLK(clknet_leaf_286_clk),
    .RESET_B(net2507),
    .D(_01626_),
    .Q_N(_13770_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[18][4] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[18][5]$_DFFE_PP_  (.CLK(clknet_leaf_286_clk),
    .RESET_B(net2508),
    .D(_01627_),
    .Q_N(_13769_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[18][5] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[18][6]$_DFFE_PP_  (.CLK(clknet_leaf_291_clk),
    .RESET_B(net2509),
    .D(_01628_),
    .Q_N(_13768_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[18][6] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[18][7]$_DFFE_PP_  (.CLK(clknet_leaf_292_clk),
    .RESET_B(net2510),
    .D(_01629_),
    .Q_N(_13767_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[18][7] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[18][8]$_DFFE_PP_  (.CLK(clknet_leaf_243_clk),
    .RESET_B(net2511),
    .D(_01630_),
    .Q_N(_13766_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[18][8] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[18][9]$_DFFE_PP_  (.CLK(clknet_leaf_245_clk),
    .RESET_B(net2512),
    .D(_01631_),
    .Q_N(_13765_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[18][9] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[19][0]$_DFFE_PP_  (.CLK(clknet_leaf_285_clk),
    .RESET_B(net2513),
    .D(_01632_),
    .Q_N(_13764_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[19][0] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[19][10]$_DFFE_PP_  (.CLK(clknet_leaf_292_clk),
    .RESET_B(net2514),
    .D(_01633_),
    .Q_N(_13763_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[19][10] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[19][11]$_DFFE_PP_  (.CLK(clknet_leaf_286_clk),
    .RESET_B(net2515),
    .D(_01634_),
    .Q_N(_13762_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[19][11] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[19][1]$_DFFE_PP_  (.CLK(clknet_leaf_290_clk),
    .RESET_B(net2516),
    .D(_01635_),
    .Q_N(_13761_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[19][1] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[19][2]$_DFFE_PP_  (.CLK(clknet_leaf_297_clk),
    .RESET_B(net2517),
    .D(_01636_),
    .Q_N(_13760_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[19][2] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[19][3]$_DFFE_PP_  (.CLK(clknet_leaf_291_clk),
    .RESET_B(net2518),
    .D(_01637_),
    .Q_N(_13759_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[19][3] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[19][4]$_DFFE_PP_  (.CLK(clknet_leaf_287_clk),
    .RESET_B(net2519),
    .D(_01638_),
    .Q_N(_13758_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[19][4] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[19][5]$_DFFE_PP_  (.CLK(clknet_leaf_287_clk),
    .RESET_B(net2520),
    .D(_01639_),
    .Q_N(_13757_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[19][5] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[19][6]$_DFFE_PP_  (.CLK(clknet_leaf_292_clk),
    .RESET_B(net2521),
    .D(_01640_),
    .Q_N(_13756_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[19][6] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[19][7]$_DFFE_PP_  (.CLK(clknet_leaf_294_clk),
    .RESET_B(net2522),
    .D(_01641_),
    .Q_N(_13755_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[19][7] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[19][8]$_DFFE_PP_  (.CLK(clknet_leaf_243_clk),
    .RESET_B(net2523),
    .D(_01642_),
    .Q_N(_13754_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[19][8] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[19][9]$_DFFE_PP_  (.CLK(clknet_leaf_245_clk),
    .RESET_B(net2524),
    .D(_01643_),
    .Q_N(_13753_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[19][9] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[1][0]$_DFFE_PP_  (.CLK(clknet_leaf_280_clk),
    .RESET_B(net2525),
    .D(_01644_),
    .Q_N(_13752_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[1][0] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[1][10]$_DFFE_PP_  (.CLK(clknet_leaf_275_clk),
    .RESET_B(net2526),
    .D(_01645_),
    .Q_N(_13751_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[1][10] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[1][11]$_DFFE_PP_  (.CLK(clknet_leaf_281_clk),
    .RESET_B(net2527),
    .D(_01646_),
    .Q_N(_13750_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[1][11] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[1][1]$_DFFE_PP_  (.CLK(clknet_leaf_279_clk),
    .RESET_B(net2528),
    .D(_01647_),
    .Q_N(_13749_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[1][1] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[1][2]$_DFFE_PP_  (.CLK(clknet_leaf_273_clk),
    .RESET_B(net2529),
    .D(_01648_),
    .Q_N(_13748_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[1][2] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[1][3]$_DFFE_PP_  (.CLK(clknet_leaf_279_clk),
    .RESET_B(net2530),
    .D(_01649_),
    .Q_N(_13747_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[1][3] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[1][4]$_DFFE_PP_  (.CLK(clknet_leaf_268_clk),
    .RESET_B(net2531),
    .D(_01650_),
    .Q_N(_13746_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[1][4] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[1][5]$_DFFE_PP_  (.CLK(clknet_leaf_269_clk),
    .RESET_B(net2532),
    .D(_01651_),
    .Q_N(_13745_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[1][5] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[1][6]$_DFFE_PP_  (.CLK(clknet_leaf_270_clk),
    .RESET_B(net2533),
    .D(_01652_),
    .Q_N(_13744_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[1][6] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[1][7]$_DFFE_PP_  (.CLK(clknet_leaf_275_clk),
    .RESET_B(net2534),
    .D(_01653_),
    .Q_N(_13743_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[1][7] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[1][8]$_DFFE_PP_  (.CLK(clknet_leaf_249_clk),
    .RESET_B(net2535),
    .D(_01654_),
    .Q_N(_13742_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[1][8] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[1][9]$_DFFE_PP_  (.CLK(clknet_leaf_249_clk),
    .RESET_B(net2536),
    .D(_01655_),
    .Q_N(_13741_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[1][9] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[20][0]$_DFFE_PP_  (.CLK(clknet_leaf_289_clk),
    .RESET_B(net2537),
    .D(_01656_),
    .Q_N(_13740_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[20][0] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[20][10]$_DFFE_PP_  (.CLK(clknet_leaf_293_clk),
    .RESET_B(net2538),
    .D(_01657_),
    .Q_N(_13739_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[20][10] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[20][11]$_DFFE_PP_  (.CLK(clknet_leaf_287_clk),
    .RESET_B(net2539),
    .D(_01658_),
    .Q_N(_13738_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[20][11] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[20][1]$_DFFE_PP_  (.CLK(clknet_leaf_289_clk),
    .RESET_B(net2540),
    .D(_01659_),
    .Q_N(_13737_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[20][1] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[20][2]$_DFFE_PP_  (.CLK(clknet_leaf_294_clk),
    .RESET_B(net2541),
    .D(_01660_),
    .Q_N(_13736_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[20][2] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[20][3]$_DFFE_PP_  (.CLK(clknet_leaf_290_clk),
    .RESET_B(net2542),
    .D(_01661_),
    .Q_N(_13735_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[20][3] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[20][4]$_DFFE_PP_  (.CLK(clknet_leaf_287_clk),
    .RESET_B(net2543),
    .D(_01662_),
    .Q_N(_13734_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[20][4] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[20][5]$_DFFE_PP_  (.CLK(clknet_leaf_288_clk),
    .RESET_B(net2544),
    .D(_01663_),
    .Q_N(_13733_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[20][5] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[20][6]$_DFFE_PP_  (.CLK(clknet_leaf_293_clk),
    .RESET_B(net2545),
    .D(_01664_),
    .Q_N(_13732_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[20][6] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[20][7]$_DFFE_PP_  (.CLK(clknet_leaf_293_clk),
    .RESET_B(net2546),
    .D(_01665_),
    .Q_N(_13731_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[20][7] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[20][8]$_DFFE_PP_  (.CLK(clknet_leaf_243_clk),
    .RESET_B(net2547),
    .D(_01666_),
    .Q_N(_13730_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[20][8] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[20][9]$_DFFE_PP_  (.CLK(clknet_leaf_244_clk),
    .RESET_B(net2548),
    .D(_01667_),
    .Q_N(_13729_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[20][9] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[21][0]$_DFFE_PP_  (.CLK(clknet_leaf_288_clk),
    .RESET_B(net2549),
    .D(_01668_),
    .Q_N(_13728_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[21][0] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[21][10]$_DFFE_PP_  (.CLK(clknet_leaf_293_clk),
    .RESET_B(net2550),
    .D(_01669_),
    .Q_N(_13727_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[21][10] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[21][11]$_DFFE_PP_  (.CLK(clknet_leaf_287_clk),
    .RESET_B(net2551),
    .D(_01670_),
    .Q_N(_13726_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[21][11] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[21][1]$_DFFE_PP_  (.CLK(clknet_leaf_289_clk),
    .RESET_B(net2552),
    .D(_01671_),
    .Q_N(_13725_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[21][1] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[21][2]$_DFFE_PP_  (.CLK(clknet_leaf_294_clk),
    .RESET_B(net2553),
    .D(_01672_),
    .Q_N(_13724_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[21][2] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[21][3]$_DFFE_PP_  (.CLK(clknet_leaf_290_clk),
    .RESET_B(net2554),
    .D(_01673_),
    .Q_N(_13723_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[21][3] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[21][4]$_DFFE_PP_  (.CLK(clknet_leaf_287_clk),
    .RESET_B(net2555),
    .D(_01674_),
    .Q_N(_13722_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[21][4] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[21][5]$_DFFE_PP_  (.CLK(clknet_leaf_288_clk),
    .RESET_B(net2556),
    .D(_01675_),
    .Q_N(_13721_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[21][5] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[21][6]$_DFFE_PP_  (.CLK(clknet_leaf_290_clk),
    .RESET_B(net2557),
    .D(_01676_),
    .Q_N(_13720_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[21][6] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[21][7]$_DFFE_PP_  (.CLK(clknet_leaf_294_clk),
    .RESET_B(net2558),
    .D(_01677_),
    .Q_N(_13719_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[21][7] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[21][8]$_DFFE_PP_  (.CLK(clknet_leaf_243_clk),
    .RESET_B(net2559),
    .D(_01678_),
    .Q_N(_13718_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[21][8] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[21][9]$_DFFE_PP_  (.CLK(clknet_leaf_244_clk),
    .RESET_B(net2560),
    .D(_01679_),
    .Q_N(_13717_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[21][9] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[22][0]$_DFFE_PP_  (.CLK(clknet_leaf_288_clk),
    .RESET_B(net2561),
    .D(_01680_),
    .Q_N(_13716_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[22][0] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[22][10]$_DFFE_PP_  (.CLK(clknet_leaf_293_clk),
    .RESET_B(net2562),
    .D(_01681_),
    .Q_N(_13715_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[22][10] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[22][11]$_DFFE_PP_  (.CLK(clknet_leaf_244_clk),
    .RESET_B(net2563),
    .D(_01682_),
    .Q_N(_13714_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[22][11] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[22][1]$_DFFE_PP_  (.CLK(clknet_leaf_289_clk),
    .RESET_B(net2564),
    .D(_01683_),
    .Q_N(_13713_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[22][1] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[22][2]$_DFFE_PP_  (.CLK(clknet_leaf_294_clk),
    .RESET_B(net2565),
    .D(_01684_),
    .Q_N(_13712_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[22][2] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[22][3]$_DFFE_PP_  (.CLK(clknet_leaf_289_clk),
    .RESET_B(net2566),
    .D(_01685_),
    .Q_N(_13711_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[22][3] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[22][4]$_DFFE_PP_  (.CLK(clknet_leaf_288_clk),
    .RESET_B(net2567),
    .D(_01686_),
    .Q_N(_13710_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[22][4] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[22][5]$_DFFE_PP_  (.CLK(clknet_leaf_288_clk),
    .RESET_B(net2568),
    .D(_01687_),
    .Q_N(_13709_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[22][5] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[22][6]$_DFFE_PP_  (.CLK(clknet_leaf_289_clk),
    .RESET_B(net2569),
    .D(_01688_),
    .Q_N(_13708_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[22][6] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[22][7]$_DFFE_PP_  (.CLK(clknet_leaf_293_clk),
    .RESET_B(net2570),
    .D(_01689_),
    .Q_N(_13707_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[22][7] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[22][8]$_DFFE_PP_  (.CLK(clknet_leaf_243_clk),
    .RESET_B(net2571),
    .D(_01690_),
    .Q_N(_13706_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[22][8] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[22][9]$_DFFE_PP_  (.CLK(clknet_leaf_244_clk),
    .RESET_B(net2572),
    .D(_01691_),
    .Q_N(_13705_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[22][9] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[23][0]$_DFFE_PP_  (.CLK(clknet_leaf_288_clk),
    .RESET_B(net2573),
    .D(_01692_),
    .Q_N(_13704_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[23][0] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[23][10]$_DFFE_PP_  (.CLK(clknet_leaf_293_clk),
    .RESET_B(net2574),
    .D(_01693_),
    .Q_N(_13703_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[23][10] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[23][11]$_DFFE_PP_  (.CLK(clknet_leaf_244_clk),
    .RESET_B(net2575),
    .D(_01694_),
    .Q_N(_13702_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[23][11] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[23][1]$_DFFE_PP_  (.CLK(clknet_leaf_289_clk),
    .RESET_B(net2576),
    .D(_01695_),
    .Q_N(_13701_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[23][1] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[23][2]$_DFFE_PP_  (.CLK(clknet_leaf_294_clk),
    .RESET_B(net2577),
    .D(_01696_),
    .Q_N(_13700_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[23][2] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[23][3]$_DFFE_PP_  (.CLK(clknet_leaf_290_clk),
    .RESET_B(net2578),
    .D(_01697_),
    .Q_N(_13699_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[23][3] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[23][4]$_DFFE_PP_  (.CLK(clknet_leaf_287_clk),
    .RESET_B(net2579),
    .D(_01698_),
    .Q_N(_13698_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[23][4] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[23][5]$_DFFE_PP_  (.CLK(clknet_leaf_288_clk),
    .RESET_B(net2580),
    .D(_01699_),
    .Q_N(_13697_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[23][5] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[23][6]$_DFFE_PP_  (.CLK(clknet_leaf_289_clk),
    .RESET_B(net2581),
    .D(_01700_),
    .Q_N(_13696_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[23][6] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[23][7]$_DFFE_PP_  (.CLK(clknet_leaf_293_clk),
    .RESET_B(net2582),
    .D(_01701_),
    .Q_N(_13695_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[23][7] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[23][8]$_DFFE_PP_  (.CLK(clknet_leaf_243_clk),
    .RESET_B(net2583),
    .D(_01702_),
    .Q_N(_13694_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[23][8] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[23][9]$_DFFE_PP_  (.CLK(clknet_leaf_243_clk),
    .RESET_B(net2584),
    .D(_01703_),
    .Q_N(_13693_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[23][9] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[24][0]$_DFFE_PP_  (.CLK(clknet_leaf_283_clk),
    .RESET_B(net2585),
    .D(_01704_),
    .Q_N(_13692_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[24][0] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[24][10]$_DFFE_PP_  (.CLK(clknet_leaf_297_clk),
    .RESET_B(net2586),
    .D(_01705_),
    .Q_N(_13691_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[24][10] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[24][11]$_DFFE_PP_  (.CLK(clknet_leaf_282_clk),
    .RESET_B(net2587),
    .D(_01706_),
    .Q_N(_13690_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[24][11] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[24][1]$_DFFE_PP_  (.CLK(clknet_leaf_284_clk),
    .RESET_B(net2588),
    .D(_01707_),
    .Q_N(_13689_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[24][1] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[24][2]$_DFFE_PP_  (.CLK(clknet_leaf_299_clk),
    .RESET_B(net2589),
    .D(_01708_),
    .Q_N(_13688_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[24][2] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[24][3]$_DFFE_PP_  (.CLK(clknet_leaf_278_clk),
    .RESET_B(net2590),
    .D(_01709_),
    .Q_N(_13687_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[24][3] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[24][4]$_DFFE_PP_  (.CLK(clknet_leaf_285_clk),
    .RESET_B(net2591),
    .D(_01710_),
    .Q_N(_13686_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[24][4] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[24][5]$_DFFE_PP_  (.CLK(clknet_leaf_285_clk),
    .RESET_B(net2592),
    .D(_01711_),
    .Q_N(_13685_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[24][5] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[24][6]$_DFFE_PP_  (.CLK(clknet_leaf_298_clk),
    .RESET_B(net2593),
    .D(_01712_),
    .Q_N(_13684_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[24][6] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[24][7]$_DFFE_PP_  (.CLK(clknet_leaf_299_clk),
    .RESET_B(net2594),
    .D(_01713_),
    .Q_N(_13683_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[24][7] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[24][8]$_DFFE_PP_  (.CLK(clknet_leaf_246_clk),
    .RESET_B(net2595),
    .D(_01714_),
    .Q_N(_13682_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[24][8] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[24][9]$_DFFE_PP_  (.CLK(clknet_leaf_245_clk),
    .RESET_B(net2596),
    .D(_01715_),
    .Q_N(_13681_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[24][9] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[25][0]$_DFFE_PP_  (.CLK(clknet_leaf_284_clk),
    .RESET_B(net2597),
    .D(_01716_),
    .Q_N(_13680_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[25][0] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[25][10]$_DFFE_PP_  (.CLK(clknet_leaf_297_clk),
    .RESET_B(net2598),
    .D(_01717_),
    .Q_N(_13679_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[25][10] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[25][11]$_DFFE_PP_  (.CLK(clknet_leaf_248_clk),
    .RESET_B(net2599),
    .D(_01718_),
    .Q_N(_13678_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[25][11] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[25][1]$_DFFE_PP_  (.CLK(clknet_leaf_284_clk),
    .RESET_B(net2600),
    .D(_01719_),
    .Q_N(_13677_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[25][1] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[25][2]$_DFFE_PP_  (.CLK(clknet_leaf_299_clk),
    .RESET_B(net2601),
    .D(_01720_),
    .Q_N(_13676_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[25][2] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[25][3]$_DFFE_PP_  (.CLK(clknet_leaf_276_clk),
    .RESET_B(net2602),
    .D(_01721_),
    .Q_N(_13675_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[25][3] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[25][4]$_DFFE_PP_  (.CLK(clknet_leaf_245_clk),
    .RESET_B(net2603),
    .D(_01722_),
    .Q_N(_13674_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[25][4] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[25][5]$_DFFE_PP_  (.CLK(clknet_leaf_283_clk),
    .RESET_B(net2604),
    .D(_01723_),
    .Q_N(_13673_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[25][5] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[25][6]$_DFFE_PP_  (.CLK(clknet_leaf_277_clk),
    .RESET_B(net2605),
    .D(_01724_),
    .Q_N(_13672_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[25][6] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[25][7]$_DFFE_PP_  (.CLK(clknet_leaf_275_clk),
    .RESET_B(net2606),
    .D(_01725_),
    .Q_N(_13671_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[25][7] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[25][8]$_DFFE_PP_  (.CLK(clknet_leaf_246_clk),
    .RESET_B(net2607),
    .D(_01726_),
    .Q_N(_13670_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[25][8] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[25][9]$_DFFE_PP_  (.CLK(clknet_leaf_245_clk),
    .RESET_B(net2608),
    .D(_01727_),
    .Q_N(_13669_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[25][9] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[26][0]$_DFFE_PP_  (.CLK(clknet_leaf_285_clk),
    .RESET_B(net2609),
    .D(_01728_),
    .Q_N(_13668_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[26][0] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[26][10]$_DFFE_PP_  (.CLK(clknet_leaf_298_clk),
    .RESET_B(net2610),
    .D(_01729_),
    .Q_N(_13667_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[26][10] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[26][11]$_DFFE_PP_  (.CLK(clknet_leaf_248_clk),
    .RESET_B(net2611),
    .D(_01730_),
    .Q_N(_13666_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[26][11] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[26][1]$_DFFE_PP_  (.CLK(clknet_leaf_284_clk),
    .RESET_B(net2612),
    .D(_01731_),
    .Q_N(_13665_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[26][1] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[26][2]$_DFFE_PP_  (.CLK(clknet_leaf_299_clk),
    .RESET_B(net2613),
    .D(_01732_),
    .Q_N(_13664_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[26][2] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[26][3]$_DFFE_PP_  (.CLK(clknet_leaf_277_clk),
    .RESET_B(net2614),
    .D(_01733_),
    .Q_N(_13663_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[26][3] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[26][4]$_DFFE_PP_  (.CLK(clknet_leaf_245_clk),
    .RESET_B(net2615),
    .D(_01734_),
    .Q_N(_13662_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[26][4] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[26][5]$_DFFE_PP_  (.CLK(clknet_leaf_283_clk),
    .RESET_B(net2616),
    .D(_01735_),
    .Q_N(_13661_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[26][5] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[26][6]$_DFFE_PP_  (.CLK(clknet_leaf_298_clk),
    .RESET_B(net2617),
    .D(_01736_),
    .Q_N(_13660_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[26][6] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[26][7]$_DFFE_PP_  (.CLK(clknet_leaf_277_clk),
    .RESET_B(net2618),
    .D(_01737_),
    .Q_N(_13659_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[26][7] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[26][8]$_DFFE_PP_  (.CLK(clknet_leaf_246_clk),
    .RESET_B(net2619),
    .D(_01738_),
    .Q_N(_13658_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[26][8] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[26][9]$_DFFE_PP_  (.CLK(clknet_leaf_246_clk),
    .RESET_B(net2620),
    .D(_01739_),
    .Q_N(_13657_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[26][9] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[27][0]$_DFFE_PP_  (.CLK(clknet_leaf_283_clk),
    .RESET_B(net2621),
    .D(_01740_),
    .Q_N(_13656_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[27][0] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[27][10]$_DFFE_PP_  (.CLK(clknet_leaf_298_clk),
    .RESET_B(net2622),
    .D(_01741_),
    .Q_N(_13655_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[27][10] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[27][11]$_DFFE_PP_  (.CLK(clknet_leaf_282_clk),
    .RESET_B(net2623),
    .D(_01742_),
    .Q_N(_13654_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[27][11] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[27][1]$_DFFE_PP_  (.CLK(clknet_leaf_284_clk),
    .RESET_B(net2624),
    .D(_01743_),
    .Q_N(_13653_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[27][1] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[27][2]$_DFFE_PP_  (.CLK(clknet_leaf_299_clk),
    .RESET_B(net2625),
    .D(_01744_),
    .Q_N(_13652_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[27][2] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[27][3]$_DFFE_PP_  (.CLK(clknet_leaf_276_clk),
    .RESET_B(net2626),
    .D(_01745_),
    .Q_N(_13651_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[27][3] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[27][4]$_DFFE_PP_  (.CLK(clknet_leaf_248_clk),
    .RESET_B(net2627),
    .D(_01746_),
    .Q_N(_13650_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[27][4] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[27][5]$_DFFE_PP_  (.CLK(clknet_leaf_283_clk),
    .RESET_B(net2628),
    .D(_01747_),
    .Q_N(_13649_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[27][5] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[27][6]$_DFFE_PP_  (.CLK(clknet_leaf_277_clk),
    .RESET_B(net2629),
    .D(_01748_),
    .Q_N(_13648_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[27][6] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[27][7]$_DFFE_PP_  (.CLK(clknet_leaf_275_clk),
    .RESET_B(net2630),
    .D(_01749_),
    .Q_N(_13647_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[27][7] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[27][8]$_DFFE_PP_  (.CLK(clknet_leaf_246_clk),
    .RESET_B(net2631),
    .D(_01750_),
    .Q_N(_13646_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[27][8] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[27][9]$_DFFE_PP_  (.CLK(clknet_leaf_245_clk),
    .RESET_B(net2632),
    .D(_01751_),
    .Q_N(_13645_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[27][9] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[28][0]$_DFFE_PP_  (.CLK(clknet_leaf_283_clk),
    .RESET_B(net2633),
    .D(_01752_),
    .Q_N(_13644_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[28][0] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[28][10]$_DFFE_PP_  (.CLK(clknet_leaf_298_clk),
    .RESET_B(net2634),
    .D(_01753_),
    .Q_N(_13643_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[28][10] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[28][11]$_DFFE_PP_  (.CLK(clknet_leaf_281_clk),
    .RESET_B(net2635),
    .D(_01754_),
    .Q_N(_13642_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[28][11] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[28][1]$_DFFE_PP_  (.CLK(clknet_leaf_278_clk),
    .RESET_B(net2636),
    .D(_01755_),
    .Q_N(_13641_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[28][1] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[28][2]$_DFFE_PP_  (.CLK(clknet_leaf_275_clk),
    .RESET_B(net2637),
    .D(_01756_),
    .Q_N(_13640_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[28][2] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[28][3]$_DFFE_PP_  (.CLK(clknet_leaf_278_clk),
    .RESET_B(net2638),
    .D(_01757_),
    .Q_N(_13639_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[28][3] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[28][4]$_DFFE_PP_  (.CLK(clknet_leaf_283_clk),
    .RESET_B(net2639),
    .D(_01758_),
    .Q_N(_13638_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[28][4] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[28][5]$_DFFE_PP_  (.CLK(clknet_leaf_282_clk),
    .RESET_B(net2640),
    .D(_01759_),
    .Q_N(_13637_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[28][5] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[28][6]$_DFFE_PP_  (.CLK(clknet_leaf_277_clk),
    .RESET_B(net2641),
    .D(_01760_),
    .Q_N(_13636_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[28][6] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[28][7]$_DFFE_PP_  (.CLK(clknet_leaf_277_clk),
    .RESET_B(net2642),
    .D(_01761_),
    .Q_N(_13635_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[28][7] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[28][8]$_DFFE_PP_  (.CLK(clknet_leaf_246_clk),
    .RESET_B(net2643),
    .D(_01762_),
    .Q_N(_13634_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[28][8] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[28][9]$_DFFE_PP_  (.CLK(clknet_leaf_248_clk),
    .RESET_B(net2644),
    .D(_01763_),
    .Q_N(_13633_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[28][9] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[29][0]$_DFFE_PP_  (.CLK(clknet_leaf_278_clk),
    .RESET_B(net2645),
    .D(_01764_),
    .Q_N(_13632_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[29][0] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[29][10]$_DFFE_PP_  (.CLK(clknet_leaf_298_clk),
    .RESET_B(net2646),
    .D(_01765_),
    .Q_N(_13631_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[29][10] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[29][11]$_DFFE_PP_  (.CLK(clknet_leaf_281_clk),
    .RESET_B(net2647),
    .D(_01766_),
    .Q_N(_13630_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[29][11] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[29][1]$_DFFE_PP_  (.CLK(clknet_leaf_280_clk),
    .RESET_B(net2648),
    .D(_01767_),
    .Q_N(_13629_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[29][1] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[29][2]$_DFFE_PP_  (.CLK(clknet_leaf_276_clk),
    .RESET_B(net2649),
    .D(_01768_),
    .Q_N(_13628_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[29][2] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[29][3]$_DFFE_PP_  (.CLK(clknet_leaf_279_clk),
    .RESET_B(net2650),
    .D(_01769_),
    .Q_N(_13627_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[29][3] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[29][4]$_DFFE_PP_  (.CLK(clknet_leaf_283_clk),
    .RESET_B(net2651),
    .D(_01770_),
    .Q_N(_13626_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[29][4] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[29][5]$_DFFE_PP_  (.CLK(clknet_leaf_280_clk),
    .RESET_B(net2652),
    .D(_01771_),
    .Q_N(_13625_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[29][5] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[29][6]$_DFFE_PP_  (.CLK(clknet_leaf_284_clk),
    .RESET_B(net2653),
    .D(_01772_),
    .Q_N(_13624_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[29][6] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[29][7]$_DFFE_PP_  (.CLK(clknet_leaf_277_clk),
    .RESET_B(net2654),
    .D(_01773_),
    .Q_N(_13623_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[29][7] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[29][8]$_DFFE_PP_  (.CLK(clknet_leaf_248_clk),
    .RESET_B(net2655),
    .D(_01774_),
    .Q_N(_13622_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[29][8] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[29][9]$_DFFE_PP_  (.CLK(clknet_leaf_248_clk),
    .RESET_B(net2656),
    .D(_01775_),
    .Q_N(_13621_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[29][9] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[2][0]$_DFFE_PP_  (.CLK(clknet_leaf_279_clk),
    .RESET_B(net2657),
    .D(_01776_),
    .Q_N(_13620_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[2][0] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[2][10]$_DFFE_PP_  (.CLK(clknet_leaf_273_clk),
    .RESET_B(net2658),
    .D(_01777_),
    .Q_N(_13619_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[2][10] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[2][11]$_DFFE_PP_  (.CLK(clknet_leaf_281_clk),
    .RESET_B(net2659),
    .D(_01778_),
    .Q_N(_13618_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[2][11] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[2][1]$_DFFE_PP_  (.CLK(clknet_leaf_270_clk),
    .RESET_B(net2660),
    .D(_01779_),
    .Q_N(_13617_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[2][1] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[2][2]$_DFFE_PP_  (.CLK(clknet_leaf_275_clk),
    .RESET_B(net2661),
    .D(_01780_),
    .Q_N(_13616_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[2][2] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[2][3]$_DFFE_PP_  (.CLK(clknet_leaf_279_clk),
    .RESET_B(net2662),
    .D(_01781_),
    .Q_N(_13615_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[2][3] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[2][4]$_DFFE_PP_  (.CLK(clknet_leaf_268_clk),
    .RESET_B(net2663),
    .D(_01782_),
    .Q_N(_13614_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[2][4] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[2][5]$_DFFE_PP_  (.CLK(clknet_leaf_280_clk),
    .RESET_B(net2664),
    .D(_01783_),
    .Q_N(_13613_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[2][5] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[2][6]$_DFFE_PP_  (.CLK(clknet_leaf_270_clk),
    .RESET_B(net2665),
    .D(_01784_),
    .Q_N(_13612_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[2][6] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[2][7]$_DFFE_PP_  (.CLK(clknet_leaf_272_clk),
    .RESET_B(net2666),
    .D(_01785_),
    .Q_N(_13611_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[2][7] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[2][8]$_DFFE_PP_  (.CLK(clknet_leaf_257_clk),
    .RESET_B(net2667),
    .D(_01786_),
    .Q_N(_13610_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[2][8] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[2][9]$_DFFE_PP_  (.CLK(clknet_leaf_249_clk),
    .RESET_B(net2668),
    .D(_01787_),
    .Q_N(_13609_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[2][9] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[30][0]$_DFFE_PP_  (.CLK(clknet_leaf_282_clk),
    .RESET_B(net2669),
    .D(_01788_),
    .Q_N(_13608_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[30][0] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[30][10]$_DFFE_PP_  (.CLK(clknet_leaf_298_clk),
    .RESET_B(net2670),
    .D(_01789_),
    .Q_N(_13607_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[30][10] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[30][11]$_DFFE_PP_  (.CLK(clknet_leaf_281_clk),
    .RESET_B(net2671),
    .D(_01790_),
    .Q_N(_13606_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[30][11] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[30][1]$_DFFE_PP_  (.CLK(clknet_leaf_278_clk),
    .RESET_B(net2672),
    .D(_01791_),
    .Q_N(_13605_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[30][1] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[30][2]$_DFFE_PP_  (.CLK(clknet_leaf_276_clk),
    .RESET_B(net2673),
    .D(_01792_),
    .Q_N(_13604_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[30][2] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[30][3]$_DFFE_PP_  (.CLK(clknet_leaf_278_clk),
    .RESET_B(net2674),
    .D(_01793_),
    .Q_N(_13603_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[30][3] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[30][4]$_DFFE_PP_  (.CLK(clknet_leaf_282_clk),
    .RESET_B(net2675),
    .D(_01794_),
    .Q_N(_13602_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[30][4] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[30][5]$_DFFE_PP_  (.CLK(clknet_leaf_282_clk),
    .RESET_B(net2676),
    .D(_01795_),
    .Q_N(_13601_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[30][5] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[30][6]$_DFFE_PP_  (.CLK(clknet_leaf_284_clk),
    .RESET_B(net2677),
    .D(_01796_),
    .Q_N(_13600_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[30][6] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[30][7]$_DFFE_PP_  (.CLK(clknet_leaf_276_clk),
    .RESET_B(net2678),
    .D(_01797_),
    .Q_N(_13599_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[30][7] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[30][8]$_DFFE_PP_  (.CLK(clknet_leaf_247_clk),
    .RESET_B(net2679),
    .D(_01798_),
    .Q_N(_13598_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[30][8] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[30][9]$_DFFE_PP_  (.CLK(clknet_leaf_249_clk),
    .RESET_B(net2680),
    .D(_01799_),
    .Q_N(_13597_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[30][9] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[31][0]$_DFFE_PP_  (.CLK(clknet_leaf_280_clk),
    .RESET_B(net2681),
    .D(_01800_),
    .Q_N(_13596_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[31][0] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[31][10]$_DFFE_PP_  (.CLK(clknet_leaf_298_clk),
    .RESET_B(net2682),
    .D(_01801_),
    .Q_N(_13595_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[31][10] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[31][11]$_DFFE_PP_  (.CLK(clknet_leaf_282_clk),
    .RESET_B(net2683),
    .D(_01802_),
    .Q_N(_13594_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[31][11] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[31][1]$_DFFE_PP_  (.CLK(clknet_leaf_278_clk),
    .RESET_B(net2684),
    .D(_01803_),
    .Q_N(_13593_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[31][1] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[31][2]$_DFFE_PP_  (.CLK(clknet_leaf_276_clk),
    .RESET_B(net2685),
    .D(_01804_),
    .Q_N(_13592_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[31][2] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[31][3]$_DFFE_PP_  (.CLK(clknet_leaf_278_clk),
    .RESET_B(net2686),
    .D(_01805_),
    .Q_N(_13591_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[31][3] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[31][4]$_DFFE_PP_  (.CLK(clknet_leaf_285_clk),
    .RESET_B(net2687),
    .D(_01806_),
    .Q_N(_13590_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[31][4] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[31][5]$_DFFE_PP_  (.CLK(clknet_leaf_282_clk),
    .RESET_B(net2688),
    .D(_01807_),
    .Q_N(_13589_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[31][5] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[31][6]$_DFFE_PP_  (.CLK(clknet_leaf_284_clk),
    .RESET_B(net2689),
    .D(_01808_),
    .Q_N(_13588_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[31][6] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[31][7]$_DFFE_PP_  (.CLK(clknet_leaf_277_clk),
    .RESET_B(net2690),
    .D(_01809_),
    .Q_N(_13587_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[31][7] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[31][8]$_DFFE_PP_  (.CLK(clknet_leaf_248_clk),
    .RESET_B(net2691),
    .D(_01810_),
    .Q_N(_13586_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[31][8] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[31][9]$_DFFE_PP_  (.CLK(clknet_leaf_248_clk),
    .RESET_B(net2692),
    .D(_01811_),
    .Q_N(_13585_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[31][9] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[3][0]$_DFFE_PP_  (.CLK(clknet_leaf_270_clk),
    .RESET_B(net2693),
    .D(_01812_),
    .Q_N(_13584_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[3][0] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[3][10]$_DFFE_PP_  (.CLK(clknet_leaf_273_clk),
    .RESET_B(net2694),
    .D(_01813_),
    .Q_N(_13583_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[3][10] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[3][11]$_DFFE_PP_  (.CLK(clknet_leaf_281_clk),
    .RESET_B(net2695),
    .D(_01814_),
    .Q_N(_13582_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[3][11] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[3][1]$_DFFE_PP_  (.CLK(clknet_leaf_269_clk),
    .RESET_B(net2696),
    .D(_01815_),
    .Q_N(_13581_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[3][1] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[3][2]$_DFFE_PP_  (.CLK(clknet_leaf_273_clk),
    .RESET_B(net2697),
    .D(_01816_),
    .Q_N(_13580_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[3][2] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[3][3]$_DFFE_PP_  (.CLK(clknet_leaf_279_clk),
    .RESET_B(net2698),
    .D(_01817_),
    .Q_N(_13579_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[3][3] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[3][4]$_DFFE_PP_  (.CLK(clknet_leaf_257_clk),
    .RESET_B(net2699),
    .D(_01818_),
    .Q_N(_13578_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[3][4] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[3][5]$_DFFE_PP_  (.CLK(clknet_leaf_280_clk),
    .RESET_B(net2700),
    .D(_01819_),
    .Q_N(_13577_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[3][5] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[3][6]$_DFFE_PP_  (.CLK(clknet_leaf_270_clk),
    .RESET_B(net2701),
    .D(_01820_),
    .Q_N(_13576_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[3][6] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[3][7]$_DFFE_PP_  (.CLK(clknet_leaf_273_clk),
    .RESET_B(net2702),
    .D(_01821_),
    .Q_N(_13575_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[3][7] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[3][8]$_DFFE_PP_  (.CLK(clknet_leaf_257_clk),
    .RESET_B(net2703),
    .D(_01822_),
    .Q_N(_13574_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[3][8] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[3][9]$_DFFE_PP_  (.CLK(clknet_leaf_249_clk),
    .RESET_B(net2704),
    .D(_01823_),
    .Q_N(_13573_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[3][9] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[4][0]$_DFFE_PP_  (.CLK(clknet_leaf_269_clk),
    .RESET_B(net2705),
    .D(_01824_),
    .Q_N(_13572_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[4][0] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[4][10]$_DFFE_PP_  (.CLK(clknet_leaf_272_clk),
    .RESET_B(net2706),
    .D(_01825_),
    .Q_N(_13571_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[4][10] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[4][11]$_DFFE_PP_  (.CLK(clknet_leaf_280_clk),
    .RESET_B(net2707),
    .D(_01826_),
    .Q_N(_13570_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[4][11] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[4][1]$_DFFE_PP_  (.CLK(clknet_leaf_270_clk),
    .RESET_B(net2708),
    .D(_01827_),
    .Q_N(_13569_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[4][1] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[4][2]$_DFFE_PP_  (.CLK(clknet_leaf_272_clk),
    .RESET_B(net2709),
    .D(_01828_),
    .Q_N(_13568_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[4][2] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[4][3]$_DFFE_PP_  (.CLK(clknet_leaf_276_clk),
    .RESET_B(net2710),
    .D(_01829_),
    .Q_N(_13567_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[4][3] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[4][4]$_DFFE_PP_  (.CLK(clknet_leaf_268_clk),
    .RESET_B(net2711),
    .D(_01830_),
    .Q_N(_13566_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[4][4] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[4][5]$_DFFE_PP_  (.CLK(clknet_leaf_280_clk),
    .RESET_B(net2712),
    .D(_01831_),
    .Q_N(_13565_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[4][5] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[4][6]$_DFFE_PP_  (.CLK(clknet_leaf_272_clk),
    .RESET_B(net2713),
    .D(_01832_),
    .Q_N(_13564_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[4][6] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[4][7]$_DFFE_PP_  (.CLK(clknet_leaf_272_clk),
    .RESET_B(net2714),
    .D(_01833_),
    .Q_N(_13563_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[4][7] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[4][8]$_DFFE_PP_  (.CLK(clknet_leaf_258_clk),
    .RESET_B(net2715),
    .D(_01834_),
    .Q_N(_13562_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[4][8] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[4][9]$_DFFE_PP_  (.CLK(clknet_leaf_249_clk),
    .RESET_B(net2716),
    .D(_01835_),
    .Q_N(_13561_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[4][9] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[5][0]$_DFFE_PP_  (.CLK(clknet_leaf_269_clk),
    .RESET_B(net2717),
    .D(_01836_),
    .Q_N(_13560_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[5][0] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[5][10]$_DFFE_PP_  (.CLK(clknet_leaf_272_clk),
    .RESET_B(net2718),
    .D(_01837_),
    .Q_N(_13559_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[5][10] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[5][11]$_DFFE_PP_  (.CLK(clknet_leaf_281_clk),
    .RESET_B(net2719),
    .D(_01838_),
    .Q_N(_13558_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[5][11] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[5][1]$_DFFE_PP_  (.CLK(clknet_leaf_269_clk),
    .RESET_B(net2720),
    .D(_01839_),
    .Q_N(_13557_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[5][1] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[5][2]$_DFFE_PP_  (.CLK(clknet_leaf_31_clk),
    .RESET_B(net2721),
    .D(_01840_),
    .Q_N(_13556_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[5][2] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[5][3]$_DFFE_PP_  (.CLK(clknet_leaf_273_clk),
    .RESET_B(net2722),
    .D(_01841_),
    .Q_N(_13555_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[5][3] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[5][4]$_DFFE_PP_  (.CLK(clknet_leaf_267_clk),
    .RESET_B(net2723),
    .D(_01842_),
    .Q_N(_13554_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[5][4] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[5][5]$_DFFE_PP_  (.CLK(clknet_leaf_268_clk),
    .RESET_B(net2724),
    .D(_01843_),
    .Q_N(_13553_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[5][5] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[5][6]$_DFFE_PP_  (.CLK(clknet_leaf_271_clk),
    .RESET_B(net2725),
    .D(_01844_),
    .Q_N(_13552_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[5][6] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[5][7]$_DFFE_PP_  (.CLK(clknet_leaf_271_clk),
    .RESET_B(net2726),
    .D(_01845_),
    .Q_N(_13551_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[5][7] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[5][8]$_DFFE_PP_  (.CLK(clknet_leaf_259_clk),
    .RESET_B(net2727),
    .D(_01846_),
    .Q_N(_13550_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[5][8] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[5][9]$_DFFE_PP_  (.CLK(clknet_leaf_257_clk),
    .RESET_B(net2728),
    .D(_01847_),
    .Q_N(_13549_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[5][9] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[6][0]$_DFFE_PP_  (.CLK(clknet_leaf_266_clk),
    .RESET_B(net2729),
    .D(_01848_),
    .Q_N(_13548_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[6][0] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[6][10]$_DFFE_PP_  (.CLK(clknet_leaf_273_clk),
    .RESET_B(net2730),
    .D(_01849_),
    .Q_N(_13547_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[6][10] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[6][11]$_DFFE_PP_  (.CLK(clknet_leaf_269_clk),
    .RESET_B(net2731),
    .D(_01850_),
    .Q_N(_13546_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[6][11] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[6][1]$_DFFE_PP_  (.CLK(clknet_leaf_270_clk),
    .RESET_B(net2732),
    .D(_01851_),
    .Q_N(_13545_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[6][1] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[6][2]$_DFFE_PP_  (.CLK(clknet_leaf_31_clk),
    .RESET_B(net2733),
    .D(_01852_),
    .Q_N(_13544_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[6][2] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[6][3]$_DFFE_PP_  (.CLK(clknet_leaf_276_clk),
    .RESET_B(net2734),
    .D(_01853_),
    .Q_N(_13543_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[6][3] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[6][4]$_DFFE_PP_  (.CLK(clknet_leaf_268_clk),
    .RESET_B(net2735),
    .D(_01854_),
    .Q_N(_13542_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[6][4] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[6][5]$_DFFE_PP_  (.CLK(clknet_leaf_268_clk),
    .RESET_B(net2736),
    .D(_01855_),
    .Q_N(_13541_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[6][5] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[6][6]$_DFFE_PP_  (.CLK(clknet_leaf_272_clk),
    .RESET_B(net2737),
    .D(_01856_),
    .Q_N(_13540_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[6][6] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[6][7]$_DFFE_PP_  (.CLK(clknet_leaf_271_clk),
    .RESET_B(net2738),
    .D(_01857_),
    .Q_N(_13539_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[6][7] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[6][8]$_DFFE_PP_  (.CLK(clknet_leaf_258_clk),
    .RESET_B(net2739),
    .D(_01858_),
    .Q_N(_13538_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[6][8] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[6][9]$_DFFE_PP_  (.CLK(clknet_leaf_249_clk),
    .RESET_B(net2740),
    .D(_01859_),
    .Q_N(_13537_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[6][9] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[7][0]$_DFFE_PP_  (.CLK(clknet_leaf_266_clk),
    .RESET_B(net2741),
    .D(_01860_),
    .Q_N(_13536_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[7][0] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[7][10]$_DFFE_PP_  (.CLK(clknet_leaf_272_clk),
    .RESET_B(net2742),
    .D(_01861_),
    .Q_N(_13535_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[7][10] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[7][11]$_DFFE_PP_  (.CLK(clknet_leaf_269_clk),
    .RESET_B(net2743),
    .D(_01862_),
    .Q_N(_13534_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[7][11] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[7][1]$_DFFE_PP_  (.CLK(clknet_leaf_271_clk),
    .RESET_B(net2744),
    .D(_01863_),
    .Q_N(_13533_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[7][1] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[7][2]$_DFFE_PP_  (.CLK(clknet_leaf_30_clk),
    .RESET_B(net2745),
    .D(_01864_),
    .Q_N(_13532_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[7][2] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[7][3]$_DFFE_PP_  (.CLK(clknet_leaf_270_clk),
    .RESET_B(net2746),
    .D(_01865_),
    .Q_N(_13531_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[7][3] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[7][4]$_DFFE_PP_  (.CLK(clknet_leaf_267_clk),
    .RESET_B(net2747),
    .D(_01866_),
    .Q_N(_13530_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[7][4] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[7][5]$_DFFE_PP_  (.CLK(clknet_leaf_268_clk),
    .RESET_B(net2748),
    .D(_01867_),
    .Q_N(_13529_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[7][5] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[7][6]$_DFFE_PP_  (.CLK(clknet_leaf_271_clk),
    .RESET_B(net2749),
    .D(_01868_),
    .Q_N(_13528_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[7][6] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[7][7]$_DFFE_PP_  (.CLK(clknet_leaf_31_clk),
    .RESET_B(net2750),
    .D(_01869_),
    .Q_N(_13527_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[7][7] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[7][8]$_DFFE_PP_  (.CLK(clknet_leaf_259_clk),
    .RESET_B(net2751),
    .D(_01870_),
    .Q_N(_13526_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[7][8] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[7][9]$_DFFE_PP_  (.CLK(clknet_leaf_258_clk),
    .RESET_B(net2752),
    .D(_01871_),
    .Q_N(_13525_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[7][9] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[8][0]$_DFFE_PP_  (.CLK(clknet_leaf_265_clk),
    .RESET_B(net2753),
    .D(_01872_),
    .Q_N(_13524_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[8][0] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[8][10]$_DFFE_PP_  (.CLK(clknet_leaf_31_clk),
    .RESET_B(net2754),
    .D(_01873_),
    .Q_N(_13523_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[8][10] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[8][11]$_DFFE_PP_  (.CLK(clknet_leaf_267_clk),
    .RESET_B(net2755),
    .D(_01874_),
    .Q_N(_13522_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[8][11] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[8][1]$_DFFE_PP_  (.CLK(clknet_leaf_265_clk),
    .RESET_B(net2756),
    .D(_01875_),
    .Q_N(_13521_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[8][1] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[8][2]$_DFFE_PP_  (.CLK(clknet_leaf_31_clk),
    .RESET_B(net2757),
    .D(_01876_),
    .Q_N(_13520_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[8][2] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[8][3]$_DFFE_PP_  (.CLK(clknet_leaf_265_clk),
    .RESET_B(net2758),
    .D(_01877_),
    .Q_N(_13519_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[8][3] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[8][4]$_DFFE_PP_  (.CLK(clknet_leaf_264_clk),
    .RESET_B(net2759),
    .D(_01878_),
    .Q_N(_13518_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[8][4] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[8][5]$_DFFE_PP_  (.CLK(clknet_leaf_266_clk),
    .RESET_B(net2760),
    .D(_01879_),
    .Q_N(_13517_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[8][5] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[8][6]$_DFFE_PP_  (.CLK(clknet_leaf_37_clk),
    .RESET_B(net2761),
    .D(_01880_),
    .Q_N(_13516_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[8][6] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[8][7]$_DFFE_PP_  (.CLK(clknet_leaf_36_clk),
    .RESET_B(net2762),
    .D(_01881_),
    .Q_N(_13515_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[8][7] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[8][8]$_DFFE_PP_  (.CLK(clknet_leaf_259_clk),
    .RESET_B(net2763),
    .D(_01882_),
    .Q_N(_13514_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[8][8] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[8][9]$_DFFE_PP_  (.CLK(clknet_leaf_258_clk),
    .RESET_B(net2764),
    .D(_01883_),
    .Q_N(_13513_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[8][9] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[9][0]$_DFFE_PP_  (.CLK(clknet_leaf_265_clk),
    .RESET_B(net2765),
    .D(_01884_),
    .Q_N(_13512_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[9][0] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[9][10]$_DFFE_PP_  (.CLK(clknet_leaf_30_clk),
    .RESET_B(net2766),
    .D(_01885_),
    .Q_N(_13511_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[9][10] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[9][11]$_DFFE_PP_  (.CLK(clknet_leaf_267_clk),
    .RESET_B(net2767),
    .D(_01886_),
    .Q_N(_13510_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[9][11] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[9][1]$_DFFE_PP_  (.CLK(clknet_leaf_37_clk),
    .RESET_B(net2768),
    .D(_01887_),
    .Q_N(_13509_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[9][1] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[9][2]$_DFFE_PP_  (.CLK(clknet_leaf_31_clk),
    .RESET_B(net2769),
    .D(_01888_),
    .Q_N(_13508_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[9][2] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[9][3]$_DFFE_PP_  (.CLK(clknet_leaf_265_clk),
    .RESET_B(net2770),
    .D(_01889_),
    .Q_N(_13507_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[9][3] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[9][4]$_DFFE_PP_  (.CLK(clknet_leaf_264_clk),
    .RESET_B(net2771),
    .D(_01890_),
    .Q_N(_13506_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[9][4] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[9][5]$_DFFE_PP_  (.CLK(clknet_leaf_267_clk),
    .RESET_B(net2772),
    .D(_01891_),
    .Q_N(_13505_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[9][5] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[9][6]$_DFFE_PP_  (.CLK(clknet_leaf_37_clk),
    .RESET_B(net2773),
    .D(_01892_),
    .Q_N(_13504_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[9][6] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[9][7]$_DFFE_PP_  (.CLK(clknet_leaf_31_clk),
    .RESET_B(net2774),
    .D(_01893_),
    .Q_N(_13503_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[9][7] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[9][8]$_DFFE_PP_  (.CLK(clknet_leaf_259_clk),
    .RESET_B(net2775),
    .D(_01894_),
    .Q_N(_13502_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[9][8] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[9][9]$_DFFE_PP_  (.CLK(clknet_leaf_257_clk),
    .RESET_B(net2776),
    .D(_01895_),
    .Q_N(_13501_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[9][9] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_writeable_d[0]$_DFFE_PP_  (.CLK(clknet_leaf_252_clk),
    .RESET_B(net2777),
    .D(_01896_),
    .Q_N(_13500_),
    .Q(\cpu.genblk1.mmu.r_writeable_d[0] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_writeable_d[10]$_DFFE_PP_  (.CLK(clknet_leaf_253_clk),
    .RESET_B(net2778),
    .D(_01897_),
    .Q_N(_13499_),
    .Q(\cpu.genblk1.mmu.r_writeable_d[10] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_writeable_d[11]$_DFFE_PP_  (.CLK(clknet_leaf_252_clk),
    .RESET_B(net2779),
    .D(_01898_),
    .Q_N(_13498_),
    .Q(\cpu.genblk1.mmu.r_writeable_d[11] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_writeable_d[12]$_DFFE_PP_  (.CLK(clknet_leaf_254_clk),
    .RESET_B(net2780),
    .D(_01899_),
    .Q_N(_13497_),
    .Q(\cpu.genblk1.mmu.r_writeable_d[12] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_writeable_d[13]$_DFFE_PP_  (.CLK(clknet_leaf_254_clk),
    .RESET_B(net2781),
    .D(_01900_),
    .Q_N(_13496_),
    .Q(\cpu.genblk1.mmu.r_writeable_d[13] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_writeable_d[14]$_DFFE_PP_  (.CLK(clknet_leaf_253_clk),
    .RESET_B(net2782),
    .D(_01901_),
    .Q_N(_13495_),
    .Q(\cpu.genblk1.mmu.r_writeable_d[14] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_writeable_d[15]$_DFFE_PP_  (.CLK(clknet_leaf_252_clk),
    .RESET_B(net2783),
    .D(_01902_),
    .Q_N(_13494_),
    .Q(\cpu.genblk1.mmu.r_writeable_d[15] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_writeable_d[16]$_DFFE_PP_  (.CLK(clknet_leaf_234_clk),
    .RESET_B(net2784),
    .D(_01903_),
    .Q_N(_13493_),
    .Q(\cpu.genblk1.mmu.r_writeable_d[16] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_writeable_d[17]$_DFFE_PP_  (.CLK(clknet_leaf_240_clk),
    .RESET_B(net2785),
    .D(_01904_),
    .Q_N(_13492_),
    .Q(\cpu.genblk1.mmu.r_writeable_d[17] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_writeable_d[18]$_DFFE_PP_  (.CLK(clknet_leaf_234_clk),
    .RESET_B(net2786),
    .D(_01905_),
    .Q_N(_13491_),
    .Q(\cpu.genblk1.mmu.r_writeable_d[18] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_writeable_d[19]$_DFFE_PP_  (.CLK(clknet_leaf_234_clk),
    .RESET_B(net2787),
    .D(_01906_),
    .Q_N(_13490_),
    .Q(\cpu.genblk1.mmu.r_writeable_d[19] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_writeable_d[1]$_DFFE_PP_  (.CLK(clknet_leaf_239_clk),
    .RESET_B(net2788),
    .D(_01907_),
    .Q_N(_13489_),
    .Q(\cpu.genblk1.mmu.r_writeable_d[1] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_writeable_d[20]$_DFFE_PP_  (.CLK(clknet_leaf_234_clk),
    .RESET_B(net2789),
    .D(_01908_),
    .Q_N(_13488_),
    .Q(\cpu.genblk1.mmu.r_writeable_d[20] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_writeable_d[21]$_DFFE_PP_  (.CLK(clknet_leaf_238_clk),
    .RESET_B(net2790),
    .D(_01909_),
    .Q_N(_13487_),
    .Q(\cpu.genblk1.mmu.r_writeable_d[21] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_writeable_d[22]$_DFFE_PP_  (.CLK(clknet_leaf_234_clk),
    .RESET_B(net2791),
    .D(_01910_),
    .Q_N(_13486_),
    .Q(\cpu.genblk1.mmu.r_writeable_d[22] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_writeable_d[23]$_DFFE_PP_  (.CLK(clknet_leaf_239_clk),
    .RESET_B(net2792),
    .D(_01911_),
    .Q_N(_13485_),
    .Q(\cpu.genblk1.mmu.r_writeable_d[23] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_writeable_d[24]$_DFFE_PP_  (.CLK(clknet_leaf_239_clk),
    .RESET_B(net2793),
    .D(_01912_),
    .Q_N(_13484_),
    .Q(\cpu.genblk1.mmu.r_writeable_d[24] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_writeable_d[25]$_DFFE_PP_  (.CLK(clknet_leaf_239_clk),
    .RESET_B(net2794),
    .D(_01913_),
    .Q_N(_13483_),
    .Q(\cpu.genblk1.mmu.r_writeable_d[25] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_writeable_d[26]$_DFFE_PP_  (.CLK(clknet_leaf_235_clk),
    .RESET_B(net2795),
    .D(_01914_),
    .Q_N(_13482_),
    .Q(\cpu.genblk1.mmu.r_writeable_d[26] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_writeable_d[27]$_DFFE_PP_  (.CLK(clknet_leaf_235_clk),
    .RESET_B(net2796),
    .D(_01915_),
    .Q_N(_13481_),
    .Q(\cpu.genblk1.mmu.r_writeable_d[27] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_writeable_d[28]$_DFFE_PP_  (.CLK(clknet_leaf_238_clk),
    .RESET_B(net2797),
    .D(_01916_),
    .Q_N(_13480_),
    .Q(\cpu.genblk1.mmu.r_writeable_d[28] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_writeable_d[29]$_DFFE_PP_  (.CLK(clknet_leaf_238_clk),
    .RESET_B(net2798),
    .D(_01917_),
    .Q_N(_13479_),
    .Q(\cpu.genblk1.mmu.r_writeable_d[29] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_writeable_d[2]$_DFFE_PP_  (.CLK(clknet_leaf_251_clk),
    .RESET_B(net2799),
    .D(_01918_),
    .Q_N(_13478_),
    .Q(\cpu.genblk1.mmu.r_writeable_d[2] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_writeable_d[30]$_DFFE_PP_  (.CLK(clknet_leaf_234_clk),
    .RESET_B(net2800),
    .D(_01919_),
    .Q_N(_13477_),
    .Q(\cpu.genblk1.mmu.r_writeable_d[30] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_writeable_d[31]$_DFFE_PP_  (.CLK(clknet_leaf_235_clk),
    .RESET_B(net2801),
    .D(_01920_),
    .Q_N(_13476_),
    .Q(\cpu.genblk1.mmu.r_writeable_d[31] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_writeable_d[3]$_DFFE_PP_  (.CLK(clknet_leaf_239_clk),
    .RESET_B(net2802),
    .D(_01921_),
    .Q_N(_13475_),
    .Q(\cpu.genblk1.mmu.r_writeable_d[3] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_writeable_d[4]$_DFFE_PP_  (.CLK(clknet_leaf_234_clk),
    .RESET_B(net2803),
    .D(_01922_),
    .Q_N(_13474_),
    .Q(\cpu.genblk1.mmu.r_writeable_d[4] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_writeable_d[5]$_DFFE_PP_  (.CLK(clknet_leaf_240_clk),
    .RESET_B(net2804),
    .D(_01923_),
    .Q_N(_13473_),
    .Q(\cpu.genblk1.mmu.r_writeable_d[5] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_writeable_d[6]$_DFFE_PP_  (.CLK(clknet_leaf_252_clk),
    .RESET_B(net2805),
    .D(_01924_),
    .Q_N(_13472_),
    .Q(\cpu.genblk1.mmu.r_writeable_d[6] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_writeable_d[7]$_DFFE_PP_  (.CLK(clknet_leaf_239_clk),
    .RESET_B(net2806),
    .D(_01925_),
    .Q_N(_13471_),
    .Q(\cpu.genblk1.mmu.r_writeable_d[7] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_writeable_d[8]$_DFFE_PP_  (.CLK(clknet_leaf_255_clk),
    .RESET_B(net2807),
    .D(_01926_),
    .Q_N(_13470_),
    .Q(\cpu.genblk1.mmu.r_writeable_d[8] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_writeable_d[9]$_DFFE_PP_  (.CLK(clknet_leaf_254_clk),
    .RESET_B(net2808),
    .D(_01927_),
    .Q_N(_13469_),
    .Q(\cpu.genblk1.mmu.r_writeable_d[9] ));
 sg13g2_dfrbp_1 \cpu.gpio.r_enable_in[0]$_SDFFE_PN0P_  (.CLK(clknet_leaf_84_clk),
    .RESET_B(net2809),
    .D(_01928_),
    .Q_N(_13468_),
    .Q(\cpu.gpio.r_enable_in[0] ));
 sg13g2_dfrbp_1 \cpu.gpio.r_enable_in[1]$_SDFFE_PN0P_  (.CLK(clknet_leaf_84_clk),
    .RESET_B(net2810),
    .D(_01929_),
    .Q_N(_13467_),
    .Q(\cpu.gpio.r_enable_in[1] ));
 sg13g2_dfrbp_1 \cpu.gpio.r_enable_in[2]$_SDFFE_PN0P_  (.CLK(clknet_leaf_68_clk),
    .RESET_B(net2811),
    .D(_01930_),
    .Q_N(_13466_),
    .Q(\cpu.gpio.r_enable_in[2] ));
 sg13g2_dfrbp_1 \cpu.gpio.r_enable_in[3]$_SDFFE_PN0P_  (.CLK(clknet_leaf_68_clk),
    .RESET_B(net2812),
    .D(_01931_),
    .Q_N(_13465_),
    .Q(\cpu.gpio.r_enable_in[3] ));
 sg13g2_dfrbp_1 \cpu.gpio.r_enable_in[4]$_SDFFE_PN0P_  (.CLK(clknet_leaf_68_clk),
    .RESET_B(net2813),
    .D(_01932_),
    .Q_N(_13464_),
    .Q(\cpu.gpio.r_enable_in[4] ));
 sg13g2_dfrbp_1 \cpu.gpio.r_enable_in[5]$_SDFFE_PN0P_  (.CLK(clknet_leaf_68_clk),
    .RESET_B(net2814),
    .D(_01933_),
    .Q_N(_13463_),
    .Q(\cpu.gpio.r_enable_in[5] ));
 sg13g2_dfrbp_1 \cpu.gpio.r_enable_in[6]$_SDFFE_PN0P_  (.CLK(clknet_leaf_67_clk),
    .RESET_B(net2815),
    .D(_01934_),
    .Q_N(_13462_),
    .Q(\cpu.gpio.r_enable_in[6] ));
 sg13g2_dfrbp_1 \cpu.gpio.r_enable_in[7]$_SDFFE_PN0P_  (.CLK(clknet_leaf_67_clk),
    .RESET_B(net2816),
    .D(_01935_),
    .Q_N(_13461_),
    .Q(\cpu.gpio.r_enable_in[7] ));
 sg13g2_dfrbp_1 \cpu.gpio.r_enable_io[0]$_SDFFE_PN0P_  (.CLK(clknet_leaf_65_clk),
    .RESET_B(net2817),
    .D(_01936_),
    .Q_N(_13460_),
    .Q(\cpu.gpio.r_enable_io[4] ));
 sg13g2_dfrbp_1 \cpu.gpio.r_enable_io[1]$_SDFFE_PN0P_  (.CLK(clknet_leaf_67_clk),
    .RESET_B(net2818),
    .D(_01937_),
    .Q_N(_13459_),
    .Q(\cpu.gpio.r_enable_io[5] ));
 sg13g2_dfrbp_1 \cpu.gpio.r_enable_io[2]$_SDFFE_PN0P_  (.CLK(clknet_leaf_65_clk),
    .RESET_B(net2819),
    .D(_01938_),
    .Q_N(_13458_),
    .Q(\cpu.gpio.r_enable_io[6] ));
 sg13g2_dfrbp_1 \cpu.gpio.r_enable_io[3]$_SDFFE_PN0P_  (.CLK(clknet_leaf_67_clk),
    .RESET_B(net2820),
    .D(_01939_),
    .Q_N(_13457_),
    .Q(\cpu.gpio.r_enable_io[7] ));
 sg13g2_dfrbp_1 \cpu.gpio.r_gpio_en[0]$_SDFFE_PN0P_  (.CLK(clknet_leaf_65_clk),
    .RESET_B(net2821),
    .D(_01940_),
    .Q_N(_13456_),
    .Q(net7));
 sg13g2_dfrbp_1 \cpu.gpio.r_gpio_en[1]$_SDFFE_PN0P_  (.CLK(clknet_leaf_65_clk),
    .RESET_B(net2822),
    .D(_01941_),
    .Q_N(_13455_),
    .Q(net8));
 sg13g2_dfrbp_1 \cpu.gpio.r_gpio_en[2]$_SDFFE_PN0P_  (.CLK(clknet_leaf_65_clk),
    .RESET_B(net2823),
    .D(_01942_),
    .Q_N(_13454_),
    .Q(net9));
 sg13g2_dfrbp_1 \cpu.gpio.r_gpio_en[3]$_SDFFE_PN0P_  (.CLK(clknet_leaf_65_clk),
    .RESET_B(net2824),
    .D(_01943_),
    .Q_N(_13453_),
    .Q(net10));
 sg13g2_dfrbp_1 \cpu.gpio.r_gpio_io[0]$_DFFE_PP_  (.CLK(clknet_leaf_69_clk),
    .RESET_B(net2825),
    .D(_01944_),
    .Q_N(_13452_),
    .Q(\cpu.gpio.genblk2[4].srcs_io[0] ));
 sg13g2_dfrbp_1 \cpu.gpio.r_gpio_io[1]$_DFFE_PP_  (.CLK(clknet_leaf_68_clk),
    .RESET_B(net2826),
    .D(_01945_),
    .Q_N(_13451_),
    .Q(\cpu.gpio.genblk2[5].srcs_io[0] ));
 sg13g2_dfrbp_1 \cpu.gpio.r_gpio_io[2]$_DFFE_PP_  (.CLK(clknet_leaf_63_clk),
    .RESET_B(net2827),
    .D(_01946_),
    .Q_N(_13450_),
    .Q(\cpu.gpio.genblk2[6].srcs_io[0] ));
 sg13g2_dfrbp_1 \cpu.gpio.r_gpio_io[3]$_DFFE_PP_  (.CLK(clknet_leaf_69_clk),
    .RESET_B(net2828),
    .D(_01947_),
    .Q_N(_13449_),
    .Q(\cpu.gpio.genblk2[7].srcs_io[0] ));
 sg13g2_dfrbp_1 \cpu.gpio.r_gpio_o[0]$_DFFE_PP_  (.CLK(clknet_leaf_63_clk),
    .RESET_B(net2829),
    .D(_01948_),
    .Q_N(_13448_),
    .Q(\cpu.gpio.genblk1[3].srcs_o[0] ));
 sg13g2_dfrbp_1 \cpu.gpio.r_gpio_o[1]$_DFFE_PP_  (.CLK(clknet_leaf_73_clk),
    .RESET_B(net2830),
    .D(_01949_),
    .Q_N(_13447_),
    .Q(\cpu.gpio.genblk1[4].srcs_o[0] ));
 sg13g2_dfrbp_1 \cpu.gpio.r_gpio_o[2]$_DFFE_PP_  (.CLK(clknet_leaf_77_clk),
    .RESET_B(net2831),
    .D(_01950_),
    .Q_N(_13446_),
    .Q(\cpu.gpio.genblk1[5].srcs_o[0] ));
 sg13g2_dfrbp_1 \cpu.gpio.r_gpio_o[3]$_DFFE_PP_  (.CLK(clknet_leaf_69_clk),
    .RESET_B(net2832),
    .D(_01951_),
    .Q_N(_13445_),
    .Q(\cpu.gpio.genblk1[6].srcs_o[0] ));
 sg13g2_dfrbp_1 \cpu.gpio.r_gpio_o[4]$_DFFE_PP_  (.CLK(clknet_leaf_73_clk),
    .RESET_B(net2833),
    .D(_01952_),
    .Q_N(_13444_),
    .Q(\cpu.gpio.genblk1[7].srcs_o[0] ));
 sg13g2_dfrbp_1 \cpu.gpio.r_spi_miso_src[0][0]$_DFFE_PP_  (.CLK(clknet_leaf_78_clk),
    .RESET_B(net2834),
    .D(_01953_),
    .Q_N(_13443_),
    .Q(\cpu.gpio.r_spi_miso_src[0][0] ));
 sg13g2_dfrbp_1 \cpu.gpio.r_spi_miso_src[0][1]$_DFFE_PP_  (.CLK(clknet_leaf_79_clk),
    .RESET_B(net2835),
    .D(_01954_),
    .Q_N(_00096_),
    .Q(\cpu.gpio.r_spi_miso_src[0][1] ));
 sg13g2_dfrbp_1 \cpu.gpio.r_spi_miso_src[0][2]$_DFFE_PP_  (.CLK(clknet_leaf_79_clk),
    .RESET_B(net2836),
    .D(_01955_),
    .Q_N(_00106_),
    .Q(\cpu.gpio.r_spi_miso_src[0][2] ));
 sg13g2_dfrbp_1 \cpu.gpio.r_spi_miso_src[0][3]$_DFFE_PP_  (.CLK(clknet_leaf_77_clk),
    .RESET_B(net2837),
    .D(_01956_),
    .Q_N(_00115_),
    .Q(\cpu.gpio.r_spi_miso_src[0][3] ));
 sg13g2_dfrbp_1 \cpu.gpio.r_spi_miso_src[1][0]$_DFFE_PP_  (.CLK(clknet_leaf_78_clk),
    .RESET_B(net2838),
    .D(_01957_),
    .Q_N(_13442_),
    .Q(\cpu.gpio.r_spi_miso_src[1][0] ));
 sg13g2_dfrbp_1 \cpu.gpio.r_spi_miso_src[1][1]$_DFFE_PP_  (.CLK(clknet_leaf_78_clk),
    .RESET_B(net2839),
    .D(_01958_),
    .Q_N(_00132_),
    .Q(\cpu.gpio.r_spi_miso_src[1][1] ));
 sg13g2_dfrbp_1 \cpu.gpio.r_spi_miso_src[1][2]$_DFFE_PP_  (.CLK(clknet_leaf_78_clk),
    .RESET_B(net2840),
    .D(_01959_),
    .Q_N(_00143_),
    .Q(\cpu.gpio.r_spi_miso_src[1][2] ));
 sg13g2_dfrbp_1 \cpu.gpio.r_spi_miso_src[1][3]$_DFFE_PP_  (.CLK(clknet_leaf_78_clk),
    .RESET_B(net2841),
    .D(_01960_),
    .Q_N(_00154_),
    .Q(\cpu.gpio.r_spi_miso_src[1][3] ));
 sg13g2_dfrbp_1 \cpu.gpio.r_src_io[4][0]$_DFFE_PP_  (.CLK(clknet_leaf_76_clk),
    .RESET_B(net2842),
    .D(_01961_),
    .Q_N(_13441_),
    .Q(\cpu.gpio.r_src_io[4][0] ));
 sg13g2_dfrbp_1 \cpu.gpio.r_src_io[4][1]$_DFFE_PP_  (.CLK(clknet_leaf_76_clk),
    .RESET_B(net2843),
    .D(_01962_),
    .Q_N(_13440_),
    .Q(\cpu.gpio.r_src_io[4][1] ));
 sg13g2_dfrbp_1 \cpu.gpio.r_src_io[4][2]$_DFFE_PP_  (.CLK(clknet_leaf_74_clk),
    .RESET_B(net2844),
    .D(_01963_),
    .Q_N(_00177_),
    .Q(\cpu.gpio.r_src_io[4][2] ));
 sg13g2_dfrbp_1 \cpu.gpio.r_src_io[4][3]$_DFFE_PP_  (.CLK(clknet_leaf_76_clk),
    .RESET_B(net2845),
    .D(_01964_),
    .Q_N(_13439_),
    .Q(\cpu.gpio.r_src_io[4][3] ));
 sg13g2_dfrbp_1 \cpu.gpio.r_src_io[5][0]$_DFFE_PP_  (.CLK(clknet_leaf_73_clk),
    .RESET_B(net2846),
    .D(_01965_),
    .Q_N(_13438_),
    .Q(\cpu.gpio.r_src_io[5][0] ));
 sg13g2_dfrbp_1 \cpu.gpio.r_src_io[5][1]$_DFFE_PP_  (.CLK(clknet_leaf_73_clk),
    .RESET_B(net2847),
    .D(_01966_),
    .Q_N(_13437_),
    .Q(\cpu.gpio.r_src_io[5][1] ));
 sg13g2_dfrbp_1 \cpu.gpio.r_src_io[5][2]$_DFFE_PP_  (.CLK(clknet_leaf_73_clk),
    .RESET_B(net2848),
    .D(_01967_),
    .Q_N(_00176_),
    .Q(\cpu.gpio.r_src_io[5][2] ));
 sg13g2_dfrbp_1 \cpu.gpio.r_src_io[5][3]$_DFFE_PP_  (.CLK(clknet_leaf_76_clk),
    .RESET_B(net2849),
    .D(_01968_),
    .Q_N(_13436_),
    .Q(\cpu.gpio.r_src_io[5][3] ));
 sg13g2_dfrbp_1 \cpu.gpio.r_src_io[6][0]$_DFFE_PP_  (.CLK(clknet_leaf_63_clk),
    .RESET_B(net2850),
    .D(_01969_),
    .Q_N(_13435_),
    .Q(\cpu.gpio.r_src_io[6][0] ));
 sg13g2_dfrbp_1 \cpu.gpio.r_src_io[6][1]$_DFFE_PP_  (.CLK(clknet_leaf_63_clk),
    .RESET_B(net2851),
    .D(_01970_),
    .Q_N(_00092_),
    .Q(\cpu.gpio.r_src_io[6][1] ));
 sg13g2_dfrbp_1 \cpu.gpio.r_src_io[6][2]$_DFFE_PP_  (.CLK(clknet_leaf_63_clk),
    .RESET_B(net2852),
    .D(_01971_),
    .Q_N(_00102_),
    .Q(\cpu.gpio.r_src_io[6][2] ));
 sg13g2_dfrbp_1 \cpu.gpio.r_src_io[6][3]$_DFFE_PP_  (.CLK(clknet_leaf_63_clk),
    .RESET_B(net2853),
    .D(_01972_),
    .Q_N(_00112_),
    .Q(\cpu.gpio.r_src_io[6][3] ));
 sg13g2_dfrbp_1 \cpu.gpio.r_src_io[7][0]$_DFFE_PP_  (.CLK(clknet_leaf_69_clk),
    .RESET_B(net2854),
    .D(_01973_),
    .Q_N(_13434_),
    .Q(\cpu.gpio.r_src_io[7][0] ));
 sg13g2_dfrbp_1 \cpu.gpio.r_src_io[7][1]$_DFFE_PP_  (.CLK(clknet_leaf_69_clk),
    .RESET_B(net2855),
    .D(_01974_),
    .Q_N(_00128_),
    .Q(\cpu.gpio.r_src_io[7][1] ));
 sg13g2_dfrbp_1 \cpu.gpio.r_src_io[7][2]$_DFFE_PP_  (.CLK(clknet_leaf_69_clk),
    .RESET_B(net2856),
    .D(_01975_),
    .Q_N(_00139_),
    .Q(\cpu.gpio.r_src_io[7][2] ));
 sg13g2_dfrbp_1 \cpu.gpio.r_src_io[7][3]$_DFFE_PP_  (.CLK(clknet_leaf_69_clk),
    .RESET_B(net2857),
    .D(_01976_),
    .Q_N(_00150_),
    .Q(\cpu.gpio.r_src_io[7][3] ));
 sg13g2_dfrbp_1 \cpu.gpio.r_src_o[3][0]$_DFFE_PP_  (.CLK(clknet_leaf_64_clk),
    .RESET_B(net2858),
    .D(_01977_),
    .Q_N(_13433_),
    .Q(\cpu.gpio.r_src_o[3][0] ));
 sg13g2_dfrbp_1 \cpu.gpio.r_src_o[3][1]$_DFFE_PP_  (.CLK(clknet_leaf_64_clk),
    .RESET_B(net2859),
    .D(_01978_),
    .Q_N(_00131_),
    .Q(\cpu.gpio.r_src_o[3][1] ));
 sg13g2_dfrbp_1 \cpu.gpio.r_src_o[3][2]$_DFFE_PP_  (.CLK(clknet_leaf_64_clk),
    .RESET_B(net2860),
    .D(_01979_),
    .Q_N(_00142_),
    .Q(\cpu.gpio.r_src_o[3][2] ));
 sg13g2_dfrbp_1 \cpu.gpio.r_src_o[3][3]$_DFFE_PP_  (.CLK(clknet_leaf_64_clk),
    .RESET_B(net2861),
    .D(_01980_),
    .Q_N(_00153_),
    .Q(\cpu.gpio.r_src_o[3][3] ));
 sg13g2_dfrbp_1 \cpu.gpio.r_src_o[4][0]$_DFFE_PP_  (.CLK(clknet_leaf_76_clk),
    .RESET_B(net2862),
    .D(_01981_),
    .Q_N(_13432_),
    .Q(\cpu.gpio.r_src_o[4][0] ));
 sg13g2_dfrbp_1 \cpu.gpio.r_src_o[4][1]$_DFFE_PP_  (.CLK(clknet_leaf_77_clk),
    .RESET_B(net2863),
    .D(_01982_),
    .Q_N(_00094_),
    .Q(\cpu.gpio.r_src_o[4][1] ));
 sg13g2_dfrbp_1 \cpu.gpio.r_src_o[4][2]$_DFFE_PP_  (.CLK(clknet_leaf_77_clk),
    .RESET_B(net2864),
    .D(_01983_),
    .Q_N(_00104_),
    .Q(\cpu.gpio.r_src_o[4][2] ));
 sg13g2_dfrbp_1 \cpu.gpio.r_src_o[4][3]$_DFFE_PP_  (.CLK(clknet_leaf_77_clk),
    .RESET_B(net2865),
    .D(_01984_),
    .Q_N(_00114_),
    .Q(\cpu.gpio.r_src_o[4][3] ));
 sg13g2_dfrbp_1 \cpu.gpio.r_src_o[5][0]$_DFFE_PP_  (.CLK(clknet_leaf_76_clk),
    .RESET_B(net2866),
    .D(_01985_),
    .Q_N(_13431_),
    .Q(\cpu.gpio.r_src_o[5][0] ));
 sg13g2_dfrbp_1 \cpu.gpio.r_src_o[5][1]$_DFFE_PP_  (.CLK(clknet_leaf_78_clk),
    .RESET_B(net2867),
    .D(_01986_),
    .Q_N(_00130_),
    .Q(\cpu.gpio.r_src_o[5][1] ));
 sg13g2_dfrbp_1 \cpu.gpio.r_src_o[5][2]$_DFFE_PP_  (.CLK(clknet_leaf_77_clk),
    .RESET_B(net2868),
    .D(_01987_),
    .Q_N(_00141_),
    .Q(\cpu.gpio.r_src_o[5][2] ));
 sg13g2_dfrbp_1 \cpu.gpio.r_src_o[5][3]$_DFFE_PP_  (.CLK(clknet_leaf_77_clk),
    .RESET_B(net2869),
    .D(_01988_),
    .Q_N(_00152_),
    .Q(\cpu.gpio.r_src_o[5][3] ));
 sg13g2_dfrbp_1 \cpu.gpio.r_src_o[6][0]$_SDFFE_PN1P_  (.CLK(clknet_leaf_73_clk),
    .RESET_B(net2870),
    .D(_01989_),
    .Q_N(_13430_),
    .Q(\cpu.gpio.r_src_o[6][0] ));
 sg13g2_dfrbp_1 \cpu.gpio.r_src_o[6][1]$_SDFFE_PN0P_  (.CLK(clknet_leaf_68_clk),
    .RESET_B(net2871),
    .D(_01990_),
    .Q_N(_00093_),
    .Q(\cpu.gpio.r_src_o[6][1] ));
 sg13g2_dfrbp_1 \cpu.gpio.r_src_o[6][2]$_SDFFE_PN0P_  (.CLK(clknet_leaf_68_clk),
    .RESET_B(net2872),
    .D(_01991_),
    .Q_N(_00103_),
    .Q(\cpu.gpio.r_src_o[6][2] ));
 sg13g2_dfrbp_1 \cpu.gpio.r_src_o[6][3]$_SDFFE_PN0P_  (.CLK(clknet_leaf_68_clk),
    .RESET_B(net2873),
    .D(_01992_),
    .Q_N(_00113_),
    .Q(\cpu.gpio.r_src_o[6][3] ));
 sg13g2_dfrbp_1 \cpu.gpio.r_src_o[7][0]$_DFFE_PP_  (.CLK(clknet_leaf_76_clk),
    .RESET_B(net2874),
    .D(_01993_),
    .Q_N(_13429_),
    .Q(\cpu.gpio.r_src_o[7][0] ));
 sg13g2_dfrbp_1 \cpu.gpio.r_src_o[7][1]$_DFFE_PP_  (.CLK(clknet_leaf_73_clk),
    .RESET_B(net2875),
    .D(_01994_),
    .Q_N(_00129_),
    .Q(\cpu.gpio.r_src_o[7][1] ));
 sg13g2_dfrbp_1 \cpu.gpio.r_src_o[7][2]$_DFFE_PP_  (.CLK(clknet_leaf_77_clk),
    .RESET_B(net2876),
    .D(_01995_),
    .Q_N(_00140_),
    .Q(\cpu.gpio.r_src_o[7][2] ));
 sg13g2_dfrbp_1 \cpu.gpio.r_src_o[7][3]$_DFFE_PP_  (.CLK(clknet_leaf_76_clk),
    .RESET_B(net2877),
    .D(_01996_),
    .Q_N(_00151_),
    .Q(\cpu.gpio.r_src_o[7][3] ));
 sg13g2_dfrbp_1 \cpu.gpio.r_uart_rx_src[0]$_SDFFE_PN0P_  (.CLK(clknet_leaf_83_clk),
    .RESET_B(net2878),
    .D(_01997_),
    .Q_N(_13428_),
    .Q(\cpu.gpio.r_uart_rx_src[0] ));
 sg13g2_dfrbp_1 \cpu.gpio.r_uart_rx_src[1]$_SDFFE_PN0P_  (.CLK(clknet_leaf_83_clk),
    .RESET_B(net2879),
    .D(_01998_),
    .Q_N(_00095_),
    .Q(\cpu.gpio.r_uart_rx_src[1] ));
 sg13g2_dfrbp_1 \cpu.gpio.r_uart_rx_src[2]$_SDFFE_PN0P_  (.CLK(clknet_leaf_83_clk),
    .RESET_B(net2880),
    .D(_01999_),
    .Q_N(_00105_),
    .Q(\cpu.gpio.r_uart_rx_src[2] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[0][0]$_DFFE_PP_  (.CLK(clknet_leaf_214_clk),
    .RESET_B(net2881),
    .D(_02000_),
    .Q_N(_13427_),
    .Q(\cpu.icache.r_data[0][0] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[0][10]$_DFFE_PP_  (.CLK(clknet_leaf_167_clk),
    .RESET_B(net2882),
    .D(_02001_),
    .Q_N(_00191_),
    .Q(\cpu.icache.r_data[0][10] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[0][11]$_DFFE_PP_  (.CLK(clknet_leaf_167_clk),
    .RESET_B(net2883),
    .D(_02002_),
    .Q_N(_00193_),
    .Q(\cpu.icache.r_data[0][11] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[0][12]$_DFFE_PP_  (.CLK(clknet_leaf_189_clk),
    .RESET_B(net2884),
    .D(_02003_),
    .Q_N(_00203_),
    .Q(\cpu.icache.r_data[0][12] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[0][13]$_DFFE_PP_  (.CLK(clknet_leaf_189_clk),
    .RESET_B(net2885),
    .D(_02004_),
    .Q_N(_13426_),
    .Q(\cpu.icache.r_data[0][13] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[0][14]$_DFFE_PP_  (.CLK(clknet_leaf_189_clk),
    .RESET_B(net2886),
    .D(_02005_),
    .Q_N(_00195_),
    .Q(\cpu.icache.r_data[0][14] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[0][15]$_DFFE_PP_  (.CLK(clknet_leaf_208_clk),
    .RESET_B(net2887),
    .D(_02006_),
    .Q_N(_00197_),
    .Q(\cpu.icache.r_data[0][15] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[0][16]$_DFFE_PP_  (.CLK(clknet_leaf_214_clk),
    .RESET_B(net2888),
    .D(_02007_),
    .Q_N(_13425_),
    .Q(\cpu.icache.r_data[0][16] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[0][17]$_DFFE_PP_  (.CLK(clknet_leaf_228_clk),
    .RESET_B(net2889),
    .D(_02008_),
    .Q_N(_13424_),
    .Q(\cpu.icache.r_data[0][17] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[0][18]$_DFFE_PP_  (.CLK(clknet_leaf_212_clk),
    .RESET_B(net2890),
    .D(_02009_),
    .Q_N(_00163_),
    .Q(\cpu.icache.r_data[0][18] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[0][19]$_DFFE_PP_  (.CLK(clknet_leaf_228_clk),
    .RESET_B(net2891),
    .D(_02010_),
    .Q_N(_00165_),
    .Q(\cpu.icache.r_data[0][19] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[0][1]$_DFFE_PP_  (.CLK(clknet_leaf_213_clk),
    .RESET_B(net2892),
    .D(_02011_),
    .Q_N(_13423_),
    .Q(\cpu.icache.r_data[0][1] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[0][20]$_DFFE_PP_  (.CLK(clknet_leaf_195_clk),
    .RESET_B(net2893),
    .D(_02012_),
    .Q_N(_00167_),
    .Q(\cpu.icache.r_data[0][20] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[0][21]$_DFFE_PP_  (.CLK(clknet_leaf_194_clk),
    .RESET_B(net2894),
    .D(_02013_),
    .Q_N(_00200_),
    .Q(\cpu.icache.r_data[0][21] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[0][22]$_DFFE_PP_  (.CLK(clknet_leaf_196_clk),
    .RESET_B(net2895),
    .D(_02014_),
    .Q_N(_00202_),
    .Q(\cpu.icache.r_data[0][22] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[0][23]$_DFFE_PP_  (.CLK(clknet_leaf_196_clk),
    .RESET_B(net2896),
    .D(_02015_),
    .Q_N(_00157_),
    .Q(\cpu.icache.r_data[0][23] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[0][24]$_DFFE_PP_  (.CLK(clknet_leaf_167_clk),
    .RESET_B(net2897),
    .D(_02016_),
    .Q_N(_00159_),
    .Q(\cpu.icache.r_data[0][24] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[0][25]$_DFFE_PP_  (.CLK(clknet_leaf_170_clk),
    .RESET_B(net2898),
    .D(_02017_),
    .Q_N(_00161_),
    .Q(\cpu.icache.r_data[0][25] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[0][26]$_DFFE_PP_  (.CLK(clknet_leaf_167_clk),
    .RESET_B(net2899),
    .D(_02018_),
    .Q_N(_00192_),
    .Q(\cpu.icache.r_data[0][26] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[0][27]$_DFFE_PP_  (.CLK(clknet_leaf_165_clk),
    .RESET_B(net2900),
    .D(_02019_),
    .Q_N(_00194_),
    .Q(\cpu.icache.r_data[0][27] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[0][28]$_DFFE_PP_  (.CLK(clknet_leaf_209_clk),
    .RESET_B(net2901),
    .D(_02020_),
    .Q_N(_00204_),
    .Q(\cpu.icache.r_data[0][28] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[0][29]$_DFFE_PP_  (.CLK(clknet_leaf_208_clk),
    .RESET_B(net2902),
    .D(_02021_),
    .Q_N(_13422_),
    .Q(\cpu.icache.r_data[0][29] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[0][2]$_DFFE_PP_  (.CLK(clknet_leaf_212_clk),
    .RESET_B(net2903),
    .D(_02022_),
    .Q_N(_00162_),
    .Q(\cpu.icache.r_data[0][2] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[0][30]$_DFFE_PP_  (.CLK(clknet_leaf_209_clk),
    .RESET_B(net2904),
    .D(_02023_),
    .Q_N(_00196_),
    .Q(\cpu.icache.r_data[0][30] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[0][31]$_DFFE_PP_  (.CLK(clknet_leaf_209_clk),
    .RESET_B(net2905),
    .D(_02024_),
    .Q_N(_00198_),
    .Q(\cpu.icache.r_data[0][31] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[0][3]$_DFFE_PP_  (.CLK(clknet_leaf_213_clk),
    .RESET_B(net2906),
    .D(_02025_),
    .Q_N(_00164_),
    .Q(\cpu.icache.r_data[0][3] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[0][4]$_DFFE_PP_  (.CLK(clknet_leaf_194_clk),
    .RESET_B(net2907),
    .D(_02026_),
    .Q_N(_00166_),
    .Q(\cpu.icache.r_data[0][4] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[0][5]$_DFFE_PP_  (.CLK(clknet_leaf_194_clk),
    .RESET_B(net2908),
    .D(_02027_),
    .Q_N(_00199_),
    .Q(\cpu.icache.r_data[0][5] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[0][6]$_DFFE_PP_  (.CLK(clknet_leaf_194_clk),
    .RESET_B(net2909),
    .D(_02028_),
    .Q_N(_00201_),
    .Q(\cpu.icache.r_data[0][6] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[0][7]$_DFFE_PP_  (.CLK(clknet_leaf_195_clk),
    .RESET_B(net2910),
    .D(_02029_),
    .Q_N(_00156_),
    .Q(\cpu.icache.r_data[0][7] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[0][8]$_DFFE_PP_  (.CLK(clknet_leaf_166_clk),
    .RESET_B(net2911),
    .D(_02030_),
    .Q_N(_00158_),
    .Q(\cpu.icache.r_data[0][8] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[0][9]$_DFFE_PP_  (.CLK(clknet_leaf_166_clk),
    .RESET_B(net2912),
    .D(_02031_),
    .Q_N(_00160_),
    .Q(\cpu.icache.r_data[0][9] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[1][0]$_DFFE_PP_  (.CLK(clknet_leaf_220_clk),
    .RESET_B(net2913),
    .D(_02032_),
    .Q_N(_13421_),
    .Q(\cpu.icache.r_data[1][0] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[1][10]$_DFFE_PP_  (.CLK(clknet_leaf_166_clk),
    .RESET_B(net2914),
    .D(_02033_),
    .Q_N(_13420_),
    .Q(\cpu.icache.r_data[1][10] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[1][11]$_DFFE_PP_  (.CLK(clknet_leaf_160_clk),
    .RESET_B(net2915),
    .D(_02034_),
    .Q_N(_13419_),
    .Q(\cpu.icache.r_data[1][11] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[1][12]$_DFFE_PP_  (.CLK(clknet_leaf_207_clk),
    .RESET_B(net2916),
    .D(_02035_),
    .Q_N(_13418_),
    .Q(\cpu.icache.r_data[1][12] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[1][13]$_DFFE_PP_  (.CLK(clknet_leaf_206_clk),
    .RESET_B(net2917),
    .D(_02036_),
    .Q_N(_13417_),
    .Q(\cpu.icache.r_data[1][13] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[1][14]$_DFFE_PP_  (.CLK(clknet_leaf_207_clk),
    .RESET_B(net2918),
    .D(_02037_),
    .Q_N(_13416_),
    .Q(\cpu.icache.r_data[1][14] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[1][15]$_DFFE_PP_  (.CLK(clknet_leaf_206_clk),
    .RESET_B(net2919),
    .D(_02038_),
    .Q_N(_13415_),
    .Q(\cpu.icache.r_data[1][15] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[1][16]$_DFFE_PP_  (.CLK(clknet_leaf_215_clk),
    .RESET_B(net2920),
    .D(_02039_),
    .Q_N(_13414_),
    .Q(\cpu.icache.r_data[1][16] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[1][17]$_DFFE_PP_  (.CLK(clknet_leaf_219_clk),
    .RESET_B(net2921),
    .D(_02040_),
    .Q_N(_13413_),
    .Q(\cpu.icache.r_data[1][17] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[1][18]$_DFFE_PP_  (.CLK(clknet_leaf_215_clk),
    .RESET_B(net2922),
    .D(_02041_),
    .Q_N(_13412_),
    .Q(\cpu.icache.r_data[1][18] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[1][19]$_DFFE_PP_  (.CLK(clknet_leaf_214_clk),
    .RESET_B(net2923),
    .D(_02042_),
    .Q_N(_13411_),
    .Q(\cpu.icache.r_data[1][19] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[1][1]$_DFFE_PP_  (.CLK(clknet_leaf_219_clk),
    .RESET_B(net2924),
    .D(_02043_),
    .Q_N(_13410_),
    .Q(\cpu.icache.r_data[1][1] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[1][20]$_DFFE_PP_  (.CLK(clknet_leaf_195_clk),
    .RESET_B(net2925),
    .D(_02044_),
    .Q_N(_13409_),
    .Q(\cpu.icache.r_data[1][20] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[1][21]$_DFFE_PP_  (.CLK(clknet_leaf_196_clk),
    .RESET_B(net2926),
    .D(_02045_),
    .Q_N(_13408_),
    .Q(\cpu.icache.r_data[1][21] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[1][22]$_DFFE_PP_  (.CLK(clknet_leaf_196_clk),
    .RESET_B(net2927),
    .D(_02046_),
    .Q_N(_13407_),
    .Q(\cpu.icache.r_data[1][22] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[1][23]$_DFFE_PP_  (.CLK(clknet_leaf_195_clk),
    .RESET_B(net2928),
    .D(_02047_),
    .Q_N(_13406_),
    .Q(\cpu.icache.r_data[1][23] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[1][24]$_DFFE_PP_  (.CLK(clknet_leaf_160_clk),
    .RESET_B(net2929),
    .D(_02048_),
    .Q_N(_13405_),
    .Q(\cpu.icache.r_data[1][24] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[1][25]$_DFFE_PP_  (.CLK(clknet_leaf_160_clk),
    .RESET_B(net2930),
    .D(_02049_),
    .Q_N(_13404_),
    .Q(\cpu.icache.r_data[1][25] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[1][26]$_DFFE_PP_  (.CLK(clknet_leaf_165_clk),
    .RESET_B(net2931),
    .D(_02050_),
    .Q_N(_13403_),
    .Q(\cpu.icache.r_data[1][26] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[1][27]$_DFFE_PP_  (.CLK(clknet_leaf_166_clk),
    .RESET_B(net2932),
    .D(_02051_),
    .Q_N(_13402_),
    .Q(\cpu.icache.r_data[1][27] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[1][28]$_DFFE_PP_  (.CLK(clknet_leaf_202_clk),
    .RESET_B(net2933),
    .D(_02052_),
    .Q_N(_13401_),
    .Q(\cpu.icache.r_data[1][28] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[1][29]$_DFFE_PP_  (.CLK(clknet_leaf_207_clk),
    .RESET_B(net2934),
    .D(_02053_),
    .Q_N(_13400_),
    .Q(\cpu.icache.r_data[1][29] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[1][2]$_DFFE_PP_  (.CLK(clknet_leaf_216_clk),
    .RESET_B(net2935),
    .D(_02054_),
    .Q_N(_13399_),
    .Q(\cpu.icache.r_data[1][2] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[1][30]$_DFFE_PP_  (.CLK(clknet_leaf_205_clk),
    .RESET_B(net2936),
    .D(_02055_),
    .Q_N(_13398_),
    .Q(\cpu.icache.r_data[1][30] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[1][31]$_DFFE_PP_  (.CLK(clknet_leaf_206_clk),
    .RESET_B(net2937),
    .D(_02056_),
    .Q_N(_13397_),
    .Q(\cpu.icache.r_data[1][31] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[1][3]$_DFFE_PP_  (.CLK(clknet_leaf_219_clk),
    .RESET_B(net2938),
    .D(_02057_),
    .Q_N(_13396_),
    .Q(\cpu.icache.r_data[1][3] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[1][4]$_DFFE_PP_  (.CLK(clknet_leaf_197_clk),
    .RESET_B(net2939),
    .D(_02058_),
    .Q_N(_13395_),
    .Q(\cpu.icache.r_data[1][4] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[1][5]$_DFFE_PP_  (.CLK(clknet_leaf_197_clk),
    .RESET_B(net2940),
    .D(_02059_),
    .Q_N(_13394_),
    .Q(\cpu.icache.r_data[1][5] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[1][6]$_DFFE_PP_  (.CLK(clknet_leaf_197_clk),
    .RESET_B(net2941),
    .D(_02060_),
    .Q_N(_13393_),
    .Q(\cpu.icache.r_data[1][6] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[1][7]$_DFFE_PP_  (.CLK(clknet_leaf_196_clk),
    .RESET_B(net2942),
    .D(_02061_),
    .Q_N(_13392_),
    .Q(\cpu.icache.r_data[1][7] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[1][8]$_DFFE_PP_  (.CLK(clknet_leaf_165_clk),
    .RESET_B(net2943),
    .D(_02062_),
    .Q_N(_13391_),
    .Q(\cpu.icache.r_data[1][8] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[1][9]$_DFFE_PP_  (.CLK(clknet_leaf_160_clk),
    .RESET_B(net2944),
    .D(_02063_),
    .Q_N(_13390_),
    .Q(\cpu.icache.r_data[1][9] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[2][0]$_DFFE_PP_  (.CLK(clknet_leaf_219_clk),
    .RESET_B(net2945),
    .D(_02064_),
    .Q_N(_13389_),
    .Q(\cpu.icache.r_data[2][0] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[2][10]$_DFFE_PP_  (.CLK(clknet_leaf_165_clk),
    .RESET_B(net2946),
    .D(_02065_),
    .Q_N(_13388_),
    .Q(\cpu.icache.r_data[2][10] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[2][11]$_DFFE_PP_  (.CLK(clknet_leaf_160_clk),
    .RESET_B(net2947),
    .D(_02066_),
    .Q_N(_13387_),
    .Q(\cpu.icache.r_data[2][11] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[2][12]$_DFFE_PP_  (.CLK(clknet_leaf_208_clk),
    .RESET_B(net2948),
    .D(_02067_),
    .Q_N(_13386_),
    .Q(\cpu.icache.r_data[2][12] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[2][13]$_DFFE_PP_  (.CLK(clknet_leaf_206_clk),
    .RESET_B(net2949),
    .D(_02068_),
    .Q_N(_13385_),
    .Q(\cpu.icache.r_data[2][13] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[2][14]$_DFFE_PP_  (.CLK(clknet_leaf_207_clk),
    .RESET_B(net2950),
    .D(_02069_),
    .Q_N(_13384_),
    .Q(\cpu.icache.r_data[2][14] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[2][15]$_DFFE_PP_  (.CLK(clknet_leaf_207_clk),
    .RESET_B(net2951),
    .D(_02070_),
    .Q_N(_13383_),
    .Q(\cpu.icache.r_data[2][15] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[2][16]$_DFFE_PP_  (.CLK(clknet_leaf_214_clk),
    .RESET_B(net2952),
    .D(_02071_),
    .Q_N(_13382_),
    .Q(\cpu.icache.r_data[2][16] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[2][17]$_DFFE_PP_  (.CLK(clknet_leaf_214_clk),
    .RESET_B(net2953),
    .D(_02072_),
    .Q_N(_13381_),
    .Q(\cpu.icache.r_data[2][17] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[2][18]$_DFFE_PP_  (.CLK(clknet_leaf_215_clk),
    .RESET_B(net2954),
    .D(_02073_),
    .Q_N(_13380_),
    .Q(\cpu.icache.r_data[2][18] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[2][19]$_DFFE_PP_  (.CLK(clknet_leaf_214_clk),
    .RESET_B(net2955),
    .D(_02074_),
    .Q_N(_13379_),
    .Q(\cpu.icache.r_data[2][19] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[2][1]$_DFFE_PP_  (.CLK(clknet_leaf_215_clk),
    .RESET_B(net2956),
    .D(_02075_),
    .Q_N(_13378_),
    .Q(\cpu.icache.r_data[2][1] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[2][20]$_DFFE_PP_  (.CLK(clknet_leaf_195_clk),
    .RESET_B(net2957),
    .D(_02076_),
    .Q_N(_13377_),
    .Q(\cpu.icache.r_data[2][20] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[2][21]$_DFFE_PP_  (.CLK(clknet_leaf_197_clk),
    .RESET_B(net2958),
    .D(_02077_),
    .Q_N(_13376_),
    .Q(\cpu.icache.r_data[2][21] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[2][22]$_DFFE_PP_  (.CLK(clknet_leaf_196_clk),
    .RESET_B(net2959),
    .D(_02078_),
    .Q_N(_13375_),
    .Q(\cpu.icache.r_data[2][22] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[2][23]$_DFFE_PP_  (.CLK(clknet_leaf_195_clk),
    .RESET_B(net2960),
    .D(_02079_),
    .Q_N(_13374_),
    .Q(\cpu.icache.r_data[2][23] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[2][24]$_DFFE_PP_  (.CLK(clknet_leaf_170_clk),
    .RESET_B(net2961),
    .D(_02080_),
    .Q_N(_13373_),
    .Q(\cpu.icache.r_data[2][24] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[2][25]$_DFFE_PP_  (.CLK(clknet_leaf_171_clk),
    .RESET_B(net2962),
    .D(_02081_),
    .Q_N(_13372_),
    .Q(\cpu.icache.r_data[2][25] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[2][26]$_DFFE_PP_  (.CLK(clknet_leaf_166_clk),
    .RESET_B(net2963),
    .D(_02082_),
    .Q_N(_13371_),
    .Q(\cpu.icache.r_data[2][26] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[2][27]$_DFFE_PP_  (.CLK(clknet_leaf_160_clk),
    .RESET_B(net2964),
    .D(_02083_),
    .Q_N(_13370_),
    .Q(\cpu.icache.r_data[2][27] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[2][28]$_DFFE_PP_  (.CLK(clknet_leaf_207_clk),
    .RESET_B(net2965),
    .D(_02084_),
    .Q_N(_13369_),
    .Q(\cpu.icache.r_data[2][28] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[2][29]$_DFFE_PP_  (.CLK(clknet_leaf_206_clk),
    .RESET_B(net2966),
    .D(_02085_),
    .Q_N(_13368_),
    .Q(\cpu.icache.r_data[2][29] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[2][2]$_DFFE_PP_  (.CLK(clknet_leaf_216_clk),
    .RESET_B(net2967),
    .D(_02086_),
    .Q_N(_13367_),
    .Q(\cpu.icache.r_data[2][2] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[2][30]$_DFFE_PP_  (.CLK(clknet_leaf_206_clk),
    .RESET_B(net2968),
    .D(_02087_),
    .Q_N(_13366_),
    .Q(\cpu.icache.r_data[2][30] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[2][31]$_DFFE_PP_  (.CLK(clknet_leaf_206_clk),
    .RESET_B(net2969),
    .D(_02088_),
    .Q_N(_13365_),
    .Q(\cpu.icache.r_data[2][31] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[2][3]$_DFFE_PP_  (.CLK(clknet_leaf_216_clk),
    .RESET_B(net2970),
    .D(_02089_),
    .Q_N(_13364_),
    .Q(\cpu.icache.r_data[2][3] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[2][4]$_DFFE_PP_  (.CLK(clknet_leaf_201_clk),
    .RESET_B(net2971),
    .D(_02090_),
    .Q_N(_13363_),
    .Q(\cpu.icache.r_data[2][4] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[2][5]$_DFFE_PP_  (.CLK(clknet_leaf_197_clk),
    .RESET_B(net2972),
    .D(_02091_),
    .Q_N(_13362_),
    .Q(\cpu.icache.r_data[2][5] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[2][6]$_DFFE_PP_  (.CLK(clknet_leaf_197_clk),
    .RESET_B(net2973),
    .D(_02092_),
    .Q_N(_13361_),
    .Q(\cpu.icache.r_data[2][6] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[2][7]$_DFFE_PP_  (.CLK(clknet_leaf_196_clk),
    .RESET_B(net2974),
    .D(_02093_),
    .Q_N(_13360_),
    .Q(\cpu.icache.r_data[2][7] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[2][8]$_DFFE_PP_  (.CLK(clknet_leaf_154_clk),
    .RESET_B(net2975),
    .D(_02094_),
    .Q_N(_13359_),
    .Q(\cpu.icache.r_data[2][8] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[2][9]$_DFFE_PP_  (.CLK(clknet_leaf_159_clk),
    .RESET_B(net2976),
    .D(_02095_),
    .Q_N(_13358_),
    .Q(\cpu.icache.r_data[2][9] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[3][0]$_DFFE_PP_  (.CLK(clknet_leaf_219_clk),
    .RESET_B(net2977),
    .D(_02096_),
    .Q_N(_13357_),
    .Q(\cpu.icache.r_data[3][0] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[3][10]$_DFFE_PP_  (.CLK(clknet_leaf_160_clk),
    .RESET_B(net2978),
    .D(_02097_),
    .Q_N(_13356_),
    .Q(\cpu.icache.r_data[3][10] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[3][11]$_DFFE_PP_  (.CLK(clknet_leaf_160_clk),
    .RESET_B(net2979),
    .D(_02098_),
    .Q_N(_13355_),
    .Q(\cpu.icache.r_data[3][11] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[3][12]$_DFFE_PP_  (.CLK(clknet_leaf_208_clk),
    .RESET_B(net2980),
    .D(_02099_),
    .Q_N(_13354_),
    .Q(\cpu.icache.r_data[3][12] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[3][13]$_DFFE_PP_  (.CLK(clknet_leaf_207_clk),
    .RESET_B(net2981),
    .D(_02100_),
    .Q_N(_13353_),
    .Q(\cpu.icache.r_data[3][13] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[3][14]$_DFFE_PP_  (.CLK(clknet_leaf_202_clk),
    .RESET_B(net2982),
    .D(_02101_),
    .Q_N(_13352_),
    .Q(\cpu.icache.r_data[3][14] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[3][15]$_DFFE_PP_  (.CLK(clknet_leaf_207_clk),
    .RESET_B(net2983),
    .D(_02102_),
    .Q_N(_13351_),
    .Q(\cpu.icache.r_data[3][15] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[3][16]$_DFFE_PP_  (.CLK(clknet_leaf_213_clk),
    .RESET_B(net2984),
    .D(_02103_),
    .Q_N(_13350_),
    .Q(\cpu.icache.r_data[3][16] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[3][17]$_DFFE_PP_  (.CLK(clknet_leaf_222_clk),
    .RESET_B(net2985),
    .D(_02104_),
    .Q_N(_13349_),
    .Q(\cpu.icache.r_data[3][17] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[3][18]$_DFFE_PP_  (.CLK(clknet_leaf_212_clk),
    .RESET_B(net2986),
    .D(_02105_),
    .Q_N(_13348_),
    .Q(\cpu.icache.r_data[3][18] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[3][19]$_DFFE_PP_  (.CLK(clknet_leaf_222_clk),
    .RESET_B(net2987),
    .D(_02106_),
    .Q_N(_13347_),
    .Q(\cpu.icache.r_data[3][19] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[3][1]$_DFFE_PP_  (.CLK(clknet_leaf_215_clk),
    .RESET_B(net2988),
    .D(_02107_),
    .Q_N(_13346_),
    .Q(\cpu.icache.r_data[3][1] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[3][20]$_DFFE_PP_  (.CLK(clknet_leaf_201_clk),
    .RESET_B(net2989),
    .D(_02108_),
    .Q_N(_13345_),
    .Q(\cpu.icache.r_data[3][20] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[3][21]$_DFFE_PP_  (.CLK(clknet_leaf_197_clk),
    .RESET_B(net2990),
    .D(_02109_),
    .Q_N(_13344_),
    .Q(\cpu.icache.r_data[3][21] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[3][22]$_DFFE_PP_  (.CLK(clknet_leaf_196_clk),
    .RESET_B(net2991),
    .D(_02110_),
    .Q_N(_13343_),
    .Q(\cpu.icache.r_data[3][22] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[3][23]$_DFFE_PP_  (.CLK(clknet_leaf_201_clk),
    .RESET_B(net2992),
    .D(_02111_),
    .Q_N(_13342_),
    .Q(\cpu.icache.r_data[3][23] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[3][24]$_DFFE_PP_  (.CLK(clknet_leaf_164_clk),
    .RESET_B(net2993),
    .D(_02112_),
    .Q_N(_13341_),
    .Q(\cpu.icache.r_data[3][24] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[3][25]$_DFFE_PP_  (.CLK(clknet_leaf_164_clk),
    .RESET_B(net2994),
    .D(_02113_),
    .Q_N(_13340_),
    .Q(\cpu.icache.r_data[3][25] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[3][26]$_DFFE_PP_  (.CLK(clknet_leaf_164_clk),
    .RESET_B(net2995),
    .D(_02114_),
    .Q_N(_13339_),
    .Q(\cpu.icache.r_data[3][26] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[3][27]$_DFFE_PP_  (.CLK(clknet_leaf_165_clk),
    .RESET_B(net2996),
    .D(_02115_),
    .Q_N(_13338_),
    .Q(\cpu.icache.r_data[3][27] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[3][28]$_DFFE_PP_  (.CLK(clknet_leaf_202_clk),
    .RESET_B(net2997),
    .D(_02116_),
    .Q_N(_13337_),
    .Q(\cpu.icache.r_data[3][28] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[3][29]$_DFFE_PP_  (.CLK(clknet_leaf_202_clk),
    .RESET_B(net2998),
    .D(_02117_),
    .Q_N(_13336_),
    .Q(\cpu.icache.r_data[3][29] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[3][2]$_DFFE_PP_  (.CLK(clknet_leaf_216_clk),
    .RESET_B(net2999),
    .D(_02118_),
    .Q_N(_13335_),
    .Q(\cpu.icache.r_data[3][2] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[3][30]$_DFFE_PP_  (.CLK(clknet_leaf_203_clk),
    .RESET_B(net3000),
    .D(_02119_),
    .Q_N(_13334_),
    .Q(\cpu.icache.r_data[3][30] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[3][31]$_DFFE_PP_  (.CLK(clknet_leaf_203_clk),
    .RESET_B(net3001),
    .D(_02120_),
    .Q_N(_13333_),
    .Q(\cpu.icache.r_data[3][31] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[3][3]$_DFFE_PP_  (.CLK(clknet_leaf_216_clk),
    .RESET_B(net3002),
    .D(_02121_),
    .Q_N(_13332_),
    .Q(\cpu.icache.r_data[3][3] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[3][4]$_DFFE_PP_  (.CLK(clknet_leaf_201_clk),
    .RESET_B(net3003),
    .D(_02122_),
    .Q_N(_13331_),
    .Q(\cpu.icache.r_data[3][4] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[3][5]$_DFFE_PP_  (.CLK(clknet_leaf_198_clk),
    .RESET_B(net3004),
    .D(_02123_),
    .Q_N(_13330_),
    .Q(\cpu.icache.r_data[3][5] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[3][6]$_DFFE_PP_  (.CLK(clknet_leaf_198_clk),
    .RESET_B(net3005),
    .D(_02124_),
    .Q_N(_13329_),
    .Q(\cpu.icache.r_data[3][6] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[3][7]$_DFFE_PP_  (.CLK(clknet_leaf_201_clk),
    .RESET_B(net3006),
    .D(_02125_),
    .Q_N(_13328_),
    .Q(\cpu.icache.r_data[3][7] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[3][8]$_DFFE_PP_  (.CLK(clknet_leaf_154_clk),
    .RESET_B(net3007),
    .D(_02126_),
    .Q_N(_13327_),
    .Q(\cpu.icache.r_data[3][8] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[3][9]$_DFFE_PP_  (.CLK(clknet_leaf_159_clk),
    .RESET_B(net3008),
    .D(_02127_),
    .Q_N(_13326_),
    .Q(\cpu.icache.r_data[3][9] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[4][0]$_DFFE_PP_  (.CLK(clknet_leaf_221_clk),
    .RESET_B(net3009),
    .D(_02128_),
    .Q_N(_13325_),
    .Q(\cpu.icache.r_data[4][0] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[4][10]$_DFFE_PP_  (.CLK(clknet_leaf_163_clk),
    .RESET_B(net3010),
    .D(_02129_),
    .Q_N(_13324_),
    .Q(\cpu.icache.r_data[4][10] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[4][11]$_DFFE_PP_  (.CLK(clknet_leaf_161_clk),
    .RESET_B(net3011),
    .D(_02130_),
    .Q_N(_13323_),
    .Q(\cpu.icache.r_data[4][11] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[4][12]$_DFFE_PP_  (.CLK(clknet_leaf_200_clk),
    .RESET_B(net3012),
    .D(_02131_),
    .Q_N(_13322_),
    .Q(\cpu.icache.r_data[4][12] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[4][13]$_DFFE_PP_  (.CLK(clknet_leaf_203_clk),
    .RESET_B(net3013),
    .D(_02132_),
    .Q_N(_13321_),
    .Q(\cpu.icache.r_data[4][13] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[4][14]$_DFFE_PP_  (.CLK(clknet_leaf_204_clk),
    .RESET_B(net3014),
    .D(_02133_),
    .Q_N(_13320_),
    .Q(\cpu.icache.r_data[4][14] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[4][15]$_DFFE_PP_  (.CLK(clknet_leaf_203_clk),
    .RESET_B(net3015),
    .D(_02134_),
    .Q_N(_13319_),
    .Q(\cpu.icache.r_data[4][15] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[4][16]$_DFFE_PP_  (.CLK(clknet_leaf_221_clk),
    .RESET_B(net3016),
    .D(_02135_),
    .Q_N(_13318_),
    .Q(\cpu.icache.r_data[4][16] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[4][17]$_DFFE_PP_  (.CLK(clknet_leaf_220_clk),
    .RESET_B(net3017),
    .D(_02136_),
    .Q_N(_13317_),
    .Q(\cpu.icache.r_data[4][17] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[4][18]$_DFFE_PP_  (.CLK(clknet_leaf_220_clk),
    .RESET_B(net3018),
    .D(_02137_),
    .Q_N(_13316_),
    .Q(\cpu.icache.r_data[4][18] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[4][19]$_DFFE_PP_  (.CLK(clknet_leaf_219_clk),
    .RESET_B(net3019),
    .D(_02138_),
    .Q_N(_13315_),
    .Q(\cpu.icache.r_data[4][19] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[4][1]$_DFFE_PP_  (.CLK(clknet_leaf_220_clk),
    .RESET_B(net3020),
    .D(_02139_),
    .Q_N(_13314_),
    .Q(\cpu.icache.r_data[4][1] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[4][20]$_DFFE_PP_  (.CLK(clknet_leaf_218_clk),
    .RESET_B(net3021),
    .D(_02140_),
    .Q_N(_13313_),
    .Q(\cpu.icache.r_data[4][20] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[4][21]$_DFFE_PP_  (.CLK(clknet_leaf_217_clk),
    .RESET_B(net3022),
    .D(_02141_),
    .Q_N(_13312_),
    .Q(\cpu.icache.r_data[4][21] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[4][22]$_DFFE_PP_  (.CLK(clknet_leaf_217_clk),
    .RESET_B(net3023),
    .D(_02142_),
    .Q_N(_13311_),
    .Q(\cpu.icache.r_data[4][22] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[4][23]$_DFFE_PP_  (.CLK(clknet_leaf_218_clk),
    .RESET_B(net3024),
    .D(_02143_),
    .Q_N(_13310_),
    .Q(\cpu.icache.r_data[4][23] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[4][24]$_DFFE_PP_  (.CLK(clknet_leaf_161_clk),
    .RESET_B(net3025),
    .D(_02144_),
    .Q_N(_13309_),
    .Q(\cpu.icache.r_data[4][24] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[4][25]$_DFFE_PP_  (.CLK(clknet_leaf_162_clk),
    .RESET_B(net3026),
    .D(_02145_),
    .Q_N(_13308_),
    .Q(\cpu.icache.r_data[4][25] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[4][26]$_DFFE_PP_  (.CLK(clknet_leaf_158_clk),
    .RESET_B(net3027),
    .D(_02146_),
    .Q_N(_13307_),
    .Q(\cpu.icache.r_data[4][26] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[4][27]$_DFFE_PP_  (.CLK(clknet_leaf_159_clk),
    .RESET_B(net3028),
    .D(_02147_),
    .Q_N(_13306_),
    .Q(\cpu.icache.r_data[4][27] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[4][28]$_DFFE_PP_  (.CLK(clknet_leaf_204_clk),
    .RESET_B(net3029),
    .D(_02148_),
    .Q_N(_13305_),
    .Q(\cpu.icache.r_data[4][28] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[4][29]$_DFFE_PP_  (.CLK(clknet_leaf_204_clk),
    .RESET_B(net3030),
    .D(_02149_),
    .Q_N(_13304_),
    .Q(\cpu.icache.r_data[4][29] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[4][2]$_DFFE_PP_  (.CLK(clknet_leaf_218_clk),
    .RESET_B(net3031),
    .D(_02150_),
    .Q_N(_13303_),
    .Q(\cpu.icache.r_data[4][2] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[4][30]$_DFFE_PP_  (.CLK(clknet_leaf_205_clk),
    .RESET_B(net3032),
    .D(_02151_),
    .Q_N(_13302_),
    .Q(\cpu.icache.r_data[4][30] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[4][31]$_DFFE_PP_  (.CLK(clknet_leaf_217_clk),
    .RESET_B(net3033),
    .D(_02152_),
    .Q_N(_13301_),
    .Q(\cpu.icache.r_data[4][31] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[4][3]$_DFFE_PP_  (.CLK(clknet_leaf_220_clk),
    .RESET_B(net3034),
    .D(_02153_),
    .Q_N(_13300_),
    .Q(\cpu.icache.r_data[4][3] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[4][4]$_DFFE_PP_  (.CLK(clknet_leaf_199_clk),
    .RESET_B(net3035),
    .D(_02154_),
    .Q_N(_13299_),
    .Q(\cpu.icache.r_data[4][4] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[4][5]$_DFFE_PP_  (.CLK(clknet_leaf_198_clk),
    .RESET_B(net3036),
    .D(_02155_),
    .Q_N(_13298_),
    .Q(\cpu.icache.r_data[4][5] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[4][6]$_DFFE_PP_  (.CLK(clknet_leaf_198_clk),
    .RESET_B(net3037),
    .D(_02156_),
    .Q_N(_13297_),
    .Q(\cpu.icache.r_data[4][6] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[4][7]$_DFFE_PP_  (.CLK(clknet_leaf_199_clk),
    .RESET_B(net3038),
    .D(_02157_),
    .Q_N(_13296_),
    .Q(\cpu.icache.r_data[4][7] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[4][8]$_DFFE_PP_  (.CLK(clknet_leaf_163_clk),
    .RESET_B(net3039),
    .D(_02158_),
    .Q_N(_13295_),
    .Q(\cpu.icache.r_data[4][8] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[4][9]$_DFFE_PP_  (.CLK(clknet_leaf_162_clk),
    .RESET_B(net3040),
    .D(_02159_),
    .Q_N(_13294_),
    .Q(\cpu.icache.r_data[4][9] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[5][0]$_DFFE_PP_  (.CLK(clknet_leaf_219_clk),
    .RESET_B(net3041),
    .D(_02160_),
    .Q_N(_13293_),
    .Q(\cpu.icache.r_data[5][0] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[5][10]$_DFFE_PP_  (.CLK(clknet_leaf_163_clk),
    .RESET_B(net3042),
    .D(_02161_),
    .Q_N(_13292_),
    .Q(\cpu.icache.r_data[5][10] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[5][11]$_DFFE_PP_  (.CLK(clknet_leaf_161_clk),
    .RESET_B(net3043),
    .D(_02162_),
    .Q_N(_13291_),
    .Q(\cpu.icache.r_data[5][11] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[5][12]$_DFFE_PP_  (.CLK(clknet_leaf_202_clk),
    .RESET_B(net3044),
    .D(_02163_),
    .Q_N(_13290_),
    .Q(\cpu.icache.r_data[5][12] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[5][13]$_DFFE_PP_  (.CLK(clknet_leaf_200_clk),
    .RESET_B(net3045),
    .D(_02164_),
    .Q_N(_13289_),
    .Q(\cpu.icache.r_data[5][13] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[5][14]$_DFFE_PP_  (.CLK(clknet_leaf_204_clk),
    .RESET_B(net3046),
    .D(_02165_),
    .Q_N(_13288_),
    .Q(\cpu.icache.r_data[5][14] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[5][15]$_DFFE_PP_  (.CLK(clknet_leaf_203_clk),
    .RESET_B(net3047),
    .D(_02166_),
    .Q_N(_13287_),
    .Q(\cpu.icache.r_data[5][15] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[5][16]$_DFFE_PP_  (.CLK(clknet_leaf_215_clk),
    .RESET_B(net3048),
    .D(_02167_),
    .Q_N(_13286_),
    .Q(\cpu.icache.r_data[5][16] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[5][17]$_DFFE_PP_  (.CLK(clknet_leaf_215_clk),
    .RESET_B(net3049),
    .D(_02168_),
    .Q_N(_13285_),
    .Q(\cpu.icache.r_data[5][17] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[5][18]$_DFFE_PP_  (.CLK(clknet_leaf_215_clk),
    .RESET_B(net3050),
    .D(_02169_),
    .Q_N(_13284_),
    .Q(\cpu.icache.r_data[5][18] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[5][19]$_DFFE_PP_  (.CLK(clknet_leaf_214_clk),
    .RESET_B(net3051),
    .D(_02170_),
    .Q_N(_13283_),
    .Q(\cpu.icache.r_data[5][19] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[5][1]$_DFFE_PP_  (.CLK(clknet_leaf_220_clk),
    .RESET_B(net3052),
    .D(_02171_),
    .Q_N(_13282_),
    .Q(\cpu.icache.r_data[5][1] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[5][20]$_DFFE_PP_  (.CLK(clknet_leaf_216_clk),
    .RESET_B(net3053),
    .D(_02172_),
    .Q_N(_13281_),
    .Q(\cpu.icache.r_data[5][20] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[5][21]$_DFFE_PP_  (.CLK(clknet_leaf_199_clk),
    .RESET_B(net3054),
    .D(_02173_),
    .Q_N(_13280_),
    .Q(\cpu.icache.r_data[5][21] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[5][22]$_DFFE_PP_  (.CLK(clknet_leaf_205_clk),
    .RESET_B(net3055),
    .D(_02174_),
    .Q_N(_13279_),
    .Q(\cpu.icache.r_data[5][22] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[5][23]$_DFFE_PP_  (.CLK(clknet_leaf_216_clk),
    .RESET_B(net3056),
    .D(_02175_),
    .Q_N(_13278_),
    .Q(\cpu.icache.r_data[5][23] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[5][24]$_DFFE_PP_  (.CLK(clknet_leaf_162_clk),
    .RESET_B(net3057),
    .D(_02176_),
    .Q_N(_13277_),
    .Q(\cpu.icache.r_data[5][24] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[5][25]$_DFFE_PP_  (.CLK(clknet_leaf_161_clk),
    .RESET_B(net3058),
    .D(_02177_),
    .Q_N(_13276_),
    .Q(\cpu.icache.r_data[5][25] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[5][26]$_DFFE_PP_  (.CLK(clknet_leaf_164_clk),
    .RESET_B(net3059),
    .D(_02178_),
    .Q_N(_13275_),
    .Q(\cpu.icache.r_data[5][26] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[5][27]$_DFFE_PP_  (.CLK(clknet_leaf_164_clk),
    .RESET_B(net3060),
    .D(_02179_),
    .Q_N(_13274_),
    .Q(\cpu.icache.r_data[5][27] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[5][28]$_DFFE_PP_  (.CLK(clknet_leaf_205_clk),
    .RESET_B(net3061),
    .D(_02180_),
    .Q_N(_13273_),
    .Q(\cpu.icache.r_data[5][28] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[5][29]$_DFFE_PP_  (.CLK(clknet_leaf_206_clk),
    .RESET_B(net3062),
    .D(_02181_),
    .Q_N(_13272_),
    .Q(\cpu.icache.r_data[5][29] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[5][2]$_DFFE_PP_  (.CLK(clknet_leaf_216_clk),
    .RESET_B(net3063),
    .D(_02182_),
    .Q_N(_13271_),
    .Q(\cpu.icache.r_data[5][2] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[5][30]$_DFFE_PP_  (.CLK(clknet_leaf_205_clk),
    .RESET_B(net3064),
    .D(_02183_),
    .Q_N(_13270_),
    .Q(\cpu.icache.r_data[5][30] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[5][31]$_DFFE_PP_  (.CLK(clknet_leaf_205_clk),
    .RESET_B(net3065),
    .D(_02184_),
    .Q_N(_13269_),
    .Q(\cpu.icache.r_data[5][31] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[5][3]$_DFFE_PP_  (.CLK(clknet_leaf_221_clk),
    .RESET_B(net3066),
    .D(_02185_),
    .Q_N(_13268_),
    .Q(\cpu.icache.r_data[5][3] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[5][4]$_DFFE_PP_  (.CLK(clknet_leaf_199_clk),
    .RESET_B(net3067),
    .D(_02186_),
    .Q_N(_13267_),
    .Q(\cpu.icache.r_data[5][4] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[5][5]$_DFFE_PP_  (.CLK(clknet_leaf_198_clk),
    .RESET_B(net3068),
    .D(_02187_),
    .Q_N(_13266_),
    .Q(\cpu.icache.r_data[5][5] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[5][6]$_DFFE_PP_  (.CLK(clknet_leaf_198_clk),
    .RESET_B(net3069),
    .D(_02188_),
    .Q_N(_13265_),
    .Q(\cpu.icache.r_data[5][6] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[5][7]$_DFFE_PP_  (.CLK(clknet_leaf_201_clk),
    .RESET_B(net3070),
    .D(_02189_),
    .Q_N(_13264_),
    .Q(\cpu.icache.r_data[5][7] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[5][8]$_DFFE_PP_  (.CLK(clknet_leaf_163_clk),
    .RESET_B(net3071),
    .D(_02190_),
    .Q_N(_13263_),
    .Q(\cpu.icache.r_data[5][8] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[5][9]$_DFFE_PP_  (.CLK(clknet_leaf_162_clk),
    .RESET_B(net3072),
    .D(_02191_),
    .Q_N(_13262_),
    .Q(\cpu.icache.r_data[5][9] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[6][0]$_DFFE_PP_  (.CLK(clknet_leaf_218_clk),
    .RESET_B(net3073),
    .D(_02192_),
    .Q_N(_13261_),
    .Q(\cpu.icache.r_data[6][0] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[6][10]$_DFFE_PP_  (.CLK(clknet_leaf_163_clk),
    .RESET_B(net3074),
    .D(_02193_),
    .Q_N(_13260_),
    .Q(\cpu.icache.r_data[6][10] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[6][11]$_DFFE_PP_  (.CLK(clknet_leaf_162_clk),
    .RESET_B(net3075),
    .D(_02194_),
    .Q_N(_13259_),
    .Q(\cpu.icache.r_data[6][11] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[6][12]$_DFFE_PP_  (.CLK(clknet_leaf_200_clk),
    .RESET_B(net3076),
    .D(_02195_),
    .Q_N(_13258_),
    .Q(\cpu.icache.r_data[6][12] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[6][13]$_DFFE_PP_  (.CLK(clknet_leaf_203_clk),
    .RESET_B(net3077),
    .D(_02196_),
    .Q_N(_13257_),
    .Q(\cpu.icache.r_data[6][13] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[6][14]$_DFFE_PP_  (.CLK(clknet_leaf_204_clk),
    .RESET_B(net3078),
    .D(_02197_),
    .Q_N(_13256_),
    .Q(\cpu.icache.r_data[6][14] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[6][15]$_DFFE_PP_  (.CLK(clknet_leaf_204_clk),
    .RESET_B(net3079),
    .D(_02198_),
    .Q_N(_13255_),
    .Q(\cpu.icache.r_data[6][15] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[6][16]$_DFFE_PP_  (.CLK(clknet_leaf_221_clk),
    .RESET_B(net3080),
    .D(_02199_),
    .Q_N(_13254_),
    .Q(\cpu.icache.r_data[6][16] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[6][17]$_DFFE_PP_  (.CLK(clknet_leaf_221_clk),
    .RESET_B(net3081),
    .D(_02200_),
    .Q_N(_13253_),
    .Q(\cpu.icache.r_data[6][17] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[6][18]$_DFFE_PP_  (.CLK(clknet_leaf_221_clk),
    .RESET_B(net3082),
    .D(_02201_),
    .Q_N(_13252_),
    .Q(\cpu.icache.r_data[6][18] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[6][19]$_DFFE_PP_  (.CLK(clknet_leaf_221_clk),
    .RESET_B(net3083),
    .D(_02202_),
    .Q_N(_13251_),
    .Q(\cpu.icache.r_data[6][19] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[6][1]$_DFFE_PP_  (.CLK(clknet_leaf_220_clk),
    .RESET_B(net3084),
    .D(_02203_),
    .Q_N(_13250_),
    .Q(\cpu.icache.r_data[6][1] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[6][20]$_DFFE_PP_  (.CLK(clknet_leaf_217_clk),
    .RESET_B(net3085),
    .D(_02204_),
    .Q_N(_13249_),
    .Q(\cpu.icache.r_data[6][20] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[6][21]$_DFFE_PP_  (.CLK(clknet_leaf_217_clk),
    .RESET_B(net3086),
    .D(_02205_),
    .Q_N(_13248_),
    .Q(\cpu.icache.r_data[6][21] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[6][22]$_DFFE_PP_  (.CLK(clknet_leaf_217_clk),
    .RESET_B(net3087),
    .D(_02206_),
    .Q_N(_13247_),
    .Q(\cpu.icache.r_data[6][22] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[6][23]$_DFFE_PP_  (.CLK(clknet_leaf_217_clk),
    .RESET_B(net3088),
    .D(_02207_),
    .Q_N(_13246_),
    .Q(\cpu.icache.r_data[6][23] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[6][24]$_DFFE_PP_  (.CLK(clknet_leaf_161_clk),
    .RESET_B(net3089),
    .D(_02208_),
    .Q_N(_13245_),
    .Q(\cpu.icache.r_data[6][24] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[6][25]$_DFFE_PP_  (.CLK(clknet_leaf_158_clk),
    .RESET_B(net3090),
    .D(_02209_),
    .Q_N(_13244_),
    .Q(\cpu.icache.r_data[6][25] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[6][26]$_DFFE_PP_  (.CLK(clknet_leaf_158_clk),
    .RESET_B(net3091),
    .D(_02210_),
    .Q_N(_13243_),
    .Q(\cpu.icache.r_data[6][26] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[6][27]$_DFFE_PP_  (.CLK(clknet_leaf_161_clk),
    .RESET_B(net3092),
    .D(_02211_),
    .Q_N(_13242_),
    .Q(\cpu.icache.r_data[6][27] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[6][28]$_DFFE_PP_  (.CLK(clknet_leaf_204_clk),
    .RESET_B(net3093),
    .D(_02212_),
    .Q_N(_13241_),
    .Q(\cpu.icache.r_data[6][28] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[6][29]$_DFFE_PP_  (.CLK(clknet_leaf_205_clk),
    .RESET_B(net3094),
    .D(_02213_),
    .Q_N(_13240_),
    .Q(\cpu.icache.r_data[6][29] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[6][2]$_DFFE_PP_  (.CLK(clknet_leaf_219_clk),
    .RESET_B(net3095),
    .D(_02214_),
    .Q_N(_13239_),
    .Q(\cpu.icache.r_data[6][2] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[6][30]$_DFFE_PP_  (.CLK(clknet_leaf_204_clk),
    .RESET_B(net3096),
    .D(_02215_),
    .Q_N(_13238_),
    .Q(\cpu.icache.r_data[6][30] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[6][31]$_DFFE_PP_  (.CLK(clknet_leaf_217_clk),
    .RESET_B(net3097),
    .D(_02216_),
    .Q_N(_13237_),
    .Q(\cpu.icache.r_data[6][31] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[6][3]$_DFFE_PP_  (.CLK(clknet_leaf_221_clk),
    .RESET_B(net3098),
    .D(_02217_),
    .Q_N(_13236_),
    .Q(\cpu.icache.r_data[6][3] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[6][4]$_DFFE_PP_  (.CLK(clknet_leaf_200_clk),
    .RESET_B(net3099),
    .D(_02218_),
    .Q_N(_13235_),
    .Q(\cpu.icache.r_data[6][4] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[6][5]$_DFFE_PP_  (.CLK(clknet_leaf_199_clk),
    .RESET_B(net3100),
    .D(_02219_),
    .Q_N(_13234_),
    .Q(\cpu.icache.r_data[6][5] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[6][6]$_DFFE_PP_  (.CLK(clknet_leaf_199_clk),
    .RESET_B(net3101),
    .D(_02220_),
    .Q_N(_13233_),
    .Q(\cpu.icache.r_data[6][6] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[6][7]$_DFFE_PP_  (.CLK(clknet_leaf_200_clk),
    .RESET_B(net3102),
    .D(_02221_),
    .Q_N(_13232_),
    .Q(\cpu.icache.r_data[6][7] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[6][8]$_DFFE_PP_  (.CLK(clknet_leaf_163_clk),
    .RESET_B(net3103),
    .D(_02222_),
    .Q_N(_13231_),
    .Q(\cpu.icache.r_data[6][8] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[6][9]$_DFFE_PP_  (.CLK(clknet_leaf_162_clk),
    .RESET_B(net3104),
    .D(_02223_),
    .Q_N(_13230_),
    .Q(\cpu.icache.r_data[6][9] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[7][0]$_DFFE_PP_  (.CLK(clknet_leaf_218_clk),
    .RESET_B(net3105),
    .D(_02224_),
    .Q_N(_13229_),
    .Q(\cpu.icache.r_data[7][0] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[7][10]$_DFFE_PP_  (.CLK(clknet_leaf_163_clk),
    .RESET_B(net3106),
    .D(_02225_),
    .Q_N(_13228_),
    .Q(\cpu.icache.r_data[7][10] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[7][11]$_DFFE_PP_  (.CLK(clknet_leaf_162_clk),
    .RESET_B(net3107),
    .D(_02226_),
    .Q_N(_13227_),
    .Q(\cpu.icache.r_data[7][11] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[7][12]$_DFFE_PP_  (.CLK(clknet_leaf_203_clk),
    .RESET_B(net3108),
    .D(_02227_),
    .Q_N(_13226_),
    .Q(\cpu.icache.r_data[7][12] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[7][13]$_DFFE_PP_  (.CLK(clknet_leaf_200_clk),
    .RESET_B(net3109),
    .D(_02228_),
    .Q_N(_13225_),
    .Q(\cpu.icache.r_data[7][13] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[7][14]$_DFFE_PP_  (.CLK(clknet_leaf_203_clk),
    .RESET_B(net3110),
    .D(_02229_),
    .Q_N(_13224_),
    .Q(\cpu.icache.r_data[7][14] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[7][15]$_DFFE_PP_  (.CLK(clknet_leaf_200_clk),
    .RESET_B(net3111),
    .D(_02230_),
    .Q_N(_13223_),
    .Q(\cpu.icache.r_data[7][15] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[7][16]$_DFFE_PP_  (.CLK(clknet_leaf_214_clk),
    .RESET_B(net3112),
    .D(_02231_),
    .Q_N(_13222_),
    .Q(\cpu.icache.r_data[7][16] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[7][17]$_DFFE_PP_  (.CLK(clknet_leaf_222_clk),
    .RESET_B(net3113),
    .D(_02232_),
    .Q_N(_13221_),
    .Q(\cpu.icache.r_data[7][17] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[7][18]$_DFFE_PP_  (.CLK(clknet_leaf_212_clk),
    .RESET_B(net3114),
    .D(_02233_),
    .Q_N(_13220_),
    .Q(\cpu.icache.r_data[7][18] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[7][19]$_DFFE_PP_  (.CLK(clknet_leaf_222_clk),
    .RESET_B(net3115),
    .D(_02234_),
    .Q_N(_13219_),
    .Q(\cpu.icache.r_data[7][19] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[7][1]$_DFFE_PP_  (.CLK(clknet_leaf_220_clk),
    .RESET_B(net3116),
    .D(_02235_),
    .Q_N(_13218_),
    .Q(\cpu.icache.r_data[7][1] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[7][20]$_DFFE_PP_  (.CLK(clknet_leaf_201_clk),
    .RESET_B(net3117),
    .D(_02236_),
    .Q_N(_13217_),
    .Q(\cpu.icache.r_data[7][20] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[7][21]$_DFFE_PP_  (.CLK(clknet_leaf_201_clk),
    .RESET_B(net3118),
    .D(_02237_),
    .Q_N(_13216_),
    .Q(\cpu.icache.r_data[7][21] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[7][22]$_DFFE_PP_  (.CLK(clknet_leaf_205_clk),
    .RESET_B(net3119),
    .D(_02238_),
    .Q_N(_13215_),
    .Q(\cpu.icache.r_data[7][22] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[7][23]$_DFFE_PP_  (.CLK(clknet_leaf_218_clk),
    .RESET_B(net3120),
    .D(_02239_),
    .Q_N(_13214_),
    .Q(\cpu.icache.r_data[7][23] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[7][24]$_DFFE_PP_  (.CLK(clknet_leaf_164_clk),
    .RESET_B(net3121),
    .D(_02240_),
    .Q_N(_13213_),
    .Q(\cpu.icache.r_data[7][24] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[7][25]$_DFFE_PP_  (.CLK(clknet_leaf_161_clk),
    .RESET_B(net3122),
    .D(_02241_),
    .Q_N(_13212_),
    .Q(\cpu.icache.r_data[7][25] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[7][26]$_DFFE_PP_  (.CLK(clknet_leaf_164_clk),
    .RESET_B(net3123),
    .D(_02242_),
    .Q_N(_13211_),
    .Q(\cpu.icache.r_data[7][26] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[7][27]$_DFFE_PP_  (.CLK(clknet_leaf_164_clk),
    .RESET_B(net3124),
    .D(_02243_),
    .Q_N(_13210_),
    .Q(\cpu.icache.r_data[7][27] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[7][28]$_DFFE_PP_  (.CLK(clknet_leaf_202_clk),
    .RESET_B(net3125),
    .D(_02244_),
    .Q_N(_13209_),
    .Q(\cpu.icache.r_data[7][28] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[7][29]$_DFFE_PP_  (.CLK(clknet_leaf_202_clk),
    .RESET_B(net3126),
    .D(_02245_),
    .Q_N(_13208_),
    .Q(\cpu.icache.r_data[7][29] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[7][2]$_DFFE_PP_  (.CLK(clknet_leaf_218_clk),
    .RESET_B(net3127),
    .D(_02246_),
    .Q_N(_13207_),
    .Q(\cpu.icache.r_data[7][2] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[7][30]$_DFFE_PP_  (.CLK(clknet_leaf_200_clk),
    .RESET_B(net3128),
    .D(_02247_),
    .Q_N(_13206_),
    .Q(\cpu.icache.r_data[7][30] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[7][31]$_DFFE_PP_  (.CLK(clknet_leaf_202_clk),
    .RESET_B(net3129),
    .D(_02248_),
    .Q_N(_13205_),
    .Q(\cpu.icache.r_data[7][31] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[7][3]$_DFFE_PP_  (.CLK(clknet_leaf_218_clk),
    .RESET_B(net3130),
    .D(_02249_),
    .Q_N(_13204_),
    .Q(\cpu.icache.r_data[7][3] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[7][4]$_DFFE_PP_  (.CLK(clknet_leaf_199_clk),
    .RESET_B(net3131),
    .D(_02250_),
    .Q_N(_13203_),
    .Q(\cpu.icache.r_data[7][4] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[7][5]$_DFFE_PP_  (.CLK(clknet_leaf_198_clk),
    .RESET_B(net3132),
    .D(_02251_),
    .Q_N(_13202_),
    .Q(\cpu.icache.r_data[7][5] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[7][6]$_DFFE_PP_  (.CLK(clknet_leaf_198_clk),
    .RESET_B(net3133),
    .D(_02252_),
    .Q_N(_13201_),
    .Q(\cpu.icache.r_data[7][6] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[7][7]$_DFFE_PP_  (.CLK(clknet_leaf_199_clk),
    .RESET_B(net3134),
    .D(_02253_),
    .Q_N(_13200_),
    .Q(\cpu.icache.r_data[7][7] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[7][8]$_DFFE_PP_  (.CLK(clknet_leaf_163_clk),
    .RESET_B(net3135),
    .D(_02254_),
    .Q_N(_13199_),
    .Q(\cpu.icache.r_data[7][8] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[7][9]$_DFFE_PP_  (.CLK(clknet_leaf_162_clk),
    .RESET_B(net3136),
    .D(_02255_),
    .Q_N(_13198_),
    .Q(\cpu.icache.r_data[7][9] ));
 sg13g2_dfrbp_1 \cpu.icache.r_offset[0]$_SDFF_PN0_  (.CLK(clknet_leaf_165_clk),
    .RESET_B(net3137),
    .D(_02256_),
    .Q_N(_00304_),
    .Q(\cpu.icache.r_offset[0] ));
 sg13g2_dfrbp_1 \cpu.icache.r_offset[1]$_SDFF_PN0_  (.CLK(clknet_leaf_197_clk),
    .RESET_B(net3138),
    .D(_02257_),
    .Q_N(_13197_),
    .Q(\cpu.icache.r_offset[1] ));
 sg13g2_dfrbp_1 \cpu.icache.r_offset[2]$_SDFF_PN0_  (.CLK(clknet_leaf_165_clk),
    .RESET_B(net3139),
    .D(_02258_),
    .Q_N(_00238_),
    .Q(\cpu.icache.r_offset[2] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[0][0]$_DFFE_PP_  (.CLK(clknet_leaf_152_clk),
    .RESET_B(net3140),
    .D(_02259_),
    .Q_N(_13196_),
    .Q(\cpu.icache.r_tag[0][5] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[0][10]$_DFFE_PP_  (.CLK(clknet_leaf_131_clk),
    .RESET_B(net3141),
    .D(_02260_),
    .Q_N(_13195_),
    .Q(\cpu.icache.r_tag[0][15] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[0][11]$_DFFE_PP_  (.CLK(clknet_leaf_131_clk),
    .RESET_B(net3142),
    .D(_02261_),
    .Q_N(_13194_),
    .Q(\cpu.icache.r_tag[0][16] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[0][12]$_DFFE_PP_  (.CLK(clknet_leaf_136_clk),
    .RESET_B(net3143),
    .D(_02262_),
    .Q_N(_13193_),
    .Q(\cpu.icache.r_tag[0][17] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[0][13]$_DFFE_PP_  (.CLK(clknet_leaf_137_clk),
    .RESET_B(net3144),
    .D(_02263_),
    .Q_N(_13192_),
    .Q(\cpu.icache.r_tag[0][18] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[0][14]$_DFFE_PP_  (.CLK(clknet_leaf_136_clk),
    .RESET_B(net3145),
    .D(_02264_),
    .Q_N(_13191_),
    .Q(\cpu.icache.r_tag[0][19] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[0][15]$_DFFE_PP_  (.CLK(clknet_leaf_137_clk),
    .RESET_B(net3146),
    .D(_02265_),
    .Q_N(_13190_),
    .Q(\cpu.icache.r_tag[0][20] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[0][16]$_DFFE_PP_  (.CLK(clknet_leaf_137_clk),
    .RESET_B(net3147),
    .D(_02266_),
    .Q_N(_13189_),
    .Q(\cpu.icache.r_tag[0][21] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[0][17]$_DFFE_PP_  (.CLK(clknet_leaf_137_clk),
    .RESET_B(net3148),
    .D(_02267_),
    .Q_N(_13188_),
    .Q(\cpu.icache.r_tag[0][22] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[0][18]$_DFFE_PP_  (.CLK(clknet_leaf_148_clk),
    .RESET_B(net3149),
    .D(_02268_),
    .Q_N(_13187_),
    .Q(\cpu.icache.r_tag[0][23] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[0][1]$_DFFE_PP_  (.CLK(clknet_leaf_152_clk),
    .RESET_B(net3150),
    .D(_02269_),
    .Q_N(_13186_),
    .Q(\cpu.icache.r_tag[0][6] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[0][2]$_DFFE_PP_  (.CLK(clknet_leaf_153_clk),
    .RESET_B(net3151),
    .D(_02270_),
    .Q_N(_13185_),
    .Q(\cpu.icache.r_tag[0][7] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[0][3]$_DFFE_PP_  (.CLK(clknet_leaf_152_clk),
    .RESET_B(net3152),
    .D(_02271_),
    .Q_N(_13184_),
    .Q(\cpu.icache.r_tag[0][8] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[0][4]$_DFFE_PP_  (.CLK(clknet_leaf_153_clk),
    .RESET_B(net3153),
    .D(_02272_),
    .Q_N(_13183_),
    .Q(\cpu.icache.r_tag[0][9] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[0][5]$_DFFE_PP_  (.CLK(clknet_leaf_152_clk),
    .RESET_B(net3154),
    .D(_02273_),
    .Q_N(_13182_),
    .Q(\cpu.icache.r_tag[0][10] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[0][6]$_DFFE_PP_  (.CLK(clknet_leaf_150_clk),
    .RESET_B(net3155),
    .D(_02274_),
    .Q_N(_13181_),
    .Q(\cpu.icache.r_tag[0][11] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[0][7]$_DFFE_PP_  (.CLK(clknet_leaf_150_clk),
    .RESET_B(net3156),
    .D(_02275_),
    .Q_N(_13180_),
    .Q(\cpu.icache.r_tag[0][12] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[0][8]$_DFFE_PP_  (.CLK(clknet_leaf_149_clk),
    .RESET_B(net3157),
    .D(_02276_),
    .Q_N(_13179_),
    .Q(\cpu.icache.r_tag[0][13] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[0][9]$_DFFE_PP_  (.CLK(clknet_leaf_149_clk),
    .RESET_B(net3158),
    .D(_02277_),
    .Q_N(_13178_),
    .Q(\cpu.icache.r_tag[0][14] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[1][0]$_DFFE_PP_  (.CLK(clknet_leaf_157_clk),
    .RESET_B(net3159),
    .D(_02278_),
    .Q_N(_13177_),
    .Q(\cpu.icache.r_tag[1][5] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[1][10]$_DFFE_PP_  (.CLK(clknet_leaf_146_clk),
    .RESET_B(net3160),
    .D(_02279_),
    .Q_N(_13176_),
    .Q(\cpu.icache.r_tag[1][15] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[1][11]$_DFFE_PP_  (.CLK(clknet_leaf_142_clk),
    .RESET_B(net3161),
    .D(_02280_),
    .Q_N(_13175_),
    .Q(\cpu.icache.r_tag[1][16] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[1][12]$_DFFE_PP_  (.CLK(clknet_leaf_141_clk),
    .RESET_B(net3162),
    .D(_02281_),
    .Q_N(_13174_),
    .Q(\cpu.icache.r_tag[1][17] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[1][13]$_DFFE_PP_  (.CLK(clknet_leaf_137_clk),
    .RESET_B(net3163),
    .D(_02282_),
    .Q_N(_13173_),
    .Q(\cpu.icache.r_tag[1][18] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[1][14]$_DFFE_PP_  (.CLK(clknet_leaf_142_clk),
    .RESET_B(net3164),
    .D(_02283_),
    .Q_N(_13172_),
    .Q(\cpu.icache.r_tag[1][19] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[1][15]$_DFFE_PP_  (.CLK(clknet_leaf_138_clk),
    .RESET_B(net3165),
    .D(_02284_),
    .Q_N(_13171_),
    .Q(\cpu.icache.r_tag[1][20] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[1][16]$_DFFE_PP_  (.CLK(clknet_leaf_139_clk),
    .RESET_B(net3166),
    .D(_02285_),
    .Q_N(_13170_),
    .Q(\cpu.icache.r_tag[1][21] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[1][17]$_DFFE_PP_  (.CLK(clknet_leaf_138_clk),
    .RESET_B(net3167),
    .D(_02286_),
    .Q_N(_13169_),
    .Q(\cpu.icache.r_tag[1][22] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[1][18]$_DFFE_PP_  (.CLK(clknet_leaf_155_clk),
    .RESET_B(net3168),
    .D(_02287_),
    .Q_N(_13168_),
    .Q(\cpu.icache.r_tag[1][23] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[1][1]$_DFFE_PP_  (.CLK(clknet_leaf_145_clk),
    .RESET_B(net3169),
    .D(_02288_),
    .Q_N(_13167_),
    .Q(\cpu.icache.r_tag[1][6] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[1][2]$_DFFE_PP_  (.CLK(clknet_leaf_158_clk),
    .RESET_B(net3170),
    .D(_02289_),
    .Q_N(_13166_),
    .Q(\cpu.icache.r_tag[1][7] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[1][3]$_DFFE_PP_  (.CLK(clknet_leaf_155_clk),
    .RESET_B(net3171),
    .D(_02290_),
    .Q_N(_13165_),
    .Q(\cpu.icache.r_tag[1][8] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[1][4]$_DFFE_PP_  (.CLK(clknet_leaf_158_clk),
    .RESET_B(net3172),
    .D(_02291_),
    .Q_N(_13164_),
    .Q(\cpu.icache.r_tag[1][9] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[1][5]$_DFFE_PP_  (.CLK(clknet_leaf_146_clk),
    .RESET_B(net3173),
    .D(_02292_),
    .Q_N(_13163_),
    .Q(\cpu.icache.r_tag[1][10] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[1][6]$_DFFE_PP_  (.CLK(clknet_leaf_155_clk),
    .RESET_B(net3174),
    .D(_02293_),
    .Q_N(_13162_),
    .Q(\cpu.icache.r_tag[1][11] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[1][7]$_DFFE_PP_  (.CLK(clknet_leaf_147_clk),
    .RESET_B(net3175),
    .D(_02294_),
    .Q_N(_13161_),
    .Q(\cpu.icache.r_tag[1][12] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[1][8]$_DFFE_PP_  (.CLK(clknet_leaf_154_clk),
    .RESET_B(net3176),
    .D(_02295_),
    .Q_N(_13160_),
    .Q(\cpu.icache.r_tag[1][13] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[1][9]$_DFFE_PP_  (.CLK(clknet_leaf_147_clk),
    .RESET_B(net3177),
    .D(_02296_),
    .Q_N(_13159_),
    .Q(\cpu.icache.r_tag[1][14] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[2][0]$_DFFE_PP_  (.CLK(clknet_leaf_156_clk),
    .RESET_B(net3178),
    .D(_02297_),
    .Q_N(_13158_),
    .Q(\cpu.icache.r_tag[2][5] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[2][10]$_DFFE_PP_  (.CLK(clknet_leaf_143_clk),
    .RESET_B(net3179),
    .D(_02298_),
    .Q_N(_13157_),
    .Q(\cpu.icache.r_tag[2][15] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[2][11]$_DFFE_PP_  (.CLK(clknet_leaf_142_clk),
    .RESET_B(net3180),
    .D(_02299_),
    .Q_N(_13156_),
    .Q(\cpu.icache.r_tag[2][16] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[2][12]$_DFFE_PP_  (.CLK(clknet_leaf_140_clk),
    .RESET_B(net3181),
    .D(_02300_),
    .Q_N(_13155_),
    .Q(\cpu.icache.r_tag[2][17] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[2][13]$_DFFE_PP_  (.CLK(clknet_leaf_137_clk),
    .RESET_B(net3182),
    .D(_02301_),
    .Q_N(_13154_),
    .Q(\cpu.icache.r_tag[2][18] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[2][14]$_DFFE_PP_  (.CLK(clknet_leaf_140_clk),
    .RESET_B(net3183),
    .D(_02302_),
    .Q_N(_13153_),
    .Q(\cpu.icache.r_tag[2][19] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[2][15]$_DFFE_PP_  (.CLK(clknet_leaf_140_clk),
    .RESET_B(net3184),
    .D(_02303_),
    .Q_N(_13152_),
    .Q(\cpu.icache.r_tag[2][20] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[2][16]$_DFFE_PP_  (.CLK(clknet_leaf_137_clk),
    .RESET_B(net3185),
    .D(_02304_),
    .Q_N(_13151_),
    .Q(\cpu.icache.r_tag[2][21] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[2][17]$_DFFE_PP_  (.CLK(clknet_leaf_139_clk),
    .RESET_B(net3186),
    .D(_02305_),
    .Q_N(_13150_),
    .Q(\cpu.icache.r_tag[2][22] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[2][18]$_DFFE_PP_  (.CLK(clknet_leaf_147_clk),
    .RESET_B(net3187),
    .D(_02306_),
    .Q_N(_13149_),
    .Q(\cpu.icache.r_tag[2][23] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[2][1]$_DFFE_PP_  (.CLK(clknet_leaf_156_clk),
    .RESET_B(net3188),
    .D(_02307_),
    .Q_N(_13148_),
    .Q(\cpu.icache.r_tag[2][6] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[2][2]$_DFFE_PP_  (.CLK(clknet_leaf_158_clk),
    .RESET_B(net3189),
    .D(_02308_),
    .Q_N(_13147_),
    .Q(\cpu.icache.r_tag[2][7] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[2][3]$_DFFE_PP_  (.CLK(clknet_leaf_147_clk),
    .RESET_B(net3190),
    .D(_02309_),
    .Q_N(_13146_),
    .Q(\cpu.icache.r_tag[2][8] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[2][4]$_DFFE_PP_  (.CLK(clknet_leaf_159_clk),
    .RESET_B(net3191),
    .D(_02310_),
    .Q_N(_13145_),
    .Q(\cpu.icache.r_tag[2][9] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[2][5]$_DFFE_PP_  (.CLK(clknet_leaf_156_clk),
    .RESET_B(net3192),
    .D(_02311_),
    .Q_N(_13144_),
    .Q(\cpu.icache.r_tag[2][10] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[2][6]$_DFFE_PP_  (.CLK(clknet_leaf_146_clk),
    .RESET_B(net3193),
    .D(_02312_),
    .Q_N(_13143_),
    .Q(\cpu.icache.r_tag[2][11] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[2][7]$_DFFE_PP_  (.CLK(clknet_leaf_146_clk),
    .RESET_B(net3194),
    .D(_02313_),
    .Q_N(_13142_),
    .Q(\cpu.icache.r_tag[2][12] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[2][8]$_DFFE_PP_  (.CLK(clknet_leaf_155_clk),
    .RESET_B(net3195),
    .D(_02314_),
    .Q_N(_13141_),
    .Q(\cpu.icache.r_tag[2][13] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[2][9]$_DFFE_PP_  (.CLK(clknet_leaf_143_clk),
    .RESET_B(net3196),
    .D(_02315_),
    .Q_N(_13140_),
    .Q(\cpu.icache.r_tag[2][14] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[3][0]$_DFFE_PP_  (.CLK(clknet_leaf_156_clk),
    .RESET_B(net3197),
    .D(_02316_),
    .Q_N(_13139_),
    .Q(\cpu.icache.r_tag[3][5] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[3][10]$_DFFE_PP_  (.CLK(clknet_leaf_144_clk),
    .RESET_B(net3198),
    .D(_02317_),
    .Q_N(_13138_),
    .Q(\cpu.icache.r_tag[3][15] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[3][11]$_DFFE_PP_  (.CLK(clknet_leaf_148_clk),
    .RESET_B(net3199),
    .D(_02318_),
    .Q_N(_13137_),
    .Q(\cpu.icache.r_tag[3][16] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[3][12]$_DFFE_PP_  (.CLK(clknet_leaf_141_clk),
    .RESET_B(net3200),
    .D(_02319_),
    .Q_N(_13136_),
    .Q(\cpu.icache.r_tag[3][17] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[3][13]$_DFFE_PP_  (.CLK(clknet_leaf_137_clk),
    .RESET_B(net3201),
    .D(_02320_),
    .Q_N(_13135_),
    .Q(\cpu.icache.r_tag[3][18] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[3][14]$_DFFE_PP_  (.CLK(clknet_leaf_141_clk),
    .RESET_B(net3202),
    .D(_02321_),
    .Q_N(_13134_),
    .Q(\cpu.icache.r_tag[3][19] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[3][15]$_DFFE_PP_  (.CLK(clknet_leaf_142_clk),
    .RESET_B(net3203),
    .D(_02322_),
    .Q_N(_13133_),
    .Q(\cpu.icache.r_tag[3][20] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[3][16]$_DFFE_PP_  (.CLK(clknet_leaf_142_clk),
    .RESET_B(net3204),
    .D(_02323_),
    .Q_N(_13132_),
    .Q(\cpu.icache.r_tag[3][21] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[3][17]$_DFFE_PP_  (.CLK(clknet_leaf_142_clk),
    .RESET_B(net3205),
    .D(_02324_),
    .Q_N(_13131_),
    .Q(\cpu.icache.r_tag[3][22] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[3][18]$_DFFE_PP_  (.CLK(clknet_leaf_155_clk),
    .RESET_B(net3206),
    .D(_02325_),
    .Q_N(_13130_),
    .Q(\cpu.icache.r_tag[3][23] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[3][1]$_DFFE_PP_  (.CLK(clknet_leaf_144_clk),
    .RESET_B(net3207),
    .D(_02326_),
    .Q_N(_13129_),
    .Q(\cpu.icache.r_tag[3][6] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[3][2]$_DFFE_PP_  (.CLK(clknet_leaf_158_clk),
    .RESET_B(net3208),
    .D(_02327_),
    .Q_N(_13128_),
    .Q(\cpu.icache.r_tag[3][7] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[3][3]$_DFFE_PP_  (.CLK(clknet_leaf_155_clk),
    .RESET_B(net3209),
    .D(_02328_),
    .Q_N(_13127_),
    .Q(\cpu.icache.r_tag[3][8] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[3][4]$_DFFE_PP_  (.CLK(clknet_leaf_154_clk),
    .RESET_B(net3210),
    .D(_02329_),
    .Q_N(_13126_),
    .Q(\cpu.icache.r_tag[3][9] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[3][5]$_DFFE_PP_  (.CLK(clknet_leaf_145_clk),
    .RESET_B(net3211),
    .D(_02330_),
    .Q_N(_13125_),
    .Q(\cpu.icache.r_tag[3][10] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[3][6]$_DFFE_PP_  (.CLK(clknet_leaf_147_clk),
    .RESET_B(net3212),
    .D(_02331_),
    .Q_N(_13124_),
    .Q(\cpu.icache.r_tag[3][11] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[3][7]$_DFFE_PP_  (.CLK(clknet_leaf_154_clk),
    .RESET_B(net3213),
    .D(_02332_),
    .Q_N(_13123_),
    .Q(\cpu.icache.r_tag[3][12] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[3][8]$_DFFE_PP_  (.CLK(clknet_leaf_155_clk),
    .RESET_B(net3214),
    .D(_02333_),
    .Q_N(_13122_),
    .Q(\cpu.icache.r_tag[3][13] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[3][9]$_DFFE_PP_  (.CLK(clknet_leaf_148_clk),
    .RESET_B(net3215),
    .D(_02334_),
    .Q_N(_13121_),
    .Q(\cpu.icache.r_tag[3][14] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[4][0]$_DFFE_PP_  (.CLK(clknet_leaf_157_clk),
    .RESET_B(net3216),
    .D(_02335_),
    .Q_N(_13120_),
    .Q(\cpu.icache.r_tag[4][5] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[4][10]$_DFFE_PP_  (.CLK(clknet_leaf_143_clk),
    .RESET_B(net3217),
    .D(_02336_),
    .Q_N(_13119_),
    .Q(\cpu.icache.r_tag[4][15] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[4][11]$_DFFE_PP_  (.CLK(clknet_leaf_139_clk),
    .RESET_B(net3218),
    .D(_02337_),
    .Q_N(_13118_),
    .Q(\cpu.icache.r_tag[4][16] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[4][12]$_DFFE_PP_  (.CLK(clknet_leaf_140_clk),
    .RESET_B(net3219),
    .D(_02338_),
    .Q_N(_13117_),
    .Q(\cpu.icache.r_tag[4][17] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[4][13]$_DFFE_PP_  (.CLK(clknet_leaf_135_clk),
    .RESET_B(net3220),
    .D(_02339_),
    .Q_N(_13116_),
    .Q(\cpu.icache.r_tag[4][18] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[4][14]$_DFFE_PP_  (.CLK(clknet_leaf_141_clk),
    .RESET_B(net3221),
    .D(_02340_),
    .Q_N(_13115_),
    .Q(\cpu.icache.r_tag[4][19] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[4][15]$_DFFE_PP_  (.CLK(clknet_leaf_140_clk),
    .RESET_B(net3222),
    .D(_02341_),
    .Q_N(_13114_),
    .Q(\cpu.icache.r_tag[4][20] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[4][16]$_DFFE_PP_  (.CLK(clknet_leaf_139_clk),
    .RESET_B(net3223),
    .D(_02342_),
    .Q_N(_13113_),
    .Q(\cpu.icache.r_tag[4][21] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[4][17]$_DFFE_PP_  (.CLK(clknet_leaf_140_clk),
    .RESET_B(net3224),
    .D(_02343_),
    .Q_N(_13112_),
    .Q(\cpu.icache.r_tag[4][22] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[4][18]$_DFFE_PP_  (.CLK(clknet_leaf_149_clk),
    .RESET_B(net3225),
    .D(_02344_),
    .Q_N(_13111_),
    .Q(\cpu.icache.r_tag[4][23] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[4][1]$_DFFE_PP_  (.CLK(clknet_leaf_157_clk),
    .RESET_B(net3226),
    .D(_02345_),
    .Q_N(_13110_),
    .Q(\cpu.icache.r_tag[4][6] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[4][2]$_DFFE_PP_  (.CLK(clknet_leaf_157_clk),
    .RESET_B(net3227),
    .D(_02346_),
    .Q_N(_13109_),
    .Q(\cpu.icache.r_tag[4][7] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[4][3]$_DFFE_PP_  (.CLK(clknet_leaf_148_clk),
    .RESET_B(net3228),
    .D(_02347_),
    .Q_N(_13108_),
    .Q(\cpu.icache.r_tag[4][8] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[4][4]$_DFFE_PP_  (.CLK(clknet_leaf_144_clk),
    .RESET_B(net3229),
    .D(_02348_),
    .Q_N(_13107_),
    .Q(\cpu.icache.r_tag[4][9] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[4][5]$_DFFE_PP_  (.CLK(clknet_leaf_156_clk),
    .RESET_B(net3230),
    .D(_02349_),
    .Q_N(_13106_),
    .Q(\cpu.icache.r_tag[4][10] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[4][6]$_DFFE_PP_  (.CLK(clknet_leaf_146_clk),
    .RESET_B(net3231),
    .D(_02350_),
    .Q_N(_13105_),
    .Q(\cpu.icache.r_tag[4][11] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[4][7]$_DFFE_PP_  (.CLK(clknet_leaf_154_clk),
    .RESET_B(net3232),
    .D(_02351_),
    .Q_N(_13104_),
    .Q(\cpu.icache.r_tag[4][12] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[4][8]$_DFFE_PP_  (.CLK(clknet_leaf_154_clk),
    .RESET_B(net3233),
    .D(_02352_),
    .Q_N(_13103_),
    .Q(\cpu.icache.r_tag[4][13] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[4][9]$_DFFE_PP_  (.CLK(clknet_leaf_146_clk),
    .RESET_B(net3234),
    .D(_02353_),
    .Q_N(_13102_),
    .Q(\cpu.icache.r_tag[4][14] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[5][0]$_DFFE_PP_  (.CLK(clknet_leaf_145_clk),
    .RESET_B(net3235),
    .D(_02354_),
    .Q_N(_13101_),
    .Q(\cpu.icache.r_tag[5][5] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[5][10]$_DFFE_PP_  (.CLK(clknet_leaf_143_clk),
    .RESET_B(net3236),
    .D(_02355_),
    .Q_N(_13100_),
    .Q(\cpu.icache.r_tag[5][15] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[5][11]$_DFFE_PP_  (.CLK(clknet_leaf_139_clk),
    .RESET_B(net3237),
    .D(_02356_),
    .Q_N(_13099_),
    .Q(\cpu.icache.r_tag[5][16] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[5][12]$_DFFE_PP_  (.CLK(clknet_leaf_140_clk),
    .RESET_B(net3238),
    .D(_02357_),
    .Q_N(_13098_),
    .Q(\cpu.icache.r_tag[5][17] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[5][13]$_DFFE_PP_  (.CLK(clknet_leaf_136_clk),
    .RESET_B(net3239),
    .D(_02358_),
    .Q_N(_13097_),
    .Q(\cpu.icache.r_tag[5][18] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[5][14]$_DFFE_PP_  (.CLK(clknet_leaf_138_clk),
    .RESET_B(net3240),
    .D(_02359_),
    .Q_N(_13096_),
    .Q(\cpu.icache.r_tag[5][19] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[5][15]$_DFFE_PP_  (.CLK(clknet_leaf_142_clk),
    .RESET_B(net3241),
    .D(_02360_),
    .Q_N(_13095_),
    .Q(\cpu.icache.r_tag[5][20] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[5][16]$_DFFE_PP_  (.CLK(clknet_leaf_138_clk),
    .RESET_B(net3242),
    .D(_02361_),
    .Q_N(_13094_),
    .Q(\cpu.icache.r_tag[5][21] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[5][17]$_DFFE_PP_  (.CLK(clknet_leaf_138_clk),
    .RESET_B(net3243),
    .D(_02362_),
    .Q_N(_13093_),
    .Q(\cpu.icache.r_tag[5][22] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[5][18]$_DFFE_PP_  (.CLK(clknet_leaf_149_clk),
    .RESET_B(net3244),
    .D(_02363_),
    .Q_N(_13092_),
    .Q(\cpu.icache.r_tag[5][23] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[5][1]$_DFFE_PP_  (.CLK(clknet_leaf_144_clk),
    .RESET_B(net3245),
    .D(_02364_),
    .Q_N(_13091_),
    .Q(\cpu.icache.r_tag[5][6] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[5][2]$_DFFE_PP_  (.CLK(clknet_leaf_157_clk),
    .RESET_B(net3246),
    .D(_02365_),
    .Q_N(_13090_),
    .Q(\cpu.icache.r_tag[5][7] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[5][3]$_DFFE_PP_  (.CLK(clknet_leaf_147_clk),
    .RESET_B(net3247),
    .D(_02366_),
    .Q_N(_13089_),
    .Q(\cpu.icache.r_tag[5][8] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[5][4]$_DFFE_PP_  (.CLK(clknet_leaf_145_clk),
    .RESET_B(net3248),
    .D(_02367_),
    .Q_N(_13088_),
    .Q(\cpu.icache.r_tag[5][9] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[5][5]$_DFFE_PP_  (.CLK(clknet_leaf_145_clk),
    .RESET_B(net3249),
    .D(_02368_),
    .Q_N(_13087_),
    .Q(\cpu.icache.r_tag[5][10] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[5][6]$_DFFE_PP_  (.CLK(clknet_leaf_143_clk),
    .RESET_B(net3250),
    .D(_02369_),
    .Q_N(_13086_),
    .Q(\cpu.icache.r_tag[5][11] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[5][7]$_DFFE_PP_  (.CLK(clknet_leaf_146_clk),
    .RESET_B(net3251),
    .D(_02370_),
    .Q_N(_13085_),
    .Q(\cpu.icache.r_tag[5][12] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[5][8]$_DFFE_PP_  (.CLK(clknet_leaf_155_clk),
    .RESET_B(net3252),
    .D(_02371_),
    .Q_N(_13084_),
    .Q(\cpu.icache.r_tag[5][13] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[5][9]$_DFFE_PP_  (.CLK(clknet_leaf_147_clk),
    .RESET_B(net3253),
    .D(_02372_),
    .Q_N(_13083_),
    .Q(\cpu.icache.r_tag[5][14] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[6][0]$_DFFE_PP_  (.CLK(clknet_leaf_157_clk),
    .RESET_B(net3254),
    .D(_02373_),
    .Q_N(_13082_),
    .Q(\cpu.icache.r_tag[6][5] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[6][10]$_DFFE_PP_  (.CLK(clknet_leaf_143_clk),
    .RESET_B(net3255),
    .D(_02374_),
    .Q_N(_13081_),
    .Q(\cpu.icache.r_tag[6][15] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[6][11]$_DFFE_PP_  (.CLK(clknet_leaf_139_clk),
    .RESET_B(net3256),
    .D(_02375_),
    .Q_N(_13080_),
    .Q(\cpu.icache.r_tag[6][16] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[6][12]$_DFFE_PP_  (.CLK(clknet_leaf_141_clk),
    .RESET_B(net3257),
    .D(_02376_),
    .Q_N(_13079_),
    .Q(\cpu.icache.r_tag[6][17] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[6][13]$_DFFE_PP_  (.CLK(clknet_leaf_135_clk),
    .RESET_B(net3258),
    .D(_02377_),
    .Q_N(_13078_),
    .Q(\cpu.icache.r_tag[6][18] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[6][14]$_DFFE_PP_  (.CLK(clknet_leaf_141_clk),
    .RESET_B(net3259),
    .D(_02378_),
    .Q_N(_13077_),
    .Q(\cpu.icache.r_tag[6][19] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[6][15]$_DFFE_PP_  (.CLK(clknet_leaf_140_clk),
    .RESET_B(net3260),
    .D(_02379_),
    .Q_N(_13076_),
    .Q(\cpu.icache.r_tag[6][20] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[6][16]$_DFFE_PP_  (.CLK(clknet_leaf_139_clk),
    .RESET_B(net3261),
    .D(_02380_),
    .Q_N(_13075_),
    .Q(\cpu.icache.r_tag[6][21] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[6][17]$_DFFE_PP_  (.CLK(clknet_leaf_138_clk),
    .RESET_B(net3262),
    .D(_02381_),
    .Q_N(_13074_),
    .Q(\cpu.icache.r_tag[6][22] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[6][18]$_DFFE_PP_  (.CLK(clknet_leaf_148_clk),
    .RESET_B(net3263),
    .D(_02382_),
    .Q_N(_13073_),
    .Q(\cpu.icache.r_tag[6][23] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[6][1]$_DFFE_PP_  (.CLK(clknet_leaf_144_clk),
    .RESET_B(net3264),
    .D(_02383_),
    .Q_N(_13072_),
    .Q(\cpu.icache.r_tag[6][6] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[6][2]$_DFFE_PP_  (.CLK(clknet_leaf_158_clk),
    .RESET_B(net3265),
    .D(_02384_),
    .Q_N(_13071_),
    .Q(\cpu.icache.r_tag[6][7] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[6][3]$_DFFE_PP_  (.CLK(clknet_leaf_148_clk),
    .RESET_B(net3266),
    .D(_02385_),
    .Q_N(_13070_),
    .Q(\cpu.icache.r_tag[6][8] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[6][4]$_DFFE_PP_  (.CLK(clknet_leaf_144_clk),
    .RESET_B(net3267),
    .D(_02386_),
    .Q_N(_13069_),
    .Q(\cpu.icache.r_tag[6][9] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[6][5]$_DFFE_PP_  (.CLK(clknet_leaf_145_clk),
    .RESET_B(net3268),
    .D(_02387_),
    .Q_N(_13068_),
    .Q(\cpu.icache.r_tag[6][10] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[6][6]$_DFFE_PP_  (.CLK(clknet_leaf_145_clk),
    .RESET_B(net3269),
    .D(_02388_),
    .Q_N(_13067_),
    .Q(\cpu.icache.r_tag[6][11] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[6][7]$_DFFE_PP_  (.CLK(clknet_leaf_146_clk),
    .RESET_B(net3270),
    .D(_02389_),
    .Q_N(_13066_),
    .Q(\cpu.icache.r_tag[6][12] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[6][8]$_DFFE_PP_  (.CLK(clknet_leaf_159_clk),
    .RESET_B(net3271),
    .D(_02390_),
    .Q_N(_13065_),
    .Q(\cpu.icache.r_tag[6][13] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[6][9]$_DFFE_PP_  (.CLK(clknet_leaf_143_clk),
    .RESET_B(net3272),
    .D(_02391_),
    .Q_N(_13064_),
    .Q(\cpu.icache.r_tag[6][14] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[7][0]$_DFFE_PP_  (.CLK(clknet_leaf_157_clk),
    .RESET_B(net3273),
    .D(_02392_),
    .Q_N(_13063_),
    .Q(\cpu.icache.r_tag[7][5] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[7][10]$_DFFE_PP_  (.CLK(clknet_leaf_143_clk),
    .RESET_B(net3274),
    .D(_02393_),
    .Q_N(_13062_),
    .Q(\cpu.icache.r_tag[7][15] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[7][11]$_DFFE_PP_  (.CLK(clknet_leaf_139_clk),
    .RESET_B(net3275),
    .D(_02394_),
    .Q_N(_13061_),
    .Q(\cpu.icache.r_tag[7][16] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[7][12]$_DFFE_PP_  (.CLK(clknet_leaf_141_clk),
    .RESET_B(net3276),
    .D(_02395_),
    .Q_N(_13060_),
    .Q(\cpu.icache.r_tag[7][17] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[7][13]$_DFFE_PP_  (.CLK(clknet_leaf_136_clk),
    .RESET_B(net3277),
    .D(_02396_),
    .Q_N(_13059_),
    .Q(\cpu.icache.r_tag[7][18] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[7][14]$_DFFE_PP_  (.CLK(clknet_leaf_141_clk),
    .RESET_B(net3278),
    .D(_02397_),
    .Q_N(_13058_),
    .Q(\cpu.icache.r_tag[7][19] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[7][15]$_DFFE_PP_  (.CLK(clknet_leaf_138_clk),
    .RESET_B(net3279),
    .D(_02398_),
    .Q_N(_13057_),
    .Q(\cpu.icache.r_tag[7][20] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[7][16]$_DFFE_PP_  (.CLK(clknet_leaf_138_clk),
    .RESET_B(net3280),
    .D(_02399_),
    .Q_N(_13056_),
    .Q(\cpu.icache.r_tag[7][21] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[7][17]$_DFFE_PP_  (.CLK(clknet_leaf_142_clk),
    .RESET_B(net3281),
    .D(_02400_),
    .Q_N(_13055_),
    .Q(\cpu.icache.r_tag[7][22] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[7][18]$_DFFE_PP_  (.CLK(clknet_leaf_148_clk),
    .RESET_B(net3282),
    .D(_02401_),
    .Q_N(_13054_),
    .Q(\cpu.icache.r_tag[7][23] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[7][1]$_DFFE_PP_  (.CLK(clknet_leaf_144_clk),
    .RESET_B(net3283),
    .D(_02402_),
    .Q_N(_13053_),
    .Q(\cpu.icache.r_tag[7][6] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[7][2]$_DFFE_PP_  (.CLK(clknet_leaf_157_clk),
    .RESET_B(net3284),
    .D(_02403_),
    .Q_N(_13052_),
    .Q(\cpu.icache.r_tag[7][7] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[7][3]$_DFFE_PP_  (.CLK(clknet_leaf_148_clk),
    .RESET_B(net3285),
    .D(_02404_),
    .Q_N(_13051_),
    .Q(\cpu.icache.r_tag[7][8] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[7][4]$_DFFE_PP_  (.CLK(clknet_leaf_145_clk),
    .RESET_B(net3286),
    .D(_02405_),
    .Q_N(_13050_),
    .Q(\cpu.icache.r_tag[7][9] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[7][5]$_DFFE_PP_  (.CLK(clknet_leaf_156_clk),
    .RESET_B(net3287),
    .D(_02406_),
    .Q_N(_13049_),
    .Q(\cpu.icache.r_tag[7][10] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[7][6]$_DFFE_PP_  (.CLK(clknet_leaf_144_clk),
    .RESET_B(net3288),
    .D(_02407_),
    .Q_N(_13048_),
    .Q(\cpu.icache.r_tag[7][11] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[7][7]$_DFFE_PP_  (.CLK(clknet_leaf_156_clk),
    .RESET_B(net3289),
    .D(_02408_),
    .Q_N(_13047_),
    .Q(\cpu.icache.r_tag[7][12] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[7][8]$_DFFE_PP_  (.CLK(clknet_leaf_156_clk),
    .RESET_B(net3290),
    .D(_02409_),
    .Q_N(_13046_),
    .Q(\cpu.icache.r_tag[7][13] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[7][9]$_DFFE_PP_  (.CLK(clknet_leaf_147_clk),
    .RESET_B(net3291),
    .D(_02410_),
    .Q_N(_13045_),
    .Q(\cpu.icache.r_tag[7][14] ));
 sg13g2_dfrbp_1 \cpu.icache.r_valid[0]$_SDFFE_PP0P_  (.CLK(clknet_leaf_153_clk),
    .RESET_B(net3292),
    .D(_02411_),
    .Q_N(_13044_),
    .Q(\cpu.icache.r_valid[0] ));
 sg13g2_dfrbp_1 \cpu.icache.r_valid[1]$_SDFFE_PP0P_  (.CLK(clknet_leaf_154_clk),
    .RESET_B(net3293),
    .D(_02412_),
    .Q_N(_13043_),
    .Q(\cpu.icache.r_valid[1] ));
 sg13g2_dfrbp_1 \cpu.icache.r_valid[2]$_SDFFE_PP0P_  (.CLK(clknet_leaf_153_clk),
    .RESET_B(net3294),
    .D(_02413_),
    .Q_N(_13042_),
    .Q(\cpu.icache.r_valid[2] ));
 sg13g2_dfrbp_1 \cpu.icache.r_valid[3]$_SDFFE_PP0P_  (.CLK(clknet_leaf_153_clk),
    .RESET_B(net3295),
    .D(_02414_),
    .Q_N(_13041_),
    .Q(\cpu.icache.r_valid[3] ));
 sg13g2_dfrbp_1 \cpu.icache.r_valid[4]$_SDFFE_PP0P_  (.CLK(clknet_leaf_159_clk),
    .RESET_B(net3296),
    .D(_02415_),
    .Q_N(_13040_),
    .Q(\cpu.icache.r_valid[4] ));
 sg13g2_dfrbp_1 \cpu.icache.r_valid[5]$_SDFFE_PP0P_  (.CLK(clknet_leaf_161_clk),
    .RESET_B(net3297),
    .D(_02416_),
    .Q_N(_13039_),
    .Q(\cpu.icache.r_valid[5] ));
 sg13g2_dfrbp_1 \cpu.icache.r_valid[6]$_SDFFE_PP0P_  (.CLK(clknet_leaf_159_clk),
    .RESET_B(net3298),
    .D(_02417_),
    .Q_N(_13038_),
    .Q(\cpu.icache.r_valid[6] ));
 sg13g2_dfrbp_1 \cpu.icache.r_valid[7]$_SDFFE_PP0P_  (.CLK(clknet_leaf_159_clk),
    .RESET_B(net3299),
    .D(_02418_),
    .Q_N(_13037_),
    .Q(\cpu.icache.r_valid[7] ));
 sg13g2_dfrbp_1 \cpu.intr.r_clock$_SDFFE_PN0P_  (.CLK(clknet_leaf_20_clk),
    .RESET_B(net3300),
    .D(_02419_),
    .Q_N(_13036_),
    .Q(\cpu.intr.r_clock ));
 sg13g2_dfrbp_1 \cpu.intr.r_clock_cmp[0]$_DFFE_PP_  (.CLK(clknet_leaf_6_clk),
    .RESET_B(net3301),
    .D(_02420_),
    .Q_N(_13035_),
    .Q(\cpu.intr.r_clock_cmp[0] ));
 sg13g2_dfrbp_1 \cpu.intr.r_clock_cmp[10]$_DFFE_PP_  (.CLK(clknet_leaf_310_clk),
    .RESET_B(net3302),
    .D(_02421_),
    .Q_N(_13034_),
    .Q(\cpu.intr.r_clock_cmp[10] ));
 sg13g2_dfrbp_1 \cpu.intr.r_clock_cmp[11]$_DFFE_PP_  (.CLK(clknet_leaf_310_clk),
    .RESET_B(net3303),
    .D(_02422_),
    .Q_N(_13033_),
    .Q(\cpu.intr.r_clock_cmp[11] ));
 sg13g2_dfrbp_1 \cpu.intr.r_clock_cmp[12]$_DFFE_PP_  (.CLK(clknet_leaf_311_clk),
    .RESET_B(net3304),
    .D(_02423_),
    .Q_N(_13032_),
    .Q(\cpu.intr.r_clock_cmp[12] ));
 sg13g2_dfrbp_1 \cpu.intr.r_clock_cmp[13]$_DFFE_PP_  (.CLK(clknet_leaf_310_clk),
    .RESET_B(net3305),
    .D(_02424_),
    .Q_N(_13031_),
    .Q(\cpu.intr.r_clock_cmp[13] ));
 sg13g2_dfrbp_1 \cpu.intr.r_clock_cmp[14]$_DFFE_PP_  (.CLK(clknet_leaf_309_clk),
    .RESET_B(net3306),
    .D(_02425_),
    .Q_N(_13030_),
    .Q(\cpu.intr.r_clock_cmp[14] ));
 sg13g2_dfrbp_1 \cpu.intr.r_clock_cmp[15]$_DFFE_PP_  (.CLK(clknet_leaf_1_clk),
    .RESET_B(net3307),
    .D(_02426_),
    .Q_N(_13029_),
    .Q(\cpu.intr.r_clock_cmp[15] ));
 sg13g2_dfrbp_1 \cpu.intr.r_clock_cmp[16]$_DFFE_PP_  (.CLK(clknet_leaf_5_clk),
    .RESET_B(net3308),
    .D(_02427_),
    .Q_N(_13028_),
    .Q(\cpu.intr.r_clock_cmp[16] ));
 sg13g2_dfrbp_1 \cpu.intr.r_clock_cmp[17]$_DFFE_PP_  (.CLK(clknet_leaf_12_clk),
    .RESET_B(net3309),
    .D(_02428_),
    .Q_N(_13027_),
    .Q(\cpu.intr.r_clock_cmp[17] ));
 sg13g2_dfrbp_1 \cpu.intr.r_clock_cmp[18]$_DFFE_PP_  (.CLK(clknet_leaf_16_clk),
    .RESET_B(net3310),
    .D(_02429_),
    .Q_N(_13026_),
    .Q(\cpu.intr.r_clock_cmp[18] ));
 sg13g2_dfrbp_1 \cpu.intr.r_clock_cmp[19]$_DFFE_PP_  (.CLK(clknet_leaf_3_clk),
    .RESET_B(net3311),
    .D(_02430_),
    .Q_N(_13025_),
    .Q(\cpu.intr.r_clock_cmp[19] ));
 sg13g2_dfrbp_1 \cpu.intr.r_clock_cmp[1]$_DFFE_PP_  (.CLK(clknet_leaf_12_clk),
    .RESET_B(net3312),
    .D(_02431_),
    .Q_N(_13024_),
    .Q(\cpu.intr.r_clock_cmp[1] ));
 sg13g2_dfrbp_1 \cpu.intr.r_clock_cmp[20]$_DFFE_PP_  (.CLK(clknet_leaf_5_clk),
    .RESET_B(net3313),
    .D(_02432_),
    .Q_N(_13023_),
    .Q(\cpu.intr.r_clock_cmp[20] ));
 sg13g2_dfrbp_1 \cpu.intr.r_clock_cmp[21]$_DFFE_PP_  (.CLK(clknet_leaf_2_clk),
    .RESET_B(net3314),
    .D(_02433_),
    .Q_N(_13022_),
    .Q(\cpu.intr.r_clock_cmp[21] ));
 sg13g2_dfrbp_1 \cpu.intr.r_clock_cmp[22]$_DFFE_PP_  (.CLK(clknet_leaf_6_clk),
    .RESET_B(net3315),
    .D(_02434_),
    .Q_N(_13021_),
    .Q(\cpu.intr.r_clock_cmp[22] ));
 sg13g2_dfrbp_1 \cpu.intr.r_clock_cmp[23]$_DFFE_PP_  (.CLK(clknet_leaf_5_clk),
    .RESET_B(net3316),
    .D(_02435_),
    .Q_N(_13020_),
    .Q(\cpu.intr.r_clock_cmp[23] ));
 sg13g2_dfrbp_1 \cpu.intr.r_clock_cmp[24]$_DFFE_PP_  (.CLK(clknet_leaf_1_clk),
    .RESET_B(net3317),
    .D(_02436_),
    .Q_N(_13019_),
    .Q(\cpu.intr.r_clock_cmp[24] ));
 sg13g2_dfrbp_1 \cpu.intr.r_clock_cmp[25]$_DFFE_PP_  (.CLK(clknet_leaf_0_clk),
    .RESET_B(net3318),
    .D(_02437_),
    .Q_N(_13018_),
    .Q(\cpu.intr.r_clock_cmp[25] ));
 sg13g2_dfrbp_1 \cpu.intr.r_clock_cmp[26]$_DFFE_PP_  (.CLK(clknet_leaf_1_clk),
    .RESET_B(net3319),
    .D(_02438_),
    .Q_N(_13017_),
    .Q(\cpu.intr.r_clock_cmp[26] ));
 sg13g2_dfrbp_1 \cpu.intr.r_clock_cmp[27]$_DFFE_PP_  (.CLK(clknet_leaf_309_clk),
    .RESET_B(net3320),
    .D(_02439_),
    .Q_N(_13016_),
    .Q(\cpu.intr.r_clock_cmp[27] ));
 sg13g2_dfrbp_1 \cpu.intr.r_clock_cmp[28]$_DFFE_PP_  (.CLK(clknet_leaf_310_clk),
    .RESET_B(net3321),
    .D(_02440_),
    .Q_N(_13015_),
    .Q(\cpu.intr.r_clock_cmp[28] ));
 sg13g2_dfrbp_1 \cpu.intr.r_clock_cmp[29]$_DFFE_PP_  (.CLK(clknet_leaf_311_clk),
    .RESET_B(net3322),
    .D(_02441_),
    .Q_N(_13014_),
    .Q(\cpu.intr.r_clock_cmp[29] ));
 sg13g2_dfrbp_1 \cpu.intr.r_clock_cmp[2]$_DFFE_PP_  (.CLK(clknet_leaf_13_clk),
    .RESET_B(net3323),
    .D(_02442_),
    .Q_N(_13013_),
    .Q(\cpu.intr.r_clock_cmp[2] ));
 sg13g2_dfrbp_1 \cpu.intr.r_clock_cmp[30]$_DFFE_PP_  (.CLK(clknet_leaf_1_clk),
    .RESET_B(net3324),
    .D(_02443_),
    .Q_N(_13012_),
    .Q(\cpu.intr.r_clock_cmp[30] ));
 sg13g2_dfrbp_1 \cpu.intr.r_clock_cmp[31]$_DFFE_PP_  (.CLK(clknet_leaf_1_clk),
    .RESET_B(net3325),
    .D(_02444_),
    .Q_N(_13011_),
    .Q(\cpu.intr.r_clock_cmp[31] ));
 sg13g2_dfrbp_1 \cpu.intr.r_clock_cmp[3]$_DFFE_PP_  (.CLK(clknet_leaf_2_clk),
    .RESET_B(net3326),
    .D(_02445_),
    .Q_N(_13010_),
    .Q(\cpu.intr.r_clock_cmp[3] ));
 sg13g2_dfrbp_1 \cpu.intr.r_clock_cmp[4]$_DFFE_PP_  (.CLK(clknet_leaf_1_clk),
    .RESET_B(net3327),
    .D(_02446_),
    .Q_N(_13009_),
    .Q(\cpu.intr.r_clock_cmp[4] ));
 sg13g2_dfrbp_1 \cpu.intr.r_clock_cmp[5]$_DFFE_PP_  (.CLK(clknet_leaf_1_clk),
    .RESET_B(net3328),
    .D(_02447_),
    .Q_N(_13008_),
    .Q(\cpu.intr.r_clock_cmp[5] ));
 sg13g2_dfrbp_1 \cpu.intr.r_clock_cmp[6]$_DFFE_PP_  (.CLK(clknet_leaf_6_clk),
    .RESET_B(net3329),
    .D(_02448_),
    .Q_N(_13007_),
    .Q(\cpu.intr.r_clock_cmp[6] ));
 sg13g2_dfrbp_1 \cpu.intr.r_clock_cmp[7]$_DFFE_PP_  (.CLK(clknet_leaf_5_clk),
    .RESET_B(net3330),
    .D(_02449_),
    .Q_N(_13006_),
    .Q(\cpu.intr.r_clock_cmp[7] ));
 sg13g2_dfrbp_1 \cpu.intr.r_clock_cmp[8]$_DFFE_PP_  (.CLK(clknet_leaf_309_clk),
    .RESET_B(net3331),
    .D(_02450_),
    .Q_N(_13005_),
    .Q(\cpu.intr.r_clock_cmp[8] ));
 sg13g2_dfrbp_1 \cpu.intr.r_clock_cmp[9]$_DFFE_PP_  (.CLK(clknet_leaf_1_clk),
    .RESET_B(net3332),
    .D(_02451_),
    .Q_N(_15008_),
    .Q(\cpu.intr.r_clock_cmp[9] ));
 sg13g2_dfrbp_1 \cpu.intr.r_clock_count[0]$_DFF_P_  (.CLK(clknet_leaf_12_clk),
    .RESET_B(net3333),
    .D(_00036_),
    .Q_N(_00270_),
    .Q(\cpu.intr.r_clock_count[0] ));
 sg13g2_dfrbp_1 \cpu.intr.r_clock_count[10]$_DFF_P_  (.CLK(clknet_leaf_307_clk),
    .RESET_B(net3334),
    .D(_00037_),
    .Q_N(_15009_),
    .Q(\cpu.intr.r_clock_count[10] ));
 sg13g2_dfrbp_1 \cpu.intr.r_clock_count[11]$_DFF_P_  (.CLK(clknet_leaf_308_clk),
    .RESET_B(net3335),
    .D(_00038_),
    .Q_N(_15010_),
    .Q(\cpu.intr.r_clock_count[11] ));
 sg13g2_dfrbp_1 \cpu.intr.r_clock_count[12]$_DFF_P_  (.CLK(clknet_leaf_307_clk),
    .RESET_B(net3336),
    .D(_00039_),
    .Q_N(_15011_),
    .Q(\cpu.intr.r_clock_count[12] ));
 sg13g2_dfrbp_1 \cpu.intr.r_clock_count[13]$_DFF_P_  (.CLK(clknet_leaf_308_clk),
    .RESET_B(net3337),
    .D(_00040_),
    .Q_N(_15012_),
    .Q(\cpu.intr.r_clock_count[13] ));
 sg13g2_dfrbp_1 \cpu.intr.r_clock_count[14]$_DFF_P_  (.CLK(clknet_leaf_309_clk),
    .RESET_B(net3338),
    .D(_00041_),
    .Q_N(_15013_),
    .Q(\cpu.intr.r_clock_count[14] ));
 sg13g2_dfrbp_1 \cpu.intr.r_clock_count[15]$_DFF_P_  (.CLK(clknet_leaf_303_clk),
    .RESET_B(net3339),
    .D(_00042_),
    .Q_N(_13004_),
    .Q(\cpu.intr.r_clock_count[15] ));
 sg13g2_dfrbp_1 \cpu.intr.r_clock_count[16]$_DFFE_PN_  (.CLK(clknet_leaf_6_clk),
    .RESET_B(net3340),
    .D(_02452_),
    .Q_N(_13003_),
    .Q(\cpu.intr.r_clock_count[16] ));
 sg13g2_dfrbp_1 \cpu.intr.r_clock_count[17]$_DFFE_PN_  (.CLK(clknet_leaf_12_clk),
    .RESET_B(net3341),
    .D(_02453_),
    .Q_N(_13002_),
    .Q(\cpu.intr.r_clock_count[17] ));
 sg13g2_dfrbp_1 \cpu.intr.r_clock_count[18]$_DFFE_PN_  (.CLK(clknet_leaf_12_clk),
    .RESET_B(net3342),
    .D(_02454_),
    .Q_N(_13001_),
    .Q(\cpu.intr.r_clock_count[18] ));
 sg13g2_dfrbp_1 \cpu.intr.r_clock_count[19]$_DFFE_PN_  (.CLK(clknet_leaf_6_clk),
    .RESET_B(net3343),
    .D(_02455_),
    .Q_N(_15014_),
    .Q(\cpu.intr.r_clock_count[19] ));
 sg13g2_dfrbp_1 \cpu.intr.r_clock_count[1]$_DFF_P_  (.CLK(clknet_leaf_11_clk),
    .RESET_B(net3344),
    .D(_00043_),
    .Q_N(_13000_),
    .Q(\cpu.intr.r_clock_count[1] ));
 sg13g2_dfrbp_1 \cpu.intr.r_clock_count[20]$_DFFE_PN_  (.CLK(clknet_leaf_7_clk),
    .RESET_B(net3345),
    .D(_02456_),
    .Q_N(_12999_),
    .Q(\cpu.intr.r_clock_count[20] ));
 sg13g2_dfrbp_1 \cpu.intr.r_clock_count[21]$_DFFE_PN_  (.CLK(clknet_leaf_6_clk),
    .RESET_B(net3346),
    .D(_02457_),
    .Q_N(_12998_),
    .Q(\cpu.intr.r_clock_count[21] ));
 sg13g2_dfrbp_1 \cpu.intr.r_clock_count[22]$_DFFE_PN_  (.CLK(clknet_leaf_6_clk),
    .RESET_B(net3347),
    .D(_02458_),
    .Q_N(_12997_),
    .Q(\cpu.intr.r_clock_count[22] ));
 sg13g2_dfrbp_1 \cpu.intr.r_clock_count[23]$_DFFE_PN_  (.CLK(clknet_leaf_6_clk),
    .RESET_B(net3348),
    .D(_02459_),
    .Q_N(_12996_),
    .Q(\cpu.intr.r_clock_count[23] ));
 sg13g2_dfrbp_1 \cpu.intr.r_clock_count[24]$_DFFE_PN_  (.CLK(clknet_leaf_309_clk),
    .RESET_B(net3349),
    .D(_02460_),
    .Q_N(_12995_),
    .Q(\cpu.intr.r_clock_count[24] ));
 sg13g2_dfrbp_1 \cpu.intr.r_clock_count[25]$_DFFE_PN_  (.CLK(clknet_leaf_309_clk),
    .RESET_B(net3350),
    .D(_02461_),
    .Q_N(_12994_),
    .Q(\cpu.intr.r_clock_count[25] ));
 sg13g2_dfrbp_1 \cpu.intr.r_clock_count[26]$_DFFE_PN_  (.CLK(clknet_leaf_309_clk),
    .RESET_B(net3351),
    .D(_02462_),
    .Q_N(_12993_),
    .Q(\cpu.intr.r_clock_count[26] ));
 sg13g2_dfrbp_1 \cpu.intr.r_clock_count[27]$_DFFE_PN_  (.CLK(clknet_leaf_309_clk),
    .RESET_B(net3352),
    .D(_02463_),
    .Q_N(_12992_),
    .Q(\cpu.intr.r_clock_count[27] ));
 sg13g2_dfrbp_1 \cpu.intr.r_clock_count[28]$_DFFE_PN_  (.CLK(clknet_leaf_310_clk),
    .RESET_B(net3353),
    .D(_02464_),
    .Q_N(_12991_),
    .Q(\cpu.intr.r_clock_count[28] ));
 sg13g2_dfrbp_1 \cpu.intr.r_clock_count[29]$_DFFE_PN_  (.CLK(clknet_leaf_310_clk),
    .RESET_B(net3354),
    .D(_02465_),
    .Q_N(_15015_),
    .Q(\cpu.intr.r_clock_count[29] ));
 sg13g2_dfrbp_1 \cpu.intr.r_clock_count[2]$_DFF_P_  (.CLK(clknet_leaf_12_clk),
    .RESET_B(net3355),
    .D(_00044_),
    .Q_N(_12990_),
    .Q(\cpu.intr.r_clock_count[2] ));
 sg13g2_dfrbp_1 \cpu.intr.r_clock_count[30]$_DFFE_PN_  (.CLK(clknet_leaf_310_clk),
    .RESET_B(net3356),
    .D(_02466_),
    .Q_N(_12989_),
    .Q(\cpu.intr.r_clock_count[30] ));
 sg13g2_dfrbp_1 \cpu.intr.r_clock_count[31]$_DFFE_PN_  (.CLK(clknet_leaf_310_clk),
    .RESET_B(net3357),
    .D(_02467_),
    .Q_N(_15016_),
    .Q(\cpu.intr.r_clock_count[31] ));
 sg13g2_dfrbp_1 \cpu.intr.r_clock_count[3]$_DFF_P_  (.CLK(clknet_leaf_7_clk),
    .RESET_B(net3358),
    .D(_00045_),
    .Q_N(_15017_),
    .Q(\cpu.intr.r_clock_count[3] ));
 sg13g2_dfrbp_1 \cpu.intr.r_clock_count[4]$_DFF_P_  (.CLK(clknet_leaf_10_clk),
    .RESET_B(net3359),
    .D(_00046_),
    .Q_N(_15018_),
    .Q(\cpu.intr.r_clock_count[4] ));
 sg13g2_dfrbp_1 \cpu.intr.r_clock_count[5]$_DFF_P_  (.CLK(clknet_leaf_7_clk),
    .RESET_B(net3360),
    .D(_00047_),
    .Q_N(_15019_),
    .Q(\cpu.intr.r_clock_count[5] ));
 sg13g2_dfrbp_1 \cpu.intr.r_clock_count[6]$_DFF_P_  (.CLK(clknet_leaf_8_clk),
    .RESET_B(net3361),
    .D(_00048_),
    .Q_N(_15020_),
    .Q(\cpu.intr.r_clock_count[6] ));
 sg13g2_dfrbp_1 \cpu.intr.r_clock_count[7]$_DFF_P_  (.CLK(clknet_leaf_7_clk),
    .RESET_B(net3362),
    .D(_00049_),
    .Q_N(_15021_),
    .Q(\cpu.intr.r_clock_count[7] ));
 sg13g2_dfrbp_1 \cpu.intr.r_clock_count[8]$_DFF_P_  (.CLK(clknet_leaf_308_clk),
    .RESET_B(net3363),
    .D(_00050_),
    .Q_N(_15022_),
    .Q(\cpu.intr.r_clock_count[8] ));
 sg13g2_dfrbp_1 \cpu.intr.r_clock_count[9]$_DFF_P_  (.CLK(clknet_leaf_308_clk),
    .RESET_B(net3364),
    .D(_00051_),
    .Q_N(_12988_),
    .Q(\cpu.intr.r_clock_count[9] ));
 sg13g2_dfrbp_1 \cpu.intr.r_enable[0]$_SDFFE_PN0P_  (.CLK(clknet_leaf_26_clk),
    .RESET_B(net3365),
    .D(_02468_),
    .Q_N(_12987_),
    .Q(\cpu.intr.r_enable[0] ));
 sg13g2_dfrbp_1 \cpu.intr.r_enable[1]$_SDFFE_PN0P_  (.CLK(clknet_leaf_21_clk),
    .RESET_B(net3366),
    .D(_02469_),
    .Q_N(_12986_),
    .Q(\cpu.intr.r_enable[1] ));
 sg13g2_dfrbp_1 \cpu.intr.r_enable[2]$_SDFFE_PN0P_  (.CLK(clknet_leaf_21_clk),
    .RESET_B(net3367),
    .D(_02470_),
    .Q_N(_12985_),
    .Q(\cpu.intr.r_enable[2] ));
 sg13g2_dfrbp_1 \cpu.intr.r_enable[3]$_SDFFE_PN0P_  (.CLK(clknet_leaf_16_clk),
    .RESET_B(net3368),
    .D(_02471_),
    .Q_N(_12984_),
    .Q(\cpu.intr.r_enable[3] ));
 sg13g2_dfrbp_1 \cpu.intr.r_enable[4]$_SDFFE_PN0P_  (.CLK(clknet_leaf_20_clk),
    .RESET_B(net3369),
    .D(_02472_),
    .Q_N(_12983_),
    .Q(\cpu.intr.r_enable[4] ));
 sg13g2_dfrbp_1 \cpu.intr.r_enable[5]$_SDFFE_PN0P_  (.CLK(clknet_leaf_21_clk),
    .RESET_B(net3370),
    .D(_02473_),
    .Q_N(_12982_),
    .Q(\cpu.intr.r_enable[5] ));
 sg13g2_dfrbp_1 \cpu.intr.r_timer$_SDFFE_PN0P_  (.CLK(clknet_leaf_16_clk),
    .RESET_B(net3371),
    .D(_02474_),
    .Q_N(_15023_),
    .Q(\cpu.intr.r_timer ));
 sg13g2_dfrbp_1 \cpu.intr.r_timer_count[0]$_DFF_P_  (.CLK(clknet_leaf_5_clk),
    .RESET_B(net3372),
    .D(_00055_),
    .Q_N(_00269_),
    .Q(\cpu.intr.r_timer_count[0] ));
 sg13g2_dfrbp_1 \cpu.intr.r_timer_count[10]$_DFF_P_  (.CLK(clknet_leaf_312_clk),
    .RESET_B(net3373),
    .D(_00056_),
    .Q_N(_15024_),
    .Q(\cpu.intr.r_timer_count[10] ));
 sg13g2_dfrbp_1 \cpu.intr.r_timer_count[11]$_DFF_P_  (.CLK(clknet_leaf_312_clk),
    .RESET_B(net3374),
    .D(_00057_),
    .Q_N(_15025_),
    .Q(\cpu.intr.r_timer_count[11] ));
 sg13g2_dfrbp_1 \cpu.intr.r_timer_count[12]$_DFF_P_  (.CLK(clknet_leaf_312_clk),
    .RESET_B(net3375),
    .D(_00058_),
    .Q_N(_15026_),
    .Q(\cpu.intr.r_timer_count[12] ));
 sg13g2_dfrbp_1 \cpu.intr.r_timer_count[13]$_DFF_P_  (.CLK(clknet_leaf_311_clk),
    .RESET_B(net3376),
    .D(_00059_),
    .Q_N(_15027_),
    .Q(\cpu.intr.r_timer_count[13] ));
 sg13g2_dfrbp_1 \cpu.intr.r_timer_count[14]$_DFF_P_  (.CLK(clknet_leaf_312_clk),
    .RESET_B(net3377),
    .D(_00060_),
    .Q_N(_15028_),
    .Q(\cpu.intr.r_timer_count[14] ));
 sg13g2_dfrbp_1 \cpu.intr.r_timer_count[15]$_DFF_P_  (.CLK(clknet_leaf_0_clk),
    .RESET_B(net3378),
    .D(_00061_),
    .Q_N(_15029_),
    .Q(\cpu.intr.r_timer_count[15] ));
 sg13g2_dfrbp_1 \cpu.intr.r_timer_count[16]$_DFF_P_  (.CLK(clknet_leaf_15_clk),
    .RESET_B(net3379),
    .D(_00062_),
    .Q_N(_15030_),
    .Q(\cpu.intr.r_timer_count[16] ));
 sg13g2_dfrbp_1 \cpu.intr.r_timer_count[17]$_DFF_P_  (.CLK(clknet_leaf_15_clk),
    .RESET_B(net3380),
    .D(_00063_),
    .Q_N(_15031_),
    .Q(\cpu.intr.r_timer_count[17] ));
 sg13g2_dfrbp_1 \cpu.intr.r_timer_count[18]$_DFF_P_  (.CLK(clknet_leaf_16_clk),
    .RESET_B(net3381),
    .D(_00064_),
    .Q_N(_15032_),
    .Q(\cpu.intr.r_timer_count[18] ));
 sg13g2_dfrbp_1 \cpu.intr.r_timer_count[19]$_DFF_P_  (.CLK(clknet_leaf_5_clk),
    .RESET_B(net3382),
    .D(_00065_),
    .Q_N(_15033_),
    .Q(\cpu.intr.r_timer_count[19] ));
 sg13g2_dfrbp_1 \cpu.intr.r_timer_count[1]$_DFF_P_  (.CLK(clknet_leaf_2_clk),
    .RESET_B(net3383),
    .D(_00066_),
    .Q_N(_15034_),
    .Q(\cpu.intr.r_timer_count[1] ));
 sg13g2_dfrbp_1 \cpu.intr.r_timer_count[20]$_DFF_P_  (.CLK(clknet_leaf_14_clk),
    .RESET_B(net3384),
    .D(_00067_),
    .Q_N(_15035_),
    .Q(\cpu.intr.r_timer_count[20] ));
 sg13g2_dfrbp_1 \cpu.intr.r_timer_count[21]$_DFF_P_  (.CLK(clknet_leaf_13_clk),
    .RESET_B(net3385),
    .D(_00068_),
    .Q_N(_15036_),
    .Q(\cpu.intr.r_timer_count[21] ));
 sg13g2_dfrbp_1 \cpu.intr.r_timer_count[22]$_DFF_P_  (.CLK(clknet_leaf_4_clk),
    .RESET_B(net3386),
    .D(_00069_),
    .Q_N(_15037_),
    .Q(\cpu.intr.r_timer_count[22] ));
 sg13g2_dfrbp_1 \cpu.intr.r_timer_count[23]$_DFF_P_  (.CLK(clknet_leaf_13_clk),
    .RESET_B(net3387),
    .D(_00070_),
    .Q_N(_15038_),
    .Q(\cpu.intr.r_timer_count[23] ));
 sg13g2_dfrbp_1 \cpu.intr.r_timer_count[2]$_DFF_P_  (.CLK(clknet_leaf_3_clk),
    .RESET_B(net3388),
    .D(_00071_),
    .Q_N(_15039_),
    .Q(\cpu.intr.r_timer_count[2] ));
 sg13g2_dfrbp_1 \cpu.intr.r_timer_count[3]$_DFF_P_  (.CLK(clknet_leaf_3_clk),
    .RESET_B(net3389),
    .D(_00072_),
    .Q_N(_15040_),
    .Q(\cpu.intr.r_timer_count[3] ));
 sg13g2_dfrbp_1 \cpu.intr.r_timer_count[4]$_DFF_P_  (.CLK(clknet_leaf_2_clk),
    .RESET_B(net3390),
    .D(_00073_),
    .Q_N(_15041_),
    .Q(\cpu.intr.r_timer_count[4] ));
 sg13g2_dfrbp_1 \cpu.intr.r_timer_count[5]$_DFF_P_  (.CLK(clknet_leaf_3_clk),
    .RESET_B(net3391),
    .D(_00074_),
    .Q_N(_15042_),
    .Q(\cpu.intr.r_timer_count[5] ));
 sg13g2_dfrbp_1 \cpu.intr.r_timer_count[6]$_DFF_P_  (.CLK(clknet_leaf_2_clk),
    .RESET_B(net3392),
    .D(_00075_),
    .Q_N(_15043_),
    .Q(\cpu.intr.r_timer_count[6] ));
 sg13g2_dfrbp_1 \cpu.intr.r_timer_count[7]$_DFF_P_  (.CLK(clknet_leaf_0_clk),
    .RESET_B(net3393),
    .D(_00076_),
    .Q_N(_15044_),
    .Q(\cpu.intr.r_timer_count[7] ));
 sg13g2_dfrbp_1 \cpu.intr.r_timer_count[8]$_DFF_P_  (.CLK(clknet_leaf_0_clk),
    .RESET_B(net3394),
    .D(_00077_),
    .Q_N(_15045_),
    .Q(\cpu.intr.r_timer_count[8] ));
 sg13g2_dfrbp_1 \cpu.intr.r_timer_count[9]$_DFF_P_  (.CLK(clknet_leaf_0_clk),
    .RESET_B(net3395),
    .D(_00078_),
    .Q_N(_12981_),
    .Q(\cpu.intr.r_timer_count[9] ));
 sg13g2_dfrbp_1 \cpu.intr.r_timer_reload[0]$_DFFE_PP_  (.CLK(clknet_leaf_3_clk),
    .RESET_B(net3396),
    .D(_02475_),
    .Q_N(_12980_),
    .Q(\cpu.intr.r_timer_reload[0] ));
 sg13g2_dfrbp_1 \cpu.intr.r_timer_reload[10]$_DFFE_PP_  (.CLK(clknet_leaf_311_clk),
    .RESET_B(net3397),
    .D(_02476_),
    .Q_N(_12979_),
    .Q(\cpu.intr.r_timer_reload[10] ));
 sg13g2_dfrbp_1 \cpu.intr.r_timer_reload[11]$_DFFE_PP_  (.CLK(clknet_leaf_311_clk),
    .RESET_B(net3398),
    .D(_02477_),
    .Q_N(_12978_),
    .Q(\cpu.intr.r_timer_reload[11] ));
 sg13g2_dfrbp_1 \cpu.intr.r_timer_reload[12]$_DFFE_PP_  (.CLK(clknet_leaf_311_clk),
    .RESET_B(net3399),
    .D(_02478_),
    .Q_N(_12977_),
    .Q(\cpu.intr.r_timer_reload[12] ));
 sg13g2_dfrbp_1 \cpu.intr.r_timer_reload[13]$_DFFE_PP_  (.CLK(clknet_leaf_311_clk),
    .RESET_B(net3400),
    .D(_02479_),
    .Q_N(_12976_),
    .Q(\cpu.intr.r_timer_reload[13] ));
 sg13g2_dfrbp_1 \cpu.intr.r_timer_reload[14]$_DFFE_PP_  (.CLK(clknet_leaf_0_clk),
    .RESET_B(net3401),
    .D(_02480_),
    .Q_N(_12975_),
    .Q(\cpu.intr.r_timer_reload[14] ));
 sg13g2_dfrbp_1 \cpu.intr.r_timer_reload[15]$_DFFE_PP_  (.CLK(clknet_leaf_0_clk),
    .RESET_B(net3402),
    .D(_02481_),
    .Q_N(_12974_),
    .Q(\cpu.intr.r_timer_reload[15] ));
 sg13g2_dfrbp_1 \cpu.intr.r_timer_reload[16]$_DFFE_PP_  (.CLK(clknet_leaf_12_clk),
    .RESET_B(net3403),
    .D(_02482_),
    .Q_N(_12973_),
    .Q(\cpu.intr.r_timer_reload[16] ));
 sg13g2_dfrbp_1 \cpu.intr.r_timer_reload[17]$_DFFE_PP_  (.CLK(clknet_leaf_16_clk),
    .RESET_B(net3404),
    .D(_02483_),
    .Q_N(_12972_),
    .Q(\cpu.intr.r_timer_reload[17] ));
 sg13g2_dfrbp_1 \cpu.intr.r_timer_reload[18]$_DFFE_PP_  (.CLK(clknet_leaf_16_clk),
    .RESET_B(net3405),
    .D(_02484_),
    .Q_N(_12971_),
    .Q(\cpu.intr.r_timer_reload[18] ));
 sg13g2_dfrbp_1 \cpu.intr.r_timer_reload[19]$_DFFE_PP_  (.CLK(clknet_leaf_5_clk),
    .RESET_B(net3406),
    .D(_02485_),
    .Q_N(_12970_),
    .Q(\cpu.intr.r_timer_reload[19] ));
 sg13g2_dfrbp_1 \cpu.intr.r_timer_reload[1]$_DFFE_PP_  (.CLK(clknet_leaf_4_clk),
    .RESET_B(net3407),
    .D(_02486_),
    .Q_N(_12969_),
    .Q(\cpu.intr.r_timer_reload[1] ));
 sg13g2_dfrbp_1 \cpu.intr.r_timer_reload[20]$_DFFE_PP_  (.CLK(clknet_leaf_15_clk),
    .RESET_B(net3408),
    .D(_02487_),
    .Q_N(_12968_),
    .Q(\cpu.intr.r_timer_reload[20] ));
 sg13g2_dfrbp_1 \cpu.intr.r_timer_reload[21]$_DFFE_PP_  (.CLK(clknet_leaf_4_clk),
    .RESET_B(net3409),
    .D(_02488_),
    .Q_N(_12967_),
    .Q(\cpu.intr.r_timer_reload[21] ));
 sg13g2_dfrbp_1 \cpu.intr.r_timer_reload[22]$_DFFE_PP_  (.CLK(clknet_leaf_4_clk),
    .RESET_B(net3410),
    .D(_02489_),
    .Q_N(_12966_),
    .Q(\cpu.intr.r_timer_reload[22] ));
 sg13g2_dfrbp_1 \cpu.intr.r_timer_reload[23]$_DFFE_PP_  (.CLK(clknet_leaf_13_clk),
    .RESET_B(net3411),
    .D(_02490_),
    .Q_N(_12965_),
    .Q(\cpu.intr.r_timer_reload[23] ));
 sg13g2_dfrbp_1 \cpu.intr.r_timer_reload[2]$_DFFE_PP_  (.CLK(clknet_leaf_4_clk),
    .RESET_B(net3412),
    .D(_02491_),
    .Q_N(_12964_),
    .Q(\cpu.intr.r_timer_reload[2] ));
 sg13g2_dfrbp_1 \cpu.intr.r_timer_reload[3]$_DFFE_PP_  (.CLK(clknet_leaf_2_clk),
    .RESET_B(net3413),
    .D(_02492_),
    .Q_N(_12963_),
    .Q(\cpu.intr.r_timer_reload[3] ));
 sg13g2_dfrbp_1 \cpu.intr.r_timer_reload[4]$_DFFE_PP_  (.CLK(clknet_leaf_2_clk),
    .RESET_B(net3414),
    .D(_02493_),
    .Q_N(_12962_),
    .Q(\cpu.intr.r_timer_reload[4] ));
 sg13g2_dfrbp_1 \cpu.intr.r_timer_reload[5]$_DFFE_PP_  (.CLK(clknet_leaf_3_clk),
    .RESET_B(net3415),
    .D(_02494_),
    .Q_N(_12961_),
    .Q(\cpu.intr.r_timer_reload[5] ));
 sg13g2_dfrbp_1 \cpu.intr.r_timer_reload[6]$_DFFE_PP_  (.CLK(clknet_leaf_2_clk),
    .RESET_B(net3416),
    .D(_02495_),
    .Q_N(_12960_),
    .Q(\cpu.intr.r_timer_reload[6] ));
 sg13g2_dfrbp_1 \cpu.intr.r_timer_reload[7]$_DFFE_PP_  (.CLK(clknet_leaf_5_clk),
    .RESET_B(net3417),
    .D(_02496_),
    .Q_N(_12959_),
    .Q(\cpu.intr.r_timer_reload[7] ));
 sg13g2_dfrbp_1 \cpu.intr.r_timer_reload[8]$_DFFE_PP_  (.CLK(clknet_leaf_311_clk),
    .RESET_B(net3418),
    .D(_02497_),
    .Q_N(_12958_),
    .Q(\cpu.intr.r_timer_reload[8] ));
 sg13g2_dfrbp_1 \cpu.intr.r_timer_reload[9]$_DFFE_PP_  (.CLK(clknet_leaf_0_clk),
    .RESET_B(net3419),
    .D(_02498_),
    .Q_N(_12957_),
    .Q(\cpu.intr.r_timer_reload[9] ));
 sg13g2_dfrbp_1 \cpu.qspi.r_count[0]$_DFFE_PP_  (.CLK(clknet_leaf_81_clk),
    .RESET_B(net3420),
    .D(_02499_),
    .Q_N(_00173_),
    .Q(\cpu.qspi.r_count[0] ));
 sg13g2_dfrbp_1 \cpu.qspi.r_count[1]$_DFFE_PP_  (.CLK(clknet_leaf_80_clk),
    .RESET_B(net3421),
    .D(_02500_),
    .Q_N(_12956_),
    .Q(\cpu.qspi.r_count[1] ));
 sg13g2_dfrbp_1 \cpu.qspi.r_count[2]$_DFFE_PP_  (.CLK(clknet_leaf_80_clk),
    .RESET_B(net3422),
    .D(_02501_),
    .Q_N(_00174_),
    .Q(\cpu.qspi.r_count[2] ));
 sg13g2_dfrbp_1 \cpu.qspi.r_count[3]$_DFFE_PP_  (.CLK(clknet_leaf_80_clk),
    .RESET_B(net3423),
    .D(_02502_),
    .Q_N(_12955_),
    .Q(\cpu.qspi.r_count[3] ));
 sg13g2_dfrbp_1 \cpu.qspi.r_count[4]$_DFFE_PP_  (.CLK(clknet_leaf_80_clk),
    .RESET_B(net3424),
    .D(_02503_),
    .Q_N(_00236_),
    .Q(\cpu.qspi.r_count[4] ));
 sg13g2_dfrbp_1 \cpu.qspi.r_cs[0]$_SDFFE_PN1P_  (.CLK(clknet_leaf_79_clk),
    .RESET_B(net3425),
    .D(_02504_),
    .Q_N(_12954_),
    .Q(net19));
 sg13g2_dfrbp_1 \cpu.qspi.r_cs[1]$_SDFFE_PN1P_  (.CLK(clknet_leaf_79_clk),
    .RESET_B(net3426),
    .D(_02505_),
    .Q_N(_12953_),
    .Q(net20));
 sg13g2_dfrbp_1 \cpu.qspi.r_cs[2]$_SDFFE_PN1P_  (.CLK(clknet_leaf_79_clk),
    .RESET_B(net3427),
    .D(_02506_),
    .Q_N(_12952_),
    .Q(\cpu.gpio.genblk1[3].srcs_o[11] ));
 sg13g2_dfrbp_1 \cpu.qspi.r_ind$_SDFFE_PN0N_  (.CLK(clknet_leaf_84_clk),
    .RESET_B(net3428),
    .D(_02507_),
    .Q_N(_12951_),
    .Q(\cpu.qspi.r_ind ));
 sg13g2_dfrbp_1 \cpu.qspi.r_mask[0]$_SDFFE_PN0P_  (.CLK(clknet_leaf_67_clk),
    .RESET_B(net3429),
    .D(_02508_),
    .Q_N(_12950_),
    .Q(\cpu.qspi.r_mask[0] ));
 sg13g2_dfrbp_1 \cpu.qspi.r_mask[1]$_SDFFE_PN1P_  (.CLK(clknet_leaf_67_clk),
    .RESET_B(net3430),
    .D(_02509_),
    .Q_N(_12949_),
    .Q(\cpu.qspi.r_mask[1] ));
 sg13g2_dfrbp_1 \cpu.qspi.r_mask[2]$_SDFFE_PN0P_  (.CLK(clknet_leaf_67_clk),
    .RESET_B(net3431),
    .D(_02510_),
    .Q_N(_12948_),
    .Q(\cpu.qspi.r_mask[2] ));
 sg13g2_dfrbp_1 \cpu.qspi.r_quad[0]$_SDFFE_PN1P_  (.CLK(clknet_leaf_67_clk),
    .RESET_B(net3432),
    .D(_02511_),
    .Q_N(_12947_),
    .Q(\cpu.qspi.r_quad[0] ));
 sg13g2_dfrbp_1 \cpu.qspi.r_quad[1]$_SDFFE_PN0P_  (.CLK(clknet_leaf_66_clk),
    .RESET_B(net3433),
    .D(_02512_),
    .Q_N(_12946_),
    .Q(\cpu.qspi.r_quad[1] ));
 sg13g2_dfrbp_1 \cpu.qspi.r_quad[2]$_SDFFE_PN1P_  (.CLK(clknet_leaf_66_clk),
    .RESET_B(net3434),
    .D(_02513_),
    .Q_N(_12945_),
    .Q(\cpu.qspi.r_quad[2] ));
 sg13g2_dfrbp_1 \cpu.qspi.r_read_delay[0][0]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_83_clk),
    .RESET_B(net3435),
    .D(_02514_),
    .Q_N(_12944_),
    .Q(\cpu.qspi.r_read_delay[0][0] ));
 sg13g2_dfrbp_1 \cpu.qspi.r_read_delay[0][1]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_83_clk),
    .RESET_B(net3436),
    .D(_02515_),
    .Q_N(_12943_),
    .Q(\cpu.qspi.r_read_delay[0][1] ));
 sg13g2_dfrbp_1 \cpu.qspi.r_read_delay[0][2]$_SDFFCE_PN1P_  (.CLK(clknet_leaf_84_clk),
    .RESET_B(net3437),
    .D(_02516_),
    .Q_N(_12942_),
    .Q(\cpu.qspi.r_read_delay[0][2] ));
 sg13g2_dfrbp_1 \cpu.qspi.r_read_delay[0][3]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_78_clk),
    .RESET_B(net3438),
    .D(_02517_),
    .Q_N(_12941_),
    .Q(\cpu.qspi.r_read_delay[0][3] ));
 sg13g2_dfrbp_1 \cpu.qspi.r_read_delay[1][0]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_83_clk),
    .RESET_B(net3439),
    .D(_02518_),
    .Q_N(_12940_),
    .Q(\cpu.qspi.r_read_delay[1][0] ));
 sg13g2_dfrbp_1 \cpu.qspi.r_read_delay[1][1]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_78_clk),
    .RESET_B(net3440),
    .D(_02519_),
    .Q_N(_12939_),
    .Q(\cpu.qspi.r_read_delay[1][1] ));
 sg13g2_dfrbp_1 \cpu.qspi.r_read_delay[1][2]$_SDFFCE_PN1P_  (.CLK(clknet_leaf_84_clk),
    .RESET_B(net3441),
    .D(_02520_),
    .Q_N(_12938_),
    .Q(\cpu.qspi.r_read_delay[1][2] ));
 sg13g2_dfrbp_1 \cpu.qspi.r_read_delay[1][3]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_83_clk),
    .RESET_B(net3442),
    .D(_02521_),
    .Q_N(_12937_),
    .Q(\cpu.qspi.r_read_delay[1][3] ));
 sg13g2_dfrbp_1 \cpu.qspi.r_read_delay[2][0]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_82_clk),
    .RESET_B(net3443),
    .D(_02522_),
    .Q_N(_12936_),
    .Q(\cpu.qspi.r_read_delay[2][0] ));
 sg13g2_dfrbp_1 \cpu.qspi.r_read_delay[2][1]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_84_clk),
    .RESET_B(net3444),
    .D(_02523_),
    .Q_N(_12935_),
    .Q(\cpu.qspi.r_read_delay[2][1] ));
 sg13g2_dfrbp_1 \cpu.qspi.r_read_delay[2][2]$_SDFFCE_PN1P_  (.CLK(clknet_leaf_84_clk),
    .RESET_B(net3445),
    .D(_02524_),
    .Q_N(_12934_),
    .Q(\cpu.qspi.r_read_delay[2][2] ));
 sg13g2_dfrbp_1 \cpu.qspi.r_read_delay[2][3]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_83_clk),
    .RESET_B(net3446),
    .D(_02525_),
    .Q_N(_12933_),
    .Q(\cpu.qspi.r_read_delay[2][3] ));
 sg13g2_dfrbp_1 \cpu.qspi.r_rom_mode[0]$_SDFFE_PN1P_  (.CLK(clknet_leaf_66_clk),
    .RESET_B(net3447),
    .D(_02526_),
    .Q_N(_12932_),
    .Q(\cpu.qspi.r_rom_mode[0] ));
 sg13g2_dfrbp_1 \cpu.qspi.r_rom_mode[1]$_SDFFE_PN1P_  (.CLK(clknet_leaf_66_clk),
    .RESET_B(net3448),
    .D(_02527_),
    .Q_N(_15046_),
    .Q(\cpu.qspi.r_rom_mode[1] ));
 sg13g2_dfrbp_1 \cpu.qspi.r_rstrobe_d$_DFF_P_  (.CLK(clknet_leaf_66_clk),
    .RESET_B(net3449),
    .D(\cpu.qspi.c_rstrobe_d ),
    .Q_N(_15047_),
    .Q(\cpu.d_rstrobe_d ));
 sg13g2_dfrbp_1 \cpu.qspi.r_state[0]$_DFF_P_  (.CLK(clknet_leaf_82_clk),
    .RESET_B(net3450),
    .D(_00021_),
    .Q_N(_00261_),
    .Q(\cpu.qspi.r_state[0] ));
 sg13g2_dfrbp_1 \cpu.qspi.r_state[10]$_DFF_P_  (.CLK(clknet_leaf_81_clk),
    .RESET_B(net3451),
    .D(_00008_),
    .Q_N(_15048_),
    .Q(\cpu.qspi.r_state[10] ));
 sg13g2_dfrbp_1 \cpu.qspi.r_state[11]$_DFF_P_  (.CLK(clknet_leaf_86_clk),
    .RESET_B(net3452),
    .D(_00022_),
    .Q_N(_15049_),
    .Q(\cpu.qspi.r_state[11] ));
 sg13g2_dfrbp_1 \cpu.qspi.r_state[12]$_DFF_P_  (.CLK(clknet_leaf_82_clk),
    .RESET_B(net3453),
    .D(_00023_),
    .Q_N(_15050_),
    .Q(\cpu.qspi.r_state[12] ));
 sg13g2_dfrbp_1 \cpu.qspi.r_state[13]$_DFF_P_  (.CLK(clknet_leaf_85_clk),
    .RESET_B(net3454),
    .D(_00009_),
    .Q_N(_15051_),
    .Q(\cpu.qspi.r_state[13] ));
 sg13g2_dfrbp_1 \cpu.qspi.r_state[14]$_DFF_P_  (.CLK(clknet_leaf_82_clk),
    .RESET_B(net3455),
    .D(_00024_),
    .Q_N(_15052_),
    .Q(\cpu.qspi.r_state[14] ));
 sg13g2_dfrbp_1 \cpu.qspi.r_state[15]$_DFF_P_  (.CLK(clknet_leaf_85_clk),
    .RESET_B(net3456),
    .D(_00010_),
    .Q_N(_15053_),
    .Q(\cpu.qspi.r_state[15] ));
 sg13g2_dfrbp_1 \cpu.qspi.r_state[16]$_DFF_P_  (.CLK(clknet_leaf_82_clk),
    .RESET_B(net3457),
    .D(_00025_),
    .Q_N(_15054_),
    .Q(\cpu.qspi.r_state[16] ));
 sg13g2_dfrbp_1 \cpu.qspi.r_state[17]$_DFF_P_  (.CLK(clknet_leaf_85_clk),
    .RESET_B(net3458),
    .D(_00026_),
    .Q_N(_15055_),
    .Q(\cpu.qspi.r_state[17] ));
 sg13g2_dfrbp_1 \cpu.qspi.r_state[1]$_DFF_P_  (.CLK(clknet_leaf_85_clk),
    .RESET_B(net3459),
    .D(_00001_),
    .Q_N(_15056_),
    .Q(\cpu.qspi.r_state[1] ));
 sg13g2_dfrbp_1 \cpu.qspi.r_state[2]$_DFF_P_  (.CLK(clknet_leaf_82_clk),
    .RESET_B(net3460),
    .D(_00027_),
    .Q_N(_15057_),
    .Q(\cpu.qspi.r_state[2] ));
 sg13g2_dfrbp_1 \cpu.qspi.r_state[3]$_DFF_P_  (.CLK(clknet_leaf_85_clk),
    .RESET_B(net3461),
    .D(_00002_),
    .Q_N(_15058_),
    .Q(\cpu.qspi.r_state[3] ));
 sg13g2_dfrbp_1 \cpu.qspi.r_state[4]$_DFF_P_  (.CLK(clknet_leaf_85_clk),
    .RESET_B(net3462),
    .D(_00028_),
    .Q_N(_15059_),
    .Q(\cpu.qspi.r_state[4] ));
 sg13g2_dfrbp_1 \cpu.qspi.r_state[5]$_DFF_P_  (.CLK(clknet_leaf_86_clk),
    .RESET_B(net3463),
    .D(_00003_),
    .Q_N(_15060_),
    .Q(\cpu.qspi.r_state[5] ));
 sg13g2_dfrbp_1 \cpu.qspi.r_state[6]$_DFF_P_  (.CLK(clknet_leaf_84_clk),
    .RESET_B(net3464),
    .D(_00004_),
    .Q_N(_15061_),
    .Q(\cpu.qspi.r_state[6] ));
 sg13g2_dfrbp_1 \cpu.qspi.r_state[7]$_DFF_P_  (.CLK(clknet_leaf_85_clk),
    .RESET_B(net3465),
    .D(_00005_),
    .Q_N(_15062_),
    .Q(\cpu.qspi.r_state[7] ));
 sg13g2_dfrbp_1 \cpu.qspi.r_state[8]$_DFF_P_  (.CLK(clknet_leaf_86_clk),
    .RESET_B(net3466),
    .D(_00006_),
    .Q_N(_00175_),
    .Q(\cpu.qspi.r_state[8] ));
 sg13g2_dfrbp_1 \cpu.qspi.r_state[9]$_DFF_P_  (.CLK(clknet_leaf_86_clk),
    .RESET_B(net3467),
    .D(_00007_),
    .Q_N(_12931_),
    .Q(\cpu.qspi.r_state[9] ));
 sg13g2_dfrbp_1 \cpu.qspi.r_uio_oe[0]$_SDFFE_PN0P_  (.CLK(clknet_leaf_80_clk),
    .RESET_B(net3468),
    .D(_02528_),
    .Q_N(_12930_),
    .Q(net3));
 sg13g2_dfrbp_1 \cpu.qspi.r_uio_oe[1]$_SDFFE_PN0P_  (.CLK(clknet_leaf_80_clk),
    .RESET_B(net3469),
    .D(_02529_),
    .Q_N(_12929_),
    .Q(net6));
 sg13g2_dfrbp_1 \cpu.qspi.r_uio_out[0]$_DFFE_PP_  (.CLK(clknet_leaf_80_clk),
    .RESET_B(net3470),
    .D(_02530_),
    .Q_N(_12928_),
    .Q(net11));
 sg13g2_dfrbp_1 \cpu.qspi.r_uio_out[1]$_DFFE_PP_  (.CLK(clknet_leaf_80_clk),
    .RESET_B(net3471),
    .D(_02531_),
    .Q_N(_12927_),
    .Q(net12));
 sg13g2_dfrbp_1 \cpu.qspi.r_uio_out[2]$_DFFE_PP_  (.CLK(clknet_leaf_81_clk),
    .RESET_B(net3472),
    .D(_02532_),
    .Q_N(_12926_),
    .Q(net13));
 sg13g2_dfrbp_1 \cpu.qspi.r_uio_out[3]$_DFFE_PP_  (.CLK(clknet_leaf_81_clk),
    .RESET_B(net3473),
    .D(_02533_),
    .Q_N(_15063_),
    .Q(net14));
 sg13g2_dfrbp_1 \cpu.qspi.r_wstrobe_d$_DFF_P_  (.CLK(clknet_leaf_51_clk),
    .RESET_B(net3474),
    .D(\cpu.qspi.c_wstrobe_d ),
    .Q_N(_15064_),
    .Q(\cpu.d_wstrobe_d ));
 sg13g2_dfrbp_1 \cpu.qspi.r_wstrobe_i$_DFF_P_  (.CLK(clknet_leaf_165_clk),
    .RESET_B(net3475),
    .D(\cpu.qspi.c_wstrobe_i ),
    .Q_N(_00237_),
    .Q(\cpu.i_wstrobe_d ));
 sg13g2_dfrbp_1 \cpu.r_clk_invert$_DFFE_PN_  (.CLK(clknet_leaf_79_clk),
    .RESET_B(net3476),
    .D(_02534_),
    .Q_N(_12925_),
    .Q(\cpu.r_clk_invert ));
 sg13g2_dfrbp_1 \cpu.spi.r_bits[0]$_SDFFE_PN1P_  (.CLK(clknet_leaf_19_clk),
    .RESET_B(net3477),
    .D(_02535_),
    .Q_N(_12924_),
    .Q(\cpu.spi.r_bits[0] ));
 sg13g2_dfrbp_1 \cpu.spi.r_bits[1]$_SDFFE_PN1P_  (.CLK(clknet_leaf_19_clk),
    .RESET_B(net3478),
    .D(_02536_),
    .Q_N(_12923_),
    .Q(\cpu.spi.r_bits[1] ));
 sg13g2_dfrbp_1 \cpu.spi.r_bits[2]$_SDFFE_PN1P_  (.CLK(clknet_leaf_19_clk),
    .RESET_B(net3479),
    .D(_02537_),
    .Q_N(_12922_),
    .Q(\cpu.spi.r_bits[2] ));
 sg13g2_dfrbp_1 \cpu.spi.r_clk_count[0][0]$_DFFE_PP_  (.CLK(clknet_leaf_17_clk),
    .RESET_B(net3480),
    .D(_02538_),
    .Q_N(_00298_),
    .Q(\cpu.spi.r_clk_count[0][0] ));
 sg13g2_dfrbp_1 \cpu.spi.r_clk_count[0][1]$_DFFE_PP_  (.CLK(clknet_leaf_15_clk),
    .RESET_B(net3481),
    .D(_02539_),
    .Q_N(_00091_),
    .Q(\cpu.spi.r_clk_count[0][1] ));
 sg13g2_dfrbp_1 \cpu.spi.r_clk_count[0][2]$_DFFE_PP_  (.CLK(clknet_leaf_19_clk),
    .RESET_B(net3482),
    .D(_02540_),
    .Q_N(_00101_),
    .Q(\cpu.spi.r_clk_count[0][2] ));
 sg13g2_dfrbp_1 \cpu.spi.r_clk_count[0][3]$_DFFE_PP_  (.CLK(clknet_leaf_18_clk),
    .RESET_B(net3483),
    .D(_02541_),
    .Q_N(_00111_),
    .Q(\cpu.spi.r_clk_count[0][3] ));
 sg13g2_dfrbp_1 \cpu.spi.r_clk_count[0][4]$_DFFE_PP_  (.CLK(clknet_leaf_18_clk),
    .RESET_B(net3484),
    .D(_02542_),
    .Q_N(_00121_),
    .Q(\cpu.spi.r_clk_count[0][4] ));
 sg13g2_dfrbp_1 \cpu.spi.r_clk_count[0][5]$_DFFE_PP_  (.CLK(clknet_leaf_18_clk),
    .RESET_B(net3485),
    .D(_02543_),
    .Q_N(_00127_),
    .Q(\cpu.spi.r_clk_count[0][5] ));
 sg13g2_dfrbp_1 \cpu.spi.r_clk_count[0][6]$_DFFE_PP_  (.CLK(clknet_leaf_18_clk),
    .RESET_B(net3486),
    .D(_02544_),
    .Q_N(_00138_),
    .Q(\cpu.spi.r_clk_count[0][6] ));
 sg13g2_dfrbp_1 \cpu.spi.r_clk_count[0][7]$_DFFE_PP_  (.CLK(clknet_leaf_17_clk),
    .RESET_B(net3487),
    .D(_02545_),
    .Q_N(_00149_),
    .Q(\cpu.spi.r_clk_count[0][7] ));
 sg13g2_dfrbp_1 \cpu.spi.r_clk_count[1][0]$_DFFE_PP_  (.CLK(clknet_leaf_17_clk),
    .RESET_B(net3488),
    .D(_02546_),
    .Q_N(_00297_),
    .Q(\cpu.spi.r_clk_count[1][0] ));
 sg13g2_dfrbp_1 \cpu.spi.r_clk_count[1][1]$_DFFE_PP_  (.CLK(clknet_leaf_17_clk),
    .RESET_B(net3489),
    .D(_02547_),
    .Q_N(_00302_),
    .Q(\cpu.spi.r_clk_count[1][1] ));
 sg13g2_dfrbp_1 \cpu.spi.r_clk_count[1][2]$_DFFE_PP_  (.CLK(clknet_leaf_19_clk),
    .RESET_B(net3490),
    .D(_02548_),
    .Q_N(_00100_),
    .Q(\cpu.spi.r_clk_count[1][2] ));
 sg13g2_dfrbp_1 \cpu.spi.r_clk_count[1][3]$_DFFE_PP_  (.CLK(clknet_leaf_18_clk),
    .RESET_B(net3491),
    .D(_02549_),
    .Q_N(_00110_),
    .Q(\cpu.spi.r_clk_count[1][3] ));
 sg13g2_dfrbp_1 \cpu.spi.r_clk_count[1][4]$_DFFE_PP_  (.CLK(clknet_leaf_18_clk),
    .RESET_B(net3492),
    .D(_02550_),
    .Q_N(_00120_),
    .Q(\cpu.spi.r_clk_count[1][4] ));
 sg13g2_dfrbp_1 \cpu.spi.r_clk_count[1][5]$_DFFE_PP_  (.CLK(clknet_leaf_18_clk),
    .RESET_B(net3493),
    .D(_02551_),
    .Q_N(_00126_),
    .Q(\cpu.spi.r_clk_count[1][5] ));
 sg13g2_dfrbp_1 \cpu.spi.r_clk_count[1][6]$_DFFE_PP_  (.CLK(clknet_leaf_18_clk),
    .RESET_B(net3494),
    .D(_02552_),
    .Q_N(_00137_),
    .Q(\cpu.spi.r_clk_count[1][6] ));
 sg13g2_dfrbp_1 \cpu.spi.r_clk_count[1][7]$_DFFE_PP_  (.CLK(clknet_leaf_17_clk),
    .RESET_B(net3495),
    .D(_02553_),
    .Q_N(_00148_),
    .Q(\cpu.spi.r_clk_count[1][7] ));
 sg13g2_dfrbp_1 \cpu.spi.r_clk_count[2][0]$_DFFE_PP_  (.CLK(clknet_leaf_17_clk),
    .RESET_B(net3496),
    .D(_02554_),
    .Q_N(_12921_),
    .Q(\cpu.spi.r_clk_count[2][0] ));
 sg13g2_dfrbp_1 \cpu.spi.r_clk_count[2][1]$_DFFE_PP_  (.CLK(clknet_leaf_17_clk),
    .RESET_B(net3497),
    .D(_02555_),
    .Q_N(_12920_),
    .Q(\cpu.spi.r_clk_count[2][1] ));
 sg13g2_dfrbp_1 \cpu.spi.r_clk_count[2][2]$_DFFE_PP_  (.CLK(clknet_leaf_16_clk),
    .RESET_B(net3498),
    .D(_02556_),
    .Q_N(_12919_),
    .Q(\cpu.spi.r_clk_count[2][2] ));
 sg13g2_dfrbp_1 \cpu.spi.r_clk_count[2][3]$_DFFE_PP_  (.CLK(clknet_leaf_14_clk),
    .RESET_B(net3499),
    .D(_02557_),
    .Q_N(_12918_),
    .Q(\cpu.spi.r_clk_count[2][3] ));
 sg13g2_dfrbp_1 \cpu.spi.r_clk_count[2][4]$_DFFE_PP_  (.CLK(clknet_leaf_15_clk),
    .RESET_B(net3500),
    .D(_02558_),
    .Q_N(_12917_),
    .Q(\cpu.spi.r_clk_count[2][4] ));
 sg13g2_dfrbp_1 \cpu.spi.r_clk_count[2][5]$_DFFE_PP_  (.CLK(clknet_leaf_15_clk),
    .RESET_B(net3501),
    .D(_02559_),
    .Q_N(_12916_),
    .Q(\cpu.spi.r_clk_count[2][5] ));
 sg13g2_dfrbp_1 \cpu.spi.r_clk_count[2][6]$_DFFE_PP_  (.CLK(clknet_leaf_15_clk),
    .RESET_B(net3502),
    .D(_02560_),
    .Q_N(_12915_),
    .Q(\cpu.spi.r_clk_count[2][6] ));
 sg13g2_dfrbp_1 \cpu.spi.r_clk_count[2][7]$_DFFE_PP_  (.CLK(clknet_leaf_17_clk),
    .RESET_B(net3503),
    .D(_02561_),
    .Q_N(_12914_),
    .Q(\cpu.spi.r_clk_count[2][7] ));
 sg13g2_dfrbp_1 \cpu.spi.r_count[0]$_DFFE_PP_  (.CLK(clknet_leaf_57_clk),
    .RESET_B(net3504),
    .D(_02562_),
    .Q_N(_12913_),
    .Q(\cpu.spi.r_count[0] ));
 sg13g2_dfrbp_1 \cpu.spi.r_count[1]$_DFFE_PP_  (.CLK(clknet_leaf_58_clk),
    .RESET_B(net3505),
    .D(_02563_),
    .Q_N(_12912_),
    .Q(\cpu.spi.r_count[1] ));
 sg13g2_dfrbp_1 \cpu.spi.r_count[2]$_DFFE_PP_  (.CLK(clknet_leaf_58_clk),
    .RESET_B(net3506),
    .D(_02564_),
    .Q_N(_12911_),
    .Q(\cpu.spi.r_count[2] ));
 sg13g2_dfrbp_1 \cpu.spi.r_count[3]$_DFFE_PP_  (.CLK(clknet_leaf_57_clk),
    .RESET_B(net3507),
    .D(_02565_),
    .Q_N(_12910_),
    .Q(\cpu.spi.r_count[3] ));
 sg13g2_dfrbp_1 \cpu.spi.r_count[4]$_DFFE_PP_  (.CLK(clknet_leaf_58_clk),
    .RESET_B(net3508),
    .D(_02566_),
    .Q_N(_12909_),
    .Q(\cpu.spi.r_count[4] ));
 sg13g2_dfrbp_1 \cpu.spi.r_count[5]$_DFFE_PP_  (.CLK(clknet_leaf_58_clk),
    .RESET_B(net3509),
    .D(_02567_),
    .Q_N(_12908_),
    .Q(\cpu.spi.r_count[5] ));
 sg13g2_dfrbp_1 \cpu.spi.r_count[6]$_DFFE_PP_  (.CLK(clknet_leaf_58_clk),
    .RESET_B(net3510),
    .D(_02568_),
    .Q_N(_12907_),
    .Q(\cpu.spi.r_count[6] ));
 sg13g2_dfrbp_1 \cpu.spi.r_count[7]$_DFFE_PP_  (.CLK(clknet_leaf_58_clk),
    .RESET_B(net3511),
    .D(_02569_),
    .Q_N(_12906_),
    .Q(\cpu.spi.r_count[7] ));
 sg13g2_dfrbp_1 \cpu.spi.r_cs[0]$_SDFFE_PN1P_  (.CLK(clknet_leaf_60_clk),
    .RESET_B(net3512),
    .D(_02570_),
    .Q_N(_12905_),
    .Q(\cpu.gpio.genblk1[3].srcs_o[6] ));
 sg13g2_dfrbp_1 \cpu.spi.r_cs[1]$_SDFFE_PN1P_  (.CLK(clknet_leaf_60_clk),
    .RESET_B(net3513),
    .D(_02571_),
    .Q_N(_12904_),
    .Q(\cpu.gpio.genblk1[3].srcs_o[7] ));
 sg13g2_dfrbp_1 \cpu.spi.r_cs[2]$_SDFFE_PN1P_  (.CLK(clknet_leaf_60_clk),
    .RESET_B(net3514),
    .D(_02572_),
    .Q_N(_12903_),
    .Q(\cpu.gpio.genblk1[3].srcs_o[8] ));
 sg13g2_dfrbp_1 \cpu.spi.r_in[0]$_DFFE_PP_  (.CLK(clknet_leaf_60_clk),
    .RESET_B(net3515),
    .D(_02573_),
    .Q_N(_12902_),
    .Q(\cpu.spi.r_in[0] ));
 sg13g2_dfrbp_1 \cpu.spi.r_in[1]$_DFFE_PP_  (.CLK(clknet_leaf_60_clk),
    .RESET_B(net3516),
    .D(_02574_),
    .Q_N(_12901_),
    .Q(\cpu.spi.r_in[1] ));
 sg13g2_dfrbp_1 \cpu.spi.r_in[2]$_DFFE_PP_  (.CLK(clknet_leaf_60_clk),
    .RESET_B(net3517),
    .D(_02575_),
    .Q_N(_12900_),
    .Q(\cpu.spi.r_in[2] ));
 sg13g2_dfrbp_1 \cpu.spi.r_in[3]$_DFFE_PP_  (.CLK(clknet_leaf_61_clk),
    .RESET_B(net3518),
    .D(_02576_),
    .Q_N(_12899_),
    .Q(\cpu.spi.r_in[3] ));
 sg13g2_dfrbp_1 \cpu.spi.r_in[4]$_DFFE_PP_  (.CLK(clknet_leaf_58_clk),
    .RESET_B(net3519),
    .D(_02577_),
    .Q_N(_12898_),
    .Q(\cpu.spi.r_in[4] ));
 sg13g2_dfrbp_1 \cpu.spi.r_in[5]$_DFFE_PP_  (.CLK(clknet_leaf_61_clk),
    .RESET_B(net3520),
    .D(_02578_),
    .Q_N(_12897_),
    .Q(\cpu.spi.r_in[5] ));
 sg13g2_dfrbp_1 \cpu.spi.r_in[6]$_DFFE_PP_  (.CLK(clknet_leaf_61_clk),
    .RESET_B(net3521),
    .D(_02579_),
    .Q_N(_12896_),
    .Q(\cpu.spi.r_in[6] ));
 sg13g2_dfrbp_1 \cpu.spi.r_in[7]$_DFFE_PP_  (.CLK(clknet_leaf_58_clk),
    .RESET_B(net3522),
    .D(_02580_),
    .Q_N(_00206_),
    .Q(\cpu.spi.r_in[7] ));
 sg13g2_dfrbp_1 \cpu.spi.r_interrupt$_SDFFE_PN0P_  (.CLK(clknet_leaf_56_clk),
    .RESET_B(net3523),
    .D(_02581_),
    .Q_N(_12895_),
    .Q(\cpu.intr.spi_intr ));
 sg13g2_dfrbp_1 \cpu.spi.r_mode[0][0]$_DFFE_PP_  (.CLK(clknet_leaf_20_clk),
    .RESET_B(net3524),
    .D(_02582_),
    .Q_N(_00209_),
    .Q(\cpu.spi.r_mode[0][0] ));
 sg13g2_dfrbp_1 \cpu.spi.r_mode[0][1]$_DFFE_PP_  (.CLK(clknet_leaf_22_clk),
    .RESET_B(net3525),
    .D(_02583_),
    .Q_N(_12894_),
    .Q(\cpu.spi.r_mode[0][1] ));
 sg13g2_dfrbp_1 \cpu.spi.r_mode[1][0]$_DFFE_PP_  (.CLK(clknet_leaf_20_clk),
    .RESET_B(net3526),
    .D(_02584_),
    .Q_N(_12893_),
    .Q(\cpu.spi.r_mode[1][0] ));
 sg13g2_dfrbp_1 \cpu.spi.r_mode[1][1]$_DFFE_PP_  (.CLK(clknet_leaf_57_clk),
    .RESET_B(net3527),
    .D(_02585_),
    .Q_N(_12892_),
    .Q(\cpu.spi.r_mode[1][1] ));
 sg13g2_dfrbp_1 \cpu.spi.r_mode[2][0]$_DFFE_PP_  (.CLK(clknet_leaf_20_clk),
    .RESET_B(net3528),
    .D(_02586_),
    .Q_N(_12891_),
    .Q(\cpu.spi.r_mode[2][0] ));
 sg13g2_dfrbp_1 \cpu.spi.r_mode[2][1]$_DFFE_PP_  (.CLK(clknet_leaf_20_clk),
    .RESET_B(net3529),
    .D(_02587_),
    .Q_N(_12890_),
    .Q(\cpu.spi.r_mode[2][1] ));
 sg13g2_dfrbp_1 \cpu.spi.r_out[0]$_DFFE_PP_  (.CLK(clknet_leaf_57_clk),
    .RESET_B(net3530),
    .D(_02588_),
    .Q_N(_12889_),
    .Q(\cpu.spi.r_out[0] ));
 sg13g2_dfrbp_1 \cpu.spi.r_out[1]$_DFFE_PP_  (.CLK(clknet_leaf_55_clk),
    .RESET_B(net3531),
    .D(_02589_),
    .Q_N(_12888_),
    .Q(\cpu.spi.r_out[1] ));
 sg13g2_dfrbp_1 \cpu.spi.r_out[2]$_DFFE_PP_  (.CLK(clknet_leaf_55_clk),
    .RESET_B(net3532),
    .D(_02590_),
    .Q_N(_12887_),
    .Q(\cpu.spi.r_out[2] ));
 sg13g2_dfrbp_1 \cpu.spi.r_out[3]$_DFFE_PP_  (.CLK(clknet_leaf_55_clk),
    .RESET_B(net3533),
    .D(_02591_),
    .Q_N(_12886_),
    .Q(\cpu.spi.r_out[3] ));
 sg13g2_dfrbp_1 \cpu.spi.r_out[4]$_DFFE_PP_  (.CLK(clknet_leaf_55_clk),
    .RESET_B(net3534),
    .D(_02592_),
    .Q_N(_12885_),
    .Q(\cpu.spi.r_out[4] ));
 sg13g2_dfrbp_1 \cpu.spi.r_out[5]$_DFFE_PP_  (.CLK(clknet_leaf_57_clk),
    .RESET_B(net3535),
    .D(_02593_),
    .Q_N(_12884_),
    .Q(\cpu.spi.r_out[5] ));
 sg13g2_dfrbp_1 \cpu.spi.r_out[6]$_DFFE_PP_  (.CLK(clknet_leaf_56_clk),
    .RESET_B(net3536),
    .D(_02594_),
    .Q_N(_12883_),
    .Q(\cpu.spi.r_out[6] ));
 sg13g2_dfrbp_1 \cpu.spi.r_out[7]$_DFFE_PP_  (.CLK(clknet_leaf_56_clk),
    .RESET_B(net3537),
    .D(_02595_),
    .Q_N(_12882_),
    .Q(\cpu.spi.r_out[7] ));
 sg13g2_dfrbp_1 \cpu.spi.r_ready$_SDFFE_PN1P_  (.CLK(clknet_leaf_19_clk),
    .RESET_B(net3538),
    .D(_02596_),
    .Q_N(_12881_),
    .Q(\cpu.spi.r_ready ));
 sg13g2_dfrbp_1 \cpu.spi.r_searching$_SDFFE_PN0P_  (.CLK(clknet_leaf_57_clk),
    .RESET_B(net3539),
    .D(_02597_),
    .Q_N(_00205_),
    .Q(\cpu.spi.r_searching ));
 sg13g2_dfrbp_1 \cpu.spi.r_sel[0]$_DFFE_PP_  (.CLK(clknet_leaf_56_clk),
    .RESET_B(net3540),
    .D(_02598_),
    .Q_N(_12880_),
    .Q(\cpu.spi.r_sel[0] ));
 sg13g2_dfrbp_1 \cpu.spi.r_sel[1]$_DFFE_PP_  (.CLK(clknet_leaf_57_clk),
    .RESET_B(net3541),
    .D(_02599_),
    .Q_N(_12879_),
    .Q(\cpu.spi.r_sel[1] ));
 sg13g2_dfrbp_1 \cpu.spi.r_src[0]$_DFFE_PP_  (.CLK(clknet_leaf_20_clk),
    .RESET_B(net3542),
    .D(_02600_),
    .Q_N(_00266_),
    .Q(\cpu.spi.r_src[0] ));
 sg13g2_dfrbp_1 \cpu.spi.r_src[1]$_DFFE_PP_  (.CLK(clknet_leaf_19_clk),
    .RESET_B(net3543),
    .D(_02601_),
    .Q_N(_00267_),
    .Q(\cpu.spi.r_src[1] ));
 sg13g2_dfrbp_1 \cpu.spi.r_src[2]$_DFFE_PP_  (.CLK(clknet_leaf_20_clk),
    .RESET_B(net3544),
    .D(_02602_),
    .Q_N(_15065_),
    .Q(\cpu.spi.r_src[2] ));
 sg13g2_dfrbp_1 \cpu.spi.r_state[0]$_DFF_P_  (.CLK(clknet_leaf_59_clk),
    .RESET_B(net3545),
    .D(_00029_),
    .Q_N(_15066_),
    .Q(\cpu.spi.r_state[0] ));
 sg13g2_dfrbp_1 \cpu.spi.r_state[1]$_DFF_P_  (.CLK(clknet_leaf_57_clk),
    .RESET_B(net3546),
    .D(_00030_),
    .Q_N(_00210_),
    .Q(\cpu.spi.r_state[1] ));
 sg13g2_dfrbp_1 \cpu.spi.r_state[2]$_DFF_P_  (.CLK(clknet_leaf_59_clk),
    .RESET_B(net3547),
    .D(_00031_),
    .Q_N(_15067_),
    .Q(\cpu.spi.r_state[2] ));
 sg13g2_dfrbp_1 \cpu.spi.r_state[3]$_DFF_P_  (.CLK(clknet_leaf_60_clk),
    .RESET_B(net3548),
    .D(_00032_),
    .Q_N(_15068_),
    .Q(\cpu.spi.r_state[3] ));
 sg13g2_dfrbp_1 \cpu.spi.r_state[4]$_DFF_P_  (.CLK(clknet_leaf_59_clk),
    .RESET_B(net3549),
    .D(_00033_),
    .Q_N(_00262_),
    .Q(\cpu.spi.r_state[4] ));
 sg13g2_dfrbp_1 \cpu.spi.r_state[5]$_DFF_P_  (.CLK(clknet_leaf_59_clk),
    .RESET_B(net3550),
    .D(_00034_),
    .Q_N(_15069_),
    .Q(\cpu.spi.r_state[5] ));
 sg13g2_dfrbp_1 \cpu.spi.r_state[6]$_DFF_P_  (.CLK(clknet_leaf_19_clk),
    .RESET_B(net3551),
    .D(_00035_),
    .Q_N(_00211_),
    .Q(\cpu.spi.r_state[6] ));
 sg13g2_dfrbp_1 \cpu.spi.r_timeout[0]$_DFFE_PP_  (.CLK(clknet_leaf_15_clk),
    .RESET_B(net3552),
    .D(_02603_),
    .Q_N(_12878_),
    .Q(\cpu.spi.r_timeout[0] ));
 sg13g2_dfrbp_1 \cpu.spi.r_timeout[1]$_DFFE_PP_  (.CLK(clknet_leaf_13_clk),
    .RESET_B(net3553),
    .D(_02604_),
    .Q_N(_12877_),
    .Q(\cpu.spi.r_timeout[1] ));
 sg13g2_dfrbp_1 \cpu.spi.r_timeout[2]$_DFFE_PP_  (.CLK(clknet_leaf_13_clk),
    .RESET_B(net3554),
    .D(_02605_),
    .Q_N(_12876_),
    .Q(\cpu.spi.r_timeout[2] ));
 sg13g2_dfrbp_1 \cpu.spi.r_timeout[3]$_DFFE_PP_  (.CLK(clknet_leaf_14_clk),
    .RESET_B(net3555),
    .D(_02606_),
    .Q_N(_12875_),
    .Q(\cpu.spi.r_timeout[3] ));
 sg13g2_dfrbp_1 \cpu.spi.r_timeout[4]$_DFFE_PP_  (.CLK(clknet_leaf_13_clk),
    .RESET_B(net3556),
    .D(_02607_),
    .Q_N(_12874_),
    .Q(\cpu.spi.r_timeout[4] ));
 sg13g2_dfrbp_1 \cpu.spi.r_timeout[5]$_DFFE_PP_  (.CLK(clknet_leaf_14_clk),
    .RESET_B(net3557),
    .D(_02608_),
    .Q_N(_12873_),
    .Q(\cpu.spi.r_timeout[5] ));
 sg13g2_dfrbp_1 \cpu.spi.r_timeout[6]$_DFFE_PP_  (.CLK(clknet_leaf_14_clk),
    .RESET_B(net3558),
    .D(_02609_),
    .Q_N(_12872_),
    .Q(\cpu.spi.r_timeout[6] ));
 sg13g2_dfrbp_1 \cpu.spi.r_timeout[7]$_DFFE_PP_  (.CLK(clknet_leaf_14_clk),
    .RESET_B(net3559),
    .D(_02610_),
    .Q_N(_12871_),
    .Q(\cpu.spi.r_timeout[7] ));
 sg13g2_dfrbp_1 \cpu.spi.r_timeout_count[0]$_DFFE_PP_  (.CLK(clknet_leaf_4_clk),
    .RESET_B(net3560),
    .D(_02611_),
    .Q_N(_00268_),
    .Q(\cpu.spi.r_timeout_count[0] ));
 sg13g2_dfrbp_1 \cpu.spi.r_timeout_count[1]$_DFFE_PP_  (.CLK(clknet_leaf_3_clk),
    .RESET_B(net3561),
    .D(_02612_),
    .Q_N(_12870_),
    .Q(\cpu.spi.r_timeout_count[1] ));
 sg13g2_dfrbp_1 \cpu.spi.r_timeout_count[2]$_DFFE_PP_  (.CLK(clknet_leaf_3_clk),
    .RESET_B(net3562),
    .D(_02613_),
    .Q_N(_12869_),
    .Q(\cpu.spi.r_timeout_count[2] ));
 sg13g2_dfrbp_1 \cpu.spi.r_timeout_count[3]$_DFFE_PP_  (.CLK(clknet_leaf_4_clk),
    .RESET_B(net3563),
    .D(_02614_),
    .Q_N(_12868_),
    .Q(\cpu.spi.r_timeout_count[3] ));
 sg13g2_dfrbp_1 \cpu.spi.r_timeout_count[4]$_DFFE_PP_  (.CLK(clknet_leaf_4_clk),
    .RESET_B(net3564),
    .D(_02615_),
    .Q_N(_12867_),
    .Q(\cpu.spi.r_timeout_count[4] ));
 sg13g2_dfrbp_1 \cpu.spi.r_timeout_count[5]$_DFFE_PP_  (.CLK(clknet_leaf_13_clk),
    .RESET_B(net3565),
    .D(_02616_),
    .Q_N(_12866_),
    .Q(\cpu.spi.r_timeout_count[5] ));
 sg13g2_dfrbp_1 \cpu.spi.r_timeout_count[6]$_DFFE_PP_  (.CLK(clknet_leaf_14_clk),
    .RESET_B(net3566),
    .D(_02617_),
    .Q_N(_12865_),
    .Q(\cpu.spi.r_timeout_count[6] ));
 sg13g2_dfrbp_1 \cpu.spi.r_timeout_count[7]$_DFFE_PP_  (.CLK(clknet_leaf_14_clk),
    .RESET_B(net3567),
    .D(_02618_),
    .Q_N(_15070_),
    .Q(\cpu.spi.r_timeout_count[7] ));
 sg13g2_dfrbp_1 \cpu.uart.r_div[0]$_DFF_P_  (.CLK(clknet_leaf_62_clk),
    .RESET_B(net3568),
    .D(_00079_),
    .Q_N(_00263_),
    .Q(\cpu.uart.r_div[0] ));
 sg13g2_dfrbp_1 \cpu.uart.r_div[10]$_DFF_P_  (.CLK(clknet_leaf_70_clk),
    .RESET_B(net3569),
    .D(_00080_),
    .Q_N(_15071_),
    .Q(\cpu.uart.r_div[10] ));
 sg13g2_dfrbp_1 \cpu.uart.r_div[11]$_DFF_P_  (.CLK(clknet_leaf_71_clk),
    .RESET_B(net3570),
    .D(_00081_),
    .Q_N(_15072_),
    .Q(\cpu.uart.r_div[11] ));
 sg13g2_dfrbp_1 \cpu.uart.r_div[1]$_DFF_P_  (.CLK(clknet_leaf_62_clk),
    .RESET_B(net3571),
    .D(_00082_),
    .Q_N(_15073_),
    .Q(\cpu.uart.r_div[1] ));
 sg13g2_dfrbp_1 \cpu.uart.r_div[2]$_DFF_P_  (.CLK(clknet_leaf_62_clk),
    .RESET_B(net3572),
    .D(_00083_),
    .Q_N(_15074_),
    .Q(\cpu.uart.r_div[2] ));
 sg13g2_dfrbp_1 \cpu.uart.r_div[3]$_DFF_P_  (.CLK(clknet_leaf_61_clk),
    .RESET_B(net3573),
    .D(_00084_),
    .Q_N(_15075_),
    .Q(\cpu.uart.r_div[3] ));
 sg13g2_dfrbp_1 \cpu.uart.r_div[4]$_DFF_P_  (.CLK(clknet_leaf_61_clk),
    .RESET_B(net3574),
    .D(_00085_),
    .Q_N(_15076_),
    .Q(\cpu.uart.r_div[4] ));
 sg13g2_dfrbp_1 \cpu.uart.r_div[5]$_DFF_P_  (.CLK(clknet_leaf_61_clk),
    .RESET_B(net3575),
    .D(_00086_),
    .Q_N(_15077_),
    .Q(\cpu.uart.r_div[5] ));
 sg13g2_dfrbp_1 \cpu.uart.r_div[6]$_DFF_P_  (.CLK(clknet_leaf_62_clk),
    .RESET_B(net3576),
    .D(_00087_),
    .Q_N(_15078_),
    .Q(\cpu.uart.r_div[6] ));
 sg13g2_dfrbp_1 \cpu.uart.r_div[7]$_DFF_P_  (.CLK(clknet_leaf_70_clk),
    .RESET_B(net3577),
    .D(_00088_),
    .Q_N(_15079_),
    .Q(\cpu.uart.r_div[7] ));
 sg13g2_dfrbp_1 \cpu.uart.r_div[8]$_DFF_P_  (.CLK(clknet_leaf_70_clk),
    .RESET_B(net3578),
    .D(_00089_),
    .Q_N(_15080_),
    .Q(\cpu.uart.r_div[8] ));
 sg13g2_dfrbp_1 \cpu.uart.r_div[9]$_DFF_P_  (.CLK(clknet_leaf_70_clk),
    .RESET_B(net3579),
    .D(_00090_),
    .Q_N(_12864_),
    .Q(\cpu.uart.r_div[9] ));
 sg13g2_dfrbp_1 \cpu.uart.r_div_value[0]$_SDFFE_PN1P_  (.CLK(clknet_leaf_63_clk),
    .RESET_B(net3580),
    .D(_02619_),
    .Q_N(_12863_),
    .Q(\cpu.uart.r_div_value[0] ));
 sg13g2_dfrbp_1 \cpu.uart.r_div_value[10]$_SDFFE_PN0P_  (.CLK(clknet_leaf_69_clk),
    .RESET_B(net3581),
    .D(_02620_),
    .Q_N(_12862_),
    .Q(\cpu.uart.r_div_value[10] ));
 sg13g2_dfrbp_1 \cpu.uart.r_div_value[11]$_SDFFE_PN0P_  (.CLK(clknet_leaf_70_clk),
    .RESET_B(net3582),
    .D(_02621_),
    .Q_N(_12861_),
    .Q(\cpu.uart.r_div_value[11] ));
 sg13g2_dfrbp_1 \cpu.uart.r_div_value[1]$_SDFFE_PN0P_  (.CLK(clknet_leaf_62_clk),
    .RESET_B(net3583),
    .D(_02622_),
    .Q_N(_12860_),
    .Q(\cpu.uart.r_div_value[1] ));
 sg13g2_dfrbp_1 \cpu.uart.r_div_value[2]$_SDFFE_PN0P_  (.CLK(clknet_leaf_61_clk),
    .RESET_B(net3584),
    .D(_02623_),
    .Q_N(_12859_),
    .Q(\cpu.uart.r_div_value[2] ));
 sg13g2_dfrbp_1 \cpu.uart.r_div_value[3]$_SDFFE_PN0P_  (.CLK(clknet_leaf_62_clk),
    .RESET_B(net3585),
    .D(_02624_),
    .Q_N(_12858_),
    .Q(\cpu.uart.r_div_value[3] ));
 sg13g2_dfrbp_1 \cpu.uart.r_div_value[4]$_SDFFE_PN0P_  (.CLK(clknet_leaf_61_clk),
    .RESET_B(net3586),
    .D(_02625_),
    .Q_N(_12857_),
    .Q(\cpu.uart.r_div_value[4] ));
 sg13g2_dfrbp_1 \cpu.uart.r_div_value[5]$_SDFFE_PN0P_  (.CLK(clknet_leaf_62_clk),
    .RESET_B(net3587),
    .D(_02626_),
    .Q_N(_12856_),
    .Q(\cpu.uart.r_div_value[5] ));
 sg13g2_dfrbp_1 \cpu.uart.r_div_value[6]$_SDFFE_PN0P_  (.CLK(clknet_leaf_62_clk),
    .RESET_B(net3588),
    .D(_02627_),
    .Q_N(_12855_),
    .Q(\cpu.uart.r_div_value[6] ));
 sg13g2_dfrbp_1 \cpu.uart.r_div_value[7]$_SDFFE_PN0P_  (.CLK(clknet_leaf_63_clk),
    .RESET_B(net3589),
    .D(_02628_),
    .Q_N(_12854_),
    .Q(\cpu.uart.r_div_value[7] ));
 sg13g2_dfrbp_1 \cpu.uart.r_div_value[8]$_SDFFE_PN0P_  (.CLK(clknet_leaf_70_clk),
    .RESET_B(net3590),
    .D(_02629_),
    .Q_N(_12853_),
    .Q(\cpu.uart.r_div_value[8] ));
 sg13g2_dfrbp_1 \cpu.uart.r_div_value[9]$_SDFFE_PN0P_  (.CLK(clknet_leaf_70_clk),
    .RESET_B(net3591),
    .D(_02630_),
    .Q_N(_12852_),
    .Q(\cpu.uart.r_div_value[9] ));
 sg13g2_dfrbp_1 \cpu.uart.r_ib[0]$_DFFE_PP_  (.CLK(clknet_leaf_71_clk),
    .RESET_B(net3592),
    .D(_02631_),
    .Q_N(_12851_),
    .Q(\cpu.uart.r_ib[0] ));
 sg13g2_dfrbp_1 \cpu.uart.r_ib[1]$_DFFE_PP_  (.CLK(clknet_leaf_71_clk),
    .RESET_B(net3593),
    .D(_02632_),
    .Q_N(_12850_),
    .Q(\cpu.uart.r_ib[1] ));
 sg13g2_dfrbp_1 \cpu.uart.r_ib[2]$_DFFE_PP_  (.CLK(clknet_leaf_71_clk),
    .RESET_B(net3594),
    .D(_02633_),
    .Q_N(_12849_),
    .Q(\cpu.uart.r_ib[2] ));
 sg13g2_dfrbp_1 \cpu.uart.r_ib[3]$_DFFE_PP_  (.CLK(clknet_leaf_71_clk),
    .RESET_B(net3595),
    .D(_02634_),
    .Q_N(_12848_),
    .Q(\cpu.uart.r_ib[3] ));
 sg13g2_dfrbp_1 \cpu.uart.r_ib[4]$_DFFE_PP_  (.CLK(clknet_leaf_72_clk),
    .RESET_B(net3596),
    .D(_02635_),
    .Q_N(_12847_),
    .Q(\cpu.uart.r_ib[4] ));
 sg13g2_dfrbp_1 \cpu.uart.r_ib[5]$_DFFE_PP_  (.CLK(clknet_leaf_74_clk),
    .RESET_B(net3597),
    .D(_02636_),
    .Q_N(_12846_),
    .Q(\cpu.uart.r_ib[5] ));
 sg13g2_dfrbp_1 \cpu.uart.r_ib[6]$_DFFE_PP_  (.CLK(clknet_leaf_72_clk),
    .RESET_B(net3598),
    .D(_02637_),
    .Q_N(_12845_),
    .Q(\cpu.uart.r_ib[6] ));
 sg13g2_dfrbp_1 \cpu.uart.r_in[0]$_DFFE_PP_  (.CLK(clknet_leaf_70_clk),
    .RESET_B(net3599),
    .D(_02638_),
    .Q_N(_12844_),
    .Q(\cpu.uart.r_in[0] ));
 sg13g2_dfrbp_1 \cpu.uart.r_in[1]$_DFFE_PP_  (.CLK(clknet_leaf_71_clk),
    .RESET_B(net3600),
    .D(_02639_),
    .Q_N(_12843_),
    .Q(\cpu.uart.r_in[1] ));
 sg13g2_dfrbp_1 \cpu.uart.r_in[2]$_DFFE_PP_  (.CLK(clknet_leaf_71_clk),
    .RESET_B(net3601),
    .D(_02640_),
    .Q_N(_12842_),
    .Q(\cpu.uart.r_in[2] ));
 sg13g2_dfrbp_1 \cpu.uart.r_in[3]$_DFFE_PP_  (.CLK(clknet_leaf_71_clk),
    .RESET_B(net3602),
    .D(_02641_),
    .Q_N(_12841_),
    .Q(\cpu.uart.r_in[3] ));
 sg13g2_dfrbp_1 \cpu.uart.r_in[4]$_DFFE_PP_  (.CLK(clknet_leaf_72_clk),
    .RESET_B(net3603),
    .D(_02642_),
    .Q_N(_12840_),
    .Q(\cpu.uart.r_in[4] ));
 sg13g2_dfrbp_1 \cpu.uart.r_in[5]$_DFFE_PP_  (.CLK(clknet_leaf_74_clk),
    .RESET_B(net3604),
    .D(_02643_),
    .Q_N(_12839_),
    .Q(\cpu.uart.r_in[5] ));
 sg13g2_dfrbp_1 \cpu.uart.r_in[6]$_DFFE_PP_  (.CLK(clknet_leaf_72_clk),
    .RESET_B(net3605),
    .D(_02644_),
    .Q_N(_12838_),
    .Q(\cpu.uart.r_in[6] ));
 sg13g2_dfrbp_1 \cpu.uart.r_in[7]$_DFFE_PP_  (.CLK(clknet_leaf_72_clk),
    .RESET_B(net3606),
    .D(_02645_),
    .Q_N(_12837_),
    .Q(\cpu.uart.r_in[7] ));
 sg13g2_dfrbp_1 \cpu.uart.r_out[0]$_DFFE_PP_  (.CLK(clknet_leaf_59_clk),
    .RESET_B(net3607),
    .D(_02646_),
    .Q_N(_12836_),
    .Q(\cpu.uart.r_out[0] ));
 sg13g2_dfrbp_1 \cpu.uart.r_out[1]$_DFFE_PP_  (.CLK(clknet_leaf_59_clk),
    .RESET_B(net3608),
    .D(_02647_),
    .Q_N(_12835_),
    .Q(\cpu.uart.r_out[1] ));
 sg13g2_dfrbp_1 \cpu.uart.r_out[2]$_DFFE_PP_  (.CLK(clknet_leaf_56_clk),
    .RESET_B(net3609),
    .D(_02648_),
    .Q_N(_12834_),
    .Q(\cpu.uart.r_out[2] ));
 sg13g2_dfrbp_1 \cpu.uart.r_out[3]$_DFFE_PP_  (.CLK(clknet_leaf_56_clk),
    .RESET_B(net3610),
    .D(_02649_),
    .Q_N(_12833_),
    .Q(\cpu.uart.r_out[3] ));
 sg13g2_dfrbp_1 \cpu.uart.r_out[4]$_DFFE_PP_  (.CLK(clknet_leaf_56_clk),
    .RESET_B(net3611),
    .D(_02650_),
    .Q_N(_12832_),
    .Q(\cpu.uart.r_out[4] ));
 sg13g2_dfrbp_1 \cpu.uart.r_out[5]$_DFFE_PP_  (.CLK(clknet_leaf_53_clk),
    .RESET_B(net3612),
    .D(_02651_),
    .Q_N(_12831_),
    .Q(\cpu.uart.r_out[5] ));
 sg13g2_dfrbp_1 \cpu.uart.r_out[6]$_DFFE_PP_  (.CLK(clknet_leaf_64_clk),
    .RESET_B(net3613),
    .D(_02652_),
    .Q_N(_12830_),
    .Q(\cpu.uart.r_out[6] ));
 sg13g2_dfrbp_1 \cpu.uart.r_out[7]$_DFFE_PP_  (.CLK(clknet_leaf_64_clk),
    .RESET_B(net3614),
    .D(_02653_),
    .Q_N(_15081_),
    .Q(\cpu.uart.r_out[7] ));
 sg13g2_dfrbp_1 \cpu.uart.r_r$_DFF_P_  (.CLK(clknet_leaf_72_clk),
    .RESET_B(net3615),
    .D(\cpu.gpio.uart_rx ),
    .Q_N(_12829_),
    .Q(\cpu.uart.r_r ));
 sg13g2_dfrbp_1 \cpu.uart.r_r_int$_SDFFE_PN0P_  (.CLK(clknet_leaf_60_clk),
    .RESET_B(net3616),
    .D(_02654_),
    .Q_N(_12828_),
    .Q(\cpu.uart.r_r_int ));
 sg13g2_dfrbp_1 \cpu.uart.r_r_invert$_SDFFE_PN0P_  (.CLK(clknet_leaf_72_clk),
    .RESET_B(net3617),
    .D(_02655_),
    .Q_N(_12827_),
    .Q(\cpu.uart.r_r_invert ));
 sg13g2_dfrbp_1 \cpu.uart.r_rcnt[0]$_DFFE_PP_  (.CLK(clknet_leaf_75_clk),
    .RESET_B(net3618),
    .D(_02656_),
    .Q_N(_12826_),
    .Q(\cpu.uart.r_rcnt[0] ));
 sg13g2_dfrbp_1 \cpu.uart.r_rcnt[1]$_DFFE_PP_  (.CLK(clknet_leaf_75_clk),
    .RESET_B(net3619),
    .D(_02657_),
    .Q_N(_12825_),
    .Q(\cpu.uart.r_rcnt[1] ));
 sg13g2_dfrbp_1 \cpu.uart.r_rstate[0]$_SDFFE_PN0P_  (.CLK(clknet_leaf_74_clk),
    .RESET_B(net3620),
    .D(_02658_),
    .Q_N(_12824_),
    .Q(\cpu.uart.r_rstate[0] ));
 sg13g2_dfrbp_1 \cpu.uart.r_rstate[1]$_SDFFE_PN0P_  (.CLK(clknet_leaf_75_clk),
    .RESET_B(net3621),
    .D(_02659_),
    .Q_N(_12823_),
    .Q(\cpu.uart.r_rstate[1] ));
 sg13g2_dfrbp_1 \cpu.uart.r_rstate[2]$_SDFFE_PN0P_  (.CLK(clknet_leaf_74_clk),
    .RESET_B(net3622),
    .D(_02660_),
    .Q_N(_12822_),
    .Q(\cpu.uart.r_rstate[2] ));
 sg13g2_dfrbp_1 \cpu.uart.r_rstate[3]$_SDFFE_PN0P_  (.CLK(clknet_leaf_75_clk),
    .RESET_B(net3623),
    .D(_02661_),
    .Q_N(_12821_),
    .Q(\cpu.uart.r_rstate[3] ));
 sg13g2_dfrbp_1 \cpu.uart.r_x$_DFFE_PP_  (.CLK(clknet_leaf_74_clk),
    .RESET_B(net3624),
    .D(_02662_),
    .Q_N(_12820_),
    .Q(\cpu.gpio.genblk1[3].srcs_o[1] ));
 sg13g2_dfrbp_1 \cpu.uart.r_x_int$_SDFFE_PN0P_  (.CLK(clknet_leaf_72_clk),
    .RESET_B(net3625),
    .D(_02663_),
    .Q_N(_12819_),
    .Q(\cpu.uart.r_x_int ));
 sg13g2_dfrbp_1 \cpu.uart.r_x_invert$_SDFFE_PN0P_  (.CLK(clknet_leaf_73_clk),
    .RESET_B(net3626),
    .D(_02664_),
    .Q_N(_00264_),
    .Q(\cpu.uart.r_x_invert ));
 sg13g2_dfrbp_1 \cpu.uart.r_xcnt[0]$_DFFE_PP_  (.CLK(clknet_leaf_75_clk),
    .RESET_B(net3627),
    .D(_02665_),
    .Q_N(_12818_),
    .Q(\cpu.uart.r_xcnt[0] ));
 sg13g2_dfrbp_1 \cpu.uart.r_xcnt[1]$_DFFE_PP_  (.CLK(clknet_leaf_74_clk),
    .RESET_B(net3628),
    .D(_02666_),
    .Q_N(_12817_),
    .Q(\cpu.uart.r_xcnt[1] ));
 sg13g2_dfrbp_1 \cpu.uart.r_xstate[0]$_SDFFE_PN0P_  (.CLK(clknet_leaf_74_clk),
    .RESET_B(net3629),
    .D(_02667_),
    .Q_N(_12816_),
    .Q(\cpu.uart.r_xstate[0] ));
 sg13g2_dfrbp_1 \cpu.uart.r_xstate[1]$_SDFFE_PN0P_  (.CLK(clknet_leaf_75_clk),
    .RESET_B(net3630),
    .D(_02668_),
    .Q_N(_12815_),
    .Q(\cpu.uart.r_xstate[1] ));
 sg13g2_dfrbp_1 \cpu.uart.r_xstate[2]$_SDFFE_PN0P_  (.CLK(clknet_leaf_75_clk),
    .RESET_B(net3631),
    .D(_02669_),
    .Q_N(_12814_),
    .Q(\cpu.uart.r_xstate[2] ));
 sg13g2_dfrbp_1 \cpu.uart.r_xstate[3]$_SDFFE_PN0P_  (.CLK(clknet_leaf_75_clk),
    .RESET_B(net3632),
    .D(_02670_),
    .Q_N(_15082_),
    .Q(\cpu.uart.r_xstate[3] ));
 sg13g2_dfrbp_1 \r_reset$_DFF_P_  (.CLK(clknet_leaf_79_clk),
    .RESET_B(net3633),
    .D(_00000_),
    .Q_N(_12813_),
    .Q(r_reset));
 sg13g2_buf_1 input1 (.A(ena),
    .X(net1));
 sg13g2_buf_1 input2 (.A(rst_n),
    .X(net2));
 sg13g2_buf_1 output3 (.A(net3),
    .X(uio_oe[0]));
 sg13g2_buf_1 output4 (.A(net4),
    .X(uio_oe[1]));
 sg13g2_buf_1 output5 (.A(net5),
    .X(uio_oe[2]));
 sg13g2_buf_1 output6 (.A(net6),
    .X(uio_oe[3]));
 sg13g2_buf_1 output7 (.A(net7),
    .X(uio_oe[4]));
 sg13g2_buf_1 output8 (.A(net8),
    .X(uio_oe[5]));
 sg13g2_buf_1 output9 (.A(net9),
    .X(uio_oe[6]));
 sg13g2_buf_1 output10 (.A(net10),
    .X(uio_oe[7]));
 sg13g2_buf_1 output11 (.A(net11),
    .X(uio_out[0]));
 sg13g2_buf_1 output12 (.A(net12),
    .X(uio_out[1]));
 sg13g2_buf_1 output13 (.A(net13),
    .X(uio_out[2]));
 sg13g2_buf_1 output14 (.A(net14),
    .X(uio_out[3]));
 sg13g2_buf_1 output15 (.A(net15),
    .X(uio_out[4]));
 sg13g2_buf_1 output16 (.A(net16),
    .X(uio_out[5]));
 sg13g2_buf_1 output17 (.A(net17),
    .X(uio_out[6]));
 sg13g2_buf_1 output18 (.A(net18),
    .X(uio_out[7]));
 sg13g2_buf_1 output19 (.A(net19),
    .X(uo_out[0]));
 sg13g2_buf_1 output20 (.A(net20),
    .X(uo_out[1]));
 sg13g2_buf_1 output21 (.A(net21),
    .X(uo_out[2]));
 sg13g2_buf_1 output22 (.A(net22),
    .X(uo_out[3]));
 sg13g2_buf_1 output23 (.A(net23),
    .X(uo_out[4]));
 sg13g2_buf_1 output24 (.A(net24),
    .X(uo_out[5]));
 sg13g2_buf_1 output25 (.A(net25),
    .X(uo_out[6]));
 sg13g2_buf_1 output26 (.A(net26),
    .X(uo_out[7]));
 sg13g2_buf_2 fanout27 (.A(_06808_),
    .X(net27));
 sg13g2_buf_2 fanout28 (.A(_03861_),
    .X(net28));
 sg13g2_buf_2 fanout29 (.A(_07413_),
    .X(net29));
 sg13g2_buf_2 fanout30 (.A(_07085_),
    .X(net30));
 sg13g2_buf_2 fanout31 (.A(_03887_),
    .X(net31));
 sg13g2_buf_2 fanout32 (.A(_03862_),
    .X(net32));
 sg13g2_buf_2 fanout33 (.A(_07332_),
    .X(net33));
 sg13g2_buf_2 fanout34 (.A(_06434_),
    .X(net34));
 sg13g2_buf_2 fanout35 (.A(_04221_),
    .X(net35));
 sg13g2_buf_2 fanout36 (.A(_03691_),
    .X(net36));
 sg13g2_buf_2 fanout37 (.A(_02884_),
    .X(net37));
 sg13g2_buf_2 fanout38 (.A(_02855_),
    .X(net38));
 sg13g2_buf_2 fanout39 (.A(_02827_),
    .X(net39));
 sg13g2_buf_2 fanout40 (.A(_02819_),
    .X(net40));
 sg13g2_buf_2 fanout41 (.A(_02764_),
    .X(net41));
 sg13g2_buf_2 fanout42 (.A(_02733_),
    .X(net42));
 sg13g2_buf_2 fanout43 (.A(_02708_),
    .X(net43));
 sg13g2_buf_2 fanout44 (.A(_02696_),
    .X(net44));
 sg13g2_buf_2 fanout45 (.A(_12777_),
    .X(net45));
 sg13g2_buf_2 fanout46 (.A(_12743_),
    .X(net46));
 sg13g2_buf_2 fanout47 (.A(_12718_),
    .X(net47));
 sg13g2_buf_2 fanout48 (.A(_12707_),
    .X(net48));
 sg13g2_buf_2 fanout49 (.A(_12627_),
    .X(net49));
 sg13g2_buf_2 fanout50 (.A(_12602_),
    .X(net50));
 sg13g2_buf_2 fanout51 (.A(_12594_),
    .X(net51));
 sg13g2_buf_2 fanout52 (.A(_12539_),
    .X(net52));
 sg13g2_buf_2 fanout53 (.A(_12511_),
    .X(net53));
 sg13g2_buf_2 fanout54 (.A(_12485_),
    .X(net54));
 sg13g2_buf_2 fanout55 (.A(_12474_),
    .X(net55));
 sg13g2_buf_2 fanout56 (.A(_12415_),
    .X(net56));
 sg13g2_buf_2 fanout57 (.A(_12383_),
    .X(net57));
 sg13g2_buf_2 fanout58 (.A(_12356_),
    .X(net58));
 sg13g2_buf_2 fanout59 (.A(_12346_),
    .X(net59));
 sg13g2_buf_2 fanout60 (.A(_12285_),
    .X(net60));
 sg13g2_buf_2 fanout61 (.A(_12248_),
    .X(net61));
 sg13g2_buf_2 fanout62 (.A(_12216_),
    .X(net62));
 sg13g2_buf_2 fanout63 (.A(_12203_),
    .X(net63));
 sg13g2_buf_2 fanout64 (.A(_10007_),
    .X(net64));
 sg13g2_buf_2 fanout65 (.A(_09994_),
    .X(net65));
 sg13g2_buf_2 fanout66 (.A(_09993_),
    .X(net66));
 sg13g2_buf_2 fanout67 (.A(_06787_),
    .X(net67));
 sg13g2_buf_2 fanout68 (.A(_06786_),
    .X(net68));
 sg13g2_buf_2 fanout69 (.A(_06770_),
    .X(net69));
 sg13g2_buf_2 fanout70 (.A(_06769_),
    .X(net70));
 sg13g2_buf_2 fanout71 (.A(_06761_),
    .X(net71));
 sg13g2_buf_2 fanout72 (.A(_06760_),
    .X(net72));
 sg13g2_buf_2 fanout73 (.A(_06447_),
    .X(net73));
 sg13g2_buf_2 fanout74 (.A(_06424_),
    .X(net74));
 sg13g2_buf_2 fanout75 (.A(_05007_),
    .X(net75));
 sg13g2_buf_2 fanout76 (.A(_03690_),
    .X(net76));
 sg13g2_buf_2 fanout77 (.A(_12660_),
    .X(net77));
 sg13g2_buf_2 fanout78 (.A(_12128_),
    .X(net78));
 sg13g2_buf_2 fanout79 (.A(_12058_),
    .X(net79));
 sg13g2_buf_2 fanout80 (.A(_10105_),
    .X(net80));
 sg13g2_buf_2 fanout81 (.A(_09863_),
    .X(net81));
 sg13g2_buf_2 fanout82 (.A(_07539_),
    .X(net82));
 sg13g2_buf_2 fanout83 (.A(_07513_),
    .X(net83));
 sg13g2_buf_2 fanout84 (.A(_07069_),
    .X(net84));
 sg13g2_buf_2 fanout85 (.A(_04284_),
    .X(net85));
 sg13g2_buf_2 fanout86 (.A(_04103_),
    .X(net86));
 sg13g2_buf_2 fanout87 (.A(_10806_),
    .X(net87));
 sg13g2_buf_2 fanout88 (.A(_10157_),
    .X(net88));
 sg13g2_buf_2 fanout89 (.A(_10098_),
    .X(net89));
 sg13g2_buf_2 fanout90 (.A(_10090_),
    .X(net90));
 sg13g2_buf_2 fanout91 (.A(_09303_),
    .X(net91));
 sg13g2_buf_2 fanout92 (.A(_07510_),
    .X(net92));
 sg13g2_buf_2 fanout93 (.A(_07322_),
    .X(net93));
 sg13g2_buf_2 fanout94 (.A(_07063_),
    .X(net94));
 sg13g2_buf_2 fanout95 (.A(_06904_),
    .X(net95));
 sg13g2_buf_2 fanout96 (.A(_06900_),
    .X(net96));
 sg13g2_buf_2 fanout97 (.A(_04209_),
    .X(net97));
 sg13g2_buf_2 fanout98 (.A(_11526_),
    .X(net98));
 sg13g2_buf_2 fanout99 (.A(_10805_),
    .X(net99));
 sg13g2_buf_2 fanout100 (.A(_09302_),
    .X(net100));
 sg13g2_buf_2 fanout101 (.A(_07977_),
    .X(net101));
 sg13g2_buf_2 fanout102 (.A(_07506_),
    .X(net102));
 sg13g2_buf_2 fanout103 (.A(_06757_),
    .X(net103));
 sg13g2_buf_2 fanout104 (.A(_05465_),
    .X(net104));
 sg13g2_buf_2 fanout105 (.A(_04360_),
    .X(net105));
 sg13g2_buf_2 fanout106 (.A(_04136_),
    .X(net106));
 sg13g2_buf_2 fanout107 (.A(_03799_),
    .X(net107));
 sg13g2_buf_2 fanout108 (.A(_11517_),
    .X(net108));
 sg13g2_buf_2 fanout109 (.A(_11453_),
    .X(net109));
 sg13g2_buf_2 fanout110 (.A(_10047_),
    .X(net110));
 sg13g2_buf_2 fanout111 (.A(_09845_),
    .X(net111));
 sg13g2_buf_2 fanout112 (.A(_06412_),
    .X(net112));
 sg13g2_buf_2 fanout113 (.A(_05772_),
    .X(net113));
 sg13g2_buf_2 fanout114 (.A(_05170_),
    .X(net114));
 sg13g2_buf_2 fanout115 (.A(_05039_),
    .X(net115));
 sg13g2_buf_2 fanout116 (.A(_05038_),
    .X(net116));
 sg13g2_buf_2 fanout117 (.A(_04253_),
    .X(net117));
 sg13g2_buf_2 fanout118 (.A(_04135_),
    .X(net118));
 sg13g2_buf_2 fanout119 (.A(_03804_),
    .X(net119));
 sg13g2_buf_2 fanout120 (.A(_03801_),
    .X(net120));
 sg13g2_buf_2 fanout121 (.A(_03689_),
    .X(net121));
 sg13g2_buf_2 fanout122 (.A(_03670_),
    .X(net122));
 sg13g2_buf_2 fanout123 (.A(_11516_),
    .X(net123));
 sg13g2_buf_2 fanout124 (.A(_11452_),
    .X(net124));
 sg13g2_buf_2 fanout125 (.A(_10046_),
    .X(net125));
 sg13g2_buf_2 fanout126 (.A(_09140_),
    .X(net126));
 sg13g2_buf_2 fanout127 (.A(_07873_),
    .X(net127));
 sg13g2_buf_2 fanout128 (.A(_07701_),
    .X(net128));
 sg13g2_buf_2 fanout129 (.A(_07384_),
    .X(net129));
 sg13g2_buf_2 fanout130 (.A(_05168_),
    .X(net130));
 sg13g2_buf_2 fanout131 (.A(_04302_),
    .X(net131));
 sg13g2_buf_2 fanout132 (.A(_04250_),
    .X(net132));
 sg13g2_buf_2 fanout133 (.A(_04248_),
    .X(net133));
 sg13g2_buf_2 fanout134 (.A(_04196_),
    .X(net134));
 sg13g2_buf_2 fanout135 (.A(_04187_),
    .X(net135));
 sg13g2_buf_2 fanout136 (.A(_04184_),
    .X(net136));
 sg13g2_buf_2 fanout137 (.A(_04173_),
    .X(net137));
 sg13g2_buf_2 fanout138 (.A(_04169_),
    .X(net138));
 sg13g2_buf_2 fanout139 (.A(_04166_),
    .X(net139));
 sg13g2_buf_2 fanout140 (.A(_03662_),
    .X(net140));
 sg13g2_buf_2 fanout141 (.A(_03553_),
    .X(net141));
 sg13g2_buf_2 fanout142 (.A(_03175_),
    .X(net142));
 sg13g2_buf_2 fanout143 (.A(_11943_),
    .X(net143));
 sg13g2_buf_2 fanout144 (.A(_11808_),
    .X(net144));
 sg13g2_buf_2 fanout145 (.A(_09897_),
    .X(net145));
 sg13g2_buf_2 fanout146 (.A(_09148_),
    .X(net146));
 sg13g2_buf_2 fanout147 (.A(_09138_),
    .X(net147));
 sg13g2_buf_2 fanout148 (.A(_09134_),
    .X(net148));
 sg13g2_buf_2 fanout149 (.A(_09123_),
    .X(net149));
 sg13g2_buf_2 fanout150 (.A(_09102_),
    .X(net150));
 sg13g2_buf_2 fanout151 (.A(_08904_),
    .X(net151));
 sg13g2_buf_2 fanout152 (.A(_05167_),
    .X(net152));
 sg13g2_buf_2 fanout153 (.A(_05165_),
    .X(net153));
 sg13g2_buf_2 fanout154 (.A(_04188_),
    .X(net154));
 sg13g2_buf_2 fanout155 (.A(_04186_),
    .X(net155));
 sg13g2_buf_2 fanout156 (.A(_04183_),
    .X(net156));
 sg13g2_buf_2 fanout157 (.A(_04172_),
    .X(net157));
 sg13g2_buf_2 fanout158 (.A(_04163_),
    .X(net158));
 sg13g2_buf_2 fanout159 (.A(_04143_),
    .X(net159));
 sg13g2_buf_2 fanout160 (.A(_03641_),
    .X(net160));
 sg13g2_buf_2 fanout161 (.A(_03567_),
    .X(net161));
 sg13g2_buf_2 fanout162 (.A(_03248_),
    .X(net162));
 sg13g2_buf_2 fanout163 (.A(_03124_),
    .X(net163));
 sg13g2_buf_2 fanout164 (.A(_03045_),
    .X(net164));
 sg13g2_buf_2 fanout165 (.A(_03042_),
    .X(net165));
 sg13g2_buf_2 fanout166 (.A(_03024_),
    .X(net166));
 sg13g2_buf_2 fanout167 (.A(_11422_),
    .X(net167));
 sg13g2_buf_2 fanout168 (.A(_11417_),
    .X(net168));
 sg13g2_buf_2 fanout169 (.A(_10523_),
    .X(net169));
 sg13g2_buf_2 fanout170 (.A(_09126_),
    .X(net170));
 sg13g2_buf_2 fanout171 (.A(_09047_),
    .X(net171));
 sg13g2_buf_2 fanout172 (.A(_08905_),
    .X(net172));
 sg13g2_buf_2 fanout173 (.A(_08903_),
    .X(net173));
 sg13g2_buf_2 fanout174 (.A(_07932_),
    .X(net174));
 sg13g2_buf_2 fanout175 (.A(_07908_),
    .X(net175));
 sg13g2_buf_2 fanout176 (.A(_07897_),
    .X(net176));
 sg13g2_buf_2 fanout177 (.A(_07880_),
    .X(net177));
 sg13g2_buf_2 fanout178 (.A(_07879_),
    .X(net178));
 sg13g2_buf_2 fanout179 (.A(_07784_),
    .X(net179));
 sg13g2_buf_2 fanout180 (.A(_07767_),
    .X(net180));
 sg13g2_buf_2 fanout181 (.A(_07719_),
    .X(net181));
 sg13g2_buf_2 fanout182 (.A(_07718_),
    .X(net182));
 sg13g2_buf_2 fanout183 (.A(_07694_),
    .X(net183));
 sg13g2_buf_2 fanout184 (.A(_04200_),
    .X(net184));
 sg13g2_buf_2 fanout185 (.A(_04174_),
    .X(net185));
 sg13g2_buf_2 fanout186 (.A(_04154_),
    .X(net186));
 sg13g2_buf_2 fanout187 (.A(_04152_),
    .X(net187));
 sg13g2_buf_2 fanout188 (.A(_04146_),
    .X(net188));
 sg13g2_buf_2 fanout189 (.A(_04132_),
    .X(net189));
 sg13g2_buf_2 fanout190 (.A(_04107_),
    .X(net190));
 sg13g2_buf_2 fanout191 (.A(_03793_),
    .X(net191));
 sg13g2_buf_2 fanout192 (.A(_03696_),
    .X(net192));
 sg13g2_buf_2 fanout193 (.A(_03566_),
    .X(net193));
 sg13g2_buf_2 fanout194 (.A(_03127_),
    .X(net194));
 sg13g2_buf_2 fanout195 (.A(_03028_),
    .X(net195));
 sg13g2_buf_2 fanout196 (.A(_03013_),
    .X(net196));
 sg13g2_buf_2 fanout197 (.A(_11795_),
    .X(net197));
 sg13g2_buf_2 fanout198 (.A(_11449_),
    .X(net198));
 sg13g2_buf_2 fanout199 (.A(_11398_),
    .X(net199));
 sg13g2_buf_2 fanout200 (.A(_10807_),
    .X(net200));
 sg13g2_buf_2 fanout201 (.A(_10486_),
    .X(net201));
 sg13g2_buf_2 fanout202 (.A(_07707_),
    .X(net202));
 sg13g2_buf_2 fanout203 (.A(_04304_),
    .X(net203));
 sg13g2_buf_2 fanout204 (.A(_04245_),
    .X(net204));
 sg13g2_buf_2 fanout205 (.A(_04144_),
    .X(net205));
 sg13g2_buf_2 fanout206 (.A(_04106_),
    .X(net206));
 sg13g2_buf_2 fanout207 (.A(_03889_),
    .X(net207));
 sg13g2_buf_2 fanout208 (.A(_03616_),
    .X(net208));
 sg13g2_buf_2 fanout209 (.A(_03568_),
    .X(net209));
 sg13g2_buf_2 fanout210 (.A(_03165_),
    .X(net210));
 sg13g2_buf_2 fanout211 (.A(_03154_),
    .X(net211));
 sg13g2_buf_2 fanout212 (.A(_03119_),
    .X(net212));
 sg13g2_buf_2 fanout213 (.A(_03033_),
    .X(net213));
 sg13g2_buf_2 fanout214 (.A(_03021_),
    .X(net214));
 sg13g2_buf_2 fanout215 (.A(_11767_),
    .X(net215));
 sg13g2_buf_2 fanout216 (.A(_11674_),
    .X(net216));
 sg13g2_buf_2 fanout217 (.A(_11540_),
    .X(net217));
 sg13g2_buf_2 fanout218 (.A(_11448_),
    .X(net218));
 sg13g2_buf_2 fanout219 (.A(_11428_),
    .X(net219));
 sg13g2_buf_2 fanout220 (.A(_10552_),
    .X(net220));
 sg13g2_buf_2 fanout221 (.A(_10422_),
    .X(net221));
 sg13g2_buf_2 fanout222 (.A(_10295_),
    .X(net222));
 sg13g2_buf_2 fanout223 (.A(_09914_),
    .X(net223));
 sg13g2_buf_2 fanout224 (.A(_09865_),
    .X(net224));
 sg13g2_buf_2 fanout225 (.A(_09027_),
    .X(net225));
 sg13g2_buf_2 fanout226 (.A(_04110_),
    .X(net226));
 sg13g2_buf_2 fanout227 (.A(_03888_),
    .X(net227));
 sg13g2_buf_2 fanout228 (.A(_03245_),
    .X(net228));
 sg13g2_buf_2 fanout229 (.A(_03238_),
    .X(net229));
 sg13g2_buf_2 fanout230 (.A(_03032_),
    .X(net230));
 sg13g2_buf_2 fanout231 (.A(_03014_),
    .X(net231));
 sg13g2_buf_2 fanout232 (.A(_11643_),
    .X(net232));
 sg13g2_buf_2 fanout233 (.A(_11625_),
    .X(net233));
 sg13g2_buf_2 fanout234 (.A(_11619_),
    .X(net234));
 sg13g2_buf_2 fanout235 (.A(_11577_),
    .X(net235));
 sg13g2_buf_2 fanout236 (.A(_11547_),
    .X(net236));
 sg13g2_buf_2 fanout237 (.A(_11539_),
    .X(net237));
 sg13g2_buf_2 fanout238 (.A(_11504_),
    .X(net238));
 sg13g2_buf_2 fanout239 (.A(_11469_),
    .X(net239));
 sg13g2_buf_2 fanout240 (.A(_11447_),
    .X(net240));
 sg13g2_buf_2 fanout241 (.A(_11186_),
    .X(net241));
 sg13g2_buf_2 fanout242 (.A(_10551_),
    .X(net242));
 sg13g2_buf_2 fanout243 (.A(_09913_),
    .X(net243));
 sg13g2_buf_2 fanout244 (.A(_06399_),
    .X(net244));
 sg13g2_buf_2 fanout245 (.A(_06378_),
    .X(net245));
 sg13g2_buf_2 fanout246 (.A(_06348_),
    .X(net246));
 sg13g2_buf_2 fanout247 (.A(_06298_),
    .X(net247));
 sg13g2_buf_2 fanout248 (.A(_06288_),
    .X(net248));
 sg13g2_buf_2 fanout249 (.A(_06245_),
    .X(net249));
 sg13g2_buf_2 fanout250 (.A(_06204_),
    .X(net250));
 sg13g2_buf_2 fanout251 (.A(_06194_),
    .X(net251));
 sg13g2_buf_2 fanout252 (.A(_06183_),
    .X(net252));
 sg13g2_buf_2 fanout253 (.A(_06148_),
    .X(net253));
 sg13g2_buf_2 fanout254 (.A(_06097_),
    .X(net254));
 sg13g2_buf_2 fanout255 (.A(_06085_),
    .X(net255));
 sg13g2_buf_2 fanout256 (.A(_06053_),
    .X(net256));
 sg13g2_buf_4 fanout257 (.X(net257),
    .A(_06044_));
 sg13g2_buf_4 fanout258 (.X(net258),
    .A(_06038_));
 sg13g2_buf_4 fanout259 (.X(net259),
    .A(_06022_));
 sg13g2_buf_4 fanout260 (.X(net260),
    .A(_06006_));
 sg13g2_buf_4 fanout261 (.X(net261),
    .A(_06001_));
 sg13g2_buf_4 fanout262 (.X(net262),
    .A(_05982_));
 sg13g2_buf_4 fanout263 (.X(net263),
    .A(_05963_));
 sg13g2_buf_4 fanout264 (.X(net264),
    .A(_05960_));
 sg13g2_buf_4 fanout265 (.X(net265),
    .A(_05955_));
 sg13g2_buf_4 fanout266 (.X(net266),
    .A(_05937_));
 sg13g2_buf_4 fanout267 (.X(net267),
    .A(_05914_));
 sg13g2_buf_4 fanout268 (.X(net268),
    .A(_05908_));
 sg13g2_buf_4 fanout269 (.X(net269),
    .A(_05887_));
 sg13g2_buf_2 fanout270 (.A(_04573_),
    .X(net270));
 sg13g2_buf_2 fanout271 (.A(_03885_),
    .X(net271));
 sg13g2_buf_2 fanout272 (.A(_03027_),
    .X(net272));
 sg13g2_buf_4 fanout273 (.X(net273),
    .A(_02996_));
 sg13g2_buf_4 fanout274 (.X(net274),
    .A(_02995_));
 sg13g2_buf_2 fanout275 (.A(_11835_),
    .X(net275));
 sg13g2_buf_2 fanout276 (.A(_11589_),
    .X(net276));
 sg13g2_buf_2 fanout277 (.A(_11554_),
    .X(net277));
 sg13g2_buf_2 fanout278 (.A(_11518_),
    .X(net278));
 sg13g2_buf_2 fanout279 (.A(_11078_),
    .X(net279));
 sg13g2_buf_2 fanout280 (.A(_10849_),
    .X(net280));
 sg13g2_buf_2 fanout281 (.A(_10798_),
    .X(net281));
 sg13g2_buf_2 fanout282 (.A(_10767_),
    .X(net282));
 sg13g2_buf_2 fanout283 (.A(_10738_),
    .X(net283));
 sg13g2_buf_2 fanout284 (.A(_10650_),
    .X(net284));
 sg13g2_buf_2 fanout285 (.A(_10618_),
    .X(net285));
 sg13g2_buf_2 fanout286 (.A(_10589_),
    .X(net286));
 sg13g2_buf_2 fanout287 (.A(_09894_),
    .X(net287));
 sg13g2_buf_2 fanout288 (.A(_09451_),
    .X(net288));
 sg13g2_buf_2 fanout289 (.A(_09397_),
    .X(net289));
 sg13g2_buf_2 fanout290 (.A(_09139_),
    .X(net290));
 sg13g2_buf_2 fanout291 (.A(_09122_),
    .X(net291));
 sg13g2_buf_2 fanout292 (.A(_09084_),
    .X(net292));
 sg13g2_buf_2 fanout293 (.A(_08987_),
    .X(net293));
 sg13g2_buf_2 fanout294 (.A(_06665_),
    .X(net294));
 sg13g2_buf_2 fanout295 (.A(_06561_),
    .X(net295));
 sg13g2_buf_2 fanout296 (.A(_06398_),
    .X(net296));
 sg13g2_buf_2 fanout297 (.A(_06389_),
    .X(net297));
 sg13g2_buf_2 fanout298 (.A(_06377_),
    .X(net298));
 sg13g2_buf_2 fanout299 (.A(_06368_),
    .X(net299));
 sg13g2_buf_2 fanout300 (.A(_06358_),
    .X(net300));
 sg13g2_buf_2 fanout301 (.A(_06347_),
    .X(net301));
 sg13g2_buf_2 fanout302 (.A(_06338_),
    .X(net302));
 sg13g2_buf_2 fanout303 (.A(_06328_),
    .X(net303));
 sg13g2_buf_2 fanout304 (.A(_06318_),
    .X(net304));
 sg13g2_buf_2 fanout305 (.A(_06308_),
    .X(net305));
 sg13g2_buf_2 fanout306 (.A(_06297_),
    .X(net306));
 sg13g2_buf_2 fanout307 (.A(_06287_),
    .X(net307));
 sg13g2_buf_2 fanout308 (.A(_06273_),
    .X(net308));
 sg13g2_buf_2 fanout309 (.A(_06262_),
    .X(net309));
 sg13g2_buf_2 fanout310 (.A(_06244_),
    .X(net310));
 sg13g2_buf_2 fanout311 (.A(_06235_),
    .X(net311));
 sg13g2_buf_2 fanout312 (.A(_06224_),
    .X(net312));
 sg13g2_buf_2 fanout313 (.A(_06214_),
    .X(net313));
 sg13g2_buf_2 fanout314 (.A(_06203_),
    .X(net314));
 sg13g2_buf_2 fanout315 (.A(_06193_),
    .X(net315));
 sg13g2_buf_2 fanout316 (.A(_06182_),
    .X(net316));
 sg13g2_buf_2 fanout317 (.A(_06173_),
    .X(net317));
 sg13g2_buf_2 fanout318 (.A(_06159_),
    .X(net318));
 sg13g2_buf_2 fanout319 (.A(_06147_),
    .X(net319));
 sg13g2_buf_2 fanout320 (.A(_06131_),
    .X(net320));
 sg13g2_buf_2 fanout321 (.A(_06119_),
    .X(net321));
 sg13g2_buf_2 fanout322 (.A(_06108_),
    .X(net322));
 sg13g2_buf_2 fanout323 (.A(_06096_),
    .X(net323));
 sg13g2_buf_2 fanout324 (.A(_06084_),
    .X(net324));
 sg13g2_buf_2 fanout325 (.A(_06074_),
    .X(net325));
 sg13g2_buf_2 fanout326 (.A(_06064_),
    .X(net326));
 sg13g2_buf_2 fanout327 (.A(_06052_),
    .X(net327));
 sg13g2_buf_4 fanout328 (.X(net328),
    .A(_06041_));
 sg13g2_buf_4 fanout329 (.X(net329),
    .A(_06033_));
 sg13g2_buf_4 fanout330 (.X(net330),
    .A(_06027_));
 sg13g2_buf_4 fanout331 (.X(net331),
    .A(_06018_));
 sg13g2_buf_4 fanout332 (.X(net332),
    .A(_06015_));
 sg13g2_buf_4 fanout333 (.X(net333),
    .A(_06012_));
 sg13g2_buf_4 fanout334 (.X(net334),
    .A(_06009_));
 sg13g2_buf_4 fanout335 (.X(net335),
    .A(_05993_));
 sg13g2_buf_4 fanout336 (.X(net336),
    .A(_05988_));
 sg13g2_buf_4 fanout337 (.X(net337),
    .A(_05979_));
 sg13g2_buf_4 fanout338 (.X(net338),
    .A(_05970_));
 sg13g2_buf_4 fanout339 (.X(net339),
    .A(_05966_));
 sg13g2_buf_4 fanout340 (.X(net340),
    .A(_05950_));
 sg13g2_buf_4 fanout341 (.X(net341),
    .A(_05942_));
 sg13g2_buf_4 fanout342 (.X(net342),
    .A(_05932_));
 sg13g2_buf_4 fanout343 (.X(net343),
    .A(_05926_));
 sg13g2_buf_4 fanout344 (.X(net344),
    .A(_05919_));
 sg13g2_buf_4 fanout345 (.X(net345),
    .A(_05903_));
 sg13g2_buf_4 fanout346 (.X(net346),
    .A(_05898_));
 sg13g2_buf_2 fanout347 (.A(_04953_),
    .X(net347));
 sg13g2_buf_2 fanout348 (.A(_04921_),
    .X(net348));
 sg13g2_buf_2 fanout349 (.A(_03896_),
    .X(net349));
 sg13g2_buf_2 fanout350 (.A(_03562_),
    .X(net350));
 sg13g2_buf_2 fanout351 (.A(_03560_),
    .X(net351));
 sg13g2_buf_2 fanout352 (.A(_03290_),
    .X(net352));
 sg13g2_buf_2 fanout353 (.A(_03026_),
    .X(net353));
 sg13g2_buf_4 fanout354 (.X(net354),
    .A(_03007_));
 sg13g2_buf_4 fanout355 (.X(net355),
    .A(_03006_));
 sg13g2_buf_4 fanout356 (.X(net356),
    .A(_03005_));
 sg13g2_buf_4 fanout357 (.X(net357),
    .A(_03004_));
 sg13g2_buf_2 fanout358 (.A(_12541_),
    .X(net358));
 sg13g2_buf_2 fanout359 (.A(_11496_),
    .X(net359));
 sg13g2_buf_2 fanout360 (.A(_10851_),
    .X(net360));
 sg13g2_buf_2 fanout361 (.A(_10818_),
    .X(net361));
 sg13g2_buf_2 fanout362 (.A(_10116_),
    .X(net362));
 sg13g2_buf_2 fanout363 (.A(_09857_),
    .X(net363));
 sg13g2_buf_2 fanout364 (.A(_09701_),
    .X(net364));
 sg13g2_buf_2 fanout365 (.A(_09679_),
    .X(net365));
 sg13g2_buf_2 fanout366 (.A(_09545_),
    .X(net366));
 sg13g2_buf_2 fanout367 (.A(_09522_),
    .X(net367));
 sg13g2_buf_2 fanout368 (.A(_09493_),
    .X(net368));
 sg13g2_buf_2 fanout369 (.A(_09142_),
    .X(net369));
 sg13g2_buf_2 fanout370 (.A(_09091_),
    .X(net370));
 sg13g2_buf_2 fanout371 (.A(_08470_),
    .X(net371));
 sg13g2_buf_2 fanout372 (.A(_06666_),
    .X(net372));
 sg13g2_buf_2 fanout373 (.A(_06651_),
    .X(net373));
 sg13g2_buf_2 fanout374 (.A(_06649_),
    .X(net374));
 sg13g2_buf_2 fanout375 (.A(_06648_),
    .X(net375));
 sg13g2_buf_2 fanout376 (.A(_06632_),
    .X(net376));
 sg13g2_buf_2 fanout377 (.A(_06630_),
    .X(net377));
 sg13g2_buf_2 fanout378 (.A(_06629_),
    .X(net378));
 sg13g2_buf_2 fanout379 (.A(_06609_),
    .X(net379));
 sg13g2_buf_2 fanout380 (.A(_06560_),
    .X(net380));
 sg13g2_buf_2 fanout381 (.A(_06498_),
    .X(net381));
 sg13g2_buf_2 fanout382 (.A(_06388_),
    .X(net382));
 sg13g2_buf_2 fanout383 (.A(_06367_),
    .X(net383));
 sg13g2_buf_2 fanout384 (.A(_06357_),
    .X(net384));
 sg13g2_buf_2 fanout385 (.A(_06337_),
    .X(net385));
 sg13g2_buf_2 fanout386 (.A(_06327_),
    .X(net386));
 sg13g2_buf_2 fanout387 (.A(_06317_),
    .X(net387));
 sg13g2_buf_2 fanout388 (.A(_06307_),
    .X(net388));
 sg13g2_buf_2 fanout389 (.A(_06272_),
    .X(net389));
 sg13g2_buf_2 fanout390 (.A(_06261_),
    .X(net390));
 sg13g2_buf_2 fanout391 (.A(_06234_),
    .X(net391));
 sg13g2_buf_2 fanout392 (.A(_06223_),
    .X(net392));
 sg13g2_buf_2 fanout393 (.A(_06213_),
    .X(net393));
 sg13g2_buf_2 fanout394 (.A(_06172_),
    .X(net394));
 sg13g2_buf_2 fanout395 (.A(_06158_),
    .X(net395));
 sg13g2_buf_2 fanout396 (.A(_06130_),
    .X(net396));
 sg13g2_buf_2 fanout397 (.A(_06118_),
    .X(net397));
 sg13g2_buf_2 fanout398 (.A(_06107_),
    .X(net398));
 sg13g2_buf_2 fanout399 (.A(_06073_),
    .X(net399));
 sg13g2_buf_2 fanout400 (.A(_06063_),
    .X(net400));
 sg13g2_buf_2 fanout401 (.A(_06003_),
    .X(net401));
 sg13g2_buf_2 fanout402 (.A(_05952_),
    .X(net402));
 sg13g2_buf_2 fanout403 (.A(_05889_),
    .X(net403));
 sg13g2_buf_2 fanout404 (.A(_05371_),
    .X(net404));
 sg13g2_buf_2 fanout405 (.A(_05153_),
    .X(net405));
 sg13g2_buf_2 fanout406 (.A(_04962_),
    .X(net406));
 sg13g2_buf_2 fanout407 (.A(_04935_),
    .X(net407));
 sg13g2_buf_2 fanout408 (.A(_04909_),
    .X(net408));
 sg13g2_buf_2 fanout409 (.A(_03519_),
    .X(net409));
 sg13g2_buf_2 fanout410 (.A(_03511_),
    .X(net410));
 sg13g2_buf_4 fanout411 (.X(net411),
    .A(_03010_));
 sg13g2_buf_4 fanout412 (.X(net412),
    .A(_03008_));
 sg13g2_buf_4 fanout413 (.X(net413),
    .A(_02999_));
 sg13g2_buf_2 fanout414 (.A(_02997_),
    .X(net414));
 sg13g2_buf_2 fanout415 (.A(_02766_),
    .X(net415));
 sg13g2_buf_2 fanout416 (.A(_12780_),
    .X(net416));
 sg13g2_buf_2 fanout417 (.A(_10115_),
    .X(net417));
 sg13g2_buf_2 fanout418 (.A(_09792_),
    .X(net418));
 sg13g2_buf_2 fanout419 (.A(_09770_),
    .X(net419));
 sg13g2_buf_2 fanout420 (.A(_09723_),
    .X(net420));
 sg13g2_buf_2 fanout421 (.A(_09658_),
    .X(net421));
 sg13g2_buf_2 fanout422 (.A(_09309_),
    .X(net422));
 sg13g2_buf_2 fanout423 (.A(_09066_),
    .X(net423));
 sg13g2_buf_2 fanout424 (.A(_08890_),
    .X(net424));
 sg13g2_buf_2 fanout425 (.A(_08869_),
    .X(net425));
 sg13g2_buf_2 fanout426 (.A(_08848_),
    .X(net426));
 sg13g2_buf_2 fanout427 (.A(_08820_),
    .X(net427));
 sg13g2_buf_2 fanout428 (.A(_08663_),
    .X(net428));
 sg13g2_buf_2 fanout429 (.A(_08603_),
    .X(net429));
 sg13g2_buf_2 fanout430 (.A(_08565_),
    .X(net430));
 sg13g2_buf_2 fanout431 (.A(_08497_),
    .X(net431));
 sg13g2_buf_2 fanout432 (.A(_06724_),
    .X(net432));
 sg13g2_buf_2 fanout433 (.A(_06722_),
    .X(net433));
 sg13g2_buf_2 fanout434 (.A(_06721_),
    .X(net434));
 sg13g2_buf_2 fanout435 (.A(_06686_),
    .X(net435));
 sg13g2_buf_2 fanout436 (.A(_06684_),
    .X(net436));
 sg13g2_buf_2 fanout437 (.A(_06683_),
    .X(net437));
 sg13g2_buf_2 fanout438 (.A(_06610_),
    .X(net438));
 sg13g2_buf_2 fanout439 (.A(_06497_),
    .X(net439));
 sg13g2_buf_2 fanout440 (.A(_06409_),
    .X(net440));
 sg13g2_buf_2 fanout441 (.A(_06408_),
    .X(net441));
 sg13g2_buf_2 fanout442 (.A(_06407_),
    .X(net442));
 sg13g2_buf_2 fanout443 (.A(_06284_),
    .X(net443));
 sg13g2_buf_2 fanout444 (.A(_06170_),
    .X(net444));
 sg13g2_buf_2 fanout445 (.A(_04998_),
    .X(net445));
 sg13g2_buf_2 fanout446 (.A(_04960_),
    .X(net446));
 sg13g2_buf_2 fanout447 (.A(_04955_),
    .X(net447));
 sg13g2_buf_2 fanout448 (.A(_04946_),
    .X(net448));
 sg13g2_buf_2 fanout449 (.A(_04938_),
    .X(net449));
 sg13g2_buf_2 fanout450 (.A(_04926_),
    .X(net450));
 sg13g2_buf_2 fanout451 (.A(_03830_),
    .X(net451));
 sg13g2_buf_4 fanout452 (.X(net452),
    .A(_03513_));
 sg13g2_buf_2 fanout453 (.A(_03510_),
    .X(net453));
 sg13g2_buf_2 fanout454 (.A(_03502_),
    .X(net454));
 sg13g2_buf_4 fanout455 (.X(net455),
    .A(_02990_));
 sg13g2_buf_2 fanout456 (.A(_02886_),
    .X(net456));
 sg13g2_buf_2 fanout457 (.A(_12657_),
    .X(net457));
 sg13g2_buf_2 fanout458 (.A(_12174_),
    .X(net458));
 sg13g2_buf_2 fanout459 (.A(_12074_),
    .X(net459));
 sg13g2_buf_2 fanout460 (.A(_11502_),
    .X(net460));
 sg13g2_buf_2 fanout461 (.A(_11497_),
    .X(net461));
 sg13g2_buf_2 fanout462 (.A(_09308_),
    .X(net462));
 sg13g2_buf_4 fanout463 (.X(net463),
    .A(_09298_));
 sg13g2_buf_2 fanout464 (.A(_08778_),
    .X(net464));
 sg13g2_buf_2 fanout465 (.A(_08758_),
    .X(net465));
 sg13g2_buf_2 fanout466 (.A(_07808_),
    .X(net466));
 sg13g2_buf_2 fanout467 (.A(_07086_),
    .X(net467));
 sg13g2_buf_2 fanout468 (.A(_06743_),
    .X(net468));
 sg13g2_buf_2 fanout469 (.A(_06741_),
    .X(net469));
 sg13g2_buf_2 fanout470 (.A(_06740_),
    .X(net470));
 sg13g2_buf_2 fanout471 (.A(_06705_),
    .X(net471));
 sg13g2_buf_2 fanout472 (.A(_06703_),
    .X(net472));
 sg13g2_buf_2 fanout473 (.A(_06702_),
    .X(net473));
 sg13g2_buf_2 fanout474 (.A(_06283_),
    .X(net474));
 sg13g2_buf_2 fanout475 (.A(_06169_),
    .X(net475));
 sg13g2_buf_2 fanout476 (.A(_06116_),
    .X(net476));
 sg13g2_buf_2 fanout477 (.A(_06061_),
    .X(net477));
 sg13g2_buf_2 fanout478 (.A(_05984_),
    .X(net478));
 sg13g2_buf_2 fanout479 (.A(_05934_),
    .X(net479));
 sg13g2_buf_2 fanout480 (.A(_05916_),
    .X(net480));
 sg13g2_buf_2 fanout481 (.A(_05890_),
    .X(net481));
 sg13g2_buf_2 fanout482 (.A(_05217_),
    .X(net482));
 sg13g2_buf_2 fanout483 (.A(_05184_),
    .X(net483));
 sg13g2_buf_2 fanout484 (.A(_05132_),
    .X(net484));
 sg13g2_buf_2 fanout485 (.A(_05129_),
    .X(net485));
 sg13g2_buf_2 fanout486 (.A(_04914_),
    .X(net486));
 sg13g2_buf_2 fanout487 (.A(_04907_),
    .X(net487));
 sg13g2_buf_2 fanout488 (.A(_03829_),
    .X(net488));
 sg13g2_buf_2 fanout489 (.A(_03551_),
    .X(net489));
 sg13g2_buf_2 fanout490 (.A(_03512_),
    .X(net490));
 sg13g2_buf_4 fanout491 (.X(net491),
    .A(_03509_));
 sg13g2_buf_2 fanout492 (.A(_03508_),
    .X(net492));
 sg13g2_buf_2 fanout493 (.A(_03501_),
    .X(net493));
 sg13g2_buf_2 fanout494 (.A(_03500_),
    .X(net494));
 sg13g2_buf_4 fanout495 (.X(net495),
    .A(_02991_));
 sg13g2_buf_4 fanout496 (.X(net496),
    .A(_02980_));
 sg13g2_buf_4 fanout497 (.X(net497),
    .A(_02978_));
 sg13g2_buf_2 fanout498 (.A(_02699_),
    .X(net498));
 sg13g2_buf_2 fanout499 (.A(_02692_),
    .X(net499));
 sg13g2_buf_2 fanout500 (.A(_12710_),
    .X(net500));
 sg13g2_buf_2 fanout501 (.A(_12418_),
    .X(net501));
 sg13g2_buf_2 fanout502 (.A(_12342_),
    .X(net502));
 sg13g2_buf_2 fanout503 (.A(_12199_),
    .X(net503));
 sg13g2_buf_2 fanout504 (.A(_12162_),
    .X(net504));
 sg13g2_buf_2 fanout505 (.A(_12117_),
    .X(net505));
 sg13g2_buf_2 fanout506 (.A(_12111_),
    .X(net506));
 sg13g2_buf_2 fanout507 (.A(_12105_),
    .X(net507));
 sg13g2_buf_2 fanout508 (.A(_12097_),
    .X(net508));
 sg13g2_buf_2 fanout509 (.A(_12085_),
    .X(net509));
 sg13g2_buf_2 fanout510 (.A(_11501_),
    .X(net510));
 sg13g2_buf_4 fanout511 (.X(net511),
    .A(_11091_));
 sg13g2_buf_2 fanout512 (.A(_10342_),
    .X(net512));
 sg13g2_buf_2 fanout513 (.A(_10339_),
    .X(net513));
 sg13g2_buf_2 fanout514 (.A(_10095_),
    .X(net514));
 sg13g2_buf_2 fanout515 (.A(_09947_),
    .X(net515));
 sg13g2_buf_4 fanout516 (.X(net516),
    .A(_09297_));
 sg13g2_buf_2 fanout517 (.A(_09286_),
    .X(net517));
 sg13g2_buf_4 fanout518 (.X(net518),
    .A(_09031_));
 sg13g2_buf_2 fanout519 (.A(_08799_),
    .X(net519));
 sg13g2_buf_2 fanout520 (.A(_08606_),
    .X(net520));
 sg13g2_buf_2 fanout521 (.A(_08509_),
    .X(net521));
 sg13g2_buf_2 fanout522 (.A(_07616_),
    .X(net522));
 sg13g2_buf_2 fanout523 (.A(_07418_),
    .X(net523));
 sg13g2_buf_2 fanout524 (.A(_07094_),
    .X(net524));
 sg13g2_buf_2 fanout525 (.A(_06275_),
    .X(net525));
 sg13g2_buf_2 fanout526 (.A(_06161_),
    .X(net526));
 sg13g2_buf_2 fanout527 (.A(_05983_),
    .X(net527));
 sg13g2_buf_2 fanout528 (.A(_05933_),
    .X(net528));
 sg13g2_buf_2 fanout529 (.A(_05172_),
    .X(net529));
 sg13g2_buf_2 fanout530 (.A(_05134_),
    .X(net530));
 sg13g2_buf_2 fanout531 (.A(_05128_),
    .X(net531));
 sg13g2_buf_2 fanout532 (.A(_04877_),
    .X(net532));
 sg13g2_buf_2 fanout533 (.A(_04842_),
    .X(net533));
 sg13g2_buf_2 fanout534 (.A(_04797_),
    .X(net534));
 sg13g2_buf_2 fanout535 (.A(_04796_),
    .X(net535));
 sg13g2_buf_2 fanout536 (.A(_04794_),
    .X(net536));
 sg13g2_buf_2 fanout537 (.A(_04787_),
    .X(net537));
 sg13g2_buf_2 fanout538 (.A(_04783_),
    .X(net538));
 sg13g2_buf_2 fanout539 (.A(_03860_),
    .X(net539));
 sg13g2_buf_2 fanout540 (.A(_03835_),
    .X(net540));
 sg13g2_buf_2 fanout541 (.A(_03831_),
    .X(net541));
 sg13g2_buf_2 fanout542 (.A(_03550_),
    .X(net542));
 sg13g2_buf_4 fanout543 (.X(net543),
    .A(_03549_));
 sg13g2_buf_4 fanout544 (.X(net544),
    .A(_03545_));
 sg13g2_buf_4 fanout545 (.X(net545),
    .A(_03537_));
 sg13g2_buf_4 fanout546 (.X(net546),
    .A(_03533_));
 sg13g2_buf_4 fanout547 (.X(net547),
    .A(_03529_));
 sg13g2_buf_4 fanout548 (.X(net548),
    .A(_03524_));
 sg13g2_buf_4 fanout549 (.X(net549),
    .A(_03517_));
 sg13g2_buf_4 fanout550 (.X(net550),
    .A(_03507_));
 sg13g2_buf_2 fanout551 (.A(_03504_),
    .X(net551));
 sg13g2_buf_2 fanout552 (.A(_03499_),
    .X(net552));
 sg13g2_buf_4 fanout553 (.X(net553),
    .A(_03497_));
 sg13g2_buf_4 fanout554 (.X(net554),
    .A(_02958_));
 sg13g2_buf_2 fanout555 (.A(_02956_),
    .X(net555));
 sg13g2_buf_2 fanout556 (.A(_02691_),
    .X(net556));
 sg13g2_buf_2 fanout557 (.A(_12703_),
    .X(net557));
 sg13g2_buf_4 fanout558 (.X(net558),
    .A(_12475_));
 sg13g2_buf_2 fanout559 (.A(_12470_),
    .X(net559));
 sg13g2_buf_2 fanout560 (.A(_12341_),
    .X(net560));
 sg13g2_buf_2 fanout561 (.A(_12287_),
    .X(net561));
 sg13g2_buf_2 fanout562 (.A(_12198_),
    .X(net562));
 sg13g2_buf_2 fanout563 (.A(_11977_),
    .X(net563));
 sg13g2_buf_2 fanout564 (.A(_11507_),
    .X(net564));
 sg13g2_buf_2 fanout565 (.A(_11500_),
    .X(net565));
 sg13g2_buf_2 fanout566 (.A(_11402_),
    .X(net566));
 sg13g2_buf_2 fanout567 (.A(_10957_),
    .X(net567));
 sg13g2_buf_2 fanout568 (.A(_10893_),
    .X(net568));
 sg13g2_buf_2 fanout569 (.A(_10286_),
    .X(net569));
 sg13g2_buf_2 fanout570 (.A(_10281_),
    .X(net570));
 sg13g2_buf_2 fanout571 (.A(_10245_),
    .X(net571));
 sg13g2_buf_2 fanout572 (.A(_10229_),
    .X(net572));
 sg13g2_buf_2 fanout573 (.A(_10094_),
    .X(net573));
 sg13g2_buf_2 fanout574 (.A(_10087_),
    .X(net574));
 sg13g2_buf_2 fanout575 (.A(_10044_),
    .X(net575));
 sg13g2_buf_2 fanout576 (.A(_09946_),
    .X(net576));
 sg13g2_buf_2 fanout577 (.A(_09448_),
    .X(net577));
 sg13g2_buf_4 fanout578 (.X(net578),
    .A(_09296_));
 sg13g2_buf_2 fanout579 (.A(_09010_),
    .X(net579));
 sg13g2_buf_2 fanout580 (.A(_08959_),
    .X(net580));
 sg13g2_buf_2 fanout581 (.A(_08800_),
    .X(net581));
 sg13g2_buf_2 fanout582 (.A(_08605_),
    .X(net582));
 sg13g2_buf_2 fanout583 (.A(_08531_),
    .X(net583));
 sg13g2_buf_2 fanout584 (.A(_08508_),
    .X(net584));
 sg13g2_buf_2 fanout585 (.A(_06276_),
    .X(net585));
 sg13g2_buf_2 fanout586 (.A(_06270_),
    .X(net586));
 sg13g2_buf_2 fanout587 (.A(_06162_),
    .X(net587));
 sg13g2_buf_2 fanout588 (.A(_06156_),
    .X(net588));
 sg13g2_buf_2 fanout589 (.A(_05994_),
    .X(net589));
 sg13g2_buf_2 fanout590 (.A(_05943_),
    .X(net590));
 sg13g2_buf_2 fanout591 (.A(_05863_),
    .X(net591));
 sg13g2_buf_2 fanout592 (.A(_05162_),
    .X(net592));
 sg13g2_buf_2 fanout593 (.A(_04994_),
    .X(net593));
 sg13g2_buf_2 fanout594 (.A(_04859_),
    .X(net594));
 sg13g2_buf_2 fanout595 (.A(_04858_),
    .X(net595));
 sg13g2_buf_2 fanout596 (.A(_04793_),
    .X(net596));
 sg13g2_buf_4 fanout597 (.X(net597),
    .A(_04781_));
 sg13g2_buf_2 fanout598 (.A(_03859_),
    .X(net598));
 sg13g2_buf_2 fanout599 (.A(_03839_),
    .X(net599));
 sg13g2_buf_2 fanout600 (.A(_03834_),
    .X(net600));
 sg13g2_buf_2 fanout601 (.A(_03832_),
    .X(net601));
 sg13g2_buf_2 fanout602 (.A(_03827_),
    .X(net602));
 sg13g2_buf_2 fanout603 (.A(_03826_),
    .X(net603));
 sg13g2_buf_4 fanout604 (.X(net604),
    .A(_03823_));
 sg13g2_buf_2 fanout605 (.A(_03503_),
    .X(net605));
 sg13g2_buf_4 fanout606 (.X(net606),
    .A(_03496_));
 sg13g2_buf_2 fanout607 (.A(_02977_),
    .X(net607));
 sg13g2_buf_2 fanout608 (.A(_12702_),
    .X(net608));
 sg13g2_buf_2 fanout609 (.A(_12469_),
    .X(net609));
 sg13g2_buf_2 fanout610 (.A(_12340_),
    .X(net610));
 sg13g2_buf_2 fanout611 (.A(_12158_),
    .X(net611));
 sg13g2_buf_2 fanout612 (.A(_12124_),
    .X(net612));
 sg13g2_buf_2 fanout613 (.A(_11976_),
    .X(net613));
 sg13g2_buf_2 fanout614 (.A(_11913_),
    .X(net614));
 sg13g2_buf_2 fanout615 (.A(_11499_),
    .X(net615));
 sg13g2_buf_2 fanout616 (.A(_10801_),
    .X(net616));
 sg13g2_buf_2 fanout617 (.A(_10341_),
    .X(net617));
 sg13g2_buf_2 fanout618 (.A(_10308_),
    .X(net618));
 sg13g2_buf_2 fanout619 (.A(_10280_),
    .X(net619));
 sg13g2_buf_2 fanout620 (.A(_10244_),
    .X(net620));
 sg13g2_buf_2 fanout621 (.A(_10086_),
    .X(net621));
 sg13g2_buf_2 fanout622 (.A(_10042_),
    .X(net622));
 sg13g2_buf_2 fanout623 (.A(_09945_),
    .X(net623));
 sg13g2_buf_2 fanout624 (.A(_09843_),
    .X(net624));
 sg13g2_buf_2 fanout625 (.A(_09705_),
    .X(net625));
 sg13g2_buf_4 fanout626 (.X(net626),
    .A(_09476_));
 sg13g2_buf_2 fanout627 (.A(_09419_),
    .X(net627));
 sg13g2_buf_2 fanout628 (.A(_09408_),
    .X(net628));
 sg13g2_buf_4 fanout629 (.X(net629),
    .A(_09388_));
 sg13g2_buf_4 fanout630 (.X(net630),
    .A(_09382_));
 sg13g2_buf_2 fanout631 (.A(_09369_),
    .X(net631));
 sg13g2_buf_4 fanout632 (.X(net632),
    .A(_09295_));
 sg13g2_buf_4 fanout633 (.X(net633),
    .A(_09234_));
 sg13g2_buf_2 fanout634 (.A(_09159_),
    .X(net634));
 sg13g2_buf_4 fanout635 (.X(net635),
    .A(_09037_));
 sg13g2_buf_4 fanout636 (.X(net636),
    .A(_09035_));
 sg13g2_buf_2 fanout637 (.A(_08958_),
    .X(net637));
 sg13g2_buf_2 fanout638 (.A(_08642_),
    .X(net638));
 sg13g2_buf_2 fanout639 (.A(_08637_),
    .X(net639));
 sg13g2_buf_2 fanout640 (.A(_08604_),
    .X(net640));
 sg13g2_buf_2 fanout641 (.A(_08530_),
    .X(net641));
 sg13g2_buf_2 fanout642 (.A(_08523_),
    .X(net642));
 sg13g2_buf_2 fanout643 (.A(_08514_),
    .X(net643));
 sg13g2_buf_2 fanout644 (.A(_08507_),
    .X(net644));
 sg13g2_buf_2 fanout645 (.A(_08180_),
    .X(net645));
 sg13g2_buf_2 fanout646 (.A(_08059_),
    .X(net646));
 sg13g2_buf_2 fanout647 (.A(_07981_),
    .X(net647));
 sg13g2_buf_2 fanout648 (.A(_07935_),
    .X(net648));
 sg13g2_buf_2 fanout649 (.A(_07911_),
    .X(net649));
 sg13g2_buf_2 fanout650 (.A(_07883_),
    .X(net650));
 sg13g2_buf_2 fanout651 (.A(_07851_),
    .X(net651));
 sg13g2_buf_2 fanout652 (.A(_07816_),
    .X(net652));
 sg13g2_buf_2 fanout653 (.A(_07756_),
    .X(net653));
 sg13g2_buf_2 fanout654 (.A(_07678_),
    .X(net654));
 sg13g2_buf_2 fanout655 (.A(_07104_),
    .X(net655));
 sg13g2_buf_2 fanout656 (.A(_06885_),
    .X(net656));
 sg13g2_buf_2 fanout657 (.A(_05971_),
    .X(net657));
 sg13g2_buf_2 fanout658 (.A(_05920_),
    .X(net658));
 sg13g2_buf_2 fanout659 (.A(_05892_),
    .X(net659));
 sg13g2_buf_2 fanout660 (.A(_05827_),
    .X(net660));
 sg13g2_buf_2 fanout661 (.A(_05161_),
    .X(net661));
 sg13g2_buf_2 fanout662 (.A(_04881_),
    .X(net662));
 sg13g2_buf_2 fanout663 (.A(_04857_),
    .X(net663));
 sg13g2_buf_2 fanout664 (.A(_04837_),
    .X(net664));
 sg13g2_buf_2 fanout665 (.A(_03950_),
    .X(net665));
 sg13g2_buf_2 fanout666 (.A(_03838_),
    .X(net666));
 sg13g2_buf_2 fanout667 (.A(_03540_),
    .X(net667));
 sg13g2_buf_2 fanout668 (.A(_02976_),
    .X(net668));
 sg13g2_buf_2 fanout669 (.A(_12348_),
    .X(net669));
 sg13g2_buf_2 fanout670 (.A(_12207_),
    .X(net670));
 sg13g2_buf_2 fanout671 (.A(_12070_),
    .X(net671));
 sg13g2_buf_2 fanout672 (.A(_12008_),
    .X(net672));
 sg13g2_buf_2 fanout673 (.A(_11975_),
    .X(net673));
 sg13g2_buf_2 fanout674 (.A(_11406_),
    .X(net674));
 sg13g2_buf_2 fanout675 (.A(_11098_),
    .X(net675));
 sg13g2_buf_2 fanout676 (.A(_10987_),
    .X(net676));
 sg13g2_buf_2 fanout677 (.A(_10903_),
    .X(net677));
 sg13g2_buf_2 fanout678 (.A(_10307_),
    .X(net678));
 sg13g2_buf_2 fanout679 (.A(_10279_),
    .X(net679));
 sg13g2_buf_2 fanout680 (.A(_10260_),
    .X(net680));
 sg13g2_buf_2 fanout681 (.A(_10253_),
    .X(net681));
 sg13g2_buf_2 fanout682 (.A(_10243_),
    .X(net682));
 sg13g2_buf_2 fanout683 (.A(_10234_),
    .X(net683));
 sg13g2_buf_2 fanout684 (.A(_10092_),
    .X(net684));
 sg13g2_buf_2 fanout685 (.A(_10041_),
    .X(net685));
 sg13g2_buf_2 fanout686 (.A(_09944_),
    .X(net686));
 sg13g2_buf_2 fanout687 (.A(_09853_),
    .X(net687));
 sg13g2_buf_2 fanout688 (.A(_09643_),
    .X(net688));
 sg13g2_buf_2 fanout689 (.A(_09560_),
    .X(net689));
 sg13g2_buf_4 fanout690 (.X(net690),
    .A(_09487_));
 sg13g2_buf_4 fanout691 (.X(net691),
    .A(_09478_));
 sg13g2_buf_4 fanout692 (.X(net692),
    .A(_09473_));
 sg13g2_buf_2 fanout693 (.A(_09468_),
    .X(net693));
 sg13g2_buf_2 fanout694 (.A(_09428_),
    .X(net694));
 sg13g2_buf_8 fanout695 (.A(_09391_),
    .X(net695));
 sg13g2_buf_2 fanout696 (.A(_09387_),
    .X(net696));
 sg13g2_buf_8 fanout697 (.A(_09385_),
    .X(net697));
 sg13g2_buf_4 fanout698 (.X(net698),
    .A(_09381_));
 sg13g2_buf_4 fanout699 (.X(net699),
    .A(_09375_));
 sg13g2_buf_4 fanout700 (.X(net700),
    .A(_09368_));
 sg13g2_buf_4 fanout701 (.X(net701),
    .A(_09366_));
 sg13g2_buf_2 fanout702 (.A(_09363_),
    .X(net702));
 sg13g2_buf_2 fanout703 (.A(_09354_),
    .X(net703));
 sg13g2_buf_2 fanout704 (.A(_09331_),
    .X(net704));
 sg13g2_buf_2 fanout705 (.A(_09323_),
    .X(net705));
 sg13g2_buf_2 fanout706 (.A(_09294_),
    .X(net706));
 sg13g2_buf_4 fanout707 (.X(net707),
    .A(_09233_));
 sg13g2_buf_2 fanout708 (.A(_09158_),
    .X(net708));
 sg13g2_buf_4 fanout709 (.X(net709),
    .A(_08835_));
 sg13g2_buf_4 fanout710 (.X(net710),
    .A(_08826_));
 sg13g2_buf_4 fanout711 (.X(net711),
    .A(_08656_));
 sg13g2_buf_2 fanout712 (.A(_08641_),
    .X(net712));
 sg13g2_buf_2 fanout713 (.A(_08636_),
    .X(net713));
 sg13g2_buf_4 fanout714 (.X(net714),
    .A(_08622_));
 sg13g2_buf_2 fanout715 (.A(_08614_),
    .X(net715));
 sg13g2_buf_4 fanout716 (.X(net716),
    .A(_08611_));
 sg13g2_buf_4 fanout717 (.X(net717),
    .A(_08591_));
 sg13g2_buf_4 fanout718 (.X(net718),
    .A(_08587_));
 sg13g2_buf_2 fanout719 (.A(_08574_),
    .X(net719));
 sg13g2_buf_2 fanout720 (.A(_08569_),
    .X(net720));
 sg13g2_buf_2 fanout721 (.A(_08536_),
    .X(net721));
 sg13g2_buf_2 fanout722 (.A(_08529_),
    .X(net722));
 sg13g2_buf_2 fanout723 (.A(_08522_),
    .X(net723));
 sg13g2_buf_2 fanout724 (.A(_08518_),
    .X(net724));
 sg13g2_buf_2 fanout725 (.A(_08513_),
    .X(net725));
 sg13g2_buf_4 fanout726 (.X(net726),
    .A(_08474_));
 sg13g2_buf_2 fanout727 (.A(_06899_),
    .X(net727));
 sg13g2_buf_2 fanout728 (.A(_06898_),
    .X(net728));
 sg13g2_buf_2 fanout729 (.A(_06257_),
    .X(net729));
 sg13g2_buf_2 fanout730 (.A(_06255_),
    .X(net730));
 sg13g2_buf_2 fanout731 (.A(_06251_),
    .X(net731));
 sg13g2_buf_2 fanout732 (.A(_06250_),
    .X(net732));
 sg13g2_buf_2 fanout733 (.A(_06248_),
    .X(net733));
 sg13g2_buf_2 fanout734 (.A(_06143_),
    .X(net734));
 sg13g2_buf_2 fanout735 (.A(_06141_),
    .X(net735));
 sg13g2_buf_2 fanout736 (.A(_06137_),
    .X(net736));
 sg13g2_buf_2 fanout737 (.A(_06136_),
    .X(net737));
 sg13g2_buf_2 fanout738 (.A(_06134_),
    .X(net738));
 sg13g2_buf_2 fanout739 (.A(_06002_),
    .X(net739));
 sg13g2_buf_2 fanout740 (.A(_05951_),
    .X(net740));
 sg13g2_buf_2 fanout741 (.A(_05888_),
    .X(net741));
 sg13g2_buf_2 fanout742 (.A(_04880_),
    .X(net742));
 sg13g2_buf_2 fanout743 (.A(_04784_),
    .X(net743));
 sg13g2_buf_2 fanout744 (.A(_04115_),
    .X(net744));
 sg13g2_buf_4 fanout745 (.X(net745),
    .A(_03539_));
 sg13g2_buf_2 fanout746 (.A(_03506_),
    .X(net746));
 sg13g2_buf_2 fanout747 (.A(_03009_),
    .X(net747));
 sg13g2_buf_2 fanout748 (.A(_02979_),
    .X(net748));
 sg13g2_buf_2 fanout749 (.A(_02975_),
    .X(net749));
 sg13g2_buf_2 fanout750 (.A(_02971_),
    .X(net750));
 sg13g2_buf_2 fanout751 (.A(_02969_),
    .X(net751));
 sg13g2_buf_2 fanout752 (.A(_02963_),
    .X(net752));
 sg13g2_buf_2 fanout753 (.A(_02961_),
    .X(net753));
 sg13g2_buf_2 fanout754 (.A(_02955_),
    .X(net754));
 sg13g2_buf_2 fanout755 (.A(_12151_),
    .X(net755));
 sg13g2_buf_2 fanout756 (.A(_12146_),
    .X(net756));
 sg13g2_buf_2 fanout757 (.A(_12138_),
    .X(net757));
 sg13g2_buf_2 fanout758 (.A(_11935_),
    .X(net758));
 sg13g2_buf_2 fanout759 (.A(_10993_),
    .X(net759));
 sg13g2_buf_2 fanout760 (.A(_10986_),
    .X(net760));
 sg13g2_buf_2 fanout761 (.A(_10983_),
    .X(net761));
 sg13g2_buf_2 fanout762 (.A(_10965_),
    .X(net762));
 sg13g2_buf_2 fanout763 (.A(_10962_),
    .X(net763));
 sg13g2_buf_2 fanout764 (.A(_10959_),
    .X(net764));
 sg13g2_buf_2 fanout765 (.A(_10945_),
    .X(net765));
 sg13g2_buf_2 fanout766 (.A(_10933_),
    .X(net766));
 sg13g2_buf_2 fanout767 (.A(_10917_),
    .X(net767));
 sg13g2_buf_2 fanout768 (.A(_10911_),
    .X(net768));
 sg13g2_buf_2 fanout769 (.A(_10902_),
    .X(net769));
 sg13g2_buf_2 fanout770 (.A(_10424_),
    .X(net770));
 sg13g2_buf_2 fanout771 (.A(_10362_),
    .X(net771));
 sg13g2_buf_2 fanout772 (.A(_10352_),
    .X(net772));
 sg13g2_buf_2 fanout773 (.A(_10306_),
    .X(net773));
 sg13g2_buf_2 fanout774 (.A(_10278_),
    .X(net774));
 sg13g2_buf_2 fanout775 (.A(_10272_),
    .X(net775));
 sg13g2_buf_2 fanout776 (.A(_10252_),
    .X(net776));
 sg13g2_buf_2 fanout777 (.A(_10248_),
    .X(net777));
 sg13g2_buf_2 fanout778 (.A(_10242_),
    .X(net778));
 sg13g2_buf_2 fanout779 (.A(_10232_),
    .X(net779));
 sg13g2_buf_2 fanout780 (.A(_10040_),
    .X(net780));
 sg13g2_buf_2 fanout781 (.A(_09943_),
    .X(net781));
 sg13g2_buf_2 fanout782 (.A(_09876_),
    .X(net782));
 sg13g2_buf_2 fanout783 (.A(_09810_),
    .X(net783));
 sg13g2_buf_8 fanout784 (.A(_09644_),
    .X(net784));
 sg13g2_buf_2 fanout785 (.A(_09547_),
    .X(net785));
 sg13g2_buf_4 fanout786 (.X(net786),
    .A(_09482_));
 sg13g2_buf_8 fanout787 (.A(_09480_),
    .X(net787));
 sg13g2_buf_8 fanout788 (.A(_09475_),
    .X(net788));
 sg13g2_buf_8 fanout789 (.A(_09472_),
    .X(net789));
 sg13g2_buf_2 fanout790 (.A(_09462_),
    .X(net790));
 sg13g2_buf_2 fanout791 (.A(_09456_),
    .X(net791));
 sg13g2_buf_2 fanout792 (.A(_09421_),
    .X(net792));
 sg13g2_buf_8 fanout793 (.A(_09384_),
    .X(net793));
 sg13g2_buf_8 fanout794 (.A(_09380_),
    .X(net794));
 sg13g2_buf_2 fanout795 (.A(_09378_),
    .X(net795));
 sg13g2_buf_4 fanout796 (.X(net796),
    .A(_09376_));
 sg13g2_buf_4 fanout797 (.X(net797),
    .A(_09374_));
 sg13g2_buf_8 fanout798 (.A(_09365_),
    .X(net798));
 sg13g2_buf_2 fanout799 (.A(_09351_),
    .X(net799));
 sg13g2_buf_2 fanout800 (.A(_09318_),
    .X(net800));
 sg13g2_buf_2 fanout801 (.A(_09293_),
    .X(net801));
 sg13g2_buf_2 fanout802 (.A(_09232_),
    .X(net802));
 sg13g2_buf_2 fanout803 (.A(_09157_),
    .X(net803));
 sg13g2_buf_2 fanout804 (.A(_09009_),
    .X(net804));
 sg13g2_buf_4 fanout805 (.X(net805),
    .A(_08950_));
 sg13g2_buf_2 fanout806 (.A(_08948_),
    .X(net806));
 sg13g2_buf_8 fanout807 (.A(_08834_),
    .X(net807));
 sg13g2_buf_4 fanout808 (.X(net808),
    .A(_08824_));
 sg13g2_buf_4 fanout809 (.X(net809),
    .A(_08745_));
 sg13g2_buf_8 fanout810 (.A(_08655_),
    .X(net810));
 sg13g2_buf_8 fanout811 (.A(_08621_),
    .X(net811));
 sg13g2_buf_2 fanout812 (.A(_08613_),
    .X(net812));
 sg13g2_buf_4 fanout813 (.X(net813),
    .A(_08610_));
 sg13g2_buf_4 fanout814 (.X(net814),
    .A(_08594_));
 sg13g2_buf_2 fanout815 (.A(_08586_),
    .X(net815));
 sg13g2_buf_8 fanout816 (.A(_08585_),
    .X(net816));
 sg13g2_buf_2 fanout817 (.A(_08575_),
    .X(net817));
 sg13g2_buf_4 fanout818 (.X(net818),
    .A(_08550_));
 sg13g2_buf_4 fanout819 (.X(net819),
    .A(_08542_));
 sg13g2_buf_2 fanout820 (.A(_08539_),
    .X(net820));
 sg13g2_buf_2 fanout821 (.A(_08535_),
    .X(net821));
 sg13g2_buf_2 fanout822 (.A(_08517_),
    .X(net822));
 sg13g2_buf_4 fanout823 (.X(net823),
    .A(_08488_));
 sg13g2_buf_4 fanout824 (.X(net824),
    .A(_08478_));
 sg13g2_buf_4 fanout825 (.X(net825),
    .A(_08473_));
 sg13g2_buf_4 fanout826 (.X(net826),
    .A(_08372_));
 sg13g2_buf_2 fanout827 (.A(_07392_),
    .X(net827));
 sg13g2_buf_2 fanout828 (.A(_07236_),
    .X(net828));
 sg13g2_buf_2 fanout829 (.A(_06897_),
    .X(net829));
 sg13g2_buf_2 fanout830 (.A(_06557_),
    .X(net830));
 sg13g2_buf_2 fanout831 (.A(_06555_),
    .X(net831));
 sg13g2_buf_2 fanout832 (.A(_06553_),
    .X(net832));
 sg13g2_buf_2 fanout833 (.A(_06543_),
    .X(net833));
 sg13g2_buf_2 fanout834 (.A(_06542_),
    .X(net834));
 sg13g2_buf_2 fanout835 (.A(_06540_),
    .X(net835));
 sg13g2_buf_2 fanout836 (.A(_06523_),
    .X(net836));
 sg13g2_buf_2 fanout837 (.A(_06519_),
    .X(net837));
 sg13g2_buf_2 fanout838 (.A(_06518_),
    .X(net838));
 sg13g2_buf_2 fanout839 (.A(_06515_),
    .X(net839));
 sg13g2_buf_2 fanout840 (.A(_06510_),
    .X(net840));
 sg13g2_buf_2 fanout841 (.A(_06505_),
    .X(net841));
 sg13g2_buf_2 fanout842 (.A(_06484_),
    .X(net842));
 sg13g2_buf_2 fanout843 (.A(_06472_),
    .X(net843));
 sg13g2_buf_2 fanout844 (.A(_06459_),
    .X(net844));
 sg13g2_buf_2 fanout845 (.A(_06426_),
    .X(net845));
 sg13g2_buf_2 fanout846 (.A(_06259_),
    .X(net846));
 sg13g2_buf_2 fanout847 (.A(_06253_),
    .X(net847));
 sg13g2_buf_2 fanout848 (.A(_06145_),
    .X(net848));
 sg13g2_buf_2 fanout849 (.A(_06139_),
    .X(net849));
 sg13g2_buf_2 fanout850 (.A(_05995_),
    .X(net850));
 sg13g2_buf_2 fanout851 (.A(_05944_),
    .X(net851));
 sg13g2_buf_2 fanout852 (.A(_05870_),
    .X(net852));
 sg13g2_buf_2 fanout853 (.A(_05807_),
    .X(net853));
 sg13g2_buf_2 fanout854 (.A(_05781_),
    .X(net854));
 sg13g2_buf_2 fanout855 (.A(_04834_),
    .X(net855));
 sg13g2_buf_2 fanout856 (.A(_04141_),
    .X(net856));
 sg13g2_buf_2 fanout857 (.A(_03542_),
    .X(net857));
 sg13g2_buf_4 fanout858 (.X(net858),
    .A(_03538_));
 sg13g2_buf_2 fanout859 (.A(_03534_),
    .X(net859));
 sg13g2_buf_2 fanout860 (.A(_03505_),
    .X(net860));
 sg13g2_buf_2 fanout861 (.A(_03490_),
    .X(net861));
 sg13g2_buf_2 fanout862 (.A(_03011_),
    .X(net862));
 sg13g2_buf_2 fanout863 (.A(_02989_),
    .X(net863));
 sg13g2_buf_2 fanout864 (.A(_02988_),
    .X(net864));
 sg13g2_buf_2 fanout865 (.A(_02986_),
    .X(net865));
 sg13g2_buf_2 fanout866 (.A(_02984_),
    .X(net866));
 sg13g2_buf_2 fanout867 (.A(_02982_),
    .X(net867));
 sg13g2_buf_2 fanout868 (.A(_02974_),
    .X(net868));
 sg13g2_buf_2 fanout869 (.A(_02968_),
    .X(net869));
 sg13g2_buf_2 fanout870 (.A(_02965_),
    .X(net870));
 sg13g2_buf_2 fanout871 (.A(_02962_),
    .X(net871));
 sg13g2_buf_2 fanout872 (.A(_02960_),
    .X(net872));
 sg13g2_buf_2 fanout873 (.A(_02954_),
    .X(net873));
 sg13g2_buf_2 fanout874 (.A(_02704_),
    .X(net874));
 sg13g2_buf_2 fanout875 (.A(_12769_),
    .X(net875));
 sg13g2_buf_2 fanout876 (.A(_12766_),
    .X(net876));
 sg13g2_buf_2 fanout877 (.A(_12761_),
    .X(net877));
 sg13g2_buf_2 fanout878 (.A(_12441_),
    .X(net878));
 sg13g2_buf_2 fanout879 (.A(_12400_),
    .X(net879));
 sg13g2_buf_2 fanout880 (.A(_12212_),
    .X(net880));
 sg13g2_buf_2 fanout881 (.A(_12150_),
    .X(net881));
 sg13g2_buf_2 fanout882 (.A(_12145_),
    .X(net882));
 sg13g2_buf_2 fanout883 (.A(_12137_),
    .X(net883));
 sg13g2_buf_2 fanout884 (.A(_12132_),
    .X(net884));
 sg13g2_buf_2 fanout885 (.A(_12130_),
    .X(net885));
 sg13g2_buf_2 fanout886 (.A(_12000_),
    .X(net886));
 sg13g2_buf_2 fanout887 (.A(_11994_),
    .X(net887));
 sg13g2_buf_2 fanout888 (.A(_11974_),
    .X(net888));
 sg13g2_buf_2 fanout889 (.A(_11225_),
    .X(net889));
 sg13g2_buf_2 fanout890 (.A(_11053_),
    .X(net890));
 sg13g2_buf_2 fanout891 (.A(_11001_),
    .X(net891));
 sg13g2_buf_2 fanout892 (.A(_10988_),
    .X(net892));
 sg13g2_buf_2 fanout893 (.A(_10970_),
    .X(net893));
 sg13g2_buf_2 fanout894 (.A(_10961_),
    .X(net894));
 sg13g2_buf_2 fanout895 (.A(_10940_),
    .X(net895));
 sg13g2_buf_2 fanout896 (.A(_10920_),
    .X(net896));
 sg13g2_buf_2 fanout897 (.A(_10916_),
    .X(net897));
 sg13g2_buf_2 fanout898 (.A(_10905_),
    .X(net898));
 sg13g2_buf_2 fanout899 (.A(_10901_),
    .X(net899));
 sg13g2_buf_2 fanout900 (.A(_10351_),
    .X(net900));
 sg13g2_buf_2 fanout901 (.A(_10298_),
    .X(net901));
 sg13g2_buf_2 fanout902 (.A(_10291_),
    .X(net902));
 sg13g2_buf_2 fanout903 (.A(_10277_),
    .X(net903));
 sg13g2_buf_2 fanout904 (.A(_10251_),
    .X(net904));
 sg13g2_buf_2 fanout905 (.A(_10241_),
    .X(net905));
 sg13g2_buf_2 fanout906 (.A(_10231_),
    .X(net906));
 sg13g2_buf_2 fanout907 (.A(_10225_),
    .X(net907));
 sg13g2_buf_2 fanout908 (.A(_10223_),
    .X(net908));
 sg13g2_buf_2 fanout909 (.A(_10206_),
    .X(net909));
 sg13g2_buf_2 fanout910 (.A(_10107_),
    .X(net910));
 sg13g2_buf_2 fanout911 (.A(_10099_),
    .X(net911));
 sg13g2_buf_2 fanout912 (.A(_10039_),
    .X(net912));
 sg13g2_buf_2 fanout913 (.A(_10034_),
    .X(net913));
 sg13g2_buf_4 fanout914 (.X(net914),
    .A(_09942_));
 sg13g2_buf_2 fanout915 (.A(_09498_),
    .X(net915));
 sg13g2_buf_2 fanout916 (.A(_09494_),
    .X(net916));
 sg13g2_buf_2 fanout917 (.A(_09431_),
    .X(net917));
 sg13g2_buf_2 fanout918 (.A(_09416_),
    .X(net918));
 sg13g2_buf_2 fanout919 (.A(_09411_),
    .X(net919));
 sg13g2_buf_2 fanout920 (.A(_09405_),
    .X(net920));
 sg13g2_buf_2 fanout921 (.A(_09402_),
    .X(net921));
 sg13g2_buf_4 fanout922 (.X(net922),
    .A(_09379_));
 sg13g2_buf_2 fanout923 (.A(_09317_),
    .X(net923));
 sg13g2_buf_2 fanout924 (.A(_09292_),
    .X(net924));
 sg13g2_buf_2 fanout925 (.A(_09290_),
    .X(net925));
 sg13g2_buf_2 fanout926 (.A(_09241_),
    .X(net926));
 sg13g2_buf_2 fanout927 (.A(_09231_),
    .X(net927));
 sg13g2_buf_2 fanout928 (.A(_09156_),
    .X(net928));
 sg13g2_buf_2 fanout929 (.A(_08968_),
    .X(net929));
 sg13g2_buf_8 fanout930 (.A(_08744_),
    .X(net930));
 sg13g2_buf_4 fanout931 (.X(net931),
    .A(_08625_));
 sg13g2_buf_4 fanout932 (.X(net932),
    .A(_08609_));
 sg13g2_buf_8 fanout933 (.A(_08590_),
    .X(net933));
 sg13g2_buf_4 fanout934 (.X(net934),
    .A(_08584_));
 sg13g2_buf_2 fanout935 (.A(_08544_),
    .X(net935));
 sg13g2_buf_2 fanout936 (.A(_08541_),
    .X(net936));
 sg13g2_buf_2 fanout937 (.A(_08538_),
    .X(net937));
 sg13g2_buf_2 fanout938 (.A(_08534_),
    .X(net938));
 sg13g2_buf_2 fanout939 (.A(_08525_),
    .X(net939));
 sg13g2_buf_4 fanout940 (.X(net940),
    .A(_08485_));
 sg13g2_buf_8 fanout941 (.A(_08484_),
    .X(net941));
 sg13g2_buf_4 fanout942 (.X(net942),
    .A(_08481_));
 sg13g2_buf_8 fanout943 (.A(_08477_),
    .X(net943));
 sg13g2_buf_2 fanout944 (.A(_08472_),
    .X(net944));
 sg13g2_buf_2 fanout945 (.A(_08436_),
    .X(net945));
 sg13g2_buf_4 fanout946 (.X(net946),
    .A(_08405_));
 sg13g2_buf_2 fanout947 (.A(_08364_),
    .X(net947));
 sg13g2_buf_2 fanout948 (.A(_08337_),
    .X(net948));
 sg13g2_buf_2 fanout949 (.A(_07374_),
    .X(net949));
 sg13g2_buf_2 fanout950 (.A(_07371_),
    .X(net950));
 sg13g2_buf_2 fanout951 (.A(_07097_),
    .X(net951));
 sg13g2_buf_2 fanout952 (.A(_07095_),
    .X(net952));
 sg13g2_buf_2 fanout953 (.A(_06937_),
    .X(net953));
 sg13g2_buf_2 fanout954 (.A(_06861_),
    .X(net954));
 sg13g2_buf_2 fanout955 (.A(_06583_),
    .X(net955));
 sg13g2_buf_2 fanout956 (.A(_06582_),
    .X(net956));
 sg13g2_buf_2 fanout957 (.A(_06581_),
    .X(net957));
 sg13g2_buf_2 fanout958 (.A(_06579_),
    .X(net958));
 sg13g2_buf_2 fanout959 (.A(_06558_),
    .X(net959));
 sg13g2_buf_2 fanout960 (.A(_06544_),
    .X(net960));
 sg13g2_buf_2 fanout961 (.A(_06520_),
    .X(net961));
 sg13g2_buf_2 fanout962 (.A(_06514_),
    .X(net962));
 sg13g2_buf_2 fanout963 (.A(_06478_),
    .X(net963));
 sg13g2_buf_2 fanout964 (.A(_06417_),
    .X(net964));
 sg13g2_buf_2 fanout965 (.A(_06127_),
    .X(net965));
 sg13g2_buf_2 fanout966 (.A(_05996_),
    .X(net966));
 sg13g2_buf_2 fanout967 (.A(_05974_),
    .X(net967));
 sg13g2_buf_2 fanout968 (.A(_05973_),
    .X(net968));
 sg13g2_buf_2 fanout969 (.A(_05972_),
    .X(net969));
 sg13g2_buf_2 fanout970 (.A(_05967_),
    .X(net970));
 sg13g2_buf_2 fanout971 (.A(_05945_),
    .X(net971));
 sg13g2_buf_2 fanout972 (.A(_05923_),
    .X(net972));
 sg13g2_buf_2 fanout973 (.A(_05922_),
    .X(net973));
 sg13g2_buf_2 fanout974 (.A(_05921_),
    .X(net974));
 sg13g2_buf_2 fanout975 (.A(_05915_),
    .X(net975));
 sg13g2_buf_2 fanout976 (.A(_05866_),
    .X(net976));
 sg13g2_buf_2 fanout977 (.A(_05865_),
    .X(net977));
 sg13g2_buf_2 fanout978 (.A(_05852_),
    .X(net978));
 sg13g2_buf_2 fanout979 (.A(_05841_),
    .X(net979));
 sg13g2_buf_2 fanout980 (.A(_05839_),
    .X(net980));
 sg13g2_buf_2 fanout981 (.A(_05156_),
    .X(net981));
 sg13g2_buf_2 fanout982 (.A(_04980_),
    .X(net982));
 sg13g2_buf_2 fanout983 (.A(_04852_),
    .X(net983));
 sg13g2_buf_2 fanout984 (.A(_04782_),
    .X(net984));
 sg13g2_buf_2 fanout985 (.A(_04774_),
    .X(net985));
 sg13g2_buf_2 fanout986 (.A(_04741_),
    .X(net986));
 sg13g2_buf_2 fanout987 (.A(_04675_),
    .X(net987));
 sg13g2_buf_2 fanout988 (.A(_04646_),
    .X(net988));
 sg13g2_buf_2 fanout989 (.A(_04612_),
    .X(net989));
 sg13g2_buf_2 fanout990 (.A(_04318_),
    .X(net990));
 sg13g2_buf_2 fanout991 (.A(_04131_),
    .X(net991));
 sg13g2_buf_2 fanout992 (.A(_03541_),
    .X(net992));
 sg13g2_buf_2 fanout993 (.A(_03489_),
    .X(net993));
 sg13g2_buf_2 fanout994 (.A(_03464_),
    .X(net994));
 sg13g2_buf_2 fanout995 (.A(_02987_),
    .X(net995));
 sg13g2_buf_2 fanout996 (.A(_02985_),
    .X(net996));
 sg13g2_buf_2 fanout997 (.A(_02983_),
    .X(net997));
 sg13g2_buf_2 fanout998 (.A(_02981_),
    .X(net998));
 sg13g2_buf_2 fanout999 (.A(_02973_),
    .X(net999));
 sg13g2_buf_2 fanout1000 (.A(_02959_),
    .X(net1000));
 sg13g2_buf_2 fanout1001 (.A(_02939_),
    .X(net1001));
 sg13g2_buf_2 fanout1002 (.A(_02861_),
    .X(net1002));
 sg13g2_buf_2 fanout1003 (.A(_02845_),
    .X(net1003));
 sg13g2_buf_2 fanout1004 (.A(_02836_),
    .X(net1004));
 sg13g2_buf_2 fanout1005 (.A(_02681_),
    .X(net1005));
 sg13g2_buf_2 fanout1006 (.A(_12788_),
    .X(net1006));
 sg13g2_buf_2 fanout1007 (.A(_12784_),
    .X(net1007));
 sg13g2_buf_2 fanout1008 (.A(_12778_),
    .X(net1008));
 sg13g2_buf_2 fanout1009 (.A(_12678_),
    .X(net1009));
 sg13g2_buf_2 fanout1010 (.A(_12564_),
    .X(net1010));
 sg13g2_buf_2 fanout1011 (.A(_12560_),
    .X(net1011));
 sg13g2_buf_2 fanout1012 (.A(_12554_),
    .X(net1012));
 sg13g2_buf_2 fanout1013 (.A(_12491_),
    .X(net1013));
 sg13g2_buf_2 fanout1014 (.A(_12371_),
    .X(net1014));
 sg13g2_buf_2 fanout1015 (.A(_12357_),
    .X(net1015));
 sg13g2_buf_2 fanout1016 (.A(_12347_),
    .X(net1016));
 sg13g2_buf_2 fanout1017 (.A(_12317_),
    .X(net1017));
 sg13g2_buf_2 fanout1018 (.A(_12281_),
    .X(net1018));
 sg13g2_buf_4 fanout1019 (.X(net1019),
    .A(_12236_));
 sg13g2_buf_4 fanout1020 (.X(net1020),
    .A(_12225_));
 sg13g2_buf_4 fanout1021 (.X(net1021),
    .A(_12218_));
 sg13g2_buf_4 fanout1022 (.X(net1022),
    .A(_12205_));
 sg13g2_buf_2 fanout1023 (.A(_12155_),
    .X(net1023));
 sg13g2_buf_2 fanout1024 (.A(_12134_),
    .X(net1024));
 sg13g2_buf_2 fanout1025 (.A(_12041_),
    .X(net1025));
 sg13g2_buf_2 fanout1026 (.A(_12038_),
    .X(net1026));
 sg13g2_buf_2 fanout1027 (.A(_12031_),
    .X(net1027));
 sg13g2_buf_2 fanout1028 (.A(_12027_),
    .X(net1028));
 sg13g2_buf_2 fanout1029 (.A(_12025_),
    .X(net1029));
 sg13g2_buf_2 fanout1030 (.A(_11973_),
    .X(net1030));
 sg13g2_buf_2 fanout1031 (.A(_11967_),
    .X(net1031));
 sg13g2_buf_2 fanout1032 (.A(_11956_),
    .X(net1032));
 sg13g2_buf_2 fanout1033 (.A(_11952_),
    .X(net1033));
 sg13g2_buf_2 fanout1034 (.A(_11662_),
    .X(net1034));
 sg13g2_buf_2 fanout1035 (.A(_11498_),
    .X(net1035));
 sg13g2_buf_2 fanout1036 (.A(_11477_),
    .X(net1036));
 sg13g2_buf_2 fanout1037 (.A(_11300_),
    .X(net1037));
 sg13g2_buf_2 fanout1038 (.A(_10915_),
    .X(net1038));
 sg13g2_buf_2 fanout1039 (.A(_10900_),
    .X(net1039));
 sg13g2_buf_2 fanout1040 (.A(_10896_),
    .X(net1040));
 sg13g2_buf_2 fanout1041 (.A(_10895_),
    .X(net1041));
 sg13g2_buf_2 fanout1042 (.A(_10813_),
    .X(net1042));
 sg13g2_buf_2 fanout1043 (.A(_10744_),
    .X(net1043));
 sg13g2_buf_2 fanout1044 (.A(_10444_),
    .X(net1044));
 sg13g2_buf_2 fanout1045 (.A(_10396_),
    .X(net1045));
 sg13g2_buf_2 fanout1046 (.A(_10297_),
    .X(net1046));
 sg13g2_buf_2 fanout1047 (.A(_10290_),
    .X(net1047));
 sg13g2_buf_2 fanout1048 (.A(_10276_),
    .X(net1048));
 sg13g2_buf_2 fanout1049 (.A(_10235_),
    .X(net1049));
 sg13g2_buf_2 fanout1050 (.A(_10224_),
    .X(net1050));
 sg13g2_buf_2 fanout1051 (.A(_10222_),
    .X(net1051));
 sg13g2_buf_2 fanout1052 (.A(_10192_),
    .X(net1052));
 sg13g2_buf_2 fanout1053 (.A(_10140_),
    .X(net1053));
 sg13g2_buf_2 fanout1054 (.A(_10121_),
    .X(net1054));
 sg13g2_buf_2 fanout1055 (.A(_10101_),
    .X(net1055));
 sg13g2_buf_2 fanout1056 (.A(_10082_),
    .X(net1056));
 sg13g2_buf_2 fanout1057 (.A(_10079_),
    .X(net1057));
 sg13g2_buf_2 fanout1058 (.A(_10073_),
    .X(net1058));
 sg13g2_buf_2 fanout1059 (.A(_10067_),
    .X(net1059));
 sg13g2_buf_2 fanout1060 (.A(_10056_),
    .X(net1060));
 sg13g2_buf_2 fanout1061 (.A(_10051_),
    .X(net1061));
 sg13g2_buf_2 fanout1062 (.A(_10033_),
    .X(net1062));
 sg13g2_buf_2 fanout1063 (.A(_09883_),
    .X(net1063));
 sg13g2_buf_2 fanout1064 (.A(_09850_),
    .X(net1064));
 sg13g2_buf_2 fanout1065 (.A(_09458_),
    .X(net1065));
 sg13g2_buf_2 fanout1066 (.A(_09430_),
    .X(net1066));
 sg13g2_buf_2 fanout1067 (.A(_09414_),
    .X(net1067));
 sg13g2_buf_2 fanout1068 (.A(_09347_),
    .X(net1068));
 sg13g2_buf_2 fanout1069 (.A(_09291_),
    .X(net1069));
 sg13g2_buf_2 fanout1070 (.A(_09289_),
    .X(net1070));
 sg13g2_buf_2 fanout1071 (.A(_09252_),
    .X(net1071));
 sg13g2_buf_2 fanout1072 (.A(_09230_),
    .X(net1072));
 sg13g2_buf_2 fanout1073 (.A(_09228_),
    .X(net1073));
 sg13g2_buf_2 fanout1074 (.A(_09214_),
    .X(net1074));
 sg13g2_buf_2 fanout1075 (.A(_08967_),
    .X(net1075));
 sg13g2_buf_2 fanout1076 (.A(_08946_),
    .X(net1076));
 sg13g2_buf_2 fanout1077 (.A(_08731_),
    .X(net1077));
 sg13g2_buf_2 fanout1078 (.A(_08709_),
    .X(net1078));
 sg13g2_buf_4 fanout1079 (.X(net1079),
    .A(_08608_));
 sg13g2_buf_2 fanout1080 (.A(_08583_),
    .X(net1080));
 sg13g2_buf_2 fanout1081 (.A(_08540_),
    .X(net1081));
 sg13g2_buf_2 fanout1082 (.A(_08533_),
    .X(net1082));
 sg13g2_buf_2 fanout1083 (.A(_08475_),
    .X(net1083));
 sg13g2_buf_2 fanout1084 (.A(_08392_),
    .X(net1084));
 sg13g2_buf_4 fanout1085 (.X(net1085),
    .A(_08390_));
 sg13g2_buf_2 fanout1086 (.A(_08384_),
    .X(net1086));
 sg13g2_buf_2 fanout1087 (.A(_08366_),
    .X(net1087));
 sg13g2_buf_4 fanout1088 (.X(net1088),
    .A(_08365_));
 sg13g2_buf_4 fanout1089 (.X(net1089),
    .A(_08351_));
 sg13g2_buf_2 fanout1090 (.A(_08336_),
    .X(net1090));
 sg13g2_buf_2 fanout1091 (.A(_08149_),
    .X(net1091));
 sg13g2_buf_2 fanout1092 (.A(_08147_),
    .X(net1092));
 sg13g2_buf_2 fanout1093 (.A(_08145_),
    .X(net1093));
 sg13g2_buf_2 fanout1094 (.A(_08090_),
    .X(net1094));
 sg13g2_buf_2 fanout1095 (.A(_07477_),
    .X(net1095));
 sg13g2_buf_2 fanout1096 (.A(_07393_),
    .X(net1096));
 sg13g2_buf_2 fanout1097 (.A(_07372_),
    .X(net1097));
 sg13g2_buf_2 fanout1098 (.A(_07370_),
    .X(net1098));
 sg13g2_buf_2 fanout1099 (.A(_02849_),
    .X(net1099));
 sg13g2_buf_1 fanout1100 (.A(_12276_),
    .X(net1100));
 sg13g2_buf_2 fanout1101 (.A(_12273_),
    .X(net1101));
 sg13g2_buf_1 fanout1102 (.A(_12266_),
    .X(net1102));
 sg13g2_buf_2 fanout1103 (.A(_12235_),
    .X(net1103));
 sg13g2_buf_2 fanout1104 (.A(_12224_),
    .X(net1104));
 sg13g2_buf_2 fanout1105 (.A(_12217_),
    .X(net1105));
 sg13g2_buf_2 fanout1106 (.A(_12204_),
    .X(net1106));
 sg13g2_buf_2 fanout1107 (.A(_12099_),
    .X(net1107));
 sg13g2_buf_2 fanout1108 (.A(_12081_),
    .X(net1108));
 sg13g2_buf_2 fanout1109 (.A(_12060_),
    .X(net1109));
 sg13g2_buf_2 fanout1110 (.A(_12021_),
    .X(net1110));
 sg13g2_buf_2 fanout1111 (.A(_12018_),
    .X(net1111));
 sg13g2_buf_2 fanout1112 (.A(_11999_),
    .X(net1112));
 sg13g2_buf_2 fanout1113 (.A(_11997_),
    .X(net1113));
 sg13g2_buf_2 fanout1114 (.A(_11990_),
    .X(net1114));
 sg13g2_buf_2 fanout1115 (.A(_11955_),
    .X(net1115));
 sg13g2_buf_2 fanout1116 (.A(_11719_),
    .X(net1116));
 sg13g2_buf_2 fanout1117 (.A(_11043_),
    .X(net1117));
 sg13g2_buf_2 fanout1118 (.A(_10888_),
    .X(net1118));
 sg13g2_buf_2 fanout1119 (.A(_10886_),
    .X(net1119));
 sg13g2_buf_2 fanout1120 (.A(_10810_),
    .X(net1120));
 sg13g2_buf_2 fanout1121 (.A(_10558_),
    .X(net1121));
 sg13g2_buf_2 fanout1122 (.A(_10379_),
    .X(net1122));
 sg13g2_buf_2 fanout1123 (.A(_10214_),
    .X(net1123));
 sg13g2_buf_2 fanout1124 (.A(_10196_),
    .X(net1124));
 sg13g2_buf_2 fanout1125 (.A(_10195_),
    .X(net1125));
 sg13g2_buf_2 fanout1126 (.A(_10190_),
    .X(net1126));
 sg13g2_buf_2 fanout1127 (.A(_10188_),
    .X(net1127));
 sg13g2_buf_2 fanout1128 (.A(_10060_),
    .X(net1128));
 sg13g2_buf_2 fanout1129 (.A(_09948_),
    .X(net1129));
 sg13g2_buf_2 fanout1130 (.A(_09891_),
    .X(net1130));
 sg13g2_buf_2 fanout1131 (.A(_09882_),
    .X(net1131));
 sg13g2_buf_2 fanout1132 (.A(_09604_),
    .X(net1132));
 sg13g2_buf_2 fanout1133 (.A(_09353_),
    .X(net1133));
 sg13g2_buf_2 fanout1134 (.A(_09313_),
    .X(net1134));
 sg13g2_buf_2 fanout1135 (.A(_09305_),
    .X(net1135));
 sg13g2_buf_2 fanout1136 (.A(_09239_),
    .X(net1136));
 sg13g2_buf_2 fanout1137 (.A(_09238_),
    .X(net1137));
 sg13g2_buf_4 fanout1138 (.X(net1138),
    .A(_09222_));
 sg13g2_buf_4 fanout1139 (.X(net1139),
    .A(_09221_));
 sg13g2_buf_2 fanout1140 (.A(_09136_),
    .X(net1140));
 sg13g2_buf_2 fanout1141 (.A(_08502_),
    .X(net1141));
 sg13g2_buf_2 fanout1142 (.A(_08499_),
    .X(net1142));
 sg13g2_buf_2 fanout1143 (.A(_08454_),
    .X(net1143));
 sg13g2_buf_2 fanout1144 (.A(_08453_),
    .X(net1144));
 sg13g2_buf_2 fanout1145 (.A(_08452_),
    .X(net1145));
 sg13g2_buf_2 fanout1146 (.A(_08403_),
    .X(net1146));
 sg13g2_buf_4 fanout1147 (.X(net1147),
    .A(_08395_));
 sg13g2_buf_4 fanout1148 (.X(net1148),
    .A(_08355_));
 sg13g2_buf_2 fanout1149 (.A(_08338_),
    .X(net1149));
 sg13g2_tiehi _27720__1150 (.L_HI(net1150));
 sg13g2_tiehi _27721__1151 (.L_HI(net1151));
 sg13g2_tiehi _27722__1152 (.L_HI(net1152));
 sg13g2_tiehi _27723__1153 (.L_HI(net1153));
 sg13g2_tiehi _27724__1154 (.L_HI(net1154));
 sg13g2_tiehi \cpu.dcache.r_data[0][0]$_DFFE_PP__1155  (.L_HI(net1155));
 sg13g2_tiehi \cpu.dcache.r_data[0][10]$_DFFE_PP__1156  (.L_HI(net1156));
 sg13g2_tiehi \cpu.dcache.r_data[0][11]$_DFFE_PP__1157  (.L_HI(net1157));
 sg13g2_tiehi \cpu.dcache.r_data[0][12]$_DFFE_PP__1158  (.L_HI(net1158));
 sg13g2_tiehi \cpu.dcache.r_data[0][13]$_DFFE_PP__1159  (.L_HI(net1159));
 sg13g2_tiehi \cpu.dcache.r_data[0][14]$_DFFE_PP__1160  (.L_HI(net1160));
 sg13g2_tiehi \cpu.dcache.r_data[0][15]$_DFFE_PP__1161  (.L_HI(net1161));
 sg13g2_tiehi \cpu.dcache.r_data[0][16]$_DFFE_PP__1162  (.L_HI(net1162));
 sg13g2_tiehi \cpu.dcache.r_data[0][17]$_DFFE_PP__1163  (.L_HI(net1163));
 sg13g2_tiehi \cpu.dcache.r_data[0][18]$_DFFE_PP__1164  (.L_HI(net1164));
 sg13g2_tiehi \cpu.dcache.r_data[0][19]$_DFFE_PP__1165  (.L_HI(net1165));
 sg13g2_tiehi \cpu.dcache.r_data[0][1]$_DFFE_PP__1166  (.L_HI(net1166));
 sg13g2_tiehi \cpu.dcache.r_data[0][20]$_DFFE_PP__1167  (.L_HI(net1167));
 sg13g2_tiehi \cpu.dcache.r_data[0][21]$_DFFE_PP__1168  (.L_HI(net1168));
 sg13g2_tiehi \cpu.dcache.r_data[0][22]$_DFFE_PP__1169  (.L_HI(net1169));
 sg13g2_tiehi \cpu.dcache.r_data[0][23]$_DFFE_PP__1170  (.L_HI(net1170));
 sg13g2_tiehi \cpu.dcache.r_data[0][24]$_DFFE_PP__1171  (.L_HI(net1171));
 sg13g2_tiehi \cpu.dcache.r_data[0][25]$_DFFE_PP__1172  (.L_HI(net1172));
 sg13g2_tiehi \cpu.dcache.r_data[0][26]$_DFFE_PP__1173  (.L_HI(net1173));
 sg13g2_tiehi \cpu.dcache.r_data[0][27]$_DFFE_PP__1174  (.L_HI(net1174));
 sg13g2_tiehi \cpu.dcache.r_data[0][28]$_DFFE_PP__1175  (.L_HI(net1175));
 sg13g2_tiehi \cpu.dcache.r_data[0][29]$_DFFE_PP__1176  (.L_HI(net1176));
 sg13g2_tiehi \cpu.dcache.r_data[0][2]$_DFFE_PP__1177  (.L_HI(net1177));
 sg13g2_tiehi \cpu.dcache.r_data[0][30]$_DFFE_PP__1178  (.L_HI(net1178));
 sg13g2_tiehi \cpu.dcache.r_data[0][31]$_DFFE_PP__1179  (.L_HI(net1179));
 sg13g2_tiehi \cpu.dcache.r_data[0][3]$_DFFE_PP__1180  (.L_HI(net1180));
 sg13g2_tiehi \cpu.dcache.r_data[0][4]$_DFFE_PP__1181  (.L_HI(net1181));
 sg13g2_tiehi \cpu.dcache.r_data[0][5]$_DFFE_PP__1182  (.L_HI(net1182));
 sg13g2_tiehi \cpu.dcache.r_data[0][6]$_DFFE_PP__1183  (.L_HI(net1183));
 sg13g2_tiehi \cpu.dcache.r_data[0][7]$_DFFE_PP__1184  (.L_HI(net1184));
 sg13g2_tiehi \cpu.dcache.r_data[0][8]$_DFFE_PP__1185  (.L_HI(net1185));
 sg13g2_tiehi \cpu.dcache.r_data[0][9]$_DFFE_PP__1186  (.L_HI(net1186));
 sg13g2_tiehi \cpu.dcache.r_data[1][0]$_DFFE_PP__1187  (.L_HI(net1187));
 sg13g2_tiehi \cpu.dcache.r_data[1][10]$_DFFE_PP__1188  (.L_HI(net1188));
 sg13g2_tiehi \cpu.dcache.r_data[1][11]$_DFFE_PP__1189  (.L_HI(net1189));
 sg13g2_tiehi \cpu.dcache.r_data[1][12]$_DFFE_PP__1190  (.L_HI(net1190));
 sg13g2_tiehi \cpu.dcache.r_data[1][13]$_DFFE_PP__1191  (.L_HI(net1191));
 sg13g2_tiehi \cpu.dcache.r_data[1][14]$_DFFE_PP__1192  (.L_HI(net1192));
 sg13g2_tiehi \cpu.dcache.r_data[1][15]$_DFFE_PP__1193  (.L_HI(net1193));
 sg13g2_tiehi \cpu.dcache.r_data[1][16]$_DFFE_PP__1194  (.L_HI(net1194));
 sg13g2_tiehi \cpu.dcache.r_data[1][17]$_DFFE_PP__1195  (.L_HI(net1195));
 sg13g2_tiehi \cpu.dcache.r_data[1][18]$_DFFE_PP__1196  (.L_HI(net1196));
 sg13g2_tiehi \cpu.dcache.r_data[1][19]$_DFFE_PP__1197  (.L_HI(net1197));
 sg13g2_tiehi \cpu.dcache.r_data[1][1]$_DFFE_PP__1198  (.L_HI(net1198));
 sg13g2_tiehi \cpu.dcache.r_data[1][20]$_DFFE_PP__1199  (.L_HI(net1199));
 sg13g2_tiehi \cpu.dcache.r_data[1][21]$_DFFE_PP__1200  (.L_HI(net1200));
 sg13g2_tiehi \cpu.dcache.r_data[1][22]$_DFFE_PP__1201  (.L_HI(net1201));
 sg13g2_tiehi \cpu.dcache.r_data[1][23]$_DFFE_PP__1202  (.L_HI(net1202));
 sg13g2_tiehi \cpu.dcache.r_data[1][24]$_DFFE_PP__1203  (.L_HI(net1203));
 sg13g2_tiehi \cpu.dcache.r_data[1][25]$_DFFE_PP__1204  (.L_HI(net1204));
 sg13g2_tiehi \cpu.dcache.r_data[1][26]$_DFFE_PP__1205  (.L_HI(net1205));
 sg13g2_tiehi \cpu.dcache.r_data[1][27]$_DFFE_PP__1206  (.L_HI(net1206));
 sg13g2_tiehi \cpu.dcache.r_data[1][28]$_DFFE_PP__1207  (.L_HI(net1207));
 sg13g2_tiehi \cpu.dcache.r_data[1][29]$_DFFE_PP__1208  (.L_HI(net1208));
 sg13g2_tiehi \cpu.dcache.r_data[1][2]$_DFFE_PP__1209  (.L_HI(net1209));
 sg13g2_tiehi \cpu.dcache.r_data[1][30]$_DFFE_PP__1210  (.L_HI(net1210));
 sg13g2_tiehi \cpu.dcache.r_data[1][31]$_DFFE_PP__1211  (.L_HI(net1211));
 sg13g2_tiehi \cpu.dcache.r_data[1][3]$_DFFE_PP__1212  (.L_HI(net1212));
 sg13g2_tiehi \cpu.dcache.r_data[1][4]$_DFFE_PP__1213  (.L_HI(net1213));
 sg13g2_tiehi \cpu.dcache.r_data[1][5]$_DFFE_PP__1214  (.L_HI(net1214));
 sg13g2_tiehi \cpu.dcache.r_data[1][6]$_DFFE_PP__1215  (.L_HI(net1215));
 sg13g2_tiehi \cpu.dcache.r_data[1][7]$_DFFE_PP__1216  (.L_HI(net1216));
 sg13g2_tiehi \cpu.dcache.r_data[1][8]$_DFFE_PP__1217  (.L_HI(net1217));
 sg13g2_tiehi \cpu.dcache.r_data[1][9]$_DFFE_PP__1218  (.L_HI(net1218));
 sg13g2_tiehi \cpu.dcache.r_data[2][0]$_DFFE_PP__1219  (.L_HI(net1219));
 sg13g2_tiehi \cpu.dcache.r_data[2][10]$_DFFE_PP__1220  (.L_HI(net1220));
 sg13g2_tiehi \cpu.dcache.r_data[2][11]$_DFFE_PP__1221  (.L_HI(net1221));
 sg13g2_tiehi \cpu.dcache.r_data[2][12]$_DFFE_PP__1222  (.L_HI(net1222));
 sg13g2_tiehi \cpu.dcache.r_data[2][13]$_DFFE_PP__1223  (.L_HI(net1223));
 sg13g2_tiehi \cpu.dcache.r_data[2][14]$_DFFE_PP__1224  (.L_HI(net1224));
 sg13g2_tiehi \cpu.dcache.r_data[2][15]$_DFFE_PP__1225  (.L_HI(net1225));
 sg13g2_tiehi \cpu.dcache.r_data[2][16]$_DFFE_PP__1226  (.L_HI(net1226));
 sg13g2_tiehi \cpu.dcache.r_data[2][17]$_DFFE_PP__1227  (.L_HI(net1227));
 sg13g2_tiehi \cpu.dcache.r_data[2][18]$_DFFE_PP__1228  (.L_HI(net1228));
 sg13g2_tiehi \cpu.dcache.r_data[2][19]$_DFFE_PP__1229  (.L_HI(net1229));
 sg13g2_tiehi \cpu.dcache.r_data[2][1]$_DFFE_PP__1230  (.L_HI(net1230));
 sg13g2_tiehi \cpu.dcache.r_data[2][20]$_DFFE_PP__1231  (.L_HI(net1231));
 sg13g2_tiehi \cpu.dcache.r_data[2][21]$_DFFE_PP__1232  (.L_HI(net1232));
 sg13g2_tiehi \cpu.dcache.r_data[2][22]$_DFFE_PP__1233  (.L_HI(net1233));
 sg13g2_tiehi \cpu.dcache.r_data[2][23]$_DFFE_PP__1234  (.L_HI(net1234));
 sg13g2_tiehi \cpu.dcache.r_data[2][24]$_DFFE_PP__1235  (.L_HI(net1235));
 sg13g2_tiehi \cpu.dcache.r_data[2][25]$_DFFE_PP__1236  (.L_HI(net1236));
 sg13g2_tiehi \cpu.dcache.r_data[2][26]$_DFFE_PP__1237  (.L_HI(net1237));
 sg13g2_tiehi \cpu.dcache.r_data[2][27]$_DFFE_PP__1238  (.L_HI(net1238));
 sg13g2_tiehi \cpu.dcache.r_data[2][28]$_DFFE_PP__1239  (.L_HI(net1239));
 sg13g2_tiehi \cpu.dcache.r_data[2][29]$_DFFE_PP__1240  (.L_HI(net1240));
 sg13g2_tiehi \cpu.dcache.r_data[2][2]$_DFFE_PP__1241  (.L_HI(net1241));
 sg13g2_tiehi \cpu.dcache.r_data[2][30]$_DFFE_PP__1242  (.L_HI(net1242));
 sg13g2_tiehi \cpu.dcache.r_data[2][31]$_DFFE_PP__1243  (.L_HI(net1243));
 sg13g2_tiehi \cpu.dcache.r_data[2][3]$_DFFE_PP__1244  (.L_HI(net1244));
 sg13g2_tiehi \cpu.dcache.r_data[2][4]$_DFFE_PP__1245  (.L_HI(net1245));
 sg13g2_tiehi \cpu.dcache.r_data[2][5]$_DFFE_PP__1246  (.L_HI(net1246));
 sg13g2_tiehi \cpu.dcache.r_data[2][6]$_DFFE_PP__1247  (.L_HI(net1247));
 sg13g2_tiehi \cpu.dcache.r_data[2][7]$_DFFE_PP__1248  (.L_HI(net1248));
 sg13g2_tiehi \cpu.dcache.r_data[2][8]$_DFFE_PP__1249  (.L_HI(net1249));
 sg13g2_tiehi \cpu.dcache.r_data[2][9]$_DFFE_PP__1250  (.L_HI(net1250));
 sg13g2_tiehi \cpu.dcache.r_data[3][0]$_DFFE_PP__1251  (.L_HI(net1251));
 sg13g2_tiehi \cpu.dcache.r_data[3][10]$_DFFE_PP__1252  (.L_HI(net1252));
 sg13g2_tiehi \cpu.dcache.r_data[3][11]$_DFFE_PP__1253  (.L_HI(net1253));
 sg13g2_tiehi \cpu.dcache.r_data[3][12]$_DFFE_PP__1254  (.L_HI(net1254));
 sg13g2_tiehi \cpu.dcache.r_data[3][13]$_DFFE_PP__1255  (.L_HI(net1255));
 sg13g2_tiehi \cpu.dcache.r_data[3][14]$_DFFE_PP__1256  (.L_HI(net1256));
 sg13g2_tiehi \cpu.dcache.r_data[3][15]$_DFFE_PP__1257  (.L_HI(net1257));
 sg13g2_tiehi \cpu.dcache.r_data[3][16]$_DFFE_PP__1258  (.L_HI(net1258));
 sg13g2_tiehi \cpu.dcache.r_data[3][17]$_DFFE_PP__1259  (.L_HI(net1259));
 sg13g2_tiehi \cpu.dcache.r_data[3][18]$_DFFE_PP__1260  (.L_HI(net1260));
 sg13g2_tiehi \cpu.dcache.r_data[3][19]$_DFFE_PP__1261  (.L_HI(net1261));
 sg13g2_tiehi \cpu.dcache.r_data[3][1]$_DFFE_PP__1262  (.L_HI(net1262));
 sg13g2_tiehi \cpu.dcache.r_data[3][20]$_DFFE_PP__1263  (.L_HI(net1263));
 sg13g2_tiehi \cpu.dcache.r_data[3][21]$_DFFE_PP__1264  (.L_HI(net1264));
 sg13g2_tiehi \cpu.dcache.r_data[3][22]$_DFFE_PP__1265  (.L_HI(net1265));
 sg13g2_tiehi \cpu.dcache.r_data[3][23]$_DFFE_PP__1266  (.L_HI(net1266));
 sg13g2_tiehi \cpu.dcache.r_data[3][24]$_DFFE_PP__1267  (.L_HI(net1267));
 sg13g2_tiehi \cpu.dcache.r_data[3][25]$_DFFE_PP__1268  (.L_HI(net1268));
 sg13g2_tiehi \cpu.dcache.r_data[3][26]$_DFFE_PP__1269  (.L_HI(net1269));
 sg13g2_tiehi \cpu.dcache.r_data[3][27]$_DFFE_PP__1270  (.L_HI(net1270));
 sg13g2_tiehi \cpu.dcache.r_data[3][28]$_DFFE_PP__1271  (.L_HI(net1271));
 sg13g2_tiehi \cpu.dcache.r_data[3][29]$_DFFE_PP__1272  (.L_HI(net1272));
 sg13g2_tiehi \cpu.dcache.r_data[3][2]$_DFFE_PP__1273  (.L_HI(net1273));
 sg13g2_tiehi \cpu.dcache.r_data[3][30]$_DFFE_PP__1274  (.L_HI(net1274));
 sg13g2_tiehi \cpu.dcache.r_data[3][31]$_DFFE_PP__1275  (.L_HI(net1275));
 sg13g2_tiehi \cpu.dcache.r_data[3][3]$_DFFE_PP__1276  (.L_HI(net1276));
 sg13g2_tiehi \cpu.dcache.r_data[3][4]$_DFFE_PP__1277  (.L_HI(net1277));
 sg13g2_tiehi \cpu.dcache.r_data[3][5]$_DFFE_PP__1278  (.L_HI(net1278));
 sg13g2_tiehi \cpu.dcache.r_data[3][6]$_DFFE_PP__1279  (.L_HI(net1279));
 sg13g2_tiehi \cpu.dcache.r_data[3][7]$_DFFE_PP__1280  (.L_HI(net1280));
 sg13g2_tiehi \cpu.dcache.r_data[3][8]$_DFFE_PP__1281  (.L_HI(net1281));
 sg13g2_tiehi \cpu.dcache.r_data[3][9]$_DFFE_PP__1282  (.L_HI(net1282));
 sg13g2_tiehi \cpu.dcache.r_data[4][0]$_DFFE_PP__1283  (.L_HI(net1283));
 sg13g2_tiehi \cpu.dcache.r_data[4][10]$_DFFE_PP__1284  (.L_HI(net1284));
 sg13g2_tiehi \cpu.dcache.r_data[4][11]$_DFFE_PP__1285  (.L_HI(net1285));
 sg13g2_tiehi \cpu.dcache.r_data[4][12]$_DFFE_PP__1286  (.L_HI(net1286));
 sg13g2_tiehi \cpu.dcache.r_data[4][13]$_DFFE_PP__1287  (.L_HI(net1287));
 sg13g2_tiehi \cpu.dcache.r_data[4][14]$_DFFE_PP__1288  (.L_HI(net1288));
 sg13g2_tiehi \cpu.dcache.r_data[4][15]$_DFFE_PP__1289  (.L_HI(net1289));
 sg13g2_tiehi \cpu.dcache.r_data[4][16]$_DFFE_PP__1290  (.L_HI(net1290));
 sg13g2_tiehi \cpu.dcache.r_data[4][17]$_DFFE_PP__1291  (.L_HI(net1291));
 sg13g2_tiehi \cpu.dcache.r_data[4][18]$_DFFE_PP__1292  (.L_HI(net1292));
 sg13g2_tiehi \cpu.dcache.r_data[4][19]$_DFFE_PP__1293  (.L_HI(net1293));
 sg13g2_tiehi \cpu.dcache.r_data[4][1]$_DFFE_PP__1294  (.L_HI(net1294));
 sg13g2_tiehi \cpu.dcache.r_data[4][20]$_DFFE_PP__1295  (.L_HI(net1295));
 sg13g2_tiehi \cpu.dcache.r_data[4][21]$_DFFE_PP__1296  (.L_HI(net1296));
 sg13g2_tiehi \cpu.dcache.r_data[4][22]$_DFFE_PP__1297  (.L_HI(net1297));
 sg13g2_tiehi \cpu.dcache.r_data[4][23]$_DFFE_PP__1298  (.L_HI(net1298));
 sg13g2_tiehi \cpu.dcache.r_data[4][24]$_DFFE_PP__1299  (.L_HI(net1299));
 sg13g2_tiehi \cpu.dcache.r_data[4][25]$_DFFE_PP__1300  (.L_HI(net1300));
 sg13g2_tiehi \cpu.dcache.r_data[4][26]$_DFFE_PP__1301  (.L_HI(net1301));
 sg13g2_tiehi \cpu.dcache.r_data[4][27]$_DFFE_PP__1302  (.L_HI(net1302));
 sg13g2_tiehi \cpu.dcache.r_data[4][28]$_DFFE_PP__1303  (.L_HI(net1303));
 sg13g2_tiehi \cpu.dcache.r_data[4][29]$_DFFE_PP__1304  (.L_HI(net1304));
 sg13g2_tiehi \cpu.dcache.r_data[4][2]$_DFFE_PP__1305  (.L_HI(net1305));
 sg13g2_tiehi \cpu.dcache.r_data[4][30]$_DFFE_PP__1306  (.L_HI(net1306));
 sg13g2_tiehi \cpu.dcache.r_data[4][31]$_DFFE_PP__1307  (.L_HI(net1307));
 sg13g2_tiehi \cpu.dcache.r_data[4][3]$_DFFE_PP__1308  (.L_HI(net1308));
 sg13g2_tiehi \cpu.dcache.r_data[4][4]$_DFFE_PP__1309  (.L_HI(net1309));
 sg13g2_tiehi \cpu.dcache.r_data[4][5]$_DFFE_PP__1310  (.L_HI(net1310));
 sg13g2_tiehi \cpu.dcache.r_data[4][6]$_DFFE_PP__1311  (.L_HI(net1311));
 sg13g2_tiehi \cpu.dcache.r_data[4][7]$_DFFE_PP__1312  (.L_HI(net1312));
 sg13g2_tiehi \cpu.dcache.r_data[4][8]$_DFFE_PP__1313  (.L_HI(net1313));
 sg13g2_tiehi \cpu.dcache.r_data[4][9]$_DFFE_PP__1314  (.L_HI(net1314));
 sg13g2_tiehi \cpu.dcache.r_data[5][0]$_DFFE_PP__1315  (.L_HI(net1315));
 sg13g2_tiehi \cpu.dcache.r_data[5][10]$_DFFE_PP__1316  (.L_HI(net1316));
 sg13g2_tiehi \cpu.dcache.r_data[5][11]$_DFFE_PP__1317  (.L_HI(net1317));
 sg13g2_tiehi \cpu.dcache.r_data[5][12]$_DFFE_PP__1318  (.L_HI(net1318));
 sg13g2_tiehi \cpu.dcache.r_data[5][13]$_DFFE_PP__1319  (.L_HI(net1319));
 sg13g2_tiehi \cpu.dcache.r_data[5][14]$_DFFE_PP__1320  (.L_HI(net1320));
 sg13g2_tiehi \cpu.dcache.r_data[5][15]$_DFFE_PP__1321  (.L_HI(net1321));
 sg13g2_tiehi \cpu.dcache.r_data[5][16]$_DFFE_PP__1322  (.L_HI(net1322));
 sg13g2_tiehi \cpu.dcache.r_data[5][17]$_DFFE_PP__1323  (.L_HI(net1323));
 sg13g2_tiehi \cpu.dcache.r_data[5][18]$_DFFE_PP__1324  (.L_HI(net1324));
 sg13g2_tiehi \cpu.dcache.r_data[5][19]$_DFFE_PP__1325  (.L_HI(net1325));
 sg13g2_tiehi \cpu.dcache.r_data[5][1]$_DFFE_PP__1326  (.L_HI(net1326));
 sg13g2_tiehi \cpu.dcache.r_data[5][20]$_DFFE_PP__1327  (.L_HI(net1327));
 sg13g2_tiehi \cpu.dcache.r_data[5][21]$_DFFE_PP__1328  (.L_HI(net1328));
 sg13g2_tiehi \cpu.dcache.r_data[5][22]$_DFFE_PP__1329  (.L_HI(net1329));
 sg13g2_tiehi \cpu.dcache.r_data[5][23]$_DFFE_PP__1330  (.L_HI(net1330));
 sg13g2_tiehi \cpu.dcache.r_data[5][24]$_DFFE_PP__1331  (.L_HI(net1331));
 sg13g2_tiehi \cpu.dcache.r_data[5][25]$_DFFE_PP__1332  (.L_HI(net1332));
 sg13g2_tiehi \cpu.dcache.r_data[5][26]$_DFFE_PP__1333  (.L_HI(net1333));
 sg13g2_tiehi \cpu.dcache.r_data[5][27]$_DFFE_PP__1334  (.L_HI(net1334));
 sg13g2_tiehi \cpu.dcache.r_data[5][28]$_DFFE_PP__1335  (.L_HI(net1335));
 sg13g2_tiehi \cpu.dcache.r_data[5][29]$_DFFE_PP__1336  (.L_HI(net1336));
 sg13g2_tiehi \cpu.dcache.r_data[5][2]$_DFFE_PP__1337  (.L_HI(net1337));
 sg13g2_tiehi \cpu.dcache.r_data[5][30]$_DFFE_PP__1338  (.L_HI(net1338));
 sg13g2_tiehi \cpu.dcache.r_data[5][31]$_DFFE_PP__1339  (.L_HI(net1339));
 sg13g2_tiehi \cpu.dcache.r_data[5][3]$_DFFE_PP__1340  (.L_HI(net1340));
 sg13g2_tiehi \cpu.dcache.r_data[5][4]$_DFFE_PP__1341  (.L_HI(net1341));
 sg13g2_tiehi \cpu.dcache.r_data[5][5]$_DFFE_PP__1342  (.L_HI(net1342));
 sg13g2_tiehi \cpu.dcache.r_data[5][6]$_DFFE_PP__1343  (.L_HI(net1343));
 sg13g2_tiehi \cpu.dcache.r_data[5][7]$_DFFE_PP__1344  (.L_HI(net1344));
 sg13g2_tiehi \cpu.dcache.r_data[5][8]$_DFFE_PP__1345  (.L_HI(net1345));
 sg13g2_tiehi \cpu.dcache.r_data[5][9]$_DFFE_PP__1346  (.L_HI(net1346));
 sg13g2_tiehi \cpu.dcache.r_data[6][0]$_DFFE_PP__1347  (.L_HI(net1347));
 sg13g2_tiehi \cpu.dcache.r_data[6][10]$_DFFE_PP__1348  (.L_HI(net1348));
 sg13g2_tiehi \cpu.dcache.r_data[6][11]$_DFFE_PP__1349  (.L_HI(net1349));
 sg13g2_tiehi \cpu.dcache.r_data[6][12]$_DFFE_PP__1350  (.L_HI(net1350));
 sg13g2_tiehi \cpu.dcache.r_data[6][13]$_DFFE_PP__1351  (.L_HI(net1351));
 sg13g2_tiehi \cpu.dcache.r_data[6][14]$_DFFE_PP__1352  (.L_HI(net1352));
 sg13g2_tiehi \cpu.dcache.r_data[6][15]$_DFFE_PP__1353  (.L_HI(net1353));
 sg13g2_tiehi \cpu.dcache.r_data[6][16]$_DFFE_PP__1354  (.L_HI(net1354));
 sg13g2_tiehi \cpu.dcache.r_data[6][17]$_DFFE_PP__1355  (.L_HI(net1355));
 sg13g2_tiehi \cpu.dcache.r_data[6][18]$_DFFE_PP__1356  (.L_HI(net1356));
 sg13g2_tiehi \cpu.dcache.r_data[6][19]$_DFFE_PP__1357  (.L_HI(net1357));
 sg13g2_tiehi \cpu.dcache.r_data[6][1]$_DFFE_PP__1358  (.L_HI(net1358));
 sg13g2_tiehi \cpu.dcache.r_data[6][20]$_DFFE_PP__1359  (.L_HI(net1359));
 sg13g2_tiehi \cpu.dcache.r_data[6][21]$_DFFE_PP__1360  (.L_HI(net1360));
 sg13g2_tiehi \cpu.dcache.r_data[6][22]$_DFFE_PP__1361  (.L_HI(net1361));
 sg13g2_tiehi \cpu.dcache.r_data[6][23]$_DFFE_PP__1362  (.L_HI(net1362));
 sg13g2_tiehi \cpu.dcache.r_data[6][24]$_DFFE_PP__1363  (.L_HI(net1363));
 sg13g2_tiehi \cpu.dcache.r_data[6][25]$_DFFE_PP__1364  (.L_HI(net1364));
 sg13g2_tiehi \cpu.dcache.r_data[6][26]$_DFFE_PP__1365  (.L_HI(net1365));
 sg13g2_tiehi \cpu.dcache.r_data[6][27]$_DFFE_PP__1366  (.L_HI(net1366));
 sg13g2_tiehi \cpu.dcache.r_data[6][28]$_DFFE_PP__1367  (.L_HI(net1367));
 sg13g2_tiehi \cpu.dcache.r_data[6][29]$_DFFE_PP__1368  (.L_HI(net1368));
 sg13g2_tiehi \cpu.dcache.r_data[6][2]$_DFFE_PP__1369  (.L_HI(net1369));
 sg13g2_tiehi \cpu.dcache.r_data[6][30]$_DFFE_PP__1370  (.L_HI(net1370));
 sg13g2_tiehi \cpu.dcache.r_data[6][31]$_DFFE_PP__1371  (.L_HI(net1371));
 sg13g2_tiehi \cpu.dcache.r_data[6][3]$_DFFE_PP__1372  (.L_HI(net1372));
 sg13g2_tiehi \cpu.dcache.r_data[6][4]$_DFFE_PP__1373  (.L_HI(net1373));
 sg13g2_tiehi \cpu.dcache.r_data[6][5]$_DFFE_PP__1374  (.L_HI(net1374));
 sg13g2_tiehi \cpu.dcache.r_data[6][6]$_DFFE_PP__1375  (.L_HI(net1375));
 sg13g2_tiehi \cpu.dcache.r_data[6][7]$_DFFE_PP__1376  (.L_HI(net1376));
 sg13g2_tiehi \cpu.dcache.r_data[6][8]$_DFFE_PP__1377  (.L_HI(net1377));
 sg13g2_tiehi \cpu.dcache.r_data[6][9]$_DFFE_PP__1378  (.L_HI(net1378));
 sg13g2_tiehi \cpu.dcache.r_data[7][0]$_DFFE_PP__1379  (.L_HI(net1379));
 sg13g2_tiehi \cpu.dcache.r_data[7][10]$_DFFE_PP__1380  (.L_HI(net1380));
 sg13g2_tiehi \cpu.dcache.r_data[7][11]$_DFFE_PP__1381  (.L_HI(net1381));
 sg13g2_tiehi \cpu.dcache.r_data[7][12]$_DFFE_PP__1382  (.L_HI(net1382));
 sg13g2_tiehi \cpu.dcache.r_data[7][13]$_DFFE_PP__1383  (.L_HI(net1383));
 sg13g2_tiehi \cpu.dcache.r_data[7][14]$_DFFE_PP__1384  (.L_HI(net1384));
 sg13g2_tiehi \cpu.dcache.r_data[7][15]$_DFFE_PP__1385  (.L_HI(net1385));
 sg13g2_tiehi \cpu.dcache.r_data[7][16]$_DFFE_PP__1386  (.L_HI(net1386));
 sg13g2_tiehi \cpu.dcache.r_data[7][17]$_DFFE_PP__1387  (.L_HI(net1387));
 sg13g2_tiehi \cpu.dcache.r_data[7][18]$_DFFE_PP__1388  (.L_HI(net1388));
 sg13g2_tiehi \cpu.dcache.r_data[7][19]$_DFFE_PP__1389  (.L_HI(net1389));
 sg13g2_tiehi \cpu.dcache.r_data[7][1]$_DFFE_PP__1390  (.L_HI(net1390));
 sg13g2_tiehi \cpu.dcache.r_data[7][20]$_DFFE_PP__1391  (.L_HI(net1391));
 sg13g2_tiehi \cpu.dcache.r_data[7][21]$_DFFE_PP__1392  (.L_HI(net1392));
 sg13g2_tiehi \cpu.dcache.r_data[7][22]$_DFFE_PP__1393  (.L_HI(net1393));
 sg13g2_tiehi \cpu.dcache.r_data[7][23]$_DFFE_PP__1394  (.L_HI(net1394));
 sg13g2_tiehi \cpu.dcache.r_data[7][24]$_DFFE_PP__1395  (.L_HI(net1395));
 sg13g2_tiehi \cpu.dcache.r_data[7][25]$_DFFE_PP__1396  (.L_HI(net1396));
 sg13g2_tiehi \cpu.dcache.r_data[7][26]$_DFFE_PP__1397  (.L_HI(net1397));
 sg13g2_tiehi \cpu.dcache.r_data[7][27]$_DFFE_PP__1398  (.L_HI(net1398));
 sg13g2_tiehi \cpu.dcache.r_data[7][28]$_DFFE_PP__1399  (.L_HI(net1399));
 sg13g2_tiehi \cpu.dcache.r_data[7][29]$_DFFE_PP__1400  (.L_HI(net1400));
 sg13g2_tiehi \cpu.dcache.r_data[7][2]$_DFFE_PP__1401  (.L_HI(net1401));
 sg13g2_tiehi \cpu.dcache.r_data[7][30]$_DFFE_PP__1402  (.L_HI(net1402));
 sg13g2_tiehi \cpu.dcache.r_data[7][31]$_DFFE_PP__1403  (.L_HI(net1403));
 sg13g2_tiehi \cpu.dcache.r_data[7][3]$_DFFE_PP__1404  (.L_HI(net1404));
 sg13g2_tiehi \cpu.dcache.r_data[7][4]$_DFFE_PP__1405  (.L_HI(net1405));
 sg13g2_tiehi \cpu.dcache.r_data[7][5]$_DFFE_PP__1406  (.L_HI(net1406));
 sg13g2_tiehi \cpu.dcache.r_data[7][6]$_DFFE_PP__1407  (.L_HI(net1407));
 sg13g2_tiehi \cpu.dcache.r_data[7][7]$_DFFE_PP__1408  (.L_HI(net1408));
 sg13g2_tiehi \cpu.dcache.r_data[7][8]$_DFFE_PP__1409  (.L_HI(net1409));
 sg13g2_tiehi \cpu.dcache.r_data[7][9]$_DFFE_PP__1410  (.L_HI(net1410));
 sg13g2_tiehi \cpu.dcache.r_dirty[0]$_SDFFCE_PP1P__1411  (.L_HI(net1411));
 sg13g2_tiehi \cpu.dcache.r_dirty[1]$_SDFFCE_PP1P__1412  (.L_HI(net1412));
 sg13g2_tiehi \cpu.dcache.r_dirty[2]$_SDFFCE_PP1P__1413  (.L_HI(net1413));
 sg13g2_tiehi \cpu.dcache.r_dirty[3]$_SDFFCE_PP1P__1414  (.L_HI(net1414));
 sg13g2_tiehi \cpu.dcache.r_dirty[4]$_SDFFCE_PP1P__1415  (.L_HI(net1415));
 sg13g2_tiehi \cpu.dcache.r_dirty[5]$_SDFFCE_PP1P__1416  (.L_HI(net1416));
 sg13g2_tiehi \cpu.dcache.r_dirty[6]$_SDFFCE_PP1P__1417  (.L_HI(net1417));
 sg13g2_tiehi \cpu.dcache.r_dirty[7]$_SDFFCE_PP1P__1418  (.L_HI(net1418));
 sg13g2_tiehi \cpu.dcache.r_offset[0]$_SDFF_PN0__1419  (.L_HI(net1419));
 sg13g2_tiehi \cpu.dcache.r_offset[1]$_SDFF_PN0__1420  (.L_HI(net1420));
 sg13g2_tiehi \cpu.dcache.r_offset[2]$_SDFF_PN0__1421  (.L_HI(net1421));
 sg13g2_tiehi \cpu.dcache.r_tag[0][0]$_DFFE_PP__1422  (.L_HI(net1422));
 sg13g2_tiehi \cpu.dcache.r_tag[0][10]$_DFFE_PP__1423  (.L_HI(net1423));
 sg13g2_tiehi \cpu.dcache.r_tag[0][11]$_DFFE_PP__1424  (.L_HI(net1424));
 sg13g2_tiehi \cpu.dcache.r_tag[0][12]$_DFFE_PP__1425  (.L_HI(net1425));
 sg13g2_tiehi \cpu.dcache.r_tag[0][13]$_DFFE_PP__1426  (.L_HI(net1426));
 sg13g2_tiehi \cpu.dcache.r_tag[0][14]$_DFFE_PP__1427  (.L_HI(net1427));
 sg13g2_tiehi \cpu.dcache.r_tag[0][15]$_DFFE_PP__1428  (.L_HI(net1428));
 sg13g2_tiehi \cpu.dcache.r_tag[0][16]$_DFFE_PP__1429  (.L_HI(net1429));
 sg13g2_tiehi \cpu.dcache.r_tag[0][17]$_DFFE_PP__1430  (.L_HI(net1430));
 sg13g2_tiehi \cpu.dcache.r_tag[0][18]$_DFFE_PP__1431  (.L_HI(net1431));
 sg13g2_tiehi \cpu.dcache.r_tag[0][1]$_DFFE_PP__1432  (.L_HI(net1432));
 sg13g2_tiehi \cpu.dcache.r_tag[0][2]$_DFFE_PP__1433  (.L_HI(net1433));
 sg13g2_tiehi \cpu.dcache.r_tag[0][3]$_DFFE_PP__1434  (.L_HI(net1434));
 sg13g2_tiehi \cpu.dcache.r_tag[0][4]$_DFFE_PP__1435  (.L_HI(net1435));
 sg13g2_tiehi \cpu.dcache.r_tag[0][5]$_DFFE_PP__1436  (.L_HI(net1436));
 sg13g2_tiehi \cpu.dcache.r_tag[0][6]$_DFFE_PP__1437  (.L_HI(net1437));
 sg13g2_tiehi \cpu.dcache.r_tag[0][7]$_DFFE_PP__1438  (.L_HI(net1438));
 sg13g2_tiehi \cpu.dcache.r_tag[0][8]$_DFFE_PP__1439  (.L_HI(net1439));
 sg13g2_tiehi \cpu.dcache.r_tag[0][9]$_DFFE_PP__1440  (.L_HI(net1440));
 sg13g2_tiehi \cpu.dcache.r_tag[1][0]$_DFFE_PP__1441  (.L_HI(net1441));
 sg13g2_tiehi \cpu.dcache.r_tag[1][10]$_DFFE_PP__1442  (.L_HI(net1442));
 sg13g2_tiehi \cpu.dcache.r_tag[1][11]$_DFFE_PP__1443  (.L_HI(net1443));
 sg13g2_tiehi \cpu.dcache.r_tag[1][12]$_DFFE_PP__1444  (.L_HI(net1444));
 sg13g2_tiehi \cpu.dcache.r_tag[1][13]$_DFFE_PP__1445  (.L_HI(net1445));
 sg13g2_tiehi \cpu.dcache.r_tag[1][14]$_DFFE_PP__1446  (.L_HI(net1446));
 sg13g2_tiehi \cpu.dcache.r_tag[1][15]$_DFFE_PP__1447  (.L_HI(net1447));
 sg13g2_tiehi \cpu.dcache.r_tag[1][16]$_DFFE_PP__1448  (.L_HI(net1448));
 sg13g2_tiehi \cpu.dcache.r_tag[1][17]$_DFFE_PP__1449  (.L_HI(net1449));
 sg13g2_tiehi \cpu.dcache.r_tag[1][18]$_DFFE_PP__1450  (.L_HI(net1450));
 sg13g2_tiehi \cpu.dcache.r_tag[1][1]$_DFFE_PP__1451  (.L_HI(net1451));
 sg13g2_tiehi \cpu.dcache.r_tag[1][2]$_DFFE_PP__1452  (.L_HI(net1452));
 sg13g2_tiehi \cpu.dcache.r_tag[1][3]$_DFFE_PP__1453  (.L_HI(net1453));
 sg13g2_tiehi \cpu.dcache.r_tag[1][4]$_DFFE_PP__1454  (.L_HI(net1454));
 sg13g2_tiehi \cpu.dcache.r_tag[1][5]$_DFFE_PP__1455  (.L_HI(net1455));
 sg13g2_tiehi \cpu.dcache.r_tag[1][6]$_DFFE_PP__1456  (.L_HI(net1456));
 sg13g2_tiehi \cpu.dcache.r_tag[1][7]$_DFFE_PP__1457  (.L_HI(net1457));
 sg13g2_tiehi \cpu.dcache.r_tag[1][8]$_DFFE_PP__1458  (.L_HI(net1458));
 sg13g2_tiehi \cpu.dcache.r_tag[1][9]$_DFFE_PP__1459  (.L_HI(net1459));
 sg13g2_tiehi \cpu.dcache.r_tag[2][0]$_DFFE_PP__1460  (.L_HI(net1460));
 sg13g2_tiehi \cpu.dcache.r_tag[2][10]$_DFFE_PP__1461  (.L_HI(net1461));
 sg13g2_tiehi \cpu.dcache.r_tag[2][11]$_DFFE_PP__1462  (.L_HI(net1462));
 sg13g2_tiehi \cpu.dcache.r_tag[2][12]$_DFFE_PP__1463  (.L_HI(net1463));
 sg13g2_tiehi \cpu.dcache.r_tag[2][13]$_DFFE_PP__1464  (.L_HI(net1464));
 sg13g2_tiehi \cpu.dcache.r_tag[2][14]$_DFFE_PP__1465  (.L_HI(net1465));
 sg13g2_tiehi \cpu.dcache.r_tag[2][15]$_DFFE_PP__1466  (.L_HI(net1466));
 sg13g2_tiehi \cpu.dcache.r_tag[2][16]$_DFFE_PP__1467  (.L_HI(net1467));
 sg13g2_tiehi \cpu.dcache.r_tag[2][17]$_DFFE_PP__1468  (.L_HI(net1468));
 sg13g2_tiehi \cpu.dcache.r_tag[2][18]$_DFFE_PP__1469  (.L_HI(net1469));
 sg13g2_tiehi \cpu.dcache.r_tag[2][1]$_DFFE_PP__1470  (.L_HI(net1470));
 sg13g2_tiehi \cpu.dcache.r_tag[2][2]$_DFFE_PP__1471  (.L_HI(net1471));
 sg13g2_tiehi \cpu.dcache.r_tag[2][3]$_DFFE_PP__1472  (.L_HI(net1472));
 sg13g2_tiehi \cpu.dcache.r_tag[2][4]$_DFFE_PP__1473  (.L_HI(net1473));
 sg13g2_tiehi \cpu.dcache.r_tag[2][5]$_DFFE_PP__1474  (.L_HI(net1474));
 sg13g2_tiehi \cpu.dcache.r_tag[2][6]$_DFFE_PP__1475  (.L_HI(net1475));
 sg13g2_tiehi \cpu.dcache.r_tag[2][7]$_DFFE_PP__1476  (.L_HI(net1476));
 sg13g2_tiehi \cpu.dcache.r_tag[2][8]$_DFFE_PP__1477  (.L_HI(net1477));
 sg13g2_tiehi \cpu.dcache.r_tag[2][9]$_DFFE_PP__1478  (.L_HI(net1478));
 sg13g2_tiehi \cpu.dcache.r_tag[3][0]$_DFFE_PP__1479  (.L_HI(net1479));
 sg13g2_tiehi \cpu.dcache.r_tag[3][10]$_DFFE_PP__1480  (.L_HI(net1480));
 sg13g2_tiehi \cpu.dcache.r_tag[3][11]$_DFFE_PP__1481  (.L_HI(net1481));
 sg13g2_tiehi \cpu.dcache.r_tag[3][12]$_DFFE_PP__1482  (.L_HI(net1482));
 sg13g2_tiehi \cpu.dcache.r_tag[3][13]$_DFFE_PP__1483  (.L_HI(net1483));
 sg13g2_tiehi \cpu.dcache.r_tag[3][14]$_DFFE_PP__1484  (.L_HI(net1484));
 sg13g2_tiehi \cpu.dcache.r_tag[3][15]$_DFFE_PP__1485  (.L_HI(net1485));
 sg13g2_tiehi \cpu.dcache.r_tag[3][16]$_DFFE_PP__1486  (.L_HI(net1486));
 sg13g2_tiehi \cpu.dcache.r_tag[3][17]$_DFFE_PP__1487  (.L_HI(net1487));
 sg13g2_tiehi \cpu.dcache.r_tag[3][18]$_DFFE_PP__1488  (.L_HI(net1488));
 sg13g2_tiehi \cpu.dcache.r_tag[3][1]$_DFFE_PP__1489  (.L_HI(net1489));
 sg13g2_tiehi \cpu.dcache.r_tag[3][2]$_DFFE_PP__1490  (.L_HI(net1490));
 sg13g2_tiehi \cpu.dcache.r_tag[3][3]$_DFFE_PP__1491  (.L_HI(net1491));
 sg13g2_tiehi \cpu.dcache.r_tag[3][4]$_DFFE_PP__1492  (.L_HI(net1492));
 sg13g2_tiehi \cpu.dcache.r_tag[3][5]$_DFFE_PP__1493  (.L_HI(net1493));
 sg13g2_tiehi \cpu.dcache.r_tag[3][6]$_DFFE_PP__1494  (.L_HI(net1494));
 sg13g2_tiehi \cpu.dcache.r_tag[3][7]$_DFFE_PP__1495  (.L_HI(net1495));
 sg13g2_tiehi \cpu.dcache.r_tag[3][8]$_DFFE_PP__1496  (.L_HI(net1496));
 sg13g2_tiehi \cpu.dcache.r_tag[3][9]$_DFFE_PP__1497  (.L_HI(net1497));
 sg13g2_tiehi \cpu.dcache.r_tag[4][0]$_DFFE_PP__1498  (.L_HI(net1498));
 sg13g2_tiehi \cpu.dcache.r_tag[4][10]$_DFFE_PP__1499  (.L_HI(net1499));
 sg13g2_tiehi \cpu.dcache.r_tag[4][11]$_DFFE_PP__1500  (.L_HI(net1500));
 sg13g2_tiehi \cpu.dcache.r_tag[4][12]$_DFFE_PP__1501  (.L_HI(net1501));
 sg13g2_tiehi \cpu.dcache.r_tag[4][13]$_DFFE_PP__1502  (.L_HI(net1502));
 sg13g2_tiehi \cpu.dcache.r_tag[4][14]$_DFFE_PP__1503  (.L_HI(net1503));
 sg13g2_tiehi \cpu.dcache.r_tag[4][15]$_DFFE_PP__1504  (.L_HI(net1504));
 sg13g2_tiehi \cpu.dcache.r_tag[4][16]$_DFFE_PP__1505  (.L_HI(net1505));
 sg13g2_tiehi \cpu.dcache.r_tag[4][17]$_DFFE_PP__1506  (.L_HI(net1506));
 sg13g2_tiehi \cpu.dcache.r_tag[4][18]$_DFFE_PP__1507  (.L_HI(net1507));
 sg13g2_tiehi \cpu.dcache.r_tag[4][1]$_DFFE_PP__1508  (.L_HI(net1508));
 sg13g2_tiehi \cpu.dcache.r_tag[4][2]$_DFFE_PP__1509  (.L_HI(net1509));
 sg13g2_tiehi \cpu.dcache.r_tag[4][3]$_DFFE_PP__1510  (.L_HI(net1510));
 sg13g2_tiehi \cpu.dcache.r_tag[4][4]$_DFFE_PP__1511  (.L_HI(net1511));
 sg13g2_tiehi \cpu.dcache.r_tag[4][5]$_DFFE_PP__1512  (.L_HI(net1512));
 sg13g2_tiehi \cpu.dcache.r_tag[4][6]$_DFFE_PP__1513  (.L_HI(net1513));
 sg13g2_tiehi \cpu.dcache.r_tag[4][7]$_DFFE_PP__1514  (.L_HI(net1514));
 sg13g2_tiehi \cpu.dcache.r_tag[4][8]$_DFFE_PP__1515  (.L_HI(net1515));
 sg13g2_tiehi \cpu.dcache.r_tag[4][9]$_DFFE_PP__1516  (.L_HI(net1516));
 sg13g2_tiehi \cpu.dcache.r_tag[5][0]$_DFFE_PP__1517  (.L_HI(net1517));
 sg13g2_tiehi \cpu.dcache.r_tag[5][10]$_DFFE_PP__1518  (.L_HI(net1518));
 sg13g2_tiehi \cpu.dcache.r_tag[5][11]$_DFFE_PP__1519  (.L_HI(net1519));
 sg13g2_tiehi \cpu.dcache.r_tag[5][12]$_DFFE_PP__1520  (.L_HI(net1520));
 sg13g2_tiehi \cpu.dcache.r_tag[5][13]$_DFFE_PP__1521  (.L_HI(net1521));
 sg13g2_tiehi \cpu.dcache.r_tag[5][14]$_DFFE_PP__1522  (.L_HI(net1522));
 sg13g2_tiehi \cpu.dcache.r_tag[5][15]$_DFFE_PP__1523  (.L_HI(net1523));
 sg13g2_tiehi \cpu.dcache.r_tag[5][16]$_DFFE_PP__1524  (.L_HI(net1524));
 sg13g2_tiehi \cpu.dcache.r_tag[5][17]$_DFFE_PP__1525  (.L_HI(net1525));
 sg13g2_tiehi \cpu.dcache.r_tag[5][18]$_DFFE_PP__1526  (.L_HI(net1526));
 sg13g2_tiehi \cpu.dcache.r_tag[5][1]$_DFFE_PP__1527  (.L_HI(net1527));
 sg13g2_tiehi \cpu.dcache.r_tag[5][2]$_DFFE_PP__1528  (.L_HI(net1528));
 sg13g2_tiehi \cpu.dcache.r_tag[5][3]$_DFFE_PP__1529  (.L_HI(net1529));
 sg13g2_tiehi \cpu.dcache.r_tag[5][4]$_DFFE_PP__1530  (.L_HI(net1530));
 sg13g2_tiehi \cpu.dcache.r_tag[5][5]$_DFFE_PP__1531  (.L_HI(net1531));
 sg13g2_tiehi \cpu.dcache.r_tag[5][6]$_DFFE_PP__1532  (.L_HI(net1532));
 sg13g2_tiehi \cpu.dcache.r_tag[5][7]$_DFFE_PP__1533  (.L_HI(net1533));
 sg13g2_tiehi \cpu.dcache.r_tag[5][8]$_DFFE_PP__1534  (.L_HI(net1534));
 sg13g2_tiehi \cpu.dcache.r_tag[5][9]$_DFFE_PP__1535  (.L_HI(net1535));
 sg13g2_tiehi \cpu.dcache.r_tag[6][0]$_DFFE_PP__1536  (.L_HI(net1536));
 sg13g2_tiehi \cpu.dcache.r_tag[6][10]$_DFFE_PP__1537  (.L_HI(net1537));
 sg13g2_tiehi \cpu.dcache.r_tag[6][11]$_DFFE_PP__1538  (.L_HI(net1538));
 sg13g2_tiehi \cpu.dcache.r_tag[6][12]$_DFFE_PP__1539  (.L_HI(net1539));
 sg13g2_tiehi \cpu.dcache.r_tag[6][13]$_DFFE_PP__1540  (.L_HI(net1540));
 sg13g2_tiehi \cpu.dcache.r_tag[6][14]$_DFFE_PP__1541  (.L_HI(net1541));
 sg13g2_tiehi \cpu.dcache.r_tag[6][15]$_DFFE_PP__1542  (.L_HI(net1542));
 sg13g2_tiehi \cpu.dcache.r_tag[6][16]$_DFFE_PP__1543  (.L_HI(net1543));
 sg13g2_tiehi \cpu.dcache.r_tag[6][17]$_DFFE_PP__1544  (.L_HI(net1544));
 sg13g2_tiehi \cpu.dcache.r_tag[6][18]$_DFFE_PP__1545  (.L_HI(net1545));
 sg13g2_tiehi \cpu.dcache.r_tag[6][1]$_DFFE_PP__1546  (.L_HI(net1546));
 sg13g2_tiehi \cpu.dcache.r_tag[6][2]$_DFFE_PP__1547  (.L_HI(net1547));
 sg13g2_tiehi \cpu.dcache.r_tag[6][3]$_DFFE_PP__1548  (.L_HI(net1548));
 sg13g2_tiehi \cpu.dcache.r_tag[6][4]$_DFFE_PP__1549  (.L_HI(net1549));
 sg13g2_tiehi \cpu.dcache.r_tag[6][5]$_DFFE_PP__1550  (.L_HI(net1550));
 sg13g2_tiehi \cpu.dcache.r_tag[6][6]$_DFFE_PP__1551  (.L_HI(net1551));
 sg13g2_tiehi \cpu.dcache.r_tag[6][7]$_DFFE_PP__1552  (.L_HI(net1552));
 sg13g2_tiehi \cpu.dcache.r_tag[6][8]$_DFFE_PP__1553  (.L_HI(net1553));
 sg13g2_tiehi \cpu.dcache.r_tag[6][9]$_DFFE_PP__1554  (.L_HI(net1554));
 sg13g2_tiehi \cpu.dcache.r_tag[7][0]$_DFFE_PP__1555  (.L_HI(net1555));
 sg13g2_tiehi \cpu.dcache.r_tag[7][10]$_DFFE_PP__1556  (.L_HI(net1556));
 sg13g2_tiehi \cpu.dcache.r_tag[7][11]$_DFFE_PP__1557  (.L_HI(net1557));
 sg13g2_tiehi \cpu.dcache.r_tag[7][12]$_DFFE_PP__1558  (.L_HI(net1558));
 sg13g2_tiehi \cpu.dcache.r_tag[7][13]$_DFFE_PP__1559  (.L_HI(net1559));
 sg13g2_tiehi \cpu.dcache.r_tag[7][14]$_DFFE_PP__1560  (.L_HI(net1560));
 sg13g2_tiehi \cpu.dcache.r_tag[7][15]$_DFFE_PP__1561  (.L_HI(net1561));
 sg13g2_tiehi \cpu.dcache.r_tag[7][16]$_DFFE_PP__1562  (.L_HI(net1562));
 sg13g2_tiehi \cpu.dcache.r_tag[7][17]$_DFFE_PP__1563  (.L_HI(net1563));
 sg13g2_tiehi \cpu.dcache.r_tag[7][18]$_DFFE_PP__1564  (.L_HI(net1564));
 sg13g2_tiehi \cpu.dcache.r_tag[7][1]$_DFFE_PP__1565  (.L_HI(net1565));
 sg13g2_tiehi \cpu.dcache.r_tag[7][2]$_DFFE_PP__1566  (.L_HI(net1566));
 sg13g2_tiehi \cpu.dcache.r_tag[7][3]$_DFFE_PP__1567  (.L_HI(net1567));
 sg13g2_tiehi \cpu.dcache.r_tag[7][4]$_DFFE_PP__1568  (.L_HI(net1568));
 sg13g2_tiehi \cpu.dcache.r_tag[7][5]$_DFFE_PP__1569  (.L_HI(net1569));
 sg13g2_tiehi \cpu.dcache.r_tag[7][6]$_DFFE_PP__1570  (.L_HI(net1570));
 sg13g2_tiehi \cpu.dcache.r_tag[7][7]$_DFFE_PP__1571  (.L_HI(net1571));
 sg13g2_tiehi \cpu.dcache.r_tag[7][8]$_DFFE_PP__1572  (.L_HI(net1572));
 sg13g2_tiehi \cpu.dcache.r_tag[7][9]$_DFFE_PP__1573  (.L_HI(net1573));
 sg13g2_tiehi \cpu.dcache.r_valid[0]$_SDFFE_PP0P__1574  (.L_HI(net1574));
 sg13g2_tiehi \cpu.dcache.r_valid[1]$_SDFFE_PP0P__1575  (.L_HI(net1575));
 sg13g2_tiehi \cpu.dcache.r_valid[2]$_SDFFE_PP0P__1576  (.L_HI(net1576));
 sg13g2_tiehi \cpu.dcache.r_valid[3]$_SDFFE_PP0P__1577  (.L_HI(net1577));
 sg13g2_tiehi \cpu.dcache.r_valid[4]$_SDFFE_PP0P__1578  (.L_HI(net1578));
 sg13g2_tiehi \cpu.dcache.r_valid[5]$_SDFFE_PP0P__1579  (.L_HI(net1579));
 sg13g2_tiehi \cpu.dcache.r_valid[6]$_SDFFE_PP0P__1580  (.L_HI(net1580));
 sg13g2_tiehi \cpu.dcache.r_valid[7]$_SDFFE_PP0P__1581  (.L_HI(net1581));
 sg13g2_tiehi \cpu.dec.r_br$_DFFE_PP__1582  (.L_HI(net1582));
 sg13g2_tiehi \cpu.dec.r_cond[0]$_DFFE_PP__1583  (.L_HI(net1583));
 sg13g2_tiehi \cpu.dec.r_cond[1]$_DFFE_PP__1584  (.L_HI(net1584));
 sg13g2_tiehi \cpu.dec.r_cond[2]$_DFFE_PP__1585  (.L_HI(net1585));
 sg13g2_tiehi \cpu.dec.r_div$_DFFE_PP__1586  (.L_HI(net1586));
 sg13g2_tiehi \cpu.dec.r_flush_all$_DFFE_PP__1587  (.L_HI(net1587));
 sg13g2_tiehi \cpu.dec.r_flush_write$_DFFE_PP__1588  (.L_HI(net1588));
 sg13g2_tiehi \cpu.dec.r_imm[0]$_DFFE_PP__1589  (.L_HI(net1589));
 sg13g2_tiehi \cpu.dec.r_imm[10]$_DFFE_PP__1590  (.L_HI(net1590));
 sg13g2_tiehi \cpu.dec.r_imm[11]$_DFFE_PP__1591  (.L_HI(net1591));
 sg13g2_tiehi \cpu.dec.r_imm[12]$_DFFE_PP__1592  (.L_HI(net1592));
 sg13g2_tiehi \cpu.dec.r_imm[13]$_DFFE_PP__1593  (.L_HI(net1593));
 sg13g2_tiehi \cpu.dec.r_imm[14]$_DFFE_PP__1594  (.L_HI(net1594));
 sg13g2_tiehi \cpu.dec.r_imm[15]$_DFFE_PP__1595  (.L_HI(net1595));
 sg13g2_tiehi \cpu.dec.r_imm[1]$_DFFE_PP__1596  (.L_HI(net1596));
 sg13g2_tiehi \cpu.dec.r_imm[2]$_DFFE_PP__1597  (.L_HI(net1597));
 sg13g2_tiehi \cpu.dec.r_imm[3]$_DFFE_PP__1598  (.L_HI(net1598));
 sg13g2_tiehi \cpu.dec.r_imm[4]$_DFFE_PP__1599  (.L_HI(net1599));
 sg13g2_tiehi \cpu.dec.r_imm[5]$_DFFE_PP__1600  (.L_HI(net1600));
 sg13g2_tiehi \cpu.dec.r_imm[6]$_DFFE_PP__1601  (.L_HI(net1601));
 sg13g2_tiehi \cpu.dec.r_imm[7]$_DFFE_PP__1602  (.L_HI(net1602));
 sg13g2_tiehi \cpu.dec.r_imm[8]$_DFFE_PP__1603  (.L_HI(net1603));
 sg13g2_tiehi \cpu.dec.r_imm[9]$_DFFE_PP__1604  (.L_HI(net1604));
 sg13g2_tiehi \cpu.dec.r_inv_mmu$_DFFE_PP__1605  (.L_HI(net1605));
 sg13g2_tiehi \cpu.dec.r_io$_DFFE_PP__1606  (.L_HI(net1606));
 sg13g2_tiehi \cpu.dec.r_jmp$_SDFFCE_PP0P__1607  (.L_HI(net1607));
 sg13g2_tiehi \cpu.dec.r_load$_DFFE_PP__1608  (.L_HI(net1608));
 sg13g2_tiehi \cpu.dec.r_mult$_DFFE_PP__1609  (.L_HI(net1609));
 sg13g2_tiehi \cpu.dec.r_needs_rs2$_DFFE_PP__1610  (.L_HI(net1610));
 sg13g2_tiehi \cpu.dec.r_op[10]$_DFF_P__1611  (.L_HI(net1611));
 sg13g2_tiehi \cpu.dec.r_op[1]$_DFF_P__1612  (.L_HI(net1612));
 sg13g2_tiehi \cpu.dec.r_op[2]$_DFF_P__1613  (.L_HI(net1613));
 sg13g2_tiehi \cpu.dec.r_op[3]$_DFF_P__1614  (.L_HI(net1614));
 sg13g2_tiehi \cpu.dec.r_op[4]$_DFF_P__1615  (.L_HI(net1615));
 sg13g2_tiehi \cpu.dec.r_op[5]$_DFF_P__1616  (.L_HI(net1616));
 sg13g2_tiehi \cpu.dec.r_op[6]$_DFF_P__1617  (.L_HI(net1617));
 sg13g2_tiehi \cpu.dec.r_op[7]$_DFF_P__1618  (.L_HI(net1618));
 sg13g2_tiehi \cpu.dec.r_op[8]$_DFF_P__1619  (.L_HI(net1619));
 sg13g2_tiehi \cpu.dec.r_op[9]$_DFF_P__1620  (.L_HI(net1620));
 sg13g2_tiehi \cpu.dec.r_rd[0]$_DFFE_PP__1621  (.L_HI(net1621));
 sg13g2_tiehi \cpu.dec.r_rd[1]$_DFFE_PP__1622  (.L_HI(net1622));
 sg13g2_tiehi \cpu.dec.r_rd[2]$_DFFE_PP__1623  (.L_HI(net1623));
 sg13g2_tiehi \cpu.dec.r_rd[3]$_DFFE_PP__1624  (.L_HI(net1624));
 sg13g2_tiehi \cpu.dec.r_ready$_DFF_P__1625  (.L_HI(net1625));
 sg13g2_tiehi \cpu.dec.r_rs1[0]$_DFFE_PP__1626  (.L_HI(net1626));
 sg13g2_tiehi \cpu.dec.r_rs1[1]$_DFFE_PP__1627  (.L_HI(net1627));
 sg13g2_tiehi \cpu.dec.r_rs1[2]$_DFFE_PP__1628  (.L_HI(net1628));
 sg13g2_tiehi \cpu.dec.r_rs1[3]$_DFFE_PP__1629  (.L_HI(net1629));
 sg13g2_tiehi \cpu.dec.r_rs2[0]$_DFFE_PP__1630  (.L_HI(net1630));
 sg13g2_tiehi \cpu.dec.r_rs2[1]$_DFFE_PP__1631  (.L_HI(net1631));
 sg13g2_tiehi \cpu.dec.r_rs2[2]$_DFFE_PP__1632  (.L_HI(net1632));
 sg13g2_tiehi \cpu.dec.r_rs2[3]$_DFFE_PP__1633  (.L_HI(net1633));
 sg13g2_tiehi \cpu.dec.r_rs2_pc$_DFFE_PP__1634  (.L_HI(net1634));
 sg13g2_tiehi \cpu.dec.r_set_cc$_SDFFCE_PP0P__1635  (.L_HI(net1635));
 sg13g2_tiehi \cpu.dec.r_store$_DFFE_PP__1636  (.L_HI(net1636));
 sg13g2_tiehi \cpu.dec.r_swapsp$_DFFE_PP__1637  (.L_HI(net1637));
 sg13g2_tiehi \cpu.dec.r_sys_call$_DFFE_PP__1638  (.L_HI(net1638));
 sg13g2_tiehi \cpu.dec.r_trap$_DFFE_PP__1639  (.L_HI(net1639));
 sg13g2_tiehi \cpu.ex.genblk3.r_mmu_d_proxy$_SDFFE_PP0P__1640  (.L_HI(net1640));
 sg13g2_tiehi \cpu.ex.genblk3.r_mmu_enable$_SDFFE_PN0P__1641  (.L_HI(net1641));
 sg13g2_tiehi \cpu.ex.genblk3.r_prev_supmode$_SDFFE_PN1P__1642  (.L_HI(net1642));
 sg13g2_tiehi \cpu.ex.genblk3.r_supmode$_DFF_P__1643  (.L_HI(net1643));
 sg13g2_tiehi \cpu.ex.genblk3.r_user_io$_SDFFE_PN0P__1644  (.L_HI(net1644));
 sg13g2_tiehi \cpu.ex.r_10[0]$_DFFE_PP__1645  (.L_HI(net1645));
 sg13g2_tiehi \cpu.ex.r_10[10]$_DFFE_PP__1646  (.L_HI(net1646));
 sg13g2_tiehi \cpu.ex.r_10[11]$_DFFE_PP__1647  (.L_HI(net1647));
 sg13g2_tiehi \cpu.ex.r_10[12]$_DFFE_PP__1648  (.L_HI(net1648));
 sg13g2_tiehi \cpu.ex.r_10[13]$_DFFE_PP__1649  (.L_HI(net1649));
 sg13g2_tiehi \cpu.ex.r_10[14]$_DFFE_PP__1650  (.L_HI(net1650));
 sg13g2_tiehi \cpu.ex.r_10[15]$_DFFE_PP__1651  (.L_HI(net1651));
 sg13g2_tiehi \cpu.ex.r_10[1]$_DFFE_PP__1652  (.L_HI(net1652));
 sg13g2_tiehi \cpu.ex.r_10[2]$_DFFE_PP__1653  (.L_HI(net1653));
 sg13g2_tiehi \cpu.ex.r_10[3]$_DFFE_PP__1654  (.L_HI(net1654));
 sg13g2_tiehi \cpu.ex.r_10[4]$_DFFE_PP__1655  (.L_HI(net1655));
 sg13g2_tiehi \cpu.ex.r_10[5]$_DFFE_PP__1656  (.L_HI(net1656));
 sg13g2_tiehi \cpu.ex.r_10[6]$_DFFE_PP__1657  (.L_HI(net1657));
 sg13g2_tiehi \cpu.ex.r_10[7]$_DFFE_PP__1658  (.L_HI(net1658));
 sg13g2_tiehi \cpu.ex.r_10[8]$_DFFE_PP__1659  (.L_HI(net1659));
 sg13g2_tiehi \cpu.ex.r_10[9]$_DFFE_PP__1660  (.L_HI(net1660));
 sg13g2_tiehi \cpu.ex.r_11[0]$_DFFE_PP__1661  (.L_HI(net1661));
 sg13g2_tiehi \cpu.ex.r_11[10]$_DFFE_PP__1662  (.L_HI(net1662));
 sg13g2_tiehi \cpu.ex.r_11[11]$_DFFE_PP__1663  (.L_HI(net1663));
 sg13g2_tiehi \cpu.ex.r_11[12]$_DFFE_PP__1664  (.L_HI(net1664));
 sg13g2_tiehi \cpu.ex.r_11[13]$_DFFE_PP__1665  (.L_HI(net1665));
 sg13g2_tiehi \cpu.ex.r_11[14]$_DFFE_PP__1666  (.L_HI(net1666));
 sg13g2_tiehi \cpu.ex.r_11[15]$_DFFE_PP__1667  (.L_HI(net1667));
 sg13g2_tiehi \cpu.ex.r_11[1]$_DFFE_PP__1668  (.L_HI(net1668));
 sg13g2_tiehi \cpu.ex.r_11[2]$_DFFE_PP__1669  (.L_HI(net1669));
 sg13g2_tiehi \cpu.ex.r_11[3]$_DFFE_PP__1670  (.L_HI(net1670));
 sg13g2_tiehi \cpu.ex.r_11[4]$_DFFE_PP__1671  (.L_HI(net1671));
 sg13g2_tiehi \cpu.ex.r_11[5]$_DFFE_PP__1672  (.L_HI(net1672));
 sg13g2_tiehi \cpu.ex.r_11[6]$_DFFE_PP__1673  (.L_HI(net1673));
 sg13g2_tiehi \cpu.ex.r_11[7]$_DFFE_PP__1674  (.L_HI(net1674));
 sg13g2_tiehi \cpu.ex.r_11[8]$_DFFE_PP__1675  (.L_HI(net1675));
 sg13g2_tiehi \cpu.ex.r_11[9]$_DFFE_PP__1676  (.L_HI(net1676));
 sg13g2_tiehi \cpu.ex.r_12[0]$_DFFE_PP__1677  (.L_HI(net1677));
 sg13g2_tiehi \cpu.ex.r_12[10]$_DFFE_PP__1678  (.L_HI(net1678));
 sg13g2_tiehi \cpu.ex.r_12[11]$_DFFE_PP__1679  (.L_HI(net1679));
 sg13g2_tiehi \cpu.ex.r_12[12]$_DFFE_PP__1680  (.L_HI(net1680));
 sg13g2_tiehi \cpu.ex.r_12[13]$_DFFE_PP__1681  (.L_HI(net1681));
 sg13g2_tiehi \cpu.ex.r_12[14]$_DFFE_PP__1682  (.L_HI(net1682));
 sg13g2_tiehi \cpu.ex.r_12[15]$_DFFE_PP__1683  (.L_HI(net1683));
 sg13g2_tiehi \cpu.ex.r_12[1]$_DFFE_PP__1684  (.L_HI(net1684));
 sg13g2_tiehi \cpu.ex.r_12[2]$_DFFE_PP__1685  (.L_HI(net1685));
 sg13g2_tiehi \cpu.ex.r_12[3]$_DFFE_PP__1686  (.L_HI(net1686));
 sg13g2_tiehi \cpu.ex.r_12[4]$_DFFE_PP__1687  (.L_HI(net1687));
 sg13g2_tiehi \cpu.ex.r_12[5]$_DFFE_PP__1688  (.L_HI(net1688));
 sg13g2_tiehi \cpu.ex.r_12[6]$_DFFE_PP__1689  (.L_HI(net1689));
 sg13g2_tiehi \cpu.ex.r_12[7]$_DFFE_PP__1690  (.L_HI(net1690));
 sg13g2_tiehi \cpu.ex.r_12[8]$_DFFE_PP__1691  (.L_HI(net1691));
 sg13g2_tiehi \cpu.ex.r_12[9]$_DFFE_PP__1692  (.L_HI(net1692));
 sg13g2_tiehi \cpu.ex.r_13[0]$_DFFE_PP__1693  (.L_HI(net1693));
 sg13g2_tiehi \cpu.ex.r_13[10]$_DFFE_PP__1694  (.L_HI(net1694));
 sg13g2_tiehi \cpu.ex.r_13[11]$_DFFE_PP__1695  (.L_HI(net1695));
 sg13g2_tiehi \cpu.ex.r_13[12]$_DFFE_PP__1696  (.L_HI(net1696));
 sg13g2_tiehi \cpu.ex.r_13[13]$_DFFE_PP__1697  (.L_HI(net1697));
 sg13g2_tiehi \cpu.ex.r_13[14]$_DFFE_PP__1698  (.L_HI(net1698));
 sg13g2_tiehi \cpu.ex.r_13[15]$_DFFE_PP__1699  (.L_HI(net1699));
 sg13g2_tiehi \cpu.ex.r_13[1]$_DFFE_PP__1700  (.L_HI(net1700));
 sg13g2_tiehi \cpu.ex.r_13[2]$_DFFE_PP__1701  (.L_HI(net1701));
 sg13g2_tiehi \cpu.ex.r_13[3]$_DFFE_PP__1702  (.L_HI(net1702));
 sg13g2_tiehi \cpu.ex.r_13[4]$_DFFE_PP__1703  (.L_HI(net1703));
 sg13g2_tiehi \cpu.ex.r_13[5]$_DFFE_PP__1704  (.L_HI(net1704));
 sg13g2_tiehi \cpu.ex.r_13[6]$_DFFE_PP__1705  (.L_HI(net1705));
 sg13g2_tiehi \cpu.ex.r_13[7]$_DFFE_PP__1706  (.L_HI(net1706));
 sg13g2_tiehi \cpu.ex.r_13[8]$_DFFE_PP__1707  (.L_HI(net1707));
 sg13g2_tiehi \cpu.ex.r_13[9]$_DFFE_PP__1708  (.L_HI(net1708));
 sg13g2_tiehi \cpu.ex.r_14[0]$_DFFE_PP__1709  (.L_HI(net1709));
 sg13g2_tiehi \cpu.ex.r_14[10]$_DFFE_PP__1710  (.L_HI(net1710));
 sg13g2_tiehi \cpu.ex.r_14[11]$_DFFE_PP__1711  (.L_HI(net1711));
 sg13g2_tiehi \cpu.ex.r_14[12]$_DFFE_PP__1712  (.L_HI(net1712));
 sg13g2_tiehi \cpu.ex.r_14[13]$_DFFE_PP__1713  (.L_HI(net1713));
 sg13g2_tiehi \cpu.ex.r_14[14]$_DFFE_PP__1714  (.L_HI(net1714));
 sg13g2_tiehi \cpu.ex.r_14[15]$_DFFE_PP__1715  (.L_HI(net1715));
 sg13g2_tiehi \cpu.ex.r_14[1]$_DFFE_PP__1716  (.L_HI(net1716));
 sg13g2_tiehi \cpu.ex.r_14[2]$_DFFE_PP__1717  (.L_HI(net1717));
 sg13g2_tiehi \cpu.ex.r_14[3]$_DFFE_PP__1718  (.L_HI(net1718));
 sg13g2_tiehi \cpu.ex.r_14[4]$_DFFE_PP__1719  (.L_HI(net1719));
 sg13g2_tiehi \cpu.ex.r_14[5]$_DFFE_PP__1720  (.L_HI(net1720));
 sg13g2_tiehi \cpu.ex.r_14[6]$_DFFE_PP__1721  (.L_HI(net1721));
 sg13g2_tiehi \cpu.ex.r_14[7]$_DFFE_PP__1722  (.L_HI(net1722));
 sg13g2_tiehi \cpu.ex.r_14[8]$_DFFE_PP__1723  (.L_HI(net1723));
 sg13g2_tiehi \cpu.ex.r_14[9]$_DFFE_PP__1724  (.L_HI(net1724));
 sg13g2_tiehi \cpu.ex.r_15[0]$_DFFE_PP__1725  (.L_HI(net1725));
 sg13g2_tiehi \cpu.ex.r_15[10]$_DFFE_PP__1726  (.L_HI(net1726));
 sg13g2_tiehi \cpu.ex.r_15[11]$_DFFE_PP__1727  (.L_HI(net1727));
 sg13g2_tiehi \cpu.ex.r_15[12]$_DFFE_PP__1728  (.L_HI(net1728));
 sg13g2_tiehi \cpu.ex.r_15[13]$_DFFE_PP__1729  (.L_HI(net1729));
 sg13g2_tiehi \cpu.ex.r_15[14]$_DFFE_PP__1730  (.L_HI(net1730));
 sg13g2_tiehi \cpu.ex.r_15[15]$_DFFE_PP__1731  (.L_HI(net1731));
 sg13g2_tiehi \cpu.ex.r_15[1]$_DFFE_PP__1732  (.L_HI(net1732));
 sg13g2_tiehi \cpu.ex.r_15[2]$_DFFE_PP__1733  (.L_HI(net1733));
 sg13g2_tiehi \cpu.ex.r_15[3]$_DFFE_PP__1734  (.L_HI(net1734));
 sg13g2_tiehi \cpu.ex.r_15[4]$_DFFE_PP__1735  (.L_HI(net1735));
 sg13g2_tiehi \cpu.ex.r_15[5]$_DFFE_PP__1736  (.L_HI(net1736));
 sg13g2_tiehi \cpu.ex.r_15[6]$_DFFE_PP__1737  (.L_HI(net1737));
 sg13g2_tiehi \cpu.ex.r_15[7]$_DFFE_PP__1738  (.L_HI(net1738));
 sg13g2_tiehi \cpu.ex.r_15[8]$_DFFE_PP__1739  (.L_HI(net1739));
 sg13g2_tiehi \cpu.ex.r_15[9]$_DFFE_PP__1740  (.L_HI(net1740));
 sg13g2_tiehi \cpu.ex.r_8[0]$_DFFE_PP__1741  (.L_HI(net1741));
 sg13g2_tiehi \cpu.ex.r_8[10]$_DFFE_PP__1742  (.L_HI(net1742));
 sg13g2_tiehi \cpu.ex.r_8[11]$_DFFE_PP__1743  (.L_HI(net1743));
 sg13g2_tiehi \cpu.ex.r_8[12]$_DFFE_PP__1744  (.L_HI(net1744));
 sg13g2_tiehi \cpu.ex.r_8[13]$_DFFE_PP__1745  (.L_HI(net1745));
 sg13g2_tiehi \cpu.ex.r_8[14]$_DFFE_PP__1746  (.L_HI(net1746));
 sg13g2_tiehi \cpu.ex.r_8[15]$_DFFE_PP__1747  (.L_HI(net1747));
 sg13g2_tiehi \cpu.ex.r_8[1]$_DFFE_PP__1748  (.L_HI(net1748));
 sg13g2_tiehi \cpu.ex.r_8[2]$_DFFE_PP__1749  (.L_HI(net1749));
 sg13g2_tiehi \cpu.ex.r_8[3]$_DFFE_PP__1750  (.L_HI(net1750));
 sg13g2_tiehi \cpu.ex.r_8[4]$_DFFE_PP__1751  (.L_HI(net1751));
 sg13g2_tiehi \cpu.ex.r_8[5]$_DFFE_PP__1752  (.L_HI(net1752));
 sg13g2_tiehi \cpu.ex.r_8[6]$_DFFE_PP__1753  (.L_HI(net1753));
 sg13g2_tiehi \cpu.ex.r_8[7]$_DFFE_PP__1754  (.L_HI(net1754));
 sg13g2_tiehi \cpu.ex.r_8[8]$_DFFE_PP__1755  (.L_HI(net1755));
 sg13g2_tiehi \cpu.ex.r_8[9]$_DFFE_PP__1756  (.L_HI(net1756));
 sg13g2_tiehi \cpu.ex.r_9[0]$_DFFE_PP__1757  (.L_HI(net1757));
 sg13g2_tiehi \cpu.ex.r_9[10]$_DFFE_PP__1758  (.L_HI(net1758));
 sg13g2_tiehi \cpu.ex.r_9[11]$_DFFE_PP__1759  (.L_HI(net1759));
 sg13g2_tiehi \cpu.ex.r_9[12]$_DFFE_PP__1760  (.L_HI(net1760));
 sg13g2_tiehi \cpu.ex.r_9[13]$_DFFE_PP__1761  (.L_HI(net1761));
 sg13g2_tiehi \cpu.ex.r_9[14]$_DFFE_PP__1762  (.L_HI(net1762));
 sg13g2_tiehi \cpu.ex.r_9[15]$_DFFE_PP__1763  (.L_HI(net1763));
 sg13g2_tiehi \cpu.ex.r_9[1]$_DFFE_PP__1764  (.L_HI(net1764));
 sg13g2_tiehi \cpu.ex.r_9[2]$_DFFE_PP__1765  (.L_HI(net1765));
 sg13g2_tiehi \cpu.ex.r_9[3]$_DFFE_PP__1766  (.L_HI(net1766));
 sg13g2_tiehi \cpu.ex.r_9[4]$_DFFE_PP__1767  (.L_HI(net1767));
 sg13g2_tiehi \cpu.ex.r_9[5]$_DFFE_PP__1768  (.L_HI(net1768));
 sg13g2_tiehi \cpu.ex.r_9[6]$_DFFE_PP__1769  (.L_HI(net1769));
 sg13g2_tiehi \cpu.ex.r_9[7]$_DFFE_PP__1770  (.L_HI(net1770));
 sg13g2_tiehi \cpu.ex.r_9[8]$_DFFE_PP__1771  (.L_HI(net1771));
 sg13g2_tiehi \cpu.ex.r_9[9]$_DFFE_PP__1772  (.L_HI(net1772));
 sg13g2_tiehi \cpu.ex.r_branch_stall$_DFF_P__1773  (.L_HI(net1773));
 sg13g2_tiehi \cpu.ex.r_cc$_DFFE_PP__1774  (.L_HI(net1774));
 sg13g2_tiehi \cpu.ex.r_d_flush_all$_SDFF_PP0__1775  (.L_HI(net1775));
 sg13g2_tiehi \cpu.ex.r_div_running$_DFF_P__1776  (.L_HI(net1776));
 sg13g2_tiehi \cpu.ex.r_epc[0]$_DFFE_PP__1777  (.L_HI(net1777));
 sg13g2_tiehi \cpu.ex.r_epc[10]$_DFFE_PP__1778  (.L_HI(net1778));
 sg13g2_tiehi \cpu.ex.r_epc[11]$_DFFE_PP__1779  (.L_HI(net1779));
 sg13g2_tiehi \cpu.ex.r_epc[12]$_DFFE_PP__1780  (.L_HI(net1780));
 sg13g2_tiehi \cpu.ex.r_epc[13]$_DFFE_PP__1781  (.L_HI(net1781));
 sg13g2_tiehi \cpu.ex.r_epc[14]$_DFFE_PP__1782  (.L_HI(net1782));
 sg13g2_tiehi \cpu.ex.r_epc[1]$_DFFE_PP__1783  (.L_HI(net1783));
 sg13g2_tiehi \cpu.ex.r_epc[2]$_DFFE_PP__1784  (.L_HI(net1784));
 sg13g2_tiehi \cpu.ex.r_epc[3]$_DFFE_PP__1785  (.L_HI(net1785));
 sg13g2_tiehi \cpu.ex.r_epc[4]$_DFFE_PP__1786  (.L_HI(net1786));
 sg13g2_tiehi \cpu.ex.r_epc[5]$_DFFE_PP__1787  (.L_HI(net1787));
 sg13g2_tiehi \cpu.ex.r_epc[6]$_DFFE_PP__1788  (.L_HI(net1788));
 sg13g2_tiehi \cpu.ex.r_epc[7]$_DFFE_PP__1789  (.L_HI(net1789));
 sg13g2_tiehi \cpu.ex.r_epc[8]$_DFFE_PP__1790  (.L_HI(net1790));
 sg13g2_tiehi \cpu.ex.r_epc[9]$_DFFE_PP__1791  (.L_HI(net1791));
 sg13g2_tiehi \cpu.ex.r_fetch$_SDFF_PN1__1792  (.L_HI(net1792));
 sg13g2_tiehi \cpu.ex.r_flush_write$_SDFFE_PN0P__1793  (.L_HI(net1793));
 sg13g2_tiehi \cpu.ex.r_i_flush_all$_SDFF_PP0__1794  (.L_HI(net1794));
 sg13g2_tiehi \cpu.ex.r_ie$_SDFFE_PP0P__1795  (.L_HI(net1795));
 sg13g2_tiehi \cpu.ex.r_io_access$_SDFFE_PN0P__1796  (.L_HI(net1796));
 sg13g2_tiehi \cpu.ex.r_lr[0]$_DFFE_PP__1797  (.L_HI(net1797));
 sg13g2_tiehi \cpu.ex.r_lr[10]$_DFFE_PP__1798  (.L_HI(net1798));
 sg13g2_tiehi \cpu.ex.r_lr[11]$_DFFE_PP__1799  (.L_HI(net1799));
 sg13g2_tiehi \cpu.ex.r_lr[12]$_DFFE_PP__1800  (.L_HI(net1800));
 sg13g2_tiehi \cpu.ex.r_lr[13]$_DFFE_PP__1801  (.L_HI(net1801));
 sg13g2_tiehi \cpu.ex.r_lr[14]$_DFFE_PP__1802  (.L_HI(net1802));
 sg13g2_tiehi \cpu.ex.r_lr[1]$_DFFE_PP__1803  (.L_HI(net1803));
 sg13g2_tiehi \cpu.ex.r_lr[2]$_DFFE_PP__1804  (.L_HI(net1804));
 sg13g2_tiehi \cpu.ex.r_lr[3]$_DFFE_PP__1805  (.L_HI(net1805));
 sg13g2_tiehi \cpu.ex.r_lr[4]$_DFFE_PP__1806  (.L_HI(net1806));
 sg13g2_tiehi \cpu.ex.r_lr[5]$_DFFE_PP__1807  (.L_HI(net1807));
 sg13g2_tiehi \cpu.ex.r_lr[6]$_DFFE_PP__1808  (.L_HI(net1808));
 sg13g2_tiehi \cpu.ex.r_lr[7]$_DFFE_PP__1809  (.L_HI(net1809));
 sg13g2_tiehi \cpu.ex.r_lr[8]$_DFFE_PP__1810  (.L_HI(net1810));
 sg13g2_tiehi \cpu.ex.r_lr[9]$_DFFE_PP__1811  (.L_HI(net1811));
 sg13g2_tiehi \cpu.ex.r_mult[0]$_DFF_P__1812  (.L_HI(net1812));
 sg13g2_tiehi \cpu.ex.r_mult[10]$_DFF_P__1813  (.L_HI(net1813));
 sg13g2_tiehi \cpu.ex.r_mult[11]$_DFF_P__1814  (.L_HI(net1814));
 sg13g2_tiehi \cpu.ex.r_mult[12]$_DFF_P__1815  (.L_HI(net1815));
 sg13g2_tiehi \cpu.ex.r_mult[13]$_DFF_P__1816  (.L_HI(net1816));
 sg13g2_tiehi \cpu.ex.r_mult[14]$_DFF_P__1817  (.L_HI(net1817));
 sg13g2_tiehi \cpu.ex.r_mult[15]$_DFF_P__1818  (.L_HI(net1818));
 sg13g2_tiehi \cpu.ex.r_mult[16]$_DFFE_PP__1819  (.L_HI(net1819));
 sg13g2_tiehi \cpu.ex.r_mult[17]$_DFFE_PP__1820  (.L_HI(net1820));
 sg13g2_tiehi \cpu.ex.r_mult[18]$_DFFE_PP__1821  (.L_HI(net1821));
 sg13g2_tiehi \cpu.ex.r_mult[19]$_DFFE_PP__1822  (.L_HI(net1822));
 sg13g2_tiehi \cpu.ex.r_mult[1]$_DFF_P__1823  (.L_HI(net1823));
 sg13g2_tiehi \cpu.ex.r_mult[20]$_DFFE_PP__1824  (.L_HI(net1824));
 sg13g2_tiehi \cpu.ex.r_mult[21]$_DFFE_PP__1825  (.L_HI(net1825));
 sg13g2_tiehi \cpu.ex.r_mult[22]$_DFFE_PP__1826  (.L_HI(net1826));
 sg13g2_tiehi \cpu.ex.r_mult[23]$_DFFE_PP__1827  (.L_HI(net1827));
 sg13g2_tiehi \cpu.ex.r_mult[24]$_DFFE_PP__1828  (.L_HI(net1828));
 sg13g2_tiehi \cpu.ex.r_mult[25]$_DFFE_PP__1829  (.L_HI(net1829));
 sg13g2_tiehi \cpu.ex.r_mult[26]$_DFFE_PP__1830  (.L_HI(net1830));
 sg13g2_tiehi \cpu.ex.r_mult[27]$_DFFE_PP__1831  (.L_HI(net1831));
 sg13g2_tiehi \cpu.ex.r_mult[28]$_DFFE_PP__1832  (.L_HI(net1832));
 sg13g2_tiehi \cpu.ex.r_mult[29]$_DFFE_PP__1833  (.L_HI(net1833));
 sg13g2_tiehi \cpu.ex.r_mult[2]$_DFF_P__1834  (.L_HI(net1834));
 sg13g2_tiehi \cpu.ex.r_mult[30]$_DFFE_PP__1835  (.L_HI(net1835));
 sg13g2_tiehi \cpu.ex.r_mult[31]$_DFFE_PP__1836  (.L_HI(net1836));
 sg13g2_tiehi \cpu.ex.r_mult[3]$_DFF_P__1837  (.L_HI(net1837));
 sg13g2_tiehi \cpu.ex.r_mult[4]$_DFF_P__1838  (.L_HI(net1838));
 sg13g2_tiehi \cpu.ex.r_mult[5]$_DFF_P__1839  (.L_HI(net1839));
 sg13g2_tiehi \cpu.ex.r_mult[6]$_DFF_P__1840  (.L_HI(net1840));
 sg13g2_tiehi \cpu.ex.r_mult[7]$_DFF_P__1841  (.L_HI(net1841));
 sg13g2_tiehi \cpu.ex.r_mult[8]$_DFF_P__1842  (.L_HI(net1842));
 sg13g2_tiehi \cpu.ex.r_mult[9]$_DFF_P__1843  (.L_HI(net1843));
 sg13g2_tiehi \cpu.ex.r_mult_off[0]$_DFF_P__1844  (.L_HI(net1844));
 sg13g2_tiehi \cpu.ex.r_mult_off[1]$_DFF_P__1845  (.L_HI(net1845));
 sg13g2_tiehi \cpu.ex.r_mult_off[2]$_DFF_P__1846  (.L_HI(net1846));
 sg13g2_tiehi \cpu.ex.r_mult_off[3]$_DFF_P__1847  (.L_HI(net1847));
 sg13g2_tiehi \cpu.ex.r_mult_running$_DFF_P__1848  (.L_HI(net1848));
 sg13g2_tiehi \cpu.ex.r_pc[0]$_DFFE_PP__1849  (.L_HI(net1849));
 sg13g2_tiehi \cpu.ex.r_pc[10]$_DFFE_PP__1850  (.L_HI(net1850));
 sg13g2_tiehi \cpu.ex.r_pc[11]$_DFFE_PP__1851  (.L_HI(net1851));
 sg13g2_tiehi \cpu.ex.r_pc[12]$_DFFE_PP__1852  (.L_HI(net1852));
 sg13g2_tiehi \cpu.ex.r_pc[13]$_DFFE_PP__1853  (.L_HI(net1853));
 sg13g2_tiehi \cpu.ex.r_pc[14]$_DFFE_PP__1854  (.L_HI(net1854));
 sg13g2_tiehi \cpu.ex.r_pc[1]$_DFFE_PP__1855  (.L_HI(net1855));
 sg13g2_tiehi \cpu.ex.r_pc[2]$_DFFE_PP__1856  (.L_HI(net1856));
 sg13g2_tiehi \cpu.ex.r_pc[3]$_DFFE_PP__1857  (.L_HI(net1857));
 sg13g2_tiehi \cpu.ex.r_pc[4]$_DFFE_PP__1858  (.L_HI(net1858));
 sg13g2_tiehi \cpu.ex.r_pc[5]$_DFFE_PP__1859  (.L_HI(net1859));
 sg13g2_tiehi \cpu.ex.r_pc[6]$_DFFE_PP__1860  (.L_HI(net1860));
 sg13g2_tiehi \cpu.ex.r_pc[7]$_DFFE_PP__1861  (.L_HI(net1861));
 sg13g2_tiehi \cpu.ex.r_pc[8]$_DFFE_PP__1862  (.L_HI(net1862));
 sg13g2_tiehi \cpu.ex.r_pc[9]$_DFFE_PP__1863  (.L_HI(net1863));
 sg13g2_tiehi \cpu.ex.r_prev_ie$_SDFFE_PN0P__1864  (.L_HI(net1864));
 sg13g2_tiehi \cpu.ex.r_read_stall$_SDFFE_PN0P__1865  (.L_HI(net1865));
 sg13g2_tiehi \cpu.ex.r_set_cc$_DFFE_PP__1866  (.L_HI(net1866));
 sg13g2_tiehi \cpu.ex.r_sp[0]$_DFFE_PP__1867  (.L_HI(net1867));
 sg13g2_tiehi \cpu.ex.r_sp[10]$_DFFE_PP__1868  (.L_HI(net1868));
 sg13g2_tiehi \cpu.ex.r_sp[11]$_DFFE_PP__1869  (.L_HI(net1869));
 sg13g2_tiehi \cpu.ex.r_sp[12]$_DFFE_PP__1870  (.L_HI(net1870));
 sg13g2_tiehi \cpu.ex.r_sp[13]$_DFFE_PP__1871  (.L_HI(net1871));
 sg13g2_tiehi \cpu.ex.r_sp[14]$_DFFE_PP__1872  (.L_HI(net1872));
 sg13g2_tiehi \cpu.ex.r_sp[1]$_DFFE_PP__1873  (.L_HI(net1873));
 sg13g2_tiehi \cpu.ex.r_sp[2]$_DFFE_PP__1874  (.L_HI(net1874));
 sg13g2_tiehi \cpu.ex.r_sp[3]$_DFFE_PP__1875  (.L_HI(net1875));
 sg13g2_tiehi \cpu.ex.r_sp[4]$_DFFE_PP__1876  (.L_HI(net1876));
 sg13g2_tiehi \cpu.ex.r_sp[5]$_DFFE_PP__1877  (.L_HI(net1877));
 sg13g2_tiehi \cpu.ex.r_sp[6]$_DFFE_PP__1878  (.L_HI(net1878));
 sg13g2_tiehi \cpu.ex.r_sp[7]$_DFFE_PP__1879  (.L_HI(net1879));
 sg13g2_tiehi \cpu.ex.r_sp[8]$_DFFE_PP__1880  (.L_HI(net1880));
 sg13g2_tiehi \cpu.ex.r_sp[9]$_DFFE_PP__1881  (.L_HI(net1881));
 sg13g2_tiehi \cpu.ex.r_stmp[0]$_SDFFCE_PN0P__1882  (.L_HI(net1882));
 sg13g2_tiehi \cpu.ex.r_stmp[10]$_DFFE_PP__1883  (.L_HI(net1883));
 sg13g2_tiehi \cpu.ex.r_stmp[11]$_DFFE_PP__1884  (.L_HI(net1884));
 sg13g2_tiehi \cpu.ex.r_stmp[12]$_DFFE_PP__1885  (.L_HI(net1885));
 sg13g2_tiehi \cpu.ex.r_stmp[13]$_DFFE_PP__1886  (.L_HI(net1886));
 sg13g2_tiehi \cpu.ex.r_stmp[14]$_DFFE_PP__1887  (.L_HI(net1887));
 sg13g2_tiehi \cpu.ex.r_stmp[15]$_DFFE_PP__1888  (.L_HI(net1888));
 sg13g2_tiehi \cpu.ex.r_stmp[1]$_DFFE_PP__1889  (.L_HI(net1889));
 sg13g2_tiehi \cpu.ex.r_stmp[2]$_DFFE_PP__1890  (.L_HI(net1890));
 sg13g2_tiehi \cpu.ex.r_stmp[3]$_DFFE_PP__1891  (.L_HI(net1891));
 sg13g2_tiehi \cpu.ex.r_stmp[4]$_DFFE_PP__1892  (.L_HI(net1892));
 sg13g2_tiehi \cpu.ex.r_stmp[5]$_DFFE_PP__1893  (.L_HI(net1893));
 sg13g2_tiehi \cpu.ex.r_stmp[6]$_DFFE_PP__1894  (.L_HI(net1894));
 sg13g2_tiehi \cpu.ex.r_stmp[7]$_DFFE_PP__1895  (.L_HI(net1895));
 sg13g2_tiehi \cpu.ex.r_stmp[8]$_DFFE_PP__1896  (.L_HI(net1896));
 sg13g2_tiehi \cpu.ex.r_stmp[9]$_DFFE_PP__1897  (.L_HI(net1897));
 sg13g2_tiehi \cpu.ex.r_wb[0]$_DFFE_PP__1898  (.L_HI(net1898));
 sg13g2_tiehi \cpu.ex.r_wb[10]$_DFFE_PP__1899  (.L_HI(net1899));
 sg13g2_tiehi \cpu.ex.r_wb[11]$_DFFE_PP__1900  (.L_HI(net1900));
 sg13g2_tiehi \cpu.ex.r_wb[12]$_DFFE_PP__1901  (.L_HI(net1901));
 sg13g2_tiehi \cpu.ex.r_wb[13]$_DFFE_PP__1902  (.L_HI(net1902));
 sg13g2_tiehi \cpu.ex.r_wb[14]$_DFFE_PP__1903  (.L_HI(net1903));
 sg13g2_tiehi \cpu.ex.r_wb[15]$_DFFE_PP__1904  (.L_HI(net1904));
 sg13g2_tiehi \cpu.ex.r_wb[1]$_DFFE_PP__1905  (.L_HI(net1905));
 sg13g2_tiehi \cpu.ex.r_wb[2]$_DFFE_PP__1906  (.L_HI(net1906));
 sg13g2_tiehi \cpu.ex.r_wb[3]$_DFFE_PP__1907  (.L_HI(net1907));
 sg13g2_tiehi \cpu.ex.r_wb[4]$_DFFE_PP__1908  (.L_HI(net1908));
 sg13g2_tiehi \cpu.ex.r_wb[5]$_DFFE_PP__1909  (.L_HI(net1909));
 sg13g2_tiehi \cpu.ex.r_wb[6]$_DFFE_PP__1910  (.L_HI(net1910));
 sg13g2_tiehi \cpu.ex.r_wb[7]$_DFFE_PP__1911  (.L_HI(net1911));
 sg13g2_tiehi \cpu.ex.r_wb[8]$_DFFE_PP__1912  (.L_HI(net1912));
 sg13g2_tiehi \cpu.ex.r_wb[9]$_DFFE_PP__1913  (.L_HI(net1913));
 sg13g2_tiehi \cpu.ex.r_wb_addr[0]$_SDFFCE_PN0P__1914  (.L_HI(net1914));
 sg13g2_tiehi \cpu.ex.r_wb_addr[1]$_SDFFCE_PN0P__1915  (.L_HI(net1915));
 sg13g2_tiehi \cpu.ex.r_wb_addr[2]$_SDFFCE_PP0P__1916  (.L_HI(net1916));
 sg13g2_tiehi \cpu.ex.r_wb_addr[3]$_SDFFCE_PP0P__1917  (.L_HI(net1917));
 sg13g2_tiehi \cpu.ex.r_wb_swapsp$_DFFE_PP__1918  (.L_HI(net1918));
 sg13g2_tiehi \cpu.ex.r_wb_valid$_DFF_P__1919  (.L_HI(net1919));
 sg13g2_tiehi \cpu.ex.r_wdata[0]$_DFFE_PP__1920  (.L_HI(net1920));
 sg13g2_tiehi \cpu.ex.r_wdata[10]$_DFFE_PP__1921  (.L_HI(net1921));
 sg13g2_tiehi \cpu.ex.r_wdata[11]$_DFFE_PP__1922  (.L_HI(net1922));
 sg13g2_tiehi \cpu.ex.r_wdata[12]$_DFFE_PP__1923  (.L_HI(net1923));
 sg13g2_tiehi \cpu.ex.r_wdata[13]$_DFFE_PP__1924  (.L_HI(net1924));
 sg13g2_tiehi \cpu.ex.r_wdata[14]$_DFFE_PP__1925  (.L_HI(net1925));
 sg13g2_tiehi \cpu.ex.r_wdata[15]$_DFFE_PP__1926  (.L_HI(net1926));
 sg13g2_tiehi \cpu.ex.r_wdata[1]$_DFFE_PP__1927  (.L_HI(net1927));
 sg13g2_tiehi \cpu.ex.r_wdata[2]$_DFFE_PP__1928  (.L_HI(net1928));
 sg13g2_tiehi \cpu.ex.r_wdata[3]$_DFFE_PP__1929  (.L_HI(net1929));
 sg13g2_tiehi \cpu.ex.r_wdata[4]$_DFFE_PP__1930  (.L_HI(net1930));
 sg13g2_tiehi \cpu.ex.r_wdata[5]$_DFFE_PP__1931  (.L_HI(net1931));
 sg13g2_tiehi \cpu.ex.r_wdata[6]$_DFFE_PP__1932  (.L_HI(net1932));
 sg13g2_tiehi \cpu.ex.r_wdata[7]$_DFFE_PP__1933  (.L_HI(net1933));
 sg13g2_tiehi \cpu.ex.r_wdata[8]$_DFFE_PP__1934  (.L_HI(net1934));
 sg13g2_tiehi \cpu.ex.r_wdata[9]$_DFFE_PP__1935  (.L_HI(net1935));
 sg13g2_tiehi \cpu.ex.r_wmask[0]$_SDFFE_PP0P__1936  (.L_HI(net1936));
 sg13g2_tiehi \cpu.ex.r_wmask[1]$_SDFFE_PP0P__1937  (.L_HI(net1937));
 sg13g2_tiehi \cpu.genblk1.mmu.r_fault_address[0]$_DFFE_PP__1938  (.L_HI(net1938));
 sg13g2_tiehi \cpu.genblk1.mmu.r_fault_address[1]$_DFFE_PP__1939  (.L_HI(net1939));
 sg13g2_tiehi \cpu.genblk1.mmu.r_fault_address[2]$_DFFE_PP__1940  (.L_HI(net1940));
 sg13g2_tiehi \cpu.genblk1.mmu.r_fault_address[3]$_DFFE_PP__1941  (.L_HI(net1941));
 sg13g2_tiehi \cpu.genblk1.mmu.r_fault_ins$_SDFFE_PN0P__1942  (.L_HI(net1942));
 sg13g2_tiehi \cpu.genblk1.mmu.r_fault_sup$_SDFFE_PN0P__1943  (.L_HI(net1943));
 sg13g2_tiehi \cpu.genblk1.mmu.r_fault_type$_SDFFE_PN0P__1944  (.L_HI(net1944));
 sg13g2_tiehi \cpu.genblk1.mmu.r_valid_d[0]$_SDFFE_PN0P__1945  (.L_HI(net1945));
 sg13g2_tiehi \cpu.genblk1.mmu.r_valid_d[10]$_SDFFE_PN0P__1946  (.L_HI(net1946));
 sg13g2_tiehi \cpu.genblk1.mmu.r_valid_d[11]$_SDFFE_PN0P__1947  (.L_HI(net1947));
 sg13g2_tiehi \cpu.genblk1.mmu.r_valid_d[12]$_SDFFE_PN0P__1948  (.L_HI(net1948));
 sg13g2_tiehi \cpu.genblk1.mmu.r_valid_d[13]$_SDFFE_PN0P__1949  (.L_HI(net1949));
 sg13g2_tiehi \cpu.genblk1.mmu.r_valid_d[14]$_SDFFE_PN0P__1950  (.L_HI(net1950));
 sg13g2_tiehi \cpu.genblk1.mmu.r_valid_d[15]$_SDFFE_PN0P__1951  (.L_HI(net1951));
 sg13g2_tiehi \cpu.genblk1.mmu.r_valid_d[16]$_SDFFE_PN0P__1952  (.L_HI(net1952));
 sg13g2_tiehi \cpu.genblk1.mmu.r_valid_d[17]$_SDFFE_PN0P__1953  (.L_HI(net1953));
 sg13g2_tiehi \cpu.genblk1.mmu.r_valid_d[18]$_SDFFE_PN0P__1954  (.L_HI(net1954));
 sg13g2_tiehi \cpu.genblk1.mmu.r_valid_d[19]$_SDFFE_PN0P__1955  (.L_HI(net1955));
 sg13g2_tiehi \cpu.genblk1.mmu.r_valid_d[1]$_SDFFE_PN0P__1956  (.L_HI(net1956));
 sg13g2_tiehi \cpu.genblk1.mmu.r_valid_d[20]$_SDFFE_PN0P__1957  (.L_HI(net1957));
 sg13g2_tiehi \cpu.genblk1.mmu.r_valid_d[21]$_SDFFE_PN0P__1958  (.L_HI(net1958));
 sg13g2_tiehi \cpu.genblk1.mmu.r_valid_d[22]$_SDFFE_PN0P__1959  (.L_HI(net1959));
 sg13g2_tiehi \cpu.genblk1.mmu.r_valid_d[23]$_SDFFE_PN0P__1960  (.L_HI(net1960));
 sg13g2_tiehi \cpu.genblk1.mmu.r_valid_d[24]$_SDFFE_PN0P__1961  (.L_HI(net1961));
 sg13g2_tiehi \cpu.genblk1.mmu.r_valid_d[25]$_SDFFE_PN0P__1962  (.L_HI(net1962));
 sg13g2_tiehi \cpu.genblk1.mmu.r_valid_d[26]$_SDFFE_PN0P__1963  (.L_HI(net1963));
 sg13g2_tiehi \cpu.genblk1.mmu.r_valid_d[27]$_SDFFE_PN0P__1964  (.L_HI(net1964));
 sg13g2_tiehi \cpu.genblk1.mmu.r_valid_d[28]$_SDFFE_PN0P__1965  (.L_HI(net1965));
 sg13g2_tiehi \cpu.genblk1.mmu.r_valid_d[29]$_SDFFE_PN0P__1966  (.L_HI(net1966));
 sg13g2_tiehi \cpu.genblk1.mmu.r_valid_d[2]$_SDFFE_PN0P__1967  (.L_HI(net1967));
 sg13g2_tiehi \cpu.genblk1.mmu.r_valid_d[30]$_SDFFE_PN0P__1968  (.L_HI(net1968));
 sg13g2_tiehi \cpu.genblk1.mmu.r_valid_d[31]$_SDFFE_PN0P__1969  (.L_HI(net1969));
 sg13g2_tiehi \cpu.genblk1.mmu.r_valid_d[3]$_SDFFE_PN0P__1970  (.L_HI(net1970));
 sg13g2_tiehi \cpu.genblk1.mmu.r_valid_d[4]$_SDFFE_PN0P__1971  (.L_HI(net1971));
 sg13g2_tiehi \cpu.genblk1.mmu.r_valid_d[5]$_SDFFE_PN0P__1972  (.L_HI(net1972));
 sg13g2_tiehi \cpu.genblk1.mmu.r_valid_d[6]$_SDFFE_PN0P__1973  (.L_HI(net1973));
 sg13g2_tiehi \cpu.genblk1.mmu.r_valid_d[7]$_SDFFE_PN0P__1974  (.L_HI(net1974));
 sg13g2_tiehi \cpu.genblk1.mmu.r_valid_d[8]$_SDFFE_PN0P__1975  (.L_HI(net1975));
 sg13g2_tiehi \cpu.genblk1.mmu.r_valid_d[9]$_SDFFE_PN0P__1976  (.L_HI(net1976));
 sg13g2_tiehi \cpu.genblk1.mmu.r_valid_i[0]$_SDFFE_PN0P__1977  (.L_HI(net1977));
 sg13g2_tiehi \cpu.genblk1.mmu.r_valid_i[10]$_SDFFE_PN0P__1978  (.L_HI(net1978));
 sg13g2_tiehi \cpu.genblk1.mmu.r_valid_i[11]$_SDFFE_PN0P__1979  (.L_HI(net1979));
 sg13g2_tiehi \cpu.genblk1.mmu.r_valid_i[12]$_SDFFE_PN0P__1980  (.L_HI(net1980));
 sg13g2_tiehi \cpu.genblk1.mmu.r_valid_i[13]$_SDFFE_PN0P__1981  (.L_HI(net1981));
 sg13g2_tiehi \cpu.genblk1.mmu.r_valid_i[14]$_SDFFE_PN0P__1982  (.L_HI(net1982));
 sg13g2_tiehi \cpu.genblk1.mmu.r_valid_i[15]$_SDFFE_PN0P__1983  (.L_HI(net1983));
 sg13g2_tiehi \cpu.genblk1.mmu.r_valid_i[16]$_SDFFE_PN0P__1984  (.L_HI(net1984));
 sg13g2_tiehi \cpu.genblk1.mmu.r_valid_i[17]$_SDFFE_PN0P__1985  (.L_HI(net1985));
 sg13g2_tiehi \cpu.genblk1.mmu.r_valid_i[18]$_SDFFE_PN0P__1986  (.L_HI(net1986));
 sg13g2_tiehi \cpu.genblk1.mmu.r_valid_i[19]$_SDFFE_PN0P__1987  (.L_HI(net1987));
 sg13g2_tiehi \cpu.genblk1.mmu.r_valid_i[1]$_SDFFE_PN0P__1988  (.L_HI(net1988));
 sg13g2_tiehi \cpu.genblk1.mmu.r_valid_i[20]$_SDFFE_PN0P__1989  (.L_HI(net1989));
 sg13g2_tiehi \cpu.genblk1.mmu.r_valid_i[21]$_SDFFE_PN0P__1990  (.L_HI(net1990));
 sg13g2_tiehi \cpu.genblk1.mmu.r_valid_i[22]$_SDFFE_PN0P__1991  (.L_HI(net1991));
 sg13g2_tiehi \cpu.genblk1.mmu.r_valid_i[23]$_SDFFE_PN0P__1992  (.L_HI(net1992));
 sg13g2_tiehi \cpu.genblk1.mmu.r_valid_i[24]$_SDFFE_PN0P__1993  (.L_HI(net1993));
 sg13g2_tiehi \cpu.genblk1.mmu.r_valid_i[25]$_SDFFE_PN0P__1994  (.L_HI(net1994));
 sg13g2_tiehi \cpu.genblk1.mmu.r_valid_i[26]$_SDFFE_PN0P__1995  (.L_HI(net1995));
 sg13g2_tiehi \cpu.genblk1.mmu.r_valid_i[27]$_SDFFE_PN0P__1996  (.L_HI(net1996));
 sg13g2_tiehi \cpu.genblk1.mmu.r_valid_i[28]$_SDFFE_PN0P__1997  (.L_HI(net1997));
 sg13g2_tiehi \cpu.genblk1.mmu.r_valid_i[29]$_SDFFE_PN0P__1998  (.L_HI(net1998));
 sg13g2_tiehi \cpu.genblk1.mmu.r_valid_i[2]$_SDFFE_PN0P__1999  (.L_HI(net1999));
 sg13g2_tiehi \cpu.genblk1.mmu.r_valid_i[30]$_SDFFE_PN0P__2000  (.L_HI(net2000));
 sg13g2_tiehi \cpu.genblk1.mmu.r_valid_i[31]$_SDFFE_PN0P__2001  (.L_HI(net2001));
 sg13g2_tiehi \cpu.genblk1.mmu.r_valid_i[3]$_SDFFE_PN0P__2002  (.L_HI(net2002));
 sg13g2_tiehi \cpu.genblk1.mmu.r_valid_i[4]$_SDFFE_PN0P__2003  (.L_HI(net2003));
 sg13g2_tiehi \cpu.genblk1.mmu.r_valid_i[5]$_SDFFE_PN0P__2004  (.L_HI(net2004));
 sg13g2_tiehi \cpu.genblk1.mmu.r_valid_i[6]$_SDFFE_PN0P__2005  (.L_HI(net2005));
 sg13g2_tiehi \cpu.genblk1.mmu.r_valid_i[7]$_SDFFE_PN0P__2006  (.L_HI(net2006));
 sg13g2_tiehi \cpu.genblk1.mmu.r_valid_i[8]$_SDFFE_PN0P__2007  (.L_HI(net2007));
 sg13g2_tiehi \cpu.genblk1.mmu.r_valid_i[9]$_SDFFE_PN0P__2008  (.L_HI(net2008));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[0][0]$_DFFE_PP__2009  (.L_HI(net2009));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[0][10]$_DFFE_PP__2010  (.L_HI(net2010));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[0][11]$_DFFE_PP__2011  (.L_HI(net2011));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[0][1]$_DFFE_PP__2012  (.L_HI(net2012));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[0][2]$_DFFE_PP__2013  (.L_HI(net2013));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[0][3]$_DFFE_PP__2014  (.L_HI(net2014));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[0][4]$_DFFE_PP__2015  (.L_HI(net2015));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[0][5]$_DFFE_PP__2016  (.L_HI(net2016));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[0][6]$_DFFE_PP__2017  (.L_HI(net2017));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[0][7]$_DFFE_PP__2018  (.L_HI(net2018));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[0][8]$_DFFE_PP__2019  (.L_HI(net2019));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[0][9]$_DFFE_PP__2020  (.L_HI(net2020));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[10][0]$_DFFE_PP__2021  (.L_HI(net2021));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[10][10]$_DFFE_PP__2022  (.L_HI(net2022));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[10][11]$_DFFE_PP__2023  (.L_HI(net2023));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[10][1]$_DFFE_PP__2024  (.L_HI(net2024));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[10][2]$_DFFE_PP__2025  (.L_HI(net2025));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[10][3]$_DFFE_PP__2026  (.L_HI(net2026));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[10][4]$_DFFE_PP__2027  (.L_HI(net2027));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[10][5]$_DFFE_PP__2028  (.L_HI(net2028));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[10][6]$_DFFE_PP__2029  (.L_HI(net2029));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[10][7]$_DFFE_PP__2030  (.L_HI(net2030));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[10][8]$_DFFE_PP__2031  (.L_HI(net2031));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[10][9]$_DFFE_PP__2032  (.L_HI(net2032));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[11][0]$_DFFE_PP__2033  (.L_HI(net2033));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[11][10]$_DFFE_PP__2034  (.L_HI(net2034));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[11][11]$_DFFE_PP__2035  (.L_HI(net2035));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[11][1]$_DFFE_PP__2036  (.L_HI(net2036));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[11][2]$_DFFE_PP__2037  (.L_HI(net2037));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[11][3]$_DFFE_PP__2038  (.L_HI(net2038));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[11][4]$_DFFE_PP__2039  (.L_HI(net2039));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[11][5]$_DFFE_PP__2040  (.L_HI(net2040));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[11][6]$_DFFE_PP__2041  (.L_HI(net2041));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[11][7]$_DFFE_PP__2042  (.L_HI(net2042));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[11][8]$_DFFE_PP__2043  (.L_HI(net2043));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[11][9]$_DFFE_PP__2044  (.L_HI(net2044));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[12][0]$_DFFE_PP__2045  (.L_HI(net2045));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[12][10]$_DFFE_PP__2046  (.L_HI(net2046));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[12][11]$_DFFE_PP__2047  (.L_HI(net2047));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[12][1]$_DFFE_PP__2048  (.L_HI(net2048));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[12][2]$_DFFE_PP__2049  (.L_HI(net2049));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[12][3]$_DFFE_PP__2050  (.L_HI(net2050));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[12][4]$_DFFE_PP__2051  (.L_HI(net2051));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[12][5]$_DFFE_PP__2052  (.L_HI(net2052));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[12][6]$_DFFE_PP__2053  (.L_HI(net2053));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[12][7]$_DFFE_PP__2054  (.L_HI(net2054));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[12][8]$_DFFE_PP__2055  (.L_HI(net2055));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[12][9]$_DFFE_PP__2056  (.L_HI(net2056));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[13][0]$_DFFE_PP__2057  (.L_HI(net2057));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[13][10]$_DFFE_PP__2058  (.L_HI(net2058));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[13][11]$_DFFE_PP__2059  (.L_HI(net2059));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[13][1]$_DFFE_PP__2060  (.L_HI(net2060));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[13][2]$_DFFE_PP__2061  (.L_HI(net2061));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[13][3]$_DFFE_PP__2062  (.L_HI(net2062));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[13][4]$_DFFE_PP__2063  (.L_HI(net2063));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[13][5]$_DFFE_PP__2064  (.L_HI(net2064));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[13][6]$_DFFE_PP__2065  (.L_HI(net2065));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[13][7]$_DFFE_PP__2066  (.L_HI(net2066));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[13][8]$_DFFE_PP__2067  (.L_HI(net2067));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[13][9]$_DFFE_PP__2068  (.L_HI(net2068));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[14][0]$_DFFE_PP__2069  (.L_HI(net2069));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[14][10]$_DFFE_PP__2070  (.L_HI(net2070));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[14][11]$_DFFE_PP__2071  (.L_HI(net2071));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[14][1]$_DFFE_PP__2072  (.L_HI(net2072));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[14][2]$_DFFE_PP__2073  (.L_HI(net2073));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[14][3]$_DFFE_PP__2074  (.L_HI(net2074));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[14][4]$_DFFE_PP__2075  (.L_HI(net2075));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[14][5]$_DFFE_PP__2076  (.L_HI(net2076));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[14][6]$_DFFE_PP__2077  (.L_HI(net2077));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[14][7]$_DFFE_PP__2078  (.L_HI(net2078));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[14][8]$_DFFE_PP__2079  (.L_HI(net2079));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[14][9]$_DFFE_PP__2080  (.L_HI(net2080));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[15][0]$_DFFE_PP__2081  (.L_HI(net2081));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[15][10]$_DFFE_PP__2082  (.L_HI(net2082));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[15][11]$_DFFE_PP__2083  (.L_HI(net2083));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[15][1]$_DFFE_PP__2084  (.L_HI(net2084));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[15][2]$_DFFE_PP__2085  (.L_HI(net2085));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[15][3]$_DFFE_PP__2086  (.L_HI(net2086));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[15][4]$_DFFE_PP__2087  (.L_HI(net2087));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[15][5]$_DFFE_PP__2088  (.L_HI(net2088));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[15][6]$_DFFE_PP__2089  (.L_HI(net2089));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[15][7]$_DFFE_PP__2090  (.L_HI(net2090));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[15][8]$_DFFE_PP__2091  (.L_HI(net2091));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[15][9]$_DFFE_PP__2092  (.L_HI(net2092));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[16][0]$_DFFE_PP__2093  (.L_HI(net2093));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[16][10]$_DFFE_PP__2094  (.L_HI(net2094));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[16][11]$_DFFE_PP__2095  (.L_HI(net2095));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[16][1]$_DFFE_PP__2096  (.L_HI(net2096));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[16][2]$_DFFE_PP__2097  (.L_HI(net2097));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[16][3]$_DFFE_PP__2098  (.L_HI(net2098));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[16][4]$_DFFE_PP__2099  (.L_HI(net2099));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[16][5]$_DFFE_PP__2100  (.L_HI(net2100));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[16][6]$_DFFE_PP__2101  (.L_HI(net2101));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[16][7]$_DFFE_PP__2102  (.L_HI(net2102));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[16][8]$_DFFE_PP__2103  (.L_HI(net2103));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[16][9]$_DFFE_PP__2104  (.L_HI(net2104));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[17][0]$_DFFE_PP__2105  (.L_HI(net2105));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[17][10]$_DFFE_PP__2106  (.L_HI(net2106));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[17][11]$_DFFE_PP__2107  (.L_HI(net2107));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[17][1]$_DFFE_PP__2108  (.L_HI(net2108));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[17][2]$_DFFE_PP__2109  (.L_HI(net2109));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[17][3]$_DFFE_PP__2110  (.L_HI(net2110));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[17][4]$_DFFE_PP__2111  (.L_HI(net2111));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[17][5]$_DFFE_PP__2112  (.L_HI(net2112));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[17][6]$_DFFE_PP__2113  (.L_HI(net2113));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[17][7]$_DFFE_PP__2114  (.L_HI(net2114));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[17][8]$_DFFE_PP__2115  (.L_HI(net2115));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[17][9]$_DFFE_PP__2116  (.L_HI(net2116));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[18][0]$_DFFE_PP__2117  (.L_HI(net2117));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[18][10]$_DFFE_PP__2118  (.L_HI(net2118));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[18][11]$_DFFE_PP__2119  (.L_HI(net2119));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[18][1]$_DFFE_PP__2120  (.L_HI(net2120));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[18][2]$_DFFE_PP__2121  (.L_HI(net2121));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[18][3]$_DFFE_PP__2122  (.L_HI(net2122));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[18][4]$_DFFE_PP__2123  (.L_HI(net2123));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[18][5]$_DFFE_PP__2124  (.L_HI(net2124));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[18][6]$_DFFE_PP__2125  (.L_HI(net2125));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[18][7]$_DFFE_PP__2126  (.L_HI(net2126));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[18][8]$_DFFE_PP__2127  (.L_HI(net2127));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[18][9]$_DFFE_PP__2128  (.L_HI(net2128));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[19][0]$_DFFE_PP__2129  (.L_HI(net2129));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[19][10]$_DFFE_PP__2130  (.L_HI(net2130));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[19][11]$_DFFE_PP__2131  (.L_HI(net2131));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[19][1]$_DFFE_PP__2132  (.L_HI(net2132));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[19][2]$_DFFE_PP__2133  (.L_HI(net2133));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[19][3]$_DFFE_PP__2134  (.L_HI(net2134));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[19][4]$_DFFE_PP__2135  (.L_HI(net2135));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[19][5]$_DFFE_PP__2136  (.L_HI(net2136));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[19][6]$_DFFE_PP__2137  (.L_HI(net2137));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[19][7]$_DFFE_PP__2138  (.L_HI(net2138));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[19][8]$_DFFE_PP__2139  (.L_HI(net2139));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[19][9]$_DFFE_PP__2140  (.L_HI(net2140));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[1][0]$_DFFE_PP__2141  (.L_HI(net2141));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[1][10]$_DFFE_PP__2142  (.L_HI(net2142));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[1][11]$_DFFE_PP__2143  (.L_HI(net2143));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[1][1]$_DFFE_PP__2144  (.L_HI(net2144));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[1][2]$_DFFE_PP__2145  (.L_HI(net2145));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[1][3]$_DFFE_PP__2146  (.L_HI(net2146));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[1][4]$_DFFE_PP__2147  (.L_HI(net2147));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[1][5]$_DFFE_PP__2148  (.L_HI(net2148));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[1][6]$_DFFE_PP__2149  (.L_HI(net2149));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[1][7]$_DFFE_PP__2150  (.L_HI(net2150));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[1][8]$_DFFE_PP__2151  (.L_HI(net2151));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[1][9]$_DFFE_PP__2152  (.L_HI(net2152));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[20][0]$_DFFE_PP__2153  (.L_HI(net2153));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[20][10]$_DFFE_PP__2154  (.L_HI(net2154));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[20][11]$_DFFE_PP__2155  (.L_HI(net2155));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[20][1]$_DFFE_PP__2156  (.L_HI(net2156));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[20][2]$_DFFE_PP__2157  (.L_HI(net2157));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[20][3]$_DFFE_PP__2158  (.L_HI(net2158));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[20][4]$_DFFE_PP__2159  (.L_HI(net2159));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[20][5]$_DFFE_PP__2160  (.L_HI(net2160));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[20][6]$_DFFE_PP__2161  (.L_HI(net2161));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[20][7]$_DFFE_PP__2162  (.L_HI(net2162));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[20][8]$_DFFE_PP__2163  (.L_HI(net2163));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[20][9]$_DFFE_PP__2164  (.L_HI(net2164));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[21][0]$_DFFE_PP__2165  (.L_HI(net2165));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[21][10]$_DFFE_PP__2166  (.L_HI(net2166));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[21][11]$_DFFE_PP__2167  (.L_HI(net2167));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[21][1]$_DFFE_PP__2168  (.L_HI(net2168));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[21][2]$_DFFE_PP__2169  (.L_HI(net2169));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[21][3]$_DFFE_PP__2170  (.L_HI(net2170));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[21][4]$_DFFE_PP__2171  (.L_HI(net2171));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[21][5]$_DFFE_PP__2172  (.L_HI(net2172));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[21][6]$_DFFE_PP__2173  (.L_HI(net2173));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[21][7]$_DFFE_PP__2174  (.L_HI(net2174));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[21][8]$_DFFE_PP__2175  (.L_HI(net2175));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[21][9]$_DFFE_PP__2176  (.L_HI(net2176));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[22][0]$_DFFE_PP__2177  (.L_HI(net2177));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[22][10]$_DFFE_PP__2178  (.L_HI(net2178));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[22][11]$_DFFE_PP__2179  (.L_HI(net2179));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[22][1]$_DFFE_PP__2180  (.L_HI(net2180));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[22][2]$_DFFE_PP__2181  (.L_HI(net2181));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[22][3]$_DFFE_PP__2182  (.L_HI(net2182));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[22][4]$_DFFE_PP__2183  (.L_HI(net2183));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[22][5]$_DFFE_PP__2184  (.L_HI(net2184));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[22][6]$_DFFE_PP__2185  (.L_HI(net2185));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[22][7]$_DFFE_PP__2186  (.L_HI(net2186));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[22][8]$_DFFE_PP__2187  (.L_HI(net2187));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[22][9]$_DFFE_PP__2188  (.L_HI(net2188));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[23][0]$_DFFE_PP__2189  (.L_HI(net2189));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[23][10]$_DFFE_PP__2190  (.L_HI(net2190));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[23][11]$_DFFE_PP__2191  (.L_HI(net2191));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[23][1]$_DFFE_PP__2192  (.L_HI(net2192));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[23][2]$_DFFE_PP__2193  (.L_HI(net2193));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[23][3]$_DFFE_PP__2194  (.L_HI(net2194));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[23][4]$_DFFE_PP__2195  (.L_HI(net2195));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[23][5]$_DFFE_PP__2196  (.L_HI(net2196));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[23][6]$_DFFE_PP__2197  (.L_HI(net2197));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[23][7]$_DFFE_PP__2198  (.L_HI(net2198));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[23][8]$_DFFE_PP__2199  (.L_HI(net2199));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[23][9]$_DFFE_PP__2200  (.L_HI(net2200));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[24][0]$_DFFE_PP__2201  (.L_HI(net2201));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[24][10]$_DFFE_PP__2202  (.L_HI(net2202));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[24][11]$_DFFE_PP__2203  (.L_HI(net2203));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[24][1]$_DFFE_PP__2204  (.L_HI(net2204));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[24][2]$_DFFE_PP__2205  (.L_HI(net2205));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[24][3]$_DFFE_PP__2206  (.L_HI(net2206));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[24][4]$_DFFE_PP__2207  (.L_HI(net2207));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[24][5]$_DFFE_PP__2208  (.L_HI(net2208));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[24][6]$_DFFE_PP__2209  (.L_HI(net2209));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[24][7]$_DFFE_PP__2210  (.L_HI(net2210));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[24][8]$_DFFE_PP__2211  (.L_HI(net2211));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[24][9]$_DFFE_PP__2212  (.L_HI(net2212));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[25][0]$_DFFE_PP__2213  (.L_HI(net2213));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[25][10]$_DFFE_PP__2214  (.L_HI(net2214));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[25][11]$_DFFE_PP__2215  (.L_HI(net2215));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[25][1]$_DFFE_PP__2216  (.L_HI(net2216));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[25][2]$_DFFE_PP__2217  (.L_HI(net2217));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[25][3]$_DFFE_PP__2218  (.L_HI(net2218));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[25][4]$_DFFE_PP__2219  (.L_HI(net2219));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[25][5]$_DFFE_PP__2220  (.L_HI(net2220));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[25][6]$_DFFE_PP__2221  (.L_HI(net2221));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[25][7]$_DFFE_PP__2222  (.L_HI(net2222));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[25][8]$_DFFE_PP__2223  (.L_HI(net2223));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[25][9]$_DFFE_PP__2224  (.L_HI(net2224));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[26][0]$_DFFE_PP__2225  (.L_HI(net2225));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[26][10]$_DFFE_PP__2226  (.L_HI(net2226));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[26][11]$_DFFE_PP__2227  (.L_HI(net2227));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[26][1]$_DFFE_PP__2228  (.L_HI(net2228));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[26][2]$_DFFE_PP__2229  (.L_HI(net2229));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[26][3]$_DFFE_PP__2230  (.L_HI(net2230));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[26][4]$_DFFE_PP__2231  (.L_HI(net2231));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[26][5]$_DFFE_PP__2232  (.L_HI(net2232));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[26][6]$_DFFE_PP__2233  (.L_HI(net2233));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[26][7]$_DFFE_PP__2234  (.L_HI(net2234));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[26][8]$_DFFE_PP__2235  (.L_HI(net2235));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[26][9]$_DFFE_PP__2236  (.L_HI(net2236));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[27][0]$_DFFE_PP__2237  (.L_HI(net2237));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[27][10]$_DFFE_PP__2238  (.L_HI(net2238));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[27][11]$_DFFE_PP__2239  (.L_HI(net2239));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[27][1]$_DFFE_PP__2240  (.L_HI(net2240));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[27][2]$_DFFE_PP__2241  (.L_HI(net2241));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[27][3]$_DFFE_PP__2242  (.L_HI(net2242));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[27][4]$_DFFE_PP__2243  (.L_HI(net2243));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[27][5]$_DFFE_PP__2244  (.L_HI(net2244));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[27][6]$_DFFE_PP__2245  (.L_HI(net2245));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[27][7]$_DFFE_PP__2246  (.L_HI(net2246));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[27][8]$_DFFE_PP__2247  (.L_HI(net2247));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[27][9]$_DFFE_PP__2248  (.L_HI(net2248));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[28][0]$_DFFE_PP__2249  (.L_HI(net2249));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[28][10]$_DFFE_PP__2250  (.L_HI(net2250));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[28][11]$_DFFE_PP__2251  (.L_HI(net2251));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[28][1]$_DFFE_PP__2252  (.L_HI(net2252));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[28][2]$_DFFE_PP__2253  (.L_HI(net2253));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[28][3]$_DFFE_PP__2254  (.L_HI(net2254));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[28][4]$_DFFE_PP__2255  (.L_HI(net2255));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[28][5]$_DFFE_PP__2256  (.L_HI(net2256));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[28][6]$_DFFE_PP__2257  (.L_HI(net2257));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[28][7]$_DFFE_PP__2258  (.L_HI(net2258));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[28][8]$_DFFE_PP__2259  (.L_HI(net2259));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[28][9]$_DFFE_PP__2260  (.L_HI(net2260));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[29][0]$_DFFE_PP__2261  (.L_HI(net2261));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[29][10]$_DFFE_PP__2262  (.L_HI(net2262));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[29][11]$_DFFE_PP__2263  (.L_HI(net2263));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[29][1]$_DFFE_PP__2264  (.L_HI(net2264));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[29][2]$_DFFE_PP__2265  (.L_HI(net2265));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[29][3]$_DFFE_PP__2266  (.L_HI(net2266));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[29][4]$_DFFE_PP__2267  (.L_HI(net2267));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[29][5]$_DFFE_PP__2268  (.L_HI(net2268));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[29][6]$_DFFE_PP__2269  (.L_HI(net2269));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[29][7]$_DFFE_PP__2270  (.L_HI(net2270));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[29][8]$_DFFE_PP__2271  (.L_HI(net2271));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[29][9]$_DFFE_PP__2272  (.L_HI(net2272));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[2][0]$_DFFE_PP__2273  (.L_HI(net2273));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[2][10]$_DFFE_PP__2274  (.L_HI(net2274));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[2][11]$_DFFE_PP__2275  (.L_HI(net2275));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[2][1]$_DFFE_PP__2276  (.L_HI(net2276));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[2][2]$_DFFE_PP__2277  (.L_HI(net2277));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[2][3]$_DFFE_PP__2278  (.L_HI(net2278));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[2][4]$_DFFE_PP__2279  (.L_HI(net2279));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[2][5]$_DFFE_PP__2280  (.L_HI(net2280));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[2][6]$_DFFE_PP__2281  (.L_HI(net2281));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[2][7]$_DFFE_PP__2282  (.L_HI(net2282));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[2][8]$_DFFE_PP__2283  (.L_HI(net2283));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[2][9]$_DFFE_PP__2284  (.L_HI(net2284));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[30][0]$_DFFE_PP__2285  (.L_HI(net2285));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[30][10]$_DFFE_PP__2286  (.L_HI(net2286));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[30][11]$_DFFE_PP__2287  (.L_HI(net2287));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[30][1]$_DFFE_PP__2288  (.L_HI(net2288));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[30][2]$_DFFE_PP__2289  (.L_HI(net2289));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[30][3]$_DFFE_PP__2290  (.L_HI(net2290));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[30][4]$_DFFE_PP__2291  (.L_HI(net2291));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[30][5]$_DFFE_PP__2292  (.L_HI(net2292));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[30][6]$_DFFE_PP__2293  (.L_HI(net2293));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[30][7]$_DFFE_PP__2294  (.L_HI(net2294));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[30][8]$_DFFE_PP__2295  (.L_HI(net2295));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[30][9]$_DFFE_PP__2296  (.L_HI(net2296));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[31][0]$_DFFE_PP__2297  (.L_HI(net2297));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[31][10]$_DFFE_PP__2298  (.L_HI(net2298));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[31][11]$_DFFE_PP__2299  (.L_HI(net2299));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[31][1]$_DFFE_PP__2300  (.L_HI(net2300));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[31][2]$_DFFE_PP__2301  (.L_HI(net2301));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[31][3]$_DFFE_PP__2302  (.L_HI(net2302));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[31][4]$_DFFE_PP__2303  (.L_HI(net2303));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[31][5]$_DFFE_PP__2304  (.L_HI(net2304));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[31][6]$_DFFE_PP__2305  (.L_HI(net2305));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[31][7]$_DFFE_PP__2306  (.L_HI(net2306));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[31][8]$_DFFE_PP__2307  (.L_HI(net2307));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[31][9]$_DFFE_PP__2308  (.L_HI(net2308));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[3][0]$_DFFE_PP__2309  (.L_HI(net2309));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[3][10]$_DFFE_PP__2310  (.L_HI(net2310));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[3][11]$_DFFE_PP__2311  (.L_HI(net2311));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[3][1]$_DFFE_PP__2312  (.L_HI(net2312));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[3][2]$_DFFE_PP__2313  (.L_HI(net2313));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[3][3]$_DFFE_PP__2314  (.L_HI(net2314));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[3][4]$_DFFE_PP__2315  (.L_HI(net2315));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[3][5]$_DFFE_PP__2316  (.L_HI(net2316));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[3][6]$_DFFE_PP__2317  (.L_HI(net2317));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[3][7]$_DFFE_PP__2318  (.L_HI(net2318));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[3][8]$_DFFE_PP__2319  (.L_HI(net2319));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[3][9]$_DFFE_PP__2320  (.L_HI(net2320));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[4][0]$_DFFE_PP__2321  (.L_HI(net2321));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[4][10]$_DFFE_PP__2322  (.L_HI(net2322));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[4][11]$_DFFE_PP__2323  (.L_HI(net2323));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[4][1]$_DFFE_PP__2324  (.L_HI(net2324));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[4][2]$_DFFE_PP__2325  (.L_HI(net2325));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[4][3]$_DFFE_PP__2326  (.L_HI(net2326));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[4][4]$_DFFE_PP__2327  (.L_HI(net2327));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[4][5]$_DFFE_PP__2328  (.L_HI(net2328));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[4][6]$_DFFE_PP__2329  (.L_HI(net2329));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[4][7]$_DFFE_PP__2330  (.L_HI(net2330));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[4][8]$_DFFE_PP__2331  (.L_HI(net2331));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[4][9]$_DFFE_PP__2332  (.L_HI(net2332));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[5][0]$_DFFE_PP__2333  (.L_HI(net2333));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[5][10]$_DFFE_PP__2334  (.L_HI(net2334));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[5][11]$_DFFE_PP__2335  (.L_HI(net2335));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[5][1]$_DFFE_PP__2336  (.L_HI(net2336));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[5][2]$_DFFE_PP__2337  (.L_HI(net2337));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[5][3]$_DFFE_PP__2338  (.L_HI(net2338));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[5][4]$_DFFE_PP__2339  (.L_HI(net2339));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[5][5]$_DFFE_PP__2340  (.L_HI(net2340));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[5][6]$_DFFE_PP__2341  (.L_HI(net2341));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[5][7]$_DFFE_PP__2342  (.L_HI(net2342));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[5][8]$_DFFE_PP__2343  (.L_HI(net2343));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[5][9]$_DFFE_PP__2344  (.L_HI(net2344));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[6][0]$_DFFE_PP__2345  (.L_HI(net2345));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[6][10]$_DFFE_PP__2346  (.L_HI(net2346));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[6][11]$_DFFE_PP__2347  (.L_HI(net2347));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[6][1]$_DFFE_PP__2348  (.L_HI(net2348));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[6][2]$_DFFE_PP__2349  (.L_HI(net2349));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[6][3]$_DFFE_PP__2350  (.L_HI(net2350));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[6][4]$_DFFE_PP__2351  (.L_HI(net2351));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[6][5]$_DFFE_PP__2352  (.L_HI(net2352));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[6][6]$_DFFE_PP__2353  (.L_HI(net2353));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[6][7]$_DFFE_PP__2354  (.L_HI(net2354));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[6][8]$_DFFE_PP__2355  (.L_HI(net2355));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[6][9]$_DFFE_PP__2356  (.L_HI(net2356));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[7][0]$_DFFE_PP__2357  (.L_HI(net2357));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[7][10]$_DFFE_PP__2358  (.L_HI(net2358));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[7][11]$_DFFE_PP__2359  (.L_HI(net2359));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[7][1]$_DFFE_PP__2360  (.L_HI(net2360));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[7][2]$_DFFE_PP__2361  (.L_HI(net2361));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[7][3]$_DFFE_PP__2362  (.L_HI(net2362));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[7][4]$_DFFE_PP__2363  (.L_HI(net2363));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[7][5]$_DFFE_PP__2364  (.L_HI(net2364));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[7][6]$_DFFE_PP__2365  (.L_HI(net2365));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[7][7]$_DFFE_PP__2366  (.L_HI(net2366));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[7][8]$_DFFE_PP__2367  (.L_HI(net2367));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[7][9]$_DFFE_PP__2368  (.L_HI(net2368));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[8][0]$_DFFE_PP__2369  (.L_HI(net2369));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[8][10]$_DFFE_PP__2370  (.L_HI(net2370));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[8][11]$_DFFE_PP__2371  (.L_HI(net2371));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[8][1]$_DFFE_PP__2372  (.L_HI(net2372));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[8][2]$_DFFE_PP__2373  (.L_HI(net2373));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[8][3]$_DFFE_PP__2374  (.L_HI(net2374));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[8][4]$_DFFE_PP__2375  (.L_HI(net2375));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[8][5]$_DFFE_PP__2376  (.L_HI(net2376));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[8][6]$_DFFE_PP__2377  (.L_HI(net2377));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[8][7]$_DFFE_PP__2378  (.L_HI(net2378));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[8][8]$_DFFE_PP__2379  (.L_HI(net2379));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[8][9]$_DFFE_PP__2380  (.L_HI(net2380));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[9][0]$_DFFE_PP__2381  (.L_HI(net2381));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[9][10]$_DFFE_PP__2382  (.L_HI(net2382));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[9][11]$_DFFE_PP__2383  (.L_HI(net2383));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[9][1]$_DFFE_PP__2384  (.L_HI(net2384));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[9][2]$_DFFE_PP__2385  (.L_HI(net2385));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[9][3]$_DFFE_PP__2386  (.L_HI(net2386));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[9][4]$_DFFE_PP__2387  (.L_HI(net2387));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[9][5]$_DFFE_PP__2388  (.L_HI(net2388));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[9][6]$_DFFE_PP__2389  (.L_HI(net2389));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[9][7]$_DFFE_PP__2390  (.L_HI(net2390));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[9][8]$_DFFE_PP__2391  (.L_HI(net2391));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[9][9]$_DFFE_PP__2392  (.L_HI(net2392));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[0][0]$_DFFE_PP__2393  (.L_HI(net2393));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[0][10]$_DFFE_PP__2394  (.L_HI(net2394));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[0][11]$_DFFE_PP__2395  (.L_HI(net2395));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[0][1]$_DFFE_PP__2396  (.L_HI(net2396));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[0][2]$_DFFE_PP__2397  (.L_HI(net2397));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[0][3]$_DFFE_PP__2398  (.L_HI(net2398));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[0][4]$_DFFE_PP__2399  (.L_HI(net2399));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[0][5]$_DFFE_PP__2400  (.L_HI(net2400));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[0][6]$_DFFE_PP__2401  (.L_HI(net2401));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[0][7]$_DFFE_PP__2402  (.L_HI(net2402));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[0][8]$_DFFE_PP__2403  (.L_HI(net2403));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[0][9]$_DFFE_PP__2404  (.L_HI(net2404));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[10][0]$_DFFE_PP__2405  (.L_HI(net2405));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[10][10]$_DFFE_PP__2406  (.L_HI(net2406));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[10][11]$_DFFE_PP__2407  (.L_HI(net2407));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[10][1]$_DFFE_PP__2408  (.L_HI(net2408));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[10][2]$_DFFE_PP__2409  (.L_HI(net2409));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[10][3]$_DFFE_PP__2410  (.L_HI(net2410));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[10][4]$_DFFE_PP__2411  (.L_HI(net2411));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[10][5]$_DFFE_PP__2412  (.L_HI(net2412));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[10][6]$_DFFE_PP__2413  (.L_HI(net2413));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[10][7]$_DFFE_PP__2414  (.L_HI(net2414));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[10][8]$_DFFE_PP__2415  (.L_HI(net2415));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[10][9]$_DFFE_PP__2416  (.L_HI(net2416));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[11][0]$_DFFE_PP__2417  (.L_HI(net2417));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[11][10]$_DFFE_PP__2418  (.L_HI(net2418));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[11][11]$_DFFE_PP__2419  (.L_HI(net2419));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[11][1]$_DFFE_PP__2420  (.L_HI(net2420));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[11][2]$_DFFE_PP__2421  (.L_HI(net2421));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[11][3]$_DFFE_PP__2422  (.L_HI(net2422));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[11][4]$_DFFE_PP__2423  (.L_HI(net2423));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[11][5]$_DFFE_PP__2424  (.L_HI(net2424));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[11][6]$_DFFE_PP__2425  (.L_HI(net2425));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[11][7]$_DFFE_PP__2426  (.L_HI(net2426));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[11][8]$_DFFE_PP__2427  (.L_HI(net2427));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[11][9]$_DFFE_PP__2428  (.L_HI(net2428));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[12][0]$_DFFE_PP__2429  (.L_HI(net2429));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[12][10]$_DFFE_PP__2430  (.L_HI(net2430));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[12][11]$_DFFE_PP__2431  (.L_HI(net2431));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[12][1]$_DFFE_PP__2432  (.L_HI(net2432));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[12][2]$_DFFE_PP__2433  (.L_HI(net2433));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[12][3]$_DFFE_PP__2434  (.L_HI(net2434));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[12][4]$_DFFE_PP__2435  (.L_HI(net2435));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[12][5]$_DFFE_PP__2436  (.L_HI(net2436));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[12][6]$_DFFE_PP__2437  (.L_HI(net2437));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[12][7]$_DFFE_PP__2438  (.L_HI(net2438));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[12][8]$_DFFE_PP__2439  (.L_HI(net2439));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[12][9]$_DFFE_PP__2440  (.L_HI(net2440));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[13][0]$_DFFE_PP__2441  (.L_HI(net2441));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[13][10]$_DFFE_PP__2442  (.L_HI(net2442));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[13][11]$_DFFE_PP__2443  (.L_HI(net2443));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[13][1]$_DFFE_PP__2444  (.L_HI(net2444));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[13][2]$_DFFE_PP__2445  (.L_HI(net2445));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[13][3]$_DFFE_PP__2446  (.L_HI(net2446));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[13][4]$_DFFE_PP__2447  (.L_HI(net2447));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[13][5]$_DFFE_PP__2448  (.L_HI(net2448));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[13][6]$_DFFE_PP__2449  (.L_HI(net2449));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[13][7]$_DFFE_PP__2450  (.L_HI(net2450));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[13][8]$_DFFE_PP__2451  (.L_HI(net2451));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[13][9]$_DFFE_PP__2452  (.L_HI(net2452));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[14][0]$_DFFE_PP__2453  (.L_HI(net2453));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[14][10]$_DFFE_PP__2454  (.L_HI(net2454));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[14][11]$_DFFE_PP__2455  (.L_HI(net2455));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[14][1]$_DFFE_PP__2456  (.L_HI(net2456));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[14][2]$_DFFE_PP__2457  (.L_HI(net2457));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[14][3]$_DFFE_PP__2458  (.L_HI(net2458));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[14][4]$_DFFE_PP__2459  (.L_HI(net2459));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[14][5]$_DFFE_PP__2460  (.L_HI(net2460));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[14][6]$_DFFE_PP__2461  (.L_HI(net2461));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[14][7]$_DFFE_PP__2462  (.L_HI(net2462));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[14][8]$_DFFE_PP__2463  (.L_HI(net2463));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[14][9]$_DFFE_PP__2464  (.L_HI(net2464));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[15][0]$_DFFE_PP__2465  (.L_HI(net2465));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[15][10]$_DFFE_PP__2466  (.L_HI(net2466));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[15][11]$_DFFE_PP__2467  (.L_HI(net2467));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[15][1]$_DFFE_PP__2468  (.L_HI(net2468));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[15][2]$_DFFE_PP__2469  (.L_HI(net2469));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[15][3]$_DFFE_PP__2470  (.L_HI(net2470));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[15][4]$_DFFE_PP__2471  (.L_HI(net2471));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[15][5]$_DFFE_PP__2472  (.L_HI(net2472));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[15][6]$_DFFE_PP__2473  (.L_HI(net2473));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[15][7]$_DFFE_PP__2474  (.L_HI(net2474));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[15][8]$_DFFE_PP__2475  (.L_HI(net2475));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[15][9]$_DFFE_PP__2476  (.L_HI(net2476));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[16][0]$_DFFE_PP__2477  (.L_HI(net2477));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[16][10]$_DFFE_PP__2478  (.L_HI(net2478));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[16][11]$_DFFE_PP__2479  (.L_HI(net2479));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[16][1]$_DFFE_PP__2480  (.L_HI(net2480));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[16][2]$_DFFE_PP__2481  (.L_HI(net2481));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[16][3]$_DFFE_PP__2482  (.L_HI(net2482));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[16][4]$_DFFE_PP__2483  (.L_HI(net2483));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[16][5]$_DFFE_PP__2484  (.L_HI(net2484));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[16][6]$_DFFE_PP__2485  (.L_HI(net2485));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[16][7]$_DFFE_PP__2486  (.L_HI(net2486));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[16][8]$_DFFE_PP__2487  (.L_HI(net2487));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[16][9]$_DFFE_PP__2488  (.L_HI(net2488));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[17][0]$_DFFE_PP__2489  (.L_HI(net2489));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[17][10]$_DFFE_PP__2490  (.L_HI(net2490));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[17][11]$_DFFE_PP__2491  (.L_HI(net2491));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[17][1]$_DFFE_PP__2492  (.L_HI(net2492));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[17][2]$_DFFE_PP__2493  (.L_HI(net2493));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[17][3]$_DFFE_PP__2494  (.L_HI(net2494));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[17][4]$_DFFE_PP__2495  (.L_HI(net2495));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[17][5]$_DFFE_PP__2496  (.L_HI(net2496));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[17][6]$_DFFE_PP__2497  (.L_HI(net2497));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[17][7]$_DFFE_PP__2498  (.L_HI(net2498));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[17][8]$_DFFE_PP__2499  (.L_HI(net2499));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[17][9]$_DFFE_PP__2500  (.L_HI(net2500));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[18][0]$_DFFE_PP__2501  (.L_HI(net2501));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[18][10]$_DFFE_PP__2502  (.L_HI(net2502));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[18][11]$_DFFE_PP__2503  (.L_HI(net2503));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[18][1]$_DFFE_PP__2504  (.L_HI(net2504));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[18][2]$_DFFE_PP__2505  (.L_HI(net2505));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[18][3]$_DFFE_PP__2506  (.L_HI(net2506));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[18][4]$_DFFE_PP__2507  (.L_HI(net2507));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[18][5]$_DFFE_PP__2508  (.L_HI(net2508));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[18][6]$_DFFE_PP__2509  (.L_HI(net2509));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[18][7]$_DFFE_PP__2510  (.L_HI(net2510));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[18][8]$_DFFE_PP__2511  (.L_HI(net2511));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[18][9]$_DFFE_PP__2512  (.L_HI(net2512));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[19][0]$_DFFE_PP__2513  (.L_HI(net2513));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[19][10]$_DFFE_PP__2514  (.L_HI(net2514));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[19][11]$_DFFE_PP__2515  (.L_HI(net2515));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[19][1]$_DFFE_PP__2516  (.L_HI(net2516));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[19][2]$_DFFE_PP__2517  (.L_HI(net2517));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[19][3]$_DFFE_PP__2518  (.L_HI(net2518));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[19][4]$_DFFE_PP__2519  (.L_HI(net2519));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[19][5]$_DFFE_PP__2520  (.L_HI(net2520));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[19][6]$_DFFE_PP__2521  (.L_HI(net2521));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[19][7]$_DFFE_PP__2522  (.L_HI(net2522));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[19][8]$_DFFE_PP__2523  (.L_HI(net2523));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[19][9]$_DFFE_PP__2524  (.L_HI(net2524));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[1][0]$_DFFE_PP__2525  (.L_HI(net2525));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[1][10]$_DFFE_PP__2526  (.L_HI(net2526));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[1][11]$_DFFE_PP__2527  (.L_HI(net2527));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[1][1]$_DFFE_PP__2528  (.L_HI(net2528));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[1][2]$_DFFE_PP__2529  (.L_HI(net2529));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[1][3]$_DFFE_PP__2530  (.L_HI(net2530));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[1][4]$_DFFE_PP__2531  (.L_HI(net2531));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[1][5]$_DFFE_PP__2532  (.L_HI(net2532));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[1][6]$_DFFE_PP__2533  (.L_HI(net2533));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[1][7]$_DFFE_PP__2534  (.L_HI(net2534));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[1][8]$_DFFE_PP__2535  (.L_HI(net2535));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[1][9]$_DFFE_PP__2536  (.L_HI(net2536));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[20][0]$_DFFE_PP__2537  (.L_HI(net2537));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[20][10]$_DFFE_PP__2538  (.L_HI(net2538));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[20][11]$_DFFE_PP__2539  (.L_HI(net2539));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[20][1]$_DFFE_PP__2540  (.L_HI(net2540));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[20][2]$_DFFE_PP__2541  (.L_HI(net2541));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[20][3]$_DFFE_PP__2542  (.L_HI(net2542));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[20][4]$_DFFE_PP__2543  (.L_HI(net2543));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[20][5]$_DFFE_PP__2544  (.L_HI(net2544));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[20][6]$_DFFE_PP__2545  (.L_HI(net2545));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[20][7]$_DFFE_PP__2546  (.L_HI(net2546));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[20][8]$_DFFE_PP__2547  (.L_HI(net2547));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[20][9]$_DFFE_PP__2548  (.L_HI(net2548));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[21][0]$_DFFE_PP__2549  (.L_HI(net2549));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[21][10]$_DFFE_PP__2550  (.L_HI(net2550));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[21][11]$_DFFE_PP__2551  (.L_HI(net2551));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[21][1]$_DFFE_PP__2552  (.L_HI(net2552));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[21][2]$_DFFE_PP__2553  (.L_HI(net2553));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[21][3]$_DFFE_PP__2554  (.L_HI(net2554));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[21][4]$_DFFE_PP__2555  (.L_HI(net2555));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[21][5]$_DFFE_PP__2556  (.L_HI(net2556));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[21][6]$_DFFE_PP__2557  (.L_HI(net2557));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[21][7]$_DFFE_PP__2558  (.L_HI(net2558));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[21][8]$_DFFE_PP__2559  (.L_HI(net2559));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[21][9]$_DFFE_PP__2560  (.L_HI(net2560));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[22][0]$_DFFE_PP__2561  (.L_HI(net2561));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[22][10]$_DFFE_PP__2562  (.L_HI(net2562));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[22][11]$_DFFE_PP__2563  (.L_HI(net2563));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[22][1]$_DFFE_PP__2564  (.L_HI(net2564));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[22][2]$_DFFE_PP__2565  (.L_HI(net2565));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[22][3]$_DFFE_PP__2566  (.L_HI(net2566));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[22][4]$_DFFE_PP__2567  (.L_HI(net2567));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[22][5]$_DFFE_PP__2568  (.L_HI(net2568));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[22][6]$_DFFE_PP__2569  (.L_HI(net2569));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[22][7]$_DFFE_PP__2570  (.L_HI(net2570));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[22][8]$_DFFE_PP__2571  (.L_HI(net2571));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[22][9]$_DFFE_PP__2572  (.L_HI(net2572));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[23][0]$_DFFE_PP__2573  (.L_HI(net2573));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[23][10]$_DFFE_PP__2574  (.L_HI(net2574));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[23][11]$_DFFE_PP__2575  (.L_HI(net2575));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[23][1]$_DFFE_PP__2576  (.L_HI(net2576));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[23][2]$_DFFE_PP__2577  (.L_HI(net2577));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[23][3]$_DFFE_PP__2578  (.L_HI(net2578));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[23][4]$_DFFE_PP__2579  (.L_HI(net2579));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[23][5]$_DFFE_PP__2580  (.L_HI(net2580));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[23][6]$_DFFE_PP__2581  (.L_HI(net2581));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[23][7]$_DFFE_PP__2582  (.L_HI(net2582));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[23][8]$_DFFE_PP__2583  (.L_HI(net2583));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[23][9]$_DFFE_PP__2584  (.L_HI(net2584));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[24][0]$_DFFE_PP__2585  (.L_HI(net2585));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[24][10]$_DFFE_PP__2586  (.L_HI(net2586));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[24][11]$_DFFE_PP__2587  (.L_HI(net2587));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[24][1]$_DFFE_PP__2588  (.L_HI(net2588));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[24][2]$_DFFE_PP__2589  (.L_HI(net2589));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[24][3]$_DFFE_PP__2590  (.L_HI(net2590));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[24][4]$_DFFE_PP__2591  (.L_HI(net2591));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[24][5]$_DFFE_PP__2592  (.L_HI(net2592));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[24][6]$_DFFE_PP__2593  (.L_HI(net2593));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[24][7]$_DFFE_PP__2594  (.L_HI(net2594));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[24][8]$_DFFE_PP__2595  (.L_HI(net2595));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[24][9]$_DFFE_PP__2596  (.L_HI(net2596));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[25][0]$_DFFE_PP__2597  (.L_HI(net2597));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[25][10]$_DFFE_PP__2598  (.L_HI(net2598));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[25][11]$_DFFE_PP__2599  (.L_HI(net2599));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[25][1]$_DFFE_PP__2600  (.L_HI(net2600));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[25][2]$_DFFE_PP__2601  (.L_HI(net2601));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[25][3]$_DFFE_PP__2602  (.L_HI(net2602));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[25][4]$_DFFE_PP__2603  (.L_HI(net2603));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[25][5]$_DFFE_PP__2604  (.L_HI(net2604));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[25][6]$_DFFE_PP__2605  (.L_HI(net2605));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[25][7]$_DFFE_PP__2606  (.L_HI(net2606));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[25][8]$_DFFE_PP__2607  (.L_HI(net2607));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[25][9]$_DFFE_PP__2608  (.L_HI(net2608));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[26][0]$_DFFE_PP__2609  (.L_HI(net2609));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[26][10]$_DFFE_PP__2610  (.L_HI(net2610));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[26][11]$_DFFE_PP__2611  (.L_HI(net2611));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[26][1]$_DFFE_PP__2612  (.L_HI(net2612));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[26][2]$_DFFE_PP__2613  (.L_HI(net2613));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[26][3]$_DFFE_PP__2614  (.L_HI(net2614));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[26][4]$_DFFE_PP__2615  (.L_HI(net2615));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[26][5]$_DFFE_PP__2616  (.L_HI(net2616));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[26][6]$_DFFE_PP__2617  (.L_HI(net2617));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[26][7]$_DFFE_PP__2618  (.L_HI(net2618));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[26][8]$_DFFE_PP__2619  (.L_HI(net2619));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[26][9]$_DFFE_PP__2620  (.L_HI(net2620));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[27][0]$_DFFE_PP__2621  (.L_HI(net2621));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[27][10]$_DFFE_PP__2622  (.L_HI(net2622));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[27][11]$_DFFE_PP__2623  (.L_HI(net2623));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[27][1]$_DFFE_PP__2624  (.L_HI(net2624));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[27][2]$_DFFE_PP__2625  (.L_HI(net2625));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[27][3]$_DFFE_PP__2626  (.L_HI(net2626));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[27][4]$_DFFE_PP__2627  (.L_HI(net2627));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[27][5]$_DFFE_PP__2628  (.L_HI(net2628));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[27][6]$_DFFE_PP__2629  (.L_HI(net2629));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[27][7]$_DFFE_PP__2630  (.L_HI(net2630));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[27][8]$_DFFE_PP__2631  (.L_HI(net2631));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[27][9]$_DFFE_PP__2632  (.L_HI(net2632));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[28][0]$_DFFE_PP__2633  (.L_HI(net2633));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[28][10]$_DFFE_PP__2634  (.L_HI(net2634));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[28][11]$_DFFE_PP__2635  (.L_HI(net2635));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[28][1]$_DFFE_PP__2636  (.L_HI(net2636));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[28][2]$_DFFE_PP__2637  (.L_HI(net2637));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[28][3]$_DFFE_PP__2638  (.L_HI(net2638));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[28][4]$_DFFE_PP__2639  (.L_HI(net2639));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[28][5]$_DFFE_PP__2640  (.L_HI(net2640));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[28][6]$_DFFE_PP__2641  (.L_HI(net2641));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[28][7]$_DFFE_PP__2642  (.L_HI(net2642));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[28][8]$_DFFE_PP__2643  (.L_HI(net2643));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[28][9]$_DFFE_PP__2644  (.L_HI(net2644));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[29][0]$_DFFE_PP__2645  (.L_HI(net2645));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[29][10]$_DFFE_PP__2646  (.L_HI(net2646));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[29][11]$_DFFE_PP__2647  (.L_HI(net2647));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[29][1]$_DFFE_PP__2648  (.L_HI(net2648));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[29][2]$_DFFE_PP__2649  (.L_HI(net2649));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[29][3]$_DFFE_PP__2650  (.L_HI(net2650));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[29][4]$_DFFE_PP__2651  (.L_HI(net2651));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[29][5]$_DFFE_PP__2652  (.L_HI(net2652));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[29][6]$_DFFE_PP__2653  (.L_HI(net2653));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[29][7]$_DFFE_PP__2654  (.L_HI(net2654));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[29][8]$_DFFE_PP__2655  (.L_HI(net2655));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[29][9]$_DFFE_PP__2656  (.L_HI(net2656));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[2][0]$_DFFE_PP__2657  (.L_HI(net2657));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[2][10]$_DFFE_PP__2658  (.L_HI(net2658));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[2][11]$_DFFE_PP__2659  (.L_HI(net2659));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[2][1]$_DFFE_PP__2660  (.L_HI(net2660));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[2][2]$_DFFE_PP__2661  (.L_HI(net2661));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[2][3]$_DFFE_PP__2662  (.L_HI(net2662));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[2][4]$_DFFE_PP__2663  (.L_HI(net2663));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[2][5]$_DFFE_PP__2664  (.L_HI(net2664));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[2][6]$_DFFE_PP__2665  (.L_HI(net2665));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[2][7]$_DFFE_PP__2666  (.L_HI(net2666));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[2][8]$_DFFE_PP__2667  (.L_HI(net2667));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[2][9]$_DFFE_PP__2668  (.L_HI(net2668));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[30][0]$_DFFE_PP__2669  (.L_HI(net2669));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[30][10]$_DFFE_PP__2670  (.L_HI(net2670));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[30][11]$_DFFE_PP__2671  (.L_HI(net2671));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[30][1]$_DFFE_PP__2672  (.L_HI(net2672));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[30][2]$_DFFE_PP__2673  (.L_HI(net2673));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[30][3]$_DFFE_PP__2674  (.L_HI(net2674));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[30][4]$_DFFE_PP__2675  (.L_HI(net2675));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[30][5]$_DFFE_PP__2676  (.L_HI(net2676));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[30][6]$_DFFE_PP__2677  (.L_HI(net2677));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[30][7]$_DFFE_PP__2678  (.L_HI(net2678));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[30][8]$_DFFE_PP__2679  (.L_HI(net2679));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[30][9]$_DFFE_PP__2680  (.L_HI(net2680));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[31][0]$_DFFE_PP__2681  (.L_HI(net2681));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[31][10]$_DFFE_PP__2682  (.L_HI(net2682));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[31][11]$_DFFE_PP__2683  (.L_HI(net2683));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[31][1]$_DFFE_PP__2684  (.L_HI(net2684));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[31][2]$_DFFE_PP__2685  (.L_HI(net2685));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[31][3]$_DFFE_PP__2686  (.L_HI(net2686));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[31][4]$_DFFE_PP__2687  (.L_HI(net2687));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[31][5]$_DFFE_PP__2688  (.L_HI(net2688));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[31][6]$_DFFE_PP__2689  (.L_HI(net2689));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[31][7]$_DFFE_PP__2690  (.L_HI(net2690));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[31][8]$_DFFE_PP__2691  (.L_HI(net2691));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[31][9]$_DFFE_PP__2692  (.L_HI(net2692));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[3][0]$_DFFE_PP__2693  (.L_HI(net2693));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[3][10]$_DFFE_PP__2694  (.L_HI(net2694));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[3][11]$_DFFE_PP__2695  (.L_HI(net2695));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[3][1]$_DFFE_PP__2696  (.L_HI(net2696));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[3][2]$_DFFE_PP__2697  (.L_HI(net2697));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[3][3]$_DFFE_PP__2698  (.L_HI(net2698));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[3][4]$_DFFE_PP__2699  (.L_HI(net2699));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[3][5]$_DFFE_PP__2700  (.L_HI(net2700));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[3][6]$_DFFE_PP__2701  (.L_HI(net2701));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[3][7]$_DFFE_PP__2702  (.L_HI(net2702));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[3][8]$_DFFE_PP__2703  (.L_HI(net2703));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[3][9]$_DFFE_PP__2704  (.L_HI(net2704));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[4][0]$_DFFE_PP__2705  (.L_HI(net2705));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[4][10]$_DFFE_PP__2706  (.L_HI(net2706));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[4][11]$_DFFE_PP__2707  (.L_HI(net2707));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[4][1]$_DFFE_PP__2708  (.L_HI(net2708));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[4][2]$_DFFE_PP__2709  (.L_HI(net2709));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[4][3]$_DFFE_PP__2710  (.L_HI(net2710));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[4][4]$_DFFE_PP__2711  (.L_HI(net2711));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[4][5]$_DFFE_PP__2712  (.L_HI(net2712));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[4][6]$_DFFE_PP__2713  (.L_HI(net2713));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[4][7]$_DFFE_PP__2714  (.L_HI(net2714));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[4][8]$_DFFE_PP__2715  (.L_HI(net2715));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[4][9]$_DFFE_PP__2716  (.L_HI(net2716));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[5][0]$_DFFE_PP__2717  (.L_HI(net2717));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[5][10]$_DFFE_PP__2718  (.L_HI(net2718));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[5][11]$_DFFE_PP__2719  (.L_HI(net2719));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[5][1]$_DFFE_PP__2720  (.L_HI(net2720));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[5][2]$_DFFE_PP__2721  (.L_HI(net2721));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[5][3]$_DFFE_PP__2722  (.L_HI(net2722));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[5][4]$_DFFE_PP__2723  (.L_HI(net2723));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[5][5]$_DFFE_PP__2724  (.L_HI(net2724));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[5][6]$_DFFE_PP__2725  (.L_HI(net2725));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[5][7]$_DFFE_PP__2726  (.L_HI(net2726));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[5][8]$_DFFE_PP__2727  (.L_HI(net2727));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[5][9]$_DFFE_PP__2728  (.L_HI(net2728));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[6][0]$_DFFE_PP__2729  (.L_HI(net2729));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[6][10]$_DFFE_PP__2730  (.L_HI(net2730));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[6][11]$_DFFE_PP__2731  (.L_HI(net2731));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[6][1]$_DFFE_PP__2732  (.L_HI(net2732));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[6][2]$_DFFE_PP__2733  (.L_HI(net2733));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[6][3]$_DFFE_PP__2734  (.L_HI(net2734));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[6][4]$_DFFE_PP__2735  (.L_HI(net2735));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[6][5]$_DFFE_PP__2736  (.L_HI(net2736));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[6][6]$_DFFE_PP__2737  (.L_HI(net2737));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[6][7]$_DFFE_PP__2738  (.L_HI(net2738));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[6][8]$_DFFE_PP__2739  (.L_HI(net2739));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[6][9]$_DFFE_PP__2740  (.L_HI(net2740));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[7][0]$_DFFE_PP__2741  (.L_HI(net2741));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[7][10]$_DFFE_PP__2742  (.L_HI(net2742));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[7][11]$_DFFE_PP__2743  (.L_HI(net2743));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[7][1]$_DFFE_PP__2744  (.L_HI(net2744));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[7][2]$_DFFE_PP__2745  (.L_HI(net2745));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[7][3]$_DFFE_PP__2746  (.L_HI(net2746));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[7][4]$_DFFE_PP__2747  (.L_HI(net2747));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[7][5]$_DFFE_PP__2748  (.L_HI(net2748));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[7][6]$_DFFE_PP__2749  (.L_HI(net2749));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[7][7]$_DFFE_PP__2750  (.L_HI(net2750));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[7][8]$_DFFE_PP__2751  (.L_HI(net2751));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[7][9]$_DFFE_PP__2752  (.L_HI(net2752));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[8][0]$_DFFE_PP__2753  (.L_HI(net2753));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[8][10]$_DFFE_PP__2754  (.L_HI(net2754));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[8][11]$_DFFE_PP__2755  (.L_HI(net2755));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[8][1]$_DFFE_PP__2756  (.L_HI(net2756));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[8][2]$_DFFE_PP__2757  (.L_HI(net2757));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[8][3]$_DFFE_PP__2758  (.L_HI(net2758));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[8][4]$_DFFE_PP__2759  (.L_HI(net2759));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[8][5]$_DFFE_PP__2760  (.L_HI(net2760));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[8][6]$_DFFE_PP__2761  (.L_HI(net2761));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[8][7]$_DFFE_PP__2762  (.L_HI(net2762));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[8][8]$_DFFE_PP__2763  (.L_HI(net2763));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[8][9]$_DFFE_PP__2764  (.L_HI(net2764));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[9][0]$_DFFE_PP__2765  (.L_HI(net2765));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[9][10]$_DFFE_PP__2766  (.L_HI(net2766));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[9][11]$_DFFE_PP__2767  (.L_HI(net2767));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[9][1]$_DFFE_PP__2768  (.L_HI(net2768));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[9][2]$_DFFE_PP__2769  (.L_HI(net2769));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[9][3]$_DFFE_PP__2770  (.L_HI(net2770));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[9][4]$_DFFE_PP__2771  (.L_HI(net2771));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[9][5]$_DFFE_PP__2772  (.L_HI(net2772));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[9][6]$_DFFE_PP__2773  (.L_HI(net2773));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[9][7]$_DFFE_PP__2774  (.L_HI(net2774));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[9][8]$_DFFE_PP__2775  (.L_HI(net2775));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[9][9]$_DFFE_PP__2776  (.L_HI(net2776));
 sg13g2_tiehi \cpu.genblk1.mmu.r_writeable_d[0]$_DFFE_PP__2777  (.L_HI(net2777));
 sg13g2_tiehi \cpu.genblk1.mmu.r_writeable_d[10]$_DFFE_PP__2778  (.L_HI(net2778));
 sg13g2_tiehi \cpu.genblk1.mmu.r_writeable_d[11]$_DFFE_PP__2779  (.L_HI(net2779));
 sg13g2_tiehi \cpu.genblk1.mmu.r_writeable_d[12]$_DFFE_PP__2780  (.L_HI(net2780));
 sg13g2_tiehi \cpu.genblk1.mmu.r_writeable_d[13]$_DFFE_PP__2781  (.L_HI(net2781));
 sg13g2_tiehi \cpu.genblk1.mmu.r_writeable_d[14]$_DFFE_PP__2782  (.L_HI(net2782));
 sg13g2_tiehi \cpu.genblk1.mmu.r_writeable_d[15]$_DFFE_PP__2783  (.L_HI(net2783));
 sg13g2_tiehi \cpu.genblk1.mmu.r_writeable_d[16]$_DFFE_PP__2784  (.L_HI(net2784));
 sg13g2_tiehi \cpu.genblk1.mmu.r_writeable_d[17]$_DFFE_PP__2785  (.L_HI(net2785));
 sg13g2_tiehi \cpu.genblk1.mmu.r_writeable_d[18]$_DFFE_PP__2786  (.L_HI(net2786));
 sg13g2_tiehi \cpu.genblk1.mmu.r_writeable_d[19]$_DFFE_PP__2787  (.L_HI(net2787));
 sg13g2_tiehi \cpu.genblk1.mmu.r_writeable_d[1]$_DFFE_PP__2788  (.L_HI(net2788));
 sg13g2_tiehi \cpu.genblk1.mmu.r_writeable_d[20]$_DFFE_PP__2789  (.L_HI(net2789));
 sg13g2_tiehi \cpu.genblk1.mmu.r_writeable_d[21]$_DFFE_PP__2790  (.L_HI(net2790));
 sg13g2_tiehi \cpu.genblk1.mmu.r_writeable_d[22]$_DFFE_PP__2791  (.L_HI(net2791));
 sg13g2_tiehi \cpu.genblk1.mmu.r_writeable_d[23]$_DFFE_PP__2792  (.L_HI(net2792));
 sg13g2_tiehi \cpu.genblk1.mmu.r_writeable_d[24]$_DFFE_PP__2793  (.L_HI(net2793));
 sg13g2_tiehi \cpu.genblk1.mmu.r_writeable_d[25]$_DFFE_PP__2794  (.L_HI(net2794));
 sg13g2_tiehi \cpu.genblk1.mmu.r_writeable_d[26]$_DFFE_PP__2795  (.L_HI(net2795));
 sg13g2_tiehi \cpu.genblk1.mmu.r_writeable_d[27]$_DFFE_PP__2796  (.L_HI(net2796));
 sg13g2_tiehi \cpu.genblk1.mmu.r_writeable_d[28]$_DFFE_PP__2797  (.L_HI(net2797));
 sg13g2_tiehi \cpu.genblk1.mmu.r_writeable_d[29]$_DFFE_PP__2798  (.L_HI(net2798));
 sg13g2_tiehi \cpu.genblk1.mmu.r_writeable_d[2]$_DFFE_PP__2799  (.L_HI(net2799));
 sg13g2_tiehi \cpu.genblk1.mmu.r_writeable_d[30]$_DFFE_PP__2800  (.L_HI(net2800));
 sg13g2_tiehi \cpu.genblk1.mmu.r_writeable_d[31]$_DFFE_PP__2801  (.L_HI(net2801));
 sg13g2_tiehi \cpu.genblk1.mmu.r_writeable_d[3]$_DFFE_PP__2802  (.L_HI(net2802));
 sg13g2_tiehi \cpu.genblk1.mmu.r_writeable_d[4]$_DFFE_PP__2803  (.L_HI(net2803));
 sg13g2_tiehi \cpu.genblk1.mmu.r_writeable_d[5]$_DFFE_PP__2804  (.L_HI(net2804));
 sg13g2_tiehi \cpu.genblk1.mmu.r_writeable_d[6]$_DFFE_PP__2805  (.L_HI(net2805));
 sg13g2_tiehi \cpu.genblk1.mmu.r_writeable_d[7]$_DFFE_PP__2806  (.L_HI(net2806));
 sg13g2_tiehi \cpu.genblk1.mmu.r_writeable_d[8]$_DFFE_PP__2807  (.L_HI(net2807));
 sg13g2_tiehi \cpu.genblk1.mmu.r_writeable_d[9]$_DFFE_PP__2808  (.L_HI(net2808));
 sg13g2_tiehi \cpu.gpio.r_enable_in[0]$_SDFFE_PN0P__2809  (.L_HI(net2809));
 sg13g2_tiehi \cpu.gpio.r_enable_in[1]$_SDFFE_PN0P__2810  (.L_HI(net2810));
 sg13g2_tiehi \cpu.gpio.r_enable_in[2]$_SDFFE_PN0P__2811  (.L_HI(net2811));
 sg13g2_tiehi \cpu.gpio.r_enable_in[3]$_SDFFE_PN0P__2812  (.L_HI(net2812));
 sg13g2_tiehi \cpu.gpio.r_enable_in[4]$_SDFFE_PN0P__2813  (.L_HI(net2813));
 sg13g2_tiehi \cpu.gpio.r_enable_in[5]$_SDFFE_PN0P__2814  (.L_HI(net2814));
 sg13g2_tiehi \cpu.gpio.r_enable_in[6]$_SDFFE_PN0P__2815  (.L_HI(net2815));
 sg13g2_tiehi \cpu.gpio.r_enable_in[7]$_SDFFE_PN0P__2816  (.L_HI(net2816));
 sg13g2_tiehi \cpu.gpio.r_enable_io[0]$_SDFFE_PN0P__2817  (.L_HI(net2817));
 sg13g2_tiehi \cpu.gpio.r_enable_io[1]$_SDFFE_PN0P__2818  (.L_HI(net2818));
 sg13g2_tiehi \cpu.gpio.r_enable_io[2]$_SDFFE_PN0P__2819  (.L_HI(net2819));
 sg13g2_tiehi \cpu.gpio.r_enable_io[3]$_SDFFE_PN0P__2820  (.L_HI(net2820));
 sg13g2_tiehi \cpu.gpio.r_gpio_en[0]$_SDFFE_PN0P__2821  (.L_HI(net2821));
 sg13g2_tiehi \cpu.gpio.r_gpio_en[1]$_SDFFE_PN0P__2822  (.L_HI(net2822));
 sg13g2_tiehi \cpu.gpio.r_gpio_en[2]$_SDFFE_PN0P__2823  (.L_HI(net2823));
 sg13g2_tiehi \cpu.gpio.r_gpio_en[3]$_SDFFE_PN0P__2824  (.L_HI(net2824));
 sg13g2_tiehi \cpu.gpio.r_gpio_io[0]$_DFFE_PP__2825  (.L_HI(net2825));
 sg13g2_tiehi \cpu.gpio.r_gpio_io[1]$_DFFE_PP__2826  (.L_HI(net2826));
 sg13g2_tiehi \cpu.gpio.r_gpio_io[2]$_DFFE_PP__2827  (.L_HI(net2827));
 sg13g2_tiehi \cpu.gpio.r_gpio_io[3]$_DFFE_PP__2828  (.L_HI(net2828));
 sg13g2_tiehi \cpu.gpio.r_gpio_o[0]$_DFFE_PP__2829  (.L_HI(net2829));
 sg13g2_tiehi \cpu.gpio.r_gpio_o[1]$_DFFE_PP__2830  (.L_HI(net2830));
 sg13g2_tiehi \cpu.gpio.r_gpio_o[2]$_DFFE_PP__2831  (.L_HI(net2831));
 sg13g2_tiehi \cpu.gpio.r_gpio_o[3]$_DFFE_PP__2832  (.L_HI(net2832));
 sg13g2_tiehi \cpu.gpio.r_gpio_o[4]$_DFFE_PP__2833  (.L_HI(net2833));
 sg13g2_tiehi \cpu.gpio.r_spi_miso_src[0][0]$_DFFE_PP__2834  (.L_HI(net2834));
 sg13g2_tiehi \cpu.gpio.r_spi_miso_src[0][1]$_DFFE_PP__2835  (.L_HI(net2835));
 sg13g2_tiehi \cpu.gpio.r_spi_miso_src[0][2]$_DFFE_PP__2836  (.L_HI(net2836));
 sg13g2_tiehi \cpu.gpio.r_spi_miso_src[0][3]$_DFFE_PP__2837  (.L_HI(net2837));
 sg13g2_tiehi \cpu.gpio.r_spi_miso_src[1][0]$_DFFE_PP__2838  (.L_HI(net2838));
 sg13g2_tiehi \cpu.gpio.r_spi_miso_src[1][1]$_DFFE_PP__2839  (.L_HI(net2839));
 sg13g2_tiehi \cpu.gpio.r_spi_miso_src[1][2]$_DFFE_PP__2840  (.L_HI(net2840));
 sg13g2_tiehi \cpu.gpio.r_spi_miso_src[1][3]$_DFFE_PP__2841  (.L_HI(net2841));
 sg13g2_tiehi \cpu.gpio.r_src_io[4][0]$_DFFE_PP__2842  (.L_HI(net2842));
 sg13g2_tiehi \cpu.gpio.r_src_io[4][1]$_DFFE_PP__2843  (.L_HI(net2843));
 sg13g2_tiehi \cpu.gpio.r_src_io[4][2]$_DFFE_PP__2844  (.L_HI(net2844));
 sg13g2_tiehi \cpu.gpio.r_src_io[4][3]$_DFFE_PP__2845  (.L_HI(net2845));
 sg13g2_tiehi \cpu.gpio.r_src_io[5][0]$_DFFE_PP__2846  (.L_HI(net2846));
 sg13g2_tiehi \cpu.gpio.r_src_io[5][1]$_DFFE_PP__2847  (.L_HI(net2847));
 sg13g2_tiehi \cpu.gpio.r_src_io[5][2]$_DFFE_PP__2848  (.L_HI(net2848));
 sg13g2_tiehi \cpu.gpio.r_src_io[5][3]$_DFFE_PP__2849  (.L_HI(net2849));
 sg13g2_tiehi \cpu.gpio.r_src_io[6][0]$_DFFE_PP__2850  (.L_HI(net2850));
 sg13g2_tiehi \cpu.gpio.r_src_io[6][1]$_DFFE_PP__2851  (.L_HI(net2851));
 sg13g2_tiehi \cpu.gpio.r_src_io[6][2]$_DFFE_PP__2852  (.L_HI(net2852));
 sg13g2_tiehi \cpu.gpio.r_src_io[6][3]$_DFFE_PP__2853  (.L_HI(net2853));
 sg13g2_tiehi \cpu.gpio.r_src_io[7][0]$_DFFE_PP__2854  (.L_HI(net2854));
 sg13g2_tiehi \cpu.gpio.r_src_io[7][1]$_DFFE_PP__2855  (.L_HI(net2855));
 sg13g2_tiehi \cpu.gpio.r_src_io[7][2]$_DFFE_PP__2856  (.L_HI(net2856));
 sg13g2_tiehi \cpu.gpio.r_src_io[7][3]$_DFFE_PP__2857  (.L_HI(net2857));
 sg13g2_tiehi \cpu.gpio.r_src_o[3][0]$_DFFE_PP__2858  (.L_HI(net2858));
 sg13g2_tiehi \cpu.gpio.r_src_o[3][1]$_DFFE_PP__2859  (.L_HI(net2859));
 sg13g2_tiehi \cpu.gpio.r_src_o[3][2]$_DFFE_PP__2860  (.L_HI(net2860));
 sg13g2_tiehi \cpu.gpio.r_src_o[3][3]$_DFFE_PP__2861  (.L_HI(net2861));
 sg13g2_tiehi \cpu.gpio.r_src_o[4][0]$_DFFE_PP__2862  (.L_HI(net2862));
 sg13g2_tiehi \cpu.gpio.r_src_o[4][1]$_DFFE_PP__2863  (.L_HI(net2863));
 sg13g2_tiehi \cpu.gpio.r_src_o[4][2]$_DFFE_PP__2864  (.L_HI(net2864));
 sg13g2_tiehi \cpu.gpio.r_src_o[4][3]$_DFFE_PP__2865  (.L_HI(net2865));
 sg13g2_tiehi \cpu.gpio.r_src_o[5][0]$_DFFE_PP__2866  (.L_HI(net2866));
 sg13g2_tiehi \cpu.gpio.r_src_o[5][1]$_DFFE_PP__2867  (.L_HI(net2867));
 sg13g2_tiehi \cpu.gpio.r_src_o[5][2]$_DFFE_PP__2868  (.L_HI(net2868));
 sg13g2_tiehi \cpu.gpio.r_src_o[5][3]$_DFFE_PP__2869  (.L_HI(net2869));
 sg13g2_tiehi \cpu.gpio.r_src_o[6][0]$_SDFFE_PN1P__2870  (.L_HI(net2870));
 sg13g2_tiehi \cpu.gpio.r_src_o[6][1]$_SDFFE_PN0P__2871  (.L_HI(net2871));
 sg13g2_tiehi \cpu.gpio.r_src_o[6][2]$_SDFFE_PN0P__2872  (.L_HI(net2872));
 sg13g2_tiehi \cpu.gpio.r_src_o[6][3]$_SDFFE_PN0P__2873  (.L_HI(net2873));
 sg13g2_tiehi \cpu.gpio.r_src_o[7][0]$_DFFE_PP__2874  (.L_HI(net2874));
 sg13g2_tiehi \cpu.gpio.r_src_o[7][1]$_DFFE_PP__2875  (.L_HI(net2875));
 sg13g2_tiehi \cpu.gpio.r_src_o[7][2]$_DFFE_PP__2876  (.L_HI(net2876));
 sg13g2_tiehi \cpu.gpio.r_src_o[7][3]$_DFFE_PP__2877  (.L_HI(net2877));
 sg13g2_tiehi \cpu.gpio.r_uart_rx_src[0]$_SDFFE_PN0P__2878  (.L_HI(net2878));
 sg13g2_tiehi \cpu.gpio.r_uart_rx_src[1]$_SDFFE_PN0P__2879  (.L_HI(net2879));
 sg13g2_tiehi \cpu.gpio.r_uart_rx_src[2]$_SDFFE_PN0P__2880  (.L_HI(net2880));
 sg13g2_tiehi \cpu.icache.r_data[0][0]$_DFFE_PP__2881  (.L_HI(net2881));
 sg13g2_tiehi \cpu.icache.r_data[0][10]$_DFFE_PP__2882  (.L_HI(net2882));
 sg13g2_tiehi \cpu.icache.r_data[0][11]$_DFFE_PP__2883  (.L_HI(net2883));
 sg13g2_tiehi \cpu.icache.r_data[0][12]$_DFFE_PP__2884  (.L_HI(net2884));
 sg13g2_tiehi \cpu.icache.r_data[0][13]$_DFFE_PP__2885  (.L_HI(net2885));
 sg13g2_tiehi \cpu.icache.r_data[0][14]$_DFFE_PP__2886  (.L_HI(net2886));
 sg13g2_tiehi \cpu.icache.r_data[0][15]$_DFFE_PP__2887  (.L_HI(net2887));
 sg13g2_tiehi \cpu.icache.r_data[0][16]$_DFFE_PP__2888  (.L_HI(net2888));
 sg13g2_tiehi \cpu.icache.r_data[0][17]$_DFFE_PP__2889  (.L_HI(net2889));
 sg13g2_tiehi \cpu.icache.r_data[0][18]$_DFFE_PP__2890  (.L_HI(net2890));
 sg13g2_tiehi \cpu.icache.r_data[0][19]$_DFFE_PP__2891  (.L_HI(net2891));
 sg13g2_tiehi \cpu.icache.r_data[0][1]$_DFFE_PP__2892  (.L_HI(net2892));
 sg13g2_tiehi \cpu.icache.r_data[0][20]$_DFFE_PP__2893  (.L_HI(net2893));
 sg13g2_tiehi \cpu.icache.r_data[0][21]$_DFFE_PP__2894  (.L_HI(net2894));
 sg13g2_tiehi \cpu.icache.r_data[0][22]$_DFFE_PP__2895  (.L_HI(net2895));
 sg13g2_tiehi \cpu.icache.r_data[0][23]$_DFFE_PP__2896  (.L_HI(net2896));
 sg13g2_tiehi \cpu.icache.r_data[0][24]$_DFFE_PP__2897  (.L_HI(net2897));
 sg13g2_tiehi \cpu.icache.r_data[0][25]$_DFFE_PP__2898  (.L_HI(net2898));
 sg13g2_tiehi \cpu.icache.r_data[0][26]$_DFFE_PP__2899  (.L_HI(net2899));
 sg13g2_tiehi \cpu.icache.r_data[0][27]$_DFFE_PP__2900  (.L_HI(net2900));
 sg13g2_tiehi \cpu.icache.r_data[0][28]$_DFFE_PP__2901  (.L_HI(net2901));
 sg13g2_tiehi \cpu.icache.r_data[0][29]$_DFFE_PP__2902  (.L_HI(net2902));
 sg13g2_tiehi \cpu.icache.r_data[0][2]$_DFFE_PP__2903  (.L_HI(net2903));
 sg13g2_tiehi \cpu.icache.r_data[0][30]$_DFFE_PP__2904  (.L_HI(net2904));
 sg13g2_tiehi \cpu.icache.r_data[0][31]$_DFFE_PP__2905  (.L_HI(net2905));
 sg13g2_tiehi \cpu.icache.r_data[0][3]$_DFFE_PP__2906  (.L_HI(net2906));
 sg13g2_tiehi \cpu.icache.r_data[0][4]$_DFFE_PP__2907  (.L_HI(net2907));
 sg13g2_tiehi \cpu.icache.r_data[0][5]$_DFFE_PP__2908  (.L_HI(net2908));
 sg13g2_tiehi \cpu.icache.r_data[0][6]$_DFFE_PP__2909  (.L_HI(net2909));
 sg13g2_tiehi \cpu.icache.r_data[0][7]$_DFFE_PP__2910  (.L_HI(net2910));
 sg13g2_tiehi \cpu.icache.r_data[0][8]$_DFFE_PP__2911  (.L_HI(net2911));
 sg13g2_tiehi \cpu.icache.r_data[0][9]$_DFFE_PP__2912  (.L_HI(net2912));
 sg13g2_tiehi \cpu.icache.r_data[1][0]$_DFFE_PP__2913  (.L_HI(net2913));
 sg13g2_tiehi \cpu.icache.r_data[1][10]$_DFFE_PP__2914  (.L_HI(net2914));
 sg13g2_tiehi \cpu.icache.r_data[1][11]$_DFFE_PP__2915  (.L_HI(net2915));
 sg13g2_tiehi \cpu.icache.r_data[1][12]$_DFFE_PP__2916  (.L_HI(net2916));
 sg13g2_tiehi \cpu.icache.r_data[1][13]$_DFFE_PP__2917  (.L_HI(net2917));
 sg13g2_tiehi \cpu.icache.r_data[1][14]$_DFFE_PP__2918  (.L_HI(net2918));
 sg13g2_tiehi \cpu.icache.r_data[1][15]$_DFFE_PP__2919  (.L_HI(net2919));
 sg13g2_tiehi \cpu.icache.r_data[1][16]$_DFFE_PP__2920  (.L_HI(net2920));
 sg13g2_tiehi \cpu.icache.r_data[1][17]$_DFFE_PP__2921  (.L_HI(net2921));
 sg13g2_tiehi \cpu.icache.r_data[1][18]$_DFFE_PP__2922  (.L_HI(net2922));
 sg13g2_tiehi \cpu.icache.r_data[1][19]$_DFFE_PP__2923  (.L_HI(net2923));
 sg13g2_tiehi \cpu.icache.r_data[1][1]$_DFFE_PP__2924  (.L_HI(net2924));
 sg13g2_tiehi \cpu.icache.r_data[1][20]$_DFFE_PP__2925  (.L_HI(net2925));
 sg13g2_tiehi \cpu.icache.r_data[1][21]$_DFFE_PP__2926  (.L_HI(net2926));
 sg13g2_tiehi \cpu.icache.r_data[1][22]$_DFFE_PP__2927  (.L_HI(net2927));
 sg13g2_tiehi \cpu.icache.r_data[1][23]$_DFFE_PP__2928  (.L_HI(net2928));
 sg13g2_tiehi \cpu.icache.r_data[1][24]$_DFFE_PP__2929  (.L_HI(net2929));
 sg13g2_tiehi \cpu.icache.r_data[1][25]$_DFFE_PP__2930  (.L_HI(net2930));
 sg13g2_tiehi \cpu.icache.r_data[1][26]$_DFFE_PP__2931  (.L_HI(net2931));
 sg13g2_tiehi \cpu.icache.r_data[1][27]$_DFFE_PP__2932  (.L_HI(net2932));
 sg13g2_tiehi \cpu.icache.r_data[1][28]$_DFFE_PP__2933  (.L_HI(net2933));
 sg13g2_tiehi \cpu.icache.r_data[1][29]$_DFFE_PP__2934  (.L_HI(net2934));
 sg13g2_tiehi \cpu.icache.r_data[1][2]$_DFFE_PP__2935  (.L_HI(net2935));
 sg13g2_tiehi \cpu.icache.r_data[1][30]$_DFFE_PP__2936  (.L_HI(net2936));
 sg13g2_tiehi \cpu.icache.r_data[1][31]$_DFFE_PP__2937  (.L_HI(net2937));
 sg13g2_tiehi \cpu.icache.r_data[1][3]$_DFFE_PP__2938  (.L_HI(net2938));
 sg13g2_tiehi \cpu.icache.r_data[1][4]$_DFFE_PP__2939  (.L_HI(net2939));
 sg13g2_tiehi \cpu.icache.r_data[1][5]$_DFFE_PP__2940  (.L_HI(net2940));
 sg13g2_tiehi \cpu.icache.r_data[1][6]$_DFFE_PP__2941  (.L_HI(net2941));
 sg13g2_tiehi \cpu.icache.r_data[1][7]$_DFFE_PP__2942  (.L_HI(net2942));
 sg13g2_tiehi \cpu.icache.r_data[1][8]$_DFFE_PP__2943  (.L_HI(net2943));
 sg13g2_tiehi \cpu.icache.r_data[1][9]$_DFFE_PP__2944  (.L_HI(net2944));
 sg13g2_tiehi \cpu.icache.r_data[2][0]$_DFFE_PP__2945  (.L_HI(net2945));
 sg13g2_tiehi \cpu.icache.r_data[2][10]$_DFFE_PP__2946  (.L_HI(net2946));
 sg13g2_tiehi \cpu.icache.r_data[2][11]$_DFFE_PP__2947  (.L_HI(net2947));
 sg13g2_tiehi \cpu.icache.r_data[2][12]$_DFFE_PP__2948  (.L_HI(net2948));
 sg13g2_tiehi \cpu.icache.r_data[2][13]$_DFFE_PP__2949  (.L_HI(net2949));
 sg13g2_tiehi \cpu.icache.r_data[2][14]$_DFFE_PP__2950  (.L_HI(net2950));
 sg13g2_tiehi \cpu.icache.r_data[2][15]$_DFFE_PP__2951  (.L_HI(net2951));
 sg13g2_tiehi \cpu.icache.r_data[2][16]$_DFFE_PP__2952  (.L_HI(net2952));
 sg13g2_tiehi \cpu.icache.r_data[2][17]$_DFFE_PP__2953  (.L_HI(net2953));
 sg13g2_tiehi \cpu.icache.r_data[2][18]$_DFFE_PP__2954  (.L_HI(net2954));
 sg13g2_tiehi \cpu.icache.r_data[2][19]$_DFFE_PP__2955  (.L_HI(net2955));
 sg13g2_tiehi \cpu.icache.r_data[2][1]$_DFFE_PP__2956  (.L_HI(net2956));
 sg13g2_tiehi \cpu.icache.r_data[2][20]$_DFFE_PP__2957  (.L_HI(net2957));
 sg13g2_tiehi \cpu.icache.r_data[2][21]$_DFFE_PP__2958  (.L_HI(net2958));
 sg13g2_tiehi \cpu.icache.r_data[2][22]$_DFFE_PP__2959  (.L_HI(net2959));
 sg13g2_tiehi \cpu.icache.r_data[2][23]$_DFFE_PP__2960  (.L_HI(net2960));
 sg13g2_tiehi \cpu.icache.r_data[2][24]$_DFFE_PP__2961  (.L_HI(net2961));
 sg13g2_tiehi \cpu.icache.r_data[2][25]$_DFFE_PP__2962  (.L_HI(net2962));
 sg13g2_tiehi \cpu.icache.r_data[2][26]$_DFFE_PP__2963  (.L_HI(net2963));
 sg13g2_tiehi \cpu.icache.r_data[2][27]$_DFFE_PP__2964  (.L_HI(net2964));
 sg13g2_tiehi \cpu.icache.r_data[2][28]$_DFFE_PP__2965  (.L_HI(net2965));
 sg13g2_tiehi \cpu.icache.r_data[2][29]$_DFFE_PP__2966  (.L_HI(net2966));
 sg13g2_tiehi \cpu.icache.r_data[2][2]$_DFFE_PP__2967  (.L_HI(net2967));
 sg13g2_tiehi \cpu.icache.r_data[2][30]$_DFFE_PP__2968  (.L_HI(net2968));
 sg13g2_tiehi \cpu.icache.r_data[2][31]$_DFFE_PP__2969  (.L_HI(net2969));
 sg13g2_tiehi \cpu.icache.r_data[2][3]$_DFFE_PP__2970  (.L_HI(net2970));
 sg13g2_tiehi \cpu.icache.r_data[2][4]$_DFFE_PP__2971  (.L_HI(net2971));
 sg13g2_tiehi \cpu.icache.r_data[2][5]$_DFFE_PP__2972  (.L_HI(net2972));
 sg13g2_tiehi \cpu.icache.r_data[2][6]$_DFFE_PP__2973  (.L_HI(net2973));
 sg13g2_tiehi \cpu.icache.r_data[2][7]$_DFFE_PP__2974  (.L_HI(net2974));
 sg13g2_tiehi \cpu.icache.r_data[2][8]$_DFFE_PP__2975  (.L_HI(net2975));
 sg13g2_tiehi \cpu.icache.r_data[2][9]$_DFFE_PP__2976  (.L_HI(net2976));
 sg13g2_tiehi \cpu.icache.r_data[3][0]$_DFFE_PP__2977  (.L_HI(net2977));
 sg13g2_tiehi \cpu.icache.r_data[3][10]$_DFFE_PP__2978  (.L_HI(net2978));
 sg13g2_tiehi \cpu.icache.r_data[3][11]$_DFFE_PP__2979  (.L_HI(net2979));
 sg13g2_tiehi \cpu.icache.r_data[3][12]$_DFFE_PP__2980  (.L_HI(net2980));
 sg13g2_tiehi \cpu.icache.r_data[3][13]$_DFFE_PP__2981  (.L_HI(net2981));
 sg13g2_tiehi \cpu.icache.r_data[3][14]$_DFFE_PP__2982  (.L_HI(net2982));
 sg13g2_tiehi \cpu.icache.r_data[3][15]$_DFFE_PP__2983  (.L_HI(net2983));
 sg13g2_tiehi \cpu.icache.r_data[3][16]$_DFFE_PP__2984  (.L_HI(net2984));
 sg13g2_tiehi \cpu.icache.r_data[3][17]$_DFFE_PP__2985  (.L_HI(net2985));
 sg13g2_tiehi \cpu.icache.r_data[3][18]$_DFFE_PP__2986  (.L_HI(net2986));
 sg13g2_tiehi \cpu.icache.r_data[3][19]$_DFFE_PP__2987  (.L_HI(net2987));
 sg13g2_tiehi \cpu.icache.r_data[3][1]$_DFFE_PP__2988  (.L_HI(net2988));
 sg13g2_tiehi \cpu.icache.r_data[3][20]$_DFFE_PP__2989  (.L_HI(net2989));
 sg13g2_tiehi \cpu.icache.r_data[3][21]$_DFFE_PP__2990  (.L_HI(net2990));
 sg13g2_tiehi \cpu.icache.r_data[3][22]$_DFFE_PP__2991  (.L_HI(net2991));
 sg13g2_tiehi \cpu.icache.r_data[3][23]$_DFFE_PP__2992  (.L_HI(net2992));
 sg13g2_tiehi \cpu.icache.r_data[3][24]$_DFFE_PP__2993  (.L_HI(net2993));
 sg13g2_tiehi \cpu.icache.r_data[3][25]$_DFFE_PP__2994  (.L_HI(net2994));
 sg13g2_tiehi \cpu.icache.r_data[3][26]$_DFFE_PP__2995  (.L_HI(net2995));
 sg13g2_tiehi \cpu.icache.r_data[3][27]$_DFFE_PP__2996  (.L_HI(net2996));
 sg13g2_tiehi \cpu.icache.r_data[3][28]$_DFFE_PP__2997  (.L_HI(net2997));
 sg13g2_tiehi \cpu.icache.r_data[3][29]$_DFFE_PP__2998  (.L_HI(net2998));
 sg13g2_tiehi \cpu.icache.r_data[3][2]$_DFFE_PP__2999  (.L_HI(net2999));
 sg13g2_tiehi \cpu.icache.r_data[3][30]$_DFFE_PP__3000  (.L_HI(net3000));
 sg13g2_tiehi \cpu.icache.r_data[3][31]$_DFFE_PP__3001  (.L_HI(net3001));
 sg13g2_tiehi \cpu.icache.r_data[3][3]$_DFFE_PP__3002  (.L_HI(net3002));
 sg13g2_tiehi \cpu.icache.r_data[3][4]$_DFFE_PP__3003  (.L_HI(net3003));
 sg13g2_tiehi \cpu.icache.r_data[3][5]$_DFFE_PP__3004  (.L_HI(net3004));
 sg13g2_tiehi \cpu.icache.r_data[3][6]$_DFFE_PP__3005  (.L_HI(net3005));
 sg13g2_tiehi \cpu.icache.r_data[3][7]$_DFFE_PP__3006  (.L_HI(net3006));
 sg13g2_tiehi \cpu.icache.r_data[3][8]$_DFFE_PP__3007  (.L_HI(net3007));
 sg13g2_tiehi \cpu.icache.r_data[3][9]$_DFFE_PP__3008  (.L_HI(net3008));
 sg13g2_tiehi \cpu.icache.r_data[4][0]$_DFFE_PP__3009  (.L_HI(net3009));
 sg13g2_tiehi \cpu.icache.r_data[4][10]$_DFFE_PP__3010  (.L_HI(net3010));
 sg13g2_tiehi \cpu.icache.r_data[4][11]$_DFFE_PP__3011  (.L_HI(net3011));
 sg13g2_tiehi \cpu.icache.r_data[4][12]$_DFFE_PP__3012  (.L_HI(net3012));
 sg13g2_tiehi \cpu.icache.r_data[4][13]$_DFFE_PP__3013  (.L_HI(net3013));
 sg13g2_tiehi \cpu.icache.r_data[4][14]$_DFFE_PP__3014  (.L_HI(net3014));
 sg13g2_tiehi \cpu.icache.r_data[4][15]$_DFFE_PP__3015  (.L_HI(net3015));
 sg13g2_tiehi \cpu.icache.r_data[4][16]$_DFFE_PP__3016  (.L_HI(net3016));
 sg13g2_tiehi \cpu.icache.r_data[4][17]$_DFFE_PP__3017  (.L_HI(net3017));
 sg13g2_tiehi \cpu.icache.r_data[4][18]$_DFFE_PP__3018  (.L_HI(net3018));
 sg13g2_tiehi \cpu.icache.r_data[4][19]$_DFFE_PP__3019  (.L_HI(net3019));
 sg13g2_tiehi \cpu.icache.r_data[4][1]$_DFFE_PP__3020  (.L_HI(net3020));
 sg13g2_tiehi \cpu.icache.r_data[4][20]$_DFFE_PP__3021  (.L_HI(net3021));
 sg13g2_tiehi \cpu.icache.r_data[4][21]$_DFFE_PP__3022  (.L_HI(net3022));
 sg13g2_tiehi \cpu.icache.r_data[4][22]$_DFFE_PP__3023  (.L_HI(net3023));
 sg13g2_tiehi \cpu.icache.r_data[4][23]$_DFFE_PP__3024  (.L_HI(net3024));
 sg13g2_tiehi \cpu.icache.r_data[4][24]$_DFFE_PP__3025  (.L_HI(net3025));
 sg13g2_tiehi \cpu.icache.r_data[4][25]$_DFFE_PP__3026  (.L_HI(net3026));
 sg13g2_tiehi \cpu.icache.r_data[4][26]$_DFFE_PP__3027  (.L_HI(net3027));
 sg13g2_tiehi \cpu.icache.r_data[4][27]$_DFFE_PP__3028  (.L_HI(net3028));
 sg13g2_tiehi \cpu.icache.r_data[4][28]$_DFFE_PP__3029  (.L_HI(net3029));
 sg13g2_tiehi \cpu.icache.r_data[4][29]$_DFFE_PP__3030  (.L_HI(net3030));
 sg13g2_tiehi \cpu.icache.r_data[4][2]$_DFFE_PP__3031  (.L_HI(net3031));
 sg13g2_tiehi \cpu.icache.r_data[4][30]$_DFFE_PP__3032  (.L_HI(net3032));
 sg13g2_tiehi \cpu.icache.r_data[4][31]$_DFFE_PP__3033  (.L_HI(net3033));
 sg13g2_tiehi \cpu.icache.r_data[4][3]$_DFFE_PP__3034  (.L_HI(net3034));
 sg13g2_tiehi \cpu.icache.r_data[4][4]$_DFFE_PP__3035  (.L_HI(net3035));
 sg13g2_tiehi \cpu.icache.r_data[4][5]$_DFFE_PP__3036  (.L_HI(net3036));
 sg13g2_tiehi \cpu.icache.r_data[4][6]$_DFFE_PP__3037  (.L_HI(net3037));
 sg13g2_tiehi \cpu.icache.r_data[4][7]$_DFFE_PP__3038  (.L_HI(net3038));
 sg13g2_tiehi \cpu.icache.r_data[4][8]$_DFFE_PP__3039  (.L_HI(net3039));
 sg13g2_tiehi \cpu.icache.r_data[4][9]$_DFFE_PP__3040  (.L_HI(net3040));
 sg13g2_tiehi \cpu.icache.r_data[5][0]$_DFFE_PP__3041  (.L_HI(net3041));
 sg13g2_tiehi \cpu.icache.r_data[5][10]$_DFFE_PP__3042  (.L_HI(net3042));
 sg13g2_tiehi \cpu.icache.r_data[5][11]$_DFFE_PP__3043  (.L_HI(net3043));
 sg13g2_tiehi \cpu.icache.r_data[5][12]$_DFFE_PP__3044  (.L_HI(net3044));
 sg13g2_tiehi \cpu.icache.r_data[5][13]$_DFFE_PP__3045  (.L_HI(net3045));
 sg13g2_tiehi \cpu.icache.r_data[5][14]$_DFFE_PP__3046  (.L_HI(net3046));
 sg13g2_tiehi \cpu.icache.r_data[5][15]$_DFFE_PP__3047  (.L_HI(net3047));
 sg13g2_tiehi \cpu.icache.r_data[5][16]$_DFFE_PP__3048  (.L_HI(net3048));
 sg13g2_tiehi \cpu.icache.r_data[5][17]$_DFFE_PP__3049  (.L_HI(net3049));
 sg13g2_tiehi \cpu.icache.r_data[5][18]$_DFFE_PP__3050  (.L_HI(net3050));
 sg13g2_tiehi \cpu.icache.r_data[5][19]$_DFFE_PP__3051  (.L_HI(net3051));
 sg13g2_tiehi \cpu.icache.r_data[5][1]$_DFFE_PP__3052  (.L_HI(net3052));
 sg13g2_tiehi \cpu.icache.r_data[5][20]$_DFFE_PP__3053  (.L_HI(net3053));
 sg13g2_tiehi \cpu.icache.r_data[5][21]$_DFFE_PP__3054  (.L_HI(net3054));
 sg13g2_tiehi \cpu.icache.r_data[5][22]$_DFFE_PP__3055  (.L_HI(net3055));
 sg13g2_tiehi \cpu.icache.r_data[5][23]$_DFFE_PP__3056  (.L_HI(net3056));
 sg13g2_tiehi \cpu.icache.r_data[5][24]$_DFFE_PP__3057  (.L_HI(net3057));
 sg13g2_tiehi \cpu.icache.r_data[5][25]$_DFFE_PP__3058  (.L_HI(net3058));
 sg13g2_tiehi \cpu.icache.r_data[5][26]$_DFFE_PP__3059  (.L_HI(net3059));
 sg13g2_tiehi \cpu.icache.r_data[5][27]$_DFFE_PP__3060  (.L_HI(net3060));
 sg13g2_tiehi \cpu.icache.r_data[5][28]$_DFFE_PP__3061  (.L_HI(net3061));
 sg13g2_tiehi \cpu.icache.r_data[5][29]$_DFFE_PP__3062  (.L_HI(net3062));
 sg13g2_tiehi \cpu.icache.r_data[5][2]$_DFFE_PP__3063  (.L_HI(net3063));
 sg13g2_tiehi \cpu.icache.r_data[5][30]$_DFFE_PP__3064  (.L_HI(net3064));
 sg13g2_tiehi \cpu.icache.r_data[5][31]$_DFFE_PP__3065  (.L_HI(net3065));
 sg13g2_tiehi \cpu.icache.r_data[5][3]$_DFFE_PP__3066  (.L_HI(net3066));
 sg13g2_tiehi \cpu.icache.r_data[5][4]$_DFFE_PP__3067  (.L_HI(net3067));
 sg13g2_tiehi \cpu.icache.r_data[5][5]$_DFFE_PP__3068  (.L_HI(net3068));
 sg13g2_tiehi \cpu.icache.r_data[5][6]$_DFFE_PP__3069  (.L_HI(net3069));
 sg13g2_tiehi \cpu.icache.r_data[5][7]$_DFFE_PP__3070  (.L_HI(net3070));
 sg13g2_tiehi \cpu.icache.r_data[5][8]$_DFFE_PP__3071  (.L_HI(net3071));
 sg13g2_tiehi \cpu.icache.r_data[5][9]$_DFFE_PP__3072  (.L_HI(net3072));
 sg13g2_tiehi \cpu.icache.r_data[6][0]$_DFFE_PP__3073  (.L_HI(net3073));
 sg13g2_tiehi \cpu.icache.r_data[6][10]$_DFFE_PP__3074  (.L_HI(net3074));
 sg13g2_tiehi \cpu.icache.r_data[6][11]$_DFFE_PP__3075  (.L_HI(net3075));
 sg13g2_tiehi \cpu.icache.r_data[6][12]$_DFFE_PP__3076  (.L_HI(net3076));
 sg13g2_tiehi \cpu.icache.r_data[6][13]$_DFFE_PP__3077  (.L_HI(net3077));
 sg13g2_tiehi \cpu.icache.r_data[6][14]$_DFFE_PP__3078  (.L_HI(net3078));
 sg13g2_tiehi \cpu.icache.r_data[6][15]$_DFFE_PP__3079  (.L_HI(net3079));
 sg13g2_tiehi \cpu.icache.r_data[6][16]$_DFFE_PP__3080  (.L_HI(net3080));
 sg13g2_tiehi \cpu.icache.r_data[6][17]$_DFFE_PP__3081  (.L_HI(net3081));
 sg13g2_tiehi \cpu.icache.r_data[6][18]$_DFFE_PP__3082  (.L_HI(net3082));
 sg13g2_tiehi \cpu.icache.r_data[6][19]$_DFFE_PP__3083  (.L_HI(net3083));
 sg13g2_tiehi \cpu.icache.r_data[6][1]$_DFFE_PP__3084  (.L_HI(net3084));
 sg13g2_tiehi \cpu.icache.r_data[6][20]$_DFFE_PP__3085  (.L_HI(net3085));
 sg13g2_tiehi \cpu.icache.r_data[6][21]$_DFFE_PP__3086  (.L_HI(net3086));
 sg13g2_tiehi \cpu.icache.r_data[6][22]$_DFFE_PP__3087  (.L_HI(net3087));
 sg13g2_tiehi \cpu.icache.r_data[6][23]$_DFFE_PP__3088  (.L_HI(net3088));
 sg13g2_tiehi \cpu.icache.r_data[6][24]$_DFFE_PP__3089  (.L_HI(net3089));
 sg13g2_tiehi \cpu.icache.r_data[6][25]$_DFFE_PP__3090  (.L_HI(net3090));
 sg13g2_tiehi \cpu.icache.r_data[6][26]$_DFFE_PP__3091  (.L_HI(net3091));
 sg13g2_tiehi \cpu.icache.r_data[6][27]$_DFFE_PP__3092  (.L_HI(net3092));
 sg13g2_tiehi \cpu.icache.r_data[6][28]$_DFFE_PP__3093  (.L_HI(net3093));
 sg13g2_tiehi \cpu.icache.r_data[6][29]$_DFFE_PP__3094  (.L_HI(net3094));
 sg13g2_tiehi \cpu.icache.r_data[6][2]$_DFFE_PP__3095  (.L_HI(net3095));
 sg13g2_tiehi \cpu.icache.r_data[6][30]$_DFFE_PP__3096  (.L_HI(net3096));
 sg13g2_tiehi \cpu.icache.r_data[6][31]$_DFFE_PP__3097  (.L_HI(net3097));
 sg13g2_tiehi \cpu.icache.r_data[6][3]$_DFFE_PP__3098  (.L_HI(net3098));
 sg13g2_tiehi \cpu.icache.r_data[6][4]$_DFFE_PP__3099  (.L_HI(net3099));
 sg13g2_tiehi \cpu.icache.r_data[6][5]$_DFFE_PP__3100  (.L_HI(net3100));
 sg13g2_tiehi \cpu.icache.r_data[6][6]$_DFFE_PP__3101  (.L_HI(net3101));
 sg13g2_tiehi \cpu.icache.r_data[6][7]$_DFFE_PP__3102  (.L_HI(net3102));
 sg13g2_tiehi \cpu.icache.r_data[6][8]$_DFFE_PP__3103  (.L_HI(net3103));
 sg13g2_tiehi \cpu.icache.r_data[6][9]$_DFFE_PP__3104  (.L_HI(net3104));
 sg13g2_tiehi \cpu.icache.r_data[7][0]$_DFFE_PP__3105  (.L_HI(net3105));
 sg13g2_tiehi \cpu.icache.r_data[7][10]$_DFFE_PP__3106  (.L_HI(net3106));
 sg13g2_tiehi \cpu.icache.r_data[7][11]$_DFFE_PP__3107  (.L_HI(net3107));
 sg13g2_tiehi \cpu.icache.r_data[7][12]$_DFFE_PP__3108  (.L_HI(net3108));
 sg13g2_tiehi \cpu.icache.r_data[7][13]$_DFFE_PP__3109  (.L_HI(net3109));
 sg13g2_tiehi \cpu.icache.r_data[7][14]$_DFFE_PP__3110  (.L_HI(net3110));
 sg13g2_tiehi \cpu.icache.r_data[7][15]$_DFFE_PP__3111  (.L_HI(net3111));
 sg13g2_tiehi \cpu.icache.r_data[7][16]$_DFFE_PP__3112  (.L_HI(net3112));
 sg13g2_tiehi \cpu.icache.r_data[7][17]$_DFFE_PP__3113  (.L_HI(net3113));
 sg13g2_tiehi \cpu.icache.r_data[7][18]$_DFFE_PP__3114  (.L_HI(net3114));
 sg13g2_tiehi \cpu.icache.r_data[7][19]$_DFFE_PP__3115  (.L_HI(net3115));
 sg13g2_tiehi \cpu.icache.r_data[7][1]$_DFFE_PP__3116  (.L_HI(net3116));
 sg13g2_tiehi \cpu.icache.r_data[7][20]$_DFFE_PP__3117  (.L_HI(net3117));
 sg13g2_tiehi \cpu.icache.r_data[7][21]$_DFFE_PP__3118  (.L_HI(net3118));
 sg13g2_tiehi \cpu.icache.r_data[7][22]$_DFFE_PP__3119  (.L_HI(net3119));
 sg13g2_tiehi \cpu.icache.r_data[7][23]$_DFFE_PP__3120  (.L_HI(net3120));
 sg13g2_tiehi \cpu.icache.r_data[7][24]$_DFFE_PP__3121  (.L_HI(net3121));
 sg13g2_tiehi \cpu.icache.r_data[7][25]$_DFFE_PP__3122  (.L_HI(net3122));
 sg13g2_tiehi \cpu.icache.r_data[7][26]$_DFFE_PP__3123  (.L_HI(net3123));
 sg13g2_tiehi \cpu.icache.r_data[7][27]$_DFFE_PP__3124  (.L_HI(net3124));
 sg13g2_tiehi \cpu.icache.r_data[7][28]$_DFFE_PP__3125  (.L_HI(net3125));
 sg13g2_tiehi \cpu.icache.r_data[7][29]$_DFFE_PP__3126  (.L_HI(net3126));
 sg13g2_tiehi \cpu.icache.r_data[7][2]$_DFFE_PP__3127  (.L_HI(net3127));
 sg13g2_tiehi \cpu.icache.r_data[7][30]$_DFFE_PP__3128  (.L_HI(net3128));
 sg13g2_tiehi \cpu.icache.r_data[7][31]$_DFFE_PP__3129  (.L_HI(net3129));
 sg13g2_tiehi \cpu.icache.r_data[7][3]$_DFFE_PP__3130  (.L_HI(net3130));
 sg13g2_tiehi \cpu.icache.r_data[7][4]$_DFFE_PP__3131  (.L_HI(net3131));
 sg13g2_tiehi \cpu.icache.r_data[7][5]$_DFFE_PP__3132  (.L_HI(net3132));
 sg13g2_tiehi \cpu.icache.r_data[7][6]$_DFFE_PP__3133  (.L_HI(net3133));
 sg13g2_tiehi \cpu.icache.r_data[7][7]$_DFFE_PP__3134  (.L_HI(net3134));
 sg13g2_tiehi \cpu.icache.r_data[7][8]$_DFFE_PP__3135  (.L_HI(net3135));
 sg13g2_tiehi \cpu.icache.r_data[7][9]$_DFFE_PP__3136  (.L_HI(net3136));
 sg13g2_tiehi \cpu.icache.r_offset[0]$_SDFF_PN0__3137  (.L_HI(net3137));
 sg13g2_tiehi \cpu.icache.r_offset[1]$_SDFF_PN0__3138  (.L_HI(net3138));
 sg13g2_tiehi \cpu.icache.r_offset[2]$_SDFF_PN0__3139  (.L_HI(net3139));
 sg13g2_tiehi \cpu.icache.r_tag[0][0]$_DFFE_PP__3140  (.L_HI(net3140));
 sg13g2_tiehi \cpu.icache.r_tag[0][10]$_DFFE_PP__3141  (.L_HI(net3141));
 sg13g2_tiehi \cpu.icache.r_tag[0][11]$_DFFE_PP__3142  (.L_HI(net3142));
 sg13g2_tiehi \cpu.icache.r_tag[0][12]$_DFFE_PP__3143  (.L_HI(net3143));
 sg13g2_tiehi \cpu.icache.r_tag[0][13]$_DFFE_PP__3144  (.L_HI(net3144));
 sg13g2_tiehi \cpu.icache.r_tag[0][14]$_DFFE_PP__3145  (.L_HI(net3145));
 sg13g2_tiehi \cpu.icache.r_tag[0][15]$_DFFE_PP__3146  (.L_HI(net3146));
 sg13g2_tiehi \cpu.icache.r_tag[0][16]$_DFFE_PP__3147  (.L_HI(net3147));
 sg13g2_tiehi \cpu.icache.r_tag[0][17]$_DFFE_PP__3148  (.L_HI(net3148));
 sg13g2_tiehi \cpu.icache.r_tag[0][18]$_DFFE_PP__3149  (.L_HI(net3149));
 sg13g2_tiehi \cpu.icache.r_tag[0][1]$_DFFE_PP__3150  (.L_HI(net3150));
 sg13g2_tiehi \cpu.icache.r_tag[0][2]$_DFFE_PP__3151  (.L_HI(net3151));
 sg13g2_tiehi \cpu.icache.r_tag[0][3]$_DFFE_PP__3152  (.L_HI(net3152));
 sg13g2_tiehi \cpu.icache.r_tag[0][4]$_DFFE_PP__3153  (.L_HI(net3153));
 sg13g2_tiehi \cpu.icache.r_tag[0][5]$_DFFE_PP__3154  (.L_HI(net3154));
 sg13g2_tiehi \cpu.icache.r_tag[0][6]$_DFFE_PP__3155  (.L_HI(net3155));
 sg13g2_tiehi \cpu.icache.r_tag[0][7]$_DFFE_PP__3156  (.L_HI(net3156));
 sg13g2_tiehi \cpu.icache.r_tag[0][8]$_DFFE_PP__3157  (.L_HI(net3157));
 sg13g2_tiehi \cpu.icache.r_tag[0][9]$_DFFE_PP__3158  (.L_HI(net3158));
 sg13g2_tiehi \cpu.icache.r_tag[1][0]$_DFFE_PP__3159  (.L_HI(net3159));
 sg13g2_tiehi \cpu.icache.r_tag[1][10]$_DFFE_PP__3160  (.L_HI(net3160));
 sg13g2_tiehi \cpu.icache.r_tag[1][11]$_DFFE_PP__3161  (.L_HI(net3161));
 sg13g2_tiehi \cpu.icache.r_tag[1][12]$_DFFE_PP__3162  (.L_HI(net3162));
 sg13g2_tiehi \cpu.icache.r_tag[1][13]$_DFFE_PP__3163  (.L_HI(net3163));
 sg13g2_tiehi \cpu.icache.r_tag[1][14]$_DFFE_PP__3164  (.L_HI(net3164));
 sg13g2_tiehi \cpu.icache.r_tag[1][15]$_DFFE_PP__3165  (.L_HI(net3165));
 sg13g2_tiehi \cpu.icache.r_tag[1][16]$_DFFE_PP__3166  (.L_HI(net3166));
 sg13g2_tiehi \cpu.icache.r_tag[1][17]$_DFFE_PP__3167  (.L_HI(net3167));
 sg13g2_tiehi \cpu.icache.r_tag[1][18]$_DFFE_PP__3168  (.L_HI(net3168));
 sg13g2_tiehi \cpu.icache.r_tag[1][1]$_DFFE_PP__3169  (.L_HI(net3169));
 sg13g2_tiehi \cpu.icache.r_tag[1][2]$_DFFE_PP__3170  (.L_HI(net3170));
 sg13g2_tiehi \cpu.icache.r_tag[1][3]$_DFFE_PP__3171  (.L_HI(net3171));
 sg13g2_tiehi \cpu.icache.r_tag[1][4]$_DFFE_PP__3172  (.L_HI(net3172));
 sg13g2_tiehi \cpu.icache.r_tag[1][5]$_DFFE_PP__3173  (.L_HI(net3173));
 sg13g2_tiehi \cpu.icache.r_tag[1][6]$_DFFE_PP__3174  (.L_HI(net3174));
 sg13g2_tiehi \cpu.icache.r_tag[1][7]$_DFFE_PP__3175  (.L_HI(net3175));
 sg13g2_tiehi \cpu.icache.r_tag[1][8]$_DFFE_PP__3176  (.L_HI(net3176));
 sg13g2_tiehi \cpu.icache.r_tag[1][9]$_DFFE_PP__3177  (.L_HI(net3177));
 sg13g2_tiehi \cpu.icache.r_tag[2][0]$_DFFE_PP__3178  (.L_HI(net3178));
 sg13g2_tiehi \cpu.icache.r_tag[2][10]$_DFFE_PP__3179  (.L_HI(net3179));
 sg13g2_tiehi \cpu.icache.r_tag[2][11]$_DFFE_PP__3180  (.L_HI(net3180));
 sg13g2_tiehi \cpu.icache.r_tag[2][12]$_DFFE_PP__3181  (.L_HI(net3181));
 sg13g2_tiehi \cpu.icache.r_tag[2][13]$_DFFE_PP__3182  (.L_HI(net3182));
 sg13g2_tiehi \cpu.icache.r_tag[2][14]$_DFFE_PP__3183  (.L_HI(net3183));
 sg13g2_tiehi \cpu.icache.r_tag[2][15]$_DFFE_PP__3184  (.L_HI(net3184));
 sg13g2_tiehi \cpu.icache.r_tag[2][16]$_DFFE_PP__3185  (.L_HI(net3185));
 sg13g2_tiehi \cpu.icache.r_tag[2][17]$_DFFE_PP__3186  (.L_HI(net3186));
 sg13g2_tiehi \cpu.icache.r_tag[2][18]$_DFFE_PP__3187  (.L_HI(net3187));
 sg13g2_tiehi \cpu.icache.r_tag[2][1]$_DFFE_PP__3188  (.L_HI(net3188));
 sg13g2_tiehi \cpu.icache.r_tag[2][2]$_DFFE_PP__3189  (.L_HI(net3189));
 sg13g2_tiehi \cpu.icache.r_tag[2][3]$_DFFE_PP__3190  (.L_HI(net3190));
 sg13g2_tiehi \cpu.icache.r_tag[2][4]$_DFFE_PP__3191  (.L_HI(net3191));
 sg13g2_tiehi \cpu.icache.r_tag[2][5]$_DFFE_PP__3192  (.L_HI(net3192));
 sg13g2_tiehi \cpu.icache.r_tag[2][6]$_DFFE_PP__3193  (.L_HI(net3193));
 sg13g2_tiehi \cpu.icache.r_tag[2][7]$_DFFE_PP__3194  (.L_HI(net3194));
 sg13g2_tiehi \cpu.icache.r_tag[2][8]$_DFFE_PP__3195  (.L_HI(net3195));
 sg13g2_tiehi \cpu.icache.r_tag[2][9]$_DFFE_PP__3196  (.L_HI(net3196));
 sg13g2_tiehi \cpu.icache.r_tag[3][0]$_DFFE_PP__3197  (.L_HI(net3197));
 sg13g2_tiehi \cpu.icache.r_tag[3][10]$_DFFE_PP__3198  (.L_HI(net3198));
 sg13g2_tiehi \cpu.icache.r_tag[3][11]$_DFFE_PP__3199  (.L_HI(net3199));
 sg13g2_tiehi \cpu.icache.r_tag[3][12]$_DFFE_PP__3200  (.L_HI(net3200));
 sg13g2_tiehi \cpu.icache.r_tag[3][13]$_DFFE_PP__3201  (.L_HI(net3201));
 sg13g2_tiehi \cpu.icache.r_tag[3][14]$_DFFE_PP__3202  (.L_HI(net3202));
 sg13g2_tiehi \cpu.icache.r_tag[3][15]$_DFFE_PP__3203  (.L_HI(net3203));
 sg13g2_tiehi \cpu.icache.r_tag[3][16]$_DFFE_PP__3204  (.L_HI(net3204));
 sg13g2_tiehi \cpu.icache.r_tag[3][17]$_DFFE_PP__3205  (.L_HI(net3205));
 sg13g2_tiehi \cpu.icache.r_tag[3][18]$_DFFE_PP__3206  (.L_HI(net3206));
 sg13g2_tiehi \cpu.icache.r_tag[3][1]$_DFFE_PP__3207  (.L_HI(net3207));
 sg13g2_tiehi \cpu.icache.r_tag[3][2]$_DFFE_PP__3208  (.L_HI(net3208));
 sg13g2_tiehi \cpu.icache.r_tag[3][3]$_DFFE_PP__3209  (.L_HI(net3209));
 sg13g2_tiehi \cpu.icache.r_tag[3][4]$_DFFE_PP__3210  (.L_HI(net3210));
 sg13g2_tiehi \cpu.icache.r_tag[3][5]$_DFFE_PP__3211  (.L_HI(net3211));
 sg13g2_tiehi \cpu.icache.r_tag[3][6]$_DFFE_PP__3212  (.L_HI(net3212));
 sg13g2_tiehi \cpu.icache.r_tag[3][7]$_DFFE_PP__3213  (.L_HI(net3213));
 sg13g2_tiehi \cpu.icache.r_tag[3][8]$_DFFE_PP__3214  (.L_HI(net3214));
 sg13g2_tiehi \cpu.icache.r_tag[3][9]$_DFFE_PP__3215  (.L_HI(net3215));
 sg13g2_tiehi \cpu.icache.r_tag[4][0]$_DFFE_PP__3216  (.L_HI(net3216));
 sg13g2_tiehi \cpu.icache.r_tag[4][10]$_DFFE_PP__3217  (.L_HI(net3217));
 sg13g2_tiehi \cpu.icache.r_tag[4][11]$_DFFE_PP__3218  (.L_HI(net3218));
 sg13g2_tiehi \cpu.icache.r_tag[4][12]$_DFFE_PP__3219  (.L_HI(net3219));
 sg13g2_tiehi \cpu.icache.r_tag[4][13]$_DFFE_PP__3220  (.L_HI(net3220));
 sg13g2_tiehi \cpu.icache.r_tag[4][14]$_DFFE_PP__3221  (.L_HI(net3221));
 sg13g2_tiehi \cpu.icache.r_tag[4][15]$_DFFE_PP__3222  (.L_HI(net3222));
 sg13g2_tiehi \cpu.icache.r_tag[4][16]$_DFFE_PP__3223  (.L_HI(net3223));
 sg13g2_tiehi \cpu.icache.r_tag[4][17]$_DFFE_PP__3224  (.L_HI(net3224));
 sg13g2_tiehi \cpu.icache.r_tag[4][18]$_DFFE_PP__3225  (.L_HI(net3225));
 sg13g2_tiehi \cpu.icache.r_tag[4][1]$_DFFE_PP__3226  (.L_HI(net3226));
 sg13g2_tiehi \cpu.icache.r_tag[4][2]$_DFFE_PP__3227  (.L_HI(net3227));
 sg13g2_tiehi \cpu.icache.r_tag[4][3]$_DFFE_PP__3228  (.L_HI(net3228));
 sg13g2_tiehi \cpu.icache.r_tag[4][4]$_DFFE_PP__3229  (.L_HI(net3229));
 sg13g2_tiehi \cpu.icache.r_tag[4][5]$_DFFE_PP__3230  (.L_HI(net3230));
 sg13g2_tiehi \cpu.icache.r_tag[4][6]$_DFFE_PP__3231  (.L_HI(net3231));
 sg13g2_tiehi \cpu.icache.r_tag[4][7]$_DFFE_PP__3232  (.L_HI(net3232));
 sg13g2_tiehi \cpu.icache.r_tag[4][8]$_DFFE_PP__3233  (.L_HI(net3233));
 sg13g2_tiehi \cpu.icache.r_tag[4][9]$_DFFE_PP__3234  (.L_HI(net3234));
 sg13g2_tiehi \cpu.icache.r_tag[5][0]$_DFFE_PP__3235  (.L_HI(net3235));
 sg13g2_tiehi \cpu.icache.r_tag[5][10]$_DFFE_PP__3236  (.L_HI(net3236));
 sg13g2_tiehi \cpu.icache.r_tag[5][11]$_DFFE_PP__3237  (.L_HI(net3237));
 sg13g2_tiehi \cpu.icache.r_tag[5][12]$_DFFE_PP__3238  (.L_HI(net3238));
 sg13g2_tiehi \cpu.icache.r_tag[5][13]$_DFFE_PP__3239  (.L_HI(net3239));
 sg13g2_tiehi \cpu.icache.r_tag[5][14]$_DFFE_PP__3240  (.L_HI(net3240));
 sg13g2_tiehi \cpu.icache.r_tag[5][15]$_DFFE_PP__3241  (.L_HI(net3241));
 sg13g2_tiehi \cpu.icache.r_tag[5][16]$_DFFE_PP__3242  (.L_HI(net3242));
 sg13g2_tiehi \cpu.icache.r_tag[5][17]$_DFFE_PP__3243  (.L_HI(net3243));
 sg13g2_tiehi \cpu.icache.r_tag[5][18]$_DFFE_PP__3244  (.L_HI(net3244));
 sg13g2_tiehi \cpu.icache.r_tag[5][1]$_DFFE_PP__3245  (.L_HI(net3245));
 sg13g2_tiehi \cpu.icache.r_tag[5][2]$_DFFE_PP__3246  (.L_HI(net3246));
 sg13g2_tiehi \cpu.icache.r_tag[5][3]$_DFFE_PP__3247  (.L_HI(net3247));
 sg13g2_tiehi \cpu.icache.r_tag[5][4]$_DFFE_PP__3248  (.L_HI(net3248));
 sg13g2_tiehi \cpu.icache.r_tag[5][5]$_DFFE_PP__3249  (.L_HI(net3249));
 sg13g2_tiehi \cpu.icache.r_tag[5][6]$_DFFE_PP__3250  (.L_HI(net3250));
 sg13g2_tiehi \cpu.icache.r_tag[5][7]$_DFFE_PP__3251  (.L_HI(net3251));
 sg13g2_tiehi \cpu.icache.r_tag[5][8]$_DFFE_PP__3252  (.L_HI(net3252));
 sg13g2_tiehi \cpu.icache.r_tag[5][9]$_DFFE_PP__3253  (.L_HI(net3253));
 sg13g2_tiehi \cpu.icache.r_tag[6][0]$_DFFE_PP__3254  (.L_HI(net3254));
 sg13g2_tiehi \cpu.icache.r_tag[6][10]$_DFFE_PP__3255  (.L_HI(net3255));
 sg13g2_tiehi \cpu.icache.r_tag[6][11]$_DFFE_PP__3256  (.L_HI(net3256));
 sg13g2_tiehi \cpu.icache.r_tag[6][12]$_DFFE_PP__3257  (.L_HI(net3257));
 sg13g2_tiehi \cpu.icache.r_tag[6][13]$_DFFE_PP__3258  (.L_HI(net3258));
 sg13g2_tiehi \cpu.icache.r_tag[6][14]$_DFFE_PP__3259  (.L_HI(net3259));
 sg13g2_tiehi \cpu.icache.r_tag[6][15]$_DFFE_PP__3260  (.L_HI(net3260));
 sg13g2_tiehi \cpu.icache.r_tag[6][16]$_DFFE_PP__3261  (.L_HI(net3261));
 sg13g2_tiehi \cpu.icache.r_tag[6][17]$_DFFE_PP__3262  (.L_HI(net3262));
 sg13g2_tiehi \cpu.icache.r_tag[6][18]$_DFFE_PP__3263  (.L_HI(net3263));
 sg13g2_tiehi \cpu.icache.r_tag[6][1]$_DFFE_PP__3264  (.L_HI(net3264));
 sg13g2_tiehi \cpu.icache.r_tag[6][2]$_DFFE_PP__3265  (.L_HI(net3265));
 sg13g2_tiehi \cpu.icache.r_tag[6][3]$_DFFE_PP__3266  (.L_HI(net3266));
 sg13g2_tiehi \cpu.icache.r_tag[6][4]$_DFFE_PP__3267  (.L_HI(net3267));
 sg13g2_tiehi \cpu.icache.r_tag[6][5]$_DFFE_PP__3268  (.L_HI(net3268));
 sg13g2_tiehi \cpu.icache.r_tag[6][6]$_DFFE_PP__3269  (.L_HI(net3269));
 sg13g2_tiehi \cpu.icache.r_tag[6][7]$_DFFE_PP__3270  (.L_HI(net3270));
 sg13g2_tiehi \cpu.icache.r_tag[6][8]$_DFFE_PP__3271  (.L_HI(net3271));
 sg13g2_tiehi \cpu.icache.r_tag[6][9]$_DFFE_PP__3272  (.L_HI(net3272));
 sg13g2_tiehi \cpu.icache.r_tag[7][0]$_DFFE_PP__3273  (.L_HI(net3273));
 sg13g2_tiehi \cpu.icache.r_tag[7][10]$_DFFE_PP__3274  (.L_HI(net3274));
 sg13g2_tiehi \cpu.icache.r_tag[7][11]$_DFFE_PP__3275  (.L_HI(net3275));
 sg13g2_tiehi \cpu.icache.r_tag[7][12]$_DFFE_PP__3276  (.L_HI(net3276));
 sg13g2_tiehi \cpu.icache.r_tag[7][13]$_DFFE_PP__3277  (.L_HI(net3277));
 sg13g2_tiehi \cpu.icache.r_tag[7][14]$_DFFE_PP__3278  (.L_HI(net3278));
 sg13g2_tiehi \cpu.icache.r_tag[7][15]$_DFFE_PP__3279  (.L_HI(net3279));
 sg13g2_tiehi \cpu.icache.r_tag[7][16]$_DFFE_PP__3280  (.L_HI(net3280));
 sg13g2_tiehi \cpu.icache.r_tag[7][17]$_DFFE_PP__3281  (.L_HI(net3281));
 sg13g2_tiehi \cpu.icache.r_tag[7][18]$_DFFE_PP__3282  (.L_HI(net3282));
 sg13g2_tiehi \cpu.icache.r_tag[7][1]$_DFFE_PP__3283  (.L_HI(net3283));
 sg13g2_tiehi \cpu.icache.r_tag[7][2]$_DFFE_PP__3284  (.L_HI(net3284));
 sg13g2_tiehi \cpu.icache.r_tag[7][3]$_DFFE_PP__3285  (.L_HI(net3285));
 sg13g2_tiehi \cpu.icache.r_tag[7][4]$_DFFE_PP__3286  (.L_HI(net3286));
 sg13g2_tiehi \cpu.icache.r_tag[7][5]$_DFFE_PP__3287  (.L_HI(net3287));
 sg13g2_tiehi \cpu.icache.r_tag[7][6]$_DFFE_PP__3288  (.L_HI(net3288));
 sg13g2_tiehi \cpu.icache.r_tag[7][7]$_DFFE_PP__3289  (.L_HI(net3289));
 sg13g2_tiehi \cpu.icache.r_tag[7][8]$_DFFE_PP__3290  (.L_HI(net3290));
 sg13g2_tiehi \cpu.icache.r_tag[7][9]$_DFFE_PP__3291  (.L_HI(net3291));
 sg13g2_tiehi \cpu.icache.r_valid[0]$_SDFFE_PP0P__3292  (.L_HI(net3292));
 sg13g2_tiehi \cpu.icache.r_valid[1]$_SDFFE_PP0P__3293  (.L_HI(net3293));
 sg13g2_tiehi \cpu.icache.r_valid[2]$_SDFFE_PP0P__3294  (.L_HI(net3294));
 sg13g2_tiehi \cpu.icache.r_valid[3]$_SDFFE_PP0P__3295  (.L_HI(net3295));
 sg13g2_tiehi \cpu.icache.r_valid[4]$_SDFFE_PP0P__3296  (.L_HI(net3296));
 sg13g2_tiehi \cpu.icache.r_valid[5]$_SDFFE_PP0P__3297  (.L_HI(net3297));
 sg13g2_tiehi \cpu.icache.r_valid[6]$_SDFFE_PP0P__3298  (.L_HI(net3298));
 sg13g2_tiehi \cpu.icache.r_valid[7]$_SDFFE_PP0P__3299  (.L_HI(net3299));
 sg13g2_tiehi \cpu.intr.r_clock$_SDFFE_PN0P__3300  (.L_HI(net3300));
 sg13g2_tiehi \cpu.intr.r_clock_cmp[0]$_DFFE_PP__3301  (.L_HI(net3301));
 sg13g2_tiehi \cpu.intr.r_clock_cmp[10]$_DFFE_PP__3302  (.L_HI(net3302));
 sg13g2_tiehi \cpu.intr.r_clock_cmp[11]$_DFFE_PP__3303  (.L_HI(net3303));
 sg13g2_tiehi \cpu.intr.r_clock_cmp[12]$_DFFE_PP__3304  (.L_HI(net3304));
 sg13g2_tiehi \cpu.intr.r_clock_cmp[13]$_DFFE_PP__3305  (.L_HI(net3305));
 sg13g2_tiehi \cpu.intr.r_clock_cmp[14]$_DFFE_PP__3306  (.L_HI(net3306));
 sg13g2_tiehi \cpu.intr.r_clock_cmp[15]$_DFFE_PP__3307  (.L_HI(net3307));
 sg13g2_tiehi \cpu.intr.r_clock_cmp[16]$_DFFE_PP__3308  (.L_HI(net3308));
 sg13g2_tiehi \cpu.intr.r_clock_cmp[17]$_DFFE_PP__3309  (.L_HI(net3309));
 sg13g2_tiehi \cpu.intr.r_clock_cmp[18]$_DFFE_PP__3310  (.L_HI(net3310));
 sg13g2_tiehi \cpu.intr.r_clock_cmp[19]$_DFFE_PP__3311  (.L_HI(net3311));
 sg13g2_tiehi \cpu.intr.r_clock_cmp[1]$_DFFE_PP__3312  (.L_HI(net3312));
 sg13g2_tiehi \cpu.intr.r_clock_cmp[20]$_DFFE_PP__3313  (.L_HI(net3313));
 sg13g2_tiehi \cpu.intr.r_clock_cmp[21]$_DFFE_PP__3314  (.L_HI(net3314));
 sg13g2_tiehi \cpu.intr.r_clock_cmp[22]$_DFFE_PP__3315  (.L_HI(net3315));
 sg13g2_tiehi \cpu.intr.r_clock_cmp[23]$_DFFE_PP__3316  (.L_HI(net3316));
 sg13g2_tiehi \cpu.intr.r_clock_cmp[24]$_DFFE_PP__3317  (.L_HI(net3317));
 sg13g2_tiehi \cpu.intr.r_clock_cmp[25]$_DFFE_PP__3318  (.L_HI(net3318));
 sg13g2_tiehi \cpu.intr.r_clock_cmp[26]$_DFFE_PP__3319  (.L_HI(net3319));
 sg13g2_tiehi \cpu.intr.r_clock_cmp[27]$_DFFE_PP__3320  (.L_HI(net3320));
 sg13g2_tiehi \cpu.intr.r_clock_cmp[28]$_DFFE_PP__3321  (.L_HI(net3321));
 sg13g2_tiehi \cpu.intr.r_clock_cmp[29]$_DFFE_PP__3322  (.L_HI(net3322));
 sg13g2_tiehi \cpu.intr.r_clock_cmp[2]$_DFFE_PP__3323  (.L_HI(net3323));
 sg13g2_tiehi \cpu.intr.r_clock_cmp[30]$_DFFE_PP__3324  (.L_HI(net3324));
 sg13g2_tiehi \cpu.intr.r_clock_cmp[31]$_DFFE_PP__3325  (.L_HI(net3325));
 sg13g2_tiehi \cpu.intr.r_clock_cmp[3]$_DFFE_PP__3326  (.L_HI(net3326));
 sg13g2_tiehi \cpu.intr.r_clock_cmp[4]$_DFFE_PP__3327  (.L_HI(net3327));
 sg13g2_tiehi \cpu.intr.r_clock_cmp[5]$_DFFE_PP__3328  (.L_HI(net3328));
 sg13g2_tiehi \cpu.intr.r_clock_cmp[6]$_DFFE_PP__3329  (.L_HI(net3329));
 sg13g2_tiehi \cpu.intr.r_clock_cmp[7]$_DFFE_PP__3330  (.L_HI(net3330));
 sg13g2_tiehi \cpu.intr.r_clock_cmp[8]$_DFFE_PP__3331  (.L_HI(net3331));
 sg13g2_tiehi \cpu.intr.r_clock_cmp[9]$_DFFE_PP__3332  (.L_HI(net3332));
 sg13g2_tiehi \cpu.intr.r_clock_count[0]$_DFF_P__3333  (.L_HI(net3333));
 sg13g2_tiehi \cpu.intr.r_clock_count[10]$_DFF_P__3334  (.L_HI(net3334));
 sg13g2_tiehi \cpu.intr.r_clock_count[11]$_DFF_P__3335  (.L_HI(net3335));
 sg13g2_tiehi \cpu.intr.r_clock_count[12]$_DFF_P__3336  (.L_HI(net3336));
 sg13g2_tiehi \cpu.intr.r_clock_count[13]$_DFF_P__3337  (.L_HI(net3337));
 sg13g2_tiehi \cpu.intr.r_clock_count[14]$_DFF_P__3338  (.L_HI(net3338));
 sg13g2_tiehi \cpu.intr.r_clock_count[15]$_DFF_P__3339  (.L_HI(net3339));
 sg13g2_tiehi \cpu.intr.r_clock_count[16]$_DFFE_PN__3340  (.L_HI(net3340));
 sg13g2_tiehi \cpu.intr.r_clock_count[17]$_DFFE_PN__3341  (.L_HI(net3341));
 sg13g2_tiehi \cpu.intr.r_clock_count[18]$_DFFE_PN__3342  (.L_HI(net3342));
 sg13g2_tiehi \cpu.intr.r_clock_count[19]$_DFFE_PN__3343  (.L_HI(net3343));
 sg13g2_tiehi \cpu.intr.r_clock_count[1]$_DFF_P__3344  (.L_HI(net3344));
 sg13g2_tiehi \cpu.intr.r_clock_count[20]$_DFFE_PN__3345  (.L_HI(net3345));
 sg13g2_tiehi \cpu.intr.r_clock_count[21]$_DFFE_PN__3346  (.L_HI(net3346));
 sg13g2_tiehi \cpu.intr.r_clock_count[22]$_DFFE_PN__3347  (.L_HI(net3347));
 sg13g2_tiehi \cpu.intr.r_clock_count[23]$_DFFE_PN__3348  (.L_HI(net3348));
 sg13g2_tiehi \cpu.intr.r_clock_count[24]$_DFFE_PN__3349  (.L_HI(net3349));
 sg13g2_tiehi \cpu.intr.r_clock_count[25]$_DFFE_PN__3350  (.L_HI(net3350));
 sg13g2_tiehi \cpu.intr.r_clock_count[26]$_DFFE_PN__3351  (.L_HI(net3351));
 sg13g2_tiehi \cpu.intr.r_clock_count[27]$_DFFE_PN__3352  (.L_HI(net3352));
 sg13g2_tiehi \cpu.intr.r_clock_count[28]$_DFFE_PN__3353  (.L_HI(net3353));
 sg13g2_tiehi \cpu.intr.r_clock_count[29]$_DFFE_PN__3354  (.L_HI(net3354));
 sg13g2_tiehi \cpu.intr.r_clock_count[2]$_DFF_P__3355  (.L_HI(net3355));
 sg13g2_tiehi \cpu.intr.r_clock_count[30]$_DFFE_PN__3356  (.L_HI(net3356));
 sg13g2_tiehi \cpu.intr.r_clock_count[31]$_DFFE_PN__3357  (.L_HI(net3357));
 sg13g2_tiehi \cpu.intr.r_clock_count[3]$_DFF_P__3358  (.L_HI(net3358));
 sg13g2_tiehi \cpu.intr.r_clock_count[4]$_DFF_P__3359  (.L_HI(net3359));
 sg13g2_tiehi \cpu.intr.r_clock_count[5]$_DFF_P__3360  (.L_HI(net3360));
 sg13g2_tiehi \cpu.intr.r_clock_count[6]$_DFF_P__3361  (.L_HI(net3361));
 sg13g2_tiehi \cpu.intr.r_clock_count[7]$_DFF_P__3362  (.L_HI(net3362));
 sg13g2_tiehi \cpu.intr.r_clock_count[8]$_DFF_P__3363  (.L_HI(net3363));
 sg13g2_tiehi \cpu.intr.r_clock_count[9]$_DFF_P__3364  (.L_HI(net3364));
 sg13g2_tiehi \cpu.intr.r_enable[0]$_SDFFE_PN0P__3365  (.L_HI(net3365));
 sg13g2_tiehi \cpu.intr.r_enable[1]$_SDFFE_PN0P__3366  (.L_HI(net3366));
 sg13g2_tiehi \cpu.intr.r_enable[2]$_SDFFE_PN0P__3367  (.L_HI(net3367));
 sg13g2_tiehi \cpu.intr.r_enable[3]$_SDFFE_PN0P__3368  (.L_HI(net3368));
 sg13g2_tiehi \cpu.intr.r_enable[4]$_SDFFE_PN0P__3369  (.L_HI(net3369));
 sg13g2_tiehi \cpu.intr.r_enable[5]$_SDFFE_PN0P__3370  (.L_HI(net3370));
 sg13g2_tiehi \cpu.intr.r_timer$_SDFFE_PN0P__3371  (.L_HI(net3371));
 sg13g2_tiehi \cpu.intr.r_timer_count[0]$_DFF_P__3372  (.L_HI(net3372));
 sg13g2_tiehi \cpu.intr.r_timer_count[10]$_DFF_P__3373  (.L_HI(net3373));
 sg13g2_tiehi \cpu.intr.r_timer_count[11]$_DFF_P__3374  (.L_HI(net3374));
 sg13g2_tiehi \cpu.intr.r_timer_count[12]$_DFF_P__3375  (.L_HI(net3375));
 sg13g2_tiehi \cpu.intr.r_timer_count[13]$_DFF_P__3376  (.L_HI(net3376));
 sg13g2_tiehi \cpu.intr.r_timer_count[14]$_DFF_P__3377  (.L_HI(net3377));
 sg13g2_tiehi \cpu.intr.r_timer_count[15]$_DFF_P__3378  (.L_HI(net3378));
 sg13g2_tiehi \cpu.intr.r_timer_count[16]$_DFF_P__3379  (.L_HI(net3379));
 sg13g2_tiehi \cpu.intr.r_timer_count[17]$_DFF_P__3380  (.L_HI(net3380));
 sg13g2_tiehi \cpu.intr.r_timer_count[18]$_DFF_P__3381  (.L_HI(net3381));
 sg13g2_tiehi \cpu.intr.r_timer_count[19]$_DFF_P__3382  (.L_HI(net3382));
 sg13g2_tiehi \cpu.intr.r_timer_count[1]$_DFF_P__3383  (.L_HI(net3383));
 sg13g2_tiehi \cpu.intr.r_timer_count[20]$_DFF_P__3384  (.L_HI(net3384));
 sg13g2_tiehi \cpu.intr.r_timer_count[21]$_DFF_P__3385  (.L_HI(net3385));
 sg13g2_tiehi \cpu.intr.r_timer_count[22]$_DFF_P__3386  (.L_HI(net3386));
 sg13g2_tiehi \cpu.intr.r_timer_count[23]$_DFF_P__3387  (.L_HI(net3387));
 sg13g2_tiehi \cpu.intr.r_timer_count[2]$_DFF_P__3388  (.L_HI(net3388));
 sg13g2_tiehi \cpu.intr.r_timer_count[3]$_DFF_P__3389  (.L_HI(net3389));
 sg13g2_tiehi \cpu.intr.r_timer_count[4]$_DFF_P__3390  (.L_HI(net3390));
 sg13g2_tiehi \cpu.intr.r_timer_count[5]$_DFF_P__3391  (.L_HI(net3391));
 sg13g2_tiehi \cpu.intr.r_timer_count[6]$_DFF_P__3392  (.L_HI(net3392));
 sg13g2_tiehi \cpu.intr.r_timer_count[7]$_DFF_P__3393  (.L_HI(net3393));
 sg13g2_tiehi \cpu.intr.r_timer_count[8]$_DFF_P__3394  (.L_HI(net3394));
 sg13g2_tiehi \cpu.intr.r_timer_count[9]$_DFF_P__3395  (.L_HI(net3395));
 sg13g2_tiehi \cpu.intr.r_timer_reload[0]$_DFFE_PP__3396  (.L_HI(net3396));
 sg13g2_tiehi \cpu.intr.r_timer_reload[10]$_DFFE_PP__3397  (.L_HI(net3397));
 sg13g2_tiehi \cpu.intr.r_timer_reload[11]$_DFFE_PP__3398  (.L_HI(net3398));
 sg13g2_tiehi \cpu.intr.r_timer_reload[12]$_DFFE_PP__3399  (.L_HI(net3399));
 sg13g2_tiehi \cpu.intr.r_timer_reload[13]$_DFFE_PP__3400  (.L_HI(net3400));
 sg13g2_tiehi \cpu.intr.r_timer_reload[14]$_DFFE_PP__3401  (.L_HI(net3401));
 sg13g2_tiehi \cpu.intr.r_timer_reload[15]$_DFFE_PP__3402  (.L_HI(net3402));
 sg13g2_tiehi \cpu.intr.r_timer_reload[16]$_DFFE_PP__3403  (.L_HI(net3403));
 sg13g2_tiehi \cpu.intr.r_timer_reload[17]$_DFFE_PP__3404  (.L_HI(net3404));
 sg13g2_tiehi \cpu.intr.r_timer_reload[18]$_DFFE_PP__3405  (.L_HI(net3405));
 sg13g2_tiehi \cpu.intr.r_timer_reload[19]$_DFFE_PP__3406  (.L_HI(net3406));
 sg13g2_tiehi \cpu.intr.r_timer_reload[1]$_DFFE_PP__3407  (.L_HI(net3407));
 sg13g2_tiehi \cpu.intr.r_timer_reload[20]$_DFFE_PP__3408  (.L_HI(net3408));
 sg13g2_tiehi \cpu.intr.r_timer_reload[21]$_DFFE_PP__3409  (.L_HI(net3409));
 sg13g2_tiehi \cpu.intr.r_timer_reload[22]$_DFFE_PP__3410  (.L_HI(net3410));
 sg13g2_tiehi \cpu.intr.r_timer_reload[23]$_DFFE_PP__3411  (.L_HI(net3411));
 sg13g2_tiehi \cpu.intr.r_timer_reload[2]$_DFFE_PP__3412  (.L_HI(net3412));
 sg13g2_tiehi \cpu.intr.r_timer_reload[3]$_DFFE_PP__3413  (.L_HI(net3413));
 sg13g2_tiehi \cpu.intr.r_timer_reload[4]$_DFFE_PP__3414  (.L_HI(net3414));
 sg13g2_tiehi \cpu.intr.r_timer_reload[5]$_DFFE_PP__3415  (.L_HI(net3415));
 sg13g2_tiehi \cpu.intr.r_timer_reload[6]$_DFFE_PP__3416  (.L_HI(net3416));
 sg13g2_tiehi \cpu.intr.r_timer_reload[7]$_DFFE_PP__3417  (.L_HI(net3417));
 sg13g2_tiehi \cpu.intr.r_timer_reload[8]$_DFFE_PP__3418  (.L_HI(net3418));
 sg13g2_tiehi \cpu.intr.r_timer_reload[9]$_DFFE_PP__3419  (.L_HI(net3419));
 sg13g2_tiehi \cpu.qspi.r_count[0]$_DFFE_PP__3420  (.L_HI(net3420));
 sg13g2_tiehi \cpu.qspi.r_count[1]$_DFFE_PP__3421  (.L_HI(net3421));
 sg13g2_tiehi \cpu.qspi.r_count[2]$_DFFE_PP__3422  (.L_HI(net3422));
 sg13g2_tiehi \cpu.qspi.r_count[3]$_DFFE_PP__3423  (.L_HI(net3423));
 sg13g2_tiehi \cpu.qspi.r_count[4]$_DFFE_PP__3424  (.L_HI(net3424));
 sg13g2_tiehi \cpu.qspi.r_cs[0]$_SDFFE_PN1P__3425  (.L_HI(net3425));
 sg13g2_tiehi \cpu.qspi.r_cs[1]$_SDFFE_PN1P__3426  (.L_HI(net3426));
 sg13g2_tiehi \cpu.qspi.r_cs[2]$_SDFFE_PN1P__3427  (.L_HI(net3427));
 sg13g2_tiehi \cpu.qspi.r_ind$_SDFFE_PN0N__3428  (.L_HI(net3428));
 sg13g2_tiehi \cpu.qspi.r_mask[0]$_SDFFE_PN0P__3429  (.L_HI(net3429));
 sg13g2_tiehi \cpu.qspi.r_mask[1]$_SDFFE_PN1P__3430  (.L_HI(net3430));
 sg13g2_tiehi \cpu.qspi.r_mask[2]$_SDFFE_PN0P__3431  (.L_HI(net3431));
 sg13g2_tiehi \cpu.qspi.r_quad[0]$_SDFFE_PN1P__3432  (.L_HI(net3432));
 sg13g2_tiehi \cpu.qspi.r_quad[1]$_SDFFE_PN0P__3433  (.L_HI(net3433));
 sg13g2_tiehi \cpu.qspi.r_quad[2]$_SDFFE_PN1P__3434  (.L_HI(net3434));
 sg13g2_tiehi \cpu.qspi.r_read_delay[0][0]$_SDFFCE_PN0P__3435  (.L_HI(net3435));
 sg13g2_tiehi \cpu.qspi.r_read_delay[0][1]$_SDFFCE_PN0P__3436  (.L_HI(net3436));
 sg13g2_tiehi \cpu.qspi.r_read_delay[0][2]$_SDFFCE_PN1P__3437  (.L_HI(net3437));
 sg13g2_tiehi \cpu.qspi.r_read_delay[0][3]$_SDFFCE_PN0P__3438  (.L_HI(net3438));
 sg13g2_tiehi \cpu.qspi.r_read_delay[1][0]$_SDFFCE_PN0P__3439  (.L_HI(net3439));
 sg13g2_tiehi \cpu.qspi.r_read_delay[1][1]$_SDFFCE_PN0P__3440  (.L_HI(net3440));
 sg13g2_tiehi \cpu.qspi.r_read_delay[1][2]$_SDFFCE_PN1P__3441  (.L_HI(net3441));
 sg13g2_tiehi \cpu.qspi.r_read_delay[1][3]$_SDFFCE_PN0P__3442  (.L_HI(net3442));
 sg13g2_tiehi \cpu.qspi.r_read_delay[2][0]$_SDFFCE_PN0P__3443  (.L_HI(net3443));
 sg13g2_tiehi \cpu.qspi.r_read_delay[2][1]$_SDFFCE_PN0P__3444  (.L_HI(net3444));
 sg13g2_tiehi \cpu.qspi.r_read_delay[2][2]$_SDFFCE_PN1P__3445  (.L_HI(net3445));
 sg13g2_tiehi \cpu.qspi.r_read_delay[2][3]$_SDFFCE_PN0P__3446  (.L_HI(net3446));
 sg13g2_tiehi \cpu.qspi.r_rom_mode[0]$_SDFFE_PN1P__3447  (.L_HI(net3447));
 sg13g2_tiehi \cpu.qspi.r_rom_mode[1]$_SDFFE_PN1P__3448  (.L_HI(net3448));
 sg13g2_tiehi \cpu.qspi.r_rstrobe_d$_DFF_P__3449  (.L_HI(net3449));
 sg13g2_tiehi \cpu.qspi.r_state[0]$_DFF_P__3450  (.L_HI(net3450));
 sg13g2_tiehi \cpu.qspi.r_state[10]$_DFF_P__3451  (.L_HI(net3451));
 sg13g2_tiehi \cpu.qspi.r_state[11]$_DFF_P__3452  (.L_HI(net3452));
 sg13g2_tiehi \cpu.qspi.r_state[12]$_DFF_P__3453  (.L_HI(net3453));
 sg13g2_tiehi \cpu.qspi.r_state[13]$_DFF_P__3454  (.L_HI(net3454));
 sg13g2_tiehi \cpu.qspi.r_state[14]$_DFF_P__3455  (.L_HI(net3455));
 sg13g2_tiehi \cpu.qspi.r_state[15]$_DFF_P__3456  (.L_HI(net3456));
 sg13g2_tiehi \cpu.qspi.r_state[16]$_DFF_P__3457  (.L_HI(net3457));
 sg13g2_tiehi \cpu.qspi.r_state[17]$_DFF_P__3458  (.L_HI(net3458));
 sg13g2_tiehi \cpu.qspi.r_state[1]$_DFF_P__3459  (.L_HI(net3459));
 sg13g2_tiehi \cpu.qspi.r_state[2]$_DFF_P__3460  (.L_HI(net3460));
 sg13g2_tiehi \cpu.qspi.r_state[3]$_DFF_P__3461  (.L_HI(net3461));
 sg13g2_tiehi \cpu.qspi.r_state[4]$_DFF_P__3462  (.L_HI(net3462));
 sg13g2_tiehi \cpu.qspi.r_state[5]$_DFF_P__3463  (.L_HI(net3463));
 sg13g2_tiehi \cpu.qspi.r_state[6]$_DFF_P__3464  (.L_HI(net3464));
 sg13g2_tiehi \cpu.qspi.r_state[7]$_DFF_P__3465  (.L_HI(net3465));
 sg13g2_tiehi \cpu.qspi.r_state[8]$_DFF_P__3466  (.L_HI(net3466));
 sg13g2_tiehi \cpu.qspi.r_state[9]$_DFF_P__3467  (.L_HI(net3467));
 sg13g2_tiehi \cpu.qspi.r_uio_oe[0]$_SDFFE_PN0P__3468  (.L_HI(net3468));
 sg13g2_tiehi \cpu.qspi.r_uio_oe[1]$_SDFFE_PN0P__3469  (.L_HI(net3469));
 sg13g2_tiehi \cpu.qspi.r_uio_out[0]$_DFFE_PP__3470  (.L_HI(net3470));
 sg13g2_tiehi \cpu.qspi.r_uio_out[1]$_DFFE_PP__3471  (.L_HI(net3471));
 sg13g2_tiehi \cpu.qspi.r_uio_out[2]$_DFFE_PP__3472  (.L_HI(net3472));
 sg13g2_tiehi \cpu.qspi.r_uio_out[3]$_DFFE_PP__3473  (.L_HI(net3473));
 sg13g2_tiehi \cpu.qspi.r_wstrobe_d$_DFF_P__3474  (.L_HI(net3474));
 sg13g2_tiehi \cpu.qspi.r_wstrobe_i$_DFF_P__3475  (.L_HI(net3475));
 sg13g2_tiehi \cpu.r_clk_invert$_DFFE_PN__3476  (.L_HI(net3476));
 sg13g2_tiehi \cpu.spi.r_bits[0]$_SDFFE_PN1P__3477  (.L_HI(net3477));
 sg13g2_tiehi \cpu.spi.r_bits[1]$_SDFFE_PN1P__3478  (.L_HI(net3478));
 sg13g2_tiehi \cpu.spi.r_bits[2]$_SDFFE_PN1P__3479  (.L_HI(net3479));
 sg13g2_tiehi \cpu.spi.r_clk_count[0][0]$_DFFE_PP__3480  (.L_HI(net3480));
 sg13g2_tiehi \cpu.spi.r_clk_count[0][1]$_DFFE_PP__3481  (.L_HI(net3481));
 sg13g2_tiehi \cpu.spi.r_clk_count[0][2]$_DFFE_PP__3482  (.L_HI(net3482));
 sg13g2_tiehi \cpu.spi.r_clk_count[0][3]$_DFFE_PP__3483  (.L_HI(net3483));
 sg13g2_tiehi \cpu.spi.r_clk_count[0][4]$_DFFE_PP__3484  (.L_HI(net3484));
 sg13g2_tiehi \cpu.spi.r_clk_count[0][5]$_DFFE_PP__3485  (.L_HI(net3485));
 sg13g2_tiehi \cpu.spi.r_clk_count[0][6]$_DFFE_PP__3486  (.L_HI(net3486));
 sg13g2_tiehi \cpu.spi.r_clk_count[0][7]$_DFFE_PP__3487  (.L_HI(net3487));
 sg13g2_tiehi \cpu.spi.r_clk_count[1][0]$_DFFE_PP__3488  (.L_HI(net3488));
 sg13g2_tiehi \cpu.spi.r_clk_count[1][1]$_DFFE_PP__3489  (.L_HI(net3489));
 sg13g2_tiehi \cpu.spi.r_clk_count[1][2]$_DFFE_PP__3490  (.L_HI(net3490));
 sg13g2_tiehi \cpu.spi.r_clk_count[1][3]$_DFFE_PP__3491  (.L_HI(net3491));
 sg13g2_tiehi \cpu.spi.r_clk_count[1][4]$_DFFE_PP__3492  (.L_HI(net3492));
 sg13g2_tiehi \cpu.spi.r_clk_count[1][5]$_DFFE_PP__3493  (.L_HI(net3493));
 sg13g2_tiehi \cpu.spi.r_clk_count[1][6]$_DFFE_PP__3494  (.L_HI(net3494));
 sg13g2_tiehi \cpu.spi.r_clk_count[1][7]$_DFFE_PP__3495  (.L_HI(net3495));
 sg13g2_tiehi \cpu.spi.r_clk_count[2][0]$_DFFE_PP__3496  (.L_HI(net3496));
 sg13g2_tiehi \cpu.spi.r_clk_count[2][1]$_DFFE_PP__3497  (.L_HI(net3497));
 sg13g2_tiehi \cpu.spi.r_clk_count[2][2]$_DFFE_PP__3498  (.L_HI(net3498));
 sg13g2_tiehi \cpu.spi.r_clk_count[2][3]$_DFFE_PP__3499  (.L_HI(net3499));
 sg13g2_tiehi \cpu.spi.r_clk_count[2][4]$_DFFE_PP__3500  (.L_HI(net3500));
 sg13g2_tiehi \cpu.spi.r_clk_count[2][5]$_DFFE_PP__3501  (.L_HI(net3501));
 sg13g2_tiehi \cpu.spi.r_clk_count[2][6]$_DFFE_PP__3502  (.L_HI(net3502));
 sg13g2_tiehi \cpu.spi.r_clk_count[2][7]$_DFFE_PP__3503  (.L_HI(net3503));
 sg13g2_tiehi \cpu.spi.r_count[0]$_DFFE_PP__3504  (.L_HI(net3504));
 sg13g2_tiehi \cpu.spi.r_count[1]$_DFFE_PP__3505  (.L_HI(net3505));
 sg13g2_tiehi \cpu.spi.r_count[2]$_DFFE_PP__3506  (.L_HI(net3506));
 sg13g2_tiehi \cpu.spi.r_count[3]$_DFFE_PP__3507  (.L_HI(net3507));
 sg13g2_tiehi \cpu.spi.r_count[4]$_DFFE_PP__3508  (.L_HI(net3508));
 sg13g2_tiehi \cpu.spi.r_count[5]$_DFFE_PP__3509  (.L_HI(net3509));
 sg13g2_tiehi \cpu.spi.r_count[6]$_DFFE_PP__3510  (.L_HI(net3510));
 sg13g2_tiehi \cpu.spi.r_count[7]$_DFFE_PP__3511  (.L_HI(net3511));
 sg13g2_tiehi \cpu.spi.r_cs[0]$_SDFFE_PN1P__3512  (.L_HI(net3512));
 sg13g2_tiehi \cpu.spi.r_cs[1]$_SDFFE_PN1P__3513  (.L_HI(net3513));
 sg13g2_tiehi \cpu.spi.r_cs[2]$_SDFFE_PN1P__3514  (.L_HI(net3514));
 sg13g2_tiehi \cpu.spi.r_in[0]$_DFFE_PP__3515  (.L_HI(net3515));
 sg13g2_tiehi \cpu.spi.r_in[1]$_DFFE_PP__3516  (.L_HI(net3516));
 sg13g2_tiehi \cpu.spi.r_in[2]$_DFFE_PP__3517  (.L_HI(net3517));
 sg13g2_tiehi \cpu.spi.r_in[3]$_DFFE_PP__3518  (.L_HI(net3518));
 sg13g2_tiehi \cpu.spi.r_in[4]$_DFFE_PP__3519  (.L_HI(net3519));
 sg13g2_tiehi \cpu.spi.r_in[5]$_DFFE_PP__3520  (.L_HI(net3520));
 sg13g2_tiehi \cpu.spi.r_in[6]$_DFFE_PP__3521  (.L_HI(net3521));
 sg13g2_tiehi \cpu.spi.r_in[7]$_DFFE_PP__3522  (.L_HI(net3522));
 sg13g2_tiehi \cpu.spi.r_interrupt$_SDFFE_PN0P__3523  (.L_HI(net3523));
 sg13g2_tiehi \cpu.spi.r_mode[0][0]$_DFFE_PP__3524  (.L_HI(net3524));
 sg13g2_tiehi \cpu.spi.r_mode[0][1]$_DFFE_PP__3525  (.L_HI(net3525));
 sg13g2_tiehi \cpu.spi.r_mode[1][0]$_DFFE_PP__3526  (.L_HI(net3526));
 sg13g2_tiehi \cpu.spi.r_mode[1][1]$_DFFE_PP__3527  (.L_HI(net3527));
 sg13g2_tiehi \cpu.spi.r_mode[2][0]$_DFFE_PP__3528  (.L_HI(net3528));
 sg13g2_tiehi \cpu.spi.r_mode[2][1]$_DFFE_PP__3529  (.L_HI(net3529));
 sg13g2_tiehi \cpu.spi.r_out[0]$_DFFE_PP__3530  (.L_HI(net3530));
 sg13g2_tiehi \cpu.spi.r_out[1]$_DFFE_PP__3531  (.L_HI(net3531));
 sg13g2_tiehi \cpu.spi.r_out[2]$_DFFE_PP__3532  (.L_HI(net3532));
 sg13g2_tiehi \cpu.spi.r_out[3]$_DFFE_PP__3533  (.L_HI(net3533));
 sg13g2_tiehi \cpu.spi.r_out[4]$_DFFE_PP__3534  (.L_HI(net3534));
 sg13g2_tiehi \cpu.spi.r_out[5]$_DFFE_PP__3535  (.L_HI(net3535));
 sg13g2_tiehi \cpu.spi.r_out[6]$_DFFE_PP__3536  (.L_HI(net3536));
 sg13g2_tiehi \cpu.spi.r_out[7]$_DFFE_PP__3537  (.L_HI(net3537));
 sg13g2_tiehi \cpu.spi.r_ready$_SDFFE_PN1P__3538  (.L_HI(net3538));
 sg13g2_tiehi \cpu.spi.r_searching$_SDFFE_PN0P__3539  (.L_HI(net3539));
 sg13g2_tiehi \cpu.spi.r_sel[0]$_DFFE_PP__3540  (.L_HI(net3540));
 sg13g2_tiehi \cpu.spi.r_sel[1]$_DFFE_PP__3541  (.L_HI(net3541));
 sg13g2_tiehi \cpu.spi.r_src[0]$_DFFE_PP__3542  (.L_HI(net3542));
 sg13g2_tiehi \cpu.spi.r_src[1]$_DFFE_PP__3543  (.L_HI(net3543));
 sg13g2_tiehi \cpu.spi.r_src[2]$_DFFE_PP__3544  (.L_HI(net3544));
 sg13g2_tiehi \cpu.spi.r_state[0]$_DFF_P__3545  (.L_HI(net3545));
 sg13g2_tiehi \cpu.spi.r_state[1]$_DFF_P__3546  (.L_HI(net3546));
 sg13g2_tiehi \cpu.spi.r_state[2]$_DFF_P__3547  (.L_HI(net3547));
 sg13g2_tiehi \cpu.spi.r_state[3]$_DFF_P__3548  (.L_HI(net3548));
 sg13g2_tiehi \cpu.spi.r_state[4]$_DFF_P__3549  (.L_HI(net3549));
 sg13g2_tiehi \cpu.spi.r_state[5]$_DFF_P__3550  (.L_HI(net3550));
 sg13g2_tiehi \cpu.spi.r_state[6]$_DFF_P__3551  (.L_HI(net3551));
 sg13g2_tiehi \cpu.spi.r_timeout[0]$_DFFE_PP__3552  (.L_HI(net3552));
 sg13g2_tiehi \cpu.spi.r_timeout[1]$_DFFE_PP__3553  (.L_HI(net3553));
 sg13g2_tiehi \cpu.spi.r_timeout[2]$_DFFE_PP__3554  (.L_HI(net3554));
 sg13g2_tiehi \cpu.spi.r_timeout[3]$_DFFE_PP__3555  (.L_HI(net3555));
 sg13g2_tiehi \cpu.spi.r_timeout[4]$_DFFE_PP__3556  (.L_HI(net3556));
 sg13g2_tiehi \cpu.spi.r_timeout[5]$_DFFE_PP__3557  (.L_HI(net3557));
 sg13g2_tiehi \cpu.spi.r_timeout[6]$_DFFE_PP__3558  (.L_HI(net3558));
 sg13g2_tiehi \cpu.spi.r_timeout[7]$_DFFE_PP__3559  (.L_HI(net3559));
 sg13g2_tiehi \cpu.spi.r_timeout_count[0]$_DFFE_PP__3560  (.L_HI(net3560));
 sg13g2_tiehi \cpu.spi.r_timeout_count[1]$_DFFE_PP__3561  (.L_HI(net3561));
 sg13g2_tiehi \cpu.spi.r_timeout_count[2]$_DFFE_PP__3562  (.L_HI(net3562));
 sg13g2_tiehi \cpu.spi.r_timeout_count[3]$_DFFE_PP__3563  (.L_HI(net3563));
 sg13g2_tiehi \cpu.spi.r_timeout_count[4]$_DFFE_PP__3564  (.L_HI(net3564));
 sg13g2_tiehi \cpu.spi.r_timeout_count[5]$_DFFE_PP__3565  (.L_HI(net3565));
 sg13g2_tiehi \cpu.spi.r_timeout_count[6]$_DFFE_PP__3566  (.L_HI(net3566));
 sg13g2_tiehi \cpu.spi.r_timeout_count[7]$_DFFE_PP__3567  (.L_HI(net3567));
 sg13g2_tiehi \cpu.uart.r_div[0]$_DFF_P__3568  (.L_HI(net3568));
 sg13g2_tiehi \cpu.uart.r_div[10]$_DFF_P__3569  (.L_HI(net3569));
 sg13g2_tiehi \cpu.uart.r_div[11]$_DFF_P__3570  (.L_HI(net3570));
 sg13g2_tiehi \cpu.uart.r_div[1]$_DFF_P__3571  (.L_HI(net3571));
 sg13g2_tiehi \cpu.uart.r_div[2]$_DFF_P__3572  (.L_HI(net3572));
 sg13g2_tiehi \cpu.uart.r_div[3]$_DFF_P__3573  (.L_HI(net3573));
 sg13g2_tiehi \cpu.uart.r_div[4]$_DFF_P__3574  (.L_HI(net3574));
 sg13g2_tiehi \cpu.uart.r_div[5]$_DFF_P__3575  (.L_HI(net3575));
 sg13g2_tiehi \cpu.uart.r_div[6]$_DFF_P__3576  (.L_HI(net3576));
 sg13g2_tiehi \cpu.uart.r_div[7]$_DFF_P__3577  (.L_HI(net3577));
 sg13g2_tiehi \cpu.uart.r_div[8]$_DFF_P__3578  (.L_HI(net3578));
 sg13g2_tiehi \cpu.uart.r_div[9]$_DFF_P__3579  (.L_HI(net3579));
 sg13g2_tiehi \cpu.uart.r_div_value[0]$_SDFFE_PN1P__3580  (.L_HI(net3580));
 sg13g2_tiehi \cpu.uart.r_div_value[10]$_SDFFE_PN0P__3581  (.L_HI(net3581));
 sg13g2_tiehi \cpu.uart.r_div_value[11]$_SDFFE_PN0P__3582  (.L_HI(net3582));
 sg13g2_tiehi \cpu.uart.r_div_value[1]$_SDFFE_PN0P__3583  (.L_HI(net3583));
 sg13g2_tiehi \cpu.uart.r_div_value[2]$_SDFFE_PN0P__3584  (.L_HI(net3584));
 sg13g2_tiehi \cpu.uart.r_div_value[3]$_SDFFE_PN0P__3585  (.L_HI(net3585));
 sg13g2_tiehi \cpu.uart.r_div_value[4]$_SDFFE_PN0P__3586  (.L_HI(net3586));
 sg13g2_tiehi \cpu.uart.r_div_value[5]$_SDFFE_PN0P__3587  (.L_HI(net3587));
 sg13g2_tiehi \cpu.uart.r_div_value[6]$_SDFFE_PN0P__3588  (.L_HI(net3588));
 sg13g2_tiehi \cpu.uart.r_div_value[7]$_SDFFE_PN0P__3589  (.L_HI(net3589));
 sg13g2_tiehi \cpu.uart.r_div_value[8]$_SDFFE_PN0P__3590  (.L_HI(net3590));
 sg13g2_tiehi \cpu.uart.r_div_value[9]$_SDFFE_PN0P__3591  (.L_HI(net3591));
 sg13g2_tiehi \cpu.uart.r_ib[0]$_DFFE_PP__3592  (.L_HI(net3592));
 sg13g2_tiehi \cpu.uart.r_ib[1]$_DFFE_PP__3593  (.L_HI(net3593));
 sg13g2_tiehi \cpu.uart.r_ib[2]$_DFFE_PP__3594  (.L_HI(net3594));
 sg13g2_tiehi \cpu.uart.r_ib[3]$_DFFE_PP__3595  (.L_HI(net3595));
 sg13g2_tiehi \cpu.uart.r_ib[4]$_DFFE_PP__3596  (.L_HI(net3596));
 sg13g2_tiehi \cpu.uart.r_ib[5]$_DFFE_PP__3597  (.L_HI(net3597));
 sg13g2_tiehi \cpu.uart.r_ib[6]$_DFFE_PP__3598  (.L_HI(net3598));
 sg13g2_tiehi \cpu.uart.r_in[0]$_DFFE_PP__3599  (.L_HI(net3599));
 sg13g2_tiehi \cpu.uart.r_in[1]$_DFFE_PP__3600  (.L_HI(net3600));
 sg13g2_tiehi \cpu.uart.r_in[2]$_DFFE_PP__3601  (.L_HI(net3601));
 sg13g2_tiehi \cpu.uart.r_in[3]$_DFFE_PP__3602  (.L_HI(net3602));
 sg13g2_tiehi \cpu.uart.r_in[4]$_DFFE_PP__3603  (.L_HI(net3603));
 sg13g2_tiehi \cpu.uart.r_in[5]$_DFFE_PP__3604  (.L_HI(net3604));
 sg13g2_tiehi \cpu.uart.r_in[6]$_DFFE_PP__3605  (.L_HI(net3605));
 sg13g2_tiehi \cpu.uart.r_in[7]$_DFFE_PP__3606  (.L_HI(net3606));
 sg13g2_tiehi \cpu.uart.r_out[0]$_DFFE_PP__3607  (.L_HI(net3607));
 sg13g2_tiehi \cpu.uart.r_out[1]$_DFFE_PP__3608  (.L_HI(net3608));
 sg13g2_tiehi \cpu.uart.r_out[2]$_DFFE_PP__3609  (.L_HI(net3609));
 sg13g2_tiehi \cpu.uart.r_out[3]$_DFFE_PP__3610  (.L_HI(net3610));
 sg13g2_tiehi \cpu.uart.r_out[4]$_DFFE_PP__3611  (.L_HI(net3611));
 sg13g2_tiehi \cpu.uart.r_out[5]$_DFFE_PP__3612  (.L_HI(net3612));
 sg13g2_tiehi \cpu.uart.r_out[6]$_DFFE_PP__3613  (.L_HI(net3613));
 sg13g2_tiehi \cpu.uart.r_out[7]$_DFFE_PP__3614  (.L_HI(net3614));
 sg13g2_tiehi \cpu.uart.r_r$_DFF_P__3615  (.L_HI(net3615));
 sg13g2_tiehi \cpu.uart.r_r_int$_SDFFE_PN0P__3616  (.L_HI(net3616));
 sg13g2_tiehi \cpu.uart.r_r_invert$_SDFFE_PN0P__3617  (.L_HI(net3617));
 sg13g2_tiehi \cpu.uart.r_rcnt[0]$_DFFE_PP__3618  (.L_HI(net3618));
 sg13g2_tiehi \cpu.uart.r_rcnt[1]$_DFFE_PP__3619  (.L_HI(net3619));
 sg13g2_tiehi \cpu.uart.r_rstate[0]$_SDFFE_PN0P__3620  (.L_HI(net3620));
 sg13g2_tiehi \cpu.uart.r_rstate[1]$_SDFFE_PN0P__3621  (.L_HI(net3621));
 sg13g2_tiehi \cpu.uart.r_rstate[2]$_SDFFE_PN0P__3622  (.L_HI(net3622));
 sg13g2_tiehi \cpu.uart.r_rstate[3]$_SDFFE_PN0P__3623  (.L_HI(net3623));
 sg13g2_tiehi \cpu.uart.r_x$_DFFE_PP__3624  (.L_HI(net3624));
 sg13g2_tiehi \cpu.uart.r_x_int$_SDFFE_PN0P__3625  (.L_HI(net3625));
 sg13g2_tiehi \cpu.uart.r_x_invert$_SDFFE_PN0P__3626  (.L_HI(net3626));
 sg13g2_tiehi \cpu.uart.r_xcnt[0]$_DFFE_PP__3627  (.L_HI(net3627));
 sg13g2_tiehi \cpu.uart.r_xcnt[1]$_DFFE_PP__3628  (.L_HI(net3628));
 sg13g2_tiehi \cpu.uart.r_xstate[0]$_SDFFE_PN0P__3629  (.L_HI(net3629));
 sg13g2_tiehi \cpu.uart.r_xstate[1]$_SDFFE_PN0P__3630  (.L_HI(net3630));
 sg13g2_tiehi \cpu.uart.r_xstate[2]$_SDFFE_PN0P__3631  (.L_HI(net3631));
 sg13g2_tiehi \cpu.uart.r_xstate[3]$_SDFFE_PN0P__3632  (.L_HI(net3632));
 sg13g2_tiehi \r_reset$_DFF_P__3633  (.L_HI(net3633));
 sg13g2_buf_8 clkbuf_leaf_1_clk (.A(clknet_6_1__leaf_clk),
    .X(clknet_leaf_1_clk));
 sg13g2_buf_8 clkbuf_leaf_2_clk (.A(clknet_6_1__leaf_clk),
    .X(clknet_leaf_2_clk));
 sg13g2_buf_8 clkbuf_leaf_3_clk (.A(clknet_6_4__leaf_clk),
    .X(clknet_leaf_3_clk));
 sg13g2_buf_8 clkbuf_leaf_4_clk (.A(clknet_6_4__leaf_clk),
    .X(clknet_leaf_4_clk));
 sg13g2_buf_8 clkbuf_leaf_5_clk (.A(clknet_6_4__leaf_clk),
    .X(clknet_leaf_5_clk));
 sg13g2_buf_8 clkbuf_leaf_6_clk (.A(clknet_6_4__leaf_clk),
    .X(clknet_leaf_6_clk));
 sg13g2_buf_8 clkbuf_leaf_7_clk (.A(clknet_6_1__leaf_clk),
    .X(clknet_leaf_7_clk));
 sg13g2_buf_8 clkbuf_leaf_8_clk (.A(clknet_6_1__leaf_clk),
    .X(clknet_leaf_8_clk));
 sg13g2_buf_8 clkbuf_leaf_9_clk (.A(clknet_6_3__leaf_clk),
    .X(clknet_leaf_9_clk));
 sg13g2_buf_8 clkbuf_leaf_10_clk (.A(clknet_6_6__leaf_clk),
    .X(clknet_leaf_10_clk));
 sg13g2_buf_8 clkbuf_leaf_11_clk (.A(clknet_6_3__leaf_clk),
    .X(clknet_leaf_11_clk));
 sg13g2_buf_8 clkbuf_leaf_12_clk (.A(clknet_6_7__leaf_clk),
    .X(clknet_leaf_12_clk));
 sg13g2_buf_8 clkbuf_leaf_13_clk (.A(clknet_6_4__leaf_clk),
    .X(clknet_leaf_13_clk));
 sg13g2_buf_8 clkbuf_leaf_14_clk (.A(clknet_6_5__leaf_clk),
    .X(clknet_leaf_14_clk));
 sg13g2_buf_8 clkbuf_leaf_15_clk (.A(clknet_6_5__leaf_clk),
    .X(clknet_leaf_15_clk));
 sg13g2_buf_8 clkbuf_leaf_16_clk (.A(clknet_6_7__leaf_clk),
    .X(clknet_leaf_16_clk));
 sg13g2_buf_8 clkbuf_leaf_17_clk (.A(clknet_6_5__leaf_clk),
    .X(clknet_leaf_17_clk));
 sg13g2_buf_8 clkbuf_leaf_18_clk (.A(clknet_6_5__leaf_clk),
    .X(clknet_leaf_18_clk));
 sg13g2_buf_8 clkbuf_leaf_19_clk (.A(clknet_6_5__leaf_clk),
    .X(clknet_leaf_19_clk));
 sg13g2_buf_8 clkbuf_leaf_20_clk (.A(clknet_6_7__leaf_clk),
    .X(clknet_leaf_20_clk));
 sg13g2_buf_8 clkbuf_leaf_21_clk (.A(clknet_6_7__leaf_clk),
    .X(clknet_leaf_21_clk));
 sg13g2_buf_8 clkbuf_leaf_22_clk (.A(clknet_6_7__leaf_clk),
    .X(clknet_leaf_22_clk));
 sg13g2_buf_8 clkbuf_leaf_23_clk (.A(clknet_6_18__leaf_clk),
    .X(clknet_leaf_23_clk));
 sg13g2_buf_8 clkbuf_leaf_24_clk (.A(clknet_6_18__leaf_clk),
    .X(clknet_leaf_24_clk));
 sg13g2_buf_8 clkbuf_leaf_25_clk (.A(clknet_6_6__leaf_clk),
    .X(clknet_leaf_25_clk));
 sg13g2_buf_8 clkbuf_leaf_26_clk (.A(clknet_6_6__leaf_clk),
    .X(clknet_leaf_26_clk));
 sg13g2_buf_8 clkbuf_leaf_27_clk (.A(clknet_6_6__leaf_clk),
    .X(clknet_leaf_27_clk));
 sg13g2_buf_8 clkbuf_leaf_28_clk (.A(clknet_6_6__leaf_clk),
    .X(clknet_leaf_28_clk));
 sg13g2_buf_8 clkbuf_leaf_29_clk (.A(clknet_6_12__leaf_clk),
    .X(clknet_leaf_29_clk));
 sg13g2_buf_8 clkbuf_leaf_30_clk (.A(clknet_6_13__leaf_clk),
    .X(clknet_leaf_30_clk));
 sg13g2_buf_8 clkbuf_leaf_31_clk (.A(clknet_6_13__leaf_clk),
    .X(clknet_leaf_31_clk));
 sg13g2_buf_8 clkbuf_leaf_32_clk (.A(clknet_6_13__leaf_clk),
    .X(clknet_leaf_32_clk));
 sg13g2_buf_8 clkbuf_leaf_33_clk (.A(clknet_6_24__leaf_clk),
    .X(clknet_leaf_33_clk));
 sg13g2_buf_8 clkbuf_leaf_34_clk (.A(clknet_6_24__leaf_clk),
    .X(clknet_leaf_34_clk));
 sg13g2_buf_8 clkbuf_leaf_35_clk (.A(clknet_6_13__leaf_clk),
    .X(clknet_leaf_35_clk));
 sg13g2_buf_8 clkbuf_leaf_36_clk (.A(clknet_6_13__leaf_clk),
    .X(clknet_leaf_36_clk));
 sg13g2_buf_8 clkbuf_leaf_37_clk (.A(clknet_6_15__leaf_clk),
    .X(clknet_leaf_37_clk));
 sg13g2_buf_8 clkbuf_leaf_38_clk (.A(clknet_6_15__leaf_clk),
    .X(clknet_leaf_38_clk));
 sg13g2_buf_8 clkbuf_leaf_39_clk (.A(clknet_6_15__leaf_clk),
    .X(clknet_leaf_39_clk));
 sg13g2_buf_8 clkbuf_leaf_40_clk (.A(clknet_6_15__leaf_clk),
    .X(clknet_leaf_40_clk));
 sg13g2_buf_8 clkbuf_leaf_41_clk (.A(clknet_6_36__leaf_clk),
    .X(clknet_leaf_41_clk));
 sg13g2_buf_8 clkbuf_leaf_42_clk (.A(clknet_6_26__leaf_clk),
    .X(clknet_leaf_42_clk));
 sg13g2_buf_8 clkbuf_leaf_43_clk (.A(clknet_6_26__leaf_clk),
    .X(clknet_leaf_43_clk));
 sg13g2_buf_8 clkbuf_leaf_44_clk (.A(clknet_6_26__leaf_clk),
    .X(clknet_leaf_44_clk));
 sg13g2_buf_8 clkbuf_leaf_45_clk (.A(clknet_6_24__leaf_clk),
    .X(clknet_leaf_45_clk));
 sg13g2_buf_8 clkbuf_leaf_46_clk (.A(clknet_6_24__leaf_clk),
    .X(clknet_leaf_46_clk));
 sg13g2_buf_8 clkbuf_leaf_47_clk (.A(clknet_6_24__leaf_clk),
    .X(clknet_leaf_47_clk));
 sg13g2_buf_8 clkbuf_leaf_48_clk (.A(clknet_6_25__leaf_clk),
    .X(clknet_leaf_48_clk));
 sg13g2_buf_8 clkbuf_leaf_49_clk (.A(clknet_6_25__leaf_clk),
    .X(clknet_leaf_49_clk));
 sg13g2_buf_8 clkbuf_leaf_50_clk (.A(clknet_6_25__leaf_clk),
    .X(clknet_leaf_50_clk));
 sg13g2_buf_8 clkbuf_leaf_51_clk (.A(clknet_6_19__leaf_clk),
    .X(clknet_leaf_51_clk));
 sg13g2_buf_8 clkbuf_leaf_52_clk (.A(clknet_6_19__leaf_clk),
    .X(clknet_leaf_52_clk));
 sg13g2_buf_8 clkbuf_leaf_53_clk (.A(clknet_6_18__leaf_clk),
    .X(clknet_leaf_53_clk));
 sg13g2_buf_8 clkbuf_leaf_54_clk (.A(clknet_6_18__leaf_clk),
    .X(clknet_leaf_54_clk));
 sg13g2_buf_8 clkbuf_leaf_55_clk (.A(clknet_6_18__leaf_clk),
    .X(clknet_leaf_55_clk));
 sg13g2_buf_8 clkbuf_leaf_56_clk (.A(clknet_6_16__leaf_clk),
    .X(clknet_leaf_56_clk));
 sg13g2_buf_8 clkbuf_leaf_57_clk (.A(clknet_6_16__leaf_clk),
    .X(clknet_leaf_57_clk));
 sg13g2_buf_8 clkbuf_leaf_58_clk (.A(clknet_6_16__leaf_clk),
    .X(clknet_leaf_58_clk));
 sg13g2_buf_8 clkbuf_leaf_59_clk (.A(clknet_6_17__leaf_clk),
    .X(clknet_leaf_59_clk));
 sg13g2_buf_8 clkbuf_leaf_60_clk (.A(clknet_6_16__leaf_clk),
    .X(clknet_leaf_60_clk));
 sg13g2_buf_8 clkbuf_leaf_61_clk (.A(clknet_6_16__leaf_clk),
    .X(clknet_leaf_61_clk));
 sg13g2_buf_8 clkbuf_leaf_62_clk (.A(clknet_6_17__leaf_clk),
    .X(clknet_leaf_62_clk));
 sg13g2_buf_8 clkbuf_leaf_63_clk (.A(clknet_6_17__leaf_clk),
    .X(clknet_leaf_63_clk));
 sg13g2_buf_8 clkbuf_leaf_64_clk (.A(clknet_6_17__leaf_clk),
    .X(clknet_leaf_64_clk));
 sg13g2_buf_8 clkbuf_leaf_65_clk (.A(clknet_6_19__leaf_clk),
    .X(clknet_leaf_65_clk));
 sg13g2_buf_8 clkbuf_leaf_66_clk (.A(clknet_6_19__leaf_clk),
    .X(clknet_leaf_66_clk));
 sg13g2_buf_8 clkbuf_leaf_67_clk (.A(clknet_6_19__leaf_clk),
    .X(clknet_leaf_67_clk));
 sg13g2_buf_8 clkbuf_leaf_68_clk (.A(clknet_6_17__leaf_clk),
    .X(clknet_leaf_68_clk));
 sg13g2_buf_8 clkbuf_leaf_69_clk (.A(clknet_6_20__leaf_clk),
    .X(clknet_leaf_69_clk));
 sg13g2_buf_8 clkbuf_leaf_70_clk (.A(clknet_6_20__leaf_clk),
    .X(clknet_leaf_70_clk));
 sg13g2_buf_8 clkbuf_leaf_71_clk (.A(clknet_6_20__leaf_clk),
    .X(clknet_leaf_71_clk));
 sg13g2_buf_8 clkbuf_leaf_72_clk (.A(clknet_6_20__leaf_clk),
    .X(clknet_leaf_72_clk));
 sg13g2_buf_8 clkbuf_leaf_73_clk (.A(clknet_6_20__leaf_clk),
    .X(clknet_leaf_73_clk));
 sg13g2_buf_8 clkbuf_leaf_74_clk (.A(clknet_6_21__leaf_clk),
    .X(clknet_leaf_74_clk));
 sg13g2_buf_8 clkbuf_leaf_75_clk (.A(clknet_6_21__leaf_clk),
    .X(clknet_leaf_75_clk));
 sg13g2_buf_8 clkbuf_leaf_76_clk (.A(clknet_6_21__leaf_clk),
    .X(clknet_leaf_76_clk));
 sg13g2_buf_8 clkbuf_leaf_77_clk (.A(clknet_6_21__leaf_clk),
    .X(clknet_leaf_77_clk));
 sg13g2_buf_8 clkbuf_leaf_78_clk (.A(clknet_6_21__leaf_clk),
    .X(clknet_leaf_78_clk));
 sg13g2_buf_8 clkbuf_leaf_79_clk (.A(clknet_6_23__leaf_clk),
    .X(clknet_leaf_79_clk));
 sg13g2_buf_8 clkbuf_leaf_80_clk (.A(clknet_6_23__leaf_clk),
    .X(clknet_leaf_80_clk));
 sg13g2_buf_8 clkbuf_leaf_81_clk (.A(clknet_6_23__leaf_clk),
    .X(clknet_leaf_81_clk));
 sg13g2_buf_8 clkbuf_leaf_82_clk (.A(clknet_6_22__leaf_clk),
    .X(clknet_leaf_82_clk));
 sg13g2_buf_8 clkbuf_leaf_83_clk (.A(clknet_6_23__leaf_clk),
    .X(clknet_leaf_83_clk));
 sg13g2_buf_8 clkbuf_leaf_84_clk (.A(clknet_6_22__leaf_clk),
    .X(clknet_leaf_84_clk));
 sg13g2_buf_8 clkbuf_leaf_85_clk (.A(clknet_6_22__leaf_clk),
    .X(clknet_leaf_85_clk));
 sg13g2_buf_8 clkbuf_leaf_86_clk (.A(clknet_6_22__leaf_clk),
    .X(clknet_leaf_86_clk));
 sg13g2_buf_8 clkbuf_leaf_87_clk (.A(clknet_6_22__leaf_clk),
    .X(clknet_leaf_87_clk));
 sg13g2_buf_8 clkbuf_leaf_88_clk (.A(clknet_6_28__leaf_clk),
    .X(clknet_leaf_88_clk));
 sg13g2_buf_8 clkbuf_leaf_89_clk (.A(clknet_6_29__leaf_clk),
    .X(clknet_leaf_89_clk));
 sg13g2_buf_8 clkbuf_leaf_90_clk (.A(clknet_6_28__leaf_clk),
    .X(clknet_leaf_90_clk));
 sg13g2_buf_8 clkbuf_leaf_91_clk (.A(clknet_6_28__leaf_clk),
    .X(clknet_leaf_91_clk));
 sg13g2_buf_8 clkbuf_leaf_92_clk (.A(clknet_6_28__leaf_clk),
    .X(clknet_leaf_92_clk));
 sg13g2_buf_8 clkbuf_leaf_93_clk (.A(clknet_6_28__leaf_clk),
    .X(clknet_leaf_93_clk));
 sg13g2_buf_8 clkbuf_leaf_94_clk (.A(clknet_6_29__leaf_clk),
    .X(clknet_leaf_94_clk));
 sg13g2_buf_8 clkbuf_leaf_95_clk (.A(clknet_6_29__leaf_clk),
    .X(clknet_leaf_95_clk));
 sg13g2_buf_8 clkbuf_leaf_96_clk (.A(clknet_6_29__leaf_clk),
    .X(clknet_leaf_96_clk));
 sg13g2_buf_8 clkbuf_leaf_97_clk (.A(clknet_6_29__leaf_clk),
    .X(clknet_leaf_97_clk));
 sg13g2_buf_8 clkbuf_leaf_98_clk (.A(clknet_6_31__leaf_clk),
    .X(clknet_leaf_98_clk));
 sg13g2_buf_8 clkbuf_leaf_99_clk (.A(clknet_6_31__leaf_clk),
    .X(clknet_leaf_99_clk));
 sg13g2_buf_8 clkbuf_leaf_100_clk (.A(clknet_6_31__leaf_clk),
    .X(clknet_leaf_100_clk));
 sg13g2_buf_8 clkbuf_leaf_101_clk (.A(clknet_6_31__leaf_clk),
    .X(clknet_leaf_101_clk));
 sg13g2_buf_8 clkbuf_leaf_102_clk (.A(clknet_6_30__leaf_clk),
    .X(clknet_leaf_102_clk));
 sg13g2_buf_8 clkbuf_leaf_103_clk (.A(clknet_6_30__leaf_clk),
    .X(clknet_leaf_103_clk));
 sg13g2_buf_8 clkbuf_leaf_104_clk (.A(clknet_6_30__leaf_clk),
    .X(clknet_leaf_104_clk));
 sg13g2_buf_8 clkbuf_leaf_105_clk (.A(clknet_6_30__leaf_clk),
    .X(clknet_leaf_105_clk));
 sg13g2_buf_8 clkbuf_leaf_106_clk (.A(clknet_6_27__leaf_clk),
    .X(clknet_leaf_106_clk));
 sg13g2_buf_8 clkbuf_leaf_107_clk (.A(clknet_6_25__leaf_clk),
    .X(clknet_leaf_107_clk));
 sg13g2_buf_8 clkbuf_leaf_108_clk (.A(clknet_6_25__leaf_clk),
    .X(clknet_leaf_108_clk));
 sg13g2_buf_8 clkbuf_leaf_109_clk (.A(clknet_6_27__leaf_clk),
    .X(clknet_leaf_109_clk));
 sg13g2_buf_8 clkbuf_leaf_110_clk (.A(clknet_6_27__leaf_clk),
    .X(clknet_leaf_110_clk));
 sg13g2_buf_8 clkbuf_leaf_111_clk (.A(clknet_6_27__leaf_clk),
    .X(clknet_leaf_111_clk));
 sg13g2_buf_8 clkbuf_leaf_112_clk (.A(clknet_6_30__leaf_clk),
    .X(clknet_leaf_112_clk));
 sg13g2_buf_8 clkbuf_leaf_113_clk (.A(clknet_6_27__leaf_clk),
    .X(clknet_leaf_113_clk));
 sg13g2_buf_8 clkbuf_leaf_114_clk (.A(clknet_6_26__leaf_clk),
    .X(clknet_leaf_114_clk));
 sg13g2_buf_8 clkbuf_leaf_115_clk (.A(clknet_6_26__leaf_clk),
    .X(clknet_leaf_115_clk));
 sg13g2_buf_8 clkbuf_leaf_116_clk (.A(clknet_6_36__leaf_clk),
    .X(clknet_leaf_116_clk));
 sg13g2_buf_8 clkbuf_leaf_117_clk (.A(clknet_6_39__leaf_clk),
    .X(clknet_leaf_117_clk));
 sg13g2_buf_8 clkbuf_leaf_118_clk (.A(clknet_6_37__leaf_clk),
    .X(clknet_leaf_118_clk));
 sg13g2_buf_8 clkbuf_leaf_119_clk (.A(clknet_6_39__leaf_clk),
    .X(clknet_leaf_119_clk));
 sg13g2_buf_8 clkbuf_leaf_120_clk (.A(clknet_6_45__leaf_clk),
    .X(clknet_leaf_120_clk));
 sg13g2_buf_8 clkbuf_leaf_121_clk (.A(clknet_6_39__leaf_clk),
    .X(clknet_leaf_121_clk));
 sg13g2_buf_8 clkbuf_leaf_122_clk (.A(clknet_6_37__leaf_clk),
    .X(clknet_leaf_122_clk));
 sg13g2_buf_8 clkbuf_leaf_123_clk (.A(clknet_6_37__leaf_clk),
    .X(clknet_leaf_123_clk));
 sg13g2_buf_8 clkbuf_leaf_124_clk (.A(clknet_6_37__leaf_clk),
    .X(clknet_leaf_124_clk));
 sg13g2_buf_8 clkbuf_leaf_125_clk (.A(clknet_6_37__leaf_clk),
    .X(clknet_leaf_125_clk));
 sg13g2_buf_8 clkbuf_leaf_126_clk (.A(clknet_6_39__leaf_clk),
    .X(clknet_leaf_126_clk));
 sg13g2_buf_8 clkbuf_leaf_127_clk (.A(clknet_6_45__leaf_clk),
    .X(clknet_leaf_127_clk));
 sg13g2_buf_8 clkbuf_leaf_128_clk (.A(clknet_6_45__leaf_clk),
    .X(clknet_leaf_128_clk));
 sg13g2_buf_8 clkbuf_leaf_129_clk (.A(clknet_6_60__leaf_clk),
    .X(clknet_leaf_129_clk));
 sg13g2_buf_8 clkbuf_leaf_130_clk (.A(clknet_6_60__leaf_clk),
    .X(clknet_leaf_130_clk));
 sg13g2_buf_8 clkbuf_leaf_131_clk (.A(clknet_6_61__leaf_clk),
    .X(clknet_leaf_131_clk));
 sg13g2_buf_8 clkbuf_leaf_132_clk (.A(clknet_6_60__leaf_clk),
    .X(clknet_leaf_132_clk));
 sg13g2_buf_8 clkbuf_leaf_133_clk (.A(clknet_6_61__leaf_clk),
    .X(clknet_leaf_133_clk));
 sg13g2_buf_8 clkbuf_leaf_134_clk (.A(clknet_6_61__leaf_clk),
    .X(clknet_leaf_134_clk));
 sg13g2_buf_8 clkbuf_leaf_135_clk (.A(clknet_6_61__leaf_clk),
    .X(clknet_leaf_135_clk));
 sg13g2_buf_8 clkbuf_leaf_136_clk (.A(clknet_6_61__leaf_clk),
    .X(clknet_leaf_136_clk));
 sg13g2_buf_8 clkbuf_leaf_137_clk (.A(clknet_6_63__leaf_clk),
    .X(clknet_leaf_137_clk));
 sg13g2_buf_8 clkbuf_leaf_138_clk (.A(clknet_6_57__leaf_clk),
    .X(clknet_leaf_138_clk));
 sg13g2_buf_8 clkbuf_leaf_139_clk (.A(clknet_6_56__leaf_clk),
    .X(clknet_leaf_139_clk));
 sg13g2_buf_8 clkbuf_leaf_140_clk (.A(clknet_6_57__leaf_clk),
    .X(clknet_leaf_140_clk));
 sg13g2_buf_8 clkbuf_leaf_141_clk (.A(clknet_6_57__leaf_clk),
    .X(clknet_leaf_141_clk));
 sg13g2_buf_8 clkbuf_leaf_142_clk (.A(clknet_6_56__leaf_clk),
    .X(clknet_leaf_142_clk));
 sg13g2_buf_8 clkbuf_leaf_143_clk (.A(clknet_6_57__leaf_clk),
    .X(clknet_leaf_143_clk));
 sg13g2_buf_8 clkbuf_leaf_144_clk (.A(clknet_6_57__leaf_clk),
    .X(clknet_leaf_144_clk));
 sg13g2_buf_8 clkbuf_leaf_145_clk (.A(clknet_6_59__leaf_clk),
    .X(clknet_leaf_145_clk));
 sg13g2_buf_8 clkbuf_leaf_146_clk (.A(clknet_6_59__leaf_clk),
    .X(clknet_leaf_146_clk));
 sg13g2_buf_8 clkbuf_leaf_147_clk (.A(clknet_6_56__leaf_clk),
    .X(clknet_leaf_147_clk));
 sg13g2_buf_8 clkbuf_leaf_148_clk (.A(clknet_6_56__leaf_clk),
    .X(clknet_leaf_148_clk));
 sg13g2_buf_8 clkbuf_leaf_149_clk (.A(clknet_6_63__leaf_clk),
    .X(clknet_leaf_149_clk));
 sg13g2_buf_8 clkbuf_leaf_150_clk (.A(clknet_6_63__leaf_clk),
    .X(clknet_leaf_150_clk));
 sg13g2_buf_8 clkbuf_leaf_151_clk (.A(clknet_6_60__leaf_clk),
    .X(clknet_leaf_151_clk));
 sg13g2_buf_8 clkbuf_leaf_152_clk (.A(clknet_6_63__leaf_clk),
    .X(clknet_leaf_152_clk));
 sg13g2_buf_8 clkbuf_leaf_153_clk (.A(clknet_6_62__leaf_clk),
    .X(clknet_leaf_153_clk));
 sg13g2_buf_8 clkbuf_leaf_154_clk (.A(clknet_6_58__leaf_clk),
    .X(clknet_leaf_154_clk));
 sg13g2_buf_8 clkbuf_leaf_155_clk (.A(clknet_6_56__leaf_clk),
    .X(clknet_leaf_155_clk));
 sg13g2_buf_8 clkbuf_leaf_156_clk (.A(clknet_6_59__leaf_clk),
    .X(clknet_leaf_156_clk));
 sg13g2_buf_8 clkbuf_leaf_157_clk (.A(clknet_6_59__leaf_clk),
    .X(clknet_leaf_157_clk));
 sg13g2_buf_8 clkbuf_leaf_158_clk (.A(clknet_6_58__leaf_clk),
    .X(clknet_leaf_158_clk));
 sg13g2_buf_8 clkbuf_leaf_159_clk (.A(clknet_6_59__leaf_clk),
    .X(clknet_leaf_159_clk));
 sg13g2_buf_8 clkbuf_leaf_160_clk (.A(clknet_6_58__leaf_clk),
    .X(clknet_leaf_160_clk));
 sg13g2_buf_8 clkbuf_leaf_161_clk (.A(clknet_6_58__leaf_clk),
    .X(clknet_leaf_161_clk));
 sg13g2_buf_8 clkbuf_leaf_162_clk (.A(clknet_6_58__leaf_clk),
    .X(clknet_leaf_162_clk));
 sg13g2_buf_8 clkbuf_leaf_163_clk (.A(clknet_6_55__leaf_clk),
    .X(clknet_leaf_163_clk));
 sg13g2_buf_8 clkbuf_leaf_164_clk (.A(clknet_6_53__leaf_clk),
    .X(clknet_leaf_164_clk));
 sg13g2_buf_8 clkbuf_leaf_165_clk (.A(clknet_6_52__leaf_clk),
    .X(clknet_leaf_165_clk));
 sg13g2_buf_8 clkbuf_leaf_166_clk (.A(clknet_6_62__leaf_clk),
    .X(clknet_leaf_166_clk));
 sg13g2_buf_8 clkbuf_leaf_167_clk (.A(clknet_6_62__leaf_clk),
    .X(clknet_leaf_167_clk));
 sg13g2_buf_8 clkbuf_leaf_168_clk (.A(clknet_6_47__leaf_clk),
    .X(clknet_leaf_168_clk));
 sg13g2_buf_8 clkbuf_leaf_169_clk (.A(clknet_6_47__leaf_clk),
    .X(clknet_leaf_169_clk));
 sg13g2_buf_8 clkbuf_leaf_170_clk (.A(clknet_6_62__leaf_clk),
    .X(clknet_leaf_170_clk));
 sg13g2_buf_8 clkbuf_leaf_171_clk (.A(clknet_6_62__leaf_clk),
    .X(clknet_leaf_171_clk));
 sg13g2_buf_8 clkbuf_leaf_172_clk (.A(clknet_6_60__leaf_clk),
    .X(clknet_leaf_172_clk));
 sg13g2_buf_8 clkbuf_leaf_173_clk (.A(clknet_6_45__leaf_clk),
    .X(clknet_leaf_173_clk));
 sg13g2_buf_8 clkbuf_leaf_174_clk (.A(clknet_6_44__leaf_clk),
    .X(clknet_leaf_174_clk));
 sg13g2_buf_8 clkbuf_leaf_175_clk (.A(clknet_6_45__leaf_clk),
    .X(clknet_leaf_175_clk));
 sg13g2_buf_8 clkbuf_leaf_176_clk (.A(clknet_6_38__leaf_clk),
    .X(clknet_leaf_176_clk));
 sg13g2_buf_8 clkbuf_leaf_177_clk (.A(clknet_6_36__leaf_clk),
    .X(clknet_leaf_177_clk));
 sg13g2_buf_8 clkbuf_leaf_178_clk (.A(clknet_6_38__leaf_clk),
    .X(clknet_leaf_178_clk));
 sg13g2_buf_8 clkbuf_leaf_179_clk (.A(clknet_6_38__leaf_clk),
    .X(clknet_leaf_179_clk));
 sg13g2_buf_8 clkbuf_leaf_180_clk (.A(clknet_6_38__leaf_clk),
    .X(clknet_leaf_180_clk));
 sg13g2_buf_8 clkbuf_leaf_181_clk (.A(clknet_6_44__leaf_clk),
    .X(clknet_leaf_181_clk));
 sg13g2_buf_8 clkbuf_leaf_182_clk (.A(clknet_6_44__leaf_clk),
    .X(clknet_leaf_182_clk));
 sg13g2_buf_8 clkbuf_leaf_183_clk (.A(clknet_6_44__leaf_clk),
    .X(clknet_leaf_183_clk));
 sg13g2_buf_8 clkbuf_leaf_184_clk (.A(clknet_6_44__leaf_clk),
    .X(clknet_leaf_184_clk));
 sg13g2_buf_8 clkbuf_leaf_185_clk (.A(clknet_6_41__leaf_clk),
    .X(clknet_leaf_185_clk));
 sg13g2_buf_8 clkbuf_leaf_186_clk (.A(clknet_6_46__leaf_clk),
    .X(clknet_leaf_186_clk));
 sg13g2_buf_8 clkbuf_leaf_187_clk (.A(clknet_6_46__leaf_clk),
    .X(clknet_leaf_187_clk));
 sg13g2_buf_8 clkbuf_leaf_188_clk (.A(clknet_6_46__leaf_clk),
    .X(clknet_leaf_188_clk));
 sg13g2_buf_8 clkbuf_leaf_189_clk (.A(clknet_6_52__leaf_clk),
    .X(clknet_leaf_189_clk));
 sg13g2_buf_8 clkbuf_leaf_190_clk (.A(clknet_6_46__leaf_clk),
    .X(clknet_leaf_190_clk));
 sg13g2_buf_8 clkbuf_leaf_191_clk (.A(clknet_6_46__leaf_clk),
    .X(clknet_leaf_191_clk));
 sg13g2_buf_8 clkbuf_leaf_192_clk (.A(clknet_6_47__leaf_clk),
    .X(clknet_leaf_192_clk));
 sg13g2_buf_8 clkbuf_leaf_193_clk (.A(clknet_6_47__leaf_clk),
    .X(clknet_leaf_193_clk));
 sg13g2_buf_8 clkbuf_leaf_194_clk (.A(clknet_6_52__leaf_clk),
    .X(clknet_leaf_194_clk));
 sg13g2_buf_8 clkbuf_leaf_195_clk (.A(clknet_6_52__leaf_clk),
    .X(clknet_leaf_195_clk));
 sg13g2_buf_8 clkbuf_leaf_196_clk (.A(clknet_6_53__leaf_clk),
    .X(clknet_leaf_196_clk));
 sg13g2_buf_8 clkbuf_leaf_197_clk (.A(clknet_6_53__leaf_clk),
    .X(clknet_leaf_197_clk));
 sg13g2_buf_8 clkbuf_leaf_198_clk (.A(clknet_6_55__leaf_clk),
    .X(clknet_leaf_198_clk));
 sg13g2_buf_8 clkbuf_leaf_199_clk (.A(clknet_6_55__leaf_clk),
    .X(clknet_leaf_199_clk));
 sg13g2_buf_8 clkbuf_leaf_200_clk (.A(clknet_6_55__leaf_clk),
    .X(clknet_leaf_200_clk));
 sg13g2_buf_8 clkbuf_leaf_201_clk (.A(clknet_6_53__leaf_clk),
    .X(clknet_leaf_201_clk));
 sg13g2_buf_8 clkbuf_leaf_202_clk (.A(clknet_6_54__leaf_clk),
    .X(clknet_leaf_202_clk));
 sg13g2_buf_8 clkbuf_leaf_203_clk (.A(clknet_6_54__leaf_clk),
    .X(clknet_leaf_203_clk));
 sg13g2_buf_8 clkbuf_leaf_204_clk (.A(clknet_6_54__leaf_clk),
    .X(clknet_leaf_204_clk));
 sg13g2_buf_8 clkbuf_leaf_205_clk (.A(clknet_6_54__leaf_clk),
    .X(clknet_leaf_205_clk));
 sg13g2_buf_8 clkbuf_leaf_206_clk (.A(clknet_6_54__leaf_clk),
    .X(clknet_leaf_206_clk));
 sg13g2_buf_8 clkbuf_leaf_207_clk (.A(clknet_6_53__leaf_clk),
    .X(clknet_leaf_207_clk));
 sg13g2_buf_8 clkbuf_leaf_208_clk (.A(clknet_6_52__leaf_clk),
    .X(clknet_leaf_208_clk));
 sg13g2_buf_8 clkbuf_leaf_209_clk (.A(clknet_6_49__leaf_clk),
    .X(clknet_leaf_209_clk));
 sg13g2_buf_8 clkbuf_leaf_210_clk (.A(clknet_6_43__leaf_clk),
    .X(clknet_leaf_210_clk));
 sg13g2_buf_8 clkbuf_leaf_211_clk (.A(clknet_6_49__leaf_clk),
    .X(clknet_leaf_211_clk));
 sg13g2_buf_8 clkbuf_leaf_212_clk (.A(clknet_6_51__leaf_clk),
    .X(clknet_leaf_212_clk));
 sg13g2_buf_8 clkbuf_leaf_213_clk (.A(clknet_6_51__leaf_clk),
    .X(clknet_leaf_213_clk));
 sg13g2_buf_8 clkbuf_leaf_214_clk (.A(clknet_6_51__leaf_clk),
    .X(clknet_leaf_214_clk));
 sg13g2_buf_8 clkbuf_leaf_215_clk (.A(clknet_6_51__leaf_clk),
    .X(clknet_leaf_215_clk));
 sg13g2_buf_8 clkbuf_leaf_216_clk (.A(clknet_6_50__leaf_clk),
    .X(clknet_leaf_216_clk));
 sg13g2_buf_8 clkbuf_leaf_217_clk (.A(clknet_6_50__leaf_clk),
    .X(clknet_leaf_217_clk));
 sg13g2_buf_8 clkbuf_leaf_218_clk (.A(clknet_6_50__leaf_clk),
    .X(clknet_leaf_218_clk));
 sg13g2_buf_8 clkbuf_leaf_219_clk (.A(clknet_6_51__leaf_clk),
    .X(clknet_leaf_219_clk));
 sg13g2_buf_8 clkbuf_leaf_220_clk (.A(clknet_6_50__leaf_clk),
    .X(clknet_leaf_220_clk));
 sg13g2_buf_8 clkbuf_leaf_221_clk (.A(clknet_6_50__leaf_clk),
    .X(clknet_leaf_221_clk));
 sg13g2_buf_8 clkbuf_leaf_222_clk (.A(clknet_6_48__leaf_clk),
    .X(clknet_leaf_222_clk));
 sg13g2_buf_8 clkbuf_leaf_223_clk (.A(clknet_6_48__leaf_clk),
    .X(clknet_leaf_223_clk));
 sg13g2_buf_8 clkbuf_leaf_224_clk (.A(clknet_6_49__leaf_clk),
    .X(clknet_leaf_224_clk));
 sg13g2_buf_8 clkbuf_leaf_225_clk (.A(clknet_6_48__leaf_clk),
    .X(clknet_leaf_225_clk));
 sg13g2_buf_8 clkbuf_leaf_226_clk (.A(clknet_6_48__leaf_clk),
    .X(clknet_leaf_226_clk));
 sg13g2_buf_8 clkbuf_leaf_227_clk (.A(clknet_6_48__leaf_clk),
    .X(clknet_leaf_227_clk));
 sg13g2_buf_8 clkbuf_leaf_228_clk (.A(clknet_6_49__leaf_clk),
    .X(clknet_leaf_228_clk));
 sg13g2_buf_8 clkbuf_leaf_229_clk (.A(clknet_6_49__leaf_clk),
    .X(clknet_leaf_229_clk));
 sg13g2_buf_8 clkbuf_leaf_230_clk (.A(clknet_6_43__leaf_clk),
    .X(clknet_leaf_230_clk));
 sg13g2_buf_8 clkbuf_leaf_231_clk (.A(clknet_6_43__leaf_clk),
    .X(clknet_leaf_231_clk));
 sg13g2_buf_8 clkbuf_leaf_232_clk (.A(clknet_6_42__leaf_clk),
    .X(clknet_leaf_232_clk));
 sg13g2_buf_8 clkbuf_leaf_233_clk (.A(clknet_6_43__leaf_clk),
    .X(clknet_leaf_233_clk));
 sg13g2_buf_8 clkbuf_leaf_234_clk (.A(clknet_6_40__leaf_clk),
    .X(clknet_leaf_234_clk));
 sg13g2_buf_8 clkbuf_leaf_235_clk (.A(clknet_6_42__leaf_clk),
    .X(clknet_leaf_235_clk));
 sg13g2_buf_8 clkbuf_leaf_236_clk (.A(clknet_6_42__leaf_clk),
    .X(clknet_leaf_236_clk));
 sg13g2_buf_8 clkbuf_leaf_237_clk (.A(clknet_6_43__leaf_clk),
    .X(clknet_leaf_237_clk));
 sg13g2_buf_8 clkbuf_leaf_238_clk (.A(clknet_6_42__leaf_clk),
    .X(clknet_leaf_238_clk));
 sg13g2_buf_8 clkbuf_leaf_239_clk (.A(clknet_6_42__leaf_clk),
    .X(clknet_leaf_239_clk));
 sg13g2_buf_8 clkbuf_leaf_240_clk (.A(clknet_6_40__leaf_clk),
    .X(clknet_leaf_240_clk));
 sg13g2_buf_8 clkbuf_leaf_241_clk (.A(clknet_6_34__leaf_clk),
    .X(clknet_leaf_241_clk));
 sg13g2_buf_8 clkbuf_leaf_242_clk (.A(clknet_6_34__leaf_clk),
    .X(clknet_leaf_242_clk));
 sg13g2_buf_8 clkbuf_leaf_243_clk (.A(clknet_6_34__leaf_clk),
    .X(clknet_leaf_243_clk));
 sg13g2_buf_8 clkbuf_leaf_244_clk (.A(clknet_6_34__leaf_clk),
    .X(clknet_leaf_244_clk));
 sg13g2_buf_8 clkbuf_leaf_245_clk (.A(clknet_6_34__leaf_clk),
    .X(clknet_leaf_245_clk));
 sg13g2_buf_8 clkbuf_leaf_246_clk (.A(clknet_6_35__leaf_clk),
    .X(clknet_leaf_246_clk));
 sg13g2_buf_8 clkbuf_leaf_247_clk (.A(clknet_6_35__leaf_clk),
    .X(clknet_leaf_247_clk));
 sg13g2_buf_8 clkbuf_leaf_248_clk (.A(clknet_6_35__leaf_clk),
    .X(clknet_leaf_248_clk));
 sg13g2_buf_8 clkbuf_leaf_249_clk (.A(clknet_6_35__leaf_clk),
    .X(clknet_leaf_249_clk));
 sg13g2_buf_8 clkbuf_leaf_250_clk (.A(clknet_6_40__leaf_clk),
    .X(clknet_leaf_250_clk));
 sg13g2_buf_8 clkbuf_leaf_251_clk (.A(clknet_6_40__leaf_clk),
    .X(clknet_leaf_251_clk));
 sg13g2_buf_8 clkbuf_leaf_252_clk (.A(clknet_6_40__leaf_clk),
    .X(clknet_leaf_252_clk));
 sg13g2_buf_8 clkbuf_leaf_253_clk (.A(clknet_6_41__leaf_clk),
    .X(clknet_leaf_253_clk));
 sg13g2_buf_8 clkbuf_leaf_254_clk (.A(clknet_6_41__leaf_clk),
    .X(clknet_leaf_254_clk));
 sg13g2_buf_8 clkbuf_leaf_255_clk (.A(clknet_6_41__leaf_clk),
    .X(clknet_leaf_255_clk));
 sg13g2_buf_8 clkbuf_leaf_256_clk (.A(clknet_6_41__leaf_clk),
    .X(clknet_leaf_256_clk));
 sg13g2_buf_8 clkbuf_leaf_257_clk (.A(clknet_6_35__leaf_clk),
    .X(clknet_leaf_257_clk));
 sg13g2_buf_8 clkbuf_leaf_258_clk (.A(clknet_6_33__leaf_clk),
    .X(clknet_leaf_258_clk));
 sg13g2_buf_8 clkbuf_leaf_259_clk (.A(clknet_6_36__leaf_clk),
    .X(clknet_leaf_259_clk));
 sg13g2_buf_8 clkbuf_leaf_260_clk (.A(clknet_6_38__leaf_clk),
    .X(clknet_leaf_260_clk));
 sg13g2_buf_8 clkbuf_leaf_261_clk (.A(clknet_6_33__leaf_clk),
    .X(clknet_leaf_261_clk));
 sg13g2_buf_8 clkbuf_leaf_262_clk (.A(clknet_6_36__leaf_clk),
    .X(clknet_leaf_262_clk));
 sg13g2_buf_8 clkbuf_leaf_263_clk (.A(clknet_6_33__leaf_clk),
    .X(clknet_leaf_263_clk));
 sg13g2_buf_8 clkbuf_leaf_264_clk (.A(clknet_6_33__leaf_clk),
    .X(clknet_leaf_264_clk));
 sg13g2_buf_8 clkbuf_leaf_265_clk (.A(clknet_6_14__leaf_clk),
    .X(clknet_leaf_265_clk));
 sg13g2_buf_8 clkbuf_leaf_266_clk (.A(clknet_6_14__leaf_clk),
    .X(clknet_leaf_266_clk));
 sg13g2_buf_8 clkbuf_leaf_267_clk (.A(clknet_6_33__leaf_clk),
    .X(clknet_leaf_267_clk));
 sg13g2_buf_8 clkbuf_leaf_268_clk (.A(clknet_6_32__leaf_clk),
    .X(clknet_leaf_268_clk));
 sg13g2_buf_8 clkbuf_leaf_269_clk (.A(clknet_6_14__leaf_clk),
    .X(clknet_leaf_269_clk));
 sg13g2_buf_8 clkbuf_leaf_270_clk (.A(clknet_6_14__leaf_clk),
    .X(clknet_leaf_270_clk));
 sg13g2_buf_8 clkbuf_leaf_271_clk (.A(clknet_6_14__leaf_clk),
    .X(clknet_leaf_271_clk));
 sg13g2_buf_8 clkbuf_leaf_272_clk (.A(clknet_6_12__leaf_clk),
    .X(clknet_leaf_272_clk));
 sg13g2_buf_8 clkbuf_leaf_273_clk (.A(clknet_6_12__leaf_clk),
    .X(clknet_leaf_273_clk));
 sg13g2_buf_8 clkbuf_leaf_274_clk (.A(clknet_6_12__leaf_clk),
    .X(clknet_leaf_274_clk));
 sg13g2_buf_8 clkbuf_leaf_275_clk (.A(clknet_6_9__leaf_clk),
    .X(clknet_leaf_275_clk));
 sg13g2_buf_8 clkbuf_leaf_276_clk (.A(clknet_6_12__leaf_clk),
    .X(clknet_leaf_276_clk));
 sg13g2_buf_8 clkbuf_leaf_277_clk (.A(clknet_6_9__leaf_clk),
    .X(clknet_leaf_277_clk));
 sg13g2_buf_8 clkbuf_leaf_278_clk (.A(clknet_6_11__leaf_clk),
    .X(clknet_leaf_278_clk));
 sg13g2_buf_8 clkbuf_leaf_279_clk (.A(clknet_6_11__leaf_clk),
    .X(clknet_leaf_279_clk));
 sg13g2_buf_8 clkbuf_leaf_280_clk (.A(clknet_6_11__leaf_clk),
    .X(clknet_leaf_280_clk));
 sg13g2_buf_8 clkbuf_leaf_281_clk (.A(clknet_6_32__leaf_clk),
    .X(clknet_leaf_281_clk));
 sg13g2_buf_8 clkbuf_leaf_282_clk (.A(clknet_6_32__leaf_clk),
    .X(clknet_leaf_282_clk));
 sg13g2_buf_8 clkbuf_leaf_283_clk (.A(clknet_6_11__leaf_clk),
    .X(clknet_leaf_283_clk));
 sg13g2_buf_8 clkbuf_leaf_284_clk (.A(clknet_6_11__leaf_clk),
    .X(clknet_leaf_284_clk));
 sg13g2_buf_8 clkbuf_leaf_285_clk (.A(clknet_6_10__leaf_clk),
    .X(clknet_leaf_285_clk));
 sg13g2_buf_8 clkbuf_leaf_286_clk (.A(clknet_6_32__leaf_clk),
    .X(clknet_leaf_286_clk));
 sg13g2_buf_8 clkbuf_leaf_287_clk (.A(clknet_6_32__leaf_clk),
    .X(clknet_leaf_287_clk));
 sg13g2_buf_8 clkbuf_leaf_288_clk (.A(clknet_6_10__leaf_clk),
    .X(clknet_leaf_288_clk));
 sg13g2_buf_8 clkbuf_leaf_289_clk (.A(clknet_6_10__leaf_clk),
    .X(clknet_leaf_289_clk));
 sg13g2_buf_8 clkbuf_leaf_290_clk (.A(clknet_6_10__leaf_clk),
    .X(clknet_leaf_290_clk));
 sg13g2_buf_8 clkbuf_leaf_291_clk (.A(clknet_6_10__leaf_clk),
    .X(clknet_leaf_291_clk));
 sg13g2_buf_8 clkbuf_leaf_292_clk (.A(clknet_6_8__leaf_clk),
    .X(clknet_leaf_292_clk));
 sg13g2_buf_8 clkbuf_leaf_293_clk (.A(clknet_6_8__leaf_clk),
    .X(clknet_leaf_293_clk));
 sg13g2_buf_8 clkbuf_leaf_294_clk (.A(clknet_6_8__leaf_clk),
    .X(clknet_leaf_294_clk));
 sg13g2_buf_8 clkbuf_leaf_295_clk (.A(clknet_6_8__leaf_clk),
    .X(clknet_leaf_295_clk));
 sg13g2_buf_8 clkbuf_leaf_296_clk (.A(clknet_6_8__leaf_clk),
    .X(clknet_leaf_296_clk));
 sg13g2_buf_8 clkbuf_leaf_297_clk (.A(clknet_6_9__leaf_clk),
    .X(clknet_leaf_297_clk));
 sg13g2_buf_8 clkbuf_leaf_298_clk (.A(clknet_6_9__leaf_clk),
    .X(clknet_leaf_298_clk));
 sg13g2_buf_8 clkbuf_leaf_299_clk (.A(clknet_6_9__leaf_clk),
    .X(clknet_leaf_299_clk));
 sg13g2_buf_8 clkbuf_leaf_300_clk (.A(clknet_6_3__leaf_clk),
    .X(clknet_leaf_300_clk));
 sg13g2_buf_8 clkbuf_leaf_301_clk (.A(clknet_6_3__leaf_clk),
    .X(clknet_leaf_301_clk));
 sg13g2_buf_8 clkbuf_leaf_302_clk (.A(clknet_6_3__leaf_clk),
    .X(clknet_leaf_302_clk));
 sg13g2_buf_8 clkbuf_leaf_303_clk (.A(clknet_6_2__leaf_clk),
    .X(clknet_leaf_303_clk));
 sg13g2_buf_8 clkbuf_leaf_304_clk (.A(clknet_6_2__leaf_clk),
    .X(clknet_leaf_304_clk));
 sg13g2_buf_8 clkbuf_leaf_305_clk (.A(clknet_6_2__leaf_clk),
    .X(clknet_leaf_305_clk));
 sg13g2_buf_8 clkbuf_leaf_306_clk (.A(clknet_6_2__leaf_clk),
    .X(clknet_leaf_306_clk));
 sg13g2_buf_8 clkbuf_leaf_307_clk (.A(clknet_6_2__leaf_clk),
    .X(clknet_leaf_307_clk));
 sg13g2_buf_8 clkbuf_leaf_308_clk (.A(clknet_6_0__leaf_clk),
    .X(clknet_leaf_308_clk));
 sg13g2_buf_8 clkbuf_leaf_309_clk (.A(clknet_6_1__leaf_clk),
    .X(clknet_leaf_309_clk));
 sg13g2_buf_8 clkbuf_leaf_310_clk (.A(clknet_6_0__leaf_clk),
    .X(clknet_leaf_310_clk));
 sg13g2_buf_8 clkbuf_leaf_311_clk (.A(clknet_6_0__leaf_clk),
    .X(clknet_leaf_311_clk));
 sg13g2_buf_8 clkbuf_leaf_312_clk (.A(clknet_6_0__leaf_clk),
    .X(clknet_leaf_312_clk));
 sg13g2_buf_4 clkbuf_0_clk (.X(clknet_0_clk),
    .A(clk));
 sg13g2_buf_8 clkbuf_3_0_0_clk (.A(clknet_0_clk),
    .X(clknet_3_0_0_clk));
 sg13g2_buf_8 clkbuf_3_1_0_clk (.A(clknet_0_clk),
    .X(clknet_3_1_0_clk));
 sg13g2_buf_8 clkbuf_3_2_0_clk (.A(clknet_0_clk),
    .X(clknet_3_2_0_clk));
 sg13g2_buf_8 clkbuf_3_3_0_clk (.A(clknet_0_clk),
    .X(clknet_3_3_0_clk));
 sg13g2_buf_8 clkbuf_3_4_0_clk (.A(clknet_0_clk),
    .X(clknet_3_4_0_clk));
 sg13g2_buf_8 clkbuf_3_5_0_clk (.A(clknet_0_clk),
    .X(clknet_3_5_0_clk));
 sg13g2_buf_8 clkbuf_3_6_0_clk (.A(clknet_0_clk),
    .X(clknet_3_6_0_clk));
 sg13g2_buf_8 clkbuf_3_7_0_clk (.A(clknet_0_clk),
    .X(clknet_3_7_0_clk));
 sg13g2_buf_4 clkbuf_6_0__f_clk (.X(clknet_6_0__leaf_clk),
    .A(clknet_3_0_0_clk));
 sg13g2_buf_4 clkbuf_6_1__f_clk (.X(clknet_6_1__leaf_clk),
    .A(clknet_3_0_0_clk));
 sg13g2_buf_4 clkbuf_6_2__f_clk (.X(clknet_6_2__leaf_clk),
    .A(clknet_3_0_0_clk));
 sg13g2_buf_4 clkbuf_6_3__f_clk (.X(clknet_6_3__leaf_clk),
    .A(clknet_3_0_0_clk));
 sg13g2_buf_4 clkbuf_6_4__f_clk (.X(clknet_6_4__leaf_clk),
    .A(clknet_3_0_0_clk));
 sg13g2_buf_4 clkbuf_6_5__f_clk (.X(clknet_6_5__leaf_clk),
    .A(clknet_3_0_0_clk));
 sg13g2_buf_4 clkbuf_6_6__f_clk (.X(clknet_6_6__leaf_clk),
    .A(clknet_3_0_0_clk));
 sg13g2_buf_4 clkbuf_6_7__f_clk (.X(clknet_6_7__leaf_clk),
    .A(clknet_3_0_0_clk));
 sg13g2_buf_4 clkbuf_6_8__f_clk (.X(clknet_6_8__leaf_clk),
    .A(clknet_3_1_0_clk));
 sg13g2_buf_4 clkbuf_6_9__f_clk (.X(clknet_6_9__leaf_clk),
    .A(clknet_3_1_0_clk));
 sg13g2_buf_4 clkbuf_6_10__f_clk (.X(clknet_6_10__leaf_clk),
    .A(clknet_3_1_0_clk));
 sg13g2_buf_4 clkbuf_6_11__f_clk (.X(clknet_6_11__leaf_clk),
    .A(clknet_3_1_0_clk));
 sg13g2_buf_4 clkbuf_6_12__f_clk (.X(clknet_6_12__leaf_clk),
    .A(clknet_3_1_0_clk));
 sg13g2_buf_4 clkbuf_6_13__f_clk (.X(clknet_6_13__leaf_clk),
    .A(clknet_3_1_0_clk));
 sg13g2_buf_4 clkbuf_6_14__f_clk (.X(clknet_6_14__leaf_clk),
    .A(clknet_3_1_0_clk));
 sg13g2_buf_4 clkbuf_6_15__f_clk (.X(clknet_6_15__leaf_clk),
    .A(clknet_3_1_0_clk));
 sg13g2_buf_4 clkbuf_6_16__f_clk (.X(clknet_6_16__leaf_clk),
    .A(clknet_3_2_0_clk));
 sg13g2_buf_4 clkbuf_6_17__f_clk (.X(clknet_6_17__leaf_clk),
    .A(clknet_3_2_0_clk));
 sg13g2_buf_4 clkbuf_6_18__f_clk (.X(clknet_6_18__leaf_clk),
    .A(clknet_3_2_0_clk));
 sg13g2_buf_4 clkbuf_6_19__f_clk (.X(clknet_6_19__leaf_clk),
    .A(clknet_3_2_0_clk));
 sg13g2_buf_4 clkbuf_6_20__f_clk (.X(clknet_6_20__leaf_clk),
    .A(clknet_3_2_0_clk));
 sg13g2_buf_4 clkbuf_6_21__f_clk (.X(clknet_6_21__leaf_clk),
    .A(clknet_3_2_0_clk));
 sg13g2_buf_4 clkbuf_6_22__f_clk (.X(clknet_6_22__leaf_clk),
    .A(clknet_3_2_0_clk));
 sg13g2_buf_4 clkbuf_6_23__f_clk (.X(clknet_6_23__leaf_clk),
    .A(clknet_3_2_0_clk));
 sg13g2_buf_4 clkbuf_6_24__f_clk (.X(clknet_6_24__leaf_clk),
    .A(clknet_3_3_0_clk));
 sg13g2_buf_4 clkbuf_6_25__f_clk (.X(clknet_6_25__leaf_clk),
    .A(clknet_3_3_0_clk));
 sg13g2_buf_4 clkbuf_6_26__f_clk (.X(clknet_6_26__leaf_clk),
    .A(clknet_3_3_0_clk));
 sg13g2_buf_4 clkbuf_6_27__f_clk (.X(clknet_6_27__leaf_clk),
    .A(clknet_3_3_0_clk));
 sg13g2_buf_4 clkbuf_6_28__f_clk (.X(clknet_6_28__leaf_clk),
    .A(clknet_3_3_0_clk));
 sg13g2_buf_4 clkbuf_6_29__f_clk (.X(clknet_6_29__leaf_clk),
    .A(clknet_3_3_0_clk));
 sg13g2_buf_4 clkbuf_6_30__f_clk (.X(clknet_6_30__leaf_clk),
    .A(clknet_3_3_0_clk));
 sg13g2_buf_4 clkbuf_6_31__f_clk (.X(clknet_6_31__leaf_clk),
    .A(clknet_3_3_0_clk));
 sg13g2_buf_4 clkbuf_6_32__f_clk (.X(clknet_6_32__leaf_clk),
    .A(clknet_3_4_0_clk));
 sg13g2_buf_4 clkbuf_6_33__f_clk (.X(clknet_6_33__leaf_clk),
    .A(clknet_3_4_0_clk));
 sg13g2_buf_4 clkbuf_6_34__f_clk (.X(clknet_6_34__leaf_clk),
    .A(clknet_3_4_0_clk));
 sg13g2_buf_4 clkbuf_6_35__f_clk (.X(clknet_6_35__leaf_clk),
    .A(clknet_3_4_0_clk));
 sg13g2_buf_4 clkbuf_6_36__f_clk (.X(clknet_6_36__leaf_clk),
    .A(clknet_3_4_0_clk));
 sg13g2_buf_4 clkbuf_6_37__f_clk (.X(clknet_6_37__leaf_clk),
    .A(clknet_3_4_0_clk));
 sg13g2_buf_4 clkbuf_6_38__f_clk (.X(clknet_6_38__leaf_clk),
    .A(clknet_3_4_0_clk));
 sg13g2_buf_4 clkbuf_6_39__f_clk (.X(clknet_6_39__leaf_clk),
    .A(clknet_3_4_0_clk));
 sg13g2_buf_4 clkbuf_6_40__f_clk (.X(clknet_6_40__leaf_clk),
    .A(clknet_3_5_0_clk));
 sg13g2_buf_4 clkbuf_6_41__f_clk (.X(clknet_6_41__leaf_clk),
    .A(clknet_3_5_0_clk));
 sg13g2_buf_4 clkbuf_6_42__f_clk (.X(clknet_6_42__leaf_clk),
    .A(clknet_3_5_0_clk));
 sg13g2_buf_4 clkbuf_6_43__f_clk (.X(clknet_6_43__leaf_clk),
    .A(clknet_3_5_0_clk));
 sg13g2_buf_4 clkbuf_6_44__f_clk (.X(clknet_6_44__leaf_clk),
    .A(clknet_3_5_0_clk));
 sg13g2_buf_4 clkbuf_6_45__f_clk (.X(clknet_6_45__leaf_clk),
    .A(clknet_3_5_0_clk));
 sg13g2_buf_4 clkbuf_6_46__f_clk (.X(clknet_6_46__leaf_clk),
    .A(clknet_3_5_0_clk));
 sg13g2_buf_4 clkbuf_6_47__f_clk (.X(clknet_6_47__leaf_clk),
    .A(clknet_3_5_0_clk));
 sg13g2_buf_4 clkbuf_6_48__f_clk (.X(clknet_6_48__leaf_clk),
    .A(clknet_3_6_0_clk));
 sg13g2_buf_4 clkbuf_6_49__f_clk (.X(clknet_6_49__leaf_clk),
    .A(clknet_3_6_0_clk));
 sg13g2_buf_4 clkbuf_6_50__f_clk (.X(clknet_6_50__leaf_clk),
    .A(clknet_3_6_0_clk));
 sg13g2_buf_4 clkbuf_6_51__f_clk (.X(clknet_6_51__leaf_clk),
    .A(clknet_3_6_0_clk));
 sg13g2_buf_4 clkbuf_6_52__f_clk (.X(clknet_6_52__leaf_clk),
    .A(clknet_3_6_0_clk));
 sg13g2_buf_4 clkbuf_6_53__f_clk (.X(clknet_6_53__leaf_clk),
    .A(clknet_3_6_0_clk));
 sg13g2_buf_4 clkbuf_6_54__f_clk (.X(clknet_6_54__leaf_clk),
    .A(clknet_3_6_0_clk));
 sg13g2_buf_4 clkbuf_6_55__f_clk (.X(clknet_6_55__leaf_clk),
    .A(clknet_3_6_0_clk));
 sg13g2_buf_4 clkbuf_6_56__f_clk (.X(clknet_6_56__leaf_clk),
    .A(clknet_3_7_0_clk));
 sg13g2_buf_4 clkbuf_6_57__f_clk (.X(clknet_6_57__leaf_clk),
    .A(clknet_3_7_0_clk));
 sg13g2_buf_4 clkbuf_6_58__f_clk (.X(clknet_6_58__leaf_clk),
    .A(clknet_3_7_0_clk));
 sg13g2_buf_4 clkbuf_6_59__f_clk (.X(clknet_6_59__leaf_clk),
    .A(clknet_3_7_0_clk));
 sg13g2_buf_4 clkbuf_6_60__f_clk (.X(clknet_6_60__leaf_clk),
    .A(clknet_3_7_0_clk));
 sg13g2_buf_4 clkbuf_6_61__f_clk (.X(clknet_6_61__leaf_clk),
    .A(clknet_3_7_0_clk));
 sg13g2_buf_4 clkbuf_6_62__f_clk (.X(clknet_6_62__leaf_clk),
    .A(clknet_3_7_0_clk));
 sg13g2_buf_4 clkbuf_6_63__f_clk (.X(clknet_6_63__leaf_clk),
    .A(clknet_3_7_0_clk));
 sg13g2_buf_8 clkload0 (.A(clknet_6_15__leaf_clk));
 sg13g2_buf_8 clkload1 (.A(clknet_6_23__leaf_clk));
 sg13g2_buf_8 clkload2 (.A(clknet_6_31__leaf_clk));
 sg13g2_buf_8 clkload3 (.A(clknet_6_39__leaf_clk));
 sg13g2_buf_8 clkload4 (.A(clknet_6_47__leaf_clk));
 sg13g2_buf_8 clkload5 (.A(clknet_6_55__leaf_clk));
 sg13g2_buf_8 clkload6 (.A(clknet_6_63__leaf_clk));
 sg13g2_inv_4 clkload7 (.A(clknet_leaf_312_clk));
 sg13g2_buf_8 clkload8 (.A(clknet_leaf_115_clk));
 sg13g2_inv_2 clkload9 (.A(clknet_leaf_116_clk));
 sg13g2_inv_2 clkload10 (.A(clknet_leaf_117_clk));
 sg13g2_buf_16 clkload11 (.A(clknet_leaf_173_clk));
 sg13g2_inv_2 clkload12 (.A(clknet_leaf_172_clk));
 sg13g2_antennanp ANTENNA_1 (.A(_00207_));
 sg13g2_antennanp ANTENNA_2 (.A(_00785_));
 sg13g2_antennanp ANTENNA_3 (.A(_00977_));
 sg13g2_antennanp ANTENNA_4 (.A(_01032_));
 sg13g2_antennanp ANTENNA_5 (.A(_01047_));
 sg13g2_antennanp ANTENNA_6 (.A(_01048_));
 sg13g2_antennanp ANTENNA_7 (.A(_02836_));
 sg13g2_antennanp ANTENNA_8 (.A(_02836_));
 sg13g2_antennanp ANTENNA_9 (.A(_02836_));
 sg13g2_antennanp ANTENNA_10 (.A(_02836_));
 sg13g2_antennanp ANTENNA_11 (.A(_02845_));
 sg13g2_antennanp ANTENNA_12 (.A(_02845_));
 sg13g2_antennanp ANTENNA_13 (.A(_02845_));
 sg13g2_antennanp ANTENNA_14 (.A(_02845_));
 sg13g2_antennanp ANTENNA_15 (.A(_02845_));
 sg13g2_antennanp ANTENNA_16 (.A(_02845_));
 sg13g2_antennanp ANTENNA_17 (.A(_02845_));
 sg13g2_antennanp ANTENNA_18 (.A(_02845_));
 sg13g2_antennanp ANTENNA_19 (.A(_02845_));
 sg13g2_antennanp ANTENNA_20 (.A(_02849_));
 sg13g2_antennanp ANTENNA_21 (.A(_02849_));
 sg13g2_antennanp ANTENNA_22 (.A(_02849_));
 sg13g2_antennanp ANTENNA_23 (.A(_02849_));
 sg13g2_antennanp ANTENNA_24 (.A(_02849_));
 sg13g2_antennanp ANTENNA_25 (.A(_02849_));
 sg13g2_antennanp ANTENNA_26 (.A(_02849_));
 sg13g2_antennanp ANTENNA_27 (.A(_02849_));
 sg13g2_antennanp ANTENNA_28 (.A(_02849_));
 sg13g2_antennanp ANTENNA_29 (.A(_02861_));
 sg13g2_antennanp ANTENNA_30 (.A(_02861_));
 sg13g2_antennanp ANTENNA_31 (.A(_02861_));
 sg13g2_antennanp ANTENNA_32 (.A(_02861_));
 sg13g2_antennanp ANTENNA_33 (.A(_02954_));
 sg13g2_antennanp ANTENNA_34 (.A(_02954_));
 sg13g2_antennanp ANTENNA_35 (.A(_02954_));
 sg13g2_antennanp ANTENNA_36 (.A(_02954_));
 sg13g2_antennanp ANTENNA_37 (.A(_02954_));
 sg13g2_antennanp ANTENNA_38 (.A(_02976_));
 sg13g2_antennanp ANTENNA_39 (.A(_02976_));
 sg13g2_antennanp ANTENNA_40 (.A(_02976_));
 sg13g2_antennanp ANTENNA_41 (.A(_02976_));
 sg13g2_antennanp ANTENNA_42 (.A(_02976_));
 sg13g2_antennanp ANTENNA_43 (.A(_02976_));
 sg13g2_antennanp ANTENNA_44 (.A(_02976_));
 sg13g2_antennanp ANTENNA_45 (.A(_02976_));
 sg13g2_antennanp ANTENNA_46 (.A(_02976_));
 sg13g2_antennanp ANTENNA_47 (.A(_03081_));
 sg13g2_antennanp ANTENNA_48 (.A(_03148_));
 sg13g2_antennanp ANTENNA_49 (.A(_03237_));
 sg13g2_antennanp ANTENNA_50 (.A(_03237_));
 sg13g2_antennanp ANTENNA_51 (.A(_03237_));
 sg13g2_antennanp ANTENNA_52 (.A(_03507_));
 sg13g2_antennanp ANTENNA_53 (.A(_03507_));
 sg13g2_antennanp ANTENNA_54 (.A(_03507_));
 sg13g2_antennanp ANTENNA_55 (.A(_03507_));
 sg13g2_antennanp ANTENNA_56 (.A(_03507_));
 sg13g2_antennanp ANTENNA_57 (.A(_03507_));
 sg13g2_antennanp ANTENNA_58 (.A(_03513_));
 sg13g2_antennanp ANTENNA_59 (.A(_03513_));
 sg13g2_antennanp ANTENNA_60 (.A(_03513_));
 sg13g2_antennanp ANTENNA_61 (.A(_03513_));
 sg13g2_antennanp ANTENNA_62 (.A(_03513_));
 sg13g2_antennanp ANTENNA_63 (.A(_03513_));
 sg13g2_antennanp ANTENNA_64 (.A(_03513_));
 sg13g2_antennanp ANTENNA_65 (.A(_03513_));
 sg13g2_antennanp ANTENNA_66 (.A(_03513_));
 sg13g2_antennanp ANTENNA_67 (.A(_03513_));
 sg13g2_antennanp ANTENNA_68 (.A(_03513_));
 sg13g2_antennanp ANTENNA_69 (.A(_03513_));
 sg13g2_antennanp ANTENNA_70 (.A(_03539_));
 sg13g2_antennanp ANTENNA_71 (.A(_03539_));
 sg13g2_antennanp ANTENNA_72 (.A(_03539_));
 sg13g2_antennanp ANTENNA_73 (.A(_03539_));
 sg13g2_antennanp ANTENNA_74 (.A(_03691_));
 sg13g2_antennanp ANTENNA_75 (.A(_03691_));
 sg13g2_antennanp ANTENNA_76 (.A(_03691_));
 sg13g2_antennanp ANTENNA_77 (.A(_03691_));
 sg13g2_antennanp ANTENNA_78 (.A(_03824_));
 sg13g2_antennanp ANTENNA_79 (.A(_03835_));
 sg13g2_antennanp ANTENNA_80 (.A(_03835_));
 sg13g2_antennanp ANTENNA_81 (.A(_03835_));
 sg13g2_antennanp ANTENNA_82 (.A(_03835_));
 sg13g2_antennanp ANTENNA_83 (.A(_03838_));
 sg13g2_antennanp ANTENNA_84 (.A(_03838_));
 sg13g2_antennanp ANTENNA_85 (.A(_03838_));
 sg13g2_antennanp ANTENNA_86 (.A(_03838_));
 sg13g2_antennanp ANTENNA_87 (.A(_03838_));
 sg13g2_antennanp ANTENNA_88 (.A(_03838_));
 sg13g2_antennanp ANTENNA_89 (.A(_03838_));
 sg13g2_antennanp ANTENNA_90 (.A(_03838_));
 sg13g2_antennanp ANTENNA_91 (.A(_03838_));
 sg13g2_antennanp ANTENNA_92 (.A(_03838_));
 sg13g2_antennanp ANTENNA_93 (.A(_04834_));
 sg13g2_antennanp ANTENNA_94 (.A(_04834_));
 sg13g2_antennanp ANTENNA_95 (.A(_04834_));
 sg13g2_antennanp ANTENNA_96 (.A(_04834_));
 sg13g2_antennanp ANTENNA_97 (.A(_04834_));
 sg13g2_antennanp ANTENNA_98 (.A(_04855_));
 sg13g2_antennanp ANTENNA_99 (.A(_04980_));
 sg13g2_antennanp ANTENNA_100 (.A(_04980_));
 sg13g2_antennanp ANTENNA_101 (.A(_04980_));
 sg13g2_antennanp ANTENNA_102 (.A(_04980_));
 sg13g2_antennanp ANTENNA_103 (.A(_04980_));
 sg13g2_antennanp ANTENNA_104 (.A(_05006_));
 sg13g2_antennanp ANTENNA_105 (.A(_05157_));
 sg13g2_antennanp ANTENNA_106 (.A(_05199_));
 sg13g2_antennanp ANTENNA_107 (.A(_05229_));
 sg13g2_antennanp ANTENNA_108 (.A(_05260_));
 sg13g2_antennanp ANTENNA_109 (.A(_05270_));
 sg13g2_antennanp ANTENNA_110 (.A(_05307_));
 sg13g2_antennanp ANTENNA_111 (.A(_05314_));
 sg13g2_antennanp ANTENNA_112 (.A(_05464_));
 sg13g2_antennanp ANTENNA_113 (.A(_05525_));
 sg13g2_antennanp ANTENNA_114 (.A(_05529_));
 sg13g2_antennanp ANTENNA_115 (.A(_05607_));
 sg13g2_antennanp ANTENNA_116 (.A(_05676_));
 sg13g2_antennanp ANTENNA_117 (.A(_05756_));
 sg13g2_antennanp ANTENNA_118 (.A(_05770_));
 sg13g2_antennanp ANTENNA_119 (.A(_05780_));
 sg13g2_antennanp ANTENNA_120 (.A(_05780_));
 sg13g2_antennanp ANTENNA_121 (.A(_05780_));
 sg13g2_antennanp ANTENNA_122 (.A(_05780_));
 sg13g2_antennanp ANTENNA_123 (.A(_05796_));
 sg13g2_antennanp ANTENNA_124 (.A(_06581_));
 sg13g2_antennanp ANTENNA_125 (.A(_06581_));
 sg13g2_antennanp ANTENNA_126 (.A(_06581_));
 sg13g2_antennanp ANTENNA_127 (.A(_06581_));
 sg13g2_antennanp ANTENNA_128 (.A(_06581_));
 sg13g2_antennanp ANTENNA_129 (.A(_06581_));
 sg13g2_antennanp ANTENNA_130 (.A(_06581_));
 sg13g2_antennanp ANTENNA_131 (.A(_06581_));
 sg13g2_antennanp ANTENNA_132 (.A(_06581_));
 sg13g2_antennanp ANTENNA_133 (.A(_06582_));
 sg13g2_antennanp ANTENNA_134 (.A(_06582_));
 sg13g2_antennanp ANTENNA_135 (.A(_06582_));
 sg13g2_antennanp ANTENNA_136 (.A(_06582_));
 sg13g2_antennanp ANTENNA_137 (.A(_06885_));
 sg13g2_antennanp ANTENNA_138 (.A(_06885_));
 sg13g2_antennanp ANTENNA_139 (.A(_06885_));
 sg13g2_antennanp ANTENNA_140 (.A(_06885_));
 sg13g2_antennanp ANTENNA_141 (.A(_07626_));
 sg13g2_antennanp ANTENNA_142 (.A(_07632_));
 sg13g2_antennanp ANTENNA_143 (.A(_07634_));
 sg13g2_antennanp ANTENNA_144 (.A(_07851_));
 sg13g2_antennanp ANTENNA_145 (.A(_07851_));
 sg13g2_antennanp ANTENNA_146 (.A(_07851_));
 sg13g2_antennanp ANTENNA_147 (.A(_07851_));
 sg13g2_antennanp ANTENNA_148 (.A(_07851_));
 sg13g2_antennanp ANTENNA_149 (.A(_07851_));
 sg13g2_antennanp ANTENNA_150 (.A(_07851_));
 sg13g2_antennanp ANTENNA_151 (.A(_07851_));
 sg13g2_antennanp ANTENNA_152 (.A(_07851_));
 sg13g2_antennanp ANTENNA_153 (.A(_07851_));
 sg13g2_antennanp ANTENNA_154 (.A(_08260_));
 sg13g2_antennanp ANTENNA_155 (.A(_08260_));
 sg13g2_antennanp ANTENNA_156 (.A(_08346_));
 sg13g2_antennanp ANTENNA_157 (.A(_08346_));
 sg13g2_antennanp ANTENNA_158 (.A(_08346_));
 sg13g2_antennanp ANTENNA_159 (.A(_08346_));
 sg13g2_antennanp ANTENNA_160 (.A(_08346_));
 sg13g2_antennanp ANTENNA_161 (.A(_08346_));
 sg13g2_antennanp ANTENNA_162 (.A(_08346_));
 sg13g2_antennanp ANTENNA_163 (.A(_08346_));
 sg13g2_antennanp ANTENNA_164 (.A(_08455_));
 sg13g2_antennanp ANTENNA_165 (.A(_08455_));
 sg13g2_antennanp ANTENNA_166 (.A(_08455_));
 sg13g2_antennanp ANTENNA_167 (.A(_08455_));
 sg13g2_antennanp ANTENNA_168 (.A(_08497_));
 sg13g2_antennanp ANTENNA_169 (.A(_08497_));
 sg13g2_antennanp ANTENNA_170 (.A(_08497_));
 sg13g2_antennanp ANTENNA_171 (.A(_08565_));
 sg13g2_antennanp ANTENNA_172 (.A(_08565_));
 sg13g2_antennanp ANTENNA_173 (.A(_08565_));
 sg13g2_antennanp ANTENNA_174 (.A(_08603_));
 sg13g2_antennanp ANTENNA_175 (.A(_08603_));
 sg13g2_antennanp ANTENNA_176 (.A(_08603_));
 sg13g2_antennanp ANTENNA_177 (.A(_08633_));
 sg13g2_antennanp ANTENNA_178 (.A(_08663_));
 sg13g2_antennanp ANTENNA_179 (.A(_08663_));
 sg13g2_antennanp ANTENNA_180 (.A(_08663_));
 sg13g2_antennanp ANTENNA_181 (.A(_08663_));
 sg13g2_antennanp ANTENNA_182 (.A(_08663_));
 sg13g2_antennanp ANTENNA_183 (.A(_08663_));
 sg13g2_antennanp ANTENNA_184 (.A(_08776_));
 sg13g2_antennanp ANTENNA_185 (.A(_08777_));
 sg13g2_antennanp ANTENNA_186 (.A(_08799_));
 sg13g2_antennanp ANTENNA_187 (.A(_08799_));
 sg13g2_antennanp ANTENNA_188 (.A(_08799_));
 sg13g2_antennanp ANTENNA_189 (.A(_08799_));
 sg13g2_antennanp ANTENNA_190 (.A(_08799_));
 sg13g2_antennanp ANTENNA_191 (.A(_08799_));
 sg13g2_antennanp ANTENNA_192 (.A(_08820_));
 sg13g2_antennanp ANTENNA_193 (.A(_08820_));
 sg13g2_antennanp ANTENNA_194 (.A(_08820_));
 sg13g2_antennanp ANTENNA_195 (.A(_08820_));
 sg13g2_antennanp ANTENNA_196 (.A(_08820_));
 sg13g2_antennanp ANTENNA_197 (.A(_08820_));
 sg13g2_antennanp ANTENNA_198 (.A(_08826_));
 sg13g2_antennanp ANTENNA_199 (.A(_08826_));
 sg13g2_antennanp ANTENNA_200 (.A(_08826_));
 sg13g2_antennanp ANTENNA_201 (.A(_08826_));
 sg13g2_antennanp ANTENNA_202 (.A(_08826_));
 sg13g2_antennanp ANTENNA_203 (.A(_08826_));
 sg13g2_antennanp ANTENNA_204 (.A(_08848_));
 sg13g2_antennanp ANTENNA_205 (.A(_08848_));
 sg13g2_antennanp ANTENNA_206 (.A(_08848_));
 sg13g2_antennanp ANTENNA_207 (.A(_08868_));
 sg13g2_antennanp ANTENNA_208 (.A(_08900_));
 sg13g2_antennanp ANTENNA_209 (.A(_08900_));
 sg13g2_antennanp ANTENNA_210 (.A(_08900_));
 sg13g2_antennanp ANTENNA_211 (.A(_08950_));
 sg13g2_antennanp ANTENNA_212 (.A(_08950_));
 sg13g2_antennanp ANTENNA_213 (.A(_08950_));
 sg13g2_antennanp ANTENNA_214 (.A(_08950_));
 sg13g2_antennanp ANTENNA_215 (.A(_08950_));
 sg13g2_antennanp ANTENNA_216 (.A(_08950_));
 sg13g2_antennanp ANTENNA_217 (.A(_08970_));
 sg13g2_antennanp ANTENNA_218 (.A(_08970_));
 sg13g2_antennanp ANTENNA_219 (.A(_08986_));
 sg13g2_antennanp ANTENNA_220 (.A(_08986_));
 sg13g2_antennanp ANTENNA_221 (.A(_09002_));
 sg13g2_antennanp ANTENNA_222 (.A(_09002_));
 sg13g2_antennanp ANTENNA_223 (.A(_09065_));
 sg13g2_antennanp ANTENNA_224 (.A(_09065_));
 sg13g2_antennanp ANTENNA_225 (.A(_09091_));
 sg13g2_antennanp ANTENNA_226 (.A(_09091_));
 sg13g2_antennanp ANTENNA_227 (.A(_09091_));
 sg13g2_antennanp ANTENNA_228 (.A(_09091_));
 sg13g2_antennanp ANTENNA_229 (.A(_09091_));
 sg13g2_antennanp ANTENNA_230 (.A(_09091_));
 sg13g2_antennanp ANTENNA_231 (.A(_09091_));
 sg13g2_antennanp ANTENNA_232 (.A(_09091_));
 sg13g2_antennanp ANTENNA_233 (.A(_09091_));
 sg13g2_antennanp ANTENNA_234 (.A(_09091_));
 sg13g2_antennanp ANTENNA_235 (.A(_09099_));
 sg13g2_antennanp ANTENNA_236 (.A(_09120_));
 sg13g2_antennanp ANTENNA_237 (.A(_09120_));
 sg13g2_antennanp ANTENNA_238 (.A(_09156_));
 sg13g2_antennanp ANTENNA_239 (.A(_09156_));
 sg13g2_antennanp ANTENNA_240 (.A(_09156_));
 sg13g2_antennanp ANTENNA_241 (.A(_09156_));
 sg13g2_antennanp ANTENNA_242 (.A(_09156_));
 sg13g2_antennanp ANTENNA_243 (.A(_09156_));
 sg13g2_antennanp ANTENNA_244 (.A(_09158_));
 sg13g2_antennanp ANTENNA_245 (.A(_09158_));
 sg13g2_antennanp ANTENNA_246 (.A(_09158_));
 sg13g2_antennanp ANTENNA_247 (.A(_09173_));
 sg13g2_antennanp ANTENNA_248 (.A(_09211_));
 sg13g2_antennanp ANTENNA_249 (.A(_09211_));
 sg13g2_antennanp ANTENNA_250 (.A(_09211_));
 sg13g2_antennanp ANTENNA_251 (.A(_09211_));
 sg13g2_antennanp ANTENNA_252 (.A(_09211_));
 sg13g2_antennanp ANTENNA_253 (.A(_09218_));
 sg13g2_antennanp ANTENNA_254 (.A(_09223_));
 sg13g2_antennanp ANTENNA_255 (.A(_09223_));
 sg13g2_antennanp ANTENNA_256 (.A(_09223_));
 sg13g2_antennanp ANTENNA_257 (.A(_09223_));
 sg13g2_antennanp ANTENNA_258 (.A(_09223_));
 sg13g2_antennanp ANTENNA_259 (.A(_09223_));
 sg13g2_antennanp ANTENNA_260 (.A(_09223_));
 sg13g2_antennanp ANTENNA_261 (.A(_09223_));
 sg13g2_antennanp ANTENNA_262 (.A(_09240_));
 sg13g2_antennanp ANTENNA_263 (.A(_09240_));
 sg13g2_antennanp ANTENNA_264 (.A(_09240_));
 sg13g2_antennanp ANTENNA_265 (.A(_09240_));
 sg13g2_antennanp ANTENNA_266 (.A(_09240_));
 sg13g2_antennanp ANTENNA_267 (.A(_09240_));
 sg13g2_antennanp ANTENNA_268 (.A(_09240_));
 sg13g2_antennanp ANTENNA_269 (.A(_09240_));
 sg13g2_antennanp ANTENNA_270 (.A(_09298_));
 sg13g2_antennanp ANTENNA_271 (.A(_09298_));
 sg13g2_antennanp ANTENNA_272 (.A(_09298_));
 sg13g2_antennanp ANTENNA_273 (.A(_09298_));
 sg13g2_antennanp ANTENNA_274 (.A(_09298_));
 sg13g2_antennanp ANTENNA_275 (.A(_09298_));
 sg13g2_antennanp ANTENNA_276 (.A(_09298_));
 sg13g2_antennanp ANTENNA_277 (.A(_09298_));
 sg13g2_antennanp ANTENNA_278 (.A(_09298_));
 sg13g2_antennanp ANTENNA_279 (.A(_09298_));
 sg13g2_antennanp ANTENNA_280 (.A(_09316_));
 sg13g2_antennanp ANTENNA_281 (.A(_09316_));
 sg13g2_antennanp ANTENNA_282 (.A(_09316_));
 sg13g2_antennanp ANTENNA_283 (.A(_09316_));
 sg13g2_antennanp ANTENNA_284 (.A(_09316_));
 sg13g2_antennanp ANTENNA_285 (.A(_09316_));
 sg13g2_antennanp ANTENNA_286 (.A(_09316_));
 sg13g2_antennanp ANTENNA_287 (.A(_09316_));
 sg13g2_antennanp ANTENNA_288 (.A(_09316_));
 sg13g2_antennanp ANTENNA_289 (.A(_09316_));
 sg13g2_antennanp ANTENNA_290 (.A(_09316_));
 sg13g2_antennanp ANTENNA_291 (.A(_09316_));
 sg13g2_antennanp ANTENNA_292 (.A(_09316_));
 sg13g2_antennanp ANTENNA_293 (.A(_09316_));
 sg13g2_antennanp ANTENNA_294 (.A(_09316_));
 sg13g2_antennanp ANTENNA_295 (.A(_09316_));
 sg13g2_antennanp ANTENNA_296 (.A(_09316_));
 sg13g2_antennanp ANTENNA_297 (.A(_09316_));
 sg13g2_antennanp ANTENNA_298 (.A(_09316_));
 sg13g2_antennanp ANTENNA_299 (.A(_09316_));
 sg13g2_antennanp ANTENNA_300 (.A(_09316_));
 sg13g2_antennanp ANTENNA_301 (.A(_09316_));
 sg13g2_antennanp ANTENNA_302 (.A(_09316_));
 sg13g2_antennanp ANTENNA_303 (.A(_09316_));
 sg13g2_antennanp ANTENNA_304 (.A(_09317_));
 sg13g2_antennanp ANTENNA_305 (.A(_09317_));
 sg13g2_antennanp ANTENNA_306 (.A(_09317_));
 sg13g2_antennanp ANTENNA_307 (.A(_09317_));
 sg13g2_antennanp ANTENNA_308 (.A(_09318_));
 sg13g2_antennanp ANTENNA_309 (.A(_09318_));
 sg13g2_antennanp ANTENNA_310 (.A(_09318_));
 sg13g2_antennanp ANTENNA_311 (.A(_09323_));
 sg13g2_antennanp ANTENNA_312 (.A(_09323_));
 sg13g2_antennanp ANTENNA_313 (.A(_09323_));
 sg13g2_antennanp ANTENNA_314 (.A(_09323_));
 sg13g2_antennanp ANTENNA_315 (.A(_09323_));
 sg13g2_antennanp ANTENNA_316 (.A(_09394_));
 sg13g2_antennanp ANTENNA_317 (.A(_09396_));
 sg13g2_antennanp ANTENNA_318 (.A(_09447_));
 sg13g2_antennanp ANTENNA_319 (.A(_09448_));
 sg13g2_antennanp ANTENNA_320 (.A(_09448_));
 sg13g2_antennanp ANTENNA_321 (.A(_09448_));
 sg13g2_antennanp ANTENNA_322 (.A(_09448_));
 sg13g2_antennanp ANTENNA_323 (.A(_09450_));
 sg13g2_antennanp ANTENNA_324 (.A(_09450_));
 sg13g2_antennanp ANTENNA_325 (.A(_09492_));
 sg13g2_antennanp ANTENNA_326 (.A(_09521_));
 sg13g2_antennanp ANTENNA_327 (.A(_09544_));
 sg13g2_antennanp ANTENNA_328 (.A(_09604_));
 sg13g2_antennanp ANTENNA_329 (.A(_09604_));
 sg13g2_antennanp ANTENNA_330 (.A(_09604_));
 sg13g2_antennanp ANTENNA_331 (.A(_09657_));
 sg13g2_antennanp ANTENNA_332 (.A(_09678_));
 sg13g2_antennanp ANTENNA_333 (.A(_09722_));
 sg13g2_antennanp ANTENNA_334 (.A(_09769_));
 sg13g2_antennanp ANTENNA_335 (.A(_09791_));
 sg13g2_antennanp ANTENNA_336 (.A(_09852_));
 sg13g2_antennanp ANTENNA_337 (.A(_09852_));
 sg13g2_antennanp ANTENNA_338 (.A(_09852_));
 sg13g2_antennanp ANTENNA_339 (.A(_09852_));
 sg13g2_antennanp ANTENNA_340 (.A(_09852_));
 sg13g2_antennanp ANTENNA_341 (.A(_09852_));
 sg13g2_antennanp ANTENNA_342 (.A(_09852_));
 sg13g2_antennanp ANTENNA_343 (.A(_09852_));
 sg13g2_antennanp ANTENNA_344 (.A(_09852_));
 sg13g2_antennanp ANTENNA_345 (.A(_10042_));
 sg13g2_antennanp ANTENNA_346 (.A(_10042_));
 sg13g2_antennanp ANTENNA_347 (.A(_10042_));
 sg13g2_antennanp ANTENNA_348 (.A(_10042_));
 sg13g2_antennanp ANTENNA_349 (.A(_10107_));
 sg13g2_antennanp ANTENNA_350 (.A(_10107_));
 sg13g2_antennanp ANTENNA_351 (.A(_10107_));
 sg13g2_antennanp ANTENNA_352 (.A(_10107_));
 sg13g2_antennanp ANTENNA_353 (.A(_10107_));
 sg13g2_antennanp ANTENNA_354 (.A(_10121_));
 sg13g2_antennanp ANTENNA_355 (.A(_10121_));
 sg13g2_antennanp ANTENNA_356 (.A(_10121_));
 sg13g2_antennanp ANTENNA_357 (.A(_10121_));
 sg13g2_antennanp ANTENNA_358 (.A(_10146_));
 sg13g2_antennanp ANTENNA_359 (.A(_10146_));
 sg13g2_antennanp ANTENNA_360 (.A(_10146_));
 sg13g2_antennanp ANTENNA_361 (.A(_10146_));
 sg13g2_antennanp ANTENNA_362 (.A(_10146_));
 sg13g2_antennanp ANTENNA_363 (.A(_10146_));
 sg13g2_antennanp ANTENNA_364 (.A(_10146_));
 sg13g2_antennanp ANTENNA_365 (.A(_10146_));
 sg13g2_antennanp ANTENNA_366 (.A(_10162_));
 sg13g2_antennanp ANTENNA_367 (.A(_10162_));
 sg13g2_antennanp ANTENNA_368 (.A(_10162_));
 sg13g2_antennanp ANTENNA_369 (.A(_10162_));
 sg13g2_antennanp ANTENNA_370 (.A(_10162_));
 sg13g2_antennanp ANTENNA_371 (.A(_10162_));
 sg13g2_antennanp ANTENNA_372 (.A(_10162_));
 sg13g2_antennanp ANTENNA_373 (.A(_10162_));
 sg13g2_antennanp ANTENNA_374 (.A(_10162_));
 sg13g2_antennanp ANTENNA_375 (.A(_10162_));
 sg13g2_antennanp ANTENNA_376 (.A(_10162_));
 sg13g2_antennanp ANTENNA_377 (.A(_10162_));
 sg13g2_antennanp ANTENNA_378 (.A(_10162_));
 sg13g2_antennanp ANTENNA_379 (.A(_10379_));
 sg13g2_antennanp ANTENNA_380 (.A(_10379_));
 sg13g2_antennanp ANTENNA_381 (.A(_10379_));
 sg13g2_antennanp ANTENNA_382 (.A(_10642_));
 sg13g2_antennanp ANTENNA_383 (.A(_10642_));
 sg13g2_antennanp ANTENNA_384 (.A(_10642_));
 sg13g2_antennanp ANTENNA_385 (.A(_10642_));
 sg13g2_antennanp ANTENNA_386 (.A(_10642_));
 sg13g2_antennanp ANTENNA_387 (.A(_10642_));
 sg13g2_antennanp ANTENNA_388 (.A(_10642_));
 sg13g2_antennanp ANTENNA_389 (.A(_10744_));
 sg13g2_antennanp ANTENNA_390 (.A(_10744_));
 sg13g2_antennanp ANTENNA_391 (.A(_10744_));
 sg13g2_antennanp ANTENNA_392 (.A(_10744_));
 sg13g2_antennanp ANTENNA_393 (.A(_12205_));
 sg13g2_antennanp ANTENNA_394 (.A(_12205_));
 sg13g2_antennanp ANTENNA_395 (.A(_12205_));
 sg13g2_antennanp ANTENNA_396 (.A(_12205_));
 sg13g2_antennanp ANTENNA_397 (.A(_12205_));
 sg13g2_antennanp ANTENNA_398 (.A(_12205_));
 sg13g2_antennanp ANTENNA_399 (.A(_12205_));
 sg13g2_antennanp ANTENNA_400 (.A(_12205_));
 sg13g2_antennanp ANTENNA_401 (.A(_12205_));
 sg13g2_antennanp ANTENNA_402 (.A(_12218_));
 sg13g2_antennanp ANTENNA_403 (.A(_12218_));
 sg13g2_antennanp ANTENNA_404 (.A(_12218_));
 sg13g2_antennanp ANTENNA_405 (.A(_12218_));
 sg13g2_antennanp ANTENNA_406 (.A(_12218_));
 sg13g2_antennanp ANTENNA_407 (.A(_12218_));
 sg13g2_antennanp ANTENNA_408 (.A(_12218_));
 sg13g2_antennanp ANTENNA_409 (.A(_12218_));
 sg13g2_antennanp ANTENNA_410 (.A(_12218_));
 sg13g2_antennanp ANTENNA_411 (.A(_12218_));
 sg13g2_antennanp ANTENNA_412 (.A(_12218_));
 sg13g2_antennanp ANTENNA_413 (.A(_12218_));
 sg13g2_antennanp ANTENNA_414 (.A(_12218_));
 sg13g2_antennanp ANTENNA_415 (.A(_12218_));
 sg13g2_antennanp ANTENNA_416 (.A(_12218_));
 sg13g2_antennanp ANTENNA_417 (.A(_12218_));
 sg13g2_antennanp ANTENNA_418 (.A(_12218_));
 sg13g2_antennanp ANTENNA_419 (.A(_12218_));
 sg13g2_antennanp ANTENNA_420 (.A(_12225_));
 sg13g2_antennanp ANTENNA_421 (.A(_12225_));
 sg13g2_antennanp ANTENNA_422 (.A(_12225_));
 sg13g2_antennanp ANTENNA_423 (.A(_12225_));
 sg13g2_antennanp ANTENNA_424 (.A(_12225_));
 sg13g2_antennanp ANTENNA_425 (.A(_12225_));
 sg13g2_antennanp ANTENNA_426 (.A(_12225_));
 sg13g2_antennanp ANTENNA_427 (.A(_12225_));
 sg13g2_antennanp ANTENNA_428 (.A(_12225_));
 sg13g2_antennanp ANTENNA_429 (.A(_12236_));
 sg13g2_antennanp ANTENNA_430 (.A(_12236_));
 sg13g2_antennanp ANTENNA_431 (.A(_12236_));
 sg13g2_antennanp ANTENNA_432 (.A(_12236_));
 sg13g2_antennanp ANTENNA_433 (.A(_12236_));
 sg13g2_antennanp ANTENNA_434 (.A(_12236_));
 sg13g2_antennanp ANTENNA_435 (.A(_12236_));
 sg13g2_antennanp ANTENNA_436 (.A(_12236_));
 sg13g2_antennanp ANTENNA_437 (.A(_12236_));
 sg13g2_antennanp ANTENNA_438 (.A(clk));
 sg13g2_antennanp ANTENNA_439 (.A(clk));
 sg13g2_antennanp ANTENNA_440 (.A(\cpu.dcache.wdata[10] ));
 sg13g2_antennanp ANTENNA_441 (.A(\cpu.dcache.wdata[10] ));
 sg13g2_antennanp ANTENNA_442 (.A(\cpu.dcache.wdata[10] ));
 sg13g2_antennanp ANTENNA_443 (.A(\cpu.dcache.wdata[10] ));
 sg13g2_antennanp ANTENNA_444 (.A(\cpu.dcache.wdata[12] ));
 sg13g2_antennanp ANTENNA_445 (.A(\cpu.dcache.wdata[12] ));
 sg13g2_antennanp ANTENNA_446 (.A(\cpu.dcache.wdata[12] ));
 sg13g2_antennanp ANTENNA_447 (.A(\cpu.dcache.wdata[12] ));
 sg13g2_antennanp ANTENNA_448 (.A(\cpu.dcache.wdata[15] ));
 sg13g2_antennanp ANTENNA_449 (.A(\cpu.dcache.wdata[15] ));
 sg13g2_antennanp ANTENNA_450 (.A(\cpu.dcache.wdata[15] ));
 sg13g2_antennanp ANTENNA_451 (.A(\cpu.dcache.wdata[15] ));
 sg13g2_antennanp ANTENNA_452 (.A(\cpu.dcache.wdata[9] ));
 sg13g2_antennanp ANTENNA_453 (.A(\cpu.dcache.wdata[9] ));
 sg13g2_antennanp ANTENNA_454 (.A(\cpu.dcache.wdata[9] ));
 sg13g2_antennanp ANTENNA_455 (.A(\cpu.dcache.wdata[9] ));
 sg13g2_antennanp ANTENNA_456 (.A(\cpu.ex.pc[1] ));
 sg13g2_antennanp ANTENNA_457 (.A(\cpu.ex.pc[2] ));
 sg13g2_antennanp ANTENNA_458 (.A(\cpu.gpio.uart_rx ));
 sg13g2_antennanp ANTENNA_459 (.A(\cpu.gpio.uart_rx ));
 sg13g2_antennanp ANTENNA_460 (.A(\cpu.qspi.c_wstrobe_i ));
 sg13g2_antennanp ANTENNA_461 (.A(\cpu.qspi.c_wstrobe_i ));
 sg13g2_antennanp ANTENNA_462 (.A(net3));
 sg13g2_antennanp ANTENNA_463 (.A(net3));
 sg13g2_antennanp ANTENNA_464 (.A(net3));
 sg13g2_antennanp ANTENNA_465 (.A(net11));
 sg13g2_antennanp ANTENNA_466 (.A(net11));
 sg13g2_antennanp ANTENNA_467 (.A(net11));
 sg13g2_antennanp ANTENNA_468 (.A(net12));
 sg13g2_antennanp ANTENNA_469 (.A(net12));
 sg13g2_antennanp ANTENNA_470 (.A(net12));
 sg13g2_antennanp ANTENNA_471 (.A(net13));
 sg13g2_antennanp ANTENNA_472 (.A(net13));
 sg13g2_antennanp ANTENNA_473 (.A(net13));
 sg13g2_antennanp ANTENNA_474 (.A(net14));
 sg13g2_antennanp ANTENNA_475 (.A(net14));
 sg13g2_antennanp ANTENNA_476 (.A(net14));
 sg13g2_antennanp ANTENNA_477 (.A(net36));
 sg13g2_antennanp ANTENNA_478 (.A(net36));
 sg13g2_antennanp ANTENNA_479 (.A(net36));
 sg13g2_antennanp ANTENNA_480 (.A(net36));
 sg13g2_antennanp ANTENNA_481 (.A(net36));
 sg13g2_antennanp ANTENNA_482 (.A(net36));
 sg13g2_antennanp ANTENNA_483 (.A(net36));
 sg13g2_antennanp ANTENNA_484 (.A(net36));
 sg13g2_antennanp ANTENNA_485 (.A(net36));
 sg13g2_antennanp ANTENNA_486 (.A(net36));
 sg13g2_antennanp ANTENNA_487 (.A(net36));
 sg13g2_antennanp ANTENNA_488 (.A(net36));
 sg13g2_antennanp ANTENNA_489 (.A(net36));
 sg13g2_antennanp ANTENNA_490 (.A(net36));
 sg13g2_antennanp ANTENNA_491 (.A(net36));
 sg13g2_antennanp ANTENNA_492 (.A(net36));
 sg13g2_antennanp ANTENNA_493 (.A(net36));
 sg13g2_antennanp ANTENNA_494 (.A(net36));
 sg13g2_antennanp ANTENNA_495 (.A(net36));
 sg13g2_antennanp ANTENNA_496 (.A(net36));
 sg13g2_antennanp ANTENNA_497 (.A(net36));
 sg13g2_antennanp ANTENNA_498 (.A(net36));
 sg13g2_antennanp ANTENNA_499 (.A(net36));
 sg13g2_antennanp ANTENNA_500 (.A(net114));
 sg13g2_antennanp ANTENNA_501 (.A(net114));
 sg13g2_antennanp ANTENNA_502 (.A(net114));
 sg13g2_antennanp ANTENNA_503 (.A(net114));
 sg13g2_antennanp ANTENNA_504 (.A(net114));
 sg13g2_antennanp ANTENNA_505 (.A(net114));
 sg13g2_antennanp ANTENNA_506 (.A(net114));
 sg13g2_antennanp ANTENNA_507 (.A(net114));
 sg13g2_antennanp ANTENNA_508 (.A(net114));
 sg13g2_antennanp ANTENNA_509 (.A(net114));
 sg13g2_antennanp ANTENNA_510 (.A(net114));
 sg13g2_antennanp ANTENNA_511 (.A(net114));
 sg13g2_antennanp ANTENNA_512 (.A(net114));
 sg13g2_antennanp ANTENNA_513 (.A(net114));
 sg13g2_antennanp ANTENNA_514 (.A(net114));
 sg13g2_antennanp ANTENNA_515 (.A(net114));
 sg13g2_antennanp ANTENNA_516 (.A(net452));
 sg13g2_antennanp ANTENNA_517 (.A(net452));
 sg13g2_antennanp ANTENNA_518 (.A(net452));
 sg13g2_antennanp ANTENNA_519 (.A(net452));
 sg13g2_antennanp ANTENNA_520 (.A(net452));
 sg13g2_antennanp ANTENNA_521 (.A(net452));
 sg13g2_antennanp ANTENNA_522 (.A(net452));
 sg13g2_antennanp ANTENNA_523 (.A(net452));
 sg13g2_antennanp ANTENNA_524 (.A(net489));
 sg13g2_antennanp ANTENNA_525 (.A(net489));
 sg13g2_antennanp ANTENNA_526 (.A(net489));
 sg13g2_antennanp ANTENNA_527 (.A(net489));
 sg13g2_antennanp ANTENNA_528 (.A(net489));
 sg13g2_antennanp ANTENNA_529 (.A(net489));
 sg13g2_antennanp ANTENNA_530 (.A(net489));
 sg13g2_antennanp ANTENNA_531 (.A(net489));
 sg13g2_antennanp ANTENNA_532 (.A(net489));
 sg13g2_antennanp ANTENNA_533 (.A(net550));
 sg13g2_antennanp ANTENNA_534 (.A(net550));
 sg13g2_antennanp ANTENNA_535 (.A(net550));
 sg13g2_antennanp ANTENNA_536 (.A(net550));
 sg13g2_antennanp ANTENNA_537 (.A(net550));
 sg13g2_antennanp ANTENNA_538 (.A(net550));
 sg13g2_antennanp ANTENNA_539 (.A(net550));
 sg13g2_antennanp ANTENNA_540 (.A(net550));
 sg13g2_antennanp ANTENNA_541 (.A(net550));
 sg13g2_antennanp ANTENNA_542 (.A(net550));
 sg13g2_antennanp ANTENNA_543 (.A(net550));
 sg13g2_antennanp ANTENNA_544 (.A(net550));
 sg13g2_antennanp ANTENNA_545 (.A(net550));
 sg13g2_antennanp ANTENNA_546 (.A(net550));
 sg13g2_antennanp ANTENNA_547 (.A(net605));
 sg13g2_antennanp ANTENNA_548 (.A(net605));
 sg13g2_antennanp ANTENNA_549 (.A(net605));
 sg13g2_antennanp ANTENNA_550 (.A(net605));
 sg13g2_antennanp ANTENNA_551 (.A(net605));
 sg13g2_antennanp ANTENNA_552 (.A(net605));
 sg13g2_antennanp ANTENNA_553 (.A(net605));
 sg13g2_antennanp ANTENNA_554 (.A(net605));
 sg13g2_antennanp ANTENNA_555 (.A(net605));
 sg13g2_antennanp ANTENNA_556 (.A(net605));
 sg13g2_antennanp ANTENNA_557 (.A(net605));
 sg13g2_antennanp ANTENNA_558 (.A(net605));
 sg13g2_antennanp ANTENNA_559 (.A(net605));
 sg13g2_antennanp ANTENNA_560 (.A(net605));
 sg13g2_antennanp ANTENNA_561 (.A(net605));
 sg13g2_antennanp ANTENNA_562 (.A(net668));
 sg13g2_antennanp ANTENNA_563 (.A(net668));
 sg13g2_antennanp ANTENNA_564 (.A(net668));
 sg13g2_antennanp ANTENNA_565 (.A(net668));
 sg13g2_antennanp ANTENNA_566 (.A(net668));
 sg13g2_antennanp ANTENNA_567 (.A(net668));
 sg13g2_antennanp ANTENNA_568 (.A(net668));
 sg13g2_antennanp ANTENNA_569 (.A(net668));
 sg13g2_antennanp ANTENNA_570 (.A(net668));
 sg13g2_antennanp ANTENNA_571 (.A(net668));
 sg13g2_antennanp ANTENNA_572 (.A(net668));
 sg13g2_antennanp ANTENNA_573 (.A(net668));
 sg13g2_antennanp ANTENNA_574 (.A(net668));
 sg13g2_antennanp ANTENNA_575 (.A(net668));
 sg13g2_antennanp ANTENNA_576 (.A(net668));
 sg13g2_antennanp ANTENNA_577 (.A(net668));
 sg13g2_antennanp ANTENNA_578 (.A(net668));
 sg13g2_antennanp ANTENNA_579 (.A(net668));
 sg13g2_antennanp ANTENNA_580 (.A(net668));
 sg13g2_antennanp ANTENNA_581 (.A(net668));
 sg13g2_antennanp ANTENNA_582 (.A(net686));
 sg13g2_antennanp ANTENNA_583 (.A(net686));
 sg13g2_antennanp ANTENNA_584 (.A(net686));
 sg13g2_antennanp ANTENNA_585 (.A(net686));
 sg13g2_antennanp ANTENNA_586 (.A(net686));
 sg13g2_antennanp ANTENNA_587 (.A(net686));
 sg13g2_antennanp ANTENNA_588 (.A(net686));
 sg13g2_antennanp ANTENNA_589 (.A(net686));
 sg13g2_antennanp ANTENNA_590 (.A(net708));
 sg13g2_antennanp ANTENNA_591 (.A(net708));
 sg13g2_antennanp ANTENNA_592 (.A(net708));
 sg13g2_antennanp ANTENNA_593 (.A(net708));
 sg13g2_antennanp ANTENNA_594 (.A(net708));
 sg13g2_antennanp ANTENNA_595 (.A(net708));
 sg13g2_antennanp ANTENNA_596 (.A(net708));
 sg13g2_antennanp ANTENNA_597 (.A(net708));
 sg13g2_antennanp ANTENNA_598 (.A(net745));
 sg13g2_antennanp ANTENNA_599 (.A(net745));
 sg13g2_antennanp ANTENNA_600 (.A(net745));
 sg13g2_antennanp ANTENNA_601 (.A(net745));
 sg13g2_antennanp ANTENNA_602 (.A(net745));
 sg13g2_antennanp ANTENNA_603 (.A(net745));
 sg13g2_antennanp ANTENNA_604 (.A(net745));
 sg13g2_antennanp ANTENNA_605 (.A(net745));
 sg13g2_antennanp ANTENNA_606 (.A(net745));
 sg13g2_antennanp ANTENNA_607 (.A(net745));
 sg13g2_antennanp ANTENNA_608 (.A(net745));
 sg13g2_antennanp ANTENNA_609 (.A(net745));
 sg13g2_antennanp ANTENNA_610 (.A(net745));
 sg13g2_antennanp ANTENNA_611 (.A(net745));
 sg13g2_antennanp ANTENNA_612 (.A(net745));
 sg13g2_antennanp ANTENNA_613 (.A(net745));
 sg13g2_antennanp ANTENNA_614 (.A(net803));
 sg13g2_antennanp ANTENNA_615 (.A(net803));
 sg13g2_antennanp ANTENNA_616 (.A(net803));
 sg13g2_antennanp ANTENNA_617 (.A(net803));
 sg13g2_antennanp ANTENNA_618 (.A(net803));
 sg13g2_antennanp ANTENNA_619 (.A(net803));
 sg13g2_antennanp ANTENNA_620 (.A(net803));
 sg13g2_antennanp ANTENNA_621 (.A(net803));
 sg13g2_antennanp ANTENNA_622 (.A(net803));
 sg13g2_antennanp ANTENNA_623 (.A(net803));
 sg13g2_antennanp ANTENNA_624 (.A(net803));
 sg13g2_antennanp ANTENNA_625 (.A(net803));
 sg13g2_antennanp ANTENNA_626 (.A(net803));
 sg13g2_antennanp ANTENNA_627 (.A(net803));
 sg13g2_antennanp ANTENNA_628 (.A(net803));
 sg13g2_antennanp ANTENNA_629 (.A(net803));
 sg13g2_antennanp ANTENNA_630 (.A(net858));
 sg13g2_antennanp ANTENNA_631 (.A(net858));
 sg13g2_antennanp ANTENNA_632 (.A(net858));
 sg13g2_antennanp ANTENNA_633 (.A(net858));
 sg13g2_antennanp ANTENNA_634 (.A(net858));
 sg13g2_antennanp ANTENNA_635 (.A(net858));
 sg13g2_antennanp ANTENNA_636 (.A(net858));
 sg13g2_antennanp ANTENNA_637 (.A(net858));
 sg13g2_antennanp ANTENNA_638 (.A(net858));
 sg13g2_antennanp ANTENNA_639 (.A(net860));
 sg13g2_antennanp ANTENNA_640 (.A(net860));
 sg13g2_antennanp ANTENNA_641 (.A(net860));
 sg13g2_antennanp ANTENNA_642 (.A(net860));
 sg13g2_antennanp ANTENNA_643 (.A(net860));
 sg13g2_antennanp ANTENNA_644 (.A(net860));
 sg13g2_antennanp ANTENNA_645 (.A(net860));
 sg13g2_antennanp ANTENNA_646 (.A(net860));
 sg13g2_antennanp ANTENNA_647 (.A(net872));
 sg13g2_antennanp ANTENNA_648 (.A(net872));
 sg13g2_antennanp ANTENNA_649 (.A(net872));
 sg13g2_antennanp ANTENNA_650 (.A(net872));
 sg13g2_antennanp ANTENNA_651 (.A(net872));
 sg13g2_antennanp ANTENNA_652 (.A(net872));
 sg13g2_antennanp ANTENNA_653 (.A(net872));
 sg13g2_antennanp ANTENNA_654 (.A(net872));
 sg13g2_antennanp ANTENNA_655 (.A(net872));
 sg13g2_antennanp ANTENNA_656 (.A(net872));
 sg13g2_antennanp ANTENNA_657 (.A(net872));
 sg13g2_antennanp ANTENNA_658 (.A(net872));
 sg13g2_antennanp ANTENNA_659 (.A(net872));
 sg13g2_antennanp ANTENNA_660 (.A(net872));
 sg13g2_antennanp ANTENNA_661 (.A(net923));
 sg13g2_antennanp ANTENNA_662 (.A(net923));
 sg13g2_antennanp ANTENNA_663 (.A(net923));
 sg13g2_antennanp ANTENNA_664 (.A(net923));
 sg13g2_antennanp ANTENNA_665 (.A(net923));
 sg13g2_antennanp ANTENNA_666 (.A(net923));
 sg13g2_antennanp ANTENNA_667 (.A(net923));
 sg13g2_antennanp ANTENNA_668 (.A(net923));
 sg13g2_antennanp ANTENNA_669 (.A(net923));
 sg13g2_antennanp ANTENNA_670 (.A(net928));
 sg13g2_antennanp ANTENNA_671 (.A(net928));
 sg13g2_antennanp ANTENNA_672 (.A(net928));
 sg13g2_antennanp ANTENNA_673 (.A(net928));
 sg13g2_antennanp ANTENNA_674 (.A(net928));
 sg13g2_antennanp ANTENNA_675 (.A(net928));
 sg13g2_antennanp ANTENNA_676 (.A(net928));
 sg13g2_antennanp ANTENNA_677 (.A(net928));
 sg13g2_antennanp ANTENNA_678 (.A(net928));
 sg13g2_antennanp ANTENNA_679 (.A(net928));
 sg13g2_antennanp ANTENNA_680 (.A(net928));
 sg13g2_antennanp ANTENNA_681 (.A(net928));
 sg13g2_antennanp ANTENNA_682 (.A(net928));
 sg13g2_antennanp ANTENNA_683 (.A(net928));
 sg13g2_antennanp ANTENNA_684 (.A(net928));
 sg13g2_antennanp ANTENNA_685 (.A(net928));
 sg13g2_antennanp ANTENNA_686 (.A(net983));
 sg13g2_antennanp ANTENNA_687 (.A(net983));
 sg13g2_antennanp ANTENNA_688 (.A(net983));
 sg13g2_antennanp ANTENNA_689 (.A(net983));
 sg13g2_antennanp ANTENNA_690 (.A(net983));
 sg13g2_antennanp ANTENNA_691 (.A(net983));
 sg13g2_antennanp ANTENNA_692 (.A(net983));
 sg13g2_antennanp ANTENNA_693 (.A(net983));
 sg13g2_antennanp ANTENNA_694 (.A(net983));
 sg13g2_antennanp ANTENNA_695 (.A(net983));
 sg13g2_antennanp ANTENNA_696 (.A(net983));
 sg13g2_antennanp ANTENNA_697 (.A(net983));
 sg13g2_antennanp ANTENNA_698 (.A(net983));
 sg13g2_antennanp ANTENNA_699 (.A(net983));
 sg13g2_antennanp ANTENNA_700 (.A(net983));
 sg13g2_antennanp ANTENNA_701 (.A(net983));
 sg13g2_antennanp ANTENNA_702 (.A(net983));
 sg13g2_antennanp ANTENNA_703 (.A(net983));
 sg13g2_antennanp ANTENNA_704 (.A(net983));
 sg13g2_antennanp ANTENNA_705 (.A(net983));
 sg13g2_antennanp ANTENNA_706 (.A(net997));
 sg13g2_antennanp ANTENNA_707 (.A(net997));
 sg13g2_antennanp ANTENNA_708 (.A(net997));
 sg13g2_antennanp ANTENNA_709 (.A(net997));
 sg13g2_antennanp ANTENNA_710 (.A(net997));
 sg13g2_antennanp ANTENNA_711 (.A(net997));
 sg13g2_antennanp ANTENNA_712 (.A(net997));
 sg13g2_antennanp ANTENNA_713 (.A(net997));
 sg13g2_antennanp ANTENNA_714 (.A(net997));
 sg13g2_antennanp ANTENNA_715 (.A(net997));
 sg13g2_antennanp ANTENNA_716 (.A(net997));
 sg13g2_antennanp ANTENNA_717 (.A(net997));
 sg13g2_antennanp ANTENNA_718 (.A(net997));
 sg13g2_antennanp ANTENNA_719 (.A(net997));
 sg13g2_antennanp ANTENNA_720 (.A(net997));
 sg13g2_antennanp ANTENNA_721 (.A(net997));
 sg13g2_antennanp ANTENNA_722 (.A(net997));
 sg13g2_antennanp ANTENNA_723 (.A(net997));
 sg13g2_antennanp ANTENNA_724 (.A(net997));
 sg13g2_antennanp ANTENNA_725 (.A(net997));
 sg13g2_antennanp ANTENNA_726 (.A(net999));
 sg13g2_antennanp ANTENNA_727 (.A(net999));
 sg13g2_antennanp ANTENNA_728 (.A(net999));
 sg13g2_antennanp ANTENNA_729 (.A(net999));
 sg13g2_antennanp ANTENNA_730 (.A(net999));
 sg13g2_antennanp ANTENNA_731 (.A(net999));
 sg13g2_antennanp ANTENNA_732 (.A(net999));
 sg13g2_antennanp ANTENNA_733 (.A(net999));
 sg13g2_antennanp ANTENNA_734 (.A(net1000));
 sg13g2_antennanp ANTENNA_735 (.A(net1000));
 sg13g2_antennanp ANTENNA_736 (.A(net1000));
 sg13g2_antennanp ANTENNA_737 (.A(net1000));
 sg13g2_antennanp ANTENNA_738 (.A(net1000));
 sg13g2_antennanp ANTENNA_739 (.A(net1000));
 sg13g2_antennanp ANTENNA_740 (.A(net1000));
 sg13g2_antennanp ANTENNA_741 (.A(net1000));
 sg13g2_antennanp ANTENNA_742 (.A(net1000));
 sg13g2_antennanp ANTENNA_743 (.A(net1000));
 sg13g2_antennanp ANTENNA_744 (.A(net1000));
 sg13g2_antennanp ANTENNA_745 (.A(net1000));
 sg13g2_antennanp ANTENNA_746 (.A(net1000));
 sg13g2_antennanp ANTENNA_747 (.A(net1000));
 sg13g2_antennanp ANTENNA_748 (.A(net1000));
 sg13g2_antennanp ANTENNA_749 (.A(net1000));
 sg13g2_antennanp ANTENNA_750 (.A(net1000));
 sg13g2_antennanp ANTENNA_751 (.A(net1000));
 sg13g2_antennanp ANTENNA_752 (.A(net1002));
 sg13g2_antennanp ANTENNA_753 (.A(net1002));
 sg13g2_antennanp ANTENNA_754 (.A(net1002));
 sg13g2_antennanp ANTENNA_755 (.A(net1002));
 sg13g2_antennanp ANTENNA_756 (.A(net1002));
 sg13g2_antennanp ANTENNA_757 (.A(net1002));
 sg13g2_antennanp ANTENNA_758 (.A(net1002));
 sg13g2_antennanp ANTENNA_759 (.A(net1002));
 sg13g2_antennanp ANTENNA_760 (.A(net1002));
 sg13g2_antennanp ANTENNA_761 (.A(net1002));
 sg13g2_antennanp ANTENNA_762 (.A(net1002));
 sg13g2_antennanp ANTENNA_763 (.A(net1002));
 sg13g2_antennanp ANTENNA_764 (.A(net1002));
 sg13g2_antennanp ANTENNA_765 (.A(net1002));
 sg13g2_antennanp ANTENNA_766 (.A(net1002));
 sg13g2_antennanp ANTENNA_767 (.A(net1002));
 sg13g2_antennanp ANTENNA_768 (.A(net1002));
 sg13g2_antennanp ANTENNA_769 (.A(net1002));
 sg13g2_antennanp ANTENNA_770 (.A(net1002));
 sg13g2_antennanp ANTENNA_771 (.A(net1002));
 sg13g2_antennanp ANTENNA_772 (.A(net1002));
 sg13g2_antennanp ANTENNA_773 (.A(net1002));
 sg13g2_antennanp ANTENNA_774 (.A(net1002));
 sg13g2_antennanp ANTENNA_775 (.A(net1002));
 sg13g2_antennanp ANTENNA_776 (.A(net1002));
 sg13g2_antennanp ANTENNA_777 (.A(net1002));
 sg13g2_antennanp ANTENNA_778 (.A(net1002));
 sg13g2_antennanp ANTENNA_779 (.A(net1002));
 sg13g2_antennanp ANTENNA_780 (.A(net1002));
 sg13g2_antennanp ANTENNA_781 (.A(net1002));
 sg13g2_antennanp ANTENNA_782 (.A(net1002));
 sg13g2_antennanp ANTENNA_783 (.A(net1002));
 sg13g2_antennanp ANTENNA_784 (.A(net1004));
 sg13g2_antennanp ANTENNA_785 (.A(net1004));
 sg13g2_antennanp ANTENNA_786 (.A(net1004));
 sg13g2_antennanp ANTENNA_787 (.A(net1004));
 sg13g2_antennanp ANTENNA_788 (.A(net1004));
 sg13g2_antennanp ANTENNA_789 (.A(net1004));
 sg13g2_antennanp ANTENNA_790 (.A(net1004));
 sg13g2_antennanp ANTENNA_791 (.A(net1004));
 sg13g2_antennanp ANTENNA_792 (.A(net1004));
 sg13g2_antennanp ANTENNA_793 (.A(net1004));
 sg13g2_antennanp ANTENNA_794 (.A(net1004));
 sg13g2_antennanp ANTENNA_795 (.A(net1004));
 sg13g2_antennanp ANTENNA_796 (.A(net1004));
 sg13g2_antennanp ANTENNA_797 (.A(net1004));
 sg13g2_antennanp ANTENNA_798 (.A(net1004));
 sg13g2_antennanp ANTENNA_799 (.A(net1004));
 sg13g2_antennanp ANTENNA_800 (.A(net1021));
 sg13g2_antennanp ANTENNA_801 (.A(net1021));
 sg13g2_antennanp ANTENNA_802 (.A(net1021));
 sg13g2_antennanp ANTENNA_803 (.A(net1021));
 sg13g2_antennanp ANTENNA_804 (.A(net1021));
 sg13g2_antennanp ANTENNA_805 (.A(net1021));
 sg13g2_antennanp ANTENNA_806 (.A(net1021));
 sg13g2_antennanp ANTENNA_807 (.A(net1021));
 sg13g2_antennanp ANTENNA_808 (.A(net1021));
 sg13g2_antennanp ANTENNA_809 (.A(net1021));
 sg13g2_antennanp ANTENNA_810 (.A(net1021));
 sg13g2_antennanp ANTENNA_811 (.A(net1021));
 sg13g2_antennanp ANTENNA_812 (.A(net1021));
 sg13g2_antennanp ANTENNA_813 (.A(net1099));
 sg13g2_antennanp ANTENNA_814 (.A(net1099));
 sg13g2_antennanp ANTENNA_815 (.A(net1099));
 sg13g2_antennanp ANTENNA_816 (.A(net1099));
 sg13g2_antennanp ANTENNA_817 (.A(net1099));
 sg13g2_antennanp ANTENNA_818 (.A(net1099));
 sg13g2_antennanp ANTENNA_819 (.A(net1099));
 sg13g2_antennanp ANTENNA_820 (.A(net1099));
 sg13g2_antennanp ANTENNA_821 (.A(net1099));
 sg13g2_antennanp ANTENNA_822 (.A(net1099));
 sg13g2_antennanp ANTENNA_823 (.A(net1099));
 sg13g2_antennanp ANTENNA_824 (.A(net1099));
 sg13g2_antennanp ANTENNA_825 (.A(net1099));
 sg13g2_antennanp ANTENNA_826 (.A(net1099));
 sg13g2_antennanp ANTENNA_827 (.A(net1099));
 sg13g2_antennanp ANTENNA_828 (.A(net1099));
 sg13g2_antennanp ANTENNA_829 (.A(net1099));
 sg13g2_antennanp ANTENNA_830 (.A(net1099));
 sg13g2_antennanp ANTENNA_831 (.A(net1099));
 sg13g2_antennanp ANTENNA_832 (.A(net1099));
 sg13g2_antennanp ANTENNA_833 (.A(net1099));
 sg13g2_antennanp ANTENNA_834 (.A(net1099));
 sg13g2_antennanp ANTENNA_835 (.A(net1099));
 sg13g2_antennanp ANTENNA_836 (.A(net1099));
 sg13g2_antennanp ANTENNA_837 (.A(net1099));
 sg13g2_antennanp ANTENNA_838 (.A(net1099));
 sg13g2_antennanp ANTENNA_839 (.A(net1099));
 sg13g2_antennanp ANTENNA_840 (.A(net1099));
 sg13g2_antennanp ANTENNA_841 (.A(net1099));
 sg13g2_antennanp ANTENNA_842 (.A(net1099));
 sg13g2_antennanp ANTENNA_843 (.A(net1099));
 sg13g2_antennanp ANTENNA_844 (.A(net1099));
 sg13g2_antennanp ANTENNA_845 (.A(net1122));
 sg13g2_antennanp ANTENNA_846 (.A(net1122));
 sg13g2_antennanp ANTENNA_847 (.A(net1122));
 sg13g2_antennanp ANTENNA_848 (.A(net1122));
 sg13g2_antennanp ANTENNA_849 (.A(net1122));
 sg13g2_antennanp ANTENNA_850 (.A(net1122));
 sg13g2_antennanp ANTENNA_851 (.A(net1122));
 sg13g2_antennanp ANTENNA_852 (.A(net1122));
 sg13g2_antennanp ANTENNA_853 (.A(net1122));
 sg13g2_antennanp ANTENNA_854 (.A(net1122));
 sg13g2_antennanp ANTENNA_855 (.A(net1122));
 sg13g2_antennanp ANTENNA_856 (.A(net1122));
 sg13g2_antennanp ANTENNA_857 (.A(net1122));
 sg13g2_antennanp ANTENNA_858 (.A(net1122));
 sg13g2_antennanp ANTENNA_859 (.A(net1122));
 sg13g2_antennanp ANTENNA_860 (.A(net1122));
 sg13g2_antennanp ANTENNA_861 (.A(net1122));
 sg13g2_antennanp ANTENNA_862 (.A(net1122));
 sg13g2_antennanp ANTENNA_863 (.A(net1122));
 sg13g2_antennanp ANTENNA_864 (.A(_00207_));
 sg13g2_antennanp ANTENNA_865 (.A(_00785_));
 sg13g2_antennanp ANTENNA_866 (.A(_00977_));
 sg13g2_antennanp ANTENNA_867 (.A(_00977_));
 sg13g2_antennanp ANTENNA_868 (.A(_01032_));
 sg13g2_antennanp ANTENNA_869 (.A(_01047_));
 sg13g2_antennanp ANTENNA_870 (.A(_01048_));
 sg13g2_antennanp ANTENNA_871 (.A(_02836_));
 sg13g2_antennanp ANTENNA_872 (.A(_02836_));
 sg13g2_antennanp ANTENNA_873 (.A(_02836_));
 sg13g2_antennanp ANTENNA_874 (.A(_02836_));
 sg13g2_antennanp ANTENNA_875 (.A(_02845_));
 sg13g2_antennanp ANTENNA_876 (.A(_02845_));
 sg13g2_antennanp ANTENNA_877 (.A(_02845_));
 sg13g2_antennanp ANTENNA_878 (.A(_02845_));
 sg13g2_antennanp ANTENNA_879 (.A(_02845_));
 sg13g2_antennanp ANTENNA_880 (.A(_02845_));
 sg13g2_antennanp ANTENNA_881 (.A(_02845_));
 sg13g2_antennanp ANTENNA_882 (.A(_02845_));
 sg13g2_antennanp ANTENNA_883 (.A(_02845_));
 sg13g2_antennanp ANTENNA_884 (.A(_02849_));
 sg13g2_antennanp ANTENNA_885 (.A(_02849_));
 sg13g2_antennanp ANTENNA_886 (.A(_02849_));
 sg13g2_antennanp ANTENNA_887 (.A(_02849_));
 sg13g2_antennanp ANTENNA_888 (.A(_02849_));
 sg13g2_antennanp ANTENNA_889 (.A(_02849_));
 sg13g2_antennanp ANTENNA_890 (.A(_02849_));
 sg13g2_antennanp ANTENNA_891 (.A(_02849_));
 sg13g2_antennanp ANTENNA_892 (.A(_02849_));
 sg13g2_antennanp ANTENNA_893 (.A(_02861_));
 sg13g2_antennanp ANTENNA_894 (.A(_02861_));
 sg13g2_antennanp ANTENNA_895 (.A(_02861_));
 sg13g2_antennanp ANTENNA_896 (.A(_02861_));
 sg13g2_antennanp ANTENNA_897 (.A(_02954_));
 sg13g2_antennanp ANTENNA_898 (.A(_02954_));
 sg13g2_antennanp ANTENNA_899 (.A(_02954_));
 sg13g2_antennanp ANTENNA_900 (.A(_02954_));
 sg13g2_antennanp ANTENNA_901 (.A(_02954_));
 sg13g2_antennanp ANTENNA_902 (.A(_02954_));
 sg13g2_antennanp ANTENNA_903 (.A(_02954_));
 sg13g2_antennanp ANTENNA_904 (.A(_02954_));
 sg13g2_antennanp ANTENNA_905 (.A(_02976_));
 sg13g2_antennanp ANTENNA_906 (.A(_02976_));
 sg13g2_antennanp ANTENNA_907 (.A(_02976_));
 sg13g2_antennanp ANTENNA_908 (.A(_02976_));
 sg13g2_antennanp ANTENNA_909 (.A(_02976_));
 sg13g2_antennanp ANTENNA_910 (.A(_02976_));
 sg13g2_antennanp ANTENNA_911 (.A(_02976_));
 sg13g2_antennanp ANTENNA_912 (.A(_02976_));
 sg13g2_antennanp ANTENNA_913 (.A(_02976_));
 sg13g2_antennanp ANTENNA_914 (.A(_03081_));
 sg13g2_antennanp ANTENNA_915 (.A(_03148_));
 sg13g2_antennanp ANTENNA_916 (.A(_03148_));
 sg13g2_antennanp ANTENNA_917 (.A(_03237_));
 sg13g2_antennanp ANTENNA_918 (.A(_03237_));
 sg13g2_antennanp ANTENNA_919 (.A(_03237_));
 sg13g2_antennanp ANTENNA_920 (.A(_03507_));
 sg13g2_antennanp ANTENNA_921 (.A(_03507_));
 sg13g2_antennanp ANTENNA_922 (.A(_03507_));
 sg13g2_antennanp ANTENNA_923 (.A(_03507_));
 sg13g2_antennanp ANTENNA_924 (.A(_03507_));
 sg13g2_antennanp ANTENNA_925 (.A(_03507_));
 sg13g2_antennanp ANTENNA_926 (.A(_03513_));
 sg13g2_antennanp ANTENNA_927 (.A(_03513_));
 sg13g2_antennanp ANTENNA_928 (.A(_03513_));
 sg13g2_antennanp ANTENNA_929 (.A(_03513_));
 sg13g2_antennanp ANTENNA_930 (.A(_03513_));
 sg13g2_antennanp ANTENNA_931 (.A(_03513_));
 sg13g2_antennanp ANTENNA_932 (.A(_03513_));
 sg13g2_antennanp ANTENNA_933 (.A(_03513_));
 sg13g2_antennanp ANTENNA_934 (.A(_03513_));
 sg13g2_antennanp ANTENNA_935 (.A(_03539_));
 sg13g2_antennanp ANTENNA_936 (.A(_03539_));
 sg13g2_antennanp ANTENNA_937 (.A(_03539_));
 sg13g2_antennanp ANTENNA_938 (.A(_03539_));
 sg13g2_antennanp ANTENNA_939 (.A(_03539_));
 sg13g2_antennanp ANTENNA_940 (.A(_03539_));
 sg13g2_antennanp ANTENNA_941 (.A(_03539_));
 sg13g2_antennanp ANTENNA_942 (.A(_03539_));
 sg13g2_antennanp ANTENNA_943 (.A(_03539_));
 sg13g2_antennanp ANTENNA_944 (.A(_03691_));
 sg13g2_antennanp ANTENNA_945 (.A(_03691_));
 sg13g2_antennanp ANTENNA_946 (.A(_03691_));
 sg13g2_antennanp ANTENNA_947 (.A(_03691_));
 sg13g2_antennanp ANTENNA_948 (.A(_03824_));
 sg13g2_antennanp ANTENNA_949 (.A(_03835_));
 sg13g2_antennanp ANTENNA_950 (.A(_03835_));
 sg13g2_antennanp ANTENNA_951 (.A(_03835_));
 sg13g2_antennanp ANTENNA_952 (.A(_03838_));
 sg13g2_antennanp ANTENNA_953 (.A(_03838_));
 sg13g2_antennanp ANTENNA_954 (.A(_03838_));
 sg13g2_antennanp ANTENNA_955 (.A(_03838_));
 sg13g2_antennanp ANTENNA_956 (.A(_03838_));
 sg13g2_antennanp ANTENNA_957 (.A(_03838_));
 sg13g2_antennanp ANTENNA_958 (.A(_04855_));
 sg13g2_antennanp ANTENNA_959 (.A(_04980_));
 sg13g2_antennanp ANTENNA_960 (.A(_04980_));
 sg13g2_antennanp ANTENNA_961 (.A(_04980_));
 sg13g2_antennanp ANTENNA_962 (.A(_04980_));
 sg13g2_antennanp ANTENNA_963 (.A(_05006_));
 sg13g2_antennanp ANTENNA_964 (.A(_05157_));
 sg13g2_antennanp ANTENNA_965 (.A(_05199_));
 sg13g2_antennanp ANTENNA_966 (.A(_05260_));
 sg13g2_antennanp ANTENNA_967 (.A(_05270_));
 sg13g2_antennanp ANTENNA_968 (.A(_05287_));
 sg13g2_antennanp ANTENNA_969 (.A(_05307_));
 sg13g2_antennanp ANTENNA_970 (.A(_05314_));
 sg13g2_antennanp ANTENNA_971 (.A(_05464_));
 sg13g2_antennanp ANTENNA_972 (.A(_05525_));
 sg13g2_antennanp ANTENNA_973 (.A(_05529_));
 sg13g2_antennanp ANTENNA_974 (.A(_05607_));
 sg13g2_antennanp ANTENNA_975 (.A(_05676_));
 sg13g2_antennanp ANTENNA_976 (.A(_05754_));
 sg13g2_antennanp ANTENNA_977 (.A(_05756_));
 sg13g2_antennanp ANTENNA_978 (.A(_05770_));
 sg13g2_antennanp ANTENNA_979 (.A(_05780_));
 sg13g2_antennanp ANTENNA_980 (.A(_05780_));
 sg13g2_antennanp ANTENNA_981 (.A(_05780_));
 sg13g2_antennanp ANTENNA_982 (.A(_05780_));
 sg13g2_antennanp ANTENNA_983 (.A(_05796_));
 sg13g2_antennanp ANTENNA_984 (.A(_06579_));
 sg13g2_antennanp ANTENNA_985 (.A(_06579_));
 sg13g2_antennanp ANTENNA_986 (.A(_06579_));
 sg13g2_antennanp ANTENNA_987 (.A(_06579_));
 sg13g2_antennanp ANTENNA_988 (.A(_06579_));
 sg13g2_antennanp ANTENNA_989 (.A(_06579_));
 sg13g2_antennanp ANTENNA_990 (.A(_06579_));
 sg13g2_antennanp ANTENNA_991 (.A(_06579_));
 sg13g2_antennanp ANTENNA_992 (.A(_06579_));
 sg13g2_antennanp ANTENNA_993 (.A(_06582_));
 sg13g2_antennanp ANTENNA_994 (.A(_06582_));
 sg13g2_antennanp ANTENNA_995 (.A(_06582_));
 sg13g2_antennanp ANTENNA_996 (.A(_06582_));
 sg13g2_antennanp ANTENNA_997 (.A(_06583_));
 sg13g2_antennanp ANTENNA_998 (.A(_06583_));
 sg13g2_antennanp ANTENNA_999 (.A(_06583_));
 sg13g2_antennanp ANTENNA_1000 (.A(_06583_));
 sg13g2_antennanp ANTENNA_1001 (.A(_06583_));
 sg13g2_antennanp ANTENNA_1002 (.A(_06583_));
 sg13g2_antennanp ANTENNA_1003 (.A(_06583_));
 sg13g2_antennanp ANTENNA_1004 (.A(_06583_));
 sg13g2_antennanp ANTENNA_1005 (.A(_06583_));
 sg13g2_antennanp ANTENNA_1006 (.A(_06885_));
 sg13g2_antennanp ANTENNA_1007 (.A(_06885_));
 sg13g2_antennanp ANTENNA_1008 (.A(_06885_));
 sg13g2_antennanp ANTENNA_1009 (.A(_06885_));
 sg13g2_antennanp ANTENNA_1010 (.A(_06885_));
 sg13g2_antennanp ANTENNA_1011 (.A(_06885_));
 sg13g2_antennanp ANTENNA_1012 (.A(_06885_));
 sg13g2_antennanp ANTENNA_1013 (.A(_06885_));
 sg13g2_antennanp ANTENNA_1014 (.A(_06885_));
 sg13g2_antennanp ANTENNA_1015 (.A(_06885_));
 sg13g2_antennanp ANTENNA_1016 (.A(_07626_));
 sg13g2_antennanp ANTENNA_1017 (.A(_07626_));
 sg13g2_antennanp ANTENNA_1018 (.A(_07632_));
 sg13g2_antennanp ANTENNA_1019 (.A(_07634_));
 sg13g2_antennanp ANTENNA_1020 (.A(_07634_));
 sg13g2_antennanp ANTENNA_1021 (.A(_07851_));
 sg13g2_antennanp ANTENNA_1022 (.A(_07851_));
 sg13g2_antennanp ANTENNA_1023 (.A(_07851_));
 sg13g2_antennanp ANTENNA_1024 (.A(_07851_));
 sg13g2_antennanp ANTENNA_1025 (.A(_07851_));
 sg13g2_antennanp ANTENNA_1026 (.A(_07851_));
 sg13g2_antennanp ANTENNA_1027 (.A(_07851_));
 sg13g2_antennanp ANTENNA_1028 (.A(_07851_));
 sg13g2_antennanp ANTENNA_1029 (.A(_07851_));
 sg13g2_antennanp ANTENNA_1030 (.A(_07851_));
 sg13g2_antennanp ANTENNA_1031 (.A(_08260_));
 sg13g2_antennanp ANTENNA_1032 (.A(_08260_));
 sg13g2_antennanp ANTENNA_1033 (.A(_08260_));
 sg13g2_antennanp ANTENNA_1034 (.A(_08346_));
 sg13g2_antennanp ANTENNA_1035 (.A(_08346_));
 sg13g2_antennanp ANTENNA_1036 (.A(_08346_));
 sg13g2_antennanp ANTENNA_1037 (.A(_08346_));
 sg13g2_antennanp ANTENNA_1038 (.A(_08346_));
 sg13g2_antennanp ANTENNA_1039 (.A(_08346_));
 sg13g2_antennanp ANTENNA_1040 (.A(_08346_));
 sg13g2_antennanp ANTENNA_1041 (.A(_08346_));
 sg13g2_antennanp ANTENNA_1042 (.A(_08455_));
 sg13g2_antennanp ANTENNA_1043 (.A(_08455_));
 sg13g2_antennanp ANTENNA_1044 (.A(_08455_));
 sg13g2_antennanp ANTENNA_1045 (.A(_08455_));
 sg13g2_antennanp ANTENNA_1046 (.A(_08497_));
 sg13g2_antennanp ANTENNA_1047 (.A(_08497_));
 sg13g2_antennanp ANTENNA_1048 (.A(_08497_));
 sg13g2_antennanp ANTENNA_1049 (.A(_08565_));
 sg13g2_antennanp ANTENNA_1050 (.A(_08565_));
 sg13g2_antennanp ANTENNA_1051 (.A(_08565_));
 sg13g2_antennanp ANTENNA_1052 (.A(_08565_));
 sg13g2_antennanp ANTENNA_1053 (.A(_08565_));
 sg13g2_antennanp ANTENNA_1054 (.A(_08565_));
 sg13g2_antennanp ANTENNA_1055 (.A(_08603_));
 sg13g2_antennanp ANTENNA_1056 (.A(_08603_));
 sg13g2_antennanp ANTENNA_1057 (.A(_08603_));
 sg13g2_antennanp ANTENNA_1058 (.A(_08633_));
 sg13g2_antennanp ANTENNA_1059 (.A(_08663_));
 sg13g2_antennanp ANTENNA_1060 (.A(_08663_));
 sg13g2_antennanp ANTENNA_1061 (.A(_08663_));
 sg13g2_antennanp ANTENNA_1062 (.A(_08663_));
 sg13g2_antennanp ANTENNA_1063 (.A(_08663_));
 sg13g2_antennanp ANTENNA_1064 (.A(_08663_));
 sg13g2_antennanp ANTENNA_1065 (.A(_08663_));
 sg13g2_antennanp ANTENNA_1066 (.A(_08663_));
 sg13g2_antennanp ANTENNA_1067 (.A(_08663_));
 sg13g2_antennanp ANTENNA_1068 (.A(_08777_));
 sg13g2_antennanp ANTENNA_1069 (.A(_08799_));
 sg13g2_antennanp ANTENNA_1070 (.A(_08799_));
 sg13g2_antennanp ANTENNA_1071 (.A(_08799_));
 sg13g2_antennanp ANTENNA_1072 (.A(_08799_));
 sg13g2_antennanp ANTENNA_1073 (.A(_08799_));
 sg13g2_antennanp ANTENNA_1074 (.A(_08799_));
 sg13g2_antennanp ANTENNA_1075 (.A(_08820_));
 sg13g2_antennanp ANTENNA_1076 (.A(_08820_));
 sg13g2_antennanp ANTENNA_1077 (.A(_08820_));
 sg13g2_antennanp ANTENNA_1078 (.A(_08820_));
 sg13g2_antennanp ANTENNA_1079 (.A(_08820_));
 sg13g2_antennanp ANTENNA_1080 (.A(_08820_));
 sg13g2_antennanp ANTENNA_1081 (.A(_08826_));
 sg13g2_antennanp ANTENNA_1082 (.A(_08826_));
 sg13g2_antennanp ANTENNA_1083 (.A(_08826_));
 sg13g2_antennanp ANTENNA_1084 (.A(_08826_));
 sg13g2_antennanp ANTENNA_1085 (.A(_08826_));
 sg13g2_antennanp ANTENNA_1086 (.A(_08826_));
 sg13g2_antennanp ANTENNA_1087 (.A(_08840_));
 sg13g2_antennanp ANTENNA_1088 (.A(_08840_));
 sg13g2_antennanp ANTENNA_1089 (.A(_08840_));
 sg13g2_antennanp ANTENNA_1090 (.A(_08840_));
 sg13g2_antennanp ANTENNA_1091 (.A(_08848_));
 sg13g2_antennanp ANTENNA_1092 (.A(_08848_));
 sg13g2_antennanp ANTENNA_1093 (.A(_08848_));
 sg13g2_antennanp ANTENNA_1094 (.A(_08868_));
 sg13g2_antennanp ANTENNA_1095 (.A(_08900_));
 sg13g2_antennanp ANTENNA_1096 (.A(_08900_));
 sg13g2_antennanp ANTENNA_1097 (.A(_08900_));
 sg13g2_antennanp ANTENNA_1098 (.A(_08950_));
 sg13g2_antennanp ANTENNA_1099 (.A(_08950_));
 sg13g2_antennanp ANTENNA_1100 (.A(_08950_));
 sg13g2_antennanp ANTENNA_1101 (.A(_08950_));
 sg13g2_antennanp ANTENNA_1102 (.A(_08950_));
 sg13g2_antennanp ANTENNA_1103 (.A(_08950_));
 sg13g2_antennanp ANTENNA_1104 (.A(_08950_));
 sg13g2_antennanp ANTENNA_1105 (.A(_08950_));
 sg13g2_antennanp ANTENNA_1106 (.A(_08950_));
 sg13g2_antennanp ANTENNA_1107 (.A(_08950_));
 sg13g2_antennanp ANTENNA_1108 (.A(_08950_));
 sg13g2_antennanp ANTENNA_1109 (.A(_08950_));
 sg13g2_antennanp ANTENNA_1110 (.A(_08950_));
 sg13g2_antennanp ANTENNA_1111 (.A(_08950_));
 sg13g2_antennanp ANTENNA_1112 (.A(_08970_));
 sg13g2_antennanp ANTENNA_1113 (.A(_08970_));
 sg13g2_antennanp ANTENNA_1114 (.A(_08986_));
 sg13g2_antennanp ANTENNA_1115 (.A(_08986_));
 sg13g2_antennanp ANTENNA_1116 (.A(_09002_));
 sg13g2_antennanp ANTENNA_1117 (.A(_09002_));
 sg13g2_antennanp ANTENNA_1118 (.A(_09065_));
 sg13g2_antennanp ANTENNA_1119 (.A(_09065_));
 sg13g2_antennanp ANTENNA_1120 (.A(_09091_));
 sg13g2_antennanp ANTENNA_1121 (.A(_09091_));
 sg13g2_antennanp ANTENNA_1122 (.A(_09091_));
 sg13g2_antennanp ANTENNA_1123 (.A(_09091_));
 sg13g2_antennanp ANTENNA_1124 (.A(_09091_));
 sg13g2_antennanp ANTENNA_1125 (.A(_09091_));
 sg13g2_antennanp ANTENNA_1126 (.A(_09091_));
 sg13g2_antennanp ANTENNA_1127 (.A(_09091_));
 sg13g2_antennanp ANTENNA_1128 (.A(_09091_));
 sg13g2_antennanp ANTENNA_1129 (.A(_09120_));
 sg13g2_antennanp ANTENNA_1130 (.A(_09120_));
 sg13g2_antennanp ANTENNA_1131 (.A(_09158_));
 sg13g2_antennanp ANTENNA_1132 (.A(_09158_));
 sg13g2_antennanp ANTENNA_1133 (.A(_09158_));
 sg13g2_antennanp ANTENNA_1134 (.A(_09173_));
 sg13g2_antennanp ANTENNA_1135 (.A(_09211_));
 sg13g2_antennanp ANTENNA_1136 (.A(_09211_));
 sg13g2_antennanp ANTENNA_1137 (.A(_09211_));
 sg13g2_antennanp ANTENNA_1138 (.A(_09211_));
 sg13g2_antennanp ANTENNA_1139 (.A(_09211_));
 sg13g2_antennanp ANTENNA_1140 (.A(_09218_));
 sg13g2_antennanp ANTENNA_1141 (.A(_09220_));
 sg13g2_antennanp ANTENNA_1142 (.A(_09220_));
 sg13g2_antennanp ANTENNA_1143 (.A(_09220_));
 sg13g2_antennanp ANTENNA_1144 (.A(_09220_));
 sg13g2_antennanp ANTENNA_1145 (.A(_09220_));
 sg13g2_antennanp ANTENNA_1146 (.A(_09220_));
 sg13g2_antennanp ANTENNA_1147 (.A(_09220_));
 sg13g2_antennanp ANTENNA_1148 (.A(_09220_));
 sg13g2_antennanp ANTENNA_1149 (.A(_09220_));
 sg13g2_antennanp ANTENNA_1150 (.A(_09220_));
 sg13g2_antennanp ANTENNA_1151 (.A(_09220_));
 sg13g2_antennanp ANTENNA_1152 (.A(_09220_));
 sg13g2_antennanp ANTENNA_1153 (.A(_09220_));
 sg13g2_antennanp ANTENNA_1154 (.A(_09223_));
 sg13g2_antennanp ANTENNA_1155 (.A(_09223_));
 sg13g2_antennanp ANTENNA_1156 (.A(_09223_));
 sg13g2_antennanp ANTENNA_1157 (.A(_09223_));
 sg13g2_antennanp ANTENNA_1158 (.A(_09223_));
 sg13g2_antennanp ANTENNA_1159 (.A(_09223_));
 sg13g2_antennanp ANTENNA_1160 (.A(_09223_));
 sg13g2_antennanp ANTENNA_1161 (.A(_09223_));
 sg13g2_antennanp ANTENNA_1162 (.A(_09318_));
 sg13g2_antennanp ANTENNA_1163 (.A(_09318_));
 sg13g2_antennanp ANTENNA_1164 (.A(_09318_));
 sg13g2_antennanp ANTENNA_1165 (.A(_09361_));
 sg13g2_antennanp ANTENNA_1166 (.A(_09361_));
 sg13g2_antennanp ANTENNA_1167 (.A(_09361_));
 sg13g2_antennanp ANTENNA_1168 (.A(_09361_));
 sg13g2_antennanp ANTENNA_1169 (.A(_09361_));
 sg13g2_antennanp ANTENNA_1170 (.A(_09361_));
 sg13g2_antennanp ANTENNA_1171 (.A(_09394_));
 sg13g2_antennanp ANTENNA_1172 (.A(_09396_));
 sg13g2_antennanp ANTENNA_1173 (.A(_09447_));
 sg13g2_antennanp ANTENNA_1174 (.A(_09448_));
 sg13g2_antennanp ANTENNA_1175 (.A(_09448_));
 sg13g2_antennanp ANTENNA_1176 (.A(_09448_));
 sg13g2_antennanp ANTENNA_1177 (.A(_09448_));
 sg13g2_antennanp ANTENNA_1178 (.A(_09450_));
 sg13g2_antennanp ANTENNA_1179 (.A(_09492_));
 sg13g2_antennanp ANTENNA_1180 (.A(_09544_));
 sg13g2_antennanp ANTENNA_1181 (.A(_09657_));
 sg13g2_antennanp ANTENNA_1182 (.A(_09678_));
 sg13g2_antennanp ANTENNA_1183 (.A(_09722_));
 sg13g2_antennanp ANTENNA_1184 (.A(_09769_));
 sg13g2_antennanp ANTENNA_1185 (.A(_09791_));
 sg13g2_antennanp ANTENNA_1186 (.A(_09852_));
 sg13g2_antennanp ANTENNA_1187 (.A(_09852_));
 sg13g2_antennanp ANTENNA_1188 (.A(_09852_));
 sg13g2_antennanp ANTENNA_1189 (.A(_09852_));
 sg13g2_antennanp ANTENNA_1190 (.A(_09852_));
 sg13g2_antennanp ANTENNA_1191 (.A(_09852_));
 sg13g2_antennanp ANTENNA_1192 (.A(_09852_));
 sg13g2_antennanp ANTENNA_1193 (.A(_09852_));
 sg13g2_antennanp ANTENNA_1194 (.A(_09852_));
 sg13g2_antennanp ANTENNA_1195 (.A(_09852_));
 sg13g2_antennanp ANTENNA_1196 (.A(_09852_));
 sg13g2_antennanp ANTENNA_1197 (.A(_09852_));
 sg13g2_antennanp ANTENNA_1198 (.A(_09852_));
 sg13g2_antennanp ANTENNA_1199 (.A(_10042_));
 sg13g2_antennanp ANTENNA_1200 (.A(_10042_));
 sg13g2_antennanp ANTENNA_1201 (.A(_10042_));
 sg13g2_antennanp ANTENNA_1202 (.A(_10121_));
 sg13g2_antennanp ANTENNA_1203 (.A(_10121_));
 sg13g2_antennanp ANTENNA_1204 (.A(_10121_));
 sg13g2_antennanp ANTENNA_1205 (.A(_10146_));
 sg13g2_antennanp ANTENNA_1206 (.A(_10146_));
 sg13g2_antennanp ANTENNA_1207 (.A(_10146_));
 sg13g2_antennanp ANTENNA_1208 (.A(_10146_));
 sg13g2_antennanp ANTENNA_1209 (.A(_10146_));
 sg13g2_antennanp ANTENNA_1210 (.A(_10146_));
 sg13g2_antennanp ANTENNA_1211 (.A(_10146_));
 sg13g2_antennanp ANTENNA_1212 (.A(_10146_));
 sg13g2_antennanp ANTENNA_1213 (.A(_10162_));
 sg13g2_antennanp ANTENNA_1214 (.A(_10162_));
 sg13g2_antennanp ANTENNA_1215 (.A(_10162_));
 sg13g2_antennanp ANTENNA_1216 (.A(_10162_));
 sg13g2_antennanp ANTENNA_1217 (.A(_10162_));
 sg13g2_antennanp ANTENNA_1218 (.A(_10162_));
 sg13g2_antennanp ANTENNA_1219 (.A(_10162_));
 sg13g2_antennanp ANTENNA_1220 (.A(_10162_));
 sg13g2_antennanp ANTENNA_1221 (.A(_10379_));
 sg13g2_antennanp ANTENNA_1222 (.A(_10379_));
 sg13g2_antennanp ANTENNA_1223 (.A(_10379_));
 sg13g2_antennanp ANTENNA_1224 (.A(_10642_));
 sg13g2_antennanp ANTENNA_1225 (.A(_10642_));
 sg13g2_antennanp ANTENNA_1226 (.A(_10642_));
 sg13g2_antennanp ANTENNA_1227 (.A(_10642_));
 sg13g2_antennanp ANTENNA_1228 (.A(_10642_));
 sg13g2_antennanp ANTENNA_1229 (.A(_10642_));
 sg13g2_antennanp ANTENNA_1230 (.A(_10642_));
 sg13g2_antennanp ANTENNA_1231 (.A(_10744_));
 sg13g2_antennanp ANTENNA_1232 (.A(_10744_));
 sg13g2_antennanp ANTENNA_1233 (.A(_10744_));
 sg13g2_antennanp ANTENNA_1234 (.A(_10744_));
 sg13g2_antennanp ANTENNA_1235 (.A(_12205_));
 sg13g2_antennanp ANTENNA_1236 (.A(_12205_));
 sg13g2_antennanp ANTENNA_1237 (.A(_12205_));
 sg13g2_antennanp ANTENNA_1238 (.A(_12205_));
 sg13g2_antennanp ANTENNA_1239 (.A(_12218_));
 sg13g2_antennanp ANTENNA_1240 (.A(_12218_));
 sg13g2_antennanp ANTENNA_1241 (.A(_12218_));
 sg13g2_antennanp ANTENNA_1242 (.A(_12218_));
 sg13g2_antennanp ANTENNA_1243 (.A(_12218_));
 sg13g2_antennanp ANTENNA_1244 (.A(_12218_));
 sg13g2_antennanp ANTENNA_1245 (.A(_12218_));
 sg13g2_antennanp ANTENNA_1246 (.A(_12218_));
 sg13g2_antennanp ANTENNA_1247 (.A(_12218_));
 sg13g2_antennanp ANTENNA_1248 (.A(_12218_));
 sg13g2_antennanp ANTENNA_1249 (.A(_12218_));
 sg13g2_antennanp ANTENNA_1250 (.A(_12218_));
 sg13g2_antennanp ANTENNA_1251 (.A(_12218_));
 sg13g2_antennanp ANTENNA_1252 (.A(_12218_));
 sg13g2_antennanp ANTENNA_1253 (.A(_12218_));
 sg13g2_antennanp ANTENNA_1254 (.A(_12218_));
 sg13g2_antennanp ANTENNA_1255 (.A(_12218_));
 sg13g2_antennanp ANTENNA_1256 (.A(_12218_));
 sg13g2_antennanp ANTENNA_1257 (.A(_12225_));
 sg13g2_antennanp ANTENNA_1258 (.A(_12225_));
 sg13g2_antennanp ANTENNA_1259 (.A(_12225_));
 sg13g2_antennanp ANTENNA_1260 (.A(_12225_));
 sg13g2_antennanp ANTENNA_1261 (.A(_12225_));
 sg13g2_antennanp ANTENNA_1262 (.A(_12225_));
 sg13g2_antennanp ANTENNA_1263 (.A(_12225_));
 sg13g2_antennanp ANTENNA_1264 (.A(_12225_));
 sg13g2_antennanp ANTENNA_1265 (.A(_12225_));
 sg13g2_antennanp ANTENNA_1266 (.A(_12225_));
 sg13g2_antennanp ANTENNA_1267 (.A(_12225_));
 sg13g2_antennanp ANTENNA_1268 (.A(_12225_));
 sg13g2_antennanp ANTENNA_1269 (.A(_12225_));
 sg13g2_antennanp ANTENNA_1270 (.A(_12225_));
 sg13g2_antennanp ANTENNA_1271 (.A(_12225_));
 sg13g2_antennanp ANTENNA_1272 (.A(_12225_));
 sg13g2_antennanp ANTENNA_1273 (.A(_12225_));
 sg13g2_antennanp ANTENNA_1274 (.A(_12225_));
 sg13g2_antennanp ANTENNA_1275 (.A(_12236_));
 sg13g2_antennanp ANTENNA_1276 (.A(_12236_));
 sg13g2_antennanp ANTENNA_1277 (.A(_12236_));
 sg13g2_antennanp ANTENNA_1278 (.A(_12236_));
 sg13g2_antennanp ANTENNA_1279 (.A(_12236_));
 sg13g2_antennanp ANTENNA_1280 (.A(_12236_));
 sg13g2_antennanp ANTENNA_1281 (.A(_12236_));
 sg13g2_antennanp ANTENNA_1282 (.A(_12236_));
 sg13g2_antennanp ANTENNA_1283 (.A(_12236_));
 sg13g2_antennanp ANTENNA_1284 (.A(\cpu.dcache.wdata[10] ));
 sg13g2_antennanp ANTENNA_1285 (.A(\cpu.dcache.wdata[10] ));
 sg13g2_antennanp ANTENNA_1286 (.A(\cpu.dcache.wdata[10] ));
 sg13g2_antennanp ANTENNA_1287 (.A(\cpu.dcache.wdata[10] ));
 sg13g2_antennanp ANTENNA_1288 (.A(\cpu.dcache.wdata[12] ));
 sg13g2_antennanp ANTENNA_1289 (.A(\cpu.dcache.wdata[12] ));
 sg13g2_antennanp ANTENNA_1290 (.A(\cpu.dcache.wdata[12] ));
 sg13g2_antennanp ANTENNA_1291 (.A(\cpu.dcache.wdata[12] ));
 sg13g2_antennanp ANTENNA_1292 (.A(\cpu.dcache.wdata[9] ));
 sg13g2_antennanp ANTENNA_1293 (.A(\cpu.dcache.wdata[9] ));
 sg13g2_antennanp ANTENNA_1294 (.A(\cpu.dcache.wdata[9] ));
 sg13g2_antennanp ANTENNA_1295 (.A(\cpu.dcache.wdata[9] ));
 sg13g2_antennanp ANTENNA_1296 (.A(\cpu.ex.pc[1] ));
 sg13g2_antennanp ANTENNA_1297 (.A(\cpu.ex.pc[2] ));
 sg13g2_antennanp ANTENNA_1298 (.A(\cpu.gpio.uart_rx ));
 sg13g2_antennanp ANTENNA_1299 (.A(\cpu.gpio.uart_rx ));
 sg13g2_antennanp ANTENNA_1300 (.A(\cpu.qspi.c_wstrobe_i ));
 sg13g2_antennanp ANTENNA_1301 (.A(\cpu.qspi.c_wstrobe_i ));
 sg13g2_antennanp ANTENNA_1302 (.A(net3));
 sg13g2_antennanp ANTENNA_1303 (.A(net3));
 sg13g2_antennanp ANTENNA_1304 (.A(net3));
 sg13g2_antennanp ANTENNA_1305 (.A(net11));
 sg13g2_antennanp ANTENNA_1306 (.A(net11));
 sg13g2_antennanp ANTENNA_1307 (.A(net11));
 sg13g2_antennanp ANTENNA_1308 (.A(net12));
 sg13g2_antennanp ANTENNA_1309 (.A(net12));
 sg13g2_antennanp ANTENNA_1310 (.A(net12));
 sg13g2_antennanp ANTENNA_1311 (.A(net13));
 sg13g2_antennanp ANTENNA_1312 (.A(net13));
 sg13g2_antennanp ANTENNA_1313 (.A(net13));
 sg13g2_antennanp ANTENNA_1314 (.A(net14));
 sg13g2_antennanp ANTENNA_1315 (.A(net14));
 sg13g2_antennanp ANTENNA_1316 (.A(net14));
 sg13g2_antennanp ANTENNA_1317 (.A(net36));
 sg13g2_antennanp ANTENNA_1318 (.A(net36));
 sg13g2_antennanp ANTENNA_1319 (.A(net36));
 sg13g2_antennanp ANTENNA_1320 (.A(net36));
 sg13g2_antennanp ANTENNA_1321 (.A(net36));
 sg13g2_antennanp ANTENNA_1322 (.A(net36));
 sg13g2_antennanp ANTENNA_1323 (.A(net36));
 sg13g2_antennanp ANTENNA_1324 (.A(net36));
 sg13g2_antennanp ANTENNA_1325 (.A(net36));
 sg13g2_antennanp ANTENNA_1326 (.A(net36));
 sg13g2_antennanp ANTENNA_1327 (.A(net36));
 sg13g2_antennanp ANTENNA_1328 (.A(net36));
 sg13g2_antennanp ANTENNA_1329 (.A(net36));
 sg13g2_antennanp ANTENNA_1330 (.A(net36));
 sg13g2_antennanp ANTENNA_1331 (.A(net36));
 sg13g2_antennanp ANTENNA_1332 (.A(net36));
 sg13g2_antennanp ANTENNA_1333 (.A(net36));
 sg13g2_antennanp ANTENNA_1334 (.A(net36));
 sg13g2_antennanp ANTENNA_1335 (.A(net36));
 sg13g2_antennanp ANTENNA_1336 (.A(net36));
 sg13g2_antennanp ANTENNA_1337 (.A(net36));
 sg13g2_antennanp ANTENNA_1338 (.A(net36));
 sg13g2_antennanp ANTENNA_1339 (.A(net36));
 sg13g2_antennanp ANTENNA_1340 (.A(net114));
 sg13g2_antennanp ANTENNA_1341 (.A(net114));
 sg13g2_antennanp ANTENNA_1342 (.A(net114));
 sg13g2_antennanp ANTENNA_1343 (.A(net114));
 sg13g2_antennanp ANTENNA_1344 (.A(net114));
 sg13g2_antennanp ANTENNA_1345 (.A(net114));
 sg13g2_antennanp ANTENNA_1346 (.A(net114));
 sg13g2_antennanp ANTENNA_1347 (.A(net114));
 sg13g2_antennanp ANTENNA_1348 (.A(net114));
 sg13g2_antennanp ANTENNA_1349 (.A(net114));
 sg13g2_antennanp ANTENNA_1350 (.A(net114));
 sg13g2_antennanp ANTENNA_1351 (.A(net114));
 sg13g2_antennanp ANTENNA_1352 (.A(net114));
 sg13g2_antennanp ANTENNA_1353 (.A(net114));
 sg13g2_antennanp ANTENNA_1354 (.A(net114));
 sg13g2_antennanp ANTENNA_1355 (.A(net114));
 sg13g2_antennanp ANTENNA_1356 (.A(net452));
 sg13g2_antennanp ANTENNA_1357 (.A(net452));
 sg13g2_antennanp ANTENNA_1358 (.A(net452));
 sg13g2_antennanp ANTENNA_1359 (.A(net452));
 sg13g2_antennanp ANTENNA_1360 (.A(net452));
 sg13g2_antennanp ANTENNA_1361 (.A(net452));
 sg13g2_antennanp ANTENNA_1362 (.A(net452));
 sg13g2_antennanp ANTENNA_1363 (.A(net452));
 sg13g2_antennanp ANTENNA_1364 (.A(net489));
 sg13g2_antennanp ANTENNA_1365 (.A(net489));
 sg13g2_antennanp ANTENNA_1366 (.A(net489));
 sg13g2_antennanp ANTENNA_1367 (.A(net489));
 sg13g2_antennanp ANTENNA_1368 (.A(net489));
 sg13g2_antennanp ANTENNA_1369 (.A(net489));
 sg13g2_antennanp ANTENNA_1370 (.A(net489));
 sg13g2_antennanp ANTENNA_1371 (.A(net489));
 sg13g2_antennanp ANTENNA_1372 (.A(net489));
 sg13g2_antennanp ANTENNA_1373 (.A(net491));
 sg13g2_antennanp ANTENNA_1374 (.A(net491));
 sg13g2_antennanp ANTENNA_1375 (.A(net491));
 sg13g2_antennanp ANTENNA_1376 (.A(net491));
 sg13g2_antennanp ANTENNA_1377 (.A(net491));
 sg13g2_antennanp ANTENNA_1378 (.A(net491));
 sg13g2_antennanp ANTENNA_1379 (.A(net491));
 sg13g2_antennanp ANTENNA_1380 (.A(net491));
 sg13g2_antennanp ANTENNA_1381 (.A(net550));
 sg13g2_antennanp ANTENNA_1382 (.A(net550));
 sg13g2_antennanp ANTENNA_1383 (.A(net550));
 sg13g2_antennanp ANTENNA_1384 (.A(net550));
 sg13g2_antennanp ANTENNA_1385 (.A(net550));
 sg13g2_antennanp ANTENNA_1386 (.A(net550));
 sg13g2_antennanp ANTENNA_1387 (.A(net550));
 sg13g2_antennanp ANTENNA_1388 (.A(net550));
 sg13g2_antennanp ANTENNA_1389 (.A(net550));
 sg13g2_antennanp ANTENNA_1390 (.A(net550));
 sg13g2_antennanp ANTENNA_1391 (.A(net550));
 sg13g2_antennanp ANTENNA_1392 (.A(net550));
 sg13g2_antennanp ANTENNA_1393 (.A(net550));
 sg13g2_antennanp ANTENNA_1394 (.A(net550));
 sg13g2_antennanp ANTENNA_1395 (.A(net622));
 sg13g2_antennanp ANTENNA_1396 (.A(net622));
 sg13g2_antennanp ANTENNA_1397 (.A(net622));
 sg13g2_antennanp ANTENNA_1398 (.A(net622));
 sg13g2_antennanp ANTENNA_1399 (.A(net622));
 sg13g2_antennanp ANTENNA_1400 (.A(net622));
 sg13g2_antennanp ANTENNA_1401 (.A(net622));
 sg13g2_antennanp ANTENNA_1402 (.A(net622));
 sg13g2_antennanp ANTENNA_1403 (.A(net622));
 sg13g2_antennanp ANTENNA_1404 (.A(net622));
 sg13g2_antennanp ANTENNA_1405 (.A(net622));
 sg13g2_antennanp ANTENNA_1406 (.A(net622));
 sg13g2_antennanp ANTENNA_1407 (.A(net622));
 sg13g2_antennanp ANTENNA_1408 (.A(net686));
 sg13g2_antennanp ANTENNA_1409 (.A(net686));
 sg13g2_antennanp ANTENNA_1410 (.A(net686));
 sg13g2_antennanp ANTENNA_1411 (.A(net686));
 sg13g2_antennanp ANTENNA_1412 (.A(net686));
 sg13g2_antennanp ANTENNA_1413 (.A(net686));
 sg13g2_antennanp ANTENNA_1414 (.A(net686));
 sg13g2_antennanp ANTENNA_1415 (.A(net686));
 sg13g2_antennanp ANTENNA_1416 (.A(net745));
 sg13g2_antennanp ANTENNA_1417 (.A(net745));
 sg13g2_antennanp ANTENNA_1418 (.A(net745));
 sg13g2_antennanp ANTENNA_1419 (.A(net745));
 sg13g2_antennanp ANTENNA_1420 (.A(net745));
 sg13g2_antennanp ANTENNA_1421 (.A(net745));
 sg13g2_antennanp ANTENNA_1422 (.A(net745));
 sg13g2_antennanp ANTENNA_1423 (.A(net745));
 sg13g2_antennanp ANTENNA_1424 (.A(net800));
 sg13g2_antennanp ANTENNA_1425 (.A(net800));
 sg13g2_antennanp ANTENNA_1426 (.A(net800));
 sg13g2_antennanp ANTENNA_1427 (.A(net800));
 sg13g2_antennanp ANTENNA_1428 (.A(net800));
 sg13g2_antennanp ANTENNA_1429 (.A(net800));
 sg13g2_antennanp ANTENNA_1430 (.A(net800));
 sg13g2_antennanp ANTENNA_1431 (.A(net800));
 sg13g2_antennanp ANTENNA_1432 (.A(net800));
 sg13g2_antennanp ANTENNA_1433 (.A(net803));
 sg13g2_antennanp ANTENNA_1434 (.A(net803));
 sg13g2_antennanp ANTENNA_1435 (.A(net803));
 sg13g2_antennanp ANTENNA_1436 (.A(net803));
 sg13g2_antennanp ANTENNA_1437 (.A(net803));
 sg13g2_antennanp ANTENNA_1438 (.A(net803));
 sg13g2_antennanp ANTENNA_1439 (.A(net803));
 sg13g2_antennanp ANTENNA_1440 (.A(net803));
 sg13g2_antennanp ANTENNA_1441 (.A(net803));
 sg13g2_antennanp ANTENNA_1442 (.A(net803));
 sg13g2_antennanp ANTENNA_1443 (.A(net803));
 sg13g2_antennanp ANTENNA_1444 (.A(net803));
 sg13g2_antennanp ANTENNA_1445 (.A(net803));
 sg13g2_antennanp ANTENNA_1446 (.A(net803));
 sg13g2_antennanp ANTENNA_1447 (.A(net803));
 sg13g2_antennanp ANTENNA_1448 (.A(net803));
 sg13g2_antennanp ANTENNA_1449 (.A(net858));
 sg13g2_antennanp ANTENNA_1450 (.A(net858));
 sg13g2_antennanp ANTENNA_1451 (.A(net858));
 sg13g2_antennanp ANTENNA_1452 (.A(net858));
 sg13g2_antennanp ANTENNA_1453 (.A(net858));
 sg13g2_antennanp ANTENNA_1454 (.A(net858));
 sg13g2_antennanp ANTENNA_1455 (.A(net858));
 sg13g2_antennanp ANTENNA_1456 (.A(net858));
 sg13g2_antennanp ANTENNA_1457 (.A(net858));
 sg13g2_antennanp ANTENNA_1458 (.A(net860));
 sg13g2_antennanp ANTENNA_1459 (.A(net860));
 sg13g2_antennanp ANTENNA_1460 (.A(net860));
 sg13g2_antennanp ANTENNA_1461 (.A(net860));
 sg13g2_antennanp ANTENNA_1462 (.A(net860));
 sg13g2_antennanp ANTENNA_1463 (.A(net860));
 sg13g2_antennanp ANTENNA_1464 (.A(net860));
 sg13g2_antennanp ANTENNA_1465 (.A(net860));
 sg13g2_antennanp ANTENNA_1466 (.A(net872));
 sg13g2_antennanp ANTENNA_1467 (.A(net872));
 sg13g2_antennanp ANTENNA_1468 (.A(net872));
 sg13g2_antennanp ANTENNA_1469 (.A(net872));
 sg13g2_antennanp ANTENNA_1470 (.A(net872));
 sg13g2_antennanp ANTENNA_1471 (.A(net872));
 sg13g2_antennanp ANTENNA_1472 (.A(net872));
 sg13g2_antennanp ANTENNA_1473 (.A(net872));
 sg13g2_antennanp ANTENNA_1474 (.A(net872));
 sg13g2_antennanp ANTENNA_1475 (.A(net872));
 sg13g2_antennanp ANTENNA_1476 (.A(net872));
 sg13g2_antennanp ANTENNA_1477 (.A(net872));
 sg13g2_antennanp ANTENNA_1478 (.A(net872));
 sg13g2_antennanp ANTENNA_1479 (.A(net872));
 sg13g2_antennanp ANTENNA_1480 (.A(net872));
 sg13g2_antennanp ANTENNA_1481 (.A(net872));
 sg13g2_antennanp ANTENNA_1482 (.A(net872));
 sg13g2_antennanp ANTENNA_1483 (.A(net872));
 sg13g2_antennanp ANTENNA_1484 (.A(net872));
 sg13g2_antennanp ANTENNA_1485 (.A(net872));
 sg13g2_antennanp ANTENNA_1486 (.A(net872));
 sg13g2_antennanp ANTENNA_1487 (.A(net872));
 sg13g2_antennanp ANTENNA_1488 (.A(net872));
 sg13g2_antennanp ANTENNA_1489 (.A(net872));
 sg13g2_antennanp ANTENNA_1490 (.A(net923));
 sg13g2_antennanp ANTENNA_1491 (.A(net923));
 sg13g2_antennanp ANTENNA_1492 (.A(net923));
 sg13g2_antennanp ANTENNA_1493 (.A(net923));
 sg13g2_antennanp ANTENNA_1494 (.A(net923));
 sg13g2_antennanp ANTENNA_1495 (.A(net923));
 sg13g2_antennanp ANTENNA_1496 (.A(net923));
 sg13g2_antennanp ANTENNA_1497 (.A(net923));
 sg13g2_antennanp ANTENNA_1498 (.A(net923));
 sg13g2_antennanp ANTENNA_1499 (.A(net928));
 sg13g2_antennanp ANTENNA_1500 (.A(net928));
 sg13g2_antennanp ANTENNA_1501 (.A(net928));
 sg13g2_antennanp ANTENNA_1502 (.A(net928));
 sg13g2_antennanp ANTENNA_1503 (.A(net928));
 sg13g2_antennanp ANTENNA_1504 (.A(net928));
 sg13g2_antennanp ANTENNA_1505 (.A(net928));
 sg13g2_antennanp ANTENNA_1506 (.A(net928));
 sg13g2_antennanp ANTENNA_1507 (.A(net928));
 sg13g2_antennanp ANTENNA_1508 (.A(net928));
 sg13g2_antennanp ANTENNA_1509 (.A(net928));
 sg13g2_antennanp ANTENNA_1510 (.A(net928));
 sg13g2_antennanp ANTENNA_1511 (.A(net928));
 sg13g2_antennanp ANTENNA_1512 (.A(net928));
 sg13g2_antennanp ANTENNA_1513 (.A(net928));
 sg13g2_antennanp ANTENNA_1514 (.A(net928));
 sg13g2_antennanp ANTENNA_1515 (.A(net995));
 sg13g2_antennanp ANTENNA_1516 (.A(net995));
 sg13g2_antennanp ANTENNA_1517 (.A(net995));
 sg13g2_antennanp ANTENNA_1518 (.A(net995));
 sg13g2_antennanp ANTENNA_1519 (.A(net995));
 sg13g2_antennanp ANTENNA_1520 (.A(net995));
 sg13g2_antennanp ANTENNA_1521 (.A(net995));
 sg13g2_antennanp ANTENNA_1522 (.A(net995));
 sg13g2_antennanp ANTENNA_1523 (.A(net995));
 sg13g2_antennanp ANTENNA_1524 (.A(net995));
 sg13g2_antennanp ANTENNA_1525 (.A(net995));
 sg13g2_antennanp ANTENNA_1526 (.A(net995));
 sg13g2_antennanp ANTENNA_1527 (.A(net995));
 sg13g2_antennanp ANTENNA_1528 (.A(net995));
 sg13g2_antennanp ANTENNA_1529 (.A(net995));
 sg13g2_antennanp ANTENNA_1530 (.A(net999));
 sg13g2_antennanp ANTENNA_1531 (.A(net999));
 sg13g2_antennanp ANTENNA_1532 (.A(net999));
 sg13g2_antennanp ANTENNA_1533 (.A(net999));
 sg13g2_antennanp ANTENNA_1534 (.A(net999));
 sg13g2_antennanp ANTENNA_1535 (.A(net999));
 sg13g2_antennanp ANTENNA_1536 (.A(net999));
 sg13g2_antennanp ANTENNA_1537 (.A(net999));
 sg13g2_antennanp ANTENNA_1538 (.A(net999));
 sg13g2_antennanp ANTENNA_1539 (.A(net1002));
 sg13g2_antennanp ANTENNA_1540 (.A(net1002));
 sg13g2_antennanp ANTENNA_1541 (.A(net1002));
 sg13g2_antennanp ANTENNA_1542 (.A(net1002));
 sg13g2_antennanp ANTENNA_1543 (.A(net1002));
 sg13g2_antennanp ANTENNA_1544 (.A(net1002));
 sg13g2_antennanp ANTENNA_1545 (.A(net1002));
 sg13g2_antennanp ANTENNA_1546 (.A(net1002));
 sg13g2_antennanp ANTENNA_1547 (.A(net1002));
 sg13g2_antennanp ANTENNA_1548 (.A(net1002));
 sg13g2_antennanp ANTENNA_1549 (.A(net1002));
 sg13g2_antennanp ANTENNA_1550 (.A(net1002));
 sg13g2_antennanp ANTENNA_1551 (.A(net1002));
 sg13g2_antennanp ANTENNA_1552 (.A(net1002));
 sg13g2_antennanp ANTENNA_1553 (.A(net1002));
 sg13g2_antennanp ANTENNA_1554 (.A(net1002));
 sg13g2_antennanp ANTENNA_1555 (.A(net1002));
 sg13g2_antennanp ANTENNA_1556 (.A(net1002));
 sg13g2_antennanp ANTENNA_1557 (.A(net1002));
 sg13g2_antennanp ANTENNA_1558 (.A(net1002));
 sg13g2_antennanp ANTENNA_1559 (.A(net1004));
 sg13g2_antennanp ANTENNA_1560 (.A(net1004));
 sg13g2_antennanp ANTENNA_1561 (.A(net1004));
 sg13g2_antennanp ANTENNA_1562 (.A(net1004));
 sg13g2_antennanp ANTENNA_1563 (.A(net1004));
 sg13g2_antennanp ANTENNA_1564 (.A(net1004));
 sg13g2_antennanp ANTENNA_1565 (.A(net1004));
 sg13g2_antennanp ANTENNA_1566 (.A(net1004));
 sg13g2_antennanp ANTENNA_1567 (.A(net1004));
 sg13g2_antennanp ANTENNA_1568 (.A(net1099));
 sg13g2_antennanp ANTENNA_1569 (.A(net1099));
 sg13g2_antennanp ANTENNA_1570 (.A(net1099));
 sg13g2_antennanp ANTENNA_1571 (.A(net1099));
 sg13g2_antennanp ANTENNA_1572 (.A(net1099));
 sg13g2_antennanp ANTENNA_1573 (.A(net1099));
 sg13g2_antennanp ANTENNA_1574 (.A(net1099));
 sg13g2_antennanp ANTENNA_1575 (.A(net1099));
 sg13g2_antennanp ANTENNA_1576 (.A(net1099));
 sg13g2_antennanp ANTENNA_1577 (.A(net1099));
 sg13g2_antennanp ANTENNA_1578 (.A(net1099));
 sg13g2_antennanp ANTENNA_1579 (.A(net1099));
 sg13g2_antennanp ANTENNA_1580 (.A(net1099));
 sg13g2_antennanp ANTENNA_1581 (.A(net1099));
 sg13g2_antennanp ANTENNA_1582 (.A(net1099));
 sg13g2_antennanp ANTENNA_1583 (.A(net1099));
 sg13g2_antennanp ANTENNA_1584 (.A(net1099));
 sg13g2_antennanp ANTENNA_1585 (.A(net1099));
 sg13g2_antennanp ANTENNA_1586 (.A(net1099));
 sg13g2_antennanp ANTENNA_1587 (.A(net1099));
 sg13g2_antennanp ANTENNA_1588 (.A(_00207_));
 sg13g2_antennanp ANTENNA_1589 (.A(_00785_));
 sg13g2_antennanp ANTENNA_1590 (.A(_00977_));
 sg13g2_antennanp ANTENNA_1591 (.A(_00977_));
 sg13g2_antennanp ANTENNA_1592 (.A(_01032_));
 sg13g2_antennanp ANTENNA_1593 (.A(_01047_));
 sg13g2_antennanp ANTENNA_1594 (.A(_01048_));
 sg13g2_antennanp ANTENNA_1595 (.A(_02836_));
 sg13g2_antennanp ANTENNA_1596 (.A(_02836_));
 sg13g2_antennanp ANTENNA_1597 (.A(_02836_));
 sg13g2_antennanp ANTENNA_1598 (.A(_02836_));
 sg13g2_antennanp ANTENNA_1599 (.A(_02845_));
 sg13g2_antennanp ANTENNA_1600 (.A(_02845_));
 sg13g2_antennanp ANTENNA_1601 (.A(_02845_));
 sg13g2_antennanp ANTENNA_1602 (.A(_02845_));
 sg13g2_antennanp ANTENNA_1603 (.A(_02845_));
 sg13g2_antennanp ANTENNA_1604 (.A(_02845_));
 sg13g2_antennanp ANTENNA_1605 (.A(_02845_));
 sg13g2_antennanp ANTENNA_1606 (.A(_02845_));
 sg13g2_antennanp ANTENNA_1607 (.A(_02845_));
 sg13g2_antennanp ANTENNA_1608 (.A(_02849_));
 sg13g2_antennanp ANTENNA_1609 (.A(_02849_));
 sg13g2_antennanp ANTENNA_1610 (.A(_02849_));
 sg13g2_antennanp ANTENNA_1611 (.A(_02849_));
 sg13g2_antennanp ANTENNA_1612 (.A(_02849_));
 sg13g2_antennanp ANTENNA_1613 (.A(_02849_));
 sg13g2_antennanp ANTENNA_1614 (.A(_02849_));
 sg13g2_antennanp ANTENNA_1615 (.A(_02849_));
 sg13g2_antennanp ANTENNA_1616 (.A(_02849_));
 sg13g2_antennanp ANTENNA_1617 (.A(_02861_));
 sg13g2_antennanp ANTENNA_1618 (.A(_02861_));
 sg13g2_antennanp ANTENNA_1619 (.A(_02861_));
 sg13g2_antennanp ANTENNA_1620 (.A(_02861_));
 sg13g2_antennanp ANTENNA_1621 (.A(_02976_));
 sg13g2_antennanp ANTENNA_1622 (.A(_02976_));
 sg13g2_antennanp ANTENNA_1623 (.A(_02976_));
 sg13g2_antennanp ANTENNA_1624 (.A(_02976_));
 sg13g2_antennanp ANTENNA_1625 (.A(_02976_));
 sg13g2_antennanp ANTENNA_1626 (.A(_02976_));
 sg13g2_antennanp ANTENNA_1627 (.A(_02976_));
 sg13g2_antennanp ANTENNA_1628 (.A(_02976_));
 sg13g2_antennanp ANTENNA_1629 (.A(_02976_));
 sg13g2_antennanp ANTENNA_1630 (.A(_03081_));
 sg13g2_antennanp ANTENNA_1631 (.A(_03148_));
 sg13g2_antennanp ANTENNA_1632 (.A(_03148_));
 sg13g2_antennanp ANTENNA_1633 (.A(_03507_));
 sg13g2_antennanp ANTENNA_1634 (.A(_03507_));
 sg13g2_antennanp ANTENNA_1635 (.A(_03507_));
 sg13g2_antennanp ANTENNA_1636 (.A(_03507_));
 sg13g2_antennanp ANTENNA_1637 (.A(_03507_));
 sg13g2_antennanp ANTENNA_1638 (.A(_03507_));
 sg13g2_antennanp ANTENNA_1639 (.A(_03513_));
 sg13g2_antennanp ANTENNA_1640 (.A(_03513_));
 sg13g2_antennanp ANTENNA_1641 (.A(_03513_));
 sg13g2_antennanp ANTENNA_1642 (.A(_03513_));
 sg13g2_antennanp ANTENNA_1643 (.A(_03513_));
 sg13g2_antennanp ANTENNA_1644 (.A(_03513_));
 sg13g2_antennanp ANTENNA_1645 (.A(_03513_));
 sg13g2_antennanp ANTENNA_1646 (.A(_03513_));
 sg13g2_antennanp ANTENNA_1647 (.A(_03513_));
 sg13g2_antennanp ANTENNA_1648 (.A(_03513_));
 sg13g2_antennanp ANTENNA_1649 (.A(_03513_));
 sg13g2_antennanp ANTENNA_1650 (.A(_03513_));
 sg13g2_antennanp ANTENNA_1651 (.A(_03513_));
 sg13g2_antennanp ANTENNA_1652 (.A(_03513_));
 sg13g2_antennanp ANTENNA_1653 (.A(_03539_));
 sg13g2_antennanp ANTENNA_1654 (.A(_03539_));
 sg13g2_antennanp ANTENNA_1655 (.A(_03539_));
 sg13g2_antennanp ANTENNA_1656 (.A(_03539_));
 sg13g2_antennanp ANTENNA_1657 (.A(_03539_));
 sg13g2_antennanp ANTENNA_1658 (.A(_03539_));
 sg13g2_antennanp ANTENNA_1659 (.A(_03539_));
 sg13g2_antennanp ANTENNA_1660 (.A(_03539_));
 sg13g2_antennanp ANTENNA_1661 (.A(_03539_));
 sg13g2_antennanp ANTENNA_1662 (.A(_03824_));
 sg13g2_antennanp ANTENNA_1663 (.A(_03838_));
 sg13g2_antennanp ANTENNA_1664 (.A(_03838_));
 sg13g2_antennanp ANTENNA_1665 (.A(_03838_));
 sg13g2_antennanp ANTENNA_1666 (.A(_03838_));
 sg13g2_antennanp ANTENNA_1667 (.A(_03838_));
 sg13g2_antennanp ANTENNA_1668 (.A(_03838_));
 sg13g2_antennanp ANTENNA_1669 (.A(_04855_));
 sg13g2_antennanp ANTENNA_1670 (.A(_04980_));
 sg13g2_antennanp ANTENNA_1671 (.A(_04980_));
 sg13g2_antennanp ANTENNA_1672 (.A(_04980_));
 sg13g2_antennanp ANTENNA_1673 (.A(_04980_));
 sg13g2_antennanp ANTENNA_1674 (.A(_05006_));
 sg13g2_antennanp ANTENNA_1675 (.A(_05157_));
 sg13g2_antennanp ANTENNA_1676 (.A(_05229_));
 sg13g2_antennanp ANTENNA_1677 (.A(_05260_));
 sg13g2_antennanp ANTENNA_1678 (.A(_05270_));
 sg13g2_antennanp ANTENNA_1679 (.A(_05287_));
 sg13g2_antennanp ANTENNA_1680 (.A(_05303_));
 sg13g2_antennanp ANTENNA_1681 (.A(_05307_));
 sg13g2_antennanp ANTENNA_1682 (.A(_05314_));
 sg13g2_antennanp ANTENNA_1683 (.A(_05464_));
 sg13g2_antennanp ANTENNA_1684 (.A(_05525_));
 sg13g2_antennanp ANTENNA_1685 (.A(_05529_));
 sg13g2_antennanp ANTENNA_1686 (.A(_05607_));
 sg13g2_antennanp ANTENNA_1687 (.A(_05676_));
 sg13g2_antennanp ANTENNA_1688 (.A(_05756_));
 sg13g2_antennanp ANTENNA_1689 (.A(_05756_));
 sg13g2_antennanp ANTENNA_1690 (.A(_05770_));
 sg13g2_antennanp ANTENNA_1691 (.A(_05780_));
 sg13g2_antennanp ANTENNA_1692 (.A(_05780_));
 sg13g2_antennanp ANTENNA_1693 (.A(_05780_));
 sg13g2_antennanp ANTENNA_1694 (.A(_05780_));
 sg13g2_antennanp ANTENNA_1695 (.A(_05796_));
 sg13g2_antennanp ANTENNA_1696 (.A(_06579_));
 sg13g2_antennanp ANTENNA_1697 (.A(_06579_));
 sg13g2_antennanp ANTENNA_1698 (.A(_06579_));
 sg13g2_antennanp ANTENNA_1699 (.A(_06579_));
 sg13g2_antennanp ANTENNA_1700 (.A(_06579_));
 sg13g2_antennanp ANTENNA_1701 (.A(_06579_));
 sg13g2_antennanp ANTENNA_1702 (.A(_06579_));
 sg13g2_antennanp ANTENNA_1703 (.A(_06579_));
 sg13g2_antennanp ANTENNA_1704 (.A(_06579_));
 sg13g2_antennanp ANTENNA_1705 (.A(_06582_));
 sg13g2_antennanp ANTENNA_1706 (.A(_06582_));
 sg13g2_antennanp ANTENNA_1707 (.A(_06582_));
 sg13g2_antennanp ANTENNA_1708 (.A(_06582_));
 sg13g2_antennanp ANTENNA_1709 (.A(_06885_));
 sg13g2_antennanp ANTENNA_1710 (.A(_06885_));
 sg13g2_antennanp ANTENNA_1711 (.A(_06885_));
 sg13g2_antennanp ANTENNA_1712 (.A(_06885_));
 sg13g2_antennanp ANTENNA_1713 (.A(_06885_));
 sg13g2_antennanp ANTENNA_1714 (.A(_06885_));
 sg13g2_antennanp ANTENNA_1715 (.A(_06885_));
 sg13g2_antennanp ANTENNA_1716 (.A(_06885_));
 sg13g2_antennanp ANTENNA_1717 (.A(_06885_));
 sg13g2_antennanp ANTENNA_1718 (.A(_06885_));
 sg13g2_antennanp ANTENNA_1719 (.A(_07626_));
 sg13g2_antennanp ANTENNA_1720 (.A(_07632_));
 sg13g2_antennanp ANTENNA_1721 (.A(_07634_));
 sg13g2_antennanp ANTENNA_1722 (.A(_07851_));
 sg13g2_antennanp ANTENNA_1723 (.A(_07851_));
 sg13g2_antennanp ANTENNA_1724 (.A(_07851_));
 sg13g2_antennanp ANTENNA_1725 (.A(_07851_));
 sg13g2_antennanp ANTENNA_1726 (.A(_07851_));
 sg13g2_antennanp ANTENNA_1727 (.A(_07851_));
 sg13g2_antennanp ANTENNA_1728 (.A(_07851_));
 sg13g2_antennanp ANTENNA_1729 (.A(_07851_));
 sg13g2_antennanp ANTENNA_1730 (.A(_07851_));
 sg13g2_antennanp ANTENNA_1731 (.A(_07851_));
 sg13g2_antennanp ANTENNA_1732 (.A(_08260_));
 sg13g2_antennanp ANTENNA_1733 (.A(_08260_));
 sg13g2_antennanp ANTENNA_1734 (.A(_08260_));
 sg13g2_antennanp ANTENNA_1735 (.A(_08346_));
 sg13g2_antennanp ANTENNA_1736 (.A(_08346_));
 sg13g2_antennanp ANTENNA_1737 (.A(_08346_));
 sg13g2_antennanp ANTENNA_1738 (.A(_08346_));
 sg13g2_antennanp ANTENNA_1739 (.A(_08346_));
 sg13g2_antennanp ANTENNA_1740 (.A(_08346_));
 sg13g2_antennanp ANTENNA_1741 (.A(_08346_));
 sg13g2_antennanp ANTENNA_1742 (.A(_08346_));
 sg13g2_antennanp ANTENNA_1743 (.A(_08455_));
 sg13g2_antennanp ANTENNA_1744 (.A(_08455_));
 sg13g2_antennanp ANTENNA_1745 (.A(_08455_));
 sg13g2_antennanp ANTENNA_1746 (.A(_08497_));
 sg13g2_antennanp ANTENNA_1747 (.A(_08497_));
 sg13g2_antennanp ANTENNA_1748 (.A(_08497_));
 sg13g2_antennanp ANTENNA_1749 (.A(_08565_));
 sg13g2_antennanp ANTENNA_1750 (.A(_08565_));
 sg13g2_antennanp ANTENNA_1751 (.A(_08565_));
 sg13g2_antennanp ANTENNA_1752 (.A(_08565_));
 sg13g2_antennanp ANTENNA_1753 (.A(_08565_));
 sg13g2_antennanp ANTENNA_1754 (.A(_08565_));
 sg13g2_antennanp ANTENNA_1755 (.A(_08603_));
 sg13g2_antennanp ANTENNA_1756 (.A(_08603_));
 sg13g2_antennanp ANTENNA_1757 (.A(_08603_));
 sg13g2_antennanp ANTENNA_1758 (.A(_08603_));
 sg13g2_antennanp ANTENNA_1759 (.A(_08603_));
 sg13g2_antennanp ANTENNA_1760 (.A(_08603_));
 sg13g2_antennanp ANTENNA_1761 (.A(_08633_));
 sg13g2_antennanp ANTENNA_1762 (.A(_08663_));
 sg13g2_antennanp ANTENNA_1763 (.A(_08663_));
 sg13g2_antennanp ANTENNA_1764 (.A(_08663_));
 sg13g2_antennanp ANTENNA_1765 (.A(_08663_));
 sg13g2_antennanp ANTENNA_1766 (.A(_08663_));
 sg13g2_antennanp ANTENNA_1767 (.A(_08663_));
 sg13g2_antennanp ANTENNA_1768 (.A(_08799_));
 sg13g2_antennanp ANTENNA_1769 (.A(_08799_));
 sg13g2_antennanp ANTENNA_1770 (.A(_08799_));
 sg13g2_antennanp ANTENNA_1771 (.A(_08799_));
 sg13g2_antennanp ANTENNA_1772 (.A(_08799_));
 sg13g2_antennanp ANTENNA_1773 (.A(_08799_));
 sg13g2_antennanp ANTENNA_1774 (.A(_08820_));
 sg13g2_antennanp ANTENNA_1775 (.A(_08820_));
 sg13g2_antennanp ANTENNA_1776 (.A(_08820_));
 sg13g2_antennanp ANTENNA_1777 (.A(_08826_));
 sg13g2_antennanp ANTENNA_1778 (.A(_08826_));
 sg13g2_antennanp ANTENNA_1779 (.A(_08826_));
 sg13g2_antennanp ANTENNA_1780 (.A(_08826_));
 sg13g2_antennanp ANTENNA_1781 (.A(_08826_));
 sg13g2_antennanp ANTENNA_1782 (.A(_08826_));
 sg13g2_antennanp ANTENNA_1783 (.A(_08848_));
 sg13g2_antennanp ANTENNA_1784 (.A(_08848_));
 sg13g2_antennanp ANTENNA_1785 (.A(_08848_));
 sg13g2_antennanp ANTENNA_1786 (.A(_08868_));
 sg13g2_antennanp ANTENNA_1787 (.A(_08900_));
 sg13g2_antennanp ANTENNA_1788 (.A(_08900_));
 sg13g2_antennanp ANTENNA_1789 (.A(_08900_));
 sg13g2_antennanp ANTENNA_1790 (.A(_08950_));
 sg13g2_antennanp ANTENNA_1791 (.A(_08950_));
 sg13g2_antennanp ANTENNA_1792 (.A(_08950_));
 sg13g2_antennanp ANTENNA_1793 (.A(_08950_));
 sg13g2_antennanp ANTENNA_1794 (.A(_08950_));
 sg13g2_antennanp ANTENNA_1795 (.A(_08950_));
 sg13g2_antennanp ANTENNA_1796 (.A(_08950_));
 sg13g2_antennanp ANTENNA_1797 (.A(_08950_));
 sg13g2_antennanp ANTENNA_1798 (.A(_08950_));
 sg13g2_antennanp ANTENNA_1799 (.A(_08970_));
 sg13g2_antennanp ANTENNA_1800 (.A(_08970_));
 sg13g2_antennanp ANTENNA_1801 (.A(_08986_));
 sg13g2_antennanp ANTENNA_1802 (.A(_08986_));
 sg13g2_antennanp ANTENNA_1803 (.A(_09002_));
 sg13g2_antennanp ANTENNA_1804 (.A(_09002_));
 sg13g2_antennanp ANTENNA_1805 (.A(_09065_));
 sg13g2_antennanp ANTENNA_1806 (.A(_09065_));
 sg13g2_antennanp ANTENNA_1807 (.A(_09091_));
 sg13g2_antennanp ANTENNA_1808 (.A(_09091_));
 sg13g2_antennanp ANTENNA_1809 (.A(_09091_));
 sg13g2_antennanp ANTENNA_1810 (.A(_09120_));
 sg13g2_antennanp ANTENNA_1811 (.A(_09120_));
 sg13g2_antennanp ANTENNA_1812 (.A(_09158_));
 sg13g2_antennanp ANTENNA_1813 (.A(_09158_));
 sg13g2_antennanp ANTENNA_1814 (.A(_09158_));
 sg13g2_antennanp ANTENNA_1815 (.A(_09173_));
 sg13g2_antennanp ANTENNA_1816 (.A(_09211_));
 sg13g2_antennanp ANTENNA_1817 (.A(_09211_));
 sg13g2_antennanp ANTENNA_1818 (.A(_09211_));
 sg13g2_antennanp ANTENNA_1819 (.A(_09211_));
 sg13g2_antennanp ANTENNA_1820 (.A(_09211_));
 sg13g2_antennanp ANTENNA_1821 (.A(_09218_));
 sg13g2_antennanp ANTENNA_1822 (.A(_09220_));
 sg13g2_antennanp ANTENNA_1823 (.A(_09220_));
 sg13g2_antennanp ANTENNA_1824 (.A(_09220_));
 sg13g2_antennanp ANTENNA_1825 (.A(_09220_));
 sg13g2_antennanp ANTENNA_1826 (.A(_09220_));
 sg13g2_antennanp ANTENNA_1827 (.A(_09220_));
 sg13g2_antennanp ANTENNA_1828 (.A(_09220_));
 sg13g2_antennanp ANTENNA_1829 (.A(_09220_));
 sg13g2_antennanp ANTENNA_1830 (.A(_09220_));
 sg13g2_antennanp ANTENNA_1831 (.A(_09220_));
 sg13g2_antennanp ANTENNA_1832 (.A(_09220_));
 sg13g2_antennanp ANTENNA_1833 (.A(_09220_));
 sg13g2_antennanp ANTENNA_1834 (.A(_09220_));
 sg13g2_antennanp ANTENNA_1835 (.A(_09298_));
 sg13g2_antennanp ANTENNA_1836 (.A(_09298_));
 sg13g2_antennanp ANTENNA_1837 (.A(_09298_));
 sg13g2_antennanp ANTENNA_1838 (.A(_09318_));
 sg13g2_antennanp ANTENNA_1839 (.A(_09318_));
 sg13g2_antennanp ANTENNA_1840 (.A(_09318_));
 sg13g2_antennanp ANTENNA_1841 (.A(_09394_));
 sg13g2_antennanp ANTENNA_1842 (.A(_09396_));
 sg13g2_antennanp ANTENNA_1843 (.A(_09447_));
 sg13g2_antennanp ANTENNA_1844 (.A(_09448_));
 sg13g2_antennanp ANTENNA_1845 (.A(_09448_));
 sg13g2_antennanp ANTENNA_1846 (.A(_09448_));
 sg13g2_antennanp ANTENNA_1847 (.A(_09448_));
 sg13g2_antennanp ANTENNA_1848 (.A(_09450_));
 sg13g2_antennanp ANTENNA_1849 (.A(_09492_));
 sg13g2_antennanp ANTENNA_1850 (.A(_09521_));
 sg13g2_antennanp ANTENNA_1851 (.A(_09544_));
 sg13g2_antennanp ANTENNA_1852 (.A(_09657_));
 sg13g2_antennanp ANTENNA_1853 (.A(_09722_));
 sg13g2_antennanp ANTENNA_1854 (.A(_09769_));
 sg13g2_antennanp ANTENNA_1855 (.A(_09791_));
 sg13g2_antennanp ANTENNA_1856 (.A(_09852_));
 sg13g2_antennanp ANTENNA_1857 (.A(_09852_));
 sg13g2_antennanp ANTENNA_1858 (.A(_09852_));
 sg13g2_antennanp ANTENNA_1859 (.A(_09852_));
 sg13g2_antennanp ANTENNA_1860 (.A(_09852_));
 sg13g2_antennanp ANTENNA_1861 (.A(_09852_));
 sg13g2_antennanp ANTENNA_1862 (.A(_09852_));
 sg13g2_antennanp ANTENNA_1863 (.A(_09852_));
 sg13g2_antennanp ANTENNA_1864 (.A(_09852_));
 sg13g2_antennanp ANTENNA_1865 (.A(_09852_));
 sg13g2_antennanp ANTENNA_1866 (.A(_09852_));
 sg13g2_antennanp ANTENNA_1867 (.A(_09852_));
 sg13g2_antennanp ANTENNA_1868 (.A(_09852_));
 sg13g2_antennanp ANTENNA_1869 (.A(_09852_));
 sg13g2_antennanp ANTENNA_1870 (.A(_09852_));
 sg13g2_antennanp ANTENNA_1871 (.A(_09852_));
 sg13g2_antennanp ANTENNA_1872 (.A(_09852_));
 sg13g2_antennanp ANTENNA_1873 (.A(_10042_));
 sg13g2_antennanp ANTENNA_1874 (.A(_10042_));
 sg13g2_antennanp ANTENNA_1875 (.A(_10042_));
 sg13g2_antennanp ANTENNA_1876 (.A(_10146_));
 sg13g2_antennanp ANTENNA_1877 (.A(_10146_));
 sg13g2_antennanp ANTENNA_1878 (.A(_10146_));
 sg13g2_antennanp ANTENNA_1879 (.A(_10146_));
 sg13g2_antennanp ANTENNA_1880 (.A(_10146_));
 sg13g2_antennanp ANTENNA_1881 (.A(_10146_));
 sg13g2_antennanp ANTENNA_1882 (.A(_10146_));
 sg13g2_antennanp ANTENNA_1883 (.A(_10146_));
 sg13g2_antennanp ANTENNA_1884 (.A(_10162_));
 sg13g2_antennanp ANTENNA_1885 (.A(_10162_));
 sg13g2_antennanp ANTENNA_1886 (.A(_10162_));
 sg13g2_antennanp ANTENNA_1887 (.A(_10162_));
 sg13g2_antennanp ANTENNA_1888 (.A(_10162_));
 sg13g2_antennanp ANTENNA_1889 (.A(_10162_));
 sg13g2_antennanp ANTENNA_1890 (.A(_10162_));
 sg13g2_antennanp ANTENNA_1891 (.A(_10162_));
 sg13g2_antennanp ANTENNA_1892 (.A(_10379_));
 sg13g2_antennanp ANTENNA_1893 (.A(_10379_));
 sg13g2_antennanp ANTENNA_1894 (.A(_10379_));
 sg13g2_antennanp ANTENNA_1895 (.A(_10642_));
 sg13g2_antennanp ANTENNA_1896 (.A(_10642_));
 sg13g2_antennanp ANTENNA_1897 (.A(_10642_));
 sg13g2_antennanp ANTENNA_1898 (.A(_10642_));
 sg13g2_antennanp ANTENNA_1899 (.A(_10642_));
 sg13g2_antennanp ANTENNA_1900 (.A(_10642_));
 sg13g2_antennanp ANTENNA_1901 (.A(_10642_));
 sg13g2_antennanp ANTENNA_1902 (.A(_10744_));
 sg13g2_antennanp ANTENNA_1903 (.A(_10744_));
 sg13g2_antennanp ANTENNA_1904 (.A(_10744_));
 sg13g2_antennanp ANTENNA_1905 (.A(_10744_));
 sg13g2_antennanp ANTENNA_1906 (.A(_12205_));
 sg13g2_antennanp ANTENNA_1907 (.A(_12205_));
 sg13g2_antennanp ANTENNA_1908 (.A(_12205_));
 sg13g2_antennanp ANTENNA_1909 (.A(_12205_));
 sg13g2_antennanp ANTENNA_1910 (.A(_12205_));
 sg13g2_antennanp ANTENNA_1911 (.A(_12205_));
 sg13g2_antennanp ANTENNA_1912 (.A(_12205_));
 sg13g2_antennanp ANTENNA_1913 (.A(_12205_));
 sg13g2_antennanp ANTENNA_1914 (.A(_12205_));
 sg13g2_antennanp ANTENNA_1915 (.A(_12218_));
 sg13g2_antennanp ANTENNA_1916 (.A(_12218_));
 sg13g2_antennanp ANTENNA_1917 (.A(_12218_));
 sg13g2_antennanp ANTENNA_1918 (.A(_12218_));
 sg13g2_antennanp ANTENNA_1919 (.A(_12218_));
 sg13g2_antennanp ANTENNA_1920 (.A(_12218_));
 sg13g2_antennanp ANTENNA_1921 (.A(_12218_));
 sg13g2_antennanp ANTENNA_1922 (.A(_12218_));
 sg13g2_antennanp ANTENNA_1923 (.A(_12218_));
 sg13g2_antennanp ANTENNA_1924 (.A(_12225_));
 sg13g2_antennanp ANTENNA_1925 (.A(_12225_));
 sg13g2_antennanp ANTENNA_1926 (.A(_12225_));
 sg13g2_antennanp ANTENNA_1927 (.A(_12225_));
 sg13g2_antennanp ANTENNA_1928 (.A(_12225_));
 sg13g2_antennanp ANTENNA_1929 (.A(_12225_));
 sg13g2_antennanp ANTENNA_1930 (.A(_12225_));
 sg13g2_antennanp ANTENNA_1931 (.A(_12225_));
 sg13g2_antennanp ANTENNA_1932 (.A(_12225_));
 sg13g2_antennanp ANTENNA_1933 (.A(_12236_));
 sg13g2_antennanp ANTENNA_1934 (.A(_12236_));
 sg13g2_antennanp ANTENNA_1935 (.A(_12236_));
 sg13g2_antennanp ANTENNA_1936 (.A(_12236_));
 sg13g2_antennanp ANTENNA_1937 (.A(_12236_));
 sg13g2_antennanp ANTENNA_1938 (.A(_12236_));
 sg13g2_antennanp ANTENNA_1939 (.A(_12236_));
 sg13g2_antennanp ANTENNA_1940 (.A(_12236_));
 sg13g2_antennanp ANTENNA_1941 (.A(_12236_));
 sg13g2_antennanp ANTENNA_1942 (.A(\cpu.dcache.wdata[10] ));
 sg13g2_antennanp ANTENNA_1943 (.A(\cpu.dcache.wdata[10] ));
 sg13g2_antennanp ANTENNA_1944 (.A(\cpu.dcache.wdata[10] ));
 sg13g2_antennanp ANTENNA_1945 (.A(\cpu.dcache.wdata[10] ));
 sg13g2_antennanp ANTENNA_1946 (.A(\cpu.dcache.wdata[12] ));
 sg13g2_antennanp ANTENNA_1947 (.A(\cpu.dcache.wdata[12] ));
 sg13g2_antennanp ANTENNA_1948 (.A(\cpu.dcache.wdata[12] ));
 sg13g2_antennanp ANTENNA_1949 (.A(\cpu.dcache.wdata[12] ));
 sg13g2_antennanp ANTENNA_1950 (.A(\cpu.dcache.wdata[9] ));
 sg13g2_antennanp ANTENNA_1951 (.A(\cpu.dcache.wdata[9] ));
 sg13g2_antennanp ANTENNA_1952 (.A(\cpu.dcache.wdata[9] ));
 sg13g2_antennanp ANTENNA_1953 (.A(\cpu.dcache.wdata[9] ));
 sg13g2_antennanp ANTENNA_1954 (.A(\cpu.ex.pc[1] ));
 sg13g2_antennanp ANTENNA_1955 (.A(\cpu.ex.pc[2] ));
 sg13g2_antennanp ANTENNA_1956 (.A(\cpu.gpio.uart_rx ));
 sg13g2_antennanp ANTENNA_1957 (.A(\cpu.gpio.uart_rx ));
 sg13g2_antennanp ANTENNA_1958 (.A(\cpu.qspi.c_wstrobe_i ));
 sg13g2_antennanp ANTENNA_1959 (.A(\cpu.qspi.c_wstrobe_i ));
 sg13g2_antennanp ANTENNA_1960 (.A(net3));
 sg13g2_antennanp ANTENNA_1961 (.A(net3));
 sg13g2_antennanp ANTENNA_1962 (.A(net3));
 sg13g2_antennanp ANTENNA_1963 (.A(net11));
 sg13g2_antennanp ANTENNA_1964 (.A(net11));
 sg13g2_antennanp ANTENNA_1965 (.A(net11));
 sg13g2_antennanp ANTENNA_1966 (.A(net12));
 sg13g2_antennanp ANTENNA_1967 (.A(net12));
 sg13g2_antennanp ANTENNA_1968 (.A(net12));
 sg13g2_antennanp ANTENNA_1969 (.A(net13));
 sg13g2_antennanp ANTENNA_1970 (.A(net13));
 sg13g2_antennanp ANTENNA_1971 (.A(net13));
 sg13g2_antennanp ANTENNA_1972 (.A(net14));
 sg13g2_antennanp ANTENNA_1973 (.A(net14));
 sg13g2_antennanp ANTENNA_1974 (.A(net14));
 sg13g2_antennanp ANTENNA_1975 (.A(net114));
 sg13g2_antennanp ANTENNA_1976 (.A(net114));
 sg13g2_antennanp ANTENNA_1977 (.A(net114));
 sg13g2_antennanp ANTENNA_1978 (.A(net114));
 sg13g2_antennanp ANTENNA_1979 (.A(net114));
 sg13g2_antennanp ANTENNA_1980 (.A(net114));
 sg13g2_antennanp ANTENNA_1981 (.A(net114));
 sg13g2_antennanp ANTENNA_1982 (.A(net114));
 sg13g2_antennanp ANTENNA_1983 (.A(net114));
 sg13g2_antennanp ANTENNA_1984 (.A(net114));
 sg13g2_antennanp ANTENNA_1985 (.A(net114));
 sg13g2_antennanp ANTENNA_1986 (.A(net114));
 sg13g2_antennanp ANTENNA_1987 (.A(net114));
 sg13g2_antennanp ANTENNA_1988 (.A(net114));
 sg13g2_antennanp ANTENNA_1989 (.A(net114));
 sg13g2_antennanp ANTENNA_1990 (.A(net489));
 sg13g2_antennanp ANTENNA_1991 (.A(net489));
 sg13g2_antennanp ANTENNA_1992 (.A(net489));
 sg13g2_antennanp ANTENNA_1993 (.A(net489));
 sg13g2_antennanp ANTENNA_1994 (.A(net489));
 sg13g2_antennanp ANTENNA_1995 (.A(net489));
 sg13g2_antennanp ANTENNA_1996 (.A(net489));
 sg13g2_antennanp ANTENNA_1997 (.A(net489));
 sg13g2_antennanp ANTENNA_1998 (.A(net489));
 sg13g2_antennanp ANTENNA_1999 (.A(net491));
 sg13g2_antennanp ANTENNA_2000 (.A(net491));
 sg13g2_antennanp ANTENNA_2001 (.A(net491));
 sg13g2_antennanp ANTENNA_2002 (.A(net491));
 sg13g2_antennanp ANTENNA_2003 (.A(net491));
 sg13g2_antennanp ANTENNA_2004 (.A(net491));
 sg13g2_antennanp ANTENNA_2005 (.A(net491));
 sg13g2_antennanp ANTENNA_2006 (.A(net491));
 sg13g2_antennanp ANTENNA_2007 (.A(net617));
 sg13g2_antennanp ANTENNA_2008 (.A(net617));
 sg13g2_antennanp ANTENNA_2009 (.A(net617));
 sg13g2_antennanp ANTENNA_2010 (.A(net617));
 sg13g2_antennanp ANTENNA_2011 (.A(net617));
 sg13g2_antennanp ANTENNA_2012 (.A(net617));
 sg13g2_antennanp ANTENNA_2013 (.A(net617));
 sg13g2_antennanp ANTENNA_2014 (.A(net617));
 sg13g2_antennanp ANTENNA_2015 (.A(net617));
 sg13g2_antennanp ANTENNA_2016 (.A(net617));
 sg13g2_antennanp ANTENNA_2017 (.A(net617));
 sg13g2_antennanp ANTENNA_2018 (.A(net617));
 sg13g2_antennanp ANTENNA_2019 (.A(net617));
 sg13g2_antennanp ANTENNA_2020 (.A(net686));
 sg13g2_antennanp ANTENNA_2021 (.A(net686));
 sg13g2_antennanp ANTENNA_2022 (.A(net686));
 sg13g2_antennanp ANTENNA_2023 (.A(net686));
 sg13g2_antennanp ANTENNA_2024 (.A(net686));
 sg13g2_antennanp ANTENNA_2025 (.A(net686));
 sg13g2_antennanp ANTENNA_2026 (.A(net686));
 sg13g2_antennanp ANTENNA_2027 (.A(net686));
 sg13g2_antennanp ANTENNA_2028 (.A(net708));
 sg13g2_antennanp ANTENNA_2029 (.A(net708));
 sg13g2_antennanp ANTENNA_2030 (.A(net708));
 sg13g2_antennanp ANTENNA_2031 (.A(net708));
 sg13g2_antennanp ANTENNA_2032 (.A(net708));
 sg13g2_antennanp ANTENNA_2033 (.A(net708));
 sg13g2_antennanp ANTENNA_2034 (.A(net708));
 sg13g2_antennanp ANTENNA_2035 (.A(net708));
 sg13g2_antennanp ANTENNA_2036 (.A(net745));
 sg13g2_antennanp ANTENNA_2037 (.A(net745));
 sg13g2_antennanp ANTENNA_2038 (.A(net745));
 sg13g2_antennanp ANTENNA_2039 (.A(net745));
 sg13g2_antennanp ANTENNA_2040 (.A(net745));
 sg13g2_antennanp ANTENNA_2041 (.A(net745));
 sg13g2_antennanp ANTENNA_2042 (.A(net745));
 sg13g2_antennanp ANTENNA_2043 (.A(net745));
 sg13g2_antennanp ANTENNA_2044 (.A(net803));
 sg13g2_antennanp ANTENNA_2045 (.A(net803));
 sg13g2_antennanp ANTENNA_2046 (.A(net803));
 sg13g2_antennanp ANTENNA_2047 (.A(net803));
 sg13g2_antennanp ANTENNA_2048 (.A(net803));
 sg13g2_antennanp ANTENNA_2049 (.A(net803));
 sg13g2_antennanp ANTENNA_2050 (.A(net803));
 sg13g2_antennanp ANTENNA_2051 (.A(net803));
 sg13g2_antennanp ANTENNA_2052 (.A(net858));
 sg13g2_antennanp ANTENNA_2053 (.A(net858));
 sg13g2_antennanp ANTENNA_2054 (.A(net858));
 sg13g2_antennanp ANTENNA_2055 (.A(net858));
 sg13g2_antennanp ANTENNA_2056 (.A(net858));
 sg13g2_antennanp ANTENNA_2057 (.A(net858));
 sg13g2_antennanp ANTENNA_2058 (.A(net858));
 sg13g2_antennanp ANTENNA_2059 (.A(net858));
 sg13g2_antennanp ANTENNA_2060 (.A(net858));
 sg13g2_antennanp ANTENNA_2061 (.A(net872));
 sg13g2_antennanp ANTENNA_2062 (.A(net872));
 sg13g2_antennanp ANTENNA_2063 (.A(net872));
 sg13g2_antennanp ANTENNA_2064 (.A(net872));
 sg13g2_antennanp ANTENNA_2065 (.A(net872));
 sg13g2_antennanp ANTENNA_2066 (.A(net872));
 sg13g2_antennanp ANTENNA_2067 (.A(net872));
 sg13g2_antennanp ANTENNA_2068 (.A(net872));
 sg13g2_antennanp ANTENNA_2069 (.A(net872));
 sg13g2_antennanp ANTENNA_2070 (.A(net872));
 sg13g2_antennanp ANTENNA_2071 (.A(net872));
 sg13g2_antennanp ANTENNA_2072 (.A(net872));
 sg13g2_antennanp ANTENNA_2073 (.A(net872));
 sg13g2_antennanp ANTENNA_2074 (.A(net872));
 sg13g2_antennanp ANTENNA_2075 (.A(net872));
 sg13g2_antennanp ANTENNA_2076 (.A(net872));
 sg13g2_antennanp ANTENNA_2077 (.A(net872));
 sg13g2_antennanp ANTENNA_2078 (.A(net872));
 sg13g2_antennanp ANTENNA_2079 (.A(net872));
 sg13g2_antennanp ANTENNA_2080 (.A(net872));
 sg13g2_antennanp ANTENNA_2081 (.A(net872));
 sg13g2_antennanp ANTENNA_2082 (.A(net872));
 sg13g2_antennanp ANTENNA_2083 (.A(net872));
 sg13g2_antennanp ANTENNA_2084 (.A(net872));
 sg13g2_antennanp ANTENNA_2085 (.A(net928));
 sg13g2_antennanp ANTENNA_2086 (.A(net928));
 sg13g2_antennanp ANTENNA_2087 (.A(net928));
 sg13g2_antennanp ANTENNA_2088 (.A(net928));
 sg13g2_antennanp ANTENNA_2089 (.A(net928));
 sg13g2_antennanp ANTENNA_2090 (.A(net928));
 sg13g2_antennanp ANTENNA_2091 (.A(net928));
 sg13g2_antennanp ANTENNA_2092 (.A(net928));
 sg13g2_antennanp ANTENNA_2093 (.A(net928));
 sg13g2_antennanp ANTENNA_2094 (.A(net995));
 sg13g2_antennanp ANTENNA_2095 (.A(net995));
 sg13g2_antennanp ANTENNA_2096 (.A(net995));
 sg13g2_antennanp ANTENNA_2097 (.A(net995));
 sg13g2_antennanp ANTENNA_2098 (.A(net995));
 sg13g2_antennanp ANTENNA_2099 (.A(net995));
 sg13g2_antennanp ANTENNA_2100 (.A(net995));
 sg13g2_antennanp ANTENNA_2101 (.A(net995));
 sg13g2_antennanp ANTENNA_2102 (.A(net995));
 sg13g2_antennanp ANTENNA_2103 (.A(net995));
 sg13g2_antennanp ANTENNA_2104 (.A(net995));
 sg13g2_antennanp ANTENNA_2105 (.A(net995));
 sg13g2_antennanp ANTENNA_2106 (.A(net995));
 sg13g2_antennanp ANTENNA_2107 (.A(net995));
 sg13g2_antennanp ANTENNA_2108 (.A(net995));
 sg13g2_antennanp ANTENNA_2109 (.A(net995));
 sg13g2_antennanp ANTENNA_2110 (.A(net995));
 sg13g2_antennanp ANTENNA_2111 (.A(net995));
 sg13g2_antennanp ANTENNA_2112 (.A(net999));
 sg13g2_antennanp ANTENNA_2113 (.A(net999));
 sg13g2_antennanp ANTENNA_2114 (.A(net999));
 sg13g2_antennanp ANTENNA_2115 (.A(net999));
 sg13g2_antennanp ANTENNA_2116 (.A(net999));
 sg13g2_antennanp ANTENNA_2117 (.A(net999));
 sg13g2_antennanp ANTENNA_2118 (.A(net999));
 sg13g2_antennanp ANTENNA_2119 (.A(net999));
 sg13g2_antennanp ANTENNA_2120 (.A(net1002));
 sg13g2_antennanp ANTENNA_2121 (.A(net1002));
 sg13g2_antennanp ANTENNA_2122 (.A(net1002));
 sg13g2_antennanp ANTENNA_2123 (.A(net1002));
 sg13g2_antennanp ANTENNA_2124 (.A(net1002));
 sg13g2_antennanp ANTENNA_2125 (.A(net1002));
 sg13g2_antennanp ANTENNA_2126 (.A(net1002));
 sg13g2_antennanp ANTENNA_2127 (.A(net1002));
 sg13g2_antennanp ANTENNA_2128 (.A(net1002));
 sg13g2_antennanp ANTENNA_2129 (.A(net1004));
 sg13g2_antennanp ANTENNA_2130 (.A(net1004));
 sg13g2_antennanp ANTENNA_2131 (.A(net1004));
 sg13g2_antennanp ANTENNA_2132 (.A(net1004));
 sg13g2_antennanp ANTENNA_2133 (.A(net1004));
 sg13g2_antennanp ANTENNA_2134 (.A(net1004));
 sg13g2_antennanp ANTENNA_2135 (.A(net1004));
 sg13g2_antennanp ANTENNA_2136 (.A(net1004));
 sg13g2_antennanp ANTENNA_2137 (.A(net1004));
 sg13g2_antennanp ANTENNA_2138 (.A(net1099));
 sg13g2_antennanp ANTENNA_2139 (.A(net1099));
 sg13g2_antennanp ANTENNA_2140 (.A(net1099));
 sg13g2_antennanp ANTENNA_2141 (.A(net1099));
 sg13g2_antennanp ANTENNA_2142 (.A(net1099));
 sg13g2_antennanp ANTENNA_2143 (.A(net1099));
 sg13g2_antennanp ANTENNA_2144 (.A(net1099));
 sg13g2_antennanp ANTENNA_2145 (.A(net1099));
 sg13g2_antennanp ANTENNA_2146 (.A(net1099));
 sg13g2_antennanp ANTENNA_2147 (.A(net1099));
 sg13g2_antennanp ANTENNA_2148 (.A(net1099));
 sg13g2_antennanp ANTENNA_2149 (.A(net1099));
 sg13g2_antennanp ANTENNA_2150 (.A(net1099));
 sg13g2_antennanp ANTENNA_2151 (.A(net1099));
 sg13g2_antennanp ANTENNA_2152 (.A(net1099));
 sg13g2_antennanp ANTENNA_2153 (.A(net1099));
 sg13g2_antennanp ANTENNA_2154 (.A(net1099));
 sg13g2_antennanp ANTENNA_2155 (.A(net1099));
 sg13g2_antennanp ANTENNA_2156 (.A(net1099));
 sg13g2_antennanp ANTENNA_2157 (.A(net1099));
 sg13g2_antennanp ANTENNA_2158 (.A(net1122));
 sg13g2_antennanp ANTENNA_2159 (.A(net1122));
 sg13g2_antennanp ANTENNA_2160 (.A(net1122));
 sg13g2_antennanp ANTENNA_2161 (.A(net1122));
 sg13g2_antennanp ANTENNA_2162 (.A(net1122));
 sg13g2_antennanp ANTENNA_2163 (.A(net1122));
 sg13g2_antennanp ANTENNA_2164 (.A(net1122));
 sg13g2_antennanp ANTENNA_2165 (.A(net1122));
 sg13g2_antennanp ANTENNA_2166 (.A(net1122));
 sg13g2_antennanp ANTENNA_2167 (.A(_00207_));
 sg13g2_antennanp ANTENNA_2168 (.A(_00785_));
 sg13g2_antennanp ANTENNA_2169 (.A(_00977_));
 sg13g2_antennanp ANTENNA_2170 (.A(_00977_));
 sg13g2_antennanp ANTENNA_2171 (.A(_01032_));
 sg13g2_antennanp ANTENNA_2172 (.A(_01047_));
 sg13g2_antennanp ANTENNA_2173 (.A(_02836_));
 sg13g2_antennanp ANTENNA_2174 (.A(_02836_));
 sg13g2_antennanp ANTENNA_2175 (.A(_02836_));
 sg13g2_antennanp ANTENNA_2176 (.A(_02836_));
 sg13g2_antennanp ANTENNA_2177 (.A(_02845_));
 sg13g2_antennanp ANTENNA_2178 (.A(_02845_));
 sg13g2_antennanp ANTENNA_2179 (.A(_02845_));
 sg13g2_antennanp ANTENNA_2180 (.A(_02845_));
 sg13g2_antennanp ANTENNA_2181 (.A(_02845_));
 sg13g2_antennanp ANTENNA_2182 (.A(_02845_));
 sg13g2_antennanp ANTENNA_2183 (.A(_02845_));
 sg13g2_antennanp ANTENNA_2184 (.A(_02845_));
 sg13g2_antennanp ANTENNA_2185 (.A(_02845_));
 sg13g2_antennanp ANTENNA_2186 (.A(_02849_));
 sg13g2_antennanp ANTENNA_2187 (.A(_02849_));
 sg13g2_antennanp ANTENNA_2188 (.A(_02849_));
 sg13g2_antennanp ANTENNA_2189 (.A(_02849_));
 sg13g2_antennanp ANTENNA_2190 (.A(_02849_));
 sg13g2_antennanp ANTENNA_2191 (.A(_02849_));
 sg13g2_antennanp ANTENNA_2192 (.A(_02849_));
 sg13g2_antennanp ANTENNA_2193 (.A(_02849_));
 sg13g2_antennanp ANTENNA_2194 (.A(_02849_));
 sg13g2_antennanp ANTENNA_2195 (.A(_02861_));
 sg13g2_antennanp ANTENNA_2196 (.A(_02861_));
 sg13g2_antennanp ANTENNA_2197 (.A(_02861_));
 sg13g2_antennanp ANTENNA_2198 (.A(_02861_));
 sg13g2_antennanp ANTENNA_2199 (.A(_02976_));
 sg13g2_antennanp ANTENNA_2200 (.A(_02976_));
 sg13g2_antennanp ANTENNA_2201 (.A(_02976_));
 sg13g2_antennanp ANTENNA_2202 (.A(_02976_));
 sg13g2_antennanp ANTENNA_2203 (.A(_02976_));
 sg13g2_antennanp ANTENNA_2204 (.A(_02976_));
 sg13g2_antennanp ANTENNA_2205 (.A(_02976_));
 sg13g2_antennanp ANTENNA_2206 (.A(_02976_));
 sg13g2_antennanp ANTENNA_2207 (.A(_02976_));
 sg13g2_antennanp ANTENNA_2208 (.A(_03148_));
 sg13g2_antennanp ANTENNA_2209 (.A(_03148_));
 sg13g2_antennanp ANTENNA_2210 (.A(_03507_));
 sg13g2_antennanp ANTENNA_2211 (.A(_03507_));
 sg13g2_antennanp ANTENNA_2212 (.A(_03507_));
 sg13g2_antennanp ANTENNA_2213 (.A(_03507_));
 sg13g2_antennanp ANTENNA_2214 (.A(_03507_));
 sg13g2_antennanp ANTENNA_2215 (.A(_03507_));
 sg13g2_antennanp ANTENNA_2216 (.A(_03513_));
 sg13g2_antennanp ANTENNA_2217 (.A(_03513_));
 sg13g2_antennanp ANTENNA_2218 (.A(_03513_));
 sg13g2_antennanp ANTENNA_2219 (.A(_03513_));
 sg13g2_antennanp ANTENNA_2220 (.A(_03513_));
 sg13g2_antennanp ANTENNA_2221 (.A(_03513_));
 sg13g2_antennanp ANTENNA_2222 (.A(_03513_));
 sg13g2_antennanp ANTENNA_2223 (.A(_03513_));
 sg13g2_antennanp ANTENNA_2224 (.A(_03513_));
 sg13g2_antennanp ANTENNA_2225 (.A(_03539_));
 sg13g2_antennanp ANTENNA_2226 (.A(_03539_));
 sg13g2_antennanp ANTENNA_2227 (.A(_03539_));
 sg13g2_antennanp ANTENNA_2228 (.A(_03539_));
 sg13g2_antennanp ANTENNA_2229 (.A(_03539_));
 sg13g2_antennanp ANTENNA_2230 (.A(_03539_));
 sg13g2_antennanp ANTENNA_2231 (.A(_03539_));
 sg13g2_antennanp ANTENNA_2232 (.A(_03539_));
 sg13g2_antennanp ANTENNA_2233 (.A(_03539_));
 sg13g2_antennanp ANTENNA_2234 (.A(_03824_));
 sg13g2_antennanp ANTENNA_2235 (.A(_03835_));
 sg13g2_antennanp ANTENNA_2236 (.A(_03835_));
 sg13g2_antennanp ANTENNA_2237 (.A(_03835_));
 sg13g2_antennanp ANTENNA_2238 (.A(_03838_));
 sg13g2_antennanp ANTENNA_2239 (.A(_03838_));
 sg13g2_antennanp ANTENNA_2240 (.A(_03838_));
 sg13g2_antennanp ANTENNA_2241 (.A(_04855_));
 sg13g2_antennanp ANTENNA_2242 (.A(_04980_));
 sg13g2_antennanp ANTENNA_2243 (.A(_04980_));
 sg13g2_antennanp ANTENNA_2244 (.A(_04980_));
 sg13g2_antennanp ANTENNA_2245 (.A(_04980_));
 sg13g2_antennanp ANTENNA_2246 (.A(_05006_));
 sg13g2_antennanp ANTENNA_2247 (.A(_05157_));
 sg13g2_antennanp ANTENNA_2248 (.A(_05229_));
 sg13g2_antennanp ANTENNA_2249 (.A(_05260_));
 sg13g2_antennanp ANTENNA_2250 (.A(_05270_));
 sg13g2_antennanp ANTENNA_2251 (.A(_05287_));
 sg13g2_antennanp ANTENNA_2252 (.A(_05314_));
 sg13g2_antennanp ANTENNA_2253 (.A(_05464_));
 sg13g2_antennanp ANTENNA_2254 (.A(_05525_));
 sg13g2_antennanp ANTENNA_2255 (.A(_05529_));
 sg13g2_antennanp ANTENNA_2256 (.A(_05607_));
 sg13g2_antennanp ANTENNA_2257 (.A(_05676_));
 sg13g2_antennanp ANTENNA_2258 (.A(_05756_));
 sg13g2_antennanp ANTENNA_2259 (.A(_05756_));
 sg13g2_antennanp ANTENNA_2260 (.A(_05770_));
 sg13g2_antennanp ANTENNA_2261 (.A(_05780_));
 sg13g2_antennanp ANTENNA_2262 (.A(_05780_));
 sg13g2_antennanp ANTENNA_2263 (.A(_05780_));
 sg13g2_antennanp ANTENNA_2264 (.A(_05780_));
 sg13g2_antennanp ANTENNA_2265 (.A(_05796_));
 sg13g2_antennanp ANTENNA_2266 (.A(_06582_));
 sg13g2_antennanp ANTENNA_2267 (.A(_06582_));
 sg13g2_antennanp ANTENNA_2268 (.A(_06582_));
 sg13g2_antennanp ANTENNA_2269 (.A(_06582_));
 sg13g2_antennanp ANTENNA_2270 (.A(_06582_));
 sg13g2_antennanp ANTENNA_2271 (.A(_06582_));
 sg13g2_antennanp ANTENNA_2272 (.A(_06582_));
 sg13g2_antennanp ANTENNA_2273 (.A(_06582_));
 sg13g2_antennanp ANTENNA_2274 (.A(_06582_));
 sg13g2_antennanp ANTENNA_2275 (.A(_06885_));
 sg13g2_antennanp ANTENNA_2276 (.A(_06885_));
 sg13g2_antennanp ANTENNA_2277 (.A(_06885_));
 sg13g2_antennanp ANTENNA_2278 (.A(_06885_));
 sg13g2_antennanp ANTENNA_2279 (.A(_06885_));
 sg13g2_antennanp ANTENNA_2280 (.A(_06885_));
 sg13g2_antennanp ANTENNA_2281 (.A(_06885_));
 sg13g2_antennanp ANTENNA_2282 (.A(_06885_));
 sg13g2_antennanp ANTENNA_2283 (.A(_06885_));
 sg13g2_antennanp ANTENNA_2284 (.A(_06885_));
 sg13g2_antennanp ANTENNA_2285 (.A(_07626_));
 sg13g2_antennanp ANTENNA_2286 (.A(_07632_));
 sg13g2_antennanp ANTENNA_2287 (.A(_07634_));
 sg13g2_antennanp ANTENNA_2288 (.A(_08260_));
 sg13g2_antennanp ANTENNA_2289 (.A(_08260_));
 sg13g2_antennanp ANTENNA_2290 (.A(_08346_));
 sg13g2_antennanp ANTENNA_2291 (.A(_08346_));
 sg13g2_antennanp ANTENNA_2292 (.A(_08346_));
 sg13g2_antennanp ANTENNA_2293 (.A(_08346_));
 sg13g2_antennanp ANTENNA_2294 (.A(_08346_));
 sg13g2_antennanp ANTENNA_2295 (.A(_08346_));
 sg13g2_antennanp ANTENNA_2296 (.A(_08346_));
 sg13g2_antennanp ANTENNA_2297 (.A(_08346_));
 sg13g2_antennanp ANTENNA_2298 (.A(_08455_));
 sg13g2_antennanp ANTENNA_2299 (.A(_08455_));
 sg13g2_antennanp ANTENNA_2300 (.A(_08455_));
 sg13g2_antennanp ANTENNA_2301 (.A(_08497_));
 sg13g2_antennanp ANTENNA_2302 (.A(_08497_));
 sg13g2_antennanp ANTENNA_2303 (.A(_08497_));
 sg13g2_antennanp ANTENNA_2304 (.A(_08497_));
 sg13g2_antennanp ANTENNA_2305 (.A(_08497_));
 sg13g2_antennanp ANTENNA_2306 (.A(_08497_));
 sg13g2_antennanp ANTENNA_2307 (.A(_08497_));
 sg13g2_antennanp ANTENNA_2308 (.A(_08497_));
 sg13g2_antennanp ANTENNA_2309 (.A(_08497_));
 sg13g2_antennanp ANTENNA_2310 (.A(_08565_));
 sg13g2_antennanp ANTENNA_2311 (.A(_08565_));
 sg13g2_antennanp ANTENNA_2312 (.A(_08565_));
 sg13g2_antennanp ANTENNA_2313 (.A(_08565_));
 sg13g2_antennanp ANTENNA_2314 (.A(_08565_));
 sg13g2_antennanp ANTENNA_2315 (.A(_08565_));
 sg13g2_antennanp ANTENNA_2316 (.A(_08565_));
 sg13g2_antennanp ANTENNA_2317 (.A(_08565_));
 sg13g2_antennanp ANTENNA_2318 (.A(_08565_));
 sg13g2_antennanp ANTENNA_2319 (.A(_08603_));
 sg13g2_antennanp ANTENNA_2320 (.A(_08603_));
 sg13g2_antennanp ANTENNA_2321 (.A(_08603_));
 sg13g2_antennanp ANTENNA_2322 (.A(_08603_));
 sg13g2_antennanp ANTENNA_2323 (.A(_08603_));
 sg13g2_antennanp ANTENNA_2324 (.A(_08603_));
 sg13g2_antennanp ANTENNA_2325 (.A(_08633_));
 sg13g2_antennanp ANTENNA_2326 (.A(_08663_));
 sg13g2_antennanp ANTENNA_2327 (.A(_08663_));
 sg13g2_antennanp ANTENNA_2328 (.A(_08663_));
 sg13g2_antennanp ANTENNA_2329 (.A(_08663_));
 sg13g2_antennanp ANTENNA_2330 (.A(_08663_));
 sg13g2_antennanp ANTENNA_2331 (.A(_08663_));
 sg13g2_antennanp ANTENNA_2332 (.A(_08799_));
 sg13g2_antennanp ANTENNA_2333 (.A(_08799_));
 sg13g2_antennanp ANTENNA_2334 (.A(_08799_));
 sg13g2_antennanp ANTENNA_2335 (.A(_08799_));
 sg13g2_antennanp ANTENNA_2336 (.A(_08799_));
 sg13g2_antennanp ANTENNA_2337 (.A(_08799_));
 sg13g2_antennanp ANTENNA_2338 (.A(_08799_));
 sg13g2_antennanp ANTENNA_2339 (.A(_08799_));
 sg13g2_antennanp ANTENNA_2340 (.A(_08799_));
 sg13g2_antennanp ANTENNA_2341 (.A(_08820_));
 sg13g2_antennanp ANTENNA_2342 (.A(_08820_));
 sg13g2_antennanp ANTENNA_2343 (.A(_08820_));
 sg13g2_antennanp ANTENNA_2344 (.A(_08826_));
 sg13g2_antennanp ANTENNA_2345 (.A(_08826_));
 sg13g2_antennanp ANTENNA_2346 (.A(_08826_));
 sg13g2_antennanp ANTENNA_2347 (.A(_08826_));
 sg13g2_antennanp ANTENNA_2348 (.A(_08826_));
 sg13g2_antennanp ANTENNA_2349 (.A(_08826_));
 sg13g2_antennanp ANTENNA_2350 (.A(_08848_));
 sg13g2_antennanp ANTENNA_2351 (.A(_08848_));
 sg13g2_antennanp ANTENNA_2352 (.A(_08848_));
 sg13g2_antennanp ANTENNA_2353 (.A(_08848_));
 sg13g2_antennanp ANTENNA_2354 (.A(_08848_));
 sg13g2_antennanp ANTENNA_2355 (.A(_08848_));
 sg13g2_antennanp ANTENNA_2356 (.A(_08868_));
 sg13g2_antennanp ANTENNA_2357 (.A(_08900_));
 sg13g2_antennanp ANTENNA_2358 (.A(_08900_));
 sg13g2_antennanp ANTENNA_2359 (.A(_08900_));
 sg13g2_antennanp ANTENNA_2360 (.A(_08950_));
 sg13g2_antennanp ANTENNA_2361 (.A(_08950_));
 sg13g2_antennanp ANTENNA_2362 (.A(_08950_));
 sg13g2_antennanp ANTENNA_2363 (.A(_08950_));
 sg13g2_antennanp ANTENNA_2364 (.A(_08950_));
 sg13g2_antennanp ANTENNA_2365 (.A(_08950_));
 sg13g2_antennanp ANTENNA_2366 (.A(_08950_));
 sg13g2_antennanp ANTENNA_2367 (.A(_08950_));
 sg13g2_antennanp ANTENNA_2368 (.A(_08950_));
 sg13g2_antennanp ANTENNA_2369 (.A(_08970_));
 sg13g2_antennanp ANTENNA_2370 (.A(_08970_));
 sg13g2_antennanp ANTENNA_2371 (.A(_08986_));
 sg13g2_antennanp ANTENNA_2372 (.A(_08986_));
 sg13g2_antennanp ANTENNA_2373 (.A(_09002_));
 sg13g2_antennanp ANTENNA_2374 (.A(_09002_));
 sg13g2_antennanp ANTENNA_2375 (.A(_09065_));
 sg13g2_antennanp ANTENNA_2376 (.A(_09065_));
 sg13g2_antennanp ANTENNA_2377 (.A(_09091_));
 sg13g2_antennanp ANTENNA_2378 (.A(_09091_));
 sg13g2_antennanp ANTENNA_2379 (.A(_09091_));
 sg13g2_antennanp ANTENNA_2380 (.A(_09091_));
 sg13g2_antennanp ANTENNA_2381 (.A(_09091_));
 sg13g2_antennanp ANTENNA_2382 (.A(_09091_));
 sg13g2_antennanp ANTENNA_2383 (.A(_09091_));
 sg13g2_antennanp ANTENNA_2384 (.A(_09091_));
 sg13g2_antennanp ANTENNA_2385 (.A(_09091_));
 sg13g2_antennanp ANTENNA_2386 (.A(_09120_));
 sg13g2_antennanp ANTENNA_2387 (.A(_09120_));
 sg13g2_antennanp ANTENNA_2388 (.A(_09158_));
 sg13g2_antennanp ANTENNA_2389 (.A(_09158_));
 sg13g2_antennanp ANTENNA_2390 (.A(_09158_));
 sg13g2_antennanp ANTENNA_2391 (.A(_09158_));
 sg13g2_antennanp ANTENNA_2392 (.A(_09158_));
 sg13g2_antennanp ANTENNA_2393 (.A(_09158_));
 sg13g2_antennanp ANTENNA_2394 (.A(_09158_));
 sg13g2_antennanp ANTENNA_2395 (.A(_09158_));
 sg13g2_antennanp ANTENNA_2396 (.A(_09173_));
 sg13g2_antennanp ANTENNA_2397 (.A(_09211_));
 sg13g2_antennanp ANTENNA_2398 (.A(_09211_));
 sg13g2_antennanp ANTENNA_2399 (.A(_09211_));
 sg13g2_antennanp ANTENNA_2400 (.A(_09211_));
 sg13g2_antennanp ANTENNA_2401 (.A(_09211_));
 sg13g2_antennanp ANTENNA_2402 (.A(_09218_));
 sg13g2_antennanp ANTENNA_2403 (.A(_09298_));
 sg13g2_antennanp ANTENNA_2404 (.A(_09298_));
 sg13g2_antennanp ANTENNA_2405 (.A(_09298_));
 sg13g2_antennanp ANTENNA_2406 (.A(_09318_));
 sg13g2_antennanp ANTENNA_2407 (.A(_09318_));
 sg13g2_antennanp ANTENNA_2408 (.A(_09318_));
 sg13g2_antennanp ANTENNA_2409 (.A(_09394_));
 sg13g2_antennanp ANTENNA_2410 (.A(_09396_));
 sg13g2_antennanp ANTENNA_2411 (.A(_09447_));
 sg13g2_antennanp ANTENNA_2412 (.A(_09448_));
 sg13g2_antennanp ANTENNA_2413 (.A(_09448_));
 sg13g2_antennanp ANTENNA_2414 (.A(_09448_));
 sg13g2_antennanp ANTENNA_2415 (.A(_09448_));
 sg13g2_antennanp ANTENNA_2416 (.A(_09450_));
 sg13g2_antennanp ANTENNA_2417 (.A(_09492_));
 sg13g2_antennanp ANTENNA_2418 (.A(_09544_));
 sg13g2_antennanp ANTENNA_2419 (.A(_09657_));
 sg13g2_antennanp ANTENNA_2420 (.A(_09722_));
 sg13g2_antennanp ANTENNA_2421 (.A(_09769_));
 sg13g2_antennanp ANTENNA_2422 (.A(_09791_));
 sg13g2_antennanp ANTENNA_2423 (.A(_09852_));
 sg13g2_antennanp ANTENNA_2424 (.A(_09852_));
 sg13g2_antennanp ANTENNA_2425 (.A(_09852_));
 sg13g2_antennanp ANTENNA_2426 (.A(_09852_));
 sg13g2_antennanp ANTENNA_2427 (.A(_09852_));
 sg13g2_antennanp ANTENNA_2428 (.A(_09852_));
 sg13g2_antennanp ANTENNA_2429 (.A(_09852_));
 sg13g2_antennanp ANTENNA_2430 (.A(_09852_));
 sg13g2_antennanp ANTENNA_2431 (.A(_09852_));
 sg13g2_antennanp ANTENNA_2432 (.A(_09852_));
 sg13g2_antennanp ANTENNA_2433 (.A(_09852_));
 sg13g2_antennanp ANTENNA_2434 (.A(_09852_));
 sg13g2_antennanp ANTENNA_2435 (.A(_09852_));
 sg13g2_antennanp ANTENNA_2436 (.A(_09852_));
 sg13g2_antennanp ANTENNA_2437 (.A(_09852_));
 sg13g2_antennanp ANTENNA_2438 (.A(_09852_));
 sg13g2_antennanp ANTENNA_2439 (.A(_09852_));
 sg13g2_antennanp ANTENNA_2440 (.A(_10042_));
 sg13g2_antennanp ANTENNA_2441 (.A(_10042_));
 sg13g2_antennanp ANTENNA_2442 (.A(_10042_));
 sg13g2_antennanp ANTENNA_2443 (.A(_10146_));
 sg13g2_antennanp ANTENNA_2444 (.A(_10146_));
 sg13g2_antennanp ANTENNA_2445 (.A(_10146_));
 sg13g2_antennanp ANTENNA_2446 (.A(_10146_));
 sg13g2_antennanp ANTENNA_2447 (.A(_10146_));
 sg13g2_antennanp ANTENNA_2448 (.A(_10146_));
 sg13g2_antennanp ANTENNA_2449 (.A(_10146_));
 sg13g2_antennanp ANTENNA_2450 (.A(_10146_));
 sg13g2_antennanp ANTENNA_2451 (.A(_10379_));
 sg13g2_antennanp ANTENNA_2452 (.A(_10379_));
 sg13g2_antennanp ANTENNA_2453 (.A(_10379_));
 sg13g2_antennanp ANTENNA_2454 (.A(_10642_));
 sg13g2_antennanp ANTENNA_2455 (.A(_10642_));
 sg13g2_antennanp ANTENNA_2456 (.A(_10642_));
 sg13g2_antennanp ANTENNA_2457 (.A(_10642_));
 sg13g2_antennanp ANTENNA_2458 (.A(_10642_));
 sg13g2_antennanp ANTENNA_2459 (.A(_10642_));
 sg13g2_antennanp ANTENNA_2460 (.A(_10642_));
 sg13g2_antennanp ANTENNA_2461 (.A(_10744_));
 sg13g2_antennanp ANTENNA_2462 (.A(_10744_));
 sg13g2_antennanp ANTENNA_2463 (.A(_10744_));
 sg13g2_antennanp ANTENNA_2464 (.A(_10744_));
 sg13g2_antennanp ANTENNA_2465 (.A(_12205_));
 sg13g2_antennanp ANTENNA_2466 (.A(_12205_));
 sg13g2_antennanp ANTENNA_2467 (.A(_12205_));
 sg13g2_antennanp ANTENNA_2468 (.A(_12205_));
 sg13g2_antennanp ANTENNA_2469 (.A(_12218_));
 sg13g2_antennanp ANTENNA_2470 (.A(_12218_));
 sg13g2_antennanp ANTENNA_2471 (.A(_12218_));
 sg13g2_antennanp ANTENNA_2472 (.A(_12218_));
 sg13g2_antennanp ANTENNA_2473 (.A(_12218_));
 sg13g2_antennanp ANTENNA_2474 (.A(_12218_));
 sg13g2_antennanp ANTENNA_2475 (.A(_12218_));
 sg13g2_antennanp ANTENNA_2476 (.A(_12218_));
 sg13g2_antennanp ANTENNA_2477 (.A(_12218_));
 sg13g2_antennanp ANTENNA_2478 (.A(_12225_));
 sg13g2_antennanp ANTENNA_2479 (.A(_12225_));
 sg13g2_antennanp ANTENNA_2480 (.A(_12225_));
 sg13g2_antennanp ANTENNA_2481 (.A(_12225_));
 sg13g2_antennanp ANTENNA_2482 (.A(_12225_));
 sg13g2_antennanp ANTENNA_2483 (.A(_12225_));
 sg13g2_antennanp ANTENNA_2484 (.A(_12225_));
 sg13g2_antennanp ANTENNA_2485 (.A(_12225_));
 sg13g2_antennanp ANTENNA_2486 (.A(_12225_));
 sg13g2_antennanp ANTENNA_2487 (.A(_12236_));
 sg13g2_antennanp ANTENNA_2488 (.A(_12236_));
 sg13g2_antennanp ANTENNA_2489 (.A(_12236_));
 sg13g2_antennanp ANTENNA_2490 (.A(_12236_));
 sg13g2_antennanp ANTENNA_2491 (.A(_12236_));
 sg13g2_antennanp ANTENNA_2492 (.A(_12236_));
 sg13g2_antennanp ANTENNA_2493 (.A(_12236_));
 sg13g2_antennanp ANTENNA_2494 (.A(_12236_));
 sg13g2_antennanp ANTENNA_2495 (.A(_12236_));
 sg13g2_antennanp ANTENNA_2496 (.A(\cpu.dcache.wdata[10] ));
 sg13g2_antennanp ANTENNA_2497 (.A(\cpu.dcache.wdata[10] ));
 sg13g2_antennanp ANTENNA_2498 (.A(\cpu.dcache.wdata[10] ));
 sg13g2_antennanp ANTENNA_2499 (.A(\cpu.dcache.wdata[10] ));
 sg13g2_antennanp ANTENNA_2500 (.A(\cpu.dcache.wdata[12] ));
 sg13g2_antennanp ANTENNA_2501 (.A(\cpu.dcache.wdata[12] ));
 sg13g2_antennanp ANTENNA_2502 (.A(\cpu.dcache.wdata[12] ));
 sg13g2_antennanp ANTENNA_2503 (.A(\cpu.dcache.wdata[12] ));
 sg13g2_antennanp ANTENNA_2504 (.A(\cpu.dcache.wdata[9] ));
 sg13g2_antennanp ANTENNA_2505 (.A(\cpu.dcache.wdata[9] ));
 sg13g2_antennanp ANTENNA_2506 (.A(\cpu.dcache.wdata[9] ));
 sg13g2_antennanp ANTENNA_2507 (.A(\cpu.dcache.wdata[9] ));
 sg13g2_antennanp ANTENNA_2508 (.A(\cpu.ex.pc[1] ));
 sg13g2_antennanp ANTENNA_2509 (.A(\cpu.ex.pc[2] ));
 sg13g2_antennanp ANTENNA_2510 (.A(\cpu.gpio.uart_rx ));
 sg13g2_antennanp ANTENNA_2511 (.A(\cpu.gpio.uart_rx ));
 sg13g2_antennanp ANTENNA_2512 (.A(\cpu.qspi.c_wstrobe_i ));
 sg13g2_antennanp ANTENNA_2513 (.A(\cpu.qspi.c_wstrobe_i ));
 sg13g2_antennanp ANTENNA_2514 (.A(net3));
 sg13g2_antennanp ANTENNA_2515 (.A(net3));
 sg13g2_antennanp ANTENNA_2516 (.A(net3));
 sg13g2_antennanp ANTENNA_2517 (.A(net12));
 sg13g2_antennanp ANTENNA_2518 (.A(net12));
 sg13g2_antennanp ANTENNA_2519 (.A(net12));
 sg13g2_antennanp ANTENNA_2520 (.A(net13));
 sg13g2_antennanp ANTENNA_2521 (.A(net13));
 sg13g2_antennanp ANTENNA_2522 (.A(net13));
 sg13g2_antennanp ANTENNA_2523 (.A(net14));
 sg13g2_antennanp ANTENNA_2524 (.A(net14));
 sg13g2_antennanp ANTENNA_2525 (.A(net14));
 sg13g2_antennanp ANTENNA_2526 (.A(net489));
 sg13g2_antennanp ANTENNA_2527 (.A(net489));
 sg13g2_antennanp ANTENNA_2528 (.A(net489));
 sg13g2_antennanp ANTENNA_2529 (.A(net489));
 sg13g2_antennanp ANTENNA_2530 (.A(net489));
 sg13g2_antennanp ANTENNA_2531 (.A(net489));
 sg13g2_antennanp ANTENNA_2532 (.A(net489));
 sg13g2_antennanp ANTENNA_2533 (.A(net489));
 sg13g2_antennanp ANTENNA_2534 (.A(net489));
 sg13g2_antennanp ANTENNA_2535 (.A(net491));
 sg13g2_antennanp ANTENNA_2536 (.A(net491));
 sg13g2_antennanp ANTENNA_2537 (.A(net491));
 sg13g2_antennanp ANTENNA_2538 (.A(net491));
 sg13g2_antennanp ANTENNA_2539 (.A(net491));
 sg13g2_antennanp ANTENNA_2540 (.A(net491));
 sg13g2_antennanp ANTENNA_2541 (.A(net491));
 sg13g2_antennanp ANTENNA_2542 (.A(net491));
 sg13g2_antennanp ANTENNA_2543 (.A(net491));
 sg13g2_antennanp ANTENNA_2544 (.A(net491));
 sg13g2_antennanp ANTENNA_2545 (.A(net491));
 sg13g2_antennanp ANTENNA_2546 (.A(net491));
 sg13g2_antennanp ANTENNA_2547 (.A(net550));
 sg13g2_antennanp ANTENNA_2548 (.A(net550));
 sg13g2_antennanp ANTENNA_2549 (.A(net550));
 sg13g2_antennanp ANTENNA_2550 (.A(net550));
 sg13g2_antennanp ANTENNA_2551 (.A(net550));
 sg13g2_antennanp ANTENNA_2552 (.A(net550));
 sg13g2_antennanp ANTENNA_2553 (.A(net550));
 sg13g2_antennanp ANTENNA_2554 (.A(net550));
 sg13g2_antennanp ANTENNA_2555 (.A(net550));
 sg13g2_antennanp ANTENNA_2556 (.A(net550));
 sg13g2_antennanp ANTENNA_2557 (.A(net550));
 sg13g2_antennanp ANTENNA_2558 (.A(net686));
 sg13g2_antennanp ANTENNA_2559 (.A(net686));
 sg13g2_antennanp ANTENNA_2560 (.A(net686));
 sg13g2_antennanp ANTENNA_2561 (.A(net686));
 sg13g2_antennanp ANTENNA_2562 (.A(net686));
 sg13g2_antennanp ANTENNA_2563 (.A(net686));
 sg13g2_antennanp ANTENNA_2564 (.A(net686));
 sg13g2_antennanp ANTENNA_2565 (.A(net686));
 sg13g2_antennanp ANTENNA_2566 (.A(net708));
 sg13g2_antennanp ANTENNA_2567 (.A(net708));
 sg13g2_antennanp ANTENNA_2568 (.A(net708));
 sg13g2_antennanp ANTENNA_2569 (.A(net708));
 sg13g2_antennanp ANTENNA_2570 (.A(net708));
 sg13g2_antennanp ANTENNA_2571 (.A(net708));
 sg13g2_antennanp ANTENNA_2572 (.A(net708));
 sg13g2_antennanp ANTENNA_2573 (.A(net708));
 sg13g2_antennanp ANTENNA_2574 (.A(net745));
 sg13g2_antennanp ANTENNA_2575 (.A(net745));
 sg13g2_antennanp ANTENNA_2576 (.A(net745));
 sg13g2_antennanp ANTENNA_2577 (.A(net745));
 sg13g2_antennanp ANTENNA_2578 (.A(net745));
 sg13g2_antennanp ANTENNA_2579 (.A(net745));
 sg13g2_antennanp ANTENNA_2580 (.A(net745));
 sg13g2_antennanp ANTENNA_2581 (.A(net745));
 sg13g2_antennanp ANTENNA_2582 (.A(net803));
 sg13g2_antennanp ANTENNA_2583 (.A(net803));
 sg13g2_antennanp ANTENNA_2584 (.A(net803));
 sg13g2_antennanp ANTENNA_2585 (.A(net803));
 sg13g2_antennanp ANTENNA_2586 (.A(net803));
 sg13g2_antennanp ANTENNA_2587 (.A(net803));
 sg13g2_antennanp ANTENNA_2588 (.A(net803));
 sg13g2_antennanp ANTENNA_2589 (.A(net803));
 sg13g2_antennanp ANTENNA_2590 (.A(net858));
 sg13g2_antennanp ANTENNA_2591 (.A(net858));
 sg13g2_antennanp ANTENNA_2592 (.A(net858));
 sg13g2_antennanp ANTENNA_2593 (.A(net858));
 sg13g2_antennanp ANTENNA_2594 (.A(net858));
 sg13g2_antennanp ANTENNA_2595 (.A(net858));
 sg13g2_antennanp ANTENNA_2596 (.A(net858));
 sg13g2_antennanp ANTENNA_2597 (.A(net858));
 sg13g2_antennanp ANTENNA_2598 (.A(net858));
 sg13g2_antennanp ANTENNA_2599 (.A(net872));
 sg13g2_antennanp ANTENNA_2600 (.A(net872));
 sg13g2_antennanp ANTENNA_2601 (.A(net872));
 sg13g2_antennanp ANTENNA_2602 (.A(net872));
 sg13g2_antennanp ANTENNA_2603 (.A(net872));
 sg13g2_antennanp ANTENNA_2604 (.A(net872));
 sg13g2_antennanp ANTENNA_2605 (.A(net872));
 sg13g2_antennanp ANTENNA_2606 (.A(net872));
 sg13g2_antennanp ANTENNA_2607 (.A(net872));
 sg13g2_antennanp ANTENNA_2608 (.A(net872));
 sg13g2_antennanp ANTENNA_2609 (.A(net872));
 sg13g2_antennanp ANTENNA_2610 (.A(net872));
 sg13g2_antennanp ANTENNA_2611 (.A(net872));
 sg13g2_antennanp ANTENNA_2612 (.A(net872));
 sg13g2_antennanp ANTENNA_2613 (.A(net872));
 sg13g2_antennanp ANTENNA_2614 (.A(net872));
 sg13g2_antennanp ANTENNA_2615 (.A(net872));
 sg13g2_antennanp ANTENNA_2616 (.A(net872));
 sg13g2_antennanp ANTENNA_2617 (.A(net872));
 sg13g2_antennanp ANTENNA_2618 (.A(net872));
 sg13g2_antennanp ANTENNA_2619 (.A(net872));
 sg13g2_antennanp ANTENNA_2620 (.A(net872));
 sg13g2_antennanp ANTENNA_2621 (.A(net872));
 sg13g2_antennanp ANTENNA_2622 (.A(net872));
 sg13g2_antennanp ANTENNA_2623 (.A(net872));
 sg13g2_antennanp ANTENNA_2624 (.A(net872));
 sg13g2_antennanp ANTENNA_2625 (.A(net872));
 sg13g2_antennanp ANTENNA_2626 (.A(net872));
 sg13g2_antennanp ANTENNA_2627 (.A(net872));
 sg13g2_antennanp ANTENNA_2628 (.A(net872));
 sg13g2_antennanp ANTENNA_2629 (.A(net872));
 sg13g2_antennanp ANTENNA_2630 (.A(net872));
 sg13g2_antennanp ANTENNA_2631 (.A(net872));
 sg13g2_antennanp ANTENNA_2632 (.A(net872));
 sg13g2_antennanp ANTENNA_2633 (.A(net872));
 sg13g2_antennanp ANTENNA_2634 (.A(net872));
 sg13g2_antennanp ANTENNA_2635 (.A(net872));
 sg13g2_antennanp ANTENNA_2636 (.A(net872));
 sg13g2_antennanp ANTENNA_2637 (.A(net872));
 sg13g2_antennanp ANTENNA_2638 (.A(net872));
 sg13g2_antennanp ANTENNA_2639 (.A(net872));
 sg13g2_antennanp ANTENNA_2640 (.A(net872));
 sg13g2_antennanp ANTENNA_2641 (.A(net872));
 sg13g2_antennanp ANTENNA_2642 (.A(net872));
 sg13g2_antennanp ANTENNA_2643 (.A(net872));
 sg13g2_antennanp ANTENNA_2644 (.A(net928));
 sg13g2_antennanp ANTENNA_2645 (.A(net928));
 sg13g2_antennanp ANTENNA_2646 (.A(net928));
 sg13g2_antennanp ANTENNA_2647 (.A(net928));
 sg13g2_antennanp ANTENNA_2648 (.A(net928));
 sg13g2_antennanp ANTENNA_2649 (.A(net928));
 sg13g2_antennanp ANTENNA_2650 (.A(net928));
 sg13g2_antennanp ANTENNA_2651 (.A(net928));
 sg13g2_antennanp ANTENNA_2652 (.A(net928));
 sg13g2_antennanp ANTENNA_2653 (.A(net928));
 sg13g2_antennanp ANTENNA_2654 (.A(net928));
 sg13g2_antennanp ANTENNA_2655 (.A(net928));
 sg13g2_antennanp ANTENNA_2656 (.A(net983));
 sg13g2_antennanp ANTENNA_2657 (.A(net983));
 sg13g2_antennanp ANTENNA_2658 (.A(net983));
 sg13g2_antennanp ANTENNA_2659 (.A(net983));
 sg13g2_antennanp ANTENNA_2660 (.A(net983));
 sg13g2_antennanp ANTENNA_2661 (.A(net983));
 sg13g2_antennanp ANTENNA_2662 (.A(net983));
 sg13g2_antennanp ANTENNA_2663 (.A(net983));
 sg13g2_antennanp ANTENNA_2664 (.A(net983));
 sg13g2_antennanp ANTENNA_2665 (.A(net983));
 sg13g2_antennanp ANTENNA_2666 (.A(net983));
 sg13g2_antennanp ANTENNA_2667 (.A(net983));
 sg13g2_antennanp ANTENNA_2668 (.A(net983));
 sg13g2_antennanp ANTENNA_2669 (.A(net983));
 sg13g2_antennanp ANTENNA_2670 (.A(net983));
 sg13g2_antennanp ANTENNA_2671 (.A(net983));
 sg13g2_antennanp ANTENNA_2672 (.A(net983));
 sg13g2_antennanp ANTENNA_2673 (.A(net995));
 sg13g2_antennanp ANTENNA_2674 (.A(net995));
 sg13g2_antennanp ANTENNA_2675 (.A(net995));
 sg13g2_antennanp ANTENNA_2676 (.A(net995));
 sg13g2_antennanp ANTENNA_2677 (.A(net995));
 sg13g2_antennanp ANTENNA_2678 (.A(net995));
 sg13g2_antennanp ANTENNA_2679 (.A(net995));
 sg13g2_antennanp ANTENNA_2680 (.A(net995));
 sg13g2_antennanp ANTENNA_2681 (.A(net995));
 sg13g2_antennanp ANTENNA_2682 (.A(net995));
 sg13g2_antennanp ANTENNA_2683 (.A(net995));
 sg13g2_antennanp ANTENNA_2684 (.A(net995));
 sg13g2_antennanp ANTENNA_2685 (.A(net995));
 sg13g2_antennanp ANTENNA_2686 (.A(net995));
 sg13g2_antennanp ANTENNA_2687 (.A(net995));
 sg13g2_antennanp ANTENNA_2688 (.A(net995));
 sg13g2_antennanp ANTENNA_2689 (.A(net995));
 sg13g2_antennanp ANTENNA_2690 (.A(net995));
 sg13g2_antennanp ANTENNA_2691 (.A(net999));
 sg13g2_antennanp ANTENNA_2692 (.A(net999));
 sg13g2_antennanp ANTENNA_2693 (.A(net999));
 sg13g2_antennanp ANTENNA_2694 (.A(net999));
 sg13g2_antennanp ANTENNA_2695 (.A(net999));
 sg13g2_antennanp ANTENNA_2696 (.A(net999));
 sg13g2_antennanp ANTENNA_2697 (.A(net999));
 sg13g2_antennanp ANTENNA_2698 (.A(net999));
 sg13g2_antennanp ANTENNA_2699 (.A(net999));
 sg13g2_antennanp ANTENNA_2700 (.A(net1000));
 sg13g2_antennanp ANTENNA_2701 (.A(net1000));
 sg13g2_antennanp ANTENNA_2702 (.A(net1000));
 sg13g2_antennanp ANTENNA_2703 (.A(net1000));
 sg13g2_antennanp ANTENNA_2704 (.A(net1000));
 sg13g2_antennanp ANTENNA_2705 (.A(net1000));
 sg13g2_antennanp ANTENNA_2706 (.A(net1000));
 sg13g2_antennanp ANTENNA_2707 (.A(net1000));
 sg13g2_antennanp ANTENNA_2708 (.A(net1000));
 sg13g2_antennanp ANTENNA_2709 (.A(net1000));
 sg13g2_antennanp ANTENNA_2710 (.A(net1000));
 sg13g2_antennanp ANTENNA_2711 (.A(net1000));
 sg13g2_antennanp ANTENNA_2712 (.A(net1000));
 sg13g2_antennanp ANTENNA_2713 (.A(net1002));
 sg13g2_antennanp ANTENNA_2714 (.A(net1002));
 sg13g2_antennanp ANTENNA_2715 (.A(net1002));
 sg13g2_antennanp ANTENNA_2716 (.A(net1002));
 sg13g2_antennanp ANTENNA_2717 (.A(net1002));
 sg13g2_antennanp ANTENNA_2718 (.A(net1002));
 sg13g2_antennanp ANTENNA_2719 (.A(net1002));
 sg13g2_antennanp ANTENNA_2720 (.A(net1002));
 sg13g2_antennanp ANTENNA_2721 (.A(net1002));
 sg13g2_antennanp ANTENNA_2722 (.A(net1004));
 sg13g2_antennanp ANTENNA_2723 (.A(net1004));
 sg13g2_antennanp ANTENNA_2724 (.A(net1004));
 sg13g2_antennanp ANTENNA_2725 (.A(net1004));
 sg13g2_antennanp ANTENNA_2726 (.A(net1004));
 sg13g2_antennanp ANTENNA_2727 (.A(net1004));
 sg13g2_antennanp ANTENNA_2728 (.A(net1004));
 sg13g2_antennanp ANTENNA_2729 (.A(net1004));
 sg13g2_antennanp ANTENNA_2730 (.A(net1004));
 sg13g2_antennanp ANTENNA_2731 (.A(net1099));
 sg13g2_antennanp ANTENNA_2732 (.A(net1099));
 sg13g2_antennanp ANTENNA_2733 (.A(net1099));
 sg13g2_antennanp ANTENNA_2734 (.A(net1099));
 sg13g2_antennanp ANTENNA_2735 (.A(net1099));
 sg13g2_antennanp ANTENNA_2736 (.A(net1099));
 sg13g2_antennanp ANTENNA_2737 (.A(net1099));
 sg13g2_antennanp ANTENNA_2738 (.A(net1099));
 sg13g2_antennanp ANTENNA_2739 (.A(net1099));
 sg13g2_antennanp ANTENNA_2740 (.A(net1099));
 sg13g2_antennanp ANTENNA_2741 (.A(net1099));
 sg13g2_antennanp ANTENNA_2742 (.A(net1099));
 sg13g2_antennanp ANTENNA_2743 (.A(net1099));
 sg13g2_antennanp ANTENNA_2744 (.A(net1099));
 sg13g2_antennanp ANTENNA_2745 (.A(net1099));
 sg13g2_antennanp ANTENNA_2746 (.A(net1099));
 sg13g2_antennanp ANTENNA_2747 (.A(net1099));
 sg13g2_antennanp ANTENNA_2748 (.A(net1099));
 sg13g2_antennanp ANTENNA_2749 (.A(net1099));
 sg13g2_antennanp ANTENNA_2750 (.A(net1099));
 sg13g2_antennanp ANTENNA_2751 (.A(net1122));
 sg13g2_antennanp ANTENNA_2752 (.A(net1122));
 sg13g2_antennanp ANTENNA_2753 (.A(net1122));
 sg13g2_antennanp ANTENNA_2754 (.A(net1122));
 sg13g2_antennanp ANTENNA_2755 (.A(net1122));
 sg13g2_antennanp ANTENNA_2756 (.A(net1122));
 sg13g2_antennanp ANTENNA_2757 (.A(net1122));
 sg13g2_antennanp ANTENNA_2758 (.A(net1122));
 sg13g2_antennanp ANTENNA_2759 (.A(net1122));
 sg13g2_antennanp ANTENNA_2760 (.A(_00207_));
 sg13g2_antennanp ANTENNA_2761 (.A(_00785_));
 sg13g2_antennanp ANTENNA_2762 (.A(_00977_));
 sg13g2_antennanp ANTENNA_2763 (.A(_00977_));
 sg13g2_antennanp ANTENNA_2764 (.A(_01032_));
 sg13g2_antennanp ANTENNA_2765 (.A(_01047_));
 sg13g2_antennanp ANTENNA_2766 (.A(_02836_));
 sg13g2_antennanp ANTENNA_2767 (.A(_02836_));
 sg13g2_antennanp ANTENNA_2768 (.A(_02836_));
 sg13g2_antennanp ANTENNA_2769 (.A(_02836_));
 sg13g2_antennanp ANTENNA_2770 (.A(_02836_));
 sg13g2_antennanp ANTENNA_2771 (.A(_02836_));
 sg13g2_antennanp ANTENNA_2772 (.A(_02836_));
 sg13g2_antennanp ANTENNA_2773 (.A(_02836_));
 sg13g2_antennanp ANTENNA_2774 (.A(_02836_));
 sg13g2_antennanp ANTENNA_2775 (.A(_02845_));
 sg13g2_antennanp ANTENNA_2776 (.A(_02845_));
 sg13g2_antennanp ANTENNA_2777 (.A(_02845_));
 sg13g2_antennanp ANTENNA_2778 (.A(_02845_));
 sg13g2_antennanp ANTENNA_2779 (.A(_02845_));
 sg13g2_antennanp ANTENNA_2780 (.A(_02845_));
 sg13g2_antennanp ANTENNA_2781 (.A(_02845_));
 sg13g2_antennanp ANTENNA_2782 (.A(_02845_));
 sg13g2_antennanp ANTENNA_2783 (.A(_02845_));
 sg13g2_antennanp ANTENNA_2784 (.A(_02849_));
 sg13g2_antennanp ANTENNA_2785 (.A(_02849_));
 sg13g2_antennanp ANTENNA_2786 (.A(_02849_));
 sg13g2_antennanp ANTENNA_2787 (.A(_02849_));
 sg13g2_antennanp ANTENNA_2788 (.A(_02849_));
 sg13g2_antennanp ANTENNA_2789 (.A(_02849_));
 sg13g2_antennanp ANTENNA_2790 (.A(_02849_));
 sg13g2_antennanp ANTENNA_2791 (.A(_02849_));
 sg13g2_antennanp ANTENNA_2792 (.A(_02849_));
 sg13g2_antennanp ANTENNA_2793 (.A(_02861_));
 sg13g2_antennanp ANTENNA_2794 (.A(_02861_));
 sg13g2_antennanp ANTENNA_2795 (.A(_02861_));
 sg13g2_antennanp ANTENNA_2796 (.A(_02861_));
 sg13g2_antennanp ANTENNA_2797 (.A(_02976_));
 sg13g2_antennanp ANTENNA_2798 (.A(_02976_));
 sg13g2_antennanp ANTENNA_2799 (.A(_02976_));
 sg13g2_antennanp ANTENNA_2800 (.A(_02976_));
 sg13g2_antennanp ANTENNA_2801 (.A(_02976_));
 sg13g2_antennanp ANTENNA_2802 (.A(_02976_));
 sg13g2_antennanp ANTENNA_2803 (.A(_02976_));
 sg13g2_antennanp ANTENNA_2804 (.A(_02976_));
 sg13g2_antennanp ANTENNA_2805 (.A(_02976_));
 sg13g2_antennanp ANTENNA_2806 (.A(_02976_));
 sg13g2_antennanp ANTENNA_2807 (.A(_02976_));
 sg13g2_antennanp ANTENNA_2808 (.A(_03148_));
 sg13g2_antennanp ANTENNA_2809 (.A(_03148_));
 sg13g2_antennanp ANTENNA_2810 (.A(_03507_));
 sg13g2_antennanp ANTENNA_2811 (.A(_03507_));
 sg13g2_antennanp ANTENNA_2812 (.A(_03507_));
 sg13g2_antennanp ANTENNA_2813 (.A(_03507_));
 sg13g2_antennanp ANTENNA_2814 (.A(_03507_));
 sg13g2_antennanp ANTENNA_2815 (.A(_03507_));
 sg13g2_antennanp ANTENNA_2816 (.A(_03507_));
 sg13g2_antennanp ANTENNA_2817 (.A(_03507_));
 sg13g2_antennanp ANTENNA_2818 (.A(_03513_));
 sg13g2_antennanp ANTENNA_2819 (.A(_03513_));
 sg13g2_antennanp ANTENNA_2820 (.A(_03513_));
 sg13g2_antennanp ANTENNA_2821 (.A(_03513_));
 sg13g2_antennanp ANTENNA_2822 (.A(_03513_));
 sg13g2_antennanp ANTENNA_2823 (.A(_03513_));
 sg13g2_antennanp ANTENNA_2824 (.A(_03513_));
 sg13g2_antennanp ANTENNA_2825 (.A(_03513_));
 sg13g2_antennanp ANTENNA_2826 (.A(_03513_));
 sg13g2_antennanp ANTENNA_2827 (.A(_03513_));
 sg13g2_antennanp ANTENNA_2828 (.A(_03513_));
 sg13g2_antennanp ANTENNA_2829 (.A(_03513_));
 sg13g2_antennanp ANTENNA_2830 (.A(_03513_));
 sg13g2_antennanp ANTENNA_2831 (.A(_03513_));
 sg13g2_antennanp ANTENNA_2832 (.A(_03539_));
 sg13g2_antennanp ANTENNA_2833 (.A(_03539_));
 sg13g2_antennanp ANTENNA_2834 (.A(_03539_));
 sg13g2_antennanp ANTENNA_2835 (.A(_03539_));
 sg13g2_antennanp ANTENNA_2836 (.A(_03838_));
 sg13g2_antennanp ANTENNA_2837 (.A(_03838_));
 sg13g2_antennanp ANTENNA_2838 (.A(_03838_));
 sg13g2_antennanp ANTENNA_2839 (.A(_04855_));
 sg13g2_antennanp ANTENNA_2840 (.A(_04980_));
 sg13g2_antennanp ANTENNA_2841 (.A(_04980_));
 sg13g2_antennanp ANTENNA_2842 (.A(_04980_));
 sg13g2_antennanp ANTENNA_2843 (.A(_04980_));
 sg13g2_antennanp ANTENNA_2844 (.A(_05006_));
 sg13g2_antennanp ANTENNA_2845 (.A(_05157_));
 sg13g2_antennanp ANTENNA_2846 (.A(_05229_));
 sg13g2_antennanp ANTENNA_2847 (.A(_05260_));
 sg13g2_antennanp ANTENNA_2848 (.A(_05270_));
 sg13g2_antennanp ANTENNA_2849 (.A(_05287_));
 sg13g2_antennanp ANTENNA_2850 (.A(_05307_));
 sg13g2_antennanp ANTENNA_2851 (.A(_05307_));
 sg13g2_antennanp ANTENNA_2852 (.A(_05314_));
 sg13g2_antennanp ANTENNA_2853 (.A(_05464_));
 sg13g2_antennanp ANTENNA_2854 (.A(_05525_));
 sg13g2_antennanp ANTENNA_2855 (.A(_05529_));
 sg13g2_antennanp ANTENNA_2856 (.A(_05607_));
 sg13g2_antennanp ANTENNA_2857 (.A(_05676_));
 sg13g2_antennanp ANTENNA_2858 (.A(_05756_));
 sg13g2_antennanp ANTENNA_2859 (.A(_05770_));
 sg13g2_antennanp ANTENNA_2860 (.A(_05780_));
 sg13g2_antennanp ANTENNA_2861 (.A(_05780_));
 sg13g2_antennanp ANTENNA_2862 (.A(_05780_));
 sg13g2_antennanp ANTENNA_2863 (.A(_05780_));
 sg13g2_antennanp ANTENNA_2864 (.A(_05780_));
 sg13g2_antennanp ANTENNA_2865 (.A(_05780_));
 sg13g2_antennanp ANTENNA_2866 (.A(_05780_));
 sg13g2_antennanp ANTENNA_2867 (.A(_05780_));
 sg13g2_antennanp ANTENNA_2868 (.A(_05796_));
 sg13g2_antennanp ANTENNA_2869 (.A(_06582_));
 sg13g2_antennanp ANTENNA_2870 (.A(_06582_));
 sg13g2_antennanp ANTENNA_2871 (.A(_06582_));
 sg13g2_antennanp ANTENNA_2872 (.A(_06582_));
 sg13g2_antennanp ANTENNA_2873 (.A(_06583_));
 sg13g2_antennanp ANTENNA_2874 (.A(_06583_));
 sg13g2_antennanp ANTENNA_2875 (.A(_06583_));
 sg13g2_antennanp ANTENNA_2876 (.A(_06583_));
 sg13g2_antennanp ANTENNA_2877 (.A(_06583_));
 sg13g2_antennanp ANTENNA_2878 (.A(_06583_));
 sg13g2_antennanp ANTENNA_2879 (.A(_06583_));
 sg13g2_antennanp ANTENNA_2880 (.A(_06583_));
 sg13g2_antennanp ANTENNA_2881 (.A(_06583_));
 sg13g2_antennanp ANTENNA_2882 (.A(_06885_));
 sg13g2_antennanp ANTENNA_2883 (.A(_06885_));
 sg13g2_antennanp ANTENNA_2884 (.A(_06885_));
 sg13g2_antennanp ANTENNA_2885 (.A(_06885_));
 sg13g2_antennanp ANTENNA_2886 (.A(_06885_));
 sg13g2_antennanp ANTENNA_2887 (.A(_06885_));
 sg13g2_antennanp ANTENNA_2888 (.A(_06885_));
 sg13g2_antennanp ANTENNA_2889 (.A(_06885_));
 sg13g2_antennanp ANTENNA_2890 (.A(_06885_));
 sg13g2_antennanp ANTENNA_2891 (.A(_06885_));
 sg13g2_antennanp ANTENNA_2892 (.A(_07626_));
 sg13g2_antennanp ANTENNA_2893 (.A(_07632_));
 sg13g2_antennanp ANTENNA_2894 (.A(_07634_));
 sg13g2_antennanp ANTENNA_2895 (.A(_08260_));
 sg13g2_antennanp ANTENNA_2896 (.A(_08260_));
 sg13g2_antennanp ANTENNA_2897 (.A(_08346_));
 sg13g2_antennanp ANTENNA_2898 (.A(_08346_));
 sg13g2_antennanp ANTENNA_2899 (.A(_08346_));
 sg13g2_antennanp ANTENNA_2900 (.A(_08346_));
 sg13g2_antennanp ANTENNA_2901 (.A(_08346_));
 sg13g2_antennanp ANTENNA_2902 (.A(_08346_));
 sg13g2_antennanp ANTENNA_2903 (.A(_08346_));
 sg13g2_antennanp ANTENNA_2904 (.A(_08346_));
 sg13g2_antennanp ANTENNA_2905 (.A(_08455_));
 sg13g2_antennanp ANTENNA_2906 (.A(_08455_));
 sg13g2_antennanp ANTENNA_2907 (.A(_08455_));
 sg13g2_antennanp ANTENNA_2908 (.A(_08497_));
 sg13g2_antennanp ANTENNA_2909 (.A(_08497_));
 sg13g2_antennanp ANTENNA_2910 (.A(_08497_));
 sg13g2_antennanp ANTENNA_2911 (.A(_08565_));
 sg13g2_antennanp ANTENNA_2912 (.A(_08565_));
 sg13g2_antennanp ANTENNA_2913 (.A(_08565_));
 sg13g2_antennanp ANTENNA_2914 (.A(_08565_));
 sg13g2_antennanp ANTENNA_2915 (.A(_08565_));
 sg13g2_antennanp ANTENNA_2916 (.A(_08565_));
 sg13g2_antennanp ANTENNA_2917 (.A(_08565_));
 sg13g2_antennanp ANTENNA_2918 (.A(_08565_));
 sg13g2_antennanp ANTENNA_2919 (.A(_08565_));
 sg13g2_antennanp ANTENNA_2920 (.A(_08603_));
 sg13g2_antennanp ANTENNA_2921 (.A(_08603_));
 sg13g2_antennanp ANTENNA_2922 (.A(_08603_));
 sg13g2_antennanp ANTENNA_2923 (.A(_08603_));
 sg13g2_antennanp ANTENNA_2924 (.A(_08603_));
 sg13g2_antennanp ANTENNA_2925 (.A(_08603_));
 sg13g2_antennanp ANTENNA_2926 (.A(_08603_));
 sg13g2_antennanp ANTENNA_2927 (.A(_08603_));
 sg13g2_antennanp ANTENNA_2928 (.A(_08603_));
 sg13g2_antennanp ANTENNA_2929 (.A(_08633_));
 sg13g2_antennanp ANTENNA_2930 (.A(_08663_));
 sg13g2_antennanp ANTENNA_2931 (.A(_08663_));
 sg13g2_antennanp ANTENNA_2932 (.A(_08663_));
 sg13g2_antennanp ANTENNA_2933 (.A(_08663_));
 sg13g2_antennanp ANTENNA_2934 (.A(_08663_));
 sg13g2_antennanp ANTENNA_2935 (.A(_08663_));
 sg13g2_antennanp ANTENNA_2936 (.A(_08663_));
 sg13g2_antennanp ANTENNA_2937 (.A(_08663_));
 sg13g2_antennanp ANTENNA_2938 (.A(_08663_));
 sg13g2_antennanp ANTENNA_2939 (.A(_08799_));
 sg13g2_antennanp ANTENNA_2940 (.A(_08799_));
 sg13g2_antennanp ANTENNA_2941 (.A(_08799_));
 sg13g2_antennanp ANTENNA_2942 (.A(_08799_));
 sg13g2_antennanp ANTENNA_2943 (.A(_08799_));
 sg13g2_antennanp ANTENNA_2944 (.A(_08799_));
 sg13g2_antennanp ANTENNA_2945 (.A(_08799_));
 sg13g2_antennanp ANTENNA_2946 (.A(_08799_));
 sg13g2_antennanp ANTENNA_2947 (.A(_08799_));
 sg13g2_antennanp ANTENNA_2948 (.A(_08820_));
 sg13g2_antennanp ANTENNA_2949 (.A(_08820_));
 sg13g2_antennanp ANTENNA_2950 (.A(_08820_));
 sg13g2_antennanp ANTENNA_2951 (.A(_08820_));
 sg13g2_antennanp ANTENNA_2952 (.A(_08820_));
 sg13g2_antennanp ANTENNA_2953 (.A(_08820_));
 sg13g2_antennanp ANTENNA_2954 (.A(_08826_));
 sg13g2_antennanp ANTENNA_2955 (.A(_08826_));
 sg13g2_antennanp ANTENNA_2956 (.A(_08826_));
 sg13g2_antennanp ANTENNA_2957 (.A(_08826_));
 sg13g2_antennanp ANTENNA_2958 (.A(_08826_));
 sg13g2_antennanp ANTENNA_2959 (.A(_08826_));
 sg13g2_antennanp ANTENNA_2960 (.A(_08826_));
 sg13g2_antennanp ANTENNA_2961 (.A(_08826_));
 sg13g2_antennanp ANTENNA_2962 (.A(_08826_));
 sg13g2_antennanp ANTENNA_2963 (.A(_08848_));
 sg13g2_antennanp ANTENNA_2964 (.A(_08848_));
 sg13g2_antennanp ANTENNA_2965 (.A(_08848_));
 sg13g2_antennanp ANTENNA_2966 (.A(_08848_));
 sg13g2_antennanp ANTENNA_2967 (.A(_08848_));
 sg13g2_antennanp ANTENNA_2968 (.A(_08848_));
 sg13g2_antennanp ANTENNA_2969 (.A(_08848_));
 sg13g2_antennanp ANTENNA_2970 (.A(_08848_));
 sg13g2_antennanp ANTENNA_2971 (.A(_08848_));
 sg13g2_antennanp ANTENNA_2972 (.A(_08868_));
 sg13g2_antennanp ANTENNA_2973 (.A(_08900_));
 sg13g2_antennanp ANTENNA_2974 (.A(_08900_));
 sg13g2_antennanp ANTENNA_2975 (.A(_08900_));
 sg13g2_antennanp ANTENNA_2976 (.A(_08950_));
 sg13g2_antennanp ANTENNA_2977 (.A(_08950_));
 sg13g2_antennanp ANTENNA_2978 (.A(_08950_));
 sg13g2_antennanp ANTENNA_2979 (.A(_08950_));
 sg13g2_antennanp ANTENNA_2980 (.A(_08950_));
 sg13g2_antennanp ANTENNA_2981 (.A(_08950_));
 sg13g2_antennanp ANTENNA_2982 (.A(_08950_));
 sg13g2_antennanp ANTENNA_2983 (.A(_08950_));
 sg13g2_antennanp ANTENNA_2984 (.A(_08950_));
 sg13g2_antennanp ANTENNA_2985 (.A(_09002_));
 sg13g2_antennanp ANTENNA_2986 (.A(_09002_));
 sg13g2_antennanp ANTENNA_2987 (.A(_09065_));
 sg13g2_antennanp ANTENNA_2988 (.A(_09065_));
 sg13g2_antennanp ANTENNA_2989 (.A(_09091_));
 sg13g2_antennanp ANTENNA_2990 (.A(_09091_));
 sg13g2_antennanp ANTENNA_2991 (.A(_09091_));
 sg13g2_antennanp ANTENNA_2992 (.A(_09091_));
 sg13g2_antennanp ANTENNA_2993 (.A(_09091_));
 sg13g2_antennanp ANTENNA_2994 (.A(_09091_));
 sg13g2_antennanp ANTENNA_2995 (.A(_09091_));
 sg13g2_antennanp ANTENNA_2996 (.A(_09091_));
 sg13g2_antennanp ANTENNA_2997 (.A(_09091_));
 sg13g2_antennanp ANTENNA_2998 (.A(_09120_));
 sg13g2_antennanp ANTENNA_2999 (.A(_09120_));
 sg13g2_antennanp ANTENNA_3000 (.A(_09156_));
 sg13g2_antennanp ANTENNA_3001 (.A(_09156_));
 sg13g2_antennanp ANTENNA_3002 (.A(_09156_));
 sg13g2_antennanp ANTENNA_3003 (.A(_09156_));
 sg13g2_antennanp ANTENNA_3004 (.A(_09158_));
 sg13g2_antennanp ANTENNA_3005 (.A(_09158_));
 sg13g2_antennanp ANTENNA_3006 (.A(_09158_));
 sg13g2_antennanp ANTENNA_3007 (.A(_09173_));
 sg13g2_antennanp ANTENNA_3008 (.A(_09211_));
 sg13g2_antennanp ANTENNA_3009 (.A(_09211_));
 sg13g2_antennanp ANTENNA_3010 (.A(_09211_));
 sg13g2_antennanp ANTENNA_3011 (.A(_09211_));
 sg13g2_antennanp ANTENNA_3012 (.A(_09211_));
 sg13g2_antennanp ANTENNA_3013 (.A(_09218_));
 sg13g2_antennanp ANTENNA_3014 (.A(_09220_));
 sg13g2_antennanp ANTENNA_3015 (.A(_09220_));
 sg13g2_antennanp ANTENNA_3016 (.A(_09220_));
 sg13g2_antennanp ANTENNA_3017 (.A(_09220_));
 sg13g2_antennanp ANTENNA_3018 (.A(_09220_));
 sg13g2_antennanp ANTENNA_3019 (.A(_09220_));
 sg13g2_antennanp ANTENNA_3020 (.A(_09220_));
 sg13g2_antennanp ANTENNA_3021 (.A(_09220_));
 sg13g2_antennanp ANTENNA_3022 (.A(_09220_));
 sg13g2_antennanp ANTENNA_3023 (.A(_09220_));
 sg13g2_antennanp ANTENNA_3024 (.A(_09220_));
 sg13g2_antennanp ANTENNA_3025 (.A(_09220_));
 sg13g2_antennanp ANTENNA_3026 (.A(_09220_));
 sg13g2_antennanp ANTENNA_3027 (.A(_09240_));
 sg13g2_antennanp ANTENNA_3028 (.A(_09240_));
 sg13g2_antennanp ANTENNA_3029 (.A(_09240_));
 sg13g2_antennanp ANTENNA_3030 (.A(_09240_));
 sg13g2_antennanp ANTENNA_3031 (.A(_09240_));
 sg13g2_antennanp ANTENNA_3032 (.A(_09240_));
 sg13g2_antennanp ANTENNA_3033 (.A(_09240_));
 sg13g2_antennanp ANTENNA_3034 (.A(_09240_));
 sg13g2_antennanp ANTENNA_3035 (.A(_09298_));
 sg13g2_antennanp ANTENNA_3036 (.A(_09298_));
 sg13g2_antennanp ANTENNA_3037 (.A(_09298_));
 sg13g2_antennanp ANTENNA_3038 (.A(_09318_));
 sg13g2_antennanp ANTENNA_3039 (.A(_09318_));
 sg13g2_antennanp ANTENNA_3040 (.A(_09318_));
 sg13g2_antennanp ANTENNA_3041 (.A(_09394_));
 sg13g2_antennanp ANTENNA_3042 (.A(_09396_));
 sg13g2_antennanp ANTENNA_3043 (.A(_09447_));
 sg13g2_antennanp ANTENNA_3044 (.A(_09448_));
 sg13g2_antennanp ANTENNA_3045 (.A(_09448_));
 sg13g2_antennanp ANTENNA_3046 (.A(_09448_));
 sg13g2_antennanp ANTENNA_3047 (.A(_09448_));
 sg13g2_antennanp ANTENNA_3048 (.A(_09450_));
 sg13g2_antennanp ANTENNA_3049 (.A(_09492_));
 sg13g2_antennanp ANTENNA_3050 (.A(_09521_));
 sg13g2_antennanp ANTENNA_3051 (.A(_09544_));
 sg13g2_antennanp ANTENNA_3052 (.A(_09657_));
 sg13g2_antennanp ANTENNA_3053 (.A(_09722_));
 sg13g2_antennanp ANTENNA_3054 (.A(_09769_));
 sg13g2_antennanp ANTENNA_3055 (.A(_09791_));
 sg13g2_antennanp ANTENNA_3056 (.A(_09852_));
 sg13g2_antennanp ANTENNA_3057 (.A(_09852_));
 sg13g2_antennanp ANTENNA_3058 (.A(_09852_));
 sg13g2_antennanp ANTENNA_3059 (.A(_09852_));
 sg13g2_antennanp ANTENNA_3060 (.A(_09852_));
 sg13g2_antennanp ANTENNA_3061 (.A(_09852_));
 sg13g2_antennanp ANTENNA_3062 (.A(_09852_));
 sg13g2_antennanp ANTENNA_3063 (.A(_09852_));
 sg13g2_antennanp ANTENNA_3064 (.A(_09852_));
 sg13g2_antennanp ANTENNA_3065 (.A(_09852_));
 sg13g2_antennanp ANTENNA_3066 (.A(_09852_));
 sg13g2_antennanp ANTENNA_3067 (.A(_09852_));
 sg13g2_antennanp ANTENNA_3068 (.A(_09852_));
 sg13g2_antennanp ANTENNA_3069 (.A(_09852_));
 sg13g2_antennanp ANTENNA_3070 (.A(_09852_));
 sg13g2_antennanp ANTENNA_3071 (.A(_09852_));
 sg13g2_antennanp ANTENNA_3072 (.A(_10042_));
 sg13g2_antennanp ANTENNA_3073 (.A(_10042_));
 sg13g2_antennanp ANTENNA_3074 (.A(_10042_));
 sg13g2_antennanp ANTENNA_3075 (.A(_10121_));
 sg13g2_antennanp ANTENNA_3076 (.A(_10121_));
 sg13g2_antennanp ANTENNA_3077 (.A(_10121_));
 sg13g2_antennanp ANTENNA_3078 (.A(_10146_));
 sg13g2_antennanp ANTENNA_3079 (.A(_10146_));
 sg13g2_antennanp ANTENNA_3080 (.A(_10146_));
 sg13g2_antennanp ANTENNA_3081 (.A(_10146_));
 sg13g2_antennanp ANTENNA_3082 (.A(_10146_));
 sg13g2_antennanp ANTENNA_3083 (.A(_10146_));
 sg13g2_antennanp ANTENNA_3084 (.A(_10146_));
 sg13g2_antennanp ANTENNA_3085 (.A(_10146_));
 sg13g2_antennanp ANTENNA_3086 (.A(_10379_));
 sg13g2_antennanp ANTENNA_3087 (.A(_10379_));
 sg13g2_antennanp ANTENNA_3088 (.A(_10379_));
 sg13g2_antennanp ANTENNA_3089 (.A(_10642_));
 sg13g2_antennanp ANTENNA_3090 (.A(_10642_));
 sg13g2_antennanp ANTENNA_3091 (.A(_10642_));
 sg13g2_antennanp ANTENNA_3092 (.A(_10642_));
 sg13g2_antennanp ANTENNA_3093 (.A(_10642_));
 sg13g2_antennanp ANTENNA_3094 (.A(_10642_));
 sg13g2_antennanp ANTENNA_3095 (.A(_10642_));
 sg13g2_antennanp ANTENNA_3096 (.A(_10744_));
 sg13g2_antennanp ANTENNA_3097 (.A(_10744_));
 sg13g2_antennanp ANTENNA_3098 (.A(_10744_));
 sg13g2_antennanp ANTENNA_3099 (.A(_10744_));
 sg13g2_antennanp ANTENNA_3100 (.A(_11913_));
 sg13g2_antennanp ANTENNA_3101 (.A(_11913_));
 sg13g2_antennanp ANTENNA_3102 (.A(_11913_));
 sg13g2_antennanp ANTENNA_3103 (.A(_12205_));
 sg13g2_antennanp ANTENNA_3104 (.A(_12205_));
 sg13g2_antennanp ANTENNA_3105 (.A(_12205_));
 sg13g2_antennanp ANTENNA_3106 (.A(_12205_));
 sg13g2_antennanp ANTENNA_3107 (.A(_12218_));
 sg13g2_antennanp ANTENNA_3108 (.A(_12218_));
 sg13g2_antennanp ANTENNA_3109 (.A(_12218_));
 sg13g2_antennanp ANTENNA_3110 (.A(_12218_));
 sg13g2_antennanp ANTENNA_3111 (.A(_12218_));
 sg13g2_antennanp ANTENNA_3112 (.A(_12218_));
 sg13g2_antennanp ANTENNA_3113 (.A(_12218_));
 sg13g2_antennanp ANTENNA_3114 (.A(_12218_));
 sg13g2_antennanp ANTENNA_3115 (.A(_12218_));
 sg13g2_antennanp ANTENNA_3116 (.A(_12225_));
 sg13g2_antennanp ANTENNA_3117 (.A(_12225_));
 sg13g2_antennanp ANTENNA_3118 (.A(_12225_));
 sg13g2_antennanp ANTENNA_3119 (.A(_12225_));
 sg13g2_antennanp ANTENNA_3120 (.A(_12225_));
 sg13g2_antennanp ANTENNA_3121 (.A(_12225_));
 sg13g2_antennanp ANTENNA_3122 (.A(_12225_));
 sg13g2_antennanp ANTENNA_3123 (.A(_12225_));
 sg13g2_antennanp ANTENNA_3124 (.A(_12225_));
 sg13g2_antennanp ANTENNA_3125 (.A(_12236_));
 sg13g2_antennanp ANTENNA_3126 (.A(_12236_));
 sg13g2_antennanp ANTENNA_3127 (.A(_12236_));
 sg13g2_antennanp ANTENNA_3128 (.A(_12236_));
 sg13g2_antennanp ANTENNA_3129 (.A(_12236_));
 sg13g2_antennanp ANTENNA_3130 (.A(_12236_));
 sg13g2_antennanp ANTENNA_3131 (.A(_12236_));
 sg13g2_antennanp ANTENNA_3132 (.A(_12236_));
 sg13g2_antennanp ANTENNA_3133 (.A(_12236_));
 sg13g2_antennanp ANTENNA_3134 (.A(\cpu.dcache.wdata[9] ));
 sg13g2_antennanp ANTENNA_3135 (.A(\cpu.dcache.wdata[9] ));
 sg13g2_antennanp ANTENNA_3136 (.A(\cpu.dcache.wdata[9] ));
 sg13g2_antennanp ANTENNA_3137 (.A(\cpu.dcache.wdata[9] ));
 sg13g2_antennanp ANTENNA_3138 (.A(\cpu.ex.pc[1] ));
 sg13g2_antennanp ANTENNA_3139 (.A(\cpu.ex.pc[2] ));
 sg13g2_antennanp ANTENNA_3140 (.A(\cpu.gpio.uart_rx ));
 sg13g2_antennanp ANTENNA_3141 (.A(\cpu.gpio.uart_rx ));
 sg13g2_antennanp ANTENNA_3142 (.A(\cpu.qspi.c_wstrobe_i ));
 sg13g2_antennanp ANTENNA_3143 (.A(\cpu.qspi.c_wstrobe_i ));
 sg13g2_antennanp ANTENNA_3144 (.A(net3));
 sg13g2_antennanp ANTENNA_3145 (.A(net3));
 sg13g2_antennanp ANTENNA_3146 (.A(net3));
 sg13g2_antennanp ANTENNA_3147 (.A(net12));
 sg13g2_antennanp ANTENNA_3148 (.A(net12));
 sg13g2_antennanp ANTENNA_3149 (.A(net12));
 sg13g2_antennanp ANTENNA_3150 (.A(net13));
 sg13g2_antennanp ANTENNA_3151 (.A(net13));
 sg13g2_antennanp ANTENNA_3152 (.A(net13));
 sg13g2_antennanp ANTENNA_3153 (.A(net14));
 sg13g2_antennanp ANTENNA_3154 (.A(net14));
 sg13g2_antennanp ANTENNA_3155 (.A(net14));
 sg13g2_antennanp ANTENNA_3156 (.A(net114));
 sg13g2_antennanp ANTENNA_3157 (.A(net114));
 sg13g2_antennanp ANTENNA_3158 (.A(net114));
 sg13g2_antennanp ANTENNA_3159 (.A(net114));
 sg13g2_antennanp ANTENNA_3160 (.A(net114));
 sg13g2_antennanp ANTENNA_3161 (.A(net114));
 sg13g2_antennanp ANTENNA_3162 (.A(net114));
 sg13g2_antennanp ANTENNA_3163 (.A(net114));
 sg13g2_antennanp ANTENNA_3164 (.A(net452));
 sg13g2_antennanp ANTENNA_3165 (.A(net452));
 sg13g2_antennanp ANTENNA_3166 (.A(net452));
 sg13g2_antennanp ANTENNA_3167 (.A(net452));
 sg13g2_antennanp ANTENNA_3168 (.A(net452));
 sg13g2_antennanp ANTENNA_3169 (.A(net452));
 sg13g2_antennanp ANTENNA_3170 (.A(net452));
 sg13g2_antennanp ANTENNA_3171 (.A(net452));
 sg13g2_antennanp ANTENNA_3172 (.A(net491));
 sg13g2_antennanp ANTENNA_3173 (.A(net491));
 sg13g2_antennanp ANTENNA_3174 (.A(net491));
 sg13g2_antennanp ANTENNA_3175 (.A(net491));
 sg13g2_antennanp ANTENNA_3176 (.A(net491));
 sg13g2_antennanp ANTENNA_3177 (.A(net491));
 sg13g2_antennanp ANTENNA_3178 (.A(net491));
 sg13g2_antennanp ANTENNA_3179 (.A(net491));
 sg13g2_antennanp ANTENNA_3180 (.A(net491));
 sg13g2_antennanp ANTENNA_3181 (.A(net491));
 sg13g2_antennanp ANTENNA_3182 (.A(net491));
 sg13g2_antennanp ANTENNA_3183 (.A(net491));
 sg13g2_antennanp ANTENNA_3184 (.A(net686));
 sg13g2_antennanp ANTENNA_3185 (.A(net686));
 sg13g2_antennanp ANTENNA_3186 (.A(net686));
 sg13g2_antennanp ANTENNA_3187 (.A(net686));
 sg13g2_antennanp ANTENNA_3188 (.A(net686));
 sg13g2_antennanp ANTENNA_3189 (.A(net686));
 sg13g2_antennanp ANTENNA_3190 (.A(net686));
 sg13g2_antennanp ANTENNA_3191 (.A(net686));
 sg13g2_antennanp ANTENNA_3192 (.A(net708));
 sg13g2_antennanp ANTENNA_3193 (.A(net708));
 sg13g2_antennanp ANTENNA_3194 (.A(net708));
 sg13g2_antennanp ANTENNA_3195 (.A(net708));
 sg13g2_antennanp ANTENNA_3196 (.A(net708));
 sg13g2_antennanp ANTENNA_3197 (.A(net708));
 sg13g2_antennanp ANTENNA_3198 (.A(net708));
 sg13g2_antennanp ANTENNA_3199 (.A(net708));
 sg13g2_antennanp ANTENNA_3200 (.A(net708));
 sg13g2_antennanp ANTENNA_3201 (.A(net708));
 sg13g2_antennanp ANTENNA_3202 (.A(net708));
 sg13g2_antennanp ANTENNA_3203 (.A(net708));
 sg13g2_antennanp ANTENNA_3204 (.A(net708));
 sg13g2_antennanp ANTENNA_3205 (.A(net708));
 sg13g2_antennanp ANTENNA_3206 (.A(net708));
 sg13g2_antennanp ANTENNA_3207 (.A(net708));
 sg13g2_antennanp ANTENNA_3208 (.A(net745));
 sg13g2_antennanp ANTENNA_3209 (.A(net745));
 sg13g2_antennanp ANTENNA_3210 (.A(net745));
 sg13g2_antennanp ANTENNA_3211 (.A(net745));
 sg13g2_antennanp ANTENNA_3212 (.A(net745));
 sg13g2_antennanp ANTENNA_3213 (.A(net745));
 sg13g2_antennanp ANTENNA_3214 (.A(net745));
 sg13g2_antennanp ANTENNA_3215 (.A(net745));
 sg13g2_antennanp ANTENNA_3216 (.A(net803));
 sg13g2_antennanp ANTENNA_3217 (.A(net803));
 sg13g2_antennanp ANTENNA_3218 (.A(net803));
 sg13g2_antennanp ANTENNA_3219 (.A(net803));
 sg13g2_antennanp ANTENNA_3220 (.A(net803));
 sg13g2_antennanp ANTENNA_3221 (.A(net803));
 sg13g2_antennanp ANTENNA_3222 (.A(net803));
 sg13g2_antennanp ANTENNA_3223 (.A(net803));
 sg13g2_antennanp ANTENNA_3224 (.A(net858));
 sg13g2_antennanp ANTENNA_3225 (.A(net858));
 sg13g2_antennanp ANTENNA_3226 (.A(net858));
 sg13g2_antennanp ANTENNA_3227 (.A(net858));
 sg13g2_antennanp ANTENNA_3228 (.A(net858));
 sg13g2_antennanp ANTENNA_3229 (.A(net858));
 sg13g2_antennanp ANTENNA_3230 (.A(net858));
 sg13g2_antennanp ANTENNA_3231 (.A(net858));
 sg13g2_antennanp ANTENNA_3232 (.A(net858));
 sg13g2_antennanp ANTENNA_3233 (.A(net860));
 sg13g2_antennanp ANTENNA_3234 (.A(net860));
 sg13g2_antennanp ANTENNA_3235 (.A(net860));
 sg13g2_antennanp ANTENNA_3236 (.A(net860));
 sg13g2_antennanp ANTENNA_3237 (.A(net860));
 sg13g2_antennanp ANTENNA_3238 (.A(net860));
 sg13g2_antennanp ANTENNA_3239 (.A(net860));
 sg13g2_antennanp ANTENNA_3240 (.A(net860));
 sg13g2_antennanp ANTENNA_3241 (.A(net860));
 sg13g2_antennanp ANTENNA_3242 (.A(net872));
 sg13g2_antennanp ANTENNA_3243 (.A(net872));
 sg13g2_antennanp ANTENNA_3244 (.A(net872));
 sg13g2_antennanp ANTENNA_3245 (.A(net872));
 sg13g2_antennanp ANTENNA_3246 (.A(net872));
 sg13g2_antennanp ANTENNA_3247 (.A(net872));
 sg13g2_antennanp ANTENNA_3248 (.A(net872));
 sg13g2_antennanp ANTENNA_3249 (.A(net872));
 sg13g2_antennanp ANTENNA_3250 (.A(net872));
 sg13g2_antennanp ANTENNA_3251 (.A(net872));
 sg13g2_antennanp ANTENNA_3252 (.A(net872));
 sg13g2_antennanp ANTENNA_3253 (.A(net872));
 sg13g2_antennanp ANTENNA_3254 (.A(net872));
 sg13g2_antennanp ANTENNA_3255 (.A(net872));
 sg13g2_antennanp ANTENNA_3256 (.A(net872));
 sg13g2_antennanp ANTENNA_3257 (.A(net872));
 sg13g2_antennanp ANTENNA_3258 (.A(net872));
 sg13g2_antennanp ANTENNA_3259 (.A(net872));
 sg13g2_antennanp ANTENNA_3260 (.A(net872));
 sg13g2_antennanp ANTENNA_3261 (.A(net872));
 sg13g2_antennanp ANTENNA_3262 (.A(net872));
 sg13g2_antennanp ANTENNA_3263 (.A(net872));
 sg13g2_antennanp ANTENNA_3264 (.A(net872));
 sg13g2_antennanp ANTENNA_3265 (.A(net872));
 sg13g2_antennanp ANTENNA_3266 (.A(net872));
 sg13g2_antennanp ANTENNA_3267 (.A(net872));
 sg13g2_antennanp ANTENNA_3268 (.A(net872));
 sg13g2_antennanp ANTENNA_3269 (.A(net872));
 sg13g2_antennanp ANTENNA_3270 (.A(net872));
 sg13g2_antennanp ANTENNA_3271 (.A(net872));
 sg13g2_antennanp ANTENNA_3272 (.A(net872));
 sg13g2_antennanp ANTENNA_3273 (.A(net872));
 sg13g2_antennanp ANTENNA_3274 (.A(net872));
 sg13g2_antennanp ANTENNA_3275 (.A(net872));
 sg13g2_antennanp ANTENNA_3276 (.A(net872));
 sg13g2_antennanp ANTENNA_3277 (.A(net872));
 sg13g2_antennanp ANTENNA_3278 (.A(net872));
 sg13g2_antennanp ANTENNA_3279 (.A(net872));
 sg13g2_antennanp ANTENNA_3280 (.A(net872));
 sg13g2_antennanp ANTENNA_3281 (.A(net872));
 sg13g2_antennanp ANTENNA_3282 (.A(net872));
 sg13g2_antennanp ANTENNA_3283 (.A(net872));
 sg13g2_antennanp ANTENNA_3284 (.A(net872));
 sg13g2_antennanp ANTENNA_3285 (.A(net872));
 sg13g2_antennanp ANTENNA_3286 (.A(net872));
 sg13g2_antennanp ANTENNA_3287 (.A(net928));
 sg13g2_antennanp ANTENNA_3288 (.A(net928));
 sg13g2_antennanp ANTENNA_3289 (.A(net928));
 sg13g2_antennanp ANTENNA_3290 (.A(net928));
 sg13g2_antennanp ANTENNA_3291 (.A(net928));
 sg13g2_antennanp ANTENNA_3292 (.A(net928));
 sg13g2_antennanp ANTENNA_3293 (.A(net928));
 sg13g2_antennanp ANTENNA_3294 (.A(net928));
 sg13g2_antennanp ANTENNA_3295 (.A(net928));
 sg13g2_antennanp ANTENNA_3296 (.A(net928));
 sg13g2_antennanp ANTENNA_3297 (.A(net928));
 sg13g2_antennanp ANTENNA_3298 (.A(net928));
 sg13g2_antennanp ANTENNA_3299 (.A(net995));
 sg13g2_antennanp ANTENNA_3300 (.A(net995));
 sg13g2_antennanp ANTENNA_3301 (.A(net995));
 sg13g2_antennanp ANTENNA_3302 (.A(net995));
 sg13g2_antennanp ANTENNA_3303 (.A(net995));
 sg13g2_antennanp ANTENNA_3304 (.A(net995));
 sg13g2_antennanp ANTENNA_3305 (.A(net995));
 sg13g2_antennanp ANTENNA_3306 (.A(net995));
 sg13g2_antennanp ANTENNA_3307 (.A(net995));
 sg13g2_antennanp ANTENNA_3308 (.A(net1002));
 sg13g2_antennanp ANTENNA_3309 (.A(net1002));
 sg13g2_antennanp ANTENNA_3310 (.A(net1002));
 sg13g2_antennanp ANTENNA_3311 (.A(net1002));
 sg13g2_antennanp ANTENNA_3312 (.A(net1002));
 sg13g2_antennanp ANTENNA_3313 (.A(net1002));
 sg13g2_antennanp ANTENNA_3314 (.A(net1002));
 sg13g2_antennanp ANTENNA_3315 (.A(net1002));
 sg13g2_antennanp ANTENNA_3316 (.A(net1002));
 sg13g2_antennanp ANTENNA_3317 (.A(net1004));
 sg13g2_antennanp ANTENNA_3318 (.A(net1004));
 sg13g2_antennanp ANTENNA_3319 (.A(net1004));
 sg13g2_antennanp ANTENNA_3320 (.A(net1004));
 sg13g2_antennanp ANTENNA_3321 (.A(net1004));
 sg13g2_antennanp ANTENNA_3322 (.A(net1004));
 sg13g2_antennanp ANTENNA_3323 (.A(net1004));
 sg13g2_antennanp ANTENNA_3324 (.A(net1004));
 sg13g2_antennanp ANTENNA_3325 (.A(net1004));
 sg13g2_antennanp ANTENNA_3326 (.A(net1099));
 sg13g2_antennanp ANTENNA_3327 (.A(net1099));
 sg13g2_antennanp ANTENNA_3328 (.A(net1099));
 sg13g2_antennanp ANTENNA_3329 (.A(net1099));
 sg13g2_antennanp ANTENNA_3330 (.A(net1099));
 sg13g2_antennanp ANTENNA_3331 (.A(net1099));
 sg13g2_antennanp ANTENNA_3332 (.A(net1099));
 sg13g2_antennanp ANTENNA_3333 (.A(net1099));
 sg13g2_antennanp ANTENNA_3334 (.A(net1099));
 sg13g2_antennanp ANTENNA_3335 (.A(net1099));
 sg13g2_antennanp ANTENNA_3336 (.A(net1099));
 sg13g2_antennanp ANTENNA_3337 (.A(net1099));
 sg13g2_antennanp ANTENNA_3338 (.A(net1099));
 sg13g2_antennanp ANTENNA_3339 (.A(net1099));
 sg13g2_antennanp ANTENNA_3340 (.A(net1099));
 sg13g2_antennanp ANTENNA_3341 (.A(net1099));
 sg13g2_antennanp ANTENNA_3342 (.A(net1099));
 sg13g2_antennanp ANTENNA_3343 (.A(net1099));
 sg13g2_antennanp ANTENNA_3344 (.A(net1099));
 sg13g2_antennanp ANTENNA_3345 (.A(net1099));
 sg13g2_antennanp ANTENNA_3346 (.A(net1122));
 sg13g2_antennanp ANTENNA_3347 (.A(net1122));
 sg13g2_antennanp ANTENNA_3348 (.A(net1122));
 sg13g2_antennanp ANTENNA_3349 (.A(net1122));
 sg13g2_antennanp ANTENNA_3350 (.A(net1122));
 sg13g2_antennanp ANTENNA_3351 (.A(net1122));
 sg13g2_antennanp ANTENNA_3352 (.A(net1122));
 sg13g2_antennanp ANTENNA_3353 (.A(net1122));
 sg13g2_decap_8 FILLER_0_0 ();
 sg13g2_decap_8 FILLER_0_7 ();
 sg13g2_decap_8 FILLER_0_14 ();
 sg13g2_decap_8 FILLER_0_21 ();
 sg13g2_decap_8 FILLER_0_28 ();
 sg13g2_decap_8 FILLER_0_35 ();
 sg13g2_decap_8 FILLER_0_42 ();
 sg13g2_decap_8 FILLER_0_49 ();
 sg13g2_decap_8 FILLER_0_56 ();
 sg13g2_decap_8 FILLER_0_63 ();
 sg13g2_decap_8 FILLER_0_70 ();
 sg13g2_decap_8 FILLER_0_77 ();
 sg13g2_fill_2 FILLER_0_110 ();
 sg13g2_fill_1 FILLER_0_112 ();
 sg13g2_decap_8 FILLER_0_121 ();
 sg13g2_decap_8 FILLER_0_128 ();
 sg13g2_decap_8 FILLER_0_135 ();
 sg13g2_fill_2 FILLER_0_142 ();
 sg13g2_decap_8 FILLER_0_170 ();
 sg13g2_decap_8 FILLER_0_177 ();
 sg13g2_decap_8 FILLER_0_184 ();
 sg13g2_decap_4 FILLER_0_191 ();
 sg13g2_fill_2 FILLER_0_195 ();
 sg13g2_decap_8 FILLER_0_201 ();
 sg13g2_decap_8 FILLER_0_208 ();
 sg13g2_fill_2 FILLER_0_215 ();
 sg13g2_fill_1 FILLER_0_217 ();
 sg13g2_decap_8 FILLER_0_222 ();
 sg13g2_fill_1 FILLER_0_229 ();
 sg13g2_decap_8 FILLER_0_267 ();
 sg13g2_decap_8 FILLER_0_274 ();
 sg13g2_decap_4 FILLER_0_281 ();
 sg13g2_decap_4 FILLER_0_311 ();
 sg13g2_fill_2 FILLER_0_315 ();
 sg13g2_fill_1 FILLER_0_349 ();
 sg13g2_fill_2 FILLER_0_356 ();
 sg13g2_decap_8 FILLER_0_396 ();
 sg13g2_decap_8 FILLER_0_403 ();
 sg13g2_decap_8 FILLER_0_410 ();
 sg13g2_decap_8 FILLER_0_417 ();
 sg13g2_decap_8 FILLER_0_424 ();
 sg13g2_decap_8 FILLER_0_431 ();
 sg13g2_decap_8 FILLER_0_438 ();
 sg13g2_decap_8 FILLER_0_445 ();
 sg13g2_decap_4 FILLER_0_452 ();
 sg13g2_fill_1 FILLER_0_456 ();
 sg13g2_decap_8 FILLER_0_461 ();
 sg13g2_decap_8 FILLER_0_468 ();
 sg13g2_decap_8 FILLER_0_475 ();
 sg13g2_decap_8 FILLER_0_486 ();
 sg13g2_decap_8 FILLER_0_519 ();
 sg13g2_decap_8 FILLER_0_526 ();
 sg13g2_decap_8 FILLER_0_533 ();
 sg13g2_decap_8 FILLER_0_570 ();
 sg13g2_decap_8 FILLER_0_577 ();
 sg13g2_decap_8 FILLER_0_584 ();
 sg13g2_fill_1 FILLER_0_591 ();
 sg13g2_decap_8 FILLER_0_596 ();
 sg13g2_decap_8 FILLER_0_603 ();
 sg13g2_decap_8 FILLER_0_610 ();
 sg13g2_fill_2 FILLER_0_617 ();
 sg13g2_decap_8 FILLER_0_623 ();
 sg13g2_decap_4 FILLER_0_630 ();
 sg13g2_fill_2 FILLER_0_634 ();
 sg13g2_decap_4 FILLER_0_641 ();
 sg13g2_fill_1 FILLER_0_645 ();
 sg13g2_decap_8 FILLER_0_651 ();
 sg13g2_fill_1 FILLER_0_662 ();
 sg13g2_fill_2 FILLER_0_667 ();
 sg13g2_decap_8 FILLER_0_681 ();
 sg13g2_decap_8 FILLER_0_688 ();
 sg13g2_fill_2 FILLER_0_695 ();
 sg13g2_fill_1 FILLER_0_697 ();
 sg13g2_decap_8 FILLER_0_710 ();
 sg13g2_decap_8 FILLER_0_717 ();
 sg13g2_decap_8 FILLER_0_724 ();
 sg13g2_decap_8 FILLER_0_731 ();
 sg13g2_decap_8 FILLER_0_738 ();
 sg13g2_fill_2 FILLER_0_745 ();
 sg13g2_decap_8 FILLER_0_751 ();
 sg13g2_decap_8 FILLER_0_758 ();
 sg13g2_decap_8 FILLER_0_765 ();
 sg13g2_decap_4 FILLER_0_772 ();
 sg13g2_decap_8 FILLER_0_780 ();
 sg13g2_decap_8 FILLER_0_787 ();
 sg13g2_decap_8 FILLER_0_794 ();
 sg13g2_decap_8 FILLER_0_801 ();
 sg13g2_decap_4 FILLER_0_808 ();
 sg13g2_decap_8 FILLER_0_816 ();
 sg13g2_fill_1 FILLER_0_853 ();
 sg13g2_decap_8 FILLER_0_864 ();
 sg13g2_decap_8 FILLER_0_871 ();
 sg13g2_decap_8 FILLER_0_878 ();
 sg13g2_fill_2 FILLER_0_885 ();
 sg13g2_fill_1 FILLER_0_887 ();
 sg13g2_decap_8 FILLER_0_898 ();
 sg13g2_fill_2 FILLER_0_905 ();
 sg13g2_fill_1 FILLER_0_907 ();
 sg13g2_decap_8 FILLER_0_934 ();
 sg13g2_decap_8 FILLER_0_977 ();
 sg13g2_decap_8 FILLER_0_984 ();
 sg13g2_decap_8 FILLER_0_991 ();
 sg13g2_decap_4 FILLER_0_998 ();
 sg13g2_fill_2 FILLER_0_1002 ();
 sg13g2_fill_2 FILLER_0_1013 ();
 sg13g2_fill_1 FILLER_0_1015 ();
 sg13g2_decap_8 FILLER_0_1020 ();
 sg13g2_decap_4 FILLER_0_1027 ();
 sg13g2_decap_8 FILLER_0_1035 ();
 sg13g2_decap_4 FILLER_0_1042 ();
 sg13g2_fill_1 FILLER_0_1046 ();
 sg13g2_fill_2 FILLER_0_1051 ();
 sg13g2_decap_8 FILLER_0_1075 ();
 sg13g2_decap_8 FILLER_0_1082 ();
 sg13g2_decap_8 FILLER_0_1089 ();
 sg13g2_decap_8 FILLER_0_1096 ();
 sg13g2_fill_2 FILLER_0_1103 ();
 sg13g2_decap_4 FILLER_0_1109 ();
 sg13g2_fill_1 FILLER_0_1113 ();
 sg13g2_decap_8 FILLER_0_1144 ();
 sg13g2_decap_8 FILLER_0_1151 ();
 sg13g2_decap_4 FILLER_0_1158 ();
 sg13g2_decap_8 FILLER_0_1193 ();
 sg13g2_decap_4 FILLER_0_1200 ();
 sg13g2_fill_1 FILLER_0_1204 ();
 sg13g2_fill_2 FILLER_0_1214 ();
 sg13g2_decap_8 FILLER_0_1237 ();
 sg13g2_decap_8 FILLER_0_1244 ();
 sg13g2_fill_1 FILLER_0_1251 ();
 sg13g2_fill_2 FILLER_0_1257 ();
 sg13g2_fill_1 FILLER_0_1259 ();
 sg13g2_decap_4 FILLER_0_1264 ();
 sg13g2_fill_2 FILLER_0_1268 ();
 sg13g2_fill_2 FILLER_0_1274 ();
 sg13g2_decap_4 FILLER_0_1280 ();
 sg13g2_fill_1 FILLER_0_1284 ();
 sg13g2_decap_8 FILLER_0_1289 ();
 sg13g2_decap_8 FILLER_0_1296 ();
 sg13g2_decap_8 FILLER_0_1303 ();
 sg13g2_decap_8 FILLER_0_1310 ();
 sg13g2_fill_2 FILLER_0_1326 ();
 sg13g2_fill_1 FILLER_0_1328 ();
 sg13g2_fill_1 FILLER_0_1334 ();
 sg13g2_decap_4 FILLER_0_1339 ();
 sg13g2_fill_2 FILLER_0_1343 ();
 sg13g2_decap_8 FILLER_0_1349 ();
 sg13g2_decap_8 FILLER_0_1356 ();
 sg13g2_decap_8 FILLER_0_1363 ();
 sg13g2_decap_8 FILLER_0_1370 ();
 sg13g2_decap_8 FILLER_0_1377 ();
 sg13g2_fill_2 FILLER_0_1384 ();
 sg13g2_fill_1 FILLER_0_1386 ();
 sg13g2_decap_8 FILLER_0_1413 ();
 sg13g2_decap_8 FILLER_0_1420 ();
 sg13g2_decap_8 FILLER_0_1427 ();
 sg13g2_decap_8 FILLER_0_1434 ();
 sg13g2_decap_4 FILLER_0_1441 ();
 sg13g2_fill_1 FILLER_0_1445 ();
 sg13g2_decap_8 FILLER_0_1472 ();
 sg13g2_decap_8 FILLER_0_1505 ();
 sg13g2_decap_8 FILLER_0_1512 ();
 sg13g2_decap_8 FILLER_0_1519 ();
 sg13g2_decap_8 FILLER_0_1526 ();
 sg13g2_decap_4 FILLER_0_1533 ();
 sg13g2_decap_8 FILLER_0_1541 ();
 sg13g2_decap_8 FILLER_0_1548 ();
 sg13g2_decap_4 FILLER_0_1555 ();
 sg13g2_fill_1 FILLER_0_1559 ();
 sg13g2_decap_8 FILLER_0_1599 ();
 sg13g2_decap_8 FILLER_0_1606 ();
 sg13g2_decap_8 FILLER_0_1613 ();
 sg13g2_decap_8 FILLER_0_1620 ();
 sg13g2_decap_8 FILLER_0_1627 ();
 sg13g2_decap_8 FILLER_0_1634 ();
 sg13g2_decap_8 FILLER_0_1641 ();
 sg13g2_decap_8 FILLER_0_1648 ();
 sg13g2_decap_4 FILLER_0_1655 ();
 sg13g2_decap_8 FILLER_0_1685 ();
 sg13g2_fill_2 FILLER_0_1692 ();
 sg13g2_fill_1 FILLER_0_1694 ();
 sg13g2_decap_8 FILLER_0_1699 ();
 sg13g2_decap_8 FILLER_0_1706 ();
 sg13g2_decap_8 FILLER_0_1713 ();
 sg13g2_decap_8 FILLER_0_1720 ();
 sg13g2_decap_8 FILLER_0_1727 ();
 sg13g2_decap_4 FILLER_0_1734 ();
 sg13g2_fill_2 FILLER_0_1738 ();
 sg13g2_decap_8 FILLER_0_1744 ();
 sg13g2_decap_4 FILLER_0_1761 ();
 sg13g2_decap_8 FILLER_0_1769 ();
 sg13g2_decap_8 FILLER_0_1776 ();
 sg13g2_decap_8 FILLER_0_1783 ();
 sg13g2_decap_8 FILLER_0_1790 ();
 sg13g2_decap_8 FILLER_0_1797 ();
 sg13g2_decap_8 FILLER_0_1804 ();
 sg13g2_decap_8 FILLER_0_1811 ();
 sg13g2_decap_8 FILLER_0_1818 ();
 sg13g2_decap_8 FILLER_0_1825 ();
 sg13g2_decap_8 FILLER_0_1832 ();
 sg13g2_decap_8 FILLER_0_1839 ();
 sg13g2_decap_8 FILLER_0_1846 ();
 sg13g2_decap_8 FILLER_0_1853 ();
 sg13g2_decap_8 FILLER_0_1860 ();
 sg13g2_decap_8 FILLER_0_1867 ();
 sg13g2_decap_8 FILLER_0_1874 ();
 sg13g2_decap_8 FILLER_0_1881 ();
 sg13g2_decap_8 FILLER_0_1888 ();
 sg13g2_decap_4 FILLER_0_1895 ();
 sg13g2_fill_2 FILLER_0_1899 ();
 sg13g2_decap_8 FILLER_0_1927 ();
 sg13g2_decap_8 FILLER_0_1934 ();
 sg13g2_decap_8 FILLER_0_1941 ();
 sg13g2_decap_8 FILLER_0_1948 ();
 sg13g2_decap_8 FILLER_0_1955 ();
 sg13g2_decap_8 FILLER_0_1962 ();
 sg13g2_decap_4 FILLER_0_1969 ();
 sg13g2_fill_1 FILLER_0_1973 ();
 sg13g2_fill_2 FILLER_0_1992 ();
 sg13g2_fill_1 FILLER_0_1994 ();
 sg13g2_decap_4 FILLER_0_1999 ();
 sg13g2_fill_2 FILLER_0_2003 ();
 sg13g2_decap_8 FILLER_0_2015 ();
 sg13g2_decap_8 FILLER_0_2022 ();
 sg13g2_decap_8 FILLER_0_2029 ();
 sg13g2_decap_8 FILLER_0_2036 ();
 sg13g2_decap_8 FILLER_0_2043 ();
 sg13g2_decap_8 FILLER_0_2050 ();
 sg13g2_decap_8 FILLER_0_2057 ();
 sg13g2_decap_8 FILLER_0_2064 ();
 sg13g2_fill_2 FILLER_0_2071 ();
 sg13g2_decap_8 FILLER_0_2106 ();
 sg13g2_decap_8 FILLER_0_2113 ();
 sg13g2_decap_8 FILLER_0_2120 ();
 sg13g2_decap_8 FILLER_0_2127 ();
 sg13g2_decap_4 FILLER_0_2134 ();
 sg13g2_fill_2 FILLER_0_2138 ();
 sg13g2_decap_8 FILLER_0_2144 ();
 sg13g2_decap_8 FILLER_0_2151 ();
 sg13g2_decap_8 FILLER_0_2158 ();
 sg13g2_decap_8 FILLER_0_2165 ();
 sg13g2_decap_8 FILLER_0_2172 ();
 sg13g2_decap_4 FILLER_0_2179 ();
 sg13g2_decap_8 FILLER_0_2204 ();
 sg13g2_decap_8 FILLER_0_2211 ();
 sg13g2_decap_8 FILLER_0_2218 ();
 sg13g2_decap_8 FILLER_0_2225 ();
 sg13g2_decap_8 FILLER_0_2232 ();
 sg13g2_decap_4 FILLER_0_2239 ();
 sg13g2_fill_2 FILLER_0_2243 ();
 sg13g2_decap_8 FILLER_0_2269 ();
 sg13g2_decap_8 FILLER_0_2276 ();
 sg13g2_decap_8 FILLER_0_2283 ();
 sg13g2_decap_8 FILLER_0_2290 ();
 sg13g2_decap_8 FILLER_0_2297 ();
 sg13g2_decap_8 FILLER_0_2304 ();
 sg13g2_decap_8 FILLER_0_2311 ();
 sg13g2_decap_8 FILLER_0_2318 ();
 sg13g2_decap_8 FILLER_0_2325 ();
 sg13g2_decap_8 FILLER_0_2332 ();
 sg13g2_decap_8 FILLER_0_2339 ();
 sg13g2_decap_8 FILLER_0_2346 ();
 sg13g2_decap_8 FILLER_0_2353 ();
 sg13g2_decap_8 FILLER_0_2360 ();
 sg13g2_decap_8 FILLER_0_2367 ();
 sg13g2_decap_8 FILLER_0_2374 ();
 sg13g2_decap_8 FILLER_0_2381 ();
 sg13g2_decap_8 FILLER_0_2388 ();
 sg13g2_decap_8 FILLER_0_2395 ();
 sg13g2_decap_8 FILLER_0_2402 ();
 sg13g2_decap_8 FILLER_0_2409 ();
 sg13g2_decap_8 FILLER_0_2416 ();
 sg13g2_decap_8 FILLER_0_2423 ();
 sg13g2_decap_8 FILLER_0_2430 ();
 sg13g2_decap_8 FILLER_0_2437 ();
 sg13g2_decap_8 FILLER_0_2444 ();
 sg13g2_decap_8 FILLER_0_2451 ();
 sg13g2_decap_8 FILLER_0_2458 ();
 sg13g2_decap_8 FILLER_0_2465 ();
 sg13g2_decap_8 FILLER_0_2472 ();
 sg13g2_decap_8 FILLER_0_2479 ();
 sg13g2_decap_8 FILLER_0_2486 ();
 sg13g2_decap_8 FILLER_0_2493 ();
 sg13g2_decap_8 FILLER_0_2500 ();
 sg13g2_decap_8 FILLER_0_2507 ();
 sg13g2_decap_8 FILLER_0_2514 ();
 sg13g2_decap_8 FILLER_0_2521 ();
 sg13g2_decap_8 FILLER_0_2528 ();
 sg13g2_decap_8 FILLER_0_2535 ();
 sg13g2_decap_8 FILLER_0_2542 ();
 sg13g2_decap_8 FILLER_0_2549 ();
 sg13g2_decap_8 FILLER_0_2556 ();
 sg13g2_decap_8 FILLER_0_2563 ();
 sg13g2_decap_8 FILLER_0_2570 ();
 sg13g2_decap_8 FILLER_0_2577 ();
 sg13g2_decap_8 FILLER_0_2584 ();
 sg13g2_decap_8 FILLER_0_2591 ();
 sg13g2_decap_8 FILLER_0_2598 ();
 sg13g2_decap_8 FILLER_0_2605 ();
 sg13g2_decap_8 FILLER_0_2612 ();
 sg13g2_decap_8 FILLER_0_2619 ();
 sg13g2_decap_8 FILLER_0_2626 ();
 sg13g2_decap_8 FILLER_0_2633 ();
 sg13g2_decap_8 FILLER_0_2640 ();
 sg13g2_decap_8 FILLER_0_2647 ();
 sg13g2_decap_8 FILLER_0_2654 ();
 sg13g2_decap_8 FILLER_0_2661 ();
 sg13g2_fill_2 FILLER_0_2668 ();
 sg13g2_decap_8 FILLER_1_0 ();
 sg13g2_decap_8 FILLER_1_7 ();
 sg13g2_decap_8 FILLER_1_14 ();
 sg13g2_decap_8 FILLER_1_21 ();
 sg13g2_decap_8 FILLER_1_28 ();
 sg13g2_decap_8 FILLER_1_35 ();
 sg13g2_decap_8 FILLER_1_42 ();
 sg13g2_decap_8 FILLER_1_49 ();
 sg13g2_decap_8 FILLER_1_56 ();
 sg13g2_decap_8 FILLER_1_63 ();
 sg13g2_decap_8 FILLER_1_70 ();
 sg13g2_decap_8 FILLER_1_77 ();
 sg13g2_decap_8 FILLER_1_84 ();
 sg13g2_fill_2 FILLER_1_95 ();
 sg13g2_decap_8 FILLER_1_103 ();
 sg13g2_decap_4 FILLER_1_136 ();
 sg13g2_fill_1 FILLER_1_140 ();
 sg13g2_fill_1 FILLER_1_151 ();
 sg13g2_decap_4 FILLER_1_182 ();
 sg13g2_fill_1 FILLER_1_190 ();
 sg13g2_fill_2 FILLER_1_217 ();
 sg13g2_decap_4 FILLER_1_272 ();
 sg13g2_fill_1 FILLER_1_276 ();
 sg13g2_fill_1 FILLER_1_342 ();
 sg13g2_decap_8 FILLER_1_427 ();
 sg13g2_fill_2 FILLER_1_434 ();
 sg13g2_fill_1 FILLER_1_436 ();
 sg13g2_fill_2 FILLER_1_472 ();
 sg13g2_fill_1 FILLER_1_474 ();
 sg13g2_decap_4 FILLER_1_505 ();
 sg13g2_fill_2 FILLER_1_509 ();
 sg13g2_decap_8 FILLER_1_537 ();
 sg13g2_fill_2 FILLER_1_544 ();
 sg13g2_fill_1 FILLER_1_546 ();
 sg13g2_decap_4 FILLER_1_551 ();
 sg13g2_fill_2 FILLER_1_555 ();
 sg13g2_fill_2 FILLER_1_583 ();
 sg13g2_fill_1 FILLER_1_585 ();
 sg13g2_fill_1 FILLER_1_638 ();
 sg13g2_fill_1 FILLER_1_649 ();
 sg13g2_fill_1 FILLER_1_732 ();
 sg13g2_fill_2 FILLER_1_738 ();
 sg13g2_fill_1 FILLER_1_766 ();
 sg13g2_decap_8 FILLER_1_793 ();
 sg13g2_fill_2 FILLER_1_800 ();
 sg13g2_fill_1 FILLER_1_802 ();
 sg13g2_fill_2 FILLER_1_829 ();
 sg13g2_fill_1 FILLER_1_831 ();
 sg13g2_fill_2 FILLER_1_842 ();
 sg13g2_fill_2 FILLER_1_904 ();
 sg13g2_fill_1 FILLER_1_916 ();
 sg13g2_fill_1 FILLER_1_943 ();
 sg13g2_fill_1 FILLER_1_954 ();
 sg13g2_fill_2 FILLER_1_981 ();
 sg13g2_fill_1 FILLER_1_1039 ();
 sg13g2_decap_4 FILLER_1_1080 ();
 sg13g2_fill_2 FILLER_1_1097 ();
 sg13g2_fill_1 FILLER_1_1099 ();
 sg13g2_fill_1 FILLER_1_1109 ();
 sg13g2_fill_2 FILLER_1_1115 ();
 sg13g2_fill_2 FILLER_1_1122 ();
 sg13g2_fill_2 FILLER_1_1145 ();
 sg13g2_fill_1 FILLER_1_1147 ();
 sg13g2_fill_1 FILLER_1_1157 ();
 sg13g2_fill_1 FILLER_1_1183 ();
 sg13g2_decap_8 FILLER_1_1188 ();
 sg13g2_fill_1 FILLER_1_1195 ();
 sg13g2_fill_2 FILLER_1_1288 ();
 sg13g2_fill_1 FILLER_1_1290 ();
 sg13g2_fill_2 FILLER_1_1317 ();
 sg13g2_fill_2 FILLER_1_1323 ();
 sg13g2_fill_2 FILLER_1_1329 ();
 sg13g2_fill_1 FILLER_1_1335 ();
 sg13g2_decap_4 FILLER_1_1362 ();
 sg13g2_fill_2 FILLER_1_1366 ();
 sg13g2_fill_2 FILLER_1_1438 ();
 sg13g2_decap_8 FILLER_1_1502 ();
 sg13g2_fill_2 FILLER_1_1509 ();
 sg13g2_fill_2 FILLER_1_1541 ();
 sg13g2_fill_1 FILLER_1_1543 ();
 sg13g2_fill_2 FILLER_1_1574 ();
 sg13g2_fill_1 FILLER_1_1576 ();
 sg13g2_fill_2 FILLER_1_1629 ();
 sg13g2_decap_8 FILLER_1_1713 ();
 sg13g2_decap_8 FILLER_1_1720 ();
 sg13g2_decap_4 FILLER_1_1727 ();
 sg13g2_fill_1 FILLER_1_1783 ();
 sg13g2_decap_8 FILLER_1_1788 ();
 sg13g2_decap_8 FILLER_1_1821 ();
 sg13g2_decap_8 FILLER_1_1828 ();
 sg13g2_decap_8 FILLER_1_1835 ();
 sg13g2_decap_8 FILLER_1_1842 ();
 sg13g2_decap_4 FILLER_1_1849 ();
 sg13g2_fill_1 FILLER_1_1853 ();
 sg13g2_decap_8 FILLER_1_1936 ();
 sg13g2_decap_8 FILLER_1_1943 ();
 sg13g2_fill_2 FILLER_1_1950 ();
 sg13g2_decap_4 FILLER_1_2030 ();
 sg13g2_fill_1 FILLER_1_2034 ();
 sg13g2_fill_2 FILLER_1_2079 ();
 sg13g2_decap_8 FILLER_1_2283 ();
 sg13g2_decap_8 FILLER_1_2290 ();
 sg13g2_decap_8 FILLER_1_2297 ();
 sg13g2_decap_8 FILLER_1_2304 ();
 sg13g2_decap_8 FILLER_1_2311 ();
 sg13g2_decap_8 FILLER_1_2318 ();
 sg13g2_decap_8 FILLER_1_2325 ();
 sg13g2_decap_8 FILLER_1_2332 ();
 sg13g2_decap_8 FILLER_1_2339 ();
 sg13g2_decap_8 FILLER_1_2346 ();
 sg13g2_decap_8 FILLER_1_2353 ();
 sg13g2_decap_8 FILLER_1_2360 ();
 sg13g2_decap_8 FILLER_1_2367 ();
 sg13g2_decap_4 FILLER_1_2374 ();
 sg13g2_fill_2 FILLER_1_2378 ();
 sg13g2_fill_2 FILLER_1_2383 ();
 sg13g2_fill_1 FILLER_1_2385 ();
 sg13g2_decap_8 FILLER_1_2392 ();
 sg13g2_decap_8 FILLER_1_2399 ();
 sg13g2_decap_8 FILLER_1_2406 ();
 sg13g2_decap_8 FILLER_1_2413 ();
 sg13g2_decap_8 FILLER_1_2420 ();
 sg13g2_decap_8 FILLER_1_2427 ();
 sg13g2_decap_8 FILLER_1_2434 ();
 sg13g2_decap_8 FILLER_1_2441 ();
 sg13g2_decap_8 FILLER_1_2448 ();
 sg13g2_decap_8 FILLER_1_2455 ();
 sg13g2_decap_8 FILLER_1_2462 ();
 sg13g2_decap_8 FILLER_1_2469 ();
 sg13g2_decap_8 FILLER_1_2476 ();
 sg13g2_decap_8 FILLER_1_2483 ();
 sg13g2_decap_8 FILLER_1_2490 ();
 sg13g2_decap_8 FILLER_1_2497 ();
 sg13g2_decap_8 FILLER_1_2504 ();
 sg13g2_decap_8 FILLER_1_2511 ();
 sg13g2_decap_8 FILLER_1_2518 ();
 sg13g2_decap_8 FILLER_1_2525 ();
 sg13g2_decap_8 FILLER_1_2532 ();
 sg13g2_decap_8 FILLER_1_2539 ();
 sg13g2_decap_8 FILLER_1_2546 ();
 sg13g2_decap_8 FILLER_1_2553 ();
 sg13g2_decap_8 FILLER_1_2560 ();
 sg13g2_decap_8 FILLER_1_2567 ();
 sg13g2_decap_8 FILLER_1_2574 ();
 sg13g2_decap_8 FILLER_1_2581 ();
 sg13g2_decap_8 FILLER_1_2588 ();
 sg13g2_decap_8 FILLER_1_2595 ();
 sg13g2_decap_8 FILLER_1_2602 ();
 sg13g2_decap_8 FILLER_1_2609 ();
 sg13g2_decap_8 FILLER_1_2616 ();
 sg13g2_decap_8 FILLER_1_2623 ();
 sg13g2_decap_8 FILLER_1_2630 ();
 sg13g2_decap_8 FILLER_1_2637 ();
 sg13g2_decap_8 FILLER_1_2644 ();
 sg13g2_decap_8 FILLER_1_2651 ();
 sg13g2_decap_8 FILLER_1_2658 ();
 sg13g2_decap_4 FILLER_1_2665 ();
 sg13g2_fill_1 FILLER_1_2669 ();
 sg13g2_decap_8 FILLER_2_0 ();
 sg13g2_decap_8 FILLER_2_7 ();
 sg13g2_decap_8 FILLER_2_14 ();
 sg13g2_decap_8 FILLER_2_21 ();
 sg13g2_decap_8 FILLER_2_28 ();
 sg13g2_decap_8 FILLER_2_35 ();
 sg13g2_decap_8 FILLER_2_42 ();
 sg13g2_decap_8 FILLER_2_49 ();
 sg13g2_decap_8 FILLER_2_56 ();
 sg13g2_fill_1 FILLER_2_63 ();
 sg13g2_fill_2 FILLER_2_107 ();
 sg13g2_decap_8 FILLER_2_162 ();
 sg13g2_fill_2 FILLER_2_169 ();
 sg13g2_fill_1 FILLER_2_171 ();
 sg13g2_fill_2 FILLER_2_198 ();
 sg13g2_decap_4 FILLER_2_205 ();
 sg13g2_fill_2 FILLER_2_209 ();
 sg13g2_fill_1 FILLER_2_255 ();
 sg13g2_fill_1 FILLER_2_262 ();
 sg13g2_decap_4 FILLER_2_277 ();
 sg13g2_fill_1 FILLER_2_281 ();
 sg13g2_fill_2 FILLER_2_296 ();
 sg13g2_fill_1 FILLER_2_308 ();
 sg13g2_fill_1 FILLER_2_314 ();
 sg13g2_fill_1 FILLER_2_320 ();
 sg13g2_fill_1 FILLER_2_325 ();
 sg13g2_fill_1 FILLER_2_352 ();
 sg13g2_fill_1 FILLER_2_360 ();
 sg13g2_fill_1 FILLER_2_378 ();
 sg13g2_decap_8 FILLER_2_420 ();
 sg13g2_decap_8 FILLER_2_427 ();
 sg13g2_decap_4 FILLER_2_434 ();
 sg13g2_fill_2 FILLER_2_464 ();
 sg13g2_fill_2 FILLER_2_471 ();
 sg13g2_fill_1 FILLER_2_473 ();
 sg13g2_fill_1 FILLER_2_500 ();
 sg13g2_fill_2 FILLER_2_506 ();
 sg13g2_fill_1 FILLER_2_508 ();
 sg13g2_fill_2 FILLER_2_522 ();
 sg13g2_fill_2 FILLER_2_544 ();
 sg13g2_fill_2 FILLER_2_565 ();
 sg13g2_fill_1 FILLER_2_595 ();
 sg13g2_fill_2 FILLER_2_616 ();
 sg13g2_fill_2 FILLER_2_649 ();
 sg13g2_fill_1 FILLER_2_651 ();
 sg13g2_fill_1 FILLER_2_657 ();
 sg13g2_fill_1 FILLER_2_663 ();
 sg13g2_fill_2 FILLER_2_698 ();
 sg13g2_decap_4 FILLER_2_730 ();
 sg13g2_fill_1 FILLER_2_765 ();
 sg13g2_decap_8 FILLER_2_776 ();
 sg13g2_fill_2 FILLER_2_783 ();
 sg13g2_fill_1 FILLER_2_785 ();
 sg13g2_fill_2 FILLER_2_812 ();
 sg13g2_fill_1 FILLER_2_814 ();
 sg13g2_fill_2 FILLER_2_841 ();
 sg13g2_fill_1 FILLER_2_843 ();
 sg13g2_fill_2 FILLER_2_901 ();
 sg13g2_fill_1 FILLER_2_903 ();
 sg13g2_decap_4 FILLER_2_956 ();
 sg13g2_fill_2 FILLER_2_964 ();
 sg13g2_decap_8 FILLER_2_970 ();
 sg13g2_decap_4 FILLER_2_977 ();
 sg13g2_fill_2 FILLER_2_981 ();
 sg13g2_fill_2 FILLER_2_987 ();
 sg13g2_fill_1 FILLER_2_989 ();
 sg13g2_fill_2 FILLER_2_995 ();
 sg13g2_fill_1 FILLER_2_997 ();
 sg13g2_fill_1 FILLER_2_1002 ();
 sg13g2_fill_2 FILLER_2_1138 ();
 sg13g2_fill_2 FILLER_2_1288 ();
 sg13g2_fill_2 FILLER_2_1295 ();
 sg13g2_fill_1 FILLER_2_1297 ();
 sg13g2_fill_1 FILLER_2_1302 ();
 sg13g2_fill_1 FILLER_2_1334 ();
 sg13g2_fill_2 FILLER_2_1361 ();
 sg13g2_fill_2 FILLER_2_1368 ();
 sg13g2_fill_1 FILLER_2_1403 ();
 sg13g2_decap_4 FILLER_2_1506 ();
 sg13g2_fill_1 FILLER_2_1540 ();
 sg13g2_fill_1 FILLER_2_1567 ();
 sg13g2_decap_4 FILLER_2_1572 ();
 sg13g2_fill_2 FILLER_2_1576 ();
 sg13g2_fill_1 FILLER_2_1582 ();
 sg13g2_fill_2 FILLER_2_1587 ();
 sg13g2_fill_1 FILLER_2_1619 ();
 sg13g2_decap_8 FILLER_2_1624 ();
 sg13g2_decap_4 FILLER_2_1631 ();
 sg13g2_fill_2 FILLER_2_1651 ();
 sg13g2_fill_2 FILLER_2_1657 ();
 sg13g2_fill_1 FILLER_2_1659 ();
 sg13g2_fill_1 FILLER_2_1664 ();
 sg13g2_fill_2 FILLER_2_1669 ();
 sg13g2_decap_8 FILLER_2_1675 ();
 sg13g2_decap_4 FILLER_2_1682 ();
 sg13g2_fill_2 FILLER_2_1690 ();
 sg13g2_fill_2 FILLER_2_1722 ();
 sg13g2_fill_1 FILLER_2_1724 ();
 sg13g2_fill_2 FILLER_2_1751 ();
 sg13g2_fill_1 FILLER_2_1753 ();
 sg13g2_fill_2 FILLER_2_1767 ();
 sg13g2_decap_4 FILLER_2_1795 ();
 sg13g2_fill_1 FILLER_2_1799 ();
 sg13g2_decap_8 FILLER_2_1830 ();
 sg13g2_decap_4 FILLER_2_1837 ();
 sg13g2_fill_1 FILLER_2_1841 ();
 sg13g2_decap_8 FILLER_2_1846 ();
 sg13g2_fill_1 FILLER_2_1853 ();
 sg13g2_fill_2 FILLER_2_1946 ();
 sg13g2_fill_2 FILLER_2_1985 ();
 sg13g2_fill_1 FILLER_2_2039 ();
 sg13g2_fill_1 FILLER_2_2176 ();
 sg13g2_fill_1 FILLER_2_2203 ();
 sg13g2_fill_1 FILLER_2_2230 ();
 sg13g2_fill_2 FILLER_2_2241 ();
 sg13g2_fill_1 FILLER_2_2264 ();
 sg13g2_decap_8 FILLER_2_2291 ();
 sg13g2_decap_8 FILLER_2_2298 ();
 sg13g2_decap_8 FILLER_2_2305 ();
 sg13g2_decap_8 FILLER_2_2312 ();
 sg13g2_decap_8 FILLER_2_2319 ();
 sg13g2_decap_8 FILLER_2_2326 ();
 sg13g2_decap_8 FILLER_2_2333 ();
 sg13g2_decap_8 FILLER_2_2340 ();
 sg13g2_decap_8 FILLER_2_2347 ();
 sg13g2_decap_8 FILLER_2_2354 ();
 sg13g2_decap_8 FILLER_2_2361 ();
 sg13g2_fill_2 FILLER_2_2368 ();
 sg13g2_fill_1 FILLER_2_2373 ();
 sg13g2_fill_1 FILLER_2_2383 ();
 sg13g2_decap_8 FILLER_2_2399 ();
 sg13g2_decap_8 FILLER_2_2406 ();
 sg13g2_decap_8 FILLER_2_2413 ();
 sg13g2_decap_8 FILLER_2_2420 ();
 sg13g2_decap_8 FILLER_2_2427 ();
 sg13g2_decap_8 FILLER_2_2434 ();
 sg13g2_decap_8 FILLER_2_2441 ();
 sg13g2_decap_8 FILLER_2_2448 ();
 sg13g2_decap_8 FILLER_2_2455 ();
 sg13g2_decap_8 FILLER_2_2462 ();
 sg13g2_decap_8 FILLER_2_2469 ();
 sg13g2_decap_8 FILLER_2_2476 ();
 sg13g2_decap_8 FILLER_2_2483 ();
 sg13g2_decap_8 FILLER_2_2490 ();
 sg13g2_decap_8 FILLER_2_2497 ();
 sg13g2_decap_8 FILLER_2_2504 ();
 sg13g2_decap_8 FILLER_2_2511 ();
 sg13g2_decap_8 FILLER_2_2518 ();
 sg13g2_decap_8 FILLER_2_2525 ();
 sg13g2_decap_8 FILLER_2_2532 ();
 sg13g2_decap_8 FILLER_2_2539 ();
 sg13g2_decap_8 FILLER_2_2546 ();
 sg13g2_decap_8 FILLER_2_2553 ();
 sg13g2_decap_8 FILLER_2_2560 ();
 sg13g2_decap_8 FILLER_2_2567 ();
 sg13g2_decap_8 FILLER_2_2574 ();
 sg13g2_decap_8 FILLER_2_2581 ();
 sg13g2_decap_8 FILLER_2_2588 ();
 sg13g2_decap_8 FILLER_2_2595 ();
 sg13g2_decap_8 FILLER_2_2602 ();
 sg13g2_decap_8 FILLER_2_2609 ();
 sg13g2_decap_8 FILLER_2_2616 ();
 sg13g2_decap_8 FILLER_2_2623 ();
 sg13g2_decap_8 FILLER_2_2630 ();
 sg13g2_decap_8 FILLER_2_2637 ();
 sg13g2_decap_8 FILLER_2_2644 ();
 sg13g2_decap_8 FILLER_2_2651 ();
 sg13g2_decap_8 FILLER_2_2658 ();
 sg13g2_decap_4 FILLER_2_2665 ();
 sg13g2_fill_1 FILLER_2_2669 ();
 sg13g2_decap_8 FILLER_3_0 ();
 sg13g2_decap_8 FILLER_3_7 ();
 sg13g2_decap_8 FILLER_3_14 ();
 sg13g2_decap_8 FILLER_3_21 ();
 sg13g2_decap_8 FILLER_3_28 ();
 sg13g2_decap_8 FILLER_3_35 ();
 sg13g2_decap_8 FILLER_3_42 ();
 sg13g2_decap_8 FILLER_3_49 ();
 sg13g2_decap_8 FILLER_3_56 ();
 sg13g2_decap_8 FILLER_3_63 ();
 sg13g2_decap_4 FILLER_3_70 ();
 sg13g2_fill_2 FILLER_3_92 ();
 sg13g2_fill_1 FILLER_3_138 ();
 sg13g2_fill_1 FILLER_3_164 ();
 sg13g2_decap_4 FILLER_3_195 ();
 sg13g2_fill_1 FILLER_3_199 ();
 sg13g2_fill_1 FILLER_3_210 ();
 sg13g2_fill_2 FILLER_3_233 ();
 sg13g2_fill_1 FILLER_3_241 ();
 sg13g2_fill_1 FILLER_3_248 ();
 sg13g2_fill_2 FILLER_3_255 ();
 sg13g2_fill_1 FILLER_3_284 ();
 sg13g2_fill_1 FILLER_3_296 ();
 sg13g2_fill_1 FILLER_3_322 ();
 sg13g2_fill_1 FILLER_3_329 ();
 sg13g2_fill_1 FILLER_3_334 ();
 sg13g2_fill_1 FILLER_3_344 ();
 sg13g2_decap_8 FILLER_3_420 ();
 sg13g2_decap_8 FILLER_3_427 ();
 sg13g2_fill_2 FILLER_3_434 ();
 sg13g2_fill_1 FILLER_3_436 ();
 sg13g2_decap_4 FILLER_3_473 ();
 sg13g2_fill_1 FILLER_3_477 ();
 sg13g2_fill_1 FILLER_3_482 ();
 sg13g2_fill_1 FILLER_3_488 ();
 sg13g2_fill_1 FILLER_3_494 ();
 sg13g2_fill_1 FILLER_3_500 ();
 sg13g2_fill_2 FILLER_3_505 ();
 sg13g2_fill_2 FILLER_3_517 ();
 sg13g2_fill_2 FILLER_3_540 ();
 sg13g2_fill_1 FILLER_3_568 ();
 sg13g2_decap_4 FILLER_3_575 ();
 sg13g2_fill_2 FILLER_3_579 ();
 sg13g2_fill_1 FILLER_3_633 ();
 sg13g2_fill_1 FILLER_3_639 ();
 sg13g2_fill_2 FILLER_3_696 ();
 sg13g2_fill_1 FILLER_3_706 ();
 sg13g2_fill_2 FILLER_3_765 ();
 sg13g2_fill_1 FILLER_3_767 ();
 sg13g2_fill_1 FILLER_3_773 ();
 sg13g2_fill_1 FILLER_3_779 ();
 sg13g2_fill_2 FILLER_3_855 ();
 sg13g2_decap_8 FILLER_3_919 ();
 sg13g2_decap_8 FILLER_3_926 ();
 sg13g2_decap_8 FILLER_3_933 ();
 sg13g2_decap_8 FILLER_3_940 ();
 sg13g2_decap_8 FILLER_3_961 ();
 sg13g2_decap_8 FILLER_3_968 ();
 sg13g2_decap_8 FILLER_3_975 ();
 sg13g2_fill_2 FILLER_3_990 ();
 sg13g2_fill_1 FILLER_3_992 ();
 sg13g2_fill_2 FILLER_3_1045 ();
 sg13g2_decap_8 FILLER_3_1077 ();
 sg13g2_decap_8 FILLER_3_1084 ();
 sg13g2_fill_2 FILLER_3_1099 ();
 sg13g2_fill_2 FILLER_3_1106 ();
 sg13g2_fill_2 FILLER_3_1138 ();
 sg13g2_fill_2 FILLER_3_1145 ();
 sg13g2_fill_1 FILLER_3_1151 ();
 sg13g2_fill_1 FILLER_3_1182 ();
 sg13g2_fill_1 FILLER_3_1188 ();
 sg13g2_fill_1 FILLER_3_1193 ();
 sg13g2_fill_2 FILLER_3_1268 ();
 sg13g2_fill_1 FILLER_3_1270 ();
 sg13g2_fill_1 FILLER_3_1300 ();
 sg13g2_fill_1 FILLER_3_1305 ();
 sg13g2_fill_1 FILLER_3_1311 ();
 sg13g2_fill_2 FILLER_3_1316 ();
 sg13g2_fill_1 FILLER_3_1318 ();
 sg13g2_fill_1 FILLER_3_1323 ();
 sg13g2_fill_2 FILLER_3_1350 ();
 sg13g2_fill_2 FILLER_3_1356 ();
 sg13g2_fill_1 FILLER_3_1358 ();
 sg13g2_fill_1 FILLER_3_1364 ();
 sg13g2_fill_2 FILLER_3_1395 ();
 sg13g2_fill_1 FILLER_3_1397 ();
 sg13g2_fill_1 FILLER_3_1423 ();
 sg13g2_fill_2 FILLER_3_1428 ();
 sg13g2_fill_1 FILLER_3_1430 ();
 sg13g2_decap_4 FILLER_3_1441 ();
 sg13g2_fill_1 FILLER_3_1445 ();
 sg13g2_fill_2 FILLER_3_1454 ();
 sg13g2_fill_1 FILLER_3_1456 ();
 sg13g2_fill_1 FILLER_3_1461 ();
 sg13g2_fill_1 FILLER_3_1466 ();
 sg13g2_fill_2 FILLER_3_1477 ();
 sg13g2_decap_8 FILLER_3_1505 ();
 sg13g2_decap_4 FILLER_3_1512 ();
 sg13g2_fill_1 FILLER_3_1577 ();
 sg13g2_fill_2 FILLER_3_1607 ();
 sg13g2_fill_1 FILLER_3_1635 ();
 sg13g2_fill_1 FILLER_3_1688 ();
 sg13g2_fill_1 FILLER_3_1719 ();
 sg13g2_fill_1 FILLER_3_1724 ();
 sg13g2_fill_2 FILLER_3_1797 ();
 sg13g2_fill_1 FILLER_3_1799 ();
 sg13g2_fill_2 FILLER_3_1810 ();
 sg13g2_decap_8 FILLER_3_1826 ();
 sg13g2_decap_8 FILLER_3_1889 ();
 sg13g2_decap_8 FILLER_3_1920 ();
 sg13g2_fill_2 FILLER_3_1927 ();
 sg13g2_fill_2 FILLER_3_1955 ();
 sg13g2_fill_1 FILLER_3_1957 ();
 sg13g2_fill_1 FILLER_3_1994 ();
 sg13g2_decap_8 FILLER_3_2024 ();
 sg13g2_fill_2 FILLER_3_2031 ();
 sg13g2_fill_1 FILLER_3_2033 ();
 sg13g2_fill_2 FILLER_3_2084 ();
 sg13g2_fill_1 FILLER_3_2166 ();
 sg13g2_fill_2 FILLER_3_2180 ();
 sg13g2_fill_1 FILLER_3_2182 ();
 sg13g2_decap_8 FILLER_3_2217 ();
 sg13g2_decap_8 FILLER_3_2224 ();
 sg13g2_decap_4 FILLER_3_2231 ();
 sg13g2_fill_2 FILLER_3_2235 ();
 sg13g2_decap_4 FILLER_3_2241 ();
 sg13g2_fill_1 FILLER_3_2245 ();
 sg13g2_decap_4 FILLER_3_2256 ();
 sg13g2_fill_1 FILLER_3_2260 ();
 sg13g2_fill_2 FILLER_3_2291 ();
 sg13g2_decap_8 FILLER_3_2297 ();
 sg13g2_decap_8 FILLER_3_2304 ();
 sg13g2_decap_8 FILLER_3_2311 ();
 sg13g2_decap_8 FILLER_3_2318 ();
 sg13g2_decap_8 FILLER_3_2325 ();
 sg13g2_decap_8 FILLER_3_2332 ();
 sg13g2_decap_8 FILLER_3_2339 ();
 sg13g2_decap_8 FILLER_3_2346 ();
 sg13g2_decap_8 FILLER_3_2353 ();
 sg13g2_decap_4 FILLER_3_2360 ();
 sg13g2_fill_1 FILLER_3_2370 ();
 sg13g2_fill_1 FILLER_3_2383 ();
 sg13g2_decap_8 FILLER_3_2418 ();
 sg13g2_decap_8 FILLER_3_2425 ();
 sg13g2_decap_8 FILLER_3_2432 ();
 sg13g2_decap_8 FILLER_3_2439 ();
 sg13g2_decap_8 FILLER_3_2446 ();
 sg13g2_decap_8 FILLER_3_2453 ();
 sg13g2_decap_8 FILLER_3_2460 ();
 sg13g2_decap_8 FILLER_3_2467 ();
 sg13g2_decap_8 FILLER_3_2474 ();
 sg13g2_decap_8 FILLER_3_2481 ();
 sg13g2_decap_8 FILLER_3_2488 ();
 sg13g2_decap_8 FILLER_3_2495 ();
 sg13g2_decap_8 FILLER_3_2502 ();
 sg13g2_decap_8 FILLER_3_2509 ();
 sg13g2_decap_8 FILLER_3_2516 ();
 sg13g2_decap_8 FILLER_3_2523 ();
 sg13g2_decap_8 FILLER_3_2530 ();
 sg13g2_decap_8 FILLER_3_2537 ();
 sg13g2_decap_8 FILLER_3_2544 ();
 sg13g2_decap_8 FILLER_3_2551 ();
 sg13g2_decap_8 FILLER_3_2558 ();
 sg13g2_decap_8 FILLER_3_2565 ();
 sg13g2_decap_8 FILLER_3_2572 ();
 sg13g2_decap_8 FILLER_3_2579 ();
 sg13g2_decap_8 FILLER_3_2586 ();
 sg13g2_decap_8 FILLER_3_2593 ();
 sg13g2_decap_8 FILLER_3_2600 ();
 sg13g2_decap_8 FILLER_3_2607 ();
 sg13g2_decap_8 FILLER_3_2614 ();
 sg13g2_decap_8 FILLER_3_2621 ();
 sg13g2_decap_8 FILLER_3_2628 ();
 sg13g2_decap_8 FILLER_3_2635 ();
 sg13g2_decap_8 FILLER_3_2642 ();
 sg13g2_decap_8 FILLER_3_2649 ();
 sg13g2_decap_8 FILLER_3_2656 ();
 sg13g2_decap_8 FILLER_3_2663 ();
 sg13g2_decap_8 FILLER_4_0 ();
 sg13g2_decap_8 FILLER_4_7 ();
 sg13g2_decap_8 FILLER_4_14 ();
 sg13g2_decap_8 FILLER_4_21 ();
 sg13g2_decap_8 FILLER_4_28 ();
 sg13g2_decap_8 FILLER_4_35 ();
 sg13g2_decap_8 FILLER_4_42 ();
 sg13g2_decap_8 FILLER_4_49 ();
 sg13g2_decap_8 FILLER_4_56 ();
 sg13g2_decap_4 FILLER_4_63 ();
 sg13g2_fill_2 FILLER_4_67 ();
 sg13g2_fill_2 FILLER_4_73 ();
 sg13g2_fill_2 FILLER_4_155 ();
 sg13g2_fill_2 FILLER_4_193 ();
 sg13g2_fill_2 FILLER_4_203 ();
 sg13g2_fill_1 FILLER_4_239 ();
 sg13g2_fill_2 FILLER_4_265 ();
 sg13g2_decap_8 FILLER_4_278 ();
 sg13g2_fill_2 FILLER_4_285 ();
 sg13g2_fill_1 FILLER_4_287 ();
 sg13g2_fill_1 FILLER_4_309 ();
 sg13g2_fill_1 FILLER_4_335 ();
 sg13g2_fill_1 FILLER_4_387 ();
 sg13g2_fill_1 FILLER_4_402 ();
 sg13g2_decap_8 FILLER_4_427 ();
 sg13g2_fill_1 FILLER_4_434 ();
 sg13g2_fill_2 FILLER_4_461 ();
 sg13g2_fill_2 FILLER_4_471 ();
 sg13g2_fill_1 FILLER_4_473 ();
 sg13g2_fill_1 FILLER_4_483 ();
 sg13g2_decap_4 FILLER_4_545 ();
 sg13g2_fill_1 FILLER_4_549 ();
 sg13g2_fill_2 FILLER_4_580 ();
 sg13g2_fill_2 FILLER_4_597 ();
 sg13g2_fill_2 FILLER_4_620 ();
 sg13g2_fill_1 FILLER_4_632 ();
 sg13g2_fill_2 FILLER_4_655 ();
 sg13g2_fill_2 FILLER_4_664 ();
 sg13g2_fill_2 FILLER_4_677 ();
 sg13g2_fill_1 FILLER_4_683 ();
 sg13g2_fill_2 FILLER_4_690 ();
 sg13g2_fill_2 FILLER_4_720 ();
 sg13g2_fill_2 FILLER_4_741 ();
 sg13g2_fill_2 FILLER_4_753 ();
 sg13g2_decap_4 FILLER_4_790 ();
 sg13g2_fill_1 FILLER_4_794 ();
 sg13g2_decap_8 FILLER_4_799 ();
 sg13g2_decap_8 FILLER_4_806 ();
 sg13g2_fill_1 FILLER_4_813 ();
 sg13g2_fill_1 FILLER_4_818 ();
 sg13g2_decap_8 FILLER_4_823 ();
 sg13g2_fill_2 FILLER_4_851 ();
 sg13g2_fill_2 FILLER_4_857 ();
 sg13g2_fill_2 FILLER_4_863 ();
 sg13g2_fill_1 FILLER_4_865 ();
 sg13g2_fill_2 FILLER_4_923 ();
 sg13g2_decap_4 FILLER_4_982 ();
 sg13g2_fill_2 FILLER_4_1016 ();
 sg13g2_fill_2 FILLER_4_1039 ();
 sg13g2_fill_1 FILLER_4_1045 ();
 sg13g2_decap_4 FILLER_4_1050 ();
 sg13g2_fill_2 FILLER_4_1058 ();
 sg13g2_fill_2 FILLER_4_1064 ();
 sg13g2_fill_1 FILLER_4_1104 ();
 sg13g2_decap_8 FILLER_4_1131 ();
 sg13g2_decap_8 FILLER_4_1138 ();
 sg13g2_decap_4 FILLER_4_1145 ();
 sg13g2_fill_1 FILLER_4_1149 ();
 sg13g2_decap_8 FILLER_4_1154 ();
 sg13g2_fill_2 FILLER_4_1170 ();
 sg13g2_fill_1 FILLER_4_1172 ();
 sg13g2_decap_8 FILLER_4_1177 ();
 sg13g2_decap_8 FILLER_4_1184 ();
 sg13g2_decap_4 FILLER_4_1191 ();
 sg13g2_fill_2 FILLER_4_1195 ();
 sg13g2_fill_1 FILLER_4_1202 ();
 sg13g2_decap_4 FILLER_4_1211 ();
 sg13g2_fill_2 FILLER_4_1220 ();
 sg13g2_fill_1 FILLER_4_1222 ();
 sg13g2_decap_4 FILLER_4_1244 ();
 sg13g2_decap_4 FILLER_4_1253 ();
 sg13g2_fill_1 FILLER_4_1257 ();
 sg13g2_fill_1 FILLER_4_1288 ();
 sg13g2_fill_2 FILLER_4_1320 ();
 sg13g2_fill_2 FILLER_4_1327 ();
 sg13g2_fill_1 FILLER_4_1329 ();
 sg13g2_fill_2 FILLER_4_1351 ();
 sg13g2_decap_4 FILLER_4_1379 ();
 sg13g2_fill_1 FILLER_4_1393 ();
 sg13g2_fill_2 FILLER_4_1404 ();
 sg13g2_fill_1 FILLER_4_1406 ();
 sg13g2_decap_8 FILLER_4_1411 ();
 sg13g2_decap_8 FILLER_4_1418 ();
 sg13g2_decap_8 FILLER_4_1425 ();
 sg13g2_fill_2 FILLER_4_1432 ();
 sg13g2_fill_1 FILLER_4_1434 ();
 sg13g2_fill_1 FILLER_4_1465 ();
 sg13g2_decap_8 FILLER_4_1502 ();
 sg13g2_decap_8 FILLER_4_1509 ();
 sg13g2_decap_8 FILLER_4_1516 ();
 sg13g2_decap_4 FILLER_4_1523 ();
 sg13g2_decap_8 FILLER_4_1548 ();
 sg13g2_fill_1 FILLER_4_1555 ();
 sg13g2_fill_1 FILLER_4_1575 ();
 sg13g2_decap_4 FILLER_4_1586 ();
 sg13g2_fill_2 FILLER_4_1631 ();
 sg13g2_fill_1 FILLER_4_1633 ();
 sg13g2_fill_2 FILLER_4_1662 ();
 sg13g2_decap_4 FILLER_4_1668 ();
 sg13g2_fill_2 FILLER_4_1676 ();
 sg13g2_fill_1 FILLER_4_1678 ();
 sg13g2_decap_4 FILLER_4_1695 ();
 sg13g2_fill_1 FILLER_4_1699 ();
 sg13g2_decap_8 FILLER_4_1704 ();
 sg13g2_fill_2 FILLER_4_1711 ();
 sg13g2_decap_8 FILLER_4_1718 ();
 sg13g2_fill_1 FILLER_4_1725 ();
 sg13g2_decap_8 FILLER_4_1761 ();
 sg13g2_decap_4 FILLER_4_1768 ();
 sg13g2_fill_1 FILLER_4_1772 ();
 sg13g2_decap_4 FILLER_4_1797 ();
 sg13g2_fill_2 FILLER_4_1811 ();
 sg13g2_fill_1 FILLER_4_1813 ();
 sg13g2_fill_1 FILLER_4_1844 ();
 sg13g2_decap_4 FILLER_4_1875 ();
 sg13g2_decap_8 FILLER_4_1900 ();
 sg13g2_fill_2 FILLER_4_1907 ();
 sg13g2_fill_1 FILLER_4_1923 ();
 sg13g2_fill_1 FILLER_4_1950 ();
 sg13g2_fill_1 FILLER_4_1961 ();
 sg13g2_fill_1 FILLER_4_1966 ();
 sg13g2_decap_4 FILLER_4_1977 ();
 sg13g2_fill_2 FILLER_4_1981 ();
 sg13g2_decap_8 FILLER_4_1991 ();
 sg13g2_decap_4 FILLER_4_1998 ();
 sg13g2_fill_1 FILLER_4_2002 ();
 sg13g2_decap_8 FILLER_4_2013 ();
 sg13g2_fill_2 FILLER_4_2028 ();
 sg13g2_fill_1 FILLER_4_2060 ();
 sg13g2_decap_4 FILLER_4_2127 ();
 sg13g2_fill_1 FILLER_4_2131 ();
 sg13g2_fill_2 FILLER_4_2142 ();
 sg13g2_fill_1 FILLER_4_2144 ();
 sg13g2_fill_2 FILLER_4_2166 ();
 sg13g2_fill_1 FILLER_4_2168 ();
 sg13g2_decap_4 FILLER_4_2183 ();
 sg13g2_fill_2 FILLER_4_2187 ();
 sg13g2_decap_4 FILLER_4_2193 ();
 sg13g2_decap_8 FILLER_4_2207 ();
 sg13g2_decap_8 FILLER_4_2214 ();
 sg13g2_fill_1 FILLER_4_2251 ();
 sg13g2_fill_2 FILLER_4_2275 ();
 sg13g2_decap_8 FILLER_4_2303 ();
 sg13g2_decap_8 FILLER_4_2310 ();
 sg13g2_decap_8 FILLER_4_2317 ();
 sg13g2_decap_8 FILLER_4_2324 ();
 sg13g2_decap_8 FILLER_4_2331 ();
 sg13g2_decap_8 FILLER_4_2338 ();
 sg13g2_decap_8 FILLER_4_2345 ();
 sg13g2_fill_2 FILLER_4_2352 ();
 sg13g2_fill_1 FILLER_4_2363 ();
 sg13g2_fill_1 FILLER_4_2370 ();
 sg13g2_fill_2 FILLER_4_2386 ();
 sg13g2_fill_2 FILLER_4_2424 ();
 sg13g2_decap_8 FILLER_4_2438 ();
 sg13g2_decap_8 FILLER_4_2445 ();
 sg13g2_decap_8 FILLER_4_2452 ();
 sg13g2_decap_8 FILLER_4_2459 ();
 sg13g2_decap_8 FILLER_4_2466 ();
 sg13g2_decap_8 FILLER_4_2473 ();
 sg13g2_decap_8 FILLER_4_2480 ();
 sg13g2_decap_8 FILLER_4_2487 ();
 sg13g2_decap_8 FILLER_4_2494 ();
 sg13g2_decap_8 FILLER_4_2501 ();
 sg13g2_decap_8 FILLER_4_2508 ();
 sg13g2_decap_8 FILLER_4_2515 ();
 sg13g2_decap_8 FILLER_4_2522 ();
 sg13g2_decap_8 FILLER_4_2529 ();
 sg13g2_decap_8 FILLER_4_2536 ();
 sg13g2_decap_8 FILLER_4_2543 ();
 sg13g2_decap_8 FILLER_4_2550 ();
 sg13g2_decap_8 FILLER_4_2557 ();
 sg13g2_decap_8 FILLER_4_2564 ();
 sg13g2_decap_8 FILLER_4_2571 ();
 sg13g2_decap_8 FILLER_4_2578 ();
 sg13g2_decap_8 FILLER_4_2585 ();
 sg13g2_decap_8 FILLER_4_2592 ();
 sg13g2_decap_8 FILLER_4_2599 ();
 sg13g2_decap_8 FILLER_4_2606 ();
 sg13g2_decap_8 FILLER_4_2613 ();
 sg13g2_decap_8 FILLER_4_2620 ();
 sg13g2_decap_8 FILLER_4_2627 ();
 sg13g2_decap_8 FILLER_4_2634 ();
 sg13g2_decap_8 FILLER_4_2641 ();
 sg13g2_decap_8 FILLER_4_2648 ();
 sg13g2_decap_8 FILLER_4_2655 ();
 sg13g2_decap_8 FILLER_4_2662 ();
 sg13g2_fill_1 FILLER_4_2669 ();
 sg13g2_decap_8 FILLER_5_0 ();
 sg13g2_decap_8 FILLER_5_7 ();
 sg13g2_decap_8 FILLER_5_14 ();
 sg13g2_decap_8 FILLER_5_21 ();
 sg13g2_decap_8 FILLER_5_28 ();
 sg13g2_decap_8 FILLER_5_35 ();
 sg13g2_decap_8 FILLER_5_42 ();
 sg13g2_decap_8 FILLER_5_49 ();
 sg13g2_decap_8 FILLER_5_56 ();
 sg13g2_decap_8 FILLER_5_63 ();
 sg13g2_decap_8 FILLER_5_70 ();
 sg13g2_fill_1 FILLER_5_77 ();
 sg13g2_fill_2 FILLER_5_96 ();
 sg13g2_fill_1 FILLER_5_98 ();
 sg13g2_decap_8 FILLER_5_103 ();
 sg13g2_fill_1 FILLER_5_110 ();
 sg13g2_decap_8 FILLER_5_133 ();
 sg13g2_fill_2 FILLER_5_140 ();
 sg13g2_fill_1 FILLER_5_142 ();
 sg13g2_fill_2 FILLER_5_162 ();
 sg13g2_fill_1 FILLER_5_164 ();
 sg13g2_fill_2 FILLER_5_169 ();
 sg13g2_decap_8 FILLER_5_207 ();
 sg13g2_decap_4 FILLER_5_214 ();
 sg13g2_fill_2 FILLER_5_218 ();
 sg13g2_decap_8 FILLER_5_224 ();
 sg13g2_decap_8 FILLER_5_231 ();
 sg13g2_decap_4 FILLER_5_238 ();
 sg13g2_fill_2 FILLER_5_242 ();
 sg13g2_fill_2 FILLER_5_250 ();
 sg13g2_fill_2 FILLER_5_260 ();
 sg13g2_fill_2 FILLER_5_268 ();
 sg13g2_decap_4 FILLER_5_285 ();
 sg13g2_fill_1 FILLER_5_289 ();
 sg13g2_fill_1 FILLER_5_331 ();
 sg13g2_fill_1 FILLER_5_339 ();
 sg13g2_fill_1 FILLER_5_358 ();
 sg13g2_fill_1 FILLER_5_369 ();
 sg13g2_fill_1 FILLER_5_387 ();
 sg13g2_fill_1 FILLER_5_391 ();
 sg13g2_fill_1 FILLER_5_398 ();
 sg13g2_fill_1 FILLER_5_408 ();
 sg13g2_decap_4 FILLER_5_433 ();
 sg13g2_decap_8 FILLER_5_480 ();
 sg13g2_decap_8 FILLER_5_487 ();
 sg13g2_fill_1 FILLER_5_494 ();
 sg13g2_fill_2 FILLER_5_519 ();
 sg13g2_fill_1 FILLER_5_526 ();
 sg13g2_fill_1 FILLER_5_530 ();
 sg13g2_fill_2 FILLER_5_541 ();
 sg13g2_fill_1 FILLER_5_543 ();
 sg13g2_fill_1 FILLER_5_572 ();
 sg13g2_fill_1 FILLER_5_578 ();
 sg13g2_fill_1 FILLER_5_589 ();
 sg13g2_fill_1 FILLER_5_596 ();
 sg13g2_decap_8 FILLER_5_616 ();
 sg13g2_fill_2 FILLER_5_623 ();
 sg13g2_decap_4 FILLER_5_630 ();
 sg13g2_decap_8 FILLER_5_638 ();
 sg13g2_decap_4 FILLER_5_645 ();
 sg13g2_fill_2 FILLER_5_649 ();
 sg13g2_fill_2 FILLER_5_707 ();
 sg13g2_fill_2 FILLER_5_729 ();
 sg13g2_fill_2 FILLER_5_757 ();
 sg13g2_decap_4 FILLER_5_764 ();
 sg13g2_decap_8 FILLER_5_802 ();
 sg13g2_decap_8 FILLER_5_809 ();
 sg13g2_decap_8 FILLER_5_816 ();
 sg13g2_decap_8 FILLER_5_823 ();
 sg13g2_fill_2 FILLER_5_830 ();
 sg13g2_decap_4 FILLER_5_850 ();
 sg13g2_fill_2 FILLER_5_854 ();
 sg13g2_fill_2 FILLER_5_866 ();
 sg13g2_fill_1 FILLER_5_868 ();
 sg13g2_fill_1 FILLER_5_899 ();
 sg13g2_fill_1 FILLER_5_921 ();
 sg13g2_fill_1 FILLER_5_948 ();
 sg13g2_fill_2 FILLER_5_975 ();
 sg13g2_fill_1 FILLER_5_1048 ();
 sg13g2_decap_8 FILLER_5_1062 ();
 sg13g2_decap_8 FILLER_5_1069 ();
 sg13g2_fill_2 FILLER_5_1076 ();
 sg13g2_fill_1 FILLER_5_1078 ();
 sg13g2_fill_2 FILLER_5_1114 ();
 sg13g2_fill_1 FILLER_5_1116 ();
 sg13g2_decap_8 FILLER_5_1134 ();
 sg13g2_decap_8 FILLER_5_1180 ();
 sg13g2_decap_4 FILLER_5_1187 ();
 sg13g2_fill_1 FILLER_5_1191 ();
 sg13g2_decap_8 FILLER_5_1196 ();
 sg13g2_decap_8 FILLER_5_1203 ();
 sg13g2_decap_8 FILLER_5_1210 ();
 sg13g2_fill_1 FILLER_5_1248 ();
 sg13g2_fill_2 FILLER_5_1284 ();
 sg13g2_fill_2 FILLER_5_1342 ();
 sg13g2_decap_8 FILLER_5_1348 ();
 sg13g2_decap_4 FILLER_5_1355 ();
 sg13g2_fill_2 FILLER_5_1368 ();
 sg13g2_fill_1 FILLER_5_1370 ();
 sg13g2_fill_2 FILLER_5_1397 ();
 sg13g2_fill_1 FILLER_5_1399 ();
 sg13g2_fill_1 FILLER_5_1426 ();
 sg13g2_decap_4 FILLER_5_1477 ();
 sg13g2_decap_8 FILLER_5_1489 ();
 sg13g2_fill_2 FILLER_5_1496 ();
 sg13g2_fill_2 FILLER_5_1554 ();
 sg13g2_fill_2 FILLER_5_1585 ();
 sg13g2_decap_8 FILLER_5_1592 ();
 sg13g2_fill_1 FILLER_5_1637 ();
 sg13g2_decap_4 FILLER_5_1709 ();
 sg13g2_fill_1 FILLER_5_1713 ();
 sg13g2_decap_8 FILLER_5_1719 ();
 sg13g2_decap_8 FILLER_5_1726 ();
 sg13g2_fill_2 FILLER_5_1733 ();
 sg13g2_fill_1 FILLER_5_1735 ();
 sg13g2_decap_8 FILLER_5_1744 ();
 sg13g2_decap_8 FILLER_5_1751 ();
 sg13g2_decap_8 FILLER_5_1758 ();
 sg13g2_decap_8 FILLER_5_1765 ();
 sg13g2_decap_4 FILLER_5_1772 ();
 sg13g2_decap_4 FILLER_5_1780 ();
 sg13g2_fill_2 FILLER_5_1784 ();
 sg13g2_decap_8 FILLER_5_1794 ();
 sg13g2_decap_4 FILLER_5_1801 ();
 sg13g2_decap_8 FILLER_5_1836 ();
 sg13g2_decap_8 FILLER_5_1843 ();
 sg13g2_decap_4 FILLER_5_1850 ();
 sg13g2_fill_2 FILLER_5_1864 ();
 sg13g2_decap_4 FILLER_5_1876 ();
 sg13g2_decap_4 FILLER_5_1924 ();
 sg13g2_decap_4 FILLER_5_1942 ();
 sg13g2_fill_1 FILLER_5_1946 ();
 sg13g2_fill_2 FILLER_5_1968 ();
 sg13g2_fill_1 FILLER_5_1970 ();
 sg13g2_fill_2 FILLER_5_2005 ();
 sg13g2_fill_1 FILLER_5_2007 ();
 sg13g2_decap_4 FILLER_5_2026 ();
 sg13g2_decap_4 FILLER_5_2034 ();
 sg13g2_fill_2 FILLER_5_2038 ();
 sg13g2_fill_2 FILLER_5_2048 ();
 sg13g2_fill_1 FILLER_5_2050 ();
 sg13g2_decap_4 FILLER_5_2120 ();
 sg13g2_fill_2 FILLER_5_2134 ();
 sg13g2_decap_8 FILLER_5_2157 ();
 sg13g2_decap_8 FILLER_5_2164 ();
 sg13g2_decap_8 FILLER_5_2192 ();
 sg13g2_decap_8 FILLER_5_2199 ();
 sg13g2_decap_8 FILLER_5_2206 ();
 sg13g2_fill_1 FILLER_5_2213 ();
 sg13g2_fill_2 FILLER_5_2218 ();
 sg13g2_decap_4 FILLER_5_2246 ();
 sg13g2_decap_8 FILLER_5_2297 ();
 sg13g2_decap_4 FILLER_5_2304 ();
 sg13g2_decap_8 FILLER_5_2323 ();
 sg13g2_decap_8 FILLER_5_2330 ();
 sg13g2_decap_8 FILLER_5_2337 ();
 sg13g2_fill_2 FILLER_5_2344 ();
 sg13g2_fill_2 FILLER_5_2358 ();
 sg13g2_fill_2 FILLER_5_2432 ();
 sg13g2_fill_2 FILLER_5_2444 ();
 sg13g2_fill_2 FILLER_5_2453 ();
 sg13g2_decap_8 FILLER_5_2465 ();
 sg13g2_decap_8 FILLER_5_2472 ();
 sg13g2_decap_8 FILLER_5_2479 ();
 sg13g2_decap_8 FILLER_5_2486 ();
 sg13g2_decap_8 FILLER_5_2493 ();
 sg13g2_decap_8 FILLER_5_2500 ();
 sg13g2_decap_8 FILLER_5_2507 ();
 sg13g2_decap_8 FILLER_5_2514 ();
 sg13g2_decap_8 FILLER_5_2521 ();
 sg13g2_decap_8 FILLER_5_2528 ();
 sg13g2_decap_8 FILLER_5_2535 ();
 sg13g2_decap_8 FILLER_5_2542 ();
 sg13g2_decap_8 FILLER_5_2549 ();
 sg13g2_decap_8 FILLER_5_2556 ();
 sg13g2_decap_8 FILLER_5_2563 ();
 sg13g2_decap_8 FILLER_5_2570 ();
 sg13g2_decap_8 FILLER_5_2577 ();
 sg13g2_decap_8 FILLER_5_2584 ();
 sg13g2_decap_8 FILLER_5_2591 ();
 sg13g2_decap_8 FILLER_5_2598 ();
 sg13g2_decap_8 FILLER_5_2605 ();
 sg13g2_decap_8 FILLER_5_2612 ();
 sg13g2_decap_8 FILLER_5_2619 ();
 sg13g2_decap_8 FILLER_5_2626 ();
 sg13g2_decap_8 FILLER_5_2633 ();
 sg13g2_decap_8 FILLER_5_2640 ();
 sg13g2_decap_8 FILLER_5_2647 ();
 sg13g2_decap_8 FILLER_5_2654 ();
 sg13g2_decap_8 FILLER_5_2661 ();
 sg13g2_fill_2 FILLER_5_2668 ();
 sg13g2_decap_8 FILLER_6_0 ();
 sg13g2_decap_8 FILLER_6_7 ();
 sg13g2_decap_8 FILLER_6_14 ();
 sg13g2_decap_8 FILLER_6_21 ();
 sg13g2_decap_8 FILLER_6_28 ();
 sg13g2_decap_8 FILLER_6_35 ();
 sg13g2_decap_4 FILLER_6_42 ();
 sg13g2_fill_2 FILLER_6_46 ();
 sg13g2_decap_8 FILLER_6_91 ();
 sg13g2_fill_1 FILLER_6_98 ();
 sg13g2_decap_4 FILLER_6_132 ();
 sg13g2_fill_2 FILLER_6_136 ();
 sg13g2_fill_1 FILLER_6_168 ();
 sg13g2_fill_2 FILLER_6_188 ();
 sg13g2_fill_2 FILLER_6_194 ();
 sg13g2_decap_4 FILLER_6_263 ();
 sg13g2_decap_8 FILLER_6_285 ();
 sg13g2_fill_2 FILLER_6_326 ();
 sg13g2_fill_1 FILLER_6_354 ();
 sg13g2_fill_1 FILLER_6_365 ();
 sg13g2_fill_2 FILLER_6_378 ();
 sg13g2_fill_2 FILLER_6_389 ();
 sg13g2_fill_1 FILLER_6_394 ();
 sg13g2_fill_1 FILLER_6_400 ();
 sg13g2_fill_1 FILLER_6_427 ();
 sg13g2_fill_1 FILLER_6_487 ();
 sg13g2_decap_8 FILLER_6_495 ();
 sg13g2_fill_1 FILLER_6_555 ();
 sg13g2_decap_8 FILLER_6_570 ();
 sg13g2_decap_4 FILLER_6_577 ();
 sg13g2_decap_4 FILLER_6_622 ();
 sg13g2_fill_1 FILLER_6_626 ();
 sg13g2_fill_2 FILLER_6_631 ();
 sg13g2_fill_2 FILLER_6_642 ();
 sg13g2_fill_1 FILLER_6_648 ();
 sg13g2_decap_4 FILLER_6_657 ();
 sg13g2_decap_4 FILLER_6_665 ();
 sg13g2_fill_1 FILLER_6_669 ();
 sg13g2_decap_4 FILLER_6_675 ();
 sg13g2_fill_1 FILLER_6_679 ();
 sg13g2_decap_8 FILLER_6_689 ();
 sg13g2_fill_1 FILLER_6_696 ();
 sg13g2_fill_2 FILLER_6_721 ();
 sg13g2_fill_2 FILLER_6_728 ();
 sg13g2_decap_8 FILLER_6_745 ();
 sg13g2_decap_4 FILLER_6_752 ();
 sg13g2_fill_2 FILLER_6_756 ();
 sg13g2_decap_8 FILLER_6_783 ();
 sg13g2_fill_2 FILLER_6_790 ();
 sg13g2_decap_8 FILLER_6_796 ();
 sg13g2_decap_8 FILLER_6_803 ();
 sg13g2_fill_2 FILLER_6_810 ();
 sg13g2_fill_1 FILLER_6_812 ();
 sg13g2_decap_4 FILLER_6_839 ();
 sg13g2_fill_2 FILLER_6_843 ();
 sg13g2_decap_4 FILLER_6_855 ();
 sg13g2_fill_2 FILLER_6_863 ();
 sg13g2_fill_1 FILLER_6_865 ();
 sg13g2_fill_1 FILLER_6_881 ();
 sg13g2_fill_2 FILLER_6_886 ();
 sg13g2_fill_2 FILLER_6_898 ();
 sg13g2_fill_1 FILLER_6_904 ();
 sg13g2_fill_2 FILLER_6_956 ();
 sg13g2_fill_1 FILLER_6_958 ();
 sg13g2_decap_4 FILLER_6_963 ();
 sg13g2_fill_2 FILLER_6_967 ();
 sg13g2_fill_1 FILLER_6_1000 ();
 sg13g2_fill_1 FILLER_6_1009 ();
 sg13g2_fill_1 FILLER_6_1031 ();
 sg13g2_fill_2 FILLER_6_1037 ();
 sg13g2_fill_2 FILLER_6_1069 ();
 sg13g2_fill_2 FILLER_6_1079 ();
 sg13g2_fill_1 FILLER_6_1081 ();
 sg13g2_fill_1 FILLER_6_1200 ();
 sg13g2_fill_2 FILLER_6_1206 ();
 sg13g2_fill_1 FILLER_6_1252 ();
 sg13g2_fill_2 FILLER_6_1288 ();
 sg13g2_fill_2 FILLER_6_1324 ();
 sg13g2_fill_1 FILLER_6_1362 ();
 sg13g2_fill_2 FILLER_6_1367 ();
 sg13g2_fill_1 FILLER_6_1369 ();
 sg13g2_decap_8 FILLER_6_1401 ();
 sg13g2_decap_8 FILLER_6_1408 ();
 sg13g2_decap_8 FILLER_6_1415 ();
 sg13g2_decap_8 FILLER_6_1422 ();
 sg13g2_decap_4 FILLER_6_1429 ();
 sg13g2_decap_4 FILLER_6_1443 ();
 sg13g2_decap_8 FILLER_6_1451 ();
 sg13g2_fill_1 FILLER_6_1479 ();
 sg13g2_fill_2 FILLER_6_1488 ();
 sg13g2_decap_8 FILLER_6_1494 ();
 sg13g2_fill_2 FILLER_6_1501 ();
 sg13g2_fill_1 FILLER_6_1503 ();
 sg13g2_fill_2 FILLER_6_1538 ();
 sg13g2_fill_1 FILLER_6_1572 ();
 sg13g2_fill_2 FILLER_6_1582 ();
 sg13g2_decap_8 FILLER_6_1591 ();
 sg13g2_decap_8 FILLER_6_1598 ();
 sg13g2_fill_1 FILLER_6_1605 ();
 sg13g2_fill_1 FILLER_6_1625 ();
 sg13g2_decap_4 FILLER_6_1634 ();
 sg13g2_fill_2 FILLER_6_1638 ();
 sg13g2_fill_1 FILLER_6_1644 ();
 sg13g2_fill_1 FILLER_6_1654 ();
 sg13g2_decap_4 FILLER_6_1730 ();
 sg13g2_fill_2 FILLER_6_1734 ();
 sg13g2_fill_1 FILLER_6_1796 ();
 sg13g2_decap_4 FILLER_6_1842 ();
 sg13g2_fill_1 FILLER_6_1876 ();
 sg13g2_decap_8 FILLER_6_1891 ();
 sg13g2_decap_8 FILLER_6_1898 ();
 sg13g2_fill_2 FILLER_6_1909 ();
 sg13g2_decap_4 FILLER_6_1937 ();
 sg13g2_decap_4 FILLER_6_1967 ();
 sg13g2_fill_2 FILLER_6_1992 ();
 sg13g2_fill_2 FILLER_6_1998 ();
 sg13g2_fill_1 FILLER_6_2000 ();
 sg13g2_fill_1 FILLER_6_2022 ();
 sg13g2_fill_1 FILLER_6_2049 ();
 sg13g2_fill_2 FILLER_6_2076 ();
 sg13g2_fill_1 FILLER_6_2082 ();
 sg13g2_fill_2 FILLER_6_2109 ();
 sg13g2_decap_8 FILLER_6_2147 ();
 sg13g2_fill_2 FILLER_6_2154 ();
 sg13g2_fill_1 FILLER_6_2182 ();
 sg13g2_decap_4 FILLER_6_2186 ();
 sg13g2_decap_8 FILLER_6_2273 ();
 sg13g2_decap_4 FILLER_6_2280 ();
 sg13g2_fill_1 FILLER_6_2284 ();
 sg13g2_fill_1 FILLER_6_2289 ();
 sg13g2_fill_2 FILLER_6_2296 ();
 sg13g2_fill_2 FILLER_6_2317 ();
 sg13g2_fill_1 FILLER_6_2359 ();
 sg13g2_fill_1 FILLER_6_2385 ();
 sg13g2_fill_2 FILLER_6_2411 ();
 sg13g2_fill_2 FILLER_6_2448 ();
 sg13g2_decap_8 FILLER_6_2480 ();
 sg13g2_decap_8 FILLER_6_2487 ();
 sg13g2_decap_8 FILLER_6_2494 ();
 sg13g2_decap_8 FILLER_6_2501 ();
 sg13g2_fill_2 FILLER_6_2511 ();
 sg13g2_fill_1 FILLER_6_2513 ();
 sg13g2_decap_8 FILLER_6_2523 ();
 sg13g2_decap_8 FILLER_6_2530 ();
 sg13g2_decap_8 FILLER_6_2537 ();
 sg13g2_decap_8 FILLER_6_2544 ();
 sg13g2_decap_8 FILLER_6_2551 ();
 sg13g2_decap_8 FILLER_6_2558 ();
 sg13g2_decap_8 FILLER_6_2565 ();
 sg13g2_decap_8 FILLER_6_2572 ();
 sg13g2_decap_8 FILLER_6_2579 ();
 sg13g2_decap_8 FILLER_6_2586 ();
 sg13g2_decap_8 FILLER_6_2593 ();
 sg13g2_decap_8 FILLER_6_2600 ();
 sg13g2_decap_8 FILLER_6_2607 ();
 sg13g2_decap_8 FILLER_6_2614 ();
 sg13g2_decap_8 FILLER_6_2621 ();
 sg13g2_decap_8 FILLER_6_2628 ();
 sg13g2_decap_8 FILLER_6_2635 ();
 sg13g2_decap_8 FILLER_6_2642 ();
 sg13g2_decap_8 FILLER_6_2649 ();
 sg13g2_decap_8 FILLER_6_2656 ();
 sg13g2_decap_8 FILLER_6_2663 ();
 sg13g2_decap_8 FILLER_7_0 ();
 sg13g2_decap_8 FILLER_7_7 ();
 sg13g2_decap_8 FILLER_7_14 ();
 sg13g2_decap_8 FILLER_7_21 ();
 sg13g2_decap_8 FILLER_7_28 ();
 sg13g2_decap_8 FILLER_7_35 ();
 sg13g2_decap_8 FILLER_7_42 ();
 sg13g2_decap_8 FILLER_7_49 ();
 sg13g2_fill_1 FILLER_7_56 ();
 sg13g2_decap_4 FILLER_7_101 ();
 sg13g2_fill_2 FILLER_7_105 ();
 sg13g2_fill_2 FILLER_7_111 ();
 sg13g2_fill_2 FILLER_7_139 ();
 sg13g2_decap_8 FILLER_7_154 ();
 sg13g2_fill_1 FILLER_7_161 ();
 sg13g2_decap_4 FILLER_7_166 ();
 sg13g2_fill_1 FILLER_7_175 ();
 sg13g2_fill_1 FILLER_7_180 ();
 sg13g2_decap_8 FILLER_7_191 ();
 sg13g2_decap_8 FILLER_7_198 ();
 sg13g2_fill_2 FILLER_7_205 ();
 sg13g2_fill_1 FILLER_7_207 ();
 sg13g2_fill_1 FILLER_7_218 ();
 sg13g2_fill_1 FILLER_7_223 ();
 sg13g2_fill_2 FILLER_7_229 ();
 sg13g2_fill_1 FILLER_7_231 ();
 sg13g2_fill_2 FILLER_7_268 ();
 sg13g2_fill_1 FILLER_7_314 ();
 sg13g2_fill_1 FILLER_7_340 ();
 sg13g2_fill_2 FILLER_7_355 ();
 sg13g2_fill_2 FILLER_7_389 ();
 sg13g2_fill_2 FILLER_7_467 ();
 sg13g2_fill_2 FILLER_7_514 ();
 sg13g2_decap_8 FILLER_7_551 ();
 sg13g2_decap_8 FILLER_7_558 ();
 sg13g2_fill_1 FILLER_7_565 ();
 sg13g2_decap_8 FILLER_7_571 ();
 sg13g2_decap_8 FILLER_7_578 ();
 sg13g2_fill_2 FILLER_7_698 ();
 sg13g2_decap_4 FILLER_7_726 ();
 sg13g2_decap_4 FILLER_7_753 ();
 sg13g2_fill_2 FILLER_7_757 ();
 sg13g2_fill_1 FILLER_7_764 ();
 sg13g2_fill_1 FILLER_7_769 ();
 sg13g2_fill_2 FILLER_7_784 ();
 sg13g2_fill_1 FILLER_7_786 ();
 sg13g2_fill_1 FILLER_7_813 ();
 sg13g2_decap_4 FILLER_7_844 ();
 sg13g2_fill_1 FILLER_7_848 ();
 sg13g2_decap_8 FILLER_7_883 ();
 sg13g2_decap_8 FILLER_7_890 ();
 sg13g2_decap_8 FILLER_7_897 ();
 sg13g2_decap_8 FILLER_7_904 ();
 sg13g2_decap_8 FILLER_7_911 ();
 sg13g2_decap_8 FILLER_7_918 ();
 sg13g2_decap_4 FILLER_7_925 ();
 sg13g2_fill_1 FILLER_7_929 ();
 sg13g2_decap_8 FILLER_7_934 ();
 sg13g2_decap_8 FILLER_7_962 ();
 sg13g2_decap_8 FILLER_7_969 ();
 sg13g2_decap_4 FILLER_7_976 ();
 sg13g2_fill_1 FILLER_7_988 ();
 sg13g2_fill_1 FILLER_7_993 ();
 sg13g2_fill_1 FILLER_7_1050 ();
 sg13g2_fill_2 FILLER_7_1129 ();
 sg13g2_fill_2 FILLER_7_1140 ();
 sg13g2_fill_2 FILLER_7_1151 ();
 sg13g2_fill_1 FILLER_7_1153 ();
 sg13g2_fill_1 FILLER_7_1163 ();
 sg13g2_fill_2 FILLER_7_1224 ();
 sg13g2_fill_1 FILLER_7_1226 ();
 sg13g2_fill_1 FILLER_7_1253 ();
 sg13g2_fill_2 FILLER_7_1259 ();
 sg13g2_fill_2 FILLER_7_1295 ();
 sg13g2_fill_1 FILLER_7_1297 ();
 sg13g2_fill_2 FILLER_7_1324 ();
 sg13g2_fill_1 FILLER_7_1326 ();
 sg13g2_decap_8 FILLER_7_1348 ();
 sg13g2_decap_4 FILLER_7_1360 ();
 sg13g2_fill_1 FILLER_7_1364 ();
 sg13g2_fill_1 FILLER_7_1373 ();
 sg13g2_fill_1 FILLER_7_1378 ();
 sg13g2_fill_1 FILLER_7_1407 ();
 sg13g2_decap_8 FILLER_7_1434 ();
 sg13g2_decap_8 FILLER_7_1441 ();
 sg13g2_decap_8 FILLER_7_1448 ();
 sg13g2_decap_4 FILLER_7_1455 ();
 sg13g2_fill_1 FILLER_7_1459 ();
 sg13g2_fill_2 FILLER_7_1490 ();
 sg13g2_fill_1 FILLER_7_1492 ();
 sg13g2_decap_8 FILLER_7_1497 ();
 sg13g2_decap_8 FILLER_7_1504 ();
 sg13g2_fill_2 FILLER_7_1511 ();
 sg13g2_fill_2 FILLER_7_1517 ();
 sg13g2_fill_2 FILLER_7_1571 ();
 sg13g2_fill_2 FILLER_7_1582 ();
 sg13g2_fill_1 FILLER_7_1609 ();
 sg13g2_fill_1 FILLER_7_1614 ();
 sg13g2_fill_1 FILLER_7_1622 ();
 sg13g2_fill_1 FILLER_7_1629 ();
 sg13g2_fill_2 FILLER_7_1642 ();
 sg13g2_decap_8 FILLER_7_1650 ();
 sg13g2_fill_1 FILLER_7_1666 ();
 sg13g2_fill_2 FILLER_7_1677 ();
 sg13g2_fill_1 FILLER_7_1689 ();
 sg13g2_fill_2 FILLER_7_1721 ();
 sg13g2_fill_2 FILLER_7_1741 ();
 sg13g2_fill_1 FILLER_7_1743 ();
 sg13g2_decap_4 FILLER_7_1748 ();
 sg13g2_fill_1 FILLER_7_1760 ();
 sg13g2_fill_2 FILLER_7_1797 ();
 sg13g2_fill_2 FILLER_7_1825 ();
 sg13g2_fill_2 FILLER_7_1853 ();
 sg13g2_fill_1 FILLER_7_1855 ();
 sg13g2_decap_8 FILLER_7_1876 ();
 sg13g2_decap_8 FILLER_7_1883 ();
 sg13g2_fill_2 FILLER_7_1890 ();
 sg13g2_fill_1 FILLER_7_1892 ();
 sg13g2_decap_8 FILLER_7_1929 ();
 sg13g2_fill_2 FILLER_7_1959 ();
 sg13g2_fill_1 FILLER_7_1961 ();
 sg13g2_decap_8 FILLER_7_1998 ();
 sg13g2_fill_1 FILLER_7_2005 ();
 sg13g2_decap_4 FILLER_7_2046 ();
 sg13g2_fill_2 FILLER_7_2050 ();
 sg13g2_decap_4 FILLER_7_2108 ();
 sg13g2_fill_2 FILLER_7_2168 ();
 sg13g2_decap_4 FILLER_7_2242 ();
 sg13g2_fill_2 FILLER_7_2317 ();
 sg13g2_fill_1 FILLER_7_2352 ();
 sg13g2_fill_1 FILLER_7_2379 ();
 sg13g2_fill_1 FILLER_7_2422 ();
 sg13g2_fill_2 FILLER_7_2462 ();
 sg13g2_fill_1 FILLER_7_2464 ();
 sg13g2_fill_1 FILLER_7_2501 ();
 sg13g2_decap_8 FILLER_7_2538 ();
 sg13g2_decap_8 FILLER_7_2545 ();
 sg13g2_decap_8 FILLER_7_2552 ();
 sg13g2_decap_8 FILLER_7_2559 ();
 sg13g2_decap_8 FILLER_7_2566 ();
 sg13g2_decap_8 FILLER_7_2573 ();
 sg13g2_decap_8 FILLER_7_2580 ();
 sg13g2_decap_8 FILLER_7_2587 ();
 sg13g2_decap_8 FILLER_7_2594 ();
 sg13g2_decap_8 FILLER_7_2601 ();
 sg13g2_decap_8 FILLER_7_2608 ();
 sg13g2_decap_8 FILLER_7_2615 ();
 sg13g2_decap_8 FILLER_7_2622 ();
 sg13g2_decap_8 FILLER_7_2629 ();
 sg13g2_decap_8 FILLER_7_2636 ();
 sg13g2_decap_8 FILLER_7_2643 ();
 sg13g2_decap_8 FILLER_7_2650 ();
 sg13g2_decap_8 FILLER_7_2657 ();
 sg13g2_decap_4 FILLER_7_2664 ();
 sg13g2_fill_2 FILLER_7_2668 ();
 sg13g2_decap_8 FILLER_8_0 ();
 sg13g2_decap_8 FILLER_8_7 ();
 sg13g2_decap_8 FILLER_8_14 ();
 sg13g2_decap_8 FILLER_8_21 ();
 sg13g2_decap_8 FILLER_8_28 ();
 sg13g2_decap_8 FILLER_8_35 ();
 sg13g2_decap_8 FILLER_8_42 ();
 sg13g2_decap_8 FILLER_8_49 ();
 sg13g2_decap_8 FILLER_8_56 ();
 sg13g2_fill_2 FILLER_8_63 ();
 sg13g2_decap_8 FILLER_8_69 ();
 sg13g2_fill_2 FILLER_8_76 ();
 sg13g2_decap_4 FILLER_8_82 ();
 sg13g2_decap_8 FILLER_8_96 ();
 sg13g2_fill_2 FILLER_8_116 ();
 sg13g2_decap_4 FILLER_8_131 ();
 sg13g2_fill_1 FILLER_8_149 ();
 sg13g2_decap_4 FILLER_8_181 ();
 sg13g2_fill_2 FILLER_8_185 ();
 sg13g2_fill_1 FILLER_8_248 ();
 sg13g2_fill_2 FILLER_8_261 ();
 sg13g2_fill_1 FILLER_8_286 ();
 sg13g2_fill_1 FILLER_8_344 ();
 sg13g2_fill_1 FILLER_8_378 ();
 sg13g2_fill_2 FILLER_8_410 ();
 sg13g2_fill_1 FILLER_8_424 ();
 sg13g2_fill_2 FILLER_8_438 ();
 sg13g2_fill_2 FILLER_8_449 ();
 sg13g2_fill_2 FILLER_8_469 ();
 sg13g2_fill_1 FILLER_8_515 ();
 sg13g2_fill_1 FILLER_8_521 ();
 sg13g2_fill_2 FILLER_8_548 ();
 sg13g2_fill_1 FILLER_8_609 ();
 sg13g2_fill_1 FILLER_8_670 ();
 sg13g2_fill_2 FILLER_8_684 ();
 sg13g2_fill_2 FILLER_8_692 ();
 sg13g2_fill_1 FILLER_8_714 ();
 sg13g2_fill_2 FILLER_8_755 ();
 sg13g2_fill_1 FILLER_8_757 ();
 sg13g2_fill_1 FILLER_8_768 ();
 sg13g2_fill_2 FILLER_8_786 ();
 sg13g2_fill_1 FILLER_8_788 ();
 sg13g2_decap_8 FILLER_8_798 ();
 sg13g2_decap_8 FILLER_8_805 ();
 sg13g2_decap_4 FILLER_8_812 ();
 sg13g2_fill_2 FILLER_8_865 ();
 sg13g2_fill_1 FILLER_8_867 ();
 sg13g2_fill_2 FILLER_8_894 ();
 sg13g2_fill_1 FILLER_8_896 ();
 sg13g2_decap_8 FILLER_8_917 ();
 sg13g2_fill_2 FILLER_8_924 ();
 sg13g2_fill_1 FILLER_8_926 ();
 sg13g2_decap_8 FILLER_8_957 ();
 sg13g2_decap_8 FILLER_8_964 ();
 sg13g2_fill_1 FILLER_8_989 ();
 sg13g2_fill_2 FILLER_8_1011 ();
 sg13g2_fill_1 FILLER_8_1018 ();
 sg13g2_decap_8 FILLER_8_1078 ();
 sg13g2_fill_2 FILLER_8_1085 ();
 sg13g2_fill_1 FILLER_8_1091 ();
 sg13g2_fill_1 FILLER_8_1101 ();
 sg13g2_decap_8 FILLER_8_1106 ();
 sg13g2_decap_8 FILLER_8_1113 ();
 sg13g2_decap_8 FILLER_8_1120 ();
 sg13g2_decap_8 FILLER_8_1127 ();
 sg13g2_decap_8 FILLER_8_1134 ();
 sg13g2_fill_2 FILLER_8_1141 ();
 sg13g2_fill_1 FILLER_8_1143 ();
 sg13g2_decap_4 FILLER_8_1152 ();
 sg13g2_decap_8 FILLER_8_1181 ();
 sg13g2_fill_2 FILLER_8_1188 ();
 sg13g2_fill_2 FILLER_8_1221 ();
 sg13g2_fill_1 FILLER_8_1223 ();
 sg13g2_decap_8 FILLER_8_1236 ();
 sg13g2_decap_4 FILLER_8_1243 ();
 sg13g2_fill_1 FILLER_8_1247 ();
 sg13g2_decap_4 FILLER_8_1252 ();
 sg13g2_decap_8 FILLER_8_1260 ();
 sg13g2_fill_2 FILLER_8_1267 ();
 sg13g2_fill_2 FILLER_8_1274 ();
 sg13g2_fill_1 FILLER_8_1276 ();
 sg13g2_fill_2 FILLER_8_1314 ();
 sg13g2_fill_1 FILLER_8_1316 ();
 sg13g2_fill_1 FILLER_8_1322 ();
 sg13g2_fill_2 FILLER_8_1331 ();
 sg13g2_fill_1 FILLER_8_1359 ();
 sg13g2_decap_8 FILLER_8_1364 ();
 sg13g2_fill_1 FILLER_8_1371 ();
 sg13g2_fill_1 FILLER_8_1428 ();
 sg13g2_fill_2 FILLER_8_1500 ();
 sg13g2_fill_1 FILLER_8_1502 ();
 sg13g2_fill_1 FILLER_8_1507 ();
 sg13g2_decap_8 FILLER_8_1512 ();
 sg13g2_fill_2 FILLER_8_1519 ();
 sg13g2_fill_1 FILLER_8_1539 ();
 sg13g2_fill_1 FILLER_8_1552 ();
 sg13g2_fill_1 FILLER_8_1575 ();
 sg13g2_fill_1 FILLER_8_1602 ();
 sg13g2_decap_4 FILLER_8_1677 ();
 sg13g2_fill_2 FILLER_8_1687 ();
 sg13g2_fill_1 FILLER_8_1689 ();
 sg13g2_fill_2 FILLER_8_1720 ();
 sg13g2_decap_8 FILLER_8_1727 ();
 sg13g2_fill_2 FILLER_8_1734 ();
 sg13g2_fill_1 FILLER_8_1736 ();
 sg13g2_fill_2 FILLER_8_1767 ();
 sg13g2_decap_4 FILLER_8_1783 ();
 sg13g2_fill_2 FILLER_8_1787 ();
 sg13g2_fill_1 FILLER_8_1793 ();
 sg13g2_fill_1 FILLER_8_1812 ();
 sg13g2_fill_1 FILLER_8_1843 ();
 sg13g2_decap_8 FILLER_8_1848 ();
 sg13g2_fill_2 FILLER_8_1855 ();
 sg13g2_fill_1 FILLER_8_1857 ();
 sg13g2_decap_4 FILLER_8_1892 ();
 sg13g2_fill_2 FILLER_8_1896 ();
 sg13g2_decap_4 FILLER_8_1944 ();
 sg13g2_fill_2 FILLER_8_1948 ();
 sg13g2_fill_2 FILLER_8_1966 ();
 sg13g2_decap_8 FILLER_8_1972 ();
 sg13g2_fill_2 FILLER_8_1979 ();
 sg13g2_fill_1 FILLER_8_1981 ();
 sg13g2_fill_1 FILLER_8_1986 ();
 sg13g2_fill_1 FILLER_8_2008 ();
 sg13g2_fill_2 FILLER_8_2045 ();
 sg13g2_fill_2 FILLER_8_2057 ();
 sg13g2_fill_1 FILLER_8_2059 ();
 sg13g2_fill_2 FILLER_8_2064 ();
 sg13g2_fill_1 FILLER_8_2066 ();
 sg13g2_fill_2 FILLER_8_2071 ();
 sg13g2_fill_1 FILLER_8_2073 ();
 sg13g2_fill_1 FILLER_8_2116 ();
 sg13g2_fill_2 FILLER_8_2147 ();
 sg13g2_fill_2 FILLER_8_2217 ();
 sg13g2_fill_1 FILLER_8_2219 ();
 sg13g2_fill_2 FILLER_8_2244 ();
 sg13g2_fill_1 FILLER_8_2267 ();
 sg13g2_fill_1 FILLER_8_2292 ();
 sg13g2_fill_2 FILLER_8_2308 ();
 sg13g2_fill_1 FILLER_8_2314 ();
 sg13g2_fill_2 FILLER_8_2341 ();
 sg13g2_fill_1 FILLER_8_2365 ();
 sg13g2_fill_1 FILLER_8_2458 ();
 sg13g2_decap_8 FILLER_8_2551 ();
 sg13g2_decap_8 FILLER_8_2558 ();
 sg13g2_decap_8 FILLER_8_2565 ();
 sg13g2_decap_8 FILLER_8_2572 ();
 sg13g2_decap_8 FILLER_8_2579 ();
 sg13g2_decap_8 FILLER_8_2586 ();
 sg13g2_decap_8 FILLER_8_2593 ();
 sg13g2_decap_8 FILLER_8_2600 ();
 sg13g2_decap_8 FILLER_8_2607 ();
 sg13g2_decap_8 FILLER_8_2614 ();
 sg13g2_decap_8 FILLER_8_2621 ();
 sg13g2_decap_8 FILLER_8_2628 ();
 sg13g2_decap_8 FILLER_8_2635 ();
 sg13g2_decap_8 FILLER_8_2642 ();
 sg13g2_decap_8 FILLER_8_2649 ();
 sg13g2_decap_8 FILLER_8_2656 ();
 sg13g2_decap_8 FILLER_8_2663 ();
 sg13g2_decap_8 FILLER_9_0 ();
 sg13g2_decap_8 FILLER_9_7 ();
 sg13g2_decap_8 FILLER_9_14 ();
 sg13g2_decap_8 FILLER_9_21 ();
 sg13g2_decap_8 FILLER_9_28 ();
 sg13g2_decap_8 FILLER_9_35 ();
 sg13g2_decap_8 FILLER_9_42 ();
 sg13g2_decap_8 FILLER_9_49 ();
 sg13g2_decap_8 FILLER_9_56 ();
 sg13g2_decap_8 FILLER_9_63 ();
 sg13g2_decap_4 FILLER_9_88 ();
 sg13g2_fill_1 FILLER_9_92 ();
 sg13g2_fill_1 FILLER_9_97 ();
 sg13g2_decap_8 FILLER_9_102 ();
 sg13g2_fill_2 FILLER_9_109 ();
 sg13g2_fill_1 FILLER_9_120 ();
 sg13g2_fill_1 FILLER_9_161 ();
 sg13g2_decap_4 FILLER_9_188 ();
 sg13g2_fill_2 FILLER_9_201 ();
 sg13g2_fill_2 FILLER_9_229 ();
 sg13g2_decap_8 FILLER_9_235 ();
 sg13g2_fill_2 FILLER_9_253 ();
 sg13g2_fill_1 FILLER_9_269 ();
 sg13g2_fill_2 FILLER_9_276 ();
 sg13g2_fill_1 FILLER_9_290 ();
 sg13g2_fill_1 FILLER_9_307 ();
 sg13g2_fill_1 FILLER_9_322 ();
 sg13g2_fill_1 FILLER_9_328 ();
 sg13g2_fill_2 FILLER_9_333 ();
 sg13g2_fill_2 FILLER_9_374 ();
 sg13g2_fill_2 FILLER_9_438 ();
 sg13g2_fill_1 FILLER_9_477 ();
 sg13g2_fill_1 FILLER_9_494 ();
 sg13g2_fill_1 FILLER_9_499 ();
 sg13g2_fill_1 FILLER_9_505 ();
 sg13g2_fill_2 FILLER_9_511 ();
 sg13g2_fill_1 FILLER_9_517 ();
 sg13g2_fill_2 FILLER_9_523 ();
 sg13g2_decap_4 FILLER_9_551 ();
 sg13g2_fill_1 FILLER_9_564 ();
 sg13g2_fill_2 FILLER_9_570 ();
 sg13g2_fill_2 FILLER_9_586 ();
 sg13g2_fill_1 FILLER_9_610 ();
 sg13g2_fill_1 FILLER_9_644 ();
 sg13g2_fill_1 FILLER_9_665 ();
 sg13g2_fill_2 FILLER_9_696 ();
 sg13g2_fill_2 FILLER_9_751 ();
 sg13g2_fill_2 FILLER_9_788 ();
 sg13g2_decap_4 FILLER_9_816 ();
 sg13g2_fill_2 FILLER_9_828 ();
 sg13g2_fill_1 FILLER_9_830 ();
 sg13g2_fill_1 FILLER_9_841 ();
 sg13g2_fill_2 FILLER_9_863 ();
 sg13g2_fill_1 FILLER_9_865 ();
 sg13g2_fill_2 FILLER_9_922 ();
 sg13g2_fill_2 FILLER_9_995 ();
 sg13g2_fill_2 FILLER_9_1018 ();
 sg13g2_fill_2 FILLER_9_1024 ();
 sg13g2_fill_2 FILLER_9_1047 ();
 sg13g2_fill_2 FILLER_9_1071 ();
 sg13g2_fill_1 FILLER_9_1073 ();
 sg13g2_decap_4 FILLER_9_1079 ();
 sg13g2_decap_8 FILLER_9_1118 ();
 sg13g2_decap_8 FILLER_9_1125 ();
 sg13g2_fill_2 FILLER_9_1132 ();
 sg13g2_fill_1 FILLER_9_1134 ();
 sg13g2_decap_4 FILLER_9_1139 ();
 sg13g2_fill_1 FILLER_9_1143 ();
 sg13g2_decap_4 FILLER_9_1157 ();
 sg13g2_decap_8 FILLER_9_1182 ();
 sg13g2_decap_4 FILLER_9_1189 ();
 sg13g2_fill_2 FILLER_9_1193 ();
 sg13g2_decap_8 FILLER_9_1246 ();
 sg13g2_decap_8 FILLER_9_1253 ();
 sg13g2_fill_2 FILLER_9_1260 ();
 sg13g2_fill_2 FILLER_9_1274 ();
 sg13g2_fill_1 FILLER_9_1276 ();
 sg13g2_decap_8 FILLER_9_1281 ();
 sg13g2_decap_8 FILLER_9_1288 ();
 sg13g2_fill_2 FILLER_9_1295 ();
 sg13g2_decap_8 FILLER_9_1322 ();
 sg13g2_fill_2 FILLER_9_1329 ();
 sg13g2_fill_1 FILLER_9_1331 ();
 sg13g2_fill_2 FILLER_9_1424 ();
 sg13g2_fill_1 FILLER_9_1456 ();
 sg13g2_fill_1 FILLER_9_1482 ();
 sg13g2_fill_2 FILLER_9_1513 ();
 sg13g2_fill_1 FILLER_9_1529 ();
 sg13g2_fill_2 FILLER_9_1551 ();
 sg13g2_fill_2 FILLER_9_1627 ();
 sg13g2_fill_1 FILLER_9_1702 ();
 sg13g2_decap_8 FILLER_9_1707 ();
 sg13g2_decap_8 FILLER_9_1714 ();
 sg13g2_decap_4 FILLER_9_1721 ();
 sg13g2_fill_2 FILLER_9_1725 ();
 sg13g2_fill_2 FILLER_9_1772 ();
 sg13g2_fill_1 FILLER_9_1774 ();
 sg13g2_decap_8 FILLER_9_1779 ();
 sg13g2_fill_1 FILLER_9_1798 ();
 sg13g2_fill_2 FILLER_9_1803 ();
 sg13g2_fill_1 FILLER_9_1805 ();
 sg13g2_fill_1 FILLER_9_1821 ();
 sg13g2_fill_2 FILLER_9_1848 ();
 sg13g2_fill_2 FILLER_9_1876 ();
 sg13g2_fill_2 FILLER_9_1904 ();
 sg13g2_fill_1 FILLER_9_1942 ();
 sg13g2_decap_4 FILLER_9_1979 ();
 sg13g2_decap_8 FILLER_9_1995 ();
 sg13g2_decap_8 FILLER_9_2036 ();
 sg13g2_decap_8 FILLER_9_2043 ();
 sg13g2_fill_2 FILLER_9_2050 ();
 sg13g2_fill_1 FILLER_9_2052 ();
 sg13g2_decap_8 FILLER_9_2061 ();
 sg13g2_fill_1 FILLER_9_2068 ();
 sg13g2_decap_8 FILLER_9_2077 ();
 sg13g2_decap_8 FILLER_9_2084 ();
 sg13g2_decap_8 FILLER_9_2091 ();
 sg13g2_fill_2 FILLER_9_2098 ();
 sg13g2_decap_8 FILLER_9_2116 ();
 sg13g2_fill_2 FILLER_9_2127 ();
 sg13g2_fill_2 FILLER_9_2159 ();
 sg13g2_fill_1 FILLER_9_2184 ();
 sg13g2_fill_2 FILLER_9_2253 ();
 sg13g2_fill_2 FILLER_9_2259 ();
 sg13g2_decap_4 FILLER_9_2327 ();
 sg13g2_fill_1 FILLER_9_2357 ();
 sg13g2_fill_2 FILLER_9_2380 ();
 sg13g2_fill_1 FILLER_9_2385 ();
 sg13g2_fill_2 FILLER_9_2412 ();
 sg13g2_fill_2 FILLER_9_2473 ();
 sg13g2_fill_2 FILLER_9_2501 ();
 sg13g2_decap_8 FILLER_9_2575 ();
 sg13g2_decap_8 FILLER_9_2582 ();
 sg13g2_decap_8 FILLER_9_2589 ();
 sg13g2_decap_8 FILLER_9_2596 ();
 sg13g2_decap_8 FILLER_9_2603 ();
 sg13g2_decap_8 FILLER_9_2610 ();
 sg13g2_decap_8 FILLER_9_2617 ();
 sg13g2_decap_8 FILLER_9_2624 ();
 sg13g2_decap_8 FILLER_9_2631 ();
 sg13g2_decap_8 FILLER_9_2638 ();
 sg13g2_decap_8 FILLER_9_2645 ();
 sg13g2_decap_8 FILLER_9_2652 ();
 sg13g2_decap_8 FILLER_9_2659 ();
 sg13g2_decap_4 FILLER_9_2666 ();
 sg13g2_decap_8 FILLER_10_0 ();
 sg13g2_decap_8 FILLER_10_7 ();
 sg13g2_decap_8 FILLER_10_14 ();
 sg13g2_decap_8 FILLER_10_21 ();
 sg13g2_decap_8 FILLER_10_28 ();
 sg13g2_decap_8 FILLER_10_35 ();
 sg13g2_decap_8 FILLER_10_42 ();
 sg13g2_decap_8 FILLER_10_49 ();
 sg13g2_decap_8 FILLER_10_56 ();
 sg13g2_decap_8 FILLER_10_63 ();
 sg13g2_decap_8 FILLER_10_70 ();
 sg13g2_decap_4 FILLER_10_77 ();
 sg13g2_fill_1 FILLER_10_81 ();
 sg13g2_decap_4 FILLER_10_126 ();
 sg13g2_fill_2 FILLER_10_134 ();
 sg13g2_fill_1 FILLER_10_136 ();
 sg13g2_decap_8 FILLER_10_150 ();
 sg13g2_decap_8 FILLER_10_157 ();
 sg13g2_fill_1 FILLER_10_164 ();
 sg13g2_fill_1 FILLER_10_178 ();
 sg13g2_fill_2 FILLER_10_223 ();
 sg13g2_fill_1 FILLER_10_225 ();
 sg13g2_fill_2 FILLER_10_230 ();
 sg13g2_decap_8 FILLER_10_240 ();
 sg13g2_fill_1 FILLER_10_258 ();
 sg13g2_fill_1 FILLER_10_281 ();
 sg13g2_decap_4 FILLER_10_287 ();
 sg13g2_fill_1 FILLER_10_291 ();
 sg13g2_fill_2 FILLER_10_296 ();
 sg13g2_fill_1 FILLER_10_298 ();
 sg13g2_decap_8 FILLER_10_313 ();
 sg13g2_fill_2 FILLER_10_320 ();
 sg13g2_fill_1 FILLER_10_322 ();
 sg13g2_decap_8 FILLER_10_327 ();
 sg13g2_decap_4 FILLER_10_334 ();
 sg13g2_fill_1 FILLER_10_338 ();
 sg13g2_fill_2 FILLER_10_343 ();
 sg13g2_fill_2 FILLER_10_363 ();
 sg13g2_fill_2 FILLER_10_386 ();
 sg13g2_fill_1 FILLER_10_486 ();
 sg13g2_fill_2 FILLER_10_512 ();
 sg13g2_decap_4 FILLER_10_546 ();
 sg13g2_fill_1 FILLER_10_562 ();
 sg13g2_fill_1 FILLER_10_573 ();
 sg13g2_fill_2 FILLER_10_587 ();
 sg13g2_fill_1 FILLER_10_594 ();
 sg13g2_fill_2 FILLER_10_636 ();
 sg13g2_fill_2 FILLER_10_648 ();
 sg13g2_fill_1 FILLER_10_658 ();
 sg13g2_fill_1 FILLER_10_666 ();
 sg13g2_fill_1 FILLER_10_674 ();
 sg13g2_fill_2 FILLER_10_688 ();
 sg13g2_fill_2 FILLER_10_697 ();
 sg13g2_fill_1 FILLER_10_699 ();
 sg13g2_decap_8 FILLER_10_713 ();
 sg13g2_decap_4 FILLER_10_720 ();
 sg13g2_fill_1 FILLER_10_729 ();
 sg13g2_decap_8 FILLER_10_738 ();
 sg13g2_decap_4 FILLER_10_745 ();
 sg13g2_fill_1 FILLER_10_749 ();
 sg13g2_decap_4 FILLER_10_759 ();
 sg13g2_fill_1 FILLER_10_768 ();
 sg13g2_fill_2 FILLER_10_788 ();
 sg13g2_decap_8 FILLER_10_816 ();
 sg13g2_decap_8 FILLER_10_823 ();
 sg13g2_decap_4 FILLER_10_830 ();
 sg13g2_fill_1 FILLER_10_834 ();
 sg13g2_decap_8 FILLER_10_840 ();
 sg13g2_decap_8 FILLER_10_847 ();
 sg13g2_decap_4 FILLER_10_854 ();
 sg13g2_fill_1 FILLER_10_858 ();
 sg13g2_fill_2 FILLER_10_899 ();
 sg13g2_fill_2 FILLER_10_937 ();
 sg13g2_fill_1 FILLER_10_939 ();
 sg13g2_fill_2 FILLER_10_974 ();
 sg13g2_fill_1 FILLER_10_976 ();
 sg13g2_fill_2 FILLER_10_1011 ();
 sg13g2_fill_1 FILLER_10_1013 ();
 sg13g2_decap_4 FILLER_10_1019 ();
 sg13g2_fill_1 FILLER_10_1023 ();
 sg13g2_decap_4 FILLER_10_1050 ();
 sg13g2_fill_1 FILLER_10_1054 ();
 sg13g2_fill_1 FILLER_10_1107 ();
 sg13g2_fill_2 FILLER_10_1112 ();
 sg13g2_fill_1 FILLER_10_1118 ();
 sg13g2_fill_2 FILLER_10_1123 ();
 sg13g2_fill_1 FILLER_10_1125 ();
 sg13g2_fill_1 FILLER_10_1151 ();
 sg13g2_decap_4 FILLER_10_1232 ();
 sg13g2_fill_1 FILLER_10_1257 ();
 sg13g2_fill_1 FILLER_10_1263 ();
 sg13g2_fill_2 FILLER_10_1295 ();
 sg13g2_fill_1 FILLER_10_1297 ();
 sg13g2_fill_2 FILLER_10_1329 ();
 sg13g2_fill_2 FILLER_10_1357 ();
 sg13g2_fill_1 FILLER_10_1363 ();
 sg13g2_decap_8 FILLER_10_1378 ();
 sg13g2_decap_4 FILLER_10_1389 ();
 sg13g2_fill_1 FILLER_10_1393 ();
 sg13g2_fill_1 FILLER_10_1404 ();
 sg13g2_fill_1 FILLER_10_1457 ();
 sg13g2_decap_4 FILLER_10_1503 ();
 sg13g2_fill_2 FILLER_10_1507 ();
 sg13g2_decap_4 FILLER_10_1513 ();
 sg13g2_fill_2 FILLER_10_1555 ();
 sg13g2_fill_1 FILLER_10_1620 ();
 sg13g2_fill_2 FILLER_10_1667 ();
 sg13g2_fill_1 FILLER_10_1690 ();
 sg13g2_decap_8 FILLER_10_1695 ();
 sg13g2_decap_8 FILLER_10_1712 ();
 sg13g2_decap_4 FILLER_10_1719 ();
 sg13g2_decap_4 FILLER_10_1728 ();
 sg13g2_decap_4 FILLER_10_1736 ();
 sg13g2_fill_1 FILLER_10_1740 ();
 sg13g2_decap_4 FILLER_10_1770 ();
 sg13g2_fill_1 FILLER_10_1774 ();
 sg13g2_fill_2 FILLER_10_1780 ();
 sg13g2_fill_1 FILLER_10_1782 ();
 sg13g2_decap_4 FILLER_10_1807 ();
 sg13g2_fill_1 FILLER_10_1811 ();
 sg13g2_decap_8 FILLER_10_1816 ();
 sg13g2_fill_1 FILLER_10_1823 ();
 sg13g2_decap_8 FILLER_10_1832 ();
 sg13g2_decap_8 FILLER_10_1839 ();
 sg13g2_fill_1 FILLER_10_1938 ();
 sg13g2_decap_8 FILLER_10_1954 ();
 sg13g2_decap_8 FILLER_10_1961 ();
 sg13g2_decap_4 FILLER_10_1968 ();
 sg13g2_fill_2 FILLER_10_1982 ();
 sg13g2_decap_8 FILLER_10_2006 ();
 sg13g2_fill_2 FILLER_10_2035 ();
 sg13g2_fill_1 FILLER_10_2037 ();
 sg13g2_fill_2 FILLER_10_2068 ();
 sg13g2_fill_1 FILLER_10_2070 ();
 sg13g2_fill_2 FILLER_10_2138 ();
 sg13g2_fill_1 FILLER_10_2140 ();
 sg13g2_fill_2 FILLER_10_2172 ();
 sg13g2_fill_2 FILLER_10_2204 ();
 sg13g2_fill_2 FILLER_10_2255 ();
 sg13g2_decap_4 FILLER_10_2267 ();
 sg13g2_fill_2 FILLER_10_2271 ();
 sg13g2_fill_2 FILLER_10_2277 ();
 sg13g2_fill_2 FILLER_10_2283 ();
 sg13g2_fill_2 FILLER_10_2291 ();
 sg13g2_fill_2 FILLER_10_2322 ();
 sg13g2_fill_2 FILLER_10_2344 ();
 sg13g2_fill_2 FILLER_10_2381 ();
 sg13g2_fill_2 FILLER_10_2439 ();
 sg13g2_fill_2 FILLER_10_2474 ();
 sg13g2_fill_1 FILLER_10_2552 ();
 sg13g2_decap_8 FILLER_10_2561 ();
 sg13g2_decap_8 FILLER_10_2568 ();
 sg13g2_decap_8 FILLER_10_2575 ();
 sg13g2_decap_8 FILLER_10_2582 ();
 sg13g2_decap_8 FILLER_10_2589 ();
 sg13g2_decap_8 FILLER_10_2596 ();
 sg13g2_decap_8 FILLER_10_2603 ();
 sg13g2_decap_8 FILLER_10_2610 ();
 sg13g2_decap_8 FILLER_10_2617 ();
 sg13g2_decap_8 FILLER_10_2624 ();
 sg13g2_decap_8 FILLER_10_2631 ();
 sg13g2_decap_8 FILLER_10_2638 ();
 sg13g2_decap_8 FILLER_10_2645 ();
 sg13g2_decap_8 FILLER_10_2652 ();
 sg13g2_decap_8 FILLER_10_2659 ();
 sg13g2_decap_4 FILLER_10_2666 ();
 sg13g2_decap_8 FILLER_11_0 ();
 sg13g2_decap_8 FILLER_11_7 ();
 sg13g2_decap_8 FILLER_11_14 ();
 sg13g2_decap_8 FILLER_11_21 ();
 sg13g2_decap_8 FILLER_11_28 ();
 sg13g2_decap_8 FILLER_11_35 ();
 sg13g2_decap_8 FILLER_11_42 ();
 sg13g2_fill_2 FILLER_11_49 ();
 sg13g2_fill_1 FILLER_11_77 ();
 sg13g2_fill_2 FILLER_11_86 ();
 sg13g2_fill_2 FILLER_11_93 ();
 sg13g2_fill_2 FILLER_11_100 ();
 sg13g2_fill_1 FILLER_11_102 ();
 sg13g2_fill_2 FILLER_11_129 ();
 sg13g2_fill_1 FILLER_11_131 ();
 sg13g2_fill_2 FILLER_11_137 ();
 sg13g2_decap_8 FILLER_11_147 ();
 sg13g2_decap_4 FILLER_11_154 ();
 sg13g2_decap_8 FILLER_11_162 ();
 sg13g2_fill_1 FILLER_11_169 ();
 sg13g2_fill_2 FILLER_11_230 ();
 sg13g2_fill_2 FILLER_11_236 ();
 sg13g2_fill_2 FILLER_11_242 ();
 sg13g2_fill_2 FILLER_11_253 ();
 sg13g2_decap_8 FILLER_11_277 ();
 sg13g2_decap_4 FILLER_11_284 ();
 sg13g2_fill_1 FILLER_11_288 ();
 sg13g2_fill_1 FILLER_11_322 ();
 sg13g2_fill_2 FILLER_11_336 ();
 sg13g2_fill_2 FILLER_11_350 ();
 sg13g2_decap_4 FILLER_11_356 ();
 sg13g2_fill_1 FILLER_11_360 ();
 sg13g2_fill_1 FILLER_11_380 ();
 sg13g2_fill_2 FILLER_11_412 ();
 sg13g2_fill_1 FILLER_11_448 ();
 sg13g2_fill_2 FILLER_11_497 ();
 sg13g2_fill_1 FILLER_11_589 ();
 sg13g2_fill_2 FILLER_11_621 ();
 sg13g2_fill_2 FILLER_11_657 ();
 sg13g2_fill_1 FILLER_11_666 ();
 sg13g2_fill_2 FILLER_11_708 ();
 sg13g2_fill_1 FILLER_11_710 ();
 sg13g2_decap_8 FILLER_11_737 ();
 sg13g2_decap_8 FILLER_11_744 ();
 sg13g2_fill_1 FILLER_11_751 ();
 sg13g2_decap_4 FILLER_11_761 ();
 sg13g2_fill_1 FILLER_11_765 ();
 sg13g2_fill_2 FILLER_11_776 ();
 sg13g2_fill_1 FILLER_11_778 ();
 sg13g2_fill_2 FILLER_11_784 ();
 sg13g2_fill_1 FILLER_11_786 ();
 sg13g2_decap_4 FILLER_11_792 ();
 sg13g2_decap_8 FILLER_11_804 ();
 sg13g2_decap_8 FILLER_11_811 ();
 sg13g2_decap_8 FILLER_11_818 ();
 sg13g2_decap_8 FILLER_11_825 ();
 sg13g2_decap_4 FILLER_11_832 ();
 sg13g2_fill_1 FILLER_11_836 ();
 sg13g2_fill_2 FILLER_11_881 ();
 sg13g2_fill_1 FILLER_11_969 ();
 sg13g2_fill_1 FILLER_11_984 ();
 sg13g2_fill_1 FILLER_11_989 ();
 sg13g2_fill_2 FILLER_11_1046 ();
 sg13g2_fill_1 FILLER_11_1048 ();
 sg13g2_fill_2 FILLER_11_1053 ();
 sg13g2_fill_2 FILLER_11_1099 ();
 sg13g2_fill_1 FILLER_11_1101 ();
 sg13g2_fill_1 FILLER_11_1133 ();
 sg13g2_decap_8 FILLER_11_1174 ();
 sg13g2_fill_2 FILLER_11_1181 ();
 sg13g2_fill_1 FILLER_11_1183 ();
 sg13g2_decap_8 FILLER_11_1232 ();
 sg13g2_fill_2 FILLER_11_1239 ();
 sg13g2_fill_1 FILLER_11_1271 ();
 sg13g2_fill_1 FILLER_11_1276 ();
 sg13g2_decap_8 FILLER_11_1303 ();
 sg13g2_fill_1 FILLER_11_1310 ();
 sg13g2_decap_4 FILLER_11_1315 ();
 sg13g2_fill_1 FILLER_11_1319 ();
 sg13g2_decap_4 FILLER_11_1328 ();
 sg13g2_fill_1 FILLER_11_1332 ();
 sg13g2_fill_2 FILLER_11_1372 ();
 sg13g2_fill_2 FILLER_11_1379 ();
 sg13g2_fill_1 FILLER_11_1381 ();
 sg13g2_fill_2 FILLER_11_1395 ();
 sg13g2_fill_2 FILLER_11_1424 ();
 sg13g2_decap_8 FILLER_11_1435 ();
 sg13g2_fill_1 FILLER_11_1442 ();
 sg13g2_fill_1 FILLER_11_1453 ();
 sg13g2_fill_1 FILLER_11_1458 ();
 sg13g2_fill_2 FILLER_11_1488 ();
 sg13g2_decap_8 FILLER_11_1495 ();
 sg13g2_fill_1 FILLER_11_1532 ();
 sg13g2_fill_2 FILLER_11_1576 ();
 sg13g2_fill_1 FILLER_11_1578 ();
 sg13g2_decap_4 FILLER_11_1590 ();
 sg13g2_fill_1 FILLER_11_1594 ();
 sg13g2_fill_1 FILLER_11_1613 ();
 sg13g2_fill_2 FILLER_11_1621 ();
 sg13g2_fill_2 FILLER_11_1634 ();
 sg13g2_decap_4 FILLER_11_1667 ();
 sg13g2_fill_2 FILLER_11_1681 ();
 sg13g2_decap_8 FILLER_11_1719 ();
 sg13g2_decap_8 FILLER_11_1726 ();
 sg13g2_decap_8 FILLER_11_1733 ();
 sg13g2_decap_4 FILLER_11_1740 ();
 sg13g2_fill_1 FILLER_11_1744 ();
 sg13g2_fill_2 FILLER_11_1764 ();
 sg13g2_decap_8 FILLER_11_1830 ();
 sg13g2_decap_8 FILLER_11_1837 ();
 sg13g2_fill_2 FILLER_11_1844 ();
 sg13g2_fill_1 FILLER_11_1846 ();
 sg13g2_decap_8 FILLER_11_1868 ();
 sg13g2_fill_1 FILLER_11_1875 ();
 sg13g2_fill_2 FILLER_11_1912 ();
 sg13g2_decap_8 FILLER_11_1918 ();
 sg13g2_decap_8 FILLER_11_1925 ();
 sg13g2_decap_8 FILLER_11_1932 ();
 sg13g2_decap_4 FILLER_11_1943 ();
 sg13g2_fill_1 FILLER_11_2009 ();
 sg13g2_fill_2 FILLER_11_2031 ();
 sg13g2_fill_2 FILLER_11_2069 ();
 sg13g2_fill_1 FILLER_11_2097 ();
 sg13g2_fill_2 FILLER_11_2124 ();
 sg13g2_fill_2 FILLER_11_2181 ();
 sg13g2_fill_2 FILLER_11_2200 ();
 sg13g2_fill_2 FILLER_11_2224 ();
 sg13g2_decap_8 FILLER_11_2252 ();
 sg13g2_decap_8 FILLER_11_2259 ();
 sg13g2_decap_8 FILLER_11_2266 ();
 sg13g2_fill_2 FILLER_11_2273 ();
 sg13g2_fill_1 FILLER_11_2275 ();
 sg13g2_fill_1 FILLER_11_2338 ();
 sg13g2_fill_2 FILLER_11_2372 ();
 sg13g2_fill_2 FILLER_11_2390 ();
 sg13g2_fill_1 FILLER_11_2421 ();
 sg13g2_fill_1 FILLER_11_2458 ();
 sg13g2_fill_2 FILLER_11_2476 ();
 sg13g2_fill_1 FILLER_11_2533 ();
 sg13g2_decap_8 FILLER_11_2560 ();
 sg13g2_decap_8 FILLER_11_2567 ();
 sg13g2_decap_8 FILLER_11_2574 ();
 sg13g2_decap_8 FILLER_11_2581 ();
 sg13g2_decap_8 FILLER_11_2588 ();
 sg13g2_decap_8 FILLER_11_2595 ();
 sg13g2_decap_8 FILLER_11_2602 ();
 sg13g2_decap_8 FILLER_11_2609 ();
 sg13g2_decap_8 FILLER_11_2616 ();
 sg13g2_decap_8 FILLER_11_2623 ();
 sg13g2_decap_8 FILLER_11_2630 ();
 sg13g2_decap_8 FILLER_11_2637 ();
 sg13g2_decap_8 FILLER_11_2644 ();
 sg13g2_decap_8 FILLER_11_2651 ();
 sg13g2_decap_8 FILLER_11_2658 ();
 sg13g2_decap_4 FILLER_11_2665 ();
 sg13g2_fill_1 FILLER_11_2669 ();
 sg13g2_decap_8 FILLER_12_0 ();
 sg13g2_decap_8 FILLER_12_7 ();
 sg13g2_decap_8 FILLER_12_14 ();
 sg13g2_decap_8 FILLER_12_21 ();
 sg13g2_decap_8 FILLER_12_28 ();
 sg13g2_decap_8 FILLER_12_35 ();
 sg13g2_decap_8 FILLER_12_42 ();
 sg13g2_decap_8 FILLER_12_49 ();
 sg13g2_fill_1 FILLER_12_56 ();
 sg13g2_decap_8 FILLER_12_61 ();
 sg13g2_decap_8 FILLER_12_68 ();
 sg13g2_fill_2 FILLER_12_75 ();
 sg13g2_fill_1 FILLER_12_77 ();
 sg13g2_fill_2 FILLER_12_82 ();
 sg13g2_fill_2 FILLER_12_89 ();
 sg13g2_fill_1 FILLER_12_91 ();
 sg13g2_fill_1 FILLER_12_100 ();
 sg13g2_fill_1 FILLER_12_106 ();
 sg13g2_fill_1 FILLER_12_119 ();
 sg13g2_decap_8 FILLER_12_159 ();
 sg13g2_decap_8 FILLER_12_166 ();
 sg13g2_decap_4 FILLER_12_173 ();
 sg13g2_decap_8 FILLER_12_181 ();
 sg13g2_decap_8 FILLER_12_188 ();
 sg13g2_decap_8 FILLER_12_195 ();
 sg13g2_decap_4 FILLER_12_202 ();
 sg13g2_fill_1 FILLER_12_240 ();
 sg13g2_decap_4 FILLER_12_245 ();
 sg13g2_fill_2 FILLER_12_257 ();
 sg13g2_fill_2 FILLER_12_267 ();
 sg13g2_fill_1 FILLER_12_269 ();
 sg13g2_fill_1 FILLER_12_276 ();
 sg13g2_fill_2 FILLER_12_296 ();
 sg13g2_fill_1 FILLER_12_303 ();
 sg13g2_fill_2 FILLER_12_308 ();
 sg13g2_fill_1 FILLER_12_310 ();
 sg13g2_decap_4 FILLER_12_347 ();
 sg13g2_fill_2 FILLER_12_361 ();
 sg13g2_fill_2 FILLER_12_417 ();
 sg13g2_fill_2 FILLER_12_453 ();
 sg13g2_fill_2 FILLER_12_458 ();
 sg13g2_fill_1 FILLER_12_465 ();
 sg13g2_fill_2 FILLER_12_541 ();
 sg13g2_fill_1 FILLER_12_623 ();
 sg13g2_fill_1 FILLER_12_634 ();
 sg13g2_fill_2 FILLER_12_638 ();
 sg13g2_fill_1 FILLER_12_649 ();
 sg13g2_fill_1 FILLER_12_710 ();
 sg13g2_fill_2 FILLER_12_716 ();
 sg13g2_decap_4 FILLER_12_749 ();
 sg13g2_fill_1 FILLER_12_757 ();
 sg13g2_fill_2 FILLER_12_762 ();
 sg13g2_fill_1 FILLER_12_764 ();
 sg13g2_fill_2 FILLER_12_773 ();
 sg13g2_decap_4 FILLER_12_779 ();
 sg13g2_fill_1 FILLER_12_783 ();
 sg13g2_decap_8 FILLER_12_788 ();
 sg13g2_decap_8 FILLER_12_795 ();
 sg13g2_decap_8 FILLER_12_802 ();
 sg13g2_fill_1 FILLER_12_865 ();
 sg13g2_decap_8 FILLER_12_902 ();
 sg13g2_decap_8 FILLER_12_909 ();
 sg13g2_decap_8 FILLER_12_961 ();
 sg13g2_fill_2 FILLER_12_972 ();
 sg13g2_fill_1 FILLER_12_974 ();
 sg13g2_decap_8 FILLER_12_1010 ();
 sg13g2_fill_2 FILLER_12_1017 ();
 sg13g2_fill_1 FILLER_12_1037 ();
 sg13g2_fill_1 FILLER_12_1047 ();
 sg13g2_decap_4 FILLER_12_1077 ();
 sg13g2_fill_2 FILLER_12_1138 ();
 sg13g2_fill_1 FILLER_12_1140 ();
 sg13g2_fill_1 FILLER_12_1167 ();
 sg13g2_fill_2 FILLER_12_1212 ();
 sg13g2_fill_2 FILLER_12_1240 ();
 sg13g2_fill_1 FILLER_12_1242 ();
 sg13g2_decap_8 FILLER_12_1299 ();
 sg13g2_decap_8 FILLER_12_1306 ();
 sg13g2_decap_8 FILLER_12_1317 ();
 sg13g2_fill_2 FILLER_12_1324 ();
 sg13g2_decap_8 FILLER_12_1360 ();
 sg13g2_decap_8 FILLER_12_1367 ();
 sg13g2_decap_4 FILLER_12_1374 ();
 sg13g2_fill_2 FILLER_12_1378 ();
 sg13g2_decap_8 FILLER_12_1389 ();
 sg13g2_decap_4 FILLER_12_1409 ();
 sg13g2_fill_1 FILLER_12_1413 ();
 sg13g2_fill_2 FILLER_12_1440 ();
 sg13g2_fill_1 FILLER_12_1442 ();
 sg13g2_fill_1 FILLER_12_1469 ();
 sg13g2_decap_8 FILLER_12_1496 ();
 sg13g2_decap_4 FILLER_12_1503 ();
 sg13g2_fill_2 FILLER_12_1507 ();
 sg13g2_decap_8 FILLER_12_1513 ();
 sg13g2_decap_8 FILLER_12_1520 ();
 sg13g2_fill_2 FILLER_12_1527 ();
 sg13g2_fill_1 FILLER_12_1529 ();
 sg13g2_fill_2 FILLER_12_1540 ();
 sg13g2_fill_1 FILLER_12_1542 ();
 sg13g2_fill_1 FILLER_12_1566 ();
 sg13g2_fill_1 FILLER_12_1577 ();
 sg13g2_decap_4 FILLER_12_1586 ();
 sg13g2_fill_2 FILLER_12_1590 ();
 sg13g2_decap_8 FILLER_12_1596 ();
 sg13g2_fill_2 FILLER_12_1603 ();
 sg13g2_fill_1 FILLER_12_1620 ();
 sg13g2_fill_2 FILLER_12_1624 ();
 sg13g2_fill_1 FILLER_12_1636 ();
 sg13g2_decap_8 FILLER_12_1667 ();
 sg13g2_decap_4 FILLER_12_1674 ();
 sg13g2_fill_1 FILLER_12_1678 ();
 sg13g2_fill_2 FILLER_12_1683 ();
 sg13g2_decap_8 FILLER_12_1715 ();
 sg13g2_decap_8 FILLER_12_1722 ();
 sg13g2_decap_8 FILLER_12_1729 ();
 sg13g2_fill_1 FILLER_12_1736 ();
 sg13g2_fill_1 FILLER_12_1747 ();
 sg13g2_fill_2 FILLER_12_1755 ();
 sg13g2_fill_1 FILLER_12_1782 ();
 sg13g2_fill_2 FILLER_12_1787 ();
 sg13g2_fill_1 FILLER_12_1793 ();
 sg13g2_fill_2 FILLER_12_1804 ();
 sg13g2_decap_8 FILLER_12_1832 ();
 sg13g2_decap_8 FILLER_12_1839 ();
 sg13g2_decap_4 FILLER_12_1846 ();
 sg13g2_fill_1 FILLER_12_1850 ();
 sg13g2_fill_1 FILLER_12_1859 ();
 sg13g2_decap_8 FILLER_12_1865 ();
 sg13g2_fill_2 FILLER_12_1872 ();
 sg13g2_fill_1 FILLER_12_1874 ();
 sg13g2_decap_4 FILLER_12_1885 ();
 sg13g2_decap_8 FILLER_12_1899 ();
 sg13g2_fill_1 FILLER_12_1906 ();
 sg13g2_decap_8 FILLER_12_1911 ();
 sg13g2_decap_8 FILLER_12_1918 ();
 sg13g2_decap_8 FILLER_12_1925 ();
 sg13g2_fill_1 FILLER_12_1932 ();
 sg13g2_fill_1 FILLER_12_1943 ();
 sg13g2_fill_1 FILLER_12_1980 ();
 sg13g2_fill_1 FILLER_12_1988 ();
 sg13g2_fill_1 FILLER_12_1995 ();
 sg13g2_fill_1 FILLER_12_2003 ();
 sg13g2_fill_1 FILLER_12_2015 ();
 sg13g2_fill_1 FILLER_12_2020 ();
 sg13g2_fill_2 FILLER_12_2031 ();
 sg13g2_fill_1 FILLER_12_2041 ();
 sg13g2_fill_1 FILLER_12_2108 ();
 sg13g2_fill_2 FILLER_12_2117 ();
 sg13g2_fill_1 FILLER_12_2122 ();
 sg13g2_fill_1 FILLER_12_2149 ();
 sg13g2_fill_2 FILLER_12_2154 ();
 sg13g2_fill_1 FILLER_12_2188 ();
 sg13g2_fill_2 FILLER_12_2236 ();
 sg13g2_fill_1 FILLER_12_2238 ();
 sg13g2_decap_8 FILLER_12_2265 ();
 sg13g2_fill_2 FILLER_12_2272 ();
 sg13g2_fill_1 FILLER_12_2296 ();
 sg13g2_fill_1 FILLER_12_2302 ();
 sg13g2_fill_2 FILLER_12_2316 ();
 sg13g2_fill_1 FILLER_12_2358 ();
 sg13g2_fill_1 FILLER_12_2381 ();
 sg13g2_fill_1 FILLER_12_2386 ();
 sg13g2_fill_1 FILLER_12_2393 ();
 sg13g2_fill_2 FILLER_12_2427 ();
 sg13g2_fill_2 FILLER_12_2482 ();
 sg13g2_decap_8 FILLER_12_2562 ();
 sg13g2_decap_8 FILLER_12_2569 ();
 sg13g2_decap_8 FILLER_12_2576 ();
 sg13g2_decap_8 FILLER_12_2583 ();
 sg13g2_decap_8 FILLER_12_2590 ();
 sg13g2_decap_8 FILLER_12_2597 ();
 sg13g2_decap_8 FILLER_12_2604 ();
 sg13g2_decap_8 FILLER_12_2611 ();
 sg13g2_decap_8 FILLER_12_2618 ();
 sg13g2_decap_8 FILLER_12_2625 ();
 sg13g2_decap_8 FILLER_12_2632 ();
 sg13g2_decap_8 FILLER_12_2639 ();
 sg13g2_decap_8 FILLER_12_2646 ();
 sg13g2_decap_8 FILLER_12_2653 ();
 sg13g2_decap_8 FILLER_12_2660 ();
 sg13g2_fill_2 FILLER_12_2667 ();
 sg13g2_fill_1 FILLER_12_2669 ();
 sg13g2_decap_8 FILLER_13_0 ();
 sg13g2_decap_8 FILLER_13_7 ();
 sg13g2_decap_8 FILLER_13_14 ();
 sg13g2_decap_8 FILLER_13_21 ();
 sg13g2_decap_8 FILLER_13_28 ();
 sg13g2_decap_8 FILLER_13_35 ();
 sg13g2_fill_1 FILLER_13_68 ();
 sg13g2_decap_4 FILLER_13_74 ();
 sg13g2_fill_1 FILLER_13_78 ();
 sg13g2_fill_1 FILLER_13_111 ();
 sg13g2_fill_1 FILLER_13_130 ();
 sg13g2_fill_1 FILLER_13_135 ();
 sg13g2_decap_4 FILLER_13_162 ();
 sg13g2_fill_2 FILLER_13_166 ();
 sg13g2_fill_1 FILLER_13_198 ();
 sg13g2_fill_2 FILLER_13_204 ();
 sg13g2_fill_2 FILLER_13_216 ();
 sg13g2_fill_1 FILLER_13_218 ();
 sg13g2_fill_2 FILLER_13_245 ();
 sg13g2_fill_2 FILLER_13_255 ();
 sg13g2_fill_1 FILLER_13_257 ();
 sg13g2_fill_1 FILLER_13_266 ();
 sg13g2_fill_1 FILLER_13_273 ();
 sg13g2_fill_1 FILLER_13_300 ();
 sg13g2_fill_2 FILLER_13_312 ();
 sg13g2_fill_1 FILLER_13_314 ();
 sg13g2_fill_2 FILLER_13_328 ();
 sg13g2_fill_1 FILLER_13_330 ();
 sg13g2_fill_2 FILLER_13_340 ();
 sg13g2_fill_1 FILLER_13_342 ();
 sg13g2_decap_4 FILLER_13_347 ();
 sg13g2_decap_4 FILLER_13_363 ();
 sg13g2_fill_1 FILLER_13_367 ();
 sg13g2_decap_4 FILLER_13_376 ();
 sg13g2_fill_1 FILLER_13_380 ();
 sg13g2_fill_2 FILLER_13_385 ();
 sg13g2_fill_1 FILLER_13_398 ();
 sg13g2_fill_2 FILLER_13_460 ();
 sg13g2_fill_1 FILLER_13_470 ();
 sg13g2_fill_1 FILLER_13_497 ();
 sg13g2_fill_1 FILLER_13_503 ();
 sg13g2_fill_1 FILLER_13_509 ();
 sg13g2_fill_2 FILLER_13_521 ();
 sg13g2_fill_2 FILLER_13_574 ();
 sg13g2_fill_2 FILLER_13_589 ();
 sg13g2_fill_2 FILLER_13_608 ();
 sg13g2_fill_2 FILLER_13_623 ();
 sg13g2_fill_2 FILLER_13_630 ();
 sg13g2_fill_1 FILLER_13_640 ();
 sg13g2_fill_2 FILLER_13_652 ();
 sg13g2_fill_2 FILLER_13_691 ();
 sg13g2_fill_1 FILLER_13_693 ();
 sg13g2_fill_1 FILLER_13_704 ();
 sg13g2_fill_2 FILLER_13_787 ();
 sg13g2_fill_2 FILLER_13_793 ();
 sg13g2_fill_1 FILLER_13_795 ();
 sg13g2_fill_2 FILLER_13_827 ();
 sg13g2_fill_1 FILLER_13_829 ();
 sg13g2_fill_1 FILLER_13_844 ();
 sg13g2_decap_8 FILLER_13_849 ();
 sg13g2_fill_2 FILLER_13_856 ();
 sg13g2_fill_1 FILLER_13_858 ();
 sg13g2_fill_2 FILLER_13_869 ();
 sg13g2_fill_1 FILLER_13_871 ();
 sg13g2_decap_8 FILLER_13_893 ();
 sg13g2_decap_8 FILLER_13_900 ();
 sg13g2_fill_1 FILLER_13_907 ();
 sg13g2_decap_8 FILLER_13_968 ();
 sg13g2_decap_4 FILLER_13_975 ();
 sg13g2_decap_4 FILLER_13_988 ();
 sg13g2_fill_2 FILLER_13_992 ();
 sg13g2_fill_1 FILLER_13_1003 ();
 sg13g2_decap_8 FILLER_13_1008 ();
 sg13g2_decap_8 FILLER_13_1015 ();
 sg13g2_decap_8 FILLER_13_1022 ();
 sg13g2_decap_8 FILLER_13_1029 ();
 sg13g2_decap_4 FILLER_13_1036 ();
 sg13g2_fill_2 FILLER_13_1040 ();
 sg13g2_decap_8 FILLER_13_1047 ();
 sg13g2_decap_8 FILLER_13_1071 ();
 sg13g2_fill_2 FILLER_13_1078 ();
 sg13g2_fill_1 FILLER_13_1089 ();
 sg13g2_fill_2 FILLER_13_1110 ();
 sg13g2_fill_2 FILLER_13_1133 ();
 sg13g2_fill_1 FILLER_13_1140 ();
 sg13g2_fill_1 FILLER_13_1145 ();
 sg13g2_fill_1 FILLER_13_1150 ();
 sg13g2_fill_1 FILLER_13_1156 ();
 sg13g2_fill_1 FILLER_13_1161 ();
 sg13g2_fill_1 FILLER_13_1166 ();
 sg13g2_fill_1 FILLER_13_1172 ();
 sg13g2_fill_1 FILLER_13_1177 ();
 sg13g2_decap_8 FILLER_13_1182 ();
 sg13g2_fill_2 FILLER_13_1189 ();
 sg13g2_fill_1 FILLER_13_1191 ();
 sg13g2_decap_4 FILLER_13_1226 ();
 sg13g2_fill_1 FILLER_13_1230 ();
 sg13g2_decap_8 FILLER_13_1240 ();
 sg13g2_fill_2 FILLER_13_1247 ();
 sg13g2_decap_4 FILLER_13_1274 ();
 sg13g2_fill_1 FILLER_13_1278 ();
 sg13g2_fill_2 FILLER_13_1288 ();
 sg13g2_fill_1 FILLER_13_1290 ();
 sg13g2_fill_1 FILLER_13_1335 ();
 sg13g2_fill_1 FILLER_13_1372 ();
 sg13g2_fill_1 FILLER_13_1408 ();
 sg13g2_fill_2 FILLER_13_1449 ();
 sg13g2_fill_2 FILLER_13_1469 ();
 sg13g2_fill_2 FILLER_13_1501 ();
 sg13g2_fill_1 FILLER_13_1503 ();
 sg13g2_decap_4 FILLER_13_1530 ();
 sg13g2_fill_1 FILLER_13_1559 ();
 sg13g2_fill_1 FILLER_13_1565 ();
 sg13g2_fill_2 FILLER_13_1600 ();
 sg13g2_fill_1 FILLER_13_1602 ();
 sg13g2_fill_1 FILLER_13_1642 ();
 sg13g2_fill_2 FILLER_13_1674 ();
 sg13g2_decap_4 FILLER_13_1693 ();
 sg13g2_fill_1 FILLER_13_1697 ();
 sg13g2_fill_1 FILLER_13_1702 ();
 sg13g2_decap_4 FILLER_13_1707 ();
 sg13g2_fill_2 FILLER_13_1711 ();
 sg13g2_fill_2 FILLER_13_1757 ();
 sg13g2_decap_4 FILLER_13_1768 ();
 sg13g2_fill_2 FILLER_13_1808 ();
 sg13g2_fill_1 FILLER_13_1810 ();
 sg13g2_decap_8 FILLER_13_1837 ();
 sg13g2_decap_4 FILLER_13_1844 ();
 sg13g2_fill_1 FILLER_13_1957 ();
 sg13g2_fill_2 FILLER_13_1962 ();
 sg13g2_fill_1 FILLER_13_2102 ();
 sg13g2_fill_1 FILLER_13_2118 ();
 sg13g2_fill_1 FILLER_13_2134 ();
 sg13g2_fill_1 FILLER_13_2139 ();
 sg13g2_decap_4 FILLER_13_2171 ();
 sg13g2_fill_1 FILLER_13_2175 ();
 sg13g2_decap_8 FILLER_13_2224 ();
 sg13g2_decap_8 FILLER_13_2231 ();
 sg13g2_decap_8 FILLER_13_2238 ();
 sg13g2_decap_8 FILLER_13_2249 ();
 sg13g2_decap_4 FILLER_13_2256 ();
 sg13g2_fill_2 FILLER_13_2260 ();
 sg13g2_fill_1 FILLER_13_2288 ();
 sg13g2_decap_4 FILLER_13_2308 ();
 sg13g2_fill_1 FILLER_13_2320 ();
 sg13g2_decap_8 FILLER_13_2329 ();
 sg13g2_fill_2 FILLER_13_2359 ();
 sg13g2_fill_1 FILLER_13_2368 ();
 sg13g2_fill_1 FILLER_13_2433 ();
 sg13g2_fill_1 FILLER_13_2457 ();
 sg13g2_decap_4 FILLER_13_2526 ();
 sg13g2_fill_1 FILLER_13_2530 ();
 sg13g2_fill_2 FILLER_13_2541 ();
 sg13g2_decap_8 FILLER_13_2569 ();
 sg13g2_decap_8 FILLER_13_2576 ();
 sg13g2_decap_8 FILLER_13_2583 ();
 sg13g2_decap_8 FILLER_13_2590 ();
 sg13g2_decap_8 FILLER_13_2597 ();
 sg13g2_decap_8 FILLER_13_2604 ();
 sg13g2_decap_8 FILLER_13_2611 ();
 sg13g2_decap_8 FILLER_13_2618 ();
 sg13g2_decap_8 FILLER_13_2625 ();
 sg13g2_decap_8 FILLER_13_2632 ();
 sg13g2_decap_8 FILLER_13_2639 ();
 sg13g2_decap_8 FILLER_13_2646 ();
 sg13g2_decap_8 FILLER_13_2653 ();
 sg13g2_decap_8 FILLER_13_2660 ();
 sg13g2_fill_2 FILLER_13_2667 ();
 sg13g2_fill_1 FILLER_13_2669 ();
 sg13g2_decap_8 FILLER_14_0 ();
 sg13g2_decap_8 FILLER_14_7 ();
 sg13g2_decap_8 FILLER_14_14 ();
 sg13g2_decap_8 FILLER_14_21 ();
 sg13g2_decap_8 FILLER_14_28 ();
 sg13g2_decap_8 FILLER_14_35 ();
 sg13g2_fill_2 FILLER_14_42 ();
 sg13g2_fill_1 FILLER_14_44 ();
 sg13g2_fill_1 FILLER_14_49 ();
 sg13g2_fill_1 FILLER_14_76 ();
 sg13g2_decap_8 FILLER_14_86 ();
 sg13g2_decap_4 FILLER_14_93 ();
 sg13g2_fill_2 FILLER_14_97 ();
 sg13g2_decap_8 FILLER_14_138 ();
 sg13g2_decap_8 FILLER_14_145 ();
 sg13g2_fill_2 FILLER_14_152 ();
 sg13g2_decap_8 FILLER_14_158 ();
 sg13g2_decap_8 FILLER_14_165 ();
 sg13g2_decap_8 FILLER_14_237 ();
 sg13g2_decap_8 FILLER_14_244 ();
 sg13g2_decap_4 FILLER_14_251 ();
 sg13g2_fill_2 FILLER_14_261 ();
 sg13g2_fill_1 FILLER_14_263 ();
 sg13g2_decap_4 FILLER_14_268 ();
 sg13g2_fill_1 FILLER_14_272 ();
 sg13g2_fill_1 FILLER_14_281 ();
 sg13g2_fill_1 FILLER_14_286 ();
 sg13g2_fill_2 FILLER_14_292 ();
 sg13g2_fill_1 FILLER_14_294 ();
 sg13g2_fill_1 FILLER_14_300 ();
 sg13g2_fill_2 FILLER_14_308 ();
 sg13g2_fill_1 FILLER_14_310 ();
 sg13g2_fill_1 FILLER_14_321 ();
 sg13g2_fill_1 FILLER_14_348 ();
 sg13g2_decap_4 FILLER_14_378 ();
 sg13g2_fill_2 FILLER_14_382 ();
 sg13g2_fill_1 FILLER_14_410 ();
 sg13g2_fill_1 FILLER_14_415 ();
 sg13g2_fill_1 FILLER_14_467 ();
 sg13g2_fill_2 FILLER_14_475 ();
 sg13g2_fill_2 FILLER_14_482 ();
 sg13g2_fill_2 FILLER_14_489 ();
 sg13g2_fill_1 FILLER_14_521 ();
 sg13g2_fill_2 FILLER_14_565 ();
 sg13g2_fill_1 FILLER_14_588 ();
 sg13g2_fill_1 FILLER_14_605 ();
 sg13g2_fill_2 FILLER_14_654 ();
 sg13g2_fill_2 FILLER_14_670 ();
 sg13g2_fill_1 FILLER_14_681 ();
 sg13g2_fill_1 FILLER_14_724 ();
 sg13g2_fill_1 FILLER_14_744 ();
 sg13g2_fill_2 FILLER_14_749 ();
 sg13g2_fill_1 FILLER_14_751 ();
 sg13g2_fill_1 FILLER_14_757 ();
 sg13g2_fill_1 FILLER_14_799 ();
 sg13g2_decap_4 FILLER_14_821 ();
 sg13g2_fill_2 FILLER_14_825 ();
 sg13g2_decap_8 FILLER_14_863 ();
 sg13g2_decap_4 FILLER_14_870 ();
 sg13g2_fill_2 FILLER_14_874 ();
 sg13g2_decap_8 FILLER_14_897 ();
 sg13g2_fill_2 FILLER_14_904 ();
 sg13g2_fill_2 FILLER_14_936 ();
 sg13g2_fill_1 FILLER_14_938 ();
 sg13g2_fill_1 FILLER_14_949 ();
 sg13g2_fill_2 FILLER_14_976 ();
 sg13g2_fill_1 FILLER_14_978 ();
 sg13g2_fill_2 FILLER_14_1005 ();
 sg13g2_decap_8 FILLER_14_1012 ();
 sg13g2_decap_8 FILLER_14_1019 ();
 sg13g2_decap_8 FILLER_14_1026 ();
 sg13g2_decap_4 FILLER_14_1033 ();
 sg13g2_fill_2 FILLER_14_1041 ();
 sg13g2_fill_1 FILLER_14_1043 ();
 sg13g2_fill_2 FILLER_14_1074 ();
 sg13g2_fill_1 FILLER_14_1076 ();
 sg13g2_fill_1 FILLER_14_1094 ();
 sg13g2_decap_8 FILLER_14_1099 ();
 sg13g2_fill_1 FILLER_14_1106 ();
 sg13g2_fill_2 FILLER_14_1168 ();
 sg13g2_fill_1 FILLER_14_1170 ();
 sg13g2_decap_8 FILLER_14_1192 ();
 sg13g2_decap_8 FILLER_14_1199 ();
 sg13g2_decap_8 FILLER_14_1206 ();
 sg13g2_decap_8 FILLER_14_1213 ();
 sg13g2_decap_8 FILLER_14_1220 ();
 sg13g2_fill_1 FILLER_14_1257 ();
 sg13g2_fill_2 FILLER_14_1423 ();
 sg13g2_decap_8 FILLER_14_1429 ();
 sg13g2_decap_8 FILLER_14_1436 ();
 sg13g2_decap_4 FILLER_14_1443 ();
 sg13g2_fill_1 FILLER_14_1447 ();
 sg13g2_fill_1 FILLER_14_1461 ();
 sg13g2_decap_4 FILLER_14_1472 ();
 sg13g2_fill_1 FILLER_14_1476 ();
 sg13g2_decap_8 FILLER_14_1485 ();
 sg13g2_decap_8 FILLER_14_1492 ();
 sg13g2_decap_8 FILLER_14_1499 ();
 sg13g2_fill_2 FILLER_14_1506 ();
 sg13g2_decap_4 FILLER_14_1512 ();
 sg13g2_fill_2 FILLER_14_1520 ();
 sg13g2_fill_2 FILLER_14_1526 ();
 sg13g2_decap_8 FILLER_14_1538 ();
 sg13g2_fill_2 FILLER_14_1545 ();
 sg13g2_fill_1 FILLER_14_1547 ();
 sg13g2_fill_2 FILLER_14_1553 ();
 sg13g2_fill_1 FILLER_14_1580 ();
 sg13g2_fill_1 FILLER_14_1617 ();
 sg13g2_fill_1 FILLER_14_1634 ();
 sg13g2_fill_1 FILLER_14_1639 ();
 sg13g2_decap_8 FILLER_14_1670 ();
 sg13g2_fill_1 FILLER_14_1677 ();
 sg13g2_decap_4 FILLER_14_1689 ();
 sg13g2_fill_2 FILLER_14_1693 ();
 sg13g2_decap_8 FILLER_14_1703 ();
 sg13g2_fill_2 FILLER_14_1710 ();
 sg13g2_fill_1 FILLER_14_1712 ();
 sg13g2_decap_8 FILLER_14_1718 ();
 sg13g2_fill_2 FILLER_14_1725 ();
 sg13g2_fill_1 FILLER_14_1727 ();
 sg13g2_fill_2 FILLER_14_1737 ();
 sg13g2_decap_4 FILLER_14_1758 ();
 sg13g2_fill_2 FILLER_14_1762 ();
 sg13g2_fill_2 FILLER_14_1768 ();
 sg13g2_fill_2 FILLER_14_1774 ();
 sg13g2_fill_1 FILLER_14_1812 ();
 sg13g2_decap_8 FILLER_14_1821 ();
 sg13g2_fill_2 FILLER_14_1828 ();
 sg13g2_decap_4 FILLER_14_1876 ();
 sg13g2_fill_2 FILLER_14_1880 ();
 sg13g2_fill_2 FILLER_14_1911 ();
 sg13g2_fill_1 FILLER_14_1953 ();
 sg13g2_decap_8 FILLER_14_1957 ();
 sg13g2_fill_1 FILLER_14_1964 ();
 sg13g2_fill_2 FILLER_14_1969 ();
 sg13g2_fill_1 FILLER_14_1971 ();
 sg13g2_fill_2 FILLER_14_1980 ();
 sg13g2_fill_2 FILLER_14_2024 ();
 sg13g2_fill_2 FILLER_14_2057 ();
 sg13g2_fill_1 FILLER_14_2059 ();
 sg13g2_fill_2 FILLER_14_2078 ();
 sg13g2_fill_1 FILLER_14_2100 ();
 sg13g2_fill_2 FILLER_14_2119 ();
 sg13g2_decap_8 FILLER_14_2146 ();
 sg13g2_fill_2 FILLER_14_2153 ();
 sg13g2_fill_2 FILLER_14_2165 ();
 sg13g2_fill_2 FILLER_14_2184 ();
 sg13g2_decap_8 FILLER_14_2238 ();
 sg13g2_decap_8 FILLER_14_2245 ();
 sg13g2_decap_4 FILLER_14_2252 ();
 sg13g2_fill_2 FILLER_14_2256 ();
 sg13g2_decap_8 FILLER_14_2314 ();
 sg13g2_fill_1 FILLER_14_2347 ();
 sg13g2_fill_1 FILLER_14_2358 ();
 sg13g2_fill_1 FILLER_14_2401 ();
 sg13g2_fill_2 FILLER_14_2420 ();
 sg13g2_fill_1 FILLER_14_2451 ();
 sg13g2_fill_2 FILLER_14_2526 ();
 sg13g2_fill_1 FILLER_14_2528 ();
 sg13g2_fill_2 FILLER_14_2561 ();
 sg13g2_fill_1 FILLER_14_2563 ();
 sg13g2_fill_2 FILLER_14_2578 ();
 sg13g2_decap_8 FILLER_14_2584 ();
 sg13g2_decap_8 FILLER_14_2591 ();
 sg13g2_decap_8 FILLER_14_2598 ();
 sg13g2_decap_8 FILLER_14_2605 ();
 sg13g2_decap_8 FILLER_14_2612 ();
 sg13g2_decap_8 FILLER_14_2619 ();
 sg13g2_decap_8 FILLER_14_2626 ();
 sg13g2_decap_8 FILLER_14_2633 ();
 sg13g2_decap_8 FILLER_14_2640 ();
 sg13g2_decap_8 FILLER_14_2647 ();
 sg13g2_decap_8 FILLER_14_2654 ();
 sg13g2_decap_8 FILLER_14_2661 ();
 sg13g2_fill_2 FILLER_14_2668 ();
 sg13g2_decap_8 FILLER_15_0 ();
 sg13g2_decap_8 FILLER_15_7 ();
 sg13g2_decap_8 FILLER_15_14 ();
 sg13g2_decap_8 FILLER_15_21 ();
 sg13g2_decap_8 FILLER_15_28 ();
 sg13g2_decap_8 FILLER_15_35 ();
 sg13g2_decap_4 FILLER_15_42 ();
 sg13g2_fill_1 FILLER_15_46 ();
 sg13g2_fill_2 FILLER_15_96 ();
 sg13g2_fill_1 FILLER_15_98 ();
 sg13g2_decap_8 FILLER_15_103 ();
 sg13g2_decap_8 FILLER_15_144 ();
 sg13g2_decap_8 FILLER_15_151 ();
 sg13g2_decap_4 FILLER_15_158 ();
 sg13g2_fill_2 FILLER_15_202 ();
 sg13g2_decap_4 FILLER_15_276 ();
 sg13g2_fill_2 FILLER_15_280 ();
 sg13g2_fill_1 FILLER_15_300 ();
 sg13g2_decap_8 FILLER_15_317 ();
 sg13g2_decap_8 FILLER_15_324 ();
 sg13g2_decap_8 FILLER_15_331 ();
 sg13g2_decap_4 FILLER_15_338 ();
 sg13g2_decap_8 FILLER_15_360 ();
 sg13g2_decap_4 FILLER_15_372 ();
 sg13g2_fill_1 FILLER_15_464 ();
 sg13g2_fill_1 FILLER_15_483 ();
 sg13g2_fill_2 FILLER_15_488 ();
 sg13g2_fill_1 FILLER_15_494 ();
 sg13g2_fill_1 FILLER_15_503 ();
 sg13g2_fill_1 FILLER_15_511 ();
 sg13g2_fill_2 FILLER_15_517 ();
 sg13g2_fill_1 FILLER_15_528 ();
 sg13g2_fill_1 FILLER_15_551 ();
 sg13g2_fill_2 FILLER_15_642 ();
 sg13g2_fill_1 FILLER_15_662 ();
 sg13g2_fill_2 FILLER_15_672 ();
 sg13g2_fill_2 FILLER_15_680 ();
 sg13g2_fill_1 FILLER_15_682 ();
 sg13g2_fill_1 FILLER_15_693 ();
 sg13g2_fill_2 FILLER_15_699 ();
 sg13g2_fill_1 FILLER_15_701 ();
 sg13g2_fill_2 FILLER_15_706 ();
 sg13g2_fill_1 FILLER_15_708 ();
 sg13g2_fill_2 FILLER_15_713 ();
 sg13g2_decap_8 FILLER_15_725 ();
 sg13g2_decap_8 FILLER_15_732 ();
 sg13g2_fill_2 FILLER_15_739 ();
 sg13g2_fill_2 FILLER_15_777 ();
 sg13g2_fill_2 FILLER_15_784 ();
 sg13g2_fill_1 FILLER_15_786 ();
 sg13g2_decap_8 FILLER_15_823 ();
 sg13g2_decap_4 FILLER_15_830 ();
 sg13g2_fill_1 FILLER_15_834 ();
 sg13g2_decap_8 FILLER_15_839 ();
 sg13g2_decap_8 FILLER_15_846 ();
 sg13g2_decap_4 FILLER_15_853 ();
 sg13g2_decap_4 FILLER_15_893 ();
 sg13g2_fill_1 FILLER_15_897 ();
 sg13g2_decap_4 FILLER_15_901 ();
 sg13g2_fill_2 FILLER_15_915 ();
 sg13g2_fill_2 FILLER_15_927 ();
 sg13g2_fill_2 FILLER_15_955 ();
 sg13g2_decap_8 FILLER_15_961 ();
 sg13g2_fill_2 FILLER_15_1046 ();
 sg13g2_fill_1 FILLER_15_1048 ();
 sg13g2_fill_1 FILLER_15_1080 ();
 sg13g2_fill_2 FILLER_15_1107 ();
 sg13g2_fill_1 FILLER_15_1118 ();
 sg13g2_fill_2 FILLER_15_1140 ();
 sg13g2_decap_4 FILLER_15_1202 ();
 sg13g2_decap_8 FILLER_15_1257 ();
 sg13g2_fill_1 FILLER_15_1277 ();
 sg13g2_fill_2 FILLER_15_1317 ();
 sg13g2_fill_2 FILLER_15_1327 ();
 sg13g2_fill_1 FILLER_15_1329 ();
 sg13g2_fill_1 FILLER_15_1339 ();
 sg13g2_fill_1 FILLER_15_1365 ();
 sg13g2_decap_8 FILLER_15_1386 ();
 sg13g2_fill_2 FILLER_15_1393 ();
 sg13g2_fill_2 FILLER_15_1404 ();
 sg13g2_fill_1 FILLER_15_1406 ();
 sg13g2_decap_8 FILLER_15_1417 ();
 sg13g2_decap_4 FILLER_15_1424 ();
 sg13g2_decap_8 FILLER_15_1432 ();
 sg13g2_fill_2 FILLER_15_1439 ();
 sg13g2_fill_2 FILLER_15_1462 ();
 sg13g2_decap_8 FILLER_15_1473 ();
 sg13g2_decap_8 FILLER_15_1480 ();
 sg13g2_fill_1 FILLER_15_1487 ();
 sg13g2_decap_4 FILLER_15_1492 ();
 sg13g2_fill_1 FILLER_15_1496 ();
 sg13g2_decap_4 FILLER_15_1539 ();
 sg13g2_fill_1 FILLER_15_1543 ();
 sg13g2_decap_4 FILLER_15_1559 ();
 sg13g2_fill_1 FILLER_15_1563 ();
 sg13g2_fill_2 FILLER_15_1573 ();
 sg13g2_fill_1 FILLER_15_1624 ();
 sg13g2_fill_1 FILLER_15_1630 ();
 sg13g2_fill_1 FILLER_15_1637 ();
 sg13g2_fill_1 FILLER_15_1642 ();
 sg13g2_fill_1 FILLER_15_1669 ();
 sg13g2_fill_2 FILLER_15_1675 ();
 sg13g2_fill_2 FILLER_15_1686 ();
 sg13g2_fill_2 FILLER_15_1718 ();
 sg13g2_fill_1 FILLER_15_1720 ();
 sg13g2_decap_8 FILLER_15_1730 ();
 sg13g2_fill_2 FILLER_15_1737 ();
 sg13g2_fill_1 FILLER_15_1739 ();
 sg13g2_decap_4 FILLER_15_1750 ();
 sg13g2_fill_1 FILLER_15_1754 ();
 sg13g2_fill_2 FILLER_15_1785 ();
 sg13g2_decap_8 FILLER_15_1797 ();
 sg13g2_decap_8 FILLER_15_1817 ();
 sg13g2_decap_8 FILLER_15_1824 ();
 sg13g2_fill_1 FILLER_15_1831 ();
 sg13g2_fill_1 FILLER_15_1868 ();
 sg13g2_fill_1 FILLER_15_1948 ();
 sg13g2_fill_2 FILLER_15_2063 ();
 sg13g2_fill_1 FILLER_15_2065 ();
 sg13g2_fill_2 FILLER_15_2086 ();
 sg13g2_fill_1 FILLER_15_2107 ();
 sg13g2_fill_2 FILLER_15_2151 ();
 sg13g2_fill_1 FILLER_15_2153 ();
 sg13g2_decap_4 FILLER_15_2175 ();
 sg13g2_fill_1 FILLER_15_2179 ();
 sg13g2_fill_2 FILLER_15_2217 ();
 sg13g2_fill_1 FILLER_15_2219 ();
 sg13g2_fill_2 FILLER_15_2256 ();
 sg13g2_fill_2 FILLER_15_2262 ();
 sg13g2_fill_1 FILLER_15_2264 ();
 sg13g2_fill_2 FILLER_15_2273 ();
 sg13g2_fill_1 FILLER_15_2477 ();
 sg13g2_fill_1 FILLER_15_2510 ();
 sg13g2_decap_8 FILLER_15_2522 ();
 sg13g2_decap_8 FILLER_15_2529 ();
 sg13g2_decap_8 FILLER_15_2550 ();
 sg13g2_fill_2 FILLER_15_2557 ();
 sg13g2_fill_1 FILLER_15_2559 ();
 sg13g2_fill_1 FILLER_15_2573 ();
 sg13g2_decap_4 FILLER_15_2600 ();
 sg13g2_decap_8 FILLER_15_2608 ();
 sg13g2_decap_8 FILLER_15_2615 ();
 sg13g2_decap_8 FILLER_15_2622 ();
 sg13g2_decap_8 FILLER_15_2629 ();
 sg13g2_decap_8 FILLER_15_2636 ();
 sg13g2_decap_8 FILLER_15_2643 ();
 sg13g2_decap_8 FILLER_15_2650 ();
 sg13g2_decap_8 FILLER_15_2657 ();
 sg13g2_decap_4 FILLER_15_2664 ();
 sg13g2_fill_2 FILLER_15_2668 ();
 sg13g2_decap_8 FILLER_16_0 ();
 sg13g2_decap_8 FILLER_16_7 ();
 sg13g2_decap_8 FILLER_16_14 ();
 sg13g2_decap_8 FILLER_16_21 ();
 sg13g2_decap_8 FILLER_16_28 ();
 sg13g2_decap_8 FILLER_16_35 ();
 sg13g2_decap_8 FILLER_16_42 ();
 sg13g2_decap_8 FILLER_16_49 ();
 sg13g2_fill_2 FILLER_16_56 ();
 sg13g2_fill_1 FILLER_16_58 ();
 sg13g2_fill_2 FILLER_16_69 ();
 sg13g2_fill_2 FILLER_16_108 ();
 sg13g2_fill_1 FILLER_16_110 ();
 sg13g2_fill_2 FILLER_16_116 ();
 sg13g2_fill_1 FILLER_16_118 ();
 sg13g2_decap_8 FILLER_16_155 ();
 sg13g2_decap_4 FILLER_16_162 ();
 sg13g2_fill_1 FILLER_16_166 ();
 sg13g2_fill_1 FILLER_16_181 ();
 sg13g2_fill_1 FILLER_16_186 ();
 sg13g2_fill_1 FILLER_16_213 ();
 sg13g2_decap_4 FILLER_16_265 ();
 sg13g2_fill_2 FILLER_16_282 ();
 sg13g2_decap_4 FILLER_16_290 ();
 sg13g2_fill_1 FILLER_16_294 ();
 sg13g2_decap_4 FILLER_16_334 ();
 sg13g2_decap_8 FILLER_16_365 ();
 sg13g2_decap_8 FILLER_16_372 ();
 sg13g2_decap_4 FILLER_16_383 ();
 sg13g2_fill_1 FILLER_16_419 ();
 sg13g2_fill_1 FILLER_16_435 ();
 sg13g2_fill_1 FILLER_16_446 ();
 sg13g2_fill_1 FILLER_16_452 ();
 sg13g2_fill_1 FILLER_16_458 ();
 sg13g2_decap_8 FILLER_16_489 ();
 sg13g2_fill_2 FILLER_16_496 ();
 sg13g2_fill_1 FILLER_16_585 ();
 sg13g2_fill_1 FILLER_16_612 ();
 sg13g2_fill_1 FILLER_16_618 ();
 sg13g2_fill_2 FILLER_16_629 ();
 sg13g2_fill_2 FILLER_16_635 ();
 sg13g2_fill_1 FILLER_16_641 ();
 sg13g2_fill_1 FILLER_16_647 ();
 sg13g2_fill_1 FILLER_16_686 ();
 sg13g2_fill_2 FILLER_16_692 ();
 sg13g2_fill_1 FILLER_16_698 ();
 sg13g2_fill_2 FILLER_16_703 ();
 sg13g2_fill_2 FILLER_16_719 ();
 sg13g2_decap_4 FILLER_16_726 ();
 sg13g2_fill_2 FILLER_16_734 ();
 sg13g2_fill_1 FILLER_16_736 ();
 sg13g2_decap_8 FILLER_16_742 ();
 sg13g2_fill_1 FILLER_16_793 ();
 sg13g2_fill_2 FILLER_16_804 ();
 sg13g2_fill_2 FILLER_16_832 ();
 sg13g2_fill_1 FILLER_16_834 ();
 sg13g2_fill_2 FILLER_16_839 ();
 sg13g2_fill_1 FILLER_16_841 ();
 sg13g2_decap_8 FILLER_16_868 ();
 sg13g2_decap_4 FILLER_16_883 ();
 sg13g2_fill_1 FILLER_16_887 ();
 sg13g2_fill_2 FILLER_16_906 ();
 sg13g2_fill_1 FILLER_16_933 ();
 sg13g2_decap_4 FILLER_16_960 ();
 sg13g2_decap_8 FILLER_16_968 ();
 sg13g2_fill_1 FILLER_16_975 ();
 sg13g2_fill_2 FILLER_16_1014 ();
 sg13g2_fill_1 FILLER_16_1016 ();
 sg13g2_fill_1 FILLER_16_1069 ();
 sg13g2_decap_4 FILLER_16_1074 ();
 sg13g2_fill_1 FILLER_16_1078 ();
 sg13g2_decap_8 FILLER_16_1137 ();
 sg13g2_decap_8 FILLER_16_1144 ();
 sg13g2_fill_1 FILLER_16_1169 ();
 sg13g2_fill_1 FILLER_16_1175 ();
 sg13g2_fill_1 FILLER_16_1206 ();
 sg13g2_fill_2 FILLER_16_1212 ();
 sg13g2_fill_2 FILLER_16_1223 ();
 sg13g2_decap_8 FILLER_16_1251 ();
 sg13g2_fill_1 FILLER_16_1258 ();
 sg13g2_fill_2 FILLER_16_1264 ();
 sg13g2_fill_2 FILLER_16_1292 ();
 sg13g2_decap_4 FILLER_16_1315 ();
 sg13g2_fill_2 FILLER_16_1319 ();
 sg13g2_fill_2 FILLER_16_1334 ();
 sg13g2_fill_1 FILLER_16_1336 ();
 sg13g2_decap_4 FILLER_16_1346 ();
 sg13g2_decap_8 FILLER_16_1354 ();
 sg13g2_decap_8 FILLER_16_1361 ();
 sg13g2_decap_8 FILLER_16_1368 ();
 sg13g2_decap_8 FILLER_16_1375 ();
 sg13g2_decap_8 FILLER_16_1382 ();
 sg13g2_fill_1 FILLER_16_1389 ();
 sg13g2_fill_2 FILLER_16_1431 ();
 sg13g2_fill_2 FILLER_16_1437 ();
 sg13g2_fill_2 FILLER_16_1443 ();
 sg13g2_fill_2 FILLER_16_1457 ();
 sg13g2_fill_1 FILLER_16_1459 ();
 sg13g2_decap_8 FILLER_16_1470 ();
 sg13g2_decap_8 FILLER_16_1477 ();
 sg13g2_decap_4 FILLER_16_1484 ();
 sg13g2_fill_1 FILLER_16_1493 ();
 sg13g2_fill_1 FILLER_16_1520 ();
 sg13g2_fill_1 FILLER_16_1525 ();
 sg13g2_decap_4 FILLER_16_1553 ();
 sg13g2_fill_2 FILLER_16_1557 ();
 sg13g2_fill_1 FILLER_16_1585 ();
 sg13g2_fill_2 FILLER_16_1600 ();
 sg13g2_fill_2 FILLER_16_1606 ();
 sg13g2_fill_2 FILLER_16_1611 ();
 sg13g2_decap_8 FILLER_16_1696 ();
 sg13g2_fill_2 FILLER_16_1703 ();
 sg13g2_fill_2 FILLER_16_1723 ();
 sg13g2_fill_1 FILLER_16_1730 ();
 sg13g2_fill_2 FILLER_16_1766 ();
 sg13g2_fill_1 FILLER_16_1768 ();
 sg13g2_decap_8 FILLER_16_1803 ();
 sg13g2_decap_8 FILLER_16_1810 ();
 sg13g2_decap_4 FILLER_16_1817 ();
 sg13g2_fill_1 FILLER_16_1821 ();
 sg13g2_fill_2 FILLER_16_1858 ();
 sg13g2_decap_4 FILLER_16_1891 ();
 sg13g2_fill_2 FILLER_16_1899 ();
 sg13g2_fill_1 FILLER_16_1901 ();
 sg13g2_fill_2 FILLER_16_1932 ();
 sg13g2_fill_1 FILLER_16_1934 ();
 sg13g2_fill_1 FILLER_16_1960 ();
 sg13g2_decap_8 FILLER_16_1987 ();
 sg13g2_fill_1 FILLER_16_2056 ();
 sg13g2_fill_2 FILLER_16_2061 ();
 sg13g2_decap_4 FILLER_16_2067 ();
 sg13g2_fill_2 FILLER_16_2071 ();
 sg13g2_fill_1 FILLER_16_2125 ();
 sg13g2_fill_1 FILLER_16_2158 ();
 sg13g2_fill_1 FILLER_16_2185 ();
 sg13g2_fill_1 FILLER_16_2226 ();
 sg13g2_decap_8 FILLER_16_2253 ();
 sg13g2_decap_4 FILLER_16_2260 ();
 sg13g2_fill_1 FILLER_16_2264 ();
 sg13g2_fill_2 FILLER_16_2285 ();
 sg13g2_fill_1 FILLER_16_2307 ();
 sg13g2_fill_1 FILLER_16_2312 ();
 sg13g2_fill_1 FILLER_16_2322 ();
 sg13g2_fill_1 FILLER_16_2417 ();
 sg13g2_fill_2 FILLER_16_2425 ();
 sg13g2_fill_1 FILLER_16_2437 ();
 sg13g2_fill_1 FILLER_16_2444 ();
 sg13g2_fill_1 FILLER_16_2451 ();
 sg13g2_fill_1 FILLER_16_2458 ();
 sg13g2_fill_2 FILLER_16_2478 ();
 sg13g2_fill_1 FILLER_16_2480 ();
 sg13g2_fill_2 FILLER_16_2485 ();
 sg13g2_fill_1 FILLER_16_2487 ();
 sg13g2_fill_1 FILLER_16_2542 ();
 sg13g2_decap_8 FILLER_16_2651 ();
 sg13g2_decap_8 FILLER_16_2658 ();
 sg13g2_decap_4 FILLER_16_2665 ();
 sg13g2_fill_1 FILLER_16_2669 ();
 sg13g2_decap_8 FILLER_17_0 ();
 sg13g2_decap_8 FILLER_17_7 ();
 sg13g2_decap_8 FILLER_17_14 ();
 sg13g2_decap_4 FILLER_17_21 ();
 sg13g2_fill_2 FILLER_17_25 ();
 sg13g2_decap_8 FILLER_17_53 ();
 sg13g2_fill_2 FILLER_17_60 ();
 sg13g2_fill_1 FILLER_17_62 ();
 sg13g2_decap_4 FILLER_17_125 ();
 sg13g2_fill_2 FILLER_17_129 ();
 sg13g2_fill_1 FILLER_17_141 ();
 sg13g2_decap_8 FILLER_17_152 ();
 sg13g2_decap_8 FILLER_17_159 ();
 sg13g2_decap_8 FILLER_17_166 ();
 sg13g2_decap_8 FILLER_17_177 ();
 sg13g2_decap_8 FILLER_17_184 ();
 sg13g2_fill_2 FILLER_17_191 ();
 sg13g2_fill_2 FILLER_17_203 ();
 sg13g2_fill_1 FILLER_17_205 ();
 sg13g2_decap_4 FILLER_17_220 ();
 sg13g2_decap_8 FILLER_17_238 ();
 sg13g2_fill_2 FILLER_17_245 ();
 sg13g2_fill_1 FILLER_17_253 ();
 sg13g2_fill_1 FILLER_17_262 ();
 sg13g2_fill_1 FILLER_17_271 ();
 sg13g2_fill_2 FILLER_17_289 ();
 sg13g2_decap_8 FILLER_17_294 ();
 sg13g2_decap_4 FILLER_17_301 ();
 sg13g2_fill_2 FILLER_17_309 ();
 sg13g2_decap_4 FILLER_17_320 ();
 sg13g2_fill_2 FILLER_17_324 ();
 sg13g2_decap_4 FILLER_17_331 ();
 sg13g2_fill_2 FILLER_17_370 ();
 sg13g2_fill_2 FILLER_17_412 ();
 sg13g2_fill_1 FILLER_17_414 ();
 sg13g2_fill_1 FILLER_17_459 ();
 sg13g2_fill_1 FILLER_17_464 ();
 sg13g2_fill_2 FILLER_17_478 ();
 sg13g2_fill_1 FILLER_17_485 ();
 sg13g2_decap_4 FILLER_17_498 ();
 sg13g2_fill_1 FILLER_17_502 ();
 sg13g2_fill_2 FILLER_17_507 ();
 sg13g2_fill_1 FILLER_17_509 ();
 sg13g2_decap_4 FILLER_17_515 ();
 sg13g2_fill_2 FILLER_17_523 ();
 sg13g2_decap_4 FILLER_17_534 ();
 sg13g2_fill_1 FILLER_17_538 ();
 sg13g2_fill_2 FILLER_17_544 ();
 sg13g2_fill_1 FILLER_17_550 ();
 sg13g2_fill_2 FILLER_17_555 ();
 sg13g2_fill_1 FILLER_17_572 ();
 sg13g2_decap_8 FILLER_17_581 ();
 sg13g2_decap_4 FILLER_17_588 ();
 sg13g2_fill_2 FILLER_17_592 ();
 sg13g2_fill_1 FILLER_17_606 ();
 sg13g2_decap_4 FILLER_17_622 ();
 sg13g2_fill_2 FILLER_17_762 ();
 sg13g2_fill_2 FILLER_17_768 ();
 sg13g2_decap_8 FILLER_17_774 ();
 sg13g2_decap_4 FILLER_17_781 ();
 sg13g2_fill_1 FILLER_17_785 ();
 sg13g2_decap_8 FILLER_17_813 ();
 sg13g2_fill_2 FILLER_17_820 ();
 sg13g2_decap_8 FILLER_17_826 ();
 sg13g2_decap_8 FILLER_17_833 ();
 sg13g2_decap_8 FILLER_17_840 ();
 sg13g2_decap_8 FILLER_17_847 ();
 sg13g2_decap_4 FILLER_17_854 ();
 sg13g2_fill_1 FILLER_17_858 ();
 sg13g2_fill_2 FILLER_17_928 ();
 sg13g2_fill_1 FILLER_17_940 ();
 sg13g2_decap_8 FILLER_17_975 ();
 sg13g2_fill_2 FILLER_17_982 ();
 sg13g2_fill_1 FILLER_17_1001 ();
 sg13g2_fill_2 FILLER_17_1027 ();
 sg13g2_fill_2 FILLER_17_1033 ();
 sg13g2_fill_1 FILLER_17_1035 ();
 sg13g2_fill_1 FILLER_17_1041 ();
 sg13g2_fill_1 FILLER_17_1046 ();
 sg13g2_fill_1 FILLER_17_1052 ();
 sg13g2_fill_1 FILLER_17_1057 ();
 sg13g2_decap_8 FILLER_17_1062 ();
 sg13g2_decap_4 FILLER_17_1069 ();
 sg13g2_fill_1 FILLER_17_1073 ();
 sg13g2_decap_8 FILLER_17_1078 ();
 sg13g2_fill_1 FILLER_17_1090 ();
 sg13g2_fill_2 FILLER_17_1096 ();
 sg13g2_decap_8 FILLER_17_1128 ();
 sg13g2_decap_8 FILLER_17_1135 ();
 sg13g2_fill_1 FILLER_17_1142 ();
 sg13g2_decap_8 FILLER_17_1151 ();
 sg13g2_decap_8 FILLER_17_1158 ();
 sg13g2_decap_8 FILLER_17_1165 ();
 sg13g2_decap_4 FILLER_17_1172 ();
 sg13g2_fill_2 FILLER_17_1176 ();
 sg13g2_fill_1 FILLER_17_1187 ();
 sg13g2_decap_8 FILLER_17_1192 ();
 sg13g2_decap_8 FILLER_17_1199 ();
 sg13g2_fill_2 FILLER_17_1206 ();
 sg13g2_decap_8 FILLER_17_1247 ();
 sg13g2_decap_8 FILLER_17_1254 ();
 sg13g2_fill_2 FILLER_17_1261 ();
 sg13g2_fill_1 FILLER_17_1263 ();
 sg13g2_fill_1 FILLER_17_1290 ();
 sg13g2_decap_8 FILLER_17_1312 ();
 sg13g2_fill_1 FILLER_17_1319 ();
 sg13g2_fill_2 FILLER_17_1330 ();
 sg13g2_decap_4 FILLER_17_1336 ();
 sg13g2_fill_1 FILLER_17_1340 ();
 sg13g2_decap_8 FILLER_17_1345 ();
 sg13g2_decap_8 FILLER_17_1352 ();
 sg13g2_decap_8 FILLER_17_1359 ();
 sg13g2_fill_2 FILLER_17_1366 ();
 sg13g2_fill_1 FILLER_17_1383 ();
 sg13g2_fill_2 FILLER_17_1388 ();
 sg13g2_fill_2 FILLER_17_1435 ();
 sg13g2_fill_1 FILLER_17_1437 ();
 sg13g2_fill_1 FILLER_17_1443 ();
 sg13g2_fill_2 FILLER_17_1448 ();
 sg13g2_fill_1 FILLER_17_1450 ();
 sg13g2_fill_1 FILLER_17_1487 ();
 sg13g2_fill_1 FILLER_17_1506 ();
 sg13g2_fill_1 FILLER_17_1537 ();
 sg13g2_decap_4 FILLER_17_1543 ();
 sg13g2_fill_2 FILLER_17_1547 ();
 sg13g2_fill_2 FILLER_17_1554 ();
 sg13g2_fill_1 FILLER_17_1556 ();
 sg13g2_fill_2 FILLER_17_1562 ();
 sg13g2_fill_1 FILLER_17_1615 ();
 sg13g2_fill_1 FILLER_17_1685 ();
 sg13g2_fill_2 FILLER_17_1716 ();
 sg13g2_decap_4 FILLER_17_1757 ();
 sg13g2_fill_1 FILLER_17_1761 ();
 sg13g2_decap_4 FILLER_17_1766 ();
 sg13g2_fill_2 FILLER_17_1774 ();
 sg13g2_decap_4 FILLER_17_1822 ();
 sg13g2_decap_8 FILLER_17_1830 ();
 sg13g2_decap_4 FILLER_17_1837 ();
 sg13g2_fill_2 FILLER_17_1845 ();
 sg13g2_fill_1 FILLER_17_1847 ();
 sg13g2_fill_1 FILLER_17_1852 ();
 sg13g2_decap_8 FILLER_17_1857 ();
 sg13g2_decap_8 FILLER_17_1864 ();
 sg13g2_decap_8 FILLER_17_1871 ();
 sg13g2_decap_8 FILLER_17_1878 ();
 sg13g2_decap_4 FILLER_17_1885 ();
 sg13g2_fill_2 FILLER_17_1939 ();
 sg13g2_fill_1 FILLER_17_1950 ();
 sg13g2_decap_8 FILLER_17_1974 ();
 sg13g2_fill_1 FILLER_17_1981 ();
 sg13g2_fill_1 FILLER_17_1990 ();
 sg13g2_decap_8 FILLER_17_1995 ();
 sg13g2_decap_4 FILLER_17_2002 ();
 sg13g2_decap_4 FILLER_17_2020 ();
 sg13g2_fill_2 FILLER_17_2024 ();
 sg13g2_decap_8 FILLER_17_2039 ();
 sg13g2_fill_1 FILLER_17_2046 ();
 sg13g2_decap_8 FILLER_17_2087 ();
 sg13g2_fill_2 FILLER_17_2094 ();
 sg13g2_fill_1 FILLER_17_2096 ();
 sg13g2_fill_2 FILLER_17_2100 ();
 sg13g2_fill_1 FILLER_17_2105 ();
 sg13g2_fill_1 FILLER_17_2110 ();
 sg13g2_fill_2 FILLER_17_2121 ();
 sg13g2_fill_2 FILLER_17_2127 ();
 sg13g2_fill_2 FILLER_17_2139 ();
 sg13g2_fill_2 FILLER_17_2190 ();
 sg13g2_fill_2 FILLER_17_2204 ();
 sg13g2_fill_1 FILLER_17_2206 ();
 sg13g2_decap_8 FILLER_17_2264 ();
 sg13g2_decap_8 FILLER_17_2271 ();
 sg13g2_decap_4 FILLER_17_2278 ();
 sg13g2_decap_4 FILLER_17_2309 ();
 sg13g2_decap_8 FILLER_17_2318 ();
 sg13g2_decap_4 FILLER_17_2325 ();
 sg13g2_fill_2 FILLER_17_2329 ();
 sg13g2_fill_1 FILLER_17_2370 ();
 sg13g2_fill_1 FILLER_17_2382 ();
 sg13g2_fill_2 FILLER_17_2393 ();
 sg13g2_decap_8 FILLER_17_2526 ();
 sg13g2_decap_4 FILLER_17_2533 ();
 sg13g2_fill_2 FILLER_17_2537 ();
 sg13g2_fill_2 FILLER_17_2560 ();
 sg13g2_decap_8 FILLER_17_2566 ();
 sg13g2_decap_4 FILLER_17_2573 ();
 sg13g2_fill_1 FILLER_17_2577 ();
 sg13g2_decap_4 FILLER_17_2582 ();
 sg13g2_fill_1 FILLER_17_2586 ();
 sg13g2_fill_1 FILLER_17_2597 ();
 sg13g2_decap_4 FILLER_17_2608 ();
 sg13g2_fill_2 FILLER_17_2612 ();
 sg13g2_decap_8 FILLER_17_2640 ();
 sg13g2_decap_8 FILLER_17_2647 ();
 sg13g2_decap_8 FILLER_17_2654 ();
 sg13g2_decap_8 FILLER_17_2661 ();
 sg13g2_fill_2 FILLER_17_2668 ();
 sg13g2_decap_8 FILLER_18_0 ();
 sg13g2_decap_8 FILLER_18_7 ();
 sg13g2_decap_4 FILLER_18_14 ();
 sg13g2_fill_1 FILLER_18_18 ();
 sg13g2_fill_1 FILLER_18_52 ();
 sg13g2_decap_8 FILLER_18_56 ();
 sg13g2_decap_8 FILLER_18_63 ();
 sg13g2_fill_1 FILLER_18_70 ();
 sg13g2_fill_2 FILLER_18_89 ();
 sg13g2_decap_4 FILLER_18_95 ();
 sg13g2_decap_4 FILLER_18_103 ();
 sg13g2_fill_2 FILLER_18_111 ();
 sg13g2_fill_1 FILLER_18_113 ();
 sg13g2_fill_2 FILLER_18_124 ();
 sg13g2_fill_1 FILLER_18_126 ();
 sg13g2_decap_4 FILLER_18_130 ();
 sg13g2_fill_1 FILLER_18_134 ();
 sg13g2_fill_2 FILLER_18_142 ();
 sg13g2_fill_2 FILLER_18_148 ();
 sg13g2_fill_1 FILLER_18_150 ();
 sg13g2_decap_4 FILLER_18_177 ();
 sg13g2_fill_1 FILLER_18_181 ();
 sg13g2_fill_2 FILLER_18_203 ();
 sg13g2_fill_1 FILLER_18_205 ();
 sg13g2_fill_1 FILLER_18_211 ();
 sg13g2_fill_2 FILLER_18_224 ();
 sg13g2_decap_8 FILLER_18_236 ();
 sg13g2_fill_1 FILLER_18_243 ();
 sg13g2_fill_2 FILLER_18_269 ();
 sg13g2_fill_2 FILLER_18_301 ();
 sg13g2_fill_2 FILLER_18_333 ();
 sg13g2_fill_2 FILLER_18_366 ();
 sg13g2_fill_1 FILLER_18_368 ();
 sg13g2_fill_1 FILLER_18_439 ();
 sg13g2_decap_8 FILLER_18_444 ();
 sg13g2_decap_4 FILLER_18_451 ();
 sg13g2_fill_1 FILLER_18_460 ();
 sg13g2_decap_8 FILLER_18_468 ();
 sg13g2_fill_2 FILLER_18_475 ();
 sg13g2_decap_4 FILLER_18_481 ();
 sg13g2_decap_4 FILLER_18_490 ();
 sg13g2_fill_1 FILLER_18_494 ();
 sg13g2_decap_8 FILLER_18_499 ();
 sg13g2_decap_4 FILLER_18_506 ();
 sg13g2_fill_1 FILLER_18_514 ();
 sg13g2_fill_2 FILLER_18_519 ();
 sg13g2_fill_1 FILLER_18_531 ();
 sg13g2_decap_8 FILLER_18_540 ();
 sg13g2_fill_2 FILLER_18_547 ();
 sg13g2_fill_1 FILLER_18_568 ();
 sg13g2_decap_4 FILLER_18_575 ();
 sg13g2_decap_8 FILLER_18_583 ();
 sg13g2_fill_1 FILLER_18_607 ();
 sg13g2_fill_2 FILLER_18_612 ();
 sg13g2_decap_8 FILLER_18_618 ();
 sg13g2_fill_2 FILLER_18_629 ();
 sg13g2_fill_2 FILLER_18_671 ();
 sg13g2_fill_1 FILLER_18_686 ();
 sg13g2_fill_2 FILLER_18_692 ();
 sg13g2_decap_4 FILLER_18_731 ();
 sg13g2_fill_2 FILLER_18_735 ();
 sg13g2_decap_4 FILLER_18_742 ();
 sg13g2_fill_2 FILLER_18_746 ();
 sg13g2_decap_4 FILLER_18_762 ();
 sg13g2_fill_1 FILLER_18_766 ();
 sg13g2_decap_8 FILLER_18_772 ();
 sg13g2_decap_4 FILLER_18_779 ();
 sg13g2_fill_2 FILLER_18_792 ();
 sg13g2_decap_8 FILLER_18_809 ();
 sg13g2_fill_2 FILLER_18_816 ();
 sg13g2_decap_4 FILLER_18_844 ();
 sg13g2_fill_1 FILLER_18_848 ();
 sg13g2_decap_4 FILLER_18_863 ();
 sg13g2_fill_2 FILLER_18_867 ();
 sg13g2_decap_4 FILLER_18_904 ();
 sg13g2_fill_1 FILLER_18_908 ();
 sg13g2_decap_4 FILLER_18_913 ();
 sg13g2_decap_8 FILLER_18_979 ();
 sg13g2_decap_8 FILLER_18_986 ();
 sg13g2_decap_4 FILLER_18_993 ();
 sg13g2_fill_2 FILLER_18_997 ();
 sg13g2_decap_8 FILLER_18_1003 ();
 sg13g2_decap_4 FILLER_18_1010 ();
 sg13g2_fill_1 FILLER_18_1014 ();
 sg13g2_decap_8 FILLER_18_1019 ();
 sg13g2_decap_8 FILLER_18_1026 ();
 sg13g2_decap_8 FILLER_18_1033 ();
 sg13g2_decap_8 FILLER_18_1040 ();
 sg13g2_fill_2 FILLER_18_1047 ();
 sg13g2_fill_2 FILLER_18_1075 ();
 sg13g2_fill_1 FILLER_18_1077 ();
 sg13g2_decap_8 FILLER_18_1091 ();
 sg13g2_decap_4 FILLER_18_1098 ();
 sg13g2_fill_2 FILLER_18_1102 ();
 sg13g2_fill_2 FILLER_18_1113 ();
 sg13g2_decap_8 FILLER_18_1119 ();
 sg13g2_fill_2 FILLER_18_1126 ();
 sg13g2_fill_1 FILLER_18_1128 ();
 sg13g2_decap_8 FILLER_18_1168 ();
 sg13g2_decap_8 FILLER_18_1175 ();
 sg13g2_fill_2 FILLER_18_1182 ();
 sg13g2_fill_1 FILLER_18_1184 ();
 sg13g2_decap_4 FILLER_18_1202 ();
 sg13g2_fill_2 FILLER_18_1206 ();
 sg13g2_decap_8 FILLER_18_1212 ();
 sg13g2_fill_2 FILLER_18_1219 ();
 sg13g2_fill_1 FILLER_18_1221 ();
 sg13g2_decap_4 FILLER_18_1230 ();
 sg13g2_decap_8 FILLER_18_1238 ();
 sg13g2_decap_8 FILLER_18_1245 ();
 sg13g2_decap_8 FILLER_18_1252 ();
 sg13g2_decap_8 FILLER_18_1272 ();
 sg13g2_decap_8 FILLER_18_1279 ();
 sg13g2_decap_8 FILLER_18_1286 ();
 sg13g2_fill_1 FILLER_18_1323 ();
 sg13g2_fill_2 FILLER_18_1328 ();
 sg13g2_decap_8 FILLER_18_1356 ();
 sg13g2_fill_2 FILLER_18_1363 ();
 sg13g2_fill_2 FILLER_18_1434 ();
 sg13g2_fill_1 FILLER_18_1436 ();
 sg13g2_fill_1 FILLER_18_1443 ();
 sg13g2_fill_1 FILLER_18_1448 ();
 sg13g2_fill_1 FILLER_18_1454 ();
 sg13g2_fill_2 FILLER_18_1461 ();
 sg13g2_fill_1 FILLER_18_1467 ();
 sg13g2_decap_8 FILLER_18_1472 ();
 sg13g2_fill_2 FILLER_18_1479 ();
 sg13g2_fill_1 FILLER_18_1481 ();
 sg13g2_fill_2 FILLER_18_1491 ();
 sg13g2_fill_2 FILLER_18_1496 ();
 sg13g2_fill_1 FILLER_18_1498 ();
 sg13g2_fill_2 FILLER_18_1502 ();
 sg13g2_fill_2 FILLER_18_1513 ();
 sg13g2_fill_2 FILLER_18_1575 ();
 sg13g2_fill_1 FILLER_18_1582 ();
 sg13g2_fill_1 FILLER_18_1589 ();
 sg13g2_fill_1 FILLER_18_1610 ();
 sg13g2_fill_1 FILLER_18_1626 ();
 sg13g2_fill_2 FILLER_18_1660 ();
 sg13g2_fill_2 FILLER_18_1693 ();
 sg13g2_decap_8 FILLER_18_1702 ();
 sg13g2_fill_2 FILLER_18_1709 ();
 sg13g2_fill_1 FILLER_18_1711 ();
 sg13g2_fill_2 FILLER_18_1720 ();
 sg13g2_decap_4 FILLER_18_1745 ();
 sg13g2_decap_8 FILLER_18_1762 ();
 sg13g2_decap_8 FILLER_18_1769 ();
 sg13g2_fill_2 FILLER_18_1776 ();
 sg13g2_fill_1 FILLER_18_1778 ();
 sg13g2_fill_2 FILLER_18_1815 ();
 sg13g2_fill_1 FILLER_18_1817 ();
 sg13g2_decap_4 FILLER_18_1844 ();
 sg13g2_fill_2 FILLER_18_1848 ();
 sg13g2_fill_2 FILLER_18_1854 ();
 sg13g2_decap_8 FILLER_18_1893 ();
 sg13g2_decap_8 FILLER_18_1900 ();
 sg13g2_fill_1 FILLER_18_1907 ();
 sg13g2_fill_1 FILLER_18_1912 ();
 sg13g2_decap_8 FILLER_18_1917 ();
 sg13g2_decap_8 FILLER_18_1924 ();
 sg13g2_decap_8 FILLER_18_1931 ();
 sg13g2_fill_2 FILLER_18_1938 ();
 sg13g2_fill_1 FILLER_18_1940 ();
 sg13g2_fill_2 FILLER_18_1970 ();
 sg13g2_fill_1 FILLER_18_1976 ();
 sg13g2_fill_2 FILLER_18_2010 ();
 sg13g2_decap_4 FILLER_18_2038 ();
 sg13g2_fill_2 FILLER_18_2073 ();
 sg13g2_fill_1 FILLER_18_2075 ();
 sg13g2_decap_8 FILLER_18_2084 ();
 sg13g2_decap_8 FILLER_18_2091 ();
 sg13g2_decap_8 FILLER_18_2098 ();
 sg13g2_decap_8 FILLER_18_2105 ();
 sg13g2_decap_4 FILLER_18_2112 ();
 sg13g2_fill_1 FILLER_18_2116 ();
 sg13g2_fill_2 FILLER_18_2143 ();
 sg13g2_fill_1 FILLER_18_2145 ();
 sg13g2_fill_2 FILLER_18_2184 ();
 sg13g2_fill_1 FILLER_18_2186 ();
 sg13g2_decap_4 FILLER_18_2233 ();
 sg13g2_decap_8 FILLER_18_2241 ();
 sg13g2_fill_2 FILLER_18_2258 ();
 sg13g2_fill_1 FILLER_18_2260 ();
 sg13g2_fill_1 FILLER_18_2291 ();
 sg13g2_fill_1 FILLER_18_2314 ();
 sg13g2_fill_1 FILLER_18_2323 ();
 sg13g2_decap_4 FILLER_18_2334 ();
 sg13g2_fill_1 FILLER_18_2414 ();
 sg13g2_decap_4 FILLER_18_2457 ();
 sg13g2_fill_1 FILLER_18_2461 ();
 sg13g2_fill_2 FILLER_18_2466 ();
 sg13g2_fill_2 FILLER_18_2511 ();
 sg13g2_fill_1 FILLER_18_2513 ();
 sg13g2_fill_1 FILLER_18_2518 ();
 sg13g2_fill_1 FILLER_18_2529 ();
 sg13g2_decap_8 FILLER_18_2566 ();
 sg13g2_decap_8 FILLER_18_2573 ();
 sg13g2_decap_8 FILLER_18_2580 ();
 sg13g2_decap_8 FILLER_18_2587 ();
 sg13g2_decap_4 FILLER_18_2594 ();
 sg13g2_fill_2 FILLER_18_2635 ();
 sg13g2_decap_8 FILLER_18_2663 ();
 sg13g2_fill_2 FILLER_19_0 ();
 sg13g2_fill_2 FILLER_19_31 ();
 sg13g2_fill_1 FILLER_19_37 ();
 sg13g2_fill_1 FILLER_19_58 ();
 sg13g2_fill_1 FILLER_19_64 ();
 sg13g2_decap_8 FILLER_19_68 ();
 sg13g2_decap_4 FILLER_19_75 ();
 sg13g2_fill_1 FILLER_19_105 ();
 sg13g2_fill_1 FILLER_19_132 ();
 sg13g2_fill_1 FILLER_19_159 ();
 sg13g2_fill_2 FILLER_19_186 ();
 sg13g2_fill_1 FILLER_19_214 ();
 sg13g2_decap_8 FILLER_19_247 ();
 sg13g2_fill_2 FILLER_19_254 ();
 sg13g2_fill_1 FILLER_19_256 ();
 sg13g2_decap_4 FILLER_19_262 ();
 sg13g2_fill_1 FILLER_19_266 ();
 sg13g2_decap_8 FILLER_19_285 ();
 sg13g2_decap_4 FILLER_19_292 ();
 sg13g2_fill_2 FILLER_19_296 ();
 sg13g2_decap_4 FILLER_19_310 ();
 sg13g2_decap_8 FILLER_19_318 ();
 sg13g2_decap_4 FILLER_19_325 ();
 sg13g2_fill_2 FILLER_19_345 ();
 sg13g2_fill_1 FILLER_19_351 ();
 sg13g2_decap_8 FILLER_19_356 ();
 sg13g2_decap_8 FILLER_19_363 ();
 sg13g2_decap_8 FILLER_19_370 ();
 sg13g2_decap_8 FILLER_19_377 ();
 sg13g2_fill_1 FILLER_19_384 ();
 sg13g2_fill_1 FILLER_19_390 ();
 sg13g2_decap_4 FILLER_19_430 ();
 sg13g2_decap_4 FILLER_19_478 ();
 sg13g2_fill_1 FILLER_19_482 ();
 sg13g2_fill_1 FILLER_19_496 ();
 sg13g2_decap_4 FILLER_19_503 ();
 sg13g2_fill_2 FILLER_19_511 ();
 sg13g2_decap_4 FILLER_19_517 ();
 sg13g2_decap_4 FILLER_19_526 ();
 sg13g2_decap_8 FILLER_19_535 ();
 sg13g2_decap_4 FILLER_19_582 ();
 sg13g2_fill_2 FILLER_19_586 ();
 sg13g2_decap_4 FILLER_19_594 ();
 sg13g2_fill_1 FILLER_19_613 ();
 sg13g2_fill_2 FILLER_19_619 ();
 sg13g2_fill_2 FILLER_19_626 ();
 sg13g2_fill_1 FILLER_19_633 ();
 sg13g2_fill_1 FILLER_19_638 ();
 sg13g2_fill_2 FILLER_19_667 ();
 sg13g2_fill_2 FILLER_19_677 ();
 sg13g2_decap_8 FILLER_19_684 ();
 sg13g2_fill_1 FILLER_19_691 ();
 sg13g2_decap_4 FILLER_19_696 ();
 sg13g2_fill_2 FILLER_19_713 ();
 sg13g2_decap_8 FILLER_19_731 ();
 sg13g2_fill_2 FILLER_19_738 ();
 sg13g2_fill_2 FILLER_19_819 ();
 sg13g2_fill_1 FILLER_19_821 ();
 sg13g2_decap_4 FILLER_19_826 ();
 sg13g2_fill_2 FILLER_19_830 ();
 sg13g2_fill_1 FILLER_19_847 ();
 sg13g2_fill_2 FILLER_19_882 ();
 sg13g2_decap_8 FILLER_19_913 ();
 sg13g2_decap_4 FILLER_19_920 ();
 sg13g2_fill_1 FILLER_19_931 ();
 sg13g2_decap_4 FILLER_19_935 ();
 sg13g2_fill_2 FILLER_19_965 ();
 sg13g2_fill_1 FILLER_19_967 ();
 sg13g2_fill_2 FILLER_19_976 ();
 sg13g2_fill_1 FILLER_19_1008 ();
 sg13g2_decap_4 FILLER_19_1030 ();
 sg13g2_fill_2 FILLER_19_1034 ();
 sg13g2_fill_1 FILLER_19_1040 ();
 sg13g2_fill_2 FILLER_19_1093 ();
 sg13g2_fill_1 FILLER_19_1121 ();
 sg13g2_fill_2 FILLER_19_1178 ();
 sg13g2_fill_1 FILLER_19_1180 ();
 sg13g2_fill_1 FILLER_19_1211 ();
 sg13g2_fill_2 FILLER_19_1220 ();
 sg13g2_decap_8 FILLER_19_1227 ();
 sg13g2_decap_4 FILLER_19_1234 ();
 sg13g2_fill_1 FILLER_19_1238 ();
 sg13g2_decap_8 FILLER_19_1243 ();
 sg13g2_fill_2 FILLER_19_1281 ();
 sg13g2_decap_4 FILLER_19_1287 ();
 sg13g2_decap_8 FILLER_19_1356 ();
 sg13g2_decap_8 FILLER_19_1363 ();
 sg13g2_decap_4 FILLER_19_1370 ();
 sg13g2_decap_8 FILLER_19_1378 ();
 sg13g2_decap_4 FILLER_19_1385 ();
 sg13g2_fill_2 FILLER_19_1389 ();
 sg13g2_decap_4 FILLER_19_1426 ();
 sg13g2_fill_2 FILLER_19_1430 ();
 sg13g2_fill_2 FILLER_19_1444 ();
 sg13g2_fill_2 FILLER_19_1450 ();
 sg13g2_fill_2 FILLER_19_1457 ();
 sg13g2_decap_8 FILLER_19_1473 ();
 sg13g2_decap_4 FILLER_19_1480 ();
 sg13g2_fill_2 FILLER_19_1484 ();
 sg13g2_decap_4 FILLER_19_1497 ();
 sg13g2_fill_1 FILLER_19_1505 ();
 sg13g2_fill_2 FILLER_19_1533 ();
 sg13g2_fill_1 FILLER_19_1535 ();
 sg13g2_fill_1 FILLER_19_1552 ();
 sg13g2_fill_1 FILLER_19_1559 ();
 sg13g2_fill_1 FILLER_19_1572 ();
 sg13g2_fill_2 FILLER_19_1586 ();
 sg13g2_fill_1 FILLER_19_1594 ();
 sg13g2_fill_1 FILLER_19_1599 ();
 sg13g2_fill_1 FILLER_19_1625 ();
 sg13g2_fill_1 FILLER_19_1665 ();
 sg13g2_fill_2 FILLER_19_1691 ();
 sg13g2_decap_8 FILLER_19_1697 ();
 sg13g2_fill_2 FILLER_19_1704 ();
 sg13g2_fill_2 FILLER_19_1738 ();
 sg13g2_decap_8 FILLER_19_1758 ();
 sg13g2_fill_1 FILLER_19_1765 ();
 sg13g2_fill_1 FILLER_19_1776 ();
 sg13g2_fill_2 FILLER_19_1781 ();
 sg13g2_fill_1 FILLER_19_1797 ();
 sg13g2_decap_8 FILLER_19_1832 ();
 sg13g2_decap_4 FILLER_19_1839 ();
 sg13g2_fill_1 FILLER_19_1843 ();
 sg13g2_decap_4 FILLER_19_1873 ();
 sg13g2_fill_1 FILLER_19_1877 ();
 sg13g2_fill_2 FILLER_19_1913 ();
 sg13g2_fill_1 FILLER_19_1923 ();
 sg13g2_fill_1 FILLER_19_1976 ();
 sg13g2_fill_2 FILLER_19_2097 ();
 sg13g2_decap_4 FILLER_19_2125 ();
 sg13g2_fill_1 FILLER_19_2129 ();
 sg13g2_decap_8 FILLER_19_2186 ();
 sg13g2_decap_8 FILLER_19_2193 ();
 sg13g2_decap_8 FILLER_19_2200 ();
 sg13g2_fill_2 FILLER_19_2207 ();
 sg13g2_decap_8 FILLER_19_2213 ();
 sg13g2_decap_4 FILLER_19_2220 ();
 sg13g2_fill_2 FILLER_19_2224 ();
 sg13g2_fill_2 FILLER_19_2288 ();
 sg13g2_fill_1 FILLER_19_2290 ();
 sg13g2_fill_2 FILLER_19_2322 ();
 sg13g2_fill_1 FILLER_19_2350 ();
 sg13g2_fill_1 FILLER_19_2390 ();
 sg13g2_fill_1 FILLER_19_2407 ();
 sg13g2_fill_1 FILLER_19_2439 ();
 sg13g2_fill_1 FILLER_19_2444 ();
 sg13g2_fill_2 FILLER_19_2487 ();
 sg13g2_fill_2 FILLER_19_2544 ();
 sg13g2_fill_2 FILLER_19_2550 ();
 sg13g2_fill_1 FILLER_19_2552 ();
 sg13g2_decap_8 FILLER_19_2573 ();
 sg13g2_decap_8 FILLER_19_2580 ();
 sg13g2_fill_2 FILLER_19_2623 ();
 sg13g2_decap_8 FILLER_19_2661 ();
 sg13g2_fill_2 FILLER_19_2668 ();
 sg13g2_fill_2 FILLER_20_0 ();
 sg13g2_fill_2 FILLER_20_43 ();
 sg13g2_decap_4 FILLER_20_81 ();
 sg13g2_fill_2 FILLER_20_111 ();
 sg13g2_fill_1 FILLER_20_113 ();
 sg13g2_fill_1 FILLER_20_118 ();
 sg13g2_fill_1 FILLER_20_124 ();
 sg13g2_fill_1 FILLER_20_151 ();
 sg13g2_decap_4 FILLER_20_162 ();
 sg13g2_fill_1 FILLER_20_166 ();
 sg13g2_fill_2 FILLER_20_201 ();
 sg13g2_fill_1 FILLER_20_207 ();
 sg13g2_fill_2 FILLER_20_212 ();
 sg13g2_fill_1 FILLER_20_214 ();
 sg13g2_decap_4 FILLER_20_227 ();
 sg13g2_decap_4 FILLER_20_257 ();
 sg13g2_decap_4 FILLER_20_291 ();
 sg13g2_fill_2 FILLER_20_295 ();
 sg13g2_decap_4 FILLER_20_301 ();
 sg13g2_fill_1 FILLER_20_305 ();
 sg13g2_fill_2 FILLER_20_317 ();
 sg13g2_fill_2 FILLER_20_334 ();
 sg13g2_fill_2 FILLER_20_342 ();
 sg13g2_decap_8 FILLER_20_348 ();
 sg13g2_decap_8 FILLER_20_355 ();
 sg13g2_decap_4 FILLER_20_362 ();
 sg13g2_fill_2 FILLER_20_366 ();
 sg13g2_fill_2 FILLER_20_372 ();
 sg13g2_decap_4 FILLER_20_400 ();
 sg13g2_fill_2 FILLER_20_409 ();
 sg13g2_decap_8 FILLER_20_420 ();
 sg13g2_fill_1 FILLER_20_427 ();
 sg13g2_fill_2 FILLER_20_433 ();
 sg13g2_decap_8 FILLER_20_439 ();
 sg13g2_fill_1 FILLER_20_446 ();
 sg13g2_fill_2 FILLER_20_529 ();
 sg13g2_fill_1 FILLER_20_531 ();
 sg13g2_fill_2 FILLER_20_563 ();
 sg13g2_decap_4 FILLER_20_591 ();
 sg13g2_fill_1 FILLER_20_595 ();
 sg13g2_fill_1 FILLER_20_601 ();
 sg13g2_fill_2 FILLER_20_628 ();
 sg13g2_fill_1 FILLER_20_639 ();
 sg13g2_decap_4 FILLER_20_669 ();
 sg13g2_fill_1 FILLER_20_673 ();
 sg13g2_fill_2 FILLER_20_688 ();
 sg13g2_fill_1 FILLER_20_690 ();
 sg13g2_fill_2 FILLER_20_696 ();
 sg13g2_fill_1 FILLER_20_698 ();
 sg13g2_fill_2 FILLER_20_704 ();
 sg13g2_decap_4 FILLER_20_711 ();
 sg13g2_fill_1 FILLER_20_715 ();
 sg13g2_fill_2 FILLER_20_722 ();
 sg13g2_fill_1 FILLER_20_724 ();
 sg13g2_fill_2 FILLER_20_752 ();
 sg13g2_fill_2 FILLER_20_758 ();
 sg13g2_fill_2 FILLER_20_765 ();
 sg13g2_fill_1 FILLER_20_767 ();
 sg13g2_fill_2 FILLER_20_772 ();
 sg13g2_fill_1 FILLER_20_774 ();
 sg13g2_fill_1 FILLER_20_780 ();
 sg13g2_fill_1 FILLER_20_786 ();
 sg13g2_fill_1 FILLER_20_792 ();
 sg13g2_fill_1 FILLER_20_802 ();
 sg13g2_fill_2 FILLER_20_813 ();
 sg13g2_fill_2 FILLER_20_841 ();
 sg13g2_fill_2 FILLER_20_896 ();
 sg13g2_decap_4 FILLER_20_924 ();
 sg13g2_fill_1 FILLER_20_928 ();
 sg13g2_fill_2 FILLER_20_941 ();
 sg13g2_fill_1 FILLER_20_943 ();
 sg13g2_fill_1 FILLER_20_978 ();
 sg13g2_fill_1 FILLER_20_1015 ();
 sg13g2_fill_2 FILLER_20_1020 ();
 sg13g2_decap_4 FILLER_20_1095 ();
 sg13g2_fill_2 FILLER_20_1099 ();
 sg13g2_decap_8 FILLER_20_1109 ();
 sg13g2_decap_4 FILLER_20_1116 ();
 sg13g2_fill_2 FILLER_20_1120 ();
 sg13g2_fill_2 FILLER_20_1135 ();
 sg13g2_fill_1 FILLER_20_1137 ();
 sg13g2_fill_2 FILLER_20_1179 ();
 sg13g2_fill_1 FILLER_20_1181 ();
 sg13g2_fill_2 FILLER_20_1217 ();
 sg13g2_fill_1 FILLER_20_1297 ();
 sg13g2_fill_2 FILLER_20_1303 ();
 sg13g2_fill_2 FILLER_20_1310 ();
 sg13g2_fill_2 FILLER_20_1317 ();
 sg13g2_fill_1 FILLER_20_1319 ();
 sg13g2_decap_8 FILLER_20_1346 ();
 sg13g2_decap_4 FILLER_20_1353 ();
 sg13g2_fill_2 FILLER_20_1357 ();
 sg13g2_fill_1 FILLER_20_1399 ();
 sg13g2_decap_8 FILLER_20_1426 ();
 sg13g2_decap_8 FILLER_20_1433 ();
 sg13g2_fill_2 FILLER_20_1440 ();
 sg13g2_fill_1 FILLER_20_1446 ();
 sg13g2_decap_4 FILLER_20_1461 ();
 sg13g2_fill_1 FILLER_20_1474 ();
 sg13g2_fill_1 FILLER_20_1480 ();
 sg13g2_decap_4 FILLER_20_1485 ();
 sg13g2_fill_1 FILLER_20_1489 ();
 sg13g2_fill_2 FILLER_20_1507 ();
 sg13g2_fill_1 FILLER_20_1521 ();
 sg13g2_fill_1 FILLER_20_1537 ();
 sg13g2_fill_1 FILLER_20_1543 ();
 sg13g2_fill_2 FILLER_20_1560 ();
 sg13g2_fill_1 FILLER_20_1622 ();
 sg13g2_fill_1 FILLER_20_1732 ();
 sg13g2_fill_2 FILLER_20_1737 ();
 sg13g2_fill_1 FILLER_20_1739 ();
 sg13g2_fill_2 FILLER_20_1748 ();
 sg13g2_fill_2 FILLER_20_1754 ();
 sg13g2_fill_1 FILLER_20_1756 ();
 sg13g2_fill_2 FILLER_20_1805 ();
 sg13g2_fill_1 FILLER_20_1807 ();
 sg13g2_fill_1 FILLER_20_1976 ();
 sg13g2_decap_4 FILLER_20_2044 ();
 sg13g2_fill_1 FILLER_20_2048 ();
 sg13g2_fill_2 FILLER_20_2089 ();
 sg13g2_fill_1 FILLER_20_2121 ();
 sg13g2_fill_2 FILLER_20_2153 ();
 sg13g2_fill_2 FILLER_20_2172 ();
 sg13g2_fill_1 FILLER_20_2174 ();
 sg13g2_decap_8 FILLER_20_2179 ();
 sg13g2_fill_2 FILLER_20_2186 ();
 sg13g2_fill_2 FILLER_20_2198 ();
 sg13g2_fill_1 FILLER_20_2200 ();
 sg13g2_decap_4 FILLER_20_2237 ();
 sg13g2_fill_2 FILLER_20_2241 ();
 sg13g2_fill_1 FILLER_20_2247 ();
 sg13g2_fill_2 FILLER_20_2258 ();
 sg13g2_fill_2 FILLER_20_2286 ();
 sg13g2_fill_2 FILLER_20_2314 ();
 sg13g2_fill_1 FILLER_20_2316 ();
 sg13g2_fill_1 FILLER_20_2387 ();
 sg13g2_fill_2 FILLER_20_2392 ();
 sg13g2_fill_1 FILLER_20_2425 ();
 sg13g2_fill_2 FILLER_20_2472 ();
 sg13g2_fill_1 FILLER_20_2474 ();
 sg13g2_decap_8 FILLER_20_2479 ();
 sg13g2_fill_2 FILLER_20_2486 ();
 sg13g2_fill_1 FILLER_20_2488 ();
 sg13g2_decap_4 FILLER_20_2517 ();
 sg13g2_fill_1 FILLER_20_2521 ();
 sg13g2_decap_8 FILLER_20_2528 ();
 sg13g2_decap_4 FILLER_20_2545 ();
 sg13g2_decap_8 FILLER_20_2585 ();
 sg13g2_fill_1 FILLER_20_2626 ();
 sg13g2_decap_8 FILLER_20_2637 ();
 sg13g2_fill_1 FILLER_20_2644 ();
 sg13g2_decap_8 FILLER_20_2653 ();
 sg13g2_decap_8 FILLER_20_2660 ();
 sg13g2_fill_2 FILLER_20_2667 ();
 sg13g2_fill_1 FILLER_20_2669 ();
 sg13g2_decap_4 FILLER_21_0 ();
 sg13g2_fill_1 FILLER_21_4 ();
 sg13g2_fill_1 FILLER_21_37 ();
 sg13g2_fill_2 FILLER_21_43 ();
 sg13g2_decap_8 FILLER_21_97 ();
 sg13g2_decap_8 FILLER_21_104 ();
 sg13g2_decap_8 FILLER_21_111 ();
 sg13g2_decap_4 FILLER_21_118 ();
 sg13g2_decap_4 FILLER_21_154 ();
 sg13g2_fill_1 FILLER_21_163 ();
 sg13g2_fill_1 FILLER_21_189 ();
 sg13g2_fill_1 FILLER_21_194 ();
 sg13g2_decap_8 FILLER_21_199 ();
 sg13g2_decap_8 FILLER_21_206 ();
 sg13g2_decap_8 FILLER_21_213 ();
 sg13g2_fill_2 FILLER_21_220 ();
 sg13g2_fill_2 FILLER_21_237 ();
 sg13g2_fill_2 FILLER_21_243 ();
 sg13g2_fill_2 FILLER_21_253 ();
 sg13g2_fill_1 FILLER_21_287 ();
 sg13g2_fill_1 FILLER_21_301 ();
 sg13g2_fill_1 FILLER_21_306 ();
 sg13g2_fill_2 FILLER_21_316 ();
 sg13g2_fill_1 FILLER_21_318 ();
 sg13g2_fill_2 FILLER_21_353 ();
 sg13g2_fill_1 FILLER_21_360 ();
 sg13g2_fill_2 FILLER_21_392 ();
 sg13g2_fill_2 FILLER_21_398 ();
 sg13g2_fill_1 FILLER_21_418 ();
 sg13g2_fill_2 FILLER_21_428 ();
 sg13g2_fill_1 FILLER_21_454 ();
 sg13g2_fill_2 FILLER_21_460 ();
 sg13g2_fill_2 FILLER_21_472 ();
 sg13g2_fill_2 FILLER_21_529 ();
 sg13g2_fill_1 FILLER_21_531 ();
 sg13g2_fill_2 FILLER_21_561 ();
 sg13g2_fill_2 FILLER_21_572 ();
 sg13g2_fill_2 FILLER_21_579 ();
 sg13g2_decap_8 FILLER_21_595 ();
 sg13g2_fill_1 FILLER_21_602 ();
 sg13g2_decap_4 FILLER_21_635 ();
 sg13g2_fill_1 FILLER_21_661 ();
 sg13g2_fill_1 FILLER_21_667 ();
 sg13g2_fill_2 FILLER_21_708 ();
 sg13g2_decap_4 FILLER_21_714 ();
 sg13g2_fill_2 FILLER_21_718 ();
 sg13g2_decap_4 FILLER_21_726 ();
 sg13g2_fill_2 FILLER_21_730 ();
 sg13g2_fill_1 FILLER_21_742 ();
 sg13g2_fill_2 FILLER_21_755 ();
 sg13g2_fill_1 FILLER_21_757 ();
 sg13g2_decap_4 FILLER_21_772 ();
 sg13g2_fill_2 FILLER_21_887 ();
 sg13g2_fill_1 FILLER_21_902 ();
 sg13g2_fill_1 FILLER_21_907 ();
 sg13g2_fill_2 FILLER_21_953 ();
 sg13g2_fill_1 FILLER_21_955 ();
 sg13g2_decap_8 FILLER_21_963 ();
 sg13g2_decap_4 FILLER_21_970 ();
 sg13g2_fill_1 FILLER_21_974 ();
 sg13g2_fill_2 FILLER_21_1032 ();
 sg13g2_fill_1 FILLER_21_1034 ();
 sg13g2_decap_4 FILLER_21_1039 ();
 sg13g2_fill_1 FILLER_21_1043 ();
 sg13g2_fill_1 FILLER_21_1052 ();
 sg13g2_fill_1 FILLER_21_1058 ();
 sg13g2_fill_1 FILLER_21_1063 ();
 sg13g2_fill_1 FILLER_21_1069 ();
 sg13g2_decap_4 FILLER_21_1087 ();
 sg13g2_fill_1 FILLER_21_1091 ();
 sg13g2_fill_2 FILLER_21_1096 ();
 sg13g2_fill_1 FILLER_21_1098 ();
 sg13g2_decap_4 FILLER_21_1103 ();
 sg13g2_decap_8 FILLER_21_1120 ();
 sg13g2_fill_2 FILLER_21_1127 ();
 sg13g2_decap_8 FILLER_21_1133 ();
 sg13g2_fill_2 FILLER_21_1140 ();
 sg13g2_fill_2 FILLER_21_1146 ();
 sg13g2_decap_8 FILLER_21_1178 ();
 sg13g2_fill_2 FILLER_21_1185 ();
 sg13g2_fill_1 FILLER_21_1228 ();
 sg13g2_decap_8 FILLER_21_1233 ();
 sg13g2_decap_8 FILLER_21_1342 ();
 sg13g2_decap_8 FILLER_21_1349 ();
 sg13g2_fill_2 FILLER_21_1356 ();
 sg13g2_decap_8 FILLER_21_1363 ();
 sg13g2_decap_4 FILLER_21_1370 ();
 sg13g2_fill_1 FILLER_21_1374 ();
 sg13g2_fill_1 FILLER_21_1379 ();
 sg13g2_fill_1 FILLER_21_1390 ();
 sg13g2_fill_2 FILLER_21_1401 ();
 sg13g2_fill_2 FILLER_21_1429 ();
 sg13g2_fill_1 FILLER_21_1431 ();
 sg13g2_fill_1 FILLER_21_1436 ();
 sg13g2_decap_4 FILLER_21_1477 ();
 sg13g2_fill_1 FILLER_21_1481 ();
 sg13g2_fill_2 FILLER_21_1494 ();
 sg13g2_fill_1 FILLER_21_1496 ();
 sg13g2_fill_1 FILLER_21_1506 ();
 sg13g2_decap_4 FILLER_21_1519 ();
 sg13g2_fill_2 FILLER_21_1523 ();
 sg13g2_fill_1 FILLER_21_1543 ();
 sg13g2_fill_1 FILLER_21_1560 ();
 sg13g2_fill_2 FILLER_21_1573 ();
 sg13g2_fill_1 FILLER_21_1585 ();
 sg13g2_fill_2 FILLER_21_1599 ();
 sg13g2_fill_1 FILLER_21_1627 ();
 sg13g2_fill_2 FILLER_21_1636 ();
 sg13g2_fill_1 FILLER_21_1652 ();
 sg13g2_fill_2 FILLER_21_1658 ();
 sg13g2_fill_2 FILLER_21_1665 ();
 sg13g2_decap_4 FILLER_21_1732 ();
 sg13g2_fill_1 FILLER_21_1736 ();
 sg13g2_fill_2 FILLER_21_1742 ();
 sg13g2_fill_1 FILLER_21_1744 ();
 sg13g2_decap_8 FILLER_21_1751 ();
 sg13g2_fill_2 FILLER_21_1792 ();
 sg13g2_decap_8 FILLER_21_1813 ();
 sg13g2_fill_1 FILLER_21_1820 ();
 sg13g2_decap_8 FILLER_21_1831 ();
 sg13g2_fill_1 FILLER_21_1838 ();
 sg13g2_fill_1 FILLER_21_1849 ();
 sg13g2_fill_1 FILLER_21_1869 ();
 sg13g2_decap_4 FILLER_21_1936 ();
 sg13g2_fill_1 FILLER_21_1940 ();
 sg13g2_fill_1 FILLER_21_1962 ();
 sg13g2_fill_1 FILLER_21_2015 ();
 sg13g2_decap_8 FILLER_21_2030 ();
 sg13g2_fill_1 FILLER_21_2037 ();
 sg13g2_decap_4 FILLER_21_2055 ();
 sg13g2_fill_2 FILLER_21_2059 ();
 sg13g2_fill_1 FILLER_21_2081 ();
 sg13g2_fill_1 FILLER_21_2092 ();
 sg13g2_decap_8 FILLER_21_2225 ();
 sg13g2_decap_8 FILLER_21_2232 ();
 sg13g2_decap_8 FILLER_21_2239 ();
 sg13g2_decap_4 FILLER_21_2246 ();
 sg13g2_fill_1 FILLER_21_2250 ();
 sg13g2_fill_1 FILLER_21_2280 ();
 sg13g2_decap_4 FILLER_21_2308 ();
 sg13g2_fill_2 FILLER_21_2316 ();
 sg13g2_fill_1 FILLER_21_2318 ();
 sg13g2_fill_1 FILLER_21_2324 ();
 sg13g2_fill_1 FILLER_21_2331 ();
 sg13g2_fill_1 FILLER_21_2336 ();
 sg13g2_fill_1 FILLER_21_2342 ();
 sg13g2_fill_1 FILLER_21_2348 ();
 sg13g2_decap_4 FILLER_21_2353 ();
 sg13g2_fill_2 FILLER_21_2397 ();
 sg13g2_fill_2 FILLER_21_2433 ();
 sg13g2_fill_2 FILLER_21_2447 ();
 sg13g2_decap_8 FILLER_21_2458 ();
 sg13g2_decap_8 FILLER_21_2465 ();
 sg13g2_decap_8 FILLER_21_2472 ();
 sg13g2_decap_8 FILLER_21_2479 ();
 sg13g2_fill_1 FILLER_21_2501 ();
 sg13g2_decap_4 FILLER_21_2560 ();
 sg13g2_fill_1 FILLER_21_2568 ();
 sg13g2_fill_1 FILLER_21_2575 ();
 sg13g2_decap_4 FILLER_21_2631 ();
 sg13g2_decap_4 FILLER_21_2665 ();
 sg13g2_fill_1 FILLER_21_2669 ();
 sg13g2_fill_2 FILLER_22_0 ();
 sg13g2_fill_1 FILLER_22_28 ();
 sg13g2_decap_4 FILLER_22_44 ();
 sg13g2_fill_2 FILLER_22_48 ();
 sg13g2_decap_4 FILLER_22_55 ();
 sg13g2_fill_1 FILLER_22_59 ();
 sg13g2_decap_4 FILLER_22_68 ();
 sg13g2_decap_8 FILLER_22_82 ();
 sg13g2_decap_8 FILLER_22_93 ();
 sg13g2_fill_1 FILLER_22_126 ();
 sg13g2_fill_1 FILLER_22_137 ();
 sg13g2_fill_1 FILLER_22_146 ();
 sg13g2_fill_2 FILLER_22_187 ();
 sg13g2_decap_8 FILLER_22_204 ();
 sg13g2_fill_2 FILLER_22_211 ();
 sg13g2_fill_2 FILLER_22_227 ();
 sg13g2_fill_2 FILLER_22_235 ();
 sg13g2_decap_4 FILLER_22_251 ();
 sg13g2_fill_2 FILLER_22_255 ();
 sg13g2_decap_8 FILLER_22_278 ();
 sg13g2_decap_4 FILLER_22_285 ();
 sg13g2_fill_2 FILLER_22_289 ();
 sg13g2_fill_2 FILLER_22_300 ();
 sg13g2_fill_1 FILLER_22_307 ();
 sg13g2_fill_2 FILLER_22_317 ();
 sg13g2_fill_1 FILLER_22_330 ();
 sg13g2_fill_2 FILLER_22_335 ();
 sg13g2_fill_1 FILLER_22_345 ();
 sg13g2_fill_2 FILLER_22_362 ();
 sg13g2_fill_2 FILLER_22_369 ();
 sg13g2_fill_1 FILLER_22_371 ();
 sg13g2_decap_4 FILLER_22_405 ();
 sg13g2_fill_2 FILLER_22_409 ();
 sg13g2_decap_8 FILLER_22_421 ();
 sg13g2_fill_1 FILLER_22_428 ();
 sg13g2_fill_1 FILLER_22_506 ();
 sg13g2_fill_1 FILLER_22_512 ();
 sg13g2_fill_1 FILLER_22_517 ();
 sg13g2_fill_1 FILLER_22_544 ();
 sg13g2_fill_1 FILLER_22_582 ();
 sg13g2_decap_4 FILLER_22_588 ();
 sg13g2_fill_1 FILLER_22_592 ();
 sg13g2_decap_8 FILLER_22_602 ();
 sg13g2_fill_2 FILLER_22_617 ();
 sg13g2_decap_4 FILLER_22_629 ();
 sg13g2_fill_1 FILLER_22_633 ();
 sg13g2_fill_1 FILLER_22_639 ();
 sg13g2_fill_1 FILLER_22_644 ();
 sg13g2_fill_1 FILLER_22_671 ();
 sg13g2_fill_2 FILLER_22_703 ();
 sg13g2_fill_1 FILLER_22_705 ();
 sg13g2_fill_1 FILLER_22_711 ();
 sg13g2_decap_4 FILLER_22_717 ();
 sg13g2_fill_1 FILLER_22_721 ();
 sg13g2_fill_1 FILLER_22_732 ();
 sg13g2_fill_2 FILLER_22_773 ();
 sg13g2_fill_2 FILLER_22_790 ();
 sg13g2_fill_1 FILLER_22_792 ();
 sg13g2_fill_2 FILLER_22_829 ();
 sg13g2_fill_2 FILLER_22_870 ();
 sg13g2_fill_2 FILLER_22_882 ();
 sg13g2_fill_1 FILLER_22_887 ();
 sg13g2_fill_2 FILLER_22_891 ();
 sg13g2_fill_2 FILLER_22_900 ();
 sg13g2_decap_8 FILLER_22_932 ();
 sg13g2_decap_4 FILLER_22_939 ();
 sg13g2_decap_8 FILLER_22_960 ();
 sg13g2_decap_8 FILLER_22_967 ();
 sg13g2_decap_4 FILLER_22_974 ();
 sg13g2_fill_2 FILLER_22_978 ();
 sg13g2_fill_1 FILLER_22_997 ();
 sg13g2_fill_1 FILLER_22_1003 ();
 sg13g2_fill_2 FILLER_22_1012 ();
 sg13g2_decap_4 FILLER_22_1018 ();
 sg13g2_fill_2 FILLER_22_1022 ();
 sg13g2_fill_2 FILLER_22_1054 ();
 sg13g2_fill_1 FILLER_22_1056 ();
 sg13g2_fill_1 FILLER_22_1074 ();
 sg13g2_fill_2 FILLER_22_1080 ();
 sg13g2_fill_1 FILLER_22_1082 ();
 sg13g2_decap_4 FILLER_22_1139 ();
 sg13g2_fill_2 FILLER_22_1143 ();
 sg13g2_decap_4 FILLER_22_1149 ();
 sg13g2_fill_1 FILLER_22_1153 ();
 sg13g2_fill_1 FILLER_22_1162 ();
 sg13g2_decap_8 FILLER_22_1168 ();
 sg13g2_decap_8 FILLER_22_1175 ();
 sg13g2_decap_4 FILLER_22_1182 ();
 sg13g2_decap_4 FILLER_22_1191 ();
 sg13g2_fill_2 FILLER_22_1199 ();
 sg13g2_fill_1 FILLER_22_1201 ();
 sg13g2_fill_2 FILLER_22_1206 ();
 sg13g2_decap_8 FILLER_22_1229 ();
 sg13g2_decap_8 FILLER_22_1236 ();
 sg13g2_decap_4 FILLER_22_1248 ();
 sg13g2_fill_2 FILLER_22_1252 ();
 sg13g2_fill_1 FILLER_22_1270 ();
 sg13g2_fill_2 FILLER_22_1276 ();
 sg13g2_fill_2 FILLER_22_1282 ();
 sg13g2_fill_1 FILLER_22_1284 ();
 sg13g2_decap_8 FILLER_22_1289 ();
 sg13g2_decap_4 FILLER_22_1296 ();
 sg13g2_fill_1 FILLER_22_1300 ();
 sg13g2_fill_2 FILLER_22_1305 ();
 sg13g2_fill_1 FILLER_22_1311 ();
 sg13g2_fill_2 FILLER_22_1316 ();
 sg13g2_fill_2 FILLER_22_1322 ();
 sg13g2_decap_4 FILLER_22_1345 ();
 sg13g2_decap_8 FILLER_22_1359 ();
 sg13g2_decap_4 FILLER_22_1366 ();
 sg13g2_fill_2 FILLER_22_1370 ();
 sg13g2_fill_2 FILLER_22_1387 ();
 sg13g2_fill_2 FILLER_22_1414 ();
 sg13g2_fill_1 FILLER_22_1416 ();
 sg13g2_decap_4 FILLER_22_1421 ();
 sg13g2_fill_1 FILLER_22_1430 ();
 sg13g2_fill_2 FILLER_22_1441 ();
 sg13g2_fill_1 FILLER_22_1443 ();
 sg13g2_fill_2 FILLER_22_1454 ();
 sg13g2_fill_1 FILLER_22_1456 ();
 sg13g2_decap_8 FILLER_22_1478 ();
 sg13g2_fill_1 FILLER_22_1485 ();
 sg13g2_fill_1 FILLER_22_1499 ();
 sg13g2_fill_2 FILLER_22_1505 ();
 sg13g2_fill_2 FILLER_22_1516 ();
 sg13g2_fill_1 FILLER_22_1528 ();
 sg13g2_fill_1 FILLER_22_1534 ();
 sg13g2_fill_2 FILLER_22_1577 ();
 sg13g2_fill_2 FILLER_22_1621 ();
 sg13g2_fill_1 FILLER_22_1631 ();
 sg13g2_decap_8 FILLER_22_1714 ();
 sg13g2_decap_8 FILLER_22_1721 ();
 sg13g2_decap_8 FILLER_22_1728 ();
 sg13g2_fill_2 FILLER_22_1735 ();
 sg13g2_fill_1 FILLER_22_1737 ();
 sg13g2_decap_8 FILLER_22_1835 ();
 sg13g2_decap_4 FILLER_22_1842 ();
 sg13g2_fill_2 FILLER_22_1846 ();
 sg13g2_fill_1 FILLER_22_1884 ();
 sg13g2_fill_1 FILLER_22_1896 ();
 sg13g2_fill_2 FILLER_22_1914 ();
 sg13g2_decap_8 FILLER_22_1930 ();
 sg13g2_fill_2 FILLER_22_1937 ();
 sg13g2_fill_1 FILLER_22_1939 ();
 sg13g2_fill_2 FILLER_22_1981 ();
 sg13g2_fill_1 FILLER_22_1983 ();
 sg13g2_fill_1 FILLER_22_1988 ();
 sg13g2_fill_2 FILLER_22_2015 ();
 sg13g2_decap_4 FILLER_22_2043 ();
 sg13g2_fill_1 FILLER_22_2047 ();
 sg13g2_fill_1 FILLER_22_2056 ();
 sg13g2_fill_1 FILLER_22_2071 ();
 sg13g2_fill_2 FILLER_22_2107 ();
 sg13g2_decap_8 FILLER_22_2117 ();
 sg13g2_fill_1 FILLER_22_2124 ();
 sg13g2_decap_8 FILLER_22_2150 ();
 sg13g2_decap_4 FILLER_22_2157 ();
 sg13g2_decap_4 FILLER_22_2222 ();
 sg13g2_fill_1 FILLER_22_2226 ();
 sg13g2_fill_2 FILLER_22_2258 ();
 sg13g2_decap_8 FILLER_22_2272 ();
 sg13g2_decap_8 FILLER_22_2279 ();
 sg13g2_decap_8 FILLER_22_2286 ();
 sg13g2_fill_2 FILLER_22_2293 ();
 sg13g2_decap_4 FILLER_22_2299 ();
 sg13g2_fill_1 FILLER_22_2303 ();
 sg13g2_decap_4 FILLER_22_2309 ();
 sg13g2_fill_1 FILLER_22_2313 ();
 sg13g2_fill_2 FILLER_22_2324 ();
 sg13g2_decap_8 FILLER_22_2330 ();
 sg13g2_decap_8 FILLER_22_2337 ();
 sg13g2_decap_8 FILLER_22_2344 ();
 sg13g2_decap_8 FILLER_22_2351 ();
 sg13g2_fill_1 FILLER_22_2358 ();
 sg13g2_fill_1 FILLER_22_2363 ();
 sg13g2_fill_2 FILLER_22_2369 ();
 sg13g2_fill_1 FILLER_22_2430 ();
 sg13g2_fill_2 FILLER_22_2441 ();
 sg13g2_fill_1 FILLER_22_2473 ();
 sg13g2_decap_4 FILLER_22_2478 ();
 sg13g2_fill_2 FILLER_22_2512 ();
 sg13g2_decap_8 FILLER_22_2518 ();
 sg13g2_decap_8 FILLER_22_2525 ();
 sg13g2_decap_8 FILLER_22_2532 ();
 sg13g2_fill_2 FILLER_22_2543 ();
 sg13g2_decap_8 FILLER_22_2551 ();
 sg13g2_decap_8 FILLER_22_2558 ();
 sg13g2_fill_2 FILLER_22_2565 ();
 sg13g2_fill_1 FILLER_22_2567 ();
 sg13g2_fill_2 FILLER_22_2571 ();
 sg13g2_decap_8 FILLER_22_2583 ();
 sg13g2_fill_2 FILLER_22_2590 ();
 sg13g2_fill_2 FILLER_22_2618 ();
 sg13g2_fill_1 FILLER_22_2620 ();
 sg13g2_decap_8 FILLER_22_2657 ();
 sg13g2_decap_4 FILLER_22_2664 ();
 sg13g2_fill_2 FILLER_22_2668 ();
 sg13g2_decap_4 FILLER_23_0 ();
 sg13g2_decap_4 FILLER_23_7 ();
 sg13g2_decap_8 FILLER_23_15 ();
 sg13g2_decap_4 FILLER_23_22 ();
 sg13g2_decap_4 FILLER_23_50 ();
 sg13g2_decap_8 FILLER_23_58 ();
 sg13g2_decap_4 FILLER_23_65 ();
 sg13g2_fill_1 FILLER_23_69 ();
 sg13g2_fill_1 FILLER_23_106 ();
 sg13g2_decap_4 FILLER_23_120 ();
 sg13g2_fill_1 FILLER_23_124 ();
 sg13g2_fill_1 FILLER_23_143 ();
 sg13g2_fill_1 FILLER_23_149 ();
 sg13g2_fill_2 FILLER_23_155 ();
 sg13g2_decap_4 FILLER_23_167 ();
 sg13g2_decap_4 FILLER_23_176 ();
 sg13g2_decap_4 FILLER_23_188 ();
 sg13g2_fill_1 FILLER_23_197 ();
 sg13g2_fill_2 FILLER_23_208 ();
 sg13g2_fill_1 FILLER_23_210 ();
 sg13g2_fill_2 FILLER_23_257 ();
 sg13g2_fill_2 FILLER_23_269 ();
 sg13g2_fill_2 FILLER_23_288 ();
 sg13g2_fill_1 FILLER_23_324 ();
 sg13g2_fill_2 FILLER_23_333 ();
 sg13g2_fill_1 FILLER_23_350 ();
 sg13g2_fill_2 FILLER_23_377 ();
 sg13g2_fill_1 FILLER_23_383 ();
 sg13g2_fill_1 FILLER_23_394 ();
 sg13g2_fill_2 FILLER_23_414 ();
 sg13g2_fill_1 FILLER_23_416 ();
 sg13g2_decap_8 FILLER_23_443 ();
 sg13g2_decap_4 FILLER_23_467 ();
 sg13g2_fill_2 FILLER_23_471 ();
 sg13g2_fill_2 FILLER_23_483 ();
 sg13g2_fill_2 FILLER_23_491 ();
 sg13g2_fill_1 FILLER_23_493 ();
 sg13g2_decap_8 FILLER_23_508 ();
 sg13g2_decap_4 FILLER_23_515 ();
 sg13g2_fill_2 FILLER_23_519 ();
 sg13g2_fill_2 FILLER_23_557 ();
 sg13g2_fill_1 FILLER_23_564 ();
 sg13g2_fill_2 FILLER_23_575 ();
 sg13g2_fill_1 FILLER_23_577 ();
 sg13g2_fill_1 FILLER_23_583 ();
 sg13g2_fill_2 FILLER_23_610 ();
 sg13g2_fill_1 FILLER_23_616 ();
 sg13g2_fill_1 FILLER_23_684 ();
 sg13g2_fill_1 FILLER_23_737 ();
 sg13g2_decap_8 FILLER_23_768 ();
 sg13g2_fill_2 FILLER_23_775 ();
 sg13g2_decap_4 FILLER_23_803 ();
 sg13g2_fill_1 FILLER_23_807 ();
 sg13g2_fill_1 FILLER_23_812 ();
 sg13g2_fill_2 FILLER_23_833 ();
 sg13g2_fill_2 FILLER_23_848 ();
 sg13g2_fill_2 FILLER_23_891 ();
 sg13g2_fill_2 FILLER_23_950 ();
 sg13g2_decap_8 FILLER_23_978 ();
 sg13g2_decap_8 FILLER_23_985 ();
 sg13g2_fill_1 FILLER_23_992 ();
 sg13g2_decap_8 FILLER_23_998 ();
 sg13g2_decap_8 FILLER_23_1005 ();
 sg13g2_fill_2 FILLER_23_1012 ();
 sg13g2_fill_1 FILLER_23_1019 ();
 sg13g2_fill_1 FILLER_23_1120 ();
 sg13g2_fill_2 FILLER_23_1217 ();
 sg13g2_decap_8 FILLER_23_1223 ();
 sg13g2_fill_2 FILLER_23_1230 ();
 sg13g2_fill_1 FILLER_23_1232 ();
 sg13g2_decap_8 FILLER_23_1237 ();
 sg13g2_decap_8 FILLER_23_1244 ();
 sg13g2_fill_2 FILLER_23_1256 ();
 sg13g2_fill_1 FILLER_23_1258 ();
 sg13g2_fill_2 FILLER_23_1264 ();
 sg13g2_fill_2 FILLER_23_1274 ();
 sg13g2_fill_2 FILLER_23_1335 ();
 sg13g2_decap_8 FILLER_23_1341 ();
 sg13g2_decap_4 FILLER_23_1392 ();
 sg13g2_decap_8 FILLER_23_1417 ();
 sg13g2_fill_1 FILLER_23_1424 ();
 sg13g2_fill_2 FILLER_23_1452 ();
 sg13g2_decap_4 FILLER_23_1480 ();
 sg13g2_fill_1 FILLER_23_1484 ();
 sg13g2_decap_4 FILLER_23_1498 ();
 sg13g2_decap_8 FILLER_23_1506 ();
 sg13g2_decap_8 FILLER_23_1513 ();
 sg13g2_decap_8 FILLER_23_1520 ();
 sg13g2_fill_2 FILLER_23_1551 ();
 sg13g2_fill_2 FILLER_23_1579 ();
 sg13g2_fill_2 FILLER_23_1674 ();
 sg13g2_decap_8 FILLER_23_1712 ();
 sg13g2_decap_8 FILLER_23_1719 ();
 sg13g2_decap_4 FILLER_23_1726 ();
 sg13g2_decap_4 FILLER_23_1734 ();
 sg13g2_fill_2 FILLER_23_1738 ();
 sg13g2_decap_4 FILLER_23_1744 ();
 sg13g2_decap_4 FILLER_23_1765 ();
 sg13g2_fill_2 FILLER_23_1769 ();
 sg13g2_decap_8 FILLER_23_1775 ();
 sg13g2_decap_4 FILLER_23_1782 ();
 sg13g2_fill_2 FILLER_23_1786 ();
 sg13g2_decap_4 FILLER_23_1832 ();
 sg13g2_fill_1 FILLER_23_1836 ();
 sg13g2_fill_1 FILLER_23_1884 ();
 sg13g2_decap_8 FILLER_23_1939 ();
 sg13g2_decap_4 FILLER_23_1976 ();
 sg13g2_fill_2 FILLER_23_1980 ();
 sg13g2_fill_1 FILLER_23_1992 ();
 sg13g2_fill_1 FILLER_23_2019 ();
 sg13g2_fill_2 FILLER_23_2046 ();
 sg13g2_fill_2 FILLER_23_2087 ();
 sg13g2_fill_1 FILLER_23_2089 ();
 sg13g2_fill_2 FILLER_23_2095 ();
 sg13g2_fill_1 FILLER_23_2208 ();
 sg13g2_fill_2 FILLER_23_2235 ();
 sg13g2_fill_1 FILLER_23_2237 ();
 sg13g2_fill_2 FILLER_23_2242 ();
 sg13g2_decap_4 FILLER_23_2283 ();
 sg13g2_decap_8 FILLER_23_2297 ();
 sg13g2_fill_1 FILLER_23_2314 ();
 sg13g2_fill_2 FILLER_23_2319 ();
 sg13g2_decap_4 FILLER_23_2347 ();
 sg13g2_fill_1 FILLER_23_2351 ();
 sg13g2_fill_2 FILLER_23_2406 ();
 sg13g2_fill_2 FILLER_23_2466 ();
 sg13g2_decap_4 FILLER_23_2520 ();
 sg13g2_fill_2 FILLER_23_2524 ();
 sg13g2_fill_2 FILLER_23_2529 ();
 sg13g2_fill_1 FILLER_23_2531 ();
 sg13g2_fill_1 FILLER_23_2536 ();
 sg13g2_fill_2 FILLER_23_2543 ();
 sg13g2_decap_4 FILLER_23_2584 ();
 sg13g2_fill_1 FILLER_23_2618 ();
 sg13g2_fill_2 FILLER_23_2640 ();
 sg13g2_fill_1 FILLER_23_2642 ();
 sg13g2_decap_8 FILLER_23_2647 ();
 sg13g2_decap_8 FILLER_23_2654 ();
 sg13g2_decap_8 FILLER_23_2661 ();
 sg13g2_fill_2 FILLER_23_2668 ();
 sg13g2_decap_4 FILLER_24_0 ();
 sg13g2_fill_1 FILLER_24_4 ();
 sg13g2_fill_1 FILLER_24_31 ();
 sg13g2_fill_1 FILLER_24_40 ();
 sg13g2_fill_2 FILLER_24_44 ();
 sg13g2_decap_8 FILLER_24_51 ();
 sg13g2_decap_8 FILLER_24_58 ();
 sg13g2_decap_4 FILLER_24_65 ();
 sg13g2_fill_1 FILLER_24_73 ();
 sg13g2_decap_8 FILLER_24_114 ();
 sg13g2_decap_4 FILLER_24_121 ();
 sg13g2_decap_8 FILLER_24_142 ();
 sg13g2_decap_8 FILLER_24_149 ();
 sg13g2_fill_2 FILLER_24_161 ();
 sg13g2_fill_1 FILLER_24_163 ();
 sg13g2_fill_1 FILLER_24_168 ();
 sg13g2_fill_1 FILLER_24_179 ();
 sg13g2_decap_8 FILLER_24_232 ();
 sg13g2_decap_4 FILLER_24_249 ();
 sg13g2_fill_1 FILLER_24_261 ();
 sg13g2_fill_1 FILLER_24_275 ();
 sg13g2_fill_2 FILLER_24_284 ();
 sg13g2_decap_8 FILLER_24_290 ();
 sg13g2_fill_2 FILLER_24_297 ();
 sg13g2_fill_2 FILLER_24_303 ();
 sg13g2_fill_1 FILLER_24_305 ();
 sg13g2_fill_2 FILLER_24_320 ();
 sg13g2_fill_2 FILLER_24_339 ();
 sg13g2_fill_1 FILLER_24_352 ();
 sg13g2_fill_1 FILLER_24_356 ();
 sg13g2_fill_1 FILLER_24_363 ();
 sg13g2_fill_1 FILLER_24_369 ();
 sg13g2_decap_4 FILLER_24_396 ();
 sg13g2_fill_1 FILLER_24_430 ();
 sg13g2_fill_2 FILLER_24_441 ();
 sg13g2_fill_1 FILLER_24_443 ();
 sg13g2_fill_2 FILLER_24_460 ();
 sg13g2_fill_1 FILLER_24_462 ();
 sg13g2_fill_1 FILLER_24_471 ();
 sg13g2_decap_8 FILLER_24_477 ();
 sg13g2_fill_2 FILLER_24_484 ();
 sg13g2_fill_1 FILLER_24_517 ();
 sg13g2_fill_1 FILLER_24_522 ();
 sg13g2_fill_1 FILLER_24_528 ();
 sg13g2_fill_1 FILLER_24_533 ();
 sg13g2_fill_2 FILLER_24_540 ();
 sg13g2_fill_1 FILLER_24_547 ();
 sg13g2_fill_1 FILLER_24_553 ();
 sg13g2_decap_8 FILLER_24_563 ();
 sg13g2_fill_1 FILLER_24_580 ();
 sg13g2_fill_2 FILLER_24_587 ();
 sg13g2_fill_2 FILLER_24_602 ();
 sg13g2_fill_2 FILLER_24_631 ();
 sg13g2_fill_1 FILLER_24_633 ();
 sg13g2_fill_1 FILLER_24_660 ();
 sg13g2_fill_2 FILLER_24_677 ();
 sg13g2_fill_2 FILLER_24_694 ();
 sg13g2_fill_2 FILLER_24_711 ();
 sg13g2_fill_1 FILLER_24_713 ();
 sg13g2_fill_1 FILLER_24_719 ();
 sg13g2_fill_2 FILLER_24_724 ();
 sg13g2_fill_2 FILLER_24_741 ();
 sg13g2_fill_1 FILLER_24_743 ();
 sg13g2_decap_8 FILLER_24_785 ();
 sg13g2_decap_4 FILLER_24_792 ();
 sg13g2_fill_1 FILLER_24_840 ();
 sg13g2_fill_2 FILLER_24_844 ();
 sg13g2_fill_2 FILLER_24_912 ();
 sg13g2_fill_1 FILLER_24_914 ();
 sg13g2_decap_4 FILLER_24_981 ();
 sg13g2_fill_2 FILLER_24_1020 ();
 sg13g2_fill_1 FILLER_24_1022 ();
 sg13g2_fill_1 FILLER_24_1032 ();
 sg13g2_fill_2 FILLER_24_1037 ();
 sg13g2_fill_1 FILLER_24_1039 ();
 sg13g2_fill_2 FILLER_24_1061 ();
 sg13g2_decap_8 FILLER_24_1150 ();
 sg13g2_fill_2 FILLER_24_1157 ();
 sg13g2_fill_1 FILLER_24_1167 ();
 sg13g2_decap_4 FILLER_24_1203 ();
 sg13g2_fill_2 FILLER_24_1242 ();
 sg13g2_fill_1 FILLER_24_1244 ();
 sg13g2_fill_2 FILLER_24_1280 ();
 sg13g2_fill_1 FILLER_24_1282 ();
 sg13g2_fill_1 FILLER_24_1318 ();
 sg13g2_decap_4 FILLER_24_1349 ();
 sg13g2_fill_1 FILLER_24_1353 ();
 sg13g2_fill_1 FILLER_24_1432 ();
 sg13g2_fill_2 FILLER_24_1468 ();
 sg13g2_decap_8 FILLER_24_1506 ();
 sg13g2_decap_4 FILLER_24_1513 ();
 sg13g2_fill_1 FILLER_24_1517 ();
 sg13g2_fill_1 FILLER_24_1552 ();
 sg13g2_fill_1 FILLER_24_1608 ();
 sg13g2_fill_2 FILLER_24_1638 ();
 sg13g2_fill_1 FILLER_24_1643 ();
 sg13g2_decap_8 FILLER_24_1694 ();
 sg13g2_decap_8 FILLER_24_1701 ();
 sg13g2_fill_2 FILLER_24_1708 ();
 sg13g2_decap_8 FILLER_24_1714 ();
 sg13g2_decap_8 FILLER_24_1721 ();
 sg13g2_decap_8 FILLER_24_1728 ();
 sg13g2_decap_8 FILLER_24_1735 ();
 sg13g2_decap_8 FILLER_24_1742 ();
 sg13g2_decap_8 FILLER_24_1749 ();
 sg13g2_decap_8 FILLER_24_1756 ();
 sg13g2_decap_8 FILLER_24_1763 ();
 sg13g2_decap_8 FILLER_24_1770 ();
 sg13g2_decap_8 FILLER_24_1777 ();
 sg13g2_fill_1 FILLER_24_1784 ();
 sg13g2_fill_2 FILLER_24_1789 ();
 sg13g2_fill_1 FILLER_24_1791 ();
 sg13g2_fill_1 FILLER_24_1796 ();
 sg13g2_fill_1 FILLER_24_1807 ();
 sg13g2_fill_2 FILLER_24_1812 ();
 sg13g2_fill_1 FILLER_24_1814 ();
 sg13g2_decap_8 FILLER_24_1819 ();
 sg13g2_decap_4 FILLER_24_1846 ();
 sg13g2_fill_2 FILLER_24_1850 ();
 sg13g2_fill_2 FILLER_24_1888 ();
 sg13g2_fill_1 FILLER_24_1916 ();
 sg13g2_fill_1 FILLER_24_2031 ();
 sg13g2_fill_2 FILLER_24_2036 ();
 sg13g2_fill_2 FILLER_24_2053 ();
 sg13g2_fill_1 FILLER_24_2055 ();
 sg13g2_fill_2 FILLER_24_2074 ();
 sg13g2_fill_1 FILLER_24_2076 ();
 sg13g2_fill_2 FILLER_24_2113 ();
 sg13g2_fill_1 FILLER_24_2115 ();
 sg13g2_fill_1 FILLER_24_2126 ();
 sg13g2_fill_2 FILLER_24_2153 ();
 sg13g2_decap_4 FILLER_24_2173 ();
 sg13g2_fill_2 FILLER_24_2177 ();
 sg13g2_fill_1 FILLER_24_2183 ();
 sg13g2_decap_8 FILLER_24_2188 ();
 sg13g2_fill_2 FILLER_24_2195 ();
 sg13g2_fill_1 FILLER_24_2197 ();
 sg13g2_fill_2 FILLER_24_2218 ();
 sg13g2_fill_2 FILLER_24_2267 ();
 sg13g2_fill_1 FILLER_24_2269 ();
 sg13g2_fill_2 FILLER_24_2274 ();
 sg13g2_decap_4 FILLER_24_2302 ();
 sg13g2_fill_2 FILLER_24_2306 ();
 sg13g2_fill_2 FILLER_24_2334 ();
 sg13g2_fill_2 FILLER_24_2340 ();
 sg13g2_fill_2 FILLER_24_2346 ();
 sg13g2_decap_8 FILLER_24_2354 ();
 sg13g2_fill_1 FILLER_24_2361 ();
 sg13g2_fill_2 FILLER_24_2398 ();
 sg13g2_decap_4 FILLER_24_2462 ();
 sg13g2_fill_2 FILLER_24_2508 ();
 sg13g2_fill_2 FILLER_24_2550 ();
 sg13g2_decap_8 FILLER_24_2614 ();
 sg13g2_decap_8 FILLER_24_2621 ();
 sg13g2_decap_4 FILLER_24_2628 ();
 sg13g2_fill_2 FILLER_24_2632 ();
 sg13g2_decap_8 FILLER_24_2648 ();
 sg13g2_decap_8 FILLER_24_2655 ();
 sg13g2_decap_8 FILLER_24_2662 ();
 sg13g2_fill_1 FILLER_24_2669 ();
 sg13g2_decap_4 FILLER_25_0 ();
 sg13g2_fill_1 FILLER_25_83 ();
 sg13g2_decap_4 FILLER_25_98 ();
 sg13g2_decap_8 FILLER_25_107 ();
 sg13g2_decap_8 FILLER_25_114 ();
 sg13g2_decap_8 FILLER_25_121 ();
 sg13g2_fill_2 FILLER_25_128 ();
 sg13g2_fill_2 FILLER_25_175 ();
 sg13g2_fill_1 FILLER_25_177 ();
 sg13g2_decap_4 FILLER_25_209 ();
 sg13g2_fill_1 FILLER_25_213 ();
 sg13g2_decap_8 FILLER_25_218 ();
 sg13g2_decap_8 FILLER_25_225 ();
 sg13g2_decap_8 FILLER_25_232 ();
 sg13g2_fill_2 FILLER_25_239 ();
 sg13g2_decap_8 FILLER_25_273 ();
 sg13g2_decap_4 FILLER_25_355 ();
 sg13g2_fill_1 FILLER_25_359 ();
 sg13g2_fill_2 FILLER_25_363 ();
 sg13g2_fill_1 FILLER_25_369 ();
 sg13g2_fill_2 FILLER_25_374 ();
 sg13g2_decap_8 FILLER_25_385 ();
 sg13g2_decap_8 FILLER_25_392 ();
 sg13g2_decap_4 FILLER_25_399 ();
 sg13g2_fill_2 FILLER_25_403 ();
 sg13g2_decap_4 FILLER_25_426 ();
 sg13g2_fill_1 FILLER_25_430 ();
 sg13g2_decap_4 FILLER_25_435 ();
 sg13g2_fill_2 FILLER_25_439 ();
 sg13g2_decap_8 FILLER_25_447 ();
 sg13g2_fill_2 FILLER_25_454 ();
 sg13g2_fill_1 FILLER_25_456 ();
 sg13g2_fill_2 FILLER_25_488 ();
 sg13g2_fill_1 FILLER_25_490 ();
 sg13g2_decap_8 FILLER_25_505 ();
 sg13g2_fill_2 FILLER_25_512 ();
 sg13g2_decap_8 FILLER_25_523 ();
 sg13g2_fill_1 FILLER_25_530 ();
 sg13g2_decap_8 FILLER_25_536 ();
 sg13g2_decap_4 FILLER_25_543 ();
 sg13g2_fill_1 FILLER_25_552 ();
 sg13g2_decap_8 FILLER_25_557 ();
 sg13g2_fill_1 FILLER_25_569 ();
 sg13g2_decap_4 FILLER_25_575 ();
 sg13g2_fill_1 FILLER_25_579 ();
 sg13g2_decap_8 FILLER_25_598 ();
 sg13g2_fill_2 FILLER_25_605 ();
 sg13g2_fill_1 FILLER_25_607 ();
 sg13g2_fill_1 FILLER_25_616 ();
 sg13g2_decap_4 FILLER_25_634 ();
 sg13g2_fill_2 FILLER_25_648 ();
 sg13g2_fill_2 FILLER_25_655 ();
 sg13g2_fill_2 FILLER_25_709 ();
 sg13g2_decap_8 FILLER_25_716 ();
 sg13g2_decap_8 FILLER_25_723 ();
 sg13g2_decap_8 FILLER_25_730 ();
 sg13g2_fill_1 FILLER_25_737 ();
 sg13g2_decap_8 FILLER_25_748 ();
 sg13g2_fill_2 FILLER_25_755 ();
 sg13g2_decap_8 FILLER_25_765 ();
 sg13g2_fill_1 FILLER_25_772 ();
 sg13g2_decap_8 FILLER_25_778 ();
 sg13g2_fill_1 FILLER_25_785 ();
 sg13g2_fill_2 FILLER_25_791 ();
 sg13g2_fill_1 FILLER_25_798 ();
 sg13g2_fill_2 FILLER_25_839 ();
 sg13g2_fill_2 FILLER_25_850 ();
 sg13g2_fill_2 FILLER_25_885 ();
 sg13g2_fill_1 FILLER_25_927 ();
 sg13g2_fill_2 FILLER_25_968 ();
 sg13g2_decap_8 FILLER_25_974 ();
 sg13g2_decap_8 FILLER_25_981 ();
 sg13g2_fill_1 FILLER_25_988 ();
 sg13g2_fill_1 FILLER_25_1019 ();
 sg13g2_fill_1 FILLER_25_1024 ();
 sg13g2_fill_1 FILLER_25_1051 ();
 sg13g2_fill_1 FILLER_25_1062 ();
 sg13g2_fill_2 FILLER_25_1067 ();
 sg13g2_fill_2 FILLER_25_1073 ();
 sg13g2_decap_8 FILLER_25_1105 ();
 sg13g2_fill_2 FILLER_25_1112 ();
 sg13g2_fill_1 FILLER_25_1114 ();
 sg13g2_fill_2 FILLER_25_1129 ();
 sg13g2_fill_1 FILLER_25_1152 ();
 sg13g2_decap_8 FILLER_25_1192 ();
 sg13g2_fill_1 FILLER_25_1199 ();
 sg13g2_fill_2 FILLER_25_1204 ();
 sg13g2_fill_1 FILLER_25_1206 ();
 sg13g2_decap_4 FILLER_25_1306 ();
 sg13g2_fill_2 FILLER_25_1331 ();
 sg13g2_decap_8 FILLER_25_1390 ();
 sg13g2_fill_1 FILLER_25_1397 ();
 sg13g2_decap_4 FILLER_25_1412 ();
 sg13g2_fill_2 FILLER_25_1430 ();
 sg13g2_fill_1 FILLER_25_1432 ();
 sg13g2_fill_1 FILLER_25_1459 ();
 sg13g2_decap_4 FILLER_25_1496 ();
 sg13g2_fill_1 FILLER_25_1500 ();
 sg13g2_fill_1 FILLER_25_1555 ();
 sg13g2_fill_1 FILLER_25_1569 ();
 sg13g2_fill_1 FILLER_25_1631 ();
 sg13g2_fill_1 FILLER_25_1647 ();
 sg13g2_decap_8 FILLER_25_1663 ();
 sg13g2_decap_4 FILLER_25_1673 ();
 sg13g2_fill_1 FILLER_25_1677 ();
 sg13g2_decap_4 FILLER_25_1694 ();
 sg13g2_fill_2 FILLER_25_1737 ();
 sg13g2_fill_2 FILLER_25_1743 ();
 sg13g2_decap_8 FILLER_25_1749 ();
 sg13g2_decap_4 FILLER_25_1756 ();
 sg13g2_decap_4 FILLER_25_1793 ();
 sg13g2_fill_2 FILLER_25_1797 ();
 sg13g2_decap_8 FILLER_25_1802 ();
 sg13g2_decap_8 FILLER_25_1809 ();
 sg13g2_decap_8 FILLER_25_1816 ();
 sg13g2_decap_8 FILLER_25_1823 ();
 sg13g2_fill_2 FILLER_25_1830 ();
 sg13g2_fill_2 FILLER_25_1950 ();
 sg13g2_decap_4 FILLER_25_1976 ();
 sg13g2_fill_1 FILLER_25_1988 ();
 sg13g2_fill_2 FILLER_25_1993 ();
 sg13g2_fill_1 FILLER_25_1999 ();
 sg13g2_fill_2 FILLER_25_2005 ();
 sg13g2_fill_1 FILLER_25_2017 ();
 sg13g2_fill_2 FILLER_25_2084 ();
 sg13g2_fill_1 FILLER_25_2086 ();
 sg13g2_fill_1 FILLER_25_2113 ();
 sg13g2_fill_2 FILLER_25_2119 ();
 sg13g2_fill_1 FILLER_25_2121 ();
 sg13g2_decap_4 FILLER_25_2126 ();
 sg13g2_decap_8 FILLER_25_2140 ();
 sg13g2_decap_4 FILLER_25_2147 ();
 sg13g2_fill_1 FILLER_25_2151 ();
 sg13g2_decap_4 FILLER_25_2157 ();
 sg13g2_decap_8 FILLER_25_2165 ();
 sg13g2_decap_8 FILLER_25_2172 ();
 sg13g2_decap_4 FILLER_25_2179 ();
 sg13g2_fill_1 FILLER_25_2183 ();
 sg13g2_decap_8 FILLER_25_2194 ();
 sg13g2_decap_4 FILLER_25_2201 ();
 sg13g2_fill_2 FILLER_25_2205 ();
 sg13g2_fill_2 FILLER_25_2243 ();
 sg13g2_fill_1 FILLER_25_2245 ();
 sg13g2_decap_8 FILLER_25_2267 ();
 sg13g2_decap_8 FILLER_25_2274 ();
 sg13g2_fill_2 FILLER_25_2281 ();
 sg13g2_fill_1 FILLER_25_2283 ();
 sg13g2_fill_1 FILLER_25_2324 ();
 sg13g2_fill_1 FILLER_25_2331 ();
 sg13g2_fill_2 FILLER_25_2342 ();
 sg13g2_fill_2 FILLER_25_2370 ();
 sg13g2_fill_1 FILLER_25_2372 ();
 sg13g2_fill_2 FILLER_25_2377 ();
 sg13g2_fill_1 FILLER_25_2379 ();
 sg13g2_fill_2 FILLER_25_2386 ();
 sg13g2_fill_1 FILLER_25_2392 ();
 sg13g2_fill_2 FILLER_25_2417 ();
 sg13g2_fill_1 FILLER_25_2431 ();
 sg13g2_fill_1 FILLER_25_2438 ();
 sg13g2_fill_1 FILLER_25_2449 ();
 sg13g2_fill_1 FILLER_25_2491 ();
 sg13g2_decap_4 FILLER_25_2502 ();
 sg13g2_fill_2 FILLER_25_2506 ();
 sg13g2_fill_1 FILLER_25_2520 ();
 sg13g2_fill_1 FILLER_25_2525 ();
 sg13g2_fill_1 FILLER_25_2535 ();
 sg13g2_fill_1 FILLER_25_2546 ();
 sg13g2_fill_1 FILLER_25_2557 ();
 sg13g2_fill_2 FILLER_25_2562 ();
 sg13g2_fill_1 FILLER_25_2574 ();
 sg13g2_fill_1 FILLER_25_2589 ();
 sg13g2_decap_8 FILLER_25_2616 ();
 sg13g2_decap_4 FILLER_25_2623 ();
 sg13g2_decap_8 FILLER_25_2663 ();
 sg13g2_fill_2 FILLER_26_0 ();
 sg13g2_fill_1 FILLER_26_2 ();
 sg13g2_fill_2 FILLER_26_46 ();
 sg13g2_decap_4 FILLER_26_87 ();
 sg13g2_fill_2 FILLER_26_143 ();
 sg13g2_fill_2 FILLER_26_150 ();
 sg13g2_fill_1 FILLER_26_196 ();
 sg13g2_fill_1 FILLER_26_208 ();
 sg13g2_decap_4 FILLER_26_224 ();
 sg13g2_fill_1 FILLER_26_228 ();
 sg13g2_decap_8 FILLER_26_233 ();
 sg13g2_fill_2 FILLER_26_240 ();
 sg13g2_fill_1 FILLER_26_242 ();
 sg13g2_fill_2 FILLER_26_246 ();
 sg13g2_decap_4 FILLER_26_260 ();
 sg13g2_fill_2 FILLER_26_291 ();
 sg13g2_decap_8 FILLER_26_319 ();
 sg13g2_fill_2 FILLER_26_326 ();
 sg13g2_decap_8 FILLER_26_371 ();
 sg13g2_fill_1 FILLER_26_383 ();
 sg13g2_fill_2 FILLER_26_389 ();
 sg13g2_fill_1 FILLER_26_395 ();
 sg13g2_fill_1 FILLER_26_441 ();
 sg13g2_fill_2 FILLER_26_452 ();
 sg13g2_fill_1 FILLER_26_454 ();
 sg13g2_fill_2 FILLER_26_460 ();
 sg13g2_fill_1 FILLER_26_462 ();
 sg13g2_fill_2 FILLER_26_489 ();
 sg13g2_decap_8 FILLER_26_505 ();
 sg13g2_fill_1 FILLER_26_561 ();
 sg13g2_fill_2 FILLER_26_594 ();
 sg13g2_decap_8 FILLER_26_605 ();
 sg13g2_decap_8 FILLER_26_652 ();
 sg13g2_fill_2 FILLER_26_667 ();
 sg13g2_decap_8 FILLER_26_675 ();
 sg13g2_decap_4 FILLER_26_682 ();
 sg13g2_fill_1 FILLER_26_686 ();
 sg13g2_decap_8 FILLER_26_694 ();
 sg13g2_fill_2 FILLER_26_701 ();
 sg13g2_fill_1 FILLER_26_703 ();
 sg13g2_decap_4 FILLER_26_717 ();
 sg13g2_decap_4 FILLER_26_725 ();
 sg13g2_fill_1 FILLER_26_729 ();
 sg13g2_fill_2 FILLER_26_745 ();
 sg13g2_fill_1 FILLER_26_747 ();
 sg13g2_fill_1 FILLER_26_754 ();
 sg13g2_decap_4 FILLER_26_769 ();
 sg13g2_fill_2 FILLER_26_799 ();
 sg13g2_decap_8 FILLER_26_816 ();
 sg13g2_fill_2 FILLER_26_823 ();
 sg13g2_decap_4 FILLER_26_859 ();
 sg13g2_fill_1 FILLER_26_863 ();
 sg13g2_decap_8 FILLER_26_868 ();
 sg13g2_decap_8 FILLER_26_875 ();
 sg13g2_fill_2 FILLER_26_882 ();
 sg13g2_fill_2 FILLER_26_922 ();
 sg13g2_fill_2 FILLER_26_947 ();
 sg13g2_fill_1 FILLER_26_1015 ();
 sg13g2_fill_1 FILLER_26_1021 ();
 sg13g2_decap_4 FILLER_26_1027 ();
 sg13g2_fill_2 FILLER_26_1039 ();
 sg13g2_decap_8 FILLER_26_1050 ();
 sg13g2_fill_1 FILLER_26_1057 ();
 sg13g2_fill_2 FILLER_26_1063 ();
 sg13g2_decap_4 FILLER_26_1069 ();
 sg13g2_decap_4 FILLER_26_1078 ();
 sg13g2_decap_8 FILLER_26_1094 ();
 sg13g2_decap_8 FILLER_26_1101 ();
 sg13g2_decap_8 FILLER_26_1108 ();
 sg13g2_decap_8 FILLER_26_1115 ();
 sg13g2_decap_8 FILLER_26_1152 ();
 sg13g2_fill_2 FILLER_26_1159 ();
 sg13g2_fill_1 FILLER_26_1170 ();
 sg13g2_fill_1 FILLER_26_1175 ();
 sg13g2_decap_8 FILLER_26_1197 ();
 sg13g2_fill_2 FILLER_26_1204 ();
 sg13g2_fill_1 FILLER_26_1206 ();
 sg13g2_fill_1 FILLER_26_1211 ();
 sg13g2_decap_4 FILLER_26_1238 ();
 sg13g2_fill_1 FILLER_26_1242 ();
 sg13g2_fill_1 FILLER_26_1248 ();
 sg13g2_fill_2 FILLER_26_1300 ();
 sg13g2_decap_8 FILLER_26_1323 ();
 sg13g2_decap_4 FILLER_26_1330 ();
 sg13g2_fill_1 FILLER_26_1334 ();
 sg13g2_fill_2 FILLER_26_1339 ();
 sg13g2_fill_1 FILLER_26_1341 ();
 sg13g2_decap_8 FILLER_26_1352 ();
 sg13g2_fill_1 FILLER_26_1359 ();
 sg13g2_decap_4 FILLER_26_1364 ();
 sg13g2_fill_1 FILLER_26_1368 ();
 sg13g2_fill_2 FILLER_26_1377 ();
 sg13g2_fill_1 FILLER_26_1379 ();
 sg13g2_decap_4 FILLER_26_1419 ();
 sg13g2_decap_8 FILLER_26_1440 ();
 sg13g2_decap_8 FILLER_26_1447 ();
 sg13g2_fill_2 FILLER_26_1454 ();
 sg13g2_fill_1 FILLER_26_1456 ();
 sg13g2_decap_4 FILLER_26_1496 ();
 sg13g2_fill_2 FILLER_26_1500 ();
 sg13g2_fill_1 FILLER_26_1532 ();
 sg13g2_fill_1 FILLER_26_1541 ();
 sg13g2_fill_1 FILLER_26_1555 ();
 sg13g2_fill_1 FILLER_26_1598 ();
 sg13g2_fill_2 FILLER_26_1616 ();
 sg13g2_fill_1 FILLER_26_1618 ();
 sg13g2_decap_8 FILLER_26_1656 ();
 sg13g2_decap_8 FILLER_26_1663 ();
 sg13g2_decap_8 FILLER_26_1670 ();
 sg13g2_decap_4 FILLER_26_1677 ();
 sg13g2_fill_1 FILLER_26_1681 ();
 sg13g2_fill_1 FILLER_26_1695 ();
 sg13g2_fill_1 FILLER_26_1712 ();
 sg13g2_fill_1 FILLER_26_1731 ();
 sg13g2_fill_1 FILLER_26_1752 ();
 sg13g2_fill_1 FILLER_26_1765 ();
 sg13g2_fill_1 FILLER_26_1770 ();
 sg13g2_fill_1 FILLER_26_1775 ();
 sg13g2_fill_2 FILLER_26_1784 ();
 sg13g2_fill_1 FILLER_26_1786 ();
 sg13g2_fill_1 FILLER_26_1796 ();
 sg13g2_fill_2 FILLER_26_1801 ();
 sg13g2_decap_8 FILLER_26_1807 ();
 sg13g2_decap_8 FILLER_26_1814 ();
 sg13g2_decap_4 FILLER_26_1821 ();
 sg13g2_fill_1 FILLER_26_1832 ();
 sg13g2_fill_1 FILLER_26_1844 ();
 sg13g2_fill_2 FILLER_26_1885 ();
 sg13g2_fill_2 FILLER_26_1917 ();
 sg13g2_fill_2 FILLER_26_1936 ();
 sg13g2_fill_2 FILLER_26_1964 ();
 sg13g2_fill_1 FILLER_26_1966 ();
 sg13g2_fill_2 FILLER_26_1988 ();
 sg13g2_fill_1 FILLER_26_1990 ();
 sg13g2_fill_2 FILLER_26_1999 ();
 sg13g2_fill_1 FILLER_26_2001 ();
 sg13g2_decap_4 FILLER_26_2038 ();
 sg13g2_decap_8 FILLER_26_2046 ();
 sg13g2_decap_8 FILLER_26_2053 ();
 sg13g2_decap_8 FILLER_26_2060 ();
 sg13g2_decap_8 FILLER_26_2067 ();
 sg13g2_decap_8 FILLER_26_2074 ();
 sg13g2_decap_4 FILLER_26_2081 ();
 sg13g2_fill_2 FILLER_26_2085 ();
 sg13g2_decap_4 FILLER_26_2099 ();
 sg13g2_fill_1 FILLER_26_2103 ();
 sg13g2_fill_2 FILLER_26_2112 ();
 sg13g2_fill_1 FILLER_26_2114 ();
 sg13g2_decap_4 FILLER_26_2119 ();
 sg13g2_fill_1 FILLER_26_2123 ();
 sg13g2_decap_4 FILLER_26_2169 ();
 sg13g2_fill_2 FILLER_26_2183 ();
 sg13g2_fill_1 FILLER_26_2185 ();
 sg13g2_decap_8 FILLER_26_2212 ();
 sg13g2_decap_4 FILLER_26_2219 ();
 sg13g2_decap_8 FILLER_26_2227 ();
 sg13g2_fill_2 FILLER_26_2234 ();
 sg13g2_fill_2 FILLER_26_2272 ();
 sg13g2_fill_1 FILLER_26_2274 ();
 sg13g2_decap_4 FILLER_26_2308 ();
 sg13g2_fill_1 FILLER_26_2321 ();
 sg13g2_decap_4 FILLER_26_2327 ();
 sg13g2_fill_2 FILLER_26_2331 ();
 sg13g2_fill_2 FILLER_26_2359 ();
 sg13g2_decap_4 FILLER_26_2365 ();
 sg13g2_fill_1 FILLER_26_2421 ();
 sg13g2_fill_2 FILLER_26_2427 ();
 sg13g2_fill_2 FILLER_26_2491 ();
 sg13g2_fill_1 FILLER_26_2493 ();
 sg13g2_fill_1 FILLER_26_2530 ();
 sg13g2_fill_2 FILLER_26_2593 ();
 sg13g2_fill_1 FILLER_26_2595 ();
 sg13g2_fill_1 FILLER_26_2600 ();
 sg13g2_fill_2 FILLER_26_2605 ();
 sg13g2_fill_1 FILLER_26_2607 ();
 sg13g2_fill_2 FILLER_26_2668 ();
 sg13g2_decap_8 FILLER_27_0 ();
 sg13g2_decap_4 FILLER_27_7 ();
 sg13g2_fill_2 FILLER_27_11 ();
 sg13g2_decap_8 FILLER_27_43 ();
 sg13g2_decap_4 FILLER_27_50 ();
 sg13g2_fill_1 FILLER_27_54 ();
 sg13g2_fill_2 FILLER_27_93 ();
 sg13g2_fill_1 FILLER_27_95 ();
 sg13g2_fill_1 FILLER_27_100 ();
 sg13g2_fill_1 FILLER_27_127 ();
 sg13g2_fill_2 FILLER_27_205 ();
 sg13g2_fill_2 FILLER_27_219 ();
 sg13g2_fill_2 FILLER_27_257 ();
 sg13g2_fill_1 FILLER_27_259 ();
 sg13g2_decap_4 FILLER_27_265 ();
 sg13g2_fill_2 FILLER_27_333 ();
 sg13g2_decap_4 FILLER_27_338 ();
 sg13g2_fill_2 FILLER_27_342 ();
 sg13g2_decap_4 FILLER_27_354 ();
 sg13g2_fill_2 FILLER_27_358 ();
 sg13g2_fill_1 FILLER_27_430 ();
 sg13g2_fill_1 FILLER_27_436 ();
 sg13g2_fill_1 FILLER_27_467 ();
 sg13g2_fill_1 FILLER_27_484 ();
 sg13g2_decap_4 FILLER_27_509 ();
 sg13g2_fill_1 FILLER_27_513 ();
 sg13g2_fill_2 FILLER_27_525 ();
 sg13g2_fill_2 FILLER_27_617 ();
 sg13g2_fill_1 FILLER_27_623 ();
 sg13g2_decap_8 FILLER_27_628 ();
 sg13g2_fill_2 FILLER_27_635 ();
 sg13g2_decap_8 FILLER_27_663 ();
 sg13g2_decap_4 FILLER_27_670 ();
 sg13g2_fill_2 FILLER_27_680 ();
 sg13g2_fill_1 FILLER_27_686 ();
 sg13g2_fill_2 FILLER_27_692 ();
 sg13g2_decap_4 FILLER_27_699 ();
 sg13g2_fill_2 FILLER_27_720 ();
 sg13g2_fill_1 FILLER_27_722 ();
 sg13g2_fill_2 FILLER_27_749 ();
 sg13g2_fill_1 FILLER_27_751 ();
 sg13g2_fill_2 FILLER_27_783 ();
 sg13g2_decap_4 FILLER_27_790 ();
 sg13g2_decap_8 FILLER_27_798 ();
 sg13g2_fill_2 FILLER_27_805 ();
 sg13g2_fill_1 FILLER_27_807 ();
 sg13g2_fill_1 FILLER_27_818 ();
 sg13g2_decap_8 FILLER_27_845 ();
 sg13g2_decap_4 FILLER_27_852 ();
 sg13g2_decap_8 FILLER_27_869 ();
 sg13g2_decap_8 FILLER_27_876 ();
 sg13g2_decap_4 FILLER_27_883 ();
 sg13g2_decap_8 FILLER_27_897 ();
 sg13g2_fill_2 FILLER_27_904 ();
 sg13g2_decap_8 FILLER_27_982 ();
 sg13g2_fill_2 FILLER_27_989 ();
 sg13g2_decap_4 FILLER_27_995 ();
 sg13g2_fill_1 FILLER_27_1008 ();
 sg13g2_decap_8 FILLER_27_1043 ();
 sg13g2_decap_8 FILLER_27_1050 ();
 sg13g2_decap_8 FILLER_27_1078 ();
 sg13g2_decap_4 FILLER_27_1085 ();
 sg13g2_fill_2 FILLER_27_1089 ();
 sg13g2_decap_4 FILLER_27_1100 ();
 sg13g2_fill_1 FILLER_27_1104 ();
 sg13g2_fill_1 FILLER_27_1113 ();
 sg13g2_fill_1 FILLER_27_1127 ();
 sg13g2_decap_4 FILLER_27_1136 ();
 sg13g2_decap_8 FILLER_27_1143 ();
 sg13g2_decap_4 FILLER_27_1150 ();
 sg13g2_decap_8 FILLER_27_1162 ();
 sg13g2_fill_1 FILLER_27_1169 ();
 sg13g2_fill_2 FILLER_27_1196 ();
 sg13g2_decap_8 FILLER_27_1202 ();
 sg13g2_decap_8 FILLER_27_1209 ();
 sg13g2_fill_1 FILLER_27_1216 ();
 sg13g2_decap_8 FILLER_27_1225 ();
 sg13g2_decap_8 FILLER_27_1232 ();
 sg13g2_decap_4 FILLER_27_1239 ();
 sg13g2_decap_8 FILLER_27_1282 ();
 sg13g2_decap_8 FILLER_27_1289 ();
 sg13g2_decap_4 FILLER_27_1296 ();
 sg13g2_decap_8 FILLER_27_1308 ();
 sg13g2_decap_4 FILLER_27_1315 ();
 sg13g2_fill_2 FILLER_27_1319 ();
 sg13g2_decap_8 FILLER_27_1335 ();
 sg13g2_decap_8 FILLER_27_1342 ();
 sg13g2_decap_8 FILLER_27_1349 ();
 sg13g2_decap_8 FILLER_27_1356 ();
 sg13g2_decap_4 FILLER_27_1363 ();
 sg13g2_decap_4 FILLER_27_1371 ();
 sg13g2_fill_1 FILLER_27_1375 ();
 sg13g2_decap_8 FILLER_27_1412 ();
 sg13g2_decap_4 FILLER_27_1423 ();
 sg13g2_fill_2 FILLER_27_1431 ();
 sg13g2_fill_2 FILLER_27_1443 ();
 sg13g2_decap_8 FILLER_27_1466 ();
 sg13g2_decap_8 FILLER_27_1481 ();
 sg13g2_decap_8 FILLER_27_1488 ();
 sg13g2_fill_1 FILLER_27_1495 ();
 sg13g2_fill_2 FILLER_27_1500 ();
 sg13g2_fill_1 FILLER_27_1502 ();
 sg13g2_fill_2 FILLER_27_1507 ();
 sg13g2_fill_1 FILLER_27_1526 ();
 sg13g2_fill_1 FILLER_27_1552 ();
 sg13g2_fill_1 FILLER_27_1558 ();
 sg13g2_decap_8 FILLER_27_1571 ();
 sg13g2_decap_4 FILLER_27_1578 ();
 sg13g2_fill_2 FILLER_27_1586 ();
 sg13g2_fill_1 FILLER_27_1592 ();
 sg13g2_fill_1 FILLER_27_1597 ();
 sg13g2_decap_4 FILLER_27_1602 ();
 sg13g2_fill_2 FILLER_27_1606 ();
 sg13g2_decap_4 FILLER_27_1613 ();
 sg13g2_fill_1 FILLER_27_1631 ();
 sg13g2_fill_2 FILLER_27_1635 ();
 sg13g2_fill_2 FILLER_27_1646 ();
 sg13g2_fill_1 FILLER_27_1682 ();
 sg13g2_fill_2 FILLER_27_1690 ();
 sg13g2_fill_1 FILLER_27_1701 ();
 sg13g2_fill_1 FILLER_27_1707 ();
 sg13g2_fill_2 FILLER_27_1718 ();
 sg13g2_fill_1 FILLER_27_1748 ();
 sg13g2_fill_1 FILLER_27_1756 ();
 sg13g2_fill_1 FILLER_27_1767 ();
 sg13g2_fill_1 FILLER_27_1845 ();
 sg13g2_fill_2 FILLER_27_1850 ();
 sg13g2_fill_2 FILLER_27_1856 ();
 sg13g2_fill_2 FILLER_27_1900 ();
 sg13g2_fill_1 FILLER_27_1939 ();
 sg13g2_decap_8 FILLER_27_1966 ();
 sg13g2_fill_2 FILLER_27_1999 ();
 sg13g2_fill_1 FILLER_27_2005 ();
 sg13g2_decap_8 FILLER_27_2095 ();
 sg13g2_decap_4 FILLER_27_2102 ();
 sg13g2_fill_2 FILLER_27_2106 ();
 sg13g2_fill_2 FILLER_27_2160 ();
 sg13g2_fill_1 FILLER_27_2162 ();
 sg13g2_fill_2 FILLER_27_2225 ();
 sg13g2_decap_4 FILLER_27_2244 ();
 sg13g2_fill_1 FILLER_27_2278 ();
 sg13g2_decap_4 FILLER_27_2296 ();
 sg13g2_fill_1 FILLER_27_2300 ();
 sg13g2_decap_8 FILLER_27_2306 ();
 sg13g2_fill_2 FILLER_27_2313 ();
 sg13g2_decap_8 FILLER_27_2320 ();
 sg13g2_fill_2 FILLER_27_2327 ();
 sg13g2_fill_2 FILLER_27_2343 ();
 sg13g2_fill_2 FILLER_27_2349 ();
 sg13g2_fill_1 FILLER_27_2387 ();
 sg13g2_fill_2 FILLER_27_2420 ();
 sg13g2_fill_1 FILLER_27_2426 ();
 sg13g2_fill_1 FILLER_27_2472 ();
 sg13g2_fill_2 FILLER_27_2484 ();
 sg13g2_fill_1 FILLER_27_2497 ();
 sg13g2_fill_1 FILLER_27_2521 ();
 sg13g2_decap_4 FILLER_27_2581 ();
 sg13g2_fill_1 FILLER_27_2585 ();
 sg13g2_decap_4 FILLER_27_2596 ();
 sg13g2_fill_1 FILLER_27_2656 ();
 sg13g2_decap_8 FILLER_27_2661 ();
 sg13g2_fill_2 FILLER_27_2668 ();
 sg13g2_decap_8 FILLER_28_0 ();
 sg13g2_decap_8 FILLER_28_7 ();
 sg13g2_fill_2 FILLER_28_14 ();
 sg13g2_decap_4 FILLER_28_20 ();
 sg13g2_fill_2 FILLER_28_24 ();
 sg13g2_decap_4 FILLER_28_52 ();
 sg13g2_fill_1 FILLER_28_56 ();
 sg13g2_fill_2 FILLER_28_70 ();
 sg13g2_fill_2 FILLER_28_90 ();
 sg13g2_fill_1 FILLER_28_92 ();
 sg13g2_fill_1 FILLER_28_108 ();
 sg13g2_decap_8 FILLER_28_113 ();
 sg13g2_decap_4 FILLER_28_120 ();
 sg13g2_fill_1 FILLER_28_138 ();
 sg13g2_fill_2 FILLER_28_143 ();
 sg13g2_fill_2 FILLER_28_149 ();
 sg13g2_fill_1 FILLER_28_151 ();
 sg13g2_fill_1 FILLER_28_156 ();
 sg13g2_decap_4 FILLER_28_175 ();
 sg13g2_fill_2 FILLER_28_239 ();
 sg13g2_fill_1 FILLER_28_241 ();
 sg13g2_fill_1 FILLER_28_248 ();
 sg13g2_fill_2 FILLER_28_277 ();
 sg13g2_fill_1 FILLER_28_279 ();
 sg13g2_fill_1 FILLER_28_289 ();
 sg13g2_decap_8 FILLER_28_304 ();
 sg13g2_decap_8 FILLER_28_315 ();
 sg13g2_decap_8 FILLER_28_322 ();
 sg13g2_decap_8 FILLER_28_329 ();
 sg13g2_decap_8 FILLER_28_336 ();
 sg13g2_decap_8 FILLER_28_348 ();
 sg13g2_decap_8 FILLER_28_355 ();
 sg13g2_decap_4 FILLER_28_362 ();
 sg13g2_fill_2 FILLER_28_375 ();
 sg13g2_fill_1 FILLER_28_377 ();
 sg13g2_fill_2 FILLER_28_388 ();
 sg13g2_decap_4 FILLER_28_412 ();
 sg13g2_fill_2 FILLER_28_416 ();
 sg13g2_fill_1 FILLER_28_432 ();
 sg13g2_fill_1 FILLER_28_444 ();
 sg13g2_fill_2 FILLER_28_454 ();
 sg13g2_fill_2 FILLER_28_462 ();
 sg13g2_decap_4 FILLER_28_525 ();
 sg13g2_fill_1 FILLER_28_544 ();
 sg13g2_fill_1 FILLER_28_549 ();
 sg13g2_fill_2 FILLER_28_582 ();
 sg13g2_fill_2 FILLER_28_600 ();
 sg13g2_decap_8 FILLER_28_628 ();
 sg13g2_decap_8 FILLER_28_635 ();
 sg13g2_fill_1 FILLER_28_642 ();
 sg13g2_decap_4 FILLER_28_647 ();
 sg13g2_fill_2 FILLER_28_651 ();
 sg13g2_fill_1 FILLER_28_679 ();
 sg13g2_fill_1 FILLER_28_685 ();
 sg13g2_fill_1 FILLER_28_705 ();
 sg13g2_decap_8 FILLER_28_716 ();
 sg13g2_fill_1 FILLER_28_723 ();
 sg13g2_fill_2 FILLER_28_753 ();
 sg13g2_fill_1 FILLER_28_771 ();
 sg13g2_decap_4 FILLER_28_790 ();
 sg13g2_fill_2 FILLER_28_794 ();
 sg13g2_decap_8 FILLER_28_840 ();
 sg13g2_decap_4 FILLER_28_847 ();
 sg13g2_fill_2 FILLER_28_851 ();
 sg13g2_fill_2 FILLER_28_857 ();
 sg13g2_fill_2 FILLER_28_885 ();
 sg13g2_fill_1 FILLER_28_887 ();
 sg13g2_decap_4 FILLER_28_898 ();
 sg13g2_fill_1 FILLER_28_902 ();
 sg13g2_fill_2 FILLER_28_929 ();
 sg13g2_decap_8 FILLER_28_978 ();
 sg13g2_fill_2 FILLER_28_985 ();
 sg13g2_fill_1 FILLER_28_1002 ();
 sg13g2_fill_1 FILLER_28_1007 ();
 sg13g2_fill_2 FILLER_28_1016 ();
 sg13g2_fill_1 FILLER_28_1018 ();
 sg13g2_decap_4 FILLER_28_1028 ();
 sg13g2_fill_1 FILLER_28_1032 ();
 sg13g2_decap_8 FILLER_28_1037 ();
 sg13g2_fill_1 FILLER_28_1044 ();
 sg13g2_decap_4 FILLER_28_1049 ();
 sg13g2_fill_1 FILLER_28_1053 ();
 sg13g2_decap_4 FILLER_28_1075 ();
 sg13g2_fill_2 FILLER_28_1117 ();
 sg13g2_fill_2 FILLER_28_1144 ();
 sg13g2_fill_1 FILLER_28_1167 ();
 sg13g2_fill_1 FILLER_28_1177 ();
 sg13g2_fill_1 FILLER_28_1182 ();
 sg13g2_fill_2 FILLER_28_1187 ();
 sg13g2_fill_1 FILLER_28_1193 ();
 sg13g2_decap_4 FILLER_28_1203 ();
 sg13g2_fill_2 FILLER_28_1207 ();
 sg13g2_decap_8 FILLER_28_1272 ();
 sg13g2_fill_2 FILLER_28_1279 ();
 sg13g2_fill_1 FILLER_28_1281 ();
 sg13g2_decap_4 FILLER_28_1286 ();
 sg13g2_fill_1 FILLER_28_1290 ();
 sg13g2_fill_2 FILLER_28_1326 ();
 sg13g2_fill_2 FILLER_28_1336 ();
 sg13g2_fill_1 FILLER_28_1338 ();
 sg13g2_decap_4 FILLER_28_1357 ();
 sg13g2_fill_1 FILLER_28_1365 ();
 sg13g2_fill_2 FILLER_28_1405 ();
 sg13g2_fill_1 FILLER_28_1411 ();
 sg13g2_fill_2 FILLER_28_1489 ();
 sg13g2_fill_1 FILLER_28_1496 ();
 sg13g2_fill_1 FILLER_28_1516 ();
 sg13g2_fill_1 FILLER_28_1529 ();
 sg13g2_fill_2 FILLER_28_1557 ();
 sg13g2_decap_4 FILLER_28_1583 ();
 sg13g2_decap_8 FILLER_28_1596 ();
 sg13g2_decap_4 FILLER_28_1603 ();
 sg13g2_fill_2 FILLER_28_1607 ();
 sg13g2_fill_1 FILLER_28_1614 ();
 sg13g2_fill_1 FILLER_28_1620 ();
 sg13g2_decap_8 FILLER_28_1631 ();
 sg13g2_decap_8 FILLER_28_1638 ();
 sg13g2_fill_2 FILLER_28_1645 ();
 sg13g2_fill_1 FILLER_28_1647 ();
 sg13g2_decap_8 FILLER_28_1674 ();
 sg13g2_decap_8 FILLER_28_1681 ();
 sg13g2_fill_2 FILLER_28_1688 ();
 sg13g2_fill_1 FILLER_28_1712 ();
 sg13g2_fill_1 FILLER_28_1738 ();
 sg13g2_fill_1 FILLER_28_1756 ();
 sg13g2_fill_2 FILLER_28_1802 ();
 sg13g2_fill_2 FILLER_28_1808 ();
 sg13g2_fill_1 FILLER_28_1810 ();
 sg13g2_fill_2 FILLER_28_1815 ();
 sg13g2_fill_1 FILLER_28_1817 ();
 sg13g2_fill_1 FILLER_28_1858 ();
 sg13g2_fill_1 FILLER_28_1874 ();
 sg13g2_fill_2 FILLER_28_1897 ();
 sg13g2_fill_2 FILLER_28_1926 ();
 sg13g2_decap_4 FILLER_28_1983 ();
 sg13g2_fill_2 FILLER_28_1987 ();
 sg13g2_fill_1 FILLER_28_2003 ();
 sg13g2_fill_2 FILLER_28_2014 ();
 sg13g2_fill_1 FILLER_28_2046 ();
 sg13g2_fill_1 FILLER_28_2051 ();
 sg13g2_fill_1 FILLER_28_2062 ();
 sg13g2_fill_2 FILLER_28_2089 ();
 sg13g2_decap_8 FILLER_28_2095 ();
 sg13g2_fill_1 FILLER_28_2102 ();
 sg13g2_fill_1 FILLER_28_2150 ();
 sg13g2_decap_4 FILLER_28_2202 ();
 sg13g2_fill_1 FILLER_28_2206 ();
 sg13g2_decap_4 FILLER_28_2211 ();
 sg13g2_fill_1 FILLER_28_2215 ();
 sg13g2_decap_4 FILLER_28_2257 ();
 sg13g2_decap_8 FILLER_28_2265 ();
 sg13g2_decap_8 FILLER_28_2272 ();
 sg13g2_fill_2 FILLER_28_2279 ();
 sg13g2_fill_1 FILLER_28_2281 ();
 sg13g2_fill_2 FILLER_28_2306 ();
 sg13g2_fill_2 FILLER_28_2317 ();
 sg13g2_fill_1 FILLER_28_2335 ();
 sg13g2_fill_2 FILLER_28_2340 ();
 sg13g2_fill_1 FILLER_28_2378 ();
 sg13g2_decap_4 FILLER_28_2399 ();
 sg13g2_fill_1 FILLER_28_2425 ();
 sg13g2_decap_4 FILLER_28_2451 ();
 sg13g2_fill_2 FILLER_28_2460 ();
 sg13g2_fill_1 FILLER_28_2468 ();
 sg13g2_fill_2 FILLER_28_2475 ();
 sg13g2_fill_1 FILLER_28_2487 ();
 sg13g2_fill_1 FILLER_28_2515 ();
 sg13g2_fill_1 FILLER_28_2574 ();
 sg13g2_fill_2 FILLER_28_2581 ();
 sg13g2_fill_2 FILLER_28_2592 ();
 sg13g2_fill_1 FILLER_28_2604 ();
 sg13g2_decap_8 FILLER_28_2612 ();
 sg13g2_fill_2 FILLER_28_2619 ();
 sg13g2_fill_1 FILLER_28_2621 ();
 sg13g2_fill_2 FILLER_28_2668 ();
 sg13g2_decap_8 FILLER_29_0 ();
 sg13g2_fill_2 FILLER_29_7 ();
 sg13g2_decap_8 FILLER_29_13 ();
 sg13g2_decap_8 FILLER_29_20 ();
 sg13g2_decap_4 FILLER_29_27 ();
 sg13g2_fill_1 FILLER_29_31 ();
 sg13g2_fill_1 FILLER_29_69 ();
 sg13g2_fill_2 FILLER_29_78 ();
 sg13g2_fill_1 FILLER_29_80 ();
 sg13g2_decap_4 FILLER_29_85 ();
 sg13g2_fill_2 FILLER_29_89 ();
 sg13g2_decap_8 FILLER_29_112 ();
 sg13g2_decap_8 FILLER_29_119 ();
 sg13g2_decap_4 FILLER_29_126 ();
 sg13g2_fill_2 FILLER_29_130 ();
 sg13g2_decap_8 FILLER_29_136 ();
 sg13g2_decap_8 FILLER_29_143 ();
 sg13g2_decap_8 FILLER_29_150 ();
 sg13g2_decap_8 FILLER_29_157 ();
 sg13g2_fill_1 FILLER_29_164 ();
 sg13g2_fill_1 FILLER_29_169 ();
 sg13g2_fill_2 FILLER_29_179 ();
 sg13g2_fill_1 FILLER_29_207 ();
 sg13g2_fill_1 FILLER_29_212 ();
 sg13g2_decap_8 FILLER_29_221 ();
 sg13g2_fill_2 FILLER_29_228 ();
 sg13g2_fill_1 FILLER_29_230 ();
 sg13g2_decap_4 FILLER_29_239 ();
 sg13g2_fill_1 FILLER_29_243 ();
 sg13g2_fill_2 FILLER_29_268 ();
 sg13g2_fill_2 FILLER_29_292 ();
 sg13g2_fill_1 FILLER_29_294 ();
 sg13g2_decap_4 FILLER_29_300 ();
 sg13g2_decap_8 FILLER_29_308 ();
 sg13g2_decap_8 FILLER_29_315 ();
 sg13g2_decap_4 FILLER_29_322 ();
 sg13g2_fill_2 FILLER_29_326 ();
 sg13g2_decap_4 FILLER_29_332 ();
 sg13g2_decap_8 FILLER_29_340 ();
 sg13g2_decap_4 FILLER_29_347 ();
 sg13g2_fill_2 FILLER_29_351 ();
 sg13g2_fill_2 FILLER_29_383 ();
 sg13g2_fill_1 FILLER_29_385 ();
 sg13g2_decap_8 FILLER_29_406 ();
 sg13g2_decap_8 FILLER_29_413 ();
 sg13g2_fill_2 FILLER_29_420 ();
 sg13g2_fill_1 FILLER_29_422 ();
 sg13g2_decap_8 FILLER_29_443 ();
 sg13g2_fill_1 FILLER_29_450 ();
 sg13g2_fill_2 FILLER_29_464 ();
 sg13g2_fill_1 FILLER_29_498 ();
 sg13g2_fill_2 FILLER_29_507 ();
 sg13g2_fill_2 FILLER_29_547 ();
 sg13g2_fill_2 FILLER_29_559 ();
 sg13g2_fill_2 FILLER_29_581 ();
 sg13g2_decap_4 FILLER_29_617 ();
 sg13g2_fill_1 FILLER_29_621 ();
 sg13g2_decap_8 FILLER_29_632 ();
 sg13g2_decap_4 FILLER_29_639 ();
 sg13g2_fill_2 FILLER_29_643 ();
 sg13g2_fill_2 FILLER_29_649 ();
 sg13g2_fill_1 FILLER_29_651 ();
 sg13g2_fill_1 FILLER_29_658 ();
 sg13g2_fill_2 FILLER_29_687 ();
 sg13g2_fill_2 FILLER_29_693 ();
 sg13g2_fill_1 FILLER_29_695 ();
 sg13g2_fill_2 FILLER_29_702 ();
 sg13g2_fill_2 FILLER_29_729 ();
 sg13g2_decap_4 FILLER_29_761 ();
 sg13g2_fill_2 FILLER_29_774 ();
 sg13g2_fill_1 FILLER_29_780 ();
 sg13g2_fill_2 FILLER_29_791 ();
 sg13g2_fill_1 FILLER_29_793 ();
 sg13g2_fill_2 FILLER_29_804 ();
 sg13g2_fill_1 FILLER_29_806 ();
 sg13g2_decap_8 FILLER_29_843 ();
 sg13g2_fill_2 FILLER_29_850 ();
 sg13g2_fill_1 FILLER_29_852 ();
 sg13g2_fill_2 FILLER_29_873 ();
 sg13g2_decap_4 FILLER_29_901 ();
 sg13g2_fill_2 FILLER_29_931 ();
 sg13g2_fill_2 FILLER_29_963 ();
 sg13g2_fill_1 FILLER_29_996 ();
 sg13g2_fill_1 FILLER_29_1023 ();
 sg13g2_fill_2 FILLER_29_1050 ();
 sg13g2_fill_1 FILLER_29_1052 ();
 sg13g2_fill_2 FILLER_29_1063 ();
 sg13g2_fill_1 FILLER_29_1065 ();
 sg13g2_fill_1 FILLER_29_1092 ();
 sg13g2_fill_1 FILLER_29_1098 ();
 sg13g2_fill_1 FILLER_29_1126 ();
 sg13g2_fill_1 FILLER_29_1166 ();
 sg13g2_fill_2 FILLER_29_1188 ();
 sg13g2_fill_1 FILLER_29_1190 ();
 sg13g2_decap_8 FILLER_29_1227 ();
 sg13g2_fill_2 FILLER_29_1234 ();
 sg13g2_fill_2 FILLER_29_1241 ();
 sg13g2_decap_4 FILLER_29_1247 ();
 sg13g2_fill_1 FILLER_29_1251 ();
 sg13g2_fill_2 FILLER_29_1274 ();
 sg13g2_fill_1 FILLER_29_1276 ();
 sg13g2_decap_4 FILLER_29_1325 ();
 sg13g2_fill_1 FILLER_29_1329 ();
 sg13g2_fill_2 FILLER_29_1340 ();
 sg13g2_fill_2 FILLER_29_1346 ();
 sg13g2_fill_1 FILLER_29_1348 ();
 sg13g2_fill_2 FILLER_29_1375 ();
 sg13g2_fill_1 FILLER_29_1377 ();
 sg13g2_fill_2 FILLER_29_1404 ();
 sg13g2_fill_1 FILLER_29_1406 ();
 sg13g2_fill_1 FILLER_29_1472 ();
 sg13g2_fill_1 FILLER_29_1499 ();
 sg13g2_fill_2 FILLER_29_1519 ();
 sg13g2_fill_1 FILLER_29_1544 ();
 sg13g2_decap_8 FILLER_29_1571 ();
 sg13g2_decap_4 FILLER_29_1578 ();
 sg13g2_fill_1 FILLER_29_1582 ();
 sg13g2_decap_8 FILLER_29_1588 ();
 sg13g2_decap_4 FILLER_29_1595 ();
 sg13g2_fill_1 FILLER_29_1599 ();
 sg13g2_fill_2 FILLER_29_1614 ();
 sg13g2_decap_4 FILLER_29_1623 ();
 sg13g2_fill_2 FILLER_29_1632 ();
 sg13g2_fill_2 FILLER_29_1660 ();
 sg13g2_decap_8 FILLER_29_1666 ();
 sg13g2_decap_4 FILLER_29_1673 ();
 sg13g2_decap_4 FILLER_29_1687 ();
 sg13g2_fill_1 FILLER_29_1691 ();
 sg13g2_fill_1 FILLER_29_1697 ();
 sg13g2_fill_1 FILLER_29_1712 ();
 sg13g2_fill_1 FILLER_29_1781 ();
 sg13g2_fill_1 FILLER_29_1851 ();
 sg13g2_fill_2 FILLER_29_1857 ();
 sg13g2_fill_2 FILLER_29_1866 ();
 sg13g2_fill_1 FILLER_29_1892 ();
 sg13g2_fill_2 FILLER_29_1903 ();
 sg13g2_fill_2 FILLER_29_1954 ();
 sg13g2_decap_8 FILLER_29_1970 ();
 sg13g2_decap_8 FILLER_29_1977 ();
 sg13g2_decap_8 FILLER_29_1984 ();
 sg13g2_decap_8 FILLER_29_1991 ();
 sg13g2_decap_8 FILLER_29_1998 ();
 sg13g2_decap_8 FILLER_29_2005 ();
 sg13g2_decap_8 FILLER_29_2012 ();
 sg13g2_fill_1 FILLER_29_2019 ();
 sg13g2_decap_8 FILLER_29_2030 ();
 sg13g2_decap_4 FILLER_29_2037 ();
 sg13g2_fill_1 FILLER_29_2041 ();
 sg13g2_decap_4 FILLER_29_2052 ();
 sg13g2_fill_2 FILLER_29_2128 ();
 sg13g2_fill_1 FILLER_29_2130 ();
 sg13g2_fill_2 FILLER_29_2141 ();
 sg13g2_fill_2 FILLER_29_2147 ();
 sg13g2_fill_1 FILLER_29_2149 ();
 sg13g2_decap_8 FILLER_29_2195 ();
 sg13g2_decap_8 FILLER_29_2202 ();
 sg13g2_decap_8 FILLER_29_2209 ();
 sg13g2_decap_8 FILLER_29_2216 ();
 sg13g2_decap_8 FILLER_29_2223 ();
 sg13g2_decap_8 FILLER_29_2230 ();
 sg13g2_decap_8 FILLER_29_2237 ();
 sg13g2_fill_1 FILLER_29_2244 ();
 sg13g2_decap_8 FILLER_29_2255 ();
 sg13g2_decap_4 FILLER_29_2262 ();
 sg13g2_fill_1 FILLER_29_2266 ();
 sg13g2_decap_4 FILLER_29_2272 ();
 sg13g2_fill_1 FILLER_29_2276 ();
 sg13g2_decap_4 FILLER_29_2281 ();
 sg13g2_decap_4 FILLER_29_2316 ();
 sg13g2_fill_2 FILLER_29_2320 ();
 sg13g2_decap_8 FILLER_29_2342 ();
 sg13g2_fill_1 FILLER_29_2353 ();
 sg13g2_decap_8 FILLER_29_2358 ();
 sg13g2_decap_8 FILLER_29_2365 ();
 sg13g2_decap_4 FILLER_29_2372 ();
 sg13g2_fill_1 FILLER_29_2376 ();
 sg13g2_fill_2 FILLER_29_2383 ();
 sg13g2_decap_8 FILLER_29_2389 ();
 sg13g2_decap_8 FILLER_29_2396 ();
 sg13g2_decap_8 FILLER_29_2403 ();
 sg13g2_decap_8 FILLER_29_2410 ();
 sg13g2_fill_2 FILLER_29_2417 ();
 sg13g2_fill_2 FILLER_29_2425 ();
 sg13g2_decap_4 FILLER_29_2463 ();
 sg13g2_fill_1 FILLER_29_2506 ();
 sg13g2_fill_2 FILLER_29_2532 ();
 sg13g2_fill_2 FILLER_29_2556 ();
 sg13g2_decap_8 FILLER_29_2623 ();
 sg13g2_fill_2 FILLER_29_2630 ();
 sg13g2_fill_1 FILLER_29_2632 ();
 sg13g2_decap_8 FILLER_29_2637 ();
 sg13g2_fill_2 FILLER_29_2644 ();
 sg13g2_decap_8 FILLER_29_2650 ();
 sg13g2_decap_8 FILLER_29_2657 ();
 sg13g2_decap_4 FILLER_29_2664 ();
 sg13g2_fill_2 FILLER_29_2668 ();
 sg13g2_fill_2 FILLER_30_0 ();
 sg13g2_fill_2 FILLER_30_28 ();
 sg13g2_fill_1 FILLER_30_37 ();
 sg13g2_fill_2 FILLER_30_48 ();
 sg13g2_decap_4 FILLER_30_54 ();
 sg13g2_fill_1 FILLER_30_62 ();
 sg13g2_fill_1 FILLER_30_89 ();
 sg13g2_fill_1 FILLER_30_122 ();
 sg13g2_decap_8 FILLER_30_133 ();
 sg13g2_decap_8 FILLER_30_140 ();
 sg13g2_decap_8 FILLER_30_147 ();
 sg13g2_fill_2 FILLER_30_154 ();
 sg13g2_fill_1 FILLER_30_156 ();
 sg13g2_decap_8 FILLER_30_167 ();
 sg13g2_decap_4 FILLER_30_174 ();
 sg13g2_fill_2 FILLER_30_178 ();
 sg13g2_fill_2 FILLER_30_196 ();
 sg13g2_decap_8 FILLER_30_208 ();
 sg13g2_decap_4 FILLER_30_215 ();
 sg13g2_decap_4 FILLER_30_222 ();
 sg13g2_fill_1 FILLER_30_226 ();
 sg13g2_fill_2 FILLER_30_244 ();
 sg13g2_fill_1 FILLER_30_259 ();
 sg13g2_decap_4 FILLER_30_266 ();
 sg13g2_fill_2 FILLER_30_273 ();
 sg13g2_fill_1 FILLER_30_275 ();
 sg13g2_fill_2 FILLER_30_290 ();
 sg13g2_fill_2 FILLER_30_310 ();
 sg13g2_fill_1 FILLER_30_312 ();
 sg13g2_fill_2 FILLER_30_329 ();
 sg13g2_fill_2 FILLER_30_357 ();
 sg13g2_fill_2 FILLER_30_363 ();
 sg13g2_fill_1 FILLER_30_365 ();
 sg13g2_fill_1 FILLER_30_400 ();
 sg13g2_decap_4 FILLER_30_435 ();
 sg13g2_decap_8 FILLER_30_443 ();
 sg13g2_decap_4 FILLER_30_450 ();
 sg13g2_fill_2 FILLER_30_454 ();
 sg13g2_fill_1 FILLER_30_491 ();
 sg13g2_fill_1 FILLER_30_501 ();
 sg13g2_decap_4 FILLER_30_521 ();
 sg13g2_fill_2 FILLER_30_525 ();
 sg13g2_fill_2 FILLER_30_546 ();
 sg13g2_fill_1 FILLER_30_568 ();
 sg13g2_fill_1 FILLER_30_583 ();
 sg13g2_fill_2 FILLER_30_633 ();
 sg13g2_fill_1 FILLER_30_635 ();
 sg13g2_decap_8 FILLER_30_640 ();
 sg13g2_fill_1 FILLER_30_647 ();
 sg13g2_fill_2 FILLER_30_654 ();
 sg13g2_fill_1 FILLER_30_656 ();
 sg13g2_fill_1 FILLER_30_671 ();
 sg13g2_fill_1 FILLER_30_677 ();
 sg13g2_fill_1 FILLER_30_682 ();
 sg13g2_fill_2 FILLER_30_703 ();
 sg13g2_decap_8 FILLER_30_713 ();
 sg13g2_decap_4 FILLER_30_751 ();
 sg13g2_fill_1 FILLER_30_759 ();
 sg13g2_decap_4 FILLER_30_799 ();
 sg13g2_decap_4 FILLER_30_817 ();
 sg13g2_decap_8 FILLER_30_825 ();
 sg13g2_decap_8 FILLER_30_832 ();
 sg13g2_decap_8 FILLER_30_839 ();
 sg13g2_decap_8 FILLER_30_846 ();
 sg13g2_fill_1 FILLER_30_853 ();
 sg13g2_fill_2 FILLER_30_937 ();
 sg13g2_fill_1 FILLER_30_939 ();
 sg13g2_decap_8 FILLER_30_944 ();
 sg13g2_decap_8 FILLER_30_972 ();
 sg13g2_decap_8 FILLER_30_979 ();
 sg13g2_decap_8 FILLER_30_986 ();
 sg13g2_decap_8 FILLER_30_993 ();
 sg13g2_decap_4 FILLER_30_1000 ();
 sg13g2_fill_1 FILLER_30_1034 ();
 sg13g2_decap_4 FILLER_30_1061 ();
 sg13g2_fill_2 FILLER_30_1065 ();
 sg13g2_fill_1 FILLER_30_1088 ();
 sg13g2_fill_2 FILLER_30_1131 ();
 sg13g2_fill_1 FILLER_30_1143 ();
 sg13g2_fill_2 FILLER_30_1174 ();
 sg13g2_fill_1 FILLER_30_1176 ();
 sg13g2_fill_1 FILLER_30_1208 ();
 sg13g2_fill_2 FILLER_30_1235 ();
 sg13g2_fill_1 FILLER_30_1263 ();
 sg13g2_fill_2 FILLER_30_1290 ();
 sg13g2_decap_4 FILLER_30_1296 ();
 sg13g2_fill_1 FILLER_30_1300 ();
 sg13g2_decap_4 FILLER_30_1326 ();
 sg13g2_fill_1 FILLER_30_1356 ();
 sg13g2_fill_2 FILLER_30_1361 ();
 sg13g2_fill_2 FILLER_30_1367 ();
 sg13g2_fill_2 FILLER_30_1379 ();
 sg13g2_fill_1 FILLER_30_1391 ();
 sg13g2_fill_2 FILLER_30_1397 ();
 sg13g2_fill_2 FILLER_30_1414 ();
 sg13g2_fill_1 FILLER_30_1425 ();
 sg13g2_fill_1 FILLER_30_1475 ();
 sg13g2_fill_2 FILLER_30_1487 ();
 sg13g2_fill_1 FILLER_30_1517 ();
 sg13g2_decap_4 FILLER_30_1598 ();
 sg13g2_fill_2 FILLER_30_1644 ();
 sg13g2_decap_8 FILLER_30_1650 ();
 sg13g2_fill_2 FILLER_30_1661 ();
 sg13g2_fill_1 FILLER_30_1663 ();
 sg13g2_decap_4 FILLER_30_1671 ();
 sg13g2_fill_2 FILLER_30_1675 ();
 sg13g2_fill_1 FILLER_30_1686 ();
 sg13g2_fill_1 FILLER_30_1705 ();
 sg13g2_fill_2 FILLER_30_1711 ();
 sg13g2_fill_2 FILLER_30_1721 ();
 sg13g2_fill_1 FILLER_30_1723 ();
 sg13g2_fill_2 FILLER_30_1752 ();
 sg13g2_fill_1 FILLER_30_1757 ();
 sg13g2_fill_1 FILLER_30_1764 ();
 sg13g2_fill_2 FILLER_30_1770 ();
 sg13g2_fill_2 FILLER_30_1777 ();
 sg13g2_fill_2 FILLER_30_1784 ();
 sg13g2_fill_1 FILLER_30_1786 ();
 sg13g2_fill_1 FILLER_30_1837 ();
 sg13g2_decap_8 FILLER_30_1866 ();
 sg13g2_fill_2 FILLER_30_1902 ();
 sg13g2_fill_1 FILLER_30_1904 ();
 sg13g2_decap_4 FILLER_30_1940 ();
 sg13g2_fill_2 FILLER_30_1944 ();
 sg13g2_decap_4 FILLER_30_1954 ();
 sg13g2_decap_8 FILLER_30_1966 ();
 sg13g2_fill_2 FILLER_30_1973 ();
 sg13g2_fill_1 FILLER_30_1975 ();
 sg13g2_decap_8 FILLER_30_2026 ();
 sg13g2_decap_4 FILLER_30_2084 ();
 sg13g2_fill_2 FILLER_30_2088 ();
 sg13g2_decap_4 FILLER_30_2130 ();
 sg13g2_decap_8 FILLER_30_2170 ();
 sg13g2_decap_8 FILLER_30_2177 ();
 sg13g2_decap_8 FILLER_30_2184 ();
 sg13g2_decap_8 FILLER_30_2191 ();
 sg13g2_decap_8 FILLER_30_2198 ();
 sg13g2_decap_8 FILLER_30_2223 ();
 sg13g2_decap_8 FILLER_30_2230 ();
 sg13g2_decap_4 FILLER_30_2237 ();
 sg13g2_fill_2 FILLER_30_2267 ();
 sg13g2_fill_1 FILLER_30_2269 ();
 sg13g2_fill_2 FILLER_30_2322 ();
 sg13g2_fill_1 FILLER_30_2324 ();
 sg13g2_decap_4 FILLER_30_2335 ();
 sg13g2_fill_2 FILLER_30_2339 ();
 sg13g2_decap_8 FILLER_30_2367 ();
 sg13g2_decap_8 FILLER_30_2374 ();
 sg13g2_decap_8 FILLER_30_2381 ();
 sg13g2_decap_8 FILLER_30_2388 ();
 sg13g2_decap_8 FILLER_30_2395 ();
 sg13g2_decap_8 FILLER_30_2402 ();
 sg13g2_decap_4 FILLER_30_2409 ();
 sg13g2_fill_1 FILLER_30_2413 ();
 sg13g2_decap_8 FILLER_30_2428 ();
 sg13g2_fill_2 FILLER_30_2435 ();
 sg13g2_fill_1 FILLER_30_2437 ();
 sg13g2_decap_4 FILLER_30_2448 ();
 sg13g2_fill_1 FILLER_30_2506 ();
 sg13g2_decap_8 FILLER_30_2635 ();
 sg13g2_fill_2 FILLER_30_2668 ();
 sg13g2_decap_4 FILLER_31_0 ();
 sg13g2_fill_2 FILLER_31_4 ();
 sg13g2_fill_1 FILLER_31_10 ();
 sg13g2_fill_2 FILLER_31_37 ();
 sg13g2_fill_1 FILLER_31_52 ();
 sg13g2_fill_2 FILLER_31_63 ();
 sg13g2_decap_4 FILLER_31_75 ();
 sg13g2_fill_2 FILLER_31_125 ();
 sg13g2_decap_4 FILLER_31_153 ();
 sg13g2_decap_4 FILLER_31_187 ();
 sg13g2_fill_1 FILLER_31_191 ();
 sg13g2_decap_8 FILLER_31_197 ();
 sg13g2_decap_8 FILLER_31_204 ();
 sg13g2_decap_8 FILLER_31_211 ();
 sg13g2_decap_8 FILLER_31_218 ();
 sg13g2_decap_4 FILLER_31_225 ();
 sg13g2_fill_1 FILLER_31_263 ();
 sg13g2_decap_4 FILLER_31_356 ();
 sg13g2_fill_2 FILLER_31_360 ();
 sg13g2_decap_8 FILLER_31_365 ();
 sg13g2_fill_1 FILLER_31_372 ();
 sg13g2_decap_4 FILLER_31_377 ();
 sg13g2_fill_1 FILLER_31_381 ();
 sg13g2_fill_2 FILLER_31_395 ();
 sg13g2_fill_2 FILLER_31_410 ();
 sg13g2_fill_1 FILLER_31_412 ();
 sg13g2_decap_8 FILLER_31_417 ();
 sg13g2_decap_8 FILLER_31_424 ();
 sg13g2_fill_1 FILLER_31_431 ();
 sg13g2_decap_8 FILLER_31_437 ();
 sg13g2_decap_8 FILLER_31_444 ();
 sg13g2_decap_4 FILLER_31_451 ();
 sg13g2_decap_8 FILLER_31_460 ();
 sg13g2_decap_4 FILLER_31_482 ();
 sg13g2_fill_2 FILLER_31_496 ();
 sg13g2_fill_1 FILLER_31_498 ();
 sg13g2_fill_2 FILLER_31_503 ();
 sg13g2_decap_4 FILLER_31_521 ();
 sg13g2_fill_2 FILLER_31_525 ();
 sg13g2_fill_2 FILLER_31_564 ();
 sg13g2_fill_1 FILLER_31_577 ();
 sg13g2_fill_2 FILLER_31_584 ();
 sg13g2_fill_2 FILLER_31_591 ();
 sg13g2_fill_2 FILLER_31_598 ();
 sg13g2_fill_1 FILLER_31_600 ();
 sg13g2_fill_2 FILLER_31_611 ();
 sg13g2_fill_1 FILLER_31_613 ();
 sg13g2_decap_8 FILLER_31_618 ();
 sg13g2_decap_8 FILLER_31_625 ();
 sg13g2_decap_8 FILLER_31_632 ();
 sg13g2_fill_1 FILLER_31_660 ();
 sg13g2_fill_1 FILLER_31_677 ();
 sg13g2_fill_2 FILLER_31_714 ();
 sg13g2_fill_1 FILLER_31_716 ();
 sg13g2_fill_2 FILLER_31_726 ();
 sg13g2_fill_1 FILLER_31_728 ();
 sg13g2_fill_1 FILLER_31_737 ();
 sg13g2_fill_1 FILLER_31_742 ();
 sg13g2_fill_2 FILLER_31_749 ();
 sg13g2_fill_1 FILLER_31_755 ();
 sg13g2_fill_1 FILLER_31_761 ();
 sg13g2_fill_1 FILLER_31_767 ();
 sg13g2_fill_1 FILLER_31_773 ();
 sg13g2_fill_1 FILLER_31_778 ();
 sg13g2_decap_8 FILLER_31_791 ();
 sg13g2_decap_8 FILLER_31_798 ();
 sg13g2_decap_8 FILLER_31_805 ();
 sg13g2_fill_2 FILLER_31_812 ();
 sg13g2_decap_8 FILLER_31_840 ();
 sg13g2_fill_1 FILLER_31_847 ();
 sg13g2_decap_4 FILLER_31_878 ();
 sg13g2_decap_8 FILLER_31_886 ();
 sg13g2_fill_1 FILLER_31_893 ();
 sg13g2_fill_1 FILLER_31_915 ();
 sg13g2_decap_4 FILLER_31_920 ();
 sg13g2_fill_1 FILLER_31_924 ();
 sg13g2_decap_8 FILLER_31_935 ();
 sg13g2_decap_8 FILLER_31_942 ();
 sg13g2_decap_8 FILLER_31_949 ();
 sg13g2_decap_8 FILLER_31_956 ();
 sg13g2_decap_8 FILLER_31_963 ();
 sg13g2_decap_8 FILLER_31_970 ();
 sg13g2_decap_8 FILLER_31_977 ();
 sg13g2_decap_8 FILLER_31_984 ();
 sg13g2_decap_8 FILLER_31_991 ();
 sg13g2_decap_8 FILLER_31_998 ();
 sg13g2_decap_8 FILLER_31_1005 ();
 sg13g2_decap_4 FILLER_31_1021 ();
 sg13g2_fill_2 FILLER_31_1034 ();
 sg13g2_decap_8 FILLER_31_1065 ();
 sg13g2_decap_4 FILLER_31_1072 ();
 sg13g2_fill_2 FILLER_31_1100 ();
 sg13g2_fill_1 FILLER_31_1102 ();
 sg13g2_fill_2 FILLER_31_1120 ();
 sg13g2_fill_1 FILLER_31_1122 ();
 sg13g2_fill_1 FILLER_31_1126 ();
 sg13g2_decap_8 FILLER_31_1166 ();
 sg13g2_fill_2 FILLER_31_1173 ();
 sg13g2_fill_2 FILLER_31_1180 ();
 sg13g2_fill_1 FILLER_31_1182 ();
 sg13g2_fill_1 FILLER_31_1188 ();
 sg13g2_fill_1 FILLER_31_1193 ();
 sg13g2_fill_1 FILLER_31_1224 ();
 sg13g2_decap_8 FILLER_31_1229 ();
 sg13g2_decap_4 FILLER_31_1236 ();
 sg13g2_fill_1 FILLER_31_1240 ();
 sg13g2_fill_1 FILLER_31_1245 ();
 sg13g2_fill_1 FILLER_31_1272 ();
 sg13g2_fill_1 FILLER_31_1312 ();
 sg13g2_fill_2 FILLER_31_1325 ();
 sg13g2_decap_8 FILLER_31_1332 ();
 sg13g2_fill_1 FILLER_31_1343 ();
 sg13g2_decap_8 FILLER_31_1349 ();
 sg13g2_decap_8 FILLER_31_1356 ();
 sg13g2_decap_8 FILLER_31_1363 ();
 sg13g2_decap_8 FILLER_31_1370 ();
 sg13g2_decap_8 FILLER_31_1377 ();
 sg13g2_fill_1 FILLER_31_1384 ();
 sg13g2_decap_8 FILLER_31_1392 ();
 sg13g2_fill_2 FILLER_31_1399 ();
 sg13g2_fill_1 FILLER_31_1401 ();
 sg13g2_decap_8 FILLER_31_1412 ();
 sg13g2_decap_4 FILLER_31_1419 ();
 sg13g2_decap_4 FILLER_31_1428 ();
 sg13g2_fill_2 FILLER_31_1432 ();
 sg13g2_decap_4 FILLER_31_1438 ();
 sg13g2_fill_2 FILLER_31_1442 ();
 sg13g2_decap_8 FILLER_31_1448 ();
 sg13g2_decap_8 FILLER_31_1455 ();
 sg13g2_decap_8 FILLER_31_1462 ();
 sg13g2_fill_1 FILLER_31_1480 ();
 sg13g2_fill_1 FILLER_31_1549 ();
 sg13g2_fill_1 FILLER_31_1560 ();
 sg13g2_fill_1 FILLER_31_1566 ();
 sg13g2_fill_2 FILLER_31_1571 ();
 sg13g2_decap_8 FILLER_31_1583 ();
 sg13g2_decap_8 FILLER_31_1602 ();
 sg13g2_fill_1 FILLER_31_1639 ();
 sg13g2_decap_8 FILLER_31_1644 ();
 sg13g2_decap_4 FILLER_31_1651 ();
 sg13g2_fill_1 FILLER_31_1691 ();
 sg13g2_fill_1 FILLER_31_1701 ();
 sg13g2_fill_2 FILLER_31_1721 ();
 sg13g2_fill_1 FILLER_31_1723 ();
 sg13g2_decap_4 FILLER_31_1755 ();
 sg13g2_fill_1 FILLER_31_1784 ();
 sg13g2_decap_4 FILLER_31_1790 ();
 sg13g2_fill_1 FILLER_31_1794 ();
 sg13g2_fill_1 FILLER_31_1831 ();
 sg13g2_fill_1 FILLER_31_1836 ();
 sg13g2_fill_1 FILLER_31_1845 ();
 sg13g2_fill_1 FILLER_31_1850 ();
 sg13g2_fill_1 FILLER_31_1856 ();
 sg13g2_fill_2 FILLER_31_1865 ();
 sg13g2_decap_8 FILLER_31_1871 ();
 sg13g2_decap_8 FILLER_31_1878 ();
 sg13g2_fill_2 FILLER_31_1885 ();
 sg13g2_decap_4 FILLER_31_1913 ();
 sg13g2_fill_1 FILLER_31_1917 ();
 sg13g2_decap_8 FILLER_31_1941 ();
 sg13g2_decap_8 FILLER_31_1948 ();
 sg13g2_decap_4 FILLER_31_1955 ();
 sg13g2_fill_1 FILLER_31_1959 ();
 sg13g2_fill_2 FILLER_31_2035 ();
 sg13g2_fill_1 FILLER_31_2037 ();
 sg13g2_decap_8 FILLER_31_2051 ();
 sg13g2_decap_8 FILLER_31_2079 ();
 sg13g2_decap_8 FILLER_31_2086 ();
 sg13g2_fill_2 FILLER_31_2093 ();
 sg13g2_fill_1 FILLER_31_2095 ();
 sg13g2_decap_8 FILLER_31_2118 ();
 sg13g2_decap_8 FILLER_31_2125 ();
 sg13g2_fill_1 FILLER_31_2132 ();
 sg13g2_decap_4 FILLER_31_2137 ();
 sg13g2_decap_4 FILLER_31_2149 ();
 sg13g2_decap_8 FILLER_31_2163 ();
 sg13g2_decap_8 FILLER_31_2170 ();
 sg13g2_fill_2 FILLER_31_2177 ();
 sg13g2_decap_8 FILLER_31_2183 ();
 sg13g2_decap_8 FILLER_31_2190 ();
 sg13g2_fill_2 FILLER_31_2197 ();
 sg13g2_decap_4 FILLER_31_2235 ();
 sg13g2_fill_2 FILLER_31_2243 ();
 sg13g2_fill_1 FILLER_31_2245 ();
 sg13g2_fill_1 FILLER_31_2280 ();
 sg13g2_fill_1 FILLER_31_2291 ();
 sg13g2_fill_2 FILLER_31_2306 ();
 sg13g2_fill_1 FILLER_31_2318 ();
 sg13g2_decap_8 FILLER_31_2326 ();
 sg13g2_decap_8 FILLER_31_2333 ();
 sg13g2_decap_8 FILLER_31_2340 ();
 sg13g2_decap_8 FILLER_31_2347 ();
 sg13g2_fill_1 FILLER_31_2368 ();
 sg13g2_fill_2 FILLER_31_2374 ();
 sg13g2_decap_4 FILLER_31_2381 ();
 sg13g2_fill_1 FILLER_31_2385 ();
 sg13g2_fill_1 FILLER_31_2498 ();
 sg13g2_fill_2 FILLER_31_2578 ();
 sg13g2_fill_1 FILLER_31_2597 ();
 sg13g2_fill_1 FILLER_31_2638 ();
 sg13g2_fill_1 FILLER_31_2669 ();
 sg13g2_decap_8 FILLER_32_0 ();
 sg13g2_fill_2 FILLER_32_7 ();
 sg13g2_fill_2 FILLER_32_35 ();
 sg13g2_decap_4 FILLER_32_60 ();
 sg13g2_fill_2 FILLER_32_64 ();
 sg13g2_fill_1 FILLER_32_95 ();
 sg13g2_fill_2 FILLER_32_143 ();
 sg13g2_decap_4 FILLER_32_149 ();
 sg13g2_fill_1 FILLER_32_170 ();
 sg13g2_fill_2 FILLER_32_220 ();
 sg13g2_decap_8 FILLER_32_226 ();
 sg13g2_decap_8 FILLER_32_233 ();
 sg13g2_fill_2 FILLER_32_240 ();
 sg13g2_fill_2 FILLER_32_246 ();
 sg13g2_fill_1 FILLER_32_253 ();
 sg13g2_fill_1 FILLER_32_258 ();
 sg13g2_fill_2 FILLER_32_273 ();
 sg13g2_fill_2 FILLER_32_279 ();
 sg13g2_fill_1 FILLER_32_291 ();
 sg13g2_fill_1 FILLER_32_296 ();
 sg13g2_fill_1 FILLER_32_302 ();
 sg13g2_fill_1 FILLER_32_307 ();
 sg13g2_fill_2 FILLER_32_312 ();
 sg13g2_fill_1 FILLER_32_323 ();
 sg13g2_fill_1 FILLER_32_329 ();
 sg13g2_decap_8 FILLER_32_339 ();
 sg13g2_fill_1 FILLER_32_346 ();
 sg13g2_decap_8 FILLER_32_351 ();
 sg13g2_fill_1 FILLER_32_358 ();
 sg13g2_decap_8 FILLER_32_371 ();
 sg13g2_fill_2 FILLER_32_378 ();
 sg13g2_fill_1 FILLER_32_380 ();
 sg13g2_fill_2 FILLER_32_396 ();
 sg13g2_decap_4 FILLER_32_437 ();
 sg13g2_fill_1 FILLER_32_441 ();
 sg13g2_fill_1 FILLER_32_478 ();
 sg13g2_fill_1 FILLER_32_483 ();
 sg13g2_decap_4 FILLER_32_512 ();
 sg13g2_fill_2 FILLER_32_530 ();
 sg13g2_decap_8 FILLER_32_613 ();
 sg13g2_fill_2 FILLER_32_620 ();
 sg13g2_fill_1 FILLER_32_622 ();
 sg13g2_fill_1 FILLER_32_653 ();
 sg13g2_fill_2 FILLER_32_701 ();
 sg13g2_decap_4 FILLER_32_709 ();
 sg13g2_fill_2 FILLER_32_713 ();
 sg13g2_fill_2 FILLER_32_719 ();
 sg13g2_fill_2 FILLER_32_731 ();
 sg13g2_fill_1 FILLER_32_733 ();
 sg13g2_fill_2 FILLER_32_739 ();
 sg13g2_fill_1 FILLER_32_741 ();
 sg13g2_fill_2 FILLER_32_754 ();
 sg13g2_fill_1 FILLER_32_756 ();
 sg13g2_decap_4 FILLER_32_761 ();
 sg13g2_fill_2 FILLER_32_785 ();
 sg13g2_fill_1 FILLER_32_809 ();
 sg13g2_fill_1 FILLER_32_815 ();
 sg13g2_decap_4 FILLER_32_842 ();
 sg13g2_fill_1 FILLER_32_846 ();
 sg13g2_fill_2 FILLER_32_859 ();
 sg13g2_fill_2 FILLER_32_871 ();
 sg13g2_fill_1 FILLER_32_883 ();
 sg13g2_decap_8 FILLER_32_910 ();
 sg13g2_fill_2 FILLER_32_927 ();
 sg13g2_decap_8 FILLER_32_976 ();
 sg13g2_fill_2 FILLER_32_983 ();
 sg13g2_fill_1 FILLER_32_985 ();
 sg13g2_fill_2 FILLER_32_990 ();
 sg13g2_decap_4 FILLER_32_1013 ();
 sg13g2_decap_4 FILLER_32_1022 ();
 sg13g2_fill_2 FILLER_32_1035 ();
 sg13g2_fill_1 FILLER_32_1037 ();
 sg13g2_decap_8 FILLER_32_1074 ();
 sg13g2_decap_8 FILLER_32_1081 ();
 sg13g2_fill_1 FILLER_32_1093 ();
 sg13g2_fill_1 FILLER_32_1098 ();
 sg13g2_decap_4 FILLER_32_1103 ();
 sg13g2_fill_1 FILLER_32_1150 ();
 sg13g2_fill_2 FILLER_32_1155 ();
 sg13g2_fill_1 FILLER_32_1157 ();
 sg13g2_fill_1 FILLER_32_1162 ();
 sg13g2_decap_4 FILLER_32_1184 ();
 sg13g2_fill_2 FILLER_32_1188 ();
 sg13g2_fill_2 FILLER_32_1208 ();
 sg13g2_decap_8 FILLER_32_1218 ();
 sg13g2_decap_8 FILLER_32_1225 ();
 sg13g2_decap_8 FILLER_32_1232 ();
 sg13g2_decap_8 FILLER_32_1239 ();
 sg13g2_fill_1 FILLER_32_1256 ();
 sg13g2_fill_2 FILLER_32_1319 ();
 sg13g2_fill_1 FILLER_32_1321 ();
 sg13g2_fill_1 FILLER_32_1332 ();
 sg13g2_fill_2 FILLER_32_1359 ();
 sg13g2_fill_2 FILLER_32_1365 ();
 sg13g2_fill_2 FILLER_32_1372 ();
 sg13g2_fill_1 FILLER_32_1374 ();
 sg13g2_fill_2 FILLER_32_1401 ();
 sg13g2_decap_8 FILLER_32_1429 ();
 sg13g2_decap_8 FILLER_32_1436 ();
 sg13g2_decap_8 FILLER_32_1443 ();
 sg13g2_fill_1 FILLER_32_1450 ();
 sg13g2_fill_1 FILLER_32_1461 ();
 sg13g2_fill_1 FILLER_32_1475 ();
 sg13g2_fill_1 FILLER_32_1502 ();
 sg13g2_fill_1 FILLER_32_1540 ();
 sg13g2_fill_2 FILLER_32_1547 ();
 sg13g2_fill_1 FILLER_32_1573 ();
 sg13g2_fill_1 FILLER_32_1577 ();
 sg13g2_fill_1 FILLER_32_1615 ();
 sg13g2_decap_4 FILLER_32_1620 ();
 sg13g2_decap_8 FILLER_32_1675 ();
 sg13g2_decap_4 FILLER_32_1682 ();
 sg13g2_fill_1 FILLER_32_1686 ();
 sg13g2_fill_2 FILLER_32_1706 ();
 sg13g2_fill_2 FILLER_32_1724 ();
 sg13g2_fill_2 FILLER_32_1736 ();
 sg13g2_fill_1 FILLER_32_1755 ();
 sg13g2_decap_4 FILLER_32_1786 ();
 sg13g2_fill_1 FILLER_32_1790 ();
 sg13g2_decap_4 FILLER_32_1796 ();
 sg13g2_fill_2 FILLER_32_1855 ();
 sg13g2_decap_8 FILLER_32_1867 ();
 sg13g2_decap_8 FILLER_32_1874 ();
 sg13g2_decap_4 FILLER_32_1881 ();
 sg13g2_fill_2 FILLER_32_1897 ();
 sg13g2_fill_2 FILLER_32_1925 ();
 sg13g2_fill_2 FILLER_32_1961 ();
 sg13g2_fill_1 FILLER_32_1989 ();
 sg13g2_fill_2 FILLER_32_2000 ();
 sg13g2_decap_8 FILLER_32_2023 ();
 sg13g2_decap_8 FILLER_32_2030 ();
 sg13g2_decap_4 FILLER_32_2060 ();
 sg13g2_fill_1 FILLER_32_2172 ();
 sg13g2_fill_1 FILLER_32_2199 ();
 sg13g2_fill_2 FILLER_32_2226 ();
 sg13g2_decap_4 FILLER_32_2238 ();
 sg13g2_decap_8 FILLER_32_2272 ();
 sg13g2_decap_8 FILLER_32_2279 ();
 sg13g2_decap_8 FILLER_32_2286 ();
 sg13g2_fill_1 FILLER_32_2293 ();
 sg13g2_decap_8 FILLER_32_2298 ();
 sg13g2_decap_4 FILLER_32_2314 ();
 sg13g2_fill_2 FILLER_32_2318 ();
 sg13g2_fill_1 FILLER_32_2328 ();
 sg13g2_fill_1 FILLER_32_2339 ();
 sg13g2_fill_1 FILLER_32_2346 ();
 sg13g2_fill_1 FILLER_32_2351 ();
 sg13g2_fill_1 FILLER_32_2378 ();
 sg13g2_fill_1 FILLER_32_2411 ();
 sg13g2_fill_2 FILLER_32_2422 ();
 sg13g2_decap_8 FILLER_32_2457 ();
 sg13g2_fill_2 FILLER_32_2464 ();
 sg13g2_decap_8 FILLER_32_2490 ();
 sg13g2_fill_2 FILLER_32_2543 ();
 sg13g2_fill_2 FILLER_32_2640 ();
 sg13g2_fill_2 FILLER_32_2668 ();
 sg13g2_fill_2 FILLER_33_0 ();
 sg13g2_fill_2 FILLER_33_49 ();
 sg13g2_fill_1 FILLER_33_58 ();
 sg13g2_fill_2 FILLER_33_98 ();
 sg13g2_fill_2 FILLER_33_105 ();
 sg13g2_fill_2 FILLER_33_131 ();
 sg13g2_fill_2 FILLER_33_205 ();
 sg13g2_decap_4 FILLER_33_237 ();
 sg13g2_fill_1 FILLER_33_241 ();
 sg13g2_fill_2 FILLER_33_288 ();
 sg13g2_fill_1 FILLER_33_290 ();
 sg13g2_fill_2 FILLER_33_296 ();
 sg13g2_fill_2 FILLER_33_308 ();
 sg13g2_fill_1 FILLER_33_310 ();
 sg13g2_fill_1 FILLER_33_355 ();
 sg13g2_fill_2 FILLER_33_396 ();
 sg13g2_fill_1 FILLER_33_434 ();
 sg13g2_fill_1 FILLER_33_466 ();
 sg13g2_decap_4 FILLER_33_497 ();
 sg13g2_fill_1 FILLER_33_531 ();
 sg13g2_fill_1 FILLER_33_540 ();
 sg13g2_fill_1 FILLER_33_555 ();
 sg13g2_fill_2 FILLER_33_587 ();
 sg13g2_fill_1 FILLER_33_650 ();
 sg13g2_fill_2 FILLER_33_743 ();
 sg13g2_decap_4 FILLER_33_751 ();
 sg13g2_fill_1 FILLER_33_755 ();
 sg13g2_fill_2 FILLER_33_760 ();
 sg13g2_fill_2 FILLER_33_811 ();
 sg13g2_decap_8 FILLER_33_839 ();
 sg13g2_decap_4 FILLER_33_872 ();
 sg13g2_decap_8 FILLER_33_901 ();
 sg13g2_decap_4 FILLER_33_908 ();
 sg13g2_fill_2 FILLER_33_912 ();
 sg13g2_decap_8 FILLER_33_966 ();
 sg13g2_fill_2 FILLER_33_973 ();
 sg13g2_fill_1 FILLER_33_1010 ();
 sg13g2_decap_8 FILLER_33_1076 ();
 sg13g2_decap_4 FILLER_33_1083 ();
 sg13g2_fill_1 FILLER_33_1087 ();
 sg13g2_decap_8 FILLER_33_1118 ();
 sg13g2_fill_2 FILLER_33_1125 ();
 sg13g2_fill_1 FILLER_33_1127 ();
 sg13g2_fill_2 FILLER_33_1132 ();
 sg13g2_fill_1 FILLER_33_1134 ();
 sg13g2_fill_2 FILLER_33_1139 ();
 sg13g2_fill_2 FILLER_33_1146 ();
 sg13g2_decap_4 FILLER_33_1174 ();
 sg13g2_fill_1 FILLER_33_1178 ();
 sg13g2_decap_4 FILLER_33_1184 ();
 sg13g2_decap_8 FILLER_33_1193 ();
 sg13g2_decap_8 FILLER_33_1200 ();
 sg13g2_decap_4 FILLER_33_1207 ();
 sg13g2_fill_1 FILLER_33_1211 ();
 sg13g2_decap_8 FILLER_33_1216 ();
 sg13g2_fill_1 FILLER_33_1223 ();
 sg13g2_decap_8 FILLER_33_1234 ();
 sg13g2_decap_8 FILLER_33_1241 ();
 sg13g2_decap_8 FILLER_33_1248 ();
 sg13g2_decap_4 FILLER_33_1278 ();
 sg13g2_fill_1 FILLER_33_1282 ();
 sg13g2_fill_1 FILLER_33_1308 ();
 sg13g2_fill_2 FILLER_33_1318 ();
 sg13g2_fill_1 FILLER_33_1392 ();
 sg13g2_fill_2 FILLER_33_1479 ();
 sg13g2_decap_4 FILLER_33_1491 ();
 sg13g2_fill_1 FILLER_33_1498 ();
 sg13g2_fill_2 FILLER_33_1511 ();
 sg13g2_fill_1 FILLER_33_1536 ();
 sg13g2_fill_2 FILLER_33_1576 ();
 sg13g2_fill_2 FILLER_33_1583 ();
 sg13g2_decap_4 FILLER_33_1589 ();
 sg13g2_fill_2 FILLER_33_1603 ();
 sg13g2_decap_4 FILLER_33_1609 ();
 sg13g2_fill_2 FILLER_33_1635 ();
 sg13g2_fill_1 FILLER_33_1693 ();
 sg13g2_fill_1 FILLER_33_1700 ();
 sg13g2_decap_4 FILLER_33_1706 ();
 sg13g2_fill_1 FILLER_33_1710 ();
 sg13g2_fill_1 FILLER_33_1715 ();
 sg13g2_fill_2 FILLER_33_1721 ();
 sg13g2_fill_2 FILLER_33_1733 ();
 sg13g2_fill_1 FILLER_33_1735 ();
 sg13g2_fill_2 FILLER_33_1747 ();
 sg13g2_fill_2 FILLER_33_1757 ();
 sg13g2_fill_1 FILLER_33_1759 ();
 sg13g2_decap_4 FILLER_33_1796 ();
 sg13g2_fill_1 FILLER_33_1800 ();
 sg13g2_fill_2 FILLER_33_1806 ();
 sg13g2_fill_1 FILLER_33_1808 ();
 sg13g2_fill_1 FILLER_33_1820 ();
 sg13g2_fill_2 FILLER_33_1826 ();
 sg13g2_fill_1 FILLER_33_1832 ();
 sg13g2_fill_1 FILLER_33_1837 ();
 sg13g2_fill_1 FILLER_33_1843 ();
 sg13g2_fill_2 FILLER_33_1859 ();
 sg13g2_fill_1 FILLER_33_1877 ();
 sg13g2_decap_4 FILLER_33_1909 ();
 sg13g2_fill_1 FILLER_33_1913 ();
 sg13g2_fill_2 FILLER_33_1919 ();
 sg13g2_fill_1 FILLER_33_2049 ();
 sg13g2_fill_1 FILLER_33_2070 ();
 sg13g2_fill_2 FILLER_33_2136 ();
 sg13g2_fill_1 FILLER_33_2164 ();
 sg13g2_fill_2 FILLER_33_2185 ();
 sg13g2_decap_4 FILLER_33_2213 ();
 sg13g2_fill_1 FILLER_33_2238 ();
 sg13g2_fill_2 FILLER_33_2253 ();
 sg13g2_decap_8 FILLER_33_2281 ();
 sg13g2_decap_8 FILLER_33_2288 ();
 sg13g2_fill_2 FILLER_33_2295 ();
 sg13g2_fill_1 FILLER_33_2297 ();
 sg13g2_fill_1 FILLER_33_2412 ();
 sg13g2_fill_1 FILLER_33_2419 ();
 sg13g2_fill_1 FILLER_33_2426 ();
 sg13g2_fill_2 FILLER_33_2472 ();
 sg13g2_fill_2 FILLER_33_2481 ();
 sg13g2_fill_1 FILLER_33_2483 ();
 sg13g2_fill_2 FILLER_33_2510 ();
 sg13g2_fill_2 FILLER_33_2554 ();
 sg13g2_fill_1 FILLER_33_2588 ();
 sg13g2_fill_1 FILLER_33_2609 ();
 sg13g2_fill_1 FILLER_33_2632 ();
 sg13g2_decap_8 FILLER_33_2653 ();
 sg13g2_decap_8 FILLER_33_2660 ();
 sg13g2_fill_2 FILLER_33_2667 ();
 sg13g2_fill_1 FILLER_33_2669 ();
 sg13g2_decap_4 FILLER_34_0 ();
 sg13g2_fill_2 FILLER_34_4 ();
 sg13g2_decap_4 FILLER_34_11 ();
 sg13g2_fill_1 FILLER_34_15 ();
 sg13g2_fill_2 FILLER_34_30 ();
 sg13g2_fill_1 FILLER_34_50 ();
 sg13g2_fill_1 FILLER_34_58 ();
 sg13g2_fill_1 FILLER_34_85 ();
 sg13g2_fill_2 FILLER_34_172 ();
 sg13g2_decap_8 FILLER_34_183 ();
 sg13g2_decap_8 FILLER_34_190 ();
 sg13g2_fill_2 FILLER_34_197 ();
 sg13g2_decap_4 FILLER_34_203 ();
 sg13g2_fill_2 FILLER_34_211 ();
 sg13g2_decap_8 FILLER_34_221 ();
 sg13g2_decap_8 FILLER_34_228 ();
 sg13g2_fill_2 FILLER_34_235 ();
 sg13g2_fill_1 FILLER_34_241 ();
 sg13g2_fill_1 FILLER_34_281 ();
 sg13g2_fill_2 FILLER_34_317 ();
 sg13g2_decap_8 FILLER_34_323 ();
 sg13g2_fill_1 FILLER_34_330 ();
 sg13g2_decap_8 FILLER_34_335 ();
 sg13g2_decap_8 FILLER_34_342 ();
 sg13g2_decap_8 FILLER_34_349 ();
 sg13g2_fill_1 FILLER_34_356 ();
 sg13g2_fill_2 FILLER_34_396 ();
 sg13g2_fill_1 FILLER_34_398 ();
 sg13g2_fill_2 FILLER_34_408 ();
 sg13g2_fill_1 FILLER_34_429 ();
 sg13g2_fill_2 FILLER_34_446 ();
 sg13g2_decap_8 FILLER_34_461 ();
 sg13g2_fill_2 FILLER_34_468 ();
 sg13g2_fill_1 FILLER_34_470 ();
 sg13g2_decap_8 FILLER_34_475 ();
 sg13g2_fill_1 FILLER_34_482 ();
 sg13g2_decap_4 FILLER_34_530 ();
 sg13g2_fill_1 FILLER_34_534 ();
 sg13g2_fill_2 FILLER_34_555 ();
 sg13g2_fill_2 FILLER_34_569 ();
 sg13g2_fill_1 FILLER_34_579 ();
 sg13g2_fill_1 FILLER_34_608 ();
 sg13g2_fill_1 FILLER_34_617 ();
 sg13g2_fill_2 FILLER_34_631 ();
 sg13g2_fill_2 FILLER_34_674 ();
 sg13g2_fill_1 FILLER_34_681 ();
 sg13g2_fill_2 FILLER_34_698 ();
 sg13g2_decap_4 FILLER_34_705 ();
 sg13g2_decap_4 FILLER_34_713 ();
 sg13g2_fill_1 FILLER_34_717 ();
 sg13g2_fill_2 FILLER_34_724 ();
 sg13g2_fill_1 FILLER_34_726 ();
 sg13g2_fill_2 FILLER_34_731 ();
 sg13g2_decap_4 FILLER_34_736 ();
 sg13g2_fill_2 FILLER_34_740 ();
 sg13g2_decap_4 FILLER_34_746 ();
 sg13g2_decap_4 FILLER_34_754 ();
 sg13g2_fill_1 FILLER_34_768 ();
 sg13g2_fill_1 FILLER_34_800 ();
 sg13g2_fill_1 FILLER_34_806 ();
 sg13g2_decap_4 FILLER_34_816 ();
 sg13g2_fill_1 FILLER_34_820 ();
 sg13g2_fill_2 FILLER_34_825 ();
 sg13g2_fill_1 FILLER_34_827 ();
 sg13g2_decap_8 FILLER_34_832 ();
 sg13g2_decap_8 FILLER_34_839 ();
 sg13g2_fill_2 FILLER_34_846 ();
 sg13g2_decap_8 FILLER_34_888 ();
 sg13g2_decap_4 FILLER_34_895 ();
 sg13g2_fill_1 FILLER_34_899 ();
 sg13g2_fill_1 FILLER_34_936 ();
 sg13g2_fill_1 FILLER_34_951 ();
 sg13g2_fill_1 FILLER_34_978 ();
 sg13g2_fill_2 FILLER_34_1057 ();
 sg13g2_decap_4 FILLER_34_1085 ();
 sg13g2_fill_2 FILLER_34_1093 ();
 sg13g2_decap_8 FILLER_34_1130 ();
 sg13g2_decap_4 FILLER_34_1137 ();
 sg13g2_fill_1 FILLER_34_1141 ();
 sg13g2_fill_1 FILLER_34_1156 ();
 sg13g2_fill_2 FILLER_34_1187 ();
 sg13g2_decap_4 FILLER_34_1194 ();
 sg13g2_fill_1 FILLER_34_1203 ();
 sg13g2_fill_2 FILLER_34_1230 ();
 sg13g2_decap_8 FILLER_34_1258 ();
 sg13g2_decap_4 FILLER_34_1265 ();
 sg13g2_fill_1 FILLER_34_1470 ();
 sg13g2_fill_2 FILLER_34_1497 ();
 sg13g2_fill_1 FILLER_34_1520 ();
 sg13g2_decap_4 FILLER_34_1554 ();
 sg13g2_decap_8 FILLER_34_1562 ();
 sg13g2_decap_8 FILLER_34_1569 ();
 sg13g2_decap_4 FILLER_34_1576 ();
 sg13g2_fill_2 FILLER_34_1590 ();
 sg13g2_decap_4 FILLER_34_1638 ();
 sg13g2_decap_8 FILLER_34_1679 ();
 sg13g2_decap_8 FILLER_34_1686 ();
 sg13g2_decap_8 FILLER_34_1693 ();
 sg13g2_fill_2 FILLER_34_1742 ();
 sg13g2_fill_1 FILLER_34_1744 ();
 sg13g2_fill_1 FILLER_34_1782 ();
 sg13g2_fill_1 FILLER_34_1810 ();
 sg13g2_fill_2 FILLER_34_1816 ();
 sg13g2_fill_1 FILLER_34_1846 ();
 sg13g2_decap_8 FILLER_34_1852 ();
 sg13g2_decap_4 FILLER_34_1859 ();
 sg13g2_fill_1 FILLER_34_1919 ();
 sg13g2_fill_1 FILLER_34_1951 ();
 sg13g2_fill_1 FILLER_34_1962 ();
 sg13g2_fill_1 FILLER_34_1977 ();
 sg13g2_decap_8 FILLER_34_1982 ();
 sg13g2_decap_8 FILLER_34_1989 ();
 sg13g2_fill_1 FILLER_34_2006 ();
 sg13g2_fill_2 FILLER_34_2011 ();
 sg13g2_fill_1 FILLER_34_2023 ();
 sg13g2_fill_2 FILLER_34_2028 ();
 sg13g2_fill_1 FILLER_34_2034 ();
 sg13g2_decap_8 FILLER_34_2111 ();
 sg13g2_fill_1 FILLER_34_2118 ();
 sg13g2_fill_1 FILLER_34_2150 ();
 sg13g2_fill_2 FILLER_34_2211 ();
 sg13g2_fill_1 FILLER_34_2213 ();
 sg13g2_fill_2 FILLER_34_2240 ();
 sg13g2_fill_1 FILLER_34_2242 ();
 sg13g2_fill_1 FILLER_34_2331 ();
 sg13g2_fill_2 FILLER_34_2357 ();
 sg13g2_fill_1 FILLER_34_2393 ();
 sg13g2_fill_1 FILLER_34_2398 ();
 sg13g2_decap_8 FILLER_34_2455 ();
 sg13g2_decap_4 FILLER_34_2462 ();
 sg13g2_fill_2 FILLER_34_2466 ();
 sg13g2_fill_2 FILLER_34_2474 ();
 sg13g2_fill_1 FILLER_34_2502 ();
 sg13g2_fill_1 FILLER_34_2508 ();
 sg13g2_fill_1 FILLER_34_2521 ();
 sg13g2_fill_2 FILLER_34_2528 ();
 sg13g2_fill_1 FILLER_34_2541 ();
 sg13g2_fill_2 FILLER_34_2568 ();
 sg13g2_fill_1 FILLER_34_2608 ();
 sg13g2_fill_2 FILLER_34_2667 ();
 sg13g2_fill_1 FILLER_34_2669 ();
 sg13g2_fill_1 FILLER_35_0 ();
 sg13g2_fill_1 FILLER_35_93 ();
 sg13g2_fill_2 FILLER_35_103 ();
 sg13g2_fill_2 FILLER_35_118 ();
 sg13g2_fill_2 FILLER_35_141 ();
 sg13g2_fill_2 FILLER_35_150 ();
 sg13g2_fill_1 FILLER_35_161 ();
 sg13g2_decap_4 FILLER_35_166 ();
 sg13g2_fill_2 FILLER_35_170 ();
 sg13g2_decap_8 FILLER_35_177 ();
 sg13g2_decap_4 FILLER_35_184 ();
 sg13g2_fill_2 FILLER_35_192 ();
 sg13g2_decap_8 FILLER_35_214 ();
 sg13g2_fill_2 FILLER_35_221 ();
 sg13g2_fill_1 FILLER_35_223 ();
 sg13g2_fill_1 FILLER_35_265 ();
 sg13g2_fill_1 FILLER_35_271 ();
 sg13g2_fill_2 FILLER_35_277 ();
 sg13g2_fill_1 FILLER_35_284 ();
 sg13g2_fill_2 FILLER_35_304 ();
 sg13g2_decap_4 FILLER_35_310 ();
 sg13g2_fill_1 FILLER_35_314 ();
 sg13g2_decap_4 FILLER_35_324 ();
 sg13g2_fill_1 FILLER_35_328 ();
 sg13g2_fill_1 FILLER_35_355 ();
 sg13g2_fill_2 FILLER_35_391 ();
 sg13g2_fill_1 FILLER_35_415 ();
 sg13g2_fill_2 FILLER_35_426 ();
 sg13g2_fill_2 FILLER_35_436 ();
 sg13g2_fill_1 FILLER_35_438 ();
 sg13g2_decap_8 FILLER_35_444 ();
 sg13g2_fill_2 FILLER_35_451 ();
 sg13g2_fill_1 FILLER_35_453 ();
 sg13g2_fill_2 FILLER_35_493 ();
 sg13g2_fill_1 FILLER_35_495 ();
 sg13g2_fill_1 FILLER_35_500 ();
 sg13g2_decap_8 FILLER_35_527 ();
 sg13g2_fill_2 FILLER_35_539 ();
 sg13g2_fill_1 FILLER_35_562 ();
 sg13g2_decap_4 FILLER_35_598 ();
 sg13g2_fill_1 FILLER_35_602 ();
 sg13g2_fill_1 FILLER_35_616 ();
 sg13g2_fill_1 FILLER_35_648 ();
 sg13g2_fill_1 FILLER_35_679 ();
 sg13g2_fill_1 FILLER_35_684 ();
 sg13g2_fill_1 FILLER_35_690 ();
 sg13g2_fill_1 FILLER_35_695 ();
 sg13g2_fill_2 FILLER_35_701 ();
 sg13g2_fill_2 FILLER_35_760 ();
 sg13g2_decap_4 FILLER_35_774 ();
 sg13g2_fill_2 FILLER_35_778 ();
 sg13g2_decap_8 FILLER_35_784 ();
 sg13g2_fill_2 FILLER_35_791 ();
 sg13g2_fill_1 FILLER_35_793 ();
 sg13g2_decap_4 FILLER_35_798 ();
 sg13g2_decap_8 FILLER_35_830 ();
 sg13g2_decap_8 FILLER_35_837 ();
 sg13g2_decap_8 FILLER_35_844 ();
 sg13g2_decap_8 FILLER_35_851 ();
 sg13g2_fill_2 FILLER_35_858 ();
 sg13g2_fill_1 FILLER_35_860 ();
 sg13g2_decap_8 FILLER_35_901 ();
 sg13g2_fill_2 FILLER_35_956 ();
 sg13g2_fill_1 FILLER_35_958 ();
 sg13g2_decap_4 FILLER_35_963 ();
 sg13g2_fill_1 FILLER_35_967 ();
 sg13g2_decap_8 FILLER_35_1007 ();
 sg13g2_fill_2 FILLER_35_1014 ();
 sg13g2_fill_1 FILLER_35_1016 ();
 sg13g2_fill_1 FILLER_35_1043 ();
 sg13g2_fill_1 FILLER_35_1074 ();
 sg13g2_fill_2 FILLER_35_1110 ();
 sg13g2_decap_8 FILLER_35_1173 ();
 sg13g2_decap_8 FILLER_35_1180 ();
 sg13g2_decap_8 FILLER_35_1192 ();
 sg13g2_fill_2 FILLER_35_1199 ();
 sg13g2_fill_1 FILLER_35_1201 ();
 sg13g2_fill_2 FILLER_35_1256 ();
 sg13g2_fill_1 FILLER_35_1258 ();
 sg13g2_fill_1 FILLER_35_1274 ();
 sg13g2_decap_8 FILLER_35_1301 ();
 sg13g2_fill_1 FILLER_35_1318 ();
 sg13g2_fill_2 FILLER_35_1355 ();
 sg13g2_fill_1 FILLER_35_1357 ();
 sg13g2_fill_1 FILLER_35_1384 ();
 sg13g2_fill_2 FILLER_35_1403 ();
 sg13g2_decap_8 FILLER_35_1460 ();
 sg13g2_decap_4 FILLER_35_1467 ();
 sg13g2_fill_2 FILLER_35_1471 ();
 sg13g2_fill_1 FILLER_35_1477 ();
 sg13g2_decap_8 FILLER_35_1481 ();
 sg13g2_decap_4 FILLER_35_1488 ();
 sg13g2_fill_2 FILLER_35_1492 ();
 sg13g2_fill_2 FILLER_35_1532 ();
 sg13g2_fill_2 FILLER_35_1543 ();
 sg13g2_decap_8 FILLER_35_1571 ();
 sg13g2_fill_1 FILLER_35_1578 ();
 sg13g2_fill_1 FILLER_35_1612 ();
 sg13g2_fill_1 FILLER_35_1616 ();
 sg13g2_fill_1 FILLER_35_1624 ();
 sg13g2_fill_2 FILLER_35_1659 ();
 sg13g2_fill_1 FILLER_35_1661 ();
 sg13g2_fill_2 FILLER_35_1669 ();
 sg13g2_fill_1 FILLER_35_1671 ();
 sg13g2_decap_8 FILLER_35_1679 ();
 sg13g2_fill_2 FILLER_35_1686 ();
 sg13g2_fill_1 FILLER_35_1688 ();
 sg13g2_fill_1 FILLER_35_1699 ();
 sg13g2_fill_1 FILLER_35_1704 ();
 sg13g2_fill_1 FILLER_35_1710 ();
 sg13g2_fill_1 FILLER_35_1715 ();
 sg13g2_fill_2 FILLER_35_1722 ();
 sg13g2_fill_1 FILLER_35_1729 ();
 sg13g2_fill_1 FILLER_35_1736 ();
 sg13g2_fill_1 FILLER_35_1742 ();
 sg13g2_fill_1 FILLER_35_1762 ();
 sg13g2_fill_2 FILLER_35_1771 ();
 sg13g2_fill_1 FILLER_35_1783 ();
 sg13g2_fill_1 FILLER_35_1791 ();
 sg13g2_decap_4 FILLER_35_1796 ();
 sg13g2_fill_2 FILLER_35_1805 ();
 sg13g2_fill_2 FILLER_35_1812 ();
 sg13g2_fill_2 FILLER_35_1819 ();
 sg13g2_decap_4 FILLER_35_1840 ();
 sg13g2_fill_1 FILLER_35_1858 ();
 sg13g2_decap_8 FILLER_35_1863 ();
 sg13g2_decap_4 FILLER_35_1870 ();
 sg13g2_fill_1 FILLER_35_1878 ();
 sg13g2_fill_2 FILLER_35_1940 ();
 sg13g2_fill_2 FILLER_35_1966 ();
 sg13g2_fill_1 FILLER_35_1978 ();
 sg13g2_decap_8 FILLER_35_2021 ();
 sg13g2_decap_4 FILLER_35_2028 ();
 sg13g2_decap_8 FILLER_35_2062 ();
 sg13g2_decap_4 FILLER_35_2069 ();
 sg13g2_fill_2 FILLER_35_2073 ();
 sg13g2_decap_8 FILLER_35_2096 ();
 sg13g2_decap_8 FILLER_35_2103 ();
 sg13g2_decap_8 FILLER_35_2110 ();
 sg13g2_fill_1 FILLER_35_2117 ();
 sg13g2_decap_8 FILLER_35_2139 ();
 sg13g2_decap_8 FILLER_35_2146 ();
 sg13g2_fill_2 FILLER_35_2157 ();
 sg13g2_decap_8 FILLER_35_2205 ();
 sg13g2_decap_4 FILLER_35_2226 ();
 sg13g2_fill_2 FILLER_35_2261 ();
 sg13g2_fill_1 FILLER_35_2263 ();
 sg13g2_decap_8 FILLER_35_2268 ();
 sg13g2_fill_1 FILLER_35_2305 ();
 sg13g2_fill_2 FILLER_35_2342 ();
 sg13g2_fill_1 FILLER_35_2344 ();
 sg13g2_decap_4 FILLER_35_2358 ();
 sg13g2_fill_2 FILLER_35_2368 ();
 sg13g2_decap_4 FILLER_35_2374 ();
 sg13g2_decap_4 FILLER_35_2384 ();
 sg13g2_fill_2 FILLER_35_2393 ();
 sg13g2_fill_1 FILLER_35_2395 ();
 sg13g2_decap_8 FILLER_35_2407 ();
 sg13g2_fill_2 FILLER_35_2414 ();
 sg13g2_fill_1 FILLER_35_2416 ();
 sg13g2_fill_1 FILLER_35_2469 ();
 sg13g2_fill_1 FILLER_35_2529 ();
 sg13g2_fill_2 FILLER_35_2572 ();
 sg13g2_fill_1 FILLER_35_2633 ();
 sg13g2_decap_4 FILLER_35_2644 ();
 sg13g2_decap_8 FILLER_35_2656 ();
 sg13g2_decap_8 FILLER_35_2663 ();
 sg13g2_fill_2 FILLER_36_0 ();
 sg13g2_fill_1 FILLER_36_31 ();
 sg13g2_fill_1 FILLER_36_47 ();
 sg13g2_decap_8 FILLER_36_84 ();
 sg13g2_fill_2 FILLER_36_91 ();
 sg13g2_fill_1 FILLER_36_93 ();
 sg13g2_fill_2 FILLER_36_99 ();
 sg13g2_fill_1 FILLER_36_113 ();
 sg13g2_fill_1 FILLER_36_127 ();
 sg13g2_fill_1 FILLER_36_133 ();
 sg13g2_fill_2 FILLER_36_167 ();
 sg13g2_fill_2 FILLER_36_174 ();
 sg13g2_fill_1 FILLER_36_176 ();
 sg13g2_decap_4 FILLER_36_207 ();
 sg13g2_decap_4 FILLER_36_219 ();
 sg13g2_fill_2 FILLER_36_276 ();
 sg13g2_fill_1 FILLER_36_278 ();
 sg13g2_decap_8 FILLER_36_307 ();
 sg13g2_decap_4 FILLER_36_314 ();
 sg13g2_fill_1 FILLER_36_318 ();
 sg13g2_decap_4 FILLER_36_323 ();
 sg13g2_decap_8 FILLER_36_341 ();
 sg13g2_decap_8 FILLER_36_348 ();
 sg13g2_fill_2 FILLER_36_377 ();
 sg13g2_fill_2 FILLER_36_430 ();
 sg13g2_decap_4 FILLER_36_442 ();
 sg13g2_fill_1 FILLER_36_446 ();
 sg13g2_decap_4 FILLER_36_456 ();
 sg13g2_fill_2 FILLER_36_460 ();
 sg13g2_decap_8 FILLER_36_480 ();
 sg13g2_decap_8 FILLER_36_487 ();
 sg13g2_decap_8 FILLER_36_494 ();
 sg13g2_decap_4 FILLER_36_501 ();
 sg13g2_fill_2 FILLER_36_505 ();
 sg13g2_fill_1 FILLER_36_511 ();
 sg13g2_decap_4 FILLER_36_522 ();
 sg13g2_fill_2 FILLER_36_594 ();
 sg13g2_decap_8 FILLER_36_601 ();
 sg13g2_decap_8 FILLER_36_608 ();
 sg13g2_decap_4 FILLER_36_615 ();
 sg13g2_fill_1 FILLER_36_623 ();
 sg13g2_fill_1 FILLER_36_639 ();
 sg13g2_fill_1 FILLER_36_644 ();
 sg13g2_fill_1 FILLER_36_676 ();
 sg13g2_fill_2 FILLER_36_681 ();
 sg13g2_fill_1 FILLER_36_683 ();
 sg13g2_fill_2 FILLER_36_719 ();
 sg13g2_fill_1 FILLER_36_721 ();
 sg13g2_decap_8 FILLER_36_728 ();
 sg13g2_fill_1 FILLER_36_739 ();
 sg13g2_fill_2 FILLER_36_748 ();
 sg13g2_fill_1 FILLER_36_756 ();
 sg13g2_decap_8 FILLER_36_762 ();
 sg13g2_fill_1 FILLER_36_769 ();
 sg13g2_decap_8 FILLER_36_775 ();
 sg13g2_fill_1 FILLER_36_782 ();
 sg13g2_decap_4 FILLER_36_788 ();
 sg13g2_fill_1 FILLER_36_807 ();
 sg13g2_fill_1 FILLER_36_813 ();
 sg13g2_decap_4 FILLER_36_819 ();
 sg13g2_fill_2 FILLER_36_823 ();
 sg13g2_decap_8 FILLER_36_855 ();
 sg13g2_fill_1 FILLER_36_862 ();
 sg13g2_fill_1 FILLER_36_867 ();
 sg13g2_fill_1 FILLER_36_872 ();
 sg13g2_fill_1 FILLER_36_883 ();
 sg13g2_fill_1 FILLER_36_894 ();
 sg13g2_fill_1 FILLER_36_921 ();
 sg13g2_fill_2 FILLER_36_926 ();
 sg13g2_decap_8 FILLER_36_958 ();
 sg13g2_decap_8 FILLER_36_965 ();
 sg13g2_decap_8 FILLER_36_972 ();
 sg13g2_fill_2 FILLER_36_979 ();
 sg13g2_fill_1 FILLER_36_981 ();
 sg13g2_fill_2 FILLER_36_1000 ();
 sg13g2_fill_1 FILLER_36_1002 ();
 sg13g2_decap_8 FILLER_36_1007 ();
 sg13g2_decap_8 FILLER_36_1014 ();
 sg13g2_fill_2 FILLER_36_1021 ();
 sg13g2_fill_2 FILLER_36_1036 ();
 sg13g2_fill_1 FILLER_36_1038 ();
 sg13g2_fill_2 FILLER_36_1047 ();
 sg13g2_fill_2 FILLER_36_1054 ();
 sg13g2_fill_2 FILLER_36_1060 ();
 sg13g2_fill_1 FILLER_36_1135 ();
 sg13g2_fill_2 FILLER_36_1140 ();
 sg13g2_decap_4 FILLER_36_1147 ();
 sg13g2_decap_4 FILLER_36_1155 ();
 sg13g2_fill_1 FILLER_36_1159 ();
 sg13g2_decap_8 FILLER_36_1164 ();
 sg13g2_decap_4 FILLER_36_1171 ();
 sg13g2_fill_2 FILLER_36_1225 ();
 sg13g2_fill_2 FILLER_36_1231 ();
 sg13g2_fill_1 FILLER_36_1268 ();
 sg13g2_decap_8 FILLER_36_1290 ();
 sg13g2_fill_2 FILLER_36_1297 ();
 sg13g2_fill_2 FILLER_36_1309 ();
 sg13g2_fill_1 FILLER_36_1311 ();
 sg13g2_fill_1 FILLER_36_1332 ();
 sg13g2_fill_2 FILLER_36_1337 ();
 sg13g2_fill_1 FILLER_36_1339 ();
 sg13g2_fill_1 FILLER_36_1426 ();
 sg13g2_fill_1 FILLER_36_1454 ();
 sg13g2_fill_2 FILLER_36_1570 ();
 sg13g2_decap_8 FILLER_36_1588 ();
 sg13g2_fill_1 FILLER_36_1595 ();
 sg13g2_fill_1 FILLER_36_1620 ();
 sg13g2_decap_8 FILLER_36_1651 ();
 sg13g2_decap_8 FILLER_36_1658 ();
 sg13g2_decap_8 FILLER_36_1665 ();
 sg13g2_fill_1 FILLER_36_1672 ();
 sg13g2_fill_1 FILLER_36_1690 ();
 sg13g2_fill_1 FILLER_36_1709 ();
 sg13g2_fill_2 FILLER_36_1722 ();
 sg13g2_fill_1 FILLER_36_1742 ();
 sg13g2_fill_1 FILLER_36_1756 ();
 sg13g2_fill_1 FILLER_36_1765 ();
 sg13g2_fill_2 FILLER_36_1782 ();
 sg13g2_fill_2 FILLER_36_1788 ();
 sg13g2_fill_1 FILLER_36_1790 ();
 sg13g2_fill_2 FILLER_36_1811 ();
 sg13g2_fill_1 FILLER_36_1813 ();
 sg13g2_fill_1 FILLER_36_1834 ();
 sg13g2_fill_2 FILLER_36_1844 ();
 sg13g2_fill_1 FILLER_36_1846 ();
 sg13g2_fill_2 FILLER_36_1857 ();
 sg13g2_fill_1 FILLER_36_1859 ();
 sg13g2_decap_8 FILLER_36_1870 ();
 sg13g2_fill_1 FILLER_36_1877 ();
 sg13g2_fill_1 FILLER_36_1890 ();
 sg13g2_fill_1 FILLER_36_1917 ();
 sg13g2_fill_2 FILLER_36_1957 ();
 sg13g2_fill_2 FILLER_36_1963 ();
 sg13g2_decap_4 FILLER_36_1991 ();
 sg13g2_decap_8 FILLER_36_2021 ();
 sg13g2_decap_8 FILLER_36_2028 ();
 sg13g2_decap_4 FILLER_36_2035 ();
 sg13g2_fill_2 FILLER_36_2039 ();
 sg13g2_fill_1 FILLER_36_2067 ();
 sg13g2_decap_8 FILLER_36_2109 ();
 sg13g2_decap_8 FILLER_36_2116 ();
 sg13g2_decap_8 FILLER_36_2123 ();
 sg13g2_decap_8 FILLER_36_2130 ();
 sg13g2_fill_2 FILLER_36_2137 ();
 sg13g2_fill_2 FILLER_36_2175 ();
 sg13g2_fill_1 FILLER_36_2181 ();
 sg13g2_fill_1 FILLER_36_2208 ();
 sg13g2_fill_1 FILLER_36_2235 ();
 sg13g2_fill_1 FILLER_36_2257 ();
 sg13g2_decap_8 FILLER_36_2271 ();
 sg13g2_fill_2 FILLER_36_2278 ();
 sg13g2_fill_2 FILLER_36_2314 ();
 sg13g2_decap_8 FILLER_36_2321 ();
 sg13g2_fill_1 FILLER_36_2328 ();
 sg13g2_decap_4 FILLER_36_2355 ();
 sg13g2_fill_1 FILLER_36_2359 ();
 sg13g2_decap_8 FILLER_36_2455 ();
 sg13g2_fill_1 FILLER_36_2462 ();
 sg13g2_decap_8 FILLER_36_2497 ();
 sg13g2_fill_2 FILLER_36_2504 ();
 sg13g2_fill_1 FILLER_36_2565 ();
 sg13g2_fill_2 FILLER_36_2631 ();
 sg13g2_fill_1 FILLER_36_2643 ();
 sg13g2_decap_4 FILLER_37_0 ();
 sg13g2_fill_1 FILLER_37_4 ();
 sg13g2_fill_2 FILLER_37_62 ();
 sg13g2_decap_8 FILLER_37_88 ();
 sg13g2_fill_2 FILLER_37_95 ();
 sg13g2_fill_1 FILLER_37_97 ();
 sg13g2_fill_1 FILLER_37_123 ();
 sg13g2_fill_1 FILLER_37_130 ();
 sg13g2_fill_2 FILLER_37_139 ();
 sg13g2_fill_1 FILLER_37_141 ();
 sg13g2_fill_1 FILLER_37_147 ();
 sg13g2_fill_1 FILLER_37_152 ();
 sg13g2_fill_1 FILLER_37_158 ();
 sg13g2_decap_4 FILLER_37_164 ();
 sg13g2_fill_2 FILLER_37_168 ();
 sg13g2_fill_2 FILLER_37_210 ();
 sg13g2_fill_2 FILLER_37_266 ();
 sg13g2_fill_1 FILLER_37_338 ();
 sg13g2_fill_2 FILLER_37_349 ();
 sg13g2_fill_1 FILLER_37_368 ();
 sg13g2_fill_2 FILLER_37_434 ();
 sg13g2_fill_1 FILLER_37_436 ();
 sg13g2_fill_1 FILLER_37_441 ();
 sg13g2_fill_1 FILLER_37_473 ();
 sg13g2_decap_4 FILLER_37_488 ();
 sg13g2_decap_8 FILLER_37_496 ();
 sg13g2_fill_1 FILLER_37_503 ();
 sg13g2_fill_1 FILLER_37_532 ();
 sg13g2_fill_1 FILLER_37_561 ();
 sg13g2_fill_1 FILLER_37_567 ();
 sg13g2_decap_4 FILLER_37_598 ();
 sg13g2_fill_2 FILLER_37_602 ();
 sg13g2_fill_1 FILLER_37_648 ();
 sg13g2_fill_2 FILLER_37_723 ();
 sg13g2_decap_8 FILLER_37_849 ();
 sg13g2_decap_8 FILLER_37_882 ();
 sg13g2_fill_2 FILLER_37_889 ();
 sg13g2_fill_1 FILLER_37_891 ();
 sg13g2_fill_1 FILLER_37_912 ();
 sg13g2_fill_1 FILLER_37_923 ();
 sg13g2_fill_1 FILLER_37_934 ();
 sg13g2_decap_8 FILLER_37_949 ();
 sg13g2_decap_8 FILLER_37_956 ();
 sg13g2_fill_2 FILLER_37_963 ();
 sg13g2_decap_8 FILLER_37_1004 ();
 sg13g2_decap_4 FILLER_37_1011 ();
 sg13g2_fill_1 FILLER_37_1020 ();
 sg13g2_decap_4 FILLER_37_1025 ();
 sg13g2_fill_1 FILLER_37_1029 ();
 sg13g2_decap_4 FILLER_37_1064 ();
 sg13g2_fill_2 FILLER_37_1068 ();
 sg13g2_fill_2 FILLER_37_1096 ();
 sg13g2_fill_1 FILLER_37_1110 ();
 sg13g2_fill_2 FILLER_37_1116 ();
 sg13g2_decap_4 FILLER_37_1122 ();
 sg13g2_fill_2 FILLER_37_1126 ();
 sg13g2_decap_8 FILLER_37_1132 ();
 sg13g2_decap_4 FILLER_37_1139 ();
 sg13g2_fill_1 FILLER_37_1147 ();
 sg13g2_decap_4 FILLER_37_1152 ();
 sg13g2_decap_8 FILLER_37_1177 ();
 sg13g2_decap_8 FILLER_37_1184 ();
 sg13g2_decap_4 FILLER_37_1195 ();
 sg13g2_decap_4 FILLER_37_1203 ();
 sg13g2_decap_4 FILLER_37_1221 ();
 sg13g2_decap_8 FILLER_37_1256 ();
 sg13g2_decap_8 FILLER_37_1312 ();
 sg13g2_decap_8 FILLER_37_1326 ();
 sg13g2_decap_8 FILLER_37_1333 ();
 sg13g2_decap_8 FILLER_37_1340 ();
 sg13g2_decap_4 FILLER_37_1347 ();
 sg13g2_fill_1 FILLER_37_1351 ();
 sg13g2_fill_1 FILLER_37_1416 ();
 sg13g2_decap_8 FILLER_37_1426 ();
 sg13g2_decap_8 FILLER_37_1465 ();
 sg13g2_decap_8 FILLER_37_1472 ();
 sg13g2_decap_8 FILLER_37_1479 ();
 sg13g2_decap_4 FILLER_37_1486 ();
 sg13g2_fill_2 FILLER_37_1490 ();
 sg13g2_fill_2 FILLER_37_1525 ();
 sg13g2_fill_1 FILLER_37_1560 ();
 sg13g2_fill_1 FILLER_37_1565 ();
 sg13g2_fill_2 FILLER_37_1569 ();
 sg13g2_fill_1 FILLER_37_1615 ();
 sg13g2_fill_2 FILLER_37_1624 ();
 sg13g2_decap_4 FILLER_37_1649 ();
 sg13g2_decap_8 FILLER_37_1660 ();
 sg13g2_decap_4 FILLER_37_1667 ();
 sg13g2_fill_2 FILLER_37_1671 ();
 sg13g2_decap_4 FILLER_37_1677 ();
 sg13g2_fill_1 FILLER_37_1681 ();
 sg13g2_fill_1 FILLER_37_1702 ();
 sg13g2_decap_4 FILLER_37_1708 ();
 sg13g2_fill_1 FILLER_37_1712 ();
 sg13g2_fill_1 FILLER_37_1719 ();
 sg13g2_fill_1 FILLER_37_1769 ();
 sg13g2_fill_1 FILLER_37_1783 ();
 sg13g2_fill_1 FILLER_37_1807 ();
 sg13g2_fill_2 FILLER_37_1815 ();
 sg13g2_fill_1 FILLER_37_1821 ();
 sg13g2_fill_1 FILLER_37_1830 ();
 sg13g2_fill_1 FILLER_37_1841 ();
 sg13g2_fill_1 FILLER_37_1846 ();
 sg13g2_fill_1 FILLER_37_1857 ();
 sg13g2_fill_2 FILLER_37_1862 ();
 sg13g2_decap_8 FILLER_37_1869 ();
 sg13g2_decap_4 FILLER_37_1876 ();
 sg13g2_fill_1 FILLER_37_1919 ();
 sg13g2_decap_4 FILLER_37_1982 ();
 sg13g2_fill_2 FILLER_37_1986 ();
 sg13g2_decap_4 FILLER_37_1998 ();
 sg13g2_decap_8 FILLER_37_2006 ();
 sg13g2_decap_4 FILLER_37_2018 ();
 sg13g2_decap_8 FILLER_37_2030 ();
 sg13g2_fill_1 FILLER_37_2037 ();
 sg13g2_decap_8 FILLER_37_2104 ();
 sg13g2_decap_8 FILLER_37_2111 ();
 sg13g2_decap_8 FILLER_37_2118 ();
 sg13g2_decap_8 FILLER_37_2125 ();
 sg13g2_fill_2 FILLER_37_2158 ();
 sg13g2_fill_1 FILLER_37_2170 ();
 sg13g2_decap_8 FILLER_37_2201 ();
 sg13g2_decap_4 FILLER_37_2208 ();
 sg13g2_fill_2 FILLER_37_2248 ();
 sg13g2_decap_8 FILLER_37_2284 ();
 sg13g2_decap_8 FILLER_37_2291 ();
 sg13g2_decap_8 FILLER_37_2298 ();
 sg13g2_decap_8 FILLER_37_2305 ();
 sg13g2_decap_8 FILLER_37_2312 ();
 sg13g2_fill_2 FILLER_37_2398 ();
 sg13g2_fill_1 FILLER_37_2400 ();
 sg13g2_fill_1 FILLER_37_2411 ();
 sg13g2_fill_2 FILLER_37_2454 ();
 sg13g2_fill_1 FILLER_37_2456 ();
 sg13g2_fill_2 FILLER_37_2493 ();
 sg13g2_fill_2 FILLER_37_2507 ();
 sg13g2_fill_1 FILLER_37_2509 ();
 sg13g2_fill_2 FILLER_37_2520 ();
 sg13g2_fill_2 FILLER_37_2566 ();
 sg13g2_fill_2 FILLER_37_2593 ();
 sg13g2_fill_2 FILLER_37_2618 ();
 sg13g2_decap_4 FILLER_37_2640 ();
 sg13g2_decap_4 FILLER_38_0 ();
 sg13g2_fill_1 FILLER_38_4 ();
 sg13g2_fill_2 FILLER_38_12 ();
 sg13g2_decap_4 FILLER_38_58 ();
 sg13g2_fill_2 FILLER_38_62 ();
 sg13g2_fill_1 FILLER_38_68 ();
 sg13g2_fill_1 FILLER_38_95 ();
 sg13g2_fill_1 FILLER_38_100 ();
 sg13g2_fill_1 FILLER_38_106 ();
 sg13g2_decap_4 FILLER_38_111 ();
 sg13g2_fill_2 FILLER_38_120 ();
 sg13g2_decap_4 FILLER_38_141 ();
 sg13g2_fill_1 FILLER_38_150 ();
 sg13g2_fill_2 FILLER_38_202 ();
 sg13g2_fill_1 FILLER_38_208 ();
 sg13g2_fill_2 FILLER_38_229 ();
 sg13g2_fill_2 FILLER_38_252 ();
 sg13g2_fill_1 FILLER_38_311 ();
 sg13g2_fill_2 FILLER_38_381 ();
 sg13g2_fill_1 FILLER_38_394 ();
 sg13g2_fill_1 FILLER_38_400 ();
 sg13g2_fill_2 FILLER_38_427 ();
 sg13g2_fill_1 FILLER_38_429 ();
 sg13g2_fill_1 FILLER_38_440 ();
 sg13g2_fill_2 FILLER_38_497 ();
 sg13g2_fill_1 FILLER_38_503 ();
 sg13g2_fill_1 FILLER_38_530 ();
 sg13g2_fill_1 FILLER_38_536 ();
 sg13g2_fill_2 FILLER_38_557 ();
 sg13g2_fill_1 FILLER_38_579 ();
 sg13g2_fill_2 FILLER_38_606 ();
 sg13g2_fill_1 FILLER_38_624 ();
 sg13g2_fill_2 FILLER_38_628 ();
 sg13g2_fill_2 FILLER_38_637 ();
 sg13g2_fill_1 FILLER_38_647 ();
 sg13g2_decap_4 FILLER_38_657 ();
 sg13g2_fill_2 FILLER_38_665 ();
 sg13g2_decap_4 FILLER_38_677 ();
 sg13g2_decap_4 FILLER_38_689 ();
 sg13g2_fill_2 FILLER_38_697 ();
 sg13g2_fill_1 FILLER_38_699 ();
 sg13g2_fill_1 FILLER_38_704 ();
 sg13g2_fill_2 FILLER_38_710 ();
 sg13g2_fill_1 FILLER_38_712 ();
 sg13g2_fill_2 FILLER_38_732 ();
 sg13g2_fill_1 FILLER_38_774 ();
 sg13g2_decap_8 FILLER_38_779 ();
 sg13g2_decap_8 FILLER_38_786 ();
 sg13g2_fill_1 FILLER_38_793 ();
 sg13g2_fill_1 FILLER_38_799 ();
 sg13g2_fill_1 FILLER_38_830 ();
 sg13g2_decap_8 FILLER_38_845 ();
 sg13g2_fill_2 FILLER_38_878 ();
 sg13g2_fill_1 FILLER_38_884 ();
 sg13g2_fill_1 FILLER_38_914 ();
 sg13g2_decap_4 FILLER_38_941 ();
 sg13g2_decap_4 FILLER_38_966 ();
 sg13g2_decap_4 FILLER_38_1009 ();
 sg13g2_fill_1 FILLER_38_1013 ();
 sg13g2_fill_2 FILLER_38_1040 ();
 sg13g2_fill_1 FILLER_38_1042 ();
 sg13g2_decap_8 FILLER_38_1056 ();
 sg13g2_decap_8 FILLER_38_1063 ();
 sg13g2_decap_8 FILLER_38_1070 ();
 sg13g2_decap_4 FILLER_38_1077 ();
 sg13g2_decap_8 FILLER_38_1108 ();
 sg13g2_decap_8 FILLER_38_1177 ();
 sg13g2_fill_2 FILLER_38_1184 ();
 sg13g2_fill_1 FILLER_38_1186 ();
 sg13g2_decap_4 FILLER_38_1223 ();
 sg13g2_fill_1 FILLER_38_1227 ();
 sg13g2_decap_8 FILLER_38_1274 ();
 sg13g2_fill_1 FILLER_38_1295 ();
 sg13g2_decap_8 FILLER_38_1325 ();
 sg13g2_fill_2 FILLER_38_1332 ();
 sg13g2_fill_2 FILLER_38_1368 ();
 sg13g2_fill_1 FILLER_38_1370 ();
 sg13g2_decap_4 FILLER_38_1407 ();
 sg13g2_fill_2 FILLER_38_1437 ();
 sg13g2_fill_1 FILLER_38_1473 ();
 sg13g2_fill_2 FILLER_38_1478 ();
 sg13g2_decap_4 FILLER_38_1483 ();
 sg13g2_fill_1 FILLER_38_1487 ();
 sg13g2_decap_8 FILLER_38_1502 ();
 sg13g2_fill_1 FILLER_38_1509 ();
 sg13g2_fill_2 FILLER_38_1536 ();
 sg13g2_fill_1 FILLER_38_1538 ();
 sg13g2_fill_2 FILLER_38_1543 ();
 sg13g2_fill_2 FILLER_38_1554 ();
 sg13g2_fill_1 FILLER_38_1565 ();
 sg13g2_fill_1 FILLER_38_1611 ();
 sg13g2_fill_2 FILLER_38_1650 ();
 sg13g2_fill_1 FILLER_38_1697 ();
 sg13g2_fill_2 FILLER_38_1702 ();
 sg13g2_fill_2 FILLER_38_1708 ();
 sg13g2_fill_1 FILLER_38_1710 ();
 sg13g2_fill_2 FILLER_38_1730 ();
 sg13g2_fill_1 FILLER_38_1732 ();
 sg13g2_fill_2 FILLER_38_1743 ();
 sg13g2_fill_1 FILLER_38_1760 ();
 sg13g2_fill_1 FILLER_38_1766 ();
 sg13g2_fill_2 FILLER_38_1772 ();
 sg13g2_fill_1 FILLER_38_1774 ();
 sg13g2_fill_2 FILLER_38_1785 ();
 sg13g2_fill_2 FILLER_38_1817 ();
 sg13g2_decap_4 FILLER_38_1829 ();
 sg13g2_fill_1 FILLER_38_1852 ();
 sg13g2_fill_1 FILLER_38_1864 ();
 sg13g2_decap_8 FILLER_38_1871 ();
 sg13g2_fill_1 FILLER_38_1885 ();
 sg13g2_fill_1 FILLER_38_1893 ();
 sg13g2_fill_2 FILLER_38_1898 ();
 sg13g2_decap_4 FILLER_38_1904 ();
 sg13g2_fill_2 FILLER_38_1913 ();
 sg13g2_fill_1 FILLER_38_1915 ();
 sg13g2_fill_1 FILLER_38_1951 ();
 sg13g2_fill_2 FILLER_38_2008 ();
 sg13g2_fill_1 FILLER_38_2010 ();
 sg13g2_decap_8 FILLER_38_2016 ();
 sg13g2_decap_8 FILLER_38_2023 ();
 sg13g2_decap_4 FILLER_38_2030 ();
 sg13g2_fill_2 FILLER_38_2052 ();
 sg13g2_fill_2 FILLER_38_2103 ();
 sg13g2_fill_1 FILLER_38_2105 ();
 sg13g2_fill_1 FILLER_38_2110 ();
 sg13g2_decap_4 FILLER_38_2121 ();
 sg13g2_fill_1 FILLER_38_2166 ();
 sg13g2_decap_8 FILLER_38_2205 ();
 sg13g2_decap_4 FILLER_38_2226 ();
 sg13g2_fill_1 FILLER_38_2230 ();
 sg13g2_fill_1 FILLER_38_2235 ();
 sg13g2_fill_1 FILLER_38_2266 ();
 sg13g2_decap_4 FILLER_38_2271 ();
 sg13g2_fill_2 FILLER_38_2275 ();
 sg13g2_decap_4 FILLER_38_2348 ();
 sg13g2_fill_2 FILLER_38_2352 ();
 sg13g2_fill_1 FILLER_38_2390 ();
 sg13g2_decap_8 FILLER_38_2402 ();
 sg13g2_decap_4 FILLER_38_2409 ();
 sg13g2_fill_2 FILLER_38_2413 ();
 sg13g2_decap_4 FILLER_38_2425 ();
 sg13g2_fill_1 FILLER_38_2429 ();
 sg13g2_fill_2 FILLER_38_2467 ();
 sg13g2_fill_1 FILLER_38_2469 ();
 sg13g2_fill_1 FILLER_38_2597 ();
 sg13g2_fill_2 FILLER_38_2611 ();
 sg13g2_fill_2 FILLER_38_2617 ();
 sg13g2_fill_1 FILLER_38_2659 ();
 sg13g2_decap_4 FILLER_38_2664 ();
 sg13g2_fill_2 FILLER_38_2668 ();
 sg13g2_decap_4 FILLER_39_0 ();
 sg13g2_decap_8 FILLER_39_54 ();
 sg13g2_decap_4 FILLER_39_61 ();
 sg13g2_fill_2 FILLER_39_106 ();
 sg13g2_decap_8 FILLER_39_134 ();
 sg13g2_decap_8 FILLER_39_141 ();
 sg13g2_decap_4 FILLER_39_148 ();
 sg13g2_decap_4 FILLER_39_161 ();
 sg13g2_fill_1 FILLER_39_200 ();
 sg13g2_fill_1 FILLER_39_205 ();
 sg13g2_fill_1 FILLER_39_213 ();
 sg13g2_fill_2 FILLER_39_241 ();
 sg13g2_fill_1 FILLER_39_269 ();
 sg13g2_decap_4 FILLER_39_279 ();
 sg13g2_fill_2 FILLER_39_328 ();
 sg13g2_fill_1 FILLER_39_330 ();
 sg13g2_fill_1 FILLER_39_341 ();
 sg13g2_fill_1 FILLER_39_361 ();
 sg13g2_fill_2 FILLER_39_375 ();
 sg13g2_fill_2 FILLER_39_386 ();
 sg13g2_fill_2 FILLER_39_408 ();
 sg13g2_fill_2 FILLER_39_440 ();
 sg13g2_fill_1 FILLER_39_472 ();
 sg13g2_fill_2 FILLER_39_508 ();
 sg13g2_fill_1 FILLER_39_510 ();
 sg13g2_decap_8 FILLER_39_521 ();
 sg13g2_decap_4 FILLER_39_528 ();
 sg13g2_fill_1 FILLER_39_532 ();
 sg13g2_fill_1 FILLER_39_559 ();
 sg13g2_fill_2 FILLER_39_577 ();
 sg13g2_fill_1 FILLER_39_615 ();
 sg13g2_fill_2 FILLER_39_673 ();
 sg13g2_fill_1 FILLER_39_675 ();
 sg13g2_fill_1 FILLER_39_686 ();
 sg13g2_decap_8 FILLER_39_691 ();
 sg13g2_fill_1 FILLER_39_698 ();
 sg13g2_fill_1 FILLER_39_712 ();
 sg13g2_fill_2 FILLER_39_717 ();
 sg13g2_fill_2 FILLER_39_745 ();
 sg13g2_fill_2 FILLER_39_751 ();
 sg13g2_fill_1 FILLER_39_753 ();
 sg13g2_decap_4 FILLER_39_794 ();
 sg13g2_fill_1 FILLER_39_798 ();
 sg13g2_fill_1 FILLER_39_828 ();
 sg13g2_decap_8 FILLER_39_840 ();
 sg13g2_decap_4 FILLER_39_847 ();
 sg13g2_fill_1 FILLER_39_851 ();
 sg13g2_fill_2 FILLER_39_862 ();
 sg13g2_fill_1 FILLER_39_927 ();
 sg13g2_decap_8 FILLER_39_964 ();
 sg13g2_fill_2 FILLER_39_971 ();
 sg13g2_fill_1 FILLER_39_973 ();
 sg13g2_fill_2 FILLER_39_983 ();
 sg13g2_decap_8 FILLER_39_1010 ();
 sg13g2_fill_1 FILLER_39_1074 ();
 sg13g2_fill_2 FILLER_39_1079 ();
 sg13g2_fill_1 FILLER_39_1081 ();
 sg13g2_fill_1 FILLER_39_1108 ();
 sg13g2_fill_1 FILLER_39_1135 ();
 sg13g2_decap_8 FILLER_39_1170 ();
 sg13g2_fill_2 FILLER_39_1177 ();
 sg13g2_fill_1 FILLER_39_1179 ();
 sg13g2_fill_1 FILLER_39_1223 ();
 sg13g2_fill_2 FILLER_39_1276 ();
 sg13g2_decap_4 FILLER_39_1344 ();
 sg13g2_fill_2 FILLER_39_1348 ();
 sg13g2_decap_4 FILLER_39_1354 ();
 sg13g2_fill_1 FILLER_39_1358 ();
 sg13g2_decap_8 FILLER_39_1363 ();
 sg13g2_decap_4 FILLER_39_1370 ();
 sg13g2_fill_2 FILLER_39_1374 ();
 sg13g2_decap_4 FILLER_39_1386 ();
 sg13g2_decap_4 FILLER_39_1394 ();
 sg13g2_decap_8 FILLER_39_1402 ();
 sg13g2_decap_8 FILLER_39_1409 ();
 sg13g2_fill_2 FILLER_39_1416 ();
 sg13g2_fill_1 FILLER_39_1418 ();
 sg13g2_fill_2 FILLER_39_1428 ();
 sg13g2_fill_2 FILLER_39_1444 ();
 sg13g2_fill_1 FILLER_39_1446 ();
 sg13g2_fill_1 FILLER_39_1504 ();
 sg13g2_decap_4 FILLER_39_1510 ();
 sg13g2_fill_1 FILLER_39_1514 ();
 sg13g2_fill_1 FILLER_39_1522 ();
 sg13g2_fill_2 FILLER_39_1570 ();
 sg13g2_fill_1 FILLER_39_1583 ();
 sg13g2_decap_4 FILLER_39_1597 ();
 sg13g2_fill_2 FILLER_39_1601 ();
 sg13g2_fill_2 FILLER_39_1606 ();
 sg13g2_fill_2 FILLER_39_1616 ();
 sg13g2_fill_1 FILLER_39_1618 ();
 sg13g2_fill_1 FILLER_39_1633 ();
 sg13g2_decap_8 FILLER_39_1638 ();
 sg13g2_decap_8 FILLER_39_1645 ();
 sg13g2_fill_1 FILLER_39_1652 ();
 sg13g2_decap_8 FILLER_39_1657 ();
 sg13g2_decap_8 FILLER_39_1664 ();
 sg13g2_fill_2 FILLER_39_1671 ();
 sg13g2_decap_4 FILLER_39_1678 ();
 sg13g2_decap_8 FILLER_39_1686 ();
 sg13g2_fill_2 FILLER_39_1693 ();
 sg13g2_fill_1 FILLER_39_1695 ();
 sg13g2_decap_8 FILLER_39_1706 ();
 sg13g2_fill_2 FILLER_39_1713 ();
 sg13g2_fill_1 FILLER_39_1715 ();
 sg13g2_decap_8 FILLER_39_1738 ();
 sg13g2_decap_8 FILLER_39_1745 ();
 sg13g2_decap_4 FILLER_39_1752 ();
 sg13g2_fill_2 FILLER_39_1761 ();
 sg13g2_fill_1 FILLER_39_1804 ();
 sg13g2_decap_4 FILLER_39_1828 ();
 sg13g2_fill_2 FILLER_39_1832 ();
 sg13g2_fill_2 FILLER_39_1839 ();
 sg13g2_decap_4 FILLER_39_1846 ();
 sg13g2_fill_1 FILLER_39_1850 ();
 sg13g2_decap_4 FILLER_39_1864 ();
 sg13g2_fill_1 FILLER_39_1868 ();
 sg13g2_decap_8 FILLER_39_1879 ();
 sg13g2_decap_8 FILLER_39_1886 ();
 sg13g2_fill_2 FILLER_39_1898 ();
 sg13g2_fill_1 FILLER_39_1900 ();
 sg13g2_fill_1 FILLER_39_1963 ();
 sg13g2_decap_8 FILLER_39_1968 ();
 sg13g2_fill_2 FILLER_39_1975 ();
 sg13g2_decap_4 FILLER_39_1987 ();
 sg13g2_decap_8 FILLER_39_2027 ();
 sg13g2_decap_8 FILLER_39_2034 ();
 sg13g2_decap_8 FILLER_39_2041 ();
 sg13g2_decap_8 FILLER_39_2048 ();
 sg13g2_fill_2 FILLER_39_2055 ();
 sg13g2_fill_1 FILLER_39_2057 ();
 sg13g2_fill_2 FILLER_39_2092 ();
 sg13g2_fill_1 FILLER_39_2094 ();
 sg13g2_fill_2 FILLER_39_2151 ();
 sg13g2_fill_2 FILLER_39_2176 ();
 sg13g2_decap_8 FILLER_39_2204 ();
 sg13g2_decap_8 FILLER_39_2211 ();
 sg13g2_decap_4 FILLER_39_2218 ();
 sg13g2_fill_2 FILLER_39_2222 ();
 sg13g2_decap_8 FILLER_39_2229 ();
 sg13g2_fill_2 FILLER_39_2236 ();
 sg13g2_fill_1 FILLER_39_2238 ();
 sg13g2_decap_8 FILLER_39_2259 ();
 sg13g2_fill_2 FILLER_39_2266 ();
 sg13g2_fill_1 FILLER_39_2268 ();
 sg13g2_fill_2 FILLER_39_2307 ();
 sg13g2_fill_1 FILLER_39_2319 ();
 sg13g2_fill_1 FILLER_39_2330 ();
 sg13g2_fill_1 FILLER_39_2335 ();
 sg13g2_fill_2 FILLER_39_2346 ();
 sg13g2_fill_2 FILLER_39_2353 ();
 sg13g2_fill_2 FILLER_39_2360 ();
 sg13g2_fill_1 FILLER_39_2362 ();
 sg13g2_fill_1 FILLER_39_2369 ();
 sg13g2_fill_1 FILLER_39_2375 ();
 sg13g2_fill_1 FILLER_39_2381 ();
 sg13g2_fill_2 FILLER_39_2386 ();
 sg13g2_decap_8 FILLER_39_2393 ();
 sg13g2_decap_8 FILLER_39_2400 ();
 sg13g2_fill_2 FILLER_39_2407 ();
 sg13g2_fill_2 FILLER_39_2465 ();
 sg13g2_fill_2 FILLER_39_2483 ();
 sg13g2_fill_1 FILLER_39_2485 ();
 sg13g2_fill_1 FILLER_39_2534 ();
 sg13g2_fill_2 FILLER_39_2544 ();
 sg13g2_fill_2 FILLER_39_2555 ();
 sg13g2_decap_8 FILLER_39_2645 ();
 sg13g2_decap_8 FILLER_39_2652 ();
 sg13g2_decap_8 FILLER_39_2659 ();
 sg13g2_decap_4 FILLER_39_2666 ();
 sg13g2_fill_1 FILLER_40_26 ();
 sg13g2_fill_2 FILLER_40_35 ();
 sg13g2_decap_8 FILLER_40_57 ();
 sg13g2_decap_8 FILLER_40_64 ();
 sg13g2_fill_1 FILLER_40_81 ();
 sg13g2_fill_1 FILLER_40_99 ();
 sg13g2_fill_2 FILLER_40_105 ();
 sg13g2_decap_8 FILLER_40_124 ();
 sg13g2_decap_4 FILLER_40_135 ();
 sg13g2_fill_2 FILLER_40_170 ();
 sg13g2_fill_1 FILLER_40_172 ();
 sg13g2_fill_2 FILLER_40_191 ();
 sg13g2_fill_1 FILLER_40_193 ();
 sg13g2_fill_1 FILLER_40_236 ();
 sg13g2_fill_2 FILLER_40_260 ();
 sg13g2_fill_1 FILLER_40_262 ();
 sg13g2_fill_2 FILLER_40_268 ();
 sg13g2_fill_1 FILLER_40_279 ();
 sg13g2_fill_2 FILLER_40_330 ();
 sg13g2_fill_1 FILLER_40_332 ();
 sg13g2_fill_1 FILLER_40_345 ();
 sg13g2_fill_2 FILLER_40_367 ();
 sg13g2_fill_1 FILLER_40_372 ();
 sg13g2_fill_2 FILLER_40_381 ();
 sg13g2_fill_2 FILLER_40_426 ();
 sg13g2_fill_1 FILLER_40_468 ();
 sg13g2_fill_2 FILLER_40_482 ();
 sg13g2_decap_4 FILLER_40_488 ();
 sg13g2_fill_2 FILLER_40_502 ();
 sg13g2_fill_1 FILLER_40_504 ();
 sg13g2_fill_1 FILLER_40_510 ();
 sg13g2_fill_2 FILLER_40_515 ();
 sg13g2_fill_1 FILLER_40_517 ();
 sg13g2_decap_8 FILLER_40_522 ();
 sg13g2_decap_8 FILLER_40_529 ();
 sg13g2_fill_1 FILLER_40_536 ();
 sg13g2_decap_8 FILLER_40_541 ();
 sg13g2_decap_4 FILLER_40_552 ();
 sg13g2_fill_1 FILLER_40_556 ();
 sg13g2_decap_4 FILLER_40_565 ();
 sg13g2_fill_1 FILLER_40_569 ();
 sg13g2_fill_1 FILLER_40_574 ();
 sg13g2_fill_1 FILLER_40_580 ();
 sg13g2_fill_2 FILLER_40_586 ();
 sg13g2_fill_1 FILLER_40_588 ();
 sg13g2_fill_1 FILLER_40_602 ();
 sg13g2_fill_1 FILLER_40_640 ();
 sg13g2_decap_4 FILLER_40_645 ();
 sg13g2_fill_2 FILLER_40_649 ();
 sg13g2_decap_8 FILLER_40_711 ();
 sg13g2_fill_2 FILLER_40_718 ();
 sg13g2_fill_2 FILLER_40_734 ();
 sg13g2_fill_1 FILLER_40_736 ();
 sg13g2_decap_4 FILLER_40_747 ();
 sg13g2_decap_4 FILLER_40_755 ();
 sg13g2_fill_2 FILLER_40_759 ();
 sg13g2_fill_2 FILLER_40_807 ();
 sg13g2_fill_1 FILLER_40_809 ();
 sg13g2_fill_1 FILLER_40_856 ();
 sg13g2_fill_2 FILLER_40_864 ();
 sg13g2_fill_2 FILLER_40_881 ();
 sg13g2_decap_4 FILLER_40_963 ();
 sg13g2_fill_1 FILLER_40_967 ();
 sg13g2_fill_2 FILLER_40_1018 ();
 sg13g2_fill_1 FILLER_40_1020 ();
 sg13g2_decap_4 FILLER_40_1051 ();
 sg13g2_decap_4 FILLER_40_1059 ();
 sg13g2_fill_2 FILLER_40_1063 ();
 sg13g2_fill_2 FILLER_40_1091 ();
 sg13g2_fill_1 FILLER_40_1093 ();
 sg13g2_fill_2 FILLER_40_1124 ();
 sg13g2_fill_1 FILLER_40_1131 ();
 sg13g2_fill_1 FILLER_40_1158 ();
 sg13g2_decap_8 FILLER_40_1163 ();
 sg13g2_decap_8 FILLER_40_1170 ();
 sg13g2_fill_2 FILLER_40_1207 ();
 sg13g2_fill_1 FILLER_40_1209 ();
 sg13g2_fill_2 FILLER_40_1214 ();
 sg13g2_decap_4 FILLER_40_1229 ();
 sg13g2_fill_2 FILLER_40_1237 ();
 sg13g2_decap_4 FILLER_40_1253 ();
 sg13g2_fill_1 FILLER_40_1291 ();
 sg13g2_fill_1 FILLER_40_1302 ();
 sg13g2_fill_2 FILLER_40_1338 ();
 sg13g2_fill_1 FILLER_40_1340 ();
 sg13g2_decap_8 FILLER_40_1361 ();
 sg13g2_decap_8 FILLER_40_1368 ();
 sg13g2_decap_8 FILLER_40_1375 ();
 sg13g2_fill_2 FILLER_40_1382 ();
 sg13g2_decap_4 FILLER_40_1420 ();
 sg13g2_fill_1 FILLER_40_1483 ();
 sg13g2_decap_4 FILLER_40_1514 ();
 sg13g2_fill_2 FILLER_40_1518 ();
 sg13g2_fill_2 FILLER_40_1533 ();
 sg13g2_fill_1 FILLER_40_1539 ();
 sg13g2_fill_2 FILLER_40_1586 ();
 sg13g2_fill_1 FILLER_40_1593 ();
 sg13g2_fill_2 FILLER_40_1650 ();
 sg13g2_decap_4 FILLER_40_1657 ();
 sg13g2_fill_2 FILLER_40_1661 ();
 sg13g2_decap_8 FILLER_40_1668 ();
 sg13g2_decap_4 FILLER_40_1675 ();
 sg13g2_fill_2 FILLER_40_1679 ();
 sg13g2_decap_4 FILLER_40_1685 ();
 sg13g2_decap_8 FILLER_40_1692 ();
 sg13g2_decap_4 FILLER_40_1699 ();
 sg13g2_fill_1 FILLER_40_1703 ();
 sg13g2_decap_4 FILLER_40_1708 ();
 sg13g2_decap_4 FILLER_40_1717 ();
 sg13g2_fill_2 FILLER_40_1721 ();
 sg13g2_decap_8 FILLER_40_1733 ();
 sg13g2_decap_8 FILLER_40_1740 ();
 sg13g2_decap_8 FILLER_40_1747 ();
 sg13g2_decap_8 FILLER_40_1754 ();
 sg13g2_decap_4 FILLER_40_1761 ();
 sg13g2_fill_2 FILLER_40_1765 ();
 sg13g2_fill_1 FILLER_40_1799 ();
 sg13g2_fill_2 FILLER_40_1809 ();
 sg13g2_fill_1 FILLER_40_1811 ();
 sg13g2_decap_8 FILLER_40_1842 ();
 sg13g2_decap_8 FILLER_40_1849 ();
 sg13g2_decap_4 FILLER_40_1856 ();
 sg13g2_fill_1 FILLER_40_1860 ();
 sg13g2_decap_8 FILLER_40_1870 ();
 sg13g2_fill_1 FILLER_40_1903 ();
 sg13g2_fill_2 FILLER_40_1907 ();
 sg13g2_fill_2 FILLER_40_1968 ();
 sg13g2_fill_1 FILLER_40_1970 ();
 sg13g2_decap_8 FILLER_40_2031 ();
 sg13g2_fill_1 FILLER_40_2038 ();
 sg13g2_decap_4 FILLER_40_2049 ();
 sg13g2_fill_2 FILLER_40_2119 ();
 sg13g2_decap_8 FILLER_40_2147 ();
 sg13g2_fill_2 FILLER_40_2154 ();
 sg13g2_decap_8 FILLER_40_2222 ();
 sg13g2_decap_8 FILLER_40_2229 ();
 sg13g2_fill_1 FILLER_40_2236 ();
 sg13g2_decap_8 FILLER_40_2247 ();
 sg13g2_decap_8 FILLER_40_2254 ();
 sg13g2_decap_8 FILLER_40_2261 ();
 sg13g2_decap_8 FILLER_40_2268 ();
 sg13g2_decap_8 FILLER_40_2275 ();
 sg13g2_decap_4 FILLER_40_2286 ();
 sg13g2_fill_2 FILLER_40_2290 ();
 sg13g2_fill_1 FILLER_40_2302 ();
 sg13g2_fill_1 FILLER_40_2307 ();
 sg13g2_fill_2 FILLER_40_2313 ();
 sg13g2_fill_1 FILLER_40_2315 ();
 sg13g2_decap_8 FILLER_40_2346 ();
 sg13g2_decap_8 FILLER_40_2353 ();
 sg13g2_decap_8 FILLER_40_2360 ();
 sg13g2_fill_2 FILLER_40_2367 ();
 sg13g2_decap_8 FILLER_40_2403 ();
 sg13g2_decap_4 FILLER_40_2410 ();
 sg13g2_decap_8 FILLER_40_2418 ();
 sg13g2_fill_1 FILLER_40_2425 ();
 sg13g2_fill_2 FILLER_40_2432 ();
 sg13g2_fill_1 FILLER_40_2434 ();
 sg13g2_fill_1 FILLER_40_2451 ();
 sg13g2_decap_8 FILLER_40_2459 ();
 sg13g2_decap_8 FILLER_40_2466 ();
 sg13g2_decap_8 FILLER_40_2473 ();
 sg13g2_fill_2 FILLER_40_2480 ();
 sg13g2_fill_1 FILLER_40_2482 ();
 sg13g2_fill_1 FILLER_40_2487 ();
 sg13g2_decap_4 FILLER_40_2492 ();
 sg13g2_fill_2 FILLER_40_2512 ();
 sg13g2_fill_2 FILLER_40_2539 ();
 sg13g2_fill_2 FILLER_40_2570 ();
 sg13g2_fill_2 FILLER_40_2581 ();
 sg13g2_decap_8 FILLER_40_2652 ();
 sg13g2_decap_8 FILLER_40_2659 ();
 sg13g2_decap_4 FILLER_40_2666 ();
 sg13g2_decap_8 FILLER_41_0 ();
 sg13g2_fill_1 FILLER_41_7 ();
 sg13g2_decap_8 FILLER_41_35 ();
 sg13g2_fill_2 FILLER_41_46 ();
 sg13g2_decap_8 FILLER_41_56 ();
 sg13g2_decap_8 FILLER_41_63 ();
 sg13g2_decap_8 FILLER_41_70 ();
 sg13g2_decap_8 FILLER_41_77 ();
 sg13g2_fill_1 FILLER_41_84 ();
 sg13g2_decap_8 FILLER_41_113 ();
 sg13g2_decap_4 FILLER_41_120 ();
 sg13g2_fill_1 FILLER_41_124 ();
 sg13g2_fill_1 FILLER_41_136 ();
 sg13g2_fill_2 FILLER_41_146 ();
 sg13g2_fill_2 FILLER_41_156 ();
 sg13g2_decap_8 FILLER_41_179 ();
 sg13g2_decap_8 FILLER_41_186 ();
 sg13g2_decap_8 FILLER_41_193 ();
 sg13g2_fill_2 FILLER_41_200 ();
 sg13g2_fill_1 FILLER_41_202 ();
 sg13g2_decap_4 FILLER_41_217 ();
 sg13g2_decap_8 FILLER_41_225 ();
 sg13g2_fill_2 FILLER_41_232 ();
 sg13g2_fill_1 FILLER_41_239 ();
 sg13g2_fill_2 FILLER_41_259 ();
 sg13g2_fill_1 FILLER_41_261 ();
 sg13g2_fill_1 FILLER_41_271 ();
 sg13g2_fill_1 FILLER_41_281 ();
 sg13g2_fill_2 FILLER_41_334 ();
 sg13g2_fill_1 FILLER_41_336 ();
 sg13g2_fill_1 FILLER_41_341 ();
 sg13g2_fill_2 FILLER_41_367 ();
 sg13g2_fill_2 FILLER_41_392 ();
 sg13g2_decap_4 FILLER_41_425 ();
 sg13g2_fill_1 FILLER_41_429 ();
 sg13g2_fill_2 FILLER_41_434 ();
 sg13g2_fill_1 FILLER_41_454 ();
 sg13g2_decap_8 FILLER_41_469 ();
 sg13g2_decap_8 FILLER_41_476 ();
 sg13g2_decap_8 FILLER_41_483 ();
 sg13g2_fill_2 FILLER_41_490 ();
 sg13g2_fill_1 FILLER_41_501 ();
 sg13g2_decap_8 FILLER_41_506 ();
 sg13g2_decap_8 FILLER_41_513 ();
 sg13g2_decap_8 FILLER_41_520 ();
 sg13g2_fill_2 FILLER_41_535 ();
 sg13g2_fill_2 FILLER_41_546 ();
 sg13g2_fill_1 FILLER_41_548 ();
 sg13g2_fill_2 FILLER_41_562 ();
 sg13g2_fill_1 FILLER_41_564 ();
 sg13g2_decap_4 FILLER_41_574 ();
 sg13g2_fill_2 FILLER_41_578 ();
 sg13g2_fill_2 FILLER_41_595 ();
 sg13g2_decap_4 FILLER_41_617 ();
 sg13g2_fill_2 FILLER_41_631 ();
 sg13g2_decap_8 FILLER_41_636 ();
 sg13g2_decap_4 FILLER_41_643 ();
 sg13g2_fill_2 FILLER_41_647 ();
 sg13g2_decap_4 FILLER_41_733 ();
 sg13g2_decap_8 FILLER_41_742 ();
 sg13g2_decap_8 FILLER_41_754 ();
 sg13g2_decap_8 FILLER_41_761 ();
 sg13g2_decap_8 FILLER_41_768 ();
 sg13g2_decap_4 FILLER_41_804 ();
 sg13g2_fill_1 FILLER_41_812 ();
 sg13g2_decap_4 FILLER_41_823 ();
 sg13g2_fill_1 FILLER_41_827 ();
 sg13g2_decap_8 FILLER_41_842 ();
 sg13g2_fill_1 FILLER_41_849 ();
 sg13g2_fill_1 FILLER_41_853 ();
 sg13g2_fill_2 FILLER_41_885 ();
 sg13g2_fill_2 FILLER_41_901 ();
 sg13g2_decap_4 FILLER_41_944 ();
 sg13g2_fill_1 FILLER_41_951 ();
 sg13g2_decap_4 FILLER_41_961 ();
 sg13g2_fill_2 FILLER_41_965 ();
 sg13g2_fill_1 FILLER_41_993 ();
 sg13g2_decap_8 FILLER_41_1025 ();
 sg13g2_fill_2 FILLER_41_1036 ();
 sg13g2_decap_8 FILLER_41_1041 ();
 sg13g2_decap_8 FILLER_41_1048 ();
 sg13g2_decap_4 FILLER_41_1055 ();
 sg13g2_fill_2 FILLER_41_1059 ();
 sg13g2_fill_2 FILLER_41_1066 ();
 sg13g2_fill_1 FILLER_41_1068 ();
 sg13g2_decap_8 FILLER_41_1126 ();
 sg13g2_decap_4 FILLER_41_1133 ();
 sg13g2_fill_1 FILLER_41_1137 ();
 sg13g2_decap_8 FILLER_41_1142 ();
 sg13g2_decap_8 FILLER_41_1149 ();
 sg13g2_decap_8 FILLER_41_1156 ();
 sg13g2_decap_8 FILLER_41_1163 ();
 sg13g2_decap_8 FILLER_41_1170 ();
 sg13g2_fill_1 FILLER_41_1177 ();
 sg13g2_fill_1 FILLER_41_1182 ();
 sg13g2_fill_2 FILLER_41_1193 ();
 sg13g2_fill_2 FILLER_41_1221 ();
 sg13g2_decap_4 FILLER_41_1233 ();
 sg13g2_decap_8 FILLER_41_1247 ();
 sg13g2_decap_8 FILLER_41_1254 ();
 sg13g2_decap_8 FILLER_41_1261 ();
 sg13g2_decap_8 FILLER_41_1304 ();
 sg13g2_fill_1 FILLER_41_1311 ();
 sg13g2_fill_2 FILLER_41_1316 ();
 sg13g2_fill_1 FILLER_41_1318 ();
 sg13g2_fill_2 FILLER_41_1369 ();
 sg13g2_decap_8 FILLER_41_1397 ();
 sg13g2_decap_8 FILLER_41_1404 ();
 sg13g2_decap_8 FILLER_41_1411 ();
 sg13g2_decap_8 FILLER_41_1418 ();
 sg13g2_decap_4 FILLER_41_1425 ();
 sg13g2_fill_1 FILLER_41_1429 ();
 sg13g2_fill_1 FILLER_41_1464 ();
 sg13g2_fill_2 FILLER_41_1477 ();
 sg13g2_fill_2 FILLER_41_1487 ();
 sg13g2_fill_2 FILLER_41_1493 ();
 sg13g2_fill_2 FILLER_41_1521 ();
 sg13g2_fill_1 FILLER_41_1523 ();
 sg13g2_fill_1 FILLER_41_1569 ();
 sg13g2_fill_2 FILLER_41_1595 ();
 sg13g2_decap_8 FILLER_41_1610 ();
 sg13g2_decap_8 FILLER_41_1617 ();
 sg13g2_decap_4 FILLER_41_1624 ();
 sg13g2_fill_2 FILLER_41_1628 ();
 sg13g2_fill_2 FILLER_41_1634 ();
 sg13g2_fill_1 FILLER_41_1636 ();
 sg13g2_fill_2 FILLER_41_1642 ();
 sg13g2_fill_1 FILLER_41_1644 ();
 sg13g2_decap_4 FILLER_41_1652 ();
 sg13g2_fill_2 FILLER_41_1656 ();
 sg13g2_decap_4 FILLER_41_1666 ();
 sg13g2_fill_2 FILLER_41_1670 ();
 sg13g2_fill_2 FILLER_41_1676 ();
 sg13g2_fill_2 FILLER_41_1692 ();
 sg13g2_fill_1 FILLER_41_1698 ();
 sg13g2_fill_2 FILLER_41_1703 ();
 sg13g2_fill_2 FILLER_41_1731 ();
 sg13g2_fill_1 FILLER_41_1733 ();
 sg13g2_fill_1 FILLER_41_1760 ();
 sg13g2_fill_2 FILLER_41_1767 ();
 sg13g2_fill_1 FILLER_41_1769 ();
 sg13g2_decap_4 FILLER_41_1774 ();
 sg13g2_fill_1 FILLER_41_1778 ();
 sg13g2_fill_1 FILLER_41_1784 ();
 sg13g2_decap_4 FILLER_41_1789 ();
 sg13g2_fill_2 FILLER_41_1793 ();
 sg13g2_fill_1 FILLER_41_1798 ();
 sg13g2_fill_1 FILLER_41_1805 ();
 sg13g2_decap_8 FILLER_41_1832 ();
 sg13g2_decap_8 FILLER_41_1839 ();
 sg13g2_decap_8 FILLER_41_1846 ();
 sg13g2_decap_8 FILLER_41_1853 ();
 sg13g2_decap_4 FILLER_41_1860 ();
 sg13g2_fill_2 FILLER_41_1864 ();
 sg13g2_fill_2 FILLER_41_1899 ();
 sg13g2_fill_1 FILLER_41_1931 ();
 sg13g2_fill_2 FILLER_41_1947 ();
 sg13g2_decap_8 FILLER_41_1955 ();
 sg13g2_fill_1 FILLER_41_1962 ();
 sg13g2_decap_8 FILLER_41_1967 ();
 sg13g2_decap_4 FILLER_41_1974 ();
 sg13g2_fill_1 FILLER_41_1978 ();
 sg13g2_decap_4 FILLER_41_1983 ();
 sg13g2_fill_2 FILLER_41_1987 ();
 sg13g2_fill_1 FILLER_41_2014 ();
 sg13g2_fill_2 FILLER_41_2019 ();
 sg13g2_fill_2 FILLER_41_2047 ();
 sg13g2_fill_2 FILLER_41_2059 ();
 sg13g2_fill_1 FILLER_41_2061 ();
 sg13g2_fill_1 FILLER_41_2072 ();
 sg13g2_decap_8 FILLER_41_2077 ();
 sg13g2_decap_8 FILLER_41_2084 ();
 sg13g2_decap_4 FILLER_41_2091 ();
 sg13g2_fill_2 FILLER_41_2095 ();
 sg13g2_decap_4 FILLER_41_2101 ();
 sg13g2_fill_1 FILLER_41_2105 ();
 sg13g2_fill_1 FILLER_41_2116 ();
 sg13g2_decap_4 FILLER_41_2130 ();
 sg13g2_fill_1 FILLER_41_2160 ();
 sg13g2_decap_4 FILLER_41_2175 ();
 sg13g2_decap_4 FILLER_41_2189 ();
 sg13g2_fill_2 FILLER_41_2193 ();
 sg13g2_decap_4 FILLER_41_2199 ();
 sg13g2_fill_2 FILLER_41_2203 ();
 sg13g2_decap_4 FILLER_41_2231 ();
 sg13g2_fill_1 FILLER_41_2235 ();
 sg13g2_decap_8 FILLER_41_2261 ();
 sg13g2_fill_1 FILLER_41_2268 ();
 sg13g2_decap_8 FILLER_41_2272 ();
 sg13g2_decap_8 FILLER_41_2279 ();
 sg13g2_decap_8 FILLER_41_2286 ();
 sg13g2_fill_1 FILLER_41_2293 ();
 sg13g2_decap_4 FILLER_41_2306 ();
 sg13g2_decap_4 FILLER_41_2315 ();
 sg13g2_fill_2 FILLER_41_2319 ();
 sg13g2_decap_4 FILLER_41_2325 ();
 sg13g2_decap_8 FILLER_41_2344 ();
 sg13g2_decap_4 FILLER_41_2351 ();
 sg13g2_fill_2 FILLER_41_2355 ();
 sg13g2_fill_1 FILLER_41_2395 ();
 sg13g2_decap_8 FILLER_41_2405 ();
 sg13g2_decap_4 FILLER_41_2412 ();
 sg13g2_fill_1 FILLER_41_2416 ();
 sg13g2_decap_8 FILLER_41_2422 ();
 sg13g2_decap_8 FILLER_41_2429 ();
 sg13g2_fill_2 FILLER_41_2436 ();
 sg13g2_fill_1 FILLER_41_2438 ();
 sg13g2_fill_2 FILLER_41_2449 ();
 sg13g2_fill_1 FILLER_41_2451 ();
 sg13g2_decap_8 FILLER_41_2508 ();
 sg13g2_decap_8 FILLER_41_2515 ();
 sg13g2_decap_4 FILLER_41_2528 ();
 sg13g2_fill_1 FILLER_41_2532 ();
 sg13g2_fill_1 FILLER_41_2615 ();
 sg13g2_decap_8 FILLER_41_2657 ();
 sg13g2_decap_4 FILLER_41_2664 ();
 sg13g2_fill_2 FILLER_41_2668 ();
 sg13g2_decap_8 FILLER_42_0 ();
 sg13g2_decap_8 FILLER_42_7 ();
 sg13g2_decap_8 FILLER_42_14 ();
 sg13g2_fill_2 FILLER_42_21 ();
 sg13g2_fill_1 FILLER_42_23 ();
 sg13g2_fill_2 FILLER_42_51 ();
 sg13g2_fill_2 FILLER_42_57 ();
 sg13g2_decap_4 FILLER_42_67 ();
 sg13g2_fill_2 FILLER_42_71 ();
 sg13g2_fill_1 FILLER_42_103 ();
 sg13g2_decap_8 FILLER_42_108 ();
 sg13g2_decap_8 FILLER_42_115 ();
 sg13g2_fill_2 FILLER_42_122 ();
 sg13g2_fill_1 FILLER_42_124 ();
 sg13g2_fill_2 FILLER_42_151 ();
 sg13g2_fill_1 FILLER_42_153 ();
 sg13g2_fill_2 FILLER_42_165 ();
 sg13g2_fill_2 FILLER_42_175 ();
 sg13g2_fill_2 FILLER_42_182 ();
 sg13g2_fill_2 FILLER_42_189 ();
 sg13g2_fill_2 FILLER_42_195 ();
 sg13g2_fill_2 FILLER_42_201 ();
 sg13g2_decap_4 FILLER_42_220 ();
 sg13g2_decap_4 FILLER_42_228 ();
 sg13g2_fill_1 FILLER_42_239 ();
 sg13g2_fill_2 FILLER_42_249 ();
 sg13g2_fill_1 FILLER_42_261 ();
 sg13g2_decap_8 FILLER_42_292 ();
 sg13g2_decap_8 FILLER_42_299 ();
 sg13g2_decap_4 FILLER_42_306 ();
 sg13g2_decap_8 FILLER_42_318 ();
 sg13g2_fill_1 FILLER_42_325 ();
 sg13g2_decap_4 FILLER_42_357 ();
 sg13g2_fill_2 FILLER_42_361 ();
 sg13g2_fill_2 FILLER_42_389 ();
 sg13g2_decap_8 FILLER_42_417 ();
 sg13g2_decap_8 FILLER_42_424 ();
 sg13g2_decap_4 FILLER_42_431 ();
 sg13g2_decap_4 FILLER_42_461 ();
 sg13g2_decap_8 FILLER_42_475 ();
 sg13g2_fill_2 FILLER_42_482 ();
 sg13g2_fill_1 FILLER_42_494 ();
 sg13g2_fill_2 FILLER_42_511 ();
 sg13g2_fill_1 FILLER_42_513 ();
 sg13g2_fill_2 FILLER_42_520 ();
 sg13g2_fill_1 FILLER_42_522 ();
 sg13g2_fill_1 FILLER_42_528 ();
 sg13g2_fill_2 FILLER_42_534 ();
 sg13g2_fill_1 FILLER_42_536 ();
 sg13g2_fill_2 FILLER_42_596 ();
 sg13g2_fill_1 FILLER_42_603 ();
 sg13g2_fill_1 FILLER_42_609 ();
 sg13g2_fill_2 FILLER_42_641 ();
 sg13g2_fill_1 FILLER_42_648 ();
 sg13g2_fill_2 FILLER_42_656 ();
 sg13g2_fill_1 FILLER_42_675 ();
 sg13g2_fill_1 FILLER_42_681 ();
 sg13g2_fill_1 FILLER_42_702 ();
 sg13g2_fill_2 FILLER_42_707 ();
 sg13g2_fill_1 FILLER_42_709 ();
 sg13g2_fill_1 FILLER_42_714 ();
 sg13g2_fill_1 FILLER_42_720 ();
 sg13g2_fill_1 FILLER_42_725 ();
 sg13g2_fill_1 FILLER_42_731 ();
 sg13g2_fill_2 FILLER_42_737 ();
 sg13g2_fill_2 FILLER_42_743 ();
 sg13g2_fill_1 FILLER_42_757 ();
 sg13g2_decap_4 FILLER_42_768 ();
 sg13g2_decap_4 FILLER_42_777 ();
 sg13g2_fill_2 FILLER_42_785 ();
 sg13g2_fill_1 FILLER_42_787 ();
 sg13g2_decap_8 FILLER_42_792 ();
 sg13g2_decap_4 FILLER_42_799 ();
 sg13g2_fill_2 FILLER_42_803 ();
 sg13g2_fill_2 FILLER_42_809 ();
 sg13g2_fill_1 FILLER_42_831 ();
 sg13g2_decap_4 FILLER_42_836 ();
 sg13g2_fill_2 FILLER_42_840 ();
 sg13g2_fill_2 FILLER_42_864 ();
 sg13g2_fill_2 FILLER_42_870 ();
 sg13g2_fill_1 FILLER_42_910 ();
 sg13g2_fill_2 FILLER_42_927 ();
 sg13g2_fill_2 FILLER_42_933 ();
 sg13g2_fill_1 FILLER_42_940 ();
 sg13g2_fill_2 FILLER_42_995 ();
 sg13g2_fill_1 FILLER_42_997 ();
 sg13g2_fill_2 FILLER_42_1032 ();
 sg13g2_fill_1 FILLER_42_1034 ();
 sg13g2_decap_8 FILLER_42_1046 ();
 sg13g2_decap_8 FILLER_42_1053 ();
 sg13g2_fill_1 FILLER_42_1060 ();
 sg13g2_decap_8 FILLER_42_1069 ();
 sg13g2_decap_8 FILLER_42_1076 ();
 sg13g2_fill_2 FILLER_42_1087 ();
 sg13g2_fill_2 FILLER_42_1093 ();
 sg13g2_decap_4 FILLER_42_1099 ();
 sg13g2_fill_1 FILLER_42_1103 ();
 sg13g2_decap_8 FILLER_42_1108 ();
 sg13g2_decap_8 FILLER_42_1115 ();
 sg13g2_fill_1 FILLER_42_1122 ();
 sg13g2_decap_8 FILLER_42_1167 ();
 sg13g2_decap_8 FILLER_42_1174 ();
 sg13g2_decap_8 FILLER_42_1181 ();
 sg13g2_decap_8 FILLER_42_1188 ();
 sg13g2_decap_8 FILLER_42_1195 ();
 sg13g2_decap_8 FILLER_42_1202 ();
 sg13g2_decap_8 FILLER_42_1209 ();
 sg13g2_decap_8 FILLER_42_1216 ();
 sg13g2_fill_2 FILLER_42_1236 ();
 sg13g2_fill_1 FILLER_42_1238 ();
 sg13g2_fill_1 FILLER_42_1249 ();
 sg13g2_decap_8 FILLER_42_1263 ();
 sg13g2_decap_4 FILLER_42_1270 ();
 sg13g2_fill_2 FILLER_42_1274 ();
 sg13g2_decap_8 FILLER_42_1280 ();
 sg13g2_decap_8 FILLER_42_1287 ();
 sg13g2_decap_8 FILLER_42_1294 ();
 sg13g2_fill_1 FILLER_42_1301 ();
 sg13g2_fill_1 FILLER_42_1322 ();
 sg13g2_fill_2 FILLER_42_1336 ();
 sg13g2_fill_2 FILLER_42_1343 ();
 sg13g2_fill_1 FILLER_42_1345 ();
 sg13g2_decap_8 FILLER_42_1350 ();
 sg13g2_fill_2 FILLER_42_1361 ();
 sg13g2_fill_1 FILLER_42_1363 ();
 sg13g2_fill_2 FILLER_42_1377 ();
 sg13g2_fill_1 FILLER_42_1379 ();
 sg13g2_decap_4 FILLER_42_1385 ();
 sg13g2_fill_2 FILLER_42_1399 ();
 sg13g2_fill_1 FILLER_42_1401 ();
 sg13g2_fill_1 FILLER_42_1407 ();
 sg13g2_decap_8 FILLER_42_1413 ();
 sg13g2_decap_4 FILLER_42_1420 ();
 sg13g2_fill_1 FILLER_42_1449 ();
 sg13g2_fill_2 FILLER_42_1497 ();
 sg13g2_fill_1 FILLER_42_1499 ();
 sg13g2_decap_4 FILLER_42_1526 ();
 sg13g2_fill_1 FILLER_42_1530 ();
 sg13g2_decap_8 FILLER_42_1535 ();
 sg13g2_fill_2 FILLER_42_1542 ();
 sg13g2_fill_2 FILLER_42_1551 ();
 sg13g2_decap_8 FILLER_42_1575 ();
 sg13g2_decap_8 FILLER_42_1582 ();
 sg13g2_decap_4 FILLER_42_1589 ();
 sg13g2_decap_4 FILLER_42_1598 ();
 sg13g2_fill_1 FILLER_42_1602 ();
 sg13g2_decap_4 FILLER_42_1616 ();
 sg13g2_fill_2 FILLER_42_1620 ();
 sg13g2_fill_1 FILLER_42_1648 ();
 sg13g2_decap_4 FILLER_42_1717 ();
 sg13g2_fill_1 FILLER_42_1721 ();
 sg13g2_fill_1 FILLER_42_1748 ();
 sg13g2_fill_1 FILLER_42_1780 ();
 sg13g2_fill_1 FILLER_42_1796 ();
 sg13g2_decap_8 FILLER_42_1827 ();
 sg13g2_decap_8 FILLER_42_1834 ();
 sg13g2_decap_8 FILLER_42_1841 ();
 sg13g2_decap_8 FILLER_42_1848 ();
 sg13g2_decap_8 FILLER_42_1855 ();
 sg13g2_decap_8 FILLER_42_1862 ();
 sg13g2_fill_2 FILLER_42_1869 ();
 sg13g2_decap_4 FILLER_42_1876 ();
 sg13g2_decap_4 FILLER_42_1884 ();
 sg13g2_decap_8 FILLER_42_1892 ();
 sg13g2_fill_1 FILLER_42_1911 ();
 sg13g2_fill_1 FILLER_42_1924 ();
 sg13g2_fill_1 FILLER_42_1928 ();
 sg13g2_fill_2 FILLER_42_1944 ();
 sg13g2_fill_1 FILLER_42_1946 ();
 sg13g2_fill_1 FILLER_42_1962 ();
 sg13g2_decap_4 FILLER_42_1967 ();
 sg13g2_decap_8 FILLER_42_1975 ();
 sg13g2_decap_8 FILLER_42_1982 ();
 sg13g2_fill_1 FILLER_42_1989 ();
 sg13g2_decap_8 FILLER_42_1994 ();
 sg13g2_decap_4 FILLER_42_2001 ();
 sg13g2_fill_2 FILLER_42_2005 ();
 sg13g2_fill_2 FILLER_42_2032 ();
 sg13g2_fill_1 FILLER_42_2034 ();
 sg13g2_fill_1 FILLER_42_2061 ();
 sg13g2_fill_2 FILLER_42_2088 ();
 sg13g2_fill_2 FILLER_42_2116 ();
 sg13g2_fill_2 FILLER_42_2139 ();
 sg13g2_decap_8 FILLER_42_2145 ();
 sg13g2_decap_8 FILLER_42_2152 ();
 sg13g2_fill_2 FILLER_42_2159 ();
 sg13g2_fill_1 FILLER_42_2161 ();
 sg13g2_decap_8 FILLER_42_2188 ();
 sg13g2_decap_8 FILLER_42_2195 ();
 sg13g2_decap_8 FILLER_42_2202 ();
 sg13g2_decap_4 FILLER_42_2209 ();
 sg13g2_fill_1 FILLER_42_2213 ();
 sg13g2_fill_1 FILLER_42_2218 ();
 sg13g2_fill_1 FILLER_42_2245 ();
 sg13g2_decap_4 FILLER_42_2272 ();
 sg13g2_fill_2 FILLER_42_2276 ();
 sg13g2_fill_1 FILLER_42_2304 ();
 sg13g2_fill_2 FILLER_42_2309 ();
 sg13g2_fill_1 FILLER_42_2311 ();
 sg13g2_decap_4 FILLER_42_2317 ();
 sg13g2_fill_1 FILLER_42_2341 ();
 sg13g2_fill_1 FILLER_42_2396 ();
 sg13g2_fill_2 FILLER_42_2405 ();
 sg13g2_fill_2 FILLER_42_2421 ();
 sg13g2_fill_2 FILLER_42_2479 ();
 sg13g2_fill_1 FILLER_42_2481 ();
 sg13g2_fill_2 FILLER_42_2505 ();
 sg13g2_decap_8 FILLER_42_2512 ();
 sg13g2_fill_2 FILLER_42_2519 ();
 sg13g2_fill_1 FILLER_42_2521 ();
 sg13g2_fill_1 FILLER_42_2552 ();
 sg13g2_fill_2 FILLER_42_2557 ();
 sg13g2_fill_2 FILLER_42_2636 ();
 sg13g2_decap_4 FILLER_42_2664 ();
 sg13g2_fill_2 FILLER_42_2668 ();
 sg13g2_decap_8 FILLER_43_0 ();
 sg13g2_decap_8 FILLER_43_7 ();
 sg13g2_decap_8 FILLER_43_14 ();
 sg13g2_fill_1 FILLER_43_21 ();
 sg13g2_fill_2 FILLER_43_31 ();
 sg13g2_fill_2 FILLER_43_67 ();
 sg13g2_fill_2 FILLER_43_74 ();
 sg13g2_fill_1 FILLER_43_76 ();
 sg13g2_fill_1 FILLER_43_97 ();
 sg13g2_fill_2 FILLER_43_117 ();
 sg13g2_fill_2 FILLER_43_131 ();
 sg13g2_fill_2 FILLER_43_138 ();
 sg13g2_fill_2 FILLER_43_147 ();
 sg13g2_fill_1 FILLER_43_154 ();
 sg13g2_fill_2 FILLER_43_233 ();
 sg13g2_fill_1 FILLER_43_235 ();
 sg13g2_fill_1 FILLER_43_241 ();
 sg13g2_fill_1 FILLER_43_248 ();
 sg13g2_fill_2 FILLER_43_262 ();
 sg13g2_decap_4 FILLER_43_290 ();
 sg13g2_decap_4 FILLER_43_298 ();
 sg13g2_fill_2 FILLER_43_302 ();
 sg13g2_decap_8 FILLER_43_309 ();
 sg13g2_decap_8 FILLER_43_316 ();
 sg13g2_fill_1 FILLER_43_327 ();
 sg13g2_fill_2 FILLER_43_354 ();
 sg13g2_fill_2 FILLER_43_382 ();
 sg13g2_fill_1 FILLER_43_409 ();
 sg13g2_decap_8 FILLER_43_427 ();
 sg13g2_decap_8 FILLER_43_434 ();
 sg13g2_fill_1 FILLER_43_441 ();
 sg13g2_fill_1 FILLER_43_472 ();
 sg13g2_fill_2 FILLER_43_570 ();
 sg13g2_fill_2 FILLER_43_605 ();
 sg13g2_fill_1 FILLER_43_630 ();
 sg13g2_fill_2 FILLER_43_636 ();
 sg13g2_fill_2 FILLER_43_663 ();
 sg13g2_fill_1 FILLER_43_665 ();
 sg13g2_decap_8 FILLER_43_679 ();
 sg13g2_decap_4 FILLER_43_686 ();
 sg13g2_fill_2 FILLER_43_690 ();
 sg13g2_decap_8 FILLER_43_696 ();
 sg13g2_fill_2 FILLER_43_703 ();
 sg13g2_fill_1 FILLER_43_705 ();
 sg13g2_fill_2 FILLER_43_711 ();
 sg13g2_fill_2 FILLER_43_770 ();
 sg13g2_fill_2 FILLER_43_801 ();
 sg13g2_fill_2 FILLER_43_816 ();
 sg13g2_fill_1 FILLER_43_818 ();
 sg13g2_fill_2 FILLER_43_845 ();
 sg13g2_fill_1 FILLER_43_857 ();
 sg13g2_fill_1 FILLER_43_863 ();
 sg13g2_fill_1 FILLER_43_893 ();
 sg13g2_fill_2 FILLER_43_930 ();
 sg13g2_fill_1 FILLER_43_932 ();
 sg13g2_fill_1 FILLER_43_946 ();
 sg13g2_fill_1 FILLER_43_962 ();
 sg13g2_decap_4 FILLER_43_981 ();
 sg13g2_fill_1 FILLER_43_985 ();
 sg13g2_fill_2 FILLER_43_1012 ();
 sg13g2_fill_1 FILLER_43_1014 ();
 sg13g2_decap_8 FILLER_43_1025 ();
 sg13g2_decap_4 FILLER_43_1075 ();
 sg13g2_fill_2 FILLER_43_1079 ();
 sg13g2_fill_2 FILLER_43_1085 ();
 sg13g2_fill_1 FILLER_43_1087 ();
 sg13g2_fill_2 FILLER_43_1097 ();
 sg13g2_fill_1 FILLER_43_1099 ();
 sg13g2_fill_2 FILLER_43_1104 ();
 sg13g2_fill_1 FILLER_43_1111 ();
 sg13g2_fill_2 FILLER_43_1119 ();
 sg13g2_fill_1 FILLER_43_1121 ();
 sg13g2_fill_1 FILLER_43_1148 ();
 sg13g2_fill_2 FILLER_43_1153 ();
 sg13g2_fill_2 FILLER_43_1181 ();
 sg13g2_fill_2 FILLER_43_1187 ();
 sg13g2_decap_8 FILLER_43_1202 ();
 sg13g2_decap_8 FILLER_43_1209 ();
 sg13g2_decap_8 FILLER_43_1216 ();
 sg13g2_fill_2 FILLER_43_1223 ();
 sg13g2_decap_4 FILLER_43_1239 ();
 sg13g2_fill_1 FILLER_43_1243 ();
 sg13g2_decap_4 FILLER_43_1264 ();
 sg13g2_decap_4 FILLER_43_1278 ();
 sg13g2_fill_2 FILLER_43_1282 ();
 sg13g2_decap_4 FILLER_43_1290 ();
 sg13g2_fill_2 FILLER_43_1294 ();
 sg13g2_fill_1 FILLER_43_1306 ();
 sg13g2_decap_4 FILLER_43_1313 ();
 sg13g2_fill_2 FILLER_43_1353 ();
 sg13g2_fill_1 FILLER_43_1355 ();
 sg13g2_decap_8 FILLER_43_1372 ();
 sg13g2_decap_4 FILLER_43_1379 ();
 sg13g2_fill_2 FILLER_43_1388 ();
 sg13g2_fill_1 FILLER_43_1400 ();
 sg13g2_fill_2 FILLER_43_1415 ();
 sg13g2_fill_1 FILLER_43_1425 ();
 sg13g2_fill_2 FILLER_43_1431 ();
 sg13g2_fill_1 FILLER_43_1444 ();
 sg13g2_fill_2 FILLER_43_1455 ();
 sg13g2_fill_1 FILLER_43_1470 ();
 sg13g2_fill_2 FILLER_43_1497 ();
 sg13g2_fill_2 FILLER_43_1515 ();
 sg13g2_fill_1 FILLER_43_1517 ();
 sg13g2_decap_8 FILLER_43_1527 ();
 sg13g2_fill_2 FILLER_43_1534 ();
 sg13g2_fill_1 FILLER_43_1540 ();
 sg13g2_fill_2 FILLER_43_1596 ();
 sg13g2_fill_1 FILLER_43_1602 ();
 sg13g2_fill_1 FILLER_43_1618 ();
 sg13g2_fill_1 FILLER_43_1629 ();
 sg13g2_fill_1 FILLER_43_1634 ();
 sg13g2_fill_1 FILLER_43_1642 ();
 sg13g2_fill_1 FILLER_43_1648 ();
 sg13g2_fill_2 FILLER_43_1656 ();
 sg13g2_fill_1 FILLER_43_1662 ();
 sg13g2_fill_2 FILLER_43_1675 ();
 sg13g2_fill_1 FILLER_43_1677 ();
 sg13g2_decap_8 FILLER_43_1682 ();
 sg13g2_decap_4 FILLER_43_1689 ();
 sg13g2_fill_1 FILLER_43_1693 ();
 sg13g2_decap_8 FILLER_43_1708 ();
 sg13g2_decap_8 FILLER_43_1715 ();
 sg13g2_decap_8 FILLER_43_1722 ();
 sg13g2_fill_2 FILLER_43_1733 ();
 sg13g2_fill_1 FILLER_43_1735 ();
 sg13g2_fill_2 FILLER_43_1745 ();
 sg13g2_fill_1 FILLER_43_1747 ();
 sg13g2_decap_4 FILLER_43_1751 ();
 sg13g2_fill_2 FILLER_43_1755 ();
 sg13g2_decap_8 FILLER_43_1786 ();
 sg13g2_decap_8 FILLER_43_1793 ();
 sg13g2_fill_2 FILLER_43_1800 ();
 sg13g2_fill_1 FILLER_43_1802 ();
 sg13g2_decap_8 FILLER_43_1807 ();
 sg13g2_decap_8 FILLER_43_1814 ();
 sg13g2_decap_8 FILLER_43_1821 ();
 sg13g2_decap_8 FILLER_43_1828 ();
 sg13g2_decap_4 FILLER_43_1835 ();
 sg13g2_decap_4 FILLER_43_1844 ();
 sg13g2_fill_2 FILLER_43_1852 ();
 sg13g2_decap_8 FILLER_43_1858 ();
 sg13g2_fill_1 FILLER_43_1865 ();
 sg13g2_fill_2 FILLER_43_1870 ();
 sg13g2_decap_8 FILLER_43_1876 ();
 sg13g2_decap_8 FILLER_43_1883 ();
 sg13g2_fill_2 FILLER_43_1890 ();
 sg13g2_fill_1 FILLER_43_1892 ();
 sg13g2_fill_1 FILLER_43_1919 ();
 sg13g2_fill_1 FILLER_43_1925 ();
 sg13g2_fill_1 FILLER_43_1931 ();
 sg13g2_decap_8 FILLER_43_1957 ();
 sg13g2_fill_2 FILLER_43_1964 ();
 sg13g2_decap_4 FILLER_43_1976 ();
 sg13g2_fill_1 FILLER_43_1980 ();
 sg13g2_decap_8 FILLER_43_1991 ();
 sg13g2_decap_8 FILLER_43_1998 ();
 sg13g2_decap_8 FILLER_43_2010 ();
 sg13g2_fill_1 FILLER_43_2017 ();
 sg13g2_decap_8 FILLER_43_2022 ();
 sg13g2_decap_8 FILLER_43_2029 ();
 sg13g2_decap_4 FILLER_43_2036 ();
 sg13g2_fill_2 FILLER_43_2040 ();
 sg13g2_decap_4 FILLER_43_2046 ();
 sg13g2_fill_2 FILLER_43_2050 ();
 sg13g2_decap_8 FILLER_43_2092 ();
 sg13g2_decap_8 FILLER_43_2099 ();
 sg13g2_decap_4 FILLER_43_2106 ();
 sg13g2_fill_2 FILLER_43_2110 ();
 sg13g2_decap_8 FILLER_43_2142 ();
 sg13g2_decap_4 FILLER_43_2149 ();
 sg13g2_fill_2 FILLER_43_2153 ();
 sg13g2_decap_8 FILLER_43_2160 ();
 sg13g2_decap_4 FILLER_43_2167 ();
 sg13g2_decap_8 FILLER_43_2181 ();
 sg13g2_decap_8 FILLER_43_2188 ();
 sg13g2_decap_8 FILLER_43_2195 ();
 sg13g2_decap_8 FILLER_43_2202 ();
 sg13g2_decap_8 FILLER_43_2209 ();
 sg13g2_fill_2 FILLER_43_2226 ();
 sg13g2_decap_8 FILLER_43_2258 ();
 sg13g2_fill_1 FILLER_43_2265 ();
 sg13g2_fill_1 FILLER_43_2302 ();
 sg13g2_fill_1 FILLER_43_2318 ();
 sg13g2_fill_1 FILLER_43_2371 ();
 sg13g2_fill_1 FILLER_43_2389 ();
 sg13g2_fill_2 FILLER_43_2395 ();
 sg13g2_fill_2 FILLER_43_2428 ();
 sg13g2_fill_1 FILLER_43_2456 ();
 sg13g2_fill_1 FILLER_43_2461 ();
 sg13g2_fill_2 FILLER_43_2488 ();
 sg13g2_decap_4 FILLER_43_2520 ();
 sg13g2_decap_4 FILLER_43_2528 ();
 sg13g2_fill_1 FILLER_43_2536 ();
 sg13g2_fill_1 FILLER_43_2563 ();
 sg13g2_fill_1 FILLER_43_2616 ();
 sg13g2_fill_2 FILLER_43_2642 ();
 sg13g2_fill_2 FILLER_44_0 ();
 sg13g2_fill_2 FILLER_44_69 ();
 sg13g2_fill_1 FILLER_44_114 ();
 sg13g2_fill_1 FILLER_44_120 ();
 sg13g2_fill_1 FILLER_44_158 ();
 sg13g2_fill_1 FILLER_44_162 ();
 sg13g2_fill_1 FILLER_44_169 ();
 sg13g2_fill_1 FILLER_44_175 ();
 sg13g2_fill_1 FILLER_44_185 ();
 sg13g2_fill_2 FILLER_44_192 ();
 sg13g2_fill_1 FILLER_44_222 ();
 sg13g2_fill_2 FILLER_44_231 ();
 sg13g2_decap_4 FILLER_44_237 ();
 sg13g2_fill_2 FILLER_44_241 ();
 sg13g2_fill_1 FILLER_44_264 ();
 sg13g2_fill_2 FILLER_44_269 ();
 sg13g2_decap_8 FILLER_44_310 ();
 sg13g2_decap_8 FILLER_44_317 ();
 sg13g2_decap_8 FILLER_44_324 ();
 sg13g2_decap_8 FILLER_44_331 ();
 sg13g2_decap_4 FILLER_44_338 ();
 sg13g2_fill_1 FILLER_44_342 ();
 sg13g2_fill_1 FILLER_44_366 ();
 sg13g2_fill_1 FILLER_44_455 ();
 sg13g2_fill_1 FILLER_44_466 ();
 sg13g2_fill_2 FILLER_44_489 ();
 sg13g2_fill_2 FILLER_44_496 ();
 sg13g2_decap_4 FILLER_44_515 ();
 sg13g2_fill_1 FILLER_44_519 ();
 sg13g2_fill_2 FILLER_44_525 ();
 sg13g2_fill_1 FILLER_44_527 ();
 sg13g2_decap_8 FILLER_44_533 ();
 sg13g2_fill_1 FILLER_44_540 ();
 sg13g2_fill_2 FILLER_44_545 ();
 sg13g2_fill_1 FILLER_44_547 ();
 sg13g2_fill_1 FILLER_44_553 ();
 sg13g2_decap_4 FILLER_44_558 ();
 sg13g2_fill_2 FILLER_44_626 ();
 sg13g2_fill_2 FILLER_44_663 ();
 sg13g2_decap_8 FILLER_44_685 ();
 sg13g2_decap_8 FILLER_44_692 ();
 sg13g2_fill_1 FILLER_44_708 ();
 sg13g2_fill_2 FILLER_44_713 ();
 sg13g2_fill_1 FILLER_44_715 ();
 sg13g2_decap_4 FILLER_44_725 ();
 sg13g2_fill_1 FILLER_44_733 ();
 sg13g2_fill_1 FILLER_44_767 ();
 sg13g2_decap_4 FILLER_44_830 ();
 sg13g2_fill_1 FILLER_44_838 ();
 sg13g2_fill_2 FILLER_44_855 ();
 sg13g2_fill_2 FILLER_44_869 ();
 sg13g2_fill_1 FILLER_44_883 ();
 sg13g2_fill_1 FILLER_44_903 ();
 sg13g2_fill_1 FILLER_44_915 ();
 sg13g2_fill_1 FILLER_44_920 ();
 sg13g2_fill_1 FILLER_44_951 ();
 sg13g2_fill_2 FILLER_44_957 ();
 sg13g2_fill_2 FILLER_44_979 ();
 sg13g2_fill_1 FILLER_44_993 ();
 sg13g2_fill_2 FILLER_44_1004 ();
 sg13g2_fill_1 FILLER_44_1006 ();
 sg13g2_decap_8 FILLER_44_1011 ();
 sg13g2_fill_1 FILLER_44_1018 ();
 sg13g2_decap_8 FILLER_44_1049 ();
 sg13g2_decap_4 FILLER_44_1056 ();
 sg13g2_fill_1 FILLER_44_1060 ();
 sg13g2_fill_1 FILLER_44_1092 ();
 sg13g2_fill_2 FILLER_44_1122 ();
 sg13g2_decap_8 FILLER_44_1128 ();
 sg13g2_fill_2 FILLER_44_1145 ();
 sg13g2_fill_1 FILLER_44_1147 ();
 sg13g2_decap_4 FILLER_44_1171 ();
 sg13g2_fill_2 FILLER_44_1175 ();
 sg13g2_fill_2 FILLER_44_1230 ();
 sg13g2_decap_8 FILLER_44_1236 ();
 sg13g2_decap_4 FILLER_44_1259 ();
 sg13g2_decap_4 FILLER_44_1272 ();
 sg13g2_fill_1 FILLER_44_1280 ();
 sg13g2_decap_8 FILLER_44_1299 ();
 sg13g2_decap_4 FILLER_44_1306 ();
 sg13g2_fill_2 FILLER_44_1310 ();
 sg13g2_decap_8 FILLER_44_1352 ();
 sg13g2_fill_1 FILLER_44_1359 ();
 sg13g2_fill_1 FILLER_44_1370 ();
 sg13g2_fill_1 FILLER_44_1400 ();
 sg13g2_fill_2 FILLER_44_1495 ();
 sg13g2_fill_1 FILLER_44_1510 ();
 sg13g2_decap_4 FILLER_44_1583 ();
 sg13g2_fill_2 FILLER_44_1608 ();
 sg13g2_fill_1 FILLER_44_1610 ();
 sg13g2_fill_2 FILLER_44_1621 ();
 sg13g2_fill_2 FILLER_44_1636 ();
 sg13g2_fill_2 FILLER_44_1642 ();
 sg13g2_fill_1 FILLER_44_1657 ();
 sg13g2_fill_2 FILLER_44_1666 ();
 sg13g2_decap_4 FILLER_44_1694 ();
 sg13g2_fill_2 FILLER_44_1724 ();
 sg13g2_fill_2 FILLER_44_1731 ();
 sg13g2_fill_1 FILLER_44_1759 ();
 sg13g2_fill_2 FILLER_44_1764 ();
 sg13g2_fill_2 FILLER_44_1770 ();
 sg13g2_fill_1 FILLER_44_1772 ();
 sg13g2_fill_1 FILLER_44_1807 ();
 sg13g2_fill_2 FILLER_44_1825 ();
 sg13g2_fill_1 FILLER_44_1827 ();
 sg13g2_fill_1 FILLER_44_1854 ();
 sg13g2_fill_2 FILLER_44_1859 ();
 sg13g2_fill_2 FILLER_44_1876 ();
 sg13g2_fill_1 FILLER_44_1878 ();
 sg13g2_decap_8 FILLER_44_1887 ();
 sg13g2_decap_4 FILLER_44_1894 ();
 sg13g2_fill_1 FILLER_44_1898 ();
 sg13g2_fill_1 FILLER_44_1902 ();
 sg13g2_fill_2 FILLER_44_1908 ();
 sg13g2_decap_8 FILLER_44_1951 ();
 sg13g2_fill_2 FILLER_44_1988 ();
 sg13g2_fill_1 FILLER_44_1990 ();
 sg13g2_decap_4 FILLER_44_1995 ();
 sg13g2_decap_8 FILLER_44_2003 ();
 sg13g2_decap_4 FILLER_44_2010 ();
 sg13g2_fill_2 FILLER_44_2014 ();
 sg13g2_fill_2 FILLER_44_2020 ();
 sg13g2_fill_1 FILLER_44_2022 ();
 sg13g2_decap_8 FILLER_44_2028 ();
 sg13g2_decap_8 FILLER_44_2035 ();
 sg13g2_decap_8 FILLER_44_2042 ();
 sg13g2_decap_4 FILLER_44_2049 ();
 sg13g2_fill_1 FILLER_44_2053 ();
 sg13g2_fill_2 FILLER_44_2062 ();
 sg13g2_decap_8 FILLER_44_2100 ();
 sg13g2_decap_4 FILLER_44_2107 ();
 sg13g2_decap_8 FILLER_44_2124 ();
 sg13g2_fill_1 FILLER_44_2131 ();
 sg13g2_decap_4 FILLER_44_2153 ();
 sg13g2_fill_2 FILLER_44_2157 ();
 sg13g2_decap_8 FILLER_44_2195 ();
 sg13g2_fill_2 FILLER_44_2202 ();
 sg13g2_fill_1 FILLER_44_2204 ();
 sg13g2_decap_4 FILLER_44_2210 ();
 sg13g2_fill_2 FILLER_44_2245 ();
 sg13g2_fill_1 FILLER_44_2296 ();
 sg13g2_fill_2 FILLER_44_2327 ();
 sg13g2_fill_1 FILLER_44_2355 ();
 sg13g2_fill_2 FILLER_44_2386 ();
 sg13g2_fill_1 FILLER_44_2402 ();
 sg13g2_fill_2 FILLER_44_2411 ();
 sg13g2_fill_1 FILLER_44_2418 ();
 sg13g2_fill_1 FILLER_44_2424 ();
 sg13g2_decap_4 FILLER_44_2435 ();
 sg13g2_fill_2 FILLER_44_2443 ();
 sg13g2_fill_1 FILLER_44_2445 ();
 sg13g2_fill_1 FILLER_44_2452 ();
 sg13g2_fill_2 FILLER_44_2463 ();
 sg13g2_decap_4 FILLER_44_2484 ();
 sg13g2_fill_1 FILLER_44_2488 ();
 sg13g2_fill_2 FILLER_44_2503 ();
 sg13g2_fill_2 FILLER_44_2548 ();
 sg13g2_fill_1 FILLER_44_2589 ();
 sg13g2_fill_2 FILLER_44_2629 ();
 sg13g2_fill_1 FILLER_44_2641 ();
 sg13g2_fill_2 FILLER_44_2668 ();
 sg13g2_decap_8 FILLER_45_0 ();
 sg13g2_fill_2 FILLER_45_7 ();
 sg13g2_fill_1 FILLER_45_9 ();
 sg13g2_fill_1 FILLER_45_27 ();
 sg13g2_fill_1 FILLER_45_33 ();
 sg13g2_decap_8 FILLER_45_47 ();
 sg13g2_decap_4 FILLER_45_59 ();
 sg13g2_fill_1 FILLER_45_63 ();
 sg13g2_fill_1 FILLER_45_69 ();
 sg13g2_fill_1 FILLER_45_74 ();
 sg13g2_fill_1 FILLER_45_92 ();
 sg13g2_fill_1 FILLER_45_98 ();
 sg13g2_fill_1 FILLER_45_108 ();
 sg13g2_fill_1 FILLER_45_140 ();
 sg13g2_fill_2 FILLER_45_150 ();
 sg13g2_fill_2 FILLER_45_190 ();
 sg13g2_fill_2 FILLER_45_196 ();
 sg13g2_fill_1 FILLER_45_208 ();
 sg13g2_fill_1 FILLER_45_233 ();
 sg13g2_fill_2 FILLER_45_239 ();
 sg13g2_decap_4 FILLER_45_249 ();
 sg13g2_fill_1 FILLER_45_253 ();
 sg13g2_fill_1 FILLER_45_258 ();
 sg13g2_decap_8 FILLER_45_262 ();
 sg13g2_fill_2 FILLER_45_269 ();
 sg13g2_fill_1 FILLER_45_271 ();
 sg13g2_decap_4 FILLER_45_276 ();
 sg13g2_fill_1 FILLER_45_280 ();
 sg13g2_fill_1 FILLER_45_286 ();
 sg13g2_decap_4 FILLER_45_302 ();
 sg13g2_fill_1 FILLER_45_325 ();
 sg13g2_fill_2 FILLER_45_357 ();
 sg13g2_fill_1 FILLER_45_384 ();
 sg13g2_fill_1 FILLER_45_395 ();
 sg13g2_decap_4 FILLER_45_426 ();
 sg13g2_fill_2 FILLER_45_430 ();
 sg13g2_fill_2 FILLER_45_442 ();
 sg13g2_fill_2 FILLER_45_466 ();
 sg13g2_fill_2 FILLER_45_477 ();
 sg13g2_fill_2 FILLER_45_483 ();
 sg13g2_fill_1 FILLER_45_489 ();
 sg13g2_fill_1 FILLER_45_494 ();
 sg13g2_fill_2 FILLER_45_498 ();
 sg13g2_fill_2 FILLER_45_524 ();
 sg13g2_fill_1 FILLER_45_526 ();
 sg13g2_fill_1 FILLER_45_531 ();
 sg13g2_decap_4 FILLER_45_537 ();
 sg13g2_decap_4 FILLER_45_546 ();
 sg13g2_fill_1 FILLER_45_550 ();
 sg13g2_decap_8 FILLER_45_557 ();
 sg13g2_fill_2 FILLER_45_564 ();
 sg13g2_fill_1 FILLER_45_566 ();
 sg13g2_fill_2 FILLER_45_571 ();
 sg13g2_fill_1 FILLER_45_573 ();
 sg13g2_fill_1 FILLER_45_588 ();
 sg13g2_fill_2 FILLER_45_602 ();
 sg13g2_fill_1 FILLER_45_604 ();
 sg13g2_fill_1 FILLER_45_671 ();
 sg13g2_fill_1 FILLER_45_687 ();
 sg13g2_fill_1 FILLER_45_729 ();
 sg13g2_fill_2 FILLER_45_786 ();
 sg13g2_fill_1 FILLER_45_788 ();
 sg13g2_fill_1 FILLER_45_850 ();
 sg13g2_fill_1 FILLER_45_896 ();
 sg13g2_fill_1 FILLER_45_934 ();
 sg13g2_decap_8 FILLER_45_1022 ();
 sg13g2_decap_8 FILLER_45_1029 ();
 sg13g2_fill_1 FILLER_45_1079 ();
 sg13g2_fill_1 FILLER_45_1090 ();
 sg13g2_fill_1 FILLER_45_1127 ();
 sg13g2_fill_1 FILLER_45_1199 ();
 sg13g2_fill_2 FILLER_45_1285 ();
 sg13g2_decap_4 FILLER_45_1298 ();
 sg13g2_decap_4 FILLER_45_1308 ();
 sg13g2_fill_1 FILLER_45_1312 ();
 sg13g2_fill_2 FILLER_45_1317 ();
 sg13g2_fill_1 FILLER_45_1344 ();
 sg13g2_fill_2 FILLER_45_1351 ();
 sg13g2_decap_8 FILLER_45_1363 ();
 sg13g2_decap_4 FILLER_45_1370 ();
 sg13g2_fill_1 FILLER_45_1416 ();
 sg13g2_fill_2 FILLER_45_1426 ();
 sg13g2_fill_1 FILLER_45_1440 ();
 sg13g2_fill_2 FILLER_45_1488 ();
 sg13g2_fill_2 FILLER_45_1520 ();
 sg13g2_fill_1 FILLER_45_1531 ();
 sg13g2_fill_1 FILLER_45_1542 ();
 sg13g2_fill_2 FILLER_45_1548 ();
 sg13g2_fill_2 FILLER_45_1556 ();
 sg13g2_decap_8 FILLER_45_1575 ();
 sg13g2_fill_1 FILLER_45_1604 ();
 sg13g2_decap_4 FILLER_45_1623 ();
 sg13g2_decap_8 FILLER_45_1631 ();
 sg13g2_decap_8 FILLER_45_1638 ();
 sg13g2_decap_8 FILLER_45_1645 ();
 sg13g2_decap_4 FILLER_45_1652 ();
 sg13g2_fill_2 FILLER_45_1656 ();
 sg13g2_decap_8 FILLER_45_1694 ();
 sg13g2_decap_8 FILLER_45_1701 ();
 sg13g2_decap_4 FILLER_45_1708 ();
 sg13g2_decap_8 FILLER_45_1717 ();
 sg13g2_fill_1 FILLER_45_1724 ();
 sg13g2_decap_4 FILLER_45_1734 ();
 sg13g2_fill_1 FILLER_45_1738 ();
 sg13g2_decap_8 FILLER_45_1760 ();
 sg13g2_decap_8 FILLER_45_1767 ();
 sg13g2_decap_4 FILLER_45_1778 ();
 sg13g2_decap_8 FILLER_45_1786 ();
 sg13g2_fill_1 FILLER_45_1872 ();
 sg13g2_fill_1 FILLER_45_1877 ();
 sg13g2_fill_1 FILLER_45_1886 ();
 sg13g2_decap_8 FILLER_45_1897 ();
 sg13g2_decap_8 FILLER_45_1904 ();
 sg13g2_fill_1 FILLER_45_1916 ();
 sg13g2_fill_1 FILLER_45_1949 ();
 sg13g2_fill_2 FILLER_45_1958 ();
 sg13g2_fill_1 FILLER_45_1978 ();
 sg13g2_fill_1 FILLER_45_2001 ();
 sg13g2_fill_1 FILLER_45_2006 ();
 sg13g2_decap_8 FILLER_45_2035 ();
 sg13g2_decap_4 FILLER_45_2042 ();
 sg13g2_fill_2 FILLER_45_2046 ();
 sg13g2_decap_8 FILLER_45_2052 ();
 sg13g2_decap_4 FILLER_45_2059 ();
 sg13g2_fill_2 FILLER_45_2063 ();
 sg13g2_decap_4 FILLER_45_2119 ();
 sg13g2_fill_2 FILLER_45_2123 ();
 sg13g2_fill_2 FILLER_45_2150 ();
 sg13g2_fill_1 FILLER_45_2152 ();
 sg13g2_decap_8 FILLER_45_2188 ();
 sg13g2_fill_1 FILLER_45_2221 ();
 sg13g2_fill_2 FILLER_45_2232 ();
 sg13g2_fill_1 FILLER_45_2267 ();
 sg13g2_fill_1 FILLER_45_2272 ();
 sg13g2_fill_1 FILLER_45_2283 ();
 sg13g2_fill_1 FILLER_45_2288 ();
 sg13g2_decap_4 FILLER_45_2299 ();
 sg13g2_fill_2 FILLER_45_2303 ();
 sg13g2_fill_2 FILLER_45_2324 ();
 sg13g2_fill_2 FILLER_45_2340 ();
 sg13g2_decap_8 FILLER_45_2348 ();
 sg13g2_decap_8 FILLER_45_2355 ();
 sg13g2_fill_1 FILLER_45_2367 ();
 sg13g2_fill_2 FILLER_45_2372 ();
 sg13g2_fill_1 FILLER_45_2395 ();
 sg13g2_fill_1 FILLER_45_2404 ();
 sg13g2_decap_8 FILLER_45_2412 ();
 sg13g2_decap_4 FILLER_45_2419 ();
 sg13g2_fill_1 FILLER_45_2423 ();
 sg13g2_decap_4 FILLER_45_2470 ();
 sg13g2_fill_2 FILLER_45_2522 ();
 sg13g2_fill_1 FILLER_45_2524 ();
 sg13g2_fill_1 FILLER_45_2531 ();
 sg13g2_fill_1 FILLER_45_2548 ();
 sg13g2_fill_2 FILLER_45_2575 ();
 sg13g2_fill_2 FILLER_45_2582 ();
 sg13g2_fill_2 FILLER_45_2596 ();
 sg13g2_fill_1 FILLER_45_2625 ();
 sg13g2_fill_2 FILLER_45_2651 ();
 sg13g2_fill_1 FILLER_45_2669 ();
 sg13g2_decap_8 FILLER_46_0 ();
 sg13g2_fill_2 FILLER_46_7 ();
 sg13g2_fill_1 FILLER_46_23 ();
 sg13g2_fill_1 FILLER_46_32 ();
 sg13g2_decap_8 FILLER_46_50 ();
 sg13g2_decap_4 FILLER_46_57 ();
 sg13g2_fill_1 FILLER_46_92 ();
 sg13g2_fill_1 FILLER_46_97 ();
 sg13g2_fill_2 FILLER_46_102 ();
 sg13g2_fill_1 FILLER_46_104 ();
 sg13g2_fill_1 FILLER_46_110 ();
 sg13g2_fill_2 FILLER_46_194 ();
 sg13g2_fill_1 FILLER_46_224 ();
 sg13g2_fill_2 FILLER_46_239 ();
 sg13g2_decap_8 FILLER_46_246 ();
 sg13g2_decap_8 FILLER_46_253 ();
 sg13g2_decap_8 FILLER_46_260 ();
 sg13g2_decap_8 FILLER_46_267 ();
 sg13g2_fill_2 FILLER_46_274 ();
 sg13g2_fill_1 FILLER_46_286 ();
 sg13g2_fill_1 FILLER_46_338 ();
 sg13g2_fill_1 FILLER_46_402 ();
 sg13g2_fill_2 FILLER_46_406 ();
 sg13g2_fill_2 FILLER_46_444 ();
 sg13g2_fill_2 FILLER_46_476 ();
 sg13g2_fill_2 FILLER_46_513 ();
 sg13g2_fill_2 FILLER_46_520 ();
 sg13g2_decap_4 FILLER_46_535 ();
 sg13g2_fill_1 FILLER_46_539 ();
 sg13g2_decap_8 FILLER_46_545 ();
 sg13g2_decap_8 FILLER_46_552 ();
 sg13g2_decap_4 FILLER_46_559 ();
 sg13g2_fill_1 FILLER_46_563 ();
 sg13g2_fill_2 FILLER_46_573 ();
 sg13g2_fill_1 FILLER_46_580 ();
 sg13g2_fill_1 FILLER_46_590 ();
 sg13g2_fill_2 FILLER_46_617 ();
 sg13g2_fill_2 FILLER_46_637 ();
 sg13g2_fill_2 FILLER_46_660 ();
 sg13g2_fill_2 FILLER_46_670 ();
 sg13g2_decap_8 FILLER_46_686 ();
 sg13g2_fill_2 FILLER_46_693 ();
 sg13g2_fill_1 FILLER_46_695 ();
 sg13g2_decap_4 FILLER_46_700 ();
 sg13g2_fill_2 FILLER_46_718 ();
 sg13g2_fill_2 FILLER_46_774 ();
 sg13g2_fill_1 FILLER_46_785 ();
 sg13g2_decap_4 FILLER_46_803 ();
 sg13g2_fill_1 FILLER_46_823 ();
 sg13g2_fill_2 FILLER_46_828 ();
 sg13g2_fill_1 FILLER_46_842 ();
 sg13g2_fill_2 FILLER_46_909 ();
 sg13g2_fill_2 FILLER_46_943 ();
 sg13g2_fill_2 FILLER_46_971 ();
 sg13g2_fill_1 FILLER_46_997 ();
 sg13g2_decap_8 FILLER_46_1034 ();
 sg13g2_decap_8 FILLER_46_1041 ();
 sg13g2_decap_4 FILLER_46_1048 ();
 sg13g2_fill_1 FILLER_46_1052 ();
 sg13g2_fill_2 FILLER_46_1057 ();
 sg13g2_fill_2 FILLER_46_1064 ();
 sg13g2_fill_1 FILLER_46_1112 ();
 sg13g2_fill_2 FILLER_46_1132 ();
 sg13g2_fill_1 FILLER_46_1170 ();
 sg13g2_fill_1 FILLER_46_1229 ();
 sg13g2_fill_2 FILLER_46_1290 ();
 sg13g2_fill_2 FILLER_46_1296 ();
 sg13g2_fill_1 FILLER_46_1303 ();
 sg13g2_fill_2 FILLER_46_1314 ();
 sg13g2_fill_1 FILLER_46_1316 ();
 sg13g2_decap_8 FILLER_46_1343 ();
 sg13g2_fill_2 FILLER_46_1350 ();
 sg13g2_decap_4 FILLER_46_1364 ();
 sg13g2_fill_2 FILLER_46_1373 ();
 sg13g2_fill_1 FILLER_46_1375 ();
 sg13g2_decap_4 FILLER_46_1387 ();
 sg13g2_fill_2 FILLER_46_1391 ();
 sg13g2_decap_8 FILLER_46_1403 ();
 sg13g2_fill_2 FILLER_46_1410 ();
 sg13g2_fill_1 FILLER_46_1500 ();
 sg13g2_fill_1 FILLER_46_1513 ();
 sg13g2_fill_2 FILLER_46_1519 ();
 sg13g2_decap_8 FILLER_46_1550 ();
 sg13g2_fill_2 FILLER_46_1557 ();
 sg13g2_decap_8 FILLER_46_1563 ();
 sg13g2_fill_2 FILLER_46_1570 ();
 sg13g2_decap_8 FILLER_46_1577 ();
 sg13g2_fill_1 FILLER_46_1584 ();
 sg13g2_fill_1 FILLER_46_1589 ();
 sg13g2_fill_2 FILLER_46_1604 ();
 sg13g2_decap_8 FILLER_46_1624 ();
 sg13g2_decap_4 FILLER_46_1631 ();
 sg13g2_decap_8 FILLER_46_1640 ();
 sg13g2_fill_1 FILLER_46_1647 ();
 sg13g2_decap_4 FILLER_46_1660 ();
 sg13g2_fill_1 FILLER_46_1664 ();
 sg13g2_decap_8 FILLER_46_1694 ();
 sg13g2_fill_2 FILLER_46_1701 ();
 sg13g2_fill_1 FILLER_46_1703 ();
 sg13g2_fill_1 FILLER_46_1714 ();
 sg13g2_decap_8 FILLER_46_1719 ();
 sg13g2_decap_8 FILLER_46_1726 ();
 sg13g2_decap_8 FILLER_46_1733 ();
 sg13g2_decap_8 FILLER_46_1740 ();
 sg13g2_fill_2 FILLER_46_1747 ();
 sg13g2_fill_2 FILLER_46_1762 ();
 sg13g2_decap_4 FILLER_46_1800 ();
 sg13g2_decap_8 FILLER_46_1808 ();
 sg13g2_decap_4 FILLER_46_1815 ();
 sg13g2_fill_1 FILLER_46_1819 ();
 sg13g2_decap_8 FILLER_46_1831 ();
 sg13g2_fill_2 FILLER_46_1843 ();
 sg13g2_fill_1 FILLER_46_1857 ();
 sg13g2_decap_8 FILLER_46_1900 ();
 sg13g2_fill_1 FILLER_46_1915 ();
 sg13g2_fill_2 FILLER_46_1930 ();
 sg13g2_fill_1 FILLER_46_1932 ();
 sg13g2_decap_4 FILLER_46_1937 ();
 sg13g2_fill_1 FILLER_46_1945 ();
 sg13g2_fill_2 FILLER_46_1951 ();
 sg13g2_fill_1 FILLER_46_1953 ();
 sg13g2_fill_2 FILLER_46_1963 ();
 sg13g2_fill_1 FILLER_46_2015 ();
 sg13g2_decap_8 FILLER_46_2039 ();
 sg13g2_decap_8 FILLER_46_2046 ();
 sg13g2_decap_8 FILLER_46_2053 ();
 sg13g2_decap_8 FILLER_46_2060 ();
 sg13g2_decap_8 FILLER_46_2067 ();
 sg13g2_fill_2 FILLER_46_2074 ();
 sg13g2_decap_4 FILLER_46_2112 ();
 sg13g2_fill_2 FILLER_46_2116 ();
 sg13g2_decap_8 FILLER_46_2144 ();
 sg13g2_decap_4 FILLER_46_2151 ();
 sg13g2_fill_2 FILLER_46_2155 ();
 sg13g2_fill_1 FILLER_46_2213 ();
 sg13g2_decap_4 FILLER_46_2248 ();
 sg13g2_fill_1 FILLER_46_2252 ();
 sg13g2_fill_1 FILLER_46_2263 ();
 sg13g2_fill_1 FILLER_46_2307 ();
 sg13g2_fill_1 FILLER_46_2317 ();
 sg13g2_decap_8 FILLER_46_2329 ();
 sg13g2_decap_8 FILLER_46_2336 ();
 sg13g2_decap_8 FILLER_46_2343 ();
 sg13g2_decap_8 FILLER_46_2350 ();
 sg13g2_decap_4 FILLER_46_2357 ();
 sg13g2_fill_1 FILLER_46_2361 ();
 sg13g2_decap_4 FILLER_46_2428 ();
 sg13g2_fill_1 FILLER_46_2432 ();
 sg13g2_fill_2 FILLER_46_2438 ();
 sg13g2_decap_8 FILLER_46_2444 ();
 sg13g2_fill_2 FILLER_46_2451 ();
 sg13g2_decap_4 FILLER_46_2458 ();
 sg13g2_decap_8 FILLER_46_2488 ();
 sg13g2_decap_8 FILLER_46_2495 ();
 sg13g2_fill_1 FILLER_46_2502 ();
 sg13g2_fill_1 FILLER_46_2509 ();
 sg13g2_fill_2 FILLER_46_2530 ();
 sg13g2_fill_2 FILLER_46_2540 ();
 sg13g2_decap_8 FILLER_46_2561 ();
 sg13g2_fill_2 FILLER_46_2568 ();
 sg13g2_fill_1 FILLER_46_2594 ();
 sg13g2_fill_2 FILLER_46_2647 ();
 sg13g2_decap_8 FILLER_46_2656 ();
 sg13g2_decap_8 FILLER_46_2663 ();
 sg13g2_fill_1 FILLER_47_0 ();
 sg13g2_fill_1 FILLER_47_32 ();
 sg13g2_fill_1 FILLER_47_38 ();
 sg13g2_decap_8 FILLER_47_86 ();
 sg13g2_decap_8 FILLER_47_93 ();
 sg13g2_fill_1 FILLER_47_109 ();
 sg13g2_fill_1 FILLER_47_131 ();
 sg13g2_fill_1 FILLER_47_152 ();
 sg13g2_fill_1 FILLER_47_162 ();
 sg13g2_decap_8 FILLER_47_236 ();
 sg13g2_decap_4 FILLER_47_251 ();
 sg13g2_decap_4 FILLER_47_291 ();
 sg13g2_fill_2 FILLER_47_325 ();
 sg13g2_fill_1 FILLER_47_327 ();
 sg13g2_fill_2 FILLER_47_337 ();
 sg13g2_fill_1 FILLER_47_339 ();
 sg13g2_fill_2 FILLER_47_350 ();
 sg13g2_fill_1 FILLER_47_357 ();
 sg13g2_fill_2 FILLER_47_444 ();
 sg13g2_fill_2 FILLER_47_449 ();
 sg13g2_fill_1 FILLER_47_520 ();
 sg13g2_decap_8 FILLER_47_547 ();
 sg13g2_decap_4 FILLER_47_554 ();
 sg13g2_fill_2 FILLER_47_568 ();
 sg13g2_fill_1 FILLER_47_570 ();
 sg13g2_fill_2 FILLER_47_584 ();
 sg13g2_fill_2 FILLER_47_601 ();
 sg13g2_decap_4 FILLER_47_609 ();
 sg13g2_fill_2 FILLER_47_655 ();
 sg13g2_fill_2 FILLER_47_687 ();
 sg13g2_decap_4 FILLER_47_693 ();
 sg13g2_fill_2 FILLER_47_701 ();
 sg13g2_decap_8 FILLER_47_715 ();
 sg13g2_decap_8 FILLER_47_722 ();
 sg13g2_decap_8 FILLER_47_729 ();
 sg13g2_fill_1 FILLER_47_736 ();
 sg13g2_fill_2 FILLER_47_750 ();
 sg13g2_fill_2 FILLER_47_757 ();
 sg13g2_fill_1 FILLER_47_759 ();
 sg13g2_fill_2 FILLER_47_768 ();
 sg13g2_fill_1 FILLER_47_792 ();
 sg13g2_fill_1 FILLER_47_800 ();
 sg13g2_fill_2 FILLER_47_818 ();
 sg13g2_fill_1 FILLER_47_884 ();
 sg13g2_fill_1 FILLER_47_914 ();
 sg13g2_fill_1 FILLER_47_919 ();
 sg13g2_fill_1 FILLER_47_984 ();
 sg13g2_fill_2 FILLER_47_993 ();
 sg13g2_decap_8 FILLER_47_1036 ();
 sg13g2_fill_2 FILLER_47_1043 ();
 sg13g2_fill_1 FILLER_47_1045 ();
 sg13g2_fill_1 FILLER_47_1050 ();
 sg13g2_fill_2 FILLER_47_1090 ();
 sg13g2_fill_1 FILLER_47_1103 ();
 sg13g2_fill_2 FILLER_47_1114 ();
 sg13g2_fill_1 FILLER_47_1179 ();
 sg13g2_fill_1 FILLER_47_1188 ();
 sg13g2_fill_2 FILLER_47_1198 ();
 sg13g2_fill_2 FILLER_47_1231 ();
 sg13g2_fill_1 FILLER_47_1233 ();
 sg13g2_fill_1 FILLER_47_1240 ();
 sg13g2_fill_2 FILLER_47_1274 ();
 sg13g2_decap_4 FILLER_47_1284 ();
 sg13g2_fill_1 FILLER_47_1288 ();
 sg13g2_fill_1 FILLER_47_1299 ();
 sg13g2_fill_1 FILLER_47_1312 ();
 sg13g2_fill_1 FILLER_47_1320 ();
 sg13g2_fill_1 FILLER_47_1336 ();
 sg13g2_decap_4 FILLER_47_1342 ();
 sg13g2_fill_2 FILLER_47_1346 ();
 sg13g2_decap_4 FILLER_47_1352 ();
 sg13g2_fill_2 FILLER_47_1369 ();
 sg13g2_fill_1 FILLER_47_1371 ();
 sg13g2_fill_1 FILLER_47_1391 ();
 sg13g2_decap_8 FILLER_47_1397 ();
 sg13g2_decap_4 FILLER_47_1404 ();
 sg13g2_fill_1 FILLER_47_1408 ();
 sg13g2_fill_2 FILLER_47_1415 ();
 sg13g2_fill_1 FILLER_47_1422 ();
 sg13g2_fill_1 FILLER_47_1432 ();
 sg13g2_fill_2 FILLER_47_1446 ();
 sg13g2_fill_2 FILLER_47_1459 ();
 sg13g2_fill_1 FILLER_47_1466 ();
 sg13g2_fill_1 FILLER_47_1496 ();
 sg13g2_fill_1 FILLER_47_1503 ();
 sg13g2_fill_1 FILLER_47_1543 ();
 sg13g2_decap_8 FILLER_47_1565 ();
 sg13g2_fill_1 FILLER_47_1572 ();
 sg13g2_fill_2 FILLER_47_1579 ();
 sg13g2_fill_1 FILLER_47_1584 ();
 sg13g2_fill_1 FILLER_47_1598 ();
 sg13g2_fill_1 FILLER_47_1617 ();
 sg13g2_fill_2 FILLER_47_1644 ();
 sg13g2_fill_1 FILLER_47_1651 ();
 sg13g2_fill_1 FILLER_47_1658 ();
 sg13g2_fill_2 FILLER_47_1669 ();
 sg13g2_fill_1 FILLER_47_1671 ();
 sg13g2_fill_2 FILLER_47_1676 ();
 sg13g2_fill_1 FILLER_47_1678 ();
 sg13g2_fill_1 FILLER_47_1684 ();
 sg13g2_fill_1 FILLER_47_1696 ();
 sg13g2_fill_2 FILLER_47_1728 ();
 sg13g2_fill_1 FILLER_47_1730 ();
 sg13g2_fill_1 FILLER_47_1735 ();
 sg13g2_fill_1 FILLER_47_1751 ();
 sg13g2_fill_1 FILLER_47_1760 ();
 sg13g2_fill_1 FILLER_47_1765 ();
 sg13g2_fill_1 FILLER_47_1776 ();
 sg13g2_fill_2 FILLER_47_1787 ();
 sg13g2_decap_8 FILLER_47_1797 ();
 sg13g2_decap_8 FILLER_47_1804 ();
 sg13g2_decap_8 FILLER_47_1811 ();
 sg13g2_decap_4 FILLER_47_1818 ();
 sg13g2_decap_4 FILLER_47_1826 ();
 sg13g2_fill_2 FILLER_47_1830 ();
 sg13g2_decap_4 FILLER_47_1837 ();
 sg13g2_fill_1 FILLER_47_1841 ();
 sg13g2_fill_2 FILLER_47_1846 ();
 sg13g2_fill_2 FILLER_47_1853 ();
 sg13g2_fill_2 FILLER_47_1864 ();
 sg13g2_decap_4 FILLER_47_1876 ();
 sg13g2_fill_1 FILLER_47_1880 ();
 sg13g2_fill_2 FILLER_47_1899 ();
 sg13g2_decap_8 FILLER_47_1944 ();
 sg13g2_fill_2 FILLER_47_1951 ();
 sg13g2_fill_1 FILLER_47_1953 ();
 sg13g2_decap_8 FILLER_47_1958 ();
 sg13g2_fill_2 FILLER_47_1965 ();
 sg13g2_fill_1 FILLER_47_1995 ();
 sg13g2_fill_2 FILLER_47_2014 ();
 sg13g2_fill_1 FILLER_47_2021 ();
 sg13g2_decap_4 FILLER_47_2040 ();
 sg13g2_fill_2 FILLER_47_2048 ();
 sg13g2_fill_1 FILLER_47_2050 ();
 sg13g2_decap_4 FILLER_47_2059 ();
 sg13g2_fill_1 FILLER_47_2068 ();
 sg13g2_decap_8 FILLER_47_2077 ();
 sg13g2_decap_8 FILLER_47_2084 ();
 sg13g2_fill_2 FILLER_47_2091 ();
 sg13g2_fill_2 FILLER_47_2097 ();
 sg13g2_fill_2 FILLER_47_2156 ();
 sg13g2_fill_1 FILLER_47_2158 ();
 sg13g2_fill_1 FILLER_47_2199 ();
 sg13g2_fill_2 FILLER_47_2227 ();
 sg13g2_fill_1 FILLER_47_2259 ();
 sg13g2_fill_2 FILLER_47_2263 ();
 sg13g2_fill_1 FILLER_47_2278 ();
 sg13g2_fill_1 FILLER_47_2286 ();
 sg13g2_decap_8 FILLER_47_2340 ();
 sg13g2_fill_2 FILLER_47_2433 ();
 sg13g2_decap_4 FILLER_47_2439 ();
 sg13g2_fill_2 FILLER_47_2447 ();
 sg13g2_decap_4 FILLER_47_2466 ();
 sg13g2_fill_1 FILLER_47_2470 ();
 sg13g2_fill_2 FILLER_47_2475 ();
 sg13g2_fill_1 FILLER_47_2488 ();
 sg13g2_fill_2 FILLER_47_2503 ();
 sg13g2_fill_1 FILLER_47_2505 ();
 sg13g2_fill_1 FILLER_47_2535 ();
 sg13g2_fill_1 FILLER_47_2549 ();
 sg13g2_decap_8 FILLER_47_2566 ();
 sg13g2_decap_4 FILLER_47_2573 ();
 sg13g2_fill_1 FILLER_47_2587 ();
 sg13g2_fill_1 FILLER_47_2592 ();
 sg13g2_fill_1 FILLER_47_2596 ();
 sg13g2_fill_2 FILLER_47_2640 ();
 sg13g2_fill_2 FILLER_47_2668 ();
 sg13g2_fill_2 FILLER_48_0 ();
 sg13g2_fill_1 FILLER_48_2 ();
 sg13g2_fill_2 FILLER_48_11 ();
 sg13g2_fill_1 FILLER_48_13 ();
 sg13g2_fill_2 FILLER_48_22 ();
 sg13g2_decap_4 FILLER_48_59 ();
 sg13g2_decap_4 FILLER_48_90 ();
 sg13g2_fill_1 FILLER_48_94 ();
 sg13g2_fill_2 FILLER_48_121 ();
 sg13g2_fill_2 FILLER_48_128 ();
 sg13g2_fill_1 FILLER_48_170 ();
 sg13g2_fill_1 FILLER_48_176 ();
 sg13g2_fill_1 FILLER_48_203 ();
 sg13g2_fill_1 FILLER_48_209 ();
 sg13g2_fill_2 FILLER_48_219 ();
 sg13g2_fill_2 FILLER_48_258 ();
 sg13g2_decap_4 FILLER_48_268 ();
 sg13g2_fill_1 FILLER_48_272 ();
 sg13g2_decap_4 FILLER_48_281 ();
 sg13g2_fill_1 FILLER_48_324 ();
 sg13g2_fill_2 FILLER_48_339 ();
 sg13g2_fill_1 FILLER_48_368 ();
 sg13g2_fill_2 FILLER_48_438 ();
 sg13g2_fill_1 FILLER_48_451 ();
 sg13g2_fill_1 FILLER_48_484 ();
 sg13g2_fill_1 FILLER_48_495 ();
 sg13g2_fill_1 FILLER_48_512 ();
 sg13g2_fill_1 FILLER_48_523 ();
 sg13g2_fill_1 FILLER_48_538 ();
 sg13g2_decap_8 FILLER_48_549 ();
 sg13g2_decap_4 FILLER_48_556 ();
 sg13g2_fill_2 FILLER_48_564 ();
 sg13g2_fill_2 FILLER_48_586 ();
 sg13g2_fill_2 FILLER_48_593 ();
 sg13g2_fill_1 FILLER_48_595 ();
 sg13g2_fill_1 FILLER_48_606 ();
 sg13g2_fill_1 FILLER_48_618 ();
 sg13g2_fill_1 FILLER_48_638 ();
 sg13g2_decap_4 FILLER_48_668 ();
 sg13g2_decap_8 FILLER_48_685 ();
 sg13g2_decap_8 FILLER_48_692 ();
 sg13g2_fill_2 FILLER_48_699 ();
 sg13g2_fill_1 FILLER_48_701 ();
 sg13g2_decap_8 FILLER_48_715 ();
 sg13g2_decap_8 FILLER_48_722 ();
 sg13g2_decap_8 FILLER_48_729 ();
 sg13g2_decap_8 FILLER_48_736 ();
 sg13g2_fill_1 FILLER_48_743 ();
 sg13g2_fill_2 FILLER_48_748 ();
 sg13g2_fill_1 FILLER_48_790 ();
 sg13g2_fill_1 FILLER_48_794 ();
 sg13g2_fill_1 FILLER_48_844 ();
 sg13g2_fill_1 FILLER_48_860 ();
 sg13g2_fill_1 FILLER_48_871 ();
 sg13g2_fill_2 FILLER_48_973 ();
 sg13g2_fill_1 FILLER_48_989 ();
 sg13g2_fill_2 FILLER_48_1031 ();
 sg13g2_fill_2 FILLER_48_1043 ();
 sg13g2_fill_1 FILLER_48_1128 ();
 sg13g2_fill_2 FILLER_48_1132 ();
 sg13g2_fill_2 FILLER_48_1163 ();
 sg13g2_fill_1 FILLER_48_1165 ();
 sg13g2_decap_4 FILLER_48_1179 ();
 sg13g2_fill_2 FILLER_48_1183 ();
 sg13g2_fill_2 FILLER_48_1205 ();
 sg13g2_fill_1 FILLER_48_1207 ();
 sg13g2_fill_2 FILLER_48_1256 ();
 sg13g2_fill_1 FILLER_48_1258 ();
 sg13g2_fill_2 FILLER_48_1263 ();
 sg13g2_fill_1 FILLER_48_1265 ();
 sg13g2_fill_2 FILLER_48_1271 ();
 sg13g2_fill_1 FILLER_48_1273 ();
 sg13g2_decap_4 FILLER_48_1284 ();
 sg13g2_fill_1 FILLER_48_1288 ();
 sg13g2_fill_1 FILLER_48_1294 ();
 sg13g2_fill_2 FILLER_48_1299 ();
 sg13g2_decap_8 FILLER_48_1327 ();
 sg13g2_decap_4 FILLER_48_1334 ();
 sg13g2_fill_1 FILLER_48_1338 ();
 sg13g2_fill_2 FILLER_48_1360 ();
 sg13g2_fill_2 FILLER_48_1391 ();
 sg13g2_fill_1 FILLER_48_1398 ();
 sg13g2_fill_1 FILLER_48_1407 ();
 sg13g2_fill_1 FILLER_48_1449 ();
 sg13g2_fill_1 FILLER_48_1471 ();
 sg13g2_fill_2 FILLER_48_1512 ();
 sg13g2_decap_4 FILLER_48_1576 ();
 sg13g2_fill_1 FILLER_48_1601 ();
 sg13g2_fill_1 FILLER_48_1611 ();
 sg13g2_decap_4 FILLER_48_1627 ();
 sg13g2_fill_2 FILLER_48_1631 ();
 sg13g2_fill_1 FILLER_48_1668 ();
 sg13g2_fill_1 FILLER_48_1679 ();
 sg13g2_fill_1 FILLER_48_1723 ();
 sg13g2_fill_1 FILLER_48_1739 ();
 sg13g2_decap_4 FILLER_48_1753 ();
 sg13g2_fill_1 FILLER_48_1764 ();
 sg13g2_fill_2 FILLER_48_1770 ();
 sg13g2_fill_1 FILLER_48_1772 ();
 sg13g2_fill_2 FILLER_48_1778 ();
 sg13g2_fill_1 FILLER_48_1780 ();
 sg13g2_fill_1 FILLER_48_1807 ();
 sg13g2_fill_2 FILLER_48_1833 ();
 sg13g2_fill_1 FILLER_48_1835 ();
 sg13g2_fill_1 FILLER_48_1842 ();
 sg13g2_fill_1 FILLER_48_1852 ();
 sg13g2_fill_1 FILLER_48_1859 ();
 sg13g2_fill_2 FILLER_48_1893 ();
 sg13g2_fill_2 FILLER_48_1900 ();
 sg13g2_decap_4 FILLER_48_1926 ();
 sg13g2_fill_1 FILLER_48_1930 ();
 sg13g2_fill_2 FILLER_48_1934 ();
 sg13g2_fill_1 FILLER_48_1941 ();
 sg13g2_fill_1 FILLER_48_1966 ();
 sg13g2_fill_2 FILLER_48_1976 ();
 sg13g2_decap_4 FILLER_48_2018 ();
 sg13g2_fill_1 FILLER_48_2022 ();
 sg13g2_decap_8 FILLER_48_2032 ();
 sg13g2_decap_4 FILLER_48_2044 ();
 sg13g2_fill_1 FILLER_48_2052 ();
 sg13g2_fill_2 FILLER_48_2066 ();
 sg13g2_fill_2 FILLER_48_2078 ();
 sg13g2_fill_2 FILLER_48_2085 ();
 sg13g2_fill_1 FILLER_48_2087 ();
 sg13g2_decap_8 FILLER_48_2092 ();
 sg13g2_fill_1 FILLER_48_2099 ();
 sg13g2_decap_8 FILLER_48_2149 ();
 sg13g2_decap_4 FILLER_48_2156 ();
 sg13g2_fill_2 FILLER_48_2160 ();
 sg13g2_decap_8 FILLER_48_2166 ();
 sg13g2_fill_2 FILLER_48_2173 ();
 sg13g2_decap_8 FILLER_48_2179 ();
 sg13g2_decap_8 FILLER_48_2186 ();
 sg13g2_decap_4 FILLER_48_2193 ();
 sg13g2_fill_2 FILLER_48_2197 ();
 sg13g2_fill_2 FILLER_48_2202 ();
 sg13g2_fill_1 FILLER_48_2210 ();
 sg13g2_fill_2 FILLER_48_2258 ();
 sg13g2_fill_2 FILLER_48_2263 ();
 sg13g2_fill_1 FILLER_48_2340 ();
 sg13g2_fill_2 FILLER_48_2372 ();
 sg13g2_fill_1 FILLER_48_2380 ();
 sg13g2_decap_4 FILLER_48_2386 ();
 sg13g2_fill_2 FILLER_48_2390 ();
 sg13g2_fill_1 FILLER_48_2606 ();
 sg13g2_fill_2 FILLER_48_2668 ();
 sg13g2_fill_1 FILLER_49_0 ();
 sg13g2_decap_8 FILLER_49_27 ();
 sg13g2_fill_2 FILLER_49_34 ();
 sg13g2_fill_1 FILLER_49_36 ();
 sg13g2_decap_4 FILLER_49_41 ();
 sg13g2_fill_1 FILLER_49_45 ();
 sg13g2_fill_1 FILLER_49_80 ();
 sg13g2_fill_1 FILLER_49_101 ();
 sg13g2_fill_2 FILLER_49_110 ();
 sg13g2_fill_2 FILLER_49_159 ();
 sg13g2_decap_4 FILLER_49_211 ();
 sg13g2_fill_2 FILLER_49_215 ();
 sg13g2_decap_8 FILLER_49_269 ();
 sg13g2_decap_4 FILLER_49_276 ();
 sg13g2_decap_4 FILLER_49_285 ();
 sg13g2_fill_2 FILLER_49_294 ();
 sg13g2_fill_2 FILLER_49_301 ();
 sg13g2_fill_2 FILLER_49_308 ();
 sg13g2_fill_1 FILLER_49_315 ();
 sg13g2_fill_1 FILLER_49_396 ();
 sg13g2_fill_2 FILLER_49_410 ();
 sg13g2_fill_1 FILLER_49_418 ();
 sg13g2_fill_2 FILLER_49_450 ();
 sg13g2_fill_2 FILLER_49_480 ();
 sg13g2_fill_1 FILLER_49_489 ();
 sg13g2_fill_1 FILLER_49_501 ();
 sg13g2_decap_8 FILLER_49_528 ();
 sg13g2_decap_8 FILLER_49_535 ();
 sg13g2_decap_8 FILLER_49_542 ();
 sg13g2_fill_2 FILLER_49_596 ();
 sg13g2_fill_1 FILLER_49_598 ();
 sg13g2_fill_2 FILLER_49_604 ();
 sg13g2_fill_1 FILLER_49_639 ();
 sg13g2_fill_1 FILLER_49_645 ();
 sg13g2_fill_2 FILLER_49_656 ();
 sg13g2_fill_2 FILLER_49_678 ();
 sg13g2_fill_1 FILLER_49_688 ();
 sg13g2_fill_2 FILLER_49_697 ();
 sg13g2_decap_8 FILLER_49_728 ();
 sg13g2_decap_4 FILLER_49_735 ();
 sg13g2_fill_2 FILLER_49_799 ();
 sg13g2_fill_2 FILLER_49_875 ();
 sg13g2_fill_1 FILLER_49_912 ();
 sg13g2_fill_2 FILLER_49_933 ();
 sg13g2_fill_1 FILLER_49_939 ();
 sg13g2_fill_1 FILLER_49_974 ();
 sg13g2_fill_2 FILLER_49_1003 ();
 sg13g2_fill_2 FILLER_49_1019 ();
 sg13g2_fill_1 FILLER_49_1053 ();
 sg13g2_fill_2 FILLER_49_1069 ();
 sg13g2_fill_1 FILLER_49_1110 ();
 sg13g2_fill_1 FILLER_49_1118 ();
 sg13g2_fill_1 FILLER_49_1133 ();
 sg13g2_fill_2 FILLER_49_1142 ();
 sg13g2_fill_2 FILLER_49_1154 ();
 sg13g2_fill_2 FILLER_49_1172 ();
 sg13g2_fill_1 FILLER_49_1181 ();
 sg13g2_fill_2 FILLER_49_1221 ();
 sg13g2_fill_1 FILLER_49_1223 ();
 sg13g2_fill_2 FILLER_49_1234 ();
 sg13g2_fill_2 FILLER_49_1245 ();
 sg13g2_fill_2 FILLER_49_1264 ();
 sg13g2_fill_2 FILLER_49_1272 ();
 sg13g2_fill_1 FILLER_49_1274 ();
 sg13g2_fill_1 FILLER_49_1307 ();
 sg13g2_decap_8 FILLER_49_1328 ();
 sg13g2_fill_2 FILLER_49_1335 ();
 sg13g2_decap_4 FILLER_49_1352 ();
 sg13g2_decap_4 FILLER_49_1384 ();
 sg13g2_fill_1 FILLER_49_1388 ();
 sg13g2_fill_2 FILLER_49_1402 ();
 sg13g2_fill_1 FILLER_49_1404 ();
 sg13g2_fill_1 FILLER_49_1420 ();
 sg13g2_fill_1 FILLER_49_1443 ();
 sg13g2_fill_1 FILLER_49_1452 ();
 sg13g2_fill_2 FILLER_49_1461 ();
 sg13g2_fill_1 FILLER_49_1491 ();
 sg13g2_fill_2 FILLER_49_1495 ();
 sg13g2_fill_2 FILLER_49_1507 ();
 sg13g2_fill_2 FILLER_49_1527 ();
 sg13g2_fill_2 FILLER_49_1542 ();
 sg13g2_fill_1 FILLER_49_1549 ();
 sg13g2_fill_1 FILLER_49_1584 ();
 sg13g2_fill_1 FILLER_49_1595 ();
 sg13g2_fill_2 FILLER_49_1599 ();
 sg13g2_fill_1 FILLER_49_1601 ();
 sg13g2_fill_1 FILLER_49_1607 ();
 sg13g2_fill_1 FILLER_49_1623 ();
 sg13g2_fill_2 FILLER_49_1630 ();
 sg13g2_fill_1 FILLER_49_1636 ();
 sg13g2_fill_1 FILLER_49_1657 ();
 sg13g2_fill_1 FILLER_49_1665 ();
 sg13g2_fill_1 FILLER_49_1705 ();
 sg13g2_fill_2 FILLER_49_1710 ();
 sg13g2_fill_1 FILLER_49_1712 ();
 sg13g2_fill_2 FILLER_49_1717 ();
 sg13g2_fill_1 FILLER_49_1719 ();
 sg13g2_fill_1 FILLER_49_1733 ();
 sg13g2_fill_1 FILLER_49_1742 ();
 sg13g2_decap_4 FILLER_49_1768 ();
 sg13g2_fill_2 FILLER_49_1772 ();
 sg13g2_decap_4 FILLER_49_1778 ();
 sg13g2_fill_1 FILLER_49_1782 ();
 sg13g2_decap_4 FILLER_49_1800 ();
 sg13g2_fill_2 FILLER_49_1826 ();
 sg13g2_fill_1 FILLER_49_1838 ();
 sg13g2_fill_1 FILLER_49_1860 ();
 sg13g2_fill_2 FILLER_49_1875 ();
 sg13g2_fill_1 FILLER_49_1877 ();
 sg13g2_fill_1 FILLER_49_1899 ();
 sg13g2_fill_1 FILLER_49_1922 ();
 sg13g2_decap_4 FILLER_49_1927 ();
 sg13g2_fill_1 FILLER_49_1936 ();
 sg13g2_decap_4 FILLER_49_1950 ();
 sg13g2_fill_2 FILLER_49_1954 ();
 sg13g2_fill_2 FILLER_49_2010 ();
 sg13g2_fill_1 FILLER_49_2012 ();
 sg13g2_fill_2 FILLER_49_2027 ();
 sg13g2_decap_4 FILLER_49_2097 ();
 sg13g2_fill_2 FILLER_49_2126 ();
 sg13g2_fill_1 FILLER_49_2128 ();
 sg13g2_fill_2 FILLER_49_2134 ();
 sg13g2_fill_1 FILLER_49_2136 ();
 sg13g2_fill_2 FILLER_49_2142 ();
 sg13g2_fill_1 FILLER_49_2154 ();
 sg13g2_decap_8 FILLER_49_2181 ();
 sg13g2_fill_2 FILLER_49_2188 ();
 sg13g2_fill_1 FILLER_49_2203 ();
 sg13g2_fill_1 FILLER_49_2214 ();
 sg13g2_fill_1 FILLER_49_2254 ();
 sg13g2_decap_4 FILLER_49_2341 ();
 sg13g2_fill_1 FILLER_49_2345 ();
 sg13g2_fill_1 FILLER_49_2350 ();
 sg13g2_fill_2 FILLER_49_2365 ();
 sg13g2_fill_2 FILLER_49_2371 ();
 sg13g2_fill_1 FILLER_49_2373 ();
 sg13g2_decap_8 FILLER_49_2388 ();
 sg13g2_fill_1 FILLER_49_2395 ();
 sg13g2_decap_8 FILLER_49_2407 ();
 sg13g2_fill_2 FILLER_49_2414 ();
 sg13g2_fill_1 FILLER_49_2416 ();
 sg13g2_fill_2 FILLER_49_2462 ();
 sg13g2_decap_4 FILLER_49_2474 ();
 sg13g2_decap_4 FILLER_49_2482 ();
 sg13g2_fill_2 FILLER_49_2486 ();
 sg13g2_fill_1 FILLER_49_2494 ();
 sg13g2_decap_4 FILLER_49_2499 ();
 sg13g2_fill_1 FILLER_49_2503 ();
 sg13g2_fill_1 FILLER_49_2509 ();
 sg13g2_fill_1 FILLER_49_2518 ();
 sg13g2_fill_1 FILLER_49_2524 ();
 sg13g2_fill_2 FILLER_49_2529 ();
 sg13g2_fill_1 FILLER_49_2531 ();
 sg13g2_fill_1 FILLER_49_2535 ();
 sg13g2_decap_8 FILLER_49_2572 ();
 sg13g2_decap_4 FILLER_49_2579 ();
 sg13g2_fill_1 FILLER_49_2596 ();
 sg13g2_fill_1 FILLER_49_2600 ();
 sg13g2_fill_1 FILLER_49_2614 ();
 sg13g2_decap_4 FILLER_49_2666 ();
 sg13g2_decap_8 FILLER_50_0 ();
 sg13g2_decap_8 FILLER_50_7 ();
 sg13g2_decap_8 FILLER_50_14 ();
 sg13g2_fill_2 FILLER_50_21 ();
 sg13g2_fill_1 FILLER_50_23 ();
 sg13g2_fill_2 FILLER_50_50 ();
 sg13g2_decap_8 FILLER_50_112 ();
 sg13g2_fill_2 FILLER_50_119 ();
 sg13g2_fill_1 FILLER_50_121 ();
 sg13g2_fill_1 FILLER_50_148 ();
 sg13g2_fill_2 FILLER_50_153 ();
 sg13g2_fill_1 FILLER_50_164 ();
 sg13g2_fill_2 FILLER_50_172 ();
 sg13g2_decap_8 FILLER_50_199 ();
 sg13g2_fill_2 FILLER_50_206 ();
 sg13g2_fill_1 FILLER_50_221 ();
 sg13g2_fill_2 FILLER_50_265 ();
 sg13g2_fill_2 FILLER_50_275 ();
 sg13g2_fill_1 FILLER_50_287 ();
 sg13g2_fill_1 FILLER_50_293 ();
 sg13g2_fill_2 FILLER_50_299 ();
 sg13g2_fill_2 FILLER_50_305 ();
 sg13g2_fill_2 FILLER_50_311 ();
 sg13g2_fill_1 FILLER_50_321 ();
 sg13g2_fill_2 FILLER_50_402 ();
 sg13g2_fill_1 FILLER_50_433 ();
 sg13g2_decap_4 FILLER_50_482 ();
 sg13g2_fill_1 FILLER_50_486 ();
 sg13g2_fill_1 FILLER_50_511 ();
 sg13g2_decap_8 FILLER_50_527 ();
 sg13g2_fill_2 FILLER_50_534 ();
 sg13g2_fill_1 FILLER_50_536 ();
 sg13g2_fill_2 FILLER_50_547 ();
 sg13g2_fill_1 FILLER_50_549 ();
 sg13g2_fill_1 FILLER_50_576 ();
 sg13g2_fill_1 FILLER_50_582 ();
 sg13g2_fill_2 FILLER_50_605 ();
 sg13g2_fill_1 FILLER_50_607 ();
 sg13g2_fill_1 FILLER_50_634 ();
 sg13g2_fill_1 FILLER_50_645 ();
 sg13g2_fill_1 FILLER_50_673 ();
 sg13g2_decap_8 FILLER_50_678 ();
 sg13g2_decap_8 FILLER_50_685 ();
 sg13g2_decap_4 FILLER_50_692 ();
 sg13g2_decap_4 FILLER_50_740 ();
 sg13g2_fill_1 FILLER_50_744 ();
 sg13g2_fill_2 FILLER_50_781 ();
 sg13g2_fill_1 FILLER_50_801 ();
 sg13g2_fill_1 FILLER_50_809 ();
 sg13g2_fill_2 FILLER_50_839 ();
 sg13g2_fill_1 FILLER_50_912 ();
 sg13g2_fill_1 FILLER_50_926 ();
 sg13g2_fill_1 FILLER_50_945 ();
 sg13g2_fill_1 FILLER_50_956 ();
 sg13g2_fill_1 FILLER_50_983 ();
 sg13g2_fill_1 FILLER_50_997 ();
 sg13g2_fill_1 FILLER_50_1006 ();
 sg13g2_fill_1 FILLER_50_1020 ();
 sg13g2_fill_1 FILLER_50_1032 ();
 sg13g2_fill_2 FILLER_50_1046 ();
 sg13g2_fill_2 FILLER_50_1081 ();
 sg13g2_fill_1 FILLER_50_1091 ();
 sg13g2_decap_8 FILLER_50_1215 ();
 sg13g2_decap_8 FILLER_50_1222 ();
 sg13g2_decap_8 FILLER_50_1229 ();
 sg13g2_decap_8 FILLER_50_1236 ();
 sg13g2_fill_2 FILLER_50_1243 ();
 sg13g2_decap_8 FILLER_50_1250 ();
 sg13g2_decap_4 FILLER_50_1257 ();
 sg13g2_fill_2 FILLER_50_1261 ();
 sg13g2_fill_2 FILLER_50_1288 ();
 sg13g2_fill_1 FILLER_50_1328 ();
 sg13g2_fill_1 FILLER_50_1355 ();
 sg13g2_fill_1 FILLER_50_1375 ();
 sg13g2_decap_4 FILLER_50_1382 ();
 sg13g2_fill_1 FILLER_50_1396 ();
 sg13g2_decap_8 FILLER_50_1401 ();
 sg13g2_decap_4 FILLER_50_1411 ();
 sg13g2_fill_1 FILLER_50_1415 ();
 sg13g2_fill_2 FILLER_50_1430 ();
 sg13g2_fill_2 FILLER_50_1450 ();
 sg13g2_fill_1 FILLER_50_1544 ();
 sg13g2_fill_2 FILLER_50_1581 ();
 sg13g2_fill_1 FILLER_50_1583 ();
 sg13g2_fill_2 FILLER_50_1589 ();
 sg13g2_fill_1 FILLER_50_1595 ();
 sg13g2_fill_2 FILLER_50_1606 ();
 sg13g2_fill_1 FILLER_50_1670 ();
 sg13g2_fill_1 FILLER_50_1691 ();
 sg13g2_decap_8 FILLER_50_1705 ();
 sg13g2_fill_1 FILLER_50_1712 ();
 sg13g2_fill_1 FILLER_50_1718 ();
 sg13g2_fill_2 FILLER_50_1723 ();
 sg13g2_fill_1 FILLER_50_1774 ();
 sg13g2_fill_2 FILLER_50_1780 ();
 sg13g2_fill_1 FILLER_50_1782 ();
 sg13g2_decap_8 FILLER_50_1812 ();
 sg13g2_decap_4 FILLER_50_1833 ();
 sg13g2_decap_4 FILLER_50_1847 ();
 sg13g2_fill_1 FILLER_50_1851 ();
 sg13g2_fill_2 FILLER_50_1857 ();
 sg13g2_fill_1 FILLER_50_1859 ();
 sg13g2_fill_2 FILLER_50_1872 ();
 sg13g2_fill_1 FILLER_50_1874 ();
 sg13g2_decap_4 FILLER_50_1889 ();
 sg13g2_fill_1 FILLER_50_1893 ();
 sg13g2_decap_4 FILLER_50_1899 ();
 sg13g2_fill_1 FILLER_50_1903 ();
 sg13g2_fill_1 FILLER_50_1934 ();
 sg13g2_fill_2 FILLER_50_1943 ();
 sg13g2_decap_8 FILLER_50_1958 ();
 sg13g2_fill_1 FILLER_50_1979 ();
 sg13g2_fill_1 FILLER_50_2002 ();
 sg13g2_fill_1 FILLER_50_2013 ();
 sg13g2_fill_1 FILLER_50_2022 ();
 sg13g2_fill_1 FILLER_50_2051 ();
 sg13g2_decap_8 FILLER_50_2087 ();
 sg13g2_fill_2 FILLER_50_2094 ();
 sg13g2_fill_1 FILLER_50_2096 ();
 sg13g2_decap_4 FILLER_50_2133 ();
 sg13g2_fill_2 FILLER_50_2137 ();
 sg13g2_decap_4 FILLER_50_2160 ();
 sg13g2_decap_4 FILLER_50_2178 ();
 sg13g2_fill_1 FILLER_50_2182 ();
 sg13g2_decap_4 FILLER_50_2219 ();
 sg13g2_fill_1 FILLER_50_2223 ();
 sg13g2_fill_2 FILLER_50_2228 ();
 sg13g2_fill_1 FILLER_50_2230 ();
 sg13g2_fill_2 FILLER_50_2252 ();
 sg13g2_fill_2 FILLER_50_2287 ();
 sg13g2_fill_2 FILLER_50_2344 ();
 sg13g2_decap_4 FILLER_50_2376 ();
 sg13g2_fill_2 FILLER_50_2380 ();
 sg13g2_decap_4 FILLER_50_2417 ();
 sg13g2_fill_2 FILLER_50_2421 ();
 sg13g2_fill_2 FILLER_50_2484 ();
 sg13g2_decap_8 FILLER_50_2490 ();
 sg13g2_fill_2 FILLER_50_2497 ();
 sg13g2_decap_4 FILLER_50_2503 ();
 sg13g2_fill_2 FILLER_50_2512 ();
 sg13g2_fill_2 FILLER_50_2540 ();
 sg13g2_fill_1 FILLER_50_2542 ();
 sg13g2_fill_1 FILLER_50_2553 ();
 sg13g2_fill_2 FILLER_50_2580 ();
 sg13g2_fill_1 FILLER_50_2582 ();
 sg13g2_fill_1 FILLER_50_2609 ();
 sg13g2_fill_2 FILLER_50_2620 ();
 sg13g2_fill_1 FILLER_50_2651 ();
 sg13g2_decap_8 FILLER_50_2659 ();
 sg13g2_decap_4 FILLER_50_2666 ();
 sg13g2_decap_8 FILLER_51_0 ();
 sg13g2_decap_8 FILLER_51_7 ();
 sg13g2_decap_8 FILLER_51_14 ();
 sg13g2_decap_8 FILLER_51_21 ();
 sg13g2_fill_2 FILLER_51_28 ();
 sg13g2_fill_1 FILLER_51_30 ();
 sg13g2_decap_4 FILLER_51_35 ();
 sg13g2_fill_2 FILLER_51_65 ();
 sg13g2_decap_4 FILLER_51_101 ();
 sg13g2_fill_1 FILLER_51_105 ();
 sg13g2_decap_8 FILLER_51_116 ();
 sg13g2_decap_4 FILLER_51_123 ();
 sg13g2_fill_1 FILLER_51_127 ();
 sg13g2_fill_2 FILLER_51_132 ();
 sg13g2_fill_1 FILLER_51_137 ();
 sg13g2_fill_2 FILLER_51_142 ();
 sg13g2_fill_1 FILLER_51_144 ();
 sg13g2_fill_2 FILLER_51_183 ();
 sg13g2_decap_8 FILLER_51_216 ();
 sg13g2_decap_8 FILLER_51_223 ();
 sg13g2_decap_8 FILLER_51_230 ();
 sg13g2_fill_1 FILLER_51_237 ();
 sg13g2_fill_2 FILLER_51_242 ();
 sg13g2_decap_4 FILLER_51_253 ();
 sg13g2_fill_1 FILLER_51_257 ();
 sg13g2_fill_1 FILLER_51_263 ();
 sg13g2_fill_1 FILLER_51_305 ();
 sg13g2_fill_1 FILLER_51_353 ();
 sg13g2_fill_2 FILLER_51_359 ();
 sg13g2_fill_1 FILLER_51_366 ();
 sg13g2_fill_1 FILLER_51_380 ();
 sg13g2_fill_1 FILLER_51_418 ();
 sg13g2_fill_2 FILLER_51_428 ();
 sg13g2_fill_2 FILLER_51_441 ();
 sg13g2_decap_4 FILLER_51_447 ();
 sg13g2_fill_2 FILLER_51_455 ();
 sg13g2_fill_2 FILLER_51_465 ();
 sg13g2_fill_1 FILLER_51_467 ();
 sg13g2_fill_1 FILLER_51_478 ();
 sg13g2_decap_4 FILLER_51_482 ();
 sg13g2_fill_1 FILLER_51_486 ();
 sg13g2_decap_4 FILLER_51_497 ();
 sg13g2_fill_1 FILLER_51_501 ();
 sg13g2_fill_2 FILLER_51_507 ();
 sg13g2_fill_2 FILLER_51_513 ();
 sg13g2_fill_2 FILLER_51_546 ();
 sg13g2_fill_2 FILLER_51_563 ();
 sg13g2_fill_2 FILLER_51_626 ();
 sg13g2_fill_2 FILLER_51_641 ();
 sg13g2_fill_2 FILLER_51_656 ();
 sg13g2_decap_8 FILLER_51_668 ();
 sg13g2_fill_1 FILLER_51_746 ();
 sg13g2_fill_1 FILLER_51_752 ();
 sg13g2_fill_1 FILLER_51_779 ();
 sg13g2_fill_2 FILLER_51_825 ();
 sg13g2_fill_1 FILLER_51_831 ();
 sg13g2_fill_2 FILLER_51_843 ();
 sg13g2_fill_1 FILLER_51_852 ();
 sg13g2_fill_2 FILLER_51_893 ();
 sg13g2_fill_2 FILLER_51_924 ();
 sg13g2_fill_2 FILLER_51_989 ();
 sg13g2_fill_2 FILLER_51_1014 ();
 sg13g2_fill_2 FILLER_51_1029 ();
 sg13g2_fill_2 FILLER_51_1057 ();
 sg13g2_fill_1 FILLER_51_1073 ();
 sg13g2_fill_2 FILLER_51_1121 ();
 sg13g2_fill_2 FILLER_51_1133 ();
 sg13g2_fill_2 FILLER_51_1161 ();
 sg13g2_fill_1 FILLER_51_1193 ();
 sg13g2_fill_2 FILLER_51_1198 ();
 sg13g2_fill_1 FILLER_51_1204 ();
 sg13g2_fill_2 FILLER_51_1211 ();
 sg13g2_fill_1 FILLER_51_1216 ();
 sg13g2_decap_4 FILLER_51_1227 ();
 sg13g2_decap_8 FILLER_51_1236 ();
 sg13g2_fill_2 FILLER_51_1243 ();
 sg13g2_fill_1 FILLER_51_1320 ();
 sg13g2_decap_4 FILLER_51_1327 ();
 sg13g2_fill_1 FILLER_51_1331 ();
 sg13g2_decap_4 FILLER_51_1336 ();
 sg13g2_fill_1 FILLER_51_1344 ();
 sg13g2_fill_2 FILLER_51_1360 ();
 sg13g2_fill_2 FILLER_51_1387 ();
 sg13g2_fill_1 FILLER_51_1389 ();
 sg13g2_decap_4 FILLER_51_1403 ();
 sg13g2_fill_2 FILLER_51_1407 ();
 sg13g2_decap_4 FILLER_51_1413 ();
 sg13g2_fill_1 FILLER_51_1423 ();
 sg13g2_fill_2 FILLER_51_1433 ();
 sg13g2_fill_1 FILLER_51_1495 ();
 sg13g2_fill_1 FILLER_51_1507 ();
 sg13g2_fill_2 FILLER_51_1522 ();
 sg13g2_fill_2 FILLER_51_1565 ();
 sg13g2_fill_1 FILLER_51_1571 ();
 sg13g2_fill_1 FILLER_51_1580 ();
 sg13g2_fill_2 FILLER_51_1586 ();
 sg13g2_fill_1 FILLER_51_1588 ();
 sg13g2_fill_2 FILLER_51_1599 ();
 sg13g2_fill_1 FILLER_51_1605 ();
 sg13g2_decap_8 FILLER_51_1612 ();
 sg13g2_fill_2 FILLER_51_1619 ();
 sg13g2_fill_1 FILLER_51_1621 ();
 sg13g2_fill_1 FILLER_51_1627 ();
 sg13g2_decap_8 FILLER_51_1632 ();
 sg13g2_fill_1 FILLER_51_1667 ();
 sg13g2_decap_4 FILLER_51_1703 ();
 sg13g2_fill_2 FILLER_51_1711 ();
 sg13g2_fill_1 FILLER_51_1713 ();
 sg13g2_decap_4 FILLER_51_1719 ();
 sg13g2_fill_1 FILLER_51_1723 ();
 sg13g2_fill_2 FILLER_51_1728 ();
 sg13g2_fill_1 FILLER_51_1730 ();
 sg13g2_decap_8 FILLER_51_1751 ();
 sg13g2_fill_2 FILLER_51_1758 ();
 sg13g2_fill_1 FILLER_51_1760 ();
 sg13g2_fill_2 FILLER_51_1769 ();
 sg13g2_fill_2 FILLER_51_1791 ();
 sg13g2_decap_8 FILLER_51_1802 ();
 sg13g2_fill_2 FILLER_51_1809 ();
 sg13g2_fill_1 FILLER_51_1811 ();
 sg13g2_decap_4 FILLER_51_1852 ();
 sg13g2_decap_8 FILLER_51_1861 ();
 sg13g2_decap_8 FILLER_51_1868 ();
 sg13g2_decap_8 FILLER_51_1875 ();
 sg13g2_fill_2 FILLER_51_1882 ();
 sg13g2_fill_1 FILLER_51_1884 ();
 sg13g2_fill_2 FILLER_51_1894 ();
 sg13g2_fill_2 FILLER_51_1911 ();
 sg13g2_fill_1 FILLER_51_1913 ();
 sg13g2_fill_1 FILLER_51_1922 ();
 sg13g2_decap_4 FILLER_51_1928 ();
 sg13g2_fill_1 FILLER_51_1932 ();
 sg13g2_decap_8 FILLER_51_1938 ();
 sg13g2_fill_2 FILLER_51_1945 ();
 sg13g2_fill_1 FILLER_51_1947 ();
 sg13g2_decap_8 FILLER_51_1953 ();
 sg13g2_decap_8 FILLER_51_1960 ();
 sg13g2_fill_2 FILLER_51_1967 ();
 sg13g2_fill_1 FILLER_51_2002 ();
 sg13g2_decap_4 FILLER_51_2007 ();
 sg13g2_fill_2 FILLER_51_2015 ();
 sg13g2_fill_1 FILLER_51_2023 ();
 sg13g2_fill_1 FILLER_51_2030 ();
 sg13g2_fill_2 FILLER_51_2074 ();
 sg13g2_decap_8 FILLER_51_2080 ();
 sg13g2_decap_8 FILLER_51_2087 ();
 sg13g2_decap_4 FILLER_51_2094 ();
 sg13g2_fill_1 FILLER_51_2098 ();
 sg13g2_fill_2 FILLER_51_2104 ();
 sg13g2_decap_4 FILLER_51_2110 ();
 sg13g2_fill_1 FILLER_51_2114 ();
 sg13g2_fill_1 FILLER_51_2123 ();
 sg13g2_fill_2 FILLER_51_2164 ();
 sg13g2_fill_1 FILLER_51_2239 ();
 sg13g2_decap_8 FILLER_51_2277 ();
 sg13g2_decap_8 FILLER_51_2284 ();
 sg13g2_decap_4 FILLER_51_2291 ();
 sg13g2_fill_1 FILLER_51_2295 ();
 sg13g2_fill_1 FILLER_51_2308 ();
 sg13g2_fill_1 FILLER_51_2345 ();
 sg13g2_decap_4 FILLER_51_2353 ();
 sg13g2_fill_1 FILLER_51_2357 ();
 sg13g2_decap_4 FILLER_51_2362 ();
 sg13g2_decap_4 FILLER_51_2386 ();
 sg13g2_decap_8 FILLER_51_2394 ();
 sg13g2_fill_1 FILLER_51_2401 ();
 sg13g2_decap_4 FILLER_51_2411 ();
 sg13g2_fill_2 FILLER_51_2415 ();
 sg13g2_fill_2 FILLER_51_2427 ();
 sg13g2_fill_2 FILLER_51_2439 ();
 sg13g2_fill_2 FILLER_51_2447 ();
 sg13g2_decap_4 FILLER_51_2457 ();
 sg13g2_fill_2 FILLER_51_2461 ();
 sg13g2_fill_2 FILLER_51_2467 ();
 sg13g2_decap_8 FILLER_51_2473 ();
 sg13g2_fill_2 FILLER_51_2480 ();
 sg13g2_decap_8 FILLER_51_2550 ();
 sg13g2_decap_4 FILLER_51_2557 ();
 sg13g2_fill_2 FILLER_51_2605 ();
 sg13g2_fill_1 FILLER_51_2669 ();
 sg13g2_fill_2 FILLER_52_0 ();
 sg13g2_decap_8 FILLER_52_33 ();
 sg13g2_fill_1 FILLER_52_40 ();
 sg13g2_fill_1 FILLER_52_81 ();
 sg13g2_decap_8 FILLER_52_86 ();
 sg13g2_fill_2 FILLER_52_133 ();
 sg13g2_fill_1 FILLER_52_135 ();
 sg13g2_decap_8 FILLER_52_140 ();
 sg13g2_decap_8 FILLER_52_147 ();
 sg13g2_decap_8 FILLER_52_171 ();
 sg13g2_fill_2 FILLER_52_201 ();
 sg13g2_fill_1 FILLER_52_203 ();
 sg13g2_decap_4 FILLER_52_234 ();
 sg13g2_fill_2 FILLER_52_238 ();
 sg13g2_fill_2 FILLER_52_245 ();
 sg13g2_fill_1 FILLER_52_247 ();
 sg13g2_fill_2 FILLER_52_283 ();
 sg13g2_fill_1 FILLER_52_289 ();
 sg13g2_fill_2 FILLER_52_311 ();
 sg13g2_fill_1 FILLER_52_322 ();
 sg13g2_fill_1 FILLER_52_333 ();
 sg13g2_fill_2 FILLER_52_346 ();
 sg13g2_fill_1 FILLER_52_388 ();
 sg13g2_fill_1 FILLER_52_405 ();
 sg13g2_decap_4 FILLER_52_440 ();
 sg13g2_fill_2 FILLER_52_447 ();
 sg13g2_fill_1 FILLER_52_449 ();
 sg13g2_fill_2 FILLER_52_464 ();
 sg13g2_fill_2 FILLER_52_505 ();
 sg13g2_decap_8 FILLER_52_517 ();
 sg13g2_fill_1 FILLER_52_524 ();
 sg13g2_fill_1 FILLER_52_593 ();
 sg13g2_fill_2 FILLER_52_612 ();
 sg13g2_fill_2 FILLER_52_645 ();
 sg13g2_fill_1 FILLER_52_664 ();
 sg13g2_decap_8 FILLER_52_670 ();
 sg13g2_decap_8 FILLER_52_677 ();
 sg13g2_decap_4 FILLER_52_684 ();
 sg13g2_fill_1 FILLER_52_688 ();
 sg13g2_fill_2 FILLER_52_742 ();
 sg13g2_fill_1 FILLER_52_744 ();
 sg13g2_fill_1 FILLER_52_749 ();
 sg13g2_fill_2 FILLER_52_764 ();
 sg13g2_fill_1 FILLER_52_785 ();
 sg13g2_fill_1 FILLER_52_791 ();
 sg13g2_fill_2 FILLER_52_839 ();
 sg13g2_fill_1 FILLER_52_911 ();
 sg13g2_fill_1 FILLER_52_929 ();
 sg13g2_fill_2 FILLER_52_959 ();
 sg13g2_fill_2 FILLER_52_1024 ();
 sg13g2_fill_2 FILLER_52_1037 ();
 sg13g2_fill_1 FILLER_52_1091 ();
 sg13g2_fill_1 FILLER_52_1134 ();
 sg13g2_fill_2 FILLER_52_1173 ();
 sg13g2_fill_1 FILLER_52_1179 ();
 sg13g2_fill_1 FILLER_52_1184 ();
 sg13g2_fill_2 FILLER_52_1194 ();
 sg13g2_fill_1 FILLER_52_1196 ();
 sg13g2_fill_2 FILLER_52_1202 ();
 sg13g2_fill_1 FILLER_52_1204 ();
 sg13g2_fill_2 FILLER_52_1215 ();
 sg13g2_fill_1 FILLER_52_1225 ();
 sg13g2_decap_8 FILLER_52_1247 ();
 sg13g2_fill_1 FILLER_52_1254 ();
 sg13g2_fill_2 FILLER_52_1261 ();
 sg13g2_fill_1 FILLER_52_1263 ();
 sg13g2_fill_2 FILLER_52_1269 ();
 sg13g2_fill_1 FILLER_52_1271 ();
 sg13g2_fill_2 FILLER_52_1276 ();
 sg13g2_decap_4 FILLER_52_1323 ();
 sg13g2_fill_2 FILLER_52_1327 ();
 sg13g2_decap_4 FILLER_52_1339 ();
 sg13g2_fill_1 FILLER_52_1343 ();
 sg13g2_fill_2 FILLER_52_1355 ();
 sg13g2_fill_1 FILLER_52_1357 ();
 sg13g2_decap_8 FILLER_52_1376 ();
 sg13g2_decap_8 FILLER_52_1383 ();
 sg13g2_decap_8 FILLER_52_1390 ();
 sg13g2_decap_4 FILLER_52_1397 ();
 sg13g2_fill_1 FILLER_52_1423 ();
 sg13g2_fill_2 FILLER_52_1443 ();
 sg13g2_fill_1 FILLER_52_1453 ();
 sg13g2_fill_1 FILLER_52_1459 ();
 sg13g2_fill_1 FILLER_52_1472 ();
 sg13g2_fill_1 FILLER_52_1498 ();
 sg13g2_fill_1 FILLER_52_1558 ();
 sg13g2_decap_8 FILLER_52_1575 ();
 sg13g2_decap_4 FILLER_52_1582 ();
 sg13g2_fill_2 FILLER_52_1586 ();
 sg13g2_decap_8 FILLER_52_1599 ();
 sg13g2_decap_4 FILLER_52_1606 ();
 sg13g2_fill_1 FILLER_52_1610 ();
 sg13g2_decap_8 FILLER_52_1616 ();
 sg13g2_decap_8 FILLER_52_1623 ();
 sg13g2_fill_2 FILLER_52_1640 ();
 sg13g2_fill_1 FILLER_52_1642 ();
 sg13g2_fill_1 FILLER_52_1704 ();
 sg13g2_fill_1 FILLER_52_1709 ();
 sg13g2_decap_4 FILLER_52_1720 ();
 sg13g2_fill_2 FILLER_52_1724 ();
 sg13g2_fill_1 FILLER_52_1762 ();
 sg13g2_fill_1 FILLER_52_1768 ();
 sg13g2_fill_1 FILLER_52_1775 ();
 sg13g2_fill_1 FILLER_52_1806 ();
 sg13g2_fill_2 FILLER_52_1812 ();
 sg13g2_fill_1 FILLER_52_1814 ();
 sg13g2_fill_2 FILLER_52_1831 ();
 sg13g2_fill_1 FILLER_52_1833 ();
 sg13g2_fill_1 FILLER_52_1853 ();
 sg13g2_fill_2 FILLER_52_1863 ();
 sg13g2_fill_1 FILLER_52_1865 ();
 sg13g2_fill_2 FILLER_52_1897 ();
 sg13g2_decap_8 FILLER_52_1920 ();
 sg13g2_fill_2 FILLER_52_1927 ();
 sg13g2_decap_8 FILLER_52_1934 ();
 sg13g2_decap_8 FILLER_52_1941 ();
 sg13g2_decap_8 FILLER_52_1948 ();
 sg13g2_decap_4 FILLER_52_1955 ();
 sg13g2_fill_2 FILLER_52_1959 ();
 sg13g2_fill_2 FILLER_52_1965 ();
 sg13g2_fill_2 FILLER_52_2003 ();
 sg13g2_fill_1 FILLER_52_2005 ();
 sg13g2_fill_2 FILLER_52_2072 ();
 sg13g2_decap_8 FILLER_52_2080 ();
 sg13g2_decap_4 FILLER_52_2087 ();
 sg13g2_fill_2 FILLER_52_2091 ();
 sg13g2_decap_8 FILLER_52_2103 ();
 sg13g2_decap_8 FILLER_52_2110 ();
 sg13g2_decap_4 FILLER_52_2117 ();
 sg13g2_fill_2 FILLER_52_2121 ();
 sg13g2_fill_1 FILLER_52_2150 ();
 sg13g2_fill_2 FILLER_52_2155 ();
 sg13g2_fill_2 FILLER_52_2203 ();
 sg13g2_fill_1 FILLER_52_2205 ();
 sg13g2_fill_2 FILLER_52_2232 ();
 sg13g2_fill_1 FILLER_52_2234 ();
 sg13g2_decap_8 FILLER_52_2264 ();
 sg13g2_decap_8 FILLER_52_2271 ();
 sg13g2_decap_8 FILLER_52_2278 ();
 sg13g2_fill_1 FILLER_52_2285 ();
 sg13g2_fill_1 FILLER_52_2294 ();
 sg13g2_fill_2 FILLER_52_2307 ();
 sg13g2_fill_1 FILLER_52_2320 ();
 sg13g2_fill_2 FILLER_52_2355 ();
 sg13g2_fill_1 FILLER_52_2357 ();
 sg13g2_decap_8 FILLER_52_2388 ();
 sg13g2_decap_4 FILLER_52_2395 ();
 sg13g2_fill_2 FILLER_52_2404 ();
 sg13g2_decap_8 FILLER_52_2471 ();
 sg13g2_decap_4 FILLER_52_2478 ();
 sg13g2_fill_1 FILLER_52_2482 ();
 sg13g2_decap_8 FILLER_52_2542 ();
 sg13g2_decap_8 FILLER_52_2549 ();
 sg13g2_decap_8 FILLER_52_2556 ();
 sg13g2_decap_8 FILLER_52_2563 ();
 sg13g2_decap_8 FILLER_52_2570 ();
 sg13g2_decap_8 FILLER_52_2577 ();
 sg13g2_fill_2 FILLER_52_2588 ();
 sg13g2_decap_8 FILLER_52_2598 ();
 sg13g2_fill_1 FILLER_52_2605 ();
 sg13g2_decap_8 FILLER_52_2616 ();
 sg13g2_fill_2 FILLER_52_2627 ();
 sg13g2_fill_1 FILLER_52_2629 ();
 sg13g2_decap_8 FILLER_52_2634 ();
 sg13g2_fill_1 FILLER_52_2641 ();
 sg13g2_fill_2 FILLER_52_2668 ();
 sg13g2_fill_2 FILLER_53_0 ();
 sg13g2_decap_4 FILLER_53_44 ();
 sg13g2_decap_8 FILLER_53_65 ();
 sg13g2_decap_8 FILLER_53_72 ();
 sg13g2_decap_8 FILLER_53_79 ();
 sg13g2_decap_8 FILLER_53_86 ();
 sg13g2_fill_2 FILLER_53_93 ();
 sg13g2_fill_1 FILLER_53_95 ();
 sg13g2_decap_8 FILLER_53_100 ();
 sg13g2_fill_1 FILLER_53_111 ();
 sg13g2_fill_2 FILLER_53_178 ();
 sg13g2_fill_1 FILLER_53_180 ();
 sg13g2_fill_1 FILLER_53_193 ();
 sg13g2_fill_1 FILLER_53_220 ();
 sg13g2_fill_1 FILLER_53_231 ();
 sg13g2_fill_1 FILLER_53_258 ();
 sg13g2_decap_4 FILLER_53_263 ();
 sg13g2_fill_1 FILLER_53_267 ();
 sg13g2_decap_8 FILLER_53_277 ();
 sg13g2_decap_4 FILLER_53_284 ();
 sg13g2_fill_1 FILLER_53_288 ();
 sg13g2_fill_2 FILLER_53_327 ();
 sg13g2_fill_1 FILLER_53_337 ();
 sg13g2_fill_2 FILLER_53_342 ();
 sg13g2_fill_1 FILLER_53_349 ();
 sg13g2_fill_1 FILLER_53_355 ();
 sg13g2_fill_1 FILLER_53_381 ();
 sg13g2_fill_2 FILLER_53_400 ();
 sg13g2_fill_1 FILLER_53_418 ();
 sg13g2_fill_2 FILLER_53_430 ();
 sg13g2_fill_2 FILLER_53_456 ();
 sg13g2_fill_2 FILLER_53_461 ();
 sg13g2_fill_1 FILLER_53_490 ();
 sg13g2_fill_1 FILLER_53_527 ();
 sg13g2_fill_2 FILLER_53_532 ();
 sg13g2_fill_1 FILLER_53_544 ();
 sg13g2_fill_1 FILLER_53_580 ();
 sg13g2_fill_1 FILLER_53_590 ();
 sg13g2_fill_2 FILLER_53_606 ();
 sg13g2_fill_1 FILLER_53_622 ();
 sg13g2_fill_1 FILLER_53_640 ();
 sg13g2_decap_8 FILLER_53_682 ();
 sg13g2_decap_8 FILLER_53_689 ();
 sg13g2_fill_2 FILLER_53_696 ();
 sg13g2_fill_1 FILLER_53_705 ();
 sg13g2_fill_2 FILLER_53_719 ();
 sg13g2_fill_2 FILLER_53_725 ();
 sg13g2_fill_2 FILLER_53_737 ();
 sg13g2_fill_1 FILLER_53_739 ();
 sg13g2_fill_1 FILLER_53_745 ();
 sg13g2_fill_2 FILLER_53_750 ();
 sg13g2_fill_1 FILLER_53_752 ();
 sg13g2_fill_2 FILLER_53_757 ();
 sg13g2_fill_2 FILLER_53_771 ();
 sg13g2_fill_2 FILLER_53_784 ();
 sg13g2_fill_2 FILLER_53_847 ();
 sg13g2_fill_2 FILLER_53_879 ();
 sg13g2_fill_1 FILLER_53_937 ();
 sg13g2_fill_1 FILLER_53_942 ();
 sg13g2_fill_1 FILLER_53_953 ();
 sg13g2_fill_2 FILLER_53_1011 ();
 sg13g2_fill_1 FILLER_53_1016 ();
 sg13g2_fill_2 FILLER_53_1046 ();
 sg13g2_fill_1 FILLER_53_1146 ();
 sg13g2_fill_2 FILLER_53_1176 ();
 sg13g2_fill_1 FILLER_53_1213 ();
 sg13g2_fill_2 FILLER_53_1235 ();
 sg13g2_fill_2 FILLER_53_1252 ();
 sg13g2_fill_1 FILLER_53_1254 ();
 sg13g2_fill_1 FILLER_53_1262 ();
 sg13g2_fill_1 FILLER_53_1267 ();
 sg13g2_fill_1 FILLER_53_1273 ();
 sg13g2_fill_1 FILLER_53_1291 ();
 sg13g2_fill_2 FILLER_53_1320 ();
 sg13g2_fill_1 FILLER_53_1340 ();
 sg13g2_fill_2 FILLER_53_1371 ();
 sg13g2_decap_8 FILLER_53_1386 ();
 sg13g2_decap_8 FILLER_53_1393 ();
 sg13g2_fill_1 FILLER_53_1435 ();
 sg13g2_fill_1 FILLER_53_1470 ();
 sg13g2_fill_2 FILLER_53_1491 ();
 sg13g2_fill_1 FILLER_53_1569 ();
 sg13g2_fill_1 FILLER_53_1593 ();
 sg13g2_decap_4 FILLER_53_1624 ();
 sg13g2_fill_1 FILLER_53_1628 ();
 sg13g2_fill_2 FILLER_53_1650 ();
 sg13g2_fill_1 FILLER_53_1652 ();
 sg13g2_fill_1 FILLER_53_1669 ();
 sg13g2_fill_1 FILLER_53_1678 ();
 sg13g2_fill_2 FILLER_53_1684 ();
 sg13g2_fill_2 FILLER_53_1691 ();
 sg13g2_decap_8 FILLER_53_1696 ();
 sg13g2_fill_2 FILLER_53_1703 ();
 sg13g2_decap_8 FILLER_53_1710 ();
 sg13g2_fill_2 FILLER_53_1717 ();
 sg13g2_fill_1 FILLER_53_1719 ();
 sg13g2_fill_2 FILLER_53_1725 ();
 sg13g2_decap_8 FILLER_53_1737 ();
 sg13g2_fill_2 FILLER_53_1748 ();
 sg13g2_fill_1 FILLER_53_1754 ();
 sg13g2_fill_1 FILLER_53_1768 ();
 sg13g2_decap_8 FILLER_53_1774 ();
 sg13g2_fill_2 FILLER_53_1786 ();
 sg13g2_decap_4 FILLER_53_1792 ();
 sg13g2_decap_8 FILLER_53_1801 ();
 sg13g2_fill_1 FILLER_53_1848 ();
 sg13g2_fill_2 FILLER_53_1854 ();
 sg13g2_fill_1 FILLER_53_1856 ();
 sg13g2_decap_4 FILLER_53_1865 ();
 sg13g2_fill_1 FILLER_53_1869 ();
 sg13g2_fill_2 FILLER_53_1874 ();
 sg13g2_fill_1 FILLER_53_1882 ();
 sg13g2_decap_8 FILLER_53_1888 ();
 sg13g2_decap_4 FILLER_53_1895 ();
 sg13g2_fill_2 FILLER_53_1906 ();
 sg13g2_fill_1 FILLER_53_1908 ();
 sg13g2_fill_2 FILLER_53_1922 ();
 sg13g2_fill_2 FILLER_53_1934 ();
 sg13g2_fill_1 FILLER_53_1936 ();
 sg13g2_decap_8 FILLER_53_1952 ();
 sg13g2_decap_4 FILLER_53_1959 ();
 sg13g2_fill_1 FILLER_53_1963 ();
 sg13g2_fill_1 FILLER_53_1981 ();
 sg13g2_fill_1 FILLER_53_2024 ();
 sg13g2_fill_1 FILLER_53_2029 ();
 sg13g2_fill_1 FILLER_53_2048 ();
 sg13g2_fill_1 FILLER_53_2067 ();
 sg13g2_decap_4 FILLER_53_2089 ();
 sg13g2_fill_2 FILLER_53_2128 ();
 sg13g2_fill_1 FILLER_53_2130 ();
 sg13g2_decap_8 FILLER_53_2157 ();
 sg13g2_decap_4 FILLER_53_2164 ();
 sg13g2_fill_1 FILLER_53_2168 ();
 sg13g2_decap_8 FILLER_53_2177 ();
 sg13g2_decap_8 FILLER_53_2184 ();
 sg13g2_fill_2 FILLER_53_2191 ();
 sg13g2_fill_2 FILLER_53_2201 ();
 sg13g2_fill_1 FILLER_53_2203 ();
 sg13g2_fill_2 FILLER_53_2227 ();
 sg13g2_fill_1 FILLER_53_2229 ();
 sg13g2_decap_8 FILLER_53_2255 ();
 sg13g2_decap_8 FILLER_53_2262 ();
 sg13g2_decap_8 FILLER_53_2269 ();
 sg13g2_decap_4 FILLER_53_2276 ();
 sg13g2_fill_2 FILLER_53_2280 ();
 sg13g2_fill_2 FILLER_53_2340 ();
 sg13g2_fill_2 FILLER_53_2345 ();
 sg13g2_fill_1 FILLER_53_2347 ();
 sg13g2_fill_2 FILLER_53_2395 ();
 sg13g2_fill_1 FILLER_53_2397 ();
 sg13g2_decap_4 FILLER_53_2409 ();
 sg13g2_fill_1 FILLER_53_2421 ();
 sg13g2_fill_1 FILLER_53_2426 ();
 sg13g2_decap_8 FILLER_53_2431 ();
 sg13g2_decap_8 FILLER_53_2438 ();
 sg13g2_fill_2 FILLER_53_2457 ();
 sg13g2_fill_2 FILLER_53_2485 ();
 sg13g2_decap_4 FILLER_53_2508 ();
 sg13g2_fill_2 FILLER_53_2512 ();
 sg13g2_decap_8 FILLER_53_2530 ();
 sg13g2_decap_4 FILLER_53_2548 ();
 sg13g2_fill_2 FILLER_53_2552 ();
 sg13g2_fill_2 FILLER_53_2606 ();
 sg13g2_decap_8 FILLER_53_2625 ();
 sg13g2_decap_8 FILLER_53_2632 ();
 sg13g2_decap_8 FILLER_53_2639 ();
 sg13g2_fill_1 FILLER_53_2646 ();
 sg13g2_decap_8 FILLER_53_2651 ();
 sg13g2_decap_8 FILLER_53_2658 ();
 sg13g2_decap_4 FILLER_53_2665 ();
 sg13g2_fill_1 FILLER_53_2669 ();
 sg13g2_fill_2 FILLER_54_0 ();
 sg13g2_decap_8 FILLER_54_46 ();
 sg13g2_fill_2 FILLER_54_53 ();
 sg13g2_fill_1 FILLER_54_55 ();
 sg13g2_decap_4 FILLER_54_60 ();
 sg13g2_fill_1 FILLER_54_64 ();
 sg13g2_decap_4 FILLER_54_91 ();
 sg13g2_decap_8 FILLER_54_103 ();
 sg13g2_decap_8 FILLER_54_110 ();
 sg13g2_decap_4 FILLER_54_117 ();
 sg13g2_decap_4 FILLER_54_125 ();
 sg13g2_decap_8 FILLER_54_164 ();
 sg13g2_decap_4 FILLER_54_171 ();
 sg13g2_fill_1 FILLER_54_210 ();
 sg13g2_fill_1 FILLER_54_215 ();
 sg13g2_decap_4 FILLER_54_251 ();
 sg13g2_fill_2 FILLER_54_255 ();
 sg13g2_decap_4 FILLER_54_261 ();
 sg13g2_fill_1 FILLER_54_265 ();
 sg13g2_fill_2 FILLER_54_292 ();
 sg13g2_fill_1 FILLER_54_294 ();
 sg13g2_fill_2 FILLER_54_312 ();
 sg13g2_fill_2 FILLER_54_326 ();
 sg13g2_fill_2 FILLER_54_436 ();
 sg13g2_fill_2 FILLER_54_499 ();
 sg13g2_fill_2 FILLER_54_541 ();
 sg13g2_fill_1 FILLER_54_543 ();
 sg13g2_fill_2 FILLER_54_548 ();
 sg13g2_fill_2 FILLER_54_554 ();
 sg13g2_fill_1 FILLER_54_579 ();
 sg13g2_fill_1 FILLER_54_594 ();
 sg13g2_fill_2 FILLER_54_612 ();
 sg13g2_fill_1 FILLER_54_614 ();
 sg13g2_fill_2 FILLER_54_639 ();
 sg13g2_decap_4 FILLER_54_646 ();
 sg13g2_fill_2 FILLER_54_650 ();
 sg13g2_fill_1 FILLER_54_665 ();
 sg13g2_fill_2 FILLER_54_696 ();
 sg13g2_fill_1 FILLER_54_698 ();
 sg13g2_fill_2 FILLER_54_724 ();
 sg13g2_fill_1 FILLER_54_726 ();
 sg13g2_fill_2 FILLER_54_731 ();
 sg13g2_fill_1 FILLER_54_733 ();
 sg13g2_fill_2 FILLER_54_756 ();
 sg13g2_fill_2 FILLER_54_787 ();
 sg13g2_fill_1 FILLER_54_804 ();
 sg13g2_fill_1 FILLER_54_852 ();
 sg13g2_fill_1 FILLER_54_866 ();
 sg13g2_fill_1 FILLER_54_886 ();
 sg13g2_fill_2 FILLER_54_916 ();
 sg13g2_fill_2 FILLER_54_927 ();
 sg13g2_fill_1 FILLER_54_933 ();
 sg13g2_fill_1 FILLER_54_939 ();
 sg13g2_fill_2 FILLER_54_944 ();
 sg13g2_fill_2 FILLER_54_953 ();
 sg13g2_fill_2 FILLER_54_981 ();
 sg13g2_fill_2 FILLER_54_987 ();
 sg13g2_fill_2 FILLER_54_1044 ();
 sg13g2_fill_1 FILLER_54_1112 ();
 sg13g2_fill_2 FILLER_54_1117 ();
 sg13g2_decap_8 FILLER_54_1149 ();
 sg13g2_decap_4 FILLER_54_1160 ();
 sg13g2_fill_1 FILLER_54_1164 ();
 sg13g2_fill_2 FILLER_54_1178 ();
 sg13g2_decap_8 FILLER_54_1194 ();
 sg13g2_fill_2 FILLER_54_1201 ();
 sg13g2_fill_2 FILLER_54_1211 ();
 sg13g2_fill_2 FILLER_54_1246 ();
 sg13g2_fill_1 FILLER_54_1248 ();
 sg13g2_decap_4 FILLER_54_1255 ();
 sg13g2_fill_2 FILLER_54_1264 ();
 sg13g2_decap_8 FILLER_54_1275 ();
 sg13g2_decap_4 FILLER_54_1282 ();
 sg13g2_fill_2 FILLER_54_1300 ();
 sg13g2_decap_8 FILLER_54_1318 ();
 sg13g2_fill_2 FILLER_54_1325 ();
 sg13g2_decap_8 FILLER_54_1336 ();
 sg13g2_fill_2 FILLER_54_1343 ();
 sg13g2_decap_8 FILLER_54_1350 ();
 sg13g2_decap_8 FILLER_54_1357 ();
 sg13g2_fill_1 FILLER_54_1364 ();
 sg13g2_decap_8 FILLER_54_1369 ();
 sg13g2_decap_8 FILLER_54_1376 ();
 sg13g2_fill_2 FILLER_54_1383 ();
 sg13g2_fill_1 FILLER_54_1385 ();
 sg13g2_fill_1 FILLER_54_1399 ();
 sg13g2_fill_1 FILLER_54_1431 ();
 sg13g2_fill_1 FILLER_54_1445 ();
 sg13g2_fill_1 FILLER_54_1450 ();
 sg13g2_fill_1 FILLER_54_1473 ();
 sg13g2_fill_2 FILLER_54_1512 ();
 sg13g2_fill_1 FILLER_54_1559 ();
 sg13g2_decap_4 FILLER_54_1579 ();
 sg13g2_fill_2 FILLER_54_1583 ();
 sg13g2_decap_4 FILLER_54_1598 ();
 sg13g2_fill_1 FILLER_54_1616 ();
 sg13g2_fill_1 FILLER_54_1623 ();
 sg13g2_fill_1 FILLER_54_1628 ();
 sg13g2_fill_1 FILLER_54_1640 ();
 sg13g2_decap_4 FILLER_54_1655 ();
 sg13g2_fill_2 FILLER_54_1659 ();
 sg13g2_decap_4 FILLER_54_1667 ();
 sg13g2_fill_1 FILLER_54_1671 ();
 sg13g2_fill_1 FILLER_54_1676 ();
 sg13g2_decap_4 FILLER_54_1685 ();
 sg13g2_fill_2 FILLER_54_1699 ();
 sg13g2_fill_1 FILLER_54_1701 ();
 sg13g2_fill_2 FILLER_54_1706 ();
 sg13g2_fill_1 FILLER_54_1708 ();
 sg13g2_decap_4 FILLER_54_1714 ();
 sg13g2_fill_1 FILLER_54_1718 ();
 sg13g2_fill_1 FILLER_54_1729 ();
 sg13g2_decap_4 FILLER_54_1740 ();
 sg13g2_fill_1 FILLER_54_1744 ();
 sg13g2_decap_4 FILLER_54_1750 ();
 sg13g2_fill_1 FILLER_54_1754 ();
 sg13g2_fill_2 FILLER_54_1759 ();
 sg13g2_decap_4 FILLER_54_1777 ();
 sg13g2_decap_4 FILLER_54_1797 ();
 sg13g2_fill_1 FILLER_54_1801 ();
 sg13g2_fill_1 FILLER_54_1836 ();
 sg13g2_fill_1 FILLER_54_1842 ();
 sg13g2_decap_4 FILLER_54_1863 ();
 sg13g2_fill_2 FILLER_54_1867 ();
 sg13g2_fill_2 FILLER_54_1879 ();
 sg13g2_decap_4 FILLER_54_1889 ();
 sg13g2_decap_8 FILLER_54_1928 ();
 sg13g2_decap_4 FILLER_54_1935 ();
 sg13g2_fill_1 FILLER_54_1939 ();
 sg13g2_decap_8 FILLER_54_1952 ();
 sg13g2_fill_2 FILLER_54_1959 ();
 sg13g2_fill_1 FILLER_54_1961 ();
 sg13g2_fill_2 FILLER_54_1996 ();
 sg13g2_fill_1 FILLER_54_2003 ();
 sg13g2_fill_1 FILLER_54_2013 ();
 sg13g2_fill_1 FILLER_54_2049 ();
 sg13g2_fill_1 FILLER_54_2054 ();
 sg13g2_decap_8 FILLER_54_2086 ();
 sg13g2_decap_4 FILLER_54_2093 ();
 sg13g2_fill_2 FILLER_54_2097 ();
 sg13g2_fill_2 FILLER_54_2109 ();
 sg13g2_fill_1 FILLER_54_2111 ();
 sg13g2_fill_2 FILLER_54_2137 ();
 sg13g2_fill_1 FILLER_54_2143 ();
 sg13g2_decap_8 FILLER_54_2163 ();
 sg13g2_decap_8 FILLER_54_2170 ();
 sg13g2_decap_8 FILLER_54_2177 ();
 sg13g2_decap_8 FILLER_54_2184 ();
 sg13g2_decap_8 FILLER_54_2191 ();
 sg13g2_fill_2 FILLER_54_2198 ();
 sg13g2_fill_1 FILLER_54_2200 ();
 sg13g2_decap_8 FILLER_54_2247 ();
 sg13g2_decap_4 FILLER_54_2254 ();
 sg13g2_fill_2 FILLER_54_2258 ();
 sg13g2_fill_1 FILLER_54_2320 ();
 sg13g2_decap_8 FILLER_54_2350 ();
 sg13g2_decap_8 FILLER_54_2357 ();
 sg13g2_fill_2 FILLER_54_2364 ();
 sg13g2_decap_4 FILLER_54_2370 ();
 sg13g2_fill_1 FILLER_54_2374 ();
 sg13g2_fill_1 FILLER_54_2388 ();
 sg13g2_decap_8 FILLER_54_2433 ();
 sg13g2_decap_4 FILLER_54_2440 ();
 sg13g2_fill_2 FILLER_54_2444 ();
 sg13g2_fill_1 FILLER_54_2450 ();
 sg13g2_fill_2 FILLER_54_2455 ();
 sg13g2_fill_1 FILLER_54_2457 ();
 sg13g2_fill_1 FILLER_54_2489 ();
 sg13g2_fill_2 FILLER_54_2498 ();
 sg13g2_fill_1 FILLER_54_2500 ();
 sg13g2_decap_4 FILLER_54_2527 ();
 sg13g2_fill_1 FILLER_54_2531 ();
 sg13g2_decap_4 FILLER_54_2583 ();
 sg13g2_fill_2 FILLER_54_2639 ();
 sg13g2_fill_2 FILLER_54_2667 ();
 sg13g2_fill_1 FILLER_54_2669 ();
 sg13g2_decap_8 FILLER_55_0 ();
 sg13g2_decap_8 FILLER_55_7 ();
 sg13g2_fill_2 FILLER_55_18 ();
 sg13g2_decap_8 FILLER_55_43 ();
 sg13g2_fill_1 FILLER_55_50 ();
 sg13g2_decap_4 FILLER_55_59 ();
 sg13g2_fill_1 FILLER_55_67 ();
 sg13g2_decap_8 FILLER_55_100 ();
 sg13g2_decap_4 FILLER_55_107 ();
 sg13g2_fill_2 FILLER_55_116 ();
 sg13g2_fill_1 FILLER_55_118 ();
 sg13g2_decap_8 FILLER_55_123 ();
 sg13g2_fill_2 FILLER_55_130 ();
 sg13g2_fill_1 FILLER_55_132 ();
 sg13g2_fill_2 FILLER_55_142 ();
 sg13g2_fill_1 FILLER_55_144 ();
 sg13g2_decap_4 FILLER_55_149 ();
 sg13g2_fill_2 FILLER_55_153 ();
 sg13g2_decap_8 FILLER_55_165 ();
 sg13g2_fill_2 FILLER_55_172 ();
 sg13g2_decap_4 FILLER_55_178 ();
 sg13g2_fill_1 FILLER_55_182 ();
 sg13g2_decap_8 FILLER_55_192 ();
 sg13g2_decap_4 FILLER_55_199 ();
 sg13g2_decap_8 FILLER_55_207 ();
 sg13g2_fill_1 FILLER_55_214 ();
 sg13g2_fill_2 FILLER_55_252 ();
 sg13g2_fill_1 FILLER_55_254 ();
 sg13g2_decap_8 FILLER_55_278 ();
 sg13g2_fill_2 FILLER_55_285 ();
 sg13g2_fill_2 FILLER_55_304 ();
 sg13g2_fill_1 FILLER_55_344 ();
 sg13g2_fill_2 FILLER_55_388 ();
 sg13g2_fill_2 FILLER_55_394 ();
 sg13g2_fill_2 FILLER_55_401 ();
 sg13g2_fill_2 FILLER_55_416 ();
 sg13g2_fill_2 FILLER_55_422 ();
 sg13g2_fill_2 FILLER_55_436 ();
 sg13g2_fill_1 FILLER_55_443 ();
 sg13g2_decap_8 FILLER_55_549 ();
 sg13g2_fill_1 FILLER_55_592 ();
 sg13g2_fill_2 FILLER_55_630 ();
 sg13g2_fill_2 FILLER_55_637 ();
 sg13g2_fill_1 FILLER_55_639 ();
 sg13g2_decap_4 FILLER_55_699 ();
 sg13g2_fill_1 FILLER_55_711 ();
 sg13g2_fill_1 FILLER_55_746 ();
 sg13g2_fill_1 FILLER_55_795 ();
 sg13g2_decap_4 FILLER_55_821 ();
 sg13g2_fill_1 FILLER_55_836 ();
 sg13g2_fill_1 FILLER_55_847 ();
 sg13g2_decap_4 FILLER_55_859 ();
 sg13g2_fill_1 FILLER_55_863 ();
 sg13g2_decap_4 FILLER_55_869 ();
 sg13g2_fill_2 FILLER_55_901 ();
 sg13g2_fill_1 FILLER_55_908 ();
 sg13g2_fill_1 FILLER_55_913 ();
 sg13g2_fill_1 FILLER_55_1023 ();
 sg13g2_fill_1 FILLER_55_1029 ();
 sg13g2_fill_2 FILLER_55_1079 ();
 sg13g2_fill_2 FILLER_55_1107 ();
 sg13g2_fill_1 FILLER_55_1109 ();
 sg13g2_fill_1 FILLER_55_1133 ();
 sg13g2_decap_4 FILLER_55_1160 ();
 sg13g2_decap_8 FILLER_55_1194 ();
 sg13g2_decap_4 FILLER_55_1201 ();
 sg13g2_decap_4 FILLER_55_1209 ();
 sg13g2_decap_4 FILLER_55_1223 ();
 sg13g2_fill_1 FILLER_55_1227 ();
 sg13g2_decap_4 FILLER_55_1240 ();
 sg13g2_fill_1 FILLER_55_1260 ();
 sg13g2_decap_8 FILLER_55_1269 ();
 sg13g2_decap_4 FILLER_55_1305 ();
 sg13g2_fill_1 FILLER_55_1309 ();
 sg13g2_fill_2 FILLER_55_1315 ();
 sg13g2_decap_4 FILLER_55_1337 ();
 sg13g2_fill_1 FILLER_55_1341 ();
 sg13g2_fill_1 FILLER_55_1377 ();
 sg13g2_fill_2 FILLER_55_1414 ();
 sg13g2_fill_2 FILLER_55_1468 ();
 sg13g2_fill_1 FILLER_55_1538 ();
 sg13g2_fill_2 FILLER_55_1576 ();
 sg13g2_fill_1 FILLER_55_1578 ();
 sg13g2_fill_2 FILLER_55_1592 ();
 sg13g2_fill_2 FILLER_55_1597 ();
 sg13g2_fill_1 FILLER_55_1599 ();
 sg13g2_fill_2 FILLER_55_1611 ();
 sg13g2_fill_2 FILLER_55_1622 ();
 sg13g2_fill_1 FILLER_55_1644 ();
 sg13g2_fill_1 FILLER_55_1650 ();
 sg13g2_decap_4 FILLER_55_1659 ();
 sg13g2_fill_1 FILLER_55_1663 ();
 sg13g2_decap_4 FILLER_55_1678 ();
 sg13g2_fill_1 FILLER_55_1714 ();
 sg13g2_fill_2 FILLER_55_1723 ();
 sg13g2_fill_1 FILLER_55_1725 ();
 sg13g2_fill_1 FILLER_55_1730 ();
 sg13g2_fill_1 FILLER_55_1770 ();
 sg13g2_fill_1 FILLER_55_1780 ();
 sg13g2_fill_2 FILLER_55_1786 ();
 sg13g2_decap_8 FILLER_55_1796 ();
 sg13g2_fill_2 FILLER_55_1811 ();
 sg13g2_decap_4 FILLER_55_1821 ();
 sg13g2_fill_2 FILLER_55_1825 ();
 sg13g2_fill_1 FILLER_55_1831 ();
 sg13g2_fill_1 FILLER_55_1840 ();
 sg13g2_fill_2 FILLER_55_1846 ();
 sg13g2_decap_4 FILLER_55_1856 ();
 sg13g2_decap_4 FILLER_55_1869 ();
 sg13g2_fill_1 FILLER_55_1873 ();
 sg13g2_decap_4 FILLER_55_1879 ();
 sg13g2_fill_2 FILLER_55_1887 ();
 sg13g2_fill_1 FILLER_55_1889 ();
 sg13g2_fill_1 FILLER_55_1898 ();
 sg13g2_fill_1 FILLER_55_1904 ();
 sg13g2_fill_2 FILLER_55_1922 ();
 sg13g2_fill_2 FILLER_55_1932 ();
 sg13g2_fill_1 FILLER_55_1934 ();
 sg13g2_fill_1 FILLER_55_1940 ();
 sg13g2_fill_2 FILLER_55_1946 ();
 sg13g2_fill_1 FILLER_55_1948 ();
 sg13g2_decap_8 FILLER_55_1954 ();
 sg13g2_fill_2 FILLER_55_1961 ();
 sg13g2_decap_8 FILLER_55_1993 ();
 sg13g2_fill_2 FILLER_55_2000 ();
 sg13g2_fill_1 FILLER_55_2002 ();
 sg13g2_fill_1 FILLER_55_2008 ();
 sg13g2_fill_1 FILLER_55_2014 ();
 sg13g2_fill_1 FILLER_55_2050 ();
 sg13g2_decap_8 FILLER_55_2090 ();
 sg13g2_decap_4 FILLER_55_2185 ();
 sg13g2_fill_2 FILLER_55_2189 ();
 sg13g2_fill_2 FILLER_55_2227 ();
 sg13g2_fill_2 FILLER_55_2255 ();
 sg13g2_fill_1 FILLER_55_2257 ();
 sg13g2_decap_8 FILLER_55_2304 ();
 sg13g2_decap_8 FILLER_55_2353 ();
 sg13g2_decap_8 FILLER_55_2360 ();
 sg13g2_fill_2 FILLER_55_2367 ();
 sg13g2_fill_2 FILLER_55_2392 ();
 sg13g2_fill_2 FILLER_55_2420 ();
 sg13g2_decap_8 FILLER_55_2434 ();
 sg13g2_fill_1 FILLER_55_2441 ();
 sg13g2_fill_2 FILLER_55_2453 ();
 sg13g2_fill_1 FILLER_55_2455 ();
 sg13g2_fill_1 FILLER_55_2520 ();
 sg13g2_fill_1 FILLER_55_2562 ();
 sg13g2_decap_8 FILLER_55_2567 ();
 sg13g2_decap_8 FILLER_55_2574 ();
 sg13g2_decap_4 FILLER_55_2665 ();
 sg13g2_fill_1 FILLER_55_2669 ();
 sg13g2_fill_2 FILLER_56_0 ();
 sg13g2_fill_1 FILLER_56_33 ();
 sg13g2_fill_1 FILLER_56_39 ();
 sg13g2_decap_8 FILLER_56_45 ();
 sg13g2_decap_8 FILLER_56_52 ();
 sg13g2_fill_2 FILLER_56_106 ();
 sg13g2_fill_2 FILLER_56_134 ();
 sg13g2_fill_1 FILLER_56_136 ();
 sg13g2_decap_8 FILLER_56_147 ();
 sg13g2_decap_4 FILLER_56_154 ();
 sg13g2_fill_2 FILLER_56_158 ();
 sg13g2_decap_4 FILLER_56_180 ();
 sg13g2_decap_8 FILLER_56_189 ();
 sg13g2_fill_1 FILLER_56_196 ();
 sg13g2_fill_1 FILLER_56_202 ();
 sg13g2_fill_1 FILLER_56_224 ();
 sg13g2_fill_2 FILLER_56_262 ();
 sg13g2_decap_4 FILLER_56_294 ();
 sg13g2_fill_2 FILLER_56_334 ();
 sg13g2_fill_2 FILLER_56_366 ();
 sg13g2_fill_2 FILLER_56_376 ();
 sg13g2_fill_1 FILLER_56_408 ();
 sg13g2_decap_8 FILLER_56_419 ();
 sg13g2_fill_1 FILLER_56_426 ();
 sg13g2_fill_1 FILLER_56_467 ();
 sg13g2_fill_2 FILLER_56_501 ();
 sg13g2_fill_2 FILLER_56_523 ();
 sg13g2_fill_1 FILLER_56_525 ();
 sg13g2_fill_1 FILLER_56_536 ();
 sg13g2_fill_1 FILLER_56_547 ();
 sg13g2_fill_1 FILLER_56_574 ();
 sg13g2_decap_4 FILLER_56_579 ();
 sg13g2_fill_1 FILLER_56_583 ();
 sg13g2_fill_2 FILLER_56_635 ();
 sg13g2_fill_2 FILLER_56_663 ();
 sg13g2_decap_8 FILLER_56_872 ();
 sg13g2_fill_2 FILLER_56_879 ();
 sg13g2_fill_1 FILLER_56_881 ();
 sg13g2_fill_1 FILLER_56_890 ();
 sg13g2_fill_2 FILLER_56_895 ();
 sg13g2_fill_2 FILLER_56_902 ();
 sg13g2_fill_1 FILLER_56_909 ();
 sg13g2_fill_1 FILLER_56_919 ();
 sg13g2_fill_1 FILLER_56_935 ();
 sg13g2_fill_2 FILLER_56_949 ();
 sg13g2_fill_1 FILLER_56_963 ();
 sg13g2_fill_2 FILLER_56_975 ();
 sg13g2_fill_1 FILLER_56_1013 ();
 sg13g2_fill_1 FILLER_56_1032 ();
 sg13g2_fill_2 FILLER_56_1053 ();
 sg13g2_fill_1 FILLER_56_1066 ();
 sg13g2_fill_2 FILLER_56_1092 ();
 sg13g2_fill_1 FILLER_56_1094 ();
 sg13g2_fill_2 FILLER_56_1121 ();
 sg13g2_fill_1 FILLER_56_1130 ();
 sg13g2_fill_2 FILLER_56_1193 ();
 sg13g2_fill_1 FILLER_56_1195 ();
 sg13g2_fill_1 FILLER_56_1233 ();
 sg13g2_fill_2 FILLER_56_1249 ();
 sg13g2_fill_1 FILLER_56_1251 ();
 sg13g2_fill_1 FILLER_56_1260 ();
 sg13g2_fill_2 FILLER_56_1266 ();
 sg13g2_fill_1 FILLER_56_1268 ();
 sg13g2_fill_1 FILLER_56_1275 ();
 sg13g2_fill_1 FILLER_56_1280 ();
 sg13g2_fill_1 FILLER_56_1287 ();
 sg13g2_decap_8 FILLER_56_1299 ();
 sg13g2_fill_2 FILLER_56_1310 ();
 sg13g2_fill_1 FILLER_56_1312 ();
 sg13g2_decap_8 FILLER_56_1318 ();
 sg13g2_decap_8 FILLER_56_1325 ();
 sg13g2_fill_1 FILLER_56_1332 ();
 sg13g2_fill_2 FILLER_56_1338 ();
 sg13g2_decap_4 FILLER_56_1360 ();
 sg13g2_decap_8 FILLER_56_1368 ();
 sg13g2_fill_2 FILLER_56_1375 ();
 sg13g2_fill_1 FILLER_56_1398 ();
 sg13g2_fill_2 FILLER_56_1407 ();
 sg13g2_fill_2 FILLER_56_1431 ();
 sg13g2_fill_2 FILLER_56_1440 ();
 sg13g2_fill_2 FILLER_56_1450 ();
 sg13g2_fill_1 FILLER_56_1462 ();
 sg13g2_fill_2 FILLER_56_1468 ();
 sg13g2_fill_2 FILLER_56_1478 ();
 sg13g2_fill_2 FILLER_56_1497 ();
 sg13g2_fill_1 FILLER_56_1526 ();
 sg13g2_fill_1 FILLER_56_1534 ();
 sg13g2_fill_2 FILLER_56_1543 ();
 sg13g2_fill_2 FILLER_56_1566 ();
 sg13g2_decap_4 FILLER_56_1585 ();
 sg13g2_fill_1 FILLER_56_1589 ();
 sg13g2_fill_1 FILLER_56_1612 ();
 sg13g2_fill_1 FILLER_56_1649 ();
 sg13g2_fill_1 FILLER_56_1655 ();
 sg13g2_fill_1 FILLER_56_1660 ();
 sg13g2_decap_4 FILLER_56_1674 ();
 sg13g2_fill_1 FILLER_56_1688 ();
 sg13g2_fill_2 FILLER_56_1725 ();
 sg13g2_fill_1 FILLER_56_1743 ();
 sg13g2_fill_2 FILLER_56_1758 ();
 sg13g2_decap_4 FILLER_56_1764 ();
 sg13g2_fill_2 FILLER_56_1768 ();
 sg13g2_fill_2 FILLER_56_1807 ();
 sg13g2_fill_1 FILLER_56_1809 ();
 sg13g2_fill_2 FILLER_56_1824 ();
 sg13g2_decap_4 FILLER_56_1836 ();
 sg13g2_fill_2 FILLER_56_1840 ();
 sg13g2_decap_8 FILLER_56_1847 ();
 sg13g2_decap_8 FILLER_56_1854 ();
 sg13g2_decap_8 FILLER_56_1861 ();
 sg13g2_fill_2 FILLER_56_1868 ();
 sg13g2_fill_2 FILLER_56_1879 ();
 sg13g2_fill_1 FILLER_56_1907 ();
 sg13g2_decap_8 FILLER_56_1916 ();
 sg13g2_fill_2 FILLER_56_1927 ();
 sg13g2_decap_4 FILLER_56_1934 ();
 sg13g2_decap_8 FILLER_56_1946 ();
 sg13g2_decap_8 FILLER_56_1953 ();
 sg13g2_decap_8 FILLER_56_1960 ();
 sg13g2_fill_1 FILLER_56_1967 ();
 sg13g2_fill_1 FILLER_56_1977 ();
 sg13g2_fill_2 FILLER_56_1983 ();
 sg13g2_fill_1 FILLER_56_1985 ();
 sg13g2_decap_8 FILLER_56_2002 ();
 sg13g2_fill_2 FILLER_56_2009 ();
 sg13g2_fill_1 FILLER_56_2011 ();
 sg13g2_fill_1 FILLER_56_2040 ();
 sg13g2_fill_2 FILLER_56_2046 ();
 sg13g2_decap_8 FILLER_56_2085 ();
 sg13g2_decap_4 FILLER_56_2092 ();
 sg13g2_fill_2 FILLER_56_2096 ();
 sg13g2_fill_1 FILLER_56_2177 ();
 sg13g2_fill_2 FILLER_56_2204 ();
 sg13g2_fill_1 FILLER_56_2206 ();
 sg13g2_decap_4 FILLER_56_2247 ();
 sg13g2_fill_2 FILLER_56_2251 ();
 sg13g2_decap_4 FILLER_56_2263 ();
 sg13g2_fill_2 FILLER_56_2267 ();
 sg13g2_fill_2 FILLER_56_2287 ();
 sg13g2_decap_4 FILLER_56_2331 ();
 sg13g2_fill_1 FILLER_56_2339 ();
 sg13g2_decap_8 FILLER_56_2345 ();
 sg13g2_decap_8 FILLER_56_2352 ();
 sg13g2_decap_4 FILLER_56_2359 ();
 sg13g2_fill_2 FILLER_56_2363 ();
 sg13g2_fill_1 FILLER_56_2373 ();
 sg13g2_fill_1 FILLER_56_2403 ();
 sg13g2_fill_1 FILLER_56_2515 ();
 sg13g2_decap_4 FILLER_56_2575 ();
 sg13g2_fill_1 FILLER_56_2579 ();
 sg13g2_fill_2 FILLER_56_2610 ();
 sg13g2_fill_1 FILLER_56_2616 ();
 sg13g2_decap_4 FILLER_56_2666 ();
 sg13g2_decap_8 FILLER_57_0 ();
 sg13g2_decap_4 FILLER_57_7 ();
 sg13g2_fill_1 FILLER_57_11 ();
 sg13g2_decap_8 FILLER_57_60 ();
 sg13g2_decap_4 FILLER_57_67 ();
 sg13g2_decap_4 FILLER_57_76 ();
 sg13g2_decap_4 FILLER_57_84 ();
 sg13g2_fill_1 FILLER_57_88 ();
 sg13g2_fill_1 FILLER_57_114 ();
 sg13g2_decap_4 FILLER_57_119 ();
 sg13g2_fill_2 FILLER_57_123 ();
 sg13g2_fill_1 FILLER_57_139 ();
 sg13g2_decap_4 FILLER_57_153 ();
 sg13g2_decap_4 FILLER_57_187 ();
 sg13g2_decap_4 FILLER_57_239 ();
 sg13g2_fill_1 FILLER_57_261 ();
 sg13g2_fill_1 FILLER_57_267 ();
 sg13g2_fill_1 FILLER_57_298 ();
 sg13g2_fill_1 FILLER_57_339 ();
 sg13g2_fill_2 FILLER_57_348 ();
 sg13g2_fill_2 FILLER_57_376 ();
 sg13g2_decap_8 FILLER_57_417 ();
 sg13g2_fill_2 FILLER_57_433 ();
 sg13g2_fill_1 FILLER_57_449 ();
 sg13g2_fill_1 FILLER_57_455 ();
 sg13g2_fill_2 FILLER_57_501 ();
 sg13g2_fill_2 FILLER_57_533 ();
 sg13g2_fill_2 FILLER_57_561 ();
 sg13g2_fill_2 FILLER_57_589 ();
 sg13g2_fill_1 FILLER_57_591 ();
 sg13g2_decap_4 FILLER_57_653 ();
 sg13g2_fill_1 FILLER_57_657 ();
 sg13g2_fill_1 FILLER_57_667 ();
 sg13g2_fill_2 FILLER_57_711 ();
 sg13g2_fill_1 FILLER_57_774 ();
 sg13g2_fill_1 FILLER_57_794 ();
 sg13g2_fill_2 FILLER_57_859 ();
 sg13g2_fill_2 FILLER_57_865 ();
 sg13g2_fill_2 FILLER_57_899 ();
 sg13g2_decap_8 FILLER_57_931 ();
 sg13g2_decap_8 FILLER_57_948 ();
 sg13g2_fill_2 FILLER_57_955 ();
 sg13g2_fill_1 FILLER_57_957 ();
 sg13g2_fill_2 FILLER_57_968 ();
 sg13g2_fill_2 FILLER_57_980 ();
 sg13g2_fill_1 FILLER_57_998 ();
 sg13g2_fill_2 FILLER_57_1038 ();
 sg13g2_fill_2 FILLER_57_1069 ();
 sg13g2_fill_1 FILLER_57_1071 ();
 sg13g2_decap_8 FILLER_57_1106 ();
 sg13g2_decap_8 FILLER_57_1113 ();
 sg13g2_decap_4 FILLER_57_1120 ();
 sg13g2_fill_2 FILLER_57_1124 ();
 sg13g2_fill_2 FILLER_57_1132 ();
 sg13g2_decap_8 FILLER_57_1176 ();
 sg13g2_decap_4 FILLER_57_1183 ();
 sg13g2_fill_1 FILLER_57_1187 ();
 sg13g2_fill_1 FILLER_57_1196 ();
 sg13g2_fill_1 FILLER_57_1200 ();
 sg13g2_fill_1 FILLER_57_1216 ();
 sg13g2_decap_4 FILLER_57_1234 ();
 sg13g2_fill_2 FILLER_57_1238 ();
 sg13g2_fill_1 FILLER_57_1261 ();
 sg13g2_fill_1 FILLER_57_1267 ();
 sg13g2_fill_2 FILLER_57_1273 ();
 sg13g2_fill_1 FILLER_57_1275 ();
 sg13g2_fill_2 FILLER_57_1282 ();
 sg13g2_fill_1 FILLER_57_1300 ();
 sg13g2_decap_4 FILLER_57_1306 ();
 sg13g2_fill_2 FILLER_57_1310 ();
 sg13g2_fill_2 FILLER_57_1317 ();
 sg13g2_fill_2 FILLER_57_1332 ();
 sg13g2_fill_1 FILLER_57_1334 ();
 sg13g2_fill_1 FILLER_57_1340 ();
 sg13g2_fill_1 FILLER_57_1353 ();
 sg13g2_fill_2 FILLER_57_1358 ();
 sg13g2_decap_4 FILLER_57_1375 ();
 sg13g2_decap_8 FILLER_57_1397 ();
 sg13g2_fill_2 FILLER_57_1404 ();
 sg13g2_fill_2 FILLER_57_1430 ();
 sg13g2_fill_1 FILLER_57_1443 ();
 sg13g2_fill_2 FILLER_57_1457 ();
 sg13g2_fill_1 FILLER_57_1530 ();
 sg13g2_fill_2 FILLER_57_1562 ();
 sg13g2_fill_2 FILLER_57_1571 ();
 sg13g2_fill_1 FILLER_57_1586 ();
 sg13g2_fill_1 FILLER_57_1593 ();
 sg13g2_fill_1 FILLER_57_1602 ();
 sg13g2_fill_2 FILLER_57_1650 ();
 sg13g2_decap_4 FILLER_57_1685 ();
 sg13g2_fill_2 FILLER_57_1692 ();
 sg13g2_decap_4 FILLER_57_1699 ();
 sg13g2_fill_2 FILLER_57_1703 ();
 sg13g2_decap_4 FILLER_57_1709 ();
 sg13g2_decap_8 FILLER_57_1720 ();
 sg13g2_fill_2 FILLER_57_1732 ();
 sg13g2_fill_1 FILLER_57_1734 ();
 sg13g2_decap_8 FILLER_57_1740 ();
 sg13g2_fill_2 FILLER_57_1747 ();
 sg13g2_fill_1 FILLER_57_1749 ();
 sg13g2_decap_8 FILLER_57_1755 ();
 sg13g2_fill_2 FILLER_57_1762 ();
 sg13g2_fill_2 FILLER_57_1767 ();
 sg13g2_fill_1 FILLER_57_1769 ();
 sg13g2_fill_2 FILLER_57_1785 ();
 sg13g2_fill_1 FILLER_57_1791 ();
 sg13g2_fill_2 FILLER_57_1813 ();
 sg13g2_fill_1 FILLER_57_1820 ();
 sg13g2_decap_8 FILLER_57_1826 ();
 sg13g2_decap_8 FILLER_57_1833 ();
 sg13g2_decap_4 FILLER_57_1840 ();
 sg13g2_fill_1 FILLER_57_1844 ();
 sg13g2_decap_8 FILLER_57_1855 ();
 sg13g2_decap_4 FILLER_57_1862 ();
 sg13g2_decap_8 FILLER_57_1879 ();
 sg13g2_fill_1 FILLER_57_1886 ();
 sg13g2_fill_2 FILLER_57_1904 ();
 sg13g2_fill_1 FILLER_57_1906 ();
 sg13g2_fill_2 FILLER_57_1911 ();
 sg13g2_fill_1 FILLER_57_1913 ();
 sg13g2_fill_2 FILLER_57_1918 ();
 sg13g2_fill_2 FILLER_57_1930 ();
 sg13g2_fill_1 FILLER_57_1932 ();
 sg13g2_fill_2 FILLER_57_1947 ();
 sg13g2_fill_1 FILLER_57_1949 ();
 sg13g2_decap_8 FILLER_57_1955 ();
 sg13g2_fill_2 FILLER_57_1962 ();
 sg13g2_fill_2 FILLER_57_1977 ();
 sg13g2_fill_1 FILLER_57_1985 ();
 sg13g2_decap_8 FILLER_57_2000 ();
 sg13g2_fill_1 FILLER_57_2007 ();
 sg13g2_fill_1 FILLER_57_2016 ();
 sg13g2_fill_1 FILLER_57_2023 ();
 sg13g2_fill_2 FILLER_57_2065 ();
 sg13g2_fill_1 FILLER_57_2067 ();
 sg13g2_decap_4 FILLER_57_2073 ();
 sg13g2_decap_4 FILLER_57_2082 ();
 sg13g2_fill_1 FILLER_57_2086 ();
 sg13g2_fill_2 FILLER_57_2095 ();
 sg13g2_fill_1 FILLER_57_2097 ();
 sg13g2_fill_1 FILLER_57_2109 ();
 sg13g2_fill_1 FILLER_57_2130 ();
 sg13g2_decap_4 FILLER_57_2170 ();
 sg13g2_decap_8 FILLER_57_2208 ();
 sg13g2_fill_2 FILLER_57_2215 ();
 sg13g2_fill_1 FILLER_57_2217 ();
 sg13g2_decap_4 FILLER_57_2254 ();
 sg13g2_fill_1 FILLER_57_2258 ();
 sg13g2_fill_1 FILLER_57_2263 ();
 sg13g2_fill_2 FILLER_57_2306 ();
 sg13g2_decap_4 FILLER_57_2338 ();
 sg13g2_fill_2 FILLER_57_2342 ();
 sg13g2_fill_2 FILLER_57_2353 ();
 sg13g2_fill_1 FILLER_57_2355 ();
 sg13g2_decap_4 FILLER_57_2369 ();
 sg13g2_decap_4 FILLER_57_2377 ();
 sg13g2_fill_2 FILLER_57_2381 ();
 sg13g2_decap_4 FILLER_57_2387 ();
 sg13g2_fill_1 FILLER_57_2391 ();
 sg13g2_fill_2 FILLER_57_2405 ();
 sg13g2_fill_1 FILLER_57_2407 ();
 sg13g2_fill_1 FILLER_57_2422 ();
 sg13g2_fill_1 FILLER_57_2453 ();
 sg13g2_fill_1 FILLER_57_2458 ();
 sg13g2_fill_1 FILLER_57_2464 ();
 sg13g2_fill_1 FILLER_57_2469 ();
 sg13g2_decap_8 FILLER_57_2474 ();
 sg13g2_fill_1 FILLER_57_2481 ();
 sg13g2_decap_8 FILLER_57_2488 ();
 sg13g2_fill_2 FILLER_57_2495 ();
 sg13g2_fill_1 FILLER_57_2497 ();
 sg13g2_decap_8 FILLER_57_2506 ();
 sg13g2_decap_8 FILLER_57_2513 ();
 sg13g2_decap_4 FILLER_57_2520 ();
 sg13g2_decap_4 FILLER_57_2541 ();
 sg13g2_fill_1 FILLER_57_2545 ();
 sg13g2_fill_2 FILLER_57_2572 ();
 sg13g2_decap_8 FILLER_57_2604 ();
 sg13g2_decap_8 FILLER_57_2611 ();
 sg13g2_decap_8 FILLER_57_2658 ();
 sg13g2_decap_4 FILLER_57_2665 ();
 sg13g2_fill_1 FILLER_57_2669 ();
 sg13g2_decap_4 FILLER_58_0 ();
 sg13g2_fill_1 FILLER_58_4 ();
 sg13g2_decap_4 FILLER_58_9 ();
 sg13g2_fill_2 FILLER_58_13 ();
 sg13g2_fill_2 FILLER_58_25 ();
 sg13g2_fill_1 FILLER_58_35 ();
 sg13g2_decap_8 FILLER_58_71 ();
 sg13g2_fill_1 FILLER_58_78 ();
 sg13g2_decap_4 FILLER_58_84 ();
 sg13g2_decap_4 FILLER_58_97 ();
 sg13g2_decap_4 FILLER_58_105 ();
 sg13g2_fill_1 FILLER_58_139 ();
 sg13g2_fill_2 FILLER_58_170 ();
 sg13g2_fill_1 FILLER_58_217 ();
 sg13g2_decap_4 FILLER_58_248 ();
 sg13g2_fill_2 FILLER_58_252 ();
 sg13g2_fill_1 FILLER_58_290 ();
 sg13g2_fill_1 FILLER_58_296 ();
 sg13g2_fill_1 FILLER_58_307 ();
 sg13g2_fill_1 FILLER_58_315 ();
 sg13g2_fill_1 FILLER_58_354 ();
 sg13g2_fill_1 FILLER_58_364 ();
 sg13g2_fill_1 FILLER_58_375 ();
 sg13g2_fill_2 FILLER_58_395 ();
 sg13g2_fill_2 FILLER_58_403 ();
 sg13g2_decap_8 FILLER_58_414 ();
 sg13g2_decap_4 FILLER_58_427 ();
 sg13g2_fill_1 FILLER_58_436 ();
 sg13g2_fill_2 FILLER_58_446 ();
 sg13g2_fill_2 FILLER_58_464 ();
 sg13g2_fill_2 FILLER_58_470 ();
 sg13g2_fill_1 FILLER_58_485 ();
 sg13g2_fill_2 FILLER_58_512 ();
 sg13g2_fill_1 FILLER_58_514 ();
 sg13g2_decap_4 FILLER_58_527 ();
 sg13g2_fill_2 FILLER_58_537 ();
 sg13g2_fill_2 FILLER_58_547 ();
 sg13g2_fill_1 FILLER_58_549 ();
 sg13g2_fill_2 FILLER_58_554 ();
 sg13g2_fill_1 FILLER_58_556 ();
 sg13g2_fill_2 FILLER_58_567 ();
 sg13g2_fill_1 FILLER_58_569 ();
 sg13g2_decap_8 FILLER_58_574 ();
 sg13g2_decap_8 FILLER_58_581 ();
 sg13g2_decap_8 FILLER_58_588 ();
 sg13g2_fill_1 FILLER_58_595 ();
 sg13g2_decap_4 FILLER_58_609 ();
 sg13g2_fill_1 FILLER_58_613 ();
 sg13g2_decap_8 FILLER_58_623 ();
 sg13g2_fill_2 FILLER_58_656 ();
 sg13g2_fill_1 FILLER_58_721 ();
 sg13g2_fill_1 FILLER_58_816 ();
 sg13g2_fill_2 FILLER_58_827 ();
 sg13g2_fill_1 FILLER_58_871 ();
 sg13g2_fill_1 FILLER_58_937 ();
 sg13g2_decap_8 FILLER_58_946 ();
 sg13g2_decap_4 FILLER_58_953 ();
 sg13g2_fill_2 FILLER_58_957 ();
 sg13g2_fill_2 FILLER_58_989 ();
 sg13g2_fill_1 FILLER_58_1006 ();
 sg13g2_fill_2 FILLER_58_1044 ();
 sg13g2_decap_8 FILLER_58_1074 ();
 sg13g2_fill_1 FILLER_58_1081 ();
 sg13g2_decap_8 FILLER_58_1177 ();
 sg13g2_fill_1 FILLER_58_1184 ();
 sg13g2_decap_8 FILLER_58_1196 ();
 sg13g2_fill_1 FILLER_58_1203 ();
 sg13g2_fill_2 FILLER_58_1221 ();
 sg13g2_fill_1 FILLER_58_1223 ();
 sg13g2_fill_2 FILLER_58_1229 ();
 sg13g2_fill_2 FILLER_58_1239 ();
 sg13g2_fill_1 FILLER_58_1273 ();
 sg13g2_fill_1 FILLER_58_1297 ();
 sg13g2_fill_1 FILLER_58_1315 ();
 sg13g2_fill_1 FILLER_58_1326 ();
 sg13g2_fill_2 FILLER_58_1340 ();
 sg13g2_fill_2 FILLER_58_1351 ();
 sg13g2_decap_4 FILLER_58_1383 ();
 sg13g2_fill_1 FILLER_58_1387 ();
 sg13g2_fill_2 FILLER_58_1398 ();
 sg13g2_decap_8 FILLER_58_1410 ();
 sg13g2_fill_1 FILLER_58_1417 ();
 sg13g2_fill_1 FILLER_58_1472 ();
 sg13g2_fill_1 FILLER_58_1483 ();
 sg13g2_fill_1 FILLER_58_1523 ();
 sg13g2_fill_1 FILLER_58_1554 ();
 sg13g2_fill_2 FILLER_58_1560 ();
 sg13g2_fill_1 FILLER_58_1562 ();
 sg13g2_fill_1 FILLER_58_1589 ();
 sg13g2_fill_2 FILLER_58_1594 ();
 sg13g2_fill_1 FILLER_58_1610 ();
 sg13g2_decap_8 FILLER_58_1675 ();
 sg13g2_decap_8 FILLER_58_1687 ();
 sg13g2_decap_8 FILLER_58_1698 ();
 sg13g2_decap_4 FILLER_58_1705 ();
 sg13g2_fill_1 FILLER_58_1709 ();
 sg13g2_fill_1 FILLER_58_1722 ();
 sg13g2_decap_4 FILLER_58_1727 ();
 sg13g2_fill_1 FILLER_58_1731 ();
 sg13g2_decap_4 FILLER_58_1740 ();
 sg13g2_fill_1 FILLER_58_1744 ();
 sg13g2_decap_8 FILLER_58_1780 ();
 sg13g2_fill_2 FILLER_58_1787 ();
 sg13g2_fill_1 FILLER_58_1789 ();
 sg13g2_fill_1 FILLER_58_1798 ();
 sg13g2_decap_8 FILLER_58_1806 ();
 sg13g2_fill_1 FILLER_58_1813 ();
 sg13g2_fill_2 FILLER_58_1824 ();
 sg13g2_fill_1 FILLER_58_1839 ();
 sg13g2_fill_2 FILLER_58_1874 ();
 sg13g2_fill_1 FILLER_58_1882 ();
 sg13g2_fill_1 FILLER_58_1897 ();
 sg13g2_fill_1 FILLER_58_1903 ();
 sg13g2_fill_1 FILLER_58_1909 ();
 sg13g2_fill_1 FILLER_58_1920 ();
 sg13g2_fill_1 FILLER_58_1940 ();
 sg13g2_fill_2 FILLER_58_1946 ();
 sg13g2_fill_2 FILLER_58_1952 ();
 sg13g2_fill_1 FILLER_58_1954 ();
 sg13g2_fill_2 FILLER_58_1959 ();
 sg13g2_fill_1 FILLER_58_1961 ();
 sg13g2_fill_2 FILLER_58_1967 ();
 sg13g2_decap_4 FILLER_58_1979 ();
 sg13g2_fill_1 FILLER_58_1983 ();
 sg13g2_decap_8 FILLER_58_2006 ();
 sg13g2_decap_4 FILLER_58_2013 ();
 sg13g2_fill_1 FILLER_58_2023 ();
 sg13g2_fill_1 FILLER_58_2031 ();
 sg13g2_fill_1 FILLER_58_2037 ();
 sg13g2_decap_8 FILLER_58_2071 ();
 sg13g2_decap_8 FILLER_58_2078 ();
 sg13g2_fill_1 FILLER_58_2085 ();
 sg13g2_decap_8 FILLER_58_2090 ();
 sg13g2_decap_4 FILLER_58_2097 ();
 sg13g2_fill_1 FILLER_58_2101 ();
 sg13g2_fill_1 FILLER_58_2138 ();
 sg13g2_fill_1 FILLER_58_2174 ();
 sg13g2_decap_8 FILLER_58_2196 ();
 sg13g2_decap_8 FILLER_58_2203 ();
 sg13g2_fill_1 FILLER_58_2210 ();
 sg13g2_decap_8 FILLER_58_2221 ();
 sg13g2_fill_1 FILLER_58_2228 ();
 sg13g2_decap_4 FILLER_58_2233 ();
 sg13g2_decap_8 FILLER_58_2241 ();
 sg13g2_decap_8 FILLER_58_2248 ();
 sg13g2_decap_4 FILLER_58_2255 ();
 sg13g2_fill_2 FILLER_58_2280 ();
 sg13g2_fill_1 FILLER_58_2282 ();
 sg13g2_fill_1 FILLER_58_2288 ();
 sg13g2_decap_4 FILLER_58_2302 ();
 sg13g2_decap_4 FILLER_58_2337 ();
 sg13g2_fill_1 FILLER_58_2341 ();
 sg13g2_decap_8 FILLER_58_2368 ();
 sg13g2_fill_2 FILLER_58_2379 ();
 sg13g2_fill_1 FILLER_58_2411 ();
 sg13g2_fill_2 FILLER_58_2444 ();
 sg13g2_decap_8 FILLER_58_2459 ();
 sg13g2_decap_8 FILLER_58_2466 ();
 sg13g2_fill_2 FILLER_58_2473 ();
 sg13g2_fill_1 FILLER_58_2475 ();
 sg13g2_fill_2 FILLER_58_2485 ();
 sg13g2_fill_2 FILLER_58_2529 ();
 sg13g2_fill_1 FILLER_58_2531 ();
 sg13g2_fill_2 FILLER_58_2564 ();
 sg13g2_fill_1 FILLER_58_2566 ();
 sg13g2_decap_8 FILLER_58_2577 ();
 sg13g2_decap_8 FILLER_58_2584 ();
 sg13g2_decap_8 FILLER_58_2601 ();
 sg13g2_decap_8 FILLER_58_2608 ();
 sg13g2_fill_1 FILLER_58_2615 ();
 sg13g2_fill_2 FILLER_58_2647 ();
 sg13g2_decap_8 FILLER_58_2653 ();
 sg13g2_decap_8 FILLER_58_2660 ();
 sg13g2_fill_2 FILLER_58_2667 ();
 sg13g2_fill_1 FILLER_58_2669 ();
 sg13g2_fill_1 FILLER_59_36 ();
 sg13g2_fill_2 FILLER_59_62 ();
 sg13g2_fill_2 FILLER_59_100 ();
 sg13g2_fill_1 FILLER_59_126 ();
 sg13g2_fill_1 FILLER_59_131 ();
 sg13g2_decap_8 FILLER_59_153 ();
 sg13g2_decap_8 FILLER_59_160 ();
 sg13g2_decap_4 FILLER_59_167 ();
 sg13g2_fill_1 FILLER_59_171 ();
 sg13g2_fill_2 FILLER_59_175 ();
 sg13g2_fill_1 FILLER_59_177 ();
 sg13g2_fill_2 FILLER_59_187 ();
 sg13g2_fill_1 FILLER_59_207 ();
 sg13g2_decap_8 FILLER_59_246 ();
 sg13g2_decap_8 FILLER_59_253 ();
 sg13g2_decap_4 FILLER_59_260 ();
 sg13g2_fill_1 FILLER_59_285 ();
 sg13g2_fill_2 FILLER_59_296 ();
 sg13g2_fill_1 FILLER_59_324 ();
 sg13g2_fill_1 FILLER_59_348 ();
 sg13g2_decap_4 FILLER_59_372 ();
 sg13g2_fill_1 FILLER_59_376 ();
 sg13g2_fill_1 FILLER_59_395 ();
 sg13g2_decap_8 FILLER_59_429 ();
 sg13g2_decap_8 FILLER_59_436 ();
 sg13g2_decap_4 FILLER_59_443 ();
 sg13g2_fill_1 FILLER_59_447 ();
 sg13g2_fill_2 FILLER_59_460 ();
 sg13g2_fill_1 FILLER_59_466 ();
 sg13g2_fill_2 FILLER_59_471 ();
 sg13g2_fill_2 FILLER_59_476 ();
 sg13g2_fill_1 FILLER_59_482 ();
 sg13g2_decap_4 FILLER_59_495 ();
 sg13g2_fill_1 FILLER_59_499 ();
 sg13g2_fill_2 FILLER_59_529 ();
 sg13g2_fill_2 FILLER_59_552 ();
 sg13g2_decap_8 FILLER_59_563 ();
 sg13g2_decap_8 FILLER_59_570 ();
 sg13g2_decap_8 FILLER_59_577 ();
 sg13g2_decap_8 FILLER_59_584 ();
 sg13g2_decap_8 FILLER_59_595 ();
 sg13g2_decap_4 FILLER_59_602 ();
 sg13g2_decap_8 FILLER_59_611 ();
 sg13g2_decap_8 FILLER_59_618 ();
 sg13g2_decap_4 FILLER_59_625 ();
 sg13g2_fill_2 FILLER_59_629 ();
 sg13g2_decap_4 FILLER_59_640 ();
 sg13g2_fill_1 FILLER_59_648 ();
 sg13g2_fill_2 FILLER_59_669 ();
 sg13g2_fill_2 FILLER_59_705 ();
 sg13g2_fill_1 FILLER_59_758 ();
 sg13g2_fill_2 FILLER_59_785 ();
 sg13g2_fill_1 FILLER_59_810 ();
 sg13g2_fill_2 FILLER_59_819 ();
 sg13g2_fill_2 FILLER_59_828 ();
 sg13g2_fill_2 FILLER_59_889 ();
 sg13g2_fill_2 FILLER_59_897 ();
 sg13g2_fill_1 FILLER_59_903 ();
 sg13g2_fill_2 FILLER_59_911 ();
 sg13g2_fill_1 FILLER_59_944 ();
 sg13g2_decap_4 FILLER_59_953 ();
 sg13g2_fill_2 FILLER_59_972 ();
 sg13g2_fill_2 FILLER_59_985 ();
 sg13g2_fill_1 FILLER_59_1001 ();
 sg13g2_fill_1 FILLER_59_1005 ();
 sg13g2_fill_2 FILLER_59_1019 ();
 sg13g2_fill_1 FILLER_59_1034 ();
 sg13g2_fill_2 FILLER_59_1044 ();
 sg13g2_fill_2 FILLER_59_1106 ();
 sg13g2_fill_1 FILLER_59_1108 ();
 sg13g2_fill_1 FILLER_59_1164 ();
 sg13g2_decap_4 FILLER_59_1168 ();
 sg13g2_fill_2 FILLER_59_1175 ();
 sg13g2_fill_2 FILLER_59_1181 ();
 sg13g2_fill_2 FILLER_59_1188 ();
 sg13g2_fill_1 FILLER_59_1190 ();
 sg13g2_fill_2 FILLER_59_1195 ();
 sg13g2_fill_1 FILLER_59_1197 ();
 sg13g2_fill_1 FILLER_59_1211 ();
 sg13g2_fill_2 FILLER_59_1222 ();
 sg13g2_fill_1 FILLER_59_1235 ();
 sg13g2_fill_1 FILLER_59_1249 ();
 sg13g2_decap_8 FILLER_59_1259 ();
 sg13g2_decap_4 FILLER_59_1266 ();
 sg13g2_fill_1 FILLER_59_1276 ();
 sg13g2_decap_8 FILLER_59_1282 ();
 sg13g2_decap_8 FILLER_59_1289 ();
 sg13g2_decap_8 FILLER_59_1296 ();
 sg13g2_fill_2 FILLER_59_1308 ();
 sg13g2_decap_8 FILLER_59_1325 ();
 sg13g2_decap_4 FILLER_59_1332 ();
 sg13g2_fill_2 FILLER_59_1340 ();
 sg13g2_fill_1 FILLER_59_1342 ();
 sg13g2_fill_2 FILLER_59_1353 ();
 sg13g2_fill_2 FILLER_59_1371 ();
 sg13g2_decap_4 FILLER_59_1387 ();
 sg13g2_fill_2 FILLER_59_1391 ();
 sg13g2_fill_1 FILLER_59_1410 ();
 sg13g2_decap_8 FILLER_59_1416 ();
 sg13g2_decap_4 FILLER_59_1423 ();
 sg13g2_decap_8 FILLER_59_1431 ();
 sg13g2_fill_2 FILLER_59_1445 ();
 sg13g2_fill_1 FILLER_59_1468 ();
 sg13g2_fill_1 FILLER_59_1474 ();
 sg13g2_fill_1 FILLER_59_1505 ();
 sg13g2_decap_4 FILLER_59_1553 ();
 sg13g2_fill_1 FILLER_59_1557 ();
 sg13g2_decap_4 FILLER_59_1563 ();
 sg13g2_fill_1 FILLER_59_1567 ();
 sg13g2_decap_8 FILLER_59_1580 ();
 sg13g2_fill_1 FILLER_59_1587 ();
 sg13g2_fill_2 FILLER_59_1592 ();
 sg13g2_decap_4 FILLER_59_1614 ();
 sg13g2_fill_2 FILLER_59_1618 ();
 sg13g2_decap_4 FILLER_59_1667 ();
 sg13g2_fill_1 FILLER_59_1671 ();
 sg13g2_fill_2 FILLER_59_1709 ();
 sg13g2_decap_4 FILLER_59_1715 ();
 sg13g2_fill_1 FILLER_59_1719 ();
 sg13g2_decap_8 FILLER_59_1729 ();
 sg13g2_decap_4 FILLER_59_1766 ();
 sg13g2_fill_1 FILLER_59_1770 ();
 sg13g2_fill_2 FILLER_59_1775 ();
 sg13g2_fill_1 FILLER_59_1777 ();
 sg13g2_fill_1 FILLER_59_1804 ();
 sg13g2_fill_2 FILLER_59_1814 ();
 sg13g2_decap_4 FILLER_59_1826 ();
 sg13g2_fill_1 FILLER_59_1858 ();
 sg13g2_decap_4 FILLER_59_1864 ();
 sg13g2_fill_1 FILLER_59_1880 ();
 sg13g2_fill_1 FILLER_59_1894 ();
 sg13g2_fill_1 FILLER_59_1902 ();
 sg13g2_fill_1 FILLER_59_1908 ();
 sg13g2_fill_2 FILLER_59_1917 ();
 sg13g2_fill_1 FILLER_59_1933 ();
 sg13g2_fill_2 FILLER_59_1947 ();
 sg13g2_fill_1 FILLER_59_1972 ();
 sg13g2_fill_2 FILLER_59_1986 ();
 sg13g2_fill_1 FILLER_59_1988 ();
 sg13g2_fill_1 FILLER_59_1994 ();
 sg13g2_decap_8 FILLER_59_1999 ();
 sg13g2_fill_1 FILLER_59_2015 ();
 sg13g2_fill_1 FILLER_59_2058 ();
 sg13g2_fill_1 FILLER_59_2063 ();
 sg13g2_fill_1 FILLER_59_2068 ();
 sg13g2_decap_8 FILLER_59_2074 ();
 sg13g2_decap_8 FILLER_59_2081 ();
 sg13g2_decap_8 FILLER_59_2088 ();
 sg13g2_decap_4 FILLER_59_2095 ();
 sg13g2_fill_1 FILLER_59_2099 ();
 sg13g2_fill_1 FILLER_59_2103 ();
 sg13g2_fill_1 FILLER_59_2166 ();
 sg13g2_fill_2 FILLER_59_2193 ();
 sg13g2_fill_1 FILLER_59_2195 ();
 sg13g2_fill_2 FILLER_59_2232 ();
 sg13g2_fill_1 FILLER_59_2234 ();
 sg13g2_decap_8 FILLER_59_2239 ();
 sg13g2_decap_4 FILLER_59_2246 ();
 sg13g2_fill_1 FILLER_59_2250 ();
 sg13g2_fill_1 FILLER_59_2277 ();
 sg13g2_fill_2 FILLER_59_2296 ();
 sg13g2_fill_1 FILLER_59_2303 ();
 sg13g2_fill_1 FILLER_59_2322 ();
 sg13g2_fill_2 FILLER_59_2395 ();
 sg13g2_fill_1 FILLER_59_2434 ();
 sg13g2_fill_1 FILLER_59_2536 ();
 sg13g2_fill_2 FILLER_59_2561 ();
 sg13g2_decap_8 FILLER_59_2663 ();
 sg13g2_decap_8 FILLER_60_0 ();
 sg13g2_decap_4 FILLER_60_7 ();
 sg13g2_decap_4 FILLER_60_15 ();
 sg13g2_fill_2 FILLER_60_19 ();
 sg13g2_decap_8 FILLER_60_26 ();
 sg13g2_decap_8 FILLER_60_33 ();
 sg13g2_fill_1 FILLER_60_40 ();
 sg13g2_fill_2 FILLER_60_53 ();
 sg13g2_fill_2 FILLER_60_86 ();
 sg13g2_decap_4 FILLER_60_93 ();
 sg13g2_fill_1 FILLER_60_106 ();
 sg13g2_decap_4 FILLER_60_117 ();
 sg13g2_fill_2 FILLER_60_121 ();
 sg13g2_fill_2 FILLER_60_127 ();
 sg13g2_decap_8 FILLER_60_139 ();
 sg13g2_decap_4 FILLER_60_146 ();
 sg13g2_fill_1 FILLER_60_150 ();
 sg13g2_decap_8 FILLER_60_160 ();
 sg13g2_fill_2 FILLER_60_167 ();
 sg13g2_fill_1 FILLER_60_177 ();
 sg13g2_fill_2 FILLER_60_212 ();
 sg13g2_fill_2 FILLER_60_224 ();
 sg13g2_fill_1 FILLER_60_226 ();
 sg13g2_decap_8 FILLER_60_272 ();
 sg13g2_decap_8 FILLER_60_279 ();
 sg13g2_fill_1 FILLER_60_286 ();
 sg13g2_decap_8 FILLER_60_292 ();
 sg13g2_decap_4 FILLER_60_299 ();
 sg13g2_fill_1 FILLER_60_303 ();
 sg13g2_decap_4 FILLER_60_313 ();
 sg13g2_fill_1 FILLER_60_317 ();
 sg13g2_decap_4 FILLER_60_330 ();
 sg13g2_fill_1 FILLER_60_334 ();
 sg13g2_fill_1 FILLER_60_340 ();
 sg13g2_fill_1 FILLER_60_344 ();
 sg13g2_fill_1 FILLER_60_363 ();
 sg13g2_decap_8 FILLER_60_438 ();
 sg13g2_decap_8 FILLER_60_445 ();
 sg13g2_decap_8 FILLER_60_452 ();
 sg13g2_fill_2 FILLER_60_459 ();
 sg13g2_fill_1 FILLER_60_461 ();
 sg13g2_fill_2 FILLER_60_492 ();
 sg13g2_fill_1 FILLER_60_494 ();
 sg13g2_fill_1 FILLER_60_499 ();
 sg13g2_decap_4 FILLER_60_505 ();
 sg13g2_fill_2 FILLER_60_509 ();
 sg13g2_decap_4 FILLER_60_515 ();
 sg13g2_fill_1 FILLER_60_519 ();
 sg13g2_fill_2 FILLER_60_535 ();
 sg13g2_fill_1 FILLER_60_537 ();
 sg13g2_fill_1 FILLER_60_574 ();
 sg13g2_fill_1 FILLER_60_579 ();
 sg13g2_fill_1 FILLER_60_583 ();
 sg13g2_decap_8 FILLER_60_610 ();
 sg13g2_fill_2 FILLER_60_617 ();
 sg13g2_fill_1 FILLER_60_619 ();
 sg13g2_fill_2 FILLER_60_628 ();
 sg13g2_fill_1 FILLER_60_630 ();
 sg13g2_fill_2 FILLER_60_636 ();
 sg13g2_fill_1 FILLER_60_638 ();
 sg13g2_decap_4 FILLER_60_651 ();
 sg13g2_fill_1 FILLER_60_655 ();
 sg13g2_fill_2 FILLER_60_710 ();
 sg13g2_fill_2 FILLER_60_781 ();
 sg13g2_fill_1 FILLER_60_790 ();
 sg13g2_fill_2 FILLER_60_794 ();
 sg13g2_fill_2 FILLER_60_805 ();
 sg13g2_fill_1 FILLER_60_815 ();
 sg13g2_fill_1 FILLER_60_875 ();
 sg13g2_fill_2 FILLER_60_884 ();
 sg13g2_fill_2 FILLER_60_911 ();
 sg13g2_decap_4 FILLER_60_922 ();
 sg13g2_fill_2 FILLER_60_926 ();
 sg13g2_fill_2 FILLER_60_938 ();
 sg13g2_decap_4 FILLER_60_946 ();
 sg13g2_fill_2 FILLER_60_958 ();
 sg13g2_fill_1 FILLER_60_970 ();
 sg13g2_fill_1 FILLER_60_981 ();
 sg13g2_fill_2 FILLER_60_987 ();
 sg13g2_decap_8 FILLER_60_1076 ();
 sg13g2_fill_1 FILLER_60_1083 ();
 sg13g2_fill_1 FILLER_60_1093 ();
 sg13g2_fill_1 FILLER_60_1138 ();
 sg13g2_decap_8 FILLER_60_1157 ();
 sg13g2_fill_1 FILLER_60_1164 ();
 sg13g2_decap_4 FILLER_60_1169 ();
 sg13g2_fill_1 FILLER_60_1199 ();
 sg13g2_fill_1 FILLER_60_1242 ();
 sg13g2_decap_8 FILLER_60_1248 ();
 sg13g2_decap_4 FILLER_60_1255 ();
 sg13g2_decap_8 FILLER_60_1264 ();
 sg13g2_decap_8 FILLER_60_1271 ();
 sg13g2_fill_1 FILLER_60_1278 ();
 sg13g2_decap_8 FILLER_60_1283 ();
 sg13g2_decap_4 FILLER_60_1290 ();
 sg13g2_decap_8 FILLER_60_1300 ();
 sg13g2_decap_4 FILLER_60_1307 ();
 sg13g2_decap_4 FILLER_60_1315 ();
 sg13g2_fill_1 FILLER_60_1319 ();
 sg13g2_fill_2 FILLER_60_1326 ();
 sg13g2_fill_2 FILLER_60_1333 ();
 sg13g2_decap_4 FILLER_60_1340 ();
 sg13g2_fill_1 FILLER_60_1344 ();
 sg13g2_decap_8 FILLER_60_1360 ();
 sg13g2_fill_2 FILLER_60_1378 ();
 sg13g2_fill_1 FILLER_60_1410 ();
 sg13g2_decap_8 FILLER_60_1424 ();
 sg13g2_decap_8 FILLER_60_1431 ();
 sg13g2_decap_4 FILLER_60_1438 ();
 sg13g2_fill_2 FILLER_60_1442 ();
 sg13g2_fill_1 FILLER_60_1455 ();
 sg13g2_fill_1 FILLER_60_1470 ();
 sg13g2_decap_4 FILLER_60_1560 ();
 sg13g2_decap_8 FILLER_60_1590 ();
 sg13g2_fill_2 FILLER_60_1619 ();
 sg13g2_decap_4 FILLER_60_1647 ();
 sg13g2_fill_1 FILLER_60_1651 ();
 sg13g2_fill_1 FILLER_60_1665 ();
 sg13g2_decap_8 FILLER_60_1670 ();
 sg13g2_decap_8 FILLER_60_1677 ();
 sg13g2_decap_4 FILLER_60_1684 ();
 sg13g2_fill_1 FILLER_60_1693 ();
 sg13g2_fill_2 FILLER_60_1699 ();
 sg13g2_fill_1 FILLER_60_1701 ();
 sg13g2_fill_2 FILLER_60_1710 ();
 sg13g2_decap_8 FILLER_60_1716 ();
 sg13g2_decap_4 FILLER_60_1723 ();
 sg13g2_decap_4 FILLER_60_1734 ();
 sg13g2_decap_4 FILLER_60_1747 ();
 sg13g2_fill_1 FILLER_60_1751 ();
 sg13g2_fill_1 FILLER_60_1791 ();
 sg13g2_fill_2 FILLER_60_1811 ();
 sg13g2_decap_4 FILLER_60_1820 ();
 sg13g2_fill_1 FILLER_60_1824 ();
 sg13g2_fill_2 FILLER_60_1829 ();
 sg13g2_fill_1 FILLER_60_1835 ();
 sg13g2_fill_2 FILLER_60_1878 ();
 sg13g2_fill_1 FILLER_60_1903 ();
 sg13g2_fill_2 FILLER_60_1917 ();
 sg13g2_fill_1 FILLER_60_1919 ();
 sg13g2_fill_2 FILLER_60_1943 ();
 sg13g2_decap_4 FILLER_60_1949 ();
 sg13g2_fill_1 FILLER_60_1958 ();
 sg13g2_decap_8 FILLER_60_1972 ();
 sg13g2_fill_2 FILLER_60_2003 ();
 sg13g2_fill_1 FILLER_60_2005 ();
 sg13g2_fill_1 FILLER_60_2016 ();
 sg13g2_fill_2 FILLER_60_2060 ();
 sg13g2_fill_1 FILLER_60_2062 ();
 sg13g2_fill_2 FILLER_60_2098 ();
 sg13g2_decap_4 FILLER_60_2110 ();
 sg13g2_fill_1 FILLER_60_2114 ();
 sg13g2_decap_4 FILLER_60_2120 ();
 sg13g2_fill_2 FILLER_60_2153 ();
 sg13g2_decap_8 FILLER_60_2181 ();
 sg13g2_fill_1 FILLER_60_2214 ();
 sg13g2_fill_2 FILLER_60_2219 ();
 sg13g2_fill_2 FILLER_60_2260 ();
 sg13g2_decap_8 FILLER_60_2293 ();
 sg13g2_decap_8 FILLER_60_2300 ();
 sg13g2_decap_8 FILLER_60_2307 ();
 sg13g2_decap_4 FILLER_60_2314 ();
 sg13g2_fill_1 FILLER_60_2318 ();
 sg13g2_fill_1 FILLER_60_2341 ();
 sg13g2_fill_2 FILLER_60_2390 ();
 sg13g2_fill_2 FILLER_60_2398 ();
 sg13g2_fill_1 FILLER_60_2426 ();
 sg13g2_fill_1 FILLER_60_2439 ();
 sg13g2_decap_4 FILLER_60_2457 ();
 sg13g2_fill_2 FILLER_60_2461 ();
 sg13g2_decap_4 FILLER_60_2467 ();
 sg13g2_fill_2 FILLER_60_2512 ();
 sg13g2_fill_1 FILLER_60_2514 ();
 sg13g2_fill_1 FILLER_60_2531 ();
 sg13g2_fill_2 FILLER_60_2537 ();
 sg13g2_decap_4 FILLER_60_2553 ();
 sg13g2_fill_2 FILLER_60_2557 ();
 sg13g2_decap_8 FILLER_60_2565 ();
 sg13g2_decap_8 FILLER_60_2572 ();
 sg13g2_fill_1 FILLER_60_2579 ();
 sg13g2_decap_8 FILLER_60_2584 ();
 sg13g2_decap_8 FILLER_60_2591 ();
 sg13g2_decap_8 FILLER_60_2598 ();
 sg13g2_fill_2 FILLER_60_2605 ();
 sg13g2_fill_2 FILLER_60_2661 ();
 sg13g2_fill_2 FILLER_60_2667 ();
 sg13g2_fill_1 FILLER_60_2669 ();
 sg13g2_decap_8 FILLER_61_0 ();
 sg13g2_decap_8 FILLER_61_7 ();
 sg13g2_fill_1 FILLER_61_14 ();
 sg13g2_fill_1 FILLER_61_45 ();
 sg13g2_fill_1 FILLER_61_59 ();
 sg13g2_fill_2 FILLER_61_67 ();
 sg13g2_fill_1 FILLER_61_73 ();
 sg13g2_fill_1 FILLER_61_105 ();
 sg13g2_decap_4 FILLER_61_137 ();
 sg13g2_fill_1 FILLER_61_141 ();
 sg13g2_fill_2 FILLER_61_148 ();
 sg13g2_decap_8 FILLER_61_160 ();
 sg13g2_decap_4 FILLER_61_167 ();
 sg13g2_fill_1 FILLER_61_171 ();
 sg13g2_fill_1 FILLER_61_185 ();
 sg13g2_decap_4 FILLER_61_212 ();
 sg13g2_decap_4 FILLER_61_221 ();
 sg13g2_fill_1 FILLER_61_239 ();
 sg13g2_fill_2 FILLER_61_281 ();
 sg13g2_decap_8 FILLER_61_289 ();
 sg13g2_decap_8 FILLER_61_296 ();
 sg13g2_fill_2 FILLER_61_303 ();
 sg13g2_fill_1 FILLER_61_309 ();
 sg13g2_decap_4 FILLER_61_314 ();
 sg13g2_fill_2 FILLER_61_327 ();
 sg13g2_fill_2 FILLER_61_334 ();
 sg13g2_fill_2 FILLER_61_342 ();
 sg13g2_fill_2 FILLER_61_357 ();
 sg13g2_fill_1 FILLER_61_359 ();
 sg13g2_fill_1 FILLER_61_369 ();
 sg13g2_fill_1 FILLER_61_396 ();
 sg13g2_fill_1 FILLER_61_437 ();
 sg13g2_fill_2 FILLER_61_468 ();
 sg13g2_fill_1 FILLER_61_470 ();
 sg13g2_decap_4 FILLER_61_481 ();
 sg13g2_fill_2 FILLER_61_485 ();
 sg13g2_fill_1 FILLER_61_495 ();
 sg13g2_decap_8 FILLER_61_526 ();
 sg13g2_fill_2 FILLER_61_533 ();
 sg13g2_decap_4 FILLER_61_545 ();
 sg13g2_fill_2 FILLER_61_554 ();
 sg13g2_decap_4 FILLER_61_586 ();
 sg13g2_decap_8 FILLER_61_595 ();
 sg13g2_decap_4 FILLER_61_602 ();
 sg13g2_decap_4 FILLER_61_609 ();
 sg13g2_fill_2 FILLER_61_613 ();
 sg13g2_decap_8 FILLER_61_629 ();
 sg13g2_decap_4 FILLER_61_636 ();
 sg13g2_fill_2 FILLER_61_648 ();
 sg13g2_fill_1 FILLER_61_650 ();
 sg13g2_fill_1 FILLER_61_656 ();
 sg13g2_fill_1 FILLER_61_685 ();
 sg13g2_fill_2 FILLER_61_703 ();
 sg13g2_fill_2 FILLER_61_714 ();
 sg13g2_fill_1 FILLER_61_733 ();
 sg13g2_fill_2 FILLER_61_760 ();
 sg13g2_fill_2 FILLER_61_769 ();
 sg13g2_fill_1 FILLER_61_786 ();
 sg13g2_fill_2 FILLER_61_827 ();
 sg13g2_fill_2 FILLER_61_855 ();
 sg13g2_fill_1 FILLER_61_866 ();
 sg13g2_decap_4 FILLER_61_923 ();
 sg13g2_fill_1 FILLER_61_927 ();
 sg13g2_fill_2 FILLER_61_936 ();
 sg13g2_fill_2 FILLER_61_999 ();
 sg13g2_fill_1 FILLER_61_1005 ();
 sg13g2_fill_1 FILLER_61_1012 ();
 sg13g2_decap_4 FILLER_61_1035 ();
 sg13g2_decap_8 FILLER_61_1069 ();
 sg13g2_fill_2 FILLER_61_1076 ();
 sg13g2_fill_1 FILLER_61_1088 ();
 sg13g2_fill_2 FILLER_61_1129 ();
 sg13g2_decap_8 FILLER_61_1157 ();
 sg13g2_decap_8 FILLER_61_1164 ();
 sg13g2_decap_4 FILLER_61_1171 ();
 sg13g2_decap_8 FILLER_61_1183 ();
 sg13g2_fill_2 FILLER_61_1190 ();
 sg13g2_fill_2 FILLER_61_1217 ();
 sg13g2_decap_4 FILLER_61_1252 ();
 sg13g2_fill_2 FILLER_61_1256 ();
 sg13g2_decap_4 FILLER_61_1263 ();
 sg13g2_fill_1 FILLER_61_1267 ();
 sg13g2_fill_1 FILLER_61_1273 ();
 sg13g2_decap_8 FILLER_61_1285 ();
 sg13g2_decap_4 FILLER_61_1332 ();
 sg13g2_fill_1 FILLER_61_1343 ();
 sg13g2_decap_4 FILLER_61_1349 ();
 sg13g2_fill_1 FILLER_61_1353 ();
 sg13g2_fill_1 FILLER_61_1359 ();
 sg13g2_fill_1 FILLER_61_1366 ();
 sg13g2_fill_2 FILLER_61_1372 ();
 sg13g2_fill_1 FILLER_61_1374 ();
 sg13g2_fill_2 FILLER_61_1388 ();
 sg13g2_decap_4 FILLER_61_1400 ();
 sg13g2_fill_2 FILLER_61_1415 ();
 sg13g2_decap_8 FILLER_61_1423 ();
 sg13g2_decap_8 FILLER_61_1430 ();
 sg13g2_decap_8 FILLER_61_1437 ();
 sg13g2_decap_8 FILLER_61_1444 ();
 sg13g2_fill_1 FILLER_61_1451 ();
 sg13g2_fill_2 FILLER_61_1455 ();
 sg13g2_fill_1 FILLER_61_1465 ();
 sg13g2_fill_1 FILLER_61_1474 ();
 sg13g2_fill_2 FILLER_61_1491 ();
 sg13g2_decap_8 FILLER_61_1506 ();
 sg13g2_decap_4 FILLER_61_1513 ();
 sg13g2_fill_1 FILLER_61_1517 ();
 sg13g2_fill_2 FILLER_61_1522 ();
 sg13g2_fill_1 FILLER_61_1524 ();
 sg13g2_decap_8 FILLER_61_1534 ();
 sg13g2_fill_2 FILLER_61_1541 ();
 sg13g2_fill_1 FILLER_61_1577 ();
 sg13g2_decap_4 FILLER_61_1582 ();
 sg13g2_decap_8 FILLER_61_1590 ();
 sg13g2_fill_2 FILLER_61_1597 ();
 sg13g2_fill_1 FILLER_61_1599 ();
 sg13g2_decap_8 FILLER_61_1604 ();
 sg13g2_fill_2 FILLER_61_1611 ();
 sg13g2_fill_1 FILLER_61_1613 ();
 sg13g2_fill_2 FILLER_61_1622 ();
 sg13g2_fill_2 FILLER_61_1628 ();
 sg13g2_fill_1 FILLER_61_1634 ();
 sg13g2_decap_4 FILLER_61_1655 ();
 sg13g2_decap_8 FILLER_61_1685 ();
 sg13g2_fill_2 FILLER_61_1692 ();
 sg13g2_decap_8 FILLER_61_1723 ();
 sg13g2_fill_1 FILLER_61_1730 ();
 sg13g2_fill_2 FILLER_61_1775 ();
 sg13g2_fill_1 FILLER_61_1782 ();
 sg13g2_fill_2 FILLER_61_1794 ();
 sg13g2_decap_8 FILLER_61_1805 ();
 sg13g2_fill_1 FILLER_61_1812 ();
 sg13g2_decap_8 FILLER_61_1817 ();
 sg13g2_decap_8 FILLER_61_1824 ();
 sg13g2_fill_2 FILLER_61_1831 ();
 sg13g2_decap_8 FILLER_61_1838 ();
 sg13g2_fill_2 FILLER_61_1845 ();
 sg13g2_fill_1 FILLER_61_1847 ();
 sg13g2_fill_2 FILLER_61_1856 ();
 sg13g2_fill_1 FILLER_61_1858 ();
 sg13g2_fill_1 FILLER_61_1869 ();
 sg13g2_fill_2 FILLER_61_1874 ();
 sg13g2_fill_1 FILLER_61_1881 ();
 sg13g2_fill_2 FILLER_61_1886 ();
 sg13g2_fill_1 FILLER_61_1947 ();
 sg13g2_fill_1 FILLER_61_1968 ();
 sg13g2_decap_4 FILLER_61_1974 ();
 sg13g2_fill_1 FILLER_61_1978 ();
 sg13g2_fill_2 FILLER_61_1984 ();
 sg13g2_fill_1 FILLER_61_1991 ();
 sg13g2_fill_2 FILLER_61_2047 ();
 sg13g2_fill_2 FILLER_61_2053 ();
 sg13g2_fill_2 FILLER_61_2072 ();
 sg13g2_fill_1 FILLER_61_2103 ();
 sg13g2_decap_8 FILLER_61_2107 ();
 sg13g2_decap_4 FILLER_61_2114 ();
 sg13g2_fill_2 FILLER_61_2122 ();
 sg13g2_fill_2 FILLER_61_2238 ();
 sg13g2_decap_4 FILLER_61_2244 ();
 sg13g2_fill_1 FILLER_61_2248 ();
 sg13g2_fill_1 FILLER_61_2273 ();
 sg13g2_fill_1 FILLER_61_2279 ();
 sg13g2_fill_1 FILLER_61_2288 ();
 sg13g2_fill_1 FILLER_61_2294 ();
 sg13g2_fill_2 FILLER_61_2303 ();
 sg13g2_fill_1 FILLER_61_2349 ();
 sg13g2_fill_1 FILLER_61_2355 ();
 sg13g2_fill_1 FILLER_61_2366 ();
 sg13g2_fill_1 FILLER_61_2403 ();
 sg13g2_fill_1 FILLER_61_2409 ();
 sg13g2_decap_4 FILLER_61_2414 ();
 sg13g2_fill_1 FILLER_61_2418 ();
 sg13g2_fill_1 FILLER_61_2423 ();
 sg13g2_fill_1 FILLER_61_2428 ();
 sg13g2_fill_1 FILLER_61_2493 ();
 sg13g2_decap_8 FILLER_61_2498 ();
 sg13g2_decap_8 FILLER_61_2505 ();
 sg13g2_decap_8 FILLER_61_2512 ();
 sg13g2_decap_8 FILLER_61_2523 ();
 sg13g2_fill_2 FILLER_61_2530 ();
 sg13g2_fill_1 FILLER_61_2532 ();
 sg13g2_decap_8 FILLER_61_2539 ();
 sg13g2_decap_4 FILLER_61_2546 ();
 sg13g2_fill_2 FILLER_61_2550 ();
 sg13g2_decap_8 FILLER_61_2566 ();
 sg13g2_fill_2 FILLER_61_2573 ();
 sg13g2_fill_1 FILLER_61_2575 ();
 sg13g2_fill_2 FILLER_61_2581 ();
 sg13g2_fill_2 FILLER_61_2629 ();
 sg13g2_fill_1 FILLER_61_2631 ();
 sg13g2_fill_2 FILLER_61_2668 ();
 sg13g2_fill_2 FILLER_62_0 ();
 sg13g2_fill_1 FILLER_62_28 ();
 sg13g2_decap_8 FILLER_62_47 ();
 sg13g2_fill_2 FILLER_62_54 ();
 sg13g2_decap_8 FILLER_62_67 ();
 sg13g2_decap_4 FILLER_62_74 ();
 sg13g2_fill_2 FILLER_62_78 ();
 sg13g2_decap_4 FILLER_62_106 ();
 sg13g2_fill_1 FILLER_62_118 ();
 sg13g2_decap_8 FILLER_62_133 ();
 sg13g2_decap_4 FILLER_62_140 ();
 sg13g2_fill_1 FILLER_62_144 ();
 sg13g2_fill_1 FILLER_62_180 ();
 sg13g2_fill_2 FILLER_62_189 ();
 sg13g2_fill_1 FILLER_62_201 ();
 sg13g2_fill_1 FILLER_62_223 ();
 sg13g2_fill_1 FILLER_62_229 ();
 sg13g2_fill_1 FILLER_62_235 ();
 sg13g2_fill_1 FILLER_62_241 ();
 sg13g2_fill_1 FILLER_62_255 ();
 sg13g2_fill_2 FILLER_62_266 ();
 sg13g2_fill_1 FILLER_62_310 ();
 sg13g2_fill_1 FILLER_62_402 ();
 sg13g2_fill_2 FILLER_62_418 ();
 sg13g2_fill_1 FILLER_62_432 ();
 sg13g2_decap_4 FILLER_62_481 ();
 sg13g2_decap_8 FILLER_62_528 ();
 sg13g2_decap_4 FILLER_62_535 ();
 sg13g2_fill_1 FILLER_62_549 ();
 sg13g2_decap_8 FILLER_62_565 ();
 sg13g2_decap_8 FILLER_62_576 ();
 sg13g2_fill_2 FILLER_62_583 ();
 sg13g2_fill_1 FILLER_62_585 ();
 sg13g2_decap_8 FILLER_62_594 ();
 sg13g2_fill_2 FILLER_62_601 ();
 sg13g2_fill_2 FILLER_62_649 ();
 sg13g2_fill_2 FILLER_62_658 ();
 sg13g2_fill_1 FILLER_62_676 ();
 sg13g2_fill_2 FILLER_62_738 ();
 sg13g2_fill_2 FILLER_62_759 ();
 sg13g2_fill_1 FILLER_62_786 ();
 sg13g2_fill_2 FILLER_62_812 ();
 sg13g2_fill_1 FILLER_62_829 ();
 sg13g2_fill_2 FILLER_62_892 ();
 sg13g2_fill_2 FILLER_62_942 ();
 sg13g2_fill_1 FILLER_62_944 ();
 sg13g2_fill_1 FILLER_62_948 ();
 sg13g2_fill_1 FILLER_62_957 ();
 sg13g2_fill_1 FILLER_62_962 ();
 sg13g2_fill_1 FILLER_62_968 ();
 sg13g2_fill_1 FILLER_62_973 ();
 sg13g2_fill_2 FILLER_62_978 ();
 sg13g2_fill_2 FILLER_62_991 ();
 sg13g2_fill_2 FILLER_62_1001 ();
 sg13g2_fill_2 FILLER_62_1006 ();
 sg13g2_decap_8 FILLER_62_1040 ();
 sg13g2_decap_4 FILLER_62_1047 ();
 sg13g2_fill_1 FILLER_62_1055 ();
 sg13g2_fill_2 FILLER_62_1089 ();
 sg13g2_fill_1 FILLER_62_1091 ();
 sg13g2_fill_2 FILLER_62_1133 ();
 sg13g2_fill_1 FILLER_62_1148 ();
 sg13g2_decap_8 FILLER_62_1157 ();
 sg13g2_decap_8 FILLER_62_1164 ();
 sg13g2_decap_4 FILLER_62_1171 ();
 sg13g2_fill_2 FILLER_62_1175 ();
 sg13g2_decap_8 FILLER_62_1181 ();
 sg13g2_fill_1 FILLER_62_1188 ();
 sg13g2_fill_1 FILLER_62_1217 ();
 sg13g2_fill_2 FILLER_62_1226 ();
 sg13g2_fill_1 FILLER_62_1249 ();
 sg13g2_fill_1 FILLER_62_1261 ();
 sg13g2_fill_1 FILLER_62_1273 ();
 sg13g2_fill_1 FILLER_62_1280 ();
 sg13g2_decap_4 FILLER_62_1286 ();
 sg13g2_decap_8 FILLER_62_1295 ();
 sg13g2_fill_2 FILLER_62_1302 ();
 sg13g2_fill_1 FILLER_62_1304 ();
 sg13g2_fill_1 FILLER_62_1309 ();
 sg13g2_fill_1 FILLER_62_1321 ();
 sg13g2_decap_8 FILLER_62_1349 ();
 sg13g2_decap_4 FILLER_62_1383 ();
 sg13g2_decap_4 FILLER_62_1410 ();
 sg13g2_decap_8 FILLER_62_1454 ();
 sg13g2_decap_8 FILLER_62_1461 ();
 sg13g2_decap_4 FILLER_62_1484 ();
 sg13g2_fill_2 FILLER_62_1497 ();
 sg13g2_fill_1 FILLER_62_1499 ();
 sg13g2_decap_8 FILLER_62_1513 ();
 sg13g2_decap_8 FILLER_62_1520 ();
 sg13g2_decap_8 FILLER_62_1527 ();
 sg13g2_fill_1 FILLER_62_1534 ();
 sg13g2_fill_2 FILLER_62_1544 ();
 sg13g2_fill_1 FILLER_62_1549 ();
 sg13g2_fill_2 FILLER_62_1584 ();
 sg13g2_fill_1 FILLER_62_1586 ();
 sg13g2_fill_2 FILLER_62_1592 ();
 sg13g2_decap_4 FILLER_62_1599 ();
 sg13g2_fill_1 FILLER_62_1603 ();
 sg13g2_fill_1 FILLER_62_1609 ();
 sg13g2_decap_8 FILLER_62_1629 ();
 sg13g2_decap_4 FILLER_62_1636 ();
 sg13g2_decap_4 FILLER_62_1644 ();
 sg13g2_fill_1 FILLER_62_1648 ();
 sg13g2_decap_8 FILLER_62_1666 ();
 sg13g2_decap_8 FILLER_62_1673 ();
 sg13g2_decap_8 FILLER_62_1680 ();
 sg13g2_decap_4 FILLER_62_1687 ();
 sg13g2_fill_1 FILLER_62_1691 ();
 sg13g2_decap_4 FILLER_62_1697 ();
 sg13g2_decap_8 FILLER_62_1705 ();
 sg13g2_decap_8 FILLER_62_1712 ();
 sg13g2_decap_8 FILLER_62_1723 ();
 sg13g2_decap_4 FILLER_62_1730 ();
 sg13g2_fill_1 FILLER_62_1734 ();
 sg13g2_decap_4 FILLER_62_1760 ();
 sg13g2_decap_8 FILLER_62_1771 ();
 sg13g2_decap_8 FILLER_62_1782 ();
 sg13g2_fill_1 FILLER_62_1789 ();
 sg13g2_decap_4 FILLER_62_1823 ();
 sg13g2_fill_2 FILLER_62_1831 ();
 sg13g2_fill_1 FILLER_62_1833 ();
 sg13g2_decap_8 FILLER_62_1838 ();
 sg13g2_decap_8 FILLER_62_1845 ();
 sg13g2_decap_8 FILLER_62_1852 ();
 sg13g2_fill_2 FILLER_62_1859 ();
 sg13g2_fill_2 FILLER_62_1893 ();
 sg13g2_fill_1 FILLER_62_1907 ();
 sg13g2_fill_2 FILLER_62_1922 ();
 sg13g2_fill_1 FILLER_62_1924 ();
 sg13g2_fill_2 FILLER_62_1933 ();
 sg13g2_fill_2 FILLER_62_1939 ();
 sg13g2_fill_1 FILLER_62_1946 ();
 sg13g2_fill_1 FILLER_62_1952 ();
 sg13g2_fill_2 FILLER_62_1961 ();
 sg13g2_fill_2 FILLER_62_1967 ();
 sg13g2_fill_1 FILLER_62_1969 ();
 sg13g2_fill_1 FILLER_62_1980 ();
 sg13g2_decap_8 FILLER_62_1987 ();
 sg13g2_fill_2 FILLER_62_2003 ();
 sg13g2_fill_1 FILLER_62_2005 ();
 sg13g2_fill_2 FILLER_62_2021 ();
 sg13g2_decap_4 FILLER_62_2033 ();
 sg13g2_fill_1 FILLER_62_2037 ();
 sg13g2_decap_8 FILLER_62_2042 ();
 sg13g2_decap_4 FILLER_62_2049 ();
 sg13g2_decap_8 FILLER_62_2057 ();
 sg13g2_decap_4 FILLER_62_2100 ();
 sg13g2_decap_8 FILLER_62_2107 ();
 sg13g2_decap_8 FILLER_62_2114 ();
 sg13g2_fill_2 FILLER_62_2121 ();
 sg13g2_fill_1 FILLER_62_2123 ();
 sg13g2_decap_8 FILLER_62_2127 ();
 sg13g2_fill_2 FILLER_62_2134 ();
 sg13g2_decap_4 FILLER_62_2140 ();
 sg13g2_fill_1 FILLER_62_2151 ();
 sg13g2_fill_2 FILLER_62_2200 ();
 sg13g2_fill_2 FILLER_62_2215 ();
 sg13g2_fill_1 FILLER_62_2230 ();
 sg13g2_fill_1 FILLER_62_2318 ();
 sg13g2_decap_8 FILLER_62_2369 ();
 sg13g2_decap_8 FILLER_62_2376 ();
 sg13g2_decap_4 FILLER_62_2383 ();
 sg13g2_fill_1 FILLER_62_2387 ();
 sg13g2_fill_2 FILLER_62_2412 ();
 sg13g2_fill_1 FILLER_62_2414 ();
 sg13g2_fill_2 FILLER_62_2446 ();
 sg13g2_fill_1 FILLER_62_2448 ();
 sg13g2_fill_2 FILLER_62_2459 ();
 sg13g2_fill_1 FILLER_62_2461 ();
 sg13g2_fill_2 FILLER_62_2467 ();
 sg13g2_fill_2 FILLER_62_2473 ();
 sg13g2_fill_2 FILLER_62_2515 ();
 sg13g2_decap_4 FILLER_62_2522 ();
 sg13g2_fill_2 FILLER_62_2526 ();
 sg13g2_fill_1 FILLER_62_2542 ();
 sg13g2_decap_4 FILLER_62_2547 ();
 sg13g2_fill_1 FILLER_62_2587 ();
 sg13g2_fill_2 FILLER_62_2642 ();
 sg13g2_decap_8 FILLER_62_2648 ();
 sg13g2_decap_8 FILLER_62_2655 ();
 sg13g2_decap_8 FILLER_62_2662 ();
 sg13g2_fill_1 FILLER_62_2669 ();
 sg13g2_decap_4 FILLER_63_0 ();
 sg13g2_fill_2 FILLER_63_4 ();
 sg13g2_fill_2 FILLER_63_49 ();
 sg13g2_fill_1 FILLER_63_51 ();
 sg13g2_fill_2 FILLER_63_75 ();
 sg13g2_fill_1 FILLER_63_77 ();
 sg13g2_decap_4 FILLER_63_82 ();
 sg13g2_fill_2 FILLER_63_86 ();
 sg13g2_fill_2 FILLER_63_137 ();
 sg13g2_decap_4 FILLER_63_165 ();
 sg13g2_fill_1 FILLER_63_169 ();
 sg13g2_decap_4 FILLER_63_199 ();
 sg13g2_fill_1 FILLER_63_229 ();
 sg13g2_fill_1 FILLER_63_235 ();
 sg13g2_fill_1 FILLER_63_276 ();
 sg13g2_fill_1 FILLER_63_287 ();
 sg13g2_fill_2 FILLER_63_296 ();
 sg13g2_fill_1 FILLER_63_310 ();
 sg13g2_fill_2 FILLER_63_316 ();
 sg13g2_fill_1 FILLER_63_318 ();
 sg13g2_fill_1 FILLER_63_340 ();
 sg13g2_fill_1 FILLER_63_350 ();
 sg13g2_fill_1 FILLER_63_370 ();
 sg13g2_fill_2 FILLER_63_376 ();
 sg13g2_fill_1 FILLER_63_504 ();
 sg13g2_fill_1 FILLER_63_510 ();
 sg13g2_decap_4 FILLER_63_549 ();
 sg13g2_fill_1 FILLER_63_553 ();
 sg13g2_decap_4 FILLER_63_558 ();
 sg13g2_fill_2 FILLER_63_562 ();
 sg13g2_decap_8 FILLER_63_601 ();
 sg13g2_decap_4 FILLER_63_608 ();
 sg13g2_fill_2 FILLER_63_612 ();
 sg13g2_fill_2 FILLER_63_629 ();
 sg13g2_fill_1 FILLER_63_649 ();
 sg13g2_fill_1 FILLER_63_658 ();
 sg13g2_fill_1 FILLER_63_675 ();
 sg13g2_fill_1 FILLER_63_730 ();
 sg13g2_fill_2 FILLER_63_749 ();
 sg13g2_fill_1 FILLER_63_769 ();
 sg13g2_fill_1 FILLER_63_787 ();
 sg13g2_fill_1 FILLER_63_802 ();
 sg13g2_fill_2 FILLER_63_817 ();
 sg13g2_fill_2 FILLER_63_857 ();
 sg13g2_fill_2 FILLER_63_877 ();
 sg13g2_fill_1 FILLER_63_886 ();
 sg13g2_fill_2 FILLER_63_896 ();
 sg13g2_fill_1 FILLER_63_920 ();
 sg13g2_fill_1 FILLER_63_931 ();
 sg13g2_fill_2 FILLER_63_936 ();
 sg13g2_fill_1 FILLER_63_938 ();
 sg13g2_fill_1 FILLER_63_944 ();
 sg13g2_decap_8 FILLER_63_961 ();
 sg13g2_fill_2 FILLER_63_968 ();
 sg13g2_fill_1 FILLER_63_970 ();
 sg13g2_decap_8 FILLER_63_1036 ();
 sg13g2_fill_2 FILLER_63_1043 ();
 sg13g2_fill_1 FILLER_63_1080 ();
 sg13g2_fill_2 FILLER_63_1086 ();
 sg13g2_fill_1 FILLER_63_1088 ();
 sg13g2_fill_2 FILLER_63_1126 ();
 sg13g2_decap_8 FILLER_63_1162 ();
 sg13g2_decap_8 FILLER_63_1169 ();
 sg13g2_fill_1 FILLER_63_1181 ();
 sg13g2_decap_4 FILLER_63_1191 ();
 sg13g2_fill_1 FILLER_63_1195 ();
 sg13g2_decap_8 FILLER_63_1201 ();
 sg13g2_decap_8 FILLER_63_1232 ();
 sg13g2_fill_1 FILLER_63_1239 ();
 sg13g2_fill_2 FILLER_63_1253 ();
 sg13g2_fill_2 FILLER_63_1268 ();
 sg13g2_fill_1 FILLER_63_1283 ();
 sg13g2_fill_1 FILLER_63_1300 ();
 sg13g2_fill_1 FILLER_63_1305 ();
 sg13g2_fill_1 FILLER_63_1331 ();
 sg13g2_fill_1 FILLER_63_1337 ();
 sg13g2_fill_1 FILLER_63_1345 ();
 sg13g2_fill_2 FILLER_63_1353 ();
 sg13g2_fill_1 FILLER_63_1355 ();
 sg13g2_decap_4 FILLER_63_1360 ();
 sg13g2_fill_1 FILLER_63_1364 ();
 sg13g2_decap_4 FILLER_63_1371 ();
 sg13g2_fill_2 FILLER_63_1375 ();
 sg13g2_decap_4 FILLER_63_1396 ();
 sg13g2_fill_2 FILLER_63_1456 ();
 sg13g2_fill_1 FILLER_63_1458 ();
 sg13g2_fill_1 FILLER_63_1464 ();
 sg13g2_fill_2 FILLER_63_1476 ();
 sg13g2_decap_8 FILLER_63_1483 ();
 sg13g2_fill_2 FILLER_63_1490 ();
 sg13g2_fill_1 FILLER_63_1556 ();
 sg13g2_decap_8 FILLER_63_1575 ();
 sg13g2_fill_2 FILLER_63_1582 ();
 sg13g2_fill_1 FILLER_63_1584 ();
 sg13g2_decap_8 FILLER_63_1590 ();
 sg13g2_decap_4 FILLER_63_1597 ();
 sg13g2_fill_2 FILLER_63_1624 ();
 sg13g2_fill_1 FILLER_63_1631 ();
 sg13g2_decap_8 FILLER_63_1637 ();
 sg13g2_fill_2 FILLER_63_1644 ();
 sg13g2_fill_1 FILLER_63_1696 ();
 sg13g2_fill_1 FILLER_63_1702 ();
 sg13g2_fill_1 FILLER_63_1729 ();
 sg13g2_fill_1 FILLER_63_1740 ();
 sg13g2_decap_8 FILLER_63_1767 ();
 sg13g2_decap_8 FILLER_63_1774 ();
 sg13g2_decap_8 FILLER_63_1781 ();
 sg13g2_fill_2 FILLER_63_1788 ();
 sg13g2_decap_8 FILLER_63_1853 ();
 sg13g2_decap_8 FILLER_63_1860 ();
 sg13g2_fill_2 FILLER_63_1872 ();
 sg13g2_decap_4 FILLER_63_1879 ();
 sg13g2_fill_2 FILLER_63_1883 ();
 sg13g2_fill_2 FILLER_63_1905 ();
 sg13g2_fill_1 FILLER_63_1912 ();
 sg13g2_fill_1 FILLER_63_1925 ();
 sg13g2_fill_2 FILLER_63_1934 ();
 sg13g2_fill_2 FILLER_63_1966 ();
 sg13g2_decap_4 FILLER_63_1982 ();
 sg13g2_fill_1 FILLER_63_1986 ();
 sg13g2_fill_2 FILLER_63_1999 ();
 sg13g2_fill_1 FILLER_63_2006 ();
 sg13g2_fill_1 FILLER_63_2011 ();
 sg13g2_decap_8 FILLER_63_2017 ();
 sg13g2_fill_1 FILLER_63_2024 ();
 sg13g2_decap_8 FILLER_63_2030 ();
 sg13g2_decap_8 FILLER_63_2041 ();
 sg13g2_decap_4 FILLER_63_2048 ();
 sg13g2_decap_8 FILLER_63_2092 ();
 sg13g2_decap_4 FILLER_63_2099 ();
 sg13g2_fill_1 FILLER_63_2103 ();
 sg13g2_decap_8 FILLER_63_2108 ();
 sg13g2_decap_8 FILLER_63_2115 ();
 sg13g2_decap_8 FILLER_63_2122 ();
 sg13g2_fill_2 FILLER_63_2129 ();
 sg13g2_fill_1 FILLER_63_2131 ();
 sg13g2_decap_8 FILLER_63_2136 ();
 sg13g2_fill_1 FILLER_63_2143 ();
 sg13g2_fill_2 FILLER_63_2158 ();
 sg13g2_fill_1 FILLER_63_2160 ();
 sg13g2_decap_8 FILLER_63_2171 ();
 sg13g2_decap_8 FILLER_63_2178 ();
 sg13g2_decap_4 FILLER_63_2185 ();
 sg13g2_decap_8 FILLER_63_2238 ();
 sg13g2_decap_8 FILLER_63_2245 ();
 sg13g2_fill_2 FILLER_63_2252 ();
 sg13g2_fill_2 FILLER_63_2316 ();
 sg13g2_decap_4 FILLER_63_2381 ();
 sg13g2_fill_1 FILLER_63_2385 ();
 sg13g2_fill_1 FILLER_63_2396 ();
 sg13g2_fill_2 FILLER_63_2421 ();
 sg13g2_fill_2 FILLER_63_2427 ();
 sg13g2_fill_1 FILLER_63_2429 ();
 sg13g2_fill_2 FILLER_63_2466 ();
 sg13g2_fill_1 FILLER_63_2472 ();
 sg13g2_fill_1 FILLER_63_2539 ();
 sg13g2_fill_1 FILLER_63_2576 ();
 sg13g2_fill_1 FILLER_63_2582 ();
 sg13g2_decap_4 FILLER_63_2613 ();
 sg13g2_fill_2 FILLER_63_2642 ();
 sg13g2_fill_2 FILLER_64_0 ();
 sg13g2_decap_8 FILLER_64_33 ();
 sg13g2_fill_1 FILLER_64_40 ();
 sg13g2_fill_1 FILLER_64_51 ();
 sg13g2_fill_1 FILLER_64_62 ();
 sg13g2_fill_2 FILLER_64_89 ();
 sg13g2_fill_2 FILLER_64_117 ();
 sg13g2_fill_2 FILLER_64_123 ();
 sg13g2_fill_2 FILLER_64_143 ();
 sg13g2_fill_2 FILLER_64_155 ();
 sg13g2_fill_2 FILLER_64_175 ();
 sg13g2_fill_1 FILLER_64_220 ();
 sg13g2_fill_1 FILLER_64_294 ();
 sg13g2_fill_1 FILLER_64_325 ();
 sg13g2_fill_1 FILLER_64_375 ();
 sg13g2_fill_2 FILLER_64_383 ();
 sg13g2_fill_1 FILLER_64_385 ();
 sg13g2_fill_1 FILLER_64_395 ();
 sg13g2_fill_1 FILLER_64_418 ();
 sg13g2_fill_1 FILLER_64_439 ();
 sg13g2_fill_2 FILLER_64_457 ();
 sg13g2_fill_1 FILLER_64_469 ();
 sg13g2_decap_4 FILLER_64_503 ();
 sg13g2_fill_2 FILLER_64_515 ();
 sg13g2_fill_1 FILLER_64_517 ();
 sg13g2_decap_8 FILLER_64_552 ();
 sg13g2_decap_8 FILLER_64_559 ();
 sg13g2_decap_4 FILLER_64_566 ();
 sg13g2_fill_1 FILLER_64_574 ();
 sg13g2_fill_1 FILLER_64_580 ();
 sg13g2_fill_1 FILLER_64_607 ();
 sg13g2_fill_1 FILLER_64_626 ();
 sg13g2_fill_2 FILLER_64_633 ();
 sg13g2_fill_2 FILLER_64_651 ();
 sg13g2_fill_1 FILLER_64_667 ();
 sg13g2_fill_1 FILLER_64_701 ();
 sg13g2_fill_1 FILLER_64_728 ();
 sg13g2_fill_1 FILLER_64_755 ();
 sg13g2_fill_1 FILLER_64_766 ();
 sg13g2_fill_1 FILLER_64_826 ();
 sg13g2_fill_1 FILLER_64_838 ();
 sg13g2_fill_2 FILLER_64_880 ();
 sg13g2_fill_2 FILLER_64_887 ();
 sg13g2_fill_1 FILLER_64_903 ();
 sg13g2_fill_1 FILLER_64_924 ();
 sg13g2_fill_2 FILLER_64_930 ();
 sg13g2_decap_8 FILLER_64_936 ();
 sg13g2_fill_2 FILLER_64_943 ();
 sg13g2_decap_8 FILLER_64_948 ();
 sg13g2_decap_4 FILLER_64_955 ();
 sg13g2_fill_1 FILLER_64_959 ();
 sg13g2_fill_1 FILLER_64_977 ();
 sg13g2_fill_2 FILLER_64_1017 ();
 sg13g2_fill_2 FILLER_64_1023 ();
 sg13g2_fill_1 FILLER_64_1025 ();
 sg13g2_fill_2 FILLER_64_1029 ();
 sg13g2_decap_4 FILLER_64_1035 ();
 sg13g2_fill_1 FILLER_64_1065 ();
 sg13g2_fill_1 FILLER_64_1076 ();
 sg13g2_fill_1 FILLER_64_1116 ();
 sg13g2_fill_2 FILLER_64_1154 ();
 sg13g2_fill_1 FILLER_64_1156 ();
 sg13g2_fill_1 FILLER_64_1188 ();
 sg13g2_decap_8 FILLER_64_1193 ();
 sg13g2_fill_1 FILLER_64_1200 ();
 sg13g2_fill_2 FILLER_64_1227 ();
 sg13g2_fill_1 FILLER_64_1229 ();
 sg13g2_fill_2 FILLER_64_1238 ();
 sg13g2_fill_1 FILLER_64_1252 ();
 sg13g2_fill_1 FILLER_64_1263 ();
 sg13g2_fill_2 FILLER_64_1294 ();
 sg13g2_fill_2 FILLER_64_1318 ();
 sg13g2_fill_1 FILLER_64_1320 ();
 sg13g2_decap_8 FILLER_64_1326 ();
 sg13g2_decap_4 FILLER_64_1333 ();
 sg13g2_fill_2 FILLER_64_1337 ();
 sg13g2_decap_4 FILLER_64_1349 ();
 sg13g2_fill_1 FILLER_64_1353 ();
 sg13g2_fill_2 FILLER_64_1358 ();
 sg13g2_fill_2 FILLER_64_1371 ();
 sg13g2_fill_1 FILLER_64_1378 ();
 sg13g2_fill_2 FILLER_64_1431 ();
 sg13g2_fill_1 FILLER_64_1433 ();
 sg13g2_fill_1 FILLER_64_1438 ();
 sg13g2_decap_8 FILLER_64_1443 ();
 sg13g2_decap_4 FILLER_64_1450 ();
 sg13g2_fill_2 FILLER_64_1454 ();
 sg13g2_fill_2 FILLER_64_1479 ();
 sg13g2_decap_8 FILLER_64_1485 ();
 sg13g2_decap_8 FILLER_64_1492 ();
 sg13g2_decap_8 FILLER_64_1499 ();
 sg13g2_decap_8 FILLER_64_1506 ();
 sg13g2_fill_1 FILLER_64_1513 ();
 sg13g2_decap_4 FILLER_64_1520 ();
 sg13g2_fill_1 FILLER_64_1524 ();
 sg13g2_fill_1 FILLER_64_1541 ();
 sg13g2_fill_2 FILLER_64_1549 ();
 sg13g2_fill_2 FILLER_64_1588 ();
 sg13g2_fill_1 FILLER_64_1590 ();
 sg13g2_fill_2 FILLER_64_1604 ();
 sg13g2_fill_1 FILLER_64_1606 ();
 sg13g2_fill_1 FILLER_64_1616 ();
 sg13g2_decap_8 FILLER_64_1637 ();
 sg13g2_decap_4 FILLER_64_1644 ();
 sg13g2_fill_1 FILLER_64_1648 ();
 sg13g2_fill_1 FILLER_64_1678 ();
 sg13g2_fill_2 FILLER_64_1684 ();
 sg13g2_fill_1 FILLER_64_1686 ();
 sg13g2_decap_4 FILLER_64_1703 ();
 sg13g2_fill_2 FILLER_64_1707 ();
 sg13g2_fill_1 FILLER_64_1729 ();
 sg13g2_decap_8 FILLER_64_1738 ();
 sg13g2_decap_4 FILLER_64_1745 ();
 sg13g2_fill_1 FILLER_64_1749 ();
 sg13g2_fill_2 FILLER_64_1754 ();
 sg13g2_decap_8 FILLER_64_1765 ();
 sg13g2_fill_2 FILLER_64_1772 ();
 sg13g2_fill_1 FILLER_64_1774 ();
 sg13g2_fill_1 FILLER_64_1791 ();
 sg13g2_decap_8 FILLER_64_1797 ();
 sg13g2_decap_4 FILLER_64_1804 ();
 sg13g2_fill_2 FILLER_64_1808 ();
 sg13g2_decap_8 FILLER_64_1815 ();
 sg13g2_decap_8 FILLER_64_1822 ();
 sg13g2_fill_2 FILLER_64_1829 ();
 sg13g2_decap_8 FILLER_64_1839 ();
 sg13g2_fill_2 FILLER_64_1855 ();
 sg13g2_decap_8 FILLER_64_1862 ();
 sg13g2_decap_8 FILLER_64_1869 ();
 sg13g2_fill_2 FILLER_64_1876 ();
 sg13g2_fill_1 FILLER_64_1878 ();
 sg13g2_decap_8 FILLER_64_1884 ();
 sg13g2_decap_8 FILLER_64_1891 ();
 sg13g2_decap_8 FILLER_64_1908 ();
 sg13g2_decap_4 FILLER_64_1915 ();
 sg13g2_fill_2 FILLER_64_1919 ();
 sg13g2_fill_1 FILLER_64_1925 ();
 sg13g2_decap_4 FILLER_64_1930 ();
 sg13g2_fill_1 FILLER_64_1980 ();
 sg13g2_decap_4 FILLER_64_1985 ();
 sg13g2_fill_1 FILLER_64_1989 ();
 sg13g2_fill_1 FILLER_64_2003 ();
 sg13g2_decap_8 FILLER_64_2027 ();
 sg13g2_fill_2 FILLER_64_2034 ();
 sg13g2_decap_8 FILLER_64_2040 ();
 sg13g2_decap_4 FILLER_64_2047 ();
 sg13g2_fill_2 FILLER_64_2051 ();
 sg13g2_fill_2 FILLER_64_2067 ();
 sg13g2_decap_8 FILLER_64_2073 ();
 sg13g2_decap_4 FILLER_64_2080 ();
 sg13g2_fill_1 FILLER_64_2084 ();
 sg13g2_decap_8 FILLER_64_2121 ();
 sg13g2_decap_8 FILLER_64_2128 ();
 sg13g2_decap_4 FILLER_64_2135 ();
 sg13g2_fill_1 FILLER_64_2139 ();
 sg13g2_fill_2 FILLER_64_2151 ();
 sg13g2_fill_1 FILLER_64_2156 ();
 sg13g2_fill_1 FILLER_64_2234 ();
 sg13g2_decap_8 FILLER_64_2243 ();
 sg13g2_decap_4 FILLER_64_2250 ();
 sg13g2_fill_1 FILLER_64_2337 ();
 sg13g2_fill_1 FILLER_64_2343 ();
 sg13g2_fill_1 FILLER_64_2348 ();
 sg13g2_fill_1 FILLER_64_2391 ();
 sg13g2_fill_2 FILLER_64_2435 ();
 sg13g2_fill_1 FILLER_64_2437 ();
 sg13g2_fill_2 FILLER_64_2442 ();
 sg13g2_fill_1 FILLER_64_2444 ();
 sg13g2_fill_2 FILLER_64_2451 ();
 sg13g2_fill_1 FILLER_64_2453 ();
 sg13g2_decap_8 FILLER_64_2471 ();
 sg13g2_fill_2 FILLER_64_2478 ();
 sg13g2_decap_4 FILLER_64_2484 ();
 sg13g2_fill_2 FILLER_64_2527 ();
 sg13g2_fill_1 FILLER_64_2577 ();
 sg13g2_fill_1 FILLER_64_2654 ();
 sg13g2_decap_8 FILLER_64_2659 ();
 sg13g2_decap_4 FILLER_64_2666 ();
 sg13g2_fill_2 FILLER_65_0 ();
 sg13g2_decap_4 FILLER_65_28 ();
 sg13g2_decap_4 FILLER_65_58 ();
 sg13g2_fill_2 FILLER_65_134 ();
 sg13g2_fill_1 FILLER_65_143 ();
 sg13g2_fill_2 FILLER_65_153 ();
 sg13g2_decap_8 FILLER_65_160 ();
 sg13g2_decap_8 FILLER_65_167 ();
 sg13g2_fill_2 FILLER_65_174 ();
 sg13g2_fill_1 FILLER_65_176 ();
 sg13g2_decap_8 FILLER_65_181 ();
 sg13g2_decap_4 FILLER_65_188 ();
 sg13g2_fill_1 FILLER_65_202 ();
 sg13g2_decap_4 FILLER_65_232 ();
 sg13g2_fill_2 FILLER_65_270 ();
 sg13g2_fill_1 FILLER_65_277 ();
 sg13g2_decap_4 FILLER_65_282 ();
 sg13g2_decap_4 FILLER_65_295 ();
 sg13g2_decap_8 FILLER_65_305 ();
 sg13g2_decap_4 FILLER_65_312 ();
 sg13g2_decap_4 FILLER_65_325 ();
 sg13g2_fill_2 FILLER_65_329 ();
 sg13g2_fill_1 FILLER_65_344 ();
 sg13g2_fill_1 FILLER_65_361 ();
 sg13g2_decap_8 FILLER_65_378 ();
 sg13g2_fill_1 FILLER_65_385 ();
 sg13g2_fill_2 FILLER_65_390 ();
 sg13g2_decap_4 FILLER_65_457 ();
 sg13g2_fill_2 FILLER_65_461 ();
 sg13g2_fill_2 FILLER_65_467 ();
 sg13g2_fill_2 FILLER_65_477 ();
 sg13g2_decap_4 FILLER_65_484 ();
 sg13g2_fill_1 FILLER_65_488 ();
 sg13g2_decap_4 FILLER_65_493 ();
 sg13g2_fill_1 FILLER_65_513 ();
 sg13g2_fill_2 FILLER_65_518 ();
 sg13g2_decap_8 FILLER_65_525 ();
 sg13g2_decap_4 FILLER_65_532 ();
 sg13g2_fill_2 FILLER_65_536 ();
 sg13g2_decap_8 FILLER_65_541 ();
 sg13g2_fill_1 FILLER_65_548 ();
 sg13g2_fill_2 FILLER_65_554 ();
 sg13g2_fill_2 FILLER_65_612 ();
 sg13g2_decap_8 FILLER_65_654 ();
 sg13g2_fill_2 FILLER_65_661 ();
 sg13g2_fill_1 FILLER_65_663 ();
 sg13g2_fill_1 FILLER_65_677 ();
 sg13g2_decap_4 FILLER_65_688 ();
 sg13g2_fill_2 FILLER_65_692 ();
 sg13g2_decap_4 FILLER_65_712 ();
 sg13g2_fill_2 FILLER_65_716 ();
 sg13g2_fill_1 FILLER_65_729 ();
 sg13g2_fill_1 FILLER_65_734 ();
 sg13g2_fill_1 FILLER_65_745 ();
 sg13g2_fill_2 FILLER_65_852 ();
 sg13g2_fill_2 FILLER_65_862 ();
 sg13g2_fill_2 FILLER_65_883 ();
 sg13g2_fill_1 FILLER_65_907 ();
 sg13g2_fill_1 FILLER_65_913 ();
 sg13g2_fill_1 FILLER_65_964 ();
 sg13g2_decap_8 FILLER_65_1012 ();
 sg13g2_decap_8 FILLER_65_1019 ();
 sg13g2_decap_8 FILLER_65_1026 ();
 sg13g2_fill_2 FILLER_65_1033 ();
 sg13g2_decap_8 FILLER_65_1052 ();
 sg13g2_fill_2 FILLER_65_1059 ();
 sg13g2_fill_2 FILLER_65_1066 ();
 sg13g2_decap_8 FILLER_65_1137 ();
 sg13g2_fill_2 FILLER_65_1144 ();
 sg13g2_fill_1 FILLER_65_1146 ();
 sg13g2_decap_8 FILLER_65_1151 ();
 sg13g2_fill_2 FILLER_65_1158 ();
 sg13g2_fill_2 FILLER_65_1164 ();
 sg13g2_fill_1 FILLER_65_1166 ();
 sg13g2_decap_8 FILLER_65_1193 ();
 sg13g2_fill_2 FILLER_65_1200 ();
 sg13g2_fill_1 FILLER_65_1202 ();
 sg13g2_fill_2 FILLER_65_1230 ();
 sg13g2_decap_4 FILLER_65_1236 ();
 sg13g2_decap_8 FILLER_65_1245 ();
 sg13g2_decap_4 FILLER_65_1252 ();
 sg13g2_fill_2 FILLER_65_1266 ();
 sg13g2_fill_1 FILLER_65_1273 ();
 sg13g2_fill_2 FILLER_65_1279 ();
 sg13g2_fill_2 FILLER_65_1289 ();
 sg13g2_fill_1 FILLER_65_1314 ();
 sg13g2_fill_1 FILLER_65_1320 ();
 sg13g2_decap_8 FILLER_65_1336 ();
 sg13g2_decap_4 FILLER_65_1343 ();
 sg13g2_fill_1 FILLER_65_1353 ();
 sg13g2_fill_1 FILLER_65_1359 ();
 sg13g2_fill_1 FILLER_65_1364 ();
 sg13g2_fill_1 FILLER_65_1370 ();
 sg13g2_fill_1 FILLER_65_1375 ();
 sg13g2_decap_8 FILLER_65_1402 ();
 sg13g2_decap_4 FILLER_65_1409 ();
 sg13g2_fill_2 FILLER_65_1413 ();
 sg13g2_decap_8 FILLER_65_1425 ();
 sg13g2_decap_8 FILLER_65_1432 ();
 sg13g2_decap_8 FILLER_65_1439 ();
 sg13g2_decap_8 FILLER_65_1446 ();
 sg13g2_decap_8 FILLER_65_1453 ();
 sg13g2_decap_8 FILLER_65_1480 ();
 sg13g2_fill_1 FILLER_65_1487 ();
 sg13g2_decap_4 FILLER_65_1493 ();
 sg13g2_fill_1 FILLER_65_1505 ();
 sg13g2_fill_2 FILLER_65_1522 ();
 sg13g2_fill_1 FILLER_65_1529 ();
 sg13g2_fill_1 FILLER_65_1546 ();
 sg13g2_decap_8 FILLER_65_1591 ();
 sg13g2_fill_2 FILLER_65_1598 ();
 sg13g2_decap_4 FILLER_65_1608 ();
 sg13g2_fill_1 FILLER_65_1612 ();
 sg13g2_decap_8 FILLER_65_1638 ();
 sg13g2_decap_4 FILLER_65_1645 ();
 sg13g2_fill_1 FILLER_65_1652 ();
 sg13g2_fill_1 FILLER_65_1661 ();
 sg13g2_fill_1 FILLER_65_1667 ();
 sg13g2_fill_1 FILLER_65_1678 ();
 sg13g2_fill_2 FILLER_65_1712 ();
 sg13g2_fill_1 FILLER_65_1722 ();
 sg13g2_decap_8 FILLER_65_1759 ();
 sg13g2_decap_4 FILLER_65_1766 ();
 sg13g2_fill_1 FILLER_65_1808 ();
 sg13g2_fill_2 FILLER_65_1813 ();
 sg13g2_fill_1 FILLER_65_1840 ();
 sg13g2_fill_2 FILLER_65_1868 ();
 sg13g2_fill_2 FILLER_65_1873 ();
 sg13g2_decap_8 FILLER_65_1901 ();
 sg13g2_decap_8 FILLER_65_1908 ();
 sg13g2_fill_2 FILLER_65_1915 ();
 sg13g2_fill_1 FILLER_65_1917 ();
 sg13g2_fill_2 FILLER_65_1922 ();
 sg13g2_fill_2 FILLER_65_1934 ();
 sg13g2_fill_1 FILLER_65_1936 ();
 sg13g2_fill_1 FILLER_65_2007 ();
 sg13g2_fill_1 FILLER_65_2017 ();
 sg13g2_fill_2 FILLER_65_2023 ();
 sg13g2_decap_8 FILLER_65_2029 ();
 sg13g2_decap_8 FILLER_65_2041 ();
 sg13g2_decap_4 FILLER_65_2048 ();
 sg13g2_fill_2 FILLER_65_2052 ();
 sg13g2_decap_8 FILLER_65_2077 ();
 sg13g2_decap_8 FILLER_65_2084 ();
 sg13g2_fill_2 FILLER_65_2091 ();
 sg13g2_fill_2 FILLER_65_2133 ();
 sg13g2_fill_1 FILLER_65_2160 ();
 sg13g2_fill_1 FILLER_65_2205 ();
 sg13g2_fill_2 FILLER_65_2216 ();
 sg13g2_fill_2 FILLER_65_2248 ();
 sg13g2_fill_1 FILLER_65_2286 ();
 sg13g2_fill_2 FILLER_65_2310 ();
 sg13g2_fill_1 FILLER_65_2317 ();
 sg13g2_fill_1 FILLER_65_2330 ();
 sg13g2_fill_1 FILLER_65_2336 ();
 sg13g2_fill_1 FILLER_65_2341 ();
 sg13g2_fill_2 FILLER_65_2363 ();
 sg13g2_decap_8 FILLER_65_2405 ();
 sg13g2_fill_2 FILLER_65_2412 ();
 sg13g2_decap_4 FILLER_65_2426 ();
 sg13g2_fill_1 FILLER_65_2430 ();
 sg13g2_decap_8 FILLER_65_2436 ();
 sg13g2_fill_2 FILLER_65_2443 ();
 sg13g2_fill_2 FILLER_65_2455 ();
 sg13g2_fill_1 FILLER_65_2457 ();
 sg13g2_fill_1 FILLER_65_2493 ();
 sg13g2_fill_2 FILLER_65_2524 ();
 sg13g2_fill_1 FILLER_65_2539 ();
 sg13g2_fill_2 FILLER_65_2544 ();
 sg13g2_fill_1 FILLER_65_2546 ();
 sg13g2_fill_2 FILLER_65_2555 ();
 sg13g2_decap_4 FILLER_65_2567 ();
 sg13g2_decap_4 FILLER_65_2577 ();
 sg13g2_fill_1 FILLER_65_2581 ();
 sg13g2_decap_4 FILLER_65_2587 ();
 sg13g2_decap_4 FILLER_65_2595 ();
 sg13g2_fill_1 FILLER_65_2599 ();
 sg13g2_decap_4 FILLER_65_2604 ();
 sg13g2_decap_4 FILLER_66_0 ();
 sg13g2_fill_2 FILLER_66_4 ();
 sg13g2_fill_2 FILLER_66_10 ();
 sg13g2_decap_4 FILLER_66_32 ();
 sg13g2_fill_2 FILLER_66_70 ();
 sg13g2_fill_1 FILLER_66_72 ();
 sg13g2_decap_8 FILLER_66_77 ();
 sg13g2_decap_8 FILLER_66_84 ();
 sg13g2_fill_2 FILLER_66_91 ();
 sg13g2_fill_1 FILLER_66_93 ();
 sg13g2_fill_2 FILLER_66_129 ();
 sg13g2_decap_4 FILLER_66_147 ();
 sg13g2_decap_8 FILLER_66_159 ();
 sg13g2_fill_2 FILLER_66_166 ();
 sg13g2_decap_8 FILLER_66_174 ();
 sg13g2_decap_4 FILLER_66_181 ();
 sg13g2_fill_2 FILLER_66_185 ();
 sg13g2_decap_4 FILLER_66_196 ();
 sg13g2_fill_2 FILLER_66_210 ();
 sg13g2_decap_8 FILLER_66_234 ();
 sg13g2_decap_4 FILLER_66_241 ();
 sg13g2_fill_1 FILLER_66_245 ();
 sg13g2_fill_2 FILLER_66_249 ();
 sg13g2_decap_8 FILLER_66_255 ();
 sg13g2_fill_2 FILLER_66_262 ();
 sg13g2_fill_1 FILLER_66_264 ();
 sg13g2_decap_4 FILLER_66_286 ();
 sg13g2_fill_2 FILLER_66_290 ();
 sg13g2_decap_8 FILLER_66_297 ();
 sg13g2_decap_8 FILLER_66_304 ();
 sg13g2_decap_4 FILLER_66_311 ();
 sg13g2_fill_1 FILLER_66_315 ();
 sg13g2_fill_2 FILLER_66_321 ();
 sg13g2_fill_1 FILLER_66_323 ();
 sg13g2_fill_1 FILLER_66_329 ();
 sg13g2_decap_8 FILLER_66_335 ();
 sg13g2_decap_4 FILLER_66_342 ();
 sg13g2_fill_1 FILLER_66_346 ();
 sg13g2_fill_1 FILLER_66_375 ();
 sg13g2_fill_1 FILLER_66_388 ();
 sg13g2_fill_1 FILLER_66_394 ();
 sg13g2_fill_1 FILLER_66_400 ();
 sg13g2_fill_2 FILLER_66_406 ();
 sg13g2_decap_8 FILLER_66_412 ();
 sg13g2_fill_1 FILLER_66_436 ();
 sg13g2_fill_2 FILLER_66_442 ();
 sg13g2_fill_2 FILLER_66_474 ();
 sg13g2_fill_1 FILLER_66_476 ();
 sg13g2_fill_1 FILLER_66_481 ();
 sg13g2_decap_4 FILLER_66_487 ();
 sg13g2_fill_2 FILLER_66_495 ();
 sg13g2_decap_8 FILLER_66_501 ();
 sg13g2_fill_1 FILLER_66_508 ();
 sg13g2_decap_8 FILLER_66_524 ();
 sg13g2_decap_8 FILLER_66_531 ();
 sg13g2_fill_2 FILLER_66_543 ();
 sg13g2_fill_2 FILLER_66_587 ();
 sg13g2_fill_2 FILLER_66_595 ();
 sg13g2_fill_2 FILLER_66_603 ();
 sg13g2_decap_8 FILLER_66_625 ();
 sg13g2_decap_8 FILLER_66_641 ();
 sg13g2_fill_2 FILLER_66_648 ();
 sg13g2_fill_1 FILLER_66_650 ();
 sg13g2_fill_2 FILLER_66_660 ();
 sg13g2_fill_1 FILLER_66_662 ();
 sg13g2_decap_8 FILLER_66_705 ();
 sg13g2_fill_1 FILLER_66_712 ();
 sg13g2_fill_1 FILLER_66_765 ();
 sg13g2_fill_1 FILLER_66_862 ();
 sg13g2_fill_1 FILLER_66_901 ();
 sg13g2_fill_2 FILLER_66_976 ();
 sg13g2_fill_1 FILLER_66_978 ();
 sg13g2_fill_2 FILLER_66_988 ();
 sg13g2_fill_1 FILLER_66_1001 ();
 sg13g2_fill_2 FILLER_66_1038 ();
 sg13g2_fill_1 FILLER_66_1066 ();
 sg13g2_fill_1 FILLER_66_1084 ();
 sg13g2_decap_4 FILLER_66_1144 ();
 sg13g2_fill_2 FILLER_66_1148 ();
 sg13g2_fill_2 FILLER_66_1165 ();
 sg13g2_fill_1 FILLER_66_1167 ();
 sg13g2_fill_1 FILLER_66_1184 ();
 sg13g2_decap_8 FILLER_66_1190 ();
 sg13g2_decap_8 FILLER_66_1197 ();
 sg13g2_decap_4 FILLER_66_1204 ();
 sg13g2_fill_1 FILLER_66_1208 ();
 sg13g2_decap_4 FILLER_66_1214 ();
 sg13g2_fill_2 FILLER_66_1218 ();
 sg13g2_fill_2 FILLER_66_1226 ();
 sg13g2_decap_8 FILLER_66_1238 ();
 sg13g2_fill_1 FILLER_66_1250 ();
 sg13g2_fill_2 FILLER_66_1291 ();
 sg13g2_fill_2 FILLER_66_1304 ();
 sg13g2_fill_2 FILLER_66_1330 ();
 sg13g2_fill_2 FILLER_66_1383 ();
 sg13g2_fill_1 FILLER_66_1385 ();
 sg13g2_fill_2 FILLER_66_1391 ();
 sg13g2_fill_1 FILLER_66_1393 ();
 sg13g2_fill_2 FILLER_66_1446 ();
 sg13g2_fill_1 FILLER_66_1452 ();
 sg13g2_fill_1 FILLER_66_1466 ();
 sg13g2_decap_8 FILLER_66_1493 ();
 sg13g2_decap_8 FILLER_66_1500 ();
 sg13g2_decap_4 FILLER_66_1507 ();
 sg13g2_fill_2 FILLER_66_1511 ();
 sg13g2_decap_4 FILLER_66_1517 ();
 sg13g2_fill_2 FILLER_66_1526 ();
 sg13g2_fill_1 FILLER_66_1566 ();
 sg13g2_fill_2 FILLER_66_1587 ();
 sg13g2_fill_1 FILLER_66_1589 ();
 sg13g2_fill_2 FILLER_66_1600 ();
 sg13g2_fill_2 FILLER_66_1606 ();
 sg13g2_fill_1 FILLER_66_1608 ();
 sg13g2_fill_1 FILLER_66_1614 ();
 sg13g2_decap_8 FILLER_66_1641 ();
 sg13g2_decap_4 FILLER_66_1648 ();
 sg13g2_fill_1 FILLER_66_1652 ();
 sg13g2_decap_4 FILLER_66_1657 ();
 sg13g2_fill_2 FILLER_66_1661 ();
 sg13g2_fill_1 FILLER_66_1673 ();
 sg13g2_fill_2 FILLER_66_1678 ();
 sg13g2_fill_1 FILLER_66_1680 ();
 sg13g2_fill_2 FILLER_66_1686 ();
 sg13g2_decap_4 FILLER_66_1697 ();
 sg13g2_fill_2 FILLER_66_1701 ();
 sg13g2_decap_4 FILLER_66_1713 ();
 sg13g2_decap_4 FILLER_66_1721 ();
 sg13g2_fill_2 FILLER_66_1725 ();
 sg13g2_decap_8 FILLER_66_1737 ();
 sg13g2_decap_4 FILLER_66_1744 ();
 sg13g2_fill_1 FILLER_66_1748 ();
 sg13g2_fill_1 FILLER_66_1759 ();
 sg13g2_decap_8 FILLER_66_1764 ();
 sg13g2_decap_8 FILLER_66_1775 ();
 sg13g2_fill_1 FILLER_66_1782 ();
 sg13g2_fill_1 FILLER_66_1797 ();
 sg13g2_fill_2 FILLER_66_1802 ();
 sg13g2_fill_1 FILLER_66_1804 ();
 sg13g2_fill_2 FILLER_66_1810 ();
 sg13g2_fill_1 FILLER_66_1812 ();
 sg13g2_fill_2 FILLER_66_1834 ();
 sg13g2_fill_1 FILLER_66_1846 ();
 sg13g2_fill_2 FILLER_66_1861 ();
 sg13g2_fill_2 FILLER_66_1889 ();
 sg13g2_decap_8 FILLER_66_1896 ();
 sg13g2_decap_8 FILLER_66_1903 ();
 sg13g2_decap_8 FILLER_66_1910 ();
 sg13g2_decap_8 FILLER_66_1917 ();
 sg13g2_decap_4 FILLER_66_1924 ();
 sg13g2_fill_1 FILLER_66_1928 ();
 sg13g2_fill_1 FILLER_66_1937 ();
 sg13g2_decap_4 FILLER_66_1942 ();
 sg13g2_fill_2 FILLER_66_1958 ();
 sg13g2_fill_2 FILLER_66_1980 ();
 sg13g2_fill_1 FILLER_66_2010 ();
 sg13g2_decap_4 FILLER_66_2016 ();
 sg13g2_decap_8 FILLER_66_2024 ();
 sg13g2_decap_8 FILLER_66_2031 ();
 sg13g2_decap_8 FILLER_66_2038 ();
 sg13g2_fill_2 FILLER_66_2045 ();
 sg13g2_decap_4 FILLER_66_2077 ();
 sg13g2_fill_1 FILLER_66_2081 ();
 sg13g2_fill_2 FILLER_66_2138 ();
 sg13g2_fill_1 FILLER_66_2192 ();
 sg13g2_fill_2 FILLER_66_2327 ();
 sg13g2_fill_1 FILLER_66_2362 ();
 sg13g2_fill_1 FILLER_66_2372 ();
 sg13g2_fill_1 FILLER_66_2377 ();
 sg13g2_fill_1 FILLER_66_2382 ();
 sg13g2_fill_2 FILLER_66_2409 ();
 sg13g2_fill_2 FILLER_66_2416 ();
 sg13g2_fill_2 FILLER_66_2422 ();
 sg13g2_fill_1 FILLER_66_2424 ();
 sg13g2_fill_1 FILLER_66_2455 ();
 sg13g2_fill_1 FILLER_66_2469 ();
 sg13g2_decap_8 FILLER_66_2528 ();
 sg13g2_decap_8 FILLER_66_2535 ();
 sg13g2_decap_8 FILLER_66_2593 ();
 sg13g2_decap_8 FILLER_66_2600 ();
 sg13g2_decap_8 FILLER_66_2607 ();
 sg13g2_decap_8 FILLER_66_2614 ();
 sg13g2_fill_2 FILLER_66_2621 ();
 sg13g2_fill_1 FILLER_66_2623 ();
 sg13g2_decap_8 FILLER_66_2638 ();
 sg13g2_fill_2 FILLER_66_2645 ();
 sg13g2_fill_1 FILLER_66_2647 ();
 sg13g2_fill_1 FILLER_66_2652 ();
 sg13g2_decap_8 FILLER_66_2657 ();
 sg13g2_decap_4 FILLER_66_2664 ();
 sg13g2_fill_2 FILLER_66_2668 ();
 sg13g2_decap_8 FILLER_67_0 ();
 sg13g2_decap_8 FILLER_67_7 ();
 sg13g2_decap_4 FILLER_67_14 ();
 sg13g2_decap_8 FILLER_67_71 ();
 sg13g2_decap_8 FILLER_67_78 ();
 sg13g2_fill_2 FILLER_67_85 ();
 sg13g2_fill_1 FILLER_67_87 ();
 sg13g2_decap_4 FILLER_67_100 ();
 sg13g2_decap_4 FILLER_67_164 ();
 sg13g2_fill_1 FILLER_67_168 ();
 sg13g2_fill_2 FILLER_67_195 ();
 sg13g2_fill_1 FILLER_67_197 ();
 sg13g2_decap_8 FILLER_67_233 ();
 sg13g2_fill_2 FILLER_67_240 ();
 sg13g2_fill_1 FILLER_67_242 ();
 sg13g2_decap_8 FILLER_67_246 ();
 sg13g2_decap_8 FILLER_67_253 ();
 sg13g2_decap_8 FILLER_67_260 ();
 sg13g2_decap_8 FILLER_67_267 ();
 sg13g2_decap_8 FILLER_67_274 ();
 sg13g2_fill_2 FILLER_67_291 ();
 sg13g2_fill_1 FILLER_67_302 ();
 sg13g2_decap_4 FILLER_67_307 ();
 sg13g2_fill_1 FILLER_67_311 ();
 sg13g2_fill_2 FILLER_67_356 ();
 sg13g2_fill_1 FILLER_67_358 ();
 sg13g2_decap_8 FILLER_67_388 ();
 sg13g2_decap_4 FILLER_67_395 ();
 sg13g2_fill_1 FILLER_67_399 ();
 sg13g2_fill_1 FILLER_67_404 ();
 sg13g2_decap_8 FILLER_67_410 ();
 sg13g2_fill_2 FILLER_67_417 ();
 sg13g2_decap_8 FILLER_67_463 ();
 sg13g2_fill_1 FILLER_67_470 ();
 sg13g2_decap_8 FILLER_67_475 ();
 sg13g2_fill_1 FILLER_67_482 ();
 sg13g2_fill_1 FILLER_67_522 ();
 sg13g2_fill_2 FILLER_67_554 ();
 sg13g2_fill_2 FILLER_67_568 ();
 sg13g2_fill_1 FILLER_67_573 ();
 sg13g2_fill_2 FILLER_67_631 ();
 sg13g2_fill_1 FILLER_67_633 ();
 sg13g2_decap_4 FILLER_67_664 ();
 sg13g2_fill_1 FILLER_67_668 ();
 sg13g2_decap_8 FILLER_67_705 ();
 sg13g2_decap_4 FILLER_67_712 ();
 sg13g2_fill_2 FILLER_67_766 ();
 sg13g2_fill_2 FILLER_67_805 ();
 sg13g2_fill_2 FILLER_67_815 ();
 sg13g2_fill_1 FILLER_67_821 ();
 sg13g2_fill_1 FILLER_67_980 ();
 sg13g2_fill_1 FILLER_67_994 ();
 sg13g2_fill_2 FILLER_67_1014 ();
 sg13g2_decap_8 FILLER_67_1020 ();
 sg13g2_decap_8 FILLER_67_1027 ();
 sg13g2_decap_8 FILLER_67_1034 ();
 sg13g2_fill_1 FILLER_67_1041 ();
 sg13g2_decap_8 FILLER_67_1051 ();
 sg13g2_fill_2 FILLER_67_1058 ();
 sg13g2_fill_1 FILLER_67_1060 ();
 sg13g2_decap_4 FILLER_67_1121 ();
 sg13g2_fill_1 FILLER_67_1125 ();
 sg13g2_decap_8 FILLER_67_1130 ();
 sg13g2_decap_8 FILLER_67_1137 ();
 sg13g2_decap_8 FILLER_67_1144 ();
 sg13g2_fill_2 FILLER_67_1151 ();
 sg13g2_fill_1 FILLER_67_1153 ();
 sg13g2_fill_1 FILLER_67_1159 ();
 sg13g2_fill_2 FILLER_67_1170 ();
 sg13g2_fill_1 FILLER_67_1172 ();
 sg13g2_decap_8 FILLER_67_1195 ();
 sg13g2_decap_4 FILLER_67_1206 ();
 sg13g2_decap_8 FILLER_67_1225 ();
 sg13g2_fill_1 FILLER_67_1232 ();
 sg13g2_fill_1 FILLER_67_1269 ();
 sg13g2_decap_8 FILLER_67_1289 ();
 sg13g2_fill_1 FILLER_67_1296 ();
 sg13g2_fill_1 FILLER_67_1307 ();
 sg13g2_fill_1 FILLER_67_1342 ();
 sg13g2_decap_4 FILLER_67_1364 ();
 sg13g2_fill_1 FILLER_67_1381 ();
 sg13g2_fill_1 FILLER_67_1415 ();
 sg13g2_fill_1 FILLER_67_1450 ();
 sg13g2_decap_4 FILLER_67_1475 ();
 sg13g2_fill_2 FILLER_67_1479 ();
 sg13g2_fill_1 FILLER_67_1507 ();
 sg13g2_fill_1 FILLER_67_1512 ();
 sg13g2_fill_2 FILLER_67_1521 ();
 sg13g2_fill_2 FILLER_67_1528 ();
 sg13g2_fill_1 FILLER_67_1547 ();
 sg13g2_fill_2 FILLER_67_1576 ();
 sg13g2_fill_2 FILLER_67_1609 ();
 sg13g2_fill_2 FILLER_67_1616 ();
 sg13g2_fill_1 FILLER_67_1618 ();
 sg13g2_fill_1 FILLER_67_1624 ();
 sg13g2_decap_4 FILLER_67_1648 ();
 sg13g2_fill_1 FILLER_67_1652 ();
 sg13g2_fill_1 FILLER_67_1681 ();
 sg13g2_fill_2 FILLER_67_1686 ();
 sg13g2_decap_8 FILLER_67_1696 ();
 sg13g2_decap_4 FILLER_67_1703 ();
 sg13g2_fill_1 FILLER_67_1707 ();
 sg13g2_decap_8 FILLER_67_1732 ();
 sg13g2_decap_8 FILLER_67_1739 ();
 sg13g2_fill_1 FILLER_67_1746 ();
 sg13g2_fill_2 FILLER_67_1752 ();
 sg13g2_fill_1 FILLER_67_1754 ();
 sg13g2_decap_8 FILLER_67_1763 ();
 sg13g2_decap_8 FILLER_67_1770 ();
 sg13g2_decap_4 FILLER_67_1777 ();
 sg13g2_fill_2 FILLER_67_1781 ();
 sg13g2_fill_1 FILLER_67_1810 ();
 sg13g2_fill_2 FILLER_67_1865 ();
 sg13g2_fill_1 FILLER_67_1867 ();
 sg13g2_decap_4 FILLER_67_1890 ();
 sg13g2_fill_2 FILLER_67_1894 ();
 sg13g2_decap_8 FILLER_67_1900 ();
 sg13g2_decap_8 FILLER_67_1907 ();
 sg13g2_fill_1 FILLER_67_1914 ();
 sg13g2_fill_2 FILLER_67_1920 ();
 sg13g2_fill_1 FILLER_67_1922 ();
 sg13g2_fill_1 FILLER_67_1944 ();
 sg13g2_fill_1 FILLER_67_1949 ();
 sg13g2_fill_2 FILLER_67_1958 ();
 sg13g2_fill_2 FILLER_67_1964 ();
 sg13g2_fill_1 FILLER_67_2004 ();
 sg13g2_decap_8 FILLER_67_2027 ();
 sg13g2_fill_2 FILLER_67_2034 ();
 sg13g2_decap_4 FILLER_67_2098 ();
 sg13g2_fill_1 FILLER_67_2102 ();
 sg13g2_decap_4 FILLER_67_2127 ();
 sg13g2_fill_1 FILLER_67_2180 ();
 sg13g2_fill_2 FILLER_67_2227 ();
 sg13g2_fill_2 FILLER_67_2250 ();
 sg13g2_fill_1 FILLER_67_2271 ();
 sg13g2_fill_1 FILLER_67_2285 ();
 sg13g2_fill_1 FILLER_67_2292 ();
 sg13g2_fill_1 FILLER_67_2298 ();
 sg13g2_fill_1 FILLER_67_2408 ();
 sg13g2_fill_1 FILLER_67_2467 ();
 sg13g2_fill_2 FILLER_67_2477 ();
 sg13g2_decap_8 FILLER_67_2485 ();
 sg13g2_fill_2 FILLER_67_2497 ();
 sg13g2_fill_1 FILLER_67_2499 ();
 sg13g2_fill_1 FILLER_67_2574 ();
 sg13g2_fill_1 FILLER_67_2589 ();
 sg13g2_decap_8 FILLER_67_2620 ();
 sg13g2_decap_8 FILLER_67_2627 ();
 sg13g2_decap_8 FILLER_67_2634 ();
 sg13g2_decap_8 FILLER_67_2641 ();
 sg13g2_decap_8 FILLER_67_2648 ();
 sg13g2_decap_8 FILLER_67_2655 ();
 sg13g2_decap_8 FILLER_67_2662 ();
 sg13g2_fill_1 FILLER_67_2669 ();
 sg13g2_decap_8 FILLER_68_0 ();
 sg13g2_decap_4 FILLER_68_7 ();
 sg13g2_fill_1 FILLER_68_11 ();
 sg13g2_decap_4 FILLER_68_32 ();
 sg13g2_fill_1 FILLER_68_80 ();
 sg13g2_fill_2 FILLER_68_97 ();
 sg13g2_fill_1 FILLER_68_130 ();
 sg13g2_fill_1 FILLER_68_136 ();
 sg13g2_fill_1 FILLER_68_168 ();
 sg13g2_fill_2 FILLER_68_173 ();
 sg13g2_decap_8 FILLER_68_237 ();
 sg13g2_decap_8 FILLER_68_244 ();
 sg13g2_decap_8 FILLER_68_251 ();
 sg13g2_fill_2 FILLER_68_262 ();
 sg13g2_fill_1 FILLER_68_264 ();
 sg13g2_fill_1 FILLER_68_286 ();
 sg13g2_fill_1 FILLER_68_292 ();
 sg13g2_fill_1 FILLER_68_319 ();
 sg13g2_fill_1 FILLER_68_325 ();
 sg13g2_fill_2 FILLER_68_352 ();
 sg13g2_fill_1 FILLER_68_359 ();
 sg13g2_fill_1 FILLER_68_366 ();
 sg13g2_fill_2 FILLER_68_388 ();
 sg13g2_fill_1 FILLER_68_390 ();
 sg13g2_fill_2 FILLER_68_418 ();
 sg13g2_fill_1 FILLER_68_429 ();
 sg13g2_fill_1 FILLER_68_434 ();
 sg13g2_decap_4 FILLER_68_465 ();
 sg13g2_fill_2 FILLER_68_469 ();
 sg13g2_fill_1 FILLER_68_476 ();
 sg13g2_fill_2 FILLER_68_503 ();
 sg13g2_fill_2 FILLER_68_531 ();
 sg13g2_fill_2 FILLER_68_537 ();
 sg13g2_fill_1 FILLER_68_539 ();
 sg13g2_fill_1 FILLER_68_544 ();
 sg13g2_fill_1 FILLER_68_568 ();
 sg13g2_fill_1 FILLER_68_581 ();
 sg13g2_decap_8 FILLER_68_651 ();
 sg13g2_decap_8 FILLER_68_658 ();
 sg13g2_decap_8 FILLER_68_665 ();
 sg13g2_fill_1 FILLER_68_672 ();
 sg13g2_fill_2 FILLER_68_677 ();
 sg13g2_fill_1 FILLER_68_679 ();
 sg13g2_decap_4 FILLER_68_690 ();
 sg13g2_fill_1 FILLER_68_694 ();
 sg13g2_fill_1 FILLER_68_738 ();
 sg13g2_fill_1 FILLER_68_811 ();
 sg13g2_fill_1 FILLER_68_815 ();
 sg13g2_fill_2 FILLER_68_833 ();
 sg13g2_fill_2 FILLER_68_844 ();
 sg13g2_fill_2 FILLER_68_861 ();
 sg13g2_fill_2 FILLER_68_867 ();
 sg13g2_fill_2 FILLER_68_949 ();
 sg13g2_fill_1 FILLER_68_982 ();
 sg13g2_fill_1 FILLER_68_1009 ();
 sg13g2_fill_1 FILLER_68_1036 ();
 sg13g2_fill_2 FILLER_68_1055 ();
 sg13g2_fill_2 FILLER_68_1074 ();
 sg13g2_fill_1 FILLER_68_1106 ();
 sg13g2_decap_4 FILLER_68_1133 ();
 sg13g2_fill_2 FILLER_68_1147 ();
 sg13g2_fill_1 FILLER_68_1149 ();
 sg13g2_fill_2 FILLER_68_1180 ();
 sg13g2_decap_4 FILLER_68_1213 ();
 sg13g2_fill_1 FILLER_68_1238 ();
 sg13g2_fill_1 FILLER_68_1245 ();
 sg13g2_fill_1 FILLER_68_1267 ();
 sg13g2_fill_1 FILLER_68_1271 ();
 sg13g2_decap_8 FILLER_68_1281 ();
 sg13g2_fill_2 FILLER_68_1288 ();
 sg13g2_decap_4 FILLER_68_1294 ();
 sg13g2_fill_2 FILLER_68_1298 ();
 sg13g2_fill_1 FILLER_68_1304 ();
 sg13g2_fill_1 FILLER_68_1343 ();
 sg13g2_decap_8 FILLER_68_1358 ();
 sg13g2_fill_2 FILLER_68_1365 ();
 sg13g2_fill_2 FILLER_68_1371 ();
 sg13g2_fill_1 FILLER_68_1373 ();
 sg13g2_decap_4 FILLER_68_1403 ();
 sg13g2_decap_4 FILLER_68_1411 ();
 sg13g2_decap_4 FILLER_68_1423 ();
 sg13g2_decap_8 FILLER_68_1467 ();
 sg13g2_decap_8 FILLER_68_1474 ();
 sg13g2_fill_2 FILLER_68_1481 ();
 sg13g2_fill_1 FILLER_68_1483 ();
 sg13g2_fill_1 FILLER_68_1515 ();
 sg13g2_fill_1 FILLER_68_1520 ();
 sg13g2_fill_1 FILLER_68_1529 ();
 sg13g2_fill_1 FILLER_68_1547 ();
 sg13g2_fill_1 FILLER_68_1598 ();
 sg13g2_fill_2 FILLER_68_1650 ();
 sg13g2_fill_1 FILLER_68_1652 ();
 sg13g2_fill_2 FILLER_68_1660 ();
 sg13g2_fill_2 FILLER_68_1669 ();
 sg13g2_fill_1 FILLER_68_1671 ();
 sg13g2_fill_1 FILLER_68_1677 ();
 sg13g2_decap_8 FILLER_68_1683 ();
 sg13g2_fill_2 FILLER_68_1690 ();
 sg13g2_fill_1 FILLER_68_1692 ();
 sg13g2_fill_2 FILLER_68_1700 ();
 sg13g2_decap_4 FILLER_68_1706 ();
 sg13g2_fill_2 FILLER_68_1746 ();
 sg13g2_fill_2 FILLER_68_1752 ();
 sg13g2_fill_1 FILLER_68_1754 ();
 sg13g2_decap_8 FILLER_68_1760 ();
 sg13g2_decap_8 FILLER_68_1767 ();
 sg13g2_decap_8 FILLER_68_1774 ();
 sg13g2_decap_4 FILLER_68_1781 ();
 sg13g2_fill_2 FILLER_68_1785 ();
 sg13g2_decap_4 FILLER_68_1805 ();
 sg13g2_fill_1 FILLER_68_1822 ();
 sg13g2_fill_2 FILLER_68_1829 ();
 sg13g2_fill_1 FILLER_68_1836 ();
 sg13g2_decap_4 FILLER_68_1841 ();
 sg13g2_fill_1 FILLER_68_1860 ();
 sg13g2_fill_1 FILLER_68_1874 ();
 sg13g2_fill_2 FILLER_68_1880 ();
 sg13g2_fill_2 FILLER_68_1888 ();
 sg13g2_decap_8 FILLER_68_1896 ();
 sg13g2_decap_8 FILLER_68_1903 ();
 sg13g2_decap_8 FILLER_68_1910 ();
 sg13g2_decap_4 FILLER_68_1917 ();
 sg13g2_fill_2 FILLER_68_1921 ();
 sg13g2_fill_2 FILLER_68_1931 ();
 sg13g2_fill_1 FILLER_68_1933 ();
 sg13g2_fill_1 FILLER_68_1939 ();
 sg13g2_decap_8 FILLER_68_1947 ();
 sg13g2_fill_2 FILLER_68_1954 ();
 sg13g2_fill_1 FILLER_68_1960 ();
 sg13g2_decap_4 FILLER_68_1975 ();
 sg13g2_fill_2 FILLER_68_1979 ();
 sg13g2_fill_1 FILLER_68_1989 ();
 sg13g2_fill_1 FILLER_68_2004 ();
 sg13g2_fill_1 FILLER_68_2011 ();
 sg13g2_fill_1 FILLER_68_2023 ();
 sg13g2_decap_4 FILLER_68_2028 ();
 sg13g2_fill_1 FILLER_68_2032 ();
 sg13g2_fill_2 FILLER_68_2038 ();
 sg13g2_fill_1 FILLER_68_2040 ();
 sg13g2_fill_1 FILLER_68_2051 ();
 sg13g2_fill_1 FILLER_68_2077 ();
 sg13g2_decap_8 FILLER_68_2082 ();
 sg13g2_fill_1 FILLER_68_2089 ();
 sg13g2_fill_1 FILLER_68_2110 ();
 sg13g2_fill_1 FILLER_68_2115 ();
 sg13g2_fill_1 FILLER_68_2134 ();
 sg13g2_fill_1 FILLER_68_2156 ();
 sg13g2_fill_2 FILLER_68_2203 ();
 sg13g2_fill_2 FILLER_68_2248 ();
 sg13g2_fill_1 FILLER_68_2280 ();
 sg13g2_fill_1 FILLER_68_2289 ();
 sg13g2_fill_1 FILLER_68_2295 ();
 sg13g2_fill_2 FILLER_68_2302 ();
 sg13g2_fill_2 FILLER_68_2318 ();
 sg13g2_fill_2 FILLER_68_2324 ();
 sg13g2_fill_2 FILLER_68_2340 ();
 sg13g2_fill_1 FILLER_68_2356 ();
 sg13g2_fill_1 FILLER_68_2363 ();
 sg13g2_fill_2 FILLER_68_2378 ();
 sg13g2_fill_1 FILLER_68_2385 ();
 sg13g2_fill_1 FILLER_68_2479 ();
 sg13g2_fill_2 FILLER_68_2485 ();
 sg13g2_fill_1 FILLER_68_2491 ();
 sg13g2_decap_8 FILLER_68_2569 ();
 sg13g2_fill_2 FILLER_68_2576 ();
 sg13g2_fill_1 FILLER_68_2578 ();
 sg13g2_decap_8 FILLER_68_2622 ();
 sg13g2_decap_8 FILLER_68_2629 ();
 sg13g2_decap_8 FILLER_68_2636 ();
 sg13g2_decap_8 FILLER_68_2643 ();
 sg13g2_decap_8 FILLER_68_2650 ();
 sg13g2_decap_8 FILLER_68_2657 ();
 sg13g2_decap_4 FILLER_68_2664 ();
 sg13g2_fill_2 FILLER_68_2668 ();
 sg13g2_decap_4 FILLER_69_0 ();
 sg13g2_fill_2 FILLER_69_4 ();
 sg13g2_decap_8 FILLER_69_36 ();
 sg13g2_decap_4 FILLER_69_47 ();
 sg13g2_fill_1 FILLER_69_51 ();
 sg13g2_fill_1 FILLER_69_147 ();
 sg13g2_decap_4 FILLER_69_172 ();
 sg13g2_fill_2 FILLER_69_185 ();
 sg13g2_fill_1 FILLER_69_192 ();
 sg13g2_fill_1 FILLER_69_206 ();
 sg13g2_fill_2 FILLER_69_225 ();
 sg13g2_fill_2 FILLER_69_232 ();
 sg13g2_fill_1 FILLER_69_291 ();
 sg13g2_fill_1 FILLER_69_297 ();
 sg13g2_fill_1 FILLER_69_309 ();
 sg13g2_fill_2 FILLER_69_350 ();
 sg13g2_fill_1 FILLER_69_358 ();
 sg13g2_fill_1 FILLER_69_366 ();
 sg13g2_fill_2 FILLER_69_424 ();
 sg13g2_decap_4 FILLER_69_431 ();
 sg13g2_fill_2 FILLER_69_435 ();
 sg13g2_fill_2 FILLER_69_445 ();
 sg13g2_fill_1 FILLER_69_447 ();
 sg13g2_decap_8 FILLER_69_452 ();
 sg13g2_decap_8 FILLER_69_459 ();
 sg13g2_fill_2 FILLER_69_479 ();
 sg13g2_fill_1 FILLER_69_481 ();
 sg13g2_fill_1 FILLER_69_486 ();
 sg13g2_fill_2 FILLER_69_495 ();
 sg13g2_decap_8 FILLER_69_536 ();
 sg13g2_fill_1 FILLER_69_543 ();
 sg13g2_fill_2 FILLER_69_555 ();
 sg13g2_fill_1 FILLER_69_557 ();
 sg13g2_fill_2 FILLER_69_574 ();
 sg13g2_fill_1 FILLER_69_576 ();
 sg13g2_fill_2 FILLER_69_581 ();
 sg13g2_fill_2 FILLER_69_589 ();
 sg13g2_decap_8 FILLER_69_595 ();
 sg13g2_fill_1 FILLER_69_602 ();
 sg13g2_fill_1 FILLER_69_608 ();
 sg13g2_fill_1 FILLER_69_635 ();
 sg13g2_fill_2 FILLER_69_662 ();
 sg13g2_fill_1 FILLER_69_664 ();
 sg13g2_decap_4 FILLER_69_695 ();
 sg13g2_fill_1 FILLER_69_710 ();
 sg13g2_fill_1 FILLER_69_756 ();
 sg13g2_fill_1 FILLER_69_768 ();
 sg13g2_fill_1 FILLER_69_843 ();
 sg13g2_decap_8 FILLER_69_854 ();
 sg13g2_fill_1 FILLER_69_861 ();
 sg13g2_decap_4 FILLER_69_868 ();
 sg13g2_decap_8 FILLER_69_876 ();
 sg13g2_fill_1 FILLER_69_892 ();
 sg13g2_fill_2 FILLER_69_904 ();
 sg13g2_decap_8 FILLER_69_941 ();
 sg13g2_fill_2 FILLER_69_948 ();
 sg13g2_fill_1 FILLER_69_950 ();
 sg13g2_fill_2 FILLER_69_965 ();
 sg13g2_fill_1 FILLER_69_1001 ();
 sg13g2_decap_4 FILLER_69_1012 ();
 sg13g2_fill_2 FILLER_69_1061 ();
 sg13g2_fill_1 FILLER_69_1063 ();
 sg13g2_fill_2 FILLER_69_1072 ();
 sg13g2_fill_2 FILLER_69_1126 ();
 sg13g2_decap_4 FILLER_69_1142 ();
 sg13g2_decap_4 FILLER_69_1150 ();
 sg13g2_fill_2 FILLER_69_1154 ();
 sg13g2_decap_8 FILLER_69_1186 ();
 sg13g2_fill_2 FILLER_69_1193 ();
 sg13g2_decap_4 FILLER_69_1199 ();
 sg13g2_fill_2 FILLER_69_1225 ();
 sg13g2_fill_1 FILLER_69_1256 ();
 sg13g2_decap_8 FILLER_69_1262 ();
 sg13g2_fill_1 FILLER_69_1269 ();
 sg13g2_decap_8 FILLER_69_1276 ();
 sg13g2_fill_2 FILLER_69_1288 ();
 sg13g2_decap_8 FILLER_69_1307 ();
 sg13g2_decap_4 FILLER_69_1314 ();
 sg13g2_fill_1 FILLER_69_1318 ();
 sg13g2_fill_2 FILLER_69_1325 ();
 sg13g2_fill_1 FILLER_69_1335 ();
 sg13g2_fill_2 FILLER_69_1339 ();
 sg13g2_fill_1 FILLER_69_1346 ();
 sg13g2_decap_8 FILLER_69_1365 ();
 sg13g2_fill_1 FILLER_69_1372 ();
 sg13g2_decap_4 FILLER_69_1376 ();
 sg13g2_decap_4 FILLER_69_1394 ();
 sg13g2_fill_1 FILLER_69_1398 ();
 sg13g2_decap_4 FILLER_69_1435 ();
 sg13g2_decap_8 FILLER_69_1449 ();
 sg13g2_decap_8 FILLER_69_1460 ();
 sg13g2_fill_2 FILLER_69_1467 ();
 sg13g2_fill_1 FILLER_69_1469 ();
 sg13g2_decap_4 FILLER_69_1480 ();
 sg13g2_fill_2 FILLER_69_1484 ();
 sg13g2_decap_4 FILLER_69_1494 ();
 sg13g2_fill_2 FILLER_69_1498 ();
 sg13g2_fill_2 FILLER_69_1512 ();
 sg13g2_fill_1 FILLER_69_1522 ();
 sg13g2_fill_2 FILLER_69_1576 ();
 sg13g2_fill_2 FILLER_69_1583 ();
 sg13g2_fill_1 FILLER_69_1613 ();
 sg13g2_fill_1 FILLER_69_1627 ();
 sg13g2_fill_2 FILLER_69_1654 ();
 sg13g2_fill_1 FILLER_69_1656 ();
 sg13g2_fill_2 FILLER_69_1661 ();
 sg13g2_fill_2 FILLER_69_1668 ();
 sg13g2_fill_2 FILLER_69_1675 ();
 sg13g2_fill_1 FILLER_69_1677 ();
 sg13g2_decap_4 FILLER_69_1704 ();
 sg13g2_decap_4 FILLER_69_1712 ();
 sg13g2_fill_1 FILLER_69_1716 ();
 sg13g2_decap_8 FILLER_69_1750 ();
 sg13g2_decap_8 FILLER_69_1757 ();
 sg13g2_decap_8 FILLER_69_1764 ();
 sg13g2_decap_8 FILLER_69_1771 ();
 sg13g2_fill_1 FILLER_69_1778 ();
 sg13g2_decap_4 FILLER_69_1790 ();
 sg13g2_fill_1 FILLER_69_1794 ();
 sg13g2_fill_1 FILLER_69_1828 ();
 sg13g2_fill_1 FILLER_69_1833 ();
 sg13g2_fill_1 FILLER_69_1839 ();
 sg13g2_decap_4 FILLER_69_1846 ();
 sg13g2_fill_2 FILLER_69_1850 ();
 sg13g2_fill_1 FILLER_69_1857 ();
 sg13g2_decap_4 FILLER_69_1873 ();
 sg13g2_fill_2 FILLER_69_1881 ();
 sg13g2_fill_1 FILLER_69_1896 ();
 sg13g2_decap_8 FILLER_69_1927 ();
 sg13g2_decap_8 FILLER_69_1934 ();
 sg13g2_decap_4 FILLER_69_1941 ();
 sg13g2_fill_1 FILLER_69_1945 ();
 sg13g2_fill_2 FILLER_69_1950 ();
 sg13g2_fill_1 FILLER_69_1968 ();
 sg13g2_fill_1 FILLER_69_2020 ();
 sg13g2_decap_8 FILLER_69_2029 ();
 sg13g2_fill_2 FILLER_69_2036 ();
 sg13g2_decap_4 FILLER_69_2042 ();
 sg13g2_fill_2 FILLER_69_2046 ();
 sg13g2_decap_4 FILLER_69_2057 ();
 sg13g2_fill_2 FILLER_69_2065 ();
 sg13g2_decap_4 FILLER_69_2088 ();
 sg13g2_fill_1 FILLER_69_2123 ();
 sg13g2_decap_8 FILLER_69_2153 ();
 sg13g2_fill_2 FILLER_69_2160 ();
 sg13g2_fill_1 FILLER_69_2177 ();
 sg13g2_fill_2 FILLER_69_2184 ();
 sg13g2_fill_1 FILLER_69_2196 ();
 sg13g2_fill_2 FILLER_69_2243 ();
 sg13g2_fill_1 FILLER_69_2245 ();
 sg13g2_fill_1 FILLER_69_2273 ();
 sg13g2_decap_8 FILLER_69_2401 ();
 sg13g2_fill_1 FILLER_69_2416 ();
 sg13g2_fill_1 FILLER_69_2442 ();
 sg13g2_fill_2 FILLER_69_2474 ();
 sg13g2_fill_2 FILLER_69_2502 ();
 sg13g2_fill_2 FILLER_69_2522 ();
 sg13g2_fill_1 FILLER_69_2546 ();
 sg13g2_fill_2 FILLER_69_2570 ();
 sg13g2_decap_8 FILLER_69_2622 ();
 sg13g2_decap_8 FILLER_69_2629 ();
 sg13g2_decap_8 FILLER_69_2636 ();
 sg13g2_decap_8 FILLER_69_2643 ();
 sg13g2_decap_8 FILLER_69_2650 ();
 sg13g2_decap_8 FILLER_69_2657 ();
 sg13g2_decap_4 FILLER_69_2664 ();
 sg13g2_fill_2 FILLER_69_2668 ();
 sg13g2_decap_4 FILLER_70_0 ();
 sg13g2_fill_2 FILLER_70_4 ();
 sg13g2_decap_4 FILLER_70_32 ();
 sg13g2_decap_4 FILLER_70_62 ();
 sg13g2_fill_1 FILLER_70_66 ();
 sg13g2_fill_1 FILLER_70_100 ();
 sg13g2_fill_2 FILLER_70_132 ();
 sg13g2_fill_1 FILLER_70_156 ();
 sg13g2_decap_8 FILLER_70_173 ();
 sg13g2_decap_8 FILLER_70_180 ();
 sg13g2_decap_4 FILLER_70_187 ();
 sg13g2_decap_8 FILLER_70_200 ();
 sg13g2_fill_2 FILLER_70_207 ();
 sg13g2_fill_1 FILLER_70_209 ();
 sg13g2_fill_1 FILLER_70_218 ();
 sg13g2_fill_1 FILLER_70_245 ();
 sg13g2_fill_1 FILLER_70_272 ();
 sg13g2_fill_1 FILLER_70_277 ();
 sg13g2_fill_1 FILLER_70_288 ();
 sg13g2_fill_2 FILLER_70_302 ();
 sg13g2_fill_1 FILLER_70_304 ();
 sg13g2_decap_8 FILLER_70_310 ();
 sg13g2_decap_4 FILLER_70_321 ();
 sg13g2_fill_2 FILLER_70_325 ();
 sg13g2_decap_8 FILLER_70_348 ();
 sg13g2_decap_8 FILLER_70_355 ();
 sg13g2_fill_2 FILLER_70_362 ();
 sg13g2_decap_8 FILLER_70_369 ();
 sg13g2_decap_8 FILLER_70_376 ();
 sg13g2_fill_2 FILLER_70_393 ();
 sg13g2_fill_1 FILLER_70_395 ();
 sg13g2_decap_8 FILLER_70_422 ();
 sg13g2_decap_4 FILLER_70_429 ();
 sg13g2_fill_1 FILLER_70_433 ();
 sg13g2_decap_8 FILLER_70_438 ();
 sg13g2_decap_8 FILLER_70_445 ();
 sg13g2_fill_2 FILLER_70_452 ();
 sg13g2_fill_1 FILLER_70_493 ();
 sg13g2_fill_1 FILLER_70_506 ();
 sg13g2_fill_2 FILLER_70_519 ();
 sg13g2_decap_4 FILLER_70_527 ();
 sg13g2_decap_4 FILLER_70_580 ();
 sg13g2_fill_1 FILLER_70_584 ();
 sg13g2_decap_4 FILLER_70_604 ();
 sg13g2_fill_1 FILLER_70_612 ();
 sg13g2_fill_2 FILLER_70_621 ();
 sg13g2_decap_4 FILLER_70_657 ();
 sg13g2_fill_1 FILLER_70_708 ();
 sg13g2_fill_2 FILLER_70_717 ();
 sg13g2_fill_1 FILLER_70_719 ();
 sg13g2_decap_4 FILLER_70_734 ();
 sg13g2_fill_1 FILLER_70_738 ();
 sg13g2_fill_1 FILLER_70_749 ();
 sg13g2_fill_2 FILLER_70_753 ();
 sg13g2_fill_2 FILLER_70_761 ();
 sg13g2_fill_1 FILLER_70_808 ();
 sg13g2_fill_1 FILLER_70_819 ();
 sg13g2_fill_2 FILLER_70_846 ();
 sg13g2_fill_2 FILLER_70_874 ();
 sg13g2_fill_2 FILLER_70_898 ();
 sg13g2_decap_8 FILLER_70_930 ();
 sg13g2_decap_4 FILLER_70_937 ();
 sg13g2_fill_1 FILLER_70_941 ();
 sg13g2_decap_4 FILLER_70_951 ();
 sg13g2_fill_2 FILLER_70_955 ();
 sg13g2_fill_1 FILLER_70_961 ();
 sg13g2_decap_8 FILLER_70_1028 ();
 sg13g2_decap_4 FILLER_70_1035 ();
 sg13g2_fill_1 FILLER_70_1043 ();
 sg13g2_fill_2 FILLER_70_1091 ();
 sg13g2_decap_8 FILLER_70_1097 ();
 sg13g2_fill_1 FILLER_70_1104 ();
 sg13g2_fill_1 FILLER_70_1109 ();
 sg13g2_fill_1 FILLER_70_1136 ();
 sg13g2_fill_1 FILLER_70_1173 ();
 sg13g2_decap_8 FILLER_70_1178 ();
 sg13g2_decap_8 FILLER_70_1185 ();
 sg13g2_decap_8 FILLER_70_1192 ();
 sg13g2_fill_2 FILLER_70_1199 ();
 sg13g2_fill_2 FILLER_70_1226 ();
 sg13g2_fill_1 FILLER_70_1228 ();
 sg13g2_fill_2 FILLER_70_1243 ();
 sg13g2_decap_4 FILLER_70_1253 ();
 sg13g2_fill_2 FILLER_70_1257 ();
 sg13g2_fill_2 FILLER_70_1264 ();
 sg13g2_fill_1 FILLER_70_1266 ();
 sg13g2_fill_1 FILLER_70_1293 ();
 sg13g2_fill_1 FILLER_70_1304 ();
 sg13g2_decap_4 FILLER_70_1313 ();
 sg13g2_fill_1 FILLER_70_1317 ();
 sg13g2_decap_4 FILLER_70_1341 ();
 sg13g2_fill_1 FILLER_70_1350 ();
 sg13g2_decap_8 FILLER_70_1374 ();
 sg13g2_fill_1 FILLER_70_1381 ();
 sg13g2_decap_8 FILLER_70_1392 ();
 sg13g2_fill_2 FILLER_70_1399 ();
 sg13g2_decap_8 FILLER_70_1411 ();
 sg13g2_decap_8 FILLER_70_1418 ();
 sg13g2_decap_8 FILLER_70_1425 ();
 sg13g2_decap_8 FILLER_70_1432 ();
 sg13g2_decap_8 FILLER_70_1439 ();
 sg13g2_decap_8 FILLER_70_1451 ();
 sg13g2_decap_8 FILLER_70_1458 ();
 sg13g2_decap_8 FILLER_70_1465 ();
 sg13g2_decap_8 FILLER_70_1472 ();
 sg13g2_decap_4 FILLER_70_1479 ();
 sg13g2_fill_1 FILLER_70_1483 ();
 sg13g2_decap_4 FILLER_70_1488 ();
 sg13g2_fill_2 FILLER_70_1492 ();
 sg13g2_fill_1 FILLER_70_1539 ();
 sg13g2_fill_1 FILLER_70_1544 ();
 sg13g2_fill_2 FILLER_70_1548 ();
 sg13g2_fill_1 FILLER_70_1563 ();
 sg13g2_fill_2 FILLER_70_1568 ();
 sg13g2_fill_1 FILLER_70_1575 ();
 sg13g2_fill_2 FILLER_70_1582 ();
 sg13g2_decap_4 FILLER_70_1625 ();
 sg13g2_fill_1 FILLER_70_1629 ();
 sg13g2_fill_2 FILLER_70_1635 ();
 sg13g2_fill_2 FILLER_70_1641 ();
 sg13g2_fill_1 FILLER_70_1643 ();
 sg13g2_decap_4 FILLER_70_1658 ();
 sg13g2_decap_4 FILLER_70_1689 ();
 sg13g2_fill_1 FILLER_70_1693 ();
 sg13g2_fill_2 FILLER_70_1703 ();
 sg13g2_fill_1 FILLER_70_1705 ();
 sg13g2_fill_1 FILLER_70_1748 ();
 sg13g2_fill_1 FILLER_70_1763 ();
 sg13g2_decap_8 FILLER_70_1769 ();
 sg13g2_decap_8 FILLER_70_1776 ();
 sg13g2_fill_2 FILLER_70_1783 ();
 sg13g2_fill_1 FILLER_70_1785 ();
 sg13g2_fill_2 FILLER_70_1790 ();
 sg13g2_fill_1 FILLER_70_1792 ();
 sg13g2_fill_1 FILLER_70_1798 ();
 sg13g2_fill_1 FILLER_70_1818 ();
 sg13g2_fill_2 FILLER_70_1833 ();
 sg13g2_fill_1 FILLER_70_1835 ();
 sg13g2_fill_2 FILLER_70_1841 ();
 sg13g2_fill_1 FILLER_70_1843 ();
 sg13g2_fill_2 FILLER_70_1863 ();
 sg13g2_fill_1 FILLER_70_1865 ();
 sg13g2_fill_1 FILLER_70_1891 ();
 sg13g2_decap_8 FILLER_70_1897 ();
 sg13g2_decap_4 FILLER_70_1904 ();
 sg13g2_decap_4 FILLER_70_1913 ();
 sg13g2_fill_1 FILLER_70_1917 ();
 sg13g2_fill_1 FILLER_70_1950 ();
 sg13g2_decap_4 FILLER_70_1955 ();
 sg13g2_fill_2 FILLER_70_1959 ();
 sg13g2_fill_2 FILLER_70_1994 ();
 sg13g2_fill_2 FILLER_70_2004 ();
 sg13g2_decap_4 FILLER_70_2011 ();
 sg13g2_fill_1 FILLER_70_2023 ();
 sg13g2_decap_4 FILLER_70_2060 ();
 sg13g2_fill_1 FILLER_70_2064 ();
 sg13g2_decap_8 FILLER_70_2085 ();
 sg13g2_decap_4 FILLER_70_2102 ();
 sg13g2_decap_8 FILLER_70_2110 ();
 sg13g2_decap_4 FILLER_70_2117 ();
 sg13g2_fill_1 FILLER_70_2131 ();
 sg13g2_fill_1 FILLER_70_2136 ();
 sg13g2_fill_2 FILLER_70_2169 ();
 sg13g2_fill_1 FILLER_70_2171 ();
 sg13g2_fill_2 FILLER_70_2208 ();
 sg13g2_fill_2 FILLER_70_2259 ();
 sg13g2_fill_1 FILLER_70_2295 ();
 sg13g2_fill_2 FILLER_70_2310 ();
 sg13g2_fill_1 FILLER_70_2329 ();
 sg13g2_fill_2 FILLER_70_2356 ();
 sg13g2_fill_1 FILLER_70_2383 ();
 sg13g2_fill_2 FILLER_70_2457 ();
 sg13g2_fill_2 FILLER_70_2516 ();
 sg13g2_fill_1 FILLER_70_2518 ();
 sg13g2_fill_2 FILLER_70_2528 ();
 sg13g2_decap_4 FILLER_70_2570 ();
 sg13g2_fill_2 FILLER_70_2574 ();
 sg13g2_decap_8 FILLER_70_2612 ();
 sg13g2_decap_8 FILLER_70_2619 ();
 sg13g2_decap_8 FILLER_70_2626 ();
 sg13g2_decap_8 FILLER_70_2633 ();
 sg13g2_decap_8 FILLER_70_2640 ();
 sg13g2_decap_8 FILLER_70_2647 ();
 sg13g2_decap_8 FILLER_70_2654 ();
 sg13g2_decap_8 FILLER_70_2661 ();
 sg13g2_fill_2 FILLER_70_2668 ();
 sg13g2_fill_2 FILLER_71_0 ();
 sg13g2_decap_4 FILLER_71_64 ();
 sg13g2_fill_1 FILLER_71_129 ();
 sg13g2_fill_1 FILLER_71_146 ();
 sg13g2_fill_1 FILLER_71_158 ();
 sg13g2_decap_8 FILLER_71_181 ();
 sg13g2_decap_8 FILLER_71_188 ();
 sg13g2_fill_2 FILLER_71_195 ();
 sg13g2_fill_1 FILLER_71_218 ();
 sg13g2_decap_4 FILLER_71_224 ();
 sg13g2_decap_8 FILLER_71_232 ();
 sg13g2_decap_8 FILLER_71_265 ();
 sg13g2_decap_8 FILLER_71_285 ();
 sg13g2_decap_8 FILLER_71_292 ();
 sg13g2_decap_4 FILLER_71_299 ();
 sg13g2_fill_1 FILLER_71_303 ();
 sg13g2_decap_8 FILLER_71_330 ();
 sg13g2_fill_1 FILLER_71_351 ();
 sg13g2_fill_1 FILLER_71_361 ();
 sg13g2_fill_2 FILLER_71_366 ();
 sg13g2_fill_1 FILLER_71_368 ();
 sg13g2_decap_8 FILLER_71_376 ();
 sg13g2_decap_4 FILLER_71_383 ();
 sg13g2_decap_4 FILLER_71_392 ();
 sg13g2_fill_2 FILLER_71_396 ();
 sg13g2_fill_1 FILLER_71_401 ();
 sg13g2_decap_8 FILLER_71_432 ();
 sg13g2_decap_4 FILLER_71_439 ();
 sg13g2_fill_1 FILLER_71_443 ();
 sg13g2_fill_1 FILLER_71_457 ();
 sg13g2_fill_1 FILLER_71_467 ();
 sg13g2_fill_1 FILLER_71_472 ();
 sg13g2_fill_2 FILLER_71_481 ();
 sg13g2_fill_1 FILLER_71_483 ();
 sg13g2_decap_4 FILLER_71_488 ();
 sg13g2_fill_1 FILLER_71_492 ();
 sg13g2_fill_1 FILLER_71_506 ();
 sg13g2_fill_1 FILLER_71_525 ();
 sg13g2_decap_4 FILLER_71_531 ();
 sg13g2_fill_1 FILLER_71_535 ();
 sg13g2_fill_1 FILLER_71_596 ();
 sg13g2_fill_2 FILLER_71_602 ();
 sg13g2_fill_1 FILLER_71_604 ();
 sg13g2_decap_8 FILLER_71_608 ();
 sg13g2_fill_1 FILLER_71_615 ();
 sg13g2_fill_1 FILLER_71_646 ();
 sg13g2_fill_2 FILLER_71_673 ();
 sg13g2_fill_1 FILLER_71_684 ();
 sg13g2_fill_1 FILLER_71_731 ();
 sg13g2_decap_4 FILLER_71_758 ();
 sg13g2_fill_2 FILLER_71_762 ();
 sg13g2_fill_1 FILLER_71_768 ();
 sg13g2_decap_8 FILLER_71_774 ();
 sg13g2_fill_2 FILLER_71_788 ();
 sg13g2_fill_1 FILLER_71_818 ();
 sg13g2_fill_2 FILLER_71_823 ();
 sg13g2_fill_2 FILLER_71_831 ();
 sg13g2_decap_8 FILLER_71_837 ();
 sg13g2_fill_1 FILLER_71_844 ();
 sg13g2_fill_1 FILLER_71_854 ();
 sg13g2_fill_2 FILLER_71_871 ();
 sg13g2_fill_1 FILLER_71_873 ();
 sg13g2_fill_1 FILLER_71_900 ();
 sg13g2_decap_4 FILLER_71_910 ();
 sg13g2_decap_4 FILLER_71_924 ();
 sg13g2_fill_2 FILLER_71_928 ();
 sg13g2_fill_2 FILLER_71_935 ();
 sg13g2_fill_2 FILLER_71_941 ();
 sg13g2_fill_2 FILLER_71_953 ();
 sg13g2_fill_1 FILLER_71_999 ();
 sg13g2_decap_8 FILLER_71_1014 ();
 sg13g2_decap_8 FILLER_71_1021 ();
 sg13g2_decap_8 FILLER_71_1028 ();
 sg13g2_decap_8 FILLER_71_1061 ();
 sg13g2_decap_4 FILLER_71_1078 ();
 sg13g2_fill_2 FILLER_71_1082 ();
 sg13g2_fill_1 FILLER_71_1090 ();
 sg13g2_decap_8 FILLER_71_1101 ();
 sg13g2_decap_8 FILLER_71_1108 ();
 sg13g2_fill_2 FILLER_71_1123 ();
 sg13g2_fill_2 FILLER_71_1151 ();
 sg13g2_fill_1 FILLER_71_1153 ();
 sg13g2_decap_4 FILLER_71_1190 ();
 sg13g2_fill_1 FILLER_71_1194 ();
 sg13g2_fill_2 FILLER_71_1254 ();
 sg13g2_fill_2 FILLER_71_1301 ();
 sg13g2_fill_1 FILLER_71_1303 ();
 sg13g2_fill_1 FILLER_71_1314 ();
 sg13g2_fill_2 FILLER_71_1333 ();
 sg13g2_fill_1 FILLER_71_1335 ();
 sg13g2_fill_1 FILLER_71_1342 ();
 sg13g2_fill_2 FILLER_71_1349 ();
 sg13g2_fill_1 FILLER_71_1351 ();
 sg13g2_fill_1 FILLER_71_1359 ();
 sg13g2_decap_4 FILLER_71_1367 ();
 sg13g2_fill_2 FILLER_71_1398 ();
 sg13g2_decap_8 FILLER_71_1426 ();
 sg13g2_fill_2 FILLER_71_1443 ();
 sg13g2_decap_8 FILLER_71_1449 ();
 sg13g2_decap_8 FILLER_71_1456 ();
 sg13g2_decap_8 FILLER_71_1463 ();
 sg13g2_decap_4 FILLER_71_1470 ();
 sg13g2_fill_2 FILLER_71_1474 ();
 sg13g2_fill_1 FILLER_71_1512 ();
 sg13g2_fill_2 FILLER_71_1521 ();
 sg13g2_fill_2 FILLER_71_1539 ();
 sg13g2_fill_1 FILLER_71_1561 ();
 sg13g2_fill_1 FILLER_71_1574 ();
 sg13g2_fill_2 FILLER_71_1583 ();
 sg13g2_fill_2 FILLER_71_1590 ();
 sg13g2_fill_2 FILLER_71_1597 ();
 sg13g2_fill_2 FILLER_71_1609 ();
 sg13g2_fill_1 FILLER_71_1611 ();
 sg13g2_fill_1 FILLER_71_1632 ();
 sg13g2_decap_4 FILLER_71_1654 ();
 sg13g2_fill_1 FILLER_71_1658 ();
 sg13g2_fill_2 FILLER_71_1667 ();
 sg13g2_decap_8 FILLER_71_1675 ();
 sg13g2_decap_8 FILLER_71_1682 ();
 sg13g2_decap_8 FILLER_71_1689 ();
 sg13g2_decap_8 FILLER_71_1696 ();
 sg13g2_fill_2 FILLER_71_1707 ();
 sg13g2_fill_1 FILLER_71_1713 ();
 sg13g2_fill_2 FILLER_71_1739 ();
 sg13g2_fill_1 FILLER_71_1741 ();
 sg13g2_fill_1 FILLER_71_1754 ();
 sg13g2_decap_4 FILLER_71_1760 ();
 sg13g2_fill_2 FILLER_71_1773 ();
 sg13g2_decap_4 FILLER_71_1781 ();
 sg13g2_fill_1 FILLER_71_1790 ();
 sg13g2_fill_2 FILLER_71_1800 ();
 sg13g2_decap_4 FILLER_71_1822 ();
 sg13g2_fill_1 FILLER_71_1847 ();
 sg13g2_fill_1 FILLER_71_1863 ();
 sg13g2_fill_2 FILLER_71_1896 ();
 sg13g2_fill_1 FILLER_71_1902 ();
 sg13g2_decap_8 FILLER_71_1907 ();
 sg13g2_decap_4 FILLER_71_1914 ();
 sg13g2_fill_1 FILLER_71_1918 ();
 sg13g2_fill_2 FILLER_71_1941 ();
 sg13g2_fill_2 FILLER_71_1961 ();
 sg13g2_fill_1 FILLER_71_1988 ();
 sg13g2_fill_1 FILLER_71_2005 ();
 sg13g2_decap_8 FILLER_71_2011 ();
 sg13g2_decap_8 FILLER_71_2018 ();
 sg13g2_decap_8 FILLER_71_2025 ();
 sg13g2_decap_4 FILLER_71_2032 ();
 sg13g2_fill_2 FILLER_71_2036 ();
 sg13g2_fill_2 FILLER_71_2068 ();
 sg13g2_fill_1 FILLER_71_2070 ();
 sg13g2_fill_1 FILLER_71_2076 ();
 sg13g2_fill_1 FILLER_71_2111 ();
 sg13g2_fill_2 FILLER_71_2138 ();
 sg13g2_fill_1 FILLER_71_2140 ();
 sg13g2_fill_1 FILLER_71_2172 ();
 sg13g2_fill_2 FILLER_71_2177 ();
 sg13g2_fill_2 FILLER_71_2243 ();
 sg13g2_fill_1 FILLER_71_2245 ();
 sg13g2_fill_2 FILLER_71_2266 ();
 sg13g2_fill_2 FILLER_71_2272 ();
 sg13g2_fill_2 FILLER_71_2285 ();
 sg13g2_fill_1 FILLER_71_2314 ();
 sg13g2_fill_1 FILLER_71_2320 ();
 sg13g2_fill_1 FILLER_71_2341 ();
 sg13g2_fill_2 FILLER_71_2352 ();
 sg13g2_fill_1 FILLER_71_2373 ();
 sg13g2_fill_1 FILLER_71_2382 ();
 sg13g2_fill_1 FILLER_71_2398 ();
 sg13g2_decap_4 FILLER_71_2403 ();
 sg13g2_fill_2 FILLER_71_2447 ();
 sg13g2_decap_8 FILLER_71_2496 ();
 sg13g2_decap_8 FILLER_71_2503 ();
 sg13g2_decap_4 FILLER_71_2510 ();
 sg13g2_fill_1 FILLER_71_2514 ();
 sg13g2_fill_1 FILLER_71_2538 ();
 sg13g2_decap_8 FILLER_71_2565 ();
 sg13g2_decap_8 FILLER_71_2572 ();
 sg13g2_decap_8 FILLER_71_2579 ();
 sg13g2_decap_8 FILLER_71_2586 ();
 sg13g2_decap_8 FILLER_71_2597 ();
 sg13g2_decap_8 FILLER_71_2604 ();
 sg13g2_decap_8 FILLER_71_2611 ();
 sg13g2_decap_8 FILLER_71_2618 ();
 sg13g2_decap_8 FILLER_71_2625 ();
 sg13g2_decap_8 FILLER_71_2632 ();
 sg13g2_decap_8 FILLER_71_2639 ();
 sg13g2_decap_8 FILLER_71_2646 ();
 sg13g2_decap_8 FILLER_71_2653 ();
 sg13g2_decap_8 FILLER_71_2660 ();
 sg13g2_fill_2 FILLER_71_2667 ();
 sg13g2_fill_1 FILLER_71_2669 ();
 sg13g2_decap_8 FILLER_72_0 ();
 sg13g2_fill_2 FILLER_72_7 ();
 sg13g2_fill_2 FILLER_72_17 ();
 sg13g2_fill_1 FILLER_72_19 ();
 sg13g2_decap_4 FILLER_72_30 ();
 sg13g2_fill_2 FILLER_72_34 ();
 sg13g2_fill_2 FILLER_72_41 ();
 sg13g2_fill_1 FILLER_72_43 ();
 sg13g2_fill_2 FILLER_72_49 ();
 sg13g2_decap_8 FILLER_72_61 ();
 sg13g2_decap_4 FILLER_72_68 ();
 sg13g2_fill_2 FILLER_72_72 ();
 sg13g2_decap_8 FILLER_72_78 ();
 sg13g2_decap_8 FILLER_72_85 ();
 sg13g2_decap_8 FILLER_72_92 ();
 sg13g2_decap_4 FILLER_72_99 ();
 sg13g2_fill_2 FILLER_72_156 ();
 sg13g2_fill_2 FILLER_72_167 ();
 sg13g2_fill_2 FILLER_72_198 ();
 sg13g2_fill_1 FILLER_72_200 ();
 sg13g2_fill_1 FILLER_72_210 ();
 sg13g2_decap_4 FILLER_72_216 ();
 sg13g2_decap_4 FILLER_72_241 ();
 sg13g2_fill_1 FILLER_72_245 ();
 sg13g2_decap_8 FILLER_72_251 ();
 sg13g2_decap_8 FILLER_72_258 ();
 sg13g2_fill_2 FILLER_72_265 ();
 sg13g2_fill_1 FILLER_72_267 ();
 sg13g2_fill_1 FILLER_72_302 ();
 sg13g2_decap_4 FILLER_72_307 ();
 sg13g2_decap_8 FILLER_72_315 ();
 sg13g2_fill_2 FILLER_72_322 ();
 sg13g2_fill_2 FILLER_72_350 ();
 sg13g2_fill_2 FILLER_72_391 ();
 sg13g2_fill_1 FILLER_72_393 ();
 sg13g2_decap_8 FILLER_72_403 ();
 sg13g2_fill_2 FILLER_72_410 ();
 sg13g2_fill_1 FILLER_72_412 ();
 sg13g2_decap_8 FILLER_72_417 ();
 sg13g2_decap_8 FILLER_72_424 ();
 sg13g2_decap_8 FILLER_72_431 ();
 sg13g2_fill_1 FILLER_72_438 ();
 sg13g2_fill_1 FILLER_72_472 ();
 sg13g2_fill_2 FILLER_72_476 ();
 sg13g2_fill_1 FILLER_72_478 ();
 sg13g2_fill_1 FILLER_72_498 ();
 sg13g2_decap_4 FILLER_72_525 ();
 sg13g2_fill_2 FILLER_72_529 ();
 sg13g2_decap_4 FILLER_72_543 ();
 sg13g2_fill_1 FILLER_72_551 ();
 sg13g2_fill_1 FILLER_72_558 ();
 sg13g2_fill_2 FILLER_72_565 ();
 sg13g2_fill_1 FILLER_72_567 ();
 sg13g2_fill_1 FILLER_72_631 ();
 sg13g2_fill_1 FILLER_72_636 ();
 sg13g2_decap_4 FILLER_72_642 ();
 sg13g2_fill_1 FILLER_72_646 ();
 sg13g2_decap_8 FILLER_72_707 ();
 sg13g2_decap_8 FILLER_72_718 ();
 sg13g2_fill_1 FILLER_72_725 ();
 sg13g2_decap_4 FILLER_72_731 ();
 sg13g2_fill_2 FILLER_72_735 ();
 sg13g2_decap_4 FILLER_72_741 ();
 sg13g2_fill_2 FILLER_72_745 ();
 sg13g2_fill_1 FILLER_72_799 ();
 sg13g2_decap_8 FILLER_72_806 ();
 sg13g2_fill_1 FILLER_72_813 ();
 sg13g2_fill_1 FILLER_72_820 ();
 sg13g2_decap_8 FILLER_72_824 ();
 sg13g2_fill_1 FILLER_72_842 ();
 sg13g2_decap_4 FILLER_72_907 ();
 sg13g2_fill_1 FILLER_72_937 ();
 sg13g2_fill_2 FILLER_72_967 ();
 sg13g2_decap_4 FILLER_72_995 ();
 sg13g2_fill_1 FILLER_72_1025 ();
 sg13g2_fill_2 FILLER_72_1052 ();
 sg13g2_fill_1 FILLER_72_1080 ();
 sg13g2_fill_2 FILLER_72_1107 ();
 sg13g2_decap_4 FILLER_72_1135 ();
 sg13g2_fill_2 FILLER_72_1139 ();
 sg13g2_fill_1 FILLER_72_1168 ();
 sg13g2_decap_4 FILLER_72_1195 ();
 sg13g2_fill_1 FILLER_72_1241 ();
 sg13g2_decap_4 FILLER_72_1247 ();
 sg13g2_fill_1 FILLER_72_1251 ();
 sg13g2_fill_2 FILLER_72_1257 ();
 sg13g2_fill_2 FILLER_72_1264 ();
 sg13g2_fill_1 FILLER_72_1266 ();
 sg13g2_fill_2 FILLER_72_1283 ();
 sg13g2_fill_1 FILLER_72_1285 ();
 sg13g2_decap_4 FILLER_72_1295 ();
 sg13g2_decap_8 FILLER_72_1319 ();
 sg13g2_fill_2 FILLER_72_1326 ();
 sg13g2_fill_2 FILLER_72_1336 ();
 sg13g2_decap_4 FILLER_72_1342 ();
 sg13g2_fill_2 FILLER_72_1366 ();
 sg13g2_fill_1 FILLER_72_1368 ();
 sg13g2_fill_2 FILLER_72_1382 ();
 sg13g2_fill_1 FILLER_72_1384 ();
 sg13g2_decap_8 FILLER_72_1426 ();
 sg13g2_fill_1 FILLER_72_1433 ();
 sg13g2_decap_4 FILLER_72_1460 ();
 sg13g2_fill_2 FILLER_72_1464 ();
 sg13g2_fill_1 FILLER_72_1517 ();
 sg13g2_fill_2 FILLER_72_1541 ();
 sg13g2_fill_1 FILLER_72_1553 ();
 sg13g2_decap_4 FILLER_72_1558 ();
 sg13g2_fill_2 FILLER_72_1575 ();
 sg13g2_fill_2 FILLER_72_1606 ();
 sg13g2_fill_1 FILLER_72_1608 ();
 sg13g2_decap_4 FILLER_72_1638 ();
 sg13g2_fill_2 FILLER_72_1642 ();
 sg13g2_decap_8 FILLER_72_1654 ();
 sg13g2_decap_4 FILLER_72_1661 ();
 sg13g2_fill_1 FILLER_72_1665 ();
 sg13g2_decap_8 FILLER_72_1672 ();
 sg13g2_decap_8 FILLER_72_1679 ();
 sg13g2_decap_8 FILLER_72_1686 ();
 sg13g2_decap_8 FILLER_72_1693 ();
 sg13g2_fill_2 FILLER_72_1700 ();
 sg13g2_fill_1 FILLER_72_1716 ();
 sg13g2_fill_1 FILLER_72_1726 ();
 sg13g2_fill_2 FILLER_72_1755 ();
 sg13g2_fill_1 FILLER_72_1757 ();
 sg13g2_fill_1 FILLER_72_1763 ();
 sg13g2_fill_2 FILLER_72_1768 ();
 sg13g2_fill_1 FILLER_72_1770 ();
 sg13g2_fill_1 FILLER_72_1786 ();
 sg13g2_fill_2 FILLER_72_1795 ();
 sg13g2_decap_4 FILLER_72_1810 ();
 sg13g2_fill_1 FILLER_72_1821 ();
 sg13g2_fill_1 FILLER_72_1827 ();
 sg13g2_fill_2 FILLER_72_1844 ();
 sg13g2_fill_1 FILLER_72_1846 ();
 sg13g2_fill_2 FILLER_72_1888 ();
 sg13g2_decap_8 FILLER_72_1915 ();
 sg13g2_decap_8 FILLER_72_1922 ();
 sg13g2_decap_4 FILLER_72_1929 ();
 sg13g2_decap_4 FILLER_72_1937 ();
 sg13g2_fill_2 FILLER_72_1941 ();
 sg13g2_decap_4 FILLER_72_1968 ();
 sg13g2_fill_2 FILLER_72_1976 ();
 sg13g2_fill_1 FILLER_72_1978 ();
 sg13g2_decap_8 FILLER_72_1984 ();
 sg13g2_decap_8 FILLER_72_1991 ();
 sg13g2_decap_8 FILLER_72_1998 ();
 sg13g2_decap_8 FILLER_72_2005 ();
 sg13g2_decap_8 FILLER_72_2012 ();
 sg13g2_decap_4 FILLER_72_2019 ();
 sg13g2_fill_1 FILLER_72_2023 ();
 sg13g2_decap_4 FILLER_72_2060 ();
 sg13g2_fill_2 FILLER_72_2064 ();
 sg13g2_fill_1 FILLER_72_2127 ();
 sg13g2_fill_2 FILLER_72_2132 ();
 sg13g2_fill_1 FILLER_72_2138 ();
 sg13g2_fill_2 FILLER_72_2160 ();
 sg13g2_fill_1 FILLER_72_2175 ();
 sg13g2_fill_1 FILLER_72_2189 ();
 sg13g2_fill_1 FILLER_72_2206 ();
 sg13g2_decap_4 FILLER_72_2220 ();
 sg13g2_fill_2 FILLER_72_2224 ();
 sg13g2_fill_1 FILLER_72_2372 ();
 sg13g2_fill_2 FILLER_72_2382 ();
 sg13g2_fill_1 FILLER_72_2388 ();
 sg13g2_decap_8 FILLER_72_2395 ();
 sg13g2_decap_4 FILLER_72_2402 ();
 sg13g2_fill_1 FILLER_72_2406 ();
 sg13g2_fill_2 FILLER_72_2417 ();
 sg13g2_fill_1 FILLER_72_2432 ();
 sg13g2_fill_2 FILLER_72_2463 ();
 sg13g2_fill_1 FILLER_72_2470 ();
 sg13g2_fill_1 FILLER_72_2555 ();
 sg13g2_decap_8 FILLER_72_2582 ();
 sg13g2_decap_8 FILLER_72_2589 ();
 sg13g2_decap_8 FILLER_72_2596 ();
 sg13g2_decap_8 FILLER_72_2603 ();
 sg13g2_decap_8 FILLER_72_2610 ();
 sg13g2_decap_8 FILLER_72_2617 ();
 sg13g2_decap_8 FILLER_72_2624 ();
 sg13g2_decap_8 FILLER_72_2631 ();
 sg13g2_decap_8 FILLER_72_2638 ();
 sg13g2_decap_8 FILLER_72_2645 ();
 sg13g2_decap_8 FILLER_72_2652 ();
 sg13g2_decap_8 FILLER_72_2659 ();
 sg13g2_decap_4 FILLER_72_2666 ();
 sg13g2_decap_4 FILLER_73_0 ();
 sg13g2_fill_2 FILLER_73_35 ();
 sg13g2_fill_1 FILLER_73_37 ();
 sg13g2_fill_2 FILLER_73_46 ();
 sg13g2_fill_2 FILLER_73_53 ();
 sg13g2_decap_4 FILLER_73_72 ();
 sg13g2_fill_2 FILLER_73_76 ();
 sg13g2_fill_2 FILLER_73_108 ();
 sg13g2_fill_1 FILLER_73_163 ();
 sg13g2_fill_1 FILLER_73_168 ();
 sg13g2_decap_4 FILLER_73_214 ();
 sg13g2_fill_1 FILLER_73_290 ();
 sg13g2_decap_8 FILLER_73_326 ();
 sg13g2_decap_8 FILLER_73_337 ();
 sg13g2_decap_8 FILLER_73_344 ();
 sg13g2_fill_1 FILLER_73_351 ();
 sg13g2_fill_1 FILLER_73_361 ();
 sg13g2_fill_1 FILLER_73_388 ();
 sg13g2_fill_1 FILLER_73_394 ();
 sg13g2_decap_4 FILLER_73_425 ();
 sg13g2_fill_2 FILLER_73_463 ();
 sg13g2_decap_4 FILLER_73_557 ();
 sg13g2_fill_2 FILLER_73_586 ();
 sg13g2_fill_2 FILLER_73_597 ();
 sg13g2_fill_1 FILLER_73_599 ();
 sg13g2_fill_1 FILLER_73_604 ();
 sg13g2_decap_8 FILLER_73_636 ();
 sg13g2_decap_8 FILLER_73_643 ();
 sg13g2_decap_8 FILLER_73_650 ();
 sg13g2_fill_2 FILLER_73_657 ();
 sg13g2_decap_4 FILLER_73_663 ();
 sg13g2_fill_2 FILLER_73_667 ();
 sg13g2_decap_8 FILLER_73_709 ();
 sg13g2_decap_8 FILLER_73_716 ();
 sg13g2_decap_4 FILLER_73_723 ();
 sg13g2_fill_2 FILLER_73_727 ();
 sg13g2_fill_1 FILLER_73_764 ();
 sg13g2_decap_4 FILLER_73_770 ();
 sg13g2_fill_1 FILLER_73_774 ();
 sg13g2_decap_8 FILLER_73_805 ();
 sg13g2_fill_2 FILLER_73_812 ();
 sg13g2_fill_1 FILLER_73_814 ();
 sg13g2_decap_4 FILLER_73_825 ();
 sg13g2_fill_1 FILLER_73_855 ();
 sg13g2_fill_2 FILLER_73_861 ();
 sg13g2_fill_1 FILLER_73_889 ();
 sg13g2_fill_2 FILLER_73_916 ();
 sg13g2_fill_2 FILLER_73_948 ();
 sg13g2_fill_1 FILLER_73_950 ();
 sg13g2_fill_2 FILLER_73_979 ();
 sg13g2_decap_8 FILLER_73_985 ();
 sg13g2_fill_2 FILLER_73_992 ();
 sg13g2_fill_1 FILLER_73_994 ();
 sg13g2_decap_4 FILLER_73_1027 ();
 sg13g2_fill_2 FILLER_73_1031 ();
 sg13g2_fill_1 FILLER_73_1059 ();
 sg13g2_fill_1 FILLER_73_1067 ();
 sg13g2_fill_2 FILLER_73_1074 ();
 sg13g2_fill_1 FILLER_73_1086 ();
 sg13g2_fill_1 FILLER_73_1095 ();
 sg13g2_fill_2 FILLER_73_1199 ();
 sg13g2_fill_1 FILLER_73_1211 ();
 sg13g2_fill_1 FILLER_73_1217 ();
 sg13g2_fill_1 FILLER_73_1223 ();
 sg13g2_fill_1 FILLER_73_1240 ();
 sg13g2_decap_4 FILLER_73_1262 ();
 sg13g2_decap_8 FILLER_73_1276 ();
 sg13g2_fill_2 FILLER_73_1314 ();
 sg13g2_fill_1 FILLER_73_1316 ();
 sg13g2_fill_2 FILLER_73_1329 ();
 sg13g2_fill_1 FILLER_73_1331 ();
 sg13g2_decap_4 FILLER_73_1337 ();
 sg13g2_fill_1 FILLER_73_1346 ();
 sg13g2_fill_2 FILLER_73_1357 ();
 sg13g2_decap_8 FILLER_73_1372 ();
 sg13g2_fill_2 FILLER_73_1387 ();
 sg13g2_fill_1 FILLER_73_1465 ();
 sg13g2_fill_2 FILLER_73_1504 ();
 sg13g2_fill_1 FILLER_73_1517 ();
 sg13g2_fill_1 FILLER_73_1552 ();
 sg13g2_decap_8 FILLER_73_1598 ();
 sg13g2_fill_1 FILLER_73_1605 ();
 sg13g2_fill_1 FILLER_73_1616 ();
 sg13g2_decap_8 FILLER_73_1625 ();
 sg13g2_fill_2 FILLER_73_1632 ();
 sg13g2_fill_2 FILLER_73_1639 ();
 sg13g2_fill_1 FILLER_73_1645 ();
 sg13g2_decap_4 FILLER_73_1659 ();
 sg13g2_fill_1 FILLER_73_1663 ();
 sg13g2_fill_2 FILLER_73_1669 ();
 sg13g2_fill_1 FILLER_73_1671 ();
 sg13g2_fill_1 FILLER_73_1689 ();
 sg13g2_fill_2 FILLER_73_1716 ();
 sg13g2_fill_1 FILLER_73_1718 ();
 sg13g2_fill_2 FILLER_73_1736 ();
 sg13g2_fill_1 FILLER_73_1762 ();
 sg13g2_fill_1 FILLER_73_1773 ();
 sg13g2_fill_1 FILLER_73_1782 ();
 sg13g2_decap_4 FILLER_73_1788 ();
 sg13g2_fill_1 FILLER_73_1792 ();
 sg13g2_fill_2 FILLER_73_1798 ();
 sg13g2_fill_1 FILLER_73_1800 ();
 sg13g2_decap_4 FILLER_73_1806 ();
 sg13g2_fill_1 FILLER_73_1810 ();
 sg13g2_fill_1 FILLER_73_1835 ();
 sg13g2_fill_1 FILLER_73_1878 ();
 sg13g2_fill_2 FILLER_73_1909 ();
 sg13g2_fill_1 FILLER_73_1911 ();
 sg13g2_decap_4 FILLER_73_1919 ();
 sg13g2_fill_2 FILLER_73_1954 ();
 sg13g2_decap_8 FILLER_73_1969 ();
 sg13g2_decap_8 FILLER_73_1976 ();
 sg13g2_decap_8 FILLER_73_1983 ();
 sg13g2_decap_8 FILLER_73_1990 ();
 sg13g2_decap_8 FILLER_73_1997 ();
 sg13g2_decap_8 FILLER_73_2004 ();
 sg13g2_fill_1 FILLER_73_2011 ();
 sg13g2_fill_1 FILLER_73_2033 ();
 sg13g2_fill_2 FILLER_73_2038 ();
 sg13g2_fill_1 FILLER_73_2040 ();
 sg13g2_fill_2 FILLER_73_2049 ();
 sg13g2_decap_8 FILLER_73_2061 ();
 sg13g2_fill_1 FILLER_73_2128 ();
 sg13g2_decap_4 FILLER_73_2185 ();
 sg13g2_fill_1 FILLER_73_2189 ();
 sg13g2_decap_4 FILLER_73_2240 ();
 sg13g2_fill_1 FILLER_73_2244 ();
 sg13g2_fill_1 FILLER_73_2324 ();
 sg13g2_decap_4 FILLER_73_2364 ();
 sg13g2_decap_8 FILLER_73_2398 ();
 sg13g2_decap_8 FILLER_73_2405 ();
 sg13g2_decap_4 FILLER_73_2412 ();
 sg13g2_fill_1 FILLER_73_2416 ();
 sg13g2_fill_1 FILLER_73_2422 ();
 sg13g2_fill_1 FILLER_73_2452 ();
 sg13g2_decap_4 FILLER_73_2486 ();
 sg13g2_fill_1 FILLER_73_2490 ();
 sg13g2_fill_1 FILLER_73_2496 ();
 sg13g2_fill_1 FILLER_73_2501 ();
 sg13g2_fill_1 FILLER_73_2508 ();
 sg13g2_fill_1 FILLER_73_2513 ();
 sg13g2_fill_1 FILLER_73_2525 ();
 sg13g2_fill_1 FILLER_73_2541 ();
 sg13g2_decap_8 FILLER_73_2585 ();
 sg13g2_decap_8 FILLER_73_2592 ();
 sg13g2_decap_8 FILLER_73_2599 ();
 sg13g2_decap_8 FILLER_73_2606 ();
 sg13g2_decap_8 FILLER_73_2613 ();
 sg13g2_decap_8 FILLER_73_2620 ();
 sg13g2_decap_8 FILLER_73_2627 ();
 sg13g2_decap_8 FILLER_73_2634 ();
 sg13g2_decap_8 FILLER_73_2641 ();
 sg13g2_decap_8 FILLER_73_2648 ();
 sg13g2_decap_8 FILLER_73_2655 ();
 sg13g2_decap_8 FILLER_73_2662 ();
 sg13g2_fill_1 FILLER_73_2669 ();
 sg13g2_decap_8 FILLER_74_0 ();
 sg13g2_decap_8 FILLER_74_7 ();
 sg13g2_decap_8 FILLER_74_14 ();
 sg13g2_decap_8 FILLER_74_21 ();
 sg13g2_decap_4 FILLER_74_28 ();
 sg13g2_fill_1 FILLER_74_36 ();
 sg13g2_fill_2 FILLER_74_119 ();
 sg13g2_fill_1 FILLER_74_134 ();
 sg13g2_fill_1 FILLER_74_150 ();
 sg13g2_fill_2 FILLER_74_203 ();
 sg13g2_fill_1 FILLER_74_205 ();
 sg13g2_fill_2 FILLER_74_216 ();
 sg13g2_decap_8 FILLER_74_253 ();
 sg13g2_fill_2 FILLER_74_260 ();
 sg13g2_fill_2 FILLER_74_283 ();
 sg13g2_fill_1 FILLER_74_285 ();
 sg13g2_fill_1 FILLER_74_318 ();
 sg13g2_decap_8 FILLER_74_323 ();
 sg13g2_fill_2 FILLER_74_330 ();
 sg13g2_fill_1 FILLER_74_335 ();
 sg13g2_decap_4 FILLER_74_339 ();
 sg13g2_fill_1 FILLER_74_343 ();
 sg13g2_fill_2 FILLER_74_349 ();
 sg13g2_fill_1 FILLER_74_351 ();
 sg13g2_fill_1 FILLER_74_361 ();
 sg13g2_decap_4 FILLER_74_423 ();
 sg13g2_fill_2 FILLER_74_467 ();
 sg13g2_decap_8 FILLER_74_514 ();
 sg13g2_fill_2 FILLER_74_521 ();
 sg13g2_fill_1 FILLER_74_523 ();
 sg13g2_fill_2 FILLER_74_528 ();
 sg13g2_fill_1 FILLER_74_530 ();
 sg13g2_fill_2 FILLER_74_536 ();
 sg13g2_fill_1 FILLER_74_538 ();
 sg13g2_fill_1 FILLER_74_548 ();
 sg13g2_decap_4 FILLER_74_553 ();
 sg13g2_fill_1 FILLER_74_557 ();
 sg13g2_fill_2 FILLER_74_574 ();
 sg13g2_fill_1 FILLER_74_576 ();
 sg13g2_fill_1 FILLER_74_586 ();
 sg13g2_fill_2 FILLER_74_600 ();
 sg13g2_fill_2 FILLER_74_613 ();
 sg13g2_fill_2 FILLER_74_644 ();
 sg13g2_decap_4 FILLER_74_672 ();
 sg13g2_decap_8 FILLER_74_690 ();
 sg13g2_fill_2 FILLER_74_759 ();
 sg13g2_fill_2 FILLER_74_837 ();
 sg13g2_decap_8 FILLER_74_884 ();
 sg13g2_decap_4 FILLER_74_891 ();
 sg13g2_fill_1 FILLER_74_895 ();
 sg13g2_decap_4 FILLER_74_900 ();
 sg13g2_fill_1 FILLER_74_904 ();
 sg13g2_fill_2 FILLER_74_915 ();
 sg13g2_fill_2 FILLER_74_927 ();
 sg13g2_fill_1 FILLER_74_929 ();
 sg13g2_fill_2 FILLER_74_934 ();
 sg13g2_fill_1 FILLER_74_936 ();
 sg13g2_fill_1 FILLER_74_947 ();
 sg13g2_fill_2 FILLER_74_952 ();
 sg13g2_fill_1 FILLER_74_979 ();
 sg13g2_decap_8 FILLER_74_984 ();
 sg13g2_decap_4 FILLER_74_991 ();
 sg13g2_fill_2 FILLER_74_995 ();
 sg13g2_fill_1 FILLER_74_1011 ();
 sg13g2_fill_2 FILLER_74_1039 ();
 sg13g2_fill_2 FILLER_74_1049 ();
 sg13g2_fill_1 FILLER_74_1070 ();
 sg13g2_fill_2 FILLER_74_1075 ();
 sg13g2_decap_8 FILLER_74_1113 ();
 sg13g2_decap_8 FILLER_74_1120 ();
 sg13g2_fill_1 FILLER_74_1127 ();
 sg13g2_fill_2 FILLER_74_1138 ();
 sg13g2_fill_1 FILLER_74_1176 ();
 sg13g2_decap_8 FILLER_74_1195 ();
 sg13g2_fill_2 FILLER_74_1217 ();
 sg13g2_fill_1 FILLER_74_1219 ();
 sg13g2_decap_4 FILLER_74_1225 ();
 sg13g2_fill_1 FILLER_74_1229 ();
 sg13g2_fill_2 FILLER_74_1235 ();
 sg13g2_fill_1 FILLER_74_1237 ();
 sg13g2_decap_4 FILLER_74_1243 ();
 sg13g2_fill_2 FILLER_74_1268 ();
 sg13g2_decap_8 FILLER_74_1276 ();
 sg13g2_decap_8 FILLER_74_1283 ();
 sg13g2_decap_8 FILLER_74_1290 ();
 sg13g2_fill_2 FILLER_74_1297 ();
 sg13g2_decap_8 FILLER_74_1306 ();
 sg13g2_decap_4 FILLER_74_1313 ();
 sg13g2_decap_8 FILLER_74_1326 ();
 sg13g2_decap_8 FILLER_74_1333 ();
 sg13g2_fill_1 FILLER_74_1353 ();
 sg13g2_fill_2 FILLER_74_1369 ();
 sg13g2_fill_2 FILLER_74_1411 ();
 sg13g2_decap_4 FILLER_74_1417 ();
 sg13g2_decap_8 FILLER_74_1426 ();
 sg13g2_fill_1 FILLER_74_1433 ();
 sg13g2_fill_2 FILLER_74_1470 ();
 sg13g2_fill_1 FILLER_74_1472 ();
 sg13g2_fill_2 FILLER_74_1477 ();
 sg13g2_fill_1 FILLER_74_1495 ();
 sg13g2_fill_1 FILLER_74_1517 ();
 sg13g2_fill_2 FILLER_74_1539 ();
 sg13g2_decap_8 FILLER_74_1551 ();
 sg13g2_fill_1 FILLER_74_1558 ();
 sg13g2_decap_8 FILLER_74_1563 ();
 sg13g2_decap_4 FILLER_74_1570 ();
 sg13g2_fill_2 FILLER_74_1589 ();
 sg13g2_decap_8 FILLER_74_1600 ();
 sg13g2_fill_2 FILLER_74_1607 ();
 sg13g2_decap_4 FILLER_74_1613 ();
 sg13g2_fill_2 FILLER_74_1617 ();
 sg13g2_fill_2 FILLER_74_1624 ();
 sg13g2_fill_1 FILLER_74_1626 ();
 sg13g2_fill_2 FILLER_74_1631 ();
 sg13g2_fill_1 FILLER_74_1633 ();
 sg13g2_fill_2 FILLER_74_1638 ();
 sg13g2_decap_4 FILLER_74_1653 ();
 sg13g2_fill_2 FILLER_74_1657 ();
 sg13g2_decap_4 FILLER_74_1664 ();
 sg13g2_fill_1 FILLER_74_1668 ();
 sg13g2_fill_2 FILLER_74_1679 ();
 sg13g2_fill_1 FILLER_74_1681 ();
 sg13g2_decap_4 FILLER_74_1686 ();
 sg13g2_fill_2 FILLER_74_1693 ();
 sg13g2_fill_1 FILLER_74_1695 ();
 sg13g2_fill_2 FILLER_74_1700 ();
 sg13g2_fill_2 FILLER_74_1710 ();
 sg13g2_fill_1 FILLER_74_1712 ();
 sg13g2_fill_2 FILLER_74_1717 ();
 sg13g2_fill_1 FILLER_74_1719 ();
 sg13g2_fill_2 FILLER_74_1735 ();
 sg13g2_fill_1 FILLER_74_1737 ();
 sg13g2_fill_2 FILLER_74_1741 ();
 sg13g2_fill_1 FILLER_74_1748 ();
 sg13g2_fill_2 FILLER_74_1753 ();
 sg13g2_fill_1 FILLER_74_1755 ();
 sg13g2_fill_2 FILLER_74_1761 ();
 sg13g2_fill_1 FILLER_74_1763 ();
 sg13g2_decap_8 FILLER_74_1772 ();
 sg13g2_decap_8 FILLER_74_1779 ();
 sg13g2_fill_2 FILLER_74_1786 ();
 sg13g2_fill_1 FILLER_74_1788 ();
 sg13g2_fill_2 FILLER_74_1825 ();
 sg13g2_fill_1 FILLER_74_1827 ();
 sg13g2_fill_1 FILLER_74_1837 ();
 sg13g2_decap_8 FILLER_74_1850 ();
 sg13g2_fill_2 FILLER_74_1873 ();
 sg13g2_decap_4 FILLER_74_1900 ();
 sg13g2_fill_1 FILLER_74_1904 ();
 sg13g2_decap_8 FILLER_74_1909 ();
 sg13g2_fill_1 FILLER_74_1916 ();
 sg13g2_fill_1 FILLER_74_1947 ();
 sg13g2_decap_8 FILLER_74_1966 ();
 sg13g2_decap_8 FILLER_74_1973 ();
 sg13g2_decap_8 FILLER_74_1980 ();
 sg13g2_decap_4 FILLER_74_1987 ();
 sg13g2_fill_1 FILLER_74_1991 ();
 sg13g2_fill_1 FILLER_74_2018 ();
 sg13g2_decap_8 FILLER_74_2049 ();
 sg13g2_decap_8 FILLER_74_2056 ();
 sg13g2_decap_4 FILLER_74_2063 ();
 sg13g2_fill_1 FILLER_74_2067 ();
 sg13g2_decap_4 FILLER_74_2078 ();
 sg13g2_fill_1 FILLER_74_2082 ();
 sg13g2_decap_4 FILLER_74_2087 ();
 sg13g2_fill_1 FILLER_74_2091 ();
 sg13g2_decap_4 FILLER_74_2098 ();
 sg13g2_decap_8 FILLER_74_2121 ();
 sg13g2_decap_8 FILLER_74_2128 ();
 sg13g2_fill_1 FILLER_74_2135 ();
 sg13g2_fill_2 FILLER_74_2146 ();
 sg13g2_fill_1 FILLER_74_2148 ();
 sg13g2_decap_8 FILLER_74_2167 ();
 sg13g2_decap_4 FILLER_74_2174 ();
 sg13g2_fill_2 FILLER_74_2214 ();
 sg13g2_fill_1 FILLER_74_2216 ();
 sg13g2_decap_8 FILLER_74_2227 ();
 sg13g2_decap_8 FILLER_74_2234 ();
 sg13g2_decap_8 FILLER_74_2241 ();
 sg13g2_fill_1 FILLER_74_2308 ();
 sg13g2_fill_1 FILLER_74_2322 ();
 sg13g2_fill_1 FILLER_74_2328 ();
 sg13g2_decap_8 FILLER_74_2376 ();
 sg13g2_decap_8 FILLER_74_2383 ();
 sg13g2_fill_2 FILLER_74_2390 ();
 sg13g2_fill_1 FILLER_74_2392 ();
 sg13g2_decap_8 FILLER_74_2419 ();
 sg13g2_fill_1 FILLER_74_2434 ();
 sg13g2_fill_2 FILLER_74_2457 ();
 sg13g2_fill_2 FILLER_74_2485 ();
 sg13g2_fill_1 FILLER_74_2487 ();
 sg13g2_fill_1 FILLER_74_2493 ();
 sg13g2_fill_1 FILLER_74_2520 ();
 sg13g2_fill_2 FILLER_74_2533 ();
 sg13g2_decap_8 FILLER_74_2590 ();
 sg13g2_decap_8 FILLER_74_2597 ();
 sg13g2_decap_8 FILLER_74_2604 ();
 sg13g2_decap_8 FILLER_74_2611 ();
 sg13g2_decap_8 FILLER_74_2618 ();
 sg13g2_decap_8 FILLER_74_2625 ();
 sg13g2_decap_8 FILLER_74_2632 ();
 sg13g2_decap_8 FILLER_74_2639 ();
 sg13g2_decap_8 FILLER_74_2646 ();
 sg13g2_decap_8 FILLER_74_2653 ();
 sg13g2_decap_8 FILLER_74_2660 ();
 sg13g2_fill_2 FILLER_74_2667 ();
 sg13g2_fill_1 FILLER_74_2669 ();
 sg13g2_fill_2 FILLER_75_0 ();
 sg13g2_fill_1 FILLER_75_28 ();
 sg13g2_fill_2 FILLER_75_87 ();
 sg13g2_fill_1 FILLER_75_114 ();
 sg13g2_fill_2 FILLER_75_129 ();
 sg13g2_fill_1 FILLER_75_140 ();
 sg13g2_fill_2 FILLER_75_200 ();
 sg13g2_fill_2 FILLER_75_217 ();
 sg13g2_decap_8 FILLER_75_247 ();
 sg13g2_decap_8 FILLER_75_254 ();
 sg13g2_fill_1 FILLER_75_261 ();
 sg13g2_fill_1 FILLER_75_283 ();
 sg13g2_fill_1 FILLER_75_289 ();
 sg13g2_decap_8 FILLER_75_341 ();
 sg13g2_decap_8 FILLER_75_348 ();
 sg13g2_decap_8 FILLER_75_379 ();
 sg13g2_fill_2 FILLER_75_386 ();
 sg13g2_fill_1 FILLER_75_401 ();
 sg13g2_decap_8 FILLER_75_406 ();
 sg13g2_decap_8 FILLER_75_413 ();
 sg13g2_decap_8 FILLER_75_420 ();
 sg13g2_decap_8 FILLER_75_427 ();
 sg13g2_fill_2 FILLER_75_434 ();
 sg13g2_fill_1 FILLER_75_443 ();
 sg13g2_fill_1 FILLER_75_451 ();
 sg13g2_fill_1 FILLER_75_472 ();
 sg13g2_fill_1 FILLER_75_477 ();
 sg13g2_decap_4 FILLER_75_523 ();
 sg13g2_fill_2 FILLER_75_537 ();
 sg13g2_decap_4 FILLER_75_543 ();
 sg13g2_fill_1 FILLER_75_552 ();
 sg13g2_fill_1 FILLER_75_558 ();
 sg13g2_fill_1 FILLER_75_564 ();
 sg13g2_fill_2 FILLER_75_569 ();
 sg13g2_fill_2 FILLER_75_579 ();
 sg13g2_fill_1 FILLER_75_581 ();
 sg13g2_fill_1 FILLER_75_587 ();
 sg13g2_fill_1 FILLER_75_593 ();
 sg13g2_fill_1 FILLER_75_607 ();
 sg13g2_fill_2 FILLER_75_626 ();
 sg13g2_fill_2 FILLER_75_644 ();
 sg13g2_decap_8 FILLER_75_676 ();
 sg13g2_decap_4 FILLER_75_693 ();
 sg13g2_fill_1 FILLER_75_697 ();
 sg13g2_decap_8 FILLER_75_708 ();
 sg13g2_fill_1 FILLER_75_715 ();
 sg13g2_decap_4 FILLER_75_722 ();
 sg13g2_fill_1 FILLER_75_726 ();
 sg13g2_fill_2 FILLER_75_741 ();
 sg13g2_decap_8 FILLER_75_803 ();
 sg13g2_decap_4 FILLER_75_810 ();
 sg13g2_fill_1 FILLER_75_814 ();
 sg13g2_decap_4 FILLER_75_825 ();
 sg13g2_fill_2 FILLER_75_829 ();
 sg13g2_fill_1 FILLER_75_845 ();
 sg13g2_fill_2 FILLER_75_856 ();
 sg13g2_decap_8 FILLER_75_868 ();
 sg13g2_decap_4 FILLER_75_875 ();
 sg13g2_fill_2 FILLER_75_879 ();
 sg13g2_decap_8 FILLER_75_891 ();
 sg13g2_decap_8 FILLER_75_898 ();
 sg13g2_decap_8 FILLER_75_905 ();
 sg13g2_decap_4 FILLER_75_912 ();
 sg13g2_fill_2 FILLER_75_916 ();
 sg13g2_decap_8 FILLER_75_930 ();
 sg13g2_decap_4 FILLER_75_1006 ();
 sg13g2_fill_2 FILLER_75_1010 ();
 sg13g2_fill_2 FILLER_75_1016 ();
 sg13g2_decap_4 FILLER_75_1021 ();
 sg13g2_fill_1 FILLER_75_1025 ();
 sg13g2_decap_8 FILLER_75_1036 ();
 sg13g2_fill_2 FILLER_75_1053 ();
 sg13g2_fill_2 FILLER_75_1068 ();
 sg13g2_fill_1 FILLER_75_1088 ();
 sg13g2_decap_8 FILLER_75_1109 ();
 sg13g2_decap_8 FILLER_75_1116 ();
 sg13g2_decap_8 FILLER_75_1123 ();
 sg13g2_decap_4 FILLER_75_1162 ();
 sg13g2_fill_2 FILLER_75_1166 ();
 sg13g2_fill_2 FILLER_75_1182 ();
 sg13g2_fill_1 FILLER_75_1184 ();
 sg13g2_decap_8 FILLER_75_1231 ();
 sg13g2_decap_8 FILLER_75_1238 ();
 sg13g2_decap_8 FILLER_75_1245 ();
 sg13g2_decap_8 FILLER_75_1252 ();
 sg13g2_decap_8 FILLER_75_1259 ();
 sg13g2_decap_4 FILLER_75_1266 ();
 sg13g2_decap_8 FILLER_75_1273 ();
 sg13g2_fill_2 FILLER_75_1280 ();
 sg13g2_decap_8 FILLER_75_1318 ();
 sg13g2_fill_2 FILLER_75_1325 ();
 sg13g2_fill_1 FILLER_75_1327 ();
 sg13g2_decap_8 FILLER_75_1364 ();
 sg13g2_decap_4 FILLER_75_1381 ();
 sg13g2_fill_2 FILLER_75_1385 ();
 sg13g2_decap_8 FILLER_75_1391 ();
 sg13g2_decap_4 FILLER_75_1398 ();
 sg13g2_fill_1 FILLER_75_1402 ();
 sg13g2_fill_1 FILLER_75_1420 ();
 sg13g2_decap_4 FILLER_75_1461 ();
 sg13g2_fill_2 FILLER_75_1465 ();
 sg13g2_fill_1 FILLER_75_1508 ();
 sg13g2_fill_2 FILLER_75_1517 ();
 sg13g2_fill_2 FILLER_75_1542 ();
 sg13g2_fill_2 FILLER_75_1556 ();
 sg13g2_fill_1 FILLER_75_1558 ();
 sg13g2_fill_1 FILLER_75_1563 ();
 sg13g2_fill_1 FILLER_75_1577 ();
 sg13g2_fill_2 FILLER_75_1583 ();
 sg13g2_decap_4 FILLER_75_1601 ();
 sg13g2_fill_2 FILLER_75_1605 ();
 sg13g2_decap_8 FILLER_75_1641 ();
 sg13g2_decap_8 FILLER_75_1648 ();
 sg13g2_decap_8 FILLER_75_1655 ();
 sg13g2_decap_8 FILLER_75_1662 ();
 sg13g2_decap_8 FILLER_75_1669 ();
 sg13g2_fill_2 FILLER_75_1676 ();
 sg13g2_fill_1 FILLER_75_1678 ();
 sg13g2_decap_8 FILLER_75_1689 ();
 sg13g2_fill_2 FILLER_75_1700 ();
 sg13g2_fill_1 FILLER_75_1702 ();
 sg13g2_fill_1 FILLER_75_1707 ();
 sg13g2_fill_1 FILLER_75_1717 ();
 sg13g2_fill_1 FILLER_75_1745 ();
 sg13g2_fill_1 FILLER_75_1751 ();
 sg13g2_fill_2 FILLER_75_1757 ();
 sg13g2_decap_4 FILLER_75_1765 ();
 sg13g2_fill_2 FILLER_75_1769 ();
 sg13g2_decap_4 FILLER_75_1782 ();
 sg13g2_fill_1 FILLER_75_1790 ();
 sg13g2_decap_4 FILLER_75_1796 ();
 sg13g2_fill_1 FILLER_75_1800 ();
 sg13g2_fill_2 FILLER_75_1805 ();
 sg13g2_fill_2 FILLER_75_1836 ();
 sg13g2_fill_2 FILLER_75_1846 ();
 sg13g2_decap_4 FILLER_75_1853 ();
 sg13g2_fill_1 FILLER_75_1857 ();
 sg13g2_fill_2 FILLER_75_1879 ();
 sg13g2_decap_8 FILLER_75_1912 ();
 sg13g2_decap_4 FILLER_75_1919 ();
 sg13g2_decap_4 FILLER_75_1927 ();
 sg13g2_fill_2 FILLER_75_1931 ();
 sg13g2_decap_4 FILLER_75_1937 ();
 sg13g2_fill_1 FILLER_75_1941 ();
 sg13g2_fill_2 FILLER_75_1968 ();
 sg13g2_fill_1 FILLER_75_1970 ();
 sg13g2_fill_1 FILLER_75_2032 ();
 sg13g2_decap_8 FILLER_75_2037 ();
 sg13g2_fill_2 FILLER_75_2044 ();
 sg13g2_fill_1 FILLER_75_2046 ();
 sg13g2_decap_8 FILLER_75_2071 ();
 sg13g2_decap_4 FILLER_75_2172 ();
 sg13g2_fill_1 FILLER_75_2176 ();
 sg13g2_decap_8 FILLER_75_2203 ();
 sg13g2_decap_4 FILLER_75_2210 ();
 sg13g2_fill_2 FILLER_75_2276 ();
 sg13g2_fill_1 FILLER_75_2292 ();
 sg13g2_fill_1 FILLER_75_2306 ();
 sg13g2_fill_1 FILLER_75_2332 ();
 sg13g2_fill_2 FILLER_75_2343 ();
 sg13g2_fill_1 FILLER_75_2345 ();
 sg13g2_decap_8 FILLER_75_2350 ();
 sg13g2_fill_2 FILLER_75_2357 ();
 sg13g2_fill_2 FILLER_75_2385 ();
 sg13g2_fill_1 FILLER_75_2387 ();
 sg13g2_fill_2 FILLER_75_2414 ();
 sg13g2_decap_4 FILLER_75_2513 ();
 sg13g2_fill_1 FILLER_75_2532 ();
 sg13g2_fill_2 FILLER_75_2542 ();
 sg13g2_decap_8 FILLER_75_2594 ();
 sg13g2_decap_8 FILLER_75_2601 ();
 sg13g2_decap_8 FILLER_75_2608 ();
 sg13g2_decap_8 FILLER_75_2615 ();
 sg13g2_decap_8 FILLER_75_2622 ();
 sg13g2_decap_8 FILLER_75_2629 ();
 sg13g2_decap_8 FILLER_75_2636 ();
 sg13g2_decap_8 FILLER_75_2643 ();
 sg13g2_decap_8 FILLER_75_2650 ();
 sg13g2_decap_8 FILLER_75_2657 ();
 sg13g2_decap_4 FILLER_75_2664 ();
 sg13g2_fill_2 FILLER_75_2668 ();
 sg13g2_decap_8 FILLER_76_0 ();
 sg13g2_fill_2 FILLER_76_7 ();
 sg13g2_decap_8 FILLER_76_13 ();
 sg13g2_fill_2 FILLER_76_75 ();
 sg13g2_fill_2 FILLER_76_158 ();
 sg13g2_fill_1 FILLER_76_196 ();
 sg13g2_fill_2 FILLER_76_202 ();
 sg13g2_fill_2 FILLER_76_223 ();
 sg13g2_fill_2 FILLER_76_240 ();
 sg13g2_fill_1 FILLER_76_242 ();
 sg13g2_decap_4 FILLER_76_247 ();
 sg13g2_fill_2 FILLER_76_251 ();
 sg13g2_fill_2 FILLER_76_258 ();
 sg13g2_fill_2 FILLER_76_264 ();
 sg13g2_decap_4 FILLER_76_271 ();
 sg13g2_fill_1 FILLER_76_275 ();
 sg13g2_fill_1 FILLER_76_281 ();
 sg13g2_fill_1 FILLER_76_287 ();
 sg13g2_fill_2 FILLER_76_293 ();
 sg13g2_fill_1 FILLER_76_295 ();
 sg13g2_fill_2 FILLER_76_309 ();
 sg13g2_fill_1 FILLER_76_311 ();
 sg13g2_decap_8 FILLER_76_352 ();
 sg13g2_fill_1 FILLER_76_359 ();
 sg13g2_decap_4 FILLER_76_365 ();
 sg13g2_fill_1 FILLER_76_369 ();
 sg13g2_decap_4 FILLER_76_375 ();
 sg13g2_fill_2 FILLER_76_379 ();
 sg13g2_fill_2 FILLER_76_422 ();
 sg13g2_fill_1 FILLER_76_424 ();
 sg13g2_decap_8 FILLER_76_430 ();
 sg13g2_decap_8 FILLER_76_437 ();
 sg13g2_fill_2 FILLER_76_481 ();
 sg13g2_fill_1 FILLER_76_495 ();
 sg13g2_fill_2 FILLER_76_502 ();
 sg13g2_fill_1 FILLER_76_520 ();
 sg13g2_fill_1 FILLER_76_530 ();
 sg13g2_fill_1 FILLER_76_541 ();
 sg13g2_fill_2 FILLER_76_572 ();
 sg13g2_fill_1 FILLER_76_574 ();
 sg13g2_fill_2 FILLER_76_611 ();
 sg13g2_fill_1 FILLER_76_619 ();
 sg13g2_fill_1 FILLER_76_626 ();
 sg13g2_decap_8 FILLER_76_644 ();
 sg13g2_decap_4 FILLER_76_651 ();
 sg13g2_fill_1 FILLER_76_655 ();
 sg13g2_decap_4 FILLER_76_660 ();
 sg13g2_fill_2 FILLER_76_664 ();
 sg13g2_decap_4 FILLER_76_676 ();
 sg13g2_decap_8 FILLER_76_704 ();
 sg13g2_decap_8 FILLER_76_711 ();
 sg13g2_decap_8 FILLER_76_718 ();
 sg13g2_fill_2 FILLER_76_734 ();
 sg13g2_fill_1 FILLER_76_772 ();
 sg13g2_fill_2 FILLER_76_783 ();
 sg13g2_fill_2 FILLER_76_789 ();
 sg13g2_fill_2 FILLER_76_801 ();
 sg13g2_decap_8 FILLER_76_806 ();
 sg13g2_decap_8 FILLER_76_823 ();
 sg13g2_decap_8 FILLER_76_830 ();
 sg13g2_fill_1 FILLER_76_837 ();
 sg13g2_fill_1 FILLER_76_842 ();
 sg13g2_fill_1 FILLER_76_869 ();
 sg13g2_fill_2 FILLER_76_880 ();
 sg13g2_decap_8 FILLER_76_902 ();
 sg13g2_fill_2 FILLER_76_909 ();
 sg13g2_fill_1 FILLER_76_911 ();
 sg13g2_fill_2 FILLER_76_962 ();
 sg13g2_fill_1 FILLER_76_964 ();
 sg13g2_decap_8 FILLER_76_970 ();
 sg13g2_fill_1 FILLER_76_977 ();
 sg13g2_fill_2 FILLER_76_983 ();
 sg13g2_fill_1 FILLER_76_994 ();
 sg13g2_decap_8 FILLER_76_1001 ();
 sg13g2_decap_8 FILLER_76_1008 ();
 sg13g2_decap_4 FILLER_76_1015 ();
 sg13g2_decap_8 FILLER_76_1033 ();
 sg13g2_fill_1 FILLER_76_1070 ();
 sg13g2_fill_1 FILLER_76_1138 ();
 sg13g2_fill_2 FILLER_76_1152 ();
 sg13g2_fill_1 FILLER_76_1154 ();
 sg13g2_decap_8 FILLER_76_1185 ();
 sg13g2_decap_8 FILLER_76_1192 ();
 sg13g2_decap_4 FILLER_76_1199 ();
 sg13g2_decap_8 FILLER_76_1207 ();
 sg13g2_decap_8 FILLER_76_1214 ();
 sg13g2_decap_8 FILLER_76_1221 ();
 sg13g2_decap_8 FILLER_76_1228 ();
 sg13g2_fill_2 FILLER_76_1235 ();
 sg13g2_fill_1 FILLER_76_1237 ();
 sg13g2_decap_8 FILLER_76_1274 ();
 sg13g2_decap_8 FILLER_76_1307 ();
 sg13g2_decap_4 FILLER_76_1314 ();
 sg13g2_fill_2 FILLER_76_1318 ();
 sg13g2_decap_8 FILLER_76_1330 ();
 sg13g2_decap_8 FILLER_76_1337 ();
 sg13g2_fill_1 FILLER_76_1344 ();
 sg13g2_decap_8 FILLER_76_1349 ();
 sg13g2_decap_8 FILLER_76_1356 ();
 sg13g2_decap_4 FILLER_76_1363 ();
 sg13g2_fill_2 FILLER_76_1367 ();
 sg13g2_decap_8 FILLER_76_1373 ();
 sg13g2_decap_8 FILLER_76_1380 ();
 sg13g2_decap_8 FILLER_76_1387 ();
 sg13g2_decap_4 FILLER_76_1394 ();
 sg13g2_decap_8 FILLER_76_1424 ();
 sg13g2_decap_8 FILLER_76_1445 ();
 sg13g2_decap_8 FILLER_76_1452 ();
 sg13g2_decap_8 FILLER_76_1459 ();
 sg13g2_fill_1 FILLER_76_1466 ();
 sg13g2_fill_2 FILLER_76_1486 ();
 sg13g2_fill_2 FILLER_76_1497 ();
 sg13g2_fill_1 FILLER_76_1540 ();
 sg13g2_decap_4 FILLER_76_1573 ();
 sg13g2_fill_1 FILLER_76_1577 ();
 sg13g2_fill_1 FILLER_76_1585 ();
 sg13g2_fill_2 FILLER_76_1621 ();
 sg13g2_fill_1 FILLER_76_1627 ();
 sg13g2_decap_4 FILLER_76_1650 ();
 sg13g2_fill_1 FILLER_76_1654 ();
 sg13g2_fill_1 FILLER_76_1660 ();
 sg13g2_fill_2 FILLER_76_1675 ();
 sg13g2_fill_2 FILLER_76_1710 ();
 sg13g2_fill_1 FILLER_76_1716 ();
 sg13g2_fill_1 FILLER_76_1722 ();
 sg13g2_fill_1 FILLER_76_1743 ();
 sg13g2_fill_2 FILLER_76_1750 ();
 sg13g2_fill_2 FILLER_76_1767 ();
 sg13g2_fill_1 FILLER_76_1769 ();
 sg13g2_fill_2 FILLER_76_1801 ();
 sg13g2_fill_1 FILLER_76_1803 ();
 sg13g2_fill_2 FILLER_76_1809 ();
 sg13g2_fill_2 FILLER_76_1816 ();
 sg13g2_fill_2 FILLER_76_1856 ();
 sg13g2_fill_1 FILLER_76_1858 ();
 sg13g2_decap_8 FILLER_76_1863 ();
 sg13g2_decap_4 FILLER_76_1870 ();
 sg13g2_fill_2 FILLER_76_1879 ();
 sg13g2_fill_1 FILLER_76_1881 ();
 sg13g2_fill_2 FILLER_76_1890 ();
 sg13g2_fill_1 FILLER_76_1892 ();
 sg13g2_fill_1 FILLER_76_1911 ();
 sg13g2_fill_2 FILLER_76_1921 ();
 sg13g2_decap_4 FILLER_76_1926 ();
 sg13g2_fill_2 FILLER_76_1930 ();
 sg13g2_fill_2 FILLER_76_1936 ();
 sg13g2_fill_1 FILLER_76_1942 ();
 sg13g2_fill_1 FILLER_76_1955 ();
 sg13g2_decap_8 FILLER_76_1969 ();
 sg13g2_decap_8 FILLER_76_1976 ();
 sg13g2_decap_4 FILLER_76_1983 ();
 sg13g2_fill_1 FILLER_76_1991 ();
 sg13g2_decap_8 FILLER_76_2018 ();
 sg13g2_fill_1 FILLER_76_2025 ();
 sg13g2_fill_1 FILLER_76_2075 ();
 sg13g2_fill_2 FILLER_76_2079 ();
 sg13g2_fill_1 FILLER_76_2088 ();
 sg13g2_fill_1 FILLER_76_2152 ();
 sg13g2_fill_1 FILLER_76_2185 ();
 sg13g2_fill_1 FILLER_76_2212 ();
 sg13g2_decap_4 FILLER_76_2223 ();
 sg13g2_fill_1 FILLER_76_2253 ();
 sg13g2_fill_2 FILLER_76_2267 ();
 sg13g2_decap_8 FILLER_76_2299 ();
 sg13g2_decap_8 FILLER_76_2344 ();
 sg13g2_decap_8 FILLER_76_2416 ();
 sg13g2_fill_2 FILLER_76_2423 ();
 sg13g2_fill_1 FILLER_76_2425 ();
 sg13g2_decap_4 FILLER_76_2430 ();
 sg13g2_fill_1 FILLER_76_2434 ();
 sg13g2_fill_1 FILLER_76_2449 ();
 sg13g2_fill_1 FILLER_76_2454 ();
 sg13g2_fill_2 FILLER_76_2469 ();
 sg13g2_fill_1 FILLER_76_2475 ();
 sg13g2_decap_4 FILLER_76_2481 ();
 sg13g2_fill_1 FILLER_76_2485 ();
 sg13g2_decap_4 FILLER_76_2495 ();
 sg13g2_fill_2 FILLER_76_2499 ();
 sg13g2_decap_4 FILLER_76_2514 ();
 sg13g2_fill_2 FILLER_76_2524 ();
 sg13g2_fill_1 FILLER_76_2526 ();
 sg13g2_fill_2 FILLER_76_2540 ();
 sg13g2_decap_8 FILLER_76_2568 ();
 sg13g2_decap_8 FILLER_76_2575 ();
 sg13g2_decap_8 FILLER_76_2582 ();
 sg13g2_decap_8 FILLER_76_2589 ();
 sg13g2_decap_8 FILLER_76_2596 ();
 sg13g2_decap_8 FILLER_76_2603 ();
 sg13g2_decap_8 FILLER_76_2610 ();
 sg13g2_decap_8 FILLER_76_2617 ();
 sg13g2_decap_8 FILLER_76_2624 ();
 sg13g2_decap_8 FILLER_76_2631 ();
 sg13g2_decap_8 FILLER_76_2638 ();
 sg13g2_decap_8 FILLER_76_2645 ();
 sg13g2_decap_8 FILLER_76_2652 ();
 sg13g2_decap_8 FILLER_76_2659 ();
 sg13g2_decap_4 FILLER_76_2666 ();
 sg13g2_decap_8 FILLER_77_0 ();
 sg13g2_fill_2 FILLER_77_7 ();
 sg13g2_fill_1 FILLER_77_9 ();
 sg13g2_fill_1 FILLER_77_34 ();
 sg13g2_fill_1 FILLER_77_48 ();
 sg13g2_fill_1 FILLER_77_134 ();
 sg13g2_fill_1 FILLER_77_178 ();
 sg13g2_decap_8 FILLER_77_222 ();
 sg13g2_fill_2 FILLER_77_229 ();
 sg13g2_fill_1 FILLER_77_231 ();
 sg13g2_fill_1 FILLER_77_268 ();
 sg13g2_fill_2 FILLER_77_283 ();
 sg13g2_fill_1 FILLER_77_285 ();
 sg13g2_fill_1 FILLER_77_296 ();
 sg13g2_decap_8 FILLER_77_312 ();
 sg13g2_decap_4 FILLER_77_319 ();
 sg13g2_fill_1 FILLER_77_323 ();
 sg13g2_fill_1 FILLER_77_328 ();
 sg13g2_fill_1 FILLER_77_333 ();
 sg13g2_fill_1 FILLER_77_391 ();
 sg13g2_fill_2 FILLER_77_405 ();
 sg13g2_fill_1 FILLER_77_407 ();
 sg13g2_fill_2 FILLER_77_412 ();
 sg13g2_decap_8 FILLER_77_440 ();
 sg13g2_decap_4 FILLER_77_447 ();
 sg13g2_fill_1 FILLER_77_451 ();
 sg13g2_decap_8 FILLER_77_467 ();
 sg13g2_fill_2 FILLER_77_479 ();
 sg13g2_fill_2 FILLER_77_491 ();
 sg13g2_fill_2 FILLER_77_514 ();
 sg13g2_fill_1 FILLER_77_516 ();
 sg13g2_fill_1 FILLER_77_525 ();
 sg13g2_fill_1 FILLER_77_540 ();
 sg13g2_fill_1 FILLER_77_551 ();
 sg13g2_fill_2 FILLER_77_574 ();
 sg13g2_fill_1 FILLER_77_606 ();
 sg13g2_fill_2 FILLER_77_633 ();
 sg13g2_fill_2 FILLER_77_648 ();
 sg13g2_decap_8 FILLER_77_654 ();
 sg13g2_decap_8 FILLER_77_661 ();
 sg13g2_decap_4 FILLER_77_668 ();
 sg13g2_decap_8 FILLER_77_698 ();
 sg13g2_decap_8 FILLER_77_741 ();
 sg13g2_decap_4 FILLER_77_748 ();
 sg13g2_fill_2 FILLER_77_798 ();
 sg13g2_fill_1 FILLER_77_800 ();
 sg13g2_decap_4 FILLER_77_807 ();
 sg13g2_fill_2 FILLER_77_811 ();
 sg13g2_fill_1 FILLER_77_839 ();
 sg13g2_fill_1 FILLER_77_850 ();
 sg13g2_fill_2 FILLER_77_964 ();
 sg13g2_decap_8 FILLER_77_997 ();
 sg13g2_fill_2 FILLER_77_1004 ();
 sg13g2_decap_8 FILLER_77_1042 ();
 sg13g2_fill_2 FILLER_77_1078 ();
 sg13g2_fill_1 FILLER_77_1083 ();
 sg13g2_decap_8 FILLER_77_1124 ();
 sg13g2_fill_1 FILLER_77_1131 ();
 sg13g2_fill_2 FILLER_77_1158 ();
 sg13g2_fill_1 FILLER_77_1160 ();
 sg13g2_decap_8 FILLER_77_1165 ();
 sg13g2_decap_4 FILLER_77_1172 ();
 sg13g2_fill_2 FILLER_77_1242 ();
 sg13g2_fill_1 FILLER_77_1244 ();
 sg13g2_fill_2 FILLER_77_1249 ();
 sg13g2_fill_1 FILLER_77_1251 ();
 sg13g2_fill_2 FILLER_77_1317 ();
 sg13g2_fill_1 FILLER_77_1345 ();
 sg13g2_decap_4 FILLER_77_1356 ();
 sg13g2_fill_1 FILLER_77_1360 ();
 sg13g2_fill_2 FILLER_77_1449 ();
 sg13g2_fill_1 FILLER_77_1455 ();
 sg13g2_fill_1 FILLER_77_1466 ();
 sg13g2_decap_4 FILLER_77_1471 ();
 sg13g2_fill_1 FILLER_77_1475 ();
 sg13g2_fill_1 FILLER_77_1482 ();
 sg13g2_fill_1 FILLER_77_1498 ();
 sg13g2_fill_1 FILLER_77_1512 ();
 sg13g2_fill_1 FILLER_77_1519 ();
 sg13g2_decap_4 FILLER_77_1559 ();
 sg13g2_fill_2 FILLER_77_1569 ();
 sg13g2_fill_1 FILLER_77_1599 ();
 sg13g2_fill_1 FILLER_77_1615 ();
 sg13g2_fill_1 FILLER_77_1621 ();
 sg13g2_fill_1 FILLER_77_1628 ();
 sg13g2_fill_1 FILLER_77_1633 ();
 sg13g2_decap_4 FILLER_77_1658 ();
 sg13g2_fill_2 FILLER_77_1666 ();
 sg13g2_fill_1 FILLER_77_1668 ();
 sg13g2_fill_2 FILLER_77_1713 ();
 sg13g2_fill_1 FILLER_77_1730 ();
 sg13g2_fill_1 FILLER_77_1779 ();
 sg13g2_fill_1 FILLER_77_1795 ();
 sg13g2_fill_2 FILLER_77_1831 ();
 sg13g2_fill_1 FILLER_77_1833 ();
 sg13g2_fill_1 FILLER_77_1844 ();
 sg13g2_fill_1 FILLER_77_1850 ();
 sg13g2_fill_2 FILLER_77_1859 ();
 sg13g2_fill_1 FILLER_77_1869 ();
 sg13g2_fill_1 FILLER_77_1880 ();
 sg13g2_fill_1 FILLER_77_1886 ();
 sg13g2_fill_1 FILLER_77_1919 ();
 sg13g2_fill_1 FILLER_77_1977 ();
 sg13g2_decap_4 FILLER_77_2003 ();
 sg13g2_fill_1 FILLER_77_2007 ();
 sg13g2_fill_2 FILLER_77_2018 ();
 sg13g2_fill_1 FILLER_77_2020 ();
 sg13g2_fill_2 FILLER_77_2031 ();
 sg13g2_fill_1 FILLER_77_2033 ();
 sg13g2_decap_4 FILLER_77_2070 ();
 sg13g2_fill_2 FILLER_77_2074 ();
 sg13g2_fill_1 FILLER_77_2183 ();
 sg13g2_fill_1 FILLER_77_2194 ();
 sg13g2_fill_2 FILLER_77_2199 ();
 sg13g2_fill_1 FILLER_77_2211 ();
 sg13g2_decap_8 FILLER_77_2247 ();
 sg13g2_fill_2 FILLER_77_2254 ();
 sg13g2_fill_1 FILLER_77_2260 ();
 sg13g2_decap_8 FILLER_77_2281 ();
 sg13g2_decap_8 FILLER_77_2288 ();
 sg13g2_decap_8 FILLER_77_2295 ();
 sg13g2_fill_1 FILLER_77_2302 ();
 sg13g2_decap_4 FILLER_77_2338 ();
 sg13g2_fill_1 FILLER_77_2342 ();
 sg13g2_fill_2 FILLER_77_2348 ();
 sg13g2_fill_2 FILLER_77_2399 ();
 sg13g2_fill_1 FILLER_77_2401 ();
 sg13g2_fill_2 FILLER_77_2412 ();
 sg13g2_fill_2 FILLER_77_2450 ();
 sg13g2_fill_1 FILLER_77_2452 ();
 sg13g2_decap_4 FILLER_77_2459 ();
 sg13g2_fill_1 FILLER_77_2463 ();
 sg13g2_decap_8 FILLER_77_2480 ();
 sg13g2_decap_8 FILLER_77_2491 ();
 sg13g2_fill_1 FILLER_77_2498 ();
 sg13g2_fill_2 FILLER_77_2544 ();
 sg13g2_fill_1 FILLER_77_2549 ();
 sg13g2_decap_8 FILLER_77_2563 ();
 sg13g2_decap_8 FILLER_77_2570 ();
 sg13g2_decap_8 FILLER_77_2577 ();
 sg13g2_decap_8 FILLER_77_2584 ();
 sg13g2_decap_8 FILLER_77_2591 ();
 sg13g2_decap_8 FILLER_77_2598 ();
 sg13g2_decap_8 FILLER_77_2605 ();
 sg13g2_decap_8 FILLER_77_2612 ();
 sg13g2_decap_8 FILLER_77_2619 ();
 sg13g2_decap_8 FILLER_77_2626 ();
 sg13g2_decap_8 FILLER_77_2633 ();
 sg13g2_decap_8 FILLER_77_2640 ();
 sg13g2_decap_8 FILLER_77_2647 ();
 sg13g2_decap_8 FILLER_77_2654 ();
 sg13g2_decap_8 FILLER_77_2661 ();
 sg13g2_fill_2 FILLER_77_2668 ();
 sg13g2_fill_2 FILLER_78_0 ();
 sg13g2_fill_2 FILLER_78_28 ();
 sg13g2_fill_2 FILLER_78_72 ();
 sg13g2_fill_1 FILLER_78_116 ();
 sg13g2_fill_2 FILLER_78_125 ();
 sg13g2_fill_2 FILLER_78_170 ();
 sg13g2_fill_2 FILLER_78_214 ();
 sg13g2_fill_1 FILLER_78_246 ();
 sg13g2_fill_2 FILLER_78_273 ();
 sg13g2_decap_8 FILLER_78_301 ();
 sg13g2_fill_2 FILLER_78_308 ();
 sg13g2_decap_8 FILLER_78_336 ();
 sg13g2_decap_8 FILLER_78_343 ();
 sg13g2_fill_1 FILLER_78_350 ();
 sg13g2_fill_1 FILLER_78_370 ();
 sg13g2_fill_2 FILLER_78_389 ();
 sg13g2_fill_1 FILLER_78_391 ();
 sg13g2_decap_4 FILLER_78_396 ();
 sg13g2_fill_1 FILLER_78_429 ();
 sg13g2_decap_4 FILLER_78_444 ();
 sg13g2_fill_2 FILLER_78_478 ();
 sg13g2_fill_1 FILLER_78_489 ();
 sg13g2_fill_1 FILLER_78_509 ();
 sg13g2_fill_1 FILLER_78_552 ();
 sg13g2_fill_1 FILLER_78_565 ();
 sg13g2_fill_1 FILLER_78_578 ();
 sg13g2_fill_1 FILLER_78_582 ();
 sg13g2_fill_2 FILLER_78_587 ();
 sg13g2_fill_2 FILLER_78_705 ();
 sg13g2_decap_4 FILLER_78_769 ();
 sg13g2_fill_2 FILLER_78_773 ();
 sg13g2_fill_2 FILLER_78_811 ();
 sg13g2_fill_2 FILLER_78_865 ();
 sg13g2_fill_1 FILLER_78_867 ();
 sg13g2_fill_2 FILLER_78_904 ();
 sg13g2_fill_1 FILLER_78_906 ();
 sg13g2_fill_1 FILLER_78_947 ();
 sg13g2_fill_1 FILLER_78_974 ();
 sg13g2_fill_2 FILLER_78_1053 ();
 sg13g2_fill_1 FILLER_78_1060 ();
 sg13g2_fill_1 FILLER_78_1095 ();
 sg13g2_fill_1 FILLER_78_1106 ();
 sg13g2_fill_1 FILLER_78_1133 ();
 sg13g2_fill_1 FILLER_78_1138 ();
 sg13g2_fill_1 FILLER_78_1165 ();
 sg13g2_fill_2 FILLER_78_1192 ();
 sg13g2_fill_2 FILLER_78_1220 ();
 sg13g2_fill_2 FILLER_78_1248 ();
 sg13g2_fill_2 FILLER_78_1276 ();
 sg13g2_fill_1 FILLER_78_1278 ();
 sg13g2_fill_2 FILLER_78_1289 ();
 sg13g2_fill_1 FILLER_78_1291 ();
 sg13g2_fill_2 FILLER_78_1378 ();
 sg13g2_fill_2 FILLER_78_1390 ();
 sg13g2_fill_1 FILLER_78_1392 ();
 sg13g2_fill_1 FILLER_78_1403 ();
 sg13g2_fill_2 FILLER_78_1466 ();
 sg13g2_fill_2 FILLER_78_1494 ();
 sg13g2_fill_1 FILLER_78_1522 ();
 sg13g2_fill_1 FILLER_78_1528 ();
 sg13g2_fill_1 FILLER_78_1570 ();
 sg13g2_fill_1 FILLER_78_1623 ();
 sg13g2_decap_8 FILLER_78_1649 ();
 sg13g2_decap_8 FILLER_78_1656 ();
 sg13g2_decap_4 FILLER_78_1663 ();
 sg13g2_fill_1 FILLER_78_1667 ();
 sg13g2_fill_2 FILLER_78_1683 ();
 sg13g2_fill_1 FILLER_78_1718 ();
 sg13g2_fill_1 FILLER_78_1754 ();
 sg13g2_fill_2 FILLER_78_1793 ();
 sg13g2_fill_2 FILLER_78_1830 ();
 sg13g2_decap_8 FILLER_78_1835 ();
 sg13g2_fill_1 FILLER_78_1842 ();
 sg13g2_fill_1 FILLER_78_1847 ();
 sg13g2_fill_1 FILLER_78_1900 ();
 sg13g2_fill_1 FILLER_78_1910 ();
 sg13g2_fill_1 FILLER_78_1916 ();
 sg13g2_fill_1 FILLER_78_1924 ();
 sg13g2_fill_1 FILLER_78_1951 ();
 sg13g2_fill_1 FILLER_78_1963 ();
 sg13g2_decap_8 FILLER_78_2000 ();
 sg13g2_decap_4 FILLER_78_2007 ();
 sg13g2_fill_2 FILLER_78_2021 ();
 sg13g2_fill_1 FILLER_78_2023 ();
 sg13g2_decap_4 FILLER_78_2082 ();
 sg13g2_fill_2 FILLER_78_2086 ();
 sg13g2_fill_1 FILLER_78_2110 ();
 sg13g2_decap_4 FILLER_78_2186 ();
 sg13g2_fill_1 FILLER_78_2190 ();
 sg13g2_fill_1 FILLER_78_2195 ();
 sg13g2_fill_2 FILLER_78_2206 ();
 sg13g2_decap_8 FILLER_78_2238 ();
 sg13g2_decap_8 FILLER_78_2245 ();
 sg13g2_decap_8 FILLER_78_2252 ();
 sg13g2_fill_2 FILLER_78_2259 ();
 sg13g2_fill_2 FILLER_78_2267 ();
 sg13g2_decap_8 FILLER_78_2281 ();
 sg13g2_decap_4 FILLER_78_2288 ();
 sg13g2_fill_1 FILLER_78_2292 ();
 sg13g2_fill_2 FILLER_78_2387 ();
 sg13g2_decap_8 FILLER_78_2415 ();
 sg13g2_fill_1 FILLER_78_2422 ();
 sg13g2_fill_2 FILLER_78_2454 ();
 sg13g2_decap_8 FILLER_78_2487 ();
 sg13g2_fill_2 FILLER_78_2494 ();
 sg13g2_fill_2 FILLER_78_2527 ();
 sg13g2_decap_8 FILLER_78_2560 ();
 sg13g2_decap_8 FILLER_78_2567 ();
 sg13g2_decap_8 FILLER_78_2574 ();
 sg13g2_decap_8 FILLER_78_2581 ();
 sg13g2_decap_8 FILLER_78_2588 ();
 sg13g2_decap_8 FILLER_78_2595 ();
 sg13g2_decap_8 FILLER_78_2602 ();
 sg13g2_decap_8 FILLER_78_2609 ();
 sg13g2_decap_8 FILLER_78_2616 ();
 sg13g2_decap_8 FILLER_78_2623 ();
 sg13g2_decap_8 FILLER_78_2630 ();
 sg13g2_decap_8 FILLER_78_2637 ();
 sg13g2_decap_8 FILLER_78_2644 ();
 sg13g2_decap_8 FILLER_78_2651 ();
 sg13g2_decap_8 FILLER_78_2658 ();
 sg13g2_decap_4 FILLER_78_2665 ();
 sg13g2_fill_1 FILLER_78_2669 ();
 sg13g2_fill_2 FILLER_79_0 ();
 sg13g2_fill_2 FILLER_79_35 ();
 sg13g2_fill_1 FILLER_79_37 ();
 sg13g2_fill_1 FILLER_79_67 ();
 sg13g2_fill_2 FILLER_79_107 ();
 sg13g2_fill_1 FILLER_79_139 ();
 sg13g2_fill_1 FILLER_79_147 ();
 sg13g2_fill_1 FILLER_79_178 ();
 sg13g2_fill_1 FILLER_79_185 ();
 sg13g2_fill_1 FILLER_79_212 ();
 sg13g2_decap_8 FILLER_79_247 ();
 sg13g2_decap_8 FILLER_79_334 ();
 sg13g2_decap_8 FILLER_79_341 ();
 sg13g2_decap_8 FILLER_79_348 ();
 sg13g2_decap_8 FILLER_79_355 ();
 sg13g2_fill_1 FILLER_79_362 ();
 sg13g2_decap_4 FILLER_79_370 ();
 sg13g2_fill_1 FILLER_79_374 ();
 sg13g2_fill_1 FILLER_79_409 ();
 sg13g2_fill_1 FILLER_79_462 ();
 sg13g2_decap_8 FILLER_79_489 ();
 sg13g2_decap_4 FILLER_79_496 ();
 sg13g2_decap_8 FILLER_79_503 ();
 sg13g2_fill_2 FILLER_79_510 ();
 sg13g2_fill_1 FILLER_79_542 ();
 sg13g2_fill_2 FILLER_79_569 ();
 sg13g2_fill_1 FILLER_79_597 ();
 sg13g2_fill_2 FILLER_79_624 ();
 sg13g2_fill_2 FILLER_79_630 ();
 sg13g2_fill_2 FILLER_79_658 ();
 sg13g2_fill_1 FILLER_79_660 ();
 sg13g2_fill_1 FILLER_79_675 ();
 sg13g2_fill_2 FILLER_79_680 ();
 sg13g2_fill_2 FILLER_79_692 ();
 sg13g2_fill_2 FILLER_79_704 ();
 sg13g2_fill_1 FILLER_79_706 ();
 sg13g2_fill_2 FILLER_79_711 ();
 sg13g2_fill_1 FILLER_79_713 ();
 sg13g2_decap_8 FILLER_79_718 ();
 sg13g2_decap_4 FILLER_79_738 ();
 sg13g2_fill_1 FILLER_79_742 ();
 sg13g2_decap_4 FILLER_79_773 ();
 sg13g2_fill_1 FILLER_79_777 ();
 sg13g2_fill_2 FILLER_79_814 ();
 sg13g2_fill_1 FILLER_79_838 ();
 sg13g2_fill_1 FILLER_79_865 ();
 sg13g2_decap_8 FILLER_79_902 ();
 sg13g2_decap_4 FILLER_79_909 ();
 sg13g2_fill_1 FILLER_79_913 ();
 sg13g2_decap_4 FILLER_79_963 ();
 sg13g2_fill_1 FILLER_79_967 ();
 sg13g2_decap_4 FILLER_79_1026 ();
 sg13g2_fill_1 FILLER_79_1034 ();
 sg13g2_decap_4 FILLER_79_1039 ();
 sg13g2_fill_1 FILLER_79_1043 ();
 sg13g2_fill_1 FILLER_79_1064 ();
 sg13g2_fill_1 FILLER_79_1094 ();
 sg13g2_fill_2 FILLER_79_1109 ();
 sg13g2_fill_1 FILLER_79_1111 ();
 sg13g2_fill_2 FILLER_79_1116 ();
 sg13g2_fill_1 FILLER_79_1118 ();
 sg13g2_fill_2 FILLER_79_1123 ();
 sg13g2_fill_1 FILLER_79_1125 ();
 sg13g2_fill_1 FILLER_79_1152 ();
 sg13g2_fill_1 FILLER_79_1157 ();
 sg13g2_fill_1 FILLER_79_1168 ();
 sg13g2_fill_1 FILLER_79_1179 ();
 sg13g2_fill_2 FILLER_79_1210 ();
 sg13g2_fill_1 FILLER_79_1252 ();
 sg13g2_fill_1 FILLER_79_1257 ();
 sg13g2_fill_1 FILLER_79_1262 ();
 sg13g2_fill_2 FILLER_79_1273 ();
 sg13g2_decap_4 FILLER_79_1301 ();
 sg13g2_fill_1 FILLER_79_1305 ();
 sg13g2_fill_1 FILLER_79_1332 ();
 sg13g2_fill_1 FILLER_79_1338 ();
 sg13g2_fill_2 FILLER_79_1385 ();
 sg13g2_decap_8 FILLER_79_1413 ();
 sg13g2_fill_1 FILLER_79_1420 ();
 sg13g2_fill_2 FILLER_79_1425 ();
 sg13g2_fill_1 FILLER_79_1427 ();
 sg13g2_fill_2 FILLER_79_1441 ();
 sg13g2_fill_1 FILLER_79_1443 ();
 sg13g2_fill_2 FILLER_79_1474 ();
 sg13g2_decap_8 FILLER_79_1484 ();
 sg13g2_fill_1 FILLER_79_1491 ();
 sg13g2_decap_8 FILLER_79_1526 ();
 sg13g2_fill_2 FILLER_79_1533 ();
 sg13g2_fill_1 FILLER_79_1535 ();
 sg13g2_fill_2 FILLER_79_1543 ();
 sg13g2_fill_2 FILLER_79_1553 ();
 sg13g2_fill_2 FILLER_79_1587 ();
 sg13g2_decap_8 FILLER_79_1598 ();
 sg13g2_decap_8 FILLER_79_1605 ();
 sg13g2_fill_1 FILLER_79_1612 ();
 sg13g2_decap_8 FILLER_79_1646 ();
 sg13g2_decap_8 FILLER_79_1653 ();
 sg13g2_decap_8 FILLER_79_1660 ();
 sg13g2_decap_4 FILLER_79_1667 ();
 sg13g2_fill_1 FILLER_79_1671 ();
 sg13g2_fill_1 FILLER_79_1682 ();
 sg13g2_decap_8 FILLER_79_1738 ();
 sg13g2_decap_4 FILLER_79_1745 ();
 sg13g2_fill_1 FILLER_79_1749 ();
 sg13g2_decap_4 FILLER_79_1779 ();
 sg13g2_fill_2 FILLER_79_1792 ();
 sg13g2_decap_8 FILLER_79_1807 ();
 sg13g2_decap_8 FILLER_79_1814 ();
 sg13g2_decap_8 FILLER_79_1821 ();
 sg13g2_fill_2 FILLER_79_1828 ();
 sg13g2_decap_8 FILLER_79_1849 ();
 sg13g2_fill_1 FILLER_79_1856 ();
 sg13g2_fill_1 FILLER_79_1862 ();
 sg13g2_fill_1 FILLER_79_1872 ();
 sg13g2_decap_4 FILLER_79_1877 ();
 sg13g2_fill_1 FILLER_79_1881 ();
 sg13g2_fill_2 FILLER_79_1886 ();
 sg13g2_fill_1 FILLER_79_1888 ();
 sg13g2_fill_2 FILLER_79_1906 ();
 sg13g2_fill_2 FILLER_79_1960 ();
 sg13g2_fill_2 FILLER_79_2040 ();
 sg13g2_decap_4 FILLER_79_2068 ();
 sg13g2_decap_8 FILLER_79_2092 ();
 sg13g2_fill_1 FILLER_79_2142 ();
 sg13g2_decap_4 FILLER_79_2179 ();
 sg13g2_fill_1 FILLER_79_2183 ();
 sg13g2_decap_8 FILLER_79_2188 ();
 sg13g2_fill_1 FILLER_79_2195 ();
 sg13g2_decap_8 FILLER_79_2235 ();
 sg13g2_decap_8 FILLER_79_2242 ();
 sg13g2_decap_8 FILLER_79_2249 ();
 sg13g2_decap_8 FILLER_79_2256 ();
 sg13g2_decap_8 FILLER_79_2263 ();
 sg13g2_decap_8 FILLER_79_2270 ();
 sg13g2_decap_8 FILLER_79_2277 ();
 sg13g2_decap_8 FILLER_79_2284 ();
 sg13g2_decap_8 FILLER_79_2291 ();
 sg13g2_fill_1 FILLER_79_2298 ();
 sg13g2_fill_1 FILLER_79_2303 ();
 sg13g2_fill_1 FILLER_79_2334 ();
 sg13g2_fill_1 FILLER_79_2340 ();
 sg13g2_fill_1 FILLER_79_2383 ();
 sg13g2_decap_8 FILLER_79_2414 ();
 sg13g2_decap_8 FILLER_79_2564 ();
 sg13g2_decap_8 FILLER_79_2571 ();
 sg13g2_decap_8 FILLER_79_2578 ();
 sg13g2_decap_8 FILLER_79_2585 ();
 sg13g2_decap_8 FILLER_79_2592 ();
 sg13g2_decap_8 FILLER_79_2599 ();
 sg13g2_decap_8 FILLER_79_2606 ();
 sg13g2_decap_8 FILLER_79_2613 ();
 sg13g2_decap_8 FILLER_79_2620 ();
 sg13g2_decap_8 FILLER_79_2627 ();
 sg13g2_decap_8 FILLER_79_2634 ();
 sg13g2_decap_8 FILLER_79_2641 ();
 sg13g2_decap_8 FILLER_79_2648 ();
 sg13g2_decap_8 FILLER_79_2655 ();
 sg13g2_decap_8 FILLER_79_2662 ();
 sg13g2_fill_1 FILLER_79_2669 ();
 sg13g2_decap_4 FILLER_80_0 ();
 sg13g2_fill_1 FILLER_80_4 ();
 sg13g2_fill_2 FILLER_80_43 ();
 sg13g2_fill_1 FILLER_80_54 ();
 sg13g2_fill_2 FILLER_80_76 ();
 sg13g2_fill_1 FILLER_80_117 ();
 sg13g2_fill_2 FILLER_80_122 ();
 sg13g2_fill_2 FILLER_80_152 ();
 sg13g2_fill_1 FILLER_80_186 ();
 sg13g2_decap_8 FILLER_80_245 ();
 sg13g2_fill_1 FILLER_80_252 ();
 sg13g2_decap_4 FILLER_80_261 ();
 sg13g2_decap_4 FILLER_80_269 ();
 sg13g2_fill_1 FILLER_80_281 ();
 sg13g2_fill_2 FILLER_80_301 ();
 sg13g2_fill_1 FILLER_80_303 ();
 sg13g2_decap_8 FILLER_80_309 ();
 sg13g2_decap_4 FILLER_80_328 ();
 sg13g2_fill_2 FILLER_80_332 ();
 sg13g2_fill_1 FILLER_80_339 ();
 sg13g2_fill_2 FILLER_80_345 ();
 sg13g2_fill_1 FILLER_80_347 ();
 sg13g2_decap_4 FILLER_80_353 ();
 sg13g2_fill_2 FILLER_80_357 ();
 sg13g2_fill_2 FILLER_80_374 ();
 sg13g2_fill_1 FILLER_80_376 ();
 sg13g2_decap_4 FILLER_80_382 ();
 sg13g2_decap_8 FILLER_80_395 ();
 sg13g2_decap_8 FILLER_80_406 ();
 sg13g2_fill_2 FILLER_80_413 ();
 sg13g2_decap_8 FILLER_80_423 ();
 sg13g2_fill_1 FILLER_80_430 ();
 sg13g2_decap_4 FILLER_80_436 ();
 sg13g2_fill_2 FILLER_80_440 ();
 sg13g2_decap_8 FILLER_80_446 ();
 sg13g2_fill_2 FILLER_80_453 ();
 sg13g2_fill_1 FILLER_80_455 ();
 sg13g2_decap_8 FILLER_80_460 ();
 sg13g2_decap_4 FILLER_80_467 ();
 sg13g2_fill_1 FILLER_80_471 ();
 sg13g2_decap_8 FILLER_80_476 ();
 sg13g2_decap_8 FILLER_80_483 ();
 sg13g2_decap_8 FILLER_80_542 ();
 sg13g2_fill_1 FILLER_80_549 ();
 sg13g2_decap_8 FILLER_80_567 ();
 sg13g2_fill_2 FILLER_80_574 ();
 sg13g2_fill_1 FILLER_80_576 ();
 sg13g2_decap_8 FILLER_80_581 ();
 sg13g2_decap_8 FILLER_80_588 ();
 sg13g2_decap_4 FILLER_80_614 ();
 sg13g2_decap_8 FILLER_80_648 ();
 sg13g2_decap_4 FILLER_80_655 ();
 sg13g2_decap_8 FILLER_80_685 ();
 sg13g2_decap_8 FILLER_80_692 ();
 sg13g2_decap_8 FILLER_80_699 ();
 sg13g2_decap_8 FILLER_80_706 ();
 sg13g2_decap_8 FILLER_80_713 ();
 sg13g2_fill_2 FILLER_80_720 ();
 sg13g2_fill_1 FILLER_80_722 ();
 sg13g2_decap_8 FILLER_80_761 ();
 sg13g2_decap_8 FILLER_80_768 ();
 sg13g2_decap_8 FILLER_80_775 ();
 sg13g2_decap_8 FILLER_80_782 ();
 sg13g2_decap_4 FILLER_80_789 ();
 sg13g2_fill_1 FILLER_80_793 ();
 sg13g2_decap_8 FILLER_80_802 ();
 sg13g2_decap_4 FILLER_80_809 ();
 sg13g2_fill_2 FILLER_80_813 ();
 sg13g2_decap_8 FILLER_80_819 ();
 sg13g2_decap_8 FILLER_80_826 ();
 sg13g2_fill_2 FILLER_80_833 ();
 sg13g2_decap_4 FILLER_80_839 ();
 sg13g2_decap_8 FILLER_80_857 ();
 sg13g2_decap_4 FILLER_80_864 ();
 sg13g2_fill_1 FILLER_80_868 ();
 sg13g2_decap_8 FILLER_80_873 ();
 sg13g2_decap_4 FILLER_80_880 ();
 sg13g2_fill_1 FILLER_80_884 ();
 sg13g2_decap_8 FILLER_80_893 ();
 sg13g2_decap_8 FILLER_80_900 ();
 sg13g2_decap_8 FILLER_80_907 ();
 sg13g2_fill_2 FILLER_80_914 ();
 sg13g2_fill_1 FILLER_80_916 ();
 sg13g2_decap_4 FILLER_80_931 ();
 sg13g2_decap_8 FILLER_80_939 ();
 sg13g2_decap_8 FILLER_80_946 ();
 sg13g2_decap_8 FILLER_80_953 ();
 sg13g2_decap_8 FILLER_80_960 ();
 sg13g2_decap_8 FILLER_80_967 ();
 sg13g2_decap_4 FILLER_80_974 ();
 sg13g2_decap_8 FILLER_80_1002 ();
 sg13g2_decap_8 FILLER_80_1009 ();
 sg13g2_decap_8 FILLER_80_1016 ();
 sg13g2_fill_1 FILLER_80_1023 ();
 sg13g2_decap_4 FILLER_80_1050 ();
 sg13g2_fill_1 FILLER_80_1054 ();
 sg13g2_fill_2 FILLER_80_1075 ();
 sg13g2_decap_8 FILLER_80_1096 ();
 sg13g2_decap_4 FILLER_80_1103 ();
 sg13g2_fill_1 FILLER_80_1107 ();
 sg13g2_decap_4 FILLER_80_1134 ();
 sg13g2_decap_8 FILLER_80_1148 ();
 sg13g2_decap_8 FILLER_80_1155 ();
 sg13g2_decap_8 FILLER_80_1162 ();
 sg13g2_decap_4 FILLER_80_1169 ();
 sg13g2_fill_2 FILLER_80_1173 ();
 sg13g2_decap_8 FILLER_80_1179 ();
 sg13g2_fill_2 FILLER_80_1186 ();
 sg13g2_fill_1 FILLER_80_1188 ();
 sg13g2_decap_8 FILLER_80_1193 ();
 sg13g2_fill_2 FILLER_80_1200 ();
 sg13g2_fill_1 FILLER_80_1202 ();
 sg13g2_decap_8 FILLER_80_1207 ();
 sg13g2_decap_8 FILLER_80_1214 ();
 sg13g2_decap_8 FILLER_80_1221 ();
 sg13g2_decap_8 FILLER_80_1249 ();
 sg13g2_decap_8 FILLER_80_1256 ();
 sg13g2_fill_2 FILLER_80_1263 ();
 sg13g2_fill_1 FILLER_80_1265 ();
 sg13g2_fill_2 FILLER_80_1286 ();
 sg13g2_decap_8 FILLER_80_1296 ();
 sg13g2_decap_8 FILLER_80_1303 ();
 sg13g2_decap_4 FILLER_80_1310 ();
 sg13g2_decap_8 FILLER_80_1318 ();
 sg13g2_fill_1 FILLER_80_1325 ();
 sg13g2_decap_4 FILLER_80_1330 ();
 sg13g2_fill_1 FILLER_80_1334 ();
 sg13g2_decap_4 FILLER_80_1339 ();
 sg13g2_fill_1 FILLER_80_1343 ();
 sg13g2_decap_8 FILLER_80_1362 ();
 sg13g2_decap_8 FILLER_80_1369 ();
 sg13g2_decap_8 FILLER_80_1376 ();
 sg13g2_decap_8 FILLER_80_1383 ();
 sg13g2_fill_1 FILLER_80_1390 ();
 sg13g2_decap_8 FILLER_80_1399 ();
 sg13g2_decap_8 FILLER_80_1406 ();
 sg13g2_decap_8 FILLER_80_1413 ();
 sg13g2_decap_4 FILLER_80_1420 ();
 sg13g2_fill_1 FILLER_80_1424 ();
 sg13g2_fill_2 FILLER_80_1429 ();
 sg13g2_decap_8 FILLER_80_1441 ();
 sg13g2_fill_2 FILLER_80_1448 ();
 sg13g2_decap_4 FILLER_80_1454 ();
 sg13g2_decap_8 FILLER_80_1484 ();
 sg13g2_decap_4 FILLER_80_1491 ();
 sg13g2_fill_2 FILLER_80_1495 ();
 sg13g2_fill_2 FILLER_80_1501 ();
 sg13g2_decap_8 FILLER_80_1507 ();
 sg13g2_decap_8 FILLER_80_1514 ();
 sg13g2_decap_8 FILLER_80_1521 ();
 sg13g2_decap_8 FILLER_80_1528 ();
 sg13g2_decap_8 FILLER_80_1535 ();
 sg13g2_decap_8 FILLER_80_1542 ();
 sg13g2_decap_8 FILLER_80_1549 ();
 sg13g2_fill_2 FILLER_80_1556 ();
 sg13g2_fill_1 FILLER_80_1558 ();
 sg13g2_decap_8 FILLER_80_1563 ();
 sg13g2_decap_8 FILLER_80_1570 ();
 sg13g2_decap_8 FILLER_80_1577 ();
 sg13g2_decap_8 FILLER_80_1584 ();
 sg13g2_decap_8 FILLER_80_1591 ();
 sg13g2_decap_8 FILLER_80_1598 ();
 sg13g2_decap_8 FILLER_80_1605 ();
 sg13g2_decap_8 FILLER_80_1612 ();
 sg13g2_fill_2 FILLER_80_1619 ();
 sg13g2_fill_2 FILLER_80_1631 ();
 sg13g2_decap_8 FILLER_80_1637 ();
 sg13g2_decap_8 FILLER_80_1644 ();
 sg13g2_decap_8 FILLER_80_1651 ();
 sg13g2_decap_8 FILLER_80_1658 ();
 sg13g2_decap_8 FILLER_80_1665 ();
 sg13g2_decap_8 FILLER_80_1672 ();
 sg13g2_decap_4 FILLER_80_1679 ();
 sg13g2_fill_1 FILLER_80_1683 ();
 sg13g2_decap_8 FILLER_80_1697 ();
 sg13g2_decap_8 FILLER_80_1704 ();
 sg13g2_fill_2 FILLER_80_1711 ();
 sg13g2_fill_1 FILLER_80_1713 ();
 sg13g2_decap_4 FILLER_80_1718 ();
 sg13g2_decap_8 FILLER_80_1730 ();
 sg13g2_decap_8 FILLER_80_1737 ();
 sg13g2_decap_8 FILLER_80_1744 ();
 sg13g2_decap_8 FILLER_80_1751 ();
 sg13g2_fill_2 FILLER_80_1758 ();
 sg13g2_decap_8 FILLER_80_1768 ();
 sg13g2_decap_8 FILLER_80_1775 ();
 sg13g2_decap_8 FILLER_80_1782 ();
 sg13g2_decap_4 FILLER_80_1789 ();
 sg13g2_decap_8 FILLER_80_1797 ();
 sg13g2_decap_8 FILLER_80_1804 ();
 sg13g2_decap_8 FILLER_80_1811 ();
 sg13g2_decap_8 FILLER_80_1818 ();
 sg13g2_decap_8 FILLER_80_1825 ();
 sg13g2_decap_8 FILLER_80_1832 ();
 sg13g2_decap_8 FILLER_80_1839 ();
 sg13g2_decap_8 FILLER_80_1846 ();
 sg13g2_decap_8 FILLER_80_1853 ();
 sg13g2_decap_8 FILLER_80_1860 ();
 sg13g2_decap_8 FILLER_80_1867 ();
 sg13g2_decap_4 FILLER_80_1874 ();
 sg13g2_fill_1 FILLER_80_1878 ();
 sg13g2_decap_8 FILLER_80_1909 ();
 sg13g2_decap_8 FILLER_80_1920 ();
 sg13g2_fill_2 FILLER_80_1927 ();
 sg13g2_fill_1 FILLER_80_1929 ();
 sg13g2_decap_8 FILLER_80_1934 ();
 sg13g2_fill_1 FILLER_80_1941 ();
 sg13g2_decap_8 FILLER_80_1946 ();
 sg13g2_decap_8 FILLER_80_1953 ();
 sg13g2_decap_4 FILLER_80_1966 ();
 sg13g2_fill_1 FILLER_80_1970 ();
 sg13g2_decap_8 FILLER_80_1979 ();
 sg13g2_decap_8 FILLER_80_1986 ();
 sg13g2_decap_4 FILLER_80_1993 ();
 sg13g2_decap_8 FILLER_80_2001 ();
 sg13g2_decap_8 FILLER_80_2008 ();
 sg13g2_fill_2 FILLER_80_2015 ();
 sg13g2_decap_4 FILLER_80_2026 ();
 sg13g2_fill_1 FILLER_80_2030 ();
 sg13g2_decap_4 FILLER_80_2035 ();
 sg13g2_fill_2 FILLER_80_2039 ();
 sg13g2_decap_8 FILLER_80_2063 ();
 sg13g2_decap_8 FILLER_80_2070 ();
 sg13g2_fill_2 FILLER_80_2077 ();
 sg13g2_fill_2 FILLER_80_2086 ();
 sg13g2_fill_1 FILLER_80_2088 ();
 sg13g2_fill_1 FILLER_80_2145 ();
 sg13g2_fill_1 FILLER_80_2153 ();
 sg13g2_fill_1 FILLER_80_2164 ();
 sg13g2_fill_2 FILLER_80_2201 ();
 sg13g2_decap_8 FILLER_80_2207 ();
 sg13g2_decap_8 FILLER_80_2214 ();
 sg13g2_fill_1 FILLER_80_2221 ();
 sg13g2_decap_8 FILLER_80_2226 ();
 sg13g2_decap_8 FILLER_80_2233 ();
 sg13g2_decap_8 FILLER_80_2240 ();
 sg13g2_decap_8 FILLER_80_2247 ();
 sg13g2_decap_8 FILLER_80_2254 ();
 sg13g2_decap_8 FILLER_80_2261 ();
 sg13g2_decap_8 FILLER_80_2268 ();
 sg13g2_decap_8 FILLER_80_2275 ();
 sg13g2_decap_8 FILLER_80_2282 ();
 sg13g2_decap_8 FILLER_80_2289 ();
 sg13g2_decap_8 FILLER_80_2296 ();
 sg13g2_decap_8 FILLER_80_2303 ();
 sg13g2_fill_1 FILLER_80_2310 ();
 sg13g2_fill_2 FILLER_80_2324 ();
 sg13g2_decap_8 FILLER_80_2330 ();
 sg13g2_decap_8 FILLER_80_2337 ();
 sg13g2_decap_4 FILLER_80_2344 ();
 sg13g2_decap_8 FILLER_80_2374 ();
 sg13g2_decap_8 FILLER_80_2381 ();
 sg13g2_decap_8 FILLER_80_2388 ();
 sg13g2_decap_8 FILLER_80_2403 ();
 sg13g2_decap_8 FILLER_80_2410 ();
 sg13g2_decap_8 FILLER_80_2417 ();
 sg13g2_fill_2 FILLER_80_2424 ();
 sg13g2_fill_2 FILLER_80_2430 ();
 sg13g2_fill_1 FILLER_80_2432 ();
 sg13g2_decap_8 FILLER_80_2437 ();
 sg13g2_decap_4 FILLER_80_2444 ();
 sg13g2_decap_4 FILLER_80_2452 ();
 sg13g2_decap_4 FILLER_80_2464 ();
 sg13g2_decap_8 FILLER_80_2472 ();
 sg13g2_decap_4 FILLER_80_2479 ();
 sg13g2_fill_1 FILLER_80_2483 ();
 sg13g2_fill_1 FILLER_80_2488 ();
 sg13g2_fill_2 FILLER_80_2506 ();
 sg13g2_fill_1 FILLER_80_2512 ();
 sg13g2_decap_8 FILLER_80_2521 ();
 sg13g2_decap_8 FILLER_80_2528 ();
 sg13g2_decap_4 FILLER_80_2535 ();
 sg13g2_fill_2 FILLER_80_2539 ();
 sg13g2_decap_8 FILLER_80_2549 ();
 sg13g2_decap_8 FILLER_80_2556 ();
 sg13g2_decap_8 FILLER_80_2563 ();
 sg13g2_decap_8 FILLER_80_2570 ();
 sg13g2_decap_8 FILLER_80_2577 ();
 sg13g2_decap_8 FILLER_80_2584 ();
 sg13g2_decap_8 FILLER_80_2591 ();
 sg13g2_decap_8 FILLER_80_2598 ();
 sg13g2_decap_8 FILLER_80_2605 ();
 sg13g2_decap_8 FILLER_80_2612 ();
 sg13g2_decap_8 FILLER_80_2619 ();
 sg13g2_decap_8 FILLER_80_2626 ();
 sg13g2_decap_8 FILLER_80_2633 ();
 sg13g2_decap_8 FILLER_80_2640 ();
 sg13g2_decap_8 FILLER_80_2647 ();
 sg13g2_decap_8 FILLER_80_2654 ();
 sg13g2_decap_8 FILLER_80_2661 ();
 sg13g2_fill_2 FILLER_80_2668 ();
endmodule
