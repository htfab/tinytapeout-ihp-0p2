module tt_um_rejunity_vga_logo (clk,
    ena,
    rst_n,
    ui_in,
    uio_in,
    uio_oe,
    uio_out,
    uo_out);
 input clk;
 input ena;
 input rst_n;
 input [7:0] ui_in;
 input [7:0] uio_in;
 output [7:0] uio_oe;
 output [7:0] uio_out;
 output [7:0] uo_out;

 wire _0000_;
 wire _0001_;
 wire _0002_;
 wire _0003_;
 wire _0004_;
 wire _0005_;
 wire _0006_;
 wire _0007_;
 wire _0008_;
 wire _0009_;
 wire _0010_;
 wire _0011_;
 wire _0012_;
 wire _0013_;
 wire _0014_;
 wire _0015_;
 wire _0016_;
 wire _0017_;
 wire _0018_;
 wire _0019_;
 wire _0020_;
 wire _0021_;
 wire _0022_;
 wire _0023_;
 wire _0024_;
 wire _0025_;
 wire _0026_;
 wire _0027_;
 wire _0028_;
 wire _0029_;
 wire _0030_;
 wire _0031_;
 wire _0032_;
 wire _0033_;
 wire _0034_;
 wire _0035_;
 wire _0036_;
 wire _0037_;
 wire _0038_;
 wire _0039_;
 wire _0040_;
 wire _0041_;
 wire _0042_;
 wire _0043_;
 wire _0044_;
 wire _0045_;
 wire _0046_;
 wire _0047_;
 wire _0048_;
 wire _0049_;
 wire _0050_;
 wire _0051_;
 wire _0052_;
 wire _0053_;
 wire _0054_;
 wire _0055_;
 wire _0056_;
 wire _0057_;
 wire _0058_;
 wire _0059_;
 wire _0060_;
 wire _0061_;
 wire _0062_;
 wire _0063_;
 wire _0064_;
 wire _0065_;
 wire _0066_;
 wire _0067_;
 wire _0068_;
 wire _0069_;
 wire _0070_;
 wire _0071_;
 wire _0072_;
 wire _0073_;
 wire _0074_;
 wire _0075_;
 wire _0076_;
 wire _0077_;
 wire _0078_;
 wire _0079_;
 wire _0080_;
 wire _0081_;
 wire _0082_;
 wire _0083_;
 wire _0084_;
 wire _0085_;
 wire _0086_;
 wire _0087_;
 wire _0088_;
 wire _0089_;
 wire _0090_;
 wire _0091_;
 wire _0092_;
 wire _0093_;
 wire _0094_;
 wire _0095_;
 wire _0096_;
 wire _0097_;
 wire _0098_;
 wire _0099_;
 wire _0100_;
 wire _0101_;
 wire _0102_;
 wire _0103_;
 wire _0104_;
 wire _0105_;
 wire _0106_;
 wire _0107_;
 wire _0108_;
 wire _0109_;
 wire _0110_;
 wire _0111_;
 wire _0112_;
 wire _0113_;
 wire _0114_;
 wire _0115_;
 wire _0116_;
 wire _0117_;
 wire _0118_;
 wire _0119_;
 wire _0120_;
 wire _0121_;
 wire _0122_;
 wire _0123_;
 wire _0124_;
 wire _0125_;
 wire _0126_;
 wire _0127_;
 wire _0128_;
 wire _0129_;
 wire _0130_;
 wire _0131_;
 wire _0132_;
 wire _0133_;
 wire _0134_;
 wire _0135_;
 wire _0136_;
 wire _0137_;
 wire _0138_;
 wire _0139_;
 wire _0140_;
 wire _0141_;
 wire _0142_;
 wire _0143_;
 wire _0144_;
 wire _0145_;
 wire _0146_;
 wire _0147_;
 wire _0148_;
 wire _0149_;
 wire _0150_;
 wire _0151_;
 wire _0152_;
 wire _0153_;
 wire _0154_;
 wire _0155_;
 wire _0156_;
 wire _0157_;
 wire _0158_;
 wire _0159_;
 wire _0160_;
 wire _0161_;
 wire _0162_;
 wire _0163_;
 wire _0164_;
 wire _0165_;
 wire _0166_;
 wire _0167_;
 wire _0168_;
 wire _0169_;
 wire _0170_;
 wire _0171_;
 wire _0172_;
 wire _0173_;
 wire _0174_;
 wire _0175_;
 wire _0176_;
 wire _0177_;
 wire _0178_;
 wire _0179_;
 wire _0180_;
 wire _0181_;
 wire _0182_;
 wire _0183_;
 wire _0184_;
 wire _0185_;
 wire _0186_;
 wire _0187_;
 wire _0188_;
 wire _0189_;
 wire _0190_;
 wire _0191_;
 wire _0192_;
 wire _0193_;
 wire _0194_;
 wire _0195_;
 wire _0196_;
 wire _0197_;
 wire _0198_;
 wire _0199_;
 wire _0200_;
 wire _0201_;
 wire _0202_;
 wire _0203_;
 wire _0204_;
 wire _0205_;
 wire _0206_;
 wire _0207_;
 wire _0208_;
 wire _0209_;
 wire _0210_;
 wire _0211_;
 wire _0212_;
 wire _0213_;
 wire _0214_;
 wire _0215_;
 wire _0216_;
 wire _0217_;
 wire _0218_;
 wire _0219_;
 wire _0220_;
 wire _0221_;
 wire _0222_;
 wire _0223_;
 wire _0224_;
 wire _0225_;
 wire _0226_;
 wire _0227_;
 wire _0228_;
 wire _0229_;
 wire _0230_;
 wire _0231_;
 wire _0232_;
 wire _0233_;
 wire _0234_;
 wire _0235_;
 wire _0236_;
 wire _0237_;
 wire _0238_;
 wire _0239_;
 wire _0240_;
 wire _0241_;
 wire _0242_;
 wire _0243_;
 wire _0244_;
 wire _0245_;
 wire _0246_;
 wire _0247_;
 wire _0248_;
 wire _0249_;
 wire _0250_;
 wire _0251_;
 wire _0252_;
 wire _0253_;
 wire _0254_;
 wire _0255_;
 wire _0256_;
 wire _0257_;
 wire _0258_;
 wire _0259_;
 wire _0260_;
 wire _0261_;
 wire _0262_;
 wire _0263_;
 wire _0264_;
 wire _0265_;
 wire _0266_;
 wire _0267_;
 wire _0268_;
 wire _0269_;
 wire _0270_;
 wire _0271_;
 wire _0272_;
 wire _0273_;
 wire _0274_;
 wire _0275_;
 wire _0276_;
 wire _0277_;
 wire _0278_;
 wire _0279_;
 wire _0280_;
 wire _0281_;
 wire _0282_;
 wire _0283_;
 wire _0284_;
 wire _0285_;
 wire _0286_;
 wire _0287_;
 wire _0288_;
 wire _0289_;
 wire _0290_;
 wire _0291_;
 wire _0292_;
 wire _0293_;
 wire _0294_;
 wire _0295_;
 wire _0296_;
 wire _0297_;
 wire _0298_;
 wire _0299_;
 wire _0300_;
 wire _0301_;
 wire _0302_;
 wire _0303_;
 wire _0304_;
 wire _0305_;
 wire _0306_;
 wire _0307_;
 wire _0308_;
 wire _0309_;
 wire _0310_;
 wire _0311_;
 wire _0312_;
 wire _0313_;
 wire _0314_;
 wire _0315_;
 wire _0316_;
 wire _0317_;
 wire _0318_;
 wire _0319_;
 wire _0320_;
 wire _0321_;
 wire _0322_;
 wire _0323_;
 wire _0324_;
 wire _0325_;
 wire _0326_;
 wire _0327_;
 wire _0328_;
 wire _0329_;
 wire _0330_;
 wire _0331_;
 wire _0332_;
 wire _0333_;
 wire _0334_;
 wire _0335_;
 wire _0336_;
 wire _0337_;
 wire _0338_;
 wire _0339_;
 wire _0340_;
 wire _0341_;
 wire _0342_;
 wire _0343_;
 wire _0344_;
 wire _0345_;
 wire _0346_;
 wire _0347_;
 wire _0348_;
 wire _0349_;
 wire _0350_;
 wire _0351_;
 wire _0352_;
 wire _0353_;
 wire _0354_;
 wire _0355_;
 wire _0356_;
 wire _0357_;
 wire _0358_;
 wire _0359_;
 wire _0360_;
 wire _0361_;
 wire _0362_;
 wire _0363_;
 wire _0364_;
 wire _0365_;
 wire _0366_;
 wire _0367_;
 wire _0368_;
 wire _0369_;
 wire _0370_;
 wire _0371_;
 wire _0372_;
 wire _0373_;
 wire _0374_;
 wire _0375_;
 wire _0376_;
 wire _0377_;
 wire _0378_;
 wire _0379_;
 wire _0380_;
 wire _0381_;
 wire _0382_;
 wire _0383_;
 wire _0384_;
 wire _0385_;
 wire _0386_;
 wire _0387_;
 wire _0388_;
 wire _0389_;
 wire _0390_;
 wire _0391_;
 wire _0392_;
 wire _0393_;
 wire _0394_;
 wire _0395_;
 wire _0396_;
 wire _0397_;
 wire _0398_;
 wire _0399_;
 wire _0400_;
 wire _0401_;
 wire _0402_;
 wire _0403_;
 wire _0404_;
 wire _0405_;
 wire _0406_;
 wire _0407_;
 wire _0408_;
 wire _0409_;
 wire _0410_;
 wire _0411_;
 wire _0412_;
 wire _0413_;
 wire _0414_;
 wire _0415_;
 wire _0416_;
 wire _0417_;
 wire _0418_;
 wire _0419_;
 wire _0420_;
 wire _0421_;
 wire _0422_;
 wire _0423_;
 wire _0424_;
 wire _0425_;
 wire _0426_;
 wire _0427_;
 wire _0428_;
 wire _0429_;
 wire _0430_;
 wire _0431_;
 wire _0432_;
 wire _0433_;
 wire _0434_;
 wire _0435_;
 wire _0436_;
 wire _0437_;
 wire _0438_;
 wire _0439_;
 wire _0440_;
 wire _0441_;
 wire _0442_;
 wire _0443_;
 wire _0444_;
 wire _0445_;
 wire _0446_;
 wire _0447_;
 wire _0448_;
 wire _0449_;
 wire _0450_;
 wire _0451_;
 wire _0452_;
 wire _0453_;
 wire _0454_;
 wire _0455_;
 wire _0456_;
 wire _0457_;
 wire _0458_;
 wire _0459_;
 wire _0460_;
 wire _0461_;
 wire _0462_;
 wire _0463_;
 wire _0464_;
 wire _0465_;
 wire _0466_;
 wire _0467_;
 wire _0468_;
 wire _0469_;
 wire _0470_;
 wire _0471_;
 wire _0472_;
 wire _0473_;
 wire _0474_;
 wire _0475_;
 wire _0476_;
 wire _0477_;
 wire _0478_;
 wire _0479_;
 wire _0480_;
 wire _0481_;
 wire _0482_;
 wire _0483_;
 wire _0484_;
 wire _0485_;
 wire _0486_;
 wire _0487_;
 wire _0488_;
 wire _0489_;
 wire _0490_;
 wire _0491_;
 wire _0492_;
 wire _0493_;
 wire _0494_;
 wire _0495_;
 wire _0496_;
 wire _0497_;
 wire _0498_;
 wire _0499_;
 wire _0500_;
 wire _0501_;
 wire _0502_;
 wire _0503_;
 wire _0504_;
 wire _0505_;
 wire _0506_;
 wire _0507_;
 wire _0508_;
 wire _0509_;
 wire _0510_;
 wire _0511_;
 wire _0512_;
 wire _0513_;
 wire _0514_;
 wire _0515_;
 wire _0516_;
 wire _0517_;
 wire _0518_;
 wire _0519_;
 wire _0520_;
 wire _0521_;
 wire _0522_;
 wire _0523_;
 wire _0524_;
 wire _0525_;
 wire _0526_;
 wire _0527_;
 wire _0528_;
 wire _0529_;
 wire _0530_;
 wire _0531_;
 wire _0532_;
 wire _0533_;
 wire _0534_;
 wire _0535_;
 wire _0536_;
 wire _0537_;
 wire _0538_;
 wire _0539_;
 wire _0540_;
 wire _0541_;
 wire _0542_;
 wire _0543_;
 wire _0544_;
 wire _0545_;
 wire _0546_;
 wire _0547_;
 wire _0548_;
 wire _0549_;
 wire _0550_;
 wire _0551_;
 wire _0552_;
 wire _0553_;
 wire _0554_;
 wire _0555_;
 wire _0556_;
 wire _0557_;
 wire _0558_;
 wire _0559_;
 wire _0560_;
 wire _0561_;
 wire _0562_;
 wire _0563_;
 wire _0564_;
 wire _0565_;
 wire _0566_;
 wire _0567_;
 wire _0568_;
 wire _0569_;
 wire _0570_;
 wire _0571_;
 wire _0572_;
 wire _0573_;
 wire _0574_;
 wire _0575_;
 wire _0576_;
 wire _0577_;
 wire _0578_;
 wire _0579_;
 wire _0580_;
 wire _0581_;
 wire _0582_;
 wire _0583_;
 wire _0584_;
 wire _0585_;
 wire _0586_;
 wire _0587_;
 wire _0588_;
 wire _0589_;
 wire _0590_;
 wire _0591_;
 wire _0592_;
 wire _0593_;
 wire _0594_;
 wire _0595_;
 wire _0596_;
 wire _0597_;
 wire _0598_;
 wire _0599_;
 wire _0600_;
 wire _0601_;
 wire _0602_;
 wire _0603_;
 wire _0604_;
 wire _0605_;
 wire _0606_;
 wire _0607_;
 wire _0608_;
 wire _0609_;
 wire _0610_;
 wire _0611_;
 wire _0612_;
 wire _0613_;
 wire _0614_;
 wire _0615_;
 wire _0616_;
 wire _0617_;
 wire _0618_;
 wire _0619_;
 wire _0620_;
 wire _0621_;
 wire _0622_;
 wire _0623_;
 wire _0624_;
 wire _0625_;
 wire _0626_;
 wire _0627_;
 wire _0628_;
 wire _0629_;
 wire _0630_;
 wire _0631_;
 wire _0632_;
 wire _0633_;
 wire _0634_;
 wire _0635_;
 wire _0636_;
 wire _0637_;
 wire _0638_;
 wire _0639_;
 wire _0640_;
 wire _0641_;
 wire _0642_;
 wire _0643_;
 wire _0644_;
 wire _0645_;
 wire _0646_;
 wire _0647_;
 wire _0648_;
 wire _0649_;
 wire _0650_;
 wire _0651_;
 wire _0652_;
 wire _0653_;
 wire _0654_;
 wire _0655_;
 wire _0656_;
 wire _0657_;
 wire _0658_;
 wire _0659_;
 wire _0660_;
 wire _0661_;
 wire _0662_;
 wire _0663_;
 wire _0664_;
 wire _0665_;
 wire _0666_;
 wire _0667_;
 wire _0668_;
 wire _0669_;
 wire _0670_;
 wire _0671_;
 wire _0672_;
 wire _0673_;
 wire _0674_;
 wire _0675_;
 wire _0676_;
 wire _0677_;
 wire _0678_;
 wire _0679_;
 wire _0680_;
 wire _0681_;
 wire _0682_;
 wire _0683_;
 wire _0684_;
 wire _0685_;
 wire _0686_;
 wire _0687_;
 wire _0688_;
 wire _0689_;
 wire _0690_;
 wire _0691_;
 wire _0692_;
 wire _0693_;
 wire _0694_;
 wire _0695_;
 wire _0696_;
 wire _0697_;
 wire _0698_;
 wire _0699_;
 wire _0700_;
 wire _0701_;
 wire _0702_;
 wire _0703_;
 wire _0704_;
 wire _0705_;
 wire _0706_;
 wire _0707_;
 wire _0708_;
 wire _0709_;
 wire _0710_;
 wire _0711_;
 wire _0712_;
 wire _0713_;
 wire _0714_;
 wire _0715_;
 wire _0716_;
 wire _0717_;
 wire _0718_;
 wire _0719_;
 wire _0720_;
 wire _0721_;
 wire _0722_;
 wire _0723_;
 wire _0724_;
 wire _0725_;
 wire _0726_;
 wire _0727_;
 wire _0728_;
 wire _0729_;
 wire _0730_;
 wire _0731_;
 wire _0732_;
 wire _0733_;
 wire _0734_;
 wire _0735_;
 wire _0736_;
 wire _0737_;
 wire _0738_;
 wire _0739_;
 wire _0740_;
 wire _0741_;
 wire _0742_;
 wire _0743_;
 wire _0744_;
 wire _0745_;
 wire _0746_;
 wire _0747_;
 wire _0748_;
 wire _0749_;
 wire _0750_;
 wire _0751_;
 wire _0752_;
 wire _0753_;
 wire _0754_;
 wire _0755_;
 wire _0756_;
 wire _0757_;
 wire _0758_;
 wire _0759_;
 wire _0760_;
 wire _0761_;
 wire _0762_;
 wire _0763_;
 wire _0764_;
 wire _0765_;
 wire _0766_;
 wire _0767_;
 wire _0768_;
 wire _0769_;
 wire _0770_;
 wire _0771_;
 wire _0772_;
 wire _0773_;
 wire _0774_;
 wire _0775_;
 wire _0776_;
 wire _0777_;
 wire _0778_;
 wire _0779_;
 wire _0780_;
 wire _0781_;
 wire _0782_;
 wire _0783_;
 wire _0784_;
 wire _0785_;
 wire _0786_;
 wire _0787_;
 wire _0788_;
 wire _0789_;
 wire _0790_;
 wire _0791_;
 wire _0792_;
 wire _0793_;
 wire _0794_;
 wire _0795_;
 wire _0796_;
 wire _0797_;
 wire _0798_;
 wire _0799_;
 wire _0800_;
 wire _0801_;
 wire _0802_;
 wire _0803_;
 wire _0804_;
 wire _0805_;
 wire _0806_;
 wire _0807_;
 wire _0808_;
 wire _0809_;
 wire _0810_;
 wire _0811_;
 wire _0812_;
 wire _0813_;
 wire _0814_;
 wire _0815_;
 wire _0816_;
 wire _0817_;
 wire _0818_;
 wire _0819_;
 wire _0820_;
 wire _0821_;
 wire _0822_;
 wire _0823_;
 wire _0824_;
 wire _0825_;
 wire _0826_;
 wire _0827_;
 wire _0828_;
 wire _0829_;
 wire _0830_;
 wire _0831_;
 wire _0832_;
 wire _0833_;
 wire _0834_;
 wire _0835_;
 wire _0836_;
 wire _0837_;
 wire _0838_;
 wire _0839_;
 wire _0840_;
 wire _0841_;
 wire _0842_;
 wire _0843_;
 wire _0844_;
 wire _0845_;
 wire _0846_;
 wire _0847_;
 wire _0848_;
 wire _0849_;
 wire _0850_;
 wire _0851_;
 wire _0852_;
 wire _0853_;
 wire _0854_;
 wire _0855_;
 wire _0856_;
 wire _0857_;
 wire _0858_;
 wire _0859_;
 wire _0860_;
 wire _0861_;
 wire _0862_;
 wire _0863_;
 wire _0864_;
 wire _0865_;
 wire _0866_;
 wire _0867_;
 wire _0868_;
 wire _0869_;
 wire _0870_;
 wire _0871_;
 wire _0872_;
 wire _0873_;
 wire _0874_;
 wire _0875_;
 wire _0876_;
 wire _0877_;
 wire _0878_;
 wire _0879_;
 wire _0880_;
 wire _0881_;
 wire _0882_;
 wire _0883_;
 wire _0884_;
 wire _0885_;
 wire _0886_;
 wire _0887_;
 wire _0888_;
 wire _0889_;
 wire _0890_;
 wire _0891_;
 wire _0892_;
 wire _0893_;
 wire _0894_;
 wire _0895_;
 wire _0896_;
 wire _0897_;
 wire _0898_;
 wire _0899_;
 wire _0900_;
 wire _0901_;
 wire _0902_;
 wire _0903_;
 wire _0904_;
 wire _0905_;
 wire _0906_;
 wire _0907_;
 wire _0908_;
 wire _0909_;
 wire _0910_;
 wire _0911_;
 wire _0912_;
 wire _0913_;
 wire _0914_;
 wire _0915_;
 wire _0916_;
 wire _0917_;
 wire _0918_;
 wire _0919_;
 wire _0920_;
 wire _0921_;
 wire _0922_;
 wire _0923_;
 wire _0924_;
 wire _0925_;
 wire _0926_;
 wire _0927_;
 wire _0928_;
 wire _0929_;
 wire _0930_;
 wire _0931_;
 wire _0932_;
 wire _0933_;
 wire _0934_;
 wire _0935_;
 wire _0936_;
 wire _0937_;
 wire _0938_;
 wire _0939_;
 wire _0940_;
 wire _0941_;
 wire _0942_;
 wire _0943_;
 wire _0944_;
 wire _0945_;
 wire _0946_;
 wire _0947_;
 wire _0948_;
 wire _0949_;
 wire _0950_;
 wire _0951_;
 wire _0952_;
 wire _0953_;
 wire _0954_;
 wire _0955_;
 wire _0956_;
 wire _0957_;
 wire _0958_;
 wire _0959_;
 wire _0960_;
 wire _0961_;
 wire _0962_;
 wire _0963_;
 wire _0964_;
 wire _0965_;
 wire _0966_;
 wire _0967_;
 wire _0968_;
 wire _0969_;
 wire _0970_;
 wire _0971_;
 wire _0972_;
 wire _0973_;
 wire _0974_;
 wire _0975_;
 wire _0976_;
 wire _0977_;
 wire _0978_;
 wire _0979_;
 wire _0980_;
 wire _0981_;
 wire _0982_;
 wire _0983_;
 wire _0984_;
 wire _0985_;
 wire _0986_;
 wire _0987_;
 wire _0988_;
 wire _0989_;
 wire _0990_;
 wire _0991_;
 wire _0992_;
 wire _0993_;
 wire _0994_;
 wire _0995_;
 wire _0996_;
 wire _0997_;
 wire _0998_;
 wire _0999_;
 wire _1000_;
 wire _1001_;
 wire _1002_;
 wire _1003_;
 wire _1004_;
 wire _1005_;
 wire _1006_;
 wire _1007_;
 wire _1008_;
 wire _1009_;
 wire _1010_;
 wire _1011_;
 wire _1012_;
 wire _1013_;
 wire _1014_;
 wire _1015_;
 wire _1016_;
 wire _1017_;
 wire _1018_;
 wire _1019_;
 wire _1020_;
 wire _1021_;
 wire _1022_;
 wire _1023_;
 wire _1024_;
 wire _1025_;
 wire _1026_;
 wire _1027_;
 wire _1028_;
 wire _1029_;
 wire _1030_;
 wire _1031_;
 wire _1032_;
 wire _1033_;
 wire _1034_;
 wire _1035_;
 wire _1036_;
 wire _1037_;
 wire _1038_;
 wire _1039_;
 wire _1040_;
 wire _1041_;
 wire _1042_;
 wire _1043_;
 wire _1044_;
 wire _1045_;
 wire _1046_;
 wire _1047_;
 wire _1048_;
 wire _1049_;
 wire _1050_;
 wire _1051_;
 wire _1052_;
 wire _1053_;
 wire _1054_;
 wire _1055_;
 wire _1056_;
 wire _1057_;
 wire _1058_;
 wire _1059_;
 wire _1060_;
 wire _1061_;
 wire _1062_;
 wire _1063_;
 wire _1064_;
 wire _1065_;
 wire _1066_;
 wire _1067_;
 wire _1068_;
 wire _1069_;
 wire _1070_;
 wire _1071_;
 wire _1072_;
 wire _1073_;
 wire _1074_;
 wire _1075_;
 wire _1076_;
 wire _1077_;
 wire _1078_;
 wire _1079_;
 wire _1080_;
 wire _1081_;
 wire _1082_;
 wire _1083_;
 wire _1084_;
 wire _1085_;
 wire _1086_;
 wire _1087_;
 wire _1088_;
 wire _1089_;
 wire _1090_;
 wire _1091_;
 wire _1092_;
 wire _1093_;
 wire _1094_;
 wire _1095_;
 wire _1096_;
 wire _1097_;
 wire _1098_;
 wire _1099_;
 wire _1100_;
 wire _1101_;
 wire _1102_;
 wire _1103_;
 wire _1104_;
 wire _1105_;
 wire _1106_;
 wire _1107_;
 wire _1108_;
 wire _1109_;
 wire _1110_;
 wire _1111_;
 wire _1112_;
 wire _1113_;
 wire _1114_;
 wire _1115_;
 wire _1116_;
 wire _1117_;
 wire _1118_;
 wire _1119_;
 wire _1120_;
 wire _1121_;
 wire _1122_;
 wire _1123_;
 wire _1124_;
 wire _1125_;
 wire _1126_;
 wire _1127_;
 wire _1128_;
 wire _1129_;
 wire _1130_;
 wire _1131_;
 wire _1132_;
 wire _1133_;
 wire _1134_;
 wire _1135_;
 wire _1136_;
 wire _1137_;
 wire _1138_;
 wire _1139_;
 wire _1140_;
 wire _1141_;
 wire _1142_;
 wire _1143_;
 wire _1144_;
 wire _1145_;
 wire _1146_;
 wire _1147_;
 wire _1148_;
 wire _1149_;
 wire _1150_;
 wire _1151_;
 wire _1152_;
 wire _1153_;
 wire _1154_;
 wire _1155_;
 wire _1156_;
 wire _1157_;
 wire _1158_;
 wire _1159_;
 wire _1160_;
 wire _1161_;
 wire _1162_;
 wire _1163_;
 wire _1164_;
 wire _1165_;
 wire _1166_;
 wire _1167_;
 wire _1168_;
 wire _1169_;
 wire _1170_;
 wire _1171_;
 wire _1172_;
 wire _1173_;
 wire _1174_;
 wire _1175_;
 wire _1176_;
 wire _1177_;
 wire _1178_;
 wire _1179_;
 wire _1180_;
 wire _1181_;
 wire _1182_;
 wire _1183_;
 wire _1184_;
 wire _1185_;
 wire _1186_;
 wire _1187_;
 wire _1188_;
 wire _1189_;
 wire _1190_;
 wire _1191_;
 wire _1192_;
 wire _1193_;
 wire _1194_;
 wire _1195_;
 wire _1196_;
 wire _1197_;
 wire _1198_;
 wire _1199_;
 wire _1200_;
 wire _1201_;
 wire _1202_;
 wire _1203_;
 wire _1204_;
 wire _1205_;
 wire _1206_;
 wire _1207_;
 wire _1208_;
 wire _1209_;
 wire _1210_;
 wire _1211_;
 wire _1212_;
 wire _1213_;
 wire _1214_;
 wire _1215_;
 wire _1216_;
 wire _1217_;
 wire _1218_;
 wire _1219_;
 wire _1220_;
 wire _1221_;
 wire _1222_;
 wire _1223_;
 wire _1224_;
 wire _1225_;
 wire _1226_;
 wire _1227_;
 wire _1228_;
 wire _1229_;
 wire _1230_;
 wire _1231_;
 wire _1232_;
 wire _1233_;
 wire _1234_;
 wire _1235_;
 wire _1236_;
 wire _1237_;
 wire _1238_;
 wire _1239_;
 wire _1240_;
 wire _1241_;
 wire _1242_;
 wire _1243_;
 wire _1244_;
 wire _1245_;
 wire _1246_;
 wire _1247_;
 wire _1248_;
 wire _1249_;
 wire _1250_;
 wire _1251_;
 wire _1252_;
 wire _1253_;
 wire _1254_;
 wire _1255_;
 wire _1256_;
 wire _1257_;
 wire _1258_;
 wire _1259_;
 wire _1260_;
 wire _1261_;
 wire _1262_;
 wire clknet_0_clk;
 wire net92;
 wire \counter[0] ;
 wire \counter[1] ;
 wire \counter[2] ;
 wire \counter[3] ;
 wire \counter[4] ;
 wire \counter[5] ;
 wire \grad1.acc[0] ;
 wire \grad1.acc[1] ;
 wire \grad1.acc[2] ;
 wire \grad1.acc[3] ;
 wire \grad1.acc[4] ;
 wire \grad1.acc[5] ;
 wire \grad1.acc[6] ;
 wire \grad1.acc[7] ;
 wire \grad1.acc[8] ;
 wire \grad1.lfsr[0] ;
 wire \grad1.lfsr[10] ;
 wire \grad1.lfsr[11] ;
 wire \grad1.lfsr[12] ;
 wire \grad1.lfsr[13] ;
 wire \grad1.lfsr[14] ;
 wire \grad1.lfsr[15] ;
 wire \grad1.lfsr[16] ;
 wire \grad1.lfsr[17] ;
 wire \grad1.lfsr[18] ;
 wire \grad1.lfsr[19] ;
 wire \grad1.lfsr[1] ;
 wire \grad1.lfsr[2] ;
 wire \grad1.lfsr[3] ;
 wire \grad1.lfsr[4] ;
 wire \grad1.lfsr[5] ;
 wire \grad1.lfsr[6] ;
 wire \grad1.lfsr[7] ;
 wire \grad1.lfsr[8] ;
 wire \grad1.lfsr[9] ;
 wire hsync;
 wire \hvsync_gen.hpos[0] ;
 wire \hvsync_gen.hpos[1] ;
 wire \hvsync_gen.hpos[2] ;
 wire \hvsync_gen.hpos[3] ;
 wire \hvsync_gen.hpos[4] ;
 wire \hvsync_gen.hpos[5] ;
 wire \hvsync_gen.hpos[6] ;
 wire \hvsync_gen.hpos[7] ;
 wire \hvsync_gen.hpos[8] ;
 wire \hvsync_gen.hpos[9] ;
 wire \hvsync_gen.vpos[0] ;
 wire \hvsync_gen.vpos[1] ;
 wire \hvsync_gen.vpos[2] ;
 wire \hvsync_gen.vpos[3] ;
 wire \hvsync_gen.vpos[4] ;
 wire \hvsync_gen.vpos[5] ;
 wire \hvsync_gen.vpos[6] ;
 wire \hvsync_gen.vpos[7] ;
 wire \hvsync_gen.vpos[8] ;
 wire \hvsync_gen.vpos[9] ;
 wire \hvsync_gen.vsync ;
 wire \r[0] ;
 wire \r[10] ;
 wire \r[11] ;
 wire \r[12] ;
 wire \r[13] ;
 wire \r[14] ;
 wire \r[15] ;
 wire \r[16] ;
 wire \r[1] ;
 wire \r[2] ;
 wire \r[3] ;
 wire \r[4] ;
 wire \r[5] ;
 wire \r[6] ;
 wire \r[7] ;
 wire \r[8] ;
 wire \r[9] ;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire clknet_4_0_0_clk;
 wire clknet_4_1_0_clk;
 wire clknet_4_2_0_clk;
 wire clknet_4_3_0_clk;
 wire clknet_4_4_0_clk;
 wire clknet_4_5_0_clk;
 wire clknet_4_6_0_clk;
 wire clknet_4_7_0_clk;
 wire clknet_4_8_0_clk;
 wire clknet_4_9_0_clk;
 wire clknet_4_10_0_clk;
 wire clknet_4_11_0_clk;
 wire clknet_4_12_0_clk;
 wire clknet_4_13_0_clk;
 wire clknet_4_14_0_clk;
 wire clknet_4_15_0_clk;

 sg13g2_dfrbp_1 \UO_OUT[0]$_SDFF_PN0_  (.CLK(clknet_4_13_0_clk),
    .RESET_B(net92),
    .D(_0077_),
    .Q_N(_1259_),
    .Q(net2));
 sg13g2_dfrbp_1 \UO_OUT[1]$_SDFF_PN0_  (.CLK(clknet_4_13_0_clk),
    .RESET_B(net93),
    .D(_0078_),
    .Q_N(_1258_),
    .Q(net3));
 sg13g2_dfrbp_1 \UO_OUT[2]$_SDFF_PN0_  (.CLK(clknet_4_13_0_clk),
    .RESET_B(net94),
    .D(_0079_),
    .Q_N(_1260_),
    .Q(net4));
 sg13g2_dfrbp_1 \UO_OUT[3]$_DFF_P_  (.CLK(clknet_4_13_0_clk),
    .RESET_B(net95),
    .D(\hvsync_gen.vsync ),
    .Q_N(_1257_),
    .Q(net5));
 sg13g2_dfrbp_1 \UO_OUT[4]$_SDFF_PN0_  (.CLK(clknet_4_13_0_clk),
    .RESET_B(net96),
    .D(_0080_),
    .Q_N(_1256_),
    .Q(net6));
 sg13g2_dfrbp_1 \UO_OUT[5]$_SDFF_PN0_  (.CLK(clknet_4_7_0_clk),
    .RESET_B(net97),
    .D(_0081_),
    .Q_N(_1255_),
    .Q(net7));
 sg13g2_dfrbp_1 \UO_OUT[6]$_SDFF_PN0_  (.CLK(clknet_4_12_0_clk),
    .RESET_B(net98),
    .D(_0082_),
    .Q_N(_1261_),
    .Q(net8));
 sg13g2_dfrbp_1 \UO_OUT[7]$_DFF_P_  (.CLK(clknet_4_3_0_clk),
    .RESET_B(net99),
    .D(hsync),
    .Q_N(_1254_),
    .Q(net9));
 sg13g2_buf_1 _1265_ (.A(\hvsync_gen.vpos[9] ),
    .X(_0435_));
 sg13g2_buf_1 _1266_ (.A(_0435_),
    .X(_0436_));
 sg13g2_buf_1 _1267_ (.A(\hvsync_gen.vpos[3] ),
    .X(_0437_));
 sg13g2_buf_1 _1268_ (.A(net73),
    .X(_0438_));
 sg13g2_buf_1 _1269_ (.A(\hvsync_gen.vpos[2] ),
    .X(_0439_));
 sg13g2_buf_1 _1270_ (.A(net72),
    .X(_0440_));
 sg13g2_inv_1 _1271_ (.Y(_0441_),
    .A(net49));
 sg13g2_buf_1 _1272_ (.A(\hvsync_gen.vpos[1] ),
    .X(_0442_));
 sg13g2_buf_1 _1273_ (.A(\hvsync_gen.vpos[0] ),
    .X(_0443_));
 sg13g2_nand2_1 _1274_ (.Y(_0444_),
    .A(net71),
    .B(net70));
 sg13g2_nand2_1 _1275_ (.Y(_0445_),
    .A(_0441_),
    .B(_0444_));
 sg13g2_buf_2 _1276_ (.A(\hvsync_gen.vpos[4] ),
    .X(_0446_));
 sg13g2_buf_1 _1277_ (.A(_0446_),
    .X(_0447_));
 sg13g2_buf_1 _1278_ (.A(net48),
    .X(_0448_));
 sg13g2_inv_2 _1279_ (.Y(_0449_),
    .A(_0442_));
 sg13g2_nor4_1 _1280_ (.A(net51),
    .B(net28),
    .C(_0449_),
    .D(net70),
    .Y(_0450_));
 sg13g2_a21oi_1 _1281_ (.A1(_0438_),
    .A2(_0445_),
    .Y(_0451_),
    .B1(_0450_));
 sg13g2_buf_8 _1282_ (.A(\hvsync_gen.vpos[6] ),
    .X(_0452_));
 sg13g2_buf_1 _1283_ (.A(_0452_),
    .X(_0453_));
 sg13g2_buf_1 _1284_ (.A(net47),
    .X(_0454_));
 sg13g2_buf_2 _1285_ (.A(\hvsync_gen.vpos[5] ),
    .X(_0455_));
 sg13g2_buf_1 _1286_ (.A(_0455_),
    .X(_0456_));
 sg13g2_buf_1 _1287_ (.A(net46),
    .X(_0457_));
 sg13g2_buf_2 _1288_ (.A(\hvsync_gen.vpos[8] ),
    .X(_0458_));
 sg13g2_buf_1 _1289_ (.A(_0458_),
    .X(_0459_));
 sg13g2_buf_2 _1290_ (.A(\hvsync_gen.vpos[7] ),
    .X(_0460_));
 sg13g2_buf_1 _1291_ (.A(_0460_),
    .X(_0461_));
 sg13g2_and2_1 _1292_ (.A(net45),
    .B(net44),
    .X(_0462_));
 sg13g2_nand3_1 _1293_ (.B(net26),
    .C(_0462_),
    .A(net27),
    .Y(_0463_));
 sg13g2_nand2_2 _1294_ (.Y(_0464_),
    .A(net46),
    .B(net48));
 sg13g2_nand3_1 _1295_ (.B(_0441_),
    .C(_0464_),
    .A(net50),
    .Y(_0465_));
 sg13g2_nor4_1 _1296_ (.A(net51),
    .B(_0451_),
    .C(_0463_),
    .D(_0465_),
    .Y(_0001_));
 sg13g2_buf_1 _1297_ (.A(_0008_),
    .X(_0466_));
 sg13g2_buf_1 _1298_ (.A(_0466_),
    .X(_0467_));
 sg13g2_inv_1 _1299_ (.Y(_0468_),
    .A(net43));
 sg13g2_buf_1 _1300_ (.A(\hvsync_gen.hpos[7] ),
    .X(_0469_));
 sg13g2_buf_1 _1301_ (.A(\hvsync_gen.hpos[6] ),
    .X(_0470_));
 sg13g2_nand2_2 _1302_ (.Y(_0471_),
    .A(net69),
    .B(net68));
 sg13g2_buf_8 _1303_ (.A(\hvsync_gen.hpos[4] ),
    .X(_0472_));
 sg13g2_buf_1 _1304_ (.A(_0472_),
    .X(_0473_));
 sg13g2_buf_1 _1305_ (.A(\hvsync_gen.hpos[5] ),
    .X(_0474_));
 sg13g2_buf_1 _1306_ (.A(_0474_),
    .X(_0475_));
 sg13g2_nand2_1 _1307_ (.Y(_0476_),
    .A(net42),
    .B(net41));
 sg13g2_buf_2 _1308_ (.A(\hvsync_gen.hpos[8] ),
    .X(_0477_));
 sg13g2_inv_1 _1309_ (.Y(_0478_),
    .A(_0477_));
 sg13g2_buf_1 _1310_ (.A(_0478_),
    .X(_0479_));
 sg13g2_o21ai_1 _1311_ (.B1(net25),
    .Y(_0480_),
    .A1(_0471_),
    .A2(_0476_));
 sg13g2_buf_1 _1312_ (.A(net68),
    .X(_0481_));
 sg13g2_inv_2 _1313_ (.Y(_0482_),
    .A(net42));
 sg13g2_inv_1 _1314_ (.Y(_0483_),
    .A(_0474_));
 sg13g2_nand2_1 _1315_ (.Y(_0484_),
    .A(_0482_),
    .B(net39));
 sg13g2_o21ai_1 _1316_ (.B1(_0469_),
    .Y(_0485_),
    .A1(net40),
    .A2(_0484_));
 sg13g2_buf_1 _1317_ (.A(\hvsync_gen.hpos[9] ),
    .X(_0486_));
 sg13g2_inv_2 _1318_ (.Y(_0487_),
    .A(_0486_));
 sg13g2_a221oi_1 _1319_ (.B2(net25),
    .C1(_0487_),
    .B1(_0485_),
    .A1(_0468_),
    .Y(_0000_),
    .A2(_0480_));
 sg13g2_inv_2 _1320_ (.Y(_0488_),
    .A(net1));
 sg13g2_buf_1 _1321_ (.A(\hvsync_gen.hpos[1] ),
    .X(_0489_));
 sg13g2_buf_1 _1322_ (.A(_0489_),
    .X(_0490_));
 sg13g2_buf_1 _1323_ (.A(\hvsync_gen.hpos[0] ),
    .X(_0491_));
 sg13g2_buf_1 _1324_ (.A(_0491_),
    .X(_0492_));
 sg13g2_nand2_1 _1325_ (.Y(_0493_),
    .A(net38),
    .B(net37));
 sg13g2_buf_1 _1326_ (.A(\hvsync_gen.hpos[3] ),
    .X(_0494_));
 sg13g2_buf_1 _1327_ (.A(net67),
    .X(_0495_));
 sg13g2_buf_2 _1328_ (.A(\hvsync_gen.hpos[2] ),
    .X(_0496_));
 sg13g2_buf_1 _1329_ (.A(_0496_),
    .X(_0497_));
 sg13g2_nand2_1 _1330_ (.Y(_0498_),
    .A(net36),
    .B(net35));
 sg13g2_nor2_1 _1331_ (.A(_0493_),
    .B(_0498_),
    .Y(_0499_));
 sg13g2_nand2_1 _1332_ (.Y(_0500_),
    .A(net42),
    .B(_0499_));
 sg13g2_or2_1 _1333_ (.X(_0501_),
    .B(net68),
    .A(\hvsync_gen.hpos[7] ));
 sg13g2_buf_2 _1334_ (.A(_0501_),
    .X(_0502_));
 sg13g2_nand2_2 _1335_ (.Y(_0503_),
    .A(_0477_),
    .B(_0486_));
 sg13g2_nor4_2 _1336_ (.A(net41),
    .B(_0500_),
    .C(_0502_),
    .Y(_0504_),
    .D(_0503_));
 sg13g2_nor2_2 _1337_ (.A(_0488_),
    .B(_0504_),
    .Y(_0505_));
 sg13g2_buf_1 _1338_ (.A(net1),
    .X(_0506_));
 sg13g2_nor3_1 _1339_ (.A(net48),
    .B(net71),
    .C(_0443_),
    .Y(_0507_));
 sg13g2_inv_2 _1340_ (.Y(_0508_),
    .A(net47));
 sg13g2_inv_2 _1341_ (.Y(_0509_),
    .A(net46));
 sg13g2_nand3_1 _1342_ (.B(_0508_),
    .C(_0509_),
    .A(net51),
    .Y(_0510_));
 sg13g2_nand2_1 _1343_ (.Y(_0511_),
    .A(net50),
    .B(net49));
 sg13g2_or2_1 _1344_ (.X(_0512_),
    .B(net44),
    .A(net45));
 sg13g2_nor3_1 _1345_ (.A(_0510_),
    .B(_0511_),
    .C(_0512_),
    .Y(_0513_));
 sg13g2_nand2_1 _1346_ (.Y(_0514_),
    .A(_0507_),
    .B(_0513_));
 sg13g2_nand2_1 _1347_ (.Y(_0515_),
    .A(net75),
    .B(_0514_));
 sg13g2_nor2_1 _1348_ (.A(_0505_),
    .B(_0515_),
    .Y(_0516_));
 sg13g2_a22oi_1 _1349_ (.Y(_0517_),
    .B1(_0516_),
    .B2(_0023_),
    .A2(_0505_),
    .A1(net70));
 sg13g2_inv_1 _1350_ (.Y(_0050_),
    .A(_0517_));
 sg13g2_buf_1 _1351_ (.A(_0488_),
    .X(_0518_));
 sg13g2_nand2_1 _1352_ (.Y(_0519_),
    .A(net70),
    .B(_0504_));
 sg13g2_xnor2_1 _1353_ (.Y(_0520_),
    .A(_0449_),
    .B(_0519_));
 sg13g2_nor2_1 _1354_ (.A(net66),
    .B(_0520_),
    .Y(_0051_));
 sg13g2_nand2b_1 _1355_ (.Y(_0521_),
    .B(_0516_),
    .A_N(_0444_));
 sg13g2_nor2b_1 _1356_ (.A(_0515_),
    .B_N(_0444_),
    .Y(_0522_));
 sg13g2_o21ai_1 _1357_ (.B1(net49),
    .Y(_0523_),
    .A1(_0505_),
    .A2(_0522_));
 sg13g2_o21ai_1 _1358_ (.B1(_0523_),
    .Y(_0052_),
    .A1(net49),
    .A2(_0521_));
 sg13g2_nand2b_2 _1359_ (.Y(_0524_),
    .B(net75),
    .A_N(_0504_));
 sg13g2_nand3_1 _1360_ (.B(net71),
    .C(net70),
    .A(net49),
    .Y(_0525_));
 sg13g2_nand3_1 _1361_ (.B(_0514_),
    .C(_0525_),
    .A(net75),
    .Y(_0526_));
 sg13g2_inv_1 _1362_ (.Y(_0527_),
    .A(_0437_));
 sg13g2_a21oi_1 _1363_ (.A1(_0524_),
    .A2(_0526_),
    .Y(_0528_),
    .B1(_0527_));
 sg13g2_nor4_1 _1364_ (.A(net50),
    .B(_0505_),
    .C(_0515_),
    .D(_0525_),
    .Y(_0529_));
 sg13g2_or2_1 _1365_ (.X(_0053_),
    .B(_0529_),
    .A(_0528_));
 sg13g2_and2_1 _1366_ (.A(_0524_),
    .B(_0515_),
    .X(_0530_));
 sg13g2_buf_1 _1367_ (.A(_0530_),
    .X(_0531_));
 sg13g2_nor3_2 _1368_ (.A(_0444_),
    .B(_0505_),
    .C(_0511_),
    .Y(_0532_));
 sg13g2_xnor2_1 _1369_ (.Y(_0533_),
    .A(net28),
    .B(_0532_));
 sg13g2_nor2_1 _1370_ (.A(_0531_),
    .B(_0533_),
    .Y(_0054_));
 sg13g2_nand2_1 _1371_ (.Y(_0534_),
    .A(net28),
    .B(_0532_));
 sg13g2_xnor2_1 _1372_ (.Y(_0535_),
    .A(_0509_),
    .B(_0534_));
 sg13g2_nor2_1 _1373_ (.A(_0531_),
    .B(_0535_),
    .Y(_0055_));
 sg13g2_inv_1 _1374_ (.Y(_0536_),
    .A(net28));
 sg13g2_nor2_2 _1375_ (.A(_0509_),
    .B(_0536_),
    .Y(_0537_));
 sg13g2_nand2_1 _1376_ (.Y(_0538_),
    .A(_0537_),
    .B(_0532_));
 sg13g2_xnor2_1 _1377_ (.Y(_0539_),
    .A(_0508_),
    .B(_0538_));
 sg13g2_nor2_1 _1378_ (.A(_0531_),
    .B(_0539_),
    .Y(_0056_));
 sg13g2_inv_2 _1379_ (.Y(_0540_),
    .A(_0460_));
 sg13g2_nand3_1 _1380_ (.B(_0537_),
    .C(_0532_),
    .A(net27),
    .Y(_0541_));
 sg13g2_xnor2_1 _1381_ (.Y(_0542_),
    .A(_0540_),
    .B(_0541_));
 sg13g2_nor2_1 _1382_ (.A(_0531_),
    .B(_0542_),
    .Y(_0057_));
 sg13g2_nand4_1 _1383_ (.B(net27),
    .C(_0537_),
    .A(net44),
    .Y(_0543_),
    .D(_0532_));
 sg13g2_xor2_1 _1384_ (.B(_0543_),
    .A(net45),
    .X(_0544_));
 sg13g2_nor2_1 _1385_ (.A(_0531_),
    .B(_0544_),
    .Y(_0058_));
 sg13g2_nand2_1 _1386_ (.Y(_0545_),
    .A(net27),
    .B(_0462_));
 sg13g2_nor2_1 _1387_ (.A(_0545_),
    .B(_0538_),
    .Y(_0546_));
 sg13g2_xnor2_1 _1388_ (.Y(_0547_),
    .A(net51),
    .B(_0546_));
 sg13g2_nor2_1 _1389_ (.A(_0531_),
    .B(_0547_),
    .Y(_0059_));
 sg13g2_and2_1 _1390_ (.A(_0022_),
    .B(_0505_),
    .X(_0040_));
 sg13g2_xnor2_1 _1391_ (.Y(_0548_),
    .A(net38),
    .B(net37));
 sg13g2_nor2_1 _1392_ (.A(net66),
    .B(_0548_),
    .Y(_0041_));
 sg13g2_xor2_1 _1393_ (.B(_0493_),
    .A(net35),
    .X(_0549_));
 sg13g2_nor2_1 _1394_ (.A(net66),
    .B(_0549_),
    .Y(_0042_));
 sg13g2_nand3_1 _1395_ (.B(net37),
    .C(net35),
    .A(net38),
    .Y(_0550_));
 sg13g2_xor2_1 _1396_ (.B(_0550_),
    .A(net36),
    .X(_0551_));
 sg13g2_nor2_1 _1397_ (.A(net66),
    .B(_0551_),
    .Y(_0043_));
 sg13g2_xnor2_1 _1398_ (.Y(_0552_),
    .A(_0473_),
    .B(_0499_));
 sg13g2_nor2_1 _1399_ (.A(net66),
    .B(_0552_),
    .Y(_0044_));
 sg13g2_xnor2_1 _1400_ (.Y(_0553_),
    .A(net39),
    .B(_0500_));
 sg13g2_nor2_1 _1401_ (.A(_0524_),
    .B(_0553_),
    .Y(_0045_));
 sg13g2_nor4_2 _1402_ (.A(_0482_),
    .B(net39),
    .C(_0493_),
    .Y(_0554_),
    .D(_0498_));
 sg13g2_xnor2_1 _1403_ (.Y(_0555_),
    .A(net40),
    .B(_0554_));
 sg13g2_nor2_1 _1404_ (.A(_0524_),
    .B(_0555_),
    .Y(_0046_));
 sg13g2_buf_1 _1405_ (.A(net75),
    .X(_0556_));
 sg13g2_nand2_1 _1406_ (.Y(_0557_),
    .A(net40),
    .B(_0554_));
 sg13g2_xnor2_1 _1407_ (.Y(_0558_),
    .A(net69),
    .B(_0557_));
 sg13g2_and2_1 _1408_ (.A(net65),
    .B(_0558_),
    .X(_0047_));
 sg13g2_nand2b_1 _1409_ (.Y(_0559_),
    .B(_0554_),
    .A_N(_0471_));
 sg13g2_xnor2_1 _1410_ (.Y(_0560_),
    .A(net25),
    .B(_0559_));
 sg13g2_nor2_1 _1411_ (.A(_0524_),
    .B(_0560_),
    .Y(_0048_));
 sg13g2_or2_1 _1412_ (.X(_0561_),
    .B(_0559_),
    .A(net25));
 sg13g2_xnor2_1 _1413_ (.Y(_0562_),
    .A(_0487_),
    .B(_0561_));
 sg13g2_nor2_1 _1414_ (.A(_0524_),
    .B(_0562_),
    .Y(_0049_));
 sg13g2_and2_1 _1415_ (.A(net65),
    .B(\grad1.lfsr[14] ),
    .X(_0026_));
 sg13g2_and2_1 _1416_ (.A(_0556_),
    .B(\grad1.lfsr[15] ),
    .X(_0027_));
 sg13g2_and2_1 _1417_ (.A(net65),
    .B(\grad1.lfsr[16] ),
    .X(_0028_));
 sg13g2_and2_1 _1418_ (.A(net65),
    .B(\grad1.lfsr[17] ),
    .X(_0029_));
 sg13g2_and2_1 _1419_ (.A(net65),
    .B(\grad1.lfsr[18] ),
    .X(_0030_));
 sg13g2_and2_1 _1420_ (.A(_0556_),
    .B(\grad1.lfsr[0] ),
    .X(_0031_));
 sg13g2_and2_1 _1421_ (.A(net65),
    .B(\grad1.lfsr[1] ),
    .X(_0032_));
 sg13g2_and2_1 _1422_ (.A(net65),
    .B(\grad1.lfsr[2] ),
    .X(_0033_));
 sg13g2_inv_1 _1423_ (.Y(_0563_),
    .A(\grad1.lfsr[3] ));
 sg13g2_nor2_1 _1424_ (.A(net66),
    .B(_0563_),
    .Y(_0034_));
 sg13g2_buf_1 _1425_ (.A(\grad1.lfsr[4] ),
    .X(_0564_));
 sg13g2_and2_1 _1426_ (.A(net65),
    .B(_0564_),
    .X(_0035_));
 sg13g2_inv_1 _1427_ (.Y(_0565_),
    .A(\grad1.lfsr[5] ));
 sg13g2_nor2_1 _1428_ (.A(net66),
    .B(_0565_),
    .Y(_0036_));
 sg13g2_inv_1 _1429_ (.Y(_0566_),
    .A(\grad1.lfsr[6] ));
 sg13g2_nor2_1 _1430_ (.A(net66),
    .B(_0566_),
    .Y(_0037_));
 sg13g2_buf_1 _1431_ (.A(net75),
    .X(_0567_));
 sg13g2_and2_1 _1432_ (.A(net64),
    .B(\grad1.lfsr[7] ),
    .X(_0038_));
 sg13g2_and2_1 _1433_ (.A(net64),
    .B(\grad1.lfsr[8] ),
    .X(_0039_));
 sg13g2_buf_2 _1434_ (.A(\r[0] ),
    .X(_0568_));
 sg13g2_buf_1 _1435_ (.A(_0477_),
    .X(_0569_));
 sg13g2_buf_1 _1436_ (.A(_0486_),
    .X(_0570_));
 sg13g2_o21ai_1 _1437_ (.B1(net33),
    .Y(_0571_),
    .A1(net34),
    .A2(net69));
 sg13g2_nand3b_1 _1438_ (.B(_0463_),
    .C(_0571_),
    .Y(_0572_),
    .A_N(net51));
 sg13g2_buf_1 _1439_ (.A(_0572_),
    .X(_0573_));
 sg13g2_nor2b_1 _1440_ (.A(net74),
    .B_N(_0573_),
    .Y(_0574_));
 sg13g2_buf_2 _1441_ (.A(_0574_),
    .X(_0575_));
 sg13g2_buf_1 _1442_ (.A(net22),
    .X(_0576_));
 sg13g2_nor2_1 _1443_ (.A(_0568_),
    .B(net20),
    .Y(_0577_));
 sg13g2_a21oi_1 _1444_ (.A1(_0568_),
    .A2(_0575_),
    .Y(_0578_),
    .B1(_0577_));
 sg13g2_nor2_1 _1445_ (.A(_0518_),
    .B(_0578_),
    .Y(_0060_));
 sg13g2_nor4_1 _1446_ (.A(net38),
    .B(_0492_),
    .C(net36),
    .D(net35),
    .Y(_0579_));
 sg13g2_nor4_1 _1447_ (.A(_0569_),
    .B(net33),
    .C(_0484_),
    .D(_0502_),
    .Y(_0580_));
 sg13g2_nand2_1 _1448_ (.Y(_0581_),
    .A(_0579_),
    .B(_0580_));
 sg13g2_buf_1 _1449_ (.A(_0581_),
    .X(_0582_));
 sg13g2_nor2_1 _1450_ (.A(net22),
    .B(net19),
    .Y(_0583_));
 sg13g2_buf_1 _1451_ (.A(_0583_),
    .X(_0584_));
 sg13g2_buf_2 _1452_ (.A(_0003_),
    .X(_0585_));
 sg13g2_nand4_1 _1453_ (.B(net47),
    .C(net46),
    .A(_0460_),
    .Y(_0586_),
    .D(_0446_));
 sg13g2_buf_2 _1454_ (.A(_0586_),
    .X(_0587_));
 sg13g2_o21ai_1 _1455_ (.B1(_0013_),
    .Y(_0588_),
    .A1(_0458_),
    .A2(_0587_));
 sg13g2_xor2_1 _1456_ (.B(_0588_),
    .A(_0435_),
    .X(_0589_));
 sg13g2_xor2_1 _1457_ (.B(_0589_),
    .A(_0585_),
    .X(_0590_));
 sg13g2_inv_1 _1458_ (.Y(_0591_),
    .A(\r[9] ));
 sg13g2_buf_2 _1459_ (.A(\r[3] ),
    .X(_0592_));
 sg13g2_buf_1 _1460_ (.A(\r[2] ),
    .X(_0593_));
 sg13g2_nor2_1 _1461_ (.A(net71),
    .B(net63),
    .Y(_0594_));
 sg13g2_buf_2 _1462_ (.A(\r[1] ),
    .X(_0595_));
 sg13g2_nor2_2 _1463_ (.A(_0595_),
    .B(_0568_),
    .Y(_0596_));
 sg13g2_a21oi_1 _1464_ (.A1(_0595_),
    .A2(_0568_),
    .Y(_0597_),
    .B1(net70));
 sg13g2_nor3_1 _1465_ (.A(_0594_),
    .B(_0596_),
    .C(_0597_),
    .Y(_0598_));
 sg13g2_a221oi_1 _1466_ (.B2(net71),
    .C1(_0598_),
    .B1(net63),
    .A1(_0439_),
    .Y(_0599_),
    .A2(_0592_));
 sg13g2_nor2_1 _1467_ (.A(_0439_),
    .B(_0592_),
    .Y(_0600_));
 sg13g2_buf_2 _1468_ (.A(\r[4] ),
    .X(_0601_));
 sg13g2_nand2_1 _1469_ (.Y(_0602_),
    .A(net73),
    .B(_0601_));
 sg13g2_o21ai_1 _1470_ (.B1(_0602_),
    .Y(_0603_),
    .A1(_0599_),
    .A2(_0600_));
 sg13g2_nor2_1 _1471_ (.A(net73),
    .B(_0601_),
    .Y(_0604_));
 sg13g2_buf_2 _1472_ (.A(_0012_),
    .X(_0605_));
 sg13g2_xor2_1 _1473_ (.B(_0002_),
    .A(_0605_),
    .X(_0606_));
 sg13g2_and3_1 _1474_ (.X(_0607_),
    .A(net46),
    .B(net48),
    .C(\r[7] ));
 sg13g2_a21o_1 _1475_ (.A2(net48),
    .A1(net46),
    .B1(\r[7] ),
    .X(_0608_));
 sg13g2_o21ai_1 _1476_ (.B1(_0608_),
    .Y(_0609_),
    .A1(net47),
    .A2(_0607_));
 sg13g2_and2_1 _1477_ (.A(_0606_),
    .B(_0609_),
    .X(_0610_));
 sg13g2_nand3_1 _1478_ (.B(net46),
    .C(net48),
    .A(net47),
    .Y(_0611_));
 sg13g2_nor2_1 _1479_ (.A(_0611_),
    .B(_0606_),
    .Y(_0612_));
 sg13g2_inv_1 _1480_ (.Y(_0613_),
    .A(\r[6] ));
 sg13g2_nand2_1 _1481_ (.Y(_0614_),
    .A(net48),
    .B(\r[5] ));
 sg13g2_nand3_1 _1482_ (.B(_0613_),
    .C(_0614_),
    .A(_0509_),
    .Y(_0615_));
 sg13g2_buf_1 _1483_ (.A(\r[6] ),
    .X(_0616_));
 sg13g2_and2_1 _1484_ (.A(net62),
    .B(\r[5] ),
    .X(_0617_));
 sg13g2_a21oi_1 _1485_ (.A1(_0464_),
    .A2(_0615_),
    .Y(_0618_),
    .B1(_0617_));
 sg13g2_nor4_1 _1486_ (.A(_0604_),
    .B(_0610_),
    .C(_0612_),
    .D(_0618_),
    .Y(_0619_));
 sg13g2_or2_1 _1487_ (.X(_0620_),
    .B(\r[5] ),
    .A(_0447_));
 sg13g2_a21oi_1 _1488_ (.A1(net62),
    .A2(_0620_),
    .Y(_0621_),
    .B1(_0456_));
 sg13g2_buf_1 _1489_ (.A(\r[5] ),
    .X(_0622_));
 sg13g2_o21ai_1 _1490_ (.B1(_0464_),
    .Y(_0623_),
    .A1(net62),
    .A2(net61));
 sg13g2_nor2_1 _1491_ (.A(_0621_),
    .B(_0623_),
    .Y(_0624_));
 sg13g2_a21oi_1 _1492_ (.A1(_0606_),
    .A2(_0609_),
    .Y(_0625_),
    .B1(_0612_));
 sg13g2_mux2_1 _1493_ (.A0(_0464_),
    .A1(_0607_),
    .S(_0606_),
    .X(_0626_));
 sg13g2_buf_1 _1494_ (.A(\r[7] ),
    .X(_0627_));
 sg13g2_a21oi_1 _1495_ (.A1(_0456_),
    .A2(_0447_),
    .Y(_0628_),
    .B1(net60));
 sg13g2_nor3_1 _1496_ (.A(_0453_),
    .B(_0606_),
    .C(_0628_),
    .Y(_0629_));
 sg13g2_a21o_1 _1497_ (.A2(_0626_),
    .A1(_0453_),
    .B1(_0629_),
    .X(_0630_));
 sg13g2_a21o_1 _1498_ (.A2(_0625_),
    .A1(_0624_),
    .B1(_0630_),
    .X(_0631_));
 sg13g2_a21o_1 _1499_ (.A2(_0619_),
    .A1(_0603_),
    .B1(_0631_),
    .X(_0632_));
 sg13g2_buf_1 _1500_ (.A(_0632_),
    .X(_0633_));
 sg13g2_buf_1 _1501_ (.A(\r[8] ),
    .X(_0634_));
 sg13g2_inv_2 _1502_ (.Y(_0635_),
    .A(_0605_));
 sg13g2_xnor2_1 _1503_ (.Y(_0636_),
    .A(_0635_),
    .B(_0611_));
 sg13g2_or2_1 _1504_ (.X(_0637_),
    .B(_0636_),
    .A(_0634_));
 sg13g2_xor2_1 _1505_ (.B(_0587_),
    .A(net45),
    .X(_0638_));
 sg13g2_or2_1 _1506_ (.X(_0639_),
    .B(_0638_),
    .A(_0637_));
 sg13g2_and2_1 _1507_ (.A(_0637_),
    .B(_0638_),
    .X(_0640_));
 sg13g2_a21oi_1 _1508_ (.A1(_0633_),
    .A2(_0639_),
    .Y(_0641_),
    .B1(_0640_));
 sg13g2_nand2_1 _1509_ (.Y(_0642_),
    .A(_0637_),
    .B(_0638_));
 sg13g2_nor2_1 _1510_ (.A(_0591_),
    .B(_0642_),
    .Y(_0643_));
 sg13g2_nor2_1 _1511_ (.A(_0633_),
    .B(_0639_),
    .Y(_0644_));
 sg13g2_a221oi_1 _1512_ (.B2(_0633_),
    .C1(_0644_),
    .B1(_0643_),
    .A1(_0591_),
    .Y(_0645_),
    .A2(_0641_));
 sg13g2_xnor2_1 _1513_ (.Y(_0646_),
    .A(_0590_),
    .B(_0645_));
 sg13g2_nand2_1 _1514_ (.Y(_0647_),
    .A(net12),
    .B(_0646_));
 sg13g2_buf_1 _1515_ (.A(\r[10] ),
    .X(_0648_));
 sg13g2_nor2b_1 _1516_ (.A(net22),
    .B_N(net19),
    .Y(_0649_));
 sg13g2_buf_2 _1517_ (.A(_0649_),
    .X(_0650_));
 sg13g2_xor2_1 _1518_ (.B(\r[10] ),
    .A(_0466_),
    .X(_0651_));
 sg13g2_nor2_2 _1519_ (.A(_0469_),
    .B(net68),
    .Y(_0652_));
 sg13g2_and2_1 _1520_ (.A(net38),
    .B(net63),
    .X(_0653_));
 sg13g2_nor2_1 _1521_ (.A(net38),
    .B(net63),
    .Y(_0654_));
 sg13g2_a21oi_1 _1522_ (.A1(_0595_),
    .A2(_0568_),
    .Y(_0655_),
    .B1(_0491_));
 sg13g2_nor3_1 _1523_ (.A(_0596_),
    .B(_0654_),
    .C(_0655_),
    .Y(_0656_));
 sg13g2_nand2_1 _1524_ (.Y(_0657_),
    .A(_0494_),
    .B(_0601_));
 sg13g2_nand2_1 _1525_ (.Y(_0658_),
    .A(net35),
    .B(_0592_));
 sg13g2_nand2_1 _1526_ (.Y(_0659_),
    .A(_0657_),
    .B(_0658_));
 sg13g2_nor3_1 _1527_ (.A(_0653_),
    .B(_0656_),
    .C(_0659_),
    .Y(_0660_));
 sg13g2_nor2_1 _1528_ (.A(net35),
    .B(_0592_),
    .Y(_0661_));
 sg13g2_nor2_1 _1529_ (.A(_0494_),
    .B(_0601_),
    .Y(_0662_));
 sg13g2_a21oi_1 _1530_ (.A1(_0657_),
    .A2(_0661_),
    .Y(_0663_),
    .B1(_0662_));
 sg13g2_inv_1 _1531_ (.Y(_0664_),
    .A(_0663_));
 sg13g2_nor2_2 _1532_ (.A(_0660_),
    .B(_0664_),
    .Y(_0665_));
 sg13g2_xor2_1 _1533_ (.B(_0634_),
    .A(\hvsync_gen.hpos[7] ),
    .X(_0666_));
 sg13g2_or2_1 _1534_ (.X(_0667_),
    .B(_0666_),
    .A(net68));
 sg13g2_nor2_1 _1535_ (.A(net41),
    .B(net62),
    .Y(_0668_));
 sg13g2_nor2_1 _1536_ (.A(_0472_),
    .B(net61),
    .Y(_0669_));
 sg13g2_nor3_1 _1537_ (.A(_0667_),
    .B(_0668_),
    .C(_0669_),
    .Y(_0670_));
 sg13g2_nand2_1 _1538_ (.Y(_0671_),
    .A(_0665_),
    .B(_0670_));
 sg13g2_or2_1 _1539_ (.X(_0672_),
    .B(\r[6] ),
    .A(_0474_));
 sg13g2_nand3_1 _1540_ (.B(_0666_),
    .C(_0672_),
    .A(net68),
    .Y(_0673_));
 sg13g2_nand2_1 _1541_ (.Y(_0674_),
    .A(net41),
    .B(net62));
 sg13g2_and2_1 _1542_ (.A(_0470_),
    .B(_0674_),
    .X(_0675_));
 sg13g2_inv_1 _1543_ (.Y(_0676_),
    .A(_0627_));
 sg13g2_a221oi_1 _1544_ (.B2(_0675_),
    .C1(_0676_),
    .B1(_0669_),
    .A1(_0667_),
    .Y(_0677_),
    .A2(_0673_));
 sg13g2_nand2_1 _1545_ (.Y(_0678_),
    .A(_0470_),
    .B(_0674_));
 sg13g2_a21oi_1 _1546_ (.A1(net42),
    .A2(net61),
    .Y(_0679_),
    .B1(_0678_));
 sg13g2_o21ai_1 _1547_ (.B1(_0679_),
    .Y(_0680_),
    .A1(_0660_),
    .A2(_0664_));
 sg13g2_nand3_1 _1548_ (.B(net61),
    .C(_0672_),
    .A(_0472_),
    .Y(_0681_));
 sg13g2_a21oi_1 _1549_ (.A1(_0674_),
    .A2(_0681_),
    .Y(_0682_),
    .B1(_0667_));
 sg13g2_a21oi_1 _1550_ (.A1(_0471_),
    .A2(_0502_),
    .Y(_0683_),
    .B1(_0002_));
 sg13g2_or2_1 _1551_ (.X(_0684_),
    .B(_0683_),
    .A(_0682_));
 sg13g2_a21oi_1 _1552_ (.A1(_0677_),
    .A2(_0680_),
    .Y(_0685_),
    .B1(_0684_));
 sg13g2_and2_1 _1553_ (.A(_0671_),
    .B(_0685_),
    .X(_0686_));
 sg13g2_buf_1 _1554_ (.A(_0686_),
    .X(_0687_));
 sg13g2_and2_1 _1555_ (.A(_0591_),
    .B(_0687_),
    .X(_0688_));
 sg13g2_buf_1 _1556_ (.A(\r[9] ),
    .X(_0689_));
 sg13g2_nor2_2 _1557_ (.A(_0478_),
    .B(_0652_),
    .Y(_0690_));
 sg13g2_nand2_1 _1558_ (.Y(_0691_),
    .A(net58),
    .B(_0690_));
 sg13g2_a21oi_1 _1559_ (.A1(_0671_),
    .A2(_0685_),
    .Y(_0692_),
    .B1(_0691_));
 sg13g2_a21oi_1 _1560_ (.A1(_0652_),
    .A2(_0688_),
    .Y(_0693_),
    .B1(_0692_));
 sg13g2_nor2_1 _1561_ (.A(_0591_),
    .B(_0687_),
    .Y(_0694_));
 sg13g2_nor2_1 _1562_ (.A(_0502_),
    .B(_0694_),
    .Y(_0695_));
 sg13g2_o21ai_1 _1563_ (.B1(net25),
    .Y(_0696_),
    .A1(_0688_),
    .A2(_0695_));
 sg13g2_nand2_1 _1564_ (.Y(_0697_),
    .A(_0693_),
    .B(_0696_));
 sg13g2_xnor2_1 _1565_ (.Y(_0698_),
    .A(_0651_),
    .B(_0697_));
 sg13g2_a22oi_1 _1566_ (.Y(_0699_),
    .B1(_0650_),
    .B2(_0698_),
    .A2(_0575_),
    .A1(net59));
 sg13g2_buf_1 _1567_ (.A(_0488_),
    .X(_0700_));
 sg13g2_a21oi_1 _1568_ (.A1(_0647_),
    .A2(_0699_),
    .Y(_0061_),
    .B1(net57));
 sg13g2_buf_1 _1569_ (.A(\r[11] ),
    .X(_0701_));
 sg13g2_buf_1 _1570_ (.A(_0701_),
    .X(_0702_));
 sg13g2_or2_1 _1571_ (.X(_0703_),
    .B(net19),
    .A(net22));
 sg13g2_buf_2 _1572_ (.A(_0703_),
    .X(_0704_));
 sg13g2_nor2_1 _1573_ (.A(_0591_),
    .B(_0590_),
    .Y(_0705_));
 sg13g2_nor3_1 _1574_ (.A(_0634_),
    .B(_0636_),
    .C(_0638_),
    .Y(_0706_));
 sg13g2_nor2_1 _1575_ (.A(_0590_),
    .B(_0706_),
    .Y(_0707_));
 sg13g2_o21ai_1 _1576_ (.B1(_0633_),
    .Y(_0708_),
    .A1(_0705_),
    .A2(_0707_));
 sg13g2_nand2b_1 _1577_ (.Y(_0709_),
    .B(\r[9] ),
    .A_N(_0706_));
 sg13g2_a21oi_1 _1578_ (.A1(_0642_),
    .A2(_0709_),
    .Y(_0710_),
    .B1(_0590_));
 sg13g2_a21oi_1 _1579_ (.A1(_0633_),
    .A2(_0643_),
    .Y(_0711_),
    .B1(_0710_));
 sg13g2_nand2_1 _1580_ (.Y(_0712_),
    .A(_0708_),
    .B(_0711_));
 sg13g2_nor2_2 _1581_ (.A(_0459_),
    .B(_0436_),
    .Y(_0713_));
 sg13g2_and2_1 _1582_ (.A(_0587_),
    .B(_0713_),
    .X(_0714_));
 sg13g2_buf_1 _1583_ (.A(_0714_),
    .X(_0715_));
 sg13g2_buf_1 _1584_ (.A(_0715_),
    .X(_0716_));
 sg13g2_nor2b_1 _1585_ (.A(_0648_),
    .B_N(_0589_),
    .Y(_0717_));
 sg13g2_xnor2_1 _1586_ (.Y(_0718_),
    .A(net18),
    .B(_0717_));
 sg13g2_xnor2_1 _1587_ (.Y(_0719_),
    .A(_0712_),
    .B(_0718_));
 sg13g2_nand2b_1 _1588_ (.Y(_0720_),
    .B(_0573_),
    .A_N(net74));
 sg13g2_buf_1 _1589_ (.A(_0720_),
    .X(_0721_));
 sg13g2_o21ai_1 _1590_ (.B1(net16),
    .Y(_0722_),
    .A1(_0704_),
    .A2(_0719_));
 sg13g2_nor2_1 _1591_ (.A(net32),
    .B(_0704_),
    .Y(_0723_));
 sg13g2_nand2b_1 _1592_ (.Y(_0724_),
    .B(net19),
    .A_N(net22));
 sg13g2_buf_1 _1593_ (.A(_0724_),
    .X(_0725_));
 sg13g2_xnor2_1 _1594_ (.Y(_0726_),
    .A(net43),
    .B(_0690_));
 sg13g2_nor2_1 _1595_ (.A(_0585_),
    .B(_0726_),
    .Y(_0727_));
 sg13g2_nor2b_1 _1596_ (.A(_0651_),
    .B_N(_0692_),
    .Y(_0728_));
 sg13g2_xnor2_1 _1597_ (.Y(_0729_),
    .A(net34),
    .B(_0652_));
 sg13g2_nand3_1 _1598_ (.B(_0651_),
    .C(_0729_),
    .A(net58),
    .Y(_0730_));
 sg13g2_inv_1 _1599_ (.Y(_0731_),
    .A(_0730_));
 sg13g2_nand2_1 _1600_ (.Y(_0732_),
    .A(_0651_),
    .B(_0729_));
 sg13g2_nand3_1 _1601_ (.B(net58),
    .C(_0651_),
    .A(_0479_),
    .Y(_0733_));
 sg13g2_a21oi_1 _1602_ (.A1(_0732_),
    .A2(_0733_),
    .Y(_0734_),
    .B1(_0687_));
 sg13g2_or4_1 _1603_ (.A(_0727_),
    .B(_0728_),
    .C(_0731_),
    .D(_0734_),
    .X(_0735_));
 sg13g2_buf_1 _1604_ (.A(_0735_),
    .X(_0736_));
 sg13g2_buf_1 _1605_ (.A(_0004_),
    .X(_0737_));
 sg13g2_buf_1 _1606_ (.A(_0737_),
    .X(_0738_));
 sg13g2_nand2_2 _1607_ (.Y(_0739_),
    .A(_0477_),
    .B(_0502_));
 sg13g2_o21ai_1 _1608_ (.B1(net43),
    .Y(_0740_),
    .A1(_0570_),
    .A2(_0739_));
 sg13g2_buf_1 _1609_ (.A(_0740_),
    .X(_0741_));
 sg13g2_xor2_1 _1610_ (.B(net21),
    .A(net31),
    .X(_0742_));
 sg13g2_xnor2_1 _1611_ (.Y(_0743_),
    .A(net59),
    .B(_0739_));
 sg13g2_and4_1 _1612_ (.A(_0487_),
    .B(net43),
    .C(net59),
    .D(_0690_),
    .X(_0744_));
 sg13g2_a21oi_1 _1613_ (.A1(_0468_),
    .A2(_0743_),
    .Y(_0745_),
    .B1(_0744_));
 sg13g2_nand3_1 _1614_ (.B(net59),
    .C(_0690_),
    .A(_0570_),
    .Y(_0746_));
 sg13g2_o21ai_1 _1615_ (.B1(_0746_),
    .Y(_0747_),
    .A1(net59),
    .A2(_0690_));
 sg13g2_nand3_1 _1616_ (.B(net31),
    .C(_0747_),
    .A(net43),
    .Y(_0748_));
 sg13g2_o21ai_1 _1617_ (.B1(_0748_),
    .Y(_0749_),
    .A1(net31),
    .A2(_0745_));
 sg13g2_inv_1 _1618_ (.Y(_0750_),
    .A(_0729_));
 sg13g2_a21oi_1 _1619_ (.A1(_0591_),
    .A2(_0687_),
    .Y(_0751_),
    .B1(_0750_));
 sg13g2_or2_1 _1620_ (.X(_0752_),
    .B(_0751_),
    .A(_0694_));
 sg13g2_nand3_1 _1621_ (.B(net31),
    .C(_0739_),
    .A(_0467_),
    .Y(_0753_));
 sg13g2_or3_1 _1622_ (.A(_0467_),
    .B(_0737_),
    .C(_0739_),
    .X(_0754_));
 sg13g2_a21oi_1 _1623_ (.A1(_0753_),
    .A2(_0754_),
    .Y(_0755_),
    .B1(_0585_));
 sg13g2_a21oi_1 _1624_ (.A1(_0749_),
    .A2(_0752_),
    .Y(_0756_),
    .B1(_0755_));
 sg13g2_o21ai_1 _1625_ (.B1(_0756_),
    .Y(_0757_),
    .A1(_0736_),
    .A2(_0742_));
 sg13g2_nor2_1 _1626_ (.A(net11),
    .B(_0757_),
    .Y(_0758_));
 sg13g2_a221oi_1 _1627_ (.B2(_0719_),
    .C1(_0758_),
    .B1(_0723_),
    .A1(net32),
    .Y(_0759_),
    .A2(_0722_));
 sg13g2_nor2_1 _1628_ (.A(_0518_),
    .B(_0759_),
    .Y(_0062_));
 sg13g2_buf_1 _1629_ (.A(\r[12] ),
    .X(_0760_));
 sg13g2_nand3_1 _1630_ (.B(_0711_),
    .C(_0717_),
    .A(_0708_),
    .Y(_0761_));
 sg13g2_buf_1 _1631_ (.A(_0761_),
    .X(_0762_));
 sg13g2_nand2_2 _1632_ (.Y(_0763_),
    .A(_0587_),
    .B(_0713_));
 sg13g2_a21o_1 _1633_ (.A2(_0711_),
    .A1(_0708_),
    .B1(_0717_),
    .X(_0764_));
 sg13g2_buf_1 _1634_ (.A(_0764_),
    .X(_0765_));
 sg13g2_nand3_1 _1635_ (.B(_0763_),
    .C(_0765_),
    .A(net32),
    .Y(_0766_));
 sg13g2_nand2_1 _1636_ (.Y(_0767_),
    .A(_0762_),
    .B(_0766_));
 sg13g2_mux2_1 _1637_ (.A0(_0762_),
    .A1(_0765_),
    .S(net18),
    .X(_0768_));
 sg13g2_and2_1 _1638_ (.A(_0762_),
    .B(_0765_),
    .X(_0769_));
 sg13g2_a22oi_1 _1639_ (.Y(_0770_),
    .B1(_0769_),
    .B2(net32),
    .A2(_0763_),
    .A1(net31));
 sg13g2_a22oi_1 _1640_ (.Y(_0771_),
    .B1(_0768_),
    .B2(_0770_),
    .A2(_0767_),
    .A1(net31));
 sg13g2_a21oi_1 _1641_ (.A1(net12),
    .A2(_0771_),
    .Y(_0772_),
    .B1(_0575_));
 sg13g2_nor2_1 _1642_ (.A(net56),
    .B(_0772_),
    .Y(_0773_));
 sg13g2_inv_1 _1643_ (.Y(_0774_),
    .A(net56));
 sg13g2_nor3_1 _1644_ (.A(_0774_),
    .B(_0704_),
    .C(_0771_),
    .Y(_0775_));
 sg13g2_buf_2 _1645_ (.A(_0005_),
    .X(_0776_));
 sg13g2_nor2_1 _1646_ (.A(_0702_),
    .B(net21),
    .Y(_0777_));
 sg13g2_mux2_1 _1647_ (.A0(net21),
    .A1(_0777_),
    .S(_0756_),
    .X(_0778_));
 sg13g2_xnor2_1 _1648_ (.Y(_0779_),
    .A(_0776_),
    .B(_0778_));
 sg13g2_o21ai_1 _1649_ (.B1(net75),
    .Y(_0780_),
    .A1(net11),
    .A2(_0779_));
 sg13g2_nor3_1 _1650_ (.A(_0773_),
    .B(_0775_),
    .C(_0780_),
    .Y(_0063_));
 sg13g2_a21o_1 _1651_ (.A2(net31),
    .A1(net56),
    .B1(_0765_),
    .X(_0781_));
 sg13g2_and2_1 _1652_ (.A(net32),
    .B(_0715_),
    .X(_0782_));
 sg13g2_nor3_1 _1653_ (.A(net56),
    .B(net32),
    .C(_0715_),
    .Y(_0783_));
 sg13g2_o21ai_1 _1654_ (.B1(_0762_),
    .Y(_0784_),
    .A1(_0782_),
    .A2(_0783_));
 sg13g2_nor3_1 _1655_ (.A(_0774_),
    .B(_0702_),
    .C(net31),
    .Y(_0785_));
 sg13g2_nor2_1 _1656_ (.A(net56),
    .B(_0737_),
    .Y(_0786_));
 sg13g2_and2_1 _1657_ (.A(_0763_),
    .B(_0786_),
    .X(_0787_));
 sg13g2_a221oi_1 _1658_ (.B2(_0785_),
    .C1(_0787_),
    .B1(_0762_),
    .A1(net56),
    .Y(_0788_),
    .A2(_0715_));
 sg13g2_nand3_1 _1659_ (.B(_0784_),
    .C(_0788_),
    .A(_0781_),
    .Y(_0789_));
 sg13g2_buf_2 _1660_ (.A(\r[13] ),
    .X(_0790_));
 sg13g2_nor2_1 _1661_ (.A(_0776_),
    .B(_0716_),
    .Y(_0791_));
 sg13g2_xnor2_1 _1662_ (.Y(_0792_),
    .A(_0790_),
    .B(_0791_));
 sg13g2_xnor2_1 _1663_ (.Y(_0793_),
    .A(_0789_),
    .B(_0792_));
 sg13g2_buf_1 _1664_ (.A(_0006_),
    .X(_0794_));
 sg13g2_inv_2 _1665_ (.Y(_0795_),
    .A(_0794_));
 sg13g2_nand2_1 _1666_ (.Y(_0796_),
    .A(_0479_),
    .B(net58));
 sg13g2_a22oi_1 _1667_ (.Y(_0797_),
    .B1(_0750_),
    .B2(_0796_),
    .A2(_0685_),
    .A1(_0671_));
 sg13g2_nor2b_1 _1668_ (.A(_0466_),
    .B_N(\r[10] ),
    .Y(_0798_));
 sg13g2_o21ai_1 _1669_ (.B1(_0798_),
    .Y(_0799_),
    .A1(_0585_),
    .A2(_0739_));
 sg13g2_nand2b_1 _1670_ (.Y(_0800_),
    .B(_0739_),
    .A_N(_0585_));
 sg13g2_nand3b_1 _1671_ (.B(_0800_),
    .C(_0466_),
    .Y(_0801_),
    .A_N(net59));
 sg13g2_a221oi_1 _1672_ (.B2(_0801_),
    .C1(_0701_),
    .B1(_0799_),
    .A1(net58),
    .Y(_0802_),
    .A2(_0729_));
 sg13g2_nor2b_1 _1673_ (.A(_0797_),
    .B_N(_0802_),
    .Y(_0803_));
 sg13g2_nand3_1 _1674_ (.B(net59),
    .C(_0800_),
    .A(_0466_),
    .Y(_0804_));
 sg13g2_nor2_1 _1675_ (.A(_0466_),
    .B(\r[10] ),
    .Y(_0805_));
 sg13g2_o21ai_1 _1676_ (.B1(_0805_),
    .Y(_0806_),
    .A1(_0585_),
    .A2(_0739_));
 sg13g2_a21oi_1 _1677_ (.A1(_0804_),
    .A2(_0806_),
    .Y(_0807_),
    .B1(_0701_));
 sg13g2_inv_1 _1678_ (.Y(_0808_),
    .A(_0807_));
 sg13g2_nor2_1 _1679_ (.A(_0701_),
    .B(_0737_),
    .Y(_0809_));
 sg13g2_nor2b_1 _1680_ (.A(_0809_),
    .B_N(_0776_),
    .Y(_0810_));
 sg13g2_o21ai_1 _1681_ (.B1(_0810_),
    .Y(_0811_),
    .A1(_0692_),
    .A2(_0808_));
 sg13g2_o21ai_1 _1682_ (.B1(_0774_),
    .Y(_0812_),
    .A1(_0803_),
    .A2(_0811_));
 sg13g2_nor2_1 _1683_ (.A(_0738_),
    .B(_0776_),
    .Y(_0813_));
 sg13g2_nand3_1 _1684_ (.B(net21),
    .C(_0813_),
    .A(_0736_),
    .Y(_0814_));
 sg13g2_o21ai_1 _1685_ (.B1(_0814_),
    .Y(_0815_),
    .A1(net21),
    .A2(_0812_));
 sg13g2_xnor2_1 _1686_ (.Y(_0816_),
    .A(_0795_),
    .B(_0815_));
 sg13g2_o21ai_1 _1687_ (.B1(net75),
    .Y(_0817_),
    .A1(_0790_),
    .A2(net16));
 sg13g2_a221oi_1 _1688_ (.B2(_0650_),
    .C1(_0817_),
    .B1(_0816_),
    .A1(net12),
    .Y(_0064_),
    .A2(_0793_));
 sg13g2_buf_1 _1689_ (.A(\r[14] ),
    .X(_0818_));
 sg13g2_inv_1 _1690_ (.Y(_0819_),
    .A(_0818_));
 sg13g2_xnor2_1 _1691_ (.Y(_0820_),
    .A(net32),
    .B(_0763_));
 sg13g2_nand2_1 _1692_ (.Y(_0821_),
    .A(_0765_),
    .B(_0820_));
 sg13g2_nor2_1 _1693_ (.A(_0790_),
    .B(_0776_),
    .Y(_0822_));
 sg13g2_nor3_1 _1694_ (.A(_0715_),
    .B(_0786_),
    .C(_0822_),
    .Y(_0823_));
 sg13g2_nor3_1 _1695_ (.A(_0790_),
    .B(net56),
    .C(_0763_),
    .Y(_0824_));
 sg13g2_nor2_1 _1696_ (.A(_0823_),
    .B(_0824_),
    .Y(_0825_));
 sg13g2_a21oi_1 _1697_ (.A1(_0762_),
    .A2(_0821_),
    .Y(_0826_),
    .B1(_0825_));
 sg13g2_inv_1 _1698_ (.Y(_0827_),
    .A(_0790_));
 sg13g2_a21oi_1 _1699_ (.A1(_0760_),
    .A2(_0737_),
    .Y(_0828_),
    .B1(_0776_));
 sg13g2_nand3_1 _1700_ (.B(_0738_),
    .C(_0776_),
    .A(_0760_),
    .Y(_0829_));
 sg13g2_o21ai_1 _1701_ (.B1(_0829_),
    .Y(_0830_),
    .A1(_0827_),
    .A2(_0828_));
 sg13g2_o21ai_1 _1702_ (.B1(_0763_),
    .Y(_0831_),
    .A1(_0795_),
    .A2(_0830_));
 sg13g2_nor2b_1 _1703_ (.A(_0826_),
    .B_N(_0831_),
    .Y(_0832_));
 sg13g2_nor2_1 _1704_ (.A(_0794_),
    .B(_0716_),
    .Y(_0833_));
 sg13g2_o21ai_1 _1705_ (.B1(_0833_),
    .Y(_0834_),
    .A1(_0826_),
    .A2(_0830_));
 sg13g2_nor2b_1 _1706_ (.A(_0832_),
    .B_N(_0834_),
    .Y(_0835_));
 sg13g2_o21ai_1 _1707_ (.B1(net16),
    .Y(_0836_),
    .A1(_0704_),
    .A2(_0835_));
 sg13g2_nor2_1 _1708_ (.A(_0819_),
    .B(_0704_),
    .Y(_0837_));
 sg13g2_buf_1 _1709_ (.A(_0009_),
    .X(_0838_));
 sg13g2_and2_1 _1710_ (.A(_0795_),
    .B(net21),
    .X(_0839_));
 sg13g2_and3_1 _1711_ (.X(_0840_),
    .A(_0736_),
    .B(_0813_),
    .C(_0839_));
 sg13g2_nor4_2 _1712_ (.A(_0795_),
    .B(net21),
    .C(_0803_),
    .Y(_0841_),
    .D(_0811_));
 sg13g2_o21ai_1 _1713_ (.B1(_0827_),
    .Y(_0842_),
    .A1(_0774_),
    .A2(_0795_));
 sg13g2_nor3_1 _1714_ (.A(_0741_),
    .B(_0841_),
    .C(_0842_),
    .Y(_0843_));
 sg13g2_nor2_1 _1715_ (.A(_0840_),
    .B(_0843_),
    .Y(_0844_));
 sg13g2_xor2_1 _1716_ (.B(_0844_),
    .A(_0838_),
    .X(_0845_));
 sg13g2_o21ai_1 _1717_ (.B1(net75),
    .Y(_0846_),
    .A1(_0725_),
    .A2(_0845_));
 sg13g2_a221oi_1 _1718_ (.B2(_0835_),
    .C1(_0846_),
    .B1(_0837_),
    .A1(_0819_),
    .Y(_0065_),
    .A2(_0836_));
 sg13g2_buf_1 _1719_ (.A(\r[15] ),
    .X(_0847_));
 sg13g2_nor2_1 _1720_ (.A(_0838_),
    .B(net18),
    .Y(_0848_));
 sg13g2_xnor2_1 _1721_ (.Y(_0849_),
    .A(_0847_),
    .B(_0848_));
 sg13g2_nor2_1 _1722_ (.A(_0790_),
    .B(net55),
    .Y(_0850_));
 sg13g2_or2_1 _1723_ (.X(_0851_),
    .B(_0794_),
    .A(net55));
 sg13g2_buf_1 _1724_ (.A(_0851_),
    .X(_0852_));
 sg13g2_nand2b_1 _1725_ (.Y(_0853_),
    .B(_0852_),
    .A_N(_0822_));
 sg13g2_nor2_1 _1726_ (.A(_0715_),
    .B(_0853_),
    .Y(_0854_));
 sg13g2_a21oi_1 _1727_ (.A1(net18),
    .A2(_0850_),
    .Y(_0855_),
    .B1(_0854_));
 sg13g2_and2_1 _1728_ (.A(_0790_),
    .B(_0852_),
    .X(_0856_));
 sg13g2_a22oi_1 _1729_ (.Y(_0857_),
    .B1(_0856_),
    .B2(_0776_),
    .A2(_0794_),
    .A1(net55));
 sg13g2_or2_1 _1730_ (.X(_0858_),
    .B(_0857_),
    .A(net18));
 sg13g2_o21ai_1 _1731_ (.B1(_0858_),
    .Y(_0859_),
    .A1(_0789_),
    .A2(_0855_));
 sg13g2_xnor2_1 _1732_ (.Y(_0860_),
    .A(_0849_),
    .B(_0859_));
 sg13g2_nor2_1 _1733_ (.A(net55),
    .B(net21),
    .Y(_0861_));
 sg13g2_a21o_1 _1734_ (.A2(_0839_),
    .A1(_0813_),
    .B1(_0861_),
    .X(_0862_));
 sg13g2_nor3_1 _1735_ (.A(_0727_),
    .B(_0728_),
    .C(_0861_),
    .Y(_0863_));
 sg13g2_nand3b_1 _1736_ (.B(_0863_),
    .C(_0730_),
    .Y(_0864_),
    .A_N(_0734_));
 sg13g2_nand4_1 _1737_ (.B(_0736_),
    .C(_0813_),
    .A(net54),
    .Y(_0865_),
    .D(_0839_));
 sg13g2_o21ai_1 _1738_ (.B1(net54),
    .Y(_0866_),
    .A1(_0841_),
    .A2(_0842_));
 sg13g2_nand4_1 _1739_ (.B(_0864_),
    .C(_0865_),
    .A(_0862_),
    .Y(_0867_),
    .D(_0866_));
 sg13g2_xor2_1 _1740_ (.B(_0867_),
    .A(_0007_),
    .X(_0868_));
 sg13g2_a221oi_1 _1741_ (.B2(_0650_),
    .C1(_0575_),
    .B1(_0868_),
    .A1(net12),
    .Y(_0869_),
    .A2(_0860_));
 sg13g2_o21ai_1 _1742_ (.B1(_0506_),
    .Y(_0870_),
    .A1(_0847_),
    .A2(net16));
 sg13g2_nor2_1 _1743_ (.A(_0869_),
    .B(_0870_),
    .Y(_0066_));
 sg13g2_nor2_1 _1744_ (.A(net54),
    .B(_0007_),
    .Y(_0871_));
 sg13g2_nor2_1 _1745_ (.A(_0847_),
    .B(_0741_),
    .Y(_0872_));
 sg13g2_o21ai_1 _1746_ (.B1(_0007_),
    .Y(_0873_),
    .A1(net54),
    .A2(net55));
 sg13g2_nor2_1 _1747_ (.A(_0774_),
    .B(_0795_),
    .Y(_0874_));
 sg13g2_nand2_1 _1748_ (.Y(_0875_),
    .A(_0850_),
    .B(_0872_));
 sg13g2_nor3_1 _1749_ (.A(_0841_),
    .B(_0874_),
    .C(_0875_),
    .Y(_0876_));
 sg13g2_a221oi_1 _1750_ (.B2(_0873_),
    .C1(_0876_),
    .B1(_0872_),
    .A1(_0840_),
    .Y(_0877_),
    .A2(_0871_));
 sg13g2_xnor2_1 _1751_ (.Y(_0878_),
    .A(\r[16] ),
    .B(_0877_));
 sg13g2_a22oi_1 _1752_ (.Y(_0879_),
    .B1(_0650_),
    .B2(_0878_),
    .A2(_0575_),
    .A1(\r[16] ));
 sg13g2_inv_1 _1753_ (.Y(_0880_),
    .A(_0847_));
 sg13g2_nand3_1 _1754_ (.B(_0818_),
    .C(_0794_),
    .A(_0009_),
    .Y(_0881_));
 sg13g2_a21oi_1 _1755_ (.A1(net55),
    .A2(_0794_),
    .Y(_0882_),
    .B1(net54));
 sg13g2_a21oi_1 _1756_ (.A1(_0880_),
    .A2(_0881_),
    .Y(_0883_),
    .B1(_0882_));
 sg13g2_nor2_1 _1757_ (.A(_0830_),
    .B(_0883_),
    .Y(_0884_));
 sg13g2_nor2_1 _1758_ (.A(net18),
    .B(_0884_),
    .Y(_0885_));
 sg13g2_o21ai_1 _1759_ (.B1(_0763_),
    .Y(_0886_),
    .A1(net54),
    .A2(_0852_));
 sg13g2_a221oi_1 _1760_ (.B2(net54),
    .C1(_0847_),
    .B1(_0852_),
    .A1(_0587_),
    .Y(_0887_),
    .A2(_0713_));
 sg13g2_a221oi_1 _1761_ (.B2(_0847_),
    .C1(_0887_),
    .B1(_0886_),
    .A1(net55),
    .Y(_0888_),
    .A2(net18));
 sg13g2_o21ai_1 _1762_ (.B1(_0888_),
    .Y(_0889_),
    .A1(_0826_),
    .A2(_0885_));
 sg13g2_nor2_1 _1763_ (.A(_0007_),
    .B(net18),
    .Y(_0890_));
 sg13g2_xnor2_1 _1764_ (.Y(_0891_),
    .A(_0011_),
    .B(_0890_));
 sg13g2_xnor2_1 _1765_ (.Y(_0892_),
    .A(_0889_),
    .B(_0891_));
 sg13g2_nand2_1 _1766_ (.Y(_0893_),
    .A(net12),
    .B(_0892_));
 sg13g2_a21oi_1 _1767_ (.A1(_0879_),
    .A2(_0893_),
    .Y(_0067_),
    .B1(net57));
 sg13g2_inv_1 _1768_ (.Y(_0894_),
    .A(_0595_));
 sg13g2_xor2_1 _1769_ (.B(_0010_),
    .A(net70),
    .X(_0895_));
 sg13g2_a21oi_1 _1770_ (.A1(_0583_),
    .A2(_0895_),
    .Y(_0896_),
    .B1(_0575_));
 sg13g2_xnor2_1 _1771_ (.Y(_0897_),
    .A(_0595_),
    .B(_0568_));
 sg13g2_xnor2_1 _1772_ (.Y(_0898_),
    .A(net37),
    .B(_0897_));
 sg13g2_nor2_1 _1773_ (.A(_0595_),
    .B(_0895_),
    .Y(_0899_));
 sg13g2_a22oi_1 _1774_ (.Y(_0900_),
    .B1(_0899_),
    .B2(net12),
    .A2(_0898_),
    .A1(_0650_));
 sg13g2_o21ai_1 _1775_ (.B1(_0900_),
    .Y(_0901_),
    .A1(_0894_),
    .A2(_0896_));
 sg13g2_and2_1 _1776_ (.A(_0567_),
    .B(_0901_),
    .X(_0068_));
 sg13g2_buf_1 _1777_ (.A(_0488_),
    .X(_0902_));
 sg13g2_nor2_1 _1778_ (.A(_0596_),
    .B(_0655_),
    .Y(_0903_));
 sg13g2_xnor2_1 _1779_ (.Y(_0904_),
    .A(net38),
    .B(_0903_));
 sg13g2_nor2_1 _1780_ (.A(_0596_),
    .B(_0597_),
    .Y(_0905_));
 sg13g2_xnor2_1 _1781_ (.Y(_0906_),
    .A(_0449_),
    .B(_0905_));
 sg13g2_nor2_1 _1782_ (.A(net19),
    .B(_0906_),
    .Y(_0907_));
 sg13g2_a21oi_1 _1783_ (.A1(net19),
    .A2(_0904_),
    .Y(_0908_),
    .B1(_0907_));
 sg13g2_o21ai_1 _1784_ (.B1(net16),
    .Y(_0909_),
    .A1(net22),
    .A2(_0908_));
 sg13g2_nor2_1 _1785_ (.A(net63),
    .B(net20),
    .Y(_0910_));
 sg13g2_a22oi_1 _1786_ (.Y(_0911_),
    .B1(_0910_),
    .B2(_0908_),
    .A2(_0909_),
    .A1(net63));
 sg13g2_nor2_1 _1787_ (.A(_0902_),
    .B(_0911_),
    .Y(_0069_));
 sg13g2_nor2_1 _1788_ (.A(_0653_),
    .B(_0656_),
    .Y(_0912_));
 sg13g2_xor2_1 _1789_ (.B(_0592_),
    .A(net35),
    .X(_0913_));
 sg13g2_xnor2_1 _1790_ (.Y(_0914_),
    .A(_0912_),
    .B(_0913_));
 sg13g2_and2_1 _1791_ (.A(net71),
    .B(net63),
    .X(_0915_));
 sg13g2_nor3_1 _1792_ (.A(_0441_),
    .B(_0915_),
    .C(_0598_),
    .Y(_0916_));
 sg13g2_o21ai_1 _1793_ (.B1(_0441_),
    .Y(_0917_),
    .A1(_0915_),
    .A2(_0598_));
 sg13g2_nor2b_1 _1794_ (.A(_0916_),
    .B_N(_0917_),
    .Y(_0918_));
 sg13g2_a21oi_1 _1795_ (.A1(_0583_),
    .A2(_0918_),
    .Y(_0919_),
    .B1(_0575_));
 sg13g2_nand2_1 _1796_ (.Y(_0920_),
    .A(_0592_),
    .B(_0919_));
 sg13g2_inv_1 _1797_ (.Y(_0921_),
    .A(_0592_));
 sg13g2_o21ai_1 _1798_ (.B1(_0921_),
    .Y(_0922_),
    .A1(_0704_),
    .A2(_0918_));
 sg13g2_a22oi_1 _1799_ (.Y(_0923_),
    .B1(_0920_),
    .B2(_0922_),
    .A2(_0914_),
    .A1(_0650_));
 sg13g2_nor2_1 _1800_ (.A(_0902_),
    .B(_0923_),
    .Y(_0070_));
 sg13g2_a21oi_1 _1801_ (.A1(_0912_),
    .A2(_0658_),
    .Y(_0924_),
    .B1(_0661_));
 sg13g2_xor2_1 _1802_ (.B(_0924_),
    .A(net36),
    .X(_0925_));
 sg13g2_nor3_1 _1803_ (.A(_0527_),
    .B(_0599_),
    .C(_0600_),
    .Y(_0926_));
 sg13g2_o21ai_1 _1804_ (.B1(_0527_),
    .Y(_0927_),
    .A1(_0599_),
    .A2(_0600_));
 sg13g2_nand2b_1 _1805_ (.Y(_0928_),
    .B(_0927_),
    .A_N(_0926_));
 sg13g2_nor2_1 _1806_ (.A(net19),
    .B(_0928_),
    .Y(_0929_));
 sg13g2_a21oi_1 _1807_ (.A1(net19),
    .A2(_0925_),
    .Y(_0930_),
    .B1(_0929_));
 sg13g2_nor2b_1 _1808_ (.A(net22),
    .B_N(_0930_),
    .Y(_0931_));
 sg13g2_o21ai_1 _1809_ (.B1(_0601_),
    .Y(_0932_),
    .A1(_0575_),
    .A2(_0931_));
 sg13g2_or3_1 _1810_ (.A(_0601_),
    .B(net20),
    .C(_0930_),
    .X(_0933_));
 sg13g2_a21oi_1 _1811_ (.A1(_0932_),
    .A2(_0933_),
    .Y(_0071_),
    .B1(net57));
 sg13g2_o21ai_1 _1812_ (.B1(_0603_),
    .Y(_0934_),
    .A1(net50),
    .A2(_0601_));
 sg13g2_xnor2_1 _1813_ (.Y(_0935_),
    .A(net28),
    .B(_0934_));
 sg13g2_xnor2_1 _1814_ (.Y(_0936_),
    .A(_0482_),
    .B(_0665_));
 sg13g2_nand2_1 _1815_ (.Y(_0937_),
    .A(_0582_),
    .B(_0936_));
 sg13g2_o21ai_1 _1816_ (.B1(_0937_),
    .Y(_0938_),
    .A1(_0582_),
    .A2(_0935_));
 sg13g2_o21ai_1 _1817_ (.B1(net16),
    .Y(_0939_),
    .A1(net22),
    .A2(_0938_));
 sg13g2_nor2_1 _1818_ (.A(net61),
    .B(net20),
    .Y(_0940_));
 sg13g2_a22oi_1 _1819_ (.Y(_0941_),
    .B1(_0940_),
    .B2(_0938_),
    .A2(_0939_),
    .A1(net61));
 sg13g2_nor2_1 _1820_ (.A(net53),
    .B(_0941_),
    .Y(_0072_));
 sg13g2_a21o_1 _1821_ (.A2(_0665_),
    .A1(net61),
    .B1(net42),
    .X(_0942_));
 sg13g2_o21ai_1 _1822_ (.B1(_0942_),
    .Y(_0943_),
    .A1(net61),
    .A2(_0665_));
 sg13g2_xnor2_1 _1823_ (.Y(_0944_),
    .A(net41),
    .B(_0943_));
 sg13g2_o21ai_1 _1824_ (.B1(net16),
    .Y(_0945_),
    .A1(net11),
    .A2(_0944_));
 sg13g2_nor2_1 _1825_ (.A(net62),
    .B(net11),
    .Y(_0946_));
 sg13g2_a22oi_1 _1826_ (.Y(_0947_),
    .B1(_0946_),
    .B2(_0944_),
    .A2(_0945_),
    .A1(net62));
 sg13g2_mux2_1 _1827_ (.A0(_0614_),
    .A1(_0620_),
    .S(_0934_),
    .X(_0948_));
 sg13g2_xnor2_1 _1828_ (.Y(_0949_),
    .A(_0457_),
    .B(net62));
 sg13g2_xnor2_1 _1829_ (.Y(_0950_),
    .A(_0948_),
    .B(_0949_));
 sg13g2_nand2_1 _1830_ (.Y(_0951_),
    .A(net12),
    .B(_0950_));
 sg13g2_a21oi_1 _1831_ (.A1(_0947_),
    .A2(_0951_),
    .Y(_0073_),
    .B1(_0700_));
 sg13g2_a21oi_1 _1832_ (.A1(_0674_),
    .A2(_0943_),
    .Y(_0952_),
    .B1(_0668_));
 sg13g2_xnor2_1 _1833_ (.Y(_0953_),
    .A(net40),
    .B(_0952_));
 sg13g2_o21ai_1 _1834_ (.B1(net16),
    .Y(_0954_),
    .A1(net11),
    .A2(_0953_));
 sg13g2_nand2_1 _1835_ (.Y(_0955_),
    .A(net60),
    .B(_0954_));
 sg13g2_inv_1 _1836_ (.Y(_0956_),
    .A(_0624_));
 sg13g2_a21oi_2 _1837_ (.B1(_0618_),
    .Y(_0957_),
    .A2(_0934_),
    .A1(_0956_));
 sg13g2_xor2_1 _1838_ (.B(net60),
    .A(_0454_),
    .X(_0958_));
 sg13g2_xnor2_1 _1839_ (.Y(_0959_),
    .A(_0464_),
    .B(_0958_));
 sg13g2_xnor2_1 _1840_ (.Y(_0960_),
    .A(_0957_),
    .B(_0959_));
 sg13g2_nor2_1 _1841_ (.A(net60),
    .B(net11),
    .Y(_0961_));
 sg13g2_a22oi_1 _1842_ (.Y(_0962_),
    .B1(_0953_),
    .B2(_0961_),
    .A2(_0960_),
    .A1(net12));
 sg13g2_a21oi_1 _1843_ (.A1(_0955_),
    .A2(_0962_),
    .Y(_0074_),
    .B1(_0700_));
 sg13g2_or2_1 _1844_ (.X(_0963_),
    .B(_0952_),
    .A(_0481_));
 sg13g2_nand3_1 _1845_ (.B(_0627_),
    .C(_0952_),
    .A(_0481_),
    .Y(_0964_));
 sg13g2_o21ai_1 _1846_ (.B1(_0964_),
    .Y(_0965_),
    .A1(net60),
    .A2(_0963_));
 sg13g2_xnor2_1 _1847_ (.Y(_0966_),
    .A(_0666_),
    .B(_0965_));
 sg13g2_nand2_1 _1848_ (.Y(_0967_),
    .A(_0537_),
    .B(_0957_));
 sg13g2_o21ai_1 _1849_ (.B1(net60),
    .Y(_0968_),
    .A1(_0537_),
    .A2(_0957_));
 sg13g2_nand2_1 _1850_ (.Y(_0969_),
    .A(_0967_),
    .B(_0968_));
 sg13g2_nor4_1 _1851_ (.A(_0454_),
    .B(net60),
    .C(_0537_),
    .D(_0957_),
    .Y(_0970_));
 sg13g2_a221oi_1 _1852_ (.B2(net27),
    .C1(_0970_),
    .B1(_0969_),
    .A1(_0607_),
    .Y(_0971_),
    .A2(_0957_));
 sg13g2_xor2_1 _1853_ (.B(_0971_),
    .A(_0606_),
    .X(_0972_));
 sg13g2_o21ai_1 _1854_ (.B1(_0506_),
    .Y(_0973_),
    .A1(_0634_),
    .A2(_0721_));
 sg13g2_a221oi_1 _1855_ (.B2(_0584_),
    .C1(_0973_),
    .B1(_0972_),
    .A1(_0650_),
    .Y(_0075_),
    .A2(_0966_));
 sg13g2_xnor2_1 _1856_ (.Y(_0974_),
    .A(_0687_),
    .B(_0729_));
 sg13g2_o21ai_1 _1857_ (.B1(_0721_),
    .Y(_0975_),
    .A1(net11),
    .A2(_0974_));
 sg13g2_nand2_1 _1858_ (.Y(_0976_),
    .A(net58),
    .B(_0975_));
 sg13g2_nor2_1 _1859_ (.A(_0706_),
    .B(_0640_),
    .Y(_0977_));
 sg13g2_xnor2_1 _1860_ (.Y(_0978_),
    .A(_0689_),
    .B(_0977_));
 sg13g2_xnor2_1 _1861_ (.Y(_0979_),
    .A(_0633_),
    .B(_0978_));
 sg13g2_nor2_1 _1862_ (.A(_0689_),
    .B(net11),
    .Y(_0980_));
 sg13g2_a22oi_1 _1863_ (.Y(_0981_),
    .B1(_0974_),
    .B2(_0980_),
    .A2(_0979_),
    .A1(_0584_));
 sg13g2_a21oi_1 _1864_ (.A1(_0976_),
    .A2(_0981_),
    .Y(_0076_),
    .B1(_0488_));
 sg13g2_buf_2 _1865_ (.A(\counter[5] ),
    .X(_0982_));
 sg13g2_buf_1 _1866_ (.A(\counter[4] ),
    .X(_0983_));
 sg13g2_a22oi_1 _1867_ (.Y(_0984_),
    .B1(_0491_),
    .B2(\hvsync_gen.vpos[2] ),
    .A2(_0489_),
    .A1(net73));
 sg13g2_nor2_1 _1868_ (.A(net73),
    .B(_0489_),
    .Y(_0985_));
 sg13g2_nand2_1 _1869_ (.Y(_0986_),
    .A(_0446_),
    .B(_0496_));
 sg13g2_o21ai_1 _1870_ (.B1(_0986_),
    .Y(_0987_),
    .A1(_0984_),
    .A2(_0985_));
 sg13g2_xnor2_1 _1871_ (.Y(_0988_),
    .A(_0452_),
    .B(_0472_));
 sg13g2_nor2_1 _1872_ (.A(_0446_),
    .B(_0496_),
    .Y(_0989_));
 sg13g2_xnor2_1 _1873_ (.Y(_0990_),
    .A(_0455_),
    .B(net67));
 sg13g2_nor3_2 _1874_ (.A(_0988_),
    .B(_0989_),
    .C(_0990_),
    .Y(_0991_));
 sg13g2_a21o_1 _1875_ (.A2(net67),
    .A1(_0455_),
    .B1(_0472_),
    .X(_0992_));
 sg13g2_buf_1 _1876_ (.A(_0992_),
    .X(_0993_));
 sg13g2_and3_1 _1877_ (.X(_0994_),
    .A(_0455_),
    .B(net67),
    .C(_0472_));
 sg13g2_or2_1 _1878_ (.X(_0995_),
    .B(_0994_),
    .A(_0452_));
 sg13g2_buf_1 _1879_ (.A(_0995_),
    .X(_0996_));
 sg13g2_a221oi_1 _1880_ (.B2(_0996_),
    .C1(net41),
    .B1(_0993_),
    .A1(_0987_),
    .Y(_0997_),
    .A2(_0991_));
 sg13g2_buf_1 _1881_ (.A(_0987_),
    .X(_0998_));
 sg13g2_a221oi_1 _1882_ (.B2(_0996_),
    .C1(_0460_),
    .B1(_0993_),
    .A1(net23),
    .Y(_0999_),
    .A2(_0991_));
 sg13g2_nor2_1 _1883_ (.A(_0460_),
    .B(_0474_),
    .Y(_1000_));
 sg13g2_nor2_1 _1884_ (.A(\hvsync_gen.hpos[7] ),
    .B(_0435_),
    .Y(_1001_));
 sg13g2_inv_1 _1885_ (.Y(_1002_),
    .A(_1001_));
 sg13g2_o21ai_1 _1886_ (.B1(_1002_),
    .Y(_1003_),
    .A1(_0458_),
    .A2(net68));
 sg13g2_or4_1 _1887_ (.A(_0997_),
    .B(_0999_),
    .C(_1000_),
    .D(_1003_),
    .X(_1004_));
 sg13g2_buf_2 _1888_ (.A(_1004_),
    .X(_1005_));
 sg13g2_nand2_1 _1889_ (.Y(_1006_),
    .A(_0458_),
    .B(\hvsync_gen.hpos[6] ));
 sg13g2_nand2_1 _1890_ (.Y(_1007_),
    .A(net69),
    .B(_0435_));
 sg13g2_o21ai_1 _1891_ (.B1(_1007_),
    .Y(_1008_),
    .A1(_1006_),
    .A2(_1001_));
 sg13g2_inv_1 _1892_ (.Y(_1009_),
    .A(_1008_));
 sg13g2_nand2_1 _1893_ (.Y(_1010_),
    .A(_1005_),
    .B(_1009_));
 sg13g2_nand2_1 _1894_ (.Y(_1011_),
    .A(_0503_),
    .B(_1010_));
 sg13g2_xor2_1 _1895_ (.B(_1011_),
    .A(_0014_),
    .X(_1012_));
 sg13g2_nand2b_1 _1896_ (.Y(_1013_),
    .B(_1010_),
    .A_N(_0503_));
 sg13g2_nand2_1 _1897_ (.Y(_1014_),
    .A(net39),
    .B(_1006_));
 sg13g2_a221oi_1 _1898_ (.B2(_0996_),
    .C1(_1014_),
    .B1(_0993_),
    .A1(net23),
    .Y(_1015_),
    .A2(_0991_));
 sg13g2_nand2_1 _1899_ (.Y(_1016_),
    .A(_0540_),
    .B(_1006_));
 sg13g2_a221oi_1 _1900_ (.B2(_0996_),
    .C1(_1016_),
    .B1(_0993_),
    .A1(net23),
    .Y(_1017_),
    .A2(_0991_));
 sg13g2_nand2_1 _1901_ (.Y(_1018_),
    .A(_1006_),
    .B(_1000_));
 sg13g2_o21ai_1 _1902_ (.B1(_1018_),
    .Y(_1019_),
    .A1(_0458_),
    .A2(net68));
 sg13g2_nor3_2 _1903_ (.A(_1015_),
    .B(_1017_),
    .C(_1019_),
    .Y(_1020_));
 sg13g2_xor2_1 _1904_ (.B(_0435_),
    .A(net69),
    .X(_1021_));
 sg13g2_and2_1 _1905_ (.A(_0477_),
    .B(_1021_),
    .X(_1022_));
 sg13g2_nor2_1 _1906_ (.A(_0014_),
    .B(_1007_),
    .Y(_1023_));
 sg13g2_a21oi_2 _1907_ (.B1(_1023_),
    .Y(_1024_),
    .A2(_1022_),
    .A1(_1020_));
 sg13g2_xnor2_1 _1908_ (.Y(_1025_),
    .A(_0487_),
    .B(_1024_));
 sg13g2_xnor2_1 _1909_ (.Y(_1026_),
    .A(_1020_),
    .B(_1021_));
 sg13g2_buf_1 _1910_ (.A(_1026_),
    .X(_1027_));
 sg13g2_xor2_1 _1911_ (.B(\hvsync_gen.hpos[6] ),
    .A(_0458_),
    .X(_1028_));
 sg13g2_nand2_1 _1912_ (.Y(_1029_),
    .A(net41),
    .B(_1028_));
 sg13g2_nand2_1 _1913_ (.Y(_1030_),
    .A(net44),
    .B(_1028_));
 sg13g2_a21oi_1 _1914_ (.A1(net47),
    .A2(_0993_),
    .Y(_1031_),
    .B1(_0994_));
 sg13g2_a21oi_1 _1915_ (.A1(_1029_),
    .A2(_1030_),
    .Y(_1032_),
    .B1(_1031_));
 sg13g2_a21o_1 _1916_ (.A2(_0491_),
    .A1(\hvsync_gen.vpos[2] ),
    .B1(_0489_),
    .X(_1033_));
 sg13g2_and3_1 _1917_ (.X(_1034_),
    .A(net72),
    .B(_0489_),
    .C(_0491_));
 sg13g2_a221oi_1 _1918_ (.B2(net73),
    .C1(_1034_),
    .B1(_1033_),
    .A1(_0446_),
    .Y(_1035_),
    .A2(_0496_));
 sg13g2_buf_2 _1919_ (.A(_1035_),
    .X(_1036_));
 sg13g2_xor2_1 _1920_ (.B(_0472_),
    .A(_0452_),
    .X(_1037_));
 sg13g2_or2_1 _1921_ (.X(_1038_),
    .B(_0496_),
    .A(_0446_));
 sg13g2_buf_2 _1922_ (.A(_1038_),
    .X(_1039_));
 sg13g2_xor2_1 _1923_ (.B(net67),
    .A(_0455_),
    .X(_1040_));
 sg13g2_nand3_1 _1924_ (.B(_1039_),
    .C(_1040_),
    .A(_1037_),
    .Y(_1041_));
 sg13g2_nor3_1 _1925_ (.A(_1036_),
    .B(_1041_),
    .C(_1029_),
    .Y(_1042_));
 sg13g2_nor3_1 _1926_ (.A(_1036_),
    .B(_1041_),
    .C(_1030_),
    .Y(_1043_));
 sg13g2_xnor2_1 _1927_ (.Y(_1044_),
    .A(_0458_),
    .B(\hvsync_gen.hpos[6] ));
 sg13g2_nand2_1 _1928_ (.Y(_1045_),
    .A(net39),
    .B(_1044_));
 sg13g2_a221oi_1 _1929_ (.B2(_0996_),
    .C1(_1045_),
    .B1(_0993_),
    .A1(_0998_),
    .Y(_1046_),
    .A2(_0991_));
 sg13g2_nor4_2 _1930_ (.A(_1032_),
    .B(_1042_),
    .C(_1043_),
    .Y(_1047_),
    .D(_1046_));
 sg13g2_nand2_1 _1931_ (.Y(_1048_),
    .A(_0540_),
    .B(_1044_));
 sg13g2_a221oi_1 _1932_ (.B2(_0996_),
    .C1(_1048_),
    .B1(_0993_),
    .A1(_0998_),
    .Y(_1049_),
    .A2(_0991_));
 sg13g2_nand3_1 _1933_ (.B(net41),
    .C(_1028_),
    .A(net44),
    .Y(_1050_));
 sg13g2_nand2_1 _1934_ (.Y(_1051_),
    .A(_1000_),
    .B(_1044_));
 sg13g2_nand2_1 _1935_ (.Y(_1052_),
    .A(_1050_),
    .B(_1051_));
 sg13g2_nor2_2 _1936_ (.A(_1049_),
    .B(_1052_),
    .Y(_1053_));
 sg13g2_o21ai_1 _1937_ (.B1(_1031_),
    .Y(_1054_),
    .A1(_1036_),
    .A2(_1041_));
 sg13g2_xnor2_1 _1938_ (.Y(_1055_),
    .A(_0460_),
    .B(_0474_));
 sg13g2_xnor2_1 _1939_ (.Y(_1056_),
    .A(_1054_),
    .B(_1055_));
 sg13g2_nand3_1 _1940_ (.B(net36),
    .C(_1037_),
    .A(net26),
    .Y(_1057_));
 sg13g2_a21oi_1 _1941_ (.A1(net23),
    .A2(_1039_),
    .Y(_1058_),
    .B1(_1057_));
 sg13g2_nand2b_1 _1942_ (.Y(_1059_),
    .B(net26),
    .A_N(net36));
 sg13g2_nor4_1 _1943_ (.A(_1036_),
    .B(_0988_),
    .C(_0989_),
    .D(_1059_),
    .Y(_1060_));
 sg13g2_or3_1 _1944_ (.A(net46),
    .B(net67),
    .C(_1037_),
    .X(_1061_));
 sg13g2_a21oi_1 _1945_ (.A1(net23),
    .A2(_1039_),
    .Y(_1062_),
    .B1(_1061_));
 sg13g2_nand2_1 _1946_ (.Y(_1063_),
    .A(net67),
    .B(_1039_));
 sg13g2_nor4_1 _1947_ (.A(net26),
    .B(_1036_),
    .C(_0988_),
    .D(_1063_),
    .Y(_1064_));
 sg13g2_nor4_2 _1948_ (.A(_1058_),
    .B(_1060_),
    .C(_1062_),
    .Y(_1065_),
    .D(_1064_));
 sg13g2_nand4_1 _1949_ (.B(_1053_),
    .C(_1056_),
    .A(_1047_),
    .Y(_1066_),
    .D(_1065_));
 sg13g2_and2_1 _1950_ (.A(net15),
    .B(_1066_),
    .X(_1067_));
 sg13g2_nand2_1 _1951_ (.Y(_1068_),
    .A(_1025_),
    .B(_1067_));
 sg13g2_mux2_1 _1952_ (.A0(_1012_),
    .A1(_1013_),
    .S(_1068_),
    .X(_1069_));
 sg13g2_nand2b_1 _1953_ (.Y(_1070_),
    .B(_1069_),
    .A_N(_0983_));
 sg13g2_buf_1 _1954_ (.A(_1024_),
    .X(_1071_));
 sg13g2_a21oi_2 _1955_ (.B1(_0503_),
    .Y(_1072_),
    .A2(_1009_),
    .A1(_1005_));
 sg13g2_nand2_1 _1956_ (.Y(_1073_),
    .A(net14),
    .B(_1072_));
 sg13g2_inv_1 _1957_ (.Y(_1074_),
    .A(_0021_));
 sg13g2_nand3_1 _1958_ (.B(_1005_),
    .C(_1009_),
    .A(_0477_),
    .Y(_1075_));
 sg13g2_nor4_2 _1959_ (.A(_0997_),
    .B(_0999_),
    .C(_1000_),
    .Y(_1076_),
    .D(_1003_));
 sg13g2_o21ai_1 _1960_ (.B1(_0478_),
    .Y(_1077_),
    .A1(_1076_),
    .A2(_1008_));
 sg13g2_and2_1 _1961_ (.A(_1075_),
    .B(_1077_),
    .X(_1078_));
 sg13g2_a21oi_1 _1962_ (.A1(_1067_),
    .A2(_1078_),
    .Y(_1079_),
    .B1(net43));
 sg13g2_o21ai_1 _1963_ (.B1(_1072_),
    .Y(_1080_),
    .A1(net14),
    .A2(_1079_));
 sg13g2_nor2_1 _1964_ (.A(_1074_),
    .B(_1080_),
    .Y(_1081_));
 sg13g2_o21ai_1 _1965_ (.B1(_1081_),
    .Y(_1082_),
    .A1(_0982_),
    .A2(_1073_));
 sg13g2_o21ai_1 _1966_ (.B1(_1082_),
    .Y(_1083_),
    .A1(_0982_),
    .A2(_1070_));
 sg13g2_buf_1 _1967_ (.A(\counter[2] ),
    .X(_1084_));
 sg13g2_buf_1 _1968_ (.A(\counter[0] ),
    .X(_1085_));
 sg13g2_nor2_1 _1969_ (.A(net29),
    .B(_1066_),
    .Y(_1086_));
 sg13g2_buf_2 _1970_ (.A(\counter[1] ),
    .X(_1087_));
 sg13g2_nor2_1 _1971_ (.A(_1087_),
    .B(net15),
    .Y(_1088_));
 sg13g2_a22oi_1 _1972_ (.Y(_1089_),
    .B1(_1056_),
    .B2(_1065_),
    .A2(_1053_),
    .A1(_1047_));
 sg13g2_a22oi_1 _1973_ (.Y(_1090_),
    .B1(_1089_),
    .B2(net29),
    .A2(net15),
    .A1(_1087_));
 sg13g2_o21ai_1 _1974_ (.B1(_1090_),
    .Y(_1091_),
    .A1(_1086_),
    .A2(_1088_));
 sg13g2_xnor2_1 _1975_ (.Y(_1092_),
    .A(_0486_),
    .B(_1024_));
 sg13g2_inv_2 _1976_ (.Y(_1093_),
    .A(_1087_));
 sg13g2_inv_1 _1977_ (.Y(_1094_),
    .A(_1085_));
 sg13g2_nor2_2 _1978_ (.A(net24),
    .B(_1094_),
    .Y(_1095_));
 sg13g2_nand3_1 _1979_ (.B(_1089_),
    .C(_1095_),
    .A(net15),
    .Y(_1096_));
 sg13g2_nand2_2 _1980_ (.Y(_1097_),
    .A(_1075_),
    .B(_1077_));
 sg13g2_a21oi_1 _1981_ (.A1(_1092_),
    .A2(_1096_),
    .Y(_1098_),
    .B1(_1097_));
 sg13g2_a21o_1 _1982_ (.A2(_1091_),
    .A1(_1025_),
    .B1(_1098_),
    .X(_1099_));
 sg13g2_buf_2 _1983_ (.A(\counter[3] ),
    .X(_1100_));
 sg13g2_a21oi_1 _1984_ (.A1(net30),
    .A2(_1099_),
    .Y(_1101_),
    .B1(_1100_));
 sg13g2_xor2_1 _1985_ (.B(_1021_),
    .A(_1020_),
    .X(_1102_));
 sg13g2_buf_8 _1986_ (.A(_1102_),
    .X(_1103_));
 sg13g2_nand2b_1 _1987_ (.Y(_1104_),
    .B(net15),
    .A_N(_1089_));
 sg13g2_a22oi_1 _1988_ (.Y(_1105_),
    .B1(_1104_),
    .B2(net29),
    .A2(_1066_),
    .A1(net13));
 sg13g2_and2_1 _1989_ (.A(_1085_),
    .B(_1089_),
    .X(_1106_));
 sg13g2_nor2_1 _1990_ (.A(_1087_),
    .B(net29),
    .Y(_1107_));
 sg13g2_nor3_1 _1991_ (.A(net13),
    .B(_1066_),
    .C(_1107_),
    .Y(_1108_));
 sg13g2_a21oi_1 _1992_ (.A1(net13),
    .A2(_1106_),
    .Y(_1109_),
    .B1(_1108_));
 sg13g2_o21ai_1 _1993_ (.B1(_1109_),
    .Y(_1110_),
    .A1(net24),
    .A2(_1105_));
 sg13g2_nand2b_1 _1994_ (.Y(_1111_),
    .B(_1097_),
    .A_N(_1067_));
 sg13g2_nor2_1 _1995_ (.A(_1110_),
    .B(_1111_),
    .Y(_1112_));
 sg13g2_o21ai_1 _1996_ (.B1(_1092_),
    .Y(_1113_),
    .A1(_1101_),
    .A2(_1112_));
 sg13g2_nand3_1 _1997_ (.B(_1067_),
    .C(_1078_),
    .A(_1025_),
    .Y(_1114_));
 sg13g2_a21oi_1 _1998_ (.A1(_1100_),
    .A2(_1110_),
    .Y(_1115_),
    .B1(_1114_));
 sg13g2_nand2_1 _1999_ (.Y(_1116_),
    .A(_1092_),
    .B(_1096_));
 sg13g2_a21o_1 _2000_ (.A2(_1091_),
    .A1(_1078_),
    .B1(_1116_),
    .X(_1117_));
 sg13g2_a21oi_1 _2001_ (.A1(_1114_),
    .A2(_1117_),
    .Y(_1118_),
    .B1(net30));
 sg13g2_a221oi_1 _2002_ (.B2(_1110_),
    .C1(_1100_),
    .B1(_1111_),
    .A1(net30),
    .Y(_1119_),
    .A2(_1099_));
 sg13g2_nor3_1 _2003_ (.A(_1115_),
    .B(_1118_),
    .C(_1119_),
    .Y(_1120_));
 sg13g2_buf_2 _2004_ (.A(_0018_),
    .X(_1121_));
 sg13g2_inv_1 _2005_ (.Y(_1122_),
    .A(_1121_));
 sg13g2_xnor2_1 _2006_ (.Y(_1123_),
    .A(_1122_),
    .B(_1069_));
 sg13g2_xor2_1 _2007_ (.B(_1080_),
    .A(_0982_),
    .X(_1124_));
 sg13g2_nand2_1 _2008_ (.Y(_1125_),
    .A(_1123_),
    .B(_1124_));
 sg13g2_a21oi_1 _2009_ (.A1(_1113_),
    .A2(_1120_),
    .Y(_1126_),
    .B1(_1125_));
 sg13g2_nand2_1 _2010_ (.Y(_1127_),
    .A(_1121_),
    .B(net14));
 sg13g2_or2_1 _2011_ (.X(_1128_),
    .B(net14),
    .A(_1121_));
 sg13g2_a21o_1 _2012_ (.A2(_1039_),
    .A1(net23),
    .B1(net36),
    .X(_1129_));
 sg13g2_o21ai_1 _2013_ (.B1(_0509_),
    .Y(_1130_),
    .A1(_1036_),
    .A2(_1063_));
 sg13g2_nand2_1 _2014_ (.Y(_1131_),
    .A(_1129_),
    .B(_1130_));
 sg13g2_nor2_1 _2015_ (.A(_0988_),
    .B(_1055_),
    .Y(_1132_));
 sg13g2_a21oi_1 _2016_ (.A1(net23),
    .A2(_1039_),
    .Y(_1133_),
    .B1(net36));
 sg13g2_and2_1 _2017_ (.A(net67),
    .B(_1039_),
    .X(_1134_));
 sg13g2_a21oi_1 _2018_ (.A1(net23),
    .A2(_1134_),
    .Y(_1135_),
    .B1(net26));
 sg13g2_nor3_1 _2019_ (.A(net47),
    .B(net42),
    .C(_1055_),
    .Y(_1136_));
 sg13g2_nand3_1 _2020_ (.B(_0472_),
    .C(_1055_),
    .A(net47),
    .Y(_1137_));
 sg13g2_nor2b_1 _2021_ (.A(_1136_),
    .B_N(_1137_),
    .Y(_1138_));
 sg13g2_nor3_1 _2022_ (.A(_1133_),
    .B(_1135_),
    .C(_1138_),
    .Y(_1139_));
 sg13g2_a221oi_1 _2023_ (.B2(_1132_),
    .C1(_1139_),
    .B1(_1131_),
    .A1(_1047_),
    .Y(_1140_),
    .A2(_1053_));
 sg13g2_a22oi_1 _2024_ (.Y(_1141_),
    .B1(_1140_),
    .B2(net15),
    .A2(_1077_),
    .A1(_1075_));
 sg13g2_buf_2 _2025_ (.A(_1141_),
    .X(_1142_));
 sg13g2_mux2_1 _2026_ (.A0(_1127_),
    .A1(_1128_),
    .S(_1142_),
    .X(_1143_));
 sg13g2_nand3b_1 _2027_ (.B(_1013_),
    .C(_1121_),
    .Y(_1144_),
    .A_N(net14));
 sg13g2_nand2_1 _2028_ (.Y(_1145_),
    .A(_1122_),
    .B(net14));
 sg13g2_mux2_1 _2029_ (.A0(_1144_),
    .A1(_1145_),
    .S(_1142_),
    .X(_1146_));
 sg13g2_nor2_1 _2030_ (.A(_1013_),
    .B(_1128_),
    .Y(_1147_));
 sg13g2_nor2_1 _2031_ (.A(_0487_),
    .B(_1147_),
    .Y(_1148_));
 sg13g2_a22oi_1 _2032_ (.Y(_1149_),
    .B1(_1146_),
    .B2(_1148_),
    .A2(_1143_),
    .A1(_0487_));
 sg13g2_buf_2 _2033_ (.A(_0019_),
    .X(_1150_));
 sg13g2_buf_1 _2034_ (.A(_0020_),
    .X(_1151_));
 sg13g2_nand2_2 _2035_ (.Y(_1152_),
    .A(_1047_),
    .B(_1053_));
 sg13g2_a21oi_1 _2036_ (.A1(_1131_),
    .A2(_1132_),
    .Y(_1153_),
    .B1(_1139_));
 sg13g2_o21ai_1 _2037_ (.B1(net29),
    .Y(_1154_),
    .A1(_1152_),
    .A2(_1153_));
 sg13g2_and3_1 _2038_ (.X(_1155_),
    .A(_1151_),
    .B(net24),
    .C(_1154_));
 sg13g2_a21oi_1 _2039_ (.A1(_1047_),
    .A2(_1053_),
    .Y(_1156_),
    .B1(_1094_));
 sg13g2_or2_1 _2040_ (.X(_1157_),
    .B(_1156_),
    .A(_1153_));
 sg13g2_nand3_1 _2041_ (.B(_1047_),
    .C(_1053_),
    .A(_1094_),
    .Y(_1158_));
 sg13g2_and2_1 _2042_ (.A(_1087_),
    .B(_1158_),
    .X(_1159_));
 sg13g2_nand2_1 _2043_ (.Y(_1160_),
    .A(_1151_),
    .B(net13));
 sg13g2_a21oi_1 _2044_ (.A1(_1157_),
    .A2(_1159_),
    .Y(_1161_),
    .B1(_1160_));
 sg13g2_xnor2_1 _2045_ (.Y(_1162_),
    .A(_0014_),
    .B(_1010_));
 sg13g2_and3_1 _2046_ (.X(_1163_),
    .A(_1027_),
    .B(_1140_),
    .C(_1162_));
 sg13g2_inv_1 _2047_ (.Y(_1164_),
    .A(_1151_));
 sg13g2_nor2_1 _2048_ (.A(net24),
    .B(net13),
    .Y(_1165_));
 sg13g2_a21o_1 _2049_ (.A2(_1158_),
    .A1(_1153_),
    .B1(_1156_),
    .X(_1166_));
 sg13g2_a21oi_1 _2050_ (.A1(net24),
    .A2(_1103_),
    .Y(_1167_),
    .B1(_1151_));
 sg13g2_a221oi_1 _2051_ (.B2(_1167_),
    .C1(_1162_),
    .B1(_1166_),
    .A1(_1164_),
    .Y(_1168_),
    .A2(_1165_));
 sg13g2_nor4_2 _2052_ (.A(_1155_),
    .B(_1161_),
    .C(_1163_),
    .Y(_1169_),
    .D(_1168_));
 sg13g2_o21ai_1 _2053_ (.B1(_1100_),
    .Y(_1170_),
    .A1(_1150_),
    .A2(_1169_));
 sg13g2_nand2_1 _2054_ (.Y(_1171_),
    .A(_0468_),
    .B(_1142_));
 sg13g2_nor3_1 _2055_ (.A(_0487_),
    .B(net14),
    .C(_1072_),
    .Y(_1172_));
 sg13g2_nand2_1 _2056_ (.Y(_1173_),
    .A(net43),
    .B(_1142_));
 sg13g2_and2_1 _2057_ (.A(_0487_),
    .B(_1071_),
    .X(_1174_));
 sg13g2_and2_1 _2058_ (.A(_1071_),
    .B(_1072_),
    .X(_1175_));
 sg13g2_a221oi_1 _2059_ (.B2(_1174_),
    .C1(_1175_),
    .B1(_1173_),
    .A1(_1171_),
    .Y(_1176_),
    .A2(_1172_));
 sg13g2_xnor2_1 _2060_ (.Y(_1177_),
    .A(_1025_),
    .B(_1142_));
 sg13g2_nand3_1 _2061_ (.B(_1150_),
    .C(_1177_),
    .A(_1122_),
    .Y(_1178_));
 sg13g2_o21ai_1 _2062_ (.B1(_0983_),
    .Y(_1179_),
    .A1(_1169_),
    .A2(_1178_));
 sg13g2_nand3_1 _2063_ (.B(_1150_),
    .C(_1177_),
    .A(_1121_),
    .Y(_1180_));
 sg13g2_nor3_1 _2064_ (.A(_1169_),
    .B(_1176_),
    .C(_1180_),
    .Y(_1181_));
 sg13g2_a221oi_1 _2065_ (.B2(_1179_),
    .C1(_1181_),
    .B1(_1176_),
    .A1(_1149_),
    .Y(_1182_),
    .A2(_1170_));
 sg13g2_a21o_1 _2066_ (.A2(_1073_),
    .A1(_0982_),
    .B1(_1182_),
    .X(_1183_));
 sg13g2_o21ai_1 _2067_ (.B1(_1183_),
    .Y(_1184_),
    .A1(_1083_),
    .A2(_1126_));
 sg13g2_nor2b_1 _2068_ (.A(_0790_),
    .B_N(net55),
    .Y(_1185_));
 sg13g2_nor2_1 _2069_ (.A(_0601_),
    .B(_0592_),
    .Y(_1186_));
 sg13g2_inv_1 _2070_ (.Y(_1187_),
    .A(_0010_));
 sg13g2_o21ai_1 _2071_ (.B1(net63),
    .Y(_1188_),
    .A1(_0595_),
    .A2(_1187_));
 sg13g2_nand2_1 _2072_ (.Y(_1189_),
    .A(_1186_),
    .B(_1188_));
 sg13g2_o21ai_1 _2073_ (.B1(_0616_),
    .Y(_1190_),
    .A1(_0622_),
    .A2(_1189_));
 sg13g2_nand2_1 _2074_ (.Y(_1191_),
    .A(_0676_),
    .B(_1190_));
 sg13g2_a21o_1 _2075_ (.A2(_1191_),
    .A1(_0634_),
    .B1(net58),
    .X(_1192_));
 sg13g2_nand4_1 _2076_ (.B(net32),
    .C(_0648_),
    .A(net56),
    .Y(_1193_),
    .D(_1192_));
 sg13g2_a21oi_1 _2077_ (.A1(_1185_),
    .A2(_1193_),
    .Y(_1194_),
    .B1(net54));
 sg13g2_nand4_1 _2078_ (.B(_0701_),
    .C(net59),
    .A(\r[12] ),
    .Y(_1195_),
    .D(_0634_));
 sg13g2_nand4_1 _2079_ (.B(_0616_),
    .C(_0593_),
    .A(_0676_),
    .Y(_1196_),
    .D(_0011_));
 sg13g2_nor2_1 _2080_ (.A(net58),
    .B(_0622_),
    .Y(_1197_));
 sg13g2_nand4_1 _2081_ (.B(_1185_),
    .C(_1186_),
    .A(_0596_),
    .Y(_1198_),
    .D(_1197_));
 sg13g2_nor3_1 _2082_ (.A(_1195_),
    .B(_1196_),
    .C(_1198_),
    .Y(_1199_));
 sg13g2_nor3_1 _2083_ (.A(_0880_),
    .B(\r[16] ),
    .C(_1199_),
    .Y(_1200_));
 sg13g2_a21oi_1 _2084_ (.A1(_0617_),
    .A2(_1189_),
    .Y(_1201_),
    .B1(net60));
 sg13g2_or2_1 _2085_ (.X(_1202_),
    .B(_1195_),
    .A(_0591_));
 sg13g2_o21ai_1 _2086_ (.B1(_0850_),
    .Y(_1203_),
    .A1(_1201_),
    .A2(_1202_));
 sg13g2_nand2_1 _2087_ (.Y(_0103_),
    .A(net40),
    .B(_0484_));
 sg13g2_nand2_1 _2088_ (.Y(_0104_),
    .A(_0475_),
    .B(net40));
 sg13g2_nand2_1 _2089_ (.Y(_0105_),
    .A(net69),
    .B(_0104_));
 sg13g2_o21ai_1 _2090_ (.B1(_0105_),
    .Y(_0106_),
    .A1(net69),
    .A2(_0103_));
 sg13g2_or2_1 _2091_ (.X(_0107_),
    .B(net51),
    .A(net45));
 sg13g2_buf_1 _2092_ (.A(_0107_),
    .X(_0108_));
 sg13g2_nand2_1 _2093_ (.Y(_0109_),
    .A(net44),
    .B(_0508_));
 sg13g2_nor4_1 _2094_ (.A(net34),
    .B(net33),
    .C(_0108_),
    .D(_0109_),
    .Y(_0110_));
 sg13g2_o21ai_1 _2095_ (.B1(_0527_),
    .Y(_0111_),
    .A1(_0441_),
    .A2(_0449_));
 sg13g2_nor2_1 _2096_ (.A(_0635_),
    .B(_0108_),
    .Y(_0112_));
 sg13g2_o21ai_1 _2097_ (.B1(_0112_),
    .Y(_0113_),
    .A1(net50),
    .A2(_0443_));
 sg13g2_nand3_1 _2098_ (.B(_0111_),
    .C(_0113_),
    .A(_0537_),
    .Y(_0114_));
 sg13g2_nor3_1 _2099_ (.A(net28),
    .B(_0437_),
    .C(net49),
    .Y(_0115_));
 sg13g2_nand2b_1 _2100_ (.Y(_0116_),
    .B(net26),
    .A_N(_0115_));
 sg13g2_nand4_1 _2101_ (.B(_0527_),
    .C(net49),
    .A(net26),
    .Y(_0117_),
    .D(_0507_));
 sg13g2_o21ai_1 _2102_ (.B1(_0117_),
    .Y(_0118_),
    .A1(_0112_),
    .A2(_0116_));
 sg13g2_nand4_1 _2103_ (.B(_0110_),
    .C(_0114_),
    .A(_0106_),
    .Y(_0119_),
    .D(_0118_));
 sg13g2_nand3_1 _2104_ (.B(_1203_),
    .C(_0119_),
    .A(_1200_),
    .Y(_0120_));
 sg13g2_a21oi_1 _2105_ (.A1(_0482_),
    .A2(_0498_),
    .Y(_0121_),
    .B1(net39));
 sg13g2_inv_1 _2106_ (.Y(_0122_),
    .A(net69));
 sg13g2_nor2_1 _2107_ (.A(net25),
    .B(_0122_),
    .Y(_0123_));
 sg13g2_o21ai_1 _2108_ (.B1(_0123_),
    .Y(_0124_),
    .A1(net40),
    .A2(_0121_));
 sg13g2_nor2_1 _2109_ (.A(net33),
    .B(_0436_),
    .Y(_0125_));
 sg13g2_nand3_1 _2110_ (.B(_0124_),
    .C(_0125_),
    .A(_0463_),
    .Y(_0126_));
 sg13g2_a21oi_1 _2111_ (.A1(net38),
    .A2(_0497_),
    .Y(_0127_),
    .B1(_0495_));
 sg13g2_nor2_1 _2112_ (.A(_0475_),
    .B(net40),
    .Y(_0128_));
 sg13g2_o21ai_1 _2113_ (.B1(_0128_),
    .Y(_0129_),
    .A1(_0482_),
    .A2(_0127_));
 sg13g2_a21oi_1 _2114_ (.A1(_0123_),
    .A2(_0129_),
    .Y(_0130_),
    .B1(net33));
 sg13g2_nand4_1 _2115_ (.B(_0438_),
    .C(_0440_),
    .A(_0448_),
    .Y(_0131_),
    .D(net71));
 sg13g2_nand4_1 _2116_ (.B(_0508_),
    .C(_0509_),
    .A(_0540_),
    .Y(_0132_),
    .D(_0131_));
 sg13g2_a21oi_1 _2117_ (.A1(_0459_),
    .A2(_0132_),
    .Y(_0133_),
    .B1(net51));
 sg13g2_nor3_1 _2118_ (.A(_0126_),
    .B(_0130_),
    .C(_0133_),
    .Y(_0134_));
 sg13g2_nor3_1 _2119_ (.A(_1194_),
    .B(_0120_),
    .C(_0134_),
    .Y(_0135_));
 sg13g2_nor2_1 _2120_ (.A(_0540_),
    .B(net27),
    .Y(_0136_));
 sg13g2_a21oi_1 _2121_ (.A1(_0136_),
    .A2(_0116_),
    .Y(_0137_),
    .B1(_0605_));
 sg13g2_nor2_1 _2122_ (.A(_0109_),
    .B(_0117_),
    .Y(_0138_));
 sg13g2_nor4_1 _2123_ (.A(net33),
    .B(_0108_),
    .C(_0137_),
    .D(_0138_),
    .Y(_0139_));
 sg13g2_inv_1 _2124_ (.Y(_0140_),
    .A(_0490_));
 sg13g2_nor3_1 _2125_ (.A(_0140_),
    .B(_0498_),
    .C(_0104_),
    .Y(_0141_));
 sg13g2_mux2_1 _2126_ (.A0(net34),
    .A1(net42),
    .S(_0141_),
    .X(_0142_));
 sg13g2_a21oi_1 _2127_ (.A1(net34),
    .A2(_0492_),
    .Y(_0143_),
    .B1(_0142_));
 sg13g2_nand2_1 _2128_ (.Y(_0144_),
    .A(_0122_),
    .B(_0143_));
 sg13g2_nor2_1 _2129_ (.A(net42),
    .B(_0499_),
    .Y(_0145_));
 sg13g2_o21ai_1 _2130_ (.B1(_0122_),
    .Y(_0146_),
    .A1(_0104_),
    .A2(_0145_));
 sg13g2_nand2_1 _2131_ (.Y(_0147_),
    .A(net34),
    .B(_0146_));
 sg13g2_nand3_1 _2132_ (.B(_0144_),
    .C(_0147_),
    .A(_0139_),
    .Y(_0148_));
 sg13g2_nor3_1 _2133_ (.A(_0457_),
    .B(_0448_),
    .C(net50),
    .Y(_0149_));
 sg13g2_o21ai_1 _2134_ (.B1(_0540_),
    .Y(_0150_),
    .A1(_0508_),
    .A2(_0149_));
 sg13g2_a21oi_1 _2135_ (.A1(_0482_),
    .A2(_0127_),
    .Y(_0151_),
    .B1(net39));
 sg13g2_nor2_1 _2136_ (.A(_0502_),
    .B(_0151_),
    .Y(_0152_));
 sg13g2_nor3_1 _2137_ (.A(net34),
    .B(net39),
    .C(_0471_),
    .Y(_0153_));
 sg13g2_a21oi_1 _2138_ (.A1(net34),
    .A2(_0152_),
    .Y(_0154_),
    .B1(_0153_));
 sg13g2_a21oi_1 _2139_ (.A1(net45),
    .A2(_0150_),
    .Y(_0155_),
    .B1(_0154_));
 sg13g2_nand2_1 _2140_ (.Y(_0156_),
    .A(_0125_),
    .B(_0155_));
 sg13g2_nor2_1 _2141_ (.A(_0508_),
    .B(_0116_),
    .Y(_0157_));
 sg13g2_nor3_1 _2142_ (.A(net44),
    .B(_0108_),
    .C(_0157_),
    .Y(_0158_));
 sg13g2_a21oi_1 _2143_ (.A1(_0148_),
    .A2(_0156_),
    .Y(_0159_),
    .B1(_0158_));
 sg13g2_nand2_1 _2144_ (.Y(_0160_),
    .A(_0509_),
    .B(_0131_));
 sg13g2_nand3_1 _2145_ (.B(net27),
    .C(_0160_),
    .A(_0461_),
    .Y(_0161_));
 sg13g2_nor2_1 _2146_ (.A(net26),
    .B(net28),
    .Y(_0162_));
 sg13g2_nand3_1 _2147_ (.B(_0440_),
    .C(net71),
    .A(net50),
    .Y(_0163_));
 sg13g2_a21oi_1 _2148_ (.A1(_0162_),
    .A2(_0163_),
    .Y(_0164_),
    .B1(_0545_));
 sg13g2_a21oi_1 _2149_ (.A1(_0122_),
    .A2(_0103_),
    .Y(_0165_),
    .B1(net25));
 sg13g2_nor2_1 _2150_ (.A(net33),
    .B(_0165_),
    .Y(_0166_));
 sg13g2_nor3_1 _2151_ (.A(net51),
    .B(_0164_),
    .C(_0166_),
    .Y(_0167_));
 sg13g2_nand4_1 _2152_ (.B(_0495_),
    .C(_0497_),
    .A(_0490_),
    .Y(_0168_),
    .D(_0473_));
 sg13g2_a21o_1 _2153_ (.A2(_0168_),
    .A1(_0483_),
    .B1(_0471_),
    .X(_0169_));
 sg13g2_a21oi_1 _2154_ (.A1(_0569_),
    .A2(_0169_),
    .Y(_0170_),
    .B1(_0153_));
 sg13g2_nor2_1 _2155_ (.A(net33),
    .B(_0170_),
    .Y(_0171_));
 sg13g2_a22oi_1 _2156_ (.Y(_0172_),
    .B1(_0171_),
    .B2(_0133_),
    .A2(_0167_),
    .A1(_0130_));
 sg13g2_a21oi_1 _2157_ (.A1(_0713_),
    .A2(_0161_),
    .Y(_0173_),
    .B1(_0172_));
 sg13g2_nor3_1 _2158_ (.A(_0135_),
    .B(_0159_),
    .C(_0173_),
    .Y(_0174_));
 sg13g2_buf_1 _2159_ (.A(_0174_),
    .X(_0175_));
 sg13g2_xnor2_1 _2160_ (.Y(_0176_),
    .A(_0021_),
    .B(_1072_));
 sg13g2_xor2_1 _2161_ (.B(_0176_),
    .A(_0983_),
    .X(_0177_));
 sg13g2_and2_1 _2162_ (.A(_1092_),
    .B(_0177_),
    .X(_0178_));
 sg13g2_nor2_1 _2163_ (.A(_1092_),
    .B(_0176_),
    .Y(_0179_));
 sg13g2_and2_1 _2164_ (.A(_1047_),
    .B(_1053_),
    .X(_0180_));
 sg13g2_nor4_1 _2165_ (.A(_1151_),
    .B(_1094_),
    .C(_0180_),
    .D(_1056_),
    .Y(_0181_));
 sg13g2_nor3_1 _2166_ (.A(_1151_),
    .B(net24),
    .C(_0180_),
    .Y(_0182_));
 sg13g2_xor2_1 _2167_ (.B(_1055_),
    .A(_1054_),
    .X(_0183_));
 sg13g2_nand4_1 _2168_ (.B(_1087_),
    .C(net29),
    .A(_1164_),
    .Y(_0184_),
    .D(_0183_));
 sg13g2_o21ai_1 _2169_ (.B1(_0184_),
    .Y(_0185_),
    .A1(_1151_),
    .A2(net30));
 sg13g2_nor4_2 _2170_ (.A(net15),
    .B(_0181_),
    .C(_0182_),
    .Y(_0186_),
    .D(_0185_));
 sg13g2_nor4_2 _2171_ (.A(_0478_),
    .B(_1150_),
    .C(_1076_),
    .Y(_0187_),
    .D(_1008_));
 sg13g2_inv_1 _2172_ (.Y(_0188_),
    .A(_1150_));
 sg13g2_nor4_2 _2173_ (.A(_0477_),
    .B(_0188_),
    .C(_1076_),
    .Y(_0189_),
    .D(_1008_));
 sg13g2_nand2_1 _2174_ (.Y(_0190_),
    .A(net25),
    .B(_0188_));
 sg13g2_a21oi_1 _2175_ (.A1(_1005_),
    .A2(_1009_),
    .Y(_0191_),
    .B1(_0190_));
 sg13g2_nand2_1 _2176_ (.Y(_0192_),
    .A(_0477_),
    .B(_1150_));
 sg13g2_a21oi_1 _2177_ (.A1(_1005_),
    .A2(_1009_),
    .Y(_0193_),
    .B1(_0192_));
 sg13g2_or4_1 _2178_ (.A(_0187_),
    .B(_0189_),
    .C(_0191_),
    .D(_0193_),
    .X(_0194_));
 sg13g2_nand2_1 _2179_ (.Y(_0195_),
    .A(net29),
    .B(_1055_));
 sg13g2_nand2b_1 _2180_ (.Y(_0196_),
    .B(\counter[0] ),
    .A_N(_1055_));
 sg13g2_mux2_1 _2181_ (.A0(_0195_),
    .A1(_0196_),
    .S(_1054_),
    .X(_0197_));
 sg13g2_nor2_1 _2182_ (.A(net24),
    .B(_0197_),
    .Y(_0198_));
 sg13g2_a22oi_1 _2183_ (.Y(_0199_),
    .B1(_0197_),
    .B2(_1093_),
    .A2(_1053_),
    .A1(_1047_));
 sg13g2_or4_1 _2184_ (.A(_1084_),
    .B(_1103_),
    .C(_0198_),
    .D(_0199_),
    .X(_0200_));
 sg13g2_nor4_2 _2185_ (.A(_0187_),
    .B(_0189_),
    .C(_0191_),
    .Y(_0201_),
    .D(_0193_));
 sg13g2_a21o_1 _2186_ (.A2(_1077_),
    .A1(_1075_),
    .B1(_1100_),
    .X(_0202_));
 sg13g2_o21ai_1 _2187_ (.B1(_0202_),
    .Y(_0203_),
    .A1(_0200_),
    .A2(_0201_));
 sg13g2_a21oi_2 _2188_ (.B1(_0203_),
    .Y(_0204_),
    .A2(_0194_),
    .A1(_0186_));
 sg13g2_xnor2_1 _2189_ (.Y(_0205_),
    .A(_1121_),
    .B(_0204_));
 sg13g2_mux2_1 _2190_ (.A0(_0178_),
    .A1(_0179_),
    .S(_0205_),
    .X(_0206_));
 sg13g2_nor2b_1 _2191_ (.A(_0186_),
    .B_N(_0200_),
    .Y(_0207_));
 sg13g2_xnor2_1 _2192_ (.Y(_0208_),
    .A(_0207_),
    .B(_0194_));
 sg13g2_xnor2_1 _2193_ (.Y(_0209_),
    .A(net24),
    .B(_0197_));
 sg13g2_xnor2_1 _2194_ (.Y(_0210_),
    .A(_0180_),
    .B(_0209_));
 sg13g2_o21ai_1 _2195_ (.B1(_0988_),
    .Y(_0211_),
    .A1(_1133_),
    .A2(_1135_));
 sg13g2_buf_1 _2196_ (.A(_0211_),
    .X(_0212_));
 sg13g2_nand3_1 _2197_ (.B(_1129_),
    .C(_1130_),
    .A(_1037_),
    .Y(_0213_));
 sg13g2_buf_1 _2198_ (.A(_0213_),
    .X(_0214_));
 sg13g2_nand2_2 _2199_ (.Y(_0215_),
    .A(_0212_),
    .B(_0214_));
 sg13g2_inv_1 _2200_ (.Y(_0216_),
    .A(\grad1.acc[4] ));
 sg13g2_nor2_1 _2201_ (.A(_0216_),
    .B(_0017_),
    .Y(_0217_));
 sg13g2_inv_1 _2202_ (.Y(_0218_),
    .A(_0017_));
 sg13g2_nand3_1 _2203_ (.B(_1129_),
    .C(_1130_),
    .A(_0988_),
    .Y(_0219_));
 sg13g2_o21ai_1 _2204_ (.B1(_1037_),
    .Y(_0220_),
    .A1(_1133_),
    .A2(_1135_));
 sg13g2_nand2_1 _2205_ (.Y(_0221_),
    .A(_0219_),
    .B(_0220_));
 sg13g2_nor2_1 _2206_ (.A(_0218_),
    .B(_0221_),
    .Y(_0222_));
 sg13g2_inv_2 _2207_ (.Y(_0223_),
    .A(\grad1.acc[2] ));
 sg13g2_o21ai_1 _2208_ (.B1(_1033_),
    .Y(_0224_),
    .A1(net73),
    .A2(_1034_));
 sg13g2_xor2_1 _2209_ (.B(net35),
    .A(net48),
    .X(_0225_));
 sg13g2_xnor2_1 _2210_ (.Y(_0226_),
    .A(_0224_),
    .B(_0225_));
 sg13g2_nor2_1 _2211_ (.A(_0223_),
    .B(_0226_),
    .Y(_0227_));
 sg13g2_xor2_1 _2212_ (.B(_0225_),
    .A(_0224_),
    .X(_0228_));
 sg13g2_nor2_1 _2213_ (.A(\grad1.acc[2] ),
    .B(_0228_),
    .Y(_0229_));
 sg13g2_buf_2 _2214_ (.A(\grad1.acc[1] ),
    .X(_0230_));
 sg13g2_xor2_1 _2215_ (.B(_0489_),
    .A(net73),
    .X(_0231_));
 sg13g2_xnor2_1 _2216_ (.Y(_0232_),
    .A(_0230_),
    .B(_0231_));
 sg13g2_buf_2 _2217_ (.A(\grad1.acc[0] ),
    .X(_0233_));
 sg13g2_nor2b_1 _2218_ (.A(_0233_),
    .B_N(net37),
    .Y(_0234_));
 sg13g2_nor2b_1 _2219_ (.A(net37),
    .B_N(_0233_),
    .Y(_0235_));
 sg13g2_nor3_1 _2220_ (.A(net72),
    .B(_0234_),
    .C(_0235_),
    .Y(_0236_));
 sg13g2_mux2_1 _2221_ (.A0(_0234_),
    .A1(_0235_),
    .S(_0232_),
    .X(_0237_));
 sg13g2_a22oi_1 _2222_ (.Y(_0238_),
    .B1(_0237_),
    .B2(net72),
    .A2(_0236_),
    .A1(_0232_));
 sg13g2_nor3_1 _2223_ (.A(_0227_),
    .B(_0229_),
    .C(_0238_),
    .Y(_0239_));
 sg13g2_buf_1 _2224_ (.A(\grad1.acc[3] ),
    .X(_0240_));
 sg13g2_nor2_1 _2225_ (.A(_1036_),
    .B(_0989_),
    .Y(_0241_));
 sg13g2_xnor2_1 _2226_ (.Y(_0242_),
    .A(_0990_),
    .B(_0241_));
 sg13g2_xnor2_1 _2227_ (.Y(_0243_),
    .A(net52),
    .B(_0242_));
 sg13g2_or2_1 _2228_ (.X(_0244_),
    .B(_0234_),
    .A(net72));
 sg13g2_nor2_1 _2229_ (.A(_0230_),
    .B(_0235_),
    .Y(_0245_));
 sg13g2_a21o_1 _2230_ (.A2(_0245_),
    .A1(_0244_),
    .B1(_0231_),
    .X(_0246_));
 sg13g2_nor2_1 _2231_ (.A(net72),
    .B(net37),
    .Y(_0247_));
 sg13g2_o21ai_1 _2232_ (.B1(_0230_),
    .Y(_0248_),
    .A1(_0233_),
    .A2(_0247_));
 sg13g2_nand3_1 _2233_ (.B(net37),
    .C(_0231_),
    .A(net72),
    .Y(_0249_));
 sg13g2_and2_1 _2234_ (.A(_0248_),
    .B(_0249_),
    .X(_0250_));
 sg13g2_a22oi_1 _2235_ (.Y(_0251_),
    .B1(_0246_),
    .B2(_0250_),
    .A2(_0226_),
    .A1(_0223_));
 sg13g2_xnor2_1 _2236_ (.Y(_0252_),
    .A(_1040_),
    .B(_0241_));
 sg13g2_buf_1 _2237_ (.A(_0252_),
    .X(_0253_));
 sg13g2_o21ai_1 _2238_ (.B1(net17),
    .Y(_0254_),
    .A1(_0227_),
    .A2(_0251_));
 sg13g2_inv_1 _2239_ (.Y(_0255_),
    .A(net52));
 sg13g2_nor3_1 _2240_ (.A(_0227_),
    .B(_0253_),
    .C(_0251_),
    .Y(_0256_));
 sg13g2_a221oi_1 _2241_ (.B2(_0255_),
    .C1(_0256_),
    .B1(_0254_),
    .A1(_0239_),
    .Y(_0257_),
    .A2(_0243_));
 sg13g2_a221oi_1 _2242_ (.B2(_0243_),
    .C1(_0216_),
    .B1(_0239_),
    .A1(_0212_),
    .Y(_0258_),
    .A2(_0214_));
 sg13g2_a221oi_1 _2243_ (.B2(_0257_),
    .C1(_0258_),
    .B1(_0222_),
    .A1(_0215_),
    .Y(_0259_),
    .A2(_0217_));
 sg13g2_nor2_1 _2244_ (.A(_0017_),
    .B(_0215_),
    .Y(_0260_));
 sg13g2_xnor2_1 _2245_ (.Y(_0261_),
    .A(_0024_),
    .B(_0183_));
 sg13g2_a21oi_1 _2246_ (.A1(_0257_),
    .A2(_0260_),
    .Y(_0262_),
    .B1(_0261_));
 sg13g2_a22oi_1 _2247_ (.Y(_0263_),
    .B1(_0259_),
    .B2(_0262_),
    .A2(_0210_),
    .A1(_0016_));
 sg13g2_buf_2 _2248_ (.A(\grad1.acc[5] ),
    .X(_0264_));
 sg13g2_a21oi_1 _2249_ (.A1(_0257_),
    .A2(_0260_),
    .Y(_0265_),
    .B1(_0264_));
 sg13g2_nor2_1 _2250_ (.A(_0264_),
    .B(_0261_),
    .Y(_0266_));
 sg13g2_a21oi_1 _2251_ (.A1(_0259_),
    .A2(_0265_),
    .Y(_0267_),
    .B1(_0266_));
 sg13g2_nor2_1 _2252_ (.A(_0016_),
    .B(_0210_),
    .Y(_0268_));
 sg13g2_a21oi_2 _2253_ (.B1(_0268_),
    .Y(_0269_),
    .A2(_0267_),
    .A1(_0263_));
 sg13g2_nand2_1 _2254_ (.Y(_0270_),
    .A(_1093_),
    .B(_0197_));
 sg13g2_o21ai_1 _2255_ (.B1(_0270_),
    .Y(_0271_),
    .A1(_1152_),
    .A2(_0198_));
 sg13g2_xnor2_1 _2256_ (.Y(_0272_),
    .A(_1084_),
    .B(net15));
 sg13g2_xnor2_1 _2257_ (.Y(_0273_),
    .A(_0271_),
    .B(_0272_));
 sg13g2_nand3_1 _2258_ (.B(_0269_),
    .C(_0273_),
    .A(_0208_),
    .Y(_0274_));
 sg13g2_or3_1 _2259_ (.A(_0208_),
    .B(_0269_),
    .C(_0273_),
    .X(_0275_));
 sg13g2_and3_1 _2260_ (.X(_0276_),
    .A(_0206_),
    .B(_0274_),
    .C(_0275_));
 sg13g2_a21oi_1 _2261_ (.A1(_0244_),
    .A2(_0245_),
    .Y(_0277_),
    .B1(_0231_));
 sg13g2_nand2_1 _2262_ (.Y(_0278_),
    .A(_0248_),
    .B(_0249_));
 sg13g2_o21ai_1 _2263_ (.B1(_0228_),
    .Y(_0279_),
    .A1(_0277_),
    .A2(_0278_));
 sg13g2_nand2_1 _2264_ (.Y(_0280_),
    .A(_0223_),
    .B(_0279_));
 sg13g2_nor3_2 _2265_ (.A(_0228_),
    .B(_0277_),
    .C(_0278_),
    .Y(_0281_));
 sg13g2_nor2_1 _2266_ (.A(_0255_),
    .B(_0281_),
    .Y(_0282_));
 sg13g2_a21oi_1 _2267_ (.A1(_0280_),
    .A2(_0282_),
    .Y(_0283_),
    .B1(_0215_));
 sg13g2_a21oi_2 _2268_ (.B1(_0281_),
    .Y(_0284_),
    .A2(_0279_),
    .A1(_0223_));
 sg13g2_o21ai_1 _2269_ (.B1(_0218_),
    .Y(_0285_),
    .A1(net52),
    .A2(_0284_));
 sg13g2_nor2_1 _2270_ (.A(_0221_),
    .B(net17),
    .Y(_0286_));
 sg13g2_a22oi_1 _2271_ (.Y(_0287_),
    .B1(_0285_),
    .B2(_0286_),
    .A2(_0283_),
    .A1(net17));
 sg13g2_nand3_1 _2272_ (.B(_0280_),
    .C(_0282_),
    .A(_0215_),
    .Y(_0288_));
 sg13g2_nor2_1 _2273_ (.A(net17),
    .B(_0281_),
    .Y(_0289_));
 sg13g2_a221oi_1 _2274_ (.B2(_0289_),
    .C1(_0218_),
    .B1(_0280_),
    .A1(net52),
    .Y(_0290_),
    .A2(_0242_));
 sg13g2_inv_1 _2275_ (.Y(_0291_),
    .A(_0264_));
 sg13g2_a21oi_1 _2276_ (.A1(_0288_),
    .A2(_0290_),
    .Y(_0292_),
    .B1(_0291_));
 sg13g2_a21oi_1 _2277_ (.A1(_0219_),
    .A2(_0220_),
    .Y(_0293_),
    .B1(net17));
 sg13g2_xnor2_1 _2278_ (.Y(_0294_),
    .A(_1056_),
    .B(_0293_));
 sg13g2_nor2_1 _2279_ (.A(_0255_),
    .B(_0017_),
    .Y(_0295_));
 sg13g2_a21oi_1 _2280_ (.A1(_0212_),
    .A2(_0214_),
    .Y(_0296_),
    .B1(_0017_));
 sg13g2_o21ai_1 _2281_ (.B1(_0284_),
    .Y(_0297_),
    .A1(_0295_),
    .A2(_0296_));
 sg13g2_and4_1 _2282_ (.A(net52),
    .B(_0219_),
    .C(_0220_),
    .D(net17),
    .X(_0298_));
 sg13g2_and4_1 _2283_ (.A(_0218_),
    .B(_0212_),
    .C(_0214_),
    .D(_0242_),
    .X(_0299_));
 sg13g2_a221oi_1 _2284_ (.B2(_0284_),
    .C1(_0299_),
    .B1(_0298_),
    .A1(_0215_),
    .Y(_0300_),
    .A2(_0295_));
 sg13g2_nor2_1 _2285_ (.A(_0255_),
    .B(net17),
    .Y(_0301_));
 sg13g2_and4_1 _2286_ (.A(_0218_),
    .B(_0219_),
    .C(_0220_),
    .D(net17),
    .X(_0302_));
 sg13g2_a221oi_1 _2287_ (.B2(_0293_),
    .C1(_0302_),
    .B1(_0284_),
    .A1(_0221_),
    .Y(_0303_),
    .A2(_0301_));
 sg13g2_nand4_1 _2288_ (.B(_0297_),
    .C(_0300_),
    .A(_0291_),
    .Y(_0304_),
    .D(_0303_));
 sg13g2_buf_2 _2289_ (.A(\grad1.acc[6] ),
    .X(_0305_));
 sg13g2_nand4_1 _2290_ (.B(_0212_),
    .C(_0214_),
    .A(_1056_),
    .Y(_0306_),
    .D(_0242_));
 sg13g2_xnor2_1 _2291_ (.Y(_0307_),
    .A(_1152_),
    .B(_0306_));
 sg13g2_and2_1 _2292_ (.A(_0305_),
    .B(_0307_),
    .X(_0308_));
 sg13g2_a221oi_1 _2293_ (.B2(_0304_),
    .C1(_0308_),
    .B1(_0294_),
    .A1(_0287_),
    .Y(_0309_),
    .A2(_0292_));
 sg13g2_inv_1 _2294_ (.Y(_0310_),
    .A(\grad1.acc[7] ));
 sg13g2_nor2_2 _2295_ (.A(_1152_),
    .B(_0306_),
    .Y(_0311_));
 sg13g2_nor2_2 _2296_ (.A(net13),
    .B(_0311_),
    .Y(_0312_));
 sg13g2_xnor2_1 _2297_ (.Y(_0313_),
    .A(_0015_),
    .B(_1097_));
 sg13g2_nor2_1 _2298_ (.A(_0305_),
    .B(_0016_),
    .Y(_0314_));
 sg13g2_mux2_1 _2299_ (.A0(_0016_),
    .A1(_0314_),
    .S(_0307_),
    .X(_0315_));
 sg13g2_nor4_1 _2300_ (.A(_0310_),
    .B(_0312_),
    .C(_0313_),
    .D(_0315_),
    .Y(_0316_));
 sg13g2_nor2b_1 _2301_ (.A(_0309_),
    .B_N(_0316_),
    .Y(_0317_));
 sg13g2_xnor2_1 _2302_ (.Y(_0318_),
    .A(net13),
    .B(_0311_));
 sg13g2_nor3_1 _2303_ (.A(_0310_),
    .B(_0313_),
    .C(_0318_),
    .Y(_0319_));
 sg13g2_nor4_1 _2304_ (.A(_0313_),
    .B(_0309_),
    .C(_0315_),
    .D(_0318_),
    .Y(_0320_));
 sg13g2_nor3_1 _2305_ (.A(_0317_),
    .B(_0319_),
    .C(_0320_),
    .Y(_0321_));
 sg13g2_xnor2_1 _2306_ (.Y(_0322_),
    .A(_1097_),
    .B(_0312_));
 sg13g2_nand2_1 _2307_ (.Y(_0323_),
    .A(\grad1.acc[7] ),
    .B(_0312_));
 sg13g2_nor3_1 _2308_ (.A(_0309_),
    .B(_0315_),
    .C(_0323_),
    .Y(_0324_));
 sg13g2_a22oi_1 _2309_ (.Y(_0325_),
    .B1(_0313_),
    .B2(_0324_),
    .A2(_0322_),
    .A1(\grad1.acc[8] ));
 sg13g2_xnor2_1 _2310_ (.Y(_0326_),
    .A(net43),
    .B(net14));
 sg13g2_o21ai_1 _2311_ (.B1(_1097_),
    .Y(_0327_),
    .A1(_1092_),
    .A2(_1162_));
 sg13g2_a21oi_1 _2312_ (.A1(_0312_),
    .A2(_0327_),
    .Y(_0328_),
    .B1(_1072_));
 sg13g2_nor2_1 _2313_ (.A(_1092_),
    .B(_1162_),
    .Y(_0329_));
 sg13g2_xnor2_1 _2314_ (.Y(_0330_),
    .A(_1072_),
    .B(_0329_));
 sg13g2_nor4_1 _2315_ (.A(net13),
    .B(_1097_),
    .C(_0311_),
    .D(_0326_),
    .Y(_0331_));
 sg13g2_a22oi_1 _2316_ (.Y(_0332_),
    .B1(_0330_),
    .B2(_0331_),
    .A2(_0328_),
    .A1(_0326_));
 sg13g2_a21oi_1 _2317_ (.A1(_0321_),
    .A2(_0325_),
    .Y(_0333_),
    .B1(_0332_));
 sg13g2_nor3_1 _2318_ (.A(net10),
    .B(_0276_),
    .C(_0333_),
    .Y(_0334_));
 sg13g2_inv_1 _2319_ (.Y(_0335_),
    .A(_0305_));
 sg13g2_nor2_1 _2320_ (.A(net49),
    .B(_0223_),
    .Y(_0336_));
 sg13g2_nor2b_1 _2321_ (.A(net70),
    .B_N(_0233_),
    .Y(_0337_));
 sg13g2_nand2_1 _2322_ (.Y(_0338_),
    .A(_0230_),
    .B(_0337_));
 sg13g2_o21ai_1 _2323_ (.B1(_0449_),
    .Y(_0339_),
    .A1(_0230_),
    .A2(_0337_));
 sg13g2_a22oi_1 _2324_ (.Y(_0340_),
    .B1(_0338_),
    .B2(_0339_),
    .A2(_0223_),
    .A1(net72));
 sg13g2_o21ai_1 _2325_ (.B1(net52),
    .Y(_0341_),
    .A1(_0336_),
    .A2(_0340_));
 sg13g2_nor3_1 _2326_ (.A(_0240_),
    .B(_0336_),
    .C(_0340_),
    .Y(_0342_));
 sg13g2_a21oi_1 _2327_ (.A1(net50),
    .A2(_0341_),
    .Y(_0343_),
    .B1(_0342_));
 sg13g2_o21ai_1 _2328_ (.B1(_0343_),
    .Y(_0344_),
    .A1(_0536_),
    .A2(\grad1.acc[4] ));
 sg13g2_o21ai_1 _2329_ (.B1(_0344_),
    .Y(_0345_),
    .A1(net28),
    .A2(_0216_));
 sg13g2_nand2_1 _2330_ (.Y(_0346_),
    .A(_0264_),
    .B(_0345_));
 sg13g2_o21ai_1 _2331_ (.B1(_0509_),
    .Y(_0347_),
    .A1(_0264_),
    .A2(_0345_));
 sg13g2_a22oi_1 _2332_ (.Y(_0348_),
    .B1(_0346_),
    .B2(_0347_),
    .A2(_0335_),
    .A1(net27));
 sg13g2_a21oi_2 _2333_ (.B1(_0348_),
    .Y(_0349_),
    .A2(_0305_),
    .A1(_0508_));
 sg13g2_and2_1 _2334_ (.A(_0462_),
    .B(_0349_),
    .X(_0350_));
 sg13g2_a221oi_1 _2335_ (.B2(net10),
    .C1(net20),
    .B1(_0350_),
    .A1(_1184_),
    .Y(_0077_),
    .A2(_0334_));
 sg13g2_or2_1 _2336_ (.X(_0351_),
    .B(_0273_),
    .A(_0269_));
 sg13g2_nand2_1 _2337_ (.Y(_0352_),
    .A(_0269_),
    .B(_0273_));
 sg13g2_nand4_1 _2338_ (.B(_0208_),
    .C(_0351_),
    .A(_0206_),
    .Y(_0353_),
    .D(_0352_));
 sg13g2_nor2b_1 _2339_ (.A(_0175_),
    .B_N(_0353_),
    .Y(_0354_));
 sg13g2_nor2_1 _2340_ (.A(_0605_),
    .B(_0013_),
    .Y(_0355_));
 sg13g2_nor2_1 _2341_ (.A(net45),
    .B(_0461_),
    .Y(_0356_));
 sg13g2_nor3_1 _2342_ (.A(_0635_),
    .B(_0462_),
    .C(_0356_),
    .Y(_0357_));
 sg13g2_mux2_1 _2343_ (.A0(_0355_),
    .A1(_0357_),
    .S(_0349_),
    .X(_0358_));
 sg13g2_or2_1 _2344_ (.X(_0359_),
    .B(_0358_),
    .A(_0350_));
 sg13g2_a221oi_1 _2345_ (.B2(net10),
    .C1(net20),
    .B1(_0359_),
    .A1(_1184_),
    .Y(_0078_),
    .A2(_0354_));
 sg13g2_nor2_1 _2346_ (.A(net10),
    .B(_0333_),
    .Y(_0360_));
 sg13g2_a21oi_1 _2347_ (.A1(_1184_),
    .A2(_0360_),
    .Y(_0079_),
    .B1(net20));
 sg13g2_a21o_1 _2348_ (.A2(_0325_),
    .A1(_0321_),
    .B1(_0332_),
    .X(_0361_));
 sg13g2_nor4_1 _2349_ (.A(_1122_),
    .B(_1092_),
    .C(_0176_),
    .D(_0204_),
    .Y(_0362_));
 sg13g2_nor4_1 _2350_ (.A(_1121_),
    .B(_1025_),
    .C(_0176_),
    .D(_0204_),
    .Y(_0363_));
 sg13g2_nor2_1 _2351_ (.A(_0362_),
    .B(_0363_),
    .Y(_0364_));
 sg13g2_nor3_1 _2352_ (.A(_1122_),
    .B(_1025_),
    .C(_0177_),
    .Y(_0365_));
 sg13g2_and3_1 _2353_ (.X(_0366_),
    .A(_1122_),
    .B(_1025_),
    .C(_0176_));
 sg13g2_o21ai_1 _2354_ (.B1(_0204_),
    .Y(_0367_),
    .A1(_0365_),
    .A2(_0366_));
 sg13g2_a21oi_1 _2355_ (.A1(_0364_),
    .A2(_0367_),
    .Y(_0368_),
    .B1(_0275_));
 sg13g2_and3_1 _2356_ (.X(_0369_),
    .A(_0206_),
    .B(_0208_),
    .C(_0351_));
 sg13g2_nor4_1 _2357_ (.A(net10),
    .B(_0361_),
    .C(_0368_),
    .D(_0369_),
    .Y(_0370_));
 sg13g2_a221oi_1 _2358_ (.B2(_1184_),
    .C1(net20),
    .B1(_0370_),
    .A1(_0175_),
    .Y(_0080_),
    .A2(_0358_));
 sg13g2_xnor2_1 _2359_ (.Y(_0371_),
    .A(_0207_),
    .B(_0201_));
 sg13g2_nand3_1 _2360_ (.B(_0269_),
    .C(_0273_),
    .A(_0371_),
    .Y(_0372_));
 sg13g2_o21ai_1 _2361_ (.B1(_0372_),
    .Y(_0373_),
    .A1(_0371_),
    .A2(_0351_));
 sg13g2_a21oi_1 _2362_ (.A1(_0206_),
    .A2(_0373_),
    .Y(_0374_),
    .B1(net10));
 sg13g2_o21ai_1 _2363_ (.B1(net45),
    .Y(_0375_),
    .A1(net44),
    .A2(_0635_));
 sg13g2_o21ai_1 _2364_ (.B1(_0375_),
    .Y(_0376_),
    .A1(_0540_),
    .A2(_0605_));
 sg13g2_nor3_1 _2365_ (.A(_0635_),
    .B(_0013_),
    .C(_0349_),
    .Y(_0377_));
 sg13g2_a21o_1 _2366_ (.A2(_0376_),
    .A1(_0349_),
    .B1(_0377_),
    .X(_0378_));
 sg13g2_a221oi_1 _2367_ (.B2(net10),
    .C1(_0576_),
    .B1(_0378_),
    .A1(_1184_),
    .Y(_0081_),
    .A2(_0374_));
 sg13g2_nand2_1 _2368_ (.Y(_0379_),
    .A(_0605_),
    .B(_0013_));
 sg13g2_nand2b_1 _2369_ (.Y(_0380_),
    .B(_0635_),
    .A_N(_0512_));
 sg13g2_mux2_1 _2370_ (.A0(_0379_),
    .A1(_0380_),
    .S(_0349_),
    .X(_0381_));
 sg13g2_mux2_1 _2371_ (.A0(_0333_),
    .A1(_0381_),
    .S(net10),
    .X(_0382_));
 sg13g2_nor2_1 _2372_ (.A(_0576_),
    .B(_0382_),
    .Y(_0082_));
 sg13g2_and2_1 _2373_ (.A(net64),
    .B(_0024_),
    .X(_0083_));
 sg13g2_xnor2_1 _2374_ (.Y(_0383_),
    .A(_1087_),
    .B(net29));
 sg13g2_nor2_1 _2375_ (.A(net53),
    .B(_0383_),
    .Y(_0084_));
 sg13g2_xnor2_1 _2376_ (.Y(_0384_),
    .A(net30),
    .B(_1095_));
 sg13g2_nor2_1 _2377_ (.A(net53),
    .B(_0384_),
    .Y(_0085_));
 sg13g2_nand2_1 _2378_ (.Y(_0385_),
    .A(net30),
    .B(_1095_));
 sg13g2_xnor2_1 _2379_ (.Y(_0386_),
    .A(_1100_),
    .B(_0385_));
 sg13g2_and2_1 _2380_ (.A(_0567_),
    .B(_0386_),
    .X(_0086_));
 sg13g2_nand3_1 _2381_ (.B(net30),
    .C(_1095_),
    .A(_1100_),
    .Y(_0387_));
 sg13g2_xor2_1 _2382_ (.B(_0387_),
    .A(_0983_),
    .X(_0388_));
 sg13g2_nor2_1 _2383_ (.A(net53),
    .B(_0388_),
    .Y(_0087_));
 sg13g2_nand4_1 _2384_ (.B(_1100_),
    .C(net30),
    .A(_0983_),
    .Y(_0389_),
    .D(_1095_));
 sg13g2_xor2_1 _2385_ (.B(_0389_),
    .A(_0982_),
    .X(_0390_));
 sg13g2_nor2_1 _2386_ (.A(net53),
    .B(_0390_),
    .Y(_0088_));
 sg13g2_xnor2_1 _2387_ (.Y(_0391_),
    .A(_0233_),
    .B(\grad1.lfsr[0] ));
 sg13g2_nor2_1 _2388_ (.A(net53),
    .B(_0391_),
    .Y(_0089_));
 sg13g2_nand2_1 _2389_ (.Y(_0392_),
    .A(_0233_),
    .B(\grad1.lfsr[0] ));
 sg13g2_xnor2_1 _2390_ (.Y(_0393_),
    .A(_0230_),
    .B(\grad1.lfsr[1] ));
 sg13g2_xnor2_1 _2391_ (.Y(_0394_),
    .A(_0392_),
    .B(_0393_));
 sg13g2_nor2_1 _2392_ (.A(net53),
    .B(_0394_),
    .Y(_0090_));
 sg13g2_inv_1 _2393_ (.Y(_0395_),
    .A(_0230_));
 sg13g2_a21oi_1 _2394_ (.A1(_0233_),
    .A2(\grad1.lfsr[0] ),
    .Y(_0396_),
    .B1(\grad1.lfsr[1] ));
 sg13g2_nand3_1 _2395_ (.B(\grad1.lfsr[1] ),
    .C(\grad1.lfsr[0] ),
    .A(_0233_),
    .Y(_0397_));
 sg13g2_o21ai_1 _2396_ (.B1(_0397_),
    .Y(_0398_),
    .A1(_0395_),
    .A2(_0396_));
 sg13g2_xor2_1 _2397_ (.B(\grad1.lfsr[2] ),
    .A(\grad1.acc[2] ),
    .X(_0399_));
 sg13g2_xnor2_1 _2398_ (.Y(_0400_),
    .A(_0398_),
    .B(_0399_));
 sg13g2_nor2_1 _2399_ (.A(net53),
    .B(_0400_),
    .Y(_0091_));
 sg13g2_nand2_1 _2400_ (.Y(_0401_),
    .A(\grad1.lfsr[2] ),
    .B(_0398_));
 sg13g2_o21ai_1 _2401_ (.B1(\grad1.acc[2] ),
    .Y(_0402_),
    .A1(\grad1.lfsr[2] ),
    .A2(_0398_));
 sg13g2_xnor2_1 _2402_ (.Y(_0403_),
    .A(net52),
    .B(\grad1.lfsr[3] ));
 sg13g2_and3_1 _2403_ (.X(_0404_),
    .A(_0401_),
    .B(_0402_),
    .C(_0403_));
 sg13g2_a21oi_1 _2404_ (.A1(_0401_),
    .A2(_0402_),
    .Y(_0405_),
    .B1(_0403_));
 sg13g2_nor3_1 _2405_ (.A(_0488_),
    .B(_0404_),
    .C(_0405_),
    .Y(_0092_));
 sg13g2_nand3_1 _2406_ (.B(_0401_),
    .C(_0402_),
    .A(_0563_),
    .Y(_0406_));
 sg13g2_a21oi_1 _2407_ (.A1(_0401_),
    .A2(_0402_),
    .Y(_0407_),
    .B1(_0563_));
 sg13g2_a21o_1 _2408_ (.A2(_0406_),
    .A1(net52),
    .B1(_0407_),
    .X(_0408_));
 sg13g2_xor2_1 _2409_ (.B(_0564_),
    .A(\grad1.acc[4] ),
    .X(_0409_));
 sg13g2_xnor2_1 _2410_ (.Y(_0410_),
    .A(_0408_),
    .B(_0409_));
 sg13g2_nor2_1 _2411_ (.A(net57),
    .B(_0410_),
    .Y(_0093_));
 sg13g2_nand2_1 _2412_ (.Y(_0411_),
    .A(_0564_),
    .B(_0408_));
 sg13g2_o21ai_1 _2413_ (.B1(\grad1.acc[4] ),
    .Y(_0412_),
    .A1(_0564_),
    .A2(_0408_));
 sg13g2_xnor2_1 _2414_ (.Y(_0413_),
    .A(_0264_),
    .B(\grad1.lfsr[5] ));
 sg13g2_and3_1 _2415_ (.X(_0414_),
    .A(_0411_),
    .B(_0412_),
    .C(_0413_));
 sg13g2_a21oi_1 _2416_ (.A1(_0411_),
    .A2(_0412_),
    .Y(_0415_),
    .B1(_0413_));
 sg13g2_nor3_1 _2417_ (.A(_0488_),
    .B(_0414_),
    .C(_0415_),
    .Y(_0094_));
 sg13g2_nand3_1 _2418_ (.B(_0411_),
    .C(_0412_),
    .A(_0565_),
    .Y(_0416_));
 sg13g2_a21oi_1 _2419_ (.A1(_0411_),
    .A2(_0412_),
    .Y(_0417_),
    .B1(_0565_));
 sg13g2_a21oi_2 _2420_ (.B1(_0417_),
    .Y(_0418_),
    .A2(_0416_),
    .A1(_0264_));
 sg13g2_xnor2_1 _2421_ (.Y(_0419_),
    .A(_0305_),
    .B(\grad1.lfsr[6] ));
 sg13g2_xnor2_1 _2422_ (.Y(_0420_),
    .A(_0418_),
    .B(_0419_));
 sg13g2_nor2_1 _2423_ (.A(net57),
    .B(_0420_),
    .Y(_0095_));
 sg13g2_nand2_1 _2424_ (.Y(_0421_),
    .A(_0566_),
    .B(_0418_));
 sg13g2_nor2_1 _2425_ (.A(_0566_),
    .B(_0418_),
    .Y(_0422_));
 sg13g2_a21oi_1 _2426_ (.A1(_0305_),
    .A2(_0421_),
    .Y(_0423_),
    .B1(_0422_));
 sg13g2_xnor2_1 _2427_ (.Y(_0424_),
    .A(\grad1.acc[7] ),
    .B(\grad1.lfsr[7] ));
 sg13g2_xnor2_1 _2428_ (.Y(_0425_),
    .A(_0423_),
    .B(_0424_));
 sg13g2_nor2_1 _2429_ (.A(net57),
    .B(_0425_),
    .Y(_0096_));
 sg13g2_nand2_1 _2430_ (.Y(_0426_),
    .A(\grad1.acc[7] ),
    .B(\grad1.lfsr[7] ));
 sg13g2_nor2_1 _2431_ (.A(\grad1.acc[7] ),
    .B(\grad1.lfsr[7] ),
    .Y(_0427_));
 sg13g2_a21oi_1 _2432_ (.A1(_0423_),
    .A2(_0426_),
    .Y(_0428_),
    .B1(_0427_));
 sg13g2_xor2_1 _2433_ (.B(_0428_),
    .A(_0015_),
    .X(_0429_));
 sg13g2_nor2_1 _2434_ (.A(net57),
    .B(_0429_),
    .Y(_0097_));
 sg13g2_xor2_1 _2435_ (.B(\grad1.lfsr[19] ),
    .A(\grad1.lfsr[15] ),
    .X(_0430_));
 sg13g2_xnor2_1 _2436_ (.Y(_0431_),
    .A(_0564_),
    .B(\grad1.lfsr[3] ));
 sg13g2_xnor2_1 _2437_ (.Y(_0432_),
    .A(\grad1.lfsr[11] ),
    .B(\grad1.lfsr[5] ));
 sg13g2_xnor2_1 _2438_ (.Y(_0433_),
    .A(_0431_),
    .B(_0432_));
 sg13g2_xnor2_1 _2439_ (.Y(_0434_),
    .A(_0430_),
    .B(_0433_));
 sg13g2_nor2_1 _2440_ (.A(net57),
    .B(_0434_),
    .Y(_0098_));
 sg13g2_and2_1 _2441_ (.A(net64),
    .B(\grad1.lfsr[9] ),
    .X(_0099_));
 sg13g2_and2_1 _2442_ (.A(net64),
    .B(\grad1.lfsr[10] ),
    .X(_0100_));
 sg13g2_and2_1 _2443_ (.A(net64),
    .B(\grad1.lfsr[11] ),
    .X(_0101_));
 sg13g2_and2_1 _2444_ (.A(net64),
    .B(\grad1.lfsr[12] ),
    .X(_0102_));
 sg13g2_and2_1 _2445_ (.A(net64),
    .B(\grad1.lfsr[13] ),
    .X(_0025_));
 sg13g2_buf_1 clkbuf_0_clk (.A(clk),
    .X(clknet_0_clk));
 sg13g2_tiehi \UO_OUT[0]$_SDFF_PN0__92  (.L_HI(net92));
 sg13g2_buf_1 _2448_ (.A(net76),
    .X(uio_oe[0]));
 sg13g2_buf_1 _2449_ (.A(net77),
    .X(uio_oe[1]));
 sg13g2_buf_1 _2450_ (.A(net78),
    .X(uio_oe[2]));
 sg13g2_buf_1 _2451_ (.A(net79),
    .X(uio_oe[3]));
 sg13g2_buf_1 _2452_ (.A(net80),
    .X(uio_oe[4]));
 sg13g2_buf_1 _2453_ (.A(net81),
    .X(uio_oe[5]));
 sg13g2_buf_1 _2454_ (.A(net82),
    .X(uio_oe[6]));
 sg13g2_buf_1 _2455_ (.A(net83),
    .X(uio_oe[7]));
 sg13g2_buf_1 _2456_ (.A(net84),
    .X(uio_out[0]));
 sg13g2_buf_1 _2457_ (.A(net85),
    .X(uio_out[1]));
 sg13g2_buf_1 _2458_ (.A(net86),
    .X(uio_out[2]));
 sg13g2_buf_1 _2459_ (.A(net87),
    .X(uio_out[3]));
 sg13g2_buf_1 _2460_ (.A(net88),
    .X(uio_out[4]));
 sg13g2_buf_1 _2461_ (.A(net89),
    .X(uio_out[5]));
 sg13g2_buf_1 _2462_ (.A(net90),
    .X(uio_out[6]));
 sg13g2_buf_1 _2463_ (.A(net91),
    .X(uio_out[7]));
 sg13g2_dfrbp_1 \counter2[0]$_SDFF_PN0_  (.CLK(net74),
    .RESET_B(net100),
    .D(_0083_),
    .Q_N(_0024_),
    .Q(\counter[0] ));
 sg13g2_dfrbp_1 \counter2[1]$_SDFF_PN0_  (.CLK(net74),
    .RESET_B(net101),
    .D(_0084_),
    .Q_N(_1253_),
    .Q(\counter[1] ));
 sg13g2_dfrbp_1 \counter2[2]$_SDFF_PN0_  (.CLK(net74),
    .RESET_B(net102),
    .D(_0085_),
    .Q_N(_0020_),
    .Q(\counter[2] ));
 sg13g2_dfrbp_1 \counter2[3]$_SDFF_PN0_  (.CLK(net74),
    .RESET_B(net103),
    .D(_0086_),
    .Q_N(_0019_),
    .Q(\counter[3] ));
 sg13g2_dfrbp_1 \counter2[4]$_SDFF_PN0_  (.CLK(net74),
    .RESET_B(net104),
    .D(_0087_),
    .Q_N(_0018_),
    .Q(\counter[4] ));
 sg13g2_dfrbp_1 \counter2[5]$_SDFF_PN0_  (.CLK(net74),
    .RESET_B(net105),
    .D(_0088_),
    .Q_N(_0021_),
    .Q(\counter[5] ));
 sg13g2_dfrbp_1 \grad1.acc[0]$_SDFF_PN0_  (.CLK(clknet_4_2_0_clk),
    .RESET_B(net106),
    .D(_0089_),
    .Q_N(_1252_),
    .Q(\grad1.acc[0] ));
 sg13g2_dfrbp_1 \grad1.acc[1]$_SDFF_PN0_  (.CLK(clknet_4_1_0_clk),
    .RESET_B(net107),
    .D(_0090_),
    .Q_N(_1251_),
    .Q(\grad1.acc[1] ));
 sg13g2_dfrbp_1 \grad1.acc[2]$_SDFF_PN0_  (.CLK(clknet_4_0_0_clk),
    .RESET_B(net108),
    .D(_0091_),
    .Q_N(_1250_),
    .Q(\grad1.acc[2] ));
 sg13g2_dfrbp_1 \grad1.acc[3]$_SDFF_PN0_  (.CLK(clknet_4_6_0_clk),
    .RESET_B(net109),
    .D(_0092_),
    .Q_N(_1249_),
    .Q(\grad1.acc[3] ));
 sg13g2_dfrbp_1 \grad1.acc[4]$_SDFF_PN0_  (.CLK(clknet_4_4_0_clk),
    .RESET_B(net110),
    .D(_0093_),
    .Q_N(_0017_),
    .Q(\grad1.acc[4] ));
 sg13g2_dfrbp_1 \grad1.acc[5]$_SDFF_PN0_  (.CLK(clknet_4_6_0_clk),
    .RESET_B(net111),
    .D(_0094_),
    .Q_N(_1248_),
    .Q(\grad1.acc[5] ));
 sg13g2_dfrbp_1 \grad1.acc[6]$_SDFF_PN0_  (.CLK(clknet_4_6_0_clk),
    .RESET_B(net112),
    .D(_0095_),
    .Q_N(_0016_),
    .Q(\grad1.acc[6] ));
 sg13g2_dfrbp_1 \grad1.acc[7]$_SDFF_PN0_  (.CLK(clknet_4_7_0_clk),
    .RESET_B(net113),
    .D(_0096_),
    .Q_N(_1247_),
    .Q(\grad1.acc[7] ));
 sg13g2_dfrbp_1 \grad1.acc[8]$_SDFF_PN0_  (.CLK(clknet_4_7_0_clk),
    .RESET_B(net114),
    .D(_0097_),
    .Q_N(_0015_),
    .Q(\grad1.acc[8] ));
 sg13g2_dfrbp_1 \grad1.lfsr[0]$_SDFF_PN0_  (.CLK(clknet_4_0_0_clk),
    .RESET_B(net115),
    .D(_0098_),
    .Q_N(_1246_),
    .Q(\grad1.lfsr[0] ));
 sg13g2_dfrbp_1 \grad1.lfsr[10]$_SDFF_PN0_  (.CLK(clknet_4_4_0_clk),
    .RESET_B(net116),
    .D(_0099_),
    .Q_N(_1245_),
    .Q(\grad1.lfsr[10] ));
 sg13g2_dfrbp_1 \grad1.lfsr[11]$_SDFF_PN0_  (.CLK(clknet_4_0_0_clk),
    .RESET_B(net117),
    .D(_0100_),
    .Q_N(_1244_),
    .Q(\grad1.lfsr[11] ));
 sg13g2_dfrbp_1 \grad1.lfsr[12]$_SDFF_PN0_  (.CLK(clknet_4_0_0_clk),
    .RESET_B(net118),
    .D(_0101_),
    .Q_N(_1243_),
    .Q(\grad1.lfsr[12] ));
 sg13g2_dfrbp_1 \grad1.lfsr[13]$_SDFF_PN0_  (.CLK(clknet_4_5_0_clk),
    .RESET_B(net119),
    .D(_0102_),
    .Q_N(_1242_),
    .Q(\grad1.lfsr[13] ));
 sg13g2_dfrbp_1 \grad1.lfsr[14]$_SDFF_PN0_  (.CLK(clknet_4_5_0_clk),
    .RESET_B(net120),
    .D(_0025_),
    .Q_N(_1241_),
    .Q(\grad1.lfsr[14] ));
 sg13g2_dfrbp_1 \grad1.lfsr[15]$_SDFF_PN0_  (.CLK(clknet_4_1_0_clk),
    .RESET_B(net121),
    .D(_0026_),
    .Q_N(_1240_),
    .Q(\grad1.lfsr[15] ));
 sg13g2_dfrbp_1 \grad1.lfsr[16]$_SDFF_PN0_  (.CLK(clknet_4_1_0_clk),
    .RESET_B(net122),
    .D(_0027_),
    .Q_N(_1239_),
    .Q(\grad1.lfsr[16] ));
 sg13g2_dfrbp_1 \grad1.lfsr[17]$_SDFF_PN0_  (.CLK(clknet_4_2_0_clk),
    .RESET_B(net123),
    .D(_0028_),
    .Q_N(_1238_),
    .Q(\grad1.lfsr[17] ));
 sg13g2_dfrbp_1 \grad1.lfsr[18]$_SDFF_PN0_  (.CLK(clknet_4_2_0_clk),
    .RESET_B(net124),
    .D(_0029_),
    .Q_N(_1237_),
    .Q(\grad1.lfsr[18] ));
 sg13g2_dfrbp_1 \grad1.lfsr[19]$_SDFF_PN0_  (.CLK(clknet_4_2_0_clk),
    .RESET_B(net125),
    .D(_0030_),
    .Q_N(_1236_),
    .Q(\grad1.lfsr[19] ));
 sg13g2_dfrbp_1 \grad1.lfsr[1]$_SDFF_PN0_  (.CLK(clknet_4_1_0_clk),
    .RESET_B(net126),
    .D(_0031_),
    .Q_N(_1235_),
    .Q(\grad1.lfsr[1] ));
 sg13g2_dfrbp_1 \grad1.lfsr[2]$_SDFF_PN0_  (.CLK(clknet_4_5_0_clk),
    .RESET_B(net127),
    .D(_0032_),
    .Q_N(_1234_),
    .Q(\grad1.lfsr[2] ));
 sg13g2_dfrbp_1 \grad1.lfsr[3]$_SDFF_PN0_  (.CLK(clknet_4_4_0_clk),
    .RESET_B(net128),
    .D(_0033_),
    .Q_N(_1233_),
    .Q(\grad1.lfsr[3] ));
 sg13g2_dfrbp_1 \grad1.lfsr[4]$_SDFF_PN0_  (.CLK(clknet_4_0_0_clk),
    .RESET_B(net129),
    .D(_0034_),
    .Q_N(_1232_),
    .Q(\grad1.lfsr[4] ));
 sg13g2_dfrbp_1 \grad1.lfsr[5]$_SDFF_PN0_  (.CLK(clknet_4_4_0_clk),
    .RESET_B(net130),
    .D(_0035_),
    .Q_N(_1231_),
    .Q(\grad1.lfsr[5] ));
 sg13g2_dfrbp_1 \grad1.lfsr[6]$_SDFF_PN0_  (.CLK(clknet_4_4_0_clk),
    .RESET_B(net131),
    .D(_0036_),
    .Q_N(_1230_),
    .Q(\grad1.lfsr[6] ));
 sg13g2_dfrbp_1 \grad1.lfsr[7]$_SDFF_PN0_  (.CLK(clknet_4_6_0_clk),
    .RESET_B(net132),
    .D(_0037_),
    .Q_N(_1229_),
    .Q(\grad1.lfsr[7] ));
 sg13g2_dfrbp_1 \grad1.lfsr[8]$_SDFF_PN0_  (.CLK(clknet_4_5_0_clk),
    .RESET_B(net133),
    .D(_0038_),
    .Q_N(_1228_),
    .Q(\grad1.lfsr[8] ));
 sg13g2_dfrbp_1 \grad1.lfsr[9]$_SDFF_PN0_  (.CLK(clknet_4_5_0_clk),
    .RESET_B(net134),
    .D(_0039_),
    .Q_N(_1227_),
    .Q(\grad1.lfsr[9] ));
 sg13g2_dfrbp_1 \hvsync_gen.hpos[0]$_SDFF_PP0_  (.CLK(clknet_4_3_0_clk),
    .RESET_B(net135),
    .D(_0040_),
    .Q_N(_0022_),
    .Q(\hvsync_gen.hpos[0] ));
 sg13g2_dfrbp_1 \hvsync_gen.hpos[1]$_SDFF_PP0_  (.CLK(clknet_4_8_0_clk),
    .RESET_B(net136),
    .D(_0041_),
    .Q_N(_1226_),
    .Q(\hvsync_gen.hpos[1] ));
 sg13g2_dfrbp_1 \hvsync_gen.hpos[2]$_SDFF_PP0_  (.CLK(clknet_4_10_0_clk),
    .RESET_B(net137),
    .D(_0042_),
    .Q_N(_1225_),
    .Q(\hvsync_gen.hpos[2] ));
 sg13g2_dfrbp_1 \hvsync_gen.hpos[3]$_SDFF_PP0_  (.CLK(clknet_4_8_0_clk),
    .RESET_B(net138),
    .D(_0043_),
    .Q_N(_1224_),
    .Q(\hvsync_gen.hpos[3] ));
 sg13g2_dfrbp_1 \hvsync_gen.hpos[4]$_SDFF_PP0_  (.CLK(clknet_4_11_0_clk),
    .RESET_B(net139),
    .D(_0044_),
    .Q_N(_1223_),
    .Q(\hvsync_gen.hpos[4] ));
 sg13g2_dfrbp_1 \hvsync_gen.hpos[5]$_SDFF_PP0_  (.CLK(clknet_4_12_0_clk),
    .RESET_B(net140),
    .D(_0045_),
    .Q_N(_1222_),
    .Q(\hvsync_gen.hpos[5] ));
 sg13g2_dfrbp_1 \hvsync_gen.hpos[6]$_SDFF_PP0_  (.CLK(clknet_4_14_0_clk),
    .RESET_B(net141),
    .D(_0046_),
    .Q_N(_1221_),
    .Q(\hvsync_gen.hpos[6] ));
 sg13g2_dfrbp_1 \hvsync_gen.hpos[7]$_SDFF_PP0_  (.CLK(clknet_4_9_0_clk),
    .RESET_B(net142),
    .D(_0047_),
    .Q_N(_1220_),
    .Q(\hvsync_gen.hpos[7] ));
 sg13g2_dfrbp_1 \hvsync_gen.hpos[8]$_SDFF_PP0_  (.CLK(clknet_4_12_0_clk),
    .RESET_B(net143),
    .D(_0048_),
    .Q_N(_0014_),
    .Q(\hvsync_gen.hpos[8] ));
 sg13g2_dfrbp_1 \hvsync_gen.hpos[9]$_SDFF_PP0_  (.CLK(clknet_4_12_0_clk),
    .RESET_B(net144),
    .D(_0049_),
    .Q_N(_0008_),
    .Q(\hvsync_gen.hpos[9] ));
 sg13g2_dfrbp_1 \hvsync_gen.hsync$_DFF_P_  (.CLK(clknet_4_7_0_clk),
    .RESET_B(net145),
    .D(_0000_),
    .Q_N(_1219_),
    .Q(hsync));
 sg13g2_dfrbp_1 \hvsync_gen.vpos[0]$_SDFFCE_PP0P_  (.CLK(clknet_4_1_0_clk),
    .RESET_B(net146),
    .D(_0050_),
    .Q_N(_0023_),
    .Q(\hvsync_gen.vpos[0] ));
 sg13g2_dfrbp_1 \hvsync_gen.vpos[1]$_SDFFCE_PP0P_  (.CLK(clknet_4_2_0_clk),
    .RESET_B(net147),
    .D(_0051_),
    .Q_N(_1218_),
    .Q(\hvsync_gen.vpos[1] ));
 sg13g2_dfrbp_1 \hvsync_gen.vpos[2]$_SDFFCE_PP0P_  (.CLK(clknet_4_3_0_clk),
    .RESET_B(net148),
    .D(_0052_),
    .Q_N(_1217_),
    .Q(\hvsync_gen.vpos[2] ));
 sg13g2_dfrbp_1 \hvsync_gen.vpos[3]$_SDFFCE_PP0P_  (.CLK(clknet_4_8_0_clk),
    .RESET_B(net149),
    .D(_0053_),
    .Q_N(_1216_),
    .Q(\hvsync_gen.vpos[3] ));
 sg13g2_dfrbp_1 \hvsync_gen.vpos[4]$_SDFFCE_PP0P_  (.CLK(clknet_4_3_0_clk),
    .RESET_B(net150),
    .D(_0054_),
    .Q_N(_1215_),
    .Q(\hvsync_gen.vpos[4] ));
 sg13g2_dfrbp_1 \hvsync_gen.vpos[5]$_SDFFCE_PP0P_  (.CLK(clknet_4_6_0_clk),
    .RESET_B(net151),
    .D(_0055_),
    .Q_N(_1214_),
    .Q(\hvsync_gen.vpos[5] ));
 sg13g2_dfrbp_1 \hvsync_gen.vpos[6]$_SDFFCE_PP0P_  (.CLK(clknet_4_9_0_clk),
    .RESET_B(net152),
    .D(_0056_),
    .Q_N(_1213_),
    .Q(\hvsync_gen.vpos[6] ));
 sg13g2_dfrbp_1 \hvsync_gen.vpos[7]$_SDFFCE_PP0P_  (.CLK(clknet_4_9_0_clk),
    .RESET_B(net153),
    .D(_0057_),
    .Q_N(_0012_),
    .Q(\hvsync_gen.vpos[7] ));
 sg13g2_dfrbp_1 \hvsync_gen.vpos[8]$_SDFFCE_PP0P_  (.CLK(clknet_4_9_0_clk),
    .RESET_B(net154),
    .D(_0058_),
    .Q_N(_0013_),
    .Q(\hvsync_gen.vpos[8] ));
 sg13g2_dfrbp_1 \hvsync_gen.vpos[9]$_SDFFCE_PP0P_  (.CLK(clknet_4_9_0_clk),
    .RESET_B(net155),
    .D(_0059_),
    .Q_N(_1262_),
    .Q(\hvsync_gen.vpos[9] ));
 sg13g2_dfrbp_1 \hvsync_gen.vsync$_DFF_P_  (.CLK(clknet_4_11_0_clk),
    .RESET_B(net156),
    .D(_0001_),
    .Q_N(_1212_),
    .Q(\hvsync_gen.vsync ));
 sg13g2_dfrbp_1 \r[0]$_SDFFE_PN0P_  (.CLK(clknet_4_8_0_clk),
    .RESET_B(net157),
    .D(_0060_),
    .Q_N(_0010_),
    .Q(\r[0] ));
 sg13g2_dfrbp_1 \r[10]$_SDFFE_PN0P_  (.CLK(clknet_4_12_0_clk),
    .RESET_B(net158),
    .D(_0061_),
    .Q_N(_0003_),
    .Q(\r[10] ));
 sg13g2_dfrbp_1 \r[11]$_SDFFE_PN0P_  (.CLK(clknet_4_14_0_clk),
    .RESET_B(net159),
    .D(_0062_),
    .Q_N(_0004_),
    .Q(\r[11] ));
 sg13g2_dfrbp_1 \r[12]$_SDFFE_PN0P_  (.CLK(clknet_4_15_0_clk),
    .RESET_B(net160),
    .D(_0063_),
    .Q_N(_0005_),
    .Q(\r[12] ));
 sg13g2_dfrbp_1 \r[13]$_SDFFE_PN0P_  (.CLK(clknet_4_15_0_clk),
    .RESET_B(net161),
    .D(_0064_),
    .Q_N(_0006_),
    .Q(\r[13] ));
 sg13g2_dfrbp_1 \r[14]$_SDFFE_PN0P_  (.CLK(clknet_4_15_0_clk),
    .RESET_B(net162),
    .D(_0065_),
    .Q_N(_0009_),
    .Q(\r[14] ));
 sg13g2_dfrbp_1 \r[15]$_SDFFE_PN0P_  (.CLK(clknet_4_15_0_clk),
    .RESET_B(net163),
    .D(_0066_),
    .Q_N(_0007_),
    .Q(\r[15] ));
 sg13g2_dfrbp_1 \r[16]$_SDFFE_PN0P_  (.CLK(clknet_4_14_0_clk),
    .RESET_B(net164),
    .D(_0067_),
    .Q_N(_0011_),
    .Q(\r[16] ));
 sg13g2_dfrbp_1 \r[1]$_SDFFE_PN0P_  (.CLK(clknet_4_8_0_clk),
    .RESET_B(net165),
    .D(_0068_),
    .Q_N(_1211_),
    .Q(\r[1] ));
 sg13g2_dfrbp_1 \r[2]$_SDFFE_PN0P_  (.CLK(clknet_4_10_0_clk),
    .RESET_B(net166),
    .D(_0069_),
    .Q_N(_1210_),
    .Q(\r[2] ));
 sg13g2_dfrbp_1 \r[3]$_SDFFE_PN0P_  (.CLK(clknet_4_10_0_clk),
    .RESET_B(net167),
    .D(_0070_),
    .Q_N(_1209_),
    .Q(\r[3] ));
 sg13g2_dfrbp_1 \r[4]$_SDFFE_PN0P_  (.CLK(clknet_4_10_0_clk),
    .RESET_B(net168),
    .D(_0071_),
    .Q_N(_1208_),
    .Q(\r[4] ));
 sg13g2_dfrbp_1 \r[5]$_SDFFE_PN0P_  (.CLK(clknet_4_10_0_clk),
    .RESET_B(net169),
    .D(_0072_),
    .Q_N(_1207_),
    .Q(\r[5] ));
 sg13g2_dfrbp_1 \r[6]$_SDFFE_PN0P_  (.CLK(clknet_4_11_0_clk),
    .RESET_B(net170),
    .D(_0073_),
    .Q_N(_1206_),
    .Q(\r[6] ));
 sg13g2_dfrbp_1 \r[7]$_SDFFE_PN0P_  (.CLK(clknet_4_11_0_clk),
    .RESET_B(net171),
    .D(_0074_),
    .Q_N(_1205_),
    .Q(\r[7] ));
 sg13g2_dfrbp_1 \r[8]$_SDFFE_PN0P_  (.CLK(clknet_4_14_0_clk),
    .RESET_B(net172),
    .D(_0075_),
    .Q_N(_0002_),
    .Q(\r[8] ));
 sg13g2_dfrbp_1 \r[9]$_SDFFE_PN0P_  (.CLK(clknet_4_14_0_clk),
    .RESET_B(net173),
    .D(_0076_),
    .Q_N(_1204_),
    .Q(\r[9] ));
 sg13g2_buf_1 input1 (.A(rst_n),
    .X(net1));
 sg13g2_buf_1 output2 (.A(net2),
    .X(uo_out[0]));
 sg13g2_buf_1 output3 (.A(net3),
    .X(uo_out[1]));
 sg13g2_buf_1 output4 (.A(net4),
    .X(uo_out[2]));
 sg13g2_buf_1 output5 (.A(net5),
    .X(uo_out[3]));
 sg13g2_buf_1 output6 (.A(net6),
    .X(uo_out[4]));
 sg13g2_buf_1 output7 (.A(net7),
    .X(uo_out[5]));
 sg13g2_buf_1 output8 (.A(net8),
    .X(uo_out[6]));
 sg13g2_buf_1 output9 (.A(net9),
    .X(uo_out[7]));
 sg13g2_buf_2 fanout10 (.A(_0175_),
    .X(net10));
 sg13g2_buf_2 fanout11 (.A(_0725_),
    .X(net11));
 sg13g2_buf_2 fanout12 (.A(_0584_),
    .X(net12));
 sg13g2_buf_2 fanout13 (.A(_1103_),
    .X(net13));
 sg13g2_buf_2 fanout14 (.A(_1071_),
    .X(net14));
 sg13g2_buf_2 fanout15 (.A(_1027_),
    .X(net15));
 sg13g2_buf_2 fanout16 (.A(_0721_),
    .X(net16));
 sg13g2_buf_2 fanout17 (.A(_0253_),
    .X(net17));
 sg13g2_buf_2 fanout18 (.A(_0716_),
    .X(net18));
 sg13g2_buf_2 fanout19 (.A(_0582_),
    .X(net19));
 sg13g2_buf_2 fanout20 (.A(_0576_),
    .X(net20));
 sg13g2_buf_2 fanout21 (.A(_0741_),
    .X(net21));
 sg13g2_buf_2 fanout22 (.A(_0573_),
    .X(net22));
 sg13g2_buf_2 fanout23 (.A(_0998_),
    .X(net23));
 sg13g2_buf_2 fanout24 (.A(_1093_),
    .X(net24));
 sg13g2_buf_2 fanout25 (.A(_0479_),
    .X(net25));
 sg13g2_buf_2 fanout26 (.A(_0457_),
    .X(net26));
 sg13g2_buf_2 fanout27 (.A(_0454_),
    .X(net27));
 sg13g2_buf_2 fanout28 (.A(_0448_),
    .X(net28));
 sg13g2_buf_2 fanout29 (.A(_1085_),
    .X(net29));
 sg13g2_buf_2 fanout30 (.A(_1084_),
    .X(net30));
 sg13g2_buf_2 fanout31 (.A(_0738_),
    .X(net31));
 sg13g2_buf_2 fanout32 (.A(_0702_),
    .X(net32));
 sg13g2_buf_2 fanout33 (.A(_0570_),
    .X(net33));
 sg13g2_buf_2 fanout34 (.A(_0569_),
    .X(net34));
 sg13g2_buf_2 fanout35 (.A(_0497_),
    .X(net35));
 sg13g2_buf_2 fanout36 (.A(_0495_),
    .X(net36));
 sg13g2_buf_2 fanout37 (.A(_0492_),
    .X(net37));
 sg13g2_buf_2 fanout38 (.A(_0490_),
    .X(net38));
 sg13g2_buf_2 fanout39 (.A(_0483_),
    .X(net39));
 sg13g2_buf_2 fanout40 (.A(_0481_),
    .X(net40));
 sg13g2_buf_2 fanout41 (.A(_0475_),
    .X(net41));
 sg13g2_buf_2 fanout42 (.A(_0473_),
    .X(net42));
 sg13g2_buf_2 fanout43 (.A(_0467_),
    .X(net43));
 sg13g2_buf_2 fanout44 (.A(_0461_),
    .X(net44));
 sg13g2_buf_2 fanout45 (.A(_0459_),
    .X(net45));
 sg13g2_buf_2 fanout46 (.A(_0456_),
    .X(net46));
 sg13g2_buf_2 fanout47 (.A(_0453_),
    .X(net47));
 sg13g2_buf_2 fanout48 (.A(_0447_),
    .X(net48));
 sg13g2_buf_2 fanout49 (.A(_0440_),
    .X(net49));
 sg13g2_buf_2 fanout50 (.A(_0438_),
    .X(net50));
 sg13g2_buf_2 fanout51 (.A(_0436_),
    .X(net51));
 sg13g2_buf_2 fanout52 (.A(_0240_),
    .X(net52));
 sg13g2_buf_2 fanout53 (.A(_0902_),
    .X(net53));
 sg13g2_buf_2 fanout54 (.A(_0838_),
    .X(net54));
 sg13g2_buf_2 fanout55 (.A(_0818_),
    .X(net55));
 sg13g2_buf_2 fanout56 (.A(_0760_),
    .X(net56));
 sg13g2_buf_2 fanout57 (.A(_0700_),
    .X(net57));
 sg13g2_buf_2 fanout58 (.A(_0689_),
    .X(net58));
 sg13g2_buf_2 fanout59 (.A(_0648_),
    .X(net59));
 sg13g2_buf_2 fanout60 (.A(_0627_),
    .X(net60));
 sg13g2_buf_2 fanout61 (.A(_0622_),
    .X(net61));
 sg13g2_buf_2 fanout62 (.A(_0616_),
    .X(net62));
 sg13g2_buf_2 fanout63 (.A(_0593_),
    .X(net63));
 sg13g2_buf_2 fanout64 (.A(_0567_),
    .X(net64));
 sg13g2_buf_2 fanout65 (.A(_0556_),
    .X(net65));
 sg13g2_buf_2 fanout66 (.A(_0518_),
    .X(net66));
 sg13g2_buf_2 fanout67 (.A(_0494_),
    .X(net67));
 sg13g2_buf_2 fanout68 (.A(_0470_),
    .X(net68));
 sg13g2_buf_2 fanout69 (.A(_0469_),
    .X(net69));
 sg13g2_buf_2 fanout70 (.A(_0443_),
    .X(net70));
 sg13g2_buf_2 fanout71 (.A(_0442_),
    .X(net71));
 sg13g2_buf_2 fanout72 (.A(_0439_),
    .X(net72));
 sg13g2_buf_2 fanout73 (.A(_0437_),
    .X(net73));
 sg13g2_buf_2 fanout74 (.A(\hvsync_gen.vsync ),
    .X(net74));
 sg13g2_buf_2 fanout75 (.A(_0506_),
    .X(net75));
 sg13g2_tielo _2448__76 (.L_LO(net76));
 sg13g2_tielo _2449__77 (.L_LO(net77));
 sg13g2_tielo _2450__78 (.L_LO(net78));
 sg13g2_tielo _2451__79 (.L_LO(net79));
 sg13g2_tielo _2452__80 (.L_LO(net80));
 sg13g2_tielo _2453__81 (.L_LO(net81));
 sg13g2_tielo _2454__82 (.L_LO(net82));
 sg13g2_tielo _2455__83 (.L_LO(net83));
 sg13g2_tielo _2456__84 (.L_LO(net84));
 sg13g2_tielo _2457__85 (.L_LO(net85));
 sg13g2_tielo _2458__86 (.L_LO(net86));
 sg13g2_tielo _2459__87 (.L_LO(net87));
 sg13g2_tielo _2460__88 (.L_LO(net88));
 sg13g2_tielo _2461__89 (.L_LO(net89));
 sg13g2_tielo _2462__90 (.L_LO(net90));
 sg13g2_tielo _2463__91 (.L_LO(net91));
 sg13g2_tiehi \UO_OUT[1]$_SDFF_PN0__93  (.L_HI(net93));
 sg13g2_tiehi \UO_OUT[2]$_SDFF_PN0__94  (.L_HI(net94));
 sg13g2_tiehi \UO_OUT[3]$_DFF_P__95  (.L_HI(net95));
 sg13g2_tiehi \UO_OUT[4]$_SDFF_PN0__96  (.L_HI(net96));
 sg13g2_tiehi \UO_OUT[5]$_SDFF_PN0__97  (.L_HI(net97));
 sg13g2_tiehi \UO_OUT[6]$_SDFF_PN0__98  (.L_HI(net98));
 sg13g2_tiehi \UO_OUT[7]$_DFF_P__99  (.L_HI(net99));
 sg13g2_tiehi \counter2[0]$_SDFF_PN0__100  (.L_HI(net100));
 sg13g2_tiehi \counter2[1]$_SDFF_PN0__101  (.L_HI(net101));
 sg13g2_tiehi \counter2[2]$_SDFF_PN0__102  (.L_HI(net102));
 sg13g2_tiehi \counter2[3]$_SDFF_PN0__103  (.L_HI(net103));
 sg13g2_tiehi \counter2[4]$_SDFF_PN0__104  (.L_HI(net104));
 sg13g2_tiehi \counter2[5]$_SDFF_PN0__105  (.L_HI(net105));
 sg13g2_tiehi \grad1.acc[0]$_SDFF_PN0__106  (.L_HI(net106));
 sg13g2_tiehi \grad1.acc[1]$_SDFF_PN0__107  (.L_HI(net107));
 sg13g2_tiehi \grad1.acc[2]$_SDFF_PN0__108  (.L_HI(net108));
 sg13g2_tiehi \grad1.acc[3]$_SDFF_PN0__109  (.L_HI(net109));
 sg13g2_tiehi \grad1.acc[4]$_SDFF_PN0__110  (.L_HI(net110));
 sg13g2_tiehi \grad1.acc[5]$_SDFF_PN0__111  (.L_HI(net111));
 sg13g2_tiehi \grad1.acc[6]$_SDFF_PN0__112  (.L_HI(net112));
 sg13g2_tiehi \grad1.acc[7]$_SDFF_PN0__113  (.L_HI(net113));
 sg13g2_tiehi \grad1.acc[8]$_SDFF_PN0__114  (.L_HI(net114));
 sg13g2_tiehi \grad1.lfsr[0]$_SDFF_PN0__115  (.L_HI(net115));
 sg13g2_tiehi \grad1.lfsr[10]$_SDFF_PN0__116  (.L_HI(net116));
 sg13g2_tiehi \grad1.lfsr[11]$_SDFF_PN0__117  (.L_HI(net117));
 sg13g2_tiehi \grad1.lfsr[12]$_SDFF_PN0__118  (.L_HI(net118));
 sg13g2_tiehi \grad1.lfsr[13]$_SDFF_PN0__119  (.L_HI(net119));
 sg13g2_tiehi \grad1.lfsr[14]$_SDFF_PN0__120  (.L_HI(net120));
 sg13g2_tiehi \grad1.lfsr[15]$_SDFF_PN0__121  (.L_HI(net121));
 sg13g2_tiehi \grad1.lfsr[16]$_SDFF_PN0__122  (.L_HI(net122));
 sg13g2_tiehi \grad1.lfsr[17]$_SDFF_PN0__123  (.L_HI(net123));
 sg13g2_tiehi \grad1.lfsr[18]$_SDFF_PN0__124  (.L_HI(net124));
 sg13g2_tiehi \grad1.lfsr[19]$_SDFF_PN0__125  (.L_HI(net125));
 sg13g2_tiehi \grad1.lfsr[1]$_SDFF_PN0__126  (.L_HI(net126));
 sg13g2_tiehi \grad1.lfsr[2]$_SDFF_PN0__127  (.L_HI(net127));
 sg13g2_tiehi \grad1.lfsr[3]$_SDFF_PN0__128  (.L_HI(net128));
 sg13g2_tiehi \grad1.lfsr[4]$_SDFF_PN0__129  (.L_HI(net129));
 sg13g2_tiehi \grad1.lfsr[5]$_SDFF_PN0__130  (.L_HI(net130));
 sg13g2_tiehi \grad1.lfsr[6]$_SDFF_PN0__131  (.L_HI(net131));
 sg13g2_tiehi \grad1.lfsr[7]$_SDFF_PN0__132  (.L_HI(net132));
 sg13g2_tiehi \grad1.lfsr[8]$_SDFF_PN0__133  (.L_HI(net133));
 sg13g2_tiehi \grad1.lfsr[9]$_SDFF_PN0__134  (.L_HI(net134));
 sg13g2_tiehi \hvsync_gen.hpos[0]$_SDFF_PP0__135  (.L_HI(net135));
 sg13g2_tiehi \hvsync_gen.hpos[1]$_SDFF_PP0__136  (.L_HI(net136));
 sg13g2_tiehi \hvsync_gen.hpos[2]$_SDFF_PP0__137  (.L_HI(net137));
 sg13g2_tiehi \hvsync_gen.hpos[3]$_SDFF_PP0__138  (.L_HI(net138));
 sg13g2_tiehi \hvsync_gen.hpos[4]$_SDFF_PP0__139  (.L_HI(net139));
 sg13g2_tiehi \hvsync_gen.hpos[5]$_SDFF_PP0__140  (.L_HI(net140));
 sg13g2_tiehi \hvsync_gen.hpos[6]$_SDFF_PP0__141  (.L_HI(net141));
 sg13g2_tiehi \hvsync_gen.hpos[7]$_SDFF_PP0__142  (.L_HI(net142));
 sg13g2_tiehi \hvsync_gen.hpos[8]$_SDFF_PP0__143  (.L_HI(net143));
 sg13g2_tiehi \hvsync_gen.hpos[9]$_SDFF_PP0__144  (.L_HI(net144));
 sg13g2_tiehi \hvsync_gen.hsync$_DFF_P__145  (.L_HI(net145));
 sg13g2_tiehi \hvsync_gen.vpos[0]$_SDFFCE_PP0P__146  (.L_HI(net146));
 sg13g2_tiehi \hvsync_gen.vpos[1]$_SDFFCE_PP0P__147  (.L_HI(net147));
 sg13g2_tiehi \hvsync_gen.vpos[2]$_SDFFCE_PP0P__148  (.L_HI(net148));
 sg13g2_tiehi \hvsync_gen.vpos[3]$_SDFFCE_PP0P__149  (.L_HI(net149));
 sg13g2_tiehi \hvsync_gen.vpos[4]$_SDFFCE_PP0P__150  (.L_HI(net150));
 sg13g2_tiehi \hvsync_gen.vpos[5]$_SDFFCE_PP0P__151  (.L_HI(net151));
 sg13g2_tiehi \hvsync_gen.vpos[6]$_SDFFCE_PP0P__152  (.L_HI(net152));
 sg13g2_tiehi \hvsync_gen.vpos[7]$_SDFFCE_PP0P__153  (.L_HI(net153));
 sg13g2_tiehi \hvsync_gen.vpos[8]$_SDFFCE_PP0P__154  (.L_HI(net154));
 sg13g2_tiehi \hvsync_gen.vpos[9]$_SDFFCE_PP0P__155  (.L_HI(net155));
 sg13g2_tiehi \hvsync_gen.vsync$_DFF_P__156  (.L_HI(net156));
 sg13g2_tiehi \r[0]$_SDFFE_PN0P__157  (.L_HI(net157));
 sg13g2_tiehi \r[10]$_SDFFE_PN0P__158  (.L_HI(net158));
 sg13g2_tiehi \r[11]$_SDFFE_PN0P__159  (.L_HI(net159));
 sg13g2_tiehi \r[12]$_SDFFE_PN0P__160  (.L_HI(net160));
 sg13g2_tiehi \r[13]$_SDFFE_PN0P__161  (.L_HI(net161));
 sg13g2_tiehi \r[14]$_SDFFE_PN0P__162  (.L_HI(net162));
 sg13g2_tiehi \r[15]$_SDFFE_PN0P__163  (.L_HI(net163));
 sg13g2_tiehi \r[16]$_SDFFE_PN0P__164  (.L_HI(net164));
 sg13g2_tiehi \r[1]$_SDFFE_PN0P__165  (.L_HI(net165));
 sg13g2_tiehi \r[2]$_SDFFE_PN0P__166  (.L_HI(net166));
 sg13g2_tiehi \r[3]$_SDFFE_PN0P__167  (.L_HI(net167));
 sg13g2_tiehi \r[4]$_SDFFE_PN0P__168  (.L_HI(net168));
 sg13g2_tiehi \r[5]$_SDFFE_PN0P__169  (.L_HI(net169));
 sg13g2_tiehi \r[6]$_SDFFE_PN0P__170  (.L_HI(net170));
 sg13g2_tiehi \r[7]$_SDFFE_PN0P__171  (.L_HI(net171));
 sg13g2_tiehi \r[8]$_SDFFE_PN0P__172  (.L_HI(net172));
 sg13g2_tiehi \r[9]$_SDFFE_PN0P__173  (.L_HI(net173));
 sg13g2_buf_2 clkbuf_4_0_0_clk (.A(clknet_0_clk),
    .X(clknet_4_0_0_clk));
 sg13g2_buf_2 clkbuf_4_1_0_clk (.A(clknet_0_clk),
    .X(clknet_4_1_0_clk));
 sg13g2_buf_2 clkbuf_4_2_0_clk (.A(clknet_0_clk),
    .X(clknet_4_2_0_clk));
 sg13g2_buf_2 clkbuf_4_3_0_clk (.A(clknet_0_clk),
    .X(clknet_4_3_0_clk));
 sg13g2_buf_2 clkbuf_4_4_0_clk (.A(clknet_0_clk),
    .X(clknet_4_4_0_clk));
 sg13g2_buf_2 clkbuf_4_5_0_clk (.A(clknet_0_clk),
    .X(clknet_4_5_0_clk));
 sg13g2_buf_2 clkbuf_4_6_0_clk (.A(clknet_0_clk),
    .X(clknet_4_6_0_clk));
 sg13g2_buf_2 clkbuf_4_7_0_clk (.A(clknet_0_clk),
    .X(clknet_4_7_0_clk));
 sg13g2_buf_2 clkbuf_4_8_0_clk (.A(clknet_0_clk),
    .X(clknet_4_8_0_clk));
 sg13g2_buf_2 clkbuf_4_9_0_clk (.A(clknet_0_clk),
    .X(clknet_4_9_0_clk));
 sg13g2_buf_2 clkbuf_4_10_0_clk (.A(clknet_0_clk),
    .X(clknet_4_10_0_clk));
 sg13g2_buf_2 clkbuf_4_11_0_clk (.A(clknet_0_clk),
    .X(clknet_4_11_0_clk));
 sg13g2_buf_2 clkbuf_4_12_0_clk (.A(clknet_0_clk),
    .X(clknet_4_12_0_clk));
 sg13g2_buf_2 clkbuf_4_13_0_clk (.A(clknet_0_clk),
    .X(clknet_4_13_0_clk));
 sg13g2_buf_2 clkbuf_4_14_0_clk (.A(clknet_0_clk),
    .X(clknet_4_14_0_clk));
 sg13g2_buf_2 clkbuf_4_15_0_clk (.A(clknet_0_clk),
    .X(clknet_4_15_0_clk));
 sg13g2_inv_1 clkload0 (.A(clknet_4_3_0_clk));
 sg13g2_inv_1 clkload1 (.A(clknet_4_7_0_clk));
 sg13g2_inv_1 clkload2 (.A(clknet_4_11_0_clk));
 sg13g2_inv_1 clkload3 (.A(clknet_4_15_0_clk));
 sg13g2_decap_8 FILLER_0_0 ();
 sg13g2_decap_8 FILLER_0_7 ();
 sg13g2_decap_8 FILLER_0_14 ();
 sg13g2_decap_8 FILLER_0_21 ();
 sg13g2_decap_8 FILLER_0_28 ();
 sg13g2_decap_8 FILLER_0_35 ();
 sg13g2_decap_8 FILLER_0_42 ();
 sg13g2_decap_8 FILLER_0_49 ();
 sg13g2_decap_8 FILLER_0_56 ();
 sg13g2_decap_8 FILLER_0_63 ();
 sg13g2_decap_8 FILLER_0_70 ();
 sg13g2_decap_8 FILLER_0_77 ();
 sg13g2_decap_8 FILLER_0_84 ();
 sg13g2_decap_8 FILLER_0_91 ();
 sg13g2_decap_8 FILLER_0_98 ();
 sg13g2_decap_8 FILLER_0_105 ();
 sg13g2_decap_8 FILLER_0_112 ();
 sg13g2_decap_8 FILLER_0_119 ();
 sg13g2_decap_8 FILLER_0_126 ();
 sg13g2_decap_8 FILLER_0_133 ();
 sg13g2_decap_8 FILLER_0_140 ();
 sg13g2_decap_8 FILLER_0_147 ();
 sg13g2_decap_8 FILLER_0_154 ();
 sg13g2_decap_8 FILLER_0_161 ();
 sg13g2_decap_8 FILLER_0_168 ();
 sg13g2_decap_8 FILLER_0_175 ();
 sg13g2_decap_8 FILLER_0_182 ();
 sg13g2_decap_8 FILLER_0_189 ();
 sg13g2_decap_8 FILLER_0_196 ();
 sg13g2_decap_8 FILLER_0_203 ();
 sg13g2_decap_8 FILLER_0_210 ();
 sg13g2_decap_8 FILLER_0_217 ();
 sg13g2_decap_8 FILLER_0_224 ();
 sg13g2_decap_8 FILLER_0_231 ();
 sg13g2_decap_8 FILLER_0_238 ();
 sg13g2_decap_8 FILLER_0_245 ();
 sg13g2_decap_8 FILLER_0_252 ();
 sg13g2_decap_8 FILLER_0_259 ();
 sg13g2_decap_8 FILLER_0_266 ();
 sg13g2_decap_8 FILLER_0_273 ();
 sg13g2_decap_8 FILLER_0_280 ();
 sg13g2_decap_8 FILLER_0_287 ();
 sg13g2_decap_8 FILLER_0_294 ();
 sg13g2_decap_8 FILLER_0_301 ();
 sg13g2_decap_8 FILLER_0_308 ();
 sg13g2_decap_8 FILLER_0_315 ();
 sg13g2_decap_8 FILLER_0_322 ();
 sg13g2_decap_8 FILLER_0_329 ();
 sg13g2_decap_8 FILLER_0_336 ();
 sg13g2_decap_8 FILLER_0_343 ();
 sg13g2_decap_8 FILLER_0_350 ();
 sg13g2_decap_8 FILLER_0_357 ();
 sg13g2_decap_8 FILLER_0_364 ();
 sg13g2_decap_8 FILLER_0_371 ();
 sg13g2_decap_8 FILLER_0_378 ();
 sg13g2_decap_8 FILLER_0_385 ();
 sg13g2_decap_8 FILLER_0_392 ();
 sg13g2_decap_8 FILLER_0_399 ();
 sg13g2_decap_8 FILLER_0_406 ();
 sg13g2_decap_8 FILLER_0_413 ();
 sg13g2_decap_8 FILLER_0_420 ();
 sg13g2_fill_2 FILLER_0_427 ();
 sg13g2_fill_1 FILLER_0_429 ();
 sg13g2_decap_8 FILLER_1_0 ();
 sg13g2_decap_8 FILLER_1_7 ();
 sg13g2_decap_8 FILLER_1_14 ();
 sg13g2_decap_8 FILLER_1_21 ();
 sg13g2_decap_8 FILLER_1_28 ();
 sg13g2_decap_8 FILLER_1_35 ();
 sg13g2_decap_8 FILLER_1_42 ();
 sg13g2_decap_8 FILLER_1_49 ();
 sg13g2_decap_8 FILLER_1_56 ();
 sg13g2_decap_8 FILLER_1_63 ();
 sg13g2_decap_8 FILLER_1_70 ();
 sg13g2_decap_8 FILLER_1_77 ();
 sg13g2_decap_8 FILLER_1_84 ();
 sg13g2_decap_8 FILLER_1_91 ();
 sg13g2_decap_8 FILLER_1_98 ();
 sg13g2_decap_8 FILLER_1_105 ();
 sg13g2_decap_8 FILLER_1_112 ();
 sg13g2_decap_8 FILLER_1_119 ();
 sg13g2_decap_8 FILLER_1_126 ();
 sg13g2_decap_8 FILLER_1_133 ();
 sg13g2_decap_8 FILLER_1_140 ();
 sg13g2_decap_8 FILLER_1_147 ();
 sg13g2_decap_8 FILLER_1_154 ();
 sg13g2_decap_8 FILLER_1_161 ();
 sg13g2_decap_8 FILLER_1_168 ();
 sg13g2_decap_8 FILLER_1_175 ();
 sg13g2_decap_8 FILLER_1_182 ();
 sg13g2_decap_8 FILLER_1_189 ();
 sg13g2_decap_8 FILLER_1_196 ();
 sg13g2_decap_8 FILLER_1_203 ();
 sg13g2_decap_8 FILLER_1_210 ();
 sg13g2_decap_8 FILLER_1_217 ();
 sg13g2_decap_8 FILLER_1_224 ();
 sg13g2_decap_8 FILLER_1_231 ();
 sg13g2_decap_8 FILLER_1_238 ();
 sg13g2_decap_8 FILLER_1_245 ();
 sg13g2_decap_8 FILLER_1_252 ();
 sg13g2_decap_8 FILLER_1_259 ();
 sg13g2_decap_8 FILLER_1_266 ();
 sg13g2_decap_8 FILLER_1_273 ();
 sg13g2_decap_8 FILLER_1_280 ();
 sg13g2_decap_8 FILLER_1_287 ();
 sg13g2_decap_8 FILLER_1_294 ();
 sg13g2_decap_8 FILLER_1_301 ();
 sg13g2_decap_8 FILLER_1_308 ();
 sg13g2_decap_8 FILLER_1_315 ();
 sg13g2_decap_8 FILLER_1_322 ();
 sg13g2_decap_8 FILLER_1_329 ();
 sg13g2_decap_8 FILLER_1_336 ();
 sg13g2_decap_8 FILLER_1_343 ();
 sg13g2_decap_8 FILLER_1_350 ();
 sg13g2_decap_8 FILLER_1_357 ();
 sg13g2_decap_8 FILLER_1_364 ();
 sg13g2_decap_8 FILLER_1_371 ();
 sg13g2_decap_8 FILLER_1_378 ();
 sg13g2_decap_8 FILLER_1_385 ();
 sg13g2_decap_8 FILLER_1_392 ();
 sg13g2_decap_8 FILLER_1_399 ();
 sg13g2_decap_8 FILLER_1_406 ();
 sg13g2_decap_8 FILLER_1_413 ();
 sg13g2_decap_8 FILLER_1_420 ();
 sg13g2_fill_2 FILLER_1_427 ();
 sg13g2_fill_1 FILLER_1_429 ();
 sg13g2_decap_8 FILLER_2_0 ();
 sg13g2_decap_8 FILLER_2_7 ();
 sg13g2_decap_8 FILLER_2_14 ();
 sg13g2_decap_8 FILLER_2_21 ();
 sg13g2_decap_8 FILLER_2_28 ();
 sg13g2_decap_8 FILLER_2_35 ();
 sg13g2_decap_8 FILLER_2_42 ();
 sg13g2_decap_8 FILLER_2_49 ();
 sg13g2_decap_8 FILLER_2_56 ();
 sg13g2_decap_8 FILLER_2_63 ();
 sg13g2_decap_8 FILLER_2_70 ();
 sg13g2_decap_8 FILLER_2_77 ();
 sg13g2_decap_8 FILLER_2_84 ();
 sg13g2_decap_8 FILLER_2_91 ();
 sg13g2_decap_8 FILLER_2_98 ();
 sg13g2_decap_8 FILLER_2_105 ();
 sg13g2_decap_8 FILLER_2_112 ();
 sg13g2_decap_8 FILLER_2_119 ();
 sg13g2_decap_8 FILLER_2_126 ();
 sg13g2_decap_8 FILLER_2_133 ();
 sg13g2_decap_8 FILLER_2_140 ();
 sg13g2_decap_8 FILLER_2_147 ();
 sg13g2_decap_8 FILLER_2_154 ();
 sg13g2_decap_8 FILLER_2_161 ();
 sg13g2_decap_8 FILLER_2_168 ();
 sg13g2_decap_8 FILLER_2_175 ();
 sg13g2_decap_8 FILLER_2_182 ();
 sg13g2_decap_8 FILLER_2_189 ();
 sg13g2_decap_8 FILLER_2_196 ();
 sg13g2_decap_8 FILLER_2_203 ();
 sg13g2_decap_8 FILLER_2_210 ();
 sg13g2_decap_8 FILLER_2_217 ();
 sg13g2_decap_8 FILLER_2_224 ();
 sg13g2_decap_8 FILLER_2_231 ();
 sg13g2_decap_8 FILLER_2_238 ();
 sg13g2_decap_8 FILLER_2_245 ();
 sg13g2_decap_8 FILLER_2_252 ();
 sg13g2_decap_8 FILLER_2_259 ();
 sg13g2_decap_8 FILLER_2_266 ();
 sg13g2_decap_8 FILLER_2_273 ();
 sg13g2_decap_8 FILLER_2_280 ();
 sg13g2_decap_8 FILLER_2_287 ();
 sg13g2_decap_8 FILLER_2_294 ();
 sg13g2_decap_8 FILLER_2_301 ();
 sg13g2_decap_8 FILLER_2_308 ();
 sg13g2_decap_8 FILLER_2_315 ();
 sg13g2_decap_8 FILLER_2_322 ();
 sg13g2_decap_8 FILLER_2_329 ();
 sg13g2_decap_8 FILLER_2_336 ();
 sg13g2_decap_8 FILLER_2_343 ();
 sg13g2_decap_8 FILLER_2_350 ();
 sg13g2_decap_8 FILLER_2_357 ();
 sg13g2_decap_8 FILLER_2_364 ();
 sg13g2_decap_8 FILLER_2_371 ();
 sg13g2_decap_8 FILLER_2_378 ();
 sg13g2_decap_8 FILLER_2_385 ();
 sg13g2_decap_8 FILLER_2_392 ();
 sg13g2_decap_8 FILLER_2_399 ();
 sg13g2_decap_8 FILLER_2_406 ();
 sg13g2_decap_8 FILLER_2_413 ();
 sg13g2_decap_8 FILLER_2_420 ();
 sg13g2_fill_2 FILLER_2_427 ();
 sg13g2_fill_1 FILLER_2_429 ();
 sg13g2_decap_8 FILLER_3_0 ();
 sg13g2_decap_8 FILLER_3_7 ();
 sg13g2_decap_8 FILLER_3_14 ();
 sg13g2_decap_8 FILLER_3_21 ();
 sg13g2_decap_8 FILLER_3_28 ();
 sg13g2_decap_4 FILLER_3_35 ();
 sg13g2_decap_8 FILLER_3_70 ();
 sg13g2_decap_4 FILLER_3_77 ();
 sg13g2_decap_8 FILLER_3_86 ();
 sg13g2_decap_8 FILLER_3_93 ();
 sg13g2_decap_4 FILLER_3_100 ();
 sg13g2_fill_2 FILLER_3_104 ();
 sg13g2_decap_8 FILLER_3_111 ();
 sg13g2_decap_8 FILLER_3_122 ();
 sg13g2_decap_4 FILLER_3_129 ();
 sg13g2_fill_1 FILLER_3_133 ();
 sg13g2_decap_4 FILLER_3_139 ();
 sg13g2_fill_1 FILLER_3_143 ();
 sg13g2_decap_8 FILLER_3_148 ();
 sg13g2_decap_8 FILLER_3_155 ();
 sg13g2_decap_8 FILLER_3_162 ();
 sg13g2_decap_8 FILLER_3_169 ();
 sg13g2_decap_8 FILLER_3_176 ();
 sg13g2_decap_8 FILLER_3_183 ();
 sg13g2_decap_8 FILLER_3_190 ();
 sg13g2_decap_8 FILLER_3_197 ();
 sg13g2_decap_8 FILLER_3_204 ();
 sg13g2_decap_8 FILLER_3_211 ();
 sg13g2_decap_8 FILLER_3_218 ();
 sg13g2_decap_8 FILLER_3_225 ();
 sg13g2_decap_8 FILLER_3_232 ();
 sg13g2_decap_8 FILLER_3_239 ();
 sg13g2_decap_8 FILLER_3_246 ();
 sg13g2_decap_8 FILLER_3_253 ();
 sg13g2_decap_8 FILLER_3_260 ();
 sg13g2_decap_8 FILLER_3_267 ();
 sg13g2_decap_8 FILLER_3_274 ();
 sg13g2_decap_8 FILLER_3_281 ();
 sg13g2_decap_8 FILLER_3_288 ();
 sg13g2_decap_8 FILLER_3_295 ();
 sg13g2_decap_8 FILLER_3_302 ();
 sg13g2_decap_8 FILLER_3_309 ();
 sg13g2_decap_8 FILLER_3_316 ();
 sg13g2_decap_8 FILLER_3_323 ();
 sg13g2_decap_8 FILLER_3_330 ();
 sg13g2_decap_8 FILLER_3_337 ();
 sg13g2_decap_8 FILLER_3_344 ();
 sg13g2_decap_8 FILLER_3_351 ();
 sg13g2_decap_8 FILLER_3_358 ();
 sg13g2_decap_8 FILLER_3_365 ();
 sg13g2_decap_8 FILLER_3_372 ();
 sg13g2_decap_8 FILLER_3_379 ();
 sg13g2_decap_8 FILLER_3_386 ();
 sg13g2_decap_8 FILLER_3_393 ();
 sg13g2_decap_8 FILLER_3_400 ();
 sg13g2_decap_8 FILLER_3_407 ();
 sg13g2_decap_8 FILLER_3_414 ();
 sg13g2_decap_8 FILLER_3_421 ();
 sg13g2_fill_2 FILLER_3_428 ();
 sg13g2_decap_8 FILLER_4_0 ();
 sg13g2_decap_8 FILLER_4_7 ();
 sg13g2_fill_2 FILLER_4_14 ();
 sg13g2_fill_1 FILLER_4_16 ();
 sg13g2_decap_4 FILLER_4_48 ();
 sg13g2_fill_1 FILLER_4_52 ();
 sg13g2_fill_2 FILLER_4_57 ();
 sg13g2_decap_4 FILLER_4_163 ();
 sg13g2_decap_8 FILLER_4_171 ();
 sg13g2_decap_8 FILLER_4_209 ();
 sg13g2_decap_4 FILLER_4_216 ();
 sg13g2_fill_1 FILLER_4_220 ();
 sg13g2_decap_8 FILLER_4_226 ();
 sg13g2_decap_8 FILLER_4_233 ();
 sg13g2_decap_8 FILLER_4_240 ();
 sg13g2_decap_8 FILLER_4_247 ();
 sg13g2_decap_8 FILLER_4_254 ();
 sg13g2_decap_8 FILLER_4_261 ();
 sg13g2_decap_8 FILLER_4_268 ();
 sg13g2_decap_8 FILLER_4_275 ();
 sg13g2_decap_8 FILLER_4_282 ();
 sg13g2_decap_8 FILLER_4_289 ();
 sg13g2_decap_8 FILLER_4_296 ();
 sg13g2_decap_8 FILLER_4_303 ();
 sg13g2_decap_8 FILLER_4_310 ();
 sg13g2_decap_8 FILLER_4_317 ();
 sg13g2_decap_8 FILLER_4_324 ();
 sg13g2_decap_8 FILLER_4_331 ();
 sg13g2_decap_8 FILLER_4_338 ();
 sg13g2_decap_8 FILLER_4_345 ();
 sg13g2_decap_8 FILLER_4_352 ();
 sg13g2_decap_8 FILLER_4_359 ();
 sg13g2_decap_8 FILLER_4_366 ();
 sg13g2_decap_8 FILLER_4_373 ();
 sg13g2_decap_8 FILLER_4_380 ();
 sg13g2_decap_8 FILLER_4_387 ();
 sg13g2_decap_8 FILLER_4_394 ();
 sg13g2_decap_8 FILLER_4_401 ();
 sg13g2_decap_8 FILLER_4_408 ();
 sg13g2_decap_8 FILLER_4_415 ();
 sg13g2_decap_8 FILLER_4_422 ();
 sg13g2_fill_1 FILLER_4_429 ();
 sg13g2_fill_2 FILLER_5_0 ();
 sg13g2_fill_1 FILLER_5_2 ();
 sg13g2_decap_8 FILLER_5_33 ();
 sg13g2_decap_8 FILLER_5_40 ();
 sg13g2_decap_8 FILLER_5_47 ();
 sg13g2_decap_4 FILLER_5_54 ();
 sg13g2_fill_2 FILLER_5_58 ();
 sg13g2_fill_2 FILLER_5_65 ();
 sg13g2_fill_1 FILLER_5_67 ();
 sg13g2_decap_8 FILLER_5_72 ();
 sg13g2_decap_8 FILLER_5_79 ();
 sg13g2_decap_8 FILLER_5_86 ();
 sg13g2_decap_8 FILLER_5_97 ();
 sg13g2_decap_8 FILLER_5_104 ();
 sg13g2_decap_8 FILLER_5_111 ();
 sg13g2_decap_8 FILLER_5_118 ();
 sg13g2_decap_4 FILLER_5_125 ();
 sg13g2_fill_2 FILLER_5_129 ();
 sg13g2_decap_8 FILLER_5_135 ();
 sg13g2_decap_8 FILLER_5_142 ();
 sg13g2_decap_8 FILLER_5_149 ();
 sg13g2_decap_4 FILLER_5_156 ();
 sg13g2_decap_4 FILLER_5_186 ();
 sg13g2_fill_1 FILLER_5_190 ();
 sg13g2_decap_4 FILLER_5_195 ();
 sg13g2_decap_8 FILLER_5_251 ();
 sg13g2_decap_8 FILLER_5_258 ();
 sg13g2_decap_8 FILLER_5_265 ();
 sg13g2_decap_8 FILLER_5_272 ();
 sg13g2_decap_8 FILLER_5_279 ();
 sg13g2_decap_8 FILLER_5_286 ();
 sg13g2_decap_8 FILLER_5_293 ();
 sg13g2_decap_8 FILLER_5_300 ();
 sg13g2_decap_8 FILLER_5_307 ();
 sg13g2_decap_8 FILLER_5_314 ();
 sg13g2_decap_8 FILLER_5_321 ();
 sg13g2_decap_8 FILLER_5_328 ();
 sg13g2_decap_8 FILLER_5_335 ();
 sg13g2_decap_8 FILLER_5_342 ();
 sg13g2_decap_8 FILLER_5_349 ();
 sg13g2_decap_8 FILLER_5_356 ();
 sg13g2_decap_8 FILLER_5_363 ();
 sg13g2_decap_8 FILLER_5_370 ();
 sg13g2_decap_8 FILLER_5_377 ();
 sg13g2_decap_8 FILLER_5_384 ();
 sg13g2_decap_8 FILLER_5_391 ();
 sg13g2_decap_8 FILLER_5_398 ();
 sg13g2_decap_8 FILLER_5_405 ();
 sg13g2_decap_8 FILLER_5_412 ();
 sg13g2_decap_8 FILLER_5_419 ();
 sg13g2_decap_4 FILLER_5_426 ();
 sg13g2_decap_8 FILLER_6_0 ();
 sg13g2_decap_4 FILLER_6_7 ();
 sg13g2_fill_1 FILLER_6_11 ();
 sg13g2_fill_1 FILLER_6_20 ();
 sg13g2_decap_8 FILLER_6_26 ();
 sg13g2_fill_2 FILLER_6_33 ();
 sg13g2_fill_1 FILLER_6_35 ();
 sg13g2_fill_2 FILLER_6_45 ();
 sg13g2_decap_8 FILLER_6_71 ();
 sg13g2_fill_1 FILLER_6_117 ();
 sg13g2_fill_1 FILLER_6_122 ();
 sg13g2_fill_1 FILLER_6_149 ();
 sg13g2_fill_2 FILLER_6_155 ();
 sg13g2_decap_8 FILLER_6_170 ();
 sg13g2_decap_8 FILLER_6_177 ();
 sg13g2_decap_8 FILLER_6_184 ();
 sg13g2_decap_8 FILLER_6_191 ();
 sg13g2_decap_4 FILLER_6_198 ();
 sg13g2_fill_1 FILLER_6_202 ();
 sg13g2_decap_8 FILLER_6_212 ();
 sg13g2_decap_8 FILLER_6_219 ();
 sg13g2_decap_8 FILLER_6_226 ();
 sg13g2_fill_1 FILLER_6_233 ();
 sg13g2_fill_2 FILLER_6_238 ();
 sg13g2_fill_1 FILLER_6_240 ();
 sg13g2_decap_8 FILLER_6_245 ();
 sg13g2_decap_8 FILLER_6_252 ();
 sg13g2_decap_8 FILLER_6_259 ();
 sg13g2_decap_8 FILLER_6_271 ();
 sg13g2_decap_4 FILLER_6_278 ();
 sg13g2_decap_8 FILLER_6_287 ();
 sg13g2_decap_8 FILLER_6_294 ();
 sg13g2_decap_8 FILLER_6_301 ();
 sg13g2_decap_8 FILLER_6_308 ();
 sg13g2_decap_8 FILLER_6_315 ();
 sg13g2_decap_8 FILLER_6_322 ();
 sg13g2_decap_8 FILLER_6_329 ();
 sg13g2_decap_8 FILLER_6_336 ();
 sg13g2_decap_8 FILLER_6_343 ();
 sg13g2_decap_8 FILLER_6_350 ();
 sg13g2_decap_8 FILLER_6_357 ();
 sg13g2_decap_8 FILLER_6_364 ();
 sg13g2_decap_8 FILLER_6_371 ();
 sg13g2_decap_8 FILLER_6_378 ();
 sg13g2_decap_8 FILLER_6_385 ();
 sg13g2_decap_8 FILLER_6_392 ();
 sg13g2_decap_8 FILLER_6_399 ();
 sg13g2_decap_8 FILLER_6_406 ();
 sg13g2_decap_8 FILLER_6_413 ();
 sg13g2_decap_8 FILLER_6_420 ();
 sg13g2_fill_2 FILLER_6_427 ();
 sg13g2_fill_1 FILLER_6_429 ();
 sg13g2_decap_8 FILLER_7_0 ();
 sg13g2_fill_1 FILLER_7_7 ();
 sg13g2_decap_4 FILLER_7_60 ();
 sg13g2_fill_1 FILLER_7_64 ();
 sg13g2_decap_8 FILLER_7_70 ();
 sg13g2_fill_1 FILLER_7_77 ();
 sg13g2_decap_8 FILLER_7_90 ();
 sg13g2_decap_8 FILLER_7_97 ();
 sg13g2_fill_1 FILLER_7_104 ();
 sg13g2_decap_4 FILLER_7_140 ();
 sg13g2_fill_1 FILLER_7_144 ();
 sg13g2_decap_8 FILLER_7_149 ();
 sg13g2_fill_1 FILLER_7_156 ();
 sg13g2_decap_4 FILLER_7_165 ();
 sg13g2_fill_2 FILLER_7_173 ();
 sg13g2_decap_8 FILLER_7_201 ();
 sg13g2_decap_8 FILLER_7_208 ();
 sg13g2_fill_1 FILLER_7_215 ();
 sg13g2_decap_8 FILLER_7_220 ();
 sg13g2_fill_2 FILLER_7_227 ();
 sg13g2_fill_1 FILLER_7_234 ();
 sg13g2_fill_1 FILLER_7_261 ();
 sg13g2_fill_1 FILLER_7_288 ();
 sg13g2_fill_1 FILLER_7_297 ();
 sg13g2_decap_8 FILLER_7_306 ();
 sg13g2_decap_8 FILLER_7_313 ();
 sg13g2_decap_8 FILLER_7_320 ();
 sg13g2_decap_8 FILLER_7_327 ();
 sg13g2_fill_1 FILLER_7_334 ();
 sg13g2_decap_8 FILLER_7_361 ();
 sg13g2_decap_8 FILLER_7_368 ();
 sg13g2_decap_8 FILLER_7_375 ();
 sg13g2_decap_8 FILLER_7_382 ();
 sg13g2_decap_8 FILLER_7_389 ();
 sg13g2_decap_8 FILLER_7_396 ();
 sg13g2_decap_8 FILLER_7_403 ();
 sg13g2_decap_8 FILLER_7_410 ();
 sg13g2_decap_8 FILLER_7_417 ();
 sg13g2_decap_4 FILLER_7_424 ();
 sg13g2_fill_2 FILLER_7_428 ();
 sg13g2_decap_8 FILLER_8_0 ();
 sg13g2_fill_1 FILLER_8_7 ();
 sg13g2_decap_4 FILLER_8_38 ();
 sg13g2_decap_4 FILLER_8_46 ();
 sg13g2_fill_1 FILLER_8_58 ();
 sg13g2_fill_1 FILLER_8_67 ();
 sg13g2_fill_1 FILLER_8_77 ();
 sg13g2_decap_8 FILLER_8_112 ();
 sg13g2_fill_2 FILLER_8_119 ();
 sg13g2_fill_1 FILLER_8_121 ();
 sg13g2_decap_4 FILLER_8_177 ();
 sg13g2_fill_1 FILLER_8_181 ();
 sg13g2_decap_8 FILLER_8_186 ();
 sg13g2_fill_2 FILLER_8_207 ();
 sg13g2_decap_8 FILLER_8_247 ();
 sg13g2_decap_8 FILLER_8_254 ();
 sg13g2_decap_8 FILLER_8_261 ();
 sg13g2_fill_1 FILLER_8_268 ();
 sg13g2_decap_4 FILLER_8_273 ();
 sg13g2_fill_2 FILLER_8_277 ();
 sg13g2_decap_4 FILLER_8_302 ();
 sg13g2_decap_8 FILLER_8_311 ();
 sg13g2_fill_2 FILLER_8_318 ();
 sg13g2_fill_1 FILLER_8_328 ();
 sg13g2_decap_4 FILLER_8_337 ();
 sg13g2_decap_8 FILLER_8_345 ();
 sg13g2_decap_8 FILLER_8_357 ();
 sg13g2_decap_8 FILLER_8_364 ();
 sg13g2_decap_8 FILLER_8_371 ();
 sg13g2_decap_8 FILLER_8_378 ();
 sg13g2_decap_8 FILLER_8_385 ();
 sg13g2_decap_8 FILLER_8_392 ();
 sg13g2_decap_8 FILLER_8_399 ();
 sg13g2_decap_8 FILLER_8_406 ();
 sg13g2_decap_8 FILLER_8_413 ();
 sg13g2_decap_8 FILLER_8_420 ();
 sg13g2_fill_2 FILLER_8_427 ();
 sg13g2_fill_1 FILLER_8_429 ();
 sg13g2_decap_8 FILLER_9_0 ();
 sg13g2_decap_4 FILLER_9_7 ();
 sg13g2_fill_1 FILLER_9_11 ();
 sg13g2_decap_8 FILLER_9_20 ();
 sg13g2_decap_8 FILLER_9_27 ();
 sg13g2_decap_8 FILLER_9_34 ();
 sg13g2_decap_8 FILLER_9_41 ();
 sg13g2_decap_4 FILLER_9_48 ();
 sg13g2_fill_1 FILLER_9_52 ();
 sg13g2_fill_2 FILLER_9_58 ();
 sg13g2_fill_1 FILLER_9_60 ();
 sg13g2_decap_8 FILLER_9_73 ();
 sg13g2_decap_4 FILLER_9_80 ();
 sg13g2_decap_4 FILLER_9_88 ();
 sg13g2_decap_8 FILLER_9_96 ();
 sg13g2_decap_8 FILLER_9_103 ();
 sg13g2_fill_2 FILLER_9_110 ();
 sg13g2_fill_1 FILLER_9_112 ();
 sg13g2_fill_1 FILLER_9_128 ();
 sg13g2_decap_8 FILLER_9_139 ();
 sg13g2_fill_2 FILLER_9_146 ();
 sg13g2_fill_1 FILLER_9_148 ();
 sg13g2_decap_4 FILLER_9_153 ();
 sg13g2_decap_8 FILLER_9_161 ();
 sg13g2_fill_2 FILLER_9_168 ();
 sg13g2_fill_1 FILLER_9_170 ();
 sg13g2_fill_2 FILLER_9_176 ();
 sg13g2_fill_2 FILLER_9_208 ();
 sg13g2_decap_8 FILLER_9_222 ();
 sg13g2_fill_2 FILLER_9_229 ();
 sg13g2_fill_1 FILLER_9_261 ();
 sg13g2_fill_2 FILLER_9_275 ();
 sg13g2_fill_1 FILLER_9_277 ();
 sg13g2_decap_8 FILLER_9_283 ();
 sg13g2_decap_8 FILLER_9_290 ();
 sg13g2_fill_1 FILLER_9_297 ();
 sg13g2_fill_1 FILLER_9_304 ();
 sg13g2_fill_2 FILLER_9_322 ();
 sg13g2_fill_2 FILLER_9_335 ();
 sg13g2_fill_1 FILLER_9_337 ();
 sg13g2_decap_8 FILLER_9_358 ();
 sg13g2_decap_8 FILLER_9_365 ();
 sg13g2_decap_8 FILLER_9_372 ();
 sg13g2_decap_8 FILLER_9_379 ();
 sg13g2_decap_8 FILLER_9_386 ();
 sg13g2_decap_8 FILLER_9_393 ();
 sg13g2_decap_8 FILLER_9_400 ();
 sg13g2_decap_8 FILLER_9_407 ();
 sg13g2_decap_8 FILLER_9_414 ();
 sg13g2_decap_8 FILLER_9_421 ();
 sg13g2_fill_2 FILLER_9_428 ();
 sg13g2_decap_4 FILLER_10_0 ();
 sg13g2_fill_2 FILLER_10_4 ();
 sg13g2_fill_2 FILLER_10_32 ();
 sg13g2_fill_1 FILLER_10_34 ();
 sg13g2_decap_8 FILLER_10_39 ();
 sg13g2_decap_8 FILLER_10_58 ();
 sg13g2_fill_1 FILLER_10_65 ();
 sg13g2_fill_1 FILLER_10_71 ();
 sg13g2_decap_8 FILLER_10_98 ();
 sg13g2_fill_2 FILLER_10_105 ();
 sg13g2_fill_2 FILLER_10_140 ();
 sg13g2_decap_8 FILLER_10_146 ();
 sg13g2_fill_2 FILLER_10_153 ();
 sg13g2_fill_1 FILLER_10_155 ();
 sg13g2_decap_8 FILLER_10_161 ();
 sg13g2_fill_1 FILLER_10_168 ();
 sg13g2_fill_2 FILLER_10_178 ();
 sg13g2_fill_1 FILLER_10_180 ();
 sg13g2_decap_4 FILLER_10_199 ();
 sg13g2_decap_8 FILLER_10_246 ();
 sg13g2_decap_4 FILLER_10_253 ();
 sg13g2_fill_1 FILLER_10_257 ();
 sg13g2_fill_1 FILLER_10_262 ();
 sg13g2_fill_1 FILLER_10_267 ();
 sg13g2_fill_2 FILLER_10_285 ();
 sg13g2_fill_1 FILLER_10_293 ();
 sg13g2_fill_2 FILLER_10_315 ();
 sg13g2_decap_8 FILLER_10_322 ();
 sg13g2_fill_2 FILLER_10_337 ();
 sg13g2_fill_2 FILLER_10_343 ();
 sg13g2_fill_1 FILLER_10_345 ();
 sg13g2_fill_1 FILLER_10_352 ();
 sg13g2_fill_2 FILLER_10_357 ();
 sg13g2_fill_1 FILLER_10_359 ();
 sg13g2_decap_8 FILLER_10_390 ();
 sg13g2_decap_8 FILLER_10_397 ();
 sg13g2_decap_8 FILLER_10_404 ();
 sg13g2_decap_8 FILLER_10_411 ();
 sg13g2_decap_8 FILLER_10_418 ();
 sg13g2_decap_4 FILLER_10_425 ();
 sg13g2_fill_1 FILLER_10_429 ();
 sg13g2_decap_8 FILLER_11_0 ();
 sg13g2_fill_1 FILLER_11_7 ();
 sg13g2_fill_1 FILLER_11_29 ();
 sg13g2_decap_4 FILLER_11_57 ();
 sg13g2_decap_8 FILLER_11_65 ();
 sg13g2_decap_8 FILLER_11_72 ();
 sg13g2_fill_2 FILLER_11_79 ();
 sg13g2_fill_2 FILLER_11_85 ();
 sg13g2_fill_1 FILLER_11_91 ();
 sg13g2_fill_1 FILLER_11_96 ();
 sg13g2_fill_1 FILLER_11_101 ();
 sg13g2_fill_1 FILLER_11_111 ();
 sg13g2_decap_4 FILLER_11_124 ();
 sg13g2_fill_1 FILLER_11_128 ();
 sg13g2_decap_4 FILLER_11_143 ();
 sg13g2_fill_1 FILLER_11_147 ();
 sg13g2_decap_8 FILLER_11_163 ();
 sg13g2_decap_8 FILLER_11_176 ();
 sg13g2_decap_4 FILLER_11_183 ();
 sg13g2_fill_2 FILLER_11_187 ();
 sg13g2_decap_8 FILLER_11_218 ();
 sg13g2_decap_8 FILLER_11_225 ();
 sg13g2_decap_8 FILLER_11_232 ();
 sg13g2_fill_2 FILLER_11_252 ();
 sg13g2_fill_2 FILLER_11_257 ();
 sg13g2_fill_2 FILLER_11_263 ();
 sg13g2_fill_1 FILLER_11_265 ();
 sg13g2_fill_2 FILLER_11_270 ();
 sg13g2_fill_1 FILLER_11_272 ();
 sg13g2_fill_2 FILLER_11_278 ();
 sg13g2_fill_2 FILLER_11_299 ();
 sg13g2_fill_1 FILLER_11_305 ();
 sg13g2_fill_1 FILLER_11_311 ();
 sg13g2_fill_1 FILLER_11_317 ();
 sg13g2_fill_1 FILLER_11_323 ();
 sg13g2_fill_1 FILLER_11_328 ();
 sg13g2_decap_4 FILLER_11_337 ();
 sg13g2_decap_8 FILLER_11_368 ();
 sg13g2_decap_4 FILLER_11_375 ();
 sg13g2_fill_1 FILLER_11_379 ();
 sg13g2_decap_8 FILLER_11_384 ();
 sg13g2_decap_8 FILLER_11_391 ();
 sg13g2_decap_8 FILLER_11_398 ();
 sg13g2_decap_8 FILLER_11_405 ();
 sg13g2_decap_8 FILLER_11_412 ();
 sg13g2_decap_8 FILLER_11_419 ();
 sg13g2_decap_4 FILLER_11_426 ();
 sg13g2_fill_2 FILLER_12_0 ();
 sg13g2_fill_1 FILLER_12_28 ();
 sg13g2_fill_2 FILLER_12_37 ();
 sg13g2_fill_2 FILLER_12_42 ();
 sg13g2_fill_2 FILLER_12_52 ();
 sg13g2_fill_2 FILLER_12_85 ();
 sg13g2_fill_2 FILLER_12_95 ();
 sg13g2_fill_1 FILLER_12_97 ();
 sg13g2_fill_2 FILLER_12_122 ();
 sg13g2_decap_8 FILLER_12_132 ();
 sg13g2_decap_4 FILLER_12_139 ();
 sg13g2_fill_1 FILLER_12_143 ();
 sg13g2_decap_8 FILLER_12_180 ();
 sg13g2_decap_4 FILLER_12_187 ();
 sg13g2_decap_8 FILLER_12_226 ();
 sg13g2_decap_4 FILLER_12_233 ();
 sg13g2_fill_1 FILLER_12_237 ();
 sg13g2_fill_2 FILLER_12_286 ();
 sg13g2_decap_8 FILLER_12_301 ();
 sg13g2_decap_8 FILLER_12_308 ();
 sg13g2_fill_2 FILLER_12_315 ();
 sg13g2_fill_1 FILLER_12_317 ();
 sg13g2_fill_2 FILLER_12_327 ();
 sg13g2_fill_1 FILLER_12_329 ();
 sg13g2_fill_1 FILLER_12_339 ();
 sg13g2_decap_8 FILLER_12_344 ();
 sg13g2_fill_2 FILLER_12_356 ();
 sg13g2_decap_4 FILLER_12_389 ();
 sg13g2_decap_8 FILLER_12_397 ();
 sg13g2_decap_8 FILLER_12_404 ();
 sg13g2_decap_8 FILLER_12_411 ();
 sg13g2_decap_8 FILLER_12_418 ();
 sg13g2_decap_4 FILLER_12_425 ();
 sg13g2_fill_1 FILLER_12_429 ();
 sg13g2_decap_8 FILLER_13_0 ();
 sg13g2_decap_4 FILLER_13_7 ();
 sg13g2_fill_2 FILLER_13_15 ();
 sg13g2_fill_1 FILLER_13_17 ();
 sg13g2_fill_2 FILLER_13_26 ();
 sg13g2_fill_1 FILLER_13_28 ();
 sg13g2_decap_8 FILLER_13_33 ();
 sg13g2_decap_8 FILLER_13_40 ();
 sg13g2_decap_8 FILLER_13_47 ();
 sg13g2_decap_8 FILLER_13_54 ();
 sg13g2_fill_1 FILLER_13_61 ();
 sg13g2_fill_1 FILLER_13_75 ();
 sg13g2_decap_4 FILLER_13_85 ();
 sg13g2_fill_1 FILLER_13_89 ();
 sg13g2_fill_2 FILLER_13_93 ();
 sg13g2_fill_1 FILLER_13_95 ();
 sg13g2_decap_4 FILLER_13_101 ();
 sg13g2_fill_1 FILLER_13_105 ();
 sg13g2_decap_8 FILLER_13_116 ();
 sg13g2_decap_4 FILLER_13_123 ();
 sg13g2_fill_1 FILLER_13_139 ();
 sg13g2_decap_8 FILLER_13_162 ();
 sg13g2_fill_1 FILLER_13_169 ();
 sg13g2_decap_8 FILLER_13_175 ();
 sg13g2_decap_8 FILLER_13_182 ();
 sg13g2_fill_1 FILLER_13_189 ();
 sg13g2_fill_1 FILLER_13_195 ();
 sg13g2_fill_1 FILLER_13_201 ();
 sg13g2_fill_1 FILLER_13_206 ();
 sg13g2_decap_4 FILLER_13_211 ();
 sg13g2_fill_2 FILLER_13_215 ();
 sg13g2_decap_4 FILLER_13_248 ();
 sg13g2_decap_4 FILLER_13_256 ();
 sg13g2_fill_1 FILLER_13_260 ();
 sg13g2_decap_4 FILLER_13_265 ();
 sg13g2_decap_8 FILLER_13_273 ();
 sg13g2_decap_8 FILLER_13_280 ();
 sg13g2_fill_1 FILLER_13_287 ();
 sg13g2_decap_4 FILLER_13_293 ();
 sg13g2_fill_2 FILLER_13_297 ();
 sg13g2_fill_1 FILLER_13_303 ();
 sg13g2_fill_1 FILLER_13_309 ();
 sg13g2_fill_1 FILLER_13_314 ();
 sg13g2_fill_1 FILLER_13_319 ();
 sg13g2_fill_2 FILLER_13_332 ();
 sg13g2_fill_1 FILLER_13_334 ();
 sg13g2_decap_8 FILLER_13_340 ();
 sg13g2_decap_4 FILLER_13_347 ();
 sg13g2_decap_8 FILLER_13_355 ();
 sg13g2_decap_4 FILLER_13_362 ();
 sg13g2_fill_1 FILLER_13_366 ();
 sg13g2_decap_8 FILLER_13_371 ();
 sg13g2_decap_8 FILLER_13_378 ();
 sg13g2_decap_8 FILLER_13_385 ();
 sg13g2_decap_8 FILLER_13_392 ();
 sg13g2_decap_8 FILLER_13_399 ();
 sg13g2_decap_8 FILLER_13_406 ();
 sg13g2_decap_8 FILLER_13_413 ();
 sg13g2_decap_8 FILLER_13_420 ();
 sg13g2_fill_2 FILLER_13_427 ();
 sg13g2_fill_1 FILLER_13_429 ();
 sg13g2_decap_8 FILLER_14_0 ();
 sg13g2_decap_4 FILLER_14_7 ();
 sg13g2_fill_2 FILLER_14_11 ();
 sg13g2_decap_4 FILLER_14_17 ();
 sg13g2_decap_8 FILLER_14_47 ();
 sg13g2_fill_2 FILLER_14_54 ();
 sg13g2_fill_1 FILLER_14_56 ();
 sg13g2_fill_1 FILLER_14_87 ();
 sg13g2_fill_1 FILLER_14_101 ();
 sg13g2_decap_4 FILLER_14_110 ();
 sg13g2_decap_8 FILLER_14_117 ();
 sg13g2_fill_2 FILLER_14_124 ();
 sg13g2_decap_8 FILLER_14_131 ();
 sg13g2_fill_1 FILLER_14_138 ();
 sg13g2_decap_8 FILLER_14_144 ();
 sg13g2_decap_8 FILLER_14_151 ();
 sg13g2_fill_2 FILLER_14_206 ();
 sg13g2_fill_2 FILLER_14_219 ();
 sg13g2_fill_1 FILLER_14_221 ();
 sg13g2_fill_1 FILLER_14_231 ();
 sg13g2_fill_2 FILLER_14_240 ();
 sg13g2_decap_4 FILLER_14_246 ();
 sg13g2_fill_2 FILLER_14_296 ();
 sg13g2_fill_1 FILLER_14_308 ();
 sg13g2_fill_2 FILLER_14_318 ();
 sg13g2_fill_1 FILLER_14_320 ();
 sg13g2_fill_2 FILLER_14_326 ();
 sg13g2_decap_8 FILLER_14_332 ();
 sg13g2_fill_2 FILLER_14_339 ();
 sg13g2_fill_2 FILLER_14_346 ();
 sg13g2_fill_2 FILLER_14_356 ();
 sg13g2_fill_1 FILLER_14_358 ();
 sg13g2_fill_2 FILLER_14_389 ();
 sg13g2_fill_1 FILLER_14_391 ();
 sg13g2_decap_8 FILLER_14_397 ();
 sg13g2_decap_8 FILLER_14_404 ();
 sg13g2_decap_8 FILLER_14_411 ();
 sg13g2_decap_8 FILLER_14_418 ();
 sg13g2_decap_4 FILLER_14_425 ();
 sg13g2_fill_1 FILLER_14_429 ();
 sg13g2_fill_2 FILLER_15_0 ();
 sg13g2_decap_8 FILLER_15_28 ();
 sg13g2_decap_4 FILLER_15_35 ();
 sg13g2_fill_2 FILLER_15_39 ();
 sg13g2_fill_1 FILLER_15_65 ();
 sg13g2_fill_2 FILLER_15_76 ();
 sg13g2_fill_1 FILLER_15_78 ();
 sg13g2_fill_2 FILLER_15_104 ();
 sg13g2_fill_1 FILLER_15_106 ();
 sg13g2_decap_4 FILLER_15_142 ();
 sg13g2_decap_4 FILLER_15_150 ();
 sg13g2_fill_1 FILLER_15_154 ();
 sg13g2_decap_8 FILLER_15_175 ();
 sg13g2_decap_4 FILLER_15_182 ();
 sg13g2_fill_2 FILLER_15_186 ();
 sg13g2_fill_2 FILLER_15_206 ();
 sg13g2_decap_8 FILLER_15_222 ();
 sg13g2_decap_4 FILLER_15_229 ();
 sg13g2_decap_4 FILLER_15_242 ();
 sg13g2_fill_1 FILLER_15_246 ();
 sg13g2_decap_4 FILLER_15_257 ();
 sg13g2_decap_4 FILLER_15_275 ();
 sg13g2_fill_1 FILLER_15_283 ();
 sg13g2_decap_8 FILLER_15_294 ();
 sg13g2_fill_2 FILLER_15_301 ();
 sg13g2_fill_1 FILLER_15_303 ();
 sg13g2_decap_8 FILLER_15_308 ();
 sg13g2_fill_1 FILLER_15_324 ();
 sg13g2_fill_1 FILLER_15_336 ();
 sg13g2_fill_1 FILLER_15_366 ();
 sg13g2_fill_1 FILLER_15_371 ();
 sg13g2_fill_2 FILLER_15_382 ();
 sg13g2_fill_1 FILLER_15_384 ();
 sg13g2_decap_8 FILLER_15_390 ();
 sg13g2_decap_8 FILLER_15_397 ();
 sg13g2_decap_8 FILLER_15_404 ();
 sg13g2_decap_8 FILLER_15_411 ();
 sg13g2_decap_8 FILLER_15_418 ();
 sg13g2_decap_4 FILLER_15_425 ();
 sg13g2_fill_1 FILLER_15_429 ();
 sg13g2_decap_8 FILLER_16_0 ();
 sg13g2_fill_1 FILLER_16_15 ();
 sg13g2_decap_8 FILLER_16_23 ();
 sg13g2_decap_8 FILLER_16_30 ();
 sg13g2_decap_4 FILLER_16_47 ();
 sg13g2_fill_1 FILLER_16_59 ();
 sg13g2_fill_1 FILLER_16_68 ();
 sg13g2_decap_8 FILLER_16_91 ();
 sg13g2_decap_8 FILLER_16_98 ();
 sg13g2_decap_8 FILLER_16_105 ();
 sg13g2_decap_8 FILLER_16_112 ();
 sg13g2_decap_8 FILLER_16_119 ();
 sg13g2_decap_8 FILLER_16_126 ();
 sg13g2_fill_2 FILLER_16_133 ();
 sg13g2_fill_1 FILLER_16_135 ();
 sg13g2_decap_4 FILLER_16_141 ();
 sg13g2_fill_2 FILLER_16_153 ();
 sg13g2_fill_1 FILLER_16_155 ();
 sg13g2_fill_2 FILLER_16_160 ();
 sg13g2_decap_8 FILLER_16_168 ();
 sg13g2_decap_8 FILLER_16_175 ();
 sg13g2_decap_4 FILLER_16_182 ();
 sg13g2_fill_1 FILLER_16_196 ();
 sg13g2_decap_4 FILLER_16_201 ();
 sg13g2_fill_2 FILLER_16_205 ();
 sg13g2_fill_2 FILLER_16_219 ();
 sg13g2_fill_1 FILLER_16_221 ();
 sg13g2_fill_2 FILLER_16_227 ();
 sg13g2_fill_1 FILLER_16_229 ();
 sg13g2_fill_2 FILLER_16_256 ();
 sg13g2_fill_1 FILLER_16_258 ();
 sg13g2_fill_1 FILLER_16_265 ();
 sg13g2_decap_4 FILLER_16_276 ();
 sg13g2_fill_2 FILLER_16_299 ();
 sg13g2_decap_8 FILLER_16_306 ();
 sg13g2_decap_4 FILLER_16_313 ();
 sg13g2_fill_1 FILLER_16_343 ();
 sg13g2_decap_4 FILLER_16_351 ();
 sg13g2_fill_1 FILLER_16_355 ();
 sg13g2_fill_1 FILLER_16_370 ();
 sg13g2_fill_1 FILLER_16_376 ();
 sg13g2_fill_1 FILLER_16_382 ();
 sg13g2_fill_2 FILLER_16_388 ();
 sg13g2_fill_1 FILLER_16_398 ();
 sg13g2_decap_8 FILLER_16_407 ();
 sg13g2_decap_8 FILLER_16_414 ();
 sg13g2_decap_8 FILLER_16_421 ();
 sg13g2_fill_2 FILLER_16_428 ();
 sg13g2_fill_2 FILLER_17_8 ();
 sg13g2_fill_1 FILLER_17_10 ();
 sg13g2_decap_4 FILLER_17_24 ();
 sg13g2_fill_2 FILLER_17_28 ();
 sg13g2_decap_8 FILLER_17_45 ();
 sg13g2_decap_4 FILLER_17_52 ();
 sg13g2_decap_8 FILLER_17_69 ();
 sg13g2_fill_2 FILLER_17_80 ();
 sg13g2_fill_1 FILLER_17_82 ();
 sg13g2_fill_2 FILLER_17_88 ();
 sg13g2_fill_2 FILLER_17_98 ();
 sg13g2_decap_4 FILLER_17_112 ();
 sg13g2_fill_1 FILLER_17_116 ();
 sg13g2_decap_4 FILLER_17_125 ();
 sg13g2_fill_1 FILLER_17_129 ();
 sg13g2_fill_1 FILLER_17_143 ();
 sg13g2_fill_2 FILLER_17_149 ();
 sg13g2_decap_4 FILLER_17_169 ();
 sg13g2_fill_2 FILLER_17_173 ();
 sg13g2_fill_1 FILLER_17_180 ();
 sg13g2_fill_2 FILLER_17_189 ();
 sg13g2_decap_8 FILLER_17_217 ();
 sg13g2_fill_1 FILLER_17_224 ();
 sg13g2_fill_2 FILLER_17_229 ();
 sg13g2_decap_4 FILLER_17_236 ();
 sg13g2_fill_1 FILLER_17_240 ();
 sg13g2_decap_8 FILLER_17_255 ();
 sg13g2_decap_8 FILLER_17_262 ();
 sg13g2_decap_4 FILLER_17_269 ();
 sg13g2_fill_1 FILLER_17_273 ();
 sg13g2_decap_4 FILLER_17_306 ();
 sg13g2_fill_1 FILLER_17_310 ();
 sg13g2_fill_2 FILLER_17_317 ();
 sg13g2_fill_1 FILLER_17_319 ();
 sg13g2_fill_2 FILLER_17_350 ();
 sg13g2_fill_1 FILLER_17_352 ();
 sg13g2_decap_8 FILLER_17_358 ();
 sg13g2_fill_2 FILLER_17_365 ();
 sg13g2_fill_1 FILLER_17_367 ();
 sg13g2_fill_2 FILLER_17_387 ();
 sg13g2_fill_1 FILLER_17_389 ();
 sg13g2_decap_4 FILLER_17_398 ();
 sg13g2_fill_1 FILLER_17_402 ();
 sg13g2_decap_8 FILLER_17_407 ();
 sg13g2_decap_8 FILLER_17_414 ();
 sg13g2_decap_8 FILLER_17_421 ();
 sg13g2_fill_2 FILLER_17_428 ();
 sg13g2_decap_8 FILLER_18_0 ();
 sg13g2_fill_2 FILLER_18_7 ();
 sg13g2_fill_2 FILLER_18_39 ();
 sg13g2_decap_8 FILLER_18_53 ();
 sg13g2_fill_1 FILLER_18_60 ();
 sg13g2_fill_2 FILLER_18_75 ();
 sg13g2_fill_1 FILLER_18_77 ();
 sg13g2_fill_2 FILLER_18_98 ();
 sg13g2_fill_1 FILLER_18_100 ();
 sg13g2_fill_2 FILLER_18_119 ();
 sg13g2_fill_1 FILLER_18_121 ();
 sg13g2_fill_2 FILLER_18_127 ();
 sg13g2_decap_4 FILLER_18_143 ();
 sg13g2_fill_2 FILLER_18_152 ();
 sg13g2_decap_8 FILLER_18_158 ();
 sg13g2_decap_4 FILLER_18_165 ();
 sg13g2_fill_1 FILLER_18_169 ();
 sg13g2_fill_2 FILLER_18_178 ();
 sg13g2_fill_1 FILLER_18_184 ();
 sg13g2_fill_1 FILLER_18_189 ();
 sg13g2_fill_2 FILLER_18_194 ();
 sg13g2_fill_2 FILLER_18_200 ();
 sg13g2_decap_4 FILLER_18_206 ();
 sg13g2_decap_4 FILLER_18_218 ();
 sg13g2_fill_2 FILLER_18_222 ();
 sg13g2_fill_2 FILLER_18_246 ();
 sg13g2_decap_8 FILLER_18_254 ();
 sg13g2_decap_8 FILLER_18_276 ();
 sg13g2_decap_4 FILLER_18_292 ();
 sg13g2_fill_1 FILLER_18_296 ();
 sg13g2_fill_1 FILLER_18_302 ();
 sg13g2_decap_4 FILLER_18_317 ();
 sg13g2_fill_1 FILLER_18_326 ();
 sg13g2_fill_2 FILLER_18_332 ();
 sg13g2_fill_2 FILLER_18_344 ();
 sg13g2_decap_8 FILLER_18_351 ();
 sg13g2_fill_2 FILLER_18_358 ();
 sg13g2_decap_8 FILLER_18_365 ();
 sg13g2_fill_1 FILLER_18_372 ();
 sg13g2_decap_4 FILLER_18_388 ();
 sg13g2_fill_2 FILLER_18_400 ();
 sg13g2_decap_4 FILLER_18_406 ();
 sg13g2_fill_1 FILLER_18_410 ();
 sg13g2_decap_8 FILLER_18_415 ();
 sg13g2_decap_8 FILLER_18_422 ();
 sg13g2_fill_1 FILLER_18_429 ();
 sg13g2_decap_8 FILLER_19_0 ();
 sg13g2_fill_1 FILLER_19_7 ();
 sg13g2_decap_8 FILLER_19_24 ();
 sg13g2_fill_2 FILLER_19_31 ();
 sg13g2_decap_8 FILLER_19_38 ();
 sg13g2_decap_4 FILLER_19_45 ();
 sg13g2_decap_4 FILLER_19_53 ();
 sg13g2_decap_8 FILLER_19_62 ();
 sg13g2_decap_8 FILLER_19_69 ();
 sg13g2_fill_2 FILLER_19_76 ();
 sg13g2_fill_1 FILLER_19_78 ();
 sg13g2_fill_1 FILLER_19_87 ();
 sg13g2_fill_1 FILLER_19_95 ();
 sg13g2_fill_2 FILLER_19_140 ();
 sg13g2_fill_1 FILLER_19_142 ();
 sg13g2_fill_2 FILLER_19_169 ();
 sg13g2_fill_1 FILLER_19_171 ();
 sg13g2_decap_4 FILLER_19_178 ();
 sg13g2_decap_8 FILLER_19_198 ();
 sg13g2_decap_8 FILLER_19_205 ();
 sg13g2_decap_8 FILLER_19_216 ();
 sg13g2_fill_2 FILLER_19_223 ();
 sg13g2_fill_1 FILLER_19_225 ();
 sg13g2_fill_2 FILLER_19_231 ();
 sg13g2_fill_1 FILLER_19_238 ();
 sg13g2_fill_1 FILLER_19_256 ();
 sg13g2_decap_4 FILLER_19_267 ();
 sg13g2_fill_2 FILLER_19_271 ();
 sg13g2_fill_2 FILLER_19_280 ();
 sg13g2_fill_1 FILLER_19_288 ();
 sg13g2_decap_4 FILLER_19_293 ();
 sg13g2_fill_1 FILLER_19_297 ();
 sg13g2_decap_8 FILLER_19_303 ();
 sg13g2_decap_8 FILLER_19_310 ();
 sg13g2_decap_8 FILLER_19_330 ();
 sg13g2_decap_8 FILLER_19_337 ();
 sg13g2_fill_1 FILLER_19_344 ();
 sg13g2_decap_4 FILLER_19_363 ();
 sg13g2_decap_4 FILLER_19_372 ();
 sg13g2_fill_1 FILLER_19_392 ();
 sg13g2_fill_1 FILLER_20_0 ();
 sg13g2_fill_2 FILLER_20_14 ();
 sg13g2_fill_2 FILLER_20_46 ();
 sg13g2_decap_8 FILLER_20_58 ();
 sg13g2_fill_1 FILLER_20_65 ();
 sg13g2_decap_4 FILLER_20_74 ();
 sg13g2_fill_1 FILLER_20_78 ();
 sg13g2_decap_4 FILLER_20_114 ();
 sg13g2_decap_8 FILLER_20_130 ();
 sg13g2_decap_8 FILLER_20_137 ();
 sg13g2_decap_4 FILLER_20_144 ();
 sg13g2_fill_1 FILLER_20_148 ();
 sg13g2_fill_1 FILLER_20_158 ();
 sg13g2_decap_4 FILLER_20_163 ();
 sg13g2_decap_4 FILLER_20_179 ();
 sg13g2_fill_2 FILLER_20_183 ();
 sg13g2_decap_4 FILLER_20_211 ();
 sg13g2_decap_8 FILLER_20_220 ();
 sg13g2_fill_1 FILLER_20_227 ();
 sg13g2_fill_1 FILLER_20_233 ();
 sg13g2_fill_2 FILLER_20_242 ();
 sg13g2_decap_4 FILLER_20_248 ();
 sg13g2_fill_1 FILLER_20_284 ();
 sg13g2_decap_8 FILLER_20_300 ();
 sg13g2_fill_2 FILLER_20_307 ();
 sg13g2_decap_4 FILLER_20_313 ();
 sg13g2_decap_8 FILLER_20_356 ();
 sg13g2_decap_8 FILLER_20_363 ();
 sg13g2_decap_4 FILLER_20_370 ();
 sg13g2_fill_2 FILLER_20_374 ();
 sg13g2_decap_4 FILLER_20_387 ();
 sg13g2_fill_1 FILLER_20_391 ();
 sg13g2_fill_2 FILLER_20_405 ();
 sg13g2_decap_8 FILLER_20_412 ();
 sg13g2_decap_8 FILLER_20_419 ();
 sg13g2_decap_4 FILLER_20_426 ();
 sg13g2_decap_8 FILLER_21_0 ();
 sg13g2_decap_8 FILLER_21_11 ();
 sg13g2_decap_8 FILLER_21_18 ();
 sg13g2_fill_1 FILLER_21_25 ();
 sg13g2_decap_8 FILLER_21_30 ();
 sg13g2_decap_8 FILLER_21_37 ();
 sg13g2_decap_4 FILLER_21_44 ();
 sg13g2_fill_1 FILLER_21_48 ();
 sg13g2_fill_2 FILLER_21_52 ();
 sg13g2_fill_1 FILLER_21_54 ();
 sg13g2_decap_4 FILLER_21_64 ();
 sg13g2_decap_8 FILLER_21_74 ();
 sg13g2_decap_8 FILLER_21_81 ();
 sg13g2_decap_8 FILLER_21_88 ();
 sg13g2_fill_1 FILLER_21_95 ();
 sg13g2_fill_2 FILLER_21_101 ();
 sg13g2_fill_1 FILLER_21_103 ();
 sg13g2_decap_4 FILLER_21_107 ();
 sg13g2_fill_2 FILLER_21_131 ();
 sg13g2_fill_2 FILLER_21_140 ();
 sg13g2_fill_1 FILLER_21_142 ();
 sg13g2_decap_8 FILLER_21_148 ();
 sg13g2_fill_2 FILLER_21_155 ();
 sg13g2_fill_1 FILLER_21_157 ();
 sg13g2_fill_2 FILLER_21_193 ();
 sg13g2_decap_4 FILLER_21_201 ();
 sg13g2_fill_2 FILLER_21_205 ();
 sg13g2_fill_2 FILLER_21_211 ();
 sg13g2_fill_1 FILLER_21_213 ();
 sg13g2_fill_1 FILLER_21_218 ();
 sg13g2_fill_1 FILLER_21_229 ();
 sg13g2_decap_8 FILLER_21_234 ();
 sg13g2_fill_2 FILLER_21_241 ();
 sg13g2_fill_1 FILLER_21_243 ();
 sg13g2_fill_1 FILLER_21_257 ();
 sg13g2_decap_4 FILLER_21_262 ();
 sg13g2_fill_2 FILLER_21_280 ();
 sg13g2_fill_1 FILLER_21_290 ();
 sg13g2_decap_8 FILLER_21_297 ();
 sg13g2_fill_1 FILLER_21_316 ();
 sg13g2_decap_8 FILLER_21_321 ();
 sg13g2_fill_2 FILLER_21_328 ();
 sg13g2_fill_1 FILLER_21_330 ();
 sg13g2_decap_4 FILLER_21_339 ();
 sg13g2_decap_8 FILLER_21_348 ();
 sg13g2_decap_8 FILLER_21_355 ();
 sg13g2_decap_8 FILLER_21_371 ();
 sg13g2_fill_2 FILLER_21_378 ();
 sg13g2_decap_4 FILLER_21_385 ();
 sg13g2_fill_2 FILLER_21_389 ();
 sg13g2_fill_2 FILLER_21_401 ();
 sg13g2_fill_1 FILLER_21_403 ();
 sg13g2_decap_8 FILLER_22_0 ();
 sg13g2_fill_1 FILLER_22_7 ();
 sg13g2_decap_8 FILLER_22_16 ();
 sg13g2_fill_1 FILLER_22_23 ();
 sg13g2_decap_8 FILLER_22_28 ();
 sg13g2_decap_8 FILLER_22_35 ();
 sg13g2_decap_4 FILLER_22_42 ();
 sg13g2_fill_1 FILLER_22_68 ();
 sg13g2_decap_8 FILLER_22_74 ();
 sg13g2_decap_4 FILLER_22_81 ();
 sg13g2_fill_1 FILLER_22_85 ();
 sg13g2_fill_2 FILLER_22_95 ();
 sg13g2_decap_8 FILLER_22_102 ();
 sg13g2_decap_8 FILLER_22_109 ();
 sg13g2_decap_4 FILLER_22_116 ();
 sg13g2_fill_1 FILLER_22_120 ();
 sg13g2_fill_2 FILLER_22_126 ();
 sg13g2_fill_1 FILLER_22_132 ();
 sg13g2_fill_2 FILLER_22_137 ();
 sg13g2_fill_1 FILLER_22_139 ();
 sg13g2_fill_1 FILLER_22_144 ();
 sg13g2_fill_2 FILLER_22_150 ();
 sg13g2_fill_1 FILLER_22_152 ();
 sg13g2_decap_8 FILLER_22_158 ();
 sg13g2_fill_2 FILLER_22_165 ();
 sg13g2_fill_1 FILLER_22_167 ();
 sg13g2_decap_4 FILLER_22_172 ();
 sg13g2_fill_1 FILLER_22_176 ();
 sg13g2_fill_2 FILLER_22_182 ();
 sg13g2_fill_1 FILLER_22_184 ();
 sg13g2_fill_1 FILLER_22_190 ();
 sg13g2_fill_1 FILLER_22_194 ();
 sg13g2_fill_2 FILLER_22_200 ();
 sg13g2_fill_1 FILLER_22_206 ();
 sg13g2_fill_1 FILLER_22_211 ();
 sg13g2_fill_1 FILLER_22_220 ();
 sg13g2_fill_1 FILLER_22_247 ();
 sg13g2_fill_1 FILLER_22_257 ();
 sg13g2_fill_2 FILLER_22_262 ();
 sg13g2_fill_1 FILLER_22_269 ();
 sg13g2_fill_2 FILLER_22_282 ();
 sg13g2_fill_2 FILLER_22_293 ();
 sg13g2_decap_8 FILLER_22_300 ();
 sg13g2_fill_2 FILLER_22_312 ();
 sg13g2_decap_4 FILLER_22_322 ();
 sg13g2_fill_2 FILLER_22_351 ();
 sg13g2_fill_1 FILLER_22_360 ();
 sg13g2_decap_4 FILLER_22_374 ();
 sg13g2_fill_2 FILLER_22_394 ();
 sg13g2_fill_1 FILLER_22_396 ();
 sg13g2_decap_8 FILLER_22_403 ();
 sg13g2_fill_1 FILLER_22_410 ();
 sg13g2_decap_8 FILLER_22_415 ();
 sg13g2_decap_8 FILLER_22_422 ();
 sg13g2_fill_1 FILLER_22_429 ();
 sg13g2_decap_8 FILLER_23_0 ();
 sg13g2_decap_4 FILLER_23_7 ();
 sg13g2_fill_2 FILLER_23_15 ();
 sg13g2_fill_2 FILLER_23_43 ();
 sg13g2_fill_2 FILLER_23_53 ();
 sg13g2_decap_8 FILLER_23_69 ();
 sg13g2_decap_8 FILLER_23_76 ();
 sg13g2_decap_8 FILLER_23_83 ();
 sg13g2_decap_4 FILLER_23_90 ();
 sg13g2_decap_4 FILLER_23_109 ();
 sg13g2_fill_1 FILLER_23_113 ();
 sg13g2_decap_8 FILLER_23_122 ();
 sg13g2_fill_1 FILLER_23_129 ();
 sg13g2_fill_2 FILLER_23_142 ();
 sg13g2_fill_1 FILLER_23_144 ();
 sg13g2_fill_2 FILLER_23_161 ();
 sg13g2_fill_1 FILLER_23_163 ();
 sg13g2_fill_1 FILLER_23_194 ();
 sg13g2_fill_2 FILLER_23_215 ();
 sg13g2_decap_8 FILLER_23_225 ();
 sg13g2_fill_2 FILLER_23_232 ();
 sg13g2_decap_8 FILLER_23_238 ();
 sg13g2_fill_2 FILLER_23_257 ();
 sg13g2_fill_1 FILLER_23_263 ();
 sg13g2_fill_1 FILLER_23_289 ();
 sg13g2_decap_8 FILLER_23_294 ();
 sg13g2_decap_8 FILLER_23_301 ();
 sg13g2_decap_4 FILLER_23_308 ();
 sg13g2_fill_1 FILLER_23_312 ();
 sg13g2_decap_8 FILLER_23_318 ();
 sg13g2_fill_1 FILLER_23_325 ();
 sg13g2_fill_1 FILLER_23_331 ();
 sg13g2_fill_1 FILLER_23_336 ();
 sg13g2_fill_1 FILLER_23_357 ();
 sg13g2_fill_2 FILLER_23_366 ();
 sg13g2_decap_8 FILLER_23_396 ();
 sg13g2_decap_8 FILLER_23_407 ();
 sg13g2_decap_8 FILLER_23_414 ();
 sg13g2_decap_8 FILLER_23_421 ();
 sg13g2_fill_2 FILLER_23_428 ();
 sg13g2_decap_8 FILLER_24_0 ();
 sg13g2_fill_2 FILLER_24_11 ();
 sg13g2_fill_1 FILLER_24_13 ();
 sg13g2_fill_2 FILLER_24_19 ();
 sg13g2_fill_2 FILLER_24_29 ();
 sg13g2_fill_1 FILLER_24_31 ();
 sg13g2_decap_8 FILLER_24_40 ();
 sg13g2_decap_8 FILLER_24_47 ();
 sg13g2_fill_2 FILLER_24_54 ();
 sg13g2_fill_1 FILLER_24_56 ();
 sg13g2_fill_2 FILLER_24_65 ();
 sg13g2_fill_1 FILLER_24_67 ();
 sg13g2_decap_4 FILLER_24_76 ();
 sg13g2_fill_1 FILLER_24_80 ();
 sg13g2_fill_1 FILLER_24_94 ();
 sg13g2_decap_8 FILLER_24_107 ();
 sg13g2_fill_2 FILLER_24_114 ();
 sg13g2_decap_4 FILLER_24_121 ();
 sg13g2_fill_2 FILLER_24_154 ();
 sg13g2_fill_1 FILLER_24_156 ();
 sg13g2_decap_8 FILLER_24_161 ();
 sg13g2_decap_8 FILLER_24_168 ();
 sg13g2_fill_1 FILLER_24_175 ();
 sg13g2_fill_2 FILLER_24_191 ();
 sg13g2_decap_4 FILLER_24_201 ();
 sg13g2_fill_2 FILLER_24_239 ();
 sg13g2_decap_8 FILLER_24_250 ();
 sg13g2_fill_1 FILLER_24_257 ();
 sg13g2_decap_4 FILLER_24_279 ();
 sg13g2_fill_2 FILLER_24_288 ();
 sg13g2_fill_1 FILLER_24_290 ();
 sg13g2_decap_8 FILLER_24_298 ();
 sg13g2_decap_8 FILLER_24_305 ();
 sg13g2_fill_1 FILLER_24_312 ();
 sg13g2_fill_2 FILLER_24_338 ();
 sg13g2_decap_4 FILLER_24_353 ();
 sg13g2_fill_2 FILLER_24_376 ();
 sg13g2_fill_1 FILLER_24_378 ();
 sg13g2_fill_2 FILLER_24_387 ();
 sg13g2_decap_4 FILLER_24_393 ();
 sg13g2_decap_8 FILLER_24_423 ();
 sg13g2_fill_1 FILLER_25_0 ();
 sg13g2_fill_1 FILLER_25_27 ();
 sg13g2_fill_1 FILLER_25_32 ();
 sg13g2_fill_2 FILLER_25_43 ();
 sg13g2_decap_8 FILLER_25_53 ();
 sg13g2_fill_1 FILLER_25_60 ();
 sg13g2_fill_2 FILLER_25_72 ();
 sg13g2_fill_1 FILLER_25_74 ();
 sg13g2_decap_8 FILLER_25_80 ();
 sg13g2_decap_8 FILLER_25_93 ();
 sg13g2_decap_8 FILLER_25_100 ();
 sg13g2_fill_2 FILLER_25_107 ();
 sg13g2_decap_4 FILLER_25_119 ();
 sg13g2_fill_2 FILLER_25_123 ();
 sg13g2_fill_1 FILLER_25_133 ();
 sg13g2_fill_1 FILLER_25_138 ();
 sg13g2_decap_8 FILLER_25_151 ();
 sg13g2_decap_8 FILLER_25_158 ();
 sg13g2_decap_8 FILLER_25_165 ();
 sg13g2_decap_8 FILLER_25_172 ();
 sg13g2_fill_2 FILLER_25_179 ();
 sg13g2_fill_1 FILLER_25_181 ();
 sg13g2_decap_4 FILLER_25_197 ();
 sg13g2_fill_2 FILLER_25_201 ();
 sg13g2_decap_8 FILLER_25_212 ();
 sg13g2_decap_8 FILLER_25_223 ();
 sg13g2_decap_4 FILLER_25_230 ();
 sg13g2_fill_1 FILLER_25_234 ();
 sg13g2_fill_1 FILLER_25_240 ();
 sg13g2_decap_4 FILLER_25_247 ();
 sg13g2_fill_1 FILLER_25_251 ();
 sg13g2_decap_4 FILLER_25_257 ();
 sg13g2_fill_2 FILLER_25_261 ();
 sg13g2_fill_2 FILLER_25_268 ();
 sg13g2_decap_8 FILLER_25_275 ();
 sg13g2_fill_2 FILLER_25_282 ();
 sg13g2_decap_8 FILLER_25_297 ();
 sg13g2_fill_1 FILLER_25_304 ();
 sg13g2_fill_2 FILLER_25_315 ();
 sg13g2_fill_1 FILLER_25_317 ();
 sg13g2_decap_4 FILLER_25_322 ();
 sg13g2_decap_8 FILLER_25_331 ();
 sg13g2_decap_8 FILLER_25_338 ();
 sg13g2_decap_8 FILLER_25_345 ();
 sg13g2_decap_4 FILLER_25_352 ();
 sg13g2_decap_8 FILLER_25_366 ();
 sg13g2_decap_8 FILLER_25_373 ();
 sg13g2_fill_1 FILLER_25_380 ();
 sg13g2_fill_2 FILLER_25_386 ();
 sg13g2_fill_1 FILLER_25_388 ();
 sg13g2_decap_8 FILLER_25_398 ();
 sg13g2_decap_4 FILLER_25_405 ();
 sg13g2_fill_2 FILLER_25_409 ();
 sg13g2_decap_8 FILLER_25_415 ();
 sg13g2_decap_8 FILLER_25_422 ();
 sg13g2_fill_1 FILLER_25_429 ();
 sg13g2_decap_8 FILLER_26_0 ();
 sg13g2_decap_8 FILLER_26_7 ();
 sg13g2_decap_8 FILLER_26_14 ();
 sg13g2_decap_8 FILLER_26_21 ();
 sg13g2_fill_1 FILLER_26_42 ();
 sg13g2_decap_4 FILLER_26_51 ();
 sg13g2_fill_1 FILLER_26_55 ();
 sg13g2_fill_2 FILLER_26_68 ();
 sg13g2_fill_2 FILLER_26_92 ();
 sg13g2_decap_8 FILLER_26_104 ();
 sg13g2_decap_8 FILLER_26_111 ();
 sg13g2_decap_8 FILLER_26_118 ();
 sg13g2_decap_4 FILLER_26_125 ();
 sg13g2_decap_4 FILLER_26_163 ();
 sg13g2_fill_1 FILLER_26_167 ();
 sg13g2_fill_2 FILLER_26_172 ();
 sg13g2_fill_1 FILLER_26_174 ();
 sg13g2_fill_2 FILLER_26_179 ();
 sg13g2_fill_1 FILLER_26_181 ();
 sg13g2_fill_2 FILLER_26_203 ();
 sg13g2_fill_1 FILLER_26_205 ();
 sg13g2_fill_1 FILLER_26_215 ();
 sg13g2_decap_4 FILLER_26_233 ();
 sg13g2_fill_1 FILLER_26_237 ();
 sg13g2_decap_8 FILLER_26_243 ();
 sg13g2_decap_8 FILLER_26_250 ();
 sg13g2_decap_4 FILLER_26_257 ();
 sg13g2_decap_8 FILLER_26_266 ();
 sg13g2_fill_1 FILLER_26_273 ();
 sg13g2_decap_8 FILLER_26_300 ();
 sg13g2_decap_8 FILLER_26_307 ();
 sg13g2_decap_8 FILLER_26_314 ();
 sg13g2_fill_2 FILLER_26_321 ();
 sg13g2_fill_2 FILLER_26_342 ();
 sg13g2_decap_8 FILLER_26_348 ();
 sg13g2_fill_1 FILLER_26_355 ();
 sg13g2_decap_4 FILLER_26_361 ();
 sg13g2_fill_1 FILLER_26_365 ();
 sg13g2_fill_2 FILLER_26_388 ();
 sg13g2_fill_1 FILLER_26_403 ();
 sg13g2_decap_8 FILLER_27_0 ();
 sg13g2_decap_8 FILLER_27_7 ();
 sg13g2_fill_2 FILLER_27_14 ();
 sg13g2_fill_2 FILLER_27_28 ();
 sg13g2_fill_1 FILLER_27_30 ();
 sg13g2_fill_2 FILLER_27_42 ();
 sg13g2_fill_1 FILLER_27_44 ();
 sg13g2_fill_2 FILLER_27_91 ();
 sg13g2_decap_8 FILLER_27_102 ();
 sg13g2_decap_8 FILLER_27_109 ();
 sg13g2_fill_2 FILLER_27_116 ();
 sg13g2_decap_4 FILLER_27_130 ();
 sg13g2_fill_2 FILLER_27_134 ();
 sg13g2_fill_1 FILLER_27_140 ();
 sg13g2_fill_1 FILLER_27_169 ();
 sg13g2_fill_1 FILLER_27_183 ();
 sg13g2_fill_1 FILLER_27_194 ();
 sg13g2_fill_1 FILLER_27_210 ();
 sg13g2_fill_2 FILLER_27_216 ();
 sg13g2_fill_1 FILLER_27_218 ();
 sg13g2_fill_2 FILLER_27_245 ();
 sg13g2_decap_4 FILLER_27_253 ();
 sg13g2_fill_1 FILLER_27_257 ();
 sg13g2_fill_2 FILLER_27_279 ();
 sg13g2_fill_1 FILLER_27_281 ();
 sg13g2_fill_1 FILLER_27_287 ();
 sg13g2_decap_8 FILLER_27_297 ();
 sg13g2_decap_8 FILLER_27_304 ();
 sg13g2_decap_8 FILLER_27_311 ();
 sg13g2_fill_2 FILLER_27_322 ();
 sg13g2_fill_1 FILLER_27_324 ();
 sg13g2_fill_2 FILLER_27_330 ();
 sg13g2_fill_1 FILLER_27_332 ();
 sg13g2_fill_1 FILLER_27_337 ();
 sg13g2_fill_1 FILLER_27_343 ();
 sg13g2_fill_2 FILLER_27_349 ();
 sg13g2_fill_2 FILLER_27_359 ();
 sg13g2_fill_1 FILLER_27_361 ();
 sg13g2_fill_1 FILLER_27_372 ();
 sg13g2_decap_8 FILLER_27_378 ();
 sg13g2_fill_2 FILLER_27_385 ();
 sg13g2_fill_2 FILLER_27_396 ();
 sg13g2_decap_4 FILLER_27_424 ();
 sg13g2_fill_2 FILLER_27_428 ();
 sg13g2_fill_1 FILLER_28_0 ();
 sg13g2_fill_1 FILLER_28_27 ();
 sg13g2_decap_4 FILLER_28_33 ();
 sg13g2_fill_2 FILLER_28_37 ();
 sg13g2_fill_1 FILLER_28_67 ();
 sg13g2_fill_1 FILLER_28_81 ();
 sg13g2_fill_1 FILLER_28_94 ();
 sg13g2_fill_1 FILLER_28_103 ();
 sg13g2_decap_8 FILLER_28_133 ();
 sg13g2_fill_2 FILLER_28_140 ();
 sg13g2_fill_1 FILLER_28_147 ();
 sg13g2_fill_1 FILLER_28_153 ();
 sg13g2_decap_4 FILLER_28_159 ();
 sg13g2_fill_2 FILLER_28_163 ();
 sg13g2_fill_2 FILLER_28_174 ();
 sg13g2_fill_1 FILLER_28_185 ();
 sg13g2_decap_8 FILLER_28_194 ();
 sg13g2_decap_8 FILLER_28_201 ();
 sg13g2_fill_2 FILLER_28_211 ();
 sg13g2_fill_1 FILLER_28_213 ();
 sg13g2_decap_4 FILLER_28_222 ();
 sg13g2_fill_2 FILLER_28_226 ();
 sg13g2_decap_8 FILLER_28_232 ();
 sg13g2_fill_2 FILLER_28_239 ();
 sg13g2_decap_8 FILLER_28_247 ();
 sg13g2_decap_4 FILLER_28_254 ();
 sg13g2_fill_1 FILLER_28_258 ();
 sg13g2_fill_1 FILLER_28_287 ();
 sg13g2_fill_2 FILLER_28_293 ();
 sg13g2_fill_1 FILLER_28_295 ();
 sg13g2_fill_2 FILLER_28_308 ();
 sg13g2_fill_1 FILLER_28_310 ();
 sg13g2_fill_2 FILLER_28_320 ();
 sg13g2_fill_1 FILLER_28_327 ();
 sg13g2_decap_8 FILLER_28_353 ();
 sg13g2_decap_8 FILLER_28_360 ();
 sg13g2_decap_8 FILLER_28_367 ();
 sg13g2_fill_2 FILLER_28_374 ();
 sg13g2_fill_2 FILLER_28_390 ();
 sg13g2_fill_1 FILLER_28_417 ();
 sg13g2_decap_4 FILLER_28_426 ();
 sg13g2_decap_8 FILLER_29_0 ();
 sg13g2_decap_8 FILLER_29_11 ();
 sg13g2_decap_4 FILLER_29_18 ();
 sg13g2_fill_1 FILLER_29_22 ();
 sg13g2_fill_2 FILLER_29_63 ();
 sg13g2_decap_4 FILLER_29_76 ();
 sg13g2_fill_1 FILLER_29_92 ();
 sg13g2_decap_8 FILLER_29_106 ();
 sg13g2_decap_8 FILLER_29_113 ();
 sg13g2_decap_8 FILLER_29_120 ();
 sg13g2_decap_8 FILLER_29_127 ();
 sg13g2_decap_8 FILLER_29_134 ();
 sg13g2_fill_2 FILLER_29_141 ();
 sg13g2_decap_4 FILLER_29_167 ();
 sg13g2_fill_1 FILLER_29_171 ();
 sg13g2_decap_4 FILLER_29_177 ();
 sg13g2_fill_2 FILLER_29_219 ();
 sg13g2_fill_1 FILLER_29_221 ();
 sg13g2_decap_4 FILLER_29_254 ();
 sg13g2_fill_1 FILLER_29_258 ();
 sg13g2_fill_2 FILLER_29_277 ();
 sg13g2_fill_1 FILLER_29_288 ();
 sg13g2_fill_2 FILLER_29_297 ();
 sg13g2_decap_4 FILLER_29_304 ();
 sg13g2_fill_1 FILLER_29_308 ();
 sg13g2_fill_1 FILLER_29_322 ();
 sg13g2_fill_2 FILLER_29_353 ();
 sg13g2_decap_8 FILLER_29_362 ();
 sg13g2_decap_8 FILLER_29_369 ();
 sg13g2_decap_8 FILLER_29_376 ();
 sg13g2_fill_1 FILLER_29_383 ();
 sg13g2_decap_8 FILLER_29_397 ();
 sg13g2_decap_8 FILLER_29_412 ();
 sg13g2_decap_8 FILLER_29_419 ();
 sg13g2_decap_4 FILLER_29_426 ();
 sg13g2_decap_4 FILLER_30_0 ();
 sg13g2_fill_2 FILLER_30_4 ();
 sg13g2_fill_2 FILLER_30_23 ();
 sg13g2_fill_2 FILLER_30_29 ();
 sg13g2_fill_2 FILLER_30_36 ();
 sg13g2_fill_1 FILLER_30_38 ();
 sg13g2_fill_2 FILLER_30_44 ();
 sg13g2_fill_1 FILLER_30_46 ();
 sg13g2_fill_2 FILLER_30_52 ();
 sg13g2_fill_2 FILLER_30_59 ();
 sg13g2_fill_1 FILLER_30_61 ();
 sg13g2_decap_4 FILLER_30_79 ();
 sg13g2_decap_4 FILLER_30_95 ();
 sg13g2_decap_4 FILLER_30_107 ();
 sg13g2_fill_1 FILLER_30_111 ();
 sg13g2_decap_4 FILLER_30_124 ();
 sg13g2_fill_1 FILLER_30_128 ();
 sg13g2_decap_4 FILLER_30_134 ();
 sg13g2_fill_1 FILLER_30_138 ();
 sg13g2_fill_1 FILLER_30_156 ();
 sg13g2_fill_1 FILLER_30_169 ();
 sg13g2_decap_8 FILLER_30_174 ();
 sg13g2_fill_2 FILLER_30_181 ();
 sg13g2_fill_1 FILLER_30_183 ();
 sg13g2_decap_4 FILLER_30_189 ();
 sg13g2_fill_1 FILLER_30_193 ();
 sg13g2_decap_4 FILLER_30_204 ();
 sg13g2_fill_1 FILLER_30_208 ();
 sg13g2_decap_8 FILLER_30_214 ();
 sg13g2_decap_4 FILLER_30_221 ();
 sg13g2_fill_1 FILLER_30_225 ();
 sg13g2_decap_8 FILLER_30_234 ();
 sg13g2_fill_2 FILLER_30_261 ();
 sg13g2_fill_2 FILLER_30_267 ();
 sg13g2_fill_2 FILLER_30_277 ();
 sg13g2_decap_8 FILLER_30_294 ();
 sg13g2_fill_2 FILLER_30_301 ();
 sg13g2_fill_1 FILLER_30_318 ();
 sg13g2_decap_4 FILLER_30_323 ();
 sg13g2_fill_2 FILLER_30_331 ();
 sg13g2_decap_8 FILLER_30_358 ();
 sg13g2_decap_4 FILLER_30_365 ();
 sg13g2_fill_2 FILLER_30_369 ();
 sg13g2_fill_1 FILLER_30_421 ();
 sg13g2_decap_4 FILLER_30_426 ();
 sg13g2_decap_8 FILLER_31_0 ();
 sg13g2_decap_4 FILLER_31_7 ();
 sg13g2_decap_4 FILLER_31_42 ();
 sg13g2_decap_8 FILLER_31_55 ();
 sg13g2_decap_8 FILLER_31_62 ();
 sg13g2_decap_8 FILLER_31_75 ();
 sg13g2_fill_1 FILLER_31_82 ();
 sg13g2_decap_8 FILLER_31_93 ();
 sg13g2_fill_1 FILLER_31_100 ();
 sg13g2_fill_1 FILLER_31_113 ();
 sg13g2_decap_4 FILLER_31_119 ();
 sg13g2_fill_1 FILLER_31_123 ();
 sg13g2_fill_2 FILLER_31_141 ();
 sg13g2_fill_1 FILLER_31_143 ();
 sg13g2_decap_8 FILLER_31_167 ();
 sg13g2_decap_8 FILLER_31_174 ();
 sg13g2_fill_2 FILLER_31_181 ();
 sg13g2_fill_1 FILLER_31_183 ();
 sg13g2_fill_1 FILLER_31_192 ();
 sg13g2_fill_2 FILLER_31_231 ();
 sg13g2_fill_2 FILLER_31_241 ();
 sg13g2_decap_4 FILLER_31_268 ();
 sg13g2_fill_1 FILLER_31_272 ();
 sg13g2_decap_8 FILLER_31_293 ();
 sg13g2_decap_4 FILLER_31_300 ();
 sg13g2_fill_2 FILLER_31_304 ();
 sg13g2_fill_2 FILLER_31_314 ();
 sg13g2_decap_8 FILLER_31_334 ();
 sg13g2_decap_4 FILLER_31_345 ();
 sg13g2_fill_1 FILLER_31_349 ();
 sg13g2_decap_8 FILLER_31_361 ();
 sg13g2_fill_1 FILLER_31_368 ();
 sg13g2_decap_4 FILLER_31_382 ();
 sg13g2_fill_1 FILLER_31_386 ();
 sg13g2_fill_2 FILLER_31_392 ();
 sg13g2_decap_4 FILLER_31_399 ();
 sg13g2_decap_4 FILLER_31_411 ();
 sg13g2_decap_8 FILLER_31_423 ();
 sg13g2_decap_8 FILLER_32_0 ();
 sg13g2_decap_8 FILLER_32_7 ();
 sg13g2_fill_2 FILLER_32_14 ();
 sg13g2_decap_8 FILLER_32_20 ();
 sg13g2_fill_1 FILLER_32_27 ();
 sg13g2_decap_4 FILLER_32_37 ();
 sg13g2_fill_1 FILLER_32_41 ();
 sg13g2_decap_8 FILLER_32_61 ();
 sg13g2_fill_1 FILLER_32_68 ();
 sg13g2_decap_8 FILLER_32_89 ();
 sg13g2_fill_1 FILLER_32_96 ();
 sg13g2_fill_1 FILLER_32_112 ();
 sg13g2_decap_4 FILLER_32_118 ();
 sg13g2_fill_1 FILLER_32_122 ();
 sg13g2_fill_2 FILLER_32_135 ();
 sg13g2_fill_1 FILLER_32_137 ();
 sg13g2_decap_8 FILLER_32_162 ();
 sg13g2_fill_1 FILLER_32_169 ();
 sg13g2_decap_8 FILLER_32_175 ();
 sg13g2_decap_8 FILLER_32_182 ();
 sg13g2_fill_2 FILLER_32_189 ();
 sg13g2_decap_4 FILLER_32_195 ();
 sg13g2_fill_1 FILLER_32_199 ();
 sg13g2_decap_8 FILLER_32_204 ();
 sg13g2_decap_4 FILLER_32_211 ();
 sg13g2_decap_8 FILLER_32_219 ();
 sg13g2_decap_8 FILLER_32_226 ();
 sg13g2_decap_8 FILLER_32_233 ();
 sg13g2_fill_2 FILLER_32_248 ();
 sg13g2_fill_1 FILLER_32_250 ();
 sg13g2_fill_1 FILLER_32_256 ();
 sg13g2_fill_2 FILLER_32_262 ();
 sg13g2_decap_4 FILLER_32_269 ();
 sg13g2_fill_2 FILLER_32_273 ();
 sg13g2_decap_4 FILLER_32_278 ();
 sg13g2_fill_2 FILLER_32_295 ();
 sg13g2_fill_1 FILLER_32_302 ();
 sg13g2_decap_8 FILLER_32_307 ();
 sg13g2_decap_8 FILLER_32_318 ();
 sg13g2_fill_1 FILLER_32_325 ();
 sg13g2_decap_4 FILLER_32_338 ();
 sg13g2_fill_1 FILLER_32_342 ();
 sg13g2_fill_2 FILLER_32_380 ();
 sg13g2_fill_2 FILLER_32_390 ();
 sg13g2_decap_8 FILLER_33_0 ();
 sg13g2_fill_1 FILLER_33_54 ();
 sg13g2_decap_4 FILLER_33_60 ();
 sg13g2_fill_2 FILLER_33_64 ();
 sg13g2_fill_1 FILLER_33_75 ();
 sg13g2_decap_8 FILLER_33_86 ();
 sg13g2_fill_2 FILLER_33_93 ();
 sg13g2_fill_1 FILLER_33_95 ();
 sg13g2_fill_1 FILLER_33_100 ();
 sg13g2_decap_8 FILLER_33_113 ();
 sg13g2_decap_4 FILLER_33_120 ();
 sg13g2_decap_8 FILLER_33_132 ();
 sg13g2_decap_8 FILLER_33_139 ();
 sg13g2_decap_4 FILLER_33_146 ();
 sg13g2_fill_1 FILLER_33_150 ();
 sg13g2_fill_2 FILLER_33_163 ();
 sg13g2_fill_2 FILLER_33_185 ();
 sg13g2_fill_2 FILLER_33_201 ();
 sg13g2_fill_1 FILLER_33_208 ();
 sg13g2_decap_8 FILLER_33_214 ();
 sg13g2_decap_8 FILLER_33_221 ();
 sg13g2_decap_8 FILLER_33_228 ();
 sg13g2_decap_8 FILLER_33_235 ();
 sg13g2_decap_8 FILLER_33_242 ();
 sg13g2_fill_1 FILLER_33_249 ();
 sg13g2_decap_4 FILLER_33_280 ();
 sg13g2_fill_2 FILLER_33_288 ();
 sg13g2_fill_1 FILLER_33_290 ();
 sg13g2_decap_4 FILLER_33_295 ();
 sg13g2_fill_2 FILLER_33_299 ();
 sg13g2_fill_1 FILLER_33_320 ();
 sg13g2_fill_2 FILLER_33_326 ();
 sg13g2_decap_4 FILLER_33_333 ();
 sg13g2_fill_2 FILLER_33_342 ();
 sg13g2_fill_1 FILLER_33_360 ();
 sg13g2_fill_2 FILLER_33_365 ();
 sg13g2_fill_1 FILLER_33_367 ();
 sg13g2_fill_2 FILLER_33_372 ();
 sg13g2_fill_1 FILLER_33_374 ();
 sg13g2_decap_8 FILLER_33_417 ();
 sg13g2_decap_4 FILLER_33_424 ();
 sg13g2_fill_2 FILLER_33_428 ();
 sg13g2_decap_4 FILLER_34_0 ();
 sg13g2_fill_1 FILLER_34_4 ();
 sg13g2_decap_4 FILLER_34_9 ();
 sg13g2_decap_8 FILLER_34_25 ();
 sg13g2_fill_1 FILLER_34_32 ();
 sg13g2_decap_8 FILLER_34_58 ();
 sg13g2_fill_2 FILLER_34_65 ();
 sg13g2_fill_1 FILLER_34_67 ();
 sg13g2_decap_8 FILLER_34_73 ();
 sg13g2_decap_8 FILLER_34_80 ();
 sg13g2_fill_2 FILLER_34_87 ();
 sg13g2_fill_1 FILLER_34_107 ();
 sg13g2_decap_8 FILLER_34_114 ();
 sg13g2_decap_8 FILLER_34_121 ();
 sg13g2_fill_1 FILLER_34_128 ();
 sg13g2_decap_4 FILLER_34_139 ();
 sg13g2_fill_2 FILLER_34_143 ();
 sg13g2_decap_4 FILLER_34_150 ();
 sg13g2_fill_2 FILLER_34_154 ();
 sg13g2_fill_2 FILLER_34_163 ();
 sg13g2_fill_1 FILLER_34_165 ();
 sg13g2_fill_1 FILLER_34_184 ();
 sg13g2_fill_1 FILLER_34_190 ();
 sg13g2_fill_1 FILLER_34_195 ();
 sg13g2_fill_1 FILLER_34_201 ();
 sg13g2_decap_8 FILLER_34_218 ();
 sg13g2_decap_4 FILLER_34_225 ();
 sg13g2_fill_2 FILLER_34_229 ();
 sg13g2_fill_1 FILLER_34_239 ();
 sg13g2_fill_1 FILLER_34_248 ();
 sg13g2_fill_2 FILLER_34_254 ();
 sg13g2_fill_2 FILLER_34_261 ();
 sg13g2_fill_2 FILLER_34_268 ();
 sg13g2_decap_4 FILLER_34_279 ();
 sg13g2_fill_2 FILLER_34_283 ();
 sg13g2_fill_1 FILLER_34_318 ();
 sg13g2_decap_8 FILLER_34_327 ();
 sg13g2_decap_4 FILLER_34_342 ();
 sg13g2_decap_4 FILLER_34_350 ();
 sg13g2_fill_1 FILLER_34_354 ();
 sg13g2_decap_8 FILLER_34_358 ();
 sg13g2_decap_4 FILLER_34_371 ();
 sg13g2_decap_4 FILLER_34_384 ();
 sg13g2_decap_8 FILLER_34_410 ();
 sg13g2_decap_8 FILLER_34_422 ();
 sg13g2_fill_1 FILLER_34_429 ();
 sg13g2_decap_8 FILLER_35_0 ();
 sg13g2_decap_8 FILLER_35_7 ();
 sg13g2_decap_8 FILLER_35_14 ();
 sg13g2_decap_8 FILLER_35_21 ();
 sg13g2_fill_1 FILLER_35_33 ();
 sg13g2_decap_4 FILLER_35_40 ();
 sg13g2_fill_2 FILLER_35_44 ();
 sg13g2_fill_1 FILLER_35_51 ();
 sg13g2_fill_2 FILLER_35_56 ();
 sg13g2_fill_2 FILLER_35_63 ();
 sg13g2_decap_8 FILLER_35_103 ();
 sg13g2_decap_4 FILLER_35_110 ();
 sg13g2_fill_1 FILLER_35_114 ();
 sg13g2_fill_1 FILLER_35_123 ();
 sg13g2_fill_2 FILLER_35_140 ();
 sg13g2_fill_1 FILLER_35_142 ();
 sg13g2_decap_8 FILLER_35_147 ();
 sg13g2_decap_8 FILLER_35_154 ();
 sg13g2_decap_8 FILLER_35_161 ();
 sg13g2_decap_8 FILLER_35_168 ();
 sg13g2_fill_2 FILLER_35_175 ();
 sg13g2_decap_8 FILLER_35_185 ();
 sg13g2_decap_8 FILLER_35_192 ();
 sg13g2_fill_2 FILLER_35_199 ();
 sg13g2_decap_4 FILLER_35_206 ();
 sg13g2_decap_8 FILLER_35_218 ();
 sg13g2_decap_8 FILLER_35_225 ();
 sg13g2_decap_4 FILLER_35_232 ();
 sg13g2_fill_2 FILLER_35_241 ();
 sg13g2_fill_1 FILLER_35_243 ();
 sg13g2_decap_4 FILLER_35_248 ();
 sg13g2_decap_8 FILLER_35_262 ();
 sg13g2_decap_8 FILLER_35_269 ();
 sg13g2_decap_8 FILLER_35_276 ();
 sg13g2_fill_1 FILLER_35_283 ();
 sg13g2_fill_2 FILLER_35_294 ();
 sg13g2_fill_1 FILLER_35_296 ();
 sg13g2_fill_1 FILLER_35_301 ();
 sg13g2_fill_2 FILLER_35_314 ();
 sg13g2_fill_2 FILLER_35_342 ();
 sg13g2_fill_1 FILLER_35_344 ();
 sg13g2_fill_1 FILLER_35_354 ();
 sg13g2_decap_8 FILLER_35_360 ();
 sg13g2_fill_1 FILLER_35_367 ();
 sg13g2_fill_1 FILLER_35_393 ();
 sg13g2_fill_2 FILLER_35_408 ();
 sg13g2_fill_1 FILLER_35_410 ();
 sg13g2_decap_8 FILLER_35_421 ();
 sg13g2_fill_2 FILLER_35_428 ();
 sg13g2_decap_8 FILLER_36_0 ();
 sg13g2_decap_8 FILLER_36_7 ();
 sg13g2_decap_8 FILLER_36_14 ();
 sg13g2_decap_4 FILLER_36_21 ();
 sg13g2_fill_2 FILLER_36_41 ();
 sg13g2_fill_1 FILLER_36_43 ();
 sg13g2_fill_2 FILLER_36_52 ();
 sg13g2_fill_2 FILLER_36_72 ();
 sg13g2_fill_1 FILLER_36_74 ();
 sg13g2_fill_2 FILLER_36_83 ();
 sg13g2_fill_1 FILLER_36_85 ();
 sg13g2_fill_2 FILLER_36_90 ();
 sg13g2_fill_1 FILLER_36_92 ();
 sg13g2_decap_4 FILLER_36_101 ();
 sg13g2_fill_2 FILLER_36_105 ();
 sg13g2_decap_4 FILLER_36_112 ();
 sg13g2_fill_1 FILLER_36_132 ();
 sg13g2_fill_2 FILLER_36_141 ();
 sg13g2_decap_8 FILLER_36_153 ();
 sg13g2_decap_4 FILLER_36_160 ();
 sg13g2_fill_2 FILLER_36_164 ();
 sg13g2_decap_4 FILLER_36_170 ();
 sg13g2_fill_2 FILLER_36_174 ();
 sg13g2_fill_1 FILLER_36_232 ();
 sg13g2_decap_8 FILLER_36_259 ();
 sg13g2_decap_8 FILLER_36_266 ();
 sg13g2_decap_8 FILLER_36_273 ();
 sg13g2_decap_8 FILLER_36_280 ();
 sg13g2_decap_4 FILLER_36_287 ();
 sg13g2_fill_1 FILLER_36_291 ();
 sg13g2_fill_1 FILLER_36_310 ();
 sg13g2_decap_4 FILLER_36_328 ();
 sg13g2_decap_4 FILLER_36_337 ();
 sg13g2_fill_1 FILLER_36_350 ();
 sg13g2_decap_8 FILLER_36_361 ();
 sg13g2_decap_4 FILLER_36_368 ();
 sg13g2_decap_4 FILLER_36_376 ();
 sg13g2_decap_4 FILLER_36_391 ();
 sg13g2_fill_1 FILLER_36_395 ();
 sg13g2_decap_8 FILLER_36_401 ();
 sg13g2_decap_8 FILLER_36_408 ();
 sg13g2_fill_1 FILLER_36_415 ();
 sg13g2_decap_8 FILLER_36_420 ();
 sg13g2_fill_2 FILLER_36_427 ();
 sg13g2_fill_1 FILLER_36_429 ();
 sg13g2_decap_8 FILLER_37_0 ();
 sg13g2_fill_1 FILLER_37_7 ();
 sg13g2_fill_1 FILLER_37_12 ();
 sg13g2_decap_8 FILLER_37_17 ();
 sg13g2_fill_2 FILLER_37_24 ();
 sg13g2_fill_2 FILLER_37_30 ();
 sg13g2_fill_1 FILLER_37_32 ();
 sg13g2_fill_2 FILLER_37_37 ();
 sg13g2_fill_1 FILLER_37_39 ();
 sg13g2_decap_8 FILLER_37_44 ();
 sg13g2_decap_4 FILLER_37_51 ();
 sg13g2_fill_1 FILLER_37_55 ();
 sg13g2_decap_8 FILLER_37_61 ();
 sg13g2_decap_8 FILLER_37_68 ();
 sg13g2_fill_2 FILLER_37_75 ();
 sg13g2_fill_1 FILLER_37_84 ();
 sg13g2_fill_1 FILLER_37_95 ();
 sg13g2_fill_1 FILLER_37_102 ();
 sg13g2_fill_1 FILLER_37_107 ();
 sg13g2_fill_1 FILLER_37_112 ();
 sg13g2_fill_1 FILLER_37_123 ();
 sg13g2_fill_1 FILLER_37_128 ();
 sg13g2_decap_4 FILLER_37_193 ();
 sg13g2_decap_4 FILLER_37_201 ();
 sg13g2_decap_4 FILLER_37_209 ();
 sg13g2_decap_4 FILLER_37_217 ();
 sg13g2_fill_2 FILLER_37_225 ();
 sg13g2_fill_1 FILLER_37_227 ();
 sg13g2_fill_1 FILLER_37_232 ();
 sg13g2_fill_1 FILLER_37_259 ();
 sg13g2_fill_1 FILLER_37_268 ();
 sg13g2_decap_8 FILLER_37_273 ();
 sg13g2_decap_8 FILLER_37_280 ();
 sg13g2_decap_8 FILLER_37_287 ();
 sg13g2_fill_2 FILLER_37_309 ();
 sg13g2_fill_1 FILLER_37_316 ();
 sg13g2_fill_2 FILLER_37_322 ();
 sg13g2_fill_2 FILLER_37_356 ();
 sg13g2_fill_1 FILLER_37_362 ();
 sg13g2_fill_2 FILLER_37_377 ();
 sg13g2_fill_1 FILLER_37_379 ();
 sg13g2_fill_2 FILLER_37_427 ();
 sg13g2_fill_1 FILLER_37_429 ();
 sg13g2_fill_2 FILLER_38_0 ();
 sg13g2_decap_4 FILLER_38_28 ();
 sg13g2_fill_1 FILLER_38_32 ();
 sg13g2_decap_4 FILLER_38_64 ();
 sg13g2_fill_2 FILLER_38_68 ();
 sg13g2_decap_8 FILLER_38_284 ();
 sg13g2_decap_4 FILLER_38_291 ();
 sg13g2_fill_1 FILLER_38_295 ();
 sg13g2_decap_8 FILLER_38_306 ();
 sg13g2_fill_2 FILLER_38_313 ();
 sg13g2_fill_1 FILLER_38_315 ();
 sg13g2_decap_4 FILLER_38_323 ();
 sg13g2_fill_1 FILLER_38_327 ();
 sg13g2_decap_8 FILLER_38_338 ();
 sg13g2_decap_8 FILLER_38_345 ();
 sg13g2_fill_1 FILLER_38_352 ();
 sg13g2_decap_8 FILLER_38_358 ();
 sg13g2_decap_8 FILLER_38_365 ();
 sg13g2_decap_8 FILLER_38_372 ();
 sg13g2_fill_2 FILLER_38_379 ();
 sg13g2_decap_4 FILLER_38_386 ();
 sg13g2_fill_2 FILLER_38_390 ();
 sg13g2_fill_2 FILLER_38_404 ();
 sg13g2_fill_1 FILLER_38_406 ();
 sg13g2_decap_8 FILLER_38_411 ();
 sg13g2_fill_2 FILLER_38_418 ();
 sg13g2_decap_4 FILLER_38_425 ();
 sg13g2_fill_1 FILLER_38_429 ();
endmodule
