module tt_um_autosel (clk,
    ena,
    rst_n,
    ui_in,
    uio_in,
    uio_oe,
    uio_out,
    uo_out);
 input clk;
 input ena;
 input rst_n;
 input [7:0] ui_in;
 input [7:0] uio_in;
 output [7:0] uio_oe;
 output [7:0] uio_out;
 output [7:0] uo_out;

 wire _0000_;
 wire _0001_;
 wire _0002_;
 wire _0003_;
 wire _0004_;
 wire _0005_;
 wire _0006_;
 wire _0007_;
 wire _0008_;
 wire _0009_;
 wire _0010_;
 wire _0011_;
 wire _0012_;
 wire _0013_;
 wire _0014_;
 wire _0015_;
 wire _0016_;
 wire _0017_;
 wire _0018_;
 wire _0019_;
 wire _0020_;
 wire _0021_;
 wire _0022_;
 wire _0023_;
 wire _0024_;
 wire _0025_;
 wire _0026_;
 wire _0027_;
 wire _0028_;
 wire _0029_;
 wire _0030_;
 wire _0031_;
 wire _0032_;
 wire _0033_;
 wire _0034_;
 wire _0035_;
 wire _0036_;
 wire _0037_;
 wire _0038_;
 wire _0039_;
 wire _0040_;
 wire _0041_;
 wire _0042_;
 wire _0043_;
 wire _0044_;
 wire _0045_;
 wire _0046_;
 wire _0047_;
 wire _0048_;
 wire _0049_;
 wire _0050_;
 wire _0051_;
 wire _0052_;
 wire _0053_;
 wire _0054_;
 wire _0055_;
 wire _0056_;
 wire _0057_;
 wire _0058_;
 wire _0059_;
 wire _0060_;
 wire _0061_;
 wire _0062_;
 wire _0063_;
 wire _0064_;
 wire _0065_;
 wire _0066_;
 wire _0067_;
 wire _0068_;
 wire _0069_;
 wire _0070_;
 wire _0071_;
 wire _0072_;
 wire _0073_;
 wire _0074_;
 wire _0075_;
 wire _0076_;
 wire _0077_;
 wire _0078_;
 wire _0079_;
 wire _0080_;
 wire _0081_;
 wire _0082_;
 wire _0083_;
 wire _0084_;
 wire _0085_;
 wire _0086_;
 wire _0087_;
 wire _0088_;
 wire _0089_;
 wire _0090_;
 wire _0091_;
 wire _0092_;
 wire _0093_;
 wire _0094_;
 wire _0095_;
 wire _0096_;
 wire _0097_;
 wire _0098_;
 wire _0099_;
 wire _0100_;
 wire _0101_;
 wire _0102_;
 wire _0103_;
 wire _0104_;
 wire _0105_;
 wire _0106_;
 wire _0107_;
 wire _0108_;
 wire _0109_;
 wire _0110_;
 wire _0111_;
 wire _0112_;
 wire _0113_;
 wire _0114_;
 wire _0115_;
 wire _0116_;
 wire _0117_;
 wire _0118_;
 wire _0119_;
 wire _0120_;
 wire _0121_;
 wire _0122_;
 wire _0123_;
 wire _0124_;
 wire _0125_;
 wire _0126_;
 wire _0127_;
 wire _0128_;
 wire _0129_;
 wire _0130_;
 wire _0131_;
 wire _0132_;
 wire _0133_;
 wire _0134_;
 wire _0135_;
 wire _0136_;
 wire _0137_;
 wire _0138_;
 wire _0139_;
 wire _0140_;
 wire _0141_;
 wire _0142_;
 wire _0143_;
 wire _0144_;
 wire _0145_;
 wire _0146_;
 wire _0147_;
 wire _0148_;
 wire _0149_;
 wire _0150_;
 wire _0151_;
 wire _0152_;
 wire _0153_;
 wire _0154_;
 wire _0155_;
 wire _0156_;
 wire _0157_;
 wire _0158_;
 wire _0159_;
 wire _0160_;
 wire _0161_;
 wire _0162_;
 wire _0163_;
 wire _0164_;
 wire _0165_;
 wire _0166_;
 wire _0167_;
 wire _0168_;
 wire _0169_;
 wire _0170_;
 wire _0171_;
 wire _0172_;
 wire _0173_;
 wire _0174_;
 wire _0175_;
 wire _0176_;
 wire _0177_;
 wire _0178_;
 wire _0179_;
 wire _0180_;
 wire _0181_;
 wire _0182_;
 wire _0183_;
 wire _0184_;
 wire _0185_;
 wire _0186_;
 wire _0187_;
 wire _0188_;
 wire _0189_;
 wire _0190_;
 wire _0191_;
 wire _0192_;
 wire _0193_;
 wire _0194_;
 wire _0195_;
 wire _0196_;
 wire _0197_;
 wire _0198_;
 wire _0199_;
 wire _0200_;
 wire _0201_;
 wire _0202_;
 wire _0203_;
 wire _0204_;
 wire _0205_;
 wire _0206_;
 wire _0207_;
 wire _0208_;
 wire _0209_;
 wire _0210_;
 wire _0211_;
 wire _0212_;
 wire _0213_;
 wire _0214_;
 wire _0215_;
 wire _0216_;
 wire _0217_;
 wire _0218_;
 wire _0219_;
 wire _0220_;
 wire _0221_;
 wire _0222_;
 wire _0223_;
 wire _0224_;
 wire _0225_;
 wire _0226_;
 wire _0227_;
 wire _0228_;
 wire _0229_;
 wire _0230_;
 wire _0231_;
 wire _0232_;
 wire _0233_;
 wire _0234_;
 wire _0235_;
 wire _0236_;
 wire _0237_;
 wire _0238_;
 wire _0239_;
 wire _0240_;
 wire _0241_;
 wire _0242_;
 wire _0243_;
 wire _0244_;
 wire _0245_;
 wire _0246_;
 wire _0247_;
 wire _0248_;
 wire _0249_;
 wire _0250_;
 wire _0251_;
 wire _0252_;
 wire _0253_;
 wire _0254_;
 wire _0255_;
 wire _0256_;
 wire _0257_;
 wire _0258_;
 wire _0259_;
 wire _0260_;
 wire _0261_;
 wire _0262_;
 wire _0263_;
 wire _0264_;
 wire _0265_;
 wire _0266_;
 wire _0267_;
 wire _0268_;
 wire _0269_;
 wire _0270_;
 wire _0271_;
 wire _0272_;
 wire _0273_;
 wire _0274_;
 wire _0275_;
 wire _0276_;
 wire _0277_;
 wire _0278_;
 wire _0279_;
 wire _0280_;
 wire _0281_;
 wire _0282_;
 wire _0283_;
 wire _0284_;
 wire _0285_;
 wire _0286_;
 wire _0287_;
 wire _0288_;
 wire _0289_;
 wire _0290_;
 wire _0291_;
 wire _0292_;
 wire _0293_;
 wire _0294_;
 wire _0295_;
 wire _0296_;
 wire _0297_;
 wire _0298_;
 wire _0299_;
 wire _0300_;
 wire _0301_;
 wire _0302_;
 wire _0303_;
 wire _0304_;
 wire _0305_;
 wire _0306_;
 wire _0307_;
 wire _0308_;
 wire _0309_;
 wire _0310_;
 wire _0311_;
 wire _0312_;
 wire _0313_;
 wire _0314_;
 wire _0315_;
 wire _0316_;
 wire _0317_;
 wire _0318_;
 wire _0319_;
 wire _0320_;
 wire _0321_;
 wire _0322_;
 wire _0323_;
 wire _0324_;
 wire _0325_;
 wire _0326_;
 wire _0327_;
 wire _0328_;
 wire _0329_;
 wire _0330_;
 wire _0331_;
 wire _0332_;
 wire _0333_;
 wire _0334_;
 wire _0335_;
 wire _0336_;
 wire _0337_;
 wire _0338_;
 wire _0339_;
 wire _0340_;
 wire _0341_;
 wire _0342_;
 wire _0343_;
 wire _0344_;
 wire _0345_;
 wire _0346_;
 wire _0347_;
 wire _0348_;
 wire _0349_;
 wire _0350_;
 wire _0351_;
 wire _0352_;
 wire _0353_;
 wire _0354_;
 wire _0355_;
 wire _0356_;
 wire _0357_;
 wire _0358_;
 wire _0359_;
 wire _0360_;
 wire _0361_;
 wire _0362_;
 wire _0363_;
 wire _0364_;
 wire _0365_;
 wire _0366_;
 wire _0367_;
 wire _0368_;
 wire _0369_;
 wire _0370_;
 wire _0371_;
 wire _0372_;
 wire _0373_;
 wire _0374_;
 wire _0375_;
 wire _0376_;
 wire _0377_;
 wire _0378_;
 wire _0379_;
 wire _0380_;
 wire _0381_;
 wire _0382_;
 wire _0383_;
 wire _0384_;
 wire _0385_;
 wire _0386_;
 wire _0387_;
 wire _0388_;
 wire _0389_;
 wire _0390_;
 wire _0391_;
 wire _0392_;
 wire _0393_;
 wire _0394_;
 wire _0395_;
 wire _0396_;
 wire _0397_;
 wire _0398_;
 wire _0399_;
 wire _0400_;
 wire _0401_;
 wire _0402_;
 wire _0403_;
 wire _0404_;
 wire _0405_;
 wire _0406_;
 wire _0407_;
 wire _0408_;
 wire _0409_;
 wire _0410_;
 wire _0411_;
 wire _0412_;
 wire _0413_;
 wire _0414_;
 wire _0415_;
 wire _0416_;
 wire _0417_;
 wire _0418_;
 wire _0419_;
 wire _0420_;
 wire _0421_;
 wire _0422_;
 wire _0423_;
 wire _0424_;
 wire _0425_;
 wire _0426_;
 wire _0427_;
 wire _0428_;
 wire _0429_;
 wire _0430_;
 wire _0431_;
 wire _0432_;
 wire _0433_;
 wire _0434_;
 wire _0435_;
 wire _0436_;
 wire _0437_;
 wire _0438_;
 wire _0439_;
 wire _0440_;
 wire _0441_;
 wire _0442_;
 wire _0443_;
 wire _0444_;
 wire _0445_;
 wire _0446_;
 wire _0447_;
 wire _0448_;
 wire _0449_;
 wire _0450_;
 wire _0451_;
 wire _0452_;
 wire _0453_;
 wire _0454_;
 wire _0455_;
 wire _0456_;
 wire _0457_;
 wire _0458_;
 wire _0459_;
 wire _0460_;
 wire _0461_;
 wire _0462_;
 wire _0463_;
 wire _0464_;
 wire _0465_;
 wire _0466_;
 wire _0467_;
 wire _0468_;
 wire _0469_;
 wire _0470_;
 wire _0471_;
 wire _0472_;
 wire _0473_;
 wire _0474_;
 wire _0475_;
 wire _0476_;
 wire _0477_;
 wire _0478_;
 wire _0479_;
 wire _0480_;
 wire _0481_;
 wire _0482_;
 wire _0483_;
 wire _0484_;
 wire _0485_;
 wire _0486_;
 wire _0487_;
 wire _0488_;
 wire _0489_;
 wire _0490_;
 wire _0491_;
 wire _0492_;
 wire _0493_;
 wire _0494_;
 wire _0495_;
 wire _0496_;
 wire _0497_;
 wire _0498_;
 wire _0499_;
 wire _0500_;
 wire _0501_;
 wire _0502_;
 wire _0503_;
 wire _0504_;
 wire _0505_;
 wire _0506_;
 wire _0507_;
 wire _0508_;
 wire _0509_;
 wire _0510_;
 wire _0511_;
 wire _0512_;
 wire _0513_;
 wire _0514_;
 wire _0515_;
 wire _0516_;
 wire _0517_;
 wire _0518_;
 wire _0519_;
 wire _0520_;
 wire _0521_;
 wire _0522_;
 wire _0523_;
 wire _0524_;
 wire _0525_;
 wire _0526_;
 wire _0527_;
 wire _0528_;
 wire _0529_;
 wire _0530_;
 wire _0531_;
 wire _0532_;
 wire _0533_;
 wire _0534_;
 wire _0535_;
 wire _0536_;
 wire _0537_;
 wire _0538_;
 wire _0539_;
 wire _0540_;
 wire _0541_;
 wire _0542_;
 wire _0543_;
 wire _0544_;
 wire _0545_;
 wire _0546_;
 wire _0547_;
 wire _0548_;
 wire _0549_;
 wire _0550_;
 wire _0551_;
 wire _0552_;
 wire _0553_;
 wire _0554_;
 wire _0555_;
 wire _0556_;
 wire _0557_;
 wire _0558_;
 wire _0559_;
 wire _0560_;
 wire _0561_;
 wire _0562_;
 wire _0563_;
 wire _0564_;
 wire _0565_;
 wire _0566_;
 wire _0567_;
 wire _0568_;
 wire _0569_;
 wire _0570_;
 wire _0571_;
 wire _0572_;
 wire _0573_;
 wire _0574_;
 wire _0575_;
 wire _0576_;
 wire _0577_;
 wire _0578_;
 wire _0579_;
 wire _0580_;
 wire _0581_;
 wire _0582_;
 wire _0583_;
 wire _0584_;
 wire _0585_;
 wire _0586_;
 wire _0587_;
 wire _0588_;
 wire _0589_;
 wire _0590_;
 wire _0591_;
 wire _0592_;
 wire _0593_;
 wire _0594_;
 wire _0595_;
 wire _0596_;
 wire _0597_;
 wire _0598_;
 wire _0599_;
 wire _0600_;
 wire _0601_;
 wire _0602_;
 wire _0603_;
 wire _0604_;
 wire _0605_;
 wire _0606_;
 wire _0607_;
 wire _0608_;
 wire _0609_;
 wire _0610_;
 wire _0611_;
 wire _0612_;
 wire _0613_;
 wire _0614_;
 wire _0615_;
 wire _0616_;
 wire _0617_;
 wire _0618_;
 wire _0619_;
 wire _0620_;
 wire _0621_;
 wire _0622_;
 wire _0623_;
 wire _0624_;
 wire _0625_;
 wire _0626_;
 wire _0627_;
 wire _0628_;
 wire _0629_;
 wire _0630_;
 wire _0631_;
 wire _0632_;
 wire _0633_;
 wire _0634_;
 wire _0635_;
 wire _0636_;
 wire _0637_;
 wire _0638_;
 wire _0639_;
 wire _0640_;
 wire _0641_;
 wire _0642_;
 wire _0643_;
 wire _0644_;
 wire _0645_;
 wire _0646_;
 wire _0647_;
 wire _0648_;
 wire _0649_;
 wire _0650_;
 wire _0651_;
 wire _0652_;
 wire _0653_;
 wire _0654_;
 wire _0655_;
 wire _0656_;
 wire _0657_;
 wire _0658_;
 wire _0659_;
 wire _0660_;
 wire _0661_;
 wire _0662_;
 wire _0663_;
 wire _0664_;
 wire _0665_;
 wire _0666_;
 wire _0667_;
 wire _0668_;
 wire _0669_;
 wire _0670_;
 wire _0671_;
 wire _0672_;
 wire _0673_;
 wire _0674_;
 wire _0675_;
 wire _0676_;
 wire _0677_;
 wire _0678_;
 wire _0679_;
 wire _0680_;
 wire _0681_;
 wire _0682_;
 wire _0683_;
 wire _0684_;
 wire _0685_;
 wire _0686_;
 wire _0687_;
 wire _0688_;
 wire _0689_;
 wire _0690_;
 wire _0691_;
 wire _0692_;
 wire _0693_;
 wire _0694_;
 wire _0695_;
 wire _0696_;
 wire _0697_;
 wire _0698_;
 wire _0699_;
 wire _0700_;
 wire _0701_;
 wire _0702_;
 wire _0703_;
 wire _0704_;
 wire _0705_;
 wire _0706_;
 wire _0707_;
 wire _0708_;
 wire _0709_;
 wire _0710_;
 wire _0711_;
 wire _0712_;
 wire _0713_;
 wire _0714_;
 wire _0715_;
 wire _0716_;
 wire _0717_;
 wire _0718_;
 wire _0719_;
 wire _0720_;
 wire _0721_;
 wire _0722_;
 wire _0723_;
 wire _0724_;
 wire _0725_;
 wire _0726_;
 wire _0727_;
 wire _0728_;
 wire _0729_;
 wire _0730_;
 wire _0731_;
 wire _0732_;
 wire _0733_;
 wire _0734_;
 wire _0735_;
 wire _0736_;
 wire _0737_;
 wire _0738_;
 wire _0739_;
 wire _0740_;
 wire _0741_;
 wire _0742_;
 wire _0743_;
 wire _0744_;
 wire _0745_;
 wire _0746_;
 wire _0747_;
 wire _0748_;
 wire _0749_;
 wire _0750_;
 wire _0751_;
 wire _0752_;
 wire _0753_;
 wire _0754_;
 wire _0755_;
 wire _0756_;
 wire _0757_;
 wire _0758_;
 wire _0759_;
 wire _0760_;
 wire _0761_;
 wire _0762_;
 wire _0763_;
 wire _0764_;
 wire _0765_;
 wire _0766_;
 wire _0767_;
 wire _0768_;
 wire _0769_;
 wire _0770_;
 wire _0771_;
 wire _0772_;
 wire _0773_;
 wire _0774_;
 wire _0775_;
 wire _0776_;
 wire _0777_;
 wire _0778_;
 wire _0779_;
 wire _0780_;
 wire _0781_;
 wire _0782_;
 wire _0783_;
 wire _0784_;
 wire _0785_;
 wire _0786_;
 wire _0787_;
 wire _0788_;
 wire _0789_;
 wire _0790_;
 wire _0791_;
 wire _0792_;
 wire _0793_;
 wire _0794_;
 wire _0795_;
 wire _0796_;
 wire _0797_;
 wire _0798_;
 wire _0799_;
 wire _0800_;
 wire _0801_;
 wire _0802_;
 wire _0803_;
 wire _0804_;
 wire _0805_;
 wire _0806_;
 wire _0807_;
 wire _0808_;
 wire _0809_;
 wire _0810_;
 wire _0811_;
 wire _0812_;
 wire _0813_;
 wire _0814_;
 wire _0815_;
 wire _0816_;
 wire _0817_;
 wire _0818_;
 wire _0819_;
 wire _0820_;
 wire _0821_;
 wire _0822_;
 wire _0823_;
 wire _0824_;
 wire _0825_;
 wire _0826_;
 wire _0827_;
 wire _0828_;
 wire _0829_;
 wire _0830_;
 wire _0831_;
 wire _0832_;
 wire _0833_;
 wire _0834_;
 wire _0835_;
 wire _0836_;
 wire _0837_;
 wire _0838_;
 wire _0839_;
 wire _0840_;
 wire _0841_;
 wire _0842_;
 wire _0843_;
 wire _0844_;
 wire _0845_;
 wire _0846_;
 wire _0847_;
 wire _0848_;
 wire _0849_;
 wire _0850_;
 wire _0851_;
 wire _0852_;
 wire _0853_;
 wire _0854_;
 wire _0855_;
 wire _0856_;
 wire _0857_;
 wire _0858_;
 wire _0859_;
 wire _0860_;
 wire _0861_;
 wire _0862_;
 wire _0863_;
 wire _0864_;
 wire _0865_;
 wire _0866_;
 wire _0867_;
 wire _0868_;
 wire _0869_;
 wire _0870_;
 wire _0871_;
 wire _0872_;
 wire _0873_;
 wire _0874_;
 wire _0875_;
 wire _0876_;
 wire _0877_;
 wire _0878_;
 wire _0879_;
 wire _0880_;
 wire _0881_;
 wire _0882_;
 wire _0883_;
 wire _0884_;
 wire _0885_;
 wire _0886_;
 wire _0887_;
 wire _0888_;
 wire _0889_;
 wire _0890_;
 wire _0891_;
 wire _0892_;
 wire _0893_;
 wire _0894_;
 wire _0895_;
 wire _0896_;
 wire _0897_;
 wire _0898_;
 wire _0899_;
 wire _0900_;
 wire _0901_;
 wire _0902_;
 wire _0903_;
 wire _0904_;
 wire _0905_;
 wire _0906_;
 wire _0907_;
 wire _0908_;
 wire _0909_;
 wire _0910_;
 wire _0911_;
 wire _0912_;
 wire _0913_;
 wire _0914_;
 wire _0915_;
 wire _0916_;
 wire _0917_;
 wire _0918_;
 wire _0919_;
 wire _0920_;
 wire _0921_;
 wire _0922_;
 wire _0923_;
 wire _0924_;
 wire _0925_;
 wire _0926_;
 wire _0927_;
 wire _0928_;
 wire _0929_;
 wire _0930_;
 wire _0931_;
 wire _0932_;
 wire _0933_;
 wire _0934_;
 wire _0935_;
 wire _0936_;
 wire _0937_;
 wire _0938_;
 wire _0939_;
 wire _0940_;
 wire _0941_;
 wire _0942_;
 wire _0943_;
 wire _0944_;
 wire _0945_;
 wire _0946_;
 wire _0947_;
 wire _0948_;
 wire _0949_;
 wire _0950_;
 wire _0951_;
 wire _0952_;
 wire _0953_;
 wire _0954_;
 wire _0955_;
 wire _0956_;
 wire _0957_;
 wire _0958_;
 wire _0959_;
 wire _0960_;
 wire _0961_;
 wire _0962_;
 wire _0963_;
 wire _0964_;
 wire _0965_;
 wire _0966_;
 wire _0967_;
 wire _0968_;
 wire _0969_;
 wire _0970_;
 wire _0971_;
 wire _0972_;
 wire _0973_;
 wire _0974_;
 wire _0975_;
 wire _0976_;
 wire _0977_;
 wire _0978_;
 wire _0979_;
 wire _0980_;
 wire _0981_;
 wire _0982_;
 wire _0983_;
 wire _0984_;
 wire _0985_;
 wire _0986_;
 wire _0987_;
 wire _0988_;
 wire _0989_;
 wire _0990_;
 wire _0991_;
 wire _0992_;
 wire _0993_;
 wire _0994_;
 wire _0995_;
 wire _0996_;
 wire _0997_;
 wire _0998_;
 wire _0999_;
 wire _1000_;
 wire _1001_;
 wire _1002_;
 wire _1003_;
 wire _1004_;
 wire _1005_;
 wire _1006_;
 wire _1007_;
 wire _1008_;
 wire _1009_;
 wire _1010_;
 wire _1011_;
 wire _1012_;
 wire _1013_;
 wire _1014_;
 wire _1015_;
 wire _1016_;
 wire _1017_;
 wire _1018_;
 wire _1019_;
 wire _1020_;
 wire _1021_;
 wire _1022_;
 wire _1023_;
 wire _1024_;
 wire _1025_;
 wire _1026_;
 wire _1027_;
 wire _1028_;
 wire _1029_;
 wire _1030_;
 wire _1031_;
 wire _1032_;
 wire _1033_;
 wire _1034_;
 wire _1035_;
 wire _1036_;
 wire _1037_;
 wire _1038_;
 wire _1039_;
 wire _1040_;
 wire _1041_;
 wire _1042_;
 wire _1043_;
 wire _1044_;
 wire _1045_;
 wire _1046_;
 wire _1047_;
 wire _1048_;
 wire _1049_;
 wire _1050_;
 wire _1051_;
 wire _1052_;
 wire _1053_;
 wire _1054_;
 wire _1055_;
 wire _1056_;
 wire _1057_;
 wire _1058_;
 wire _1059_;
 wire _1060_;
 wire _1061_;
 wire _1062_;
 wire _1063_;
 wire _1064_;
 wire _1065_;
 wire _1066_;
 wire _1067_;
 wire _1068_;
 wire _1069_;
 wire _1070_;
 wire _1071_;
 wire _1072_;
 wire _1073_;
 wire _1074_;
 wire _1075_;
 wire _1076_;
 wire _1077_;
 wire _1078_;
 wire _1079_;
 wire _1080_;
 wire _1081_;
 wire _1082_;
 wire _1083_;
 wire _1084_;
 wire _1085_;
 wire _1086_;
 wire _1087_;
 wire _1088_;
 wire _1089_;
 wire _1090_;
 wire _1091_;
 wire _1092_;
 wire _1093_;
 wire _1094_;
 wire _1095_;
 wire _1096_;
 wire _1097_;
 wire _1098_;
 wire _1099_;
 wire _1100_;
 wire _1101_;
 wire _1102_;
 wire _1103_;
 wire _1104_;
 wire _1105_;
 wire _1106_;
 wire _1107_;
 wire _1108_;
 wire _1109_;
 wire _1110_;
 wire _1111_;
 wire _1112_;
 wire _1113_;
 wire _1114_;
 wire _1115_;
 wire _1116_;
 wire _1117_;
 wire _1118_;
 wire _1119_;
 wire _1120_;
 wire _1121_;
 wire _1122_;
 wire _1123_;
 wire _1124_;
 wire _1125_;
 wire _1126_;
 wire _1127_;
 wire _1128_;
 wire _1129_;
 wire _1130_;
 wire _1131_;
 wire _1132_;
 wire _1133_;
 wire _1134_;
 wire _1135_;
 wire _1136_;
 wire _1137_;
 wire _1138_;
 wire _1139_;
 wire _1140_;
 wire _1141_;
 wire _1142_;
 wire _1143_;
 wire _1144_;
 wire _1145_;
 wire _1146_;
 wire _1147_;
 wire _1148_;
 wire _1149_;
 wire _1150_;
 wire clknet_0_clk;
 wire net81;
 wire \autosel.addr_counter[0] ;
 wire \autosel.addr_counter[1] ;
 wire \autosel.addr_counter[2] ;
 wire \autosel.addr_counter[3] ;
 wire \autosel.addr_counter[4] ;
 wire \autosel.addr_counter[5] ;
 wire \autosel.addr_counter[6] ;
 wire \autosel.addr_counter[7] ;
 wire \autosel.addr_counter[8] ;
 wire \autosel.addr_counter[9] ;
 wire \autosel.ctrl_ena ;
 wire \autosel.ctrl_sel_inc ;
 wire \autosel.ctrl_sel_rst_n ;
 wire \autosel.eeprom_busy ;
 wire \autosel.eeprom_data[0] ;
 wire \autosel.eeprom_data[10] ;
 wire \autosel.eeprom_data[11] ;
 wire \autosel.eeprom_data[12] ;
 wire \autosel.eeprom_data[13] ;
 wire \autosel.eeprom_data[14] ;
 wire \autosel.eeprom_data[15] ;
 wire \autosel.eeprom_data[1] ;
 wire \autosel.eeprom_data[2] ;
 wire \autosel.eeprom_data[3] ;
 wire \autosel.eeprom_data[4] ;
 wire \autosel.eeprom_data[5] ;
 wire \autosel.eeprom_data[6] ;
 wire \autosel.eeprom_data[7] ;
 wire \autosel.eeprom_data[8] ;
 wire \autosel.eeprom_data[9] ;
 wire \autosel.i2c.data_out_hi[0] ;
 wire \autosel.i2c.data_out_hi[1] ;
 wire \autosel.i2c.data_out_hi[2] ;
 wire \autosel.i2c.data_out_hi[3] ;
 wire \autosel.i2c.data_out_hi[4] ;
 wire \autosel.i2c.data_out_hi[5] ;
 wire \autosel.i2c.data_out_hi[6] ;
 wire \autosel.i2c.data_out_hi[7] ;
 wire \autosel.i2c.i2c.addr_reg[4] ;
 wire \autosel.i2c.i2c.bit_count_reg[0] ;
 wire \autosel.i2c.i2c.bit_count_reg[1] ;
 wire \autosel.i2c.i2c.bit_count_reg[2] ;
 wire \autosel.i2c.i2c.bit_count_reg[3] ;
 wire \autosel.i2c.i2c.bus_active_reg ;
 wire \autosel.i2c.i2c.busy_reg ;
 wire \autosel.i2c.i2c.data_reg[0] ;
 wire \autosel.i2c.i2c.data_reg[1] ;
 wire \autosel.i2c.i2c.data_reg[2] ;
 wire \autosel.i2c.i2c.data_reg[3] ;
 wire \autosel.i2c.i2c.data_reg[4] ;
 wire \autosel.i2c.i2c.data_reg[5] ;
 wire \autosel.i2c.i2c.data_reg[6] ;
 wire \autosel.i2c.i2c.data_reg[7] ;
 wire \autosel.i2c.i2c.delay_reg[0] ;
 wire \autosel.i2c.i2c.delay_reg[10] ;
 wire \autosel.i2c.i2c.delay_reg[11] ;
 wire \autosel.i2c.i2c.delay_reg[12] ;
 wire \autosel.i2c.i2c.delay_reg[13] ;
 wire \autosel.i2c.i2c.delay_reg[14] ;
 wire \autosel.i2c.i2c.delay_reg[15] ;
 wire \autosel.i2c.i2c.delay_reg[1] ;
 wire \autosel.i2c.i2c.delay_reg[2] ;
 wire \autosel.i2c.i2c.delay_reg[3] ;
 wire \autosel.i2c.i2c.delay_reg[4] ;
 wire \autosel.i2c.i2c.delay_reg[5] ;
 wire \autosel.i2c.i2c.delay_reg[6] ;
 wire \autosel.i2c.i2c.delay_reg[7] ;
 wire \autosel.i2c.i2c.delay_reg[8] ;
 wire \autosel.i2c.i2c.delay_reg[9] ;
 wire \autosel.i2c.i2c.delay_scl_reg ;
 wire \autosel.i2c.i2c.delay_sda_reg ;
 wire \autosel.i2c.i2c.last_sda_i_reg ;
 wire \autosel.i2c.i2c.m_axis_data_tdata_reg[0] ;
 wire \autosel.i2c.i2c.m_axis_data_tdata_reg[1] ;
 wire \autosel.i2c.i2c.m_axis_data_tdata_reg[2] ;
 wire \autosel.i2c.i2c.m_axis_data_tdata_reg[3] ;
 wire \autosel.i2c.i2c.m_axis_data_tdata_reg[4] ;
 wire \autosel.i2c.i2c.m_axis_data_tdata_reg[5] ;
 wire \autosel.i2c.i2c.m_axis_data_tdata_reg[6] ;
 wire \autosel.i2c.i2c.m_axis_data_tdata_reg[7] ;
 wire \autosel.i2c.i2c.m_axis_data_tvalid_reg ;
 wire \autosel.i2c.i2c.missed_ack_reg ;
 wire \autosel.i2c.i2c.mode_read_reg ;
 wire \autosel.i2c.i2c.mode_stop_reg ;
 wire \autosel.i2c.i2c.phy_rx_data_reg ;
 wire \autosel.i2c.i2c.phy_state_reg[0] ;
 wire \autosel.i2c.i2c.phy_state_reg[1] ;
 wire \autosel.i2c.i2c.phy_state_reg[2] ;
 wire \autosel.i2c.i2c.phy_state_reg[3] ;
 wire \autosel.i2c.i2c.s_axis_cmd_ready_reg ;
 wire \autosel.i2c.i2c.s_axis_data_tready_reg ;
 wire \autosel.i2c.i2c.scl_i_reg ;
 wire \autosel.i2c.i2c.scl_o_reg ;
 wire \autosel.i2c.i2c.sda_i_reg ;
 wire \autosel.i2c.i2c.sda_o_reg ;
 wire \autosel.i2c.i2c.state_reg[0] ;
 wire \autosel.i2c.i2c.state_reg[1] ;
 wire \autosel.i2c.i2c.state_reg[2] ;
 wire \autosel.i2c.i2c.state_reg[3] ;
 wire \autosel.i2c.start ;
 wire \autosel.i2c.state[0] ;
 wire \autosel.i2c.state[1] ;
 wire \autosel.i2c.state[2] ;
 wire \autosel.scl_oe ;
 wire \autosel.sda_oe ;
 wire \autosel.state[1] ;
 wire \autosel.state[2] ;
 wire \debug_out.counter[0] ;
 wire \debug_out.counter[10] ;
 wire \debug_out.counter[11] ;
 wire \debug_out.counter[12] ;
 wire \debug_out.counter[13] ;
 wire \debug_out.counter[14] ;
 wire \debug_out.counter[15] ;
 wire \debug_out.counter[16] ;
 wire \debug_out.counter[17] ;
 wire \debug_out.counter[18] ;
 wire \debug_out.counter[19] ;
 wire \debug_out.counter[1] ;
 wire \debug_out.counter[20] ;
 wire \debug_out.counter[21] ;
 wire \debug_out.counter[22] ;
 wire \debug_out.counter[23] ;
 wire \debug_out.counter[24] ;
 wire \debug_out.counter[25] ;
 wire \debug_out.counter[26] ;
 wire \debug_out.counter[27] ;
 wire \debug_out.counter[28] ;
 wire \debug_out.counter[29] ;
 wire \debug_out.counter[2] ;
 wire \debug_out.counter[30] ;
 wire \debug_out.counter[31] ;
 wire \debug_out.counter[3] ;
 wire \debug_out.counter[4] ;
 wire \debug_out.counter[5] ;
 wire \debug_out.counter[6] ;
 wire \debug_out.counter[7] ;
 wire \debug_out.counter[8] ;
 wire \debug_out.counter[9] ;
 wire \debug_out.send_index[0] ;
 wire \debug_out.send_index[1] ;
 wire \debug_out.send_index[2] ;
 wire \debug_out.tx_byte[0] ;
 wire \debug_out.tx_byte[1] ;
 wire \debug_out.tx_byte[2] ;
 wire \debug_out.tx_byte[3] ;
 wire \debug_out.tx_byte[4] ;
 wire \debug_out.tx_byte[6] ;
 wire \debug_out.tx_ready ;
 wire \debug_out.tx_valid ;
 wire \debug_out.uart_tx ;
 wire \debug_out.uart_tx_inst.bit_cnt[0] ;
 wire \debug_out.uart_tx_inst.bit_cnt[1] ;
 wire \debug_out.uart_tx_inst.bit_cnt[2] ;
 wire \debug_out.uart_tx_inst.cycle_cnt[0] ;
 wire \debug_out.uart_tx_inst.cycle_cnt[10] ;
 wire \debug_out.uart_tx_inst.cycle_cnt[11] ;
 wire \debug_out.uart_tx_inst.cycle_cnt[12] ;
 wire \debug_out.uart_tx_inst.cycle_cnt[13] ;
 wire \debug_out.uart_tx_inst.cycle_cnt[14] ;
 wire \debug_out.uart_tx_inst.cycle_cnt[15] ;
 wire \debug_out.uart_tx_inst.cycle_cnt[1] ;
 wire \debug_out.uart_tx_inst.cycle_cnt[2] ;
 wire \debug_out.uart_tx_inst.cycle_cnt[3] ;
 wire \debug_out.uart_tx_inst.cycle_cnt[4] ;
 wire \debug_out.uart_tx_inst.cycle_cnt[5] ;
 wire \debug_out.uart_tx_inst.cycle_cnt[6] ;
 wire \debug_out.uart_tx_inst.cycle_cnt[7] ;
 wire \debug_out.uart_tx_inst.cycle_cnt[8] ;
 wire \debug_out.uart_tx_inst.cycle_cnt[9] ;
 wire \debug_out.uart_tx_inst.next_state[1] ;
 wire \debug_out.uart_tx_inst.next_state[2] ;
 wire \debug_out.uart_tx_inst.state[0] ;
 wire \debug_out.uart_tx_inst.state[1] ;
 wire \debug_out.uart_tx_inst.state[2] ;
 wire \debug_out.uart_tx_inst.tx_data_latch[0] ;
 wire \debug_out.uart_tx_inst.tx_data_latch[1] ;
 wire \debug_out.uart_tx_inst.tx_data_latch[2] ;
 wire \debug_out.uart_tx_inst.tx_data_latch[3] ;
 wire \debug_out.uart_tx_inst.tx_data_latch[4] ;
 wire \debug_out.uart_tx_inst.tx_data_latch[6] ;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net180;
 wire net181;
 wire net182;
 wire net183;
 wire net184;
 wire net185;
 wire net186;
 wire net187;
 wire net188;
 wire net189;
 wire net190;
 wire net191;
 wire net192;
 wire net193;
 wire net194;
 wire net195;
 wire net196;
 wire net197;
 wire net198;
 wire net199;
 wire net200;
 wire net201;
 wire net202;
 wire net203;
 wire net204;
 wire net205;
 wire net206;
 wire net207;
 wire clknet_4_0_0_clk;
 wire clknet_4_1_0_clk;
 wire clknet_4_2_0_clk;
 wire clknet_4_3_0_clk;
 wire clknet_4_4_0_clk;
 wire clknet_4_5_0_clk;
 wire clknet_4_6_0_clk;
 wire clknet_4_7_0_clk;
 wire clknet_4_8_0_clk;
 wire clknet_4_9_0_clk;
 wire clknet_4_10_0_clk;
 wire clknet_4_11_0_clk;
 wire clknet_4_12_0_clk;
 wire clknet_4_13_0_clk;
 wire clknet_4_14_0_clk;
 wire clknet_4_15_0_clk;
 wire clknet_5_0__leaf_clk;
 wire clknet_5_1__leaf_clk;
 wire clknet_5_2__leaf_clk;
 wire clknet_5_3__leaf_clk;
 wire clknet_5_4__leaf_clk;
 wire clknet_5_5__leaf_clk;
 wire clknet_5_6__leaf_clk;
 wire clknet_5_7__leaf_clk;
 wire clknet_5_8__leaf_clk;
 wire clknet_5_9__leaf_clk;
 wire clknet_5_10__leaf_clk;
 wire clknet_5_11__leaf_clk;
 wire clknet_5_12__leaf_clk;
 wire clknet_5_13__leaf_clk;
 wire clknet_5_14__leaf_clk;
 wire clknet_5_15__leaf_clk;
 wire clknet_5_16__leaf_clk;
 wire clknet_5_17__leaf_clk;
 wire clknet_5_18__leaf_clk;
 wire clknet_5_19__leaf_clk;
 wire clknet_5_20__leaf_clk;
 wire clknet_5_21__leaf_clk;
 wire clknet_5_22__leaf_clk;
 wire clknet_5_23__leaf_clk;
 wire clknet_5_24__leaf_clk;
 wire clknet_5_25__leaf_clk;
 wire clknet_5_26__leaf_clk;
 wire clknet_5_27__leaf_clk;
 wire clknet_5_28__leaf_clk;
 wire clknet_5_29__leaf_clk;
 wire clknet_5_30__leaf_clk;
 wire clknet_5_31__leaf_clk;

 sg13g2_buf_1 _1153_ (.A(net59),
    .X(_0527_));
 sg13g2_inv_2 _1154_ (.Y(_0528_),
    .A(net55));
 sg13g2_buf_1 _1155_ (.A(_0528_),
    .X(_0000_));
 sg13g2_nor2b_1 _1156_ (.A(\autosel.eeprom_busy ),
    .B_N(\autosel.state[2] ),
    .Y(_0529_));
 sg13g2_buf_1 _1157_ (.A(net55),
    .X(_0530_));
 sg13g2_o21ai_1 _1158_ (.B1(net54),
    .Y(_0531_),
    .A1(\autosel.state[1] ),
    .A2(_0529_));
 sg13g2_inv_1 _1159_ (.Y(_0001_),
    .A(_0531_));
 sg13g2_a21oi_1 _1160_ (.A1(\autosel.eeprom_busy ),
    .A2(\autosel.state[2] ),
    .Y(_0532_),
    .B1(\autosel.i2c.start ));
 sg13g2_nor2_1 _1161_ (.A(net36),
    .B(_0532_),
    .Y(_0002_));
 sg13g2_buf_1 _1162_ (.A(\debug_out.uart_tx_inst.state[0] ),
    .X(_0533_));
 sg13g2_buf_2 _1163_ (.A(\debug_out.uart_tx_inst.cycle_cnt[9] ),
    .X(_0534_));
 sg13g2_nor4_1 _1164_ (.A(\debug_out.uart_tx_inst.cycle_cnt[1] ),
    .B(_0534_),
    .C(\debug_out.uart_tx_inst.cycle_cnt[11] ),
    .D(\debug_out.uart_tx_inst.cycle_cnt[10] ),
    .Y(_0535_));
 sg13g2_nor4_1 _1165_ (.A(\debug_out.uart_tx_inst.cycle_cnt[13] ),
    .B(\debug_out.uart_tx_inst.cycle_cnt[12] ),
    .C(\debug_out.uart_tx_inst.cycle_cnt[15] ),
    .D(\debug_out.uart_tx_inst.cycle_cnt[14] ),
    .Y(_0536_));
 sg13g2_nand2_2 _1166_ (.Y(_0537_),
    .A(_0535_),
    .B(_0536_));
 sg13g2_nor2b_1 _1167_ (.A(\debug_out.uart_tx_inst.cycle_cnt[6] ),
    .B_N(\debug_out.uart_tx_inst.cycle_cnt[7] ),
    .Y(_0538_));
 sg13g2_nor2b_1 _1168_ (.A(\debug_out.uart_tx_inst.cycle_cnt[4] ),
    .B_N(\debug_out.uart_tx_inst.cycle_cnt[5] ),
    .Y(_0539_));
 sg13g2_and2_1 _1169_ (.A(\debug_out.uart_tx_inst.cycle_cnt[3] ),
    .B(\debug_out.uart_tx_inst.cycle_cnt[2] ),
    .X(_0540_));
 sg13g2_buf_1 _1170_ (.A(\debug_out.uart_tx_inst.cycle_cnt[0] ),
    .X(_0541_));
 sg13g2_nor2_1 _1171_ (.A(_0541_),
    .B(\debug_out.uart_tx_inst.cycle_cnt[8] ),
    .Y(_0542_));
 sg13g2_nand4_1 _1172_ (.B(_0539_),
    .C(_0540_),
    .A(_0538_),
    .Y(_0543_),
    .D(_0542_));
 sg13g2_buf_1 _1173_ (.A(_0543_),
    .X(_0544_));
 sg13g2_buf_1 _1174_ (.A(_0033_),
    .X(_0545_));
 sg13g2_inv_1 _1175_ (.Y(_0546_),
    .A(_0545_));
 sg13g2_o21ai_1 _1176_ (.B1(_0546_),
    .Y(_0547_),
    .A1(_0537_),
    .A2(_0544_));
 sg13g2_nand3_1 _1177_ (.B(_0545_),
    .C(\debug_out.tx_valid ),
    .A(net53),
    .Y(_0548_));
 sg13g2_o21ai_1 _1178_ (.B1(_0548_),
    .Y(_0549_),
    .A1(net53),
    .A2(_0547_));
 sg13g2_inv_1 _1179_ (.Y(_0550_),
    .A(\debug_out.uart_tx_inst.state[2] ));
 sg13g2_nand2_1 _1180_ (.Y(_0551_),
    .A(net53),
    .B(_0550_));
 sg13g2_buf_2 _1181_ (.A(\debug_out.uart_tx_inst.bit_cnt[1] ),
    .X(_0552_));
 sg13g2_buf_2 _1182_ (.A(\debug_out.uart_tx_inst.bit_cnt[0] ),
    .X(_0553_));
 sg13g2_nor2_2 _1183_ (.A(_0537_),
    .B(_0544_),
    .Y(_0554_));
 sg13g2_nand4_1 _1184_ (.B(_0553_),
    .C(\debug_out.uart_tx_inst.bit_cnt[2] ),
    .A(_0552_),
    .Y(_0555_),
    .D(_0554_));
 sg13g2_nor2_1 _1185_ (.A(_0533_),
    .B(_0546_),
    .Y(_0556_));
 sg13g2_o21ai_1 _1186_ (.B1(_0556_),
    .Y(_0557_),
    .A1(_0537_),
    .A2(_0544_));
 sg13g2_o21ai_1 _1187_ (.B1(_0557_),
    .Y(_0558_),
    .A1(_0551_),
    .A2(_0555_));
 sg13g2_buf_1 _1188_ (.A(\debug_out.uart_tx_inst.state[1] ),
    .X(_0559_));
 sg13g2_mux2_1 _1189_ (.A0(_0549_),
    .A1(_0558_),
    .S(net52),
    .X(_0045_));
 sg13g2_inv_1 _1190_ (.Y(_0560_),
    .A(net53));
 sg13g2_nor2_1 _1191_ (.A(_0560_),
    .B(\debug_out.uart_tx_inst.state[2] ),
    .Y(_0561_));
 sg13g2_a21o_1 _1192_ (.A2(_0555_),
    .A1(_0561_),
    .B1(_0556_),
    .X(_0562_));
 sg13g2_nand2_1 _1193_ (.Y(_0563_),
    .A(_0545_),
    .B(\debug_out.tx_valid ));
 sg13g2_nand2b_1 _1194_ (.Y(_0564_),
    .B(net53),
    .A_N(net52));
 sg13g2_nor2_2 _1195_ (.A(_0563_),
    .B(_0564_),
    .Y(_0565_));
 sg13g2_a21o_1 _1196_ (.A2(_0562_),
    .A1(net52),
    .B1(_0565_),
    .X(\debug_out.uart_tx_inst.next_state[1] ));
 sg13g2_or3_1 _1197_ (.A(net52),
    .B(net53),
    .C(_0547_),
    .X(_0566_));
 sg13g2_and3_1 _1198_ (.X(_0567_),
    .A(_0552_),
    .B(_0553_),
    .C(\debug_out.uart_tx_inst.bit_cnt[2] ));
 sg13g2_nand4_1 _1199_ (.B(_0554_),
    .C(_0561_),
    .A(net52),
    .Y(_0568_),
    .D(_0567_));
 sg13g2_nand2_1 _1200_ (.Y(\debug_out.uart_tx_inst.next_state[2] ),
    .A(_0566_),
    .B(_0568_));
 sg13g2_a21oi_1 _1201_ (.A1(_0566_),
    .A2(_0568_),
    .Y(_0569_),
    .B1(\debug_out.uart_tx_inst.state[2] ));
 sg13g2_nand2_1 _1202_ (.Y(_0570_),
    .A(\debug_out.uart_tx_inst.state[1] ),
    .B(net53));
 sg13g2_nand2b_1 _1203_ (.Y(_0571_),
    .B(_0563_),
    .A_N(\debug_out.uart_tx_inst.state[1] ));
 sg13g2_o21ai_1 _1204_ (.B1(_0571_),
    .Y(_0572_),
    .A1(_0554_),
    .A2(_0570_));
 sg13g2_nand2_1 _1205_ (.Y(_0573_),
    .A(_0545_),
    .B(_0550_));
 sg13g2_o21ai_1 _1206_ (.B1(_0573_),
    .Y(_0574_),
    .A1(net52),
    .A2(_0547_));
 sg13g2_a22oi_1 _1207_ (.Y(_0575_),
    .B1(_0574_),
    .B2(_0560_),
    .A2(_0572_),
    .A1(_0550_));
 sg13g2_nand2b_1 _1208_ (.Y(_0576_),
    .B(_0545_),
    .A_N(net52));
 sg13g2_nor2_1 _1209_ (.A(_0560_),
    .B(\debug_out.tx_valid ),
    .Y(_0577_));
 sg13g2_nand2_1 _1210_ (.Y(_0578_),
    .A(_0560_),
    .B(_0554_));
 sg13g2_o21ai_1 _1211_ (.B1(_0578_),
    .Y(_0579_),
    .A1(_0576_),
    .A2(_0577_));
 sg13g2_or3_1 _1212_ (.A(_0569_),
    .B(_0575_),
    .C(_0579_),
    .X(_0580_));
 sg13g2_buf_2 _1213_ (.A(_0580_),
    .X(_0581_));
 sg13g2_buf_1 _1214_ (.A(_0581_),
    .X(_0582_));
 sg13g2_nor2_1 _1215_ (.A(_0541_),
    .B(_0582_),
    .Y(_0003_));
 sg13g2_xnor2_1 _1216_ (.Y(_0583_),
    .A(\debug_out.uart_tx_inst.cycle_cnt[1] ),
    .B(_0541_));
 sg13g2_nor2_1 _1217_ (.A(net13),
    .B(_0583_),
    .Y(_0010_));
 sg13g2_nand2_1 _1218_ (.Y(_0584_),
    .A(\debug_out.uart_tx_inst.cycle_cnt[1] ),
    .B(_0541_));
 sg13g2_xor2_1 _1219_ (.B(_0584_),
    .A(\debug_out.uart_tx_inst.cycle_cnt[2] ),
    .X(_0585_));
 sg13g2_nor2_1 _1220_ (.A(net13),
    .B(_0585_),
    .Y(_0011_));
 sg13g2_nand3_1 _1221_ (.B(_0541_),
    .C(\debug_out.uart_tx_inst.cycle_cnt[2] ),
    .A(\debug_out.uart_tx_inst.cycle_cnt[1] ),
    .Y(_0586_));
 sg13g2_xor2_1 _1222_ (.B(_0586_),
    .A(\debug_out.uart_tx_inst.cycle_cnt[3] ),
    .X(_0587_));
 sg13g2_nor2_1 _1223_ (.A(net13),
    .B(_0587_),
    .Y(_0012_));
 sg13g2_and4_1 _1224_ (.A(\debug_out.uart_tx_inst.cycle_cnt[1] ),
    .B(_0541_),
    .C(\debug_out.uart_tx_inst.cycle_cnt[3] ),
    .D(\debug_out.uart_tx_inst.cycle_cnt[2] ),
    .X(_0588_));
 sg13g2_buf_1 _1225_ (.A(_0588_),
    .X(_0589_));
 sg13g2_xnor2_1 _1226_ (.Y(_0590_),
    .A(\debug_out.uart_tx_inst.cycle_cnt[4] ),
    .B(_0589_));
 sg13g2_nor2_1 _1227_ (.A(net13),
    .B(_0590_),
    .Y(_0013_));
 sg13g2_nand2_1 _1228_ (.Y(_0591_),
    .A(\debug_out.uart_tx_inst.cycle_cnt[4] ),
    .B(_0589_));
 sg13g2_xor2_1 _1229_ (.B(_0591_),
    .A(\debug_out.uart_tx_inst.cycle_cnt[5] ),
    .X(_0592_));
 sg13g2_nor2_1 _1230_ (.A(net13),
    .B(_0592_),
    .Y(_0014_));
 sg13g2_nand3_1 _1231_ (.B(\debug_out.uart_tx_inst.cycle_cnt[5] ),
    .C(_0589_),
    .A(\debug_out.uart_tx_inst.cycle_cnt[4] ),
    .Y(_0593_));
 sg13g2_xor2_1 _1232_ (.B(_0593_),
    .A(\debug_out.uart_tx_inst.cycle_cnt[6] ),
    .X(_0594_));
 sg13g2_nor2_1 _1233_ (.A(net13),
    .B(_0594_),
    .Y(_0015_));
 sg13g2_and4_1 _1234_ (.A(\debug_out.uart_tx_inst.cycle_cnt[4] ),
    .B(\debug_out.uart_tx_inst.cycle_cnt[5] ),
    .C(\debug_out.uart_tx_inst.cycle_cnt[6] ),
    .D(_0589_),
    .X(_0595_));
 sg13g2_xnor2_1 _1235_ (.Y(_0596_),
    .A(\debug_out.uart_tx_inst.cycle_cnt[7] ),
    .B(_0595_));
 sg13g2_nor2_1 _1236_ (.A(net13),
    .B(_0596_),
    .Y(_0016_));
 sg13g2_nand2_1 _1237_ (.Y(_0597_),
    .A(\debug_out.uart_tx_inst.cycle_cnt[7] ),
    .B(_0595_));
 sg13g2_xor2_1 _1238_ (.B(_0597_),
    .A(\debug_out.uart_tx_inst.cycle_cnt[8] ),
    .X(_0598_));
 sg13g2_nor2_1 _1239_ (.A(_0582_),
    .B(_0598_),
    .Y(_0017_));
 sg13g2_nand3_1 _1240_ (.B(\debug_out.uart_tx_inst.cycle_cnt[8] ),
    .C(_0595_),
    .A(\debug_out.uart_tx_inst.cycle_cnt[7] ),
    .Y(_0599_));
 sg13g2_xor2_1 _1241_ (.B(_0599_),
    .A(_0534_),
    .X(_0600_));
 sg13g2_nor2_1 _1242_ (.A(net13),
    .B(_0600_),
    .Y(_0018_));
 sg13g2_inv_1 _1243_ (.Y(_0601_),
    .A(_0599_));
 sg13g2_nand2_1 _1244_ (.Y(_0602_),
    .A(_0534_),
    .B(_0601_));
 sg13g2_xor2_1 _1245_ (.B(_0602_),
    .A(\debug_out.uart_tx_inst.cycle_cnt[10] ),
    .X(_0603_));
 sg13g2_nor2_1 _1246_ (.A(_0581_),
    .B(_0603_),
    .Y(_0004_));
 sg13g2_nand3_1 _1247_ (.B(\debug_out.uart_tx_inst.cycle_cnt[10] ),
    .C(_0601_),
    .A(_0534_),
    .Y(_0604_));
 sg13g2_xor2_1 _1248_ (.B(_0604_),
    .A(\debug_out.uart_tx_inst.cycle_cnt[11] ),
    .X(_0605_));
 sg13g2_nor2_1 _1249_ (.A(_0581_),
    .B(_0605_),
    .Y(_0005_));
 sg13g2_nand4_1 _1250_ (.B(\debug_out.uart_tx_inst.cycle_cnt[11] ),
    .C(\debug_out.uart_tx_inst.cycle_cnt[10] ),
    .A(_0534_),
    .Y(_0606_),
    .D(_0601_));
 sg13g2_xor2_1 _1251_ (.B(_0606_),
    .A(\debug_out.uart_tx_inst.cycle_cnt[12] ),
    .X(_0607_));
 sg13g2_nor2_1 _1252_ (.A(_0581_),
    .B(_0607_),
    .Y(_0006_));
 sg13g2_nand4_1 _1253_ (.B(\debug_out.uart_tx_inst.cycle_cnt[11] ),
    .C(\debug_out.uart_tx_inst.cycle_cnt[10] ),
    .A(_0534_),
    .Y(_0608_),
    .D(\debug_out.uart_tx_inst.cycle_cnt[12] ));
 sg13g2_nor2_1 _1254_ (.A(_0599_),
    .B(_0608_),
    .Y(_0609_));
 sg13g2_xnor2_1 _1255_ (.Y(_0610_),
    .A(\debug_out.uart_tx_inst.cycle_cnt[13] ),
    .B(_0609_));
 sg13g2_nor2_1 _1256_ (.A(_0581_),
    .B(_0610_),
    .Y(_0007_));
 sg13g2_nand2_1 _1257_ (.Y(_0611_),
    .A(\debug_out.uart_tx_inst.cycle_cnt[13] ),
    .B(_0609_));
 sg13g2_xor2_1 _1258_ (.B(_0611_),
    .A(\debug_out.uart_tx_inst.cycle_cnt[14] ),
    .X(_0612_));
 sg13g2_nor2_1 _1259_ (.A(_0581_),
    .B(_0612_),
    .Y(_0008_));
 sg13g2_nand3_1 _1260_ (.B(\debug_out.uart_tx_inst.cycle_cnt[14] ),
    .C(_0609_),
    .A(\debug_out.uart_tx_inst.cycle_cnt[13] ),
    .Y(_0613_));
 sg13g2_xor2_1 _1261_ (.B(_0613_),
    .A(\debug_out.uart_tx_inst.cycle_cnt[15] ),
    .X(_0614_));
 sg13g2_nor2_1 _1262_ (.A(_0581_),
    .B(_0614_),
    .Y(_0009_));
 sg13g2_buf_2 _1263_ (.A(\autosel.i2c.state[1] ),
    .X(_0615_));
 sg13g2_buf_2 _1264_ (.A(\autosel.i2c.state[2] ),
    .X(_0616_));
 sg13g2_nor2b_1 _1265_ (.A(_0615_),
    .B_N(_0616_),
    .Y(_0617_));
 sg13g2_inv_1 _1266_ (.Y(_0618_),
    .A(\autosel.eeprom_busy ));
 sg13g2_a21oi_1 _1267_ (.A1(_0038_),
    .A2(_0617_),
    .Y(_0619_),
    .B1(_0618_));
 sg13g2_nor2b_1 _1268_ (.A(\autosel.i2c.i2c.busy_reg ),
    .B_N(\autosel.i2c.start ),
    .Y(_0620_));
 sg13g2_buf_1 _1269_ (.A(\autosel.i2c.state[0] ),
    .X(_0621_));
 sg13g2_nor2_1 _1270_ (.A(_0615_),
    .B(net51),
    .Y(_0622_));
 sg13g2_nand2_1 _1271_ (.Y(_0623_),
    .A(_0035_),
    .B(_0622_));
 sg13g2_nor2_1 _1272_ (.A(_0616_),
    .B(_0623_),
    .Y(_0624_));
 sg13g2_mux2_1 _1273_ (.A0(_0619_),
    .A1(_0620_),
    .S(_0624_),
    .X(_0065_));
 sg13g2_buf_1 _1274_ (.A(\autosel.i2c.i2c.missed_ack_reg ),
    .X(_0625_));
 sg13g2_buf_1 _1275_ (.A(net50),
    .X(_0626_));
 sg13g2_nor2b_1 _1276_ (.A(net35),
    .B_N(\autosel.i2c.i2c.m_axis_data_tdata_reg[0] ),
    .Y(_0627_));
 sg13g2_nor2b_2 _1277_ (.A(_0616_),
    .B_N(_0615_),
    .Y(_0628_));
 sg13g2_a21o_1 _1278_ (.A2(_0628_),
    .A1(net51),
    .B1(_0625_),
    .X(_0629_));
 sg13g2_nand4_1 _1279_ (.B(_0036_),
    .C(_0037_),
    .A(net51),
    .Y(_0630_),
    .D(_0628_));
 sg13g2_and2_1 _1280_ (.A(_0629_),
    .B(_0630_),
    .X(_0631_));
 sg13g2_buf_1 _1281_ (.A(_0631_),
    .X(_0632_));
 sg13g2_buf_1 _1282_ (.A(net21),
    .X(_0633_));
 sg13g2_mux2_1 _1283_ (.A0(\autosel.eeprom_data[0] ),
    .A1(_0627_),
    .S(_0633_),
    .X(_0066_));
 sg13g2_nor2b_1 _1284_ (.A(net35),
    .B_N(\autosel.i2c.data_out_hi[2] ),
    .Y(_0634_));
 sg13g2_mux2_1 _1285_ (.A0(\autosel.eeprom_data[10] ),
    .A1(_0634_),
    .S(net19),
    .X(_0067_));
 sg13g2_buf_2 _1286_ (.A(\autosel.eeprom_data[11] ),
    .X(_0635_));
 sg13g2_nor2b_1 _1287_ (.A(net35),
    .B_N(\autosel.i2c.data_out_hi[3] ),
    .Y(_0636_));
 sg13g2_mux2_1 _1288_ (.A0(_0635_),
    .A1(_0636_),
    .S(net19),
    .X(_0068_));
 sg13g2_nor2b_1 _1289_ (.A(net35),
    .B_N(\autosel.i2c.data_out_hi[4] ),
    .Y(_0637_));
 sg13g2_mux2_1 _1290_ (.A0(\autosel.eeprom_data[12] ),
    .A1(_0637_),
    .S(net19),
    .X(_0069_));
 sg13g2_inv_1 _1291_ (.Y(_0638_),
    .A(\autosel.eeprom_data[13] ));
 sg13g2_nand3b_1 _1292_ (.B(\autosel.i2c.data_out_hi[5] ),
    .C(net21),
    .Y(_0639_),
    .A_N(net50));
 sg13g2_o21ai_1 _1293_ (.B1(_0639_),
    .Y(_0070_),
    .A1(_0638_),
    .A2(net19));
 sg13g2_buf_1 _1294_ (.A(\autosel.eeprom_data[14] ),
    .X(_0640_));
 sg13g2_inv_1 _1295_ (.Y(_0641_),
    .A(_0640_));
 sg13g2_nand3b_1 _1296_ (.B(\autosel.i2c.data_out_hi[6] ),
    .C(net21),
    .Y(_0642_),
    .A_N(net50));
 sg13g2_o21ai_1 _1297_ (.B1(_0642_),
    .Y(_0071_),
    .A1(_0641_),
    .A2(net19));
 sg13g2_nor2b_1 _1298_ (.A(net35),
    .B_N(\autosel.i2c.data_out_hi[7] ),
    .Y(_0643_));
 sg13g2_mux2_1 _1299_ (.A0(\autosel.eeprom_data[15] ),
    .A1(_0643_),
    .S(net19),
    .X(_0072_));
 sg13g2_buf_2 _1300_ (.A(\autosel.eeprom_data[1] ),
    .X(_0644_));
 sg13g2_nor2b_1 _1301_ (.A(net35),
    .B_N(\autosel.i2c.i2c.m_axis_data_tdata_reg[1] ),
    .Y(_0645_));
 sg13g2_mux2_1 _1302_ (.A0(_0644_),
    .A1(_0645_),
    .S(net19),
    .X(_0073_));
 sg13g2_nor2b_1 _1303_ (.A(_0626_),
    .B_N(\autosel.i2c.i2c.m_axis_data_tdata_reg[2] ),
    .Y(_0646_));
 sg13g2_mux2_1 _1304_ (.A0(\autosel.eeprom_data[2] ),
    .A1(_0646_),
    .S(_0633_),
    .X(_0074_));
 sg13g2_buf_1 _1305_ (.A(\autosel.eeprom_data[3] ),
    .X(_0647_));
 sg13g2_nor2b_1 _1306_ (.A(net35),
    .B_N(\autosel.i2c.i2c.m_axis_data_tdata_reg[3] ),
    .Y(_0648_));
 sg13g2_mux2_1 _1307_ (.A0(net49),
    .A1(_0648_),
    .S(net19),
    .X(_0075_));
 sg13g2_nor2b_1 _1308_ (.A(net35),
    .B_N(\autosel.i2c.i2c.m_axis_data_tdata_reg[4] ),
    .Y(_0649_));
 sg13g2_mux2_1 _1309_ (.A0(\autosel.eeprom_data[4] ),
    .A1(_0649_),
    .S(net21),
    .X(_0076_));
 sg13g2_nor2b_1 _1310_ (.A(net50),
    .B_N(\autosel.i2c.i2c.m_axis_data_tdata_reg[5] ),
    .Y(_0650_));
 sg13g2_mux2_1 _1311_ (.A0(\autosel.eeprom_data[5] ),
    .A1(_0650_),
    .S(net21),
    .X(_0077_));
 sg13g2_nor2b_1 _1312_ (.A(net50),
    .B_N(\autosel.i2c.i2c.m_axis_data_tdata_reg[6] ),
    .Y(_0651_));
 sg13g2_mux2_1 _1313_ (.A0(\autosel.eeprom_data[6] ),
    .A1(_0651_),
    .S(net21),
    .X(_0078_));
 sg13g2_buf_1 _1314_ (.A(\autosel.eeprom_data[7] ),
    .X(_0652_));
 sg13g2_nor2b_1 _1315_ (.A(net50),
    .B_N(\autosel.i2c.i2c.m_axis_data_tdata_reg[7] ),
    .Y(_0653_));
 sg13g2_mux2_1 _1316_ (.A0(net48),
    .A1(_0653_),
    .S(net21),
    .X(_0079_));
 sg13g2_nor2b_1 _1317_ (.A(net50),
    .B_N(\autosel.i2c.data_out_hi[0] ),
    .Y(_0654_));
 sg13g2_mux2_1 _1318_ (.A0(\autosel.eeprom_data[8] ),
    .A1(_0654_),
    .S(net21),
    .X(_0080_));
 sg13g2_buf_2 _1319_ (.A(\autosel.eeprom_data[9] ),
    .X(_0655_));
 sg13g2_nor2b_1 _1320_ (.A(net50),
    .B_N(\autosel.i2c.data_out_hi[1] ),
    .Y(_0656_));
 sg13g2_mux2_1 _1321_ (.A0(_0655_),
    .A1(_0656_),
    .S(_0632_),
    .X(_0081_));
 sg13g2_nand2b_1 _1322_ (.Y(_0657_),
    .B(_0615_),
    .A_N(_0616_));
 sg13g2_buf_1 _1323_ (.A(_0657_),
    .X(_0658_));
 sg13g2_nor2_1 _1324_ (.A(_0621_),
    .B(net24),
    .Y(_0659_));
 sg13g2_and3_1 _1325_ (.X(_0660_),
    .A(net55),
    .B(\autosel.i2c.i2c.m_axis_data_tvalid_reg ),
    .C(_0659_));
 sg13g2_buf_4 _1326_ (.X(_0661_),
    .A(_0660_));
 sg13g2_mux2_1 _1327_ (.A0(\autosel.i2c.data_out_hi[0] ),
    .A1(\autosel.i2c.i2c.m_axis_data_tdata_reg[0] ),
    .S(_0661_),
    .X(_0082_));
 sg13g2_mux2_1 _1328_ (.A0(\autosel.i2c.data_out_hi[1] ),
    .A1(\autosel.i2c.i2c.m_axis_data_tdata_reg[1] ),
    .S(_0661_),
    .X(_0083_));
 sg13g2_mux2_1 _1329_ (.A0(\autosel.i2c.data_out_hi[2] ),
    .A1(\autosel.i2c.i2c.m_axis_data_tdata_reg[2] ),
    .S(_0661_),
    .X(_0084_));
 sg13g2_mux2_1 _1330_ (.A0(\autosel.i2c.data_out_hi[3] ),
    .A1(\autosel.i2c.i2c.m_axis_data_tdata_reg[3] ),
    .S(_0661_),
    .X(_0085_));
 sg13g2_mux2_1 _1331_ (.A0(\autosel.i2c.data_out_hi[4] ),
    .A1(\autosel.i2c.i2c.m_axis_data_tdata_reg[4] ),
    .S(_0661_),
    .X(_0086_));
 sg13g2_mux2_1 _1332_ (.A0(\autosel.i2c.data_out_hi[5] ),
    .A1(\autosel.i2c.i2c.m_axis_data_tdata_reg[5] ),
    .S(_0661_),
    .X(_0087_));
 sg13g2_mux2_1 _1333_ (.A0(\autosel.i2c.data_out_hi[6] ),
    .A1(\autosel.i2c.i2c.m_axis_data_tdata_reg[6] ),
    .S(_0661_),
    .X(_0088_));
 sg13g2_mux2_1 _1334_ (.A0(\autosel.i2c.data_out_hi[7] ),
    .A1(\autosel.i2c.i2c.m_axis_data_tdata_reg[7] ),
    .S(_0661_),
    .X(_0089_));
 sg13g2_buf_1 _1335_ (.A(\autosel.i2c.i2c.addr_reg[4] ),
    .X(_0662_));
 sg13g2_nand3b_1 _1336_ (.B(net51),
    .C(_0035_),
    .Y(_0663_),
    .A_N(_0615_));
 sg13g2_buf_2 _1337_ (.A(_0663_),
    .X(_0664_));
 sg13g2_a21o_1 _1338_ (.A2(_0664_),
    .A1(net24),
    .B1(_0040_),
    .X(_0665_));
 sg13g2_buf_8 _1339_ (.A(\autosel.i2c.i2c.phy_state_reg[1] ),
    .X(_0666_));
 sg13g2_buf_8 _1340_ (.A(\autosel.i2c.i2c.phy_state_reg[3] ),
    .X(_0667_));
 sg13g2_buf_1 _1341_ (.A(\autosel.i2c.i2c.phy_state_reg[2] ),
    .X(_0668_));
 sg13g2_nor3_1 _1342_ (.A(net47),
    .B(_0667_),
    .C(_0668_),
    .Y(_0669_));
 sg13g2_buf_1 _1343_ (.A(\autosel.i2c.i2c.state_reg[0] ),
    .X(_0670_));
 sg13g2_buf_1 _1344_ (.A(net46),
    .X(_0671_));
 sg13g2_buf_8 _1345_ (.A(\autosel.i2c.i2c.state_reg[1] ),
    .X(_0672_));
 sg13g2_buf_1 _1346_ (.A(net45),
    .X(_0673_));
 sg13g2_nand2_1 _1347_ (.Y(_0674_),
    .A(net33),
    .B(_0673_));
 sg13g2_buf_8 _1348_ (.A(\autosel.i2c.i2c.state_reg[3] ),
    .X(_0675_));
 sg13g2_buf_1 _1349_ (.A(\autosel.i2c.i2c.state_reg[2] ),
    .X(_0676_));
 sg13g2_nor2_2 _1350_ (.A(net44),
    .B(net43),
    .Y(_0677_));
 sg13g2_nand3_1 _1351_ (.B(_0674_),
    .C(_0677_),
    .A(net34),
    .Y(_0678_));
 sg13g2_nor2_1 _1352_ (.A(_0665_),
    .B(_0678_),
    .Y(_0679_));
 sg13g2_or2_1 _1353_ (.X(_0090_),
    .B(_0679_),
    .A(_0662_));
 sg13g2_buf_1 _1354_ (.A(\autosel.i2c.i2c.bit_count_reg[0] ),
    .X(_0680_));
 sg13g2_inv_1 _1355_ (.Y(_0681_),
    .A(net42));
 sg13g2_inv_1 _1356_ (.Y(_0682_),
    .A(net33));
 sg13g2_buf_1 _1357_ (.A(net43),
    .X(_0683_));
 sg13g2_nor2_1 _1358_ (.A(net31),
    .B(_0042_),
    .Y(_0684_));
 sg13g2_buf_1 _1359_ (.A(_0675_),
    .X(_0685_));
 sg13g2_a21oi_1 _1360_ (.A1(_0672_),
    .A2(_0684_),
    .Y(_0686_),
    .B1(net30));
 sg13g2_nor2_1 _1361_ (.A(net23),
    .B(_0686_),
    .Y(_0687_));
 sg13g2_nor3_2 _1362_ (.A(net45),
    .B(net44),
    .C(net43),
    .Y(_0688_));
 sg13g2_a21oi_2 _1363_ (.B1(_0040_),
    .Y(_0689_),
    .A2(_0664_),
    .A1(net24));
 sg13g2_nand2_1 _1364_ (.Y(_0690_),
    .A(_0042_),
    .B(_0689_));
 sg13g2_and3_1 _1365_ (.X(_0691_),
    .A(net23),
    .B(_0688_),
    .C(_0690_));
 sg13g2_nor2b_2 _1366_ (.A(net44),
    .B_N(net43),
    .Y(_0692_));
 sg13g2_nand2_1 _1367_ (.Y(_0693_),
    .A(net23),
    .B(\autosel.i2c.i2c.mode_read_reg ));
 sg13g2_inv_1 _1368_ (.Y(_0694_),
    .A(\autosel.i2c.i2c.s_axis_data_tready_reg ));
 sg13g2_or3_1 _1369_ (.A(_0682_),
    .B(_0694_),
    .C(_0664_),
    .X(_0695_));
 sg13g2_nand4_1 _1370_ (.B(_0692_),
    .C(_0693_),
    .A(net45),
    .Y(_0696_),
    .D(_0695_));
 sg13g2_buf_1 _1371_ (.A(\autosel.i2c.i2c.s_axis_cmd_ready_reg ),
    .X(_0697_));
 sg13g2_nor2b_2 _1372_ (.A(net46),
    .B_N(\autosel.i2c.i2c.state_reg[1] ),
    .Y(_0698_));
 sg13g2_o21ai_1 _1373_ (.B1(_0664_),
    .Y(_0699_),
    .A1(_0662_),
    .A2(net24));
 sg13g2_nand4_1 _1374_ (.B(_0677_),
    .C(_0698_),
    .A(net41),
    .Y(_0700_),
    .D(_0699_));
 sg13g2_inv_1 _1375_ (.Y(_0701_),
    .A(_0666_));
 sg13g2_nor2_1 _1376_ (.A(_0667_),
    .B(_0668_),
    .Y(_0702_));
 sg13g2_nand2_1 _1377_ (.Y(_0703_),
    .A(_0701_),
    .B(_0702_));
 sg13g2_a21oi_1 _1378_ (.A1(net30),
    .A2(net31),
    .Y(_0704_),
    .B1(net22));
 sg13g2_nand3_1 _1379_ (.B(_0700_),
    .C(_0704_),
    .A(_0696_),
    .Y(_0705_));
 sg13g2_nor2b_2 _1380_ (.A(net45),
    .B_N(net46),
    .Y(_0706_));
 sg13g2_and2_1 _1381_ (.A(_0677_),
    .B(_0706_),
    .X(_0707_));
 sg13g2_and3_1 _1382_ (.X(_0708_),
    .A(_0662_),
    .B(net24),
    .C(_0707_));
 sg13g2_o21ai_1 _1383_ (.B1(_0677_),
    .Y(_0709_),
    .A1(_0698_),
    .A2(_0706_));
 sg13g2_a21oi_1 _1384_ (.A1(net41),
    .A2(_0040_),
    .Y(_0710_),
    .B1(_0709_));
 sg13g2_inv_1 _1385_ (.Y(_0711_),
    .A(net41));
 sg13g2_a21o_1 _1386_ (.A2(_0664_),
    .A1(net24),
    .B1(_0711_),
    .X(_0712_));
 sg13g2_mux2_1 _1387_ (.A0(_0708_),
    .A1(_0710_),
    .S(_0712_),
    .X(_0713_));
 sg13g2_nor4_2 _1388_ (.A(_0687_),
    .B(_0691_),
    .C(_0705_),
    .Y(_0714_),
    .D(_0713_));
 sg13g2_nand2b_2 _1389_ (.Y(_0715_),
    .B(net44),
    .A_N(net43));
 sg13g2_nand2_1 _1390_ (.Y(_0716_),
    .A(_0692_),
    .B(_0706_));
 sg13g2_o21ai_1 _1391_ (.B1(_0716_),
    .Y(_0717_),
    .A1(net33),
    .A2(_0715_));
 sg13g2_buf_1 _1392_ (.A(_0717_),
    .X(_0718_));
 sg13g2_nand3_1 _1393_ (.B(_0714_),
    .C(_0718_),
    .A(_0047_),
    .Y(_0719_));
 sg13g2_o21ai_1 _1394_ (.B1(_0719_),
    .Y(_0091_),
    .A1(_0681_),
    .A2(_0714_));
 sg13g2_buf_1 _1395_ (.A(\autosel.i2c.i2c.bit_count_reg[1] ),
    .X(_0720_));
 sg13g2_or2_1 _1396_ (.X(_0721_),
    .B(net40),
    .A(net42));
 sg13g2_nand2_1 _1397_ (.Y(_0722_),
    .A(_0714_),
    .B(_0718_));
 sg13g2_nand2_1 _1398_ (.Y(_0723_),
    .A(_0680_),
    .B(_0718_));
 sg13g2_inv_1 _1399_ (.Y(_0724_),
    .A(net40));
 sg13g2_a21o_1 _1400_ (.A2(_0723_),
    .A1(_0714_),
    .B1(_0724_),
    .X(_0725_));
 sg13g2_o21ai_1 _1401_ (.B1(_0725_),
    .Y(_0092_),
    .A1(_0721_),
    .A2(_0722_));
 sg13g2_and2_1 _1402_ (.A(_0714_),
    .B(_0718_),
    .X(_0726_));
 sg13g2_buf_2 _1403_ (.A(\autosel.i2c.i2c.bit_count_reg[2] ),
    .X(_0727_));
 sg13g2_nor3_2 _1404_ (.A(_0727_),
    .B(_0680_),
    .C(net40),
    .Y(_0728_));
 sg13g2_nand2_1 _1405_ (.Y(_0729_),
    .A(_0718_),
    .B(_0721_));
 sg13g2_inv_1 _1406_ (.Y(_0730_),
    .A(_0727_));
 sg13g2_a21oi_1 _1407_ (.A1(_0714_),
    .A2(_0729_),
    .Y(_0731_),
    .B1(_0730_));
 sg13g2_a21o_1 _1408_ (.A2(_0728_),
    .A1(_0726_),
    .B1(_0731_),
    .X(_0093_));
 sg13g2_buf_2 _1409_ (.A(\autosel.i2c.i2c.bit_count_reg[3] ),
    .X(_0732_));
 sg13g2_inv_1 _1410_ (.Y(_0733_),
    .A(_0732_));
 sg13g2_inv_1 _1411_ (.Y(_0734_),
    .A(_0718_));
 sg13g2_o21ai_1 _1412_ (.B1(_0714_),
    .Y(_0735_),
    .A1(_0734_),
    .A2(_0728_));
 sg13g2_and2_1 _1413_ (.A(_0732_),
    .B(_0728_),
    .X(_0736_));
 sg13g2_a22oi_1 _1414_ (.Y(_0094_),
    .B1(_0736_),
    .B2(_0726_),
    .A2(_0735_),
    .A1(_0733_));
 sg13g2_inv_1 _1415_ (.Y(_0737_),
    .A(\autosel.i2c.i2c.phy_rx_data_reg ));
 sg13g2_nor2b_1 _1416_ (.A(net43),
    .B_N(net44),
    .Y(_0738_));
 sg13g2_buf_2 _1417_ (.A(_0738_),
    .X(_0739_));
 sg13g2_nand2_1 _1418_ (.Y(_0740_),
    .A(_0698_),
    .B(_0739_));
 sg13g2_nor2_1 _1419_ (.A(_0737_),
    .B(_0740_),
    .Y(_0741_));
 sg13g2_inv_1 _1420_ (.Y(_0742_),
    .A(_0705_));
 sg13g2_nor2_1 _1421_ (.A(net30),
    .B(net41),
    .Y(_0743_));
 sg13g2_inv_1 _1422_ (.Y(_0744_),
    .A(net31));
 sg13g2_o21ai_1 _1423_ (.B1(_0744_),
    .Y(_0745_),
    .A1(net33),
    .A2(_0743_));
 sg13g2_or2_1 _1424_ (.X(_0746_),
    .B(net31),
    .A(net30));
 sg13g2_buf_1 _1425_ (.A(_0746_),
    .X(_0747_));
 sg13g2_nand2b_2 _1426_ (.Y(_0748_),
    .B(\autosel.i2c.i2c.state_reg[1] ),
    .A_N(net46));
 sg13g2_nor3_2 _1427_ (.A(_0040_),
    .B(_0747_),
    .C(_0748_),
    .Y(_0749_));
 sg13g2_nand3_1 _1428_ (.B(_0664_),
    .C(_0749_),
    .A(_0658_),
    .Y(_0750_));
 sg13g2_nand4_1 _1429_ (.B(_0742_),
    .C(_0745_),
    .A(net32),
    .Y(_0751_),
    .D(_0750_));
 sg13g2_buf_4 _1430_ (.X(_0752_),
    .A(_0751_));
 sg13g2_mux2_1 _1431_ (.A0(_0741_),
    .A1(\autosel.i2c.i2c.data_reg[0] ),
    .S(_0752_),
    .X(_0097_));
 sg13g2_nor2_2 _1432_ (.A(_0748_),
    .B(_0715_),
    .Y(_0753_));
 sg13g2_and2_1 _1433_ (.A(\autosel.i2c.i2c.data_reg[0] ),
    .B(_0753_),
    .X(_0754_));
 sg13g2_mux2_1 _1434_ (.A0(_0754_),
    .A1(\autosel.i2c.i2c.data_reg[1] ),
    .S(_0752_),
    .X(_0098_));
 sg13g2_and2_1 _1435_ (.A(\autosel.i2c.i2c.data_reg[1] ),
    .B(_0753_),
    .X(_0755_));
 sg13g2_mux2_1 _1436_ (.A0(_0755_),
    .A1(\autosel.i2c.i2c.data_reg[2] ),
    .S(_0752_),
    .X(_0099_));
 sg13g2_and2_1 _1437_ (.A(\autosel.i2c.i2c.data_reg[2] ),
    .B(_0753_),
    .X(_0756_));
 sg13g2_mux2_1 _1438_ (.A0(_0756_),
    .A1(\autosel.i2c.i2c.data_reg[3] ),
    .S(_0752_),
    .X(_0100_));
 sg13g2_and2_1 _1439_ (.A(\autosel.i2c.i2c.data_reg[3] ),
    .B(_0753_),
    .X(_0757_));
 sg13g2_mux2_1 _1440_ (.A0(_0757_),
    .A1(\autosel.i2c.i2c.data_reg[4] ),
    .S(_0752_),
    .X(_0101_));
 sg13g2_and2_1 _1441_ (.A(\autosel.i2c.i2c.data_reg[4] ),
    .B(_0753_),
    .X(_0758_));
 sg13g2_mux2_1 _1442_ (.A0(_0758_),
    .A1(\autosel.i2c.i2c.data_reg[5] ),
    .S(_0752_),
    .X(_0102_));
 sg13g2_and2_1 _1443_ (.A(\autosel.i2c.i2c.data_reg[5] ),
    .B(_0753_),
    .X(_0759_));
 sg13g2_mux2_1 _1444_ (.A0(_0759_),
    .A1(\autosel.i2c.i2c.data_reg[6] ),
    .S(_0752_),
    .X(_0103_));
 sg13g2_and2_1 _1445_ (.A(\autosel.i2c.i2c.data_reg[6] ),
    .B(_0753_),
    .X(_0760_));
 sg13g2_mux2_1 _1446_ (.A0(_0760_),
    .A1(\autosel.i2c.i2c.data_reg[7] ),
    .S(_0752_),
    .X(_0104_));
 sg13g2_or4_1 _1447_ (.A(_0732_),
    .B(_0727_),
    .C(\autosel.i2c.i2c.bit_count_reg[0] ),
    .D(\autosel.i2c.i2c.bit_count_reg[1] ),
    .X(_0761_));
 sg13g2_buf_2 _1448_ (.A(_0761_),
    .X(_0762_));
 sg13g2_nor3_1 _1449_ (.A(_0748_),
    .B(_0715_),
    .C(_0762_),
    .Y(_0763_));
 sg13g2_nand2_1 _1450_ (.Y(_0764_),
    .A(net34),
    .B(_0763_));
 sg13g2_buf_1 _1451_ (.A(_0764_),
    .X(_0765_));
 sg13g2_nand2_1 _1452_ (.Y(_0766_),
    .A(\autosel.i2c.i2c.m_axis_data_tdata_reg[0] ),
    .B(_0765_));
 sg13g2_o21ai_1 _1453_ (.B1(_0766_),
    .Y(_0123_),
    .A1(_0737_),
    .A2(net18));
 sg13g2_mux2_1 _1454_ (.A0(\autosel.i2c.i2c.data_reg[0] ),
    .A1(\autosel.i2c.i2c.m_axis_data_tdata_reg[1] ),
    .S(net18),
    .X(_0124_));
 sg13g2_mux2_1 _1455_ (.A0(\autosel.i2c.i2c.data_reg[1] ),
    .A1(\autosel.i2c.i2c.m_axis_data_tdata_reg[2] ),
    .S(net18),
    .X(_0125_));
 sg13g2_mux2_1 _1456_ (.A0(\autosel.i2c.i2c.data_reg[2] ),
    .A1(\autosel.i2c.i2c.m_axis_data_tdata_reg[3] ),
    .S(net18),
    .X(_0126_));
 sg13g2_mux2_1 _1457_ (.A0(\autosel.i2c.i2c.data_reg[3] ),
    .A1(\autosel.i2c.i2c.m_axis_data_tdata_reg[4] ),
    .S(net18),
    .X(_0127_));
 sg13g2_mux2_1 _1458_ (.A0(\autosel.i2c.i2c.data_reg[4] ),
    .A1(\autosel.i2c.i2c.m_axis_data_tdata_reg[5] ),
    .S(net18),
    .X(_0128_));
 sg13g2_mux2_1 _1459_ (.A0(\autosel.i2c.i2c.data_reg[5] ),
    .A1(\autosel.i2c.i2c.m_axis_data_tdata_reg[6] ),
    .S(net18),
    .X(_0129_));
 sg13g2_mux2_1 _1460_ (.A0(\autosel.i2c.i2c.data_reg[6] ),
    .A1(\autosel.i2c.i2c.m_axis_data_tdata_reg[7] ),
    .S(net18),
    .X(_0130_));
 sg13g2_mux2_1 _1461_ (.A0(\autosel.i2c.i2c.mode_read_reg ),
    .A1(_0628_),
    .S(_0679_),
    .X(_0133_));
 sg13g2_buf_1 _1462_ (.A(\autosel.i2c.i2c.mode_stop_reg ),
    .X(_0767_));
 sg13g2_o21ai_1 _1463_ (.B1(net51),
    .Y(_0768_),
    .A1(_0617_),
    .A2(_0628_));
 sg13g2_inv_1 _1464_ (.Y(_0769_),
    .A(_0768_));
 sg13g2_mux2_1 _1465_ (.A0(_0767_),
    .A1(_0769_),
    .S(_0679_),
    .X(_0134_));
 sg13g2_buf_1 _1466_ (.A(\autosel.i2c.i2c.delay_reg[11] ),
    .X(_0770_));
 sg13g2_nor4_1 _1467_ (.A(\autosel.i2c.i2c.delay_reg[14] ),
    .B(\autosel.i2c.i2c.delay_reg[13] ),
    .C(\autosel.i2c.i2c.delay_reg[12] ),
    .D(_0770_),
    .Y(_0771_));
 sg13g2_nor2b_2 _1468_ (.A(\autosel.i2c.i2c.delay_reg[15] ),
    .B_N(_0771_),
    .Y(_0772_));
 sg13g2_nor2_2 _1469_ (.A(\autosel.i2c.i2c.delay_reg[10] ),
    .B(\autosel.i2c.i2c.delay_reg[9] ),
    .Y(_0773_));
 sg13g2_inv_1 _1470_ (.Y(_0774_),
    .A(\autosel.i2c.i2c.delay_reg[8] ));
 sg13g2_nor4_2 _1471_ (.A(\autosel.i2c.i2c.delay_reg[3] ),
    .B(\autosel.i2c.i2c.delay_reg[2] ),
    .C(\autosel.i2c.i2c.delay_reg[1] ),
    .Y(_0775_),
    .D(\autosel.i2c.i2c.delay_reg[0] ));
 sg13g2_nor2_1 _1472_ (.A(\autosel.i2c.i2c.delay_reg[4] ),
    .B(\autosel.i2c.i2c.delay_reg[5] ),
    .Y(_0776_));
 sg13g2_nor2_1 _1473_ (.A(\autosel.i2c.i2c.delay_reg[6] ),
    .B(\autosel.i2c.i2c.delay_reg[7] ),
    .Y(_0777_));
 sg13g2_and4_1 _1474_ (.A(_0774_),
    .B(_0775_),
    .C(_0776_),
    .D(_0777_),
    .X(_0778_));
 sg13g2_buf_2 _1475_ (.A(_0778_),
    .X(_0779_));
 sg13g2_nand3_1 _1476_ (.B(_0773_),
    .C(_0779_),
    .A(_0772_),
    .Y(_0780_));
 sg13g2_buf_1 _1477_ (.A(_0780_),
    .X(_0781_));
 sg13g2_buf_1 _1478_ (.A(\autosel.i2c.i2c.phy_state_reg[0] ),
    .X(_0782_));
 sg13g2_inv_2 _1479_ (.Y(_0783_),
    .A(net39));
 sg13g2_nand2_1 _1480_ (.Y(_0784_),
    .A(net47),
    .B(_0783_));
 sg13g2_buf_1 _1481_ (.A(_0668_),
    .X(_0785_));
 sg13g2_buf_1 _1482_ (.A(_0667_),
    .X(_0786_));
 sg13g2_nand3b_1 _1483_ (.B(_0039_),
    .C(net28),
    .Y(_0787_),
    .A_N(net29));
 sg13g2_nor4_1 _1484_ (.A(\autosel.i2c.i2c.delay_sda_reg ),
    .B(_0781_),
    .C(_0784_),
    .D(_0787_),
    .Y(_0788_));
 sg13g2_nand2_1 _1485_ (.Y(_0789_),
    .A(\autosel.i2c.i2c.sda_i_reg ),
    .B(_0788_));
 sg13g2_o21ai_1 _1486_ (.B1(_0789_),
    .Y(_0135_),
    .A1(_0737_),
    .A2(_0788_));
 sg13g2_inv_1 _1487_ (.Y(_0790_),
    .A(net51));
 sg13g2_inv_1 _1488_ (.Y(_0791_),
    .A(_0664_));
 sg13g2_a22oi_1 _1489_ (.Y(_0792_),
    .B1(_0791_),
    .B2(_0694_),
    .A2(_0617_),
    .A1(\autosel.i2c.i2c.busy_reg ));
 sg13g2_nand2_1 _1490_ (.Y(_0793_),
    .A(_0037_),
    .B(_0628_));
 sg13g2_o21ai_1 _1491_ (.B1(_0793_),
    .Y(_0794_),
    .A1(_0620_),
    .A2(_0623_));
 sg13g2_nand2_1 _1492_ (.Y(_0795_),
    .A(_0036_),
    .B(_0794_));
 sg13g2_o21ai_1 _1493_ (.B1(_0795_),
    .Y(_0796_),
    .A1(_0625_),
    .A2(_0792_));
 sg13g2_o21ai_1 _1494_ (.B1(_0623_),
    .Y(_0797_),
    .A1(net51),
    .A2(net24));
 sg13g2_nor3_1 _1495_ (.A(_0626_),
    .B(_0796_),
    .C(_0797_),
    .Y(_0798_));
 sg13g2_a21oi_1 _1496_ (.A1(_0790_),
    .A2(_0796_),
    .Y(_0148_),
    .B1(_0798_));
 sg13g2_nor2_1 _1497_ (.A(_0659_),
    .B(_0791_),
    .Y(_0799_));
 sg13g2_o21ai_1 _1498_ (.B1(_0793_),
    .Y(_0800_),
    .A1(_0796_),
    .A2(_0799_));
 sg13g2_and2_1 _1499_ (.A(_0036_),
    .B(_0800_),
    .X(_0149_));
 sg13g2_mux2_1 _1500_ (.A0(_0629_),
    .A1(_0616_),
    .S(_0796_),
    .X(_0150_));
 sg13g2_nand2_1 _1501_ (.Y(_0801_),
    .A(_0559_),
    .B(_0561_));
 sg13g2_xnor2_1 _1502_ (.Y(_0802_),
    .A(_0553_),
    .B(_0554_));
 sg13g2_nor2_1 _1503_ (.A(_0801_),
    .B(_0802_),
    .Y(_0193_));
 sg13g2_nand2_1 _1504_ (.Y(_0803_),
    .A(_0553_),
    .B(_0554_));
 sg13g2_xor2_1 _1505_ (.B(_0803_),
    .A(_0552_),
    .X(_0804_));
 sg13g2_nor2_1 _1506_ (.A(_0801_),
    .B(_0804_),
    .Y(_0194_));
 sg13g2_o21ai_1 _1507_ (.B1(\debug_out.uart_tx_inst.bit_cnt[2] ),
    .Y(_0805_),
    .A1(_0537_),
    .A2(_0544_));
 sg13g2_nand2_1 _1508_ (.Y(_0806_),
    .A(_0552_),
    .B(_0553_));
 sg13g2_xor2_1 _1509_ (.B(_0806_),
    .A(_0046_),
    .X(_0807_));
 sg13g2_nand2_1 _1510_ (.Y(_0808_),
    .A(_0554_),
    .B(_0807_));
 sg13g2_a21oi_1 _1511_ (.A1(_0805_),
    .A2(_0808_),
    .Y(_0195_),
    .B1(_0801_));
 sg13g2_mux2_1 _1512_ (.A0(\debug_out.uart_tx_inst.tx_data_latch[0] ),
    .A1(\debug_out.tx_byte[0] ),
    .S(_0565_),
    .X(_0196_));
 sg13g2_mux2_1 _1513_ (.A0(\debug_out.uart_tx_inst.tx_data_latch[1] ),
    .A1(\debug_out.tx_byte[1] ),
    .S(_0565_),
    .X(_0197_));
 sg13g2_mux2_1 _1514_ (.A0(\debug_out.uart_tx_inst.tx_data_latch[2] ),
    .A1(\debug_out.tx_byte[2] ),
    .S(_0565_),
    .X(_0198_));
 sg13g2_mux2_1 _1515_ (.A0(\debug_out.uart_tx_inst.tx_data_latch[3] ),
    .A1(\debug_out.tx_byte[3] ),
    .S(_0565_),
    .X(_0199_));
 sg13g2_mux2_1 _1516_ (.A0(\debug_out.uart_tx_inst.tx_data_latch[4] ),
    .A1(\debug_out.tx_byte[4] ),
    .S(_0565_),
    .X(_0200_));
 sg13g2_mux2_1 _1517_ (.A0(\debug_out.uart_tx_inst.tx_data_latch[6] ),
    .A1(\debug_out.tx_byte[6] ),
    .S(_0565_),
    .X(_0201_));
 sg13g2_nor2_1 _1518_ (.A(net53),
    .B(_0545_),
    .Y(_0809_));
 sg13g2_nor3_1 _1519_ (.A(_0560_),
    .B(_0546_),
    .C(\debug_out.tx_valid ),
    .Y(_0810_));
 sg13g2_a21oi_1 _1520_ (.A1(_0554_),
    .A2(_0809_),
    .Y(_0811_),
    .B1(_0810_));
 sg13g2_buf_2 _1521_ (.A(\debug_out.tx_ready ),
    .X(_0812_));
 sg13g2_o21ai_1 _1522_ (.B1(_0812_),
    .Y(_0813_),
    .A1(_0546_),
    .A2(_0564_));
 sg13g2_o21ai_1 _1523_ (.B1(_0813_),
    .Y(_0202_),
    .A1(net52),
    .A2(_0811_));
 sg13g2_a22oi_1 _1524_ (.Y(_0814_),
    .B1(_0706_),
    .B2(_0739_),
    .A2(_0698_),
    .A1(_0692_));
 sg13g2_nand2_1 _1525_ (.Y(_0815_),
    .A(net55),
    .B(net34));
 sg13g2_nor3_1 _1526_ (.A(_0737_),
    .B(_0814_),
    .C(_0815_),
    .Y(_0132_));
 sg13g2_nor2_1 _1527_ (.A(\autosel.i2c.i2c.m_axis_data_tvalid_reg ),
    .B(net41),
    .Y(_0816_));
 sg13g2_a21oi_1 _1528_ (.A1(_0037_),
    .A2(net41),
    .Y(_0817_),
    .B1(_0816_));
 sg13g2_nor3_1 _1529_ (.A(_0747_),
    .B(_0748_),
    .C(_0817_),
    .Y(_0818_));
 sg13g2_a22oi_1 _1530_ (.Y(_0819_),
    .B1(_0712_),
    .B2(_0818_),
    .A2(_0688_),
    .A1(_0665_));
 sg13g2_nor2_1 _1531_ (.A(_0815_),
    .B(_0819_),
    .Y(_0140_));
 sg13g2_inv_1 _1532_ (.Y(_0820_),
    .A(_0672_));
 sg13g2_nor2b_1 _1533_ (.A(_0676_),
    .B_N(net46),
    .Y(_0821_));
 sg13g2_nor2_1 _1534_ (.A(_0820_),
    .B(_0744_),
    .Y(_0822_));
 sg13g2_a21oi_1 _1535_ (.A1(_0820_),
    .A2(_0821_),
    .Y(_0823_),
    .B1(_0822_));
 sg13g2_inv_1 _1536_ (.Y(_0824_),
    .A(_0696_));
 sg13g2_a21oi_1 _1537_ (.A1(_0689_),
    .A2(_0708_),
    .Y(_0825_),
    .B1(_0824_));
 sg13g2_nor4_1 _1538_ (.A(net30),
    .B(_0815_),
    .C(_0823_),
    .D(_0825_),
    .Y(_0141_));
 sg13g2_inv_1 _1539_ (.Y(_0826_),
    .A(_0049_));
 sg13g2_nor4_1 _1540_ (.A(\debug_out.counter[12] ),
    .B(\debug_out.counter[15] ),
    .C(\debug_out.counter[14] ),
    .D(\debug_out.counter[17] ),
    .Y(_0827_));
 sg13g2_nand3b_1 _1541_ (.B(\debug_out.counter[8] ),
    .C(_0827_),
    .Y(_0828_),
    .A_N(\debug_out.counter[9] ));
 sg13g2_nor4_1 _1542_ (.A(\debug_out.counter[1] ),
    .B(\debug_out.counter[26] ),
    .C(\debug_out.counter[31] ),
    .D(\debug_out.counter[30] ),
    .Y(_0829_));
 sg13g2_nor4_1 _1543_ (.A(\debug_out.counter[19] ),
    .B(\debug_out.counter[27] ),
    .C(\debug_out.counter[29] ),
    .D(\debug_out.counter[28] ),
    .Y(_0830_));
 sg13g2_buf_1 _1544_ (.A(\debug_out.counter[4] ),
    .X(_0831_));
 sg13g2_inv_1 _1545_ (.Y(_0832_),
    .A(\debug_out.counter[16] ));
 sg13g2_nor4_1 _1546_ (.A(_0831_),
    .B(\debug_out.counter[7] ),
    .C(\debug_out.counter[6] ),
    .D(_0832_),
    .Y(_0833_));
 sg13g2_nor4_1 _1547_ (.A(\debug_out.counter[0] ),
    .B(\debug_out.counter[3] ),
    .C(\debug_out.counter[2] ),
    .D(\debug_out.counter[5] ),
    .Y(_0834_));
 sg13g2_nand4_1 _1548_ (.B(_0830_),
    .C(_0833_),
    .A(_0829_),
    .Y(_0835_),
    .D(_0834_));
 sg13g2_nor4_1 _1549_ (.A(\debug_out.counter[18] ),
    .B(\debug_out.counter[23] ),
    .C(\debug_out.counter[22] ),
    .D(\debug_out.counter[25] ),
    .Y(_0836_));
 sg13g2_and2_1 _1550_ (.A(\debug_out.counter[20] ),
    .B(\debug_out.counter[21] ),
    .X(_0837_));
 sg13g2_buf_1 _1551_ (.A(_0837_),
    .X(_0838_));
 sg13g2_and3_1 _1552_ (.X(_0839_),
    .A(\debug_out.counter[10] ),
    .B(\debug_out.counter[11] ),
    .C(\debug_out.counter[13] ));
 sg13g2_nand4_1 _1553_ (.B(_0836_),
    .C(_0838_),
    .A(\debug_out.counter[24] ),
    .Y(_0840_),
    .D(_0839_));
 sg13g2_nor3_2 _1554_ (.A(_0828_),
    .B(_0835_),
    .C(_0840_),
    .Y(_0841_));
 sg13g2_nand2b_1 _1555_ (.Y(_0842_),
    .B(net55),
    .A_N(_0841_));
 sg13g2_buf_2 _1556_ (.A(_0842_),
    .X(_0843_));
 sg13g2_buf_1 _1557_ (.A(_0843_),
    .X(_0844_));
 sg13g2_nor2_1 _1558_ (.A(_0826_),
    .B(net17),
    .Y(_0151_));
 sg13g2_and4_1 _1559_ (.A(\debug_out.counter[1] ),
    .B(\debug_out.counter[0] ),
    .C(\debug_out.counter[3] ),
    .D(\debug_out.counter[2] ),
    .X(_0845_));
 sg13g2_buf_8 _1560_ (.A(_0845_),
    .X(_0846_));
 sg13g2_and4_1 _1561_ (.A(\debug_out.counter[5] ),
    .B(_0831_),
    .C(\debug_out.counter[6] ),
    .D(_0846_),
    .X(_0847_));
 sg13g2_buf_1 _1562_ (.A(_0847_),
    .X(_0848_));
 sg13g2_and3_1 _1563_ (.X(_0849_),
    .A(\debug_out.counter[7] ),
    .B(\debug_out.counter[9] ),
    .C(\debug_out.counter[8] ));
 sg13g2_and2_1 _1564_ (.A(_0848_),
    .B(_0849_),
    .X(_0850_));
 sg13g2_buf_1 _1565_ (.A(_0850_),
    .X(_0851_));
 sg13g2_xnor2_1 _1566_ (.Y(_0852_),
    .A(\debug_out.counter[10] ),
    .B(_0851_));
 sg13g2_nor2_1 _1567_ (.A(net17),
    .B(_0852_),
    .Y(_0152_));
 sg13g2_nand2_1 _1568_ (.Y(_0853_),
    .A(\debug_out.counter[10] ),
    .B(_0851_));
 sg13g2_xor2_1 _1569_ (.B(_0853_),
    .A(\debug_out.counter[11] ),
    .X(_0854_));
 sg13g2_nor2_1 _1570_ (.A(net17),
    .B(_0854_),
    .Y(_0153_));
 sg13g2_nand3_1 _1571_ (.B(\debug_out.counter[11] ),
    .C(_0851_),
    .A(\debug_out.counter[10] ),
    .Y(_0855_));
 sg13g2_xor2_1 _1572_ (.B(_0855_),
    .A(\debug_out.counter[12] ),
    .X(_0856_));
 sg13g2_nor2_1 _1573_ (.A(net17),
    .B(_0856_),
    .Y(_0154_));
 sg13g2_nand4_1 _1574_ (.B(\debug_out.counter[11] ),
    .C(\debug_out.counter[12] ),
    .A(\debug_out.counter[10] ),
    .Y(_0857_),
    .D(_0851_));
 sg13g2_xor2_1 _1575_ (.B(_0857_),
    .A(\debug_out.counter[13] ),
    .X(_0858_));
 sg13g2_nor2_1 _1576_ (.A(net17),
    .B(_0858_),
    .Y(_0155_));
 sg13g2_and3_1 _1577_ (.X(_0859_),
    .A(\debug_out.counter[12] ),
    .B(_0839_),
    .C(_0851_));
 sg13g2_xnor2_1 _1578_ (.Y(_0860_),
    .A(\debug_out.counter[14] ),
    .B(_0859_));
 sg13g2_nor2_1 _1579_ (.A(net17),
    .B(_0860_),
    .Y(_0156_));
 sg13g2_nand2_1 _1580_ (.Y(_0861_),
    .A(\debug_out.counter[14] ),
    .B(_0859_));
 sg13g2_xor2_1 _1581_ (.B(_0861_),
    .A(\debug_out.counter[15] ),
    .X(_0862_));
 sg13g2_nor2_1 _1582_ (.A(net17),
    .B(_0862_),
    .Y(_0157_));
 sg13g2_nand4_1 _1583_ (.B(_0831_),
    .C(\debug_out.counter[6] ),
    .A(\debug_out.counter[5] ),
    .Y(_0863_),
    .D(_0846_));
 sg13g2_and2_1 _1584_ (.A(\debug_out.counter[12] ),
    .B(\debug_out.counter[15] ),
    .X(_0864_));
 sg13g2_nand4_1 _1585_ (.B(_0839_),
    .C(_0849_),
    .A(\debug_out.counter[14] ),
    .Y(_0865_),
    .D(_0864_));
 sg13g2_nor2_1 _1586_ (.A(_0863_),
    .B(_0865_),
    .Y(_0866_));
 sg13g2_xnor2_1 _1587_ (.Y(_0867_),
    .A(\debug_out.counter[16] ),
    .B(_0866_));
 sg13g2_nor2_1 _1588_ (.A(net17),
    .B(_0867_),
    .Y(_0158_));
 sg13g2_nor3_2 _1589_ (.A(_0832_),
    .B(_0863_),
    .C(_0865_),
    .Y(_0868_));
 sg13g2_xnor2_1 _1590_ (.Y(_0869_),
    .A(\debug_out.counter[17] ),
    .B(_0868_));
 sg13g2_nor2_1 _1591_ (.A(_0844_),
    .B(_0869_),
    .Y(_0159_));
 sg13g2_nand2_1 _1592_ (.Y(_0870_),
    .A(\debug_out.counter[17] ),
    .B(_0868_));
 sg13g2_xor2_1 _1593_ (.B(_0870_),
    .A(\debug_out.counter[18] ),
    .X(_0871_));
 sg13g2_nor2_1 _1594_ (.A(_0844_),
    .B(_0871_),
    .Y(_0160_));
 sg13g2_buf_1 _1595_ (.A(_0843_),
    .X(_0872_));
 sg13g2_nand3_1 _1596_ (.B(\debug_out.counter[18] ),
    .C(_0868_),
    .A(\debug_out.counter[17] ),
    .Y(_0873_));
 sg13g2_xor2_1 _1597_ (.B(_0873_),
    .A(\debug_out.counter[19] ),
    .X(_0874_));
 sg13g2_nor2_1 _1598_ (.A(net16),
    .B(_0874_),
    .Y(_0161_));
 sg13g2_xnor2_1 _1599_ (.Y(_0875_),
    .A(\debug_out.counter[1] ),
    .B(\debug_out.counter[0] ));
 sg13g2_nor2_1 _1600_ (.A(net16),
    .B(_0875_),
    .Y(_0162_));
 sg13g2_nand4_1 _1601_ (.B(\debug_out.counter[16] ),
    .C(\debug_out.counter[19] ),
    .A(\debug_out.counter[17] ),
    .Y(_0876_),
    .D(\debug_out.counter[18] ));
 sg13g2_nor3_2 _1602_ (.A(_0863_),
    .B(_0865_),
    .C(_0876_),
    .Y(_0877_));
 sg13g2_xnor2_1 _1603_ (.Y(_0878_),
    .A(\debug_out.counter[20] ),
    .B(_0877_));
 sg13g2_nor2_1 _1604_ (.A(net16),
    .B(_0878_),
    .Y(_0163_));
 sg13g2_nand2_1 _1605_ (.Y(_0879_),
    .A(\debug_out.counter[20] ),
    .B(_0877_));
 sg13g2_xor2_1 _1606_ (.B(_0879_),
    .A(\debug_out.counter[21] ),
    .X(_0880_));
 sg13g2_nor2_1 _1607_ (.A(net16),
    .B(_0880_),
    .Y(_0164_));
 sg13g2_nand2_1 _1608_ (.Y(_0881_),
    .A(_0838_),
    .B(_0877_));
 sg13g2_xor2_1 _1609_ (.B(_0881_),
    .A(\debug_out.counter[22] ),
    .X(_0882_));
 sg13g2_nor2_1 _1610_ (.A(net16),
    .B(_0882_),
    .Y(_0165_));
 sg13g2_nand3_1 _1611_ (.B(_0838_),
    .C(_0877_),
    .A(\debug_out.counter[22] ),
    .Y(_0883_));
 sg13g2_xor2_1 _1612_ (.B(_0883_),
    .A(\debug_out.counter[23] ),
    .X(_0884_));
 sg13g2_nor2_1 _1613_ (.A(net16),
    .B(_0884_),
    .Y(_0166_));
 sg13g2_and2_1 _1614_ (.A(\debug_out.counter[23] ),
    .B(\debug_out.counter[22] ),
    .X(_0885_));
 sg13g2_nand3_1 _1615_ (.B(_0877_),
    .C(_0885_),
    .A(_0838_),
    .Y(_0886_));
 sg13g2_xor2_1 _1616_ (.B(_0886_),
    .A(\debug_out.counter[24] ),
    .X(_0887_));
 sg13g2_nor2_1 _1617_ (.A(net16),
    .B(_0887_),
    .Y(_0167_));
 sg13g2_and3_1 _1618_ (.X(_0888_),
    .A(\debug_out.counter[24] ),
    .B(_0838_),
    .C(_0885_));
 sg13g2_nand2_1 _1619_ (.Y(_0889_),
    .A(_0877_),
    .B(_0888_));
 sg13g2_xor2_1 _1620_ (.B(_0889_),
    .A(\debug_out.counter[25] ),
    .X(_0890_));
 sg13g2_nor2_1 _1621_ (.A(_0872_),
    .B(_0890_),
    .Y(_0168_));
 sg13g2_nand3_1 _1622_ (.B(_0877_),
    .C(_0888_),
    .A(\debug_out.counter[25] ),
    .Y(_0891_));
 sg13g2_xor2_1 _1623_ (.B(_0891_),
    .A(\debug_out.counter[26] ),
    .X(_0892_));
 sg13g2_nor2_1 _1624_ (.A(_0872_),
    .B(_0892_),
    .Y(_0169_));
 sg13g2_and4_1 _1625_ (.A(\debug_out.counter[25] ),
    .B(\debug_out.counter[26] ),
    .C(_0877_),
    .D(_0888_),
    .X(_0893_));
 sg13g2_buf_2 _1626_ (.A(_0893_),
    .X(_0894_));
 sg13g2_xnor2_1 _1627_ (.Y(_0895_),
    .A(\debug_out.counter[27] ),
    .B(_0894_));
 sg13g2_nor2_1 _1628_ (.A(net16),
    .B(_0895_),
    .Y(_0170_));
 sg13g2_buf_1 _1629_ (.A(_0843_),
    .X(_0896_));
 sg13g2_nand2_1 _1630_ (.Y(_0897_),
    .A(\debug_out.counter[27] ),
    .B(_0894_));
 sg13g2_xor2_1 _1631_ (.B(_0897_),
    .A(\debug_out.counter[28] ),
    .X(_0898_));
 sg13g2_nor2_1 _1632_ (.A(net15),
    .B(_0898_),
    .Y(_0171_));
 sg13g2_and2_1 _1633_ (.A(\debug_out.counter[27] ),
    .B(\debug_out.counter[28] ),
    .X(_0899_));
 sg13g2_nand2_1 _1634_ (.Y(_0900_),
    .A(_0894_),
    .B(_0899_));
 sg13g2_xor2_1 _1635_ (.B(_0900_),
    .A(\debug_out.counter[29] ),
    .X(_0901_));
 sg13g2_nor2_1 _1636_ (.A(net15),
    .B(_0901_),
    .Y(_0172_));
 sg13g2_nand2_1 _1637_ (.Y(_0902_),
    .A(\debug_out.counter[1] ),
    .B(\debug_out.counter[0] ));
 sg13g2_xor2_1 _1638_ (.B(_0902_),
    .A(\debug_out.counter[2] ),
    .X(_0903_));
 sg13g2_nor2_1 _1639_ (.A(net15),
    .B(_0903_),
    .Y(_0173_));
 sg13g2_nand3_1 _1640_ (.B(_0894_),
    .C(_0899_),
    .A(\debug_out.counter[29] ),
    .Y(_0904_));
 sg13g2_xor2_1 _1641_ (.B(_0904_),
    .A(\debug_out.counter[30] ),
    .X(_0905_));
 sg13g2_nor2_1 _1642_ (.A(_0896_),
    .B(_0905_),
    .Y(_0174_));
 sg13g2_nand4_1 _1643_ (.B(\debug_out.counter[30] ),
    .C(_0894_),
    .A(\debug_out.counter[29] ),
    .Y(_0906_),
    .D(_0899_));
 sg13g2_xor2_1 _1644_ (.B(_0906_),
    .A(\debug_out.counter[31] ),
    .X(_0907_));
 sg13g2_nor2_1 _1645_ (.A(_0896_),
    .B(_0907_),
    .Y(_0175_));
 sg13g2_nand3_1 _1646_ (.B(\debug_out.counter[0] ),
    .C(\debug_out.counter[2] ),
    .A(\debug_out.counter[1] ),
    .Y(_0908_));
 sg13g2_xor2_1 _1647_ (.B(_0908_),
    .A(\debug_out.counter[3] ),
    .X(_0909_));
 sg13g2_nor2_1 _1648_ (.A(net15),
    .B(_0909_),
    .Y(_0176_));
 sg13g2_xnor2_1 _1649_ (.Y(_0910_),
    .A(_0831_),
    .B(_0846_));
 sg13g2_nor2_1 _1650_ (.A(net15),
    .B(_0910_),
    .Y(_0177_));
 sg13g2_nand2_1 _1651_ (.Y(_0911_),
    .A(_0831_),
    .B(_0846_));
 sg13g2_xor2_1 _1652_ (.B(_0911_),
    .A(\debug_out.counter[5] ),
    .X(_0912_));
 sg13g2_nor2_1 _1653_ (.A(net15),
    .B(_0912_),
    .Y(_0178_));
 sg13g2_nand3_1 _1654_ (.B(_0831_),
    .C(_0846_),
    .A(\debug_out.counter[5] ),
    .Y(_0913_));
 sg13g2_xor2_1 _1655_ (.B(_0913_),
    .A(\debug_out.counter[6] ),
    .X(_0914_));
 sg13g2_nor2_1 _1656_ (.A(net15),
    .B(_0914_),
    .Y(_0179_));
 sg13g2_xnor2_1 _1657_ (.Y(_0915_),
    .A(\debug_out.counter[7] ),
    .B(_0848_));
 sg13g2_nor2_1 _1658_ (.A(net15),
    .B(_0915_),
    .Y(_0180_));
 sg13g2_nand2_1 _1659_ (.Y(_0916_),
    .A(\debug_out.counter[7] ),
    .B(_0848_));
 sg13g2_xor2_1 _1660_ (.B(_0916_),
    .A(\debug_out.counter[8] ),
    .X(_0917_));
 sg13g2_nor2_1 _1661_ (.A(_0843_),
    .B(_0917_),
    .Y(_0181_));
 sg13g2_nand3_1 _1662_ (.B(\debug_out.counter[8] ),
    .C(_0848_),
    .A(\debug_out.counter[7] ),
    .Y(_0918_));
 sg13g2_xor2_1 _1663_ (.B(_0918_),
    .A(\debug_out.counter[9] ),
    .X(_0919_));
 sg13g2_nor2_1 _1664_ (.A(_0843_),
    .B(_0919_),
    .Y(_0182_));
 sg13g2_buf_1 _1665_ (.A(\debug_out.send_index[1] ),
    .X(_0920_));
 sg13g2_buf_1 _1666_ (.A(\debug_out.send_index[2] ),
    .X(_0921_));
 sg13g2_nand2_1 _1667_ (.Y(_0922_),
    .A(net38),
    .B(_0921_));
 sg13g2_nand3_1 _1668_ (.B(_0050_),
    .C(_0922_),
    .A(_0812_),
    .Y(_0923_));
 sg13g2_buf_1 _1669_ (.A(\debug_out.send_index[0] ),
    .X(_0924_));
 sg13g2_nand2_1 _1670_ (.Y(_0925_),
    .A(_0812_),
    .B(_0922_));
 sg13g2_nand2_1 _1671_ (.Y(_0926_),
    .A(net37),
    .B(_0925_));
 sg13g2_a21oi_1 _1672_ (.A1(_0923_),
    .A2(_0926_),
    .Y(_0183_),
    .B1(_0843_));
 sg13g2_nor2b_1 _1673_ (.A(_0921_),
    .B_N(net37),
    .Y(_0927_));
 sg13g2_and3_1 _1674_ (.X(_0928_),
    .A(net38),
    .B(_0812_),
    .C(_0927_));
 sg13g2_a21oi_1 _1675_ (.A1(net37),
    .A2(_0812_),
    .Y(_0929_),
    .B1(net38));
 sg13g2_nor3_1 _1676_ (.A(_0843_),
    .B(_0928_),
    .C(_0929_),
    .Y(_0184_));
 sg13g2_inv_1 _1677_ (.Y(_0930_),
    .A(_0921_));
 sg13g2_nand3_1 _1678_ (.B(net37),
    .C(_0812_),
    .A(net38),
    .Y(_0931_));
 sg13g2_a21oi_1 _1679_ (.A1(_0930_),
    .A2(_0931_),
    .Y(_0185_),
    .B1(_0843_));
 sg13g2_xor2_1 _1680_ (.B(\autosel.eeprom_data[6] ),
    .A(\autosel.addr_counter[6] ),
    .X(_0932_));
 sg13g2_xor2_1 _1681_ (.B(\autosel.eeprom_data[5] ),
    .A(\autosel.addr_counter[5] ),
    .X(_0933_));
 sg13g2_xnor2_1 _1682_ (.Y(_0934_),
    .A(\autosel.addr_counter[2] ),
    .B(\autosel.eeprom_data[2] ));
 sg13g2_buf_1 _1683_ (.A(\autosel.addr_counter[1] ),
    .X(_0935_));
 sg13g2_xnor2_1 _1684_ (.Y(_0936_),
    .A(_0935_),
    .B(_0644_));
 sg13g2_xnor2_1 _1685_ (.Y(_0937_),
    .A(\autosel.addr_counter[9] ),
    .B(_0655_));
 sg13g2_xnor2_1 _1686_ (.Y(_0938_),
    .A(\autosel.addr_counter[4] ),
    .B(\autosel.eeprom_data[4] ));
 sg13g2_nand4_1 _1687_ (.B(_0936_),
    .C(_0937_),
    .A(_0934_),
    .Y(_0939_),
    .D(_0938_));
 sg13g2_xnor2_1 _1688_ (.Y(_0940_),
    .A(\autosel.addr_counter[8] ),
    .B(\autosel.eeprom_data[8] ));
 sg13g2_xnor2_1 _1689_ (.Y(_0941_),
    .A(\autosel.addr_counter[3] ),
    .B(net49));
 sg13g2_xnor2_1 _1690_ (.Y(_0942_),
    .A(\autosel.addr_counter[7] ),
    .B(_0652_));
 sg13g2_buf_1 _1691_ (.A(\autosel.addr_counter[0] ),
    .X(_0943_));
 sg13g2_xnor2_1 _1692_ (.Y(_0944_),
    .A(\autosel.eeprom_data[0] ),
    .B(_0943_));
 sg13g2_nand4_1 _1693_ (.B(_0941_),
    .C(_0942_),
    .A(_0940_),
    .Y(_0945_),
    .D(_0944_));
 sg13g2_nor4_2 _1694_ (.A(_0932_),
    .B(_0933_),
    .C(_0939_),
    .Y(_0946_),
    .D(_0945_));
 sg13g2_nand2_1 _1695_ (.Y(_0947_),
    .A(\autosel.state[1] ),
    .B(_0034_));
 sg13g2_nor2_2 _1696_ (.A(_0946_),
    .B(_0947_),
    .Y(_0948_));
 sg13g2_nand2_1 _1697_ (.Y(_0949_),
    .A(_0048_),
    .B(_0948_));
 sg13g2_o21ai_1 _1698_ (.B1(_0943_),
    .Y(_0950_),
    .A1(_0946_),
    .A2(_0947_));
 sg13g2_buf_1 _1699_ (.A(_0528_),
    .X(_0951_));
 sg13g2_a21oi_1 _1700_ (.A1(_0949_),
    .A2(_0950_),
    .Y(_0052_),
    .B1(net27));
 sg13g2_nand2_1 _1701_ (.Y(_0952_),
    .A(_0943_),
    .B(_0948_));
 sg13g2_xor2_1 _1702_ (.B(_0952_),
    .A(_0935_),
    .X(_0953_));
 sg13g2_nor2_1 _1703_ (.A(net36),
    .B(_0953_),
    .Y(_0053_));
 sg13g2_nand3_1 _1704_ (.B(_0935_),
    .C(_0948_),
    .A(_0943_),
    .Y(_0954_));
 sg13g2_xor2_1 _1705_ (.B(_0954_),
    .A(\autosel.addr_counter[2] ),
    .X(_0955_));
 sg13g2_nor2_1 _1706_ (.A(net36),
    .B(_0955_),
    .Y(_0054_));
 sg13g2_nand4_1 _1707_ (.B(_0935_),
    .C(\autosel.addr_counter[2] ),
    .A(_0943_),
    .Y(_0956_),
    .D(_0948_));
 sg13g2_xor2_1 _1708_ (.B(_0956_),
    .A(\autosel.addr_counter[3] ),
    .X(_0957_));
 sg13g2_nor2_1 _1709_ (.A(net36),
    .B(_0957_),
    .Y(_0055_));
 sg13g2_nand4_1 _1710_ (.B(_0935_),
    .C(\autosel.addr_counter[2] ),
    .A(_0943_),
    .Y(_0958_),
    .D(\autosel.addr_counter[3] ));
 sg13g2_or2_1 _1711_ (.X(_0959_),
    .B(_0958_),
    .A(_0947_));
 sg13g2_buf_1 _1712_ (.A(_0959_),
    .X(_0960_));
 sg13g2_o21ai_1 _1713_ (.B1(\autosel.addr_counter[4] ),
    .Y(_0961_),
    .A1(_0946_),
    .A2(_0960_));
 sg13g2_or3_1 _1714_ (.A(\autosel.addr_counter[4] ),
    .B(_0946_),
    .C(_0960_),
    .X(_0962_));
 sg13g2_a21oi_1 _1715_ (.A1(_0961_),
    .A2(_0962_),
    .Y(_0056_),
    .B1(net27));
 sg13g2_inv_1 _1716_ (.Y(_0963_),
    .A(\autosel.addr_counter[4] ));
 sg13g2_nor3_1 _1717_ (.A(_0963_),
    .B(_0946_),
    .C(_0960_),
    .Y(_0964_));
 sg13g2_xnor2_1 _1718_ (.Y(_0965_),
    .A(\autosel.addr_counter[5] ),
    .B(_0964_));
 sg13g2_nor2_1 _1719_ (.A(net36),
    .B(_0965_),
    .Y(_0057_));
 sg13g2_nand2_1 _1720_ (.Y(_0966_),
    .A(\autosel.addr_counter[4] ),
    .B(\autosel.addr_counter[5] ));
 sg13g2_nor3_1 _1721_ (.A(_0946_),
    .B(_0960_),
    .C(_0966_),
    .Y(_0967_));
 sg13g2_xnor2_1 _1722_ (.Y(_0968_),
    .A(\autosel.addr_counter[6] ),
    .B(_0967_));
 sg13g2_nor2_1 _1723_ (.A(net36),
    .B(_0968_),
    .Y(_0058_));
 sg13g2_inv_1 _1724_ (.Y(_0969_),
    .A(\autosel.addr_counter[6] ));
 sg13g2_nor4_2 _1725_ (.A(_0969_),
    .B(_0946_),
    .C(_0960_),
    .Y(_0970_),
    .D(_0966_));
 sg13g2_xnor2_1 _1726_ (.Y(_0971_),
    .A(\autosel.addr_counter[7] ),
    .B(_0970_));
 sg13g2_nor2_1 _1727_ (.A(net36),
    .B(_0971_),
    .Y(_0059_));
 sg13g2_nand2_1 _1728_ (.Y(_0972_),
    .A(\autosel.addr_counter[7] ),
    .B(_0970_));
 sg13g2_xor2_1 _1729_ (.B(_0972_),
    .A(\autosel.addr_counter[8] ),
    .X(_0973_));
 sg13g2_nor2_1 _1730_ (.A(_0000_),
    .B(_0973_),
    .Y(_0060_));
 sg13g2_nand3_1 _1731_ (.B(\autosel.addr_counter[8] ),
    .C(_0970_),
    .A(\autosel.addr_counter[7] ),
    .Y(_0974_));
 sg13g2_xor2_1 _1732_ (.B(_0974_),
    .A(\autosel.addr_counter[9] ),
    .X(_0975_));
 sg13g2_nor2_1 _1733_ (.A(_0000_),
    .B(_0975_),
    .Y(_0061_));
 sg13g2_inv_1 _1734_ (.Y(_0976_),
    .A(\autosel.state[1] ));
 sg13g2_nor2_1 _1735_ (.A(_0976_),
    .B(\autosel.ctrl_sel_inc ),
    .Y(_0977_));
 sg13g2_a21oi_1 _1736_ (.A1(_0946_),
    .A2(_0977_),
    .Y(_0978_),
    .B1(\autosel.ctrl_ena ));
 sg13g2_nor2_1 _1737_ (.A(net27),
    .B(_0978_),
    .Y(_0062_));
 sg13g2_a21oi_1 _1738_ (.A1(_0976_),
    .A2(\autosel.ctrl_sel_inc ),
    .Y(_0979_),
    .B1(_0948_));
 sg13g2_nor2_1 _1739_ (.A(net27),
    .B(_0979_),
    .Y(_0063_));
 sg13g2_o21ai_1 _1740_ (.B1(net54),
    .Y(_0980_),
    .A1(\autosel.ctrl_sel_rst_n ),
    .A2(_0529_));
 sg13g2_inv_1 _1741_ (.Y(_0064_),
    .A(_0980_));
 sg13g2_inv_1 _1742_ (.Y(_0981_),
    .A(\autosel.i2c.i2c.sda_i_reg ));
 sg13g2_a21o_1 _1743_ (.A2(\autosel.i2c.i2c.scl_i_reg ),
    .A1(\autosel.i2c.i2c.last_sda_i_reg ),
    .B1(\autosel.i2c.i2c.bus_active_reg ),
    .X(_0982_));
 sg13g2_nand2b_1 _1744_ (.Y(_0983_),
    .B(\autosel.i2c.i2c.scl_i_reg ),
    .A_N(\autosel.i2c.i2c.last_sda_i_reg ));
 sg13g2_a22oi_1 _1745_ (.Y(_0984_),
    .B1(_0983_),
    .B2(\autosel.i2c.i2c.bus_active_reg ),
    .A2(_0982_),
    .A1(_0981_));
 sg13g2_nor2_1 _1746_ (.A(net27),
    .B(_0984_),
    .Y(_0095_));
 sg13g2_and2_1 _1747_ (.A(net54),
    .B(_0678_),
    .X(_0096_));
 sg13g2_and3_1 _1748_ (.X(_0985_),
    .A(_0772_),
    .B(_0773_),
    .C(_0779_));
 sg13g2_buf_1 _1749_ (.A(_0985_),
    .X(_0986_));
 sg13g2_nand4_1 _1750_ (.B(_0657_),
    .C(_0677_),
    .A(_0662_),
    .Y(_0987_),
    .D(_0706_));
 sg13g2_a21oi_2 _1751_ (.B1(_0711_),
    .Y(_0988_),
    .A2(_0664_),
    .A1(_0657_));
 sg13g2_inv_1 _1752_ (.Y(_0989_),
    .A(_0675_));
 sg13g2_nand2b_1 _1753_ (.Y(_0990_),
    .B(\autosel.i2c.i2c.bus_active_reg ),
    .A_N(_0670_));
 sg13g2_and4_1 _1754_ (.A(_0989_),
    .B(net34),
    .C(_0688_),
    .D(_0990_),
    .X(_0991_));
 sg13g2_and3_1 _1755_ (.X(_0992_),
    .A(_0987_),
    .B(_0988_),
    .C(_0991_));
 sg13g2_and2_1 _1756_ (.A(net45),
    .B(_0042_),
    .X(_0993_));
 sg13g2_nor2_1 _1757_ (.A(net46),
    .B(net45),
    .Y(_0994_));
 sg13g2_a22oi_1 _1758_ (.Y(_0995_),
    .B1(_0994_),
    .B2(net43),
    .A2(_0993_),
    .A1(_0821_));
 sg13g2_or2_1 _1759_ (.X(_0996_),
    .B(_0667_),
    .A(_0685_));
 sg13g2_nor2_1 _1760_ (.A(net47),
    .B(net39),
    .Y(_0997_));
 sg13g2_nand2b_1 _1761_ (.Y(_0998_),
    .B(_0668_),
    .A_N(_0667_));
 sg13g2_and2_1 _1762_ (.A(_0997_),
    .B(_0998_),
    .X(_0999_));
 sg13g2_o21ai_1 _1763_ (.B1(_0999_),
    .Y(_1000_),
    .A1(_0995_),
    .A2(_0996_));
 sg13g2_xnor2_1 _1764_ (.Y(_1001_),
    .A(net47),
    .B(_0667_));
 sg13g2_nand3_1 _1765_ (.B(_0668_),
    .C(_1001_),
    .A(_0782_),
    .Y(_1002_));
 sg13g2_o21ai_1 _1766_ (.B1(_1002_),
    .Y(_1003_),
    .A1(_0992_),
    .A2(_1000_));
 sg13g2_or2_1 _1767_ (.X(_1004_),
    .B(_0995_),
    .A(net44));
 sg13g2_nand3_1 _1768_ (.B(_0988_),
    .C(_0991_),
    .A(_0987_),
    .Y(_1005_));
 sg13g2_nand3b_1 _1769_ (.B(net43),
    .C(net46),
    .Y(_1006_),
    .A_N(net44));
 sg13g2_o21ai_1 _1770_ (.B1(_1006_),
    .Y(_0203_),
    .A1(net46),
    .A2(_0715_));
 sg13g2_nor4_2 _1771_ (.A(_0732_),
    .B(_0727_),
    .C(net42),
    .Y(_0204_),
    .D(net40));
 sg13g2_nor2_1 _1772_ (.A(net45),
    .B(_0204_),
    .Y(_0205_));
 sg13g2_mux2_1 _1773_ (.A0(net51),
    .A1(_0035_),
    .S(_0615_),
    .X(_0206_));
 sg13g2_and4_1 _1774_ (.A(net41),
    .B(_0677_),
    .C(_0698_),
    .D(_0206_),
    .X(_0207_));
 sg13g2_a221oi_1 _1775_ (.B2(_0205_),
    .C1(_0207_),
    .B1(_0203_),
    .A1(_0767_),
    .Y(_0208_),
    .A2(_0763_));
 sg13g2_nor2_1 _1776_ (.A(_0783_),
    .B(net22),
    .Y(_0209_));
 sg13g2_and4_1 _1777_ (.A(_1004_),
    .B(_1005_),
    .C(_0208_),
    .D(_0209_),
    .X(_0210_));
 sg13g2_buf_1 _1778_ (.A(_0210_),
    .X(_0211_));
 sg13g2_nand2_1 _1779_ (.Y(_0212_),
    .A(_0739_),
    .B(_0994_));
 sg13g2_a21oi_1 _1780_ (.A1(_0692_),
    .A2(_0706_),
    .Y(_0213_),
    .B1(_0762_));
 sg13g2_a221oi_1 _1781_ (.B2(_0213_),
    .C1(net22),
    .B1(_0212_),
    .A1(_0740_),
    .Y(_0214_),
    .A2(_0762_));
 sg13g2_nand2b_1 _1782_ (.Y(_0215_),
    .B(_0621_),
    .A_N(_0615_));
 sg13g2_nor3_1 _1783_ (.A(_0035_),
    .B(_0040_),
    .C(_0215_),
    .Y(_0216_));
 sg13g2_o21ai_1 _1784_ (.B1(net44),
    .Y(_0217_),
    .A1(net45),
    .A2(_0767_));
 sg13g2_nor3_1 _1785_ (.A(net23),
    .B(_0683_),
    .C(_0217_),
    .Y(_0218_));
 sg13g2_a21o_1 _1786_ (.A2(_0216_),
    .A1(_0707_),
    .B1(_0218_),
    .X(_0219_));
 sg13g2_nor3_1 _1787_ (.A(_0781_),
    .B(_0214_),
    .C(_0219_),
    .Y(_0220_));
 sg13g2_nand2b_1 _1788_ (.Y(_0221_),
    .B(_0041_),
    .A_N(\autosel.i2c.i2c.delay_scl_reg ));
 sg13g2_a221oi_1 _1789_ (.B2(_0220_),
    .C1(_0221_),
    .B1(_0211_),
    .A1(_0986_),
    .Y(_0222_),
    .A2(_1003_));
 sg13g2_buf_2 _1790_ (.A(_0222_),
    .X(_0223_));
 sg13g2_buf_8 _1791_ (.A(_0223_),
    .X(_0224_));
 sg13g2_nand2b_1 _1792_ (.Y(_0225_),
    .B(\autosel.i2c.i2c.delay_reg[0] ),
    .A_N(net12));
 sg13g2_inv_1 _1793_ (.Y(_0226_),
    .A(_0044_));
 sg13g2_nor3_1 _1794_ (.A(_0781_),
    .B(_0784_),
    .C(_0998_),
    .Y(_0227_));
 sg13g2_a21oi_1 _1795_ (.A1(_0226_),
    .A2(_0781_),
    .Y(_0228_),
    .B1(_0227_));
 sg13g2_nand2_1 _1796_ (.Y(_0229_),
    .A(net12),
    .B(_0228_));
 sg13g2_buf_1 _1797_ (.A(_0528_),
    .X(_0230_));
 sg13g2_a21oi_1 _1798_ (.A1(_0225_),
    .A2(_0229_),
    .Y(_0105_),
    .B1(net26));
 sg13g2_nor2b_1 _1799_ (.A(\autosel.i2c.i2c.delay_scl_reg ),
    .B_N(_0041_),
    .Y(_0231_));
 sg13g2_nand2_1 _1800_ (.Y(_0232_),
    .A(_0779_),
    .B(_0231_));
 sg13g2_or4_1 _1801_ (.A(\autosel.i2c.i2c.delay_reg[10] ),
    .B(\autosel.i2c.i2c.delay_reg[9] ),
    .C(_0772_),
    .D(_0232_),
    .X(_0233_));
 sg13g2_o21ai_1 _1802_ (.B1(\autosel.i2c.i2c.delay_reg[10] ),
    .Y(_0234_),
    .A1(\autosel.i2c.i2c.delay_reg[9] ),
    .A2(_0232_));
 sg13g2_a21oi_1 _1803_ (.A1(_0233_),
    .A2(_0234_),
    .Y(_0106_),
    .B1(net26));
 sg13g2_nand3_1 _1804_ (.B(_0779_),
    .C(_0231_),
    .A(_0773_),
    .Y(_0235_));
 sg13g2_buf_1 _1805_ (.A(_0235_),
    .X(_0236_));
 sg13g2_nor3_1 _1806_ (.A(_0770_),
    .B(_0772_),
    .C(_0236_),
    .Y(_0237_));
 sg13g2_a21oi_1 _1807_ (.A1(_0770_),
    .A2(_0236_),
    .Y(_0238_),
    .B1(_0237_));
 sg13g2_nor2_1 _1808_ (.A(_0951_),
    .B(_0238_),
    .Y(_0107_));
 sg13g2_or4_1 _1809_ (.A(\autosel.i2c.i2c.delay_reg[12] ),
    .B(_0770_),
    .C(_0772_),
    .D(_0236_),
    .X(_0239_));
 sg13g2_o21ai_1 _1810_ (.B1(\autosel.i2c.i2c.delay_reg[12] ),
    .Y(_0240_),
    .A1(_0770_),
    .A2(_0236_));
 sg13g2_a21oi_1 _1811_ (.A1(_0239_),
    .A2(_0240_),
    .Y(_0108_),
    .B1(net26));
 sg13g2_nor2_1 _1812_ (.A(_0770_),
    .B(_0236_),
    .Y(_0241_));
 sg13g2_nand2b_1 _1813_ (.Y(_0242_),
    .B(_0241_),
    .A_N(\autosel.i2c.i2c.delay_reg[12] ));
 sg13g2_or3_1 _1814_ (.A(\autosel.i2c.i2c.delay_reg[13] ),
    .B(_0772_),
    .C(_0242_),
    .X(_0243_));
 sg13g2_nand2_1 _1815_ (.Y(_0244_),
    .A(\autosel.i2c.i2c.delay_reg[13] ),
    .B(_0242_));
 sg13g2_a21oi_1 _1816_ (.A1(_0243_),
    .A2(_0244_),
    .Y(_0109_),
    .B1(net26));
 sg13g2_o21ai_1 _1817_ (.B1(\autosel.i2c.i2c.delay_reg[14] ),
    .Y(_0245_),
    .A1(\autosel.i2c.i2c.delay_reg[13] ),
    .A2(_0242_));
 sg13g2_or4_1 _1818_ (.A(\autosel.i2c.i2c.delay_reg[14] ),
    .B(\autosel.i2c.i2c.delay_reg[13] ),
    .C(_0986_),
    .D(_0242_),
    .X(_0246_));
 sg13g2_a21oi_1 _1819_ (.A1(_0245_),
    .A2(_0246_),
    .Y(_0110_),
    .B1(net26));
 sg13g2_nand4_1 _1820_ (.B(_0773_),
    .C(_0779_),
    .A(_0771_),
    .Y(_0247_),
    .D(_0224_));
 sg13g2_and3_1 _1821_ (.X(_0111_),
    .A(net54),
    .B(\autosel.i2c.i2c.delay_reg[15] ),
    .C(_0247_));
 sg13g2_nor2_1 _1822_ (.A(_0528_),
    .B(\autosel.i2c.i2c.delay_reg[1] ),
    .Y(_0248_));
 sg13g2_and2_1 _1823_ (.A(net55),
    .B(\autosel.i2c.i2c.delay_reg[1] ),
    .X(_0249_));
 sg13g2_nand2b_1 _1824_ (.Y(_0250_),
    .B(_0223_),
    .A_N(\autosel.i2c.i2c.delay_reg[0] ));
 sg13g2_mux2_1 _1825_ (.A0(_0248_),
    .A1(_0249_),
    .S(_0250_),
    .X(_0112_));
 sg13g2_nor2_1 _1826_ (.A(_0528_),
    .B(\autosel.i2c.i2c.delay_reg[2] ),
    .Y(_0251_));
 sg13g2_and2_1 _1827_ (.A(net55),
    .B(\autosel.i2c.i2c.delay_reg[2] ),
    .X(_0252_));
 sg13g2_nor2_1 _1828_ (.A(\autosel.i2c.i2c.delay_reg[1] ),
    .B(\autosel.i2c.i2c.delay_reg[0] ),
    .Y(_0253_));
 sg13g2_nand2_1 _1829_ (.Y(_0254_),
    .A(_0253_),
    .B(_0223_));
 sg13g2_mux2_1 _1830_ (.A0(_0251_),
    .A1(_0252_),
    .S(_0254_),
    .X(_0113_));
 sg13g2_nor3_1 _1831_ (.A(\autosel.i2c.i2c.delay_reg[2] ),
    .B(\autosel.i2c.i2c.delay_reg[1] ),
    .C(\autosel.i2c.i2c.delay_reg[0] ),
    .Y(_0255_));
 sg13g2_nand2_1 _1832_ (.Y(_0256_),
    .A(net55),
    .B(\autosel.i2c.i2c.delay_reg[3] ));
 sg13g2_a21oi_1 _1833_ (.A1(_0255_),
    .A2(net12),
    .Y(_0257_),
    .B1(_0256_));
 sg13g2_o21ai_1 _1834_ (.B1(_0986_),
    .Y(_0258_),
    .A1(_0784_),
    .A2(_0998_));
 sg13g2_nand4_1 _1835_ (.B(_0775_),
    .C(net12),
    .A(net54),
    .Y(_0259_),
    .D(_0258_));
 sg13g2_nand2b_1 _1836_ (.Y(_0114_),
    .B(_0259_),
    .A_N(_0257_));
 sg13g2_nand2_1 _1837_ (.Y(_0260_),
    .A(_0775_),
    .B(_0231_));
 sg13g2_nor2_1 _1838_ (.A(\autosel.i2c.i2c.delay_reg[4] ),
    .B(_0260_),
    .Y(_0261_));
 sg13g2_and2_1 _1839_ (.A(_0781_),
    .B(_0261_),
    .X(_0262_));
 sg13g2_a21oi_1 _1840_ (.A1(\autosel.i2c.i2c.delay_reg[4] ),
    .A2(_0260_),
    .Y(_0263_),
    .B1(_0262_));
 sg13g2_nor2_1 _1841_ (.A(net27),
    .B(_0263_),
    .Y(_0115_));
 sg13g2_nor2_1 _1842_ (.A(_0528_),
    .B(\autosel.i2c.i2c.delay_reg[5] ),
    .Y(_0264_));
 sg13g2_a22oi_1 _1843_ (.Y(_0265_),
    .B1(_0211_),
    .B2(_0220_),
    .A2(_1003_),
    .A1(_0986_));
 sg13g2_nand2_1 _1844_ (.Y(_0266_),
    .A(_0527_),
    .B(\autosel.i2c.i2c.delay_reg[5] ));
 sg13g2_a21oi_1 _1845_ (.A1(_0265_),
    .A2(_0261_),
    .Y(_0267_),
    .B1(_0266_));
 sg13g2_a21o_1 _1846_ (.A2(_0264_),
    .A1(_0262_),
    .B1(_0267_),
    .X(_0116_));
 sg13g2_nand2_1 _1847_ (.Y(_0268_),
    .A(_0775_),
    .B(_0776_));
 sg13g2_inv_1 _1848_ (.Y(_0269_),
    .A(_0268_));
 sg13g2_nor2_1 _1849_ (.A(\autosel.i2c.i2c.delay_reg[6] ),
    .B(_0227_),
    .Y(_0270_));
 sg13g2_nand3_1 _1850_ (.B(net12),
    .C(_0270_),
    .A(_0269_),
    .Y(_0271_));
 sg13g2_inv_1 _1851_ (.Y(_0272_),
    .A(\autosel.i2c.i2c.delay_reg[6] ));
 sg13g2_a21o_1 _1852_ (.A2(_0223_),
    .A1(_0269_),
    .B1(_0272_),
    .X(_0273_));
 sg13g2_a21oi_1 _1853_ (.A1(_0271_),
    .A2(_0273_),
    .Y(_0117_),
    .B1(net26));
 sg13g2_nor2_1 _1854_ (.A(\autosel.i2c.i2c.delay_reg[6] ),
    .B(_0268_),
    .Y(_0274_));
 sg13g2_inv_1 _1855_ (.Y(_0275_),
    .A(\autosel.i2c.i2c.delay_reg[7] ));
 sg13g2_a21o_1 _1856_ (.A2(net12),
    .A1(_0274_),
    .B1(_0275_),
    .X(_0276_));
 sg13g2_nor3_1 _1857_ (.A(\autosel.i2c.i2c.delay_reg[6] ),
    .B(\autosel.i2c.i2c.delay_reg[7] ),
    .C(_0268_),
    .Y(_0277_));
 sg13g2_nand2_1 _1858_ (.Y(_0278_),
    .A(_0277_),
    .B(_0224_));
 sg13g2_a21oi_1 _1859_ (.A1(_0276_),
    .A2(_0278_),
    .Y(_0118_),
    .B1(_0230_));
 sg13g2_nand2_1 _1860_ (.Y(_0279_),
    .A(_0527_),
    .B(\autosel.i2c.i2c.delay_reg[8] ));
 sg13g2_a21oi_1 _1861_ (.A1(_0277_),
    .A2(net12),
    .Y(_0280_),
    .B1(_0279_));
 sg13g2_nand4_1 _1862_ (.B(_0779_),
    .C(net12),
    .A(_0530_),
    .Y(_0281_),
    .D(_0258_));
 sg13g2_nand2b_1 _1863_ (.Y(_0119_),
    .B(_0281_),
    .A_N(_0280_));
 sg13g2_nand2_1 _1864_ (.Y(_0282_),
    .A(\autosel.i2c.i2c.delay_reg[9] ),
    .B(_0232_));
 sg13g2_nor2_1 _1865_ (.A(\autosel.i2c.i2c.delay_reg[9] ),
    .B(_0232_),
    .Y(_0283_));
 sg13g2_nand2_1 _1866_ (.Y(_0284_),
    .A(_0781_),
    .B(_0283_));
 sg13g2_a21oi_1 _1867_ (.A1(_0282_),
    .A2(_0284_),
    .Y(_0120_),
    .B1(_0230_));
 sg13g2_nor2b_1 _1868_ (.A(net47),
    .B_N(_0667_),
    .Y(_0285_));
 sg13g2_nor2_1 _1869_ (.A(net39),
    .B(net28),
    .Y(_0286_));
 sg13g2_a22oi_1 _1870_ (.Y(_0287_),
    .B1(_0286_),
    .B2(net47),
    .A2(_0285_),
    .A1(_0782_));
 sg13g2_nor2_1 _1871_ (.A(_0221_),
    .B(_0287_),
    .Y(_0288_));
 sg13g2_nor2b_1 _1872_ (.A(\autosel.i2c.i2c.scl_i_reg ),
    .B_N(\autosel.i2c.i2c.scl_o_reg ),
    .Y(_0289_));
 sg13g2_a22oi_1 _1873_ (.Y(_0290_),
    .B1(_0289_),
    .B2(\autosel.i2c.i2c.delay_scl_reg ),
    .A2(_0288_),
    .A1(_0986_));
 sg13g2_nor2_1 _1874_ (.A(_0951_),
    .B(_0290_),
    .Y(_0121_));
 sg13g2_buf_1 _1875_ (.A(_0528_),
    .X(_0291_));
 sg13g2_inv_1 _1876_ (.Y(_0292_),
    .A(\autosel.i2c.i2c.delay_sda_reg ));
 sg13g2_a21oi_1 _1877_ (.A1(_0981_),
    .A2(\autosel.i2c.i2c.sda_o_reg ),
    .Y(_0293_),
    .B1(\autosel.i2c.i2c.delay_scl_reg ));
 sg13g2_nor3_1 _1878_ (.A(net25),
    .B(_0292_),
    .C(_0293_),
    .Y(_0122_));
 sg13g2_nand2b_1 _1879_ (.Y(_0294_),
    .B(net24),
    .A_N(_0037_));
 sg13g2_a21oi_1 _1880_ (.A1(_0765_),
    .A2(_0294_),
    .Y(_0131_),
    .B1(net26));
 sg13g2_nor2_1 _1881_ (.A(\autosel.i2c.i2c.delay_sda_reg ),
    .B(\autosel.i2c.i2c.delay_scl_reg ),
    .Y(_0295_));
 sg13g2_nand4_1 _1882_ (.B(_0773_),
    .C(_0779_),
    .A(_0772_),
    .Y(_0296_),
    .D(_0295_));
 sg13g2_buf_1 _1883_ (.A(_0296_),
    .X(_0297_));
 sg13g2_nand2b_1 _1884_ (.Y(_0298_),
    .B(net22),
    .A_N(net20));
 sg13g2_or2_1 _1885_ (.X(_0299_),
    .B(net20),
    .A(_0783_));
 sg13g2_inv_1 _1886_ (.Y(_0300_),
    .A(_0299_));
 sg13g2_nor2b_1 _1887_ (.A(net28),
    .B_N(net29),
    .Y(_0301_));
 sg13g2_o21ai_1 _1888_ (.B1(_0701_),
    .Y(_0302_),
    .A1(_0301_),
    .A2(_0211_));
 sg13g2_a221oi_1 _1889_ (.B2(_0302_),
    .C1(net25),
    .B1(_0300_),
    .A1(_0783_),
    .Y(_0136_),
    .A2(_0298_));
 sg13g2_nor2_1 _1890_ (.A(net22),
    .B(_0208_),
    .Y(_0303_));
 sg13g2_nand4_1 _1891_ (.B(_0987_),
    .C(_0988_),
    .A(_0688_),
    .Y(_0304_),
    .D(_0990_));
 sg13g2_nand2_1 _1892_ (.Y(_0305_),
    .A(_0989_),
    .B(_0669_));
 sg13g2_a21oi_1 _1893_ (.A1(_0995_),
    .A2(_0304_),
    .Y(_0306_),
    .B1(_0305_));
 sg13g2_or3_1 _1894_ (.A(net28),
    .B(_0303_),
    .C(_0306_),
    .X(_0307_));
 sg13g2_nand3_1 _1895_ (.B(_0300_),
    .C(_0307_),
    .A(_0701_),
    .Y(_0308_));
 sg13g2_nand2_1 _1896_ (.Y(_0309_),
    .A(_0666_),
    .B(_0299_));
 sg13g2_a21oi_1 _1897_ (.A1(_0308_),
    .A2(_0309_),
    .Y(_0137_),
    .B1(net26));
 sg13g2_nor2_1 _1898_ (.A(net39),
    .B(_0285_),
    .Y(_0310_));
 sg13g2_o21ai_1 _1899_ (.B1(net29),
    .Y(_0311_),
    .A1(net20),
    .A2(_0310_));
 sg13g2_a21oi_1 _1900_ (.A1(_0707_),
    .A2(_0216_),
    .Y(_0312_),
    .B1(_0218_));
 sg13g2_a21oi_1 _1901_ (.A1(_0208_),
    .A2(_0312_),
    .Y(_0313_),
    .B1(net28));
 sg13g2_or3_1 _1902_ (.A(net47),
    .B(net29),
    .C(_0313_),
    .X(_0314_));
 sg13g2_nand2b_1 _1903_ (.Y(_0315_),
    .B(net29),
    .A_N(_0285_));
 sg13g2_nand3_1 _1904_ (.B(_0314_),
    .C(_0315_),
    .A(net39),
    .Y(_0316_));
 sg13g2_nand2_1 _1905_ (.Y(_0317_),
    .A(_0783_),
    .B(_0306_));
 sg13g2_and2_1 _1906_ (.A(_0317_),
    .B(_0311_),
    .X(_0318_));
 sg13g2_a221oi_1 _1907_ (.B2(_0318_),
    .C1(_0291_),
    .B1(_0316_),
    .A1(net20),
    .Y(_0138_),
    .A2(_0311_));
 sg13g2_nor2b_1 _1908_ (.A(net28),
    .B_N(net20),
    .Y(_0319_));
 sg13g2_nor2_1 _1909_ (.A(_0701_),
    .B(_0783_),
    .Y(_0320_));
 sg13g2_nand3_1 _1910_ (.B(_0785_),
    .C(_0320_),
    .A(net28),
    .Y(_0321_));
 sg13g2_nor2_1 _1911_ (.A(_0297_),
    .B(_0321_),
    .Y(_0322_));
 sg13g2_a21o_1 _1912_ (.A2(_0219_),
    .A1(net34),
    .B1(_0214_),
    .X(_0323_));
 sg13g2_o21ai_1 _1913_ (.B1(_0786_),
    .Y(_0324_),
    .A1(net39),
    .A2(_0297_));
 sg13g2_a21oi_1 _1914_ (.A1(net39),
    .A2(_0785_),
    .Y(_0325_),
    .B1(_0786_));
 sg13g2_a21oi_1 _1915_ (.A1(_0701_),
    .A2(_0324_),
    .Y(_0326_),
    .B1(_0325_));
 sg13g2_a21oi_1 _1916_ (.A1(_0211_),
    .A2(_0323_),
    .Y(_0327_),
    .B1(_0326_));
 sg13g2_nor4_1 _1917_ (.A(_0528_),
    .B(_0319_),
    .C(_0322_),
    .D(_0327_),
    .Y(_0139_));
 sg13g2_nand2_1 _1918_ (.Y(_0328_),
    .A(_0701_),
    .B(net29));
 sg13g2_a22oi_1 _1919_ (.Y(_0329_),
    .B1(_0286_),
    .B2(_0328_),
    .A2(_0285_),
    .A1(net39));
 sg13g2_o21ai_1 _1920_ (.B1(net54),
    .Y(_0330_),
    .A1(net20),
    .A2(_0329_));
 sg13g2_xor2_1 _1921_ (.B(net29),
    .A(net28),
    .X(_0331_));
 sg13g2_a22oi_1 _1922_ (.Y(_0332_),
    .B1(_0320_),
    .B2(_0331_),
    .A2(_0301_),
    .A1(_0997_));
 sg13g2_o21ai_1 _1923_ (.B1(\autosel.i2c.i2c.scl_o_reg ),
    .Y(_0333_),
    .A1(net20),
    .A2(_0332_));
 sg13g2_nand2b_1 _1924_ (.Y(_0142_),
    .B(_0333_),
    .A_N(_0330_));
 sg13g2_nor2_1 _1925_ (.A(_0214_),
    .B(_0219_),
    .Y(_0334_));
 sg13g2_nand4_1 _1926_ (.B(_0783_),
    .C(_0667_),
    .A(net47),
    .Y(_0335_),
    .D(net29));
 sg13g2_nand2_1 _1927_ (.Y(_0336_),
    .A(_0702_),
    .B(_0784_));
 sg13g2_a221oi_1 _1928_ (.B2(_0336_),
    .C1(net20),
    .B1(_0335_),
    .A1(_0211_),
    .Y(_0337_),
    .A2(_0334_));
 sg13g2_nand2b_1 _1929_ (.Y(_0338_),
    .B(net34),
    .A_N(_0208_));
 sg13g2_o21ai_1 _1930_ (.B1(_0215_),
    .Y(_0339_),
    .A1(_0662_),
    .A2(_0658_));
 sg13g2_and2_1 _1931_ (.A(_0749_),
    .B(_0339_),
    .X(_0340_));
 sg13g2_nand3_1 _1932_ (.B(\autosel.i2c.i2c.data_reg[7] ),
    .C(_0728_),
    .A(_0732_),
    .Y(_0341_));
 sg13g2_nand4_1 _1933_ (.B(_0698_),
    .C(_0739_),
    .A(_0767_),
    .Y(_0342_),
    .D(_0204_));
 sg13g2_o21ai_1 _1934_ (.B1(_0342_),
    .Y(_0343_),
    .A1(_0212_),
    .A2(_0341_));
 sg13g2_nor2_1 _1935_ (.A(_0732_),
    .B(net40),
    .Y(_0344_));
 sg13g2_nand2_1 _1936_ (.Y(_0345_),
    .A(\autosel.i2c.i2c.mode_read_reg ),
    .B(net42));
 sg13g2_or2_1 _1937_ (.X(_0346_),
    .B(_0720_),
    .A(_0727_));
 sg13g2_nand3b_1 _1938_ (.B(_0727_),
    .C(_0720_),
    .Y(_0347_),
    .A_N(_0732_));
 sg13g2_nand2b_1 _1939_ (.Y(_0348_),
    .B(_0662_),
    .A_N(net42));
 sg13g2_a21o_1 _1940_ (.A2(_0347_),
    .A1(_0346_),
    .B1(_0348_),
    .X(_0349_));
 sg13g2_nand2b_1 _1941_ (.Y(_0350_),
    .B(_0733_),
    .A_N(_0346_));
 sg13g2_a221oi_1 _1942_ (.B2(_0350_),
    .C1(_0716_),
    .B1(_0349_),
    .A1(_0344_),
    .Y(_0351_),
    .A2(_0345_));
 sg13g2_mux4_1 _1943_ (.S0(net40),
    .A0(\autosel.i2c.i2c.data_reg[3] ),
    .A1(\autosel.i2c.i2c.data_reg[5] ),
    .A2(\autosel.i2c.i2c.data_reg[4] ),
    .A3(\autosel.i2c.i2c.data_reg[6] ),
    .S1(net42),
    .X(_0352_));
 sg13g2_nor2_1 _1944_ (.A(_0730_),
    .B(_0352_),
    .Y(_0353_));
 sg13g2_mux2_1 _1945_ (.A0(\autosel.i2c.i2c.data_reg[0] ),
    .A1(\autosel.i2c.i2c.data_reg[2] ),
    .S(net40),
    .X(_0354_));
 sg13g2_nor2b_1 _1946_ (.A(net42),
    .B_N(net40),
    .Y(_0355_));
 sg13g2_a221oi_1 _1947_ (.B2(\autosel.i2c.i2c.data_reg[1] ),
    .C1(_0727_),
    .B1(_0355_),
    .A1(net42),
    .Y(_0356_),
    .A2(_0354_));
 sg13g2_nor4_1 _1948_ (.A(_0732_),
    .B(_0212_),
    .C(_0353_),
    .D(_0356_),
    .Y(_0357_));
 sg13g2_nor4_1 _1949_ (.A(_0340_),
    .B(_0343_),
    .C(_0351_),
    .D(_0357_),
    .Y(_0358_));
 sg13g2_o21ai_1 _1950_ (.B1(_0702_),
    .Y(_0359_),
    .A1(_0995_),
    .A2(_0305_));
 sg13g2_nor4_1 _1951_ (.A(_0783_),
    .B(_0992_),
    .C(_0214_),
    .D(_0359_),
    .Y(_0360_));
 sg13g2_o21ai_1 _1952_ (.B1(_0360_),
    .Y(_0361_),
    .A1(_0338_),
    .A2(_0358_));
 sg13g2_nand2_1 _1953_ (.Y(_0362_),
    .A(_0702_),
    .B(_0320_));
 sg13g2_nand4_1 _1954_ (.B(_0337_),
    .C(_0361_),
    .A(_0317_),
    .Y(_0363_),
    .D(_0362_));
 sg13g2_nand2b_1 _1955_ (.Y(_0364_),
    .B(\autosel.i2c.i2c.sda_o_reg ),
    .A_N(_0337_));
 sg13g2_nand3_1 _1956_ (.B(_0363_),
    .C(_0364_),
    .A(net54),
    .Y(_0143_));
 sg13g2_a22oi_1 _1957_ (.Y(_0365_),
    .B1(_0994_),
    .B2(_0739_),
    .A2(_0753_),
    .A1(_0767_));
 sg13g2_nand2b_1 _1958_ (.Y(_0366_),
    .B(_0204_),
    .A_N(_0365_));
 sg13g2_nor2_1 _1959_ (.A(_0673_),
    .B(net30),
    .Y(_0367_));
 sg13g2_nor2_1 _1960_ (.A(_0035_),
    .B(_0215_),
    .Y(_0368_));
 sg13g2_nand3_1 _1961_ (.B(_0367_),
    .C(_0368_),
    .A(net41),
    .Y(_0369_));
 sg13g2_nand3_1 _1962_ (.B(_0217_),
    .C(_0369_),
    .A(_0821_),
    .Y(_0370_));
 sg13g2_nand2_1 _1963_ (.Y(_0371_),
    .A(_0749_),
    .B(_0368_));
 sg13g2_nand4_1 _1964_ (.B(_0366_),
    .C(_0370_),
    .A(_0696_),
    .Y(_0372_),
    .D(_0371_));
 sg13g2_nand2_1 _1965_ (.Y(_0373_),
    .A(_0744_),
    .B(_0712_));
 sg13g2_a22oi_1 _1966_ (.Y(_0374_),
    .B1(_0373_),
    .B2(net23),
    .A2(_0762_),
    .A1(net31));
 sg13g2_nor2b_1 _1967_ (.A(_0374_),
    .B_N(_0367_),
    .Y(_0375_));
 sg13g2_a21oi_1 _1968_ (.A1(net33),
    .A2(net32),
    .Y(_0376_),
    .B1(net31));
 sg13g2_nor2_1 _1969_ (.A(_0989_),
    .B(_0376_),
    .Y(_0377_));
 sg13g2_nor2_1 _1970_ (.A(net22),
    .B(_0377_),
    .Y(_0378_));
 sg13g2_o21ai_1 _1971_ (.B1(_0378_),
    .Y(_0379_),
    .A1(_0372_),
    .A2(_0375_));
 sg13g2_nand2_1 _1972_ (.Y(_0380_),
    .A(net33),
    .B(net22));
 sg13g2_a21oi_1 _1973_ (.A1(_0379_),
    .A2(_0380_),
    .Y(_0144_),
    .B1(_0291_));
 sg13g2_o21ai_1 _1974_ (.B1(net34),
    .Y(_0381_),
    .A1(_0989_),
    .A2(_0376_));
 sg13g2_nand2_1 _1975_ (.Y(_0382_),
    .A(\autosel.i2c.i2c.s_axis_data_tready_reg ),
    .B(_0791_));
 sg13g2_inv_1 _1976_ (.Y(_0383_),
    .A(_1006_));
 sg13g2_nor2_1 _1977_ (.A(_0671_),
    .B(_0683_),
    .Y(_0384_));
 sg13g2_nand3_1 _1978_ (.B(_0697_),
    .C(_0699_),
    .A(_0989_),
    .Y(_0385_));
 sg13g2_a22oi_1 _1979_ (.Y(_0386_),
    .B1(_0384_),
    .B2(_0385_),
    .A2(_0383_),
    .A1(_0382_));
 sg13g2_o21ai_1 _1980_ (.B1(net34),
    .Y(_0387_),
    .A1(_0381_),
    .A2(_0386_));
 sg13g2_nand2_1 _1981_ (.Y(_0388_),
    .A(_0820_),
    .B(net31));
 sg13g2_nand3_1 _1982_ (.B(_0744_),
    .C(\autosel.i2c.i2c.bus_active_reg ),
    .A(net32),
    .Y(_0389_));
 sg13g2_o21ai_1 _1983_ (.B1(_0389_),
    .Y(_0390_),
    .A1(_0762_),
    .A2(_0388_));
 sg13g2_o21ai_1 _1984_ (.B1(net23),
    .Y(_0391_),
    .A1(_0820_),
    .A2(_0744_));
 sg13g2_o21ai_1 _1985_ (.B1(_0391_),
    .Y(_0392_),
    .A1(net23),
    .A2(_0390_));
 sg13g2_nor4_1 _1986_ (.A(net33),
    .B(net32),
    .C(_0042_),
    .D(_0747_),
    .Y(_0393_));
 sg13g2_o21ai_1 _1987_ (.B1(_0689_),
    .Y(_0394_),
    .A1(_0708_),
    .A2(_0393_));
 sg13g2_o21ai_1 _1988_ (.B1(_0394_),
    .Y(_0395_),
    .A1(net30),
    .A2(_0392_));
 sg13g2_a22oi_1 _1989_ (.Y(_0396_),
    .B1(_0395_),
    .B2(_0378_),
    .A2(_0387_),
    .A1(net32));
 sg13g2_nor2_1 _1990_ (.A(net27),
    .B(_0396_),
    .Y(_0145_));
 sg13g2_nor4_1 _1991_ (.A(_0671_),
    .B(net32),
    .C(\autosel.i2c.i2c.bus_active_reg ),
    .D(_0747_),
    .Y(_0397_));
 sg13g2_nand2_1 _1992_ (.Y(_0398_),
    .A(_0821_),
    .B(_0993_));
 sg13g2_a21oi_1 _1993_ (.A1(_0398_),
    .A2(_0388_),
    .Y(_0399_),
    .B1(net30));
 sg13g2_a221oi_1 _1994_ (.B2(_0689_),
    .C1(_0399_),
    .B1(_0397_),
    .A1(_0699_),
    .Y(_0400_),
    .A2(_0749_));
 sg13g2_nand2_1 _1995_ (.Y(_0401_),
    .A(_0707_),
    .B(_0988_));
 sg13g2_nand3_1 _1996_ (.B(_0400_),
    .C(_0401_),
    .A(_0696_),
    .Y(_0402_));
 sg13g2_a22oi_1 _1997_ (.Y(_0403_),
    .B1(_0378_),
    .B2(_0402_),
    .A2(net22),
    .A1(net31));
 sg13g2_nor2_1 _1998_ (.A(net27),
    .B(_0403_),
    .Y(_0146_));
 sg13g2_a21oi_1 _1999_ (.A1(_0615_),
    .A2(_0616_),
    .Y(_0404_),
    .B1(_0622_));
 sg13g2_nor2b_1 _2000_ (.A(_0699_),
    .B_N(_0749_),
    .Y(_0405_));
 sg13g2_nand3_1 _2001_ (.B(_0739_),
    .C(_0762_),
    .A(net23),
    .Y(_0406_));
 sg13g2_o21ai_1 _2002_ (.B1(_0406_),
    .Y(_0407_),
    .A1(_0382_),
    .A2(_1006_));
 sg13g2_nand3_1 _2003_ (.B(\autosel.i2c.i2c.mode_read_reg ),
    .C(_0692_),
    .A(net32),
    .Y(_0408_));
 sg13g2_o21ai_1 _2004_ (.B1(_0739_),
    .Y(_0409_),
    .A1(_0820_),
    .A2(_0767_));
 sg13g2_a21oi_1 _2005_ (.A1(_0408_),
    .A2(_0409_),
    .Y(_0410_),
    .B1(net33));
 sg13g2_a221oi_1 _2006_ (.B2(net32),
    .C1(_0410_),
    .B1(_0407_),
    .A1(_0404_),
    .Y(_0411_),
    .A2(_0405_));
 sg13g2_nand2_1 _2007_ (.Y(_0412_),
    .A(_0685_),
    .B(_0703_));
 sg13g2_o21ai_1 _2008_ (.B1(_0412_),
    .Y(_0413_),
    .A1(_0381_),
    .A2(_0411_));
 sg13g2_and2_1 _2009_ (.A(net54),
    .B(_0413_),
    .X(_0147_));
 sg13g2_o21ai_1 _2010_ (.B1(\autosel.eeprom_data[15] ),
    .Y(_0414_),
    .A1(\autosel.eeprom_data[13] ),
    .A2(_0640_));
 sg13g2_nor3_1 _2011_ (.A(\autosel.eeprom_data[12] ),
    .B(_0638_),
    .C(_0640_),
    .Y(_0415_));
 sg13g2_a21o_1 _2012_ (.A2(_0640_),
    .A1(_0020_),
    .B1(_0415_),
    .X(_0416_));
 sg13g2_nor2b_1 _2013_ (.A(net37),
    .B_N(_0043_),
    .Y(_0417_));
 sg13g2_nor2_1 _2014_ (.A(_0927_),
    .B(_0417_),
    .Y(_0418_));
 sg13g2_nor2_1 _2015_ (.A(\debug_out.send_index[1] ),
    .B(_0921_),
    .Y(_0419_));
 sg13g2_nand2_1 _2016_ (.Y(_0420_),
    .A(net37),
    .B(_0043_));
 sg13g2_a22oi_1 _2017_ (.Y(_0421_),
    .B1(_0419_),
    .B2(_0420_),
    .A2(_0418_),
    .A1(net38));
 sg13g2_buf_1 _2018_ (.A(_0421_),
    .X(_0422_));
 sg13g2_a221oi_1 _2019_ (.B2(\autosel.eeprom_data[15] ),
    .C1(_0422_),
    .B1(_0416_),
    .A1(\autosel.eeprom_data[12] ),
    .Y(_0423_),
    .A2(_0414_));
 sg13g2_inv_1 _2020_ (.Y(_0424_),
    .A(_0812_));
 sg13g2_inv_1 _2021_ (.Y(_0425_),
    .A(\debug_out.send_index[1] ));
 sg13g2_nand2_1 _2022_ (.Y(_0426_),
    .A(_0425_),
    .B(_0930_));
 sg13g2_nand2_1 _2023_ (.Y(_0427_),
    .A(net38),
    .B(_0418_));
 sg13g2_o21ai_1 _2024_ (.B1(_0427_),
    .Y(_0428_),
    .A1(_0043_),
    .A2(_0426_));
 sg13g2_nor3_1 _2025_ (.A(_0424_),
    .B(_0841_),
    .C(_0428_),
    .Y(_0429_));
 sg13g2_buf_1 _2026_ (.A(_0429_),
    .X(_0430_));
 sg13g2_nand2_1 _2027_ (.Y(_0431_),
    .A(_0425_),
    .B(_0921_));
 sg13g2_or2_1 _2028_ (.X(_0432_),
    .B(_0431_),
    .A(net37));
 sg13g2_nand2_1 _2029_ (.Y(_0433_),
    .A(net38),
    .B(_0417_));
 sg13g2_nor2_2 _2030_ (.A(\autosel.eeprom_data[5] ),
    .B(\autosel.eeprom_data[6] ),
    .Y(_0434_));
 sg13g2_xnor2_1 _2031_ (.Y(_0435_),
    .A(\autosel.eeprom_data[4] ),
    .B(_0434_));
 sg13g2_nor2_1 _2032_ (.A(net48),
    .B(_0023_),
    .Y(_0436_));
 sg13g2_a21oi_1 _2033_ (.A1(net48),
    .A2(_0435_),
    .Y(_0437_),
    .B1(_0436_));
 sg13g2_or2_1 _2034_ (.X(_0438_),
    .B(_0437_),
    .A(_0433_));
 sg13g2_and2_1 _2035_ (.A(\debug_out.send_index[1] ),
    .B(_0927_),
    .X(_0439_));
 sg13g2_buf_1 _2036_ (.A(_0439_),
    .X(_0440_));
 sg13g2_nor2_1 _2037_ (.A(_0644_),
    .B(\autosel.eeprom_data[2] ),
    .Y(_0441_));
 sg13g2_xor2_1 _2038_ (.B(_0441_),
    .A(\autosel.eeprom_data[0] ),
    .X(_0442_));
 sg13g2_nor2b_1 _2039_ (.A(net49),
    .B_N(_0021_),
    .Y(_0443_));
 sg13g2_a21oi_1 _2040_ (.A1(net49),
    .A2(_0442_),
    .Y(_0444_),
    .B1(_0443_));
 sg13g2_nor2_2 _2041_ (.A(_0920_),
    .B(_0420_),
    .Y(_0445_));
 sg13g2_nor2_1 _2042_ (.A(_0655_),
    .B(\autosel.eeprom_data[10] ),
    .Y(_0446_));
 sg13g2_xor2_1 _2043_ (.B(_0446_),
    .A(\autosel.eeprom_data[8] ),
    .X(_0447_));
 sg13g2_nor2b_1 _2044_ (.A(_0635_),
    .B_N(_0025_),
    .Y(_0448_));
 sg13g2_a21oi_1 _2045_ (.A1(_0635_),
    .A2(_0447_),
    .Y(_0449_),
    .B1(_0448_));
 sg13g2_a22oi_1 _2046_ (.Y(_0450_),
    .B1(_0445_),
    .B2(_0449_),
    .A2(_0444_),
    .A1(_0440_));
 sg13g2_nand4_1 _2047_ (.B(_0432_),
    .C(_0438_),
    .A(_0422_),
    .Y(_0451_),
    .D(_0450_));
 sg13g2_nand3b_1 _2048_ (.B(net14),
    .C(_0451_),
    .Y(_0452_),
    .A_N(_0423_));
 sg13g2_nand2b_1 _2049_ (.Y(_0453_),
    .B(\debug_out.tx_byte[0] ),
    .A_N(net14));
 sg13g2_a21oi_1 _2050_ (.A1(_0452_),
    .A2(_0453_),
    .Y(_0186_),
    .B1(net25));
 sg13g2_nand2b_1 _2051_ (.Y(_0454_),
    .B(_0640_),
    .A_N(\autosel.eeprom_data[13] ));
 sg13g2_nor2b_1 _2052_ (.A(\autosel.eeprom_data[12] ),
    .B_N(\autosel.eeprom_data[15] ),
    .Y(_0455_));
 sg13g2_mux2_1 _2053_ (.A0(_0638_),
    .A1(_0454_),
    .S(_0455_),
    .X(_0456_));
 sg13g2_nor2_1 _2054_ (.A(_0043_),
    .B(_0456_),
    .Y(_0457_));
 sg13g2_nor2_1 _2055_ (.A(_0921_),
    .B(_0457_),
    .Y(_0458_));
 sg13g2_nor2_1 _2056_ (.A(net38),
    .B(_0458_),
    .Y(_0459_));
 sg13g2_o21ai_1 _2057_ (.B1(net37),
    .Y(_0460_),
    .A1(_0930_),
    .A2(_0456_));
 sg13g2_nor2_1 _2058_ (.A(\autosel.eeprom_data[4] ),
    .B(\autosel.eeprom_data[5] ),
    .Y(_0461_));
 sg13g2_and2_1 _2059_ (.A(\autosel.eeprom_data[4] ),
    .B(\autosel.eeprom_data[5] ),
    .X(_0462_));
 sg13g2_a21oi_1 _2060_ (.A1(\autosel.eeprom_data[6] ),
    .A2(_0461_),
    .Y(_0463_),
    .B1(_0462_));
 sg13g2_nor2b_1 _2061_ (.A(net48),
    .B_N(_0029_),
    .Y(_0464_));
 sg13g2_a21oi_1 _2062_ (.A1(net48),
    .A2(_0463_),
    .Y(_0465_),
    .B1(_0464_));
 sg13g2_a21oi_1 _2063_ (.A1(_0043_),
    .A2(_0465_),
    .Y(_0466_),
    .B1(_0457_));
 sg13g2_nor2_1 _2064_ (.A(_0426_),
    .B(_0456_),
    .Y(_0467_));
 sg13g2_nor2_1 _2065_ (.A(_0924_),
    .B(_0467_),
    .Y(_0468_));
 sg13g2_o21ai_1 _2066_ (.B1(_0468_),
    .Y(_0469_),
    .A1(_0425_),
    .A2(_0466_));
 sg13g2_o21ai_1 _2067_ (.B1(_0469_),
    .Y(_0470_),
    .A1(_0459_),
    .A2(_0460_));
 sg13g2_nor2_1 _2068_ (.A(\autosel.eeprom_data[8] ),
    .B(_0655_),
    .Y(_0471_));
 sg13g2_and2_1 _2069_ (.A(\autosel.eeprom_data[8] ),
    .B(_0655_),
    .X(_0472_));
 sg13g2_a21oi_1 _2070_ (.A1(\autosel.eeprom_data[10] ),
    .A2(_0471_),
    .Y(_0473_),
    .B1(_0472_));
 sg13g2_nor2b_1 _2071_ (.A(_0635_),
    .B_N(_0031_),
    .Y(_0474_));
 sg13g2_a21oi_1 _2072_ (.A1(_0635_),
    .A2(_0473_),
    .Y(_0475_),
    .B1(_0474_));
 sg13g2_nor2_1 _2073_ (.A(\autosel.eeprom_data[0] ),
    .B(_0644_),
    .Y(_0476_));
 sg13g2_and2_1 _2074_ (.A(\autosel.eeprom_data[0] ),
    .B(_0644_),
    .X(_0477_));
 sg13g2_a21oi_1 _2075_ (.A1(\autosel.eeprom_data[2] ),
    .A2(_0476_),
    .Y(_0478_),
    .B1(_0477_));
 sg13g2_nor2b_1 _2076_ (.A(net49),
    .B_N(_0027_),
    .Y(_0479_));
 sg13g2_a21oi_1 _2077_ (.A1(net49),
    .A2(_0478_),
    .Y(_0480_),
    .B1(_0479_));
 sg13g2_a22oi_1 _2078_ (.Y(_0481_),
    .B1(_0480_),
    .B2(_0440_),
    .A2(_0475_),
    .A1(_0445_));
 sg13g2_and2_1 _2079_ (.A(_0429_),
    .B(_0481_),
    .X(_0482_));
 sg13g2_o21ai_1 _2080_ (.B1(_0530_),
    .Y(_0483_),
    .A1(\debug_out.tx_byte[1] ),
    .A2(net14));
 sg13g2_a21oi_1 _2081_ (.A1(_0470_),
    .A2(_0482_),
    .Y(_0187_),
    .B1(_0483_));
 sg13g2_nor2_1 _2082_ (.A(\debug_out.tx_byte[2] ),
    .B(net14),
    .Y(_0484_));
 sg13g2_a21oi_1 _2083_ (.A1(_0635_),
    .A2(_0471_),
    .Y(_0485_),
    .B1(_0032_));
 sg13g2_nand2_1 _2084_ (.Y(_0486_),
    .A(_0445_),
    .B(_0485_));
 sg13g2_and2_1 _2085_ (.A(_0432_),
    .B(_0486_),
    .X(_0487_));
 sg13g2_a21oi_1 _2086_ (.A1(net48),
    .A2(_0461_),
    .Y(_0488_),
    .B1(_0030_));
 sg13g2_nand2b_1 _2087_ (.Y(_0489_),
    .B(_0488_),
    .A_N(_0433_));
 sg13g2_nand2_1 _2088_ (.Y(_0490_),
    .A(_0647_),
    .B(_0476_));
 sg13g2_nand3b_1 _2089_ (.B(_0440_),
    .C(_0490_),
    .Y(_0491_),
    .A_N(_0028_));
 sg13g2_and2_1 _2090_ (.A(_0489_),
    .B(_0491_),
    .X(_0492_));
 sg13g2_a21oi_1 _2091_ (.A1(_0638_),
    .A2(_0455_),
    .Y(_0493_),
    .B1(_0641_));
 sg13g2_nand2b_1 _2092_ (.Y(_0494_),
    .B(_0493_),
    .A_N(_0422_));
 sg13g2_and4_1 _2093_ (.A(_0429_),
    .B(_0487_),
    .C(_0492_),
    .D(_0494_),
    .X(_0495_));
 sg13g2_nor3_1 _2094_ (.A(net25),
    .B(_0484_),
    .C(_0495_),
    .Y(_0188_));
 sg13g2_nand2b_1 _2095_ (.Y(_0496_),
    .B(\debug_out.tx_byte[3] ),
    .A_N(_0430_));
 sg13g2_nand3_1 _2096_ (.B(_0445_),
    .C(_0446_),
    .A(_0635_),
    .Y(_0497_));
 sg13g2_nand4_1 _2097_ (.B(_0920_),
    .C(_0417_),
    .A(net48),
    .Y(_0498_),
    .D(_0434_));
 sg13g2_nand3_1 _2098_ (.B(_0440_),
    .C(_0441_),
    .A(net49),
    .Y(_0499_));
 sg13g2_nand4_1 _2099_ (.B(_0497_),
    .C(_0498_),
    .A(_0431_),
    .Y(_0500_),
    .D(_0499_));
 sg13g2_nor4_1 _2100_ (.A(\autosel.eeprom_data[13] ),
    .B(_0640_),
    .C(_0019_),
    .D(_0422_),
    .Y(_0501_));
 sg13g2_o21ai_1 _2101_ (.B1(net14),
    .Y(_0502_),
    .A1(_0500_),
    .A2(_0501_));
 sg13g2_a21oi_1 _2102_ (.A1(_0496_),
    .A2(_0502_),
    .Y(_0189_),
    .B1(net25));
 sg13g2_nand2b_1 _2103_ (.Y(_0503_),
    .B(\debug_out.tx_byte[4] ),
    .A_N(net14));
 sg13g2_nor2b_1 _2104_ (.A(_0434_),
    .B_N(net48),
    .Y(_0504_));
 sg13g2_o21ai_1 _2105_ (.B1(net49),
    .Y(_0505_),
    .A1(_0644_),
    .A2(\autosel.eeprom_data[2] ));
 sg13g2_o21ai_1 _2106_ (.B1(_0635_),
    .Y(_0506_),
    .A1(_0655_),
    .A2(\autosel.eeprom_data[10] ));
 sg13g2_a22oi_1 _2107_ (.Y(_0507_),
    .B1(_0506_),
    .B2(_0445_),
    .A2(_0505_),
    .A1(_0440_));
 sg13g2_o21ai_1 _2108_ (.B1(_0507_),
    .Y(_0508_),
    .A1(_0433_),
    .A2(_0504_));
 sg13g2_a21oi_1 _2109_ (.A1(_0638_),
    .A2(_0641_),
    .Y(_0509_),
    .B1(_0019_));
 sg13g2_nor2_1 _2110_ (.A(_0422_),
    .B(_0509_),
    .Y(_0510_));
 sg13g2_o21ai_1 _2111_ (.B1(net14),
    .Y(_0511_),
    .A1(_0508_),
    .A2(_0510_));
 sg13g2_a21oi_1 _2112_ (.A1(_0503_),
    .A2(_0511_),
    .Y(_0190_),
    .B1(net25));
 sg13g2_nor2_1 _2113_ (.A(_0026_),
    .B(_0446_),
    .Y(_0512_));
 sg13g2_nor2_1 _2114_ (.A(_0022_),
    .B(_0441_),
    .Y(_0513_));
 sg13g2_nor3_1 _2115_ (.A(_0024_),
    .B(_0433_),
    .C(_0434_),
    .Y(_0514_));
 sg13g2_a221oi_1 _2116_ (.B2(_0440_),
    .C1(_0514_),
    .B1(_0513_),
    .A1(_0445_),
    .Y(_0515_),
    .A2(_0512_));
 sg13g2_o21ai_1 _2117_ (.B1(_0515_),
    .Y(_0516_),
    .A1(_0422_),
    .A2(_0414_));
 sg13g2_nand2_1 _2118_ (.Y(_0517_),
    .A(net14),
    .B(_0516_));
 sg13g2_nand2b_1 _2119_ (.Y(_0518_),
    .B(\debug_out.tx_byte[6] ),
    .A_N(_0430_));
 sg13g2_a21oi_1 _2120_ (.A1(_0517_),
    .A2(_0518_),
    .Y(_0191_),
    .B1(net25));
 sg13g2_nand3b_1 _2121_ (.B(_0922_),
    .C(_0812_),
    .Y(_0519_),
    .A_N(_0841_));
 sg13g2_o21ai_1 _2122_ (.B1(\debug_out.tx_valid ),
    .Y(_0520_),
    .A1(_0424_),
    .A2(_0841_));
 sg13g2_a21oi_1 _2123_ (.A1(_0519_),
    .A2(_0520_),
    .Y(_0192_),
    .B1(net25));
 sg13g2_mux4_1 _2124_ (.S0(_0553_),
    .A0(\debug_out.uart_tx_inst.tx_data_latch[0] ),
    .A1(\debug_out.uart_tx_inst.tx_data_latch[1] ),
    .A2(\debug_out.uart_tx_inst.tx_data_latch[2] ),
    .A3(\debug_out.uart_tx_inst.tx_data_latch[3] ),
    .S1(_0552_),
    .X(_0521_));
 sg13g2_nand2b_1 _2125_ (.Y(_0522_),
    .B(\debug_out.uart_tx_inst.tx_data_latch[4] ),
    .A_N(_0552_));
 sg13g2_nand3b_1 _2126_ (.B(\debug_out.uart_tx_inst.tx_data_latch[6] ),
    .C(_0552_),
    .Y(_0523_),
    .A_N(_0553_));
 sg13g2_nand3_1 _2127_ (.B(_0522_),
    .C(_0523_),
    .A(\debug_out.uart_tx_inst.bit_cnt[2] ),
    .Y(_0524_));
 sg13g2_o21ai_1 _2128_ (.B1(_0524_),
    .Y(_0525_),
    .A1(\debug_out.uart_tx_inst.bit_cnt[2] ),
    .A2(_0521_));
 sg13g2_a21oi_1 _2129_ (.A1(_0561_),
    .A2(_0525_),
    .Y(_0526_),
    .B1(_0556_));
 sg13g2_nor2b_1 _2130_ (.A(_0526_),
    .B_N(_0559_),
    .Y(_0051_));
 sg13g2_buf_1 clkbuf_0_clk (.A(clk),
    .X(clknet_0_clk));
 sg13g2_tiehi \autosel.addr_counter[0]$_SDFFE_PN0P__81  (.L_HI(net81));
 sg13g2_buf_1 _2133_ (.A(\autosel.scl_oe ),
    .X(net4));
 sg13g2_buf_1 _2134_ (.A(\autosel.sda_oe ),
    .X(net5));
 sg13g2_buf_1 _2135_ (.A(net65),
    .X(uio_oe[2]));
 sg13g2_buf_1 _2136_ (.A(net66),
    .X(uio_oe[3]));
 sg13g2_buf_1 _2137_ (.A(net67),
    .X(uio_oe[4]));
 sg13g2_buf_1 _2138_ (.A(net68),
    .X(uio_oe[5]));
 sg13g2_buf_1 _2139_ (.A(net69),
    .X(uio_oe[6]));
 sg13g2_buf_1 _2140_ (.A(net70),
    .X(uio_oe[7]));
 sg13g2_buf_1 _2141_ (.A(\autosel.i2c.i2c.scl_o_reg ),
    .X(net6));
 sg13g2_buf_1 _2142_ (.A(\autosel.i2c.i2c.sda_o_reg ),
    .X(net7));
 sg13g2_buf_1 _2143_ (.A(net71),
    .X(uio_out[2]));
 sg13g2_buf_1 _2144_ (.A(net72),
    .X(uio_out[3]));
 sg13g2_buf_1 _2145_ (.A(net73),
    .X(uio_out[4]));
 sg13g2_buf_1 _2146_ (.A(net74),
    .X(uio_out[5]));
 sg13g2_buf_1 _2147_ (.A(net75),
    .X(uio_out[6]));
 sg13g2_buf_1 _2148_ (.A(net76),
    .X(uio_out[7]));
 sg13g2_buf_1 _2149_ (.A(\autosel.ctrl_sel_rst_n ),
    .X(net8));
 sg13g2_buf_1 _2150_ (.A(\autosel.ctrl_sel_inc ),
    .X(net9));
 sg13g2_buf_1 _2151_ (.A(\autosel.ctrl_ena ),
    .X(net10));
 sg13g2_buf_1 _2152_ (.A(net77),
    .X(uo_out[3]));
 sg13g2_buf_1 _2153_ (.A(\debug_out.uart_tx ),
    .X(net11));
 sg13g2_buf_1 _2154_ (.A(net78),
    .X(uo_out[5]));
 sg13g2_buf_1 _2155_ (.A(net79),
    .X(uo_out[6]));
 sg13g2_buf_1 _2156_ (.A(net80),
    .X(uo_out[7]));
 sg13g2_dfrbp_1 \autosel.addr_counter[0]$_SDFFE_PN0P_  (.CLK(clknet_5_29__leaf_clk),
    .RESET_B(net81),
    .D(_0052_),
    .Q_N(_0048_),
    .Q(\autosel.addr_counter[0] ));
 sg13g2_dfrbp_1 \autosel.addr_counter[1]$_SDFFE_PN0P_  (.CLK(clknet_5_28__leaf_clk),
    .RESET_B(net82),
    .D(_0053_),
    .Q_N(_1129_),
    .Q(\autosel.addr_counter[1] ));
 sg13g2_dfrbp_1 \autosel.addr_counter[2]$_SDFFE_PN0P_  (.CLK(clknet_5_29__leaf_clk),
    .RESET_B(net83),
    .D(_0054_),
    .Q_N(_1128_),
    .Q(\autosel.addr_counter[2] ));
 sg13g2_dfrbp_1 \autosel.addr_counter[3]$_SDFFE_PN0P_  (.CLK(clknet_5_28__leaf_clk),
    .RESET_B(net84),
    .D(_0055_),
    .Q_N(_1127_),
    .Q(\autosel.addr_counter[3] ));
 sg13g2_dfrbp_1 \autosel.addr_counter[4]$_SDFFE_PN0P_  (.CLK(clknet_5_25__leaf_clk),
    .RESET_B(net85),
    .D(_0056_),
    .Q_N(_1126_),
    .Q(\autosel.addr_counter[4] ));
 sg13g2_dfrbp_1 \autosel.addr_counter[5]$_SDFFE_PN0P_  (.CLK(clknet_5_19__leaf_clk),
    .RESET_B(net86),
    .D(_0057_),
    .Q_N(_1125_),
    .Q(\autosel.addr_counter[5] ));
 sg13g2_dfrbp_1 \autosel.addr_counter[6]$_SDFFE_PN0P_  (.CLK(clknet_5_19__leaf_clk),
    .RESET_B(net87),
    .D(_0058_),
    .Q_N(_1124_),
    .Q(\autosel.addr_counter[6] ));
 sg13g2_dfrbp_1 \autosel.addr_counter[7]$_SDFFE_PN0P_  (.CLK(clknet_5_22__leaf_clk),
    .RESET_B(net88),
    .D(_0059_),
    .Q_N(_1123_),
    .Q(\autosel.addr_counter[7] ));
 sg13g2_dfrbp_1 \autosel.addr_counter[8]$_SDFFE_PN0P_  (.CLK(clknet_5_22__leaf_clk),
    .RESET_B(net89),
    .D(_0060_),
    .Q_N(_1122_),
    .Q(\autosel.addr_counter[8] ));
 sg13g2_dfrbp_1 \autosel.addr_counter[9]$_SDFFE_PN0P_  (.CLK(clknet_5_23__leaf_clk),
    .RESET_B(net90),
    .D(_0061_),
    .Q_N(_1121_),
    .Q(\autosel.addr_counter[9] ));
 sg13g2_dfrbp_1 \autosel.ctrl_ena$_SDFFE_PN0P_  (.CLK(clknet_5_27__leaf_clk),
    .RESET_B(net91),
    .D(_0062_),
    .Q_N(_1120_),
    .Q(\autosel.ctrl_ena ));
 sg13g2_dfrbp_1 \autosel.ctrl_sel_inc$_SDFFE_PN0P_  (.CLK(clknet_5_25__leaf_clk),
    .RESET_B(net92),
    .D(_0063_),
    .Q_N(_0034_),
    .Q(\autosel.ctrl_sel_inc ));
 sg13g2_dfrbp_1 \autosel.ctrl_sel_rst_n$_SDFFE_PN0P_  (.CLK(clknet_5_26__leaf_clk),
    .RESET_B(net93),
    .D(_0064_),
    .Q_N(_1119_),
    .Q(\autosel.ctrl_sel_rst_n ));
 sg13g2_dfrbp_1 \autosel.i2c.busy$_DFFE_PN0P_  (.CLK(clknet_5_24__leaf_clk),
    .RESET_B(net59),
    .D(_0065_),
    .Q_N(_1118_),
    .Q(\autosel.eeprom_busy ));
 sg13g2_dfrbp_1 \autosel.i2c.data_out[0]$_DFFE_PN0P_  (.CLK(clknet_5_24__leaf_clk),
    .RESET_B(net59),
    .D(_0066_),
    .Q_N(_0021_),
    .Q(\autosel.eeprom_data[0] ));
 sg13g2_dfrbp_1 \autosel.i2c.data_out[10]$_DFFE_PN0P_  (.CLK(clknet_5_13__leaf_clk),
    .RESET_B(net57),
    .D(_0067_),
    .Q_N(_0032_),
    .Q(\autosel.eeprom_data[10] ));
 sg13g2_dfrbp_1 \autosel.i2c.data_out[11]$_DFFE_PN0P_  (.CLK(clknet_5_13__leaf_clk),
    .RESET_B(net57),
    .D(_0068_),
    .Q_N(_0026_),
    .Q(\autosel.eeprom_data[11] ));
 sg13g2_dfrbp_1 \autosel.i2c.data_out[12]$_DFFE_PN0P_  (.CLK(clknet_5_6__leaf_clk),
    .RESET_B(net56),
    .D(_0069_),
    .Q_N(_0020_),
    .Q(\autosel.eeprom_data[12] ));
 sg13g2_dfrbp_1 \autosel.i2c.data_out[13]$_DFFE_PN0P_  (.CLK(clknet_5_7__leaf_clk),
    .RESET_B(net56),
    .D(_0070_),
    .Q_N(_1117_),
    .Q(\autosel.eeprom_data[13] ));
 sg13g2_dfrbp_1 \autosel.i2c.data_out[14]$_DFFE_PN0P_  (.CLK(clknet_5_7__leaf_clk),
    .RESET_B(net56),
    .D(_0071_),
    .Q_N(_1116_),
    .Q(\autosel.eeprom_data[14] ));
 sg13g2_dfrbp_1 \autosel.i2c.data_out[15]$_DFFE_PN0P_  (.CLK(clknet_5_6__leaf_clk),
    .RESET_B(net56),
    .D(_0072_),
    .Q_N(_0019_),
    .Q(\autosel.eeprom_data[15] ));
 sg13g2_dfrbp_1 \autosel.i2c.data_out[1]$_DFFE_PN0P_  (.CLK(clknet_5_25__leaf_clk),
    .RESET_B(net59),
    .D(_0073_),
    .Q_N(_0027_),
    .Q(\autosel.eeprom_data[1] ));
 sg13g2_dfrbp_1 \autosel.i2c.data_out[2]$_DFFE_PN0P_  (.CLK(clknet_5_18__leaf_clk),
    .RESET_B(net59),
    .D(_0074_),
    .Q_N(_0028_),
    .Q(\autosel.eeprom_data[2] ));
 sg13g2_dfrbp_1 \autosel.i2c.data_out[3]$_DFFE_PN0P_  (.CLK(clknet_5_24__leaf_clk),
    .RESET_B(net57),
    .D(_0075_),
    .Q_N(_0022_),
    .Q(\autosel.eeprom_data[3] ));
 sg13g2_dfrbp_1 \autosel.i2c.data_out[4]$_DFFE_PN0P_  (.CLK(clknet_5_7__leaf_clk),
    .RESET_B(net57),
    .D(_0076_),
    .Q_N(_0023_),
    .Q(\autosel.eeprom_data[4] ));
 sg13g2_dfrbp_1 \autosel.i2c.data_out[5]$_DFFE_PN0P_  (.CLK(clknet_5_6__leaf_clk),
    .RESET_B(net57),
    .D(_0077_),
    .Q_N(_0029_),
    .Q(\autosel.eeprom_data[5] ));
 sg13g2_dfrbp_1 \autosel.i2c.data_out[6]$_DFFE_PN0P_  (.CLK(clknet_5_6__leaf_clk),
    .RESET_B(net57),
    .D(_0078_),
    .Q_N(_0030_),
    .Q(\autosel.eeprom_data[6] ));
 sg13g2_dfrbp_1 \autosel.i2c.data_out[7]$_DFFE_PN0P_  (.CLK(clknet_5_18__leaf_clk),
    .RESET_B(net57),
    .D(_0079_),
    .Q_N(_0024_),
    .Q(\autosel.eeprom_data[7] ));
 sg13g2_dfrbp_1 \autosel.i2c.data_out[8]$_DFFE_PN0P_  (.CLK(clknet_5_24__leaf_clk),
    .RESET_B(net58),
    .D(_0080_),
    .Q_N(_0025_),
    .Q(\autosel.eeprom_data[8] ));
 sg13g2_dfrbp_1 \autosel.i2c.data_out[9]$_DFFE_PN0P_  (.CLK(clknet_5_13__leaf_clk),
    .RESET_B(net57),
    .D(_0081_),
    .Q_N(_0031_),
    .Q(\autosel.eeprom_data[9] ));
 sg13g2_dfrbp_1 \autosel.i2c.data_out_hi[0]$_DFFE_PP_  (.CLK(clknet_5_13__leaf_clk),
    .RESET_B(net94),
    .D(_0082_),
    .Q_N(_1115_),
    .Q(\autosel.i2c.data_out_hi[0] ));
 sg13g2_dfrbp_1 \autosel.i2c.data_out_hi[1]$_DFFE_PP_  (.CLK(clknet_5_9__leaf_clk),
    .RESET_B(net95),
    .D(_0083_),
    .Q_N(_1114_),
    .Q(\autosel.i2c.data_out_hi[1] ));
 sg13g2_dfrbp_1 \autosel.i2c.data_out_hi[2]$_DFFE_PP_  (.CLK(clknet_5_13__leaf_clk),
    .RESET_B(net96),
    .D(_0084_),
    .Q_N(_1113_),
    .Q(\autosel.i2c.data_out_hi[2] ));
 sg13g2_dfrbp_1 \autosel.i2c.data_out_hi[3]$_DFFE_PP_  (.CLK(clknet_5_12__leaf_clk),
    .RESET_B(net97),
    .D(_0085_),
    .Q_N(_1112_),
    .Q(\autosel.i2c.data_out_hi[3] ));
 sg13g2_dfrbp_1 \autosel.i2c.data_out_hi[4]$_DFFE_PP_  (.CLK(clknet_5_3__leaf_clk),
    .RESET_B(net98),
    .D(_0086_),
    .Q_N(_1111_),
    .Q(\autosel.i2c.data_out_hi[4] ));
 sg13g2_dfrbp_1 \autosel.i2c.data_out_hi[5]$_DFFE_PP_  (.CLK(clknet_5_12__leaf_clk),
    .RESET_B(net99),
    .D(_0087_),
    .Q_N(_1110_),
    .Q(\autosel.i2c.data_out_hi[5] ));
 sg13g2_dfrbp_1 \autosel.i2c.data_out_hi[6]$_DFFE_PP_  (.CLK(clknet_5_9__leaf_clk),
    .RESET_B(net100),
    .D(_0088_),
    .Q_N(_1109_),
    .Q(\autosel.i2c.data_out_hi[6] ));
 sg13g2_dfrbp_1 \autosel.i2c.data_out_hi[7]$_DFFE_PP_  (.CLK(clknet_5_12__leaf_clk),
    .RESET_B(net101),
    .D(_0089_),
    .Q_N(_1108_),
    .Q(\autosel.i2c.data_out_hi[7] ));
 sg13g2_dfrbp_1 \autosel.i2c.i2c.addr_reg[4]$_DFFE_PP_  (.CLK(clknet_5_10__leaf_clk),
    .RESET_B(net102),
    .D(_0090_),
    .Q_N(_1107_),
    .Q(\autosel.i2c.i2c.addr_reg[4] ));
 sg13g2_dfrbp_1 \autosel.i2c.i2c.bit_count_reg[0]$_SDFFCE_PN0P_  (.CLK(clknet_5_10__leaf_clk),
    .RESET_B(net103),
    .D(_0091_),
    .Q_N(_0047_),
    .Q(\autosel.i2c.i2c.bit_count_reg[0] ));
 sg13g2_dfrbp_1 \autosel.i2c.i2c.bit_count_reg[1]$_SDFFCE_PN0P_  (.CLK(clknet_5_10__leaf_clk),
    .RESET_B(net104),
    .D(_0092_),
    .Q_N(_1106_),
    .Q(\autosel.i2c.i2c.bit_count_reg[1] ));
 sg13g2_dfrbp_1 \autosel.i2c.i2c.bit_count_reg[2]$_SDFFCE_PN0P_  (.CLK(clknet_5_10__leaf_clk),
    .RESET_B(net105),
    .D(_0093_),
    .Q_N(_1105_),
    .Q(\autosel.i2c.i2c.bit_count_reg[2] ));
 sg13g2_dfrbp_1 \autosel.i2c.i2c.bit_count_reg[3]$_SDFFCE_PN1P_  (.CLK(clknet_5_10__leaf_clk),
    .RESET_B(net106),
    .D(_0094_),
    .Q_N(_1104_),
    .Q(\autosel.i2c.i2c.bit_count_reg[3] ));
 sg13g2_dfrbp_1 \autosel.i2c.i2c.bus_active_reg$_SDFFE_PN0P_  (.CLK(clknet_5_15__leaf_clk),
    .RESET_B(net107),
    .D(_0095_),
    .Q_N(_0042_),
    .Q(\autosel.i2c.i2c.bus_active_reg ));
 sg13g2_dfrbp_1 \autosel.i2c.i2c.busy_reg$_SDFF_PN0_  (.CLK(clknet_5_15__leaf_clk),
    .RESET_B(net108),
    .D(_0096_),
    .Q_N(_0038_),
    .Q(\autosel.i2c.i2c.busy_reg ));
 sg13g2_dfrbp_1 \autosel.i2c.i2c.data_reg[0]$_SDFFCE_PN0P_  (.CLK(clknet_5_12__leaf_clk),
    .RESET_B(net109),
    .D(_0097_),
    .Q_N(_1103_),
    .Q(\autosel.i2c.i2c.data_reg[0] ));
 sg13g2_dfrbp_1 \autosel.i2c.i2c.data_reg[1]$_SDFFCE_PN0P_  (.CLK(clknet_5_11__leaf_clk),
    .RESET_B(net110),
    .D(_0098_),
    .Q_N(_1102_),
    .Q(\autosel.i2c.i2c.data_reg[1] ));
 sg13g2_dfrbp_1 \autosel.i2c.i2c.data_reg[2]$_SDFFCE_PN0P_  (.CLK(clknet_5_8__leaf_clk),
    .RESET_B(net111),
    .D(_0099_),
    .Q_N(_1101_),
    .Q(\autosel.i2c.i2c.data_reg[2] ));
 sg13g2_dfrbp_1 \autosel.i2c.i2c.data_reg[3]$_SDFFCE_PN0P_  (.CLK(clknet_5_8__leaf_clk),
    .RESET_B(net112),
    .D(_0100_),
    .Q_N(_1100_),
    .Q(\autosel.i2c.i2c.data_reg[3] ));
 sg13g2_dfrbp_1 \autosel.i2c.i2c.data_reg[4]$_SDFFCE_PN0P_  (.CLK(clknet_5_8__leaf_clk),
    .RESET_B(net113),
    .D(_0101_),
    .Q_N(_1099_),
    .Q(\autosel.i2c.i2c.data_reg[4] ));
 sg13g2_dfrbp_1 \autosel.i2c.i2c.data_reg[5]$_SDFFCE_PN0P_  (.CLK(clknet_5_8__leaf_clk),
    .RESET_B(net114),
    .D(_0102_),
    .Q_N(_1098_),
    .Q(\autosel.i2c.i2c.data_reg[5] ));
 sg13g2_dfrbp_1 \autosel.i2c.i2c.data_reg[6]$_SDFFCE_PN0P_  (.CLK(clknet_5_8__leaf_clk),
    .RESET_B(net115),
    .D(_0103_),
    .Q_N(_1097_),
    .Q(\autosel.i2c.i2c.data_reg[6] ));
 sg13g2_dfrbp_1 \autosel.i2c.i2c.data_reg[7]$_SDFFCE_PN0P_  (.CLK(clknet_5_10__leaf_clk),
    .RESET_B(net116),
    .D(_0104_),
    .Q_N(_1096_),
    .Q(\autosel.i2c.i2c.data_reg[7] ));
 sg13g2_dfrbp_1 \autosel.i2c.i2c.delay_reg[0]$_SDFFE_PN0P_  (.CLK(clknet_5_28__leaf_clk),
    .RESET_B(net117),
    .D(_0105_),
    .Q_N(_0044_),
    .Q(\autosel.i2c.i2c.delay_reg[0] ));
 sg13g2_dfrbp_1 \autosel.i2c.i2c.delay_reg[10]$_SDFFE_PN0P_  (.CLK(clknet_5_31__leaf_clk),
    .RESET_B(net118),
    .D(_0106_),
    .Q_N(_1095_),
    .Q(\autosel.i2c.i2c.delay_reg[10] ));
 sg13g2_dfrbp_1 \autosel.i2c.i2c.delay_reg[11]$_SDFFE_PN0P_  (.CLK(clknet_5_29__leaf_clk),
    .RESET_B(net119),
    .D(_0107_),
    .Q_N(_1094_),
    .Q(\autosel.i2c.i2c.delay_reg[11] ));
 sg13g2_dfrbp_1 \autosel.i2c.i2c.delay_reg[12]$_SDFFE_PN0P_  (.CLK(clknet_5_31__leaf_clk),
    .RESET_B(net120),
    .D(_0108_),
    .Q_N(_1093_),
    .Q(\autosel.i2c.i2c.delay_reg[12] ));
 sg13g2_dfrbp_1 \autosel.i2c.i2c.delay_reg[13]$_SDFFE_PN0P_  (.CLK(clknet_5_31__leaf_clk),
    .RESET_B(net121),
    .D(_0109_),
    .Q_N(_1092_),
    .Q(\autosel.i2c.i2c.delay_reg[13] ));
 sg13g2_dfrbp_1 \autosel.i2c.i2c.delay_reg[14]$_SDFFE_PN0P_  (.CLK(clknet_5_31__leaf_clk),
    .RESET_B(net122),
    .D(_0110_),
    .Q_N(_1091_),
    .Q(\autosel.i2c.i2c.delay_reg[14] ));
 sg13g2_dfrbp_1 \autosel.i2c.i2c.delay_reg[15]$_SDFFE_PN0P_  (.CLK(clknet_5_30__leaf_clk),
    .RESET_B(net123),
    .D(_0111_),
    .Q_N(_1090_),
    .Q(\autosel.i2c.i2c.delay_reg[15] ));
 sg13g2_dfrbp_1 \autosel.i2c.i2c.delay_reg[1]$_SDFFE_PN0P_  (.CLK(clknet_5_29__leaf_clk),
    .RESET_B(net124),
    .D(_0112_),
    .Q_N(_1089_),
    .Q(\autosel.i2c.i2c.delay_reg[1] ));
 sg13g2_dfrbp_1 \autosel.i2c.i2c.delay_reg[2]$_SDFFE_PN0P_  (.CLK(clknet_5_27__leaf_clk),
    .RESET_B(net125),
    .D(_0113_),
    .Q_N(_1088_),
    .Q(\autosel.i2c.i2c.delay_reg[2] ));
 sg13g2_dfrbp_1 \autosel.i2c.i2c.delay_reg[3]$_SDFFE_PN0P_  (.CLK(clknet_5_29__leaf_clk),
    .RESET_B(net126),
    .D(_0114_),
    .Q_N(_1087_),
    .Q(\autosel.i2c.i2c.delay_reg[3] ));
 sg13g2_dfrbp_1 \autosel.i2c.i2c.delay_reg[4]$_SDFFE_PN0P_  (.CLK(clknet_5_30__leaf_clk),
    .RESET_B(net127),
    .D(_0115_),
    .Q_N(_1086_),
    .Q(\autosel.i2c.i2c.delay_reg[4] ));
 sg13g2_dfrbp_1 \autosel.i2c.i2c.delay_reg[5]$_SDFFE_PN0P_  (.CLK(clknet_5_27__leaf_clk),
    .RESET_B(net128),
    .D(_0116_),
    .Q_N(_1085_),
    .Q(\autosel.i2c.i2c.delay_reg[5] ));
 sg13g2_dfrbp_1 \autosel.i2c.i2c.delay_reg[6]$_SDFFE_PN0P_  (.CLK(clknet_5_28__leaf_clk),
    .RESET_B(net129),
    .D(_0117_),
    .Q_N(_1084_),
    .Q(\autosel.i2c.i2c.delay_reg[6] ));
 sg13g2_dfrbp_1 \autosel.i2c.i2c.delay_reg[7]$_SDFFE_PN0P_  (.CLK(clknet_5_31__leaf_clk),
    .RESET_B(net130),
    .D(_0118_),
    .Q_N(_1083_),
    .Q(\autosel.i2c.i2c.delay_reg[7] ));
 sg13g2_dfrbp_1 \autosel.i2c.i2c.delay_reg[8]$_SDFFE_PN0P_  (.CLK(clknet_5_28__leaf_clk),
    .RESET_B(net131),
    .D(_0119_),
    .Q_N(_1082_),
    .Q(\autosel.i2c.i2c.delay_reg[8] ));
 sg13g2_dfrbp_1 \autosel.i2c.i2c.delay_reg[9]$_SDFFE_PN0P_  (.CLK(clknet_5_30__leaf_clk),
    .RESET_B(net132),
    .D(_0120_),
    .Q_N(_1081_),
    .Q(\autosel.i2c.i2c.delay_reg[9] ));
 sg13g2_dfrbp_1 \autosel.i2c.i2c.delay_scl_reg$_SDFF_PN0_  (.CLK(clknet_5_26__leaf_clk),
    .RESET_B(net133),
    .D(_0121_),
    .Q_N(_0039_),
    .Q(\autosel.i2c.i2c.delay_scl_reg ));
 sg13g2_dfrbp_1 \autosel.i2c.i2c.delay_sda_reg$_SDFFE_PN0N_  (.CLK(clknet_5_30__leaf_clk),
    .RESET_B(net134),
    .D(_0122_),
    .Q_N(_0041_),
    .Q(\autosel.i2c.i2c.delay_sda_reg ));
 sg13g2_dfrbp_1 \autosel.i2c.i2c.last_sda_i_reg$_DFF_P_  (.CLK(clknet_5_30__leaf_clk),
    .RESET_B(net135),
    .D(\autosel.i2c.i2c.sda_i_reg ),
    .Q_N(_1080_),
    .Q(\autosel.i2c.i2c.last_sda_i_reg ));
 sg13g2_dfrbp_1 \autosel.i2c.i2c.m_axis_data_tdata_reg[0]$_DFFE_PP_  (.CLK(clknet_5_12__leaf_clk),
    .RESET_B(net136),
    .D(_0123_),
    .Q_N(_1079_),
    .Q(\autosel.i2c.i2c.m_axis_data_tdata_reg[0] ));
 sg13g2_dfrbp_1 \autosel.i2c.i2c.m_axis_data_tdata_reg[1]$_DFFE_PP_  (.CLK(clknet_5_9__leaf_clk),
    .RESET_B(net137),
    .D(_0124_),
    .Q_N(_1078_),
    .Q(\autosel.i2c.i2c.m_axis_data_tdata_reg[1] ));
 sg13g2_dfrbp_1 \autosel.i2c.i2c.m_axis_data_tdata_reg[2]$_DFFE_PP_  (.CLK(clknet_5_9__leaf_clk),
    .RESET_B(net138),
    .D(_0125_),
    .Q_N(_1077_),
    .Q(\autosel.i2c.i2c.m_axis_data_tdata_reg[2] ));
 sg13g2_dfrbp_1 \autosel.i2c.i2c.m_axis_data_tdata_reg[3]$_DFFE_PP_  (.CLK(clknet_5_9__leaf_clk),
    .RESET_B(net139),
    .D(_0126_),
    .Q_N(_1076_),
    .Q(\autosel.i2c.i2c.m_axis_data_tdata_reg[3] ));
 sg13g2_dfrbp_1 \autosel.i2c.i2c.m_axis_data_tdata_reg[4]$_DFFE_PP_  (.CLK(clknet_5_3__leaf_clk),
    .RESET_B(net140),
    .D(_0127_),
    .Q_N(_1075_),
    .Q(\autosel.i2c.i2c.m_axis_data_tdata_reg[4] ));
 sg13g2_dfrbp_1 \autosel.i2c.i2c.m_axis_data_tdata_reg[5]$_DFFE_PP_  (.CLK(clknet_5_2__leaf_clk),
    .RESET_B(net141),
    .D(_0128_),
    .Q_N(_1074_),
    .Q(\autosel.i2c.i2c.m_axis_data_tdata_reg[5] ));
 sg13g2_dfrbp_1 \autosel.i2c.i2c.m_axis_data_tdata_reg[6]$_DFFE_PP_  (.CLK(clknet_5_8__leaf_clk),
    .RESET_B(net142),
    .D(_0129_),
    .Q_N(_1073_),
    .Q(\autosel.i2c.i2c.m_axis_data_tdata_reg[6] ));
 sg13g2_dfrbp_1 \autosel.i2c.i2c.m_axis_data_tdata_reg[7]$_DFFE_PP_  (.CLK(clknet_5_2__leaf_clk),
    .RESET_B(net143),
    .D(_0130_),
    .Q_N(_1072_),
    .Q(\autosel.i2c.i2c.m_axis_data_tdata_reg[7] ));
 sg13g2_dfrbp_1 \autosel.i2c.i2c.m_axis_data_tvalid_reg$_SDFF_PN0_  (.CLK(clknet_5_14__leaf_clk),
    .RESET_B(net144),
    .D(_0131_),
    .Q_N(_0037_),
    .Q(\autosel.i2c.i2c.m_axis_data_tvalid_reg ));
 sg13g2_dfrbp_1 \autosel.i2c.i2c.missed_ack_reg$_SDFF_PP0_  (.CLK(clknet_5_12__leaf_clk),
    .RESET_B(net145),
    .D(_0132_),
    .Q_N(_0036_),
    .Q(\autosel.i2c.i2c.missed_ack_reg ));
 sg13g2_dfrbp_1 \autosel.i2c.i2c.mode_read_reg$_DFFE_PP_  (.CLK(clknet_5_11__leaf_clk),
    .RESET_B(net146),
    .D(_0133_),
    .Q_N(_1071_),
    .Q(\autosel.i2c.i2c.mode_read_reg ));
 sg13g2_dfrbp_1 \autosel.i2c.i2c.mode_stop_reg$_DFFE_PP_  (.CLK(clknet_5_11__leaf_clk),
    .RESET_B(net147),
    .D(_0134_),
    .Q_N(_1070_),
    .Q(\autosel.i2c.i2c.mode_stop_reg ));
 sg13g2_dfrbp_1 \autosel.i2c.i2c.phy_rx_data_reg$_DFFE_PP_  (.CLK(clknet_5_27__leaf_clk),
    .RESET_B(net148),
    .D(_0135_),
    .Q_N(_1069_),
    .Q(\autosel.i2c.i2c.phy_rx_data_reg ));
 sg13g2_dfrbp_1 \autosel.i2c.i2c.phy_state_reg[0]$_SDFFE_PN0P_  (.CLK(clknet_5_26__leaf_clk),
    .RESET_B(net149),
    .D(_0136_),
    .Q_N(_1068_),
    .Q(\autosel.i2c.i2c.phy_state_reg[0] ));
 sg13g2_dfrbp_1 \autosel.i2c.i2c.phy_state_reg[1]$_SDFFE_PN0P_  (.CLK(clknet_5_26__leaf_clk),
    .RESET_B(net150),
    .D(_0137_),
    .Q_N(_1067_),
    .Q(\autosel.i2c.i2c.phy_state_reg[1] ));
 sg13g2_dfrbp_1 \autosel.i2c.i2c.phy_state_reg[2]$_SDFFE_PN0P_  (.CLK(clknet_5_24__leaf_clk),
    .RESET_B(net151),
    .D(_0138_),
    .Q_N(_1066_),
    .Q(\autosel.i2c.i2c.phy_state_reg[2] ));
 sg13g2_dfrbp_1 \autosel.i2c.i2c.phy_state_reg[3]$_SDFFE_PN0P_  (.CLK(clknet_5_27__leaf_clk),
    .RESET_B(net152),
    .D(_0139_),
    .Q_N(_1065_),
    .Q(\autosel.i2c.i2c.phy_state_reg[3] ));
 sg13g2_dfrbp_1 \autosel.i2c.i2c.s_axis_cmd_ready_reg$_SDFF_PP0_  (.CLK(clknet_5_11__leaf_clk),
    .RESET_B(net153),
    .D(_0140_),
    .Q_N(_0040_),
    .Q(\autosel.i2c.i2c.s_axis_cmd_ready_reg ));
 sg13g2_dfrbp_1 \autosel.i2c.i2c.s_axis_data_tready_reg$_SDFF_PP0_  (.CLK(clknet_5_14__leaf_clk),
    .RESET_B(net154),
    .D(_0141_),
    .Q_N(_1130_),
    .Q(\autosel.i2c.i2c.s_axis_data_tready_reg ));
 sg13g2_dfrbp_1 \autosel.i2c.i2c.scl_i_reg$_DFF_P_  (.CLK(clknet_5_30__leaf_clk),
    .RESET_B(net155),
    .D(net2),
    .Q_N(_1064_),
    .Q(\autosel.i2c.i2c.scl_i_reg ));
 sg13g2_dfrbp_1 \autosel.i2c.i2c.scl_o_reg$_SDFFE_PN1P_  (.CLK(clknet_5_26__leaf_clk),
    .RESET_B(net156),
    .D(_0142_),
    .Q_N(\autosel.scl_oe ),
    .Q(\autosel.i2c.i2c.scl_o_reg ));
 sg13g2_dfrbp_1 \autosel.i2c.i2c.sda_i_reg$_DFF_P_  (.CLK(clknet_5_26__leaf_clk),
    .RESET_B(net157),
    .D(net3),
    .Q_N(_1063_),
    .Q(\autosel.i2c.i2c.sda_i_reg ));
 sg13g2_dfrbp_1 \autosel.i2c.i2c.sda_o_reg$_SDFFE_PN1P_  (.CLK(clknet_5_15__leaf_clk),
    .RESET_B(net158),
    .D(_0143_),
    .Q_N(\autosel.sda_oe ),
    .Q(\autosel.i2c.i2c.sda_o_reg ));
 sg13g2_dfrbp_1 \autosel.i2c.i2c.state_reg[0]$_SDFFE_PN0N_  (.CLK(clknet_5_15__leaf_clk),
    .RESET_B(net159),
    .D(_0144_),
    .Q_N(_1062_),
    .Q(\autosel.i2c.i2c.state_reg[0] ));
 sg13g2_dfrbp_1 \autosel.i2c.i2c.state_reg[1]$_SDFFE_PN0N_  (.CLK(clknet_5_11__leaf_clk),
    .RESET_B(net160),
    .D(_0145_),
    .Q_N(_1061_),
    .Q(\autosel.i2c.i2c.state_reg[1] ));
 sg13g2_dfrbp_1 \autosel.i2c.i2c.state_reg[2]$_SDFFE_PN0N_  (.CLK(clknet_5_14__leaf_clk),
    .RESET_B(net161),
    .D(_0146_),
    .Q_N(_1060_),
    .Q(\autosel.i2c.i2c.state_reg[2] ));
 sg13g2_dfrbp_1 \autosel.i2c.i2c.state_reg[3]$_SDFFE_PN0N_  (.CLK(clknet_5_15__leaf_clk),
    .RESET_B(net162),
    .D(_0147_),
    .Q_N(_1059_),
    .Q(\autosel.i2c.i2c.state_reg[3] ));
 sg13g2_dfrbp_1 \autosel.i2c.state[0]$_DFFE_PN0P_  (.CLK(clknet_5_14__leaf_clk),
    .RESET_B(net58),
    .D(_0148_),
    .Q_N(_1058_),
    .Q(\autosel.i2c.state[0] ));
 sg13g2_dfrbp_1 \autosel.i2c.state[1]$_DFFE_PN0P_  (.CLK(clknet_5_14__leaf_clk),
    .RESET_B(net58),
    .D(_0149_),
    .Q_N(_1057_),
    .Q(\autosel.i2c.state[1] ));
 sg13g2_dfrbp_1 \autosel.i2c.state[2]$_DFFE_PN0P_  (.CLK(clknet_5_14__leaf_clk),
    .RESET_B(net58),
    .D(_0150_),
    .Q_N(_0035_),
    .Q(\autosel.i2c.state[2] ));
 sg13g2_dfrbp_1 \autosel.state[0]$_DFF_P_  (.CLK(clknet_5_25__leaf_clk),
    .RESET_B(net163),
    .D(net36),
    .Q_N(_1131_),
    .Q(\autosel.i2c.start ));
 sg13g2_dfrbp_1 \autosel.state[1]$_DFF_P_  (.CLK(clknet_5_25__leaf_clk),
    .RESET_B(net164),
    .D(_0001_),
    .Q_N(_1132_),
    .Q(\autosel.state[1] ));
 sg13g2_dfrbp_1 \autosel.state[2]$_DFF_P_  (.CLK(clknet_5_24__leaf_clk),
    .RESET_B(net165),
    .D(_0002_),
    .Q_N(_1056_),
    .Q(\autosel.state[2] ));
 sg13g2_dfrbp_1 \debug_out.counter[0]$_SDFF_PP0_  (.CLK(clknet_5_0__leaf_clk),
    .RESET_B(net166),
    .D(_0151_),
    .Q_N(_0049_),
    .Q(\debug_out.counter[0] ));
 sg13g2_dfrbp_1 \debug_out.counter[10]$_SDFF_PP0_  (.CLK(clknet_5_2__leaf_clk),
    .RESET_B(net167),
    .D(_0152_),
    .Q_N(_1055_),
    .Q(\debug_out.counter[10] ));
 sg13g2_dfrbp_1 \debug_out.counter[11]$_SDFF_PP0_  (.CLK(clknet_5_2__leaf_clk),
    .RESET_B(net168),
    .D(_0153_),
    .Q_N(_1054_),
    .Q(\debug_out.counter[11] ));
 sg13g2_dfrbp_1 \debug_out.counter[12]$_SDFF_PP0_  (.CLK(clknet_5_2__leaf_clk),
    .RESET_B(net169),
    .D(_0154_),
    .Q_N(_1053_),
    .Q(\debug_out.counter[12] ));
 sg13g2_dfrbp_1 \debug_out.counter[13]$_SDFF_PP0_  (.CLK(clknet_5_2__leaf_clk),
    .RESET_B(net170),
    .D(_0155_),
    .Q_N(_1052_),
    .Q(\debug_out.counter[13] ));
 sg13g2_dfrbp_1 \debug_out.counter[14]$_SDFF_PP0_  (.CLK(clknet_5_3__leaf_clk),
    .RESET_B(net171),
    .D(_0156_),
    .Q_N(_1051_),
    .Q(\debug_out.counter[14] ));
 sg13g2_dfrbp_1 \debug_out.counter[15]$_SDFF_PP0_  (.CLK(clknet_5_3__leaf_clk),
    .RESET_B(net172),
    .D(_0157_),
    .Q_N(_1050_),
    .Q(\debug_out.counter[15] ));
 sg13g2_dfrbp_1 \debug_out.counter[16]$_SDFF_PP0_  (.CLK(clknet_5_0__leaf_clk),
    .RESET_B(net173),
    .D(_0158_),
    .Q_N(_1049_),
    .Q(\debug_out.counter[16] ));
 sg13g2_dfrbp_1 \debug_out.counter[17]$_SDFF_PP0_  (.CLK(clknet_5_3__leaf_clk),
    .RESET_B(net174),
    .D(_0159_),
    .Q_N(_1048_),
    .Q(\debug_out.counter[17] ));
 sg13g2_dfrbp_1 \debug_out.counter[18]$_SDFF_PP0_  (.CLK(clknet_5_1__leaf_clk),
    .RESET_B(net175),
    .D(_0160_),
    .Q_N(_1047_),
    .Q(\debug_out.counter[18] ));
 sg13g2_dfrbp_1 \debug_out.counter[19]$_SDFF_PP0_  (.CLK(clknet_5_4__leaf_clk),
    .RESET_B(net176),
    .D(_0161_),
    .Q_N(_1046_),
    .Q(\debug_out.counter[19] ));
 sg13g2_dfrbp_1 \debug_out.counter[1]$_SDFF_PP0_  (.CLK(clknet_5_1__leaf_clk),
    .RESET_B(net177),
    .D(_0162_),
    .Q_N(_1045_),
    .Q(\debug_out.counter[1] ));
 sg13g2_dfrbp_1 \debug_out.counter[20]$_SDFF_PP0_  (.CLK(clknet_5_5__leaf_clk),
    .RESET_B(net178),
    .D(_0163_),
    .Q_N(_1044_),
    .Q(\debug_out.counter[20] ));
 sg13g2_dfrbp_1 \debug_out.counter[21]$_SDFF_PP0_  (.CLK(clknet_5_5__leaf_clk),
    .RESET_B(net179),
    .D(_0164_),
    .Q_N(_1043_),
    .Q(\debug_out.counter[21] ));
 sg13g2_dfrbp_1 \debug_out.counter[22]$_SDFF_PP0_  (.CLK(clknet_5_7__leaf_clk),
    .RESET_B(net180),
    .D(_0165_),
    .Q_N(_1042_),
    .Q(\debug_out.counter[22] ));
 sg13g2_dfrbp_1 \debug_out.counter[23]$_SDFF_PP0_  (.CLK(clknet_5_5__leaf_clk),
    .RESET_B(net181),
    .D(_0166_),
    .Q_N(_1041_),
    .Q(\debug_out.counter[23] ));
 sg13g2_dfrbp_1 \debug_out.counter[24]$_SDFF_PP0_  (.CLK(clknet_5_4__leaf_clk),
    .RESET_B(net182),
    .D(_0167_),
    .Q_N(_1040_),
    .Q(\debug_out.counter[24] ));
 sg13g2_dfrbp_1 \debug_out.counter[25]$_SDFF_PP0_  (.CLK(clknet_5_5__leaf_clk),
    .RESET_B(net183),
    .D(_0168_),
    .Q_N(_1039_),
    .Q(\debug_out.counter[25] ));
 sg13g2_dfrbp_1 \debug_out.counter[26]$_SDFF_PP0_  (.CLK(clknet_5_4__leaf_clk),
    .RESET_B(net184),
    .D(_0169_),
    .Q_N(_1038_),
    .Q(\debug_out.counter[26] ));
 sg13g2_dfrbp_1 \debug_out.counter[27]$_SDFF_PP0_  (.CLK(clknet_5_4__leaf_clk),
    .RESET_B(net185),
    .D(_0170_),
    .Q_N(_1037_),
    .Q(\debug_out.counter[27] ));
 sg13g2_dfrbp_1 \debug_out.counter[28]$_SDFF_PP0_  (.CLK(clknet_5_4__leaf_clk),
    .RESET_B(net186),
    .D(_0171_),
    .Q_N(_1036_),
    .Q(\debug_out.counter[28] ));
 sg13g2_dfrbp_1 \debug_out.counter[29]$_SDFF_PP0_  (.CLK(clknet_5_4__leaf_clk),
    .RESET_B(net187),
    .D(_0172_),
    .Q_N(_1035_),
    .Q(\debug_out.counter[29] ));
 sg13g2_dfrbp_1 \debug_out.counter[2]$_SDFF_PP0_  (.CLK(clknet_5_1__leaf_clk),
    .RESET_B(net188),
    .D(_0173_),
    .Q_N(_1034_),
    .Q(\debug_out.counter[2] ));
 sg13g2_dfrbp_1 \debug_out.counter[30]$_SDFF_PP0_  (.CLK(clknet_5_1__leaf_clk),
    .RESET_B(net189),
    .D(_0174_),
    .Q_N(_1033_),
    .Q(\debug_out.counter[30] ));
 sg13g2_dfrbp_1 \debug_out.counter[31]$_SDFF_PP0_  (.CLK(clknet_5_1__leaf_clk),
    .RESET_B(net190),
    .D(_0175_),
    .Q_N(_1032_),
    .Q(\debug_out.counter[31] ));
 sg13g2_dfrbp_1 \debug_out.counter[3]$_SDFF_PP0_  (.CLK(clknet_5_0__leaf_clk),
    .RESET_B(net191),
    .D(_0176_),
    .Q_N(_1031_),
    .Q(\debug_out.counter[3] ));
 sg13g2_dfrbp_1 \debug_out.counter[4]$_SDFF_PP0_  (.CLK(clknet_5_0__leaf_clk),
    .RESET_B(net192),
    .D(_0177_),
    .Q_N(_1030_),
    .Q(\debug_out.counter[4] ));
 sg13g2_dfrbp_1 \debug_out.counter[5]$_SDFF_PP0_  (.CLK(clknet_5_0__leaf_clk),
    .RESET_B(net193),
    .D(_0178_),
    .Q_N(_1029_),
    .Q(\debug_out.counter[5] ));
 sg13g2_dfrbp_1 \debug_out.counter[6]$_SDFF_PP0_  (.CLK(clknet_5_0__leaf_clk),
    .RESET_B(net194),
    .D(_0179_),
    .Q_N(_1028_),
    .Q(\debug_out.counter[6] ));
 sg13g2_dfrbp_1 \debug_out.counter[7]$_SDFF_PP0_  (.CLK(clknet_5_1__leaf_clk),
    .RESET_B(net195),
    .D(_0180_),
    .Q_N(_1027_),
    .Q(\debug_out.counter[7] ));
 sg13g2_dfrbp_1 \debug_out.counter[8]$_SDFF_PP0_  (.CLK(clknet_5_6__leaf_clk),
    .RESET_B(net196),
    .D(_0181_),
    .Q_N(_1026_),
    .Q(\debug_out.counter[8] ));
 sg13g2_dfrbp_1 \debug_out.counter[9]$_SDFF_PP0_  (.CLK(clknet_5_6__leaf_clk),
    .RESET_B(net197),
    .D(_0182_),
    .Q_N(_1025_),
    .Q(\debug_out.counter[9] ));
 sg13g2_dfrbp_1 \debug_out.send_index[0]$_SDFFE_PP0P_  (.CLK(clknet_5_16__leaf_clk),
    .RESET_B(net198),
    .D(_0183_),
    .Q_N(_0050_),
    .Q(\debug_out.send_index[0] ));
 sg13g2_dfrbp_1 \debug_out.send_index[1]$_SDFFE_PP0P_  (.CLK(clknet_5_16__leaf_clk),
    .RESET_B(net199),
    .D(_0184_),
    .Q_N(_1024_),
    .Q(\debug_out.send_index[1] ));
 sg13g2_dfrbp_1 \debug_out.send_index[2]$_SDFFE_PP0P_  (.CLK(clknet_5_7__leaf_clk),
    .RESET_B(net200),
    .D(_0185_),
    .Q_N(_0043_),
    .Q(\debug_out.send_index[2] ));
 sg13g2_dfrbp_1 \debug_out.tx_byte[0]$_SDFFE_PN0P_  (.CLK(clknet_5_18__leaf_clk),
    .RESET_B(net201),
    .D(_0186_),
    .Q_N(_1023_),
    .Q(\debug_out.tx_byte[0] ));
 sg13g2_dfrbp_1 \debug_out.tx_byte[1]$_SDFFE_PN0P_  (.CLK(clknet_5_18__leaf_clk),
    .RESET_B(net202),
    .D(_0187_),
    .Q_N(_1022_),
    .Q(\debug_out.tx_byte[1] ));
 sg13g2_dfrbp_1 \debug_out.tx_byte[2]$_SDFFE_PN0P_  (.CLK(clknet_5_22__leaf_clk),
    .RESET_B(net203),
    .D(_0188_),
    .Q_N(_1021_),
    .Q(\debug_out.tx_byte[2] ));
 sg13g2_dfrbp_1 \debug_out.tx_byte[3]$_SDFFE_PN0P_  (.CLK(clknet_5_19__leaf_clk),
    .RESET_B(net204),
    .D(_0189_),
    .Q_N(_1020_),
    .Q(\debug_out.tx_byte[3] ));
 sg13g2_dfrbp_1 \debug_out.tx_byte[5]$_SDFFE_PN0P_  (.CLK(clknet_5_18__leaf_clk),
    .RESET_B(net205),
    .D(_0190_),
    .Q_N(_1019_),
    .Q(\debug_out.tx_byte[4] ));
 sg13g2_dfrbp_1 \debug_out.tx_byte[6]$_SDFFE_PN0P_  (.CLK(clknet_5_19__leaf_clk),
    .RESET_B(net206),
    .D(_0191_),
    .Q_N(_1018_),
    .Q(\debug_out.tx_byte[6] ));
 sg13g2_dfrbp_1 \debug_out.tx_valid$_SDFFE_PN0P_  (.CLK(clknet_5_18__leaf_clk),
    .RESET_B(net207),
    .D(_0192_),
    .Q_N(_1017_),
    .Q(\debug_out.tx_valid ));
 sg13g2_dfrbp_1 \debug_out.uart_tx_inst.bit_cnt[0]$_DFFE_PN0P_  (.CLK(clknet_5_23__leaf_clk),
    .RESET_B(net61),
    .D(_0193_),
    .Q_N(_1016_),
    .Q(\debug_out.uart_tx_inst.bit_cnt[0] ));
 sg13g2_dfrbp_1 \debug_out.uart_tx_inst.bit_cnt[1]$_DFFE_PN0P_  (.CLK(clknet_5_23__leaf_clk),
    .RESET_B(net63),
    .D(_0194_),
    .Q_N(_1015_),
    .Q(\debug_out.uart_tx_inst.bit_cnt[1] ));
 sg13g2_dfrbp_1 \debug_out.uart_tx_inst.bit_cnt[2]$_DFFE_PN0P_  (.CLK(clknet_5_21__leaf_clk),
    .RESET_B(net63),
    .D(_0195_),
    .Q_N(_0046_),
    .Q(\debug_out.uart_tx_inst.bit_cnt[2] ));
 sg13g2_dfrbp_1 \debug_out.uart_tx_inst.cycle_cnt[0]$_DFF_PN0_  (.CLK(clknet_5_17__leaf_clk),
    .RESET_B(net56),
    .D(_0003_),
    .Q_N(_1133_),
    .Q(\debug_out.uart_tx_inst.cycle_cnt[0] ));
 sg13g2_dfrbp_1 \debug_out.uart_tx_inst.cycle_cnt[10]$_DFF_PN0_  (.CLK(clknet_5_20__leaf_clk),
    .RESET_B(net62),
    .D(_0004_),
    .Q_N(_1134_),
    .Q(\debug_out.uart_tx_inst.cycle_cnt[10] ));
 sg13g2_dfrbp_1 \debug_out.uart_tx_inst.cycle_cnt[11]$_DFF_PN0_  (.CLK(clknet_5_20__leaf_clk),
    .RESET_B(net61),
    .D(_0005_),
    .Q_N(_1135_),
    .Q(\debug_out.uart_tx_inst.cycle_cnt[11] ));
 sg13g2_dfrbp_1 \debug_out.uart_tx_inst.cycle_cnt[12]$_DFF_PN0_  (.CLK(clknet_5_20__leaf_clk),
    .RESET_B(net61),
    .D(_0006_),
    .Q_N(_1136_),
    .Q(\debug_out.uart_tx_inst.cycle_cnt[12] ));
 sg13g2_dfrbp_1 \debug_out.uart_tx_inst.cycle_cnt[13]$_DFF_PN0_  (.CLK(clknet_5_21__leaf_clk),
    .RESET_B(net61),
    .D(_0007_),
    .Q_N(_1137_),
    .Q(\debug_out.uart_tx_inst.cycle_cnt[13] ));
 sg13g2_dfrbp_1 \debug_out.uart_tx_inst.cycle_cnt[14]$_DFF_PN0_  (.CLK(clknet_5_21__leaf_clk),
    .RESET_B(net61),
    .D(_0008_),
    .Q_N(_1138_),
    .Q(\debug_out.uart_tx_inst.cycle_cnt[14] ));
 sg13g2_dfrbp_1 \debug_out.uart_tx_inst.cycle_cnt[15]$_DFF_PN0_  (.CLK(clknet_5_21__leaf_clk),
    .RESET_B(net61),
    .D(_0009_),
    .Q_N(_1139_),
    .Q(\debug_out.uart_tx_inst.cycle_cnt[15] ));
 sg13g2_dfrbp_1 \debug_out.uart_tx_inst.cycle_cnt[1]$_DFF_PN0_  (.CLK(clknet_5_17__leaf_clk),
    .RESET_B(net62),
    .D(_0010_),
    .Q_N(_1140_),
    .Q(\debug_out.uart_tx_inst.cycle_cnt[1] ));
 sg13g2_dfrbp_1 \debug_out.uart_tx_inst.cycle_cnt[2]$_DFF_PN0_  (.CLK(clknet_5_16__leaf_clk),
    .RESET_B(net56),
    .D(_0011_),
    .Q_N(_1141_),
    .Q(\debug_out.uart_tx_inst.cycle_cnt[2] ));
 sg13g2_dfrbp_1 \debug_out.uart_tx_inst.cycle_cnt[3]$_DFF_PN0_  (.CLK(clknet_5_16__leaf_clk),
    .RESET_B(net60),
    .D(_0012_),
    .Q_N(_1142_),
    .Q(\debug_out.uart_tx_inst.cycle_cnt[3] ));
 sg13g2_dfrbp_1 \debug_out.uart_tx_inst.cycle_cnt[4]$_DFF_PN0_  (.CLK(clknet_5_16__leaf_clk),
    .RESET_B(net56),
    .D(_0013_),
    .Q_N(_1143_),
    .Q(\debug_out.uart_tx_inst.cycle_cnt[4] ));
 sg13g2_dfrbp_1 \debug_out.uart_tx_inst.cycle_cnt[5]$_DFF_PN0_  (.CLK(clknet_5_5__leaf_clk),
    .RESET_B(net56),
    .D(_0014_),
    .Q_N(_1144_),
    .Q(\debug_out.uart_tx_inst.cycle_cnt[5] ));
 sg13g2_dfrbp_1 \debug_out.uart_tx_inst.cycle_cnt[6]$_DFF_PN0_  (.CLK(clknet_5_16__leaf_clk),
    .RESET_B(net60),
    .D(_0015_),
    .Q_N(_1145_),
    .Q(\debug_out.uart_tx_inst.cycle_cnt[6] ));
 sg13g2_dfrbp_1 \debug_out.uart_tx_inst.cycle_cnt[7]$_DFF_PN0_  (.CLK(clknet_5_17__leaf_clk),
    .RESET_B(net62),
    .D(_0016_),
    .Q_N(_1146_),
    .Q(\debug_out.uart_tx_inst.cycle_cnt[7] ));
 sg13g2_dfrbp_1 \debug_out.uart_tx_inst.cycle_cnt[8]$_DFF_PN0_  (.CLK(clknet_5_17__leaf_clk),
    .RESET_B(net62),
    .D(_0017_),
    .Q_N(_1147_),
    .Q(\debug_out.uart_tx_inst.cycle_cnt[8] ));
 sg13g2_dfrbp_1 \debug_out.uart_tx_inst.cycle_cnt[9]$_DFF_PN0_  (.CLK(clknet_5_20__leaf_clk),
    .RESET_B(net62),
    .D(_0018_),
    .Q_N(_1014_),
    .Q(\debug_out.uart_tx_inst.cycle_cnt[9] ));
 sg13g2_dfrbp_1 \debug_out.uart_tx_inst.state[0]$_DFF_PN1_  (.CLK(clknet_5_21__leaf_clk),
    .RESET_B(net61),
    .D(_0045_),
    .Q_N(\debug_out.uart_tx_inst.state[0] ),
    .Q(_1149_));
 sg13g2_dfrbp_1 \debug_out.uart_tx_inst.state[1]$_DFF_PN0_  (.CLK(clknet_5_19__leaf_clk),
    .RESET_B(net62),
    .D(\debug_out.uart_tx_inst.next_state[1] ),
    .Q_N(_1148_),
    .Q(\debug_out.uart_tx_inst.state[1] ));
 sg13g2_dfrbp_1 \debug_out.uart_tx_inst.state[2]$_DFF_PN0_  (.CLK(clknet_5_20__leaf_clk),
    .RESET_B(net61),
    .D(\debug_out.uart_tx_inst.next_state[2] ),
    .Q_N(_0033_),
    .Q(\debug_out.uart_tx_inst.state[2] ));
 sg13g2_dfrbp_1 \debug_out.uart_tx_inst.tx_data_latch[0]$_DFFE_PN0P_  (.CLK(clknet_5_22__leaf_clk),
    .RESET_B(net64),
    .D(_0196_),
    .Q_N(_1013_),
    .Q(\debug_out.uart_tx_inst.tx_data_latch[0] ));
 sg13g2_dfrbp_1 \debug_out.uart_tx_inst.tx_data_latch[1]$_DFFE_PN0P_  (.CLK(clknet_5_22__leaf_clk),
    .RESET_B(net64),
    .D(_0197_),
    .Q_N(_1012_),
    .Q(\debug_out.uart_tx_inst.tx_data_latch[1] ));
 sg13g2_dfrbp_1 \debug_out.uart_tx_inst.tx_data_latch[2]$_DFFE_PN0P_  (.CLK(clknet_5_23__leaf_clk),
    .RESET_B(net64),
    .D(_0198_),
    .Q_N(_1011_),
    .Q(\debug_out.uart_tx_inst.tx_data_latch[2] ));
 sg13g2_dfrbp_1 \debug_out.uart_tx_inst.tx_data_latch[3]$_DFFE_PN0P_  (.CLK(clknet_5_23__leaf_clk),
    .RESET_B(net64),
    .D(_0199_),
    .Q_N(_1010_),
    .Q(\debug_out.uart_tx_inst.tx_data_latch[3] ));
 sg13g2_dfrbp_1 \debug_out.uart_tx_inst.tx_data_latch[5]$_DFFE_PN0P_  (.CLK(clknet_5_20__leaf_clk),
    .RESET_B(net62),
    .D(_0200_),
    .Q_N(_1009_),
    .Q(\debug_out.uart_tx_inst.tx_data_latch[4] ));
 sg13g2_dfrbp_1 \debug_out.uart_tx_inst.tx_data_latch[6]$_DFFE_PN0P_  (.CLK(clknet_5_22__leaf_clk),
    .RESET_B(net63),
    .D(_0201_),
    .Q_N(_1008_),
    .Q(\debug_out.uart_tx_inst.tx_data_latch[6] ));
 sg13g2_dfrbp_1 \debug_out.uart_tx_inst.tx_data_ready$_DFFE_PN0P_  (.CLK(clknet_5_17__leaf_clk),
    .RESET_B(net62),
    .D(_0202_),
    .Q_N(_1007_),
    .Q(\debug_out.tx_ready ));
 sg13g2_dfrbp_1 \debug_out.uart_tx_inst.tx_reg$_DFF_PN1_  (.CLK(clknet_5_28__leaf_clk),
    .RESET_B(net64),
    .D(_0051_),
    .Q_N(\debug_out.uart_tx ),
    .Q(_1150_));
 sg13g2_buf_1 input1 (.A(rst_n),
    .X(net1));
 sg13g2_buf_1 input2 (.A(uio_in[0]),
    .X(net2));
 sg13g2_buf_1 input3 (.A(uio_in[1]),
    .X(net3));
 sg13g2_buf_1 output4 (.A(net4),
    .X(uio_oe[0]));
 sg13g2_buf_1 output5 (.A(net5),
    .X(uio_oe[1]));
 sg13g2_buf_1 output6 (.A(net6),
    .X(uio_out[0]));
 sg13g2_buf_1 output7 (.A(net7),
    .X(uio_out[1]));
 sg13g2_buf_1 output8 (.A(net8),
    .X(uo_out[0]));
 sg13g2_buf_1 output9 (.A(net9),
    .X(uo_out[1]));
 sg13g2_buf_1 output10 (.A(net10),
    .X(uo_out[2]));
 sg13g2_buf_1 output11 (.A(net11),
    .X(uo_out[4]));
 sg13g2_buf_2 fanout12 (.A(_0224_),
    .X(net12));
 sg13g2_buf_2 fanout13 (.A(_0582_),
    .X(net13));
 sg13g2_buf_2 fanout14 (.A(_0430_),
    .X(net14));
 sg13g2_buf_2 fanout15 (.A(_0896_),
    .X(net15));
 sg13g2_buf_2 fanout16 (.A(_0872_),
    .X(net16));
 sg13g2_buf_2 fanout17 (.A(_0844_),
    .X(net17));
 sg13g2_buf_2 fanout18 (.A(_0765_),
    .X(net18));
 sg13g2_buf_2 fanout19 (.A(_0633_),
    .X(net19));
 sg13g2_buf_2 fanout20 (.A(_0297_),
    .X(net20));
 sg13g2_buf_2 fanout21 (.A(_0632_),
    .X(net21));
 sg13g2_buf_2 fanout22 (.A(_0703_),
    .X(net22));
 sg13g2_buf_2 fanout23 (.A(_0682_),
    .X(net23));
 sg13g2_buf_2 fanout24 (.A(_0658_),
    .X(net24));
 sg13g2_buf_2 fanout25 (.A(_0291_),
    .X(net25));
 sg13g2_buf_2 fanout26 (.A(_0230_),
    .X(net26));
 sg13g2_buf_2 fanout27 (.A(_0951_),
    .X(net27));
 sg13g2_buf_2 fanout28 (.A(_0786_),
    .X(net28));
 sg13g2_buf_2 fanout29 (.A(_0785_),
    .X(net29));
 sg13g2_buf_2 fanout30 (.A(_0685_),
    .X(net30));
 sg13g2_buf_2 fanout31 (.A(_0683_),
    .X(net31));
 sg13g2_buf_2 fanout32 (.A(_0673_),
    .X(net32));
 sg13g2_buf_2 fanout33 (.A(_0671_),
    .X(net33));
 sg13g2_buf_2 fanout34 (.A(_0669_),
    .X(net34));
 sg13g2_buf_2 fanout35 (.A(_0626_),
    .X(net35));
 sg13g2_buf_2 fanout36 (.A(_0000_),
    .X(net36));
 sg13g2_buf_2 fanout37 (.A(_0924_),
    .X(net37));
 sg13g2_buf_2 fanout38 (.A(_0920_),
    .X(net38));
 sg13g2_buf_2 fanout39 (.A(_0782_),
    .X(net39));
 sg13g2_buf_2 fanout40 (.A(_0720_),
    .X(net40));
 sg13g2_buf_2 fanout41 (.A(_0697_),
    .X(net41));
 sg13g2_buf_2 fanout42 (.A(_0680_),
    .X(net42));
 sg13g2_buf_2 fanout43 (.A(_0676_),
    .X(net43));
 sg13g2_buf_2 fanout44 (.A(_0675_),
    .X(net44));
 sg13g2_buf_2 fanout45 (.A(_0672_),
    .X(net45));
 sg13g2_buf_2 fanout46 (.A(_0670_),
    .X(net46));
 sg13g2_buf_2 fanout47 (.A(_0666_),
    .X(net47));
 sg13g2_buf_2 fanout48 (.A(_0652_),
    .X(net48));
 sg13g2_buf_2 fanout49 (.A(_0647_),
    .X(net49));
 sg13g2_buf_2 fanout50 (.A(_0625_),
    .X(net50));
 sg13g2_buf_2 fanout51 (.A(_0621_),
    .X(net51));
 sg13g2_buf_2 fanout52 (.A(_0559_),
    .X(net52));
 sg13g2_buf_2 fanout53 (.A(_0533_),
    .X(net53));
 sg13g2_buf_2 fanout54 (.A(_0530_),
    .X(net54));
 sg13g2_buf_2 fanout55 (.A(_0527_),
    .X(net55));
 sg13g2_buf_4 fanout56 (.X(net56),
    .A(net60));
 sg13g2_buf_4 fanout57 (.X(net57),
    .A(net59));
 sg13g2_buf_2 fanout58 (.A(net59),
    .X(net58));
 sg13g2_buf_2 fanout59 (.A(net60),
    .X(net59));
 sg13g2_buf_2 fanout60 (.A(net1),
    .X(net60));
 sg13g2_buf_4 fanout61 (.X(net61),
    .A(net63));
 sg13g2_buf_4 fanout62 (.X(net62),
    .A(net64));
 sg13g2_buf_2 fanout63 (.A(net64),
    .X(net63));
 sg13g2_buf_2 fanout64 (.A(net1),
    .X(net64));
 sg13g2_tielo _2135__65 (.L_LO(net65));
 sg13g2_tielo _2136__66 (.L_LO(net66));
 sg13g2_tielo _2137__67 (.L_LO(net67));
 sg13g2_tielo _2138__68 (.L_LO(net68));
 sg13g2_tielo _2139__69 (.L_LO(net69));
 sg13g2_tielo _2140__70 (.L_LO(net70));
 sg13g2_tielo _2143__71 (.L_LO(net71));
 sg13g2_tielo _2144__72 (.L_LO(net72));
 sg13g2_tielo _2145__73 (.L_LO(net73));
 sg13g2_tielo _2146__74 (.L_LO(net74));
 sg13g2_tielo _2147__75 (.L_LO(net75));
 sg13g2_tielo _2148__76 (.L_LO(net76));
 sg13g2_tielo _2152__77 (.L_LO(net77));
 sg13g2_tielo _2154__78 (.L_LO(net78));
 sg13g2_tielo _2155__79 (.L_LO(net79));
 sg13g2_tielo _2156__80 (.L_LO(net80));
 sg13g2_tiehi \autosel.addr_counter[1]$_SDFFE_PN0P__82  (.L_HI(net82));
 sg13g2_tiehi \autosel.addr_counter[2]$_SDFFE_PN0P__83  (.L_HI(net83));
 sg13g2_tiehi \autosel.addr_counter[3]$_SDFFE_PN0P__84  (.L_HI(net84));
 sg13g2_tiehi \autosel.addr_counter[4]$_SDFFE_PN0P__85  (.L_HI(net85));
 sg13g2_tiehi \autosel.addr_counter[5]$_SDFFE_PN0P__86  (.L_HI(net86));
 sg13g2_tiehi \autosel.addr_counter[6]$_SDFFE_PN0P__87  (.L_HI(net87));
 sg13g2_tiehi \autosel.addr_counter[7]$_SDFFE_PN0P__88  (.L_HI(net88));
 sg13g2_tiehi \autosel.addr_counter[8]$_SDFFE_PN0P__89  (.L_HI(net89));
 sg13g2_tiehi \autosel.addr_counter[9]$_SDFFE_PN0P__90  (.L_HI(net90));
 sg13g2_tiehi \autosel.ctrl_ena$_SDFFE_PN0P__91  (.L_HI(net91));
 sg13g2_tiehi \autosel.ctrl_sel_inc$_SDFFE_PN0P__92  (.L_HI(net92));
 sg13g2_tiehi \autosel.ctrl_sel_rst_n$_SDFFE_PN0P__93  (.L_HI(net93));
 sg13g2_tiehi \autosel.i2c.data_out_hi[0]$_DFFE_PP__94  (.L_HI(net94));
 sg13g2_tiehi \autosel.i2c.data_out_hi[1]$_DFFE_PP__95  (.L_HI(net95));
 sg13g2_tiehi \autosel.i2c.data_out_hi[2]$_DFFE_PP__96  (.L_HI(net96));
 sg13g2_tiehi \autosel.i2c.data_out_hi[3]$_DFFE_PP__97  (.L_HI(net97));
 sg13g2_tiehi \autosel.i2c.data_out_hi[4]$_DFFE_PP__98  (.L_HI(net98));
 sg13g2_tiehi \autosel.i2c.data_out_hi[5]$_DFFE_PP__99  (.L_HI(net99));
 sg13g2_tiehi \autosel.i2c.data_out_hi[6]$_DFFE_PP__100  (.L_HI(net100));
 sg13g2_tiehi \autosel.i2c.data_out_hi[7]$_DFFE_PP__101  (.L_HI(net101));
 sg13g2_tiehi \autosel.i2c.i2c.addr_reg[4]$_DFFE_PP__102  (.L_HI(net102));
 sg13g2_tiehi \autosel.i2c.i2c.bit_count_reg[0]$_SDFFCE_PN0P__103  (.L_HI(net103));
 sg13g2_tiehi \autosel.i2c.i2c.bit_count_reg[1]$_SDFFCE_PN0P__104  (.L_HI(net104));
 sg13g2_tiehi \autosel.i2c.i2c.bit_count_reg[2]$_SDFFCE_PN0P__105  (.L_HI(net105));
 sg13g2_tiehi \autosel.i2c.i2c.bit_count_reg[3]$_SDFFCE_PN1P__106  (.L_HI(net106));
 sg13g2_tiehi \autosel.i2c.i2c.bus_active_reg$_SDFFE_PN0P__107  (.L_HI(net107));
 sg13g2_tiehi \autosel.i2c.i2c.busy_reg$_SDFF_PN0__108  (.L_HI(net108));
 sg13g2_tiehi \autosel.i2c.i2c.data_reg[0]$_SDFFCE_PN0P__109  (.L_HI(net109));
 sg13g2_tiehi \autosel.i2c.i2c.data_reg[1]$_SDFFCE_PN0P__110  (.L_HI(net110));
 sg13g2_tiehi \autosel.i2c.i2c.data_reg[2]$_SDFFCE_PN0P__111  (.L_HI(net111));
 sg13g2_tiehi \autosel.i2c.i2c.data_reg[3]$_SDFFCE_PN0P__112  (.L_HI(net112));
 sg13g2_tiehi \autosel.i2c.i2c.data_reg[4]$_SDFFCE_PN0P__113  (.L_HI(net113));
 sg13g2_tiehi \autosel.i2c.i2c.data_reg[5]$_SDFFCE_PN0P__114  (.L_HI(net114));
 sg13g2_tiehi \autosel.i2c.i2c.data_reg[6]$_SDFFCE_PN0P__115  (.L_HI(net115));
 sg13g2_tiehi \autosel.i2c.i2c.data_reg[7]$_SDFFCE_PN0P__116  (.L_HI(net116));
 sg13g2_tiehi \autosel.i2c.i2c.delay_reg[0]$_SDFFE_PN0P__117  (.L_HI(net117));
 sg13g2_tiehi \autosel.i2c.i2c.delay_reg[10]$_SDFFE_PN0P__118  (.L_HI(net118));
 sg13g2_tiehi \autosel.i2c.i2c.delay_reg[11]$_SDFFE_PN0P__119  (.L_HI(net119));
 sg13g2_tiehi \autosel.i2c.i2c.delay_reg[12]$_SDFFE_PN0P__120  (.L_HI(net120));
 sg13g2_tiehi \autosel.i2c.i2c.delay_reg[13]$_SDFFE_PN0P__121  (.L_HI(net121));
 sg13g2_tiehi \autosel.i2c.i2c.delay_reg[14]$_SDFFE_PN0P__122  (.L_HI(net122));
 sg13g2_tiehi \autosel.i2c.i2c.delay_reg[15]$_SDFFE_PN0P__123  (.L_HI(net123));
 sg13g2_tiehi \autosel.i2c.i2c.delay_reg[1]$_SDFFE_PN0P__124  (.L_HI(net124));
 sg13g2_tiehi \autosel.i2c.i2c.delay_reg[2]$_SDFFE_PN0P__125  (.L_HI(net125));
 sg13g2_tiehi \autosel.i2c.i2c.delay_reg[3]$_SDFFE_PN0P__126  (.L_HI(net126));
 sg13g2_tiehi \autosel.i2c.i2c.delay_reg[4]$_SDFFE_PN0P__127  (.L_HI(net127));
 sg13g2_tiehi \autosel.i2c.i2c.delay_reg[5]$_SDFFE_PN0P__128  (.L_HI(net128));
 sg13g2_tiehi \autosel.i2c.i2c.delay_reg[6]$_SDFFE_PN0P__129  (.L_HI(net129));
 sg13g2_tiehi \autosel.i2c.i2c.delay_reg[7]$_SDFFE_PN0P__130  (.L_HI(net130));
 sg13g2_tiehi \autosel.i2c.i2c.delay_reg[8]$_SDFFE_PN0P__131  (.L_HI(net131));
 sg13g2_tiehi \autosel.i2c.i2c.delay_reg[9]$_SDFFE_PN0P__132  (.L_HI(net132));
 sg13g2_tiehi \autosel.i2c.i2c.delay_scl_reg$_SDFF_PN0__133  (.L_HI(net133));
 sg13g2_tiehi \autosel.i2c.i2c.delay_sda_reg$_SDFFE_PN0N__134  (.L_HI(net134));
 sg13g2_tiehi \autosel.i2c.i2c.last_sda_i_reg$_DFF_P__135  (.L_HI(net135));
 sg13g2_tiehi \autosel.i2c.i2c.m_axis_data_tdata_reg[0]$_DFFE_PP__136  (.L_HI(net136));
 sg13g2_tiehi \autosel.i2c.i2c.m_axis_data_tdata_reg[1]$_DFFE_PP__137  (.L_HI(net137));
 sg13g2_tiehi \autosel.i2c.i2c.m_axis_data_tdata_reg[2]$_DFFE_PP__138  (.L_HI(net138));
 sg13g2_tiehi \autosel.i2c.i2c.m_axis_data_tdata_reg[3]$_DFFE_PP__139  (.L_HI(net139));
 sg13g2_tiehi \autosel.i2c.i2c.m_axis_data_tdata_reg[4]$_DFFE_PP__140  (.L_HI(net140));
 sg13g2_tiehi \autosel.i2c.i2c.m_axis_data_tdata_reg[5]$_DFFE_PP__141  (.L_HI(net141));
 sg13g2_tiehi \autosel.i2c.i2c.m_axis_data_tdata_reg[6]$_DFFE_PP__142  (.L_HI(net142));
 sg13g2_tiehi \autosel.i2c.i2c.m_axis_data_tdata_reg[7]$_DFFE_PP__143  (.L_HI(net143));
 sg13g2_tiehi \autosel.i2c.i2c.m_axis_data_tvalid_reg$_SDFF_PN0__144  (.L_HI(net144));
 sg13g2_tiehi \autosel.i2c.i2c.missed_ack_reg$_SDFF_PP0__145  (.L_HI(net145));
 sg13g2_tiehi \autosel.i2c.i2c.mode_read_reg$_DFFE_PP__146  (.L_HI(net146));
 sg13g2_tiehi \autosel.i2c.i2c.mode_stop_reg$_DFFE_PP__147  (.L_HI(net147));
 sg13g2_tiehi \autosel.i2c.i2c.phy_rx_data_reg$_DFFE_PP__148  (.L_HI(net148));
 sg13g2_tiehi \autosel.i2c.i2c.phy_state_reg[0]$_SDFFE_PN0P__149  (.L_HI(net149));
 sg13g2_tiehi \autosel.i2c.i2c.phy_state_reg[1]$_SDFFE_PN0P__150  (.L_HI(net150));
 sg13g2_tiehi \autosel.i2c.i2c.phy_state_reg[2]$_SDFFE_PN0P__151  (.L_HI(net151));
 sg13g2_tiehi \autosel.i2c.i2c.phy_state_reg[3]$_SDFFE_PN0P__152  (.L_HI(net152));
 sg13g2_tiehi \autosel.i2c.i2c.s_axis_cmd_ready_reg$_SDFF_PP0__153  (.L_HI(net153));
 sg13g2_tiehi \autosel.i2c.i2c.s_axis_data_tready_reg$_SDFF_PP0__154  (.L_HI(net154));
 sg13g2_tiehi \autosel.i2c.i2c.scl_i_reg$_DFF_P__155  (.L_HI(net155));
 sg13g2_tiehi \autosel.i2c.i2c.scl_o_reg$_SDFFE_PN1P__156  (.L_HI(net156));
 sg13g2_tiehi \autosel.i2c.i2c.sda_i_reg$_DFF_P__157  (.L_HI(net157));
 sg13g2_tiehi \autosel.i2c.i2c.sda_o_reg$_SDFFE_PN1P__158  (.L_HI(net158));
 sg13g2_tiehi \autosel.i2c.i2c.state_reg[0]$_SDFFE_PN0N__159  (.L_HI(net159));
 sg13g2_tiehi \autosel.i2c.i2c.state_reg[1]$_SDFFE_PN0N__160  (.L_HI(net160));
 sg13g2_tiehi \autosel.i2c.i2c.state_reg[2]$_SDFFE_PN0N__161  (.L_HI(net161));
 sg13g2_tiehi \autosel.i2c.i2c.state_reg[3]$_SDFFE_PN0N__162  (.L_HI(net162));
 sg13g2_tiehi \autosel.state[0]$_DFF_P__163  (.L_HI(net163));
 sg13g2_tiehi \autosel.state[1]$_DFF_P__164  (.L_HI(net164));
 sg13g2_tiehi \autosel.state[2]$_DFF_P__165  (.L_HI(net165));
 sg13g2_tiehi \debug_out.counter[0]$_SDFF_PP0__166  (.L_HI(net166));
 sg13g2_tiehi \debug_out.counter[10]$_SDFF_PP0__167  (.L_HI(net167));
 sg13g2_tiehi \debug_out.counter[11]$_SDFF_PP0__168  (.L_HI(net168));
 sg13g2_tiehi \debug_out.counter[12]$_SDFF_PP0__169  (.L_HI(net169));
 sg13g2_tiehi \debug_out.counter[13]$_SDFF_PP0__170  (.L_HI(net170));
 sg13g2_tiehi \debug_out.counter[14]$_SDFF_PP0__171  (.L_HI(net171));
 sg13g2_tiehi \debug_out.counter[15]$_SDFF_PP0__172  (.L_HI(net172));
 sg13g2_tiehi \debug_out.counter[16]$_SDFF_PP0__173  (.L_HI(net173));
 sg13g2_tiehi \debug_out.counter[17]$_SDFF_PP0__174  (.L_HI(net174));
 sg13g2_tiehi \debug_out.counter[18]$_SDFF_PP0__175  (.L_HI(net175));
 sg13g2_tiehi \debug_out.counter[19]$_SDFF_PP0__176  (.L_HI(net176));
 sg13g2_tiehi \debug_out.counter[1]$_SDFF_PP0__177  (.L_HI(net177));
 sg13g2_tiehi \debug_out.counter[20]$_SDFF_PP0__178  (.L_HI(net178));
 sg13g2_tiehi \debug_out.counter[21]$_SDFF_PP0__179  (.L_HI(net179));
 sg13g2_tiehi \debug_out.counter[22]$_SDFF_PP0__180  (.L_HI(net180));
 sg13g2_tiehi \debug_out.counter[23]$_SDFF_PP0__181  (.L_HI(net181));
 sg13g2_tiehi \debug_out.counter[24]$_SDFF_PP0__182  (.L_HI(net182));
 sg13g2_tiehi \debug_out.counter[25]$_SDFF_PP0__183  (.L_HI(net183));
 sg13g2_tiehi \debug_out.counter[26]$_SDFF_PP0__184  (.L_HI(net184));
 sg13g2_tiehi \debug_out.counter[27]$_SDFF_PP0__185  (.L_HI(net185));
 sg13g2_tiehi \debug_out.counter[28]$_SDFF_PP0__186  (.L_HI(net186));
 sg13g2_tiehi \debug_out.counter[29]$_SDFF_PP0__187  (.L_HI(net187));
 sg13g2_tiehi \debug_out.counter[2]$_SDFF_PP0__188  (.L_HI(net188));
 sg13g2_tiehi \debug_out.counter[30]$_SDFF_PP0__189  (.L_HI(net189));
 sg13g2_tiehi \debug_out.counter[31]$_SDFF_PP0__190  (.L_HI(net190));
 sg13g2_tiehi \debug_out.counter[3]$_SDFF_PP0__191  (.L_HI(net191));
 sg13g2_tiehi \debug_out.counter[4]$_SDFF_PP0__192  (.L_HI(net192));
 sg13g2_tiehi \debug_out.counter[5]$_SDFF_PP0__193  (.L_HI(net193));
 sg13g2_tiehi \debug_out.counter[6]$_SDFF_PP0__194  (.L_HI(net194));
 sg13g2_tiehi \debug_out.counter[7]$_SDFF_PP0__195  (.L_HI(net195));
 sg13g2_tiehi \debug_out.counter[8]$_SDFF_PP0__196  (.L_HI(net196));
 sg13g2_tiehi \debug_out.counter[9]$_SDFF_PP0__197  (.L_HI(net197));
 sg13g2_tiehi \debug_out.send_index[0]$_SDFFE_PP0P__198  (.L_HI(net198));
 sg13g2_tiehi \debug_out.send_index[1]$_SDFFE_PP0P__199  (.L_HI(net199));
 sg13g2_tiehi \debug_out.send_index[2]$_SDFFE_PP0P__200  (.L_HI(net200));
 sg13g2_tiehi \debug_out.tx_byte[0]$_SDFFE_PN0P__201  (.L_HI(net201));
 sg13g2_tiehi \debug_out.tx_byte[1]$_SDFFE_PN0P__202  (.L_HI(net202));
 sg13g2_tiehi \debug_out.tx_byte[2]$_SDFFE_PN0P__203  (.L_HI(net203));
 sg13g2_tiehi \debug_out.tx_byte[3]$_SDFFE_PN0P__204  (.L_HI(net204));
 sg13g2_tiehi \debug_out.tx_byte[5]$_SDFFE_PN0P__205  (.L_HI(net205));
 sg13g2_tiehi \debug_out.tx_byte[6]$_SDFFE_PN0P__206  (.L_HI(net206));
 sg13g2_tiehi \debug_out.tx_valid$_SDFFE_PN0P__207  (.L_HI(net207));
 sg13g2_buf_2 clkbuf_4_0_0_clk (.A(clknet_0_clk),
    .X(clknet_4_0_0_clk));
 sg13g2_buf_2 clkbuf_4_1_0_clk (.A(clknet_0_clk),
    .X(clknet_4_1_0_clk));
 sg13g2_buf_2 clkbuf_4_2_0_clk (.A(clknet_0_clk),
    .X(clknet_4_2_0_clk));
 sg13g2_buf_2 clkbuf_4_3_0_clk (.A(clknet_0_clk),
    .X(clknet_4_3_0_clk));
 sg13g2_buf_2 clkbuf_4_4_0_clk (.A(clknet_0_clk),
    .X(clknet_4_4_0_clk));
 sg13g2_buf_2 clkbuf_4_5_0_clk (.A(clknet_0_clk),
    .X(clknet_4_5_0_clk));
 sg13g2_buf_2 clkbuf_4_6_0_clk (.A(clknet_0_clk),
    .X(clknet_4_6_0_clk));
 sg13g2_buf_2 clkbuf_4_7_0_clk (.A(clknet_0_clk),
    .X(clknet_4_7_0_clk));
 sg13g2_buf_2 clkbuf_4_8_0_clk (.A(clknet_0_clk),
    .X(clknet_4_8_0_clk));
 sg13g2_buf_2 clkbuf_4_9_0_clk (.A(clknet_0_clk),
    .X(clknet_4_9_0_clk));
 sg13g2_buf_2 clkbuf_4_10_0_clk (.A(clknet_0_clk),
    .X(clknet_4_10_0_clk));
 sg13g2_buf_2 clkbuf_4_11_0_clk (.A(clknet_0_clk),
    .X(clknet_4_11_0_clk));
 sg13g2_buf_2 clkbuf_4_12_0_clk (.A(clknet_0_clk),
    .X(clknet_4_12_0_clk));
 sg13g2_buf_2 clkbuf_4_13_0_clk (.A(clknet_0_clk),
    .X(clknet_4_13_0_clk));
 sg13g2_buf_2 clkbuf_4_14_0_clk (.A(clknet_0_clk),
    .X(clknet_4_14_0_clk));
 sg13g2_buf_2 clkbuf_4_15_0_clk (.A(clknet_0_clk),
    .X(clknet_4_15_0_clk));
 sg13g2_buf_1 clkbuf_5_0__f_clk (.A(clknet_4_0_0_clk),
    .X(clknet_5_0__leaf_clk));
 sg13g2_buf_1 clkbuf_5_1__f_clk (.A(clknet_4_0_0_clk),
    .X(clknet_5_1__leaf_clk));
 sg13g2_buf_1 clkbuf_5_2__f_clk (.A(clknet_4_1_0_clk),
    .X(clknet_5_2__leaf_clk));
 sg13g2_buf_1 clkbuf_5_3__f_clk (.A(clknet_4_1_0_clk),
    .X(clknet_5_3__leaf_clk));
 sg13g2_buf_1 clkbuf_5_4__f_clk (.A(clknet_4_2_0_clk),
    .X(clknet_5_4__leaf_clk));
 sg13g2_buf_1 clkbuf_5_5__f_clk (.A(clknet_4_2_0_clk),
    .X(clknet_5_5__leaf_clk));
 sg13g2_buf_1 clkbuf_5_6__f_clk (.A(clknet_4_3_0_clk),
    .X(clknet_5_6__leaf_clk));
 sg13g2_buf_1 clkbuf_5_7__f_clk (.A(clknet_4_3_0_clk),
    .X(clknet_5_7__leaf_clk));
 sg13g2_buf_1 clkbuf_5_8__f_clk (.A(clknet_4_4_0_clk),
    .X(clknet_5_8__leaf_clk));
 sg13g2_buf_1 clkbuf_5_9__f_clk (.A(clknet_4_4_0_clk),
    .X(clknet_5_9__leaf_clk));
 sg13g2_buf_1 clkbuf_5_10__f_clk (.A(clknet_4_5_0_clk),
    .X(clknet_5_10__leaf_clk));
 sg13g2_buf_1 clkbuf_5_11__f_clk (.A(clknet_4_5_0_clk),
    .X(clknet_5_11__leaf_clk));
 sg13g2_buf_1 clkbuf_5_12__f_clk (.A(clknet_4_6_0_clk),
    .X(clknet_5_12__leaf_clk));
 sg13g2_buf_1 clkbuf_5_13__f_clk (.A(clknet_4_6_0_clk),
    .X(clknet_5_13__leaf_clk));
 sg13g2_buf_1 clkbuf_5_14__f_clk (.A(clknet_4_7_0_clk),
    .X(clknet_5_14__leaf_clk));
 sg13g2_buf_1 clkbuf_5_15__f_clk (.A(clknet_4_7_0_clk),
    .X(clknet_5_15__leaf_clk));
 sg13g2_buf_1 clkbuf_5_16__f_clk (.A(clknet_4_8_0_clk),
    .X(clknet_5_16__leaf_clk));
 sg13g2_buf_1 clkbuf_5_17__f_clk (.A(clknet_4_8_0_clk),
    .X(clknet_5_17__leaf_clk));
 sg13g2_buf_1 clkbuf_5_18__f_clk (.A(clknet_4_9_0_clk),
    .X(clknet_5_18__leaf_clk));
 sg13g2_buf_1 clkbuf_5_19__f_clk (.A(clknet_4_9_0_clk),
    .X(clknet_5_19__leaf_clk));
 sg13g2_buf_1 clkbuf_5_20__f_clk (.A(clknet_4_10_0_clk),
    .X(clknet_5_20__leaf_clk));
 sg13g2_buf_1 clkbuf_5_21__f_clk (.A(clknet_4_10_0_clk),
    .X(clknet_5_21__leaf_clk));
 sg13g2_buf_1 clkbuf_5_22__f_clk (.A(clknet_4_11_0_clk),
    .X(clknet_5_22__leaf_clk));
 sg13g2_buf_1 clkbuf_5_23__f_clk (.A(clknet_4_11_0_clk),
    .X(clknet_5_23__leaf_clk));
 sg13g2_buf_1 clkbuf_5_24__f_clk (.A(clknet_4_12_0_clk),
    .X(clknet_5_24__leaf_clk));
 sg13g2_buf_1 clkbuf_5_25__f_clk (.A(clknet_4_12_0_clk),
    .X(clknet_5_25__leaf_clk));
 sg13g2_buf_1 clkbuf_5_26__f_clk (.A(clknet_4_13_0_clk),
    .X(clknet_5_26__leaf_clk));
 sg13g2_buf_1 clkbuf_5_27__f_clk (.A(clknet_4_13_0_clk),
    .X(clknet_5_27__leaf_clk));
 sg13g2_buf_1 clkbuf_5_28__f_clk (.A(clknet_4_14_0_clk),
    .X(clknet_5_28__leaf_clk));
 sg13g2_buf_1 clkbuf_5_29__f_clk (.A(clknet_4_14_0_clk),
    .X(clknet_5_29__leaf_clk));
 sg13g2_buf_1 clkbuf_5_30__f_clk (.A(clknet_4_15_0_clk),
    .X(clknet_5_30__leaf_clk));
 sg13g2_buf_1 clkbuf_5_31__f_clk (.A(clknet_4_15_0_clk),
    .X(clknet_5_31__leaf_clk));
 sg13g2_inv_1 clkload0 (.A(clknet_5_3__leaf_clk));
 sg13g2_inv_1 clkload1 (.A(clknet_5_5__leaf_clk));
 sg13g2_inv_1 clkload2 (.A(clknet_5_7__leaf_clk));
 sg13g2_inv_1 clkload3 (.A(clknet_5_9__leaf_clk));
 sg13g2_inv_1 clkload4 (.A(clknet_5_11__leaf_clk));
 sg13g2_inv_1 clkload5 (.A(clknet_5_13__leaf_clk));
 sg13g2_inv_1 clkload6 (.A(clknet_5_15__leaf_clk));
 sg13g2_inv_1 clkload7 (.A(clknet_5_17__leaf_clk));
 sg13g2_inv_1 clkload8 (.A(clknet_5_19__leaf_clk));
 sg13g2_inv_1 clkload9 (.A(clknet_5_21__leaf_clk));
 sg13g2_inv_1 clkload10 (.A(clknet_5_23__leaf_clk));
 sg13g2_inv_1 clkload11 (.A(clknet_5_25__leaf_clk));
 sg13g2_inv_1 clkload12 (.A(clknet_5_27__leaf_clk));
 sg13g2_inv_1 clkload13 (.A(clknet_5_29__leaf_clk));
 sg13g2_inv_1 clkload14 (.A(clknet_5_31__leaf_clk));
 sg13g2_decap_8 FILLER_0_0 ();
 sg13g2_decap_8 FILLER_0_7 ();
 sg13g2_decap_8 FILLER_0_14 ();
 sg13g2_decap_8 FILLER_0_21 ();
 sg13g2_decap_4 FILLER_0_28 ();
 sg13g2_fill_1 FILLER_0_32 ();
 sg13g2_decap_8 FILLER_0_37 ();
 sg13g2_decap_4 FILLER_0_44 ();
 sg13g2_fill_1 FILLER_0_48 ();
 sg13g2_decap_8 FILLER_0_65 ();
 sg13g2_decap_8 FILLER_0_72 ();
 sg13g2_decap_4 FILLER_0_79 ();
 sg13g2_fill_2 FILLER_0_83 ();
 sg13g2_decap_8 FILLER_0_89 ();
 sg13g2_decap_4 FILLER_0_96 ();
 sg13g2_fill_1 FILLER_0_100 ();
 sg13g2_fill_2 FILLER_0_109 ();
 sg13g2_decap_4 FILLER_0_119 ();
 sg13g2_fill_2 FILLER_0_142 ();
 sg13g2_fill_1 FILLER_0_144 ();
 sg13g2_decap_8 FILLER_0_171 ();
 sg13g2_fill_1 FILLER_0_178 ();
 sg13g2_fill_2 FILLER_0_205 ();
 sg13g2_fill_1 FILLER_0_211 ();
 sg13g2_fill_2 FILLER_0_216 ();
 sg13g2_fill_2 FILLER_0_249 ();
 sg13g2_fill_1 FILLER_0_251 ();
 sg13g2_decap_8 FILLER_0_278 ();
 sg13g2_fill_1 FILLER_0_285 ();
 sg13g2_fill_2 FILLER_0_316 ();
 sg13g2_decap_8 FILLER_0_344 ();
 sg13g2_decap_4 FILLER_0_351 ();
 sg13g2_decap_4 FILLER_0_381 ();
 sg13g2_decap_8 FILLER_0_411 ();
 sg13g2_decap_8 FILLER_0_418 ();
 sg13g2_decap_4 FILLER_0_425 ();
 sg13g2_fill_1 FILLER_0_429 ();
 sg13g2_decap_8 FILLER_1_0 ();
 sg13g2_decap_8 FILLER_1_7 ();
 sg13g2_decap_8 FILLER_1_14 ();
 sg13g2_decap_4 FILLER_1_21 ();
 sg13g2_fill_1 FILLER_1_25 ();
 sg13g2_fill_1 FILLER_1_134 ();
 sg13g2_fill_2 FILLER_1_151 ();
 sg13g2_fill_1 FILLER_1_153 ();
 sg13g2_decap_8 FILLER_1_158 ();
 sg13g2_decap_8 FILLER_1_165 ();
 sg13g2_decap_8 FILLER_1_176 ();
 sg13g2_decap_8 FILLER_1_183 ();
 sg13g2_decap_8 FILLER_1_190 ();
 sg13g2_decap_4 FILLER_1_197 ();
 sg13g2_fill_2 FILLER_1_201 ();
 sg13g2_decap_8 FILLER_1_223 ();
 sg13g2_decap_8 FILLER_1_230 ();
 sg13g2_fill_2 FILLER_1_237 ();
 sg13g2_fill_1 FILLER_1_239 ();
 sg13g2_decap_8 FILLER_1_265 ();
 sg13g2_fill_1 FILLER_1_272 ();
 sg13g2_fill_2 FILLER_1_282 ();
 sg13g2_fill_1 FILLER_1_284 ();
 sg13g2_decap_8 FILLER_1_293 ();
 sg13g2_decap_8 FILLER_1_305 ();
 sg13g2_decap_8 FILLER_1_312 ();
 sg13g2_decap_8 FILLER_1_319 ();
 sg13g2_fill_1 FILLER_1_326 ();
 sg13g2_decap_4 FILLER_1_331 ();
 sg13g2_decap_8 FILLER_1_343 ();
 sg13g2_fill_1 FILLER_1_350 ();
 sg13g2_decap_8 FILLER_1_363 ();
 sg13g2_decap_8 FILLER_1_370 ();
 sg13g2_decap_4 FILLER_1_377 ();
 sg13g2_fill_2 FILLER_1_397 ();
 sg13g2_fill_1 FILLER_1_403 ();
 sg13g2_decap_8 FILLER_2_0 ();
 sg13g2_decap_4 FILLER_2_7 ();
 sg13g2_fill_2 FILLER_2_11 ();
 sg13g2_decap_8 FILLER_2_17 ();
 sg13g2_decap_8 FILLER_2_24 ();
 sg13g2_decap_8 FILLER_2_31 ();
 sg13g2_fill_1 FILLER_2_38 ();
 sg13g2_decap_4 FILLER_2_43 ();
 sg13g2_fill_2 FILLER_2_59 ();
 sg13g2_fill_1 FILLER_2_66 ();
 sg13g2_decap_8 FILLER_2_75 ();
 sg13g2_decap_8 FILLER_2_82 ();
 sg13g2_decap_8 FILLER_2_89 ();
 sg13g2_decap_8 FILLER_2_96 ();
 sg13g2_fill_1 FILLER_2_103 ();
 sg13g2_decap_8 FILLER_2_110 ();
 sg13g2_fill_1 FILLER_2_117 ();
 sg13g2_decap_8 FILLER_2_122 ();
 sg13g2_fill_1 FILLER_2_129 ();
 sg13g2_fill_2 FILLER_2_144 ();
 sg13g2_fill_2 FILLER_2_162 ();
 sg13g2_fill_1 FILLER_2_164 ();
 sg13g2_decap_8 FILLER_2_199 ();
 sg13g2_decap_8 FILLER_2_206 ();
 sg13g2_decap_8 FILLER_2_213 ();
 sg13g2_decap_8 FILLER_2_220 ();
 sg13g2_decap_4 FILLER_2_227 ();
 sg13g2_fill_1 FILLER_2_231 ();
 sg13g2_fill_1 FILLER_2_258 ();
 sg13g2_decap_8 FILLER_2_264 ();
 sg13g2_fill_1 FILLER_2_283 ();
 sg13g2_decap_4 FILLER_2_310 ();
 sg13g2_fill_2 FILLER_2_323 ();
 sg13g2_fill_1 FILLER_2_325 ();
 sg13g2_fill_1 FILLER_2_334 ();
 sg13g2_fill_2 FILLER_2_367 ();
 sg13g2_fill_1 FILLER_2_369 ();
 sg13g2_decap_4 FILLER_2_376 ();
 sg13g2_fill_2 FILLER_2_380 ();
 sg13g2_decap_8 FILLER_2_401 ();
 sg13g2_decap_8 FILLER_2_408 ();
 sg13g2_decap_8 FILLER_2_415 ();
 sg13g2_decap_8 FILLER_2_422 ();
 sg13g2_fill_1 FILLER_2_429 ();
 sg13g2_fill_2 FILLER_3_0 ();
 sg13g2_decap_8 FILLER_3_44 ();
 sg13g2_fill_2 FILLER_3_51 ();
 sg13g2_fill_1 FILLER_3_53 ();
 sg13g2_fill_2 FILLER_3_62 ();
 sg13g2_decap_4 FILLER_3_70 ();
 sg13g2_fill_2 FILLER_3_141 ();
 sg13g2_fill_1 FILLER_3_143 ();
 sg13g2_fill_2 FILLER_3_153 ();
 sg13g2_decap_8 FILLER_3_219 ();
 sg13g2_decap_8 FILLER_3_226 ();
 sg13g2_fill_2 FILLER_3_233 ();
 sg13g2_fill_2 FILLER_3_239 ();
 sg13g2_fill_1 FILLER_3_241 ();
 sg13g2_fill_1 FILLER_3_246 ();
 sg13g2_fill_1 FILLER_3_268 ();
 sg13g2_fill_2 FILLER_3_279 ();
 sg13g2_decap_8 FILLER_3_323 ();
 sg13g2_decap_8 FILLER_3_330 ();
 sg13g2_fill_2 FILLER_3_342 ();
 sg13g2_fill_1 FILLER_3_344 ();
 sg13g2_fill_1 FILLER_3_351 ();
 sg13g2_decap_4 FILLER_3_386 ();
 sg13g2_fill_1 FILLER_3_390 ();
 sg13g2_decap_8 FILLER_3_399 ();
 sg13g2_decap_8 FILLER_3_406 ();
 sg13g2_decap_8 FILLER_3_413 ();
 sg13g2_decap_8 FILLER_3_420 ();
 sg13g2_fill_2 FILLER_3_427 ();
 sg13g2_fill_1 FILLER_3_429 ();
 sg13g2_fill_2 FILLER_4_0 ();
 sg13g2_fill_2 FILLER_4_32 ();
 sg13g2_decap_4 FILLER_4_46 ();
 sg13g2_fill_2 FILLER_4_50 ();
 sg13g2_decap_4 FILLER_4_75 ();
 sg13g2_fill_1 FILLER_4_79 ();
 sg13g2_fill_1 FILLER_4_84 ();
 sg13g2_decap_8 FILLER_4_93 ();
 sg13g2_decap_8 FILLER_4_100 ();
 sg13g2_decap_8 FILLER_4_107 ();
 sg13g2_fill_2 FILLER_4_114 ();
 sg13g2_decap_8 FILLER_4_125 ();
 sg13g2_decap_8 FILLER_4_132 ();
 sg13g2_decap_8 FILLER_4_139 ();
 sg13g2_decap_8 FILLER_4_163 ();
 sg13g2_decap_8 FILLER_4_174 ();
 sg13g2_decap_8 FILLER_4_181 ();
 sg13g2_fill_2 FILLER_4_188 ();
 sg13g2_fill_1 FILLER_4_194 ();
 sg13g2_fill_2 FILLER_4_199 ();
 sg13g2_decap_8 FILLER_4_209 ();
 sg13g2_decap_8 FILLER_4_216 ();
 sg13g2_fill_2 FILLER_4_223 ();
 sg13g2_fill_1 FILLER_4_225 ();
 sg13g2_decap_4 FILLER_4_280 ();
 sg13g2_fill_2 FILLER_4_284 ();
 sg13g2_fill_2 FILLER_4_290 ();
 sg13g2_decap_8 FILLER_4_299 ();
 sg13g2_decap_8 FILLER_4_306 ();
 sg13g2_decap_8 FILLER_4_313 ();
 sg13g2_fill_2 FILLER_4_320 ();
 sg13g2_decap_8 FILLER_4_357 ();
 sg13g2_decap_8 FILLER_4_364 ();
 sg13g2_decap_8 FILLER_4_371 ();
 sg13g2_fill_2 FILLER_4_378 ();
 sg13g2_decap_8 FILLER_4_383 ();
 sg13g2_decap_4 FILLER_4_390 ();
 sg13g2_decap_4 FILLER_4_424 ();
 sg13g2_fill_2 FILLER_4_428 ();
 sg13g2_decap_8 FILLER_5_0 ();
 sg13g2_decap_4 FILLER_5_7 ();
 sg13g2_fill_2 FILLER_5_11 ();
 sg13g2_fill_1 FILLER_5_17 ();
 sg13g2_fill_2 FILLER_5_22 ();
 sg13g2_fill_2 FILLER_5_28 ();
 sg13g2_fill_2 FILLER_5_38 ();
 sg13g2_fill_1 FILLER_5_40 ();
 sg13g2_decap_4 FILLER_5_46 ();
 sg13g2_fill_1 FILLER_5_64 ();
 sg13g2_fill_1 FILLER_5_99 ();
 sg13g2_decap_4 FILLER_5_104 ();
 sg13g2_decap_8 FILLER_5_134 ();
 sg13g2_decap_4 FILLER_5_141 ();
 sg13g2_fill_2 FILLER_5_145 ();
 sg13g2_fill_2 FILLER_5_159 ();
 sg13g2_fill_1 FILLER_5_161 ();
 sg13g2_fill_2 FILLER_5_188 ();
 sg13g2_fill_1 FILLER_5_203 ();
 sg13g2_decap_8 FILLER_5_230 ();
 sg13g2_decap_8 FILLER_5_237 ();
 sg13g2_decap_8 FILLER_5_244 ();
 sg13g2_decap_4 FILLER_5_251 ();
 sg13g2_fill_1 FILLER_5_255 ();
 sg13g2_decap_8 FILLER_5_260 ();
 sg13g2_fill_1 FILLER_5_267 ();
 sg13g2_decap_8 FILLER_5_294 ();
 sg13g2_decap_8 FILLER_5_301 ();
 sg13g2_decap_8 FILLER_5_308 ();
 sg13g2_decap_8 FILLER_5_315 ();
 sg13g2_decap_8 FILLER_5_322 ();
 sg13g2_fill_2 FILLER_5_329 ();
 sg13g2_fill_2 FILLER_5_336 ();
 sg13g2_fill_2 FILLER_5_350 ();
 sg13g2_decap_4 FILLER_5_356 ();
 sg13g2_fill_2 FILLER_5_360 ();
 sg13g2_decap_8 FILLER_5_398 ();
 sg13g2_decap_8 FILLER_5_405 ();
 sg13g2_decap_8 FILLER_5_412 ();
 sg13g2_decap_8 FILLER_5_419 ();
 sg13g2_decap_4 FILLER_5_426 ();
 sg13g2_decap_4 FILLER_6_0 ();
 sg13g2_fill_2 FILLER_6_4 ();
 sg13g2_decap_4 FILLER_6_32 ();
 sg13g2_fill_2 FILLER_6_36 ();
 sg13g2_decap_8 FILLER_6_42 ();
 sg13g2_decap_8 FILLER_6_49 ();
 sg13g2_decap_4 FILLER_6_56 ();
 sg13g2_decap_8 FILLER_6_86 ();
 sg13g2_fill_2 FILLER_6_93 ();
 sg13g2_fill_1 FILLER_6_95 ();
 sg13g2_decap_8 FILLER_6_104 ();
 sg13g2_decap_8 FILLER_6_119 ();
 sg13g2_decap_8 FILLER_6_126 ();
 sg13g2_decap_8 FILLER_6_133 ();
 sg13g2_fill_2 FILLER_6_140 ();
 sg13g2_fill_1 FILLER_6_142 ();
 sg13g2_decap_4 FILLER_6_163 ();
 sg13g2_fill_1 FILLER_6_167 ();
 sg13g2_decap_8 FILLER_6_172 ();
 sg13g2_decap_8 FILLER_6_183 ();
 sg13g2_fill_1 FILLER_6_193 ();
 sg13g2_decap_4 FILLER_6_198 ();
 sg13g2_decap_4 FILLER_6_206 ();
 sg13g2_decap_8 FILLER_6_218 ();
 sg13g2_decap_8 FILLER_6_225 ();
 sg13g2_decap_4 FILLER_6_232 ();
 sg13g2_decap_8 FILLER_6_266 ();
 sg13g2_decap_8 FILLER_6_273 ();
 sg13g2_decap_8 FILLER_6_280 ();
 sg13g2_decap_8 FILLER_6_287 ();
 sg13g2_decap_8 FILLER_6_294 ();
 sg13g2_decap_8 FILLER_6_301 ();
 sg13g2_decap_8 FILLER_6_308 ();
 sg13g2_decap_8 FILLER_6_315 ();
 sg13g2_decap_8 FILLER_6_322 ();
 sg13g2_fill_1 FILLER_6_329 ();
 sg13g2_fill_1 FILLER_6_338 ();
 sg13g2_fill_1 FILLER_6_389 ();
 sg13g2_decap_8 FILLER_6_416 ();
 sg13g2_decap_8 FILLER_6_423 ();
 sg13g2_decap_8 FILLER_7_30 ();
 sg13g2_decap_4 FILLER_7_37 ();
 sg13g2_fill_2 FILLER_7_41 ();
 sg13g2_decap_8 FILLER_7_47 ();
 sg13g2_decap_4 FILLER_7_54 ();
 sg13g2_fill_2 FILLER_7_66 ();
 sg13g2_decap_4 FILLER_7_71 ();
 sg13g2_fill_2 FILLER_7_83 ();
 sg13g2_fill_1 FILLER_7_85 ();
 sg13g2_decap_8 FILLER_7_131 ();
 sg13g2_fill_2 FILLER_7_138 ();
 sg13g2_fill_1 FILLER_7_140 ();
 sg13g2_decap_8 FILLER_7_160 ();
 sg13g2_decap_8 FILLER_7_167 ();
 sg13g2_fill_2 FILLER_7_174 ();
 sg13g2_fill_1 FILLER_7_176 ();
 sg13g2_decap_4 FILLER_7_189 ();
 sg13g2_fill_1 FILLER_7_193 ();
 sg13g2_fill_2 FILLER_7_233 ();
 sg13g2_fill_2 FILLER_7_240 ();
 sg13g2_fill_2 FILLER_7_247 ();
 sg13g2_fill_1 FILLER_7_249 ();
 sg13g2_fill_2 FILLER_7_255 ();
 sg13g2_fill_1 FILLER_7_257 ();
 sg13g2_fill_2 FILLER_7_263 ();
 sg13g2_decap_8 FILLER_7_273 ();
 sg13g2_decap_8 FILLER_7_280 ();
 sg13g2_decap_4 FILLER_7_287 ();
 sg13g2_decap_4 FILLER_7_317 ();
 sg13g2_fill_1 FILLER_7_321 ();
 sg13g2_decap_4 FILLER_7_341 ();
 sg13g2_fill_1 FILLER_7_345 ();
 sg13g2_fill_1 FILLER_7_349 ();
 sg13g2_fill_1 FILLER_7_360 ();
 sg13g2_fill_1 FILLER_7_370 ();
 sg13g2_fill_1 FILLER_7_375 ();
 sg13g2_fill_2 FILLER_7_381 ();
 sg13g2_decap_4 FILLER_7_398 ();
 sg13g2_fill_2 FILLER_7_402 ();
 sg13g2_decap_8 FILLER_7_408 ();
 sg13g2_decap_8 FILLER_7_415 ();
 sg13g2_decap_8 FILLER_7_422 ();
 sg13g2_fill_1 FILLER_7_429 ();
 sg13g2_decap_8 FILLER_8_0 ();
 sg13g2_fill_1 FILLER_8_7 ();
 sg13g2_fill_2 FILLER_8_12 ();
 sg13g2_fill_1 FILLER_8_14 ();
 sg13g2_decap_8 FILLER_8_18 ();
 sg13g2_decap_8 FILLER_8_25 ();
 sg13g2_decap_4 FILLER_8_32 ();
 sg13g2_decap_8 FILLER_8_66 ();
 sg13g2_fill_1 FILLER_8_73 ();
 sg13g2_fill_2 FILLER_8_78 ();
 sg13g2_decap_8 FILLER_8_84 ();
 sg13g2_fill_1 FILLER_8_91 ();
 sg13g2_fill_1 FILLER_8_117 ();
 sg13g2_decap_8 FILLER_8_126 ();
 sg13g2_fill_2 FILLER_8_178 ();
 sg13g2_decap_8 FILLER_8_206 ();
 sg13g2_decap_8 FILLER_8_213 ();
 sg13g2_decap_8 FILLER_8_220 ();
 sg13g2_fill_2 FILLER_8_231 ();
 sg13g2_fill_1 FILLER_8_268 ();
 sg13g2_fill_2 FILLER_8_280 ();
 sg13g2_fill_1 FILLER_8_282 ();
 sg13g2_fill_1 FILLER_8_309 ();
 sg13g2_decap_8 FILLER_8_315 ();
 sg13g2_fill_1 FILLER_8_332 ();
 sg13g2_fill_1 FILLER_8_348 ();
 sg13g2_decap_8 FILLER_8_354 ();
 sg13g2_decap_4 FILLER_8_361 ();
 sg13g2_fill_2 FILLER_8_365 ();
 sg13g2_decap_4 FILLER_8_377 ();
 sg13g2_fill_2 FILLER_8_388 ();
 sg13g2_fill_1 FILLER_8_390 ();
 sg13g2_decap_4 FILLER_8_400 ();
 sg13g2_decap_8 FILLER_8_416 ();
 sg13g2_decap_8 FILLER_8_423 ();
 sg13g2_fill_2 FILLER_9_0 ();
 sg13g2_fill_2 FILLER_9_6 ();
 sg13g2_fill_1 FILLER_9_8 ();
 sg13g2_fill_2 FILLER_9_35 ();
 sg13g2_fill_1 FILLER_9_37 ();
 sg13g2_fill_1 FILLER_9_100 ();
 sg13g2_fill_2 FILLER_9_108 ();
 sg13g2_fill_2 FILLER_9_117 ();
 sg13g2_fill_2 FILLER_9_149 ();
 sg13g2_fill_1 FILLER_9_151 ();
 sg13g2_decap_8 FILLER_9_171 ();
 sg13g2_decap_4 FILLER_9_178 ();
 sg13g2_fill_2 FILLER_9_182 ();
 sg13g2_decap_4 FILLER_9_192 ();
 sg13g2_fill_1 FILLER_9_196 ();
 sg13g2_fill_2 FILLER_9_200 ();
 sg13g2_fill_1 FILLER_9_228 ();
 sg13g2_fill_1 FILLER_9_234 ();
 sg13g2_fill_1 FILLER_9_240 ();
 sg13g2_fill_1 FILLER_9_248 ();
 sg13g2_fill_1 FILLER_9_253 ();
 sg13g2_fill_1 FILLER_9_259 ();
 sg13g2_fill_1 FILLER_9_264 ();
 sg13g2_decap_8 FILLER_9_270 ();
 sg13g2_fill_1 FILLER_9_277 ();
 sg13g2_fill_1 FILLER_9_281 ();
 sg13g2_decap_8 FILLER_9_301 ();
 sg13g2_fill_1 FILLER_9_308 ();
 sg13g2_decap_8 FILLER_9_335 ();
 sg13g2_decap_4 FILLER_9_342 ();
 sg13g2_fill_2 FILLER_9_346 ();
 sg13g2_fill_2 FILLER_9_364 ();
 sg13g2_fill_1 FILLER_9_366 ();
 sg13g2_fill_1 FILLER_9_374 ();
 sg13g2_fill_2 FILLER_9_384 ();
 sg13g2_fill_1 FILLER_9_392 ();
 sg13g2_decap_4 FILLER_9_424 ();
 sg13g2_fill_2 FILLER_9_428 ();
 sg13g2_decap_8 FILLER_10_0 ();
 sg13g2_fill_2 FILLER_10_7 ();
 sg13g2_decap_4 FILLER_10_13 ();
 sg13g2_fill_1 FILLER_10_17 ();
 sg13g2_decap_4 FILLER_10_26 ();
 sg13g2_fill_1 FILLER_10_30 ();
 sg13g2_fill_2 FILLER_10_43 ();
 sg13g2_decap_8 FILLER_10_49 ();
 sg13g2_fill_2 FILLER_10_56 ();
 sg13g2_decap_4 FILLER_10_84 ();
 sg13g2_decap_8 FILLER_10_93 ();
 sg13g2_decap_4 FILLER_10_100 ();
 sg13g2_decap_8 FILLER_10_116 ();
 sg13g2_decap_8 FILLER_10_123 ();
 sg13g2_fill_2 FILLER_10_130 ();
 sg13g2_decap_4 FILLER_10_136 ();
 sg13g2_fill_2 FILLER_10_140 ();
 sg13g2_fill_1 FILLER_10_147 ();
 sg13g2_fill_2 FILLER_10_209 ();
 sg13g2_decap_8 FILLER_10_215 ();
 sg13g2_decap_8 FILLER_10_222 ();
 sg13g2_fill_2 FILLER_10_229 ();
 sg13g2_fill_1 FILLER_10_231 ();
 sg13g2_fill_1 FILLER_10_235 ();
 sg13g2_fill_1 FILLER_10_249 ();
 sg13g2_fill_1 FILLER_10_254 ();
 sg13g2_fill_1 FILLER_10_258 ();
 sg13g2_fill_1 FILLER_10_263 ();
 sg13g2_fill_1 FILLER_10_269 ();
 sg13g2_decap_4 FILLER_10_275 ();
 sg13g2_fill_2 FILLER_10_284 ();
 sg13g2_fill_1 FILLER_10_286 ();
 sg13g2_decap_8 FILLER_10_313 ();
 sg13g2_decap_8 FILLER_10_320 ();
 sg13g2_fill_2 FILLER_10_327 ();
 sg13g2_decap_8 FILLER_10_365 ();
 sg13g2_fill_2 FILLER_10_372 ();
 sg13g2_fill_2 FILLER_10_384 ();
 sg13g2_fill_1 FILLER_10_386 ();
 sg13g2_decap_4 FILLER_10_392 ();
 sg13g2_decap_8 FILLER_10_404 ();
 sg13g2_fill_2 FILLER_10_411 ();
 sg13g2_fill_1 FILLER_10_413 ();
 sg13g2_decap_8 FILLER_10_419 ();
 sg13g2_decap_4 FILLER_10_426 ();
 sg13g2_decap_8 FILLER_11_0 ();
 sg13g2_decap_4 FILLER_11_7 ();
 sg13g2_fill_2 FILLER_11_11 ();
 sg13g2_decap_4 FILLER_11_25 ();
 sg13g2_fill_1 FILLER_11_33 ();
 sg13g2_fill_2 FILLER_11_40 ();
 sg13g2_fill_1 FILLER_11_73 ();
 sg13g2_decap_8 FILLER_11_86 ();
 sg13g2_fill_1 FILLER_11_93 ();
 sg13g2_decap_8 FILLER_11_98 ();
 sg13g2_fill_1 FILLER_11_105 ();
 sg13g2_decap_8 FILLER_11_132 ();
 sg13g2_decap_8 FILLER_11_139 ();
 sg13g2_decap_8 FILLER_11_146 ();
 sg13g2_fill_2 FILLER_11_153 ();
 sg13g2_fill_1 FILLER_11_155 ();
 sg13g2_fill_2 FILLER_11_182 ();
 sg13g2_fill_1 FILLER_11_184 ();
 sg13g2_decap_8 FILLER_11_190 ();
 sg13g2_fill_2 FILLER_11_197 ();
 sg13g2_decap_8 FILLER_11_217 ();
 sg13g2_decap_4 FILLER_11_224 ();
 sg13g2_fill_2 FILLER_11_240 ();
 sg13g2_fill_1 FILLER_11_242 ();
 sg13g2_fill_1 FILLER_11_253 ();
 sg13g2_fill_1 FILLER_11_258 ();
 sg13g2_fill_1 FILLER_11_268 ();
 sg13g2_decap_8 FILLER_11_273 ();
 sg13g2_decap_4 FILLER_11_280 ();
 sg13g2_fill_2 FILLER_11_284 ();
 sg13g2_fill_1 FILLER_11_291 ();
 sg13g2_decap_8 FILLER_11_296 ();
 sg13g2_fill_1 FILLER_11_303 ();
 sg13g2_decap_8 FILLER_11_335 ();
 sg13g2_decap_8 FILLER_11_342 ();
 sg13g2_decap_8 FILLER_11_362 ();
 sg13g2_decap_8 FILLER_11_369 ();
 sg13g2_decap_4 FILLER_11_376 ();
 sg13g2_fill_1 FILLER_11_380 ();
 sg13g2_fill_1 FILLER_11_398 ();
 sg13g2_fill_1 FILLER_11_429 ();
 sg13g2_fill_2 FILLER_12_0 ();
 sg13g2_fill_1 FILLER_12_2 ();
 sg13g2_fill_1 FILLER_12_29 ();
 sg13g2_fill_1 FILLER_12_34 ();
 sg13g2_decap_8 FILLER_12_43 ();
 sg13g2_decap_4 FILLER_12_50 ();
 sg13g2_fill_1 FILLER_12_54 ();
 sg13g2_decap_4 FILLER_12_111 ();
 sg13g2_decap_8 FILLER_12_119 ();
 sg13g2_decap_8 FILLER_12_126 ();
 sg13g2_decap_8 FILLER_12_133 ();
 sg13g2_decap_8 FILLER_12_140 ();
 sg13g2_decap_4 FILLER_12_147 ();
 sg13g2_decap_8 FILLER_12_166 ();
 sg13g2_decap_4 FILLER_12_173 ();
 sg13g2_fill_2 FILLER_12_192 ();
 sg13g2_fill_1 FILLER_12_194 ();
 sg13g2_fill_1 FILLER_12_200 ();
 sg13g2_fill_1 FILLER_12_212 ();
 sg13g2_decap_8 FILLER_12_222 ();
 sg13g2_fill_1 FILLER_12_229 ();
 sg13g2_decap_8 FILLER_12_235 ();
 sg13g2_decap_8 FILLER_12_242 ();
 sg13g2_fill_1 FILLER_12_254 ();
 sg13g2_fill_2 FILLER_12_259 ();
 sg13g2_fill_1 FILLER_12_267 ();
 sg13g2_fill_2 FILLER_12_277 ();
 sg13g2_fill_1 FILLER_12_279 ();
 sg13g2_fill_1 FILLER_12_289 ();
 sg13g2_fill_1 FILLER_12_314 ();
 sg13g2_fill_1 FILLER_12_324 ();
 sg13g2_decap_8 FILLER_12_330 ();
 sg13g2_fill_2 FILLER_12_337 ();
 sg13g2_fill_2 FILLER_12_375 ();
 sg13g2_fill_2 FILLER_12_384 ();
 sg13g2_fill_1 FILLER_12_386 ();
 sg13g2_decap_4 FILLER_12_392 ();
 sg13g2_decap_8 FILLER_12_408 ();
 sg13g2_fill_1 FILLER_12_415 ();
 sg13g2_decap_8 FILLER_12_421 ();
 sg13g2_fill_2 FILLER_12_428 ();
 sg13g2_decap_8 FILLER_13_0 ();
 sg13g2_fill_1 FILLER_13_7 ();
 sg13g2_fill_2 FILLER_13_12 ();
 sg13g2_decap_4 FILLER_13_18 ();
 sg13g2_fill_2 FILLER_13_22 ();
 sg13g2_decap_8 FILLER_13_54 ();
 sg13g2_fill_1 FILLER_13_61 ();
 sg13g2_decap_8 FILLER_13_66 ();
 sg13g2_decap_4 FILLER_13_73 ();
 sg13g2_fill_1 FILLER_13_77 ();
 sg13g2_decap_4 FILLER_13_99 ();
 sg13g2_fill_2 FILLER_13_103 ();
 sg13g2_fill_2 FILLER_13_115 ();
 sg13g2_fill_1 FILLER_13_117 ();
 sg13g2_decap_8 FILLER_13_122 ();
 sg13g2_decap_8 FILLER_13_129 ();
 sg13g2_decap_8 FILLER_13_136 ();
 sg13g2_fill_2 FILLER_13_153 ();
 sg13g2_fill_1 FILLER_13_155 ();
 sg13g2_decap_4 FILLER_13_166 ();
 sg13g2_decap_8 FILLER_13_196 ();
 sg13g2_fill_1 FILLER_13_203 ();
 sg13g2_decap_8 FILLER_13_217 ();
 sg13g2_decap_8 FILLER_13_224 ();
 sg13g2_decap_8 FILLER_13_231 ();
 sg13g2_decap_8 FILLER_13_243 ();
 sg13g2_decap_4 FILLER_13_250 ();
 sg13g2_fill_1 FILLER_13_254 ();
 sg13g2_fill_2 FILLER_13_270 ();
 sg13g2_fill_1 FILLER_13_272 ();
 sg13g2_fill_2 FILLER_13_280 ();
 sg13g2_fill_2 FILLER_13_287 ();
 sg13g2_fill_2 FILLER_13_315 ();
 sg13g2_decap_8 FILLER_13_353 ();
 sg13g2_fill_1 FILLER_13_360 ();
 sg13g2_decap_8 FILLER_13_366 ();
 sg13g2_fill_1 FILLER_13_373 ();
 sg13g2_fill_2 FILLER_13_395 ();
 sg13g2_decap_4 FILLER_13_426 ();
 sg13g2_decap_4 FILLER_14_0 ();
 sg13g2_decap_8 FILLER_14_30 ();
 sg13g2_fill_1 FILLER_14_37 ();
 sg13g2_decap_8 FILLER_14_42 ();
 sg13g2_decap_8 FILLER_14_49 ();
 sg13g2_fill_2 FILLER_14_56 ();
 sg13g2_fill_1 FILLER_14_58 ();
 sg13g2_decap_4 FILLER_14_142 ();
 sg13g2_fill_1 FILLER_14_146 ();
 sg13g2_decap_8 FILLER_14_158 ();
 sg13g2_decap_8 FILLER_14_165 ();
 sg13g2_decap_8 FILLER_14_172 ();
 sg13g2_decap_8 FILLER_14_179 ();
 sg13g2_decap_4 FILLER_14_186 ();
 sg13g2_fill_1 FILLER_14_190 ();
 sg13g2_decap_4 FILLER_14_201 ();
 sg13g2_fill_1 FILLER_14_205 ();
 sg13g2_fill_2 FILLER_14_232 ();
 sg13g2_fill_2 FILLER_14_238 ();
 sg13g2_fill_2 FILLER_14_258 ();
 sg13g2_decap_8 FILLER_14_282 ();
 sg13g2_decap_4 FILLER_14_289 ();
 sg13g2_fill_2 FILLER_14_293 ();
 sg13g2_decap_8 FILLER_14_299 ();
 sg13g2_decap_8 FILLER_14_306 ();
 sg13g2_decap_4 FILLER_14_313 ();
 sg13g2_fill_2 FILLER_14_317 ();
 sg13g2_fill_1 FILLER_14_324 ();
 sg13g2_decap_8 FILLER_14_336 ();
 sg13g2_decap_4 FILLER_14_343 ();
 sg13g2_fill_2 FILLER_14_347 ();
 sg13g2_decap_8 FILLER_14_375 ();
 sg13g2_fill_1 FILLER_14_382 ();
 sg13g2_decap_8 FILLER_14_423 ();
 sg13g2_decap_8 FILLER_15_0 ();
 sg13g2_decap_4 FILLER_15_7 ();
 sg13g2_fill_2 FILLER_15_15 ();
 sg13g2_fill_2 FILLER_15_27 ();
 sg13g2_decap_8 FILLER_15_69 ();
 sg13g2_decap_8 FILLER_15_76 ();
 sg13g2_decap_8 FILLER_15_83 ();
 sg13g2_decap_8 FILLER_15_94 ();
 sg13g2_decap_8 FILLER_15_101 ();
 sg13g2_decap_8 FILLER_15_118 ();
 sg13g2_decap_8 FILLER_15_125 ();
 sg13g2_decap_8 FILLER_15_132 ();
 sg13g2_fill_1 FILLER_15_144 ();
 sg13g2_fill_2 FILLER_15_150 ();
 sg13g2_fill_1 FILLER_15_152 ();
 sg13g2_fill_1 FILLER_15_163 ();
 sg13g2_fill_1 FILLER_15_190 ();
 sg13g2_fill_2 FILLER_15_210 ();
 sg13g2_decap_8 FILLER_15_238 ();
 sg13g2_fill_1 FILLER_15_245 ();
 sg13g2_fill_2 FILLER_15_251 ();
 sg13g2_decap_4 FILLER_15_277 ();
 sg13g2_decap_4 FILLER_15_299 ();
 sg13g2_fill_1 FILLER_15_303 ();
 sg13g2_decap_4 FILLER_15_317 ();
 sg13g2_fill_2 FILLER_15_321 ();
 sg13g2_decap_4 FILLER_15_349 ();
 sg13g2_decap_4 FILLER_15_379 ();
 sg13g2_fill_2 FILLER_15_393 ();
 sg13g2_fill_1 FILLER_15_395 ();
 sg13g2_decap_8 FILLER_15_422 ();
 sg13g2_fill_1 FILLER_15_429 ();
 sg13g2_decap_8 FILLER_16_36 ();
 sg13g2_fill_1 FILLER_16_43 ();
 sg13g2_fill_2 FILLER_16_70 ();
 sg13g2_fill_1 FILLER_16_72 ();
 sg13g2_decap_4 FILLER_16_109 ();
 sg13g2_decap_4 FILLER_16_144 ();
 sg13g2_fill_1 FILLER_16_148 ();
 sg13g2_decap_8 FILLER_16_212 ();
 sg13g2_decap_4 FILLER_16_219 ();
 sg13g2_fill_1 FILLER_16_223 ();
 sg13g2_decap_8 FILLER_16_228 ();
 sg13g2_decap_4 FILLER_16_235 ();
 sg13g2_fill_2 FILLER_16_256 ();
 sg13g2_decap_8 FILLER_16_264 ();
 sg13g2_decap_8 FILLER_16_271 ();
 sg13g2_decap_4 FILLER_16_278 ();
 sg13g2_fill_1 FILLER_16_282 ();
 sg13g2_decap_4 FILLER_16_288 ();
 sg13g2_decap_8 FILLER_16_323 ();
 sg13g2_fill_1 FILLER_16_330 ();
 sg13g2_decap_8 FILLER_16_335 ();
 sg13g2_decap_4 FILLER_16_342 ();
 sg13g2_fill_1 FILLER_16_346 ();
 sg13g2_decap_8 FILLER_16_357 ();
 sg13g2_decap_8 FILLER_16_364 ();
 sg13g2_decap_4 FILLER_16_371 ();
 sg13g2_decap_8 FILLER_16_379 ();
 sg13g2_decap_8 FILLER_16_386 ();
 sg13g2_decap_4 FILLER_16_393 ();
 sg13g2_decap_4 FILLER_16_405 ();
 sg13g2_fill_2 FILLER_16_409 ();
 sg13g2_decap_8 FILLER_16_415 ();
 sg13g2_decap_8 FILLER_16_422 ();
 sg13g2_fill_1 FILLER_16_429 ();
 sg13g2_decap_8 FILLER_17_0 ();
 sg13g2_decap_8 FILLER_17_11 ();
 sg13g2_fill_1 FILLER_17_18 ();
 sg13g2_decap_8 FILLER_17_23 ();
 sg13g2_decap_4 FILLER_17_30 ();
 sg13g2_fill_2 FILLER_17_34 ();
 sg13g2_decap_4 FILLER_17_46 ();
 sg13g2_fill_2 FILLER_17_50 ();
 sg13g2_decap_8 FILLER_17_56 ();
 sg13g2_fill_2 FILLER_17_63 ();
 sg13g2_fill_1 FILLER_17_65 ();
 sg13g2_decap_8 FILLER_17_70 ();
 sg13g2_decap_4 FILLER_17_77 ();
 sg13g2_fill_2 FILLER_17_81 ();
 sg13g2_decap_8 FILLER_17_87 ();
 sg13g2_decap_8 FILLER_17_94 ();
 sg13g2_decap_4 FILLER_17_101 ();
 sg13g2_decap_8 FILLER_17_109 ();
 sg13g2_fill_2 FILLER_17_116 ();
 sg13g2_fill_1 FILLER_17_118 ();
 sg13g2_decap_8 FILLER_17_123 ();
 sg13g2_decap_8 FILLER_17_130 ();
 sg13g2_decap_8 FILLER_17_137 ();
 sg13g2_decap_8 FILLER_17_149 ();
 sg13g2_decap_8 FILLER_17_156 ();
 sg13g2_decap_8 FILLER_17_163 ();
 sg13g2_decap_8 FILLER_17_170 ();
 sg13g2_decap_8 FILLER_17_177 ();
 sg13g2_decap_8 FILLER_17_184 ();
 sg13g2_decap_4 FILLER_17_191 ();
 sg13g2_fill_2 FILLER_17_205 ();
 sg13g2_fill_1 FILLER_17_207 ();
 sg13g2_decap_8 FILLER_17_234 ();
 sg13g2_fill_2 FILLER_17_241 ();
 sg13g2_fill_1 FILLER_17_243 ();
 sg13g2_decap_8 FILLER_17_257 ();
 sg13g2_decap_8 FILLER_17_264 ();
 sg13g2_decap_4 FILLER_17_271 ();
 sg13g2_decap_4 FILLER_17_281 ();
 sg13g2_fill_2 FILLER_17_285 ();
 sg13g2_decap_8 FILLER_17_294 ();
 sg13g2_decap_4 FILLER_17_301 ();
 sg13g2_fill_2 FILLER_17_305 ();
 sg13g2_decap_8 FILLER_17_311 ();
 sg13g2_decap_8 FILLER_17_318 ();
 sg13g2_fill_1 FILLER_17_325 ();
 sg13g2_fill_1 FILLER_17_334 ();
 sg13g2_fill_2 FILLER_17_343 ();
 sg13g2_fill_1 FILLER_17_353 ();
 sg13g2_fill_2 FILLER_17_362 ();
 sg13g2_fill_2 FILLER_17_372 ();
 sg13g2_fill_1 FILLER_17_374 ();
 sg13g2_fill_2 FILLER_17_401 ();
 sg13g2_fill_1 FILLER_17_403 ();
 sg13g2_decap_8 FILLER_18_0 ();
 sg13g2_decap_4 FILLER_18_43 ();
 sg13g2_fill_2 FILLER_18_47 ();
 sg13g2_fill_2 FILLER_18_124 ();
 sg13g2_fill_1 FILLER_18_126 ();
 sg13g2_decap_8 FILLER_18_131 ();
 sg13g2_decap_4 FILLER_18_138 ();
 sg13g2_fill_2 FILLER_18_147 ();
 sg13g2_fill_2 FILLER_18_168 ();
 sg13g2_fill_2 FILLER_18_196 ();
 sg13g2_fill_2 FILLER_18_203 ();
 sg13g2_decap_8 FILLER_18_219 ();
 sg13g2_fill_1 FILLER_18_226 ();
 sg13g2_fill_2 FILLER_18_232 ();
 sg13g2_fill_1 FILLER_18_246 ();
 sg13g2_fill_1 FILLER_18_252 ();
 sg13g2_fill_2 FILLER_18_259 ();
 sg13g2_fill_1 FILLER_18_267 ();
 sg13g2_fill_2 FILLER_18_294 ();
 sg13g2_fill_1 FILLER_18_337 ();
 sg13g2_decap_4 FILLER_18_343 ();
 sg13g2_fill_2 FILLER_18_369 ();
 sg13g2_fill_1 FILLER_18_371 ();
 sg13g2_fill_2 FILLER_18_380 ();
 sg13g2_fill_2 FILLER_18_386 ();
 sg13g2_fill_1 FILLER_18_388 ();
 sg13g2_fill_2 FILLER_18_393 ();
 sg13g2_fill_1 FILLER_18_395 ();
 sg13g2_fill_2 FILLER_18_401 ();
 sg13g2_decap_4 FILLER_18_407 ();
 sg13g2_decap_8 FILLER_18_415 ();
 sg13g2_decap_8 FILLER_18_422 ();
 sg13g2_fill_1 FILLER_18_429 ();
 sg13g2_decap_8 FILLER_19_0 ();
 sg13g2_decap_8 FILLER_19_17 ();
 sg13g2_fill_2 FILLER_19_24 ();
 sg13g2_fill_2 FILLER_19_62 ();
 sg13g2_decap_4 FILLER_19_104 ();
 sg13g2_fill_2 FILLER_19_108 ();
 sg13g2_fill_2 FILLER_19_156 ();
 sg13g2_decap_4 FILLER_19_196 ();
 sg13g2_decap_4 FILLER_19_222 ();
 sg13g2_fill_1 FILLER_19_226 ();
 sg13g2_fill_1 FILLER_19_232 ();
 sg13g2_decap_4 FILLER_19_243 ();
 sg13g2_fill_1 FILLER_19_247 ();
 sg13g2_decap_4 FILLER_19_252 ();
 sg13g2_decap_8 FILLER_19_276 ();
 sg13g2_decap_4 FILLER_19_283 ();
 sg13g2_fill_2 FILLER_19_291 ();
 sg13g2_decap_8 FILLER_19_297 ();
 sg13g2_decap_8 FILLER_19_304 ();
 sg13g2_fill_2 FILLER_19_311 ();
 sg13g2_fill_1 FILLER_19_313 ();
 sg13g2_decap_4 FILLER_19_350 ();
 sg13g2_fill_2 FILLER_19_368 ();
 sg13g2_decap_8 FILLER_19_378 ();
 sg13g2_decap_8 FILLER_19_385 ();
 sg13g2_decap_4 FILLER_20_0 ();
 sg13g2_fill_1 FILLER_20_4 ();
 sg13g2_decap_8 FILLER_20_20 ();
 sg13g2_fill_2 FILLER_20_41 ();
 sg13g2_decap_8 FILLER_20_47 ();
 sg13g2_decap_4 FILLER_20_54 ();
 sg13g2_decap_8 FILLER_20_68 ();
 sg13g2_fill_2 FILLER_20_75 ();
 sg13g2_decap_8 FILLER_20_117 ();
 sg13g2_fill_1 FILLER_20_124 ();
 sg13g2_decap_4 FILLER_20_129 ();
 sg13g2_fill_2 FILLER_20_133 ();
 sg13g2_fill_1 FILLER_20_145 ();
 sg13g2_decap_4 FILLER_20_151 ();
 sg13g2_fill_2 FILLER_20_155 ();
 sg13g2_decap_8 FILLER_20_167 ();
 sg13g2_decap_8 FILLER_20_174 ();
 sg13g2_decap_8 FILLER_20_181 ();
 sg13g2_decap_4 FILLER_20_188 ();
 sg13g2_fill_2 FILLER_20_192 ();
 sg13g2_decap_4 FILLER_20_198 ();
 sg13g2_fill_1 FILLER_20_238 ();
 sg13g2_fill_1 FILLER_20_249 ();
 sg13g2_fill_2 FILLER_20_258 ();
 sg13g2_fill_2 FILLER_20_264 ();
 sg13g2_decap_8 FILLER_20_270 ();
 sg13g2_decap_8 FILLER_20_277 ();
 sg13g2_fill_1 FILLER_20_284 ();
 sg13g2_fill_2 FILLER_20_305 ();
 sg13g2_decap_8 FILLER_20_333 ();
 sg13g2_fill_2 FILLER_20_340 ();
 sg13g2_fill_1 FILLER_20_342 ();
 sg13g2_decap_8 FILLER_20_367 ();
 sg13g2_decap_8 FILLER_20_374 ();
 sg13g2_fill_2 FILLER_20_381 ();
 sg13g2_decap_8 FILLER_20_421 ();
 sg13g2_fill_2 FILLER_20_428 ();
 sg13g2_fill_2 FILLER_21_0 ();
 sg13g2_fill_2 FILLER_21_28 ();
 sg13g2_fill_2 FILLER_21_35 ();
 sg13g2_fill_2 FILLER_21_63 ();
 sg13g2_fill_1 FILLER_21_65 ();
 sg13g2_fill_2 FILLER_21_92 ();
 sg13g2_fill_1 FILLER_21_94 ();
 sg13g2_fill_2 FILLER_21_99 ();
 sg13g2_fill_1 FILLER_21_101 ();
 sg13g2_fill_2 FILLER_21_106 ();
 sg13g2_fill_1 FILLER_21_108 ();
 sg13g2_fill_1 FILLER_21_145 ();
 sg13g2_decap_4 FILLER_21_151 ();
 sg13g2_decap_8 FILLER_21_163 ();
 sg13g2_decap_8 FILLER_21_170 ();
 sg13g2_decap_8 FILLER_21_177 ();
 sg13g2_decap_8 FILLER_21_184 ();
 sg13g2_fill_1 FILLER_21_191 ();
 sg13g2_decap_8 FILLER_21_202 ();
 sg13g2_decap_8 FILLER_21_209 ();
 sg13g2_decap_8 FILLER_21_216 ();
 sg13g2_fill_1 FILLER_21_223 ();
 sg13g2_decap_8 FILLER_21_234 ();
 sg13g2_decap_8 FILLER_21_241 ();
 sg13g2_fill_1 FILLER_21_248 ();
 sg13g2_fill_1 FILLER_21_259 ();
 sg13g2_decap_8 FILLER_21_296 ();
 sg13g2_decap_8 FILLER_21_303 ();
 sg13g2_decap_4 FILLER_21_310 ();
 sg13g2_decap_8 FILLER_21_318 ();
 sg13g2_decap_8 FILLER_21_325 ();
 sg13g2_decap_8 FILLER_21_332 ();
 sg13g2_fill_2 FILLER_21_339 ();
 sg13g2_fill_1 FILLER_21_341 ();
 sg13g2_fill_2 FILLER_21_346 ();
 sg13g2_fill_1 FILLER_21_353 ();
 sg13g2_decap_8 FILLER_21_360 ();
 sg13g2_decap_8 FILLER_21_367 ();
 sg13g2_decap_8 FILLER_21_374 ();
 sg13g2_fill_1 FILLER_21_381 ();
 sg13g2_fill_1 FILLER_21_388 ();
 sg13g2_decap_8 FILLER_21_394 ();
 sg13g2_fill_1 FILLER_21_401 ();
 sg13g2_decap_4 FILLER_21_406 ();
 sg13g2_fill_1 FILLER_21_410 ();
 sg13g2_decap_8 FILLER_21_415 ();
 sg13g2_decap_8 FILLER_21_422 ();
 sg13g2_fill_1 FILLER_21_429 ();
 sg13g2_decap_8 FILLER_22_14 ();
 sg13g2_decap_8 FILLER_22_21 ();
 sg13g2_decap_8 FILLER_22_28 ();
 sg13g2_fill_1 FILLER_22_45 ();
 sg13g2_decap_8 FILLER_22_50 ();
 sg13g2_decap_8 FILLER_22_57 ();
 sg13g2_decap_8 FILLER_22_64 ();
 sg13g2_fill_2 FILLER_22_71 ();
 sg13g2_fill_1 FILLER_22_77 ();
 sg13g2_fill_1 FILLER_22_83 ();
 sg13g2_fill_1 FILLER_22_89 ();
 sg13g2_decap_8 FILLER_22_116 ();
 sg13g2_fill_2 FILLER_22_123 ();
 sg13g2_fill_2 FILLER_22_133 ();
 sg13g2_fill_1 FILLER_22_135 ();
 sg13g2_fill_1 FILLER_22_140 ();
 sg13g2_decap_8 FILLER_22_146 ();
 sg13g2_fill_1 FILLER_22_153 ();
 sg13g2_decap_4 FILLER_22_194 ();
 sg13g2_fill_2 FILLER_22_198 ();
 sg13g2_decap_4 FILLER_22_226 ();
 sg13g2_fill_2 FILLER_22_230 ();
 sg13g2_decap_8 FILLER_22_258 ();
 sg13g2_decap_8 FILLER_22_265 ();
 sg13g2_decap_8 FILLER_22_272 ();
 sg13g2_decap_8 FILLER_22_279 ();
 sg13g2_fill_1 FILLER_22_286 ();
 sg13g2_fill_2 FILLER_22_291 ();
 sg13g2_decap_8 FILLER_22_301 ();
 sg13g2_fill_2 FILLER_22_308 ();
 sg13g2_fill_1 FILLER_22_310 ();
 sg13g2_decap_8 FILLER_22_315 ();
 sg13g2_decap_8 FILLER_22_322 ();
 sg13g2_fill_1 FILLER_22_329 ();
 sg13g2_fill_2 FILLER_22_348 ();
 sg13g2_fill_1 FILLER_22_350 ();
 sg13g2_decap_8 FILLER_22_356 ();
 sg13g2_decap_8 FILLER_22_363 ();
 sg13g2_decap_8 FILLER_22_374 ();
 sg13g2_decap_8 FILLER_22_381 ();
 sg13g2_fill_2 FILLER_22_396 ();
 sg13g2_fill_2 FILLER_22_402 ();
 sg13g2_fill_1 FILLER_23_0 ();
 sg13g2_decap_4 FILLER_23_27 ();
 sg13g2_decap_8 FILLER_23_36 ();
 sg13g2_fill_1 FILLER_23_43 ();
 sg13g2_decap_8 FILLER_23_48 ();
 sg13g2_fill_2 FILLER_23_55 ();
 sg13g2_fill_1 FILLER_23_57 ();
 sg13g2_decap_8 FILLER_23_88 ();
 sg13g2_fill_2 FILLER_23_95 ();
 sg13g2_decap_4 FILLER_23_101 ();
 sg13g2_fill_1 FILLER_23_105 ();
 sg13g2_fill_2 FILLER_23_148 ();
 sg13g2_decap_4 FILLER_23_159 ();
 sg13g2_decap_8 FILLER_23_199 ();
 sg13g2_decap_4 FILLER_23_206 ();
 sg13g2_fill_2 FILLER_23_210 ();
 sg13g2_decap_8 FILLER_23_217 ();
 sg13g2_decap_8 FILLER_23_224 ();
 sg13g2_decap_4 FILLER_23_231 ();
 sg13g2_fill_2 FILLER_23_235 ();
 sg13g2_decap_8 FILLER_23_241 ();
 sg13g2_decap_8 FILLER_23_248 ();
 sg13g2_decap_4 FILLER_23_255 ();
 sg13g2_fill_2 FILLER_23_259 ();
 sg13g2_fill_2 FILLER_23_325 ();
 sg13g2_fill_1 FILLER_23_353 ();
 sg13g2_fill_1 FILLER_23_389 ();
 sg13g2_decap_8 FILLER_23_402 ();
 sg13g2_fill_2 FILLER_23_409 ();
 sg13g2_decap_8 FILLER_23_419 ();
 sg13g2_decap_4 FILLER_23_426 ();
 sg13g2_decap_8 FILLER_24_0 ();
 sg13g2_decap_4 FILLER_24_22 ();
 sg13g2_fill_1 FILLER_24_26 ();
 sg13g2_decap_4 FILLER_24_63 ();
 sg13g2_fill_2 FILLER_24_82 ();
 sg13g2_fill_2 FILLER_24_96 ();
 sg13g2_fill_1 FILLER_24_98 ();
 sg13g2_decap_8 FILLER_24_125 ();
 sg13g2_decap_8 FILLER_24_132 ();
 sg13g2_fill_2 FILLER_24_139 ();
 sg13g2_decap_8 FILLER_24_207 ();
 sg13g2_decap_8 FILLER_24_214 ();
 sg13g2_decap_4 FILLER_24_221 ();
 sg13g2_fill_1 FILLER_24_225 ();
 sg13g2_fill_1 FILLER_24_256 ();
 sg13g2_fill_1 FILLER_24_262 ();
 sg13g2_fill_2 FILLER_24_268 ();
 sg13g2_fill_1 FILLER_24_270 ();
 sg13g2_decap_4 FILLER_24_275 ();
 sg13g2_fill_1 FILLER_24_279 ();
 sg13g2_fill_2 FILLER_24_285 ();
 sg13g2_fill_1 FILLER_24_290 ();
 sg13g2_decap_4 FILLER_24_295 ();
 sg13g2_fill_1 FILLER_24_303 ();
 sg13g2_decap_8 FILLER_24_308 ();
 sg13g2_fill_1 FILLER_24_315 ();
 sg13g2_decap_4 FILLER_24_324 ();
 sg13g2_fill_2 FILLER_24_328 ();
 sg13g2_fill_2 FILLER_24_374 ();
 sg13g2_fill_2 FILLER_24_402 ();
 sg13g2_decap_4 FILLER_25_26 ();
 sg13g2_fill_1 FILLER_25_30 ();
 sg13g2_decap_8 FILLER_25_44 ();
 sg13g2_decap_8 FILLER_25_51 ();
 sg13g2_fill_2 FILLER_25_58 ();
 sg13g2_fill_1 FILLER_25_65 ();
 sg13g2_decap_8 FILLER_25_92 ();
 sg13g2_fill_2 FILLER_25_99 ();
 sg13g2_fill_1 FILLER_25_101 ();
 sg13g2_decap_4 FILLER_25_111 ();
 sg13g2_fill_2 FILLER_25_120 ();
 sg13g2_fill_2 FILLER_25_137 ();
 sg13g2_fill_1 FILLER_25_161 ();
 sg13g2_fill_1 FILLER_25_167 ();
 sg13g2_fill_2 FILLER_25_175 ();
 sg13g2_decap_8 FILLER_25_185 ();
 sg13g2_fill_2 FILLER_25_192 ();
 sg13g2_fill_1 FILLER_25_194 ();
 sg13g2_decap_8 FILLER_25_199 ();
 sg13g2_fill_2 FILLER_25_221 ();
 sg13g2_fill_1 FILLER_25_223 ();
 sg13g2_decap_8 FILLER_25_227 ();
 sg13g2_decap_8 FILLER_25_234 ();
 sg13g2_fill_1 FILLER_25_245 ();
 sg13g2_decap_4 FILLER_25_272 ();
 sg13g2_fill_2 FILLER_25_276 ();
 sg13g2_decap_4 FILLER_25_282 ();
 sg13g2_fill_2 FILLER_25_326 ();
 sg13g2_fill_1 FILLER_25_328 ();
 sg13g2_fill_2 FILLER_25_337 ();
 sg13g2_fill_2 FILLER_25_349 ();
 sg13g2_fill_1 FILLER_25_355 ();
 sg13g2_decap_8 FILLER_25_361 ();
 sg13g2_decap_8 FILLER_25_368 ();
 sg13g2_fill_2 FILLER_25_375 ();
 sg13g2_decap_8 FILLER_25_382 ();
 sg13g2_fill_2 FILLER_25_389 ();
 sg13g2_fill_2 FILLER_25_398 ();
 sg13g2_decap_8 FILLER_25_404 ();
 sg13g2_decap_8 FILLER_25_411 ();
 sg13g2_decap_8 FILLER_25_418 ();
 sg13g2_decap_4 FILLER_25_425 ();
 sg13g2_fill_1 FILLER_25_429 ();
 sg13g2_decap_8 FILLER_26_0 ();
 sg13g2_decap_8 FILLER_26_15 ();
 sg13g2_decap_8 FILLER_26_22 ();
 sg13g2_decap_8 FILLER_26_29 ();
 sg13g2_decap_8 FILLER_26_36 ();
 sg13g2_decap_4 FILLER_26_43 ();
 sg13g2_fill_2 FILLER_26_47 ();
 sg13g2_decap_8 FILLER_26_53 ();
 sg13g2_fill_1 FILLER_26_60 ();
 sg13g2_fill_2 FILLER_26_71 ();
 sg13g2_decap_4 FILLER_26_77 ();
 sg13g2_fill_1 FILLER_26_88 ();
 sg13g2_decap_8 FILLER_26_93 ();
 sg13g2_decap_8 FILLER_26_100 ();
 sg13g2_decap_4 FILLER_26_107 ();
 sg13g2_fill_2 FILLER_26_111 ();
 sg13g2_decap_4 FILLER_26_117 ();
 sg13g2_decap_4 FILLER_26_126 ();
 sg13g2_decap_4 FILLER_26_134 ();
 sg13g2_fill_2 FILLER_26_138 ();
 sg13g2_decap_8 FILLER_26_156 ();
 sg13g2_decap_4 FILLER_26_163 ();
 sg13g2_decap_4 FILLER_26_182 ();
 sg13g2_fill_1 FILLER_26_191 ();
 sg13g2_fill_1 FILLER_26_218 ();
 sg13g2_fill_2 FILLER_26_245 ();
 sg13g2_fill_1 FILLER_26_251 ();
 sg13g2_fill_2 FILLER_26_257 ();
 sg13g2_fill_2 FILLER_26_264 ();
 sg13g2_fill_1 FILLER_26_292 ();
 sg13g2_decap_8 FILLER_26_296 ();
 sg13g2_fill_2 FILLER_26_303 ();
 sg13g2_decap_4 FILLER_26_309 ();
 sg13g2_fill_2 FILLER_26_313 ();
 sg13g2_fill_1 FILLER_26_325 ();
 sg13g2_fill_1 FILLER_26_330 ();
 sg13g2_fill_1 FILLER_26_335 ();
 sg13g2_fill_1 FILLER_26_341 ();
 sg13g2_fill_2 FILLER_26_394 ();
 sg13g2_decap_8 FILLER_26_404 ();
 sg13g2_decap_8 FILLER_26_411 ();
 sg13g2_decap_8 FILLER_26_418 ();
 sg13g2_decap_4 FILLER_26_425 ();
 sg13g2_fill_1 FILLER_26_429 ();
 sg13g2_fill_2 FILLER_27_0 ();
 sg13g2_fill_1 FILLER_27_2 ();
 sg13g2_decap_4 FILLER_27_38 ();
 sg13g2_fill_1 FILLER_27_42 ();
 sg13g2_decap_4 FILLER_27_69 ();
 sg13g2_fill_2 FILLER_27_73 ();
 sg13g2_decap_4 FILLER_27_85 ();
 sg13g2_fill_1 FILLER_27_89 ();
 sg13g2_decap_8 FILLER_27_94 ();
 sg13g2_fill_1 FILLER_27_101 ();
 sg13g2_fill_1 FILLER_27_149 ();
 sg13g2_decap_8 FILLER_27_157 ();
 sg13g2_fill_2 FILLER_27_164 ();
 sg13g2_fill_1 FILLER_27_171 ();
 sg13g2_decap_8 FILLER_27_179 ();
 sg13g2_decap_8 FILLER_27_186 ();
 sg13g2_decap_8 FILLER_27_193 ();
 sg13g2_decap_4 FILLER_27_204 ();
 sg13g2_fill_2 FILLER_27_208 ();
 sg13g2_decap_8 FILLER_27_215 ();
 sg13g2_decap_8 FILLER_27_222 ();
 sg13g2_fill_2 FILLER_27_260 ();
 sg13g2_decap_8 FILLER_27_267 ();
 sg13g2_fill_1 FILLER_27_274 ();
 sg13g2_fill_1 FILLER_27_279 ();
 sg13g2_decap_8 FILLER_27_285 ();
 sg13g2_fill_2 FILLER_27_301 ();
 sg13g2_fill_1 FILLER_27_303 ();
 sg13g2_decap_4 FILLER_27_309 ();
 sg13g2_fill_1 FILLER_27_313 ();
 sg13g2_fill_2 FILLER_27_322 ();
 sg13g2_decap_4 FILLER_27_356 ();
 sg13g2_fill_2 FILLER_27_360 ();
 sg13g2_fill_1 FILLER_27_366 ();
 sg13g2_decap_8 FILLER_27_389 ();
 sg13g2_decap_4 FILLER_27_396 ();
 sg13g2_fill_2 FILLER_28_0 ();
 sg13g2_decap_8 FILLER_28_33 ();
 sg13g2_decap_8 FILLER_28_40 ();
 sg13g2_decap_8 FILLER_28_47 ();
 sg13g2_decap_8 FILLER_28_54 ();
 sg13g2_decap_8 FILLER_28_61 ();
 sg13g2_fill_2 FILLER_28_68 ();
 sg13g2_fill_1 FILLER_28_78 ();
 sg13g2_fill_1 FILLER_28_119 ();
 sg13g2_fill_2 FILLER_28_129 ();
 sg13g2_fill_1 FILLER_28_131 ();
 sg13g2_fill_2 FILLER_28_139 ();
 sg13g2_fill_1 FILLER_28_141 ();
 sg13g2_fill_1 FILLER_28_145 ();
 sg13g2_fill_2 FILLER_28_153 ();
 sg13g2_fill_1 FILLER_28_155 ();
 sg13g2_fill_2 FILLER_28_164 ();
 sg13g2_decap_8 FILLER_28_181 ();
 sg13g2_decap_8 FILLER_28_188 ();
 sg13g2_decap_8 FILLER_28_199 ();
 sg13g2_decap_8 FILLER_28_206 ();
 sg13g2_decap_8 FILLER_28_213 ();
 sg13g2_decap_4 FILLER_28_220 ();
 sg13g2_decap_4 FILLER_28_237 ();
 sg13g2_fill_1 FILLER_28_241 ();
 sg13g2_decap_8 FILLER_28_246 ();
 sg13g2_decap_4 FILLER_28_253 ();
 sg13g2_fill_1 FILLER_28_257 ();
 sg13g2_decap_8 FILLER_28_262 ();
 sg13g2_fill_2 FILLER_28_273 ();
 sg13g2_fill_1 FILLER_28_275 ();
 sg13g2_decap_8 FILLER_28_306 ();
 sg13g2_decap_4 FILLER_28_313 ();
 sg13g2_fill_1 FILLER_28_317 ();
 sg13g2_decap_8 FILLER_28_323 ();
 sg13g2_fill_2 FILLER_28_330 ();
 sg13g2_decap_8 FILLER_28_336 ();
 sg13g2_fill_2 FILLER_28_343 ();
 sg13g2_fill_1 FILLER_28_345 ();
 sg13g2_decap_4 FILLER_28_389 ();
 sg13g2_decap_8 FILLER_28_417 ();
 sg13g2_decap_4 FILLER_28_424 ();
 sg13g2_fill_2 FILLER_28_428 ();
 sg13g2_decap_8 FILLER_29_0 ();
 sg13g2_fill_1 FILLER_29_7 ();
 sg13g2_decap_8 FILLER_29_12 ();
 sg13g2_decap_4 FILLER_29_19 ();
 sg13g2_decap_4 FILLER_29_32 ();
 sg13g2_fill_1 FILLER_29_36 ();
 sg13g2_decap_8 FILLER_29_45 ();
 sg13g2_decap_8 FILLER_29_52 ();
 sg13g2_fill_2 FILLER_29_59 ();
 sg13g2_fill_1 FILLER_29_61 ();
 sg13g2_fill_2 FILLER_29_90 ();
 sg13g2_fill_2 FILLER_29_112 ();
 sg13g2_fill_1 FILLER_29_114 ();
 sg13g2_fill_1 FILLER_29_130 ();
 sg13g2_decap_8 FILLER_29_139 ();
 sg13g2_fill_2 FILLER_29_146 ();
 sg13g2_fill_2 FILLER_29_159 ();
 sg13g2_fill_1 FILLER_29_161 ();
 sg13g2_decap_8 FILLER_29_166 ();
 sg13g2_decap_8 FILLER_29_178 ();
 sg13g2_fill_2 FILLER_29_185 ();
 sg13g2_fill_1 FILLER_29_187 ();
 sg13g2_fill_2 FILLER_29_227 ();
 sg13g2_fill_1 FILLER_29_229 ();
 sg13g2_decap_8 FILLER_29_245 ();
 sg13g2_decap_8 FILLER_29_252 ();
 sg13g2_fill_1 FILLER_29_259 ();
 sg13g2_fill_1 FILLER_29_275 ();
 sg13g2_fill_2 FILLER_29_300 ();
 sg13g2_fill_1 FILLER_29_315 ();
 sg13g2_decap_4 FILLER_29_374 ();
 sg13g2_fill_1 FILLER_29_394 ();
 sg13g2_decap_8 FILLER_29_407 ();
 sg13g2_decap_8 FILLER_29_414 ();
 sg13g2_decap_8 FILLER_29_421 ();
 sg13g2_fill_2 FILLER_29_428 ();
 sg13g2_decap_8 FILLER_30_0 ();
 sg13g2_fill_2 FILLER_30_7 ();
 sg13g2_fill_1 FILLER_30_9 ();
 sg13g2_fill_2 FILLER_30_18 ();
 sg13g2_decap_4 FILLER_30_51 ();
 sg13g2_fill_2 FILLER_30_97 ();
 sg13g2_fill_2 FILLER_30_114 ();
 sg13g2_fill_2 FILLER_30_123 ();
 sg13g2_fill_1 FILLER_30_125 ();
 sg13g2_fill_2 FILLER_30_133 ();
 sg13g2_fill_1 FILLER_30_135 ();
 sg13g2_fill_2 FILLER_30_151 ();
 sg13g2_fill_1 FILLER_30_153 ();
 sg13g2_decap_4 FILLER_30_159 ();
 sg13g2_fill_1 FILLER_30_168 ();
 sg13g2_decap_4 FILLER_30_181 ();
 sg13g2_fill_1 FILLER_30_185 ();
 sg13g2_decap_8 FILLER_30_191 ();
 sg13g2_decap_4 FILLER_30_198 ();
 sg13g2_fill_1 FILLER_30_202 ();
 sg13g2_decap_8 FILLER_30_213 ();
 sg13g2_decap_4 FILLER_30_225 ();
 sg13g2_fill_1 FILLER_30_229 ();
 sg13g2_fill_1 FILLER_30_241 ();
 sg13g2_decap_4 FILLER_30_246 ();
 sg13g2_fill_1 FILLER_30_254 ();
 sg13g2_fill_1 FILLER_30_287 ();
 sg13g2_decap_4 FILLER_30_292 ();
 sg13g2_decap_8 FILLER_30_299 ();
 sg13g2_decap_8 FILLER_30_306 ();
 sg13g2_fill_1 FILLER_30_318 ();
 sg13g2_fill_1 FILLER_30_326 ();
 sg13g2_decap_8 FILLER_30_332 ();
 sg13g2_decap_8 FILLER_30_339 ();
 sg13g2_decap_4 FILLER_30_346 ();
 sg13g2_fill_1 FILLER_30_356 ();
 sg13g2_fill_1 FILLER_30_403 ();
 sg13g2_decap_8 FILLER_31_0 ();
 sg13g2_fill_2 FILLER_31_7 ();
 sg13g2_fill_2 FILLER_31_14 ();
 sg13g2_fill_1 FILLER_31_16 ();
 sg13g2_decap_4 FILLER_31_24 ();
 sg13g2_fill_1 FILLER_31_28 ();
 sg13g2_decap_8 FILLER_31_34 ();
 sg13g2_decap_4 FILLER_31_41 ();
 sg13g2_fill_2 FILLER_31_55 ();
 sg13g2_fill_1 FILLER_31_57 ();
 sg13g2_fill_1 FILLER_31_76 ();
 sg13g2_fill_2 FILLER_31_85 ();
 sg13g2_fill_1 FILLER_31_87 ();
 sg13g2_fill_2 FILLER_31_99 ();
 sg13g2_decap_4 FILLER_31_107 ();
 sg13g2_fill_2 FILLER_31_111 ();
 sg13g2_decap_8 FILLER_31_121 ();
 sg13g2_decap_4 FILLER_31_138 ();
 sg13g2_fill_1 FILLER_31_142 ();
 sg13g2_fill_1 FILLER_31_159 ();
 sg13g2_fill_2 FILLER_31_164 ();
 sg13g2_fill_1 FILLER_31_166 ();
 sg13g2_decap_8 FILLER_31_178 ();
 sg13g2_decap_8 FILLER_31_185 ();
 sg13g2_fill_2 FILLER_31_192 ();
 sg13g2_fill_1 FILLER_31_194 ();
 sg13g2_decap_4 FILLER_31_202 ();
 sg13g2_fill_1 FILLER_31_212 ();
 sg13g2_fill_2 FILLER_31_218 ();
 sg13g2_fill_2 FILLER_31_226 ();
 sg13g2_fill_2 FILLER_31_232 ();
 sg13g2_fill_1 FILLER_31_267 ();
 sg13g2_fill_1 FILLER_31_273 ();
 sg13g2_fill_1 FILLER_31_279 ();
 sg13g2_fill_2 FILLER_31_285 ();
 sg13g2_fill_1 FILLER_31_294 ();
 sg13g2_fill_1 FILLER_31_300 ();
 sg13g2_fill_1 FILLER_31_315 ();
 sg13g2_fill_2 FILLER_31_330 ();
 sg13g2_fill_2 FILLER_31_341 ();
 sg13g2_fill_1 FILLER_31_343 ();
 sg13g2_decap_4 FILLER_31_348 ();
 sg13g2_fill_1 FILLER_31_352 ();
 sg13g2_fill_2 FILLER_31_358 ();
 sg13g2_fill_1 FILLER_31_365 ();
 sg13g2_decap_8 FILLER_31_370 ();
 sg13g2_fill_2 FILLER_31_377 ();
 sg13g2_decap_8 FILLER_31_382 ();
 sg13g2_fill_1 FILLER_31_389 ();
 sg13g2_decap_8 FILLER_31_394 ();
 sg13g2_decap_8 FILLER_31_401 ();
 sg13g2_fill_2 FILLER_31_408 ();
 sg13g2_fill_1 FILLER_31_410 ();
 sg13g2_decap_8 FILLER_31_415 ();
 sg13g2_decap_8 FILLER_31_422 ();
 sg13g2_fill_1 FILLER_31_429 ();
 sg13g2_fill_2 FILLER_32_0 ();
 sg13g2_fill_1 FILLER_32_2 ();
 sg13g2_fill_2 FILLER_32_15 ();
 sg13g2_fill_1 FILLER_32_17 ();
 sg13g2_decap_4 FILLER_32_21 ();
 sg13g2_fill_1 FILLER_32_30 ();
 sg13g2_decap_4 FILLER_32_47 ();
 sg13g2_fill_1 FILLER_32_58 ();
 sg13g2_fill_1 FILLER_32_65 ();
 sg13g2_fill_1 FILLER_32_85 ();
 sg13g2_fill_2 FILLER_32_91 ();
 sg13g2_fill_2 FILLER_32_96 ();
 sg13g2_decap_4 FILLER_32_103 ();
 sg13g2_fill_1 FILLER_32_117 ();
 sg13g2_fill_1 FILLER_32_140 ();
 sg13g2_fill_1 FILLER_32_145 ();
 sg13g2_fill_2 FILLER_32_151 ();
 sg13g2_decap_4 FILLER_32_174 ();
 sg13g2_fill_1 FILLER_32_178 ();
 sg13g2_fill_2 FILLER_32_202 ();
 sg13g2_fill_1 FILLER_32_213 ();
 sg13g2_fill_2 FILLER_32_219 ();
 sg13g2_fill_2 FILLER_32_225 ();
 sg13g2_fill_1 FILLER_32_231 ();
 sg13g2_fill_2 FILLER_32_249 ();
 sg13g2_fill_1 FILLER_32_251 ();
 sg13g2_fill_2 FILLER_32_255 ();
 sg13g2_fill_1 FILLER_32_257 ();
 sg13g2_fill_2 FILLER_32_266 ();
 sg13g2_decap_4 FILLER_32_293 ();
 sg13g2_fill_2 FILLER_32_297 ();
 sg13g2_decap_8 FILLER_32_312 ();
 sg13g2_fill_2 FILLER_32_319 ();
 sg13g2_fill_1 FILLER_32_321 ();
 sg13g2_decap_4 FILLER_32_348 ();
 sg13g2_decap_8 FILLER_32_356 ();
 sg13g2_decap_8 FILLER_32_363 ();
 sg13g2_fill_1 FILLER_32_403 ();
 sg13g2_decap_4 FILLER_33_0 ();
 sg13g2_fill_1 FILLER_33_4 ();
 sg13g2_fill_1 FILLER_33_20 ();
 sg13g2_decap_8 FILLER_33_39 ();
 sg13g2_decap_8 FILLER_33_46 ();
 sg13g2_decap_8 FILLER_33_53 ();
 sg13g2_fill_2 FILLER_33_60 ();
 sg13g2_fill_1 FILLER_33_77 ();
 sg13g2_fill_1 FILLER_33_104 ();
 sg13g2_fill_1 FILLER_33_109 ();
 sg13g2_decap_4 FILLER_33_130 ();
 sg13g2_fill_2 FILLER_33_149 ();
 sg13g2_fill_1 FILLER_33_156 ();
 sg13g2_decap_8 FILLER_33_161 ();
 sg13g2_decap_8 FILLER_33_168 ();
 sg13g2_decap_8 FILLER_33_175 ();
 sg13g2_decap_8 FILLER_33_182 ();
 sg13g2_fill_1 FILLER_33_189 ();
 sg13g2_fill_1 FILLER_33_203 ();
 sg13g2_fill_1 FILLER_33_216 ();
 sg13g2_fill_2 FILLER_33_232 ();
 sg13g2_fill_1 FILLER_33_238 ();
 sg13g2_fill_1 FILLER_33_255 ();
 sg13g2_decap_8 FILLER_33_272 ();
 sg13g2_decap_4 FILLER_33_279 ();
 sg13g2_fill_2 FILLER_33_283 ();
 sg13g2_decap_4 FILLER_33_314 ();
 sg13g2_fill_1 FILLER_33_318 ();
 sg13g2_decap_4 FILLER_33_324 ();
 sg13g2_fill_1 FILLER_33_328 ();
 sg13g2_decap_4 FILLER_33_333 ();
 sg13g2_fill_2 FILLER_33_337 ();
 sg13g2_fill_1 FILLER_33_380 ();
 sg13g2_fill_2 FILLER_33_391 ();
 sg13g2_fill_2 FILLER_33_401 ();
 sg13g2_fill_1 FILLER_33_403 ();
 sg13g2_fill_1 FILLER_33_409 ();
 sg13g2_fill_2 FILLER_33_415 ();
 sg13g2_fill_1 FILLER_33_417 ();
 sg13g2_decap_8 FILLER_33_422 ();
 sg13g2_fill_1 FILLER_33_429 ();
 sg13g2_decap_4 FILLER_34_0 ();
 sg13g2_fill_1 FILLER_34_4 ();
 sg13g2_fill_2 FILLER_34_10 ();
 sg13g2_fill_1 FILLER_34_15 ();
 sg13g2_decap_8 FILLER_34_21 ();
 sg13g2_decap_8 FILLER_34_28 ();
 sg13g2_fill_1 FILLER_34_35 ();
 sg13g2_decap_8 FILLER_34_44 ();
 sg13g2_decap_4 FILLER_34_51 ();
 sg13g2_fill_2 FILLER_34_77 ();
 sg13g2_fill_2 FILLER_34_86 ();
 sg13g2_fill_1 FILLER_34_96 ();
 sg13g2_fill_1 FILLER_34_117 ();
 sg13g2_fill_1 FILLER_34_122 ();
 sg13g2_fill_1 FILLER_34_129 ();
 sg13g2_decap_4 FILLER_34_135 ();
 sg13g2_fill_2 FILLER_34_155 ();
 sg13g2_fill_1 FILLER_34_157 ();
 sg13g2_fill_2 FILLER_34_162 ();
 sg13g2_fill_1 FILLER_34_164 ();
 sg13g2_decap_8 FILLER_34_179 ();
 sg13g2_decap_8 FILLER_34_195 ();
 sg13g2_decap_8 FILLER_34_202 ();
 sg13g2_decap_4 FILLER_34_213 ();
 sg13g2_decap_8 FILLER_34_221 ();
 sg13g2_fill_1 FILLER_34_238 ();
 sg13g2_fill_2 FILLER_34_244 ();
 sg13g2_fill_2 FILLER_34_254 ();
 sg13g2_fill_1 FILLER_34_256 ();
 sg13g2_decap_8 FILLER_34_261 ();
 sg13g2_fill_2 FILLER_34_268 ();
 sg13g2_decap_4 FILLER_34_274 ();
 sg13g2_fill_2 FILLER_34_291 ();
 sg13g2_fill_2 FILLER_34_307 ();
 sg13g2_decap_8 FILLER_34_355 ();
 sg13g2_decap_8 FILLER_34_388 ();
 sg13g2_fill_2 FILLER_34_395 ();
 sg13g2_fill_1 FILLER_34_406 ();
 sg13g2_decap_8 FILLER_34_418 ();
 sg13g2_decap_4 FILLER_34_425 ();
 sg13g2_fill_1 FILLER_34_429 ();
 sg13g2_decap_8 FILLER_35_0 ();
 sg13g2_fill_1 FILLER_35_16 ();
 sg13g2_decap_8 FILLER_35_46 ();
 sg13g2_decap_8 FILLER_35_53 ();
 sg13g2_decap_8 FILLER_35_60 ();
 sg13g2_fill_2 FILLER_35_67 ();
 sg13g2_fill_1 FILLER_35_69 ();
 sg13g2_fill_1 FILLER_35_95 ();
 sg13g2_fill_2 FILLER_35_101 ();
 sg13g2_fill_1 FILLER_35_103 ();
 sg13g2_fill_1 FILLER_35_112 ();
 sg13g2_fill_1 FILLER_35_118 ();
 sg13g2_decap_8 FILLER_35_140 ();
 sg13g2_decap_4 FILLER_35_153 ();
 sg13g2_fill_2 FILLER_35_157 ();
 sg13g2_decap_8 FILLER_35_163 ();
 sg13g2_fill_1 FILLER_35_170 ();
 sg13g2_decap_8 FILLER_35_197 ();
 sg13g2_decap_8 FILLER_35_204 ();
 sg13g2_decap_8 FILLER_35_211 ();
 sg13g2_fill_1 FILLER_35_218 ();
 sg13g2_fill_1 FILLER_35_224 ();
 sg13g2_fill_1 FILLER_35_235 ();
 sg13g2_fill_1 FILLER_35_244 ();
 sg13g2_fill_1 FILLER_35_249 ();
 sg13g2_decap_8 FILLER_35_276 ();
 sg13g2_decap_8 FILLER_35_283 ();
 sg13g2_decap_4 FILLER_35_290 ();
 sg13g2_fill_2 FILLER_35_294 ();
 sg13g2_decap_8 FILLER_35_309 ();
 sg13g2_decap_4 FILLER_35_316 ();
 sg13g2_decap_8 FILLER_35_324 ();
 sg13g2_decap_4 FILLER_35_331 ();
 sg13g2_fill_1 FILLER_35_335 ();
 sg13g2_decap_8 FILLER_35_340 ();
 sg13g2_decap_8 FILLER_35_347 ();
 sg13g2_fill_1 FILLER_35_354 ();
 sg13g2_decap_4 FILLER_35_364 ();
 sg13g2_fill_2 FILLER_35_372 ();
 sg13g2_fill_1 FILLER_35_374 ();
 sg13g2_decap_8 FILLER_35_386 ();
 sg13g2_fill_2 FILLER_35_393 ();
 sg13g2_fill_1 FILLER_35_395 ();
 sg13g2_decap_4 FILLER_36_0 ();
 sg13g2_fill_1 FILLER_36_4 ();
 sg13g2_fill_2 FILLER_36_13 ();
 sg13g2_fill_2 FILLER_36_26 ();
 sg13g2_fill_1 FILLER_36_28 ();
 sg13g2_decap_8 FILLER_36_33 ();
 sg13g2_decap_8 FILLER_36_45 ();
 sg13g2_decap_8 FILLER_36_52 ();
 sg13g2_decap_8 FILLER_36_59 ();
 sg13g2_fill_2 FILLER_36_66 ();
 sg13g2_decap_8 FILLER_36_81 ();
 sg13g2_fill_1 FILLER_36_107 ();
 sg13g2_fill_1 FILLER_36_112 ();
 sg13g2_fill_1 FILLER_36_118 ();
 sg13g2_decap_8 FILLER_36_128 ();
 sg13g2_decap_4 FILLER_36_135 ();
 sg13g2_decap_4 FILLER_36_143 ();
 sg13g2_fill_1 FILLER_36_151 ();
 sg13g2_decap_8 FILLER_36_186 ();
 sg13g2_decap_8 FILLER_36_193 ();
 sg13g2_decap_8 FILLER_36_200 ();
 sg13g2_decap_8 FILLER_36_207 ();
 sg13g2_decap_8 FILLER_36_214 ();
 sg13g2_decap_8 FILLER_36_221 ();
 sg13g2_fill_1 FILLER_36_228 ();
 sg13g2_decap_4 FILLER_36_239 ();
 sg13g2_fill_2 FILLER_36_243 ();
 sg13g2_decap_8 FILLER_36_258 ();
 sg13g2_fill_1 FILLER_36_265 ();
 sg13g2_decap_4 FILLER_36_282 ();
 sg13g2_decap_4 FILLER_36_299 ();
 sg13g2_fill_2 FILLER_36_303 ();
 sg13g2_decap_8 FILLER_36_340 ();
 sg13g2_fill_2 FILLER_36_347 ();
 sg13g2_fill_2 FILLER_36_362 ();
 sg13g2_decap_8 FILLER_36_378 ();
 sg13g2_decap_8 FILLER_36_385 ();
 sg13g2_fill_2 FILLER_36_392 ();
 sg13g2_fill_1 FILLER_36_394 ();
 sg13g2_fill_2 FILLER_36_402 ();
 sg13g2_fill_2 FILLER_36_409 ();
 sg13g2_decap_8 FILLER_36_415 ();
 sg13g2_decap_8 FILLER_36_422 ();
 sg13g2_fill_1 FILLER_36_429 ();
 sg13g2_decap_4 FILLER_37_52 ();
 sg13g2_fill_2 FILLER_37_56 ();
 sg13g2_decap_4 FILLER_37_84 ();
 sg13g2_fill_2 FILLER_37_88 ();
 sg13g2_decap_8 FILLER_37_94 ();
 sg13g2_fill_2 FILLER_37_101 ();
 sg13g2_fill_1 FILLER_37_103 ();
 sg13g2_decap_8 FILLER_37_138 ();
 sg13g2_decap_4 FILLER_37_145 ();
 sg13g2_decap_8 FILLER_37_153 ();
 sg13g2_decap_4 FILLER_37_160 ();
 sg13g2_fill_1 FILLER_37_164 ();
 sg13g2_decap_8 FILLER_37_169 ();
 sg13g2_fill_2 FILLER_37_176 ();
 sg13g2_fill_1 FILLER_37_234 ();
 sg13g2_fill_2 FILLER_37_261 ();
 sg13g2_decap_4 FILLER_37_293 ();
 sg13g2_fill_1 FILLER_37_297 ();
 sg13g2_decap_8 FILLER_37_302 ();
 sg13g2_fill_1 FILLER_37_309 ();
 sg13g2_decap_8 FILLER_37_318 ();
 sg13g2_decap_4 FILLER_37_325 ();
 sg13g2_decap_8 FILLER_37_333 ();
 sg13g2_decap_8 FILLER_37_340 ();
 sg13g2_fill_2 FILLER_37_347 ();
 sg13g2_fill_1 FILLER_37_375 ();
 sg13g2_fill_2 FILLER_37_402 ();
 sg13g2_decap_4 FILLER_38_0 ();
 sg13g2_fill_2 FILLER_38_4 ();
 sg13g2_decap_4 FILLER_38_10 ();
 sg13g2_fill_1 FILLER_38_14 ();
 sg13g2_decap_4 FILLER_38_20 ();
 sg13g2_fill_2 FILLER_38_33 ();
 sg13g2_fill_1 FILLER_38_35 ();
 sg13g2_decap_8 FILLER_38_40 ();
 sg13g2_decap_8 FILLER_38_47 ();
 sg13g2_decap_8 FILLER_38_54 ();
 sg13g2_decap_4 FILLER_38_61 ();
 sg13g2_fill_1 FILLER_38_65 ();
 sg13g2_decap_4 FILLER_38_70 ();
 sg13g2_fill_1 FILLER_38_106 ();
 sg13g2_decap_4 FILLER_38_111 ();
 sg13g2_fill_1 FILLER_38_115 ();
 sg13g2_fill_1 FILLER_38_124 ();
 sg13g2_fill_2 FILLER_38_141 ();
 sg13g2_fill_1 FILLER_38_175 ();
 sg13g2_fill_1 FILLER_38_180 ();
 sg13g2_fill_1 FILLER_38_185 ();
 sg13g2_fill_2 FILLER_38_190 ();
 sg13g2_fill_1 FILLER_38_236 ();
 sg13g2_fill_2 FILLER_38_241 ();
 sg13g2_decap_8 FILLER_38_247 ();
 sg13g2_decap_4 FILLER_38_254 ();
 sg13g2_fill_2 FILLER_38_258 ();
 sg13g2_decap_8 FILLER_38_276 ();
 sg13g2_decap_4 FILLER_38_283 ();
 sg13g2_fill_1 FILLER_38_317 ();
 sg13g2_decap_8 FILLER_38_348 ();
 sg13g2_fill_2 FILLER_38_363 ();
 sg13g2_fill_1 FILLER_38_365 ();
 sg13g2_fill_2 FILLER_38_371 ();
 sg13g2_fill_1 FILLER_38_373 ();
 sg13g2_decap_4 FILLER_38_379 ();
 sg13g2_fill_2 FILLER_38_383 ();
 sg13g2_fill_2 FILLER_38_393 ();
 sg13g2_fill_1 FILLER_38_395 ();
 sg13g2_fill_1 FILLER_38_409 ();
 sg13g2_decap_8 FILLER_38_414 ();
 sg13g2_decap_8 FILLER_38_421 ();
 sg13g2_fill_2 FILLER_38_428 ();
endmodule
