module tt_um_htfab_caterpillar (clk,
    ena,
    rst_n,
    ui_in,
    uio_in,
    uio_oe,
    uio_out,
    uo_out);
 input clk;
 input ena;
 input rst_n;
 input [7:0] ui_in;
 input [7:0] uio_in;
 output [7:0] uio_oe;
 output [7:0] uio_out;
 output [7:0] uo_out;

 wire _0000_;
 wire _0001_;
 wire _0002_;
 wire _0003_;
 wire _0004_;
 wire _0005_;
 wire _0006_;
 wire _0007_;
 wire _0008_;
 wire _0009_;
 wire _0010_;
 wire _0011_;
 wire _0012_;
 wire _0013_;
 wire _0014_;
 wire _0015_;
 wire _0016_;
 wire _0017_;
 wire _0018_;
 wire _0019_;
 wire _0020_;
 wire _0021_;
 wire _0022_;
 wire _0023_;
 wire _0024_;
 wire _0025_;
 wire _0026_;
 wire _0027_;
 wire _0028_;
 wire _0029_;
 wire _0030_;
 wire _0031_;
 wire _0032_;
 wire _0033_;
 wire _0034_;
 wire _0035_;
 wire _0036_;
 wire _0037_;
 wire _0038_;
 wire _0039_;
 wire _0040_;
 wire _0041_;
 wire _0042_;
 wire _0043_;
 wire _0044_;
 wire _0045_;
 wire _0046_;
 wire _0047_;
 wire _0048_;
 wire _0049_;
 wire _0050_;
 wire _0051_;
 wire _0052_;
 wire _0053_;
 wire _0054_;
 wire _0055_;
 wire _0056_;
 wire _0057_;
 wire _0058_;
 wire _0059_;
 wire _0060_;
 wire _0061_;
 wire _0062_;
 wire _0063_;
 wire _0064_;
 wire _0065_;
 wire _0066_;
 wire _0067_;
 wire _0068_;
 wire _0069_;
 wire _0070_;
 wire _0071_;
 wire _0072_;
 wire _0073_;
 wire _0074_;
 wire _0075_;
 wire _0076_;
 wire _0077_;
 wire _0078_;
 wire _0079_;
 wire _0080_;
 wire _0081_;
 wire _0082_;
 wire _0083_;
 wire _0084_;
 wire _0085_;
 wire _0086_;
 wire _0087_;
 wire _0088_;
 wire _0089_;
 wire _0090_;
 wire _0091_;
 wire _0092_;
 wire _0093_;
 wire _0094_;
 wire _0095_;
 wire _0096_;
 wire _0097_;
 wire _0098_;
 wire _0099_;
 wire _0100_;
 wire _0101_;
 wire _0102_;
 wire _0103_;
 wire _0104_;
 wire _0105_;
 wire _0106_;
 wire _0107_;
 wire _0108_;
 wire _0109_;
 wire _0110_;
 wire _0111_;
 wire _0112_;
 wire _0113_;
 wire _0114_;
 wire _0115_;
 wire _0116_;
 wire _0117_;
 wire _0118_;
 wire _0119_;
 wire _0120_;
 wire _0121_;
 wire _0122_;
 wire _0123_;
 wire _0124_;
 wire _0125_;
 wire _0126_;
 wire _0127_;
 wire _0128_;
 wire _0129_;
 wire _0130_;
 wire _0131_;
 wire _0132_;
 wire _0133_;
 wire _0134_;
 wire _0135_;
 wire _0136_;
 wire _0137_;
 wire _0138_;
 wire _0139_;
 wire _0140_;
 wire _0141_;
 wire _0142_;
 wire _0143_;
 wire _0144_;
 wire _0145_;
 wire _0146_;
 wire _0147_;
 wire _0148_;
 wire _0149_;
 wire _0150_;
 wire _0151_;
 wire _0152_;
 wire _0153_;
 wire _0154_;
 wire _0155_;
 wire _0156_;
 wire _0157_;
 wire _0158_;
 wire _0159_;
 wire _0160_;
 wire _0161_;
 wire _0162_;
 wire _0163_;
 wire _0164_;
 wire _0165_;
 wire _0166_;
 wire _0167_;
 wire _0168_;
 wire _0169_;
 wire _0170_;
 wire _0171_;
 wire _0172_;
 wire _0173_;
 wire _0174_;
 wire _0175_;
 wire _0176_;
 wire _0177_;
 wire _0178_;
 wire _0179_;
 wire _0180_;
 wire _0181_;
 wire _0182_;
 wire _0183_;
 wire _0184_;
 wire _0185_;
 wire _0186_;
 wire _0187_;
 wire _0188_;
 wire _0189_;
 wire _0190_;
 wire _0191_;
 wire _0192_;
 wire _0193_;
 wire _0194_;
 wire _0195_;
 wire _0196_;
 wire _0197_;
 wire _0198_;
 wire _0199_;
 wire _0200_;
 wire _0201_;
 wire _0202_;
 wire _0203_;
 wire _0204_;
 wire _0205_;
 wire _0206_;
 wire _0207_;
 wire _0208_;
 wire _0209_;
 wire _0210_;
 wire _0211_;
 wire _0212_;
 wire _0213_;
 wire _0214_;
 wire _0215_;
 wire _0216_;
 wire _0217_;
 wire _0218_;
 wire _0219_;
 wire _0220_;
 wire _0221_;
 wire _0222_;
 wire _0223_;
 wire _0224_;
 wire _0225_;
 wire _0226_;
 wire _0227_;
 wire _0228_;
 wire _0229_;
 wire _0230_;
 wire _0231_;
 wire _0232_;
 wire _0233_;
 wire _0234_;
 wire _0235_;
 wire _0236_;
 wire _0237_;
 wire _0238_;
 wire _0239_;
 wire _0240_;
 wire _0241_;
 wire _0242_;
 wire _0243_;
 wire _0244_;
 wire _0245_;
 wire _0246_;
 wire _0247_;
 wire _0248_;
 wire _0249_;
 wire _0250_;
 wire _0251_;
 wire _0252_;
 wire _0253_;
 wire _0254_;
 wire _0255_;
 wire _0256_;
 wire _0257_;
 wire _0258_;
 wire _0259_;
 wire _0260_;
 wire _0261_;
 wire _0262_;
 wire _0263_;
 wire _0264_;
 wire _0265_;
 wire _0266_;
 wire _0267_;
 wire _0268_;
 wire _0269_;
 wire _0270_;
 wire _0271_;
 wire _0272_;
 wire _0273_;
 wire _0274_;
 wire _0275_;
 wire _0276_;
 wire _0277_;
 wire _0278_;
 wire _0279_;
 wire _0280_;
 wire _0281_;
 wire _0282_;
 wire _0283_;
 wire _0284_;
 wire _0285_;
 wire _0286_;
 wire _0287_;
 wire _0288_;
 wire _0289_;
 wire _0290_;
 wire _0291_;
 wire _0292_;
 wire _0293_;
 wire _0294_;
 wire _0295_;
 wire _0296_;
 wire _0297_;
 wire _0298_;
 wire _0299_;
 wire _0300_;
 wire _0301_;
 wire _0302_;
 wire _0303_;
 wire _0304_;
 wire _0305_;
 wire _0306_;
 wire _0307_;
 wire _0308_;
 wire _0309_;
 wire _0310_;
 wire _0311_;
 wire _0312_;
 wire _0313_;
 wire _0314_;
 wire _0315_;
 wire _0316_;
 wire _0317_;
 wire _0318_;
 wire _0319_;
 wire _0320_;
 wire _0321_;
 wire _0322_;
 wire _0323_;
 wire _0324_;
 wire _0325_;
 wire _0326_;
 wire _0327_;
 wire _0328_;
 wire _0329_;
 wire _0330_;
 wire _0331_;
 wire _0332_;
 wire _0333_;
 wire _0334_;
 wire _0335_;
 wire _0336_;
 wire _0337_;
 wire _0338_;
 wire _0339_;
 wire _0340_;
 wire _0341_;
 wire _0342_;
 wire _0343_;
 wire _0344_;
 wire _0345_;
 wire _0346_;
 wire _0347_;
 wire _0348_;
 wire _0349_;
 wire _0350_;
 wire _0351_;
 wire _0352_;
 wire _0353_;
 wire _0354_;
 wire _0355_;
 wire _0356_;
 wire _0357_;
 wire _0358_;
 wire _0359_;
 wire _0360_;
 wire _0361_;
 wire _0362_;
 wire _0363_;
 wire _0364_;
 wire _0365_;
 wire _0366_;
 wire _0367_;
 wire _0368_;
 wire _0369_;
 wire _0370_;
 wire _0371_;
 wire _0372_;
 wire _0373_;
 wire _0374_;
 wire _0375_;
 wire _0376_;
 wire _0377_;
 wire _0378_;
 wire _0379_;
 wire _0380_;
 wire _0381_;
 wire _0382_;
 wire _0383_;
 wire _0384_;
 wire _0385_;
 wire _0386_;
 wire _0387_;
 wire _0388_;
 wire _0389_;
 wire _0390_;
 wire _0391_;
 wire _0392_;
 wire _0393_;
 wire _0394_;
 wire _0395_;
 wire _0396_;
 wire _0397_;
 wire _0398_;
 wire _0399_;
 wire _0400_;
 wire _0401_;
 wire _0402_;
 wire _0403_;
 wire _0404_;
 wire _0405_;
 wire _0406_;
 wire _0407_;
 wire _0408_;
 wire _0409_;
 wire _0410_;
 wire _0411_;
 wire _0412_;
 wire _0413_;
 wire _0414_;
 wire _0415_;
 wire _0416_;
 wire _0417_;
 wire _0418_;
 wire _0419_;
 wire _0420_;
 wire _0421_;
 wire _0422_;
 wire _0423_;
 wire _0424_;
 wire _0425_;
 wire _0426_;
 wire _0427_;
 wire _0428_;
 wire _0429_;
 wire _0430_;
 wire _0431_;
 wire _0432_;
 wire _0433_;
 wire _0434_;
 wire _0435_;
 wire _0436_;
 wire _0437_;
 wire _0438_;
 wire _0439_;
 wire _0440_;
 wire _0441_;
 wire _0442_;
 wire _0443_;
 wire _0444_;
 wire _0445_;
 wire _0446_;
 wire _0447_;
 wire _0448_;
 wire _0449_;
 wire _0450_;
 wire _0451_;
 wire _0452_;
 wire _0453_;
 wire _0454_;
 wire _0455_;
 wire _0456_;
 wire _0457_;
 wire _0458_;
 wire _0459_;
 wire _0460_;
 wire _0461_;
 wire _0462_;
 wire _0463_;
 wire _0464_;
 wire _0465_;
 wire _0466_;
 wire _0467_;
 wire _0468_;
 wire _0469_;
 wire _0470_;
 wire _0471_;
 wire _0472_;
 wire _0473_;
 wire _0474_;
 wire _0475_;
 wire _0476_;
 wire _0477_;
 wire _0478_;
 wire _0479_;
 wire _0480_;
 wire _0481_;
 wire _0482_;
 wire _0483_;
 wire _0484_;
 wire _0485_;
 wire _0486_;
 wire _0487_;
 wire _0488_;
 wire _0489_;
 wire _0490_;
 wire _0491_;
 wire _0492_;
 wire _0493_;
 wire _0494_;
 wire _0495_;
 wire _0496_;
 wire _0497_;
 wire _0498_;
 wire _0499_;
 wire _0500_;
 wire _0501_;
 wire _0502_;
 wire _0503_;
 wire _0504_;
 wire _0505_;
 wire _0506_;
 wire _0507_;
 wire _0508_;
 wire _0509_;
 wire _0510_;
 wire _0511_;
 wire _0512_;
 wire _0513_;
 wire _0514_;
 wire _0515_;
 wire _0516_;
 wire _0517_;
 wire _0518_;
 wire _0519_;
 wire _0520_;
 wire _0521_;
 wire _0522_;
 wire _0523_;
 wire _0524_;
 wire _0525_;
 wire _0526_;
 wire _0527_;
 wire _0528_;
 wire _0529_;
 wire _0530_;
 wire _0531_;
 wire _0532_;
 wire _0533_;
 wire _0534_;
 wire _0535_;
 wire _0536_;
 wire _0537_;
 wire _0538_;
 wire _0539_;
 wire _0540_;
 wire _0541_;
 wire _0542_;
 wire _0543_;
 wire _0544_;
 wire _0545_;
 wire _0546_;
 wire _0547_;
 wire _0548_;
 wire _0549_;
 wire _0550_;
 wire _0551_;
 wire _0552_;
 wire _0553_;
 wire _0554_;
 wire _0555_;
 wire _0556_;
 wire _0557_;
 wire _0558_;
 wire _0559_;
 wire _0560_;
 wire _0561_;
 wire _0562_;
 wire _0563_;
 wire _0564_;
 wire _0565_;
 wire _0566_;
 wire _0567_;
 wire _0568_;
 wire _0569_;
 wire _0570_;
 wire _0571_;
 wire _0572_;
 wire _0573_;
 wire _0574_;
 wire _0575_;
 wire _0576_;
 wire _0577_;
 wire _0578_;
 wire _0579_;
 wire _0580_;
 wire _0581_;
 wire _0582_;
 wire _0583_;
 wire _0584_;
 wire _0585_;
 wire _0586_;
 wire _0587_;
 wire _0588_;
 wire _0589_;
 wire _0590_;
 wire _0591_;
 wire _0592_;
 wire _0593_;
 wire _0594_;
 wire _0595_;
 wire _0596_;
 wire _0597_;
 wire _0598_;
 wire _0599_;
 wire _0600_;
 wire _0601_;
 wire _0602_;
 wire _0603_;
 wire _0604_;
 wire _0605_;
 wire _0606_;
 wire _0607_;
 wire _0608_;
 wire _0609_;
 wire _0610_;
 wire _0611_;
 wire _0612_;
 wire _0613_;
 wire _0614_;
 wire _0615_;
 wire _0616_;
 wire _0617_;
 wire _0618_;
 wire _0619_;
 wire _0620_;
 wire _0621_;
 wire _0622_;
 wire _0623_;
 wire _0624_;
 wire _0625_;
 wire _0626_;
 wire _0627_;
 wire _0628_;
 wire _0629_;
 wire _0630_;
 wire _0631_;
 wire _0632_;
 wire _0633_;
 wire _0634_;
 wire _0635_;
 wire _0636_;
 wire _0637_;
 wire _0638_;
 wire _0639_;
 wire _0640_;
 wire _0641_;
 wire _0642_;
 wire _0643_;
 wire _0644_;
 wire _0645_;
 wire _0646_;
 wire _0647_;
 wire _0648_;
 wire _0649_;
 wire _0650_;
 wire _0651_;
 wire _0652_;
 wire _0653_;
 wire _0654_;
 wire _0655_;
 wire _0656_;
 wire _0657_;
 wire _0658_;
 wire _0659_;
 wire _0660_;
 wire _0661_;
 wire _0662_;
 wire _0663_;
 wire _0664_;
 wire _0665_;
 wire _0666_;
 wire _0667_;
 wire _0668_;
 wire _0669_;
 wire _0670_;
 wire _0671_;
 wire _0672_;
 wire _0673_;
 wire _0674_;
 wire _0675_;
 wire _0676_;
 wire _0677_;
 wire _0678_;
 wire _0679_;
 wire _0680_;
 wire _0681_;
 wire _0682_;
 wire _0683_;
 wire _0684_;
 wire _0685_;
 wire _0686_;
 wire _0687_;
 wire _0688_;
 wire _0689_;
 wire _0690_;
 wire _0691_;
 wire _0692_;
 wire _0693_;
 wire _0694_;
 wire _0695_;
 wire _0696_;
 wire _0697_;
 wire _0698_;
 wire _0699_;
 wire _0700_;
 wire _0701_;
 wire _0702_;
 wire _0703_;
 wire _0704_;
 wire _0705_;
 wire _0706_;
 wire _0707_;
 wire _0708_;
 wire _0709_;
 wire _0710_;
 wire _0711_;
 wire _0712_;
 wire _0713_;
 wire _0714_;
 wire _0715_;
 wire _0716_;
 wire _0717_;
 wire _0718_;
 wire _0719_;
 wire _0720_;
 wire _0721_;
 wire _0722_;
 wire _0723_;
 wire _0724_;
 wire _0725_;
 wire _0726_;
 wire _0727_;
 wire _0728_;
 wire _0729_;
 wire _0730_;
 wire _0731_;
 wire _0732_;
 wire _0733_;
 wire _0734_;
 wire _0735_;
 wire _0736_;
 wire _0737_;
 wire _0738_;
 wire _0739_;
 wire _0740_;
 wire _0741_;
 wire _0742_;
 wire _0743_;
 wire _0744_;
 wire _0745_;
 wire _0746_;
 wire _0747_;
 wire _0748_;
 wire _0749_;
 wire _0750_;
 wire _0751_;
 wire _0752_;
 wire _0753_;
 wire _0754_;
 wire _0755_;
 wire _0756_;
 wire _0757_;
 wire _0758_;
 wire _0759_;
 wire _0760_;
 wire _0761_;
 wire _0762_;
 wire _0763_;
 wire _0764_;
 wire _0765_;
 wire _0766_;
 wire _0767_;
 wire _0768_;
 wire _0769_;
 wire _0770_;
 wire _0771_;
 wire _0772_;
 wire _0773_;
 wire _0774_;
 wire _0775_;
 wire _0776_;
 wire _0777_;
 wire _0778_;
 wire _0779_;
 wire _0780_;
 wire _0781_;
 wire _0782_;
 wire _0783_;
 wire _0784_;
 wire _0785_;
 wire _0786_;
 wire _0787_;
 wire _0788_;
 wire _0789_;
 wire _0790_;
 wire _0791_;
 wire _0792_;
 wire _0793_;
 wire _0794_;
 wire _0795_;
 wire _0796_;
 wire _0797_;
 wire _0798_;
 wire _0799_;
 wire _0800_;
 wire _0801_;
 wire _0802_;
 wire _0803_;
 wire _0804_;
 wire _0805_;
 wire _0806_;
 wire _0807_;
 wire _0808_;
 wire _0809_;
 wire _0810_;
 wire _0811_;
 wire _0812_;
 wire _0813_;
 wire _0814_;
 wire _0815_;
 wire _0816_;
 wire _0817_;
 wire _0818_;
 wire _0819_;
 wire _0820_;
 wire _0821_;
 wire _0822_;
 wire _0823_;
 wire _0824_;
 wire _0825_;
 wire _0826_;
 wire _0827_;
 wire _0828_;
 wire _0829_;
 wire _0830_;
 wire _0831_;
 wire _0832_;
 wire _0833_;
 wire _0834_;
 wire _0835_;
 wire _0836_;
 wire _0837_;
 wire _0838_;
 wire _0839_;
 wire _0840_;
 wire _0841_;
 wire _0842_;
 wire _0843_;
 wire _0844_;
 wire _0845_;
 wire _0846_;
 wire _0847_;
 wire _0848_;
 wire _0849_;
 wire _0850_;
 wire _0851_;
 wire _0852_;
 wire _0853_;
 wire _0854_;
 wire _0855_;
 wire _0856_;
 wire _0857_;
 wire _0858_;
 wire _0859_;
 wire _0860_;
 wire _0861_;
 wire _0862_;
 wire _0863_;
 wire _0864_;
 wire _0865_;
 wire _0866_;
 wire _0867_;
 wire _0868_;
 wire _0869_;
 wire _0870_;
 wire _0871_;
 wire _0872_;
 wire _0873_;
 wire _0874_;
 wire _0875_;
 wire _0876_;
 wire _0877_;
 wire _0878_;
 wire _0879_;
 wire _0880_;
 wire _0881_;
 wire _0882_;
 wire _0883_;
 wire _0884_;
 wire _0885_;
 wire _0886_;
 wire _0887_;
 wire _0888_;
 wire _0889_;
 wire _0890_;
 wire _0891_;
 wire _0892_;
 wire _0893_;
 wire _0894_;
 wire _0895_;
 wire _0896_;
 wire _0897_;
 wire _0898_;
 wire _0899_;
 wire _0900_;
 wire _0901_;
 wire _0902_;
 wire _0903_;
 wire _0904_;
 wire _0905_;
 wire _0906_;
 wire _0907_;
 wire _0908_;
 wire _0909_;
 wire _0910_;
 wire _0911_;
 wire _0912_;
 wire _0913_;
 wire _0914_;
 wire _0915_;
 wire _0916_;
 wire _0917_;
 wire _0918_;
 wire _0919_;
 wire _0920_;
 wire _0921_;
 wire _0922_;
 wire _0923_;
 wire _0924_;
 wire _0925_;
 wire _0926_;
 wire _0927_;
 wire _0928_;
 wire _0929_;
 wire _0930_;
 wire _0931_;
 wire _0932_;
 wire _0933_;
 wire _0934_;
 wire _0935_;
 wire _0936_;
 wire _0937_;
 wire _0938_;
 wire _0939_;
 wire _0940_;
 wire _0941_;
 wire _0942_;
 wire _0943_;
 wire _0944_;
 wire _0945_;
 wire _0946_;
 wire _0947_;
 wire _0948_;
 wire _0949_;
 wire _0950_;
 wire _0951_;
 wire _0952_;
 wire _0953_;
 wire _0954_;
 wire _0955_;
 wire _0956_;
 wire _0957_;
 wire _0958_;
 wire _0959_;
 wire _0960_;
 wire _0961_;
 wire _0962_;
 wire _0963_;
 wire _0964_;
 wire _0965_;
 wire _0966_;
 wire _0967_;
 wire _0968_;
 wire _0969_;
 wire _0970_;
 wire _0971_;
 wire _0972_;
 wire _0973_;
 wire _0974_;
 wire _0975_;
 wire _0976_;
 wire _0977_;
 wire _0978_;
 wire _0979_;
 wire _0980_;
 wire _0981_;
 wire _0982_;
 wire _0983_;
 wire _0984_;
 wire _0985_;
 wire _0986_;
 wire _0987_;
 wire _0988_;
 wire _0989_;
 wire _0990_;
 wire _0991_;
 wire _0992_;
 wire _0993_;
 wire _0994_;
 wire _0995_;
 wire _0996_;
 wire _0997_;
 wire _0998_;
 wire _0999_;
 wire _1000_;
 wire _1001_;
 wire _1002_;
 wire _1003_;
 wire _1004_;
 wire _1005_;
 wire _1006_;
 wire _1007_;
 wire _1008_;
 wire _1009_;
 wire _1010_;
 wire _1011_;
 wire _1012_;
 wire _1013_;
 wire _1014_;
 wire _1015_;
 wire _1016_;
 wire _1017_;
 wire _1018_;
 wire _1019_;
 wire _1020_;
 wire _1021_;
 wire _1022_;
 wire _1023_;
 wire _1024_;
 wire _1025_;
 wire _1026_;
 wire _1027_;
 wire _1028_;
 wire _1029_;
 wire _1030_;
 wire _1031_;
 wire _1032_;
 wire _1033_;
 wire _1034_;
 wire _1035_;
 wire _1036_;
 wire _1037_;
 wire _1038_;
 wire _1039_;
 wire _1040_;
 wire _1041_;
 wire _1042_;
 wire _1043_;
 wire _1044_;
 wire _1045_;
 wire _1046_;
 wire _1047_;
 wire _1048_;
 wire _1049_;
 wire _1050_;
 wire _1051_;
 wire _1052_;
 wire _1053_;
 wire _1054_;
 wire _1055_;
 wire _1056_;
 wire _1057_;
 wire _1058_;
 wire _1059_;
 wire _1060_;
 wire _1061_;
 wire _1062_;
 wire _1063_;
 wire _1064_;
 wire _1065_;
 wire _1066_;
 wire _1067_;
 wire _1068_;
 wire _1069_;
 wire _1070_;
 wire _1071_;
 wire _1072_;
 wire _1073_;
 wire _1074_;
 wire _1075_;
 wire _1076_;
 wire _1077_;
 wire _1078_;
 wire _1079_;
 wire _1080_;
 wire _1081_;
 wire _1082_;
 wire _1083_;
 wire _1084_;
 wire _1085_;
 wire _1086_;
 wire _1087_;
 wire _1088_;
 wire _1089_;
 wire _1090_;
 wire _1091_;
 wire _1092_;
 wire _1093_;
 wire _1094_;
 wire _1095_;
 wire _1096_;
 wire _1097_;
 wire _1098_;
 wire _1099_;
 wire _1100_;
 wire _1101_;
 wire _1102_;
 wire _1103_;
 wire _1104_;
 wire _1105_;
 wire _1106_;
 wire _1107_;
 wire _1108_;
 wire _1109_;
 wire _1110_;
 wire _1111_;
 wire _1112_;
 wire _1113_;
 wire _1114_;
 wire _1115_;
 wire _1116_;
 wire _1117_;
 wire _1118_;
 wire _1119_;
 wire _1120_;
 wire _1121_;
 wire _1122_;
 wire _1123_;
 wire _1124_;
 wire _1125_;
 wire _1126_;
 wire _1127_;
 wire _1128_;
 wire _1129_;
 wire _1130_;
 wire _1131_;
 wire _1132_;
 wire _1133_;
 wire _1134_;
 wire _1135_;
 wire _1136_;
 wire _1137_;
 wire _1138_;
 wire _1139_;
 wire _1140_;
 wire _1141_;
 wire _1142_;
 wire _1143_;
 wire _1144_;
 wire _1145_;
 wire _1146_;
 wire _1147_;
 wire _1148_;
 wire _1149_;
 wire _1150_;
 wire _1151_;
 wire _1152_;
 wire _1153_;
 wire _1154_;
 wire _1155_;
 wire _1156_;
 wire _1157_;
 wire _1158_;
 wire _1159_;
 wire _1160_;
 wire _1161_;
 wire _1162_;
 wire _1163_;
 wire _1164_;
 wire _1165_;
 wire _1166_;
 wire _1167_;
 wire _1168_;
 wire _1169_;
 wire _1170_;
 wire _1171_;
 wire _1172_;
 wire _1173_;
 wire _1174_;
 wire _1175_;
 wire _1176_;
 wire _1177_;
 wire _1178_;
 wire _1179_;
 wire _1180_;
 wire _1181_;
 wire _1182_;
 wire _1183_;
 wire _1184_;
 wire _1185_;
 wire _1186_;
 wire _1187_;
 wire _1188_;
 wire _1189_;
 wire _1190_;
 wire _1191_;
 wire _1192_;
 wire _1193_;
 wire _1194_;
 wire _1195_;
 wire _1196_;
 wire _1197_;
 wire _1198_;
 wire _1199_;
 wire _1200_;
 wire _1201_;
 wire _1202_;
 wire _1203_;
 wire _1204_;
 wire _1205_;
 wire _1206_;
 wire _1207_;
 wire _1208_;
 wire _1209_;
 wire _1210_;
 wire _1211_;
 wire _1212_;
 wire _1213_;
 wire _1214_;
 wire _1215_;
 wire _1216_;
 wire _1217_;
 wire _1218_;
 wire _1219_;
 wire _1220_;
 wire _1221_;
 wire _1222_;
 wire _1223_;
 wire _1224_;
 wire _1225_;
 wire _1226_;
 wire _1227_;
 wire _1228_;
 wire _1229_;
 wire _1230_;
 wire _1231_;
 wire _1232_;
 wire _1233_;
 wire _1234_;
 wire _1235_;
 wire _1236_;
 wire _1237_;
 wire _1238_;
 wire _1239_;
 wire _1240_;
 wire _1241_;
 wire _1242_;
 wire _1243_;
 wire _1244_;
 wire _1245_;
 wire _1246_;
 wire _1247_;
 wire _1248_;
 wire _1249_;
 wire _1250_;
 wire _1251_;
 wire _1252_;
 wire _1253_;
 wire _1254_;
 wire _1255_;
 wire _1256_;
 wire _1257_;
 wire _1258_;
 wire _1259_;
 wire _1260_;
 wire _1261_;
 wire _1262_;
 wire _1263_;
 wire _1264_;
 wire _1265_;
 wire _1266_;
 wire _1267_;
 wire _1268_;
 wire _1269_;
 wire _1270_;
 wire _1271_;
 wire _1272_;
 wire _1273_;
 wire _1274_;
 wire _1275_;
 wire _1276_;
 wire _1277_;
 wire _1278_;
 wire _1279_;
 wire _1280_;
 wire _1281_;
 wire _1282_;
 wire _1283_;
 wire _1284_;
 wire _1285_;
 wire _1286_;
 wire _1287_;
 wire _1288_;
 wire _1289_;
 wire _1290_;
 wire _1291_;
 wire _1292_;
 wire _1293_;
 wire _1294_;
 wire _1295_;
 wire _1296_;
 wire _1297_;
 wire _1298_;
 wire _1299_;
 wire _1300_;
 wire _1301_;
 wire _1302_;
 wire _1303_;
 wire _1304_;
 wire _1305_;
 wire _1306_;
 wire _1307_;
 wire _1308_;
 wire _1309_;
 wire _1310_;
 wire _1311_;
 wire _1312_;
 wire _1313_;
 wire _1314_;
 wire _1315_;
 wire _1316_;
 wire _1317_;
 wire _1318_;
 wire _1319_;
 wire _1320_;
 wire _1321_;
 wire _1322_;
 wire _1323_;
 wire _1324_;
 wire _1325_;
 wire _1326_;
 wire _1327_;
 wire _1328_;
 wire _1329_;
 wire _1330_;
 wire _1331_;
 wire _1332_;
 wire _1333_;
 wire _1334_;
 wire _1335_;
 wire _1336_;
 wire _1337_;
 wire _1338_;
 wire _1339_;
 wire _1340_;
 wire _1341_;
 wire _1342_;
 wire _1343_;
 wire _1344_;
 wire _1345_;
 wire _1346_;
 wire _1347_;
 wire _1348_;
 wire _1349_;
 wire _1350_;
 wire _1351_;
 wire _1352_;
 wire _1353_;
 wire _1354_;
 wire _1355_;
 wire _1356_;
 wire _1357_;
 wire _1358_;
 wire _1359_;
 wire _1360_;
 wire _1361_;
 wire _1362_;
 wire _1363_;
 wire _1364_;
 wire _1365_;
 wire _1366_;
 wire _1367_;
 wire _1368_;
 wire _1369_;
 wire _1370_;
 wire _1371_;
 wire _1372_;
 wire _1373_;
 wire _1374_;
 wire _1375_;
 wire _1376_;
 wire _1377_;
 wire _1378_;
 wire _1379_;
 wire _1380_;
 wire _1381_;
 wire _1382_;
 wire _1383_;
 wire _1384_;
 wire _1385_;
 wire _1386_;
 wire _1387_;
 wire _1388_;
 wire _1389_;
 wire _1390_;
 wire _1391_;
 wire _1392_;
 wire _1393_;
 wire _1394_;
 wire _1395_;
 wire _1396_;
 wire _1397_;
 wire _1398_;
 wire _1399_;
 wire _1400_;
 wire _1401_;
 wire _1402_;
 wire _1403_;
 wire _1404_;
 wire _1405_;
 wire _1406_;
 wire _1407_;
 wire _1408_;
 wire _1409_;
 wire _1410_;
 wire _1411_;
 wire _1412_;
 wire _1413_;
 wire _1414_;
 wire _1415_;
 wire _1416_;
 wire _1417_;
 wire _1418_;
 wire _1419_;
 wire _1420_;
 wire _1421_;
 wire _1422_;
 wire _1423_;
 wire _1424_;
 wire _1425_;
 wire _1426_;
 wire _1427_;
 wire _1428_;
 wire _1429_;
 wire _1430_;
 wire _1431_;
 wire _1432_;
 wire _1433_;
 wire _1434_;
 wire _1435_;
 wire _1436_;
 wire _1437_;
 wire _1438_;
 wire _1439_;
 wire _1440_;
 wire _1441_;
 wire _1442_;
 wire _1443_;
 wire _1444_;
 wire _1445_;
 wire _1446_;
 wire _1447_;
 wire _1448_;
 wire _1449_;
 wire _1450_;
 wire _1451_;
 wire _1452_;
 wire _1453_;
 wire _1454_;
 wire _1455_;
 wire _1456_;
 wire _1457_;
 wire _1458_;
 wire _1459_;
 wire _1460_;
 wire _1461_;
 wire _1462_;
 wire _1463_;
 wire _1464_;
 wire _1465_;
 wire _1466_;
 wire _1467_;
 wire _1468_;
 wire _1469_;
 wire _1470_;
 wire _1471_;
 wire _1472_;
 wire _1473_;
 wire _1474_;
 wire _1475_;
 wire _1476_;
 wire _1477_;
 wire _1478_;
 wire _1479_;
 wire _1480_;
 wire _1481_;
 wire _1482_;
 wire _1483_;
 wire _1484_;
 wire _1485_;
 wire _1486_;
 wire _1487_;
 wire _1488_;
 wire _1489_;
 wire _1490_;
 wire _1491_;
 wire _1492_;
 wire _1493_;
 wire _1494_;
 wire _1495_;
 wire _1496_;
 wire _1497_;
 wire _1498_;
 wire _1499_;
 wire _1500_;
 wire _1501_;
 wire _1502_;
 wire _1503_;
 wire _1504_;
 wire _1505_;
 wire _1506_;
 wire _1507_;
 wire _1508_;
 wire _1509_;
 wire _1510_;
 wire _1511_;
 wire _1512_;
 wire _1513_;
 wire _1514_;
 wire _1515_;
 wire _1516_;
 wire _1517_;
 wire _1518_;
 wire _1519_;
 wire _1520_;
 wire _1521_;
 wire _1522_;
 wire _1523_;
 wire _1524_;
 wire _1525_;
 wire _1526_;
 wire _1527_;
 wire _1528_;
 wire _1529_;
 wire _1530_;
 wire _1531_;
 wire _1532_;
 wire _1533_;
 wire _1534_;
 wire _1535_;
 wire _1536_;
 wire _1537_;
 wire _1538_;
 wire _1539_;
 wire _1540_;
 wire _1541_;
 wire _1542_;
 wire _1543_;
 wire _1544_;
 wire _1545_;
 wire _1546_;
 wire _1547_;
 wire _1548_;
 wire _1549_;
 wire _1550_;
 wire _1551_;
 wire _1552_;
 wire _1553_;
 wire _1554_;
 wire _1555_;
 wire _1556_;
 wire _1557_;
 wire _1558_;
 wire _1559_;
 wire _1560_;
 wire _1561_;
 wire _1562_;
 wire _1563_;
 wire _1564_;
 wire _1565_;
 wire _1566_;
 wire _1567_;
 wire _1568_;
 wire _1569_;
 wire _1570_;
 wire _1571_;
 wire _1572_;
 wire _1573_;
 wire _1574_;
 wire _1575_;
 wire _1576_;
 wire _1577_;
 wire _1578_;
 wire _1579_;
 wire _1580_;
 wire _1581_;
 wire _1582_;
 wire _1583_;
 wire _1584_;
 wire _1585_;
 wire _1586_;
 wire _1587_;
 wire _1588_;
 wire _1589_;
 wire _1590_;
 wire _1591_;
 wire _1592_;
 wire _1593_;
 wire _1594_;
 wire _1595_;
 wire _1596_;
 wire _1597_;
 wire _1598_;
 wire _1599_;
 wire _1600_;
 wire _1601_;
 wire _1602_;
 wire _1603_;
 wire _1604_;
 wire _1605_;
 wire _1606_;
 wire _1607_;
 wire _1608_;
 wire _1609_;
 wire _1610_;
 wire _1611_;
 wire _1612_;
 wire _1613_;
 wire _1614_;
 wire _1615_;
 wire _1616_;
 wire _1617_;
 wire _1618_;
 wire _1619_;
 wire _1620_;
 wire _1621_;
 wire _1622_;
 wire _1623_;
 wire _1624_;
 wire _1625_;
 wire _1626_;
 wire _1627_;
 wire _1628_;
 wire _1629_;
 wire _1630_;
 wire _1631_;
 wire _1632_;
 wire _1633_;
 wire _1634_;
 wire _1635_;
 wire _1636_;
 wire _1637_;
 wire _1638_;
 wire _1639_;
 wire _1640_;
 wire _1641_;
 wire _1642_;
 wire _1643_;
 wire _1644_;
 wire _1645_;
 wire _1646_;
 wire _1647_;
 wire _1648_;
 wire _1649_;
 wire _1650_;
 wire _1651_;
 wire _1652_;
 wire _1653_;
 wire _1654_;
 wire _1655_;
 wire _1656_;
 wire _1657_;
 wire _1658_;
 wire _1659_;
 wire _1660_;
 wire _1661_;
 wire _1662_;
 wire _1663_;
 wire _1664_;
 wire _1665_;
 wire _1666_;
 wire _1667_;
 wire _1668_;
 wire _1669_;
 wire _1670_;
 wire _1671_;
 wire _1672_;
 wire _1673_;
 wire _1674_;
 wire _1675_;
 wire _1676_;
 wire _1677_;
 wire _1678_;
 wire _1679_;
 wire _1680_;
 wire _1681_;
 wire _1682_;
 wire _1683_;
 wire _1684_;
 wire _1685_;
 wire _1686_;
 wire _1687_;
 wire _1688_;
 wire _1689_;
 wire _1690_;
 wire _1691_;
 wire _1692_;
 wire _1693_;
 wire _1694_;
 wire _1695_;
 wire _1696_;
 wire _1697_;
 wire _1698_;
 wire _1699_;
 wire _1700_;
 wire _1701_;
 wire _1702_;
 wire _1703_;
 wire _1704_;
 wire _1705_;
 wire _1706_;
 wire _1707_;
 wire _1708_;
 wire _1709_;
 wire _1710_;
 wire _1711_;
 wire _1712_;
 wire _1713_;
 wire _1714_;
 wire _1715_;
 wire _1716_;
 wire _1717_;
 wire _1718_;
 wire _1719_;
 wire _1720_;
 wire _1721_;
 wire _1722_;
 wire _1723_;
 wire _1724_;
 wire _1725_;
 wire _1726_;
 wire _1727_;
 wire _1728_;
 wire _1729_;
 wire _1730_;
 wire _1731_;
 wire _1732_;
 wire _1733_;
 wire _1734_;
 wire _1735_;
 wire _1736_;
 wire _1737_;
 wire _1738_;
 wire _1739_;
 wire _1740_;
 wire _1741_;
 wire _1742_;
 wire _1743_;
 wire _1744_;
 wire _1745_;
 wire _1746_;
 wire _1747_;
 wire _1748_;
 wire _1749_;
 wire _1750_;
 wire _1751_;
 wire _1752_;
 wire _1753_;
 wire _1754_;
 wire _1755_;
 wire _1756_;
 wire _1757_;
 wire _1758_;
 wire _1759_;
 wire _1760_;
 wire _1761_;
 wire _1762_;
 wire _1763_;
 wire _1764_;
 wire _1765_;
 wire _1766_;
 wire _1767_;
 wire _1768_;
 wire _1769_;
 wire _1770_;
 wire _1771_;
 wire _1772_;
 wire _1773_;
 wire _1774_;
 wire _1775_;
 wire _1776_;
 wire _1777_;
 wire _1778_;
 wire _1779_;
 wire _1780_;
 wire _1781_;
 wire _1782_;
 wire _1783_;
 wire _1784_;
 wire _1785_;
 wire _1786_;
 wire _1787_;
 wire _1788_;
 wire _1789_;
 wire _1790_;
 wire _1791_;
 wire _1792_;
 wire _1793_;
 wire _1794_;
 wire _1795_;
 wire _1796_;
 wire _1797_;
 wire _1798_;
 wire _1799_;
 wire _1800_;
 wire _1801_;
 wire _1802_;
 wire _1803_;
 wire _1804_;
 wire _1805_;
 wire _1806_;
 wire _1807_;
 wire _1808_;
 wire _1809_;
 wire _1810_;
 wire _1811_;
 wire _1812_;
 wire _1813_;
 wire _1814_;
 wire _1815_;
 wire _1816_;
 wire _1817_;
 wire _1818_;
 wire _1819_;
 wire _1820_;
 wire _1821_;
 wire _1822_;
 wire _1823_;
 wire _1824_;
 wire _1825_;
 wire _1826_;
 wire _1827_;
 wire _1828_;
 wire _1829_;
 wire _1830_;
 wire _1831_;
 wire _1832_;
 wire _1833_;
 wire _1834_;
 wire _1835_;
 wire _1836_;
 wire _1837_;
 wire _1838_;
 wire _1839_;
 wire _1840_;
 wire _1841_;
 wire _1842_;
 wire _1843_;
 wire _1844_;
 wire _1845_;
 wire _1846_;
 wire _1847_;
 wire _1848_;
 wire _1849_;
 wire _1850_;
 wire _1851_;
 wire _1852_;
 wire _1853_;
 wire _1854_;
 wire _1855_;
 wire _1856_;
 wire _1857_;
 wire _1858_;
 wire _1859_;
 wire _1860_;
 wire _1861_;
 wire _1862_;
 wire _1863_;
 wire _1864_;
 wire _1865_;
 wire _1866_;
 wire _1867_;
 wire _1868_;
 wire _1869_;
 wire _1870_;
 wire _1871_;
 wire _1872_;
 wire _1873_;
 wire _1874_;
 wire _1875_;
 wire _1876_;
 wire _1877_;
 wire _1878_;
 wire _1879_;
 wire _1880_;
 wire _1881_;
 wire _1882_;
 wire _1883_;
 wire _1884_;
 wire _1885_;
 wire _1886_;
 wire _1887_;
 wire _1888_;
 wire _1889_;
 wire _1890_;
 wire _1891_;
 wire _1892_;
 wire _1893_;
 wire _1894_;
 wire _1895_;
 wire _1896_;
 wire _1897_;
 wire _1898_;
 wire _1899_;
 wire _1900_;
 wire _1901_;
 wire _1902_;
 wire _1903_;
 wire _1904_;
 wire _1905_;
 wire _1906_;
 wire _1907_;
 wire _1908_;
 wire _1909_;
 wire _1910_;
 wire _1911_;
 wire _1912_;
 wire _1913_;
 wire _1914_;
 wire _1915_;
 wire _1916_;
 wire _1917_;
 wire _1918_;
 wire _1919_;
 wire _1920_;
 wire _1921_;
 wire _1922_;
 wire _1923_;
 wire _1924_;
 wire _1925_;
 wire _1926_;
 wire _1927_;
 wire _1928_;
 wire _1929_;
 wire _1930_;
 wire _1931_;
 wire _1932_;
 wire _1933_;
 wire _1934_;
 wire _1935_;
 wire _1936_;
 wire _1937_;
 wire _1938_;
 wire _1939_;
 wire _1940_;
 wire _1941_;
 wire _1942_;
 wire _1943_;
 wire _1944_;
 wire _1945_;
 wire _1946_;
 wire _1947_;
 wire _1948_;
 wire _1949_;
 wire _1950_;
 wire _1951_;
 wire _1952_;
 wire _1953_;
 wire _1954_;
 wire _1955_;
 wire _1956_;
 wire _1957_;
 wire _1958_;
 wire _1959_;
 wire _1960_;
 wire _1961_;
 wire _1962_;
 wire _1963_;
 wire _1964_;
 wire _1965_;
 wire _1966_;
 wire _1967_;
 wire _1968_;
 wire _1969_;
 wire _1970_;
 wire _1971_;
 wire _1972_;
 wire _1973_;
 wire _1974_;
 wire _1975_;
 wire _1976_;
 wire _1977_;
 wire _1978_;
 wire _1979_;
 wire _1980_;
 wire _1981_;
 wire _1982_;
 wire _1983_;
 wire _1984_;
 wire _1985_;
 wire _1986_;
 wire _1987_;
 wire _1988_;
 wire _1989_;
 wire _1990_;
 wire _1991_;
 wire _1992_;
 wire _1993_;
 wire _1994_;
 wire _1995_;
 wire _1996_;
 wire _1997_;
 wire _1998_;
 wire _1999_;
 wire _2000_;
 wire _2001_;
 wire _2002_;
 wire _2003_;
 wire _2004_;
 wire _2005_;
 wire _2006_;
 wire _2007_;
 wire _2008_;
 wire _2009_;
 wire _2010_;
 wire _2011_;
 wire _2012_;
 wire _2013_;
 wire _2014_;
 wire _2015_;
 wire _2016_;
 wire _2017_;
 wire _2018_;
 wire _2019_;
 wire _2020_;
 wire _2021_;
 wire _2022_;
 wire _2023_;
 wire _2024_;
 wire _2025_;
 wire _2026_;
 wire _2027_;
 wire _2028_;
 wire _2029_;
 wire _2030_;
 wire _2031_;
 wire _2032_;
 wire _2033_;
 wire _2034_;
 wire _2035_;
 wire _2036_;
 wire _2037_;
 wire _2038_;
 wire _2039_;
 wire _2040_;
 wire _2041_;
 wire _2042_;
 wire _2043_;
 wire _2044_;
 wire _2045_;
 wire _2046_;
 wire _2047_;
 wire _2048_;
 wire _2049_;
 wire _2050_;
 wire _2051_;
 wire _2052_;
 wire _2053_;
 wire _2054_;
 wire _2055_;
 wire _2056_;
 wire _2057_;
 wire _2058_;
 wire _2059_;
 wire _2060_;
 wire _2061_;
 wire _2062_;
 wire _2063_;
 wire _2064_;
 wire _2065_;
 wire _2066_;
 wire _2067_;
 wire _2068_;
 wire _2069_;
 wire _2070_;
 wire _2071_;
 wire _2072_;
 wire _2073_;
 wire _2074_;
 wire _2075_;
 wire _2076_;
 wire _2077_;
 wire _2078_;
 wire _2079_;
 wire _2080_;
 wire _2081_;
 wire _2082_;
 wire _2083_;
 wire _2084_;
 wire _2085_;
 wire _2086_;
 wire _2087_;
 wire _2088_;
 wire _2089_;
 wire _2090_;
 wire _2091_;
 wire _2092_;
 wire _2093_;
 wire _2094_;
 wire _2095_;
 wire _2096_;
 wire _2097_;
 wire _2098_;
 wire _2099_;
 wire _2100_;
 wire _2101_;
 wire _2102_;
 wire _2103_;
 wire _2104_;
 wire _2105_;
 wire _2106_;
 wire _2107_;
 wire _2108_;
 wire _2109_;
 wire _2110_;
 wire _2111_;
 wire _2112_;
 wire _2113_;
 wire _2114_;
 wire _2115_;
 wire _2116_;
 wire _2117_;
 wire _2118_;
 wire _2119_;
 wire _2120_;
 wire _2121_;
 wire _2122_;
 wire _2123_;
 wire _2124_;
 wire _2125_;
 wire _2126_;
 wire _2127_;
 wire _2128_;
 wire _2129_;
 wire _2130_;
 wire _2131_;
 wire _2132_;
 wire _2133_;
 wire _2134_;
 wire _2135_;
 wire _2136_;
 wire _2137_;
 wire _2138_;
 wire _2139_;
 wire _2140_;
 wire _2141_;
 wire _2142_;
 wire _2143_;
 wire _2144_;
 wire _2145_;
 wire _2146_;
 wire _2147_;
 wire _2148_;
 wire _2149_;
 wire _2150_;
 wire _2151_;
 wire _2152_;
 wire _2153_;
 wire _2154_;
 wire _2155_;
 wire _2156_;
 wire _2157_;
 wire _2158_;
 wire _2159_;
 wire _2160_;
 wire _2161_;
 wire _2162_;
 wire _2163_;
 wire _2164_;
 wire _2165_;
 wire _2166_;
 wire _2167_;
 wire _2168_;
 wire _2169_;
 wire _2170_;
 wire _2171_;
 wire _2172_;
 wire _2173_;
 wire _2174_;
 wire _2175_;
 wire _2176_;
 wire _2177_;
 wire _2178_;
 wire _2179_;
 wire _2180_;
 wire _2181_;
 wire _2182_;
 wire _2183_;
 wire _2184_;
 wire _2185_;
 wire _2186_;
 wire _2187_;
 wire _2188_;
 wire _2189_;
 wire _2190_;
 wire _2191_;
 wire _2192_;
 wire _2193_;
 wire _2194_;
 wire _2195_;
 wire _2196_;
 wire _2197_;
 wire _2198_;
 wire _2199_;
 wire _2200_;
 wire _2201_;
 wire _2202_;
 wire _2203_;
 wire _2204_;
 wire _2205_;
 wire _2206_;
 wire _2207_;
 wire _2208_;
 wire _2209_;
 wire _2210_;
 wire _2211_;
 wire _2212_;
 wire _2213_;
 wire _2214_;
 wire _2215_;
 wire _2216_;
 wire _2217_;
 wire _2218_;
 wire _2219_;
 wire _2220_;
 wire _2221_;
 wire _2222_;
 wire _2223_;
 wire _2224_;
 wire _2225_;
 wire _2226_;
 wire _2227_;
 wire _2228_;
 wire _2229_;
 wire _2230_;
 wire _2231_;
 wire _2232_;
 wire _2233_;
 wire _2234_;
 wire _2235_;
 wire _2236_;
 wire _2237_;
 wire _2238_;
 wire _2239_;
 wire _2240_;
 wire _2241_;
 wire _2242_;
 wire _2243_;
 wire _2244_;
 wire _2245_;
 wire _2246_;
 wire _2247_;
 wire _2248_;
 wire _2249_;
 wire _2250_;
 wire _2251_;
 wire _2252_;
 wire _2253_;
 wire _2254_;
 wire _2255_;
 wire _2256_;
 wire _2257_;
 wire _2258_;
 wire _2259_;
 wire _2260_;
 wire _2261_;
 wire _2262_;
 wire _2263_;
 wire _2264_;
 wire _2265_;
 wire _2266_;
 wire _2267_;
 wire _2268_;
 wire _2269_;
 wire _2270_;
 wire _2271_;
 wire _2272_;
 wire _2273_;
 wire _2274_;
 wire _2275_;
 wire _2276_;
 wire _2277_;
 wire _2278_;
 wire _2279_;
 wire _2280_;
 wire _2281_;
 wire _2282_;
 wire _2283_;
 wire _2284_;
 wire _2285_;
 wire _2286_;
 wire _2287_;
 wire _2288_;
 wire _2289_;
 wire _2290_;
 wire _2291_;
 wire _2292_;
 wire _2293_;
 wire _2294_;
 wire _2295_;
 wire _2296_;
 wire _2297_;
 wire _2298_;
 wire _2299_;
 wire _2300_;
 wire _2301_;
 wire _2302_;
 wire _2303_;
 wire _2304_;
 wire _2305_;
 wire _2306_;
 wire _2307_;
 wire _2308_;
 wire _2309_;
 wire _2310_;
 wire _2311_;
 wire _2312_;
 wire _2313_;
 wire _2314_;
 wire _2315_;
 wire _2316_;
 wire _2317_;
 wire _2318_;
 wire _2319_;
 wire _2320_;
 wire _2321_;
 wire _2322_;
 wire _2323_;
 wire _2324_;
 wire _2325_;
 wire _2326_;
 wire _2327_;
 wire _2328_;
 wire _2329_;
 wire _2330_;
 wire _2331_;
 wire _2332_;
 wire _2333_;
 wire _2334_;
 wire _2335_;
 wire _2336_;
 wire _2337_;
 wire _2338_;
 wire _2339_;
 wire _2340_;
 wire _2341_;
 wire _2342_;
 wire _2343_;
 wire _2344_;
 wire _2345_;
 wire _2346_;
 wire _2347_;
 wire _2348_;
 wire _2349_;
 wire _2350_;
 wire _2351_;
 wire _2352_;
 wire _2353_;
 wire _2354_;
 wire _2355_;
 wire _2356_;
 wire _2357_;
 wire _2358_;
 wire _2359_;
 wire _2360_;
 wire _2361_;
 wire _2362_;
 wire _2363_;
 wire _2364_;
 wire _2365_;
 wire _2366_;
 wire _2367_;
 wire _2368_;
 wire _2369_;
 wire _2370_;
 wire _2371_;
 wire _2372_;
 wire _2373_;
 wire _2374_;
 wire _2375_;
 wire _2376_;
 wire _2377_;
 wire _2378_;
 wire _2379_;
 wire _2380_;
 wire _2381_;
 wire _2382_;
 wire _2383_;
 wire _2384_;
 wire _2385_;
 wire _2386_;
 wire _2387_;
 wire _2388_;
 wire _2389_;
 wire _2390_;
 wire _2391_;
 wire _2392_;
 wire _2393_;
 wire _2394_;
 wire _2395_;
 wire _2396_;
 wire _2397_;
 wire _2398_;
 wire _2399_;
 wire _2400_;
 wire _2401_;
 wire _2402_;
 wire _2403_;
 wire _2404_;
 wire _2405_;
 wire _2406_;
 wire _2407_;
 wire _2408_;
 wire _2409_;
 wire _2410_;
 wire _2411_;
 wire _2412_;
 wire _2413_;
 wire _2414_;
 wire _2415_;
 wire _2416_;
 wire _2417_;
 wire _2418_;
 wire _2419_;
 wire _2420_;
 wire _2421_;
 wire _2422_;
 wire _2423_;
 wire _2424_;
 wire _2425_;
 wire _2426_;
 wire _2427_;
 wire _2428_;
 wire _2429_;
 wire _2430_;
 wire _2431_;
 wire _2432_;
 wire _2433_;
 wire _2434_;
 wire _2435_;
 wire _2436_;
 wire _2437_;
 wire _2438_;
 wire _2439_;
 wire _2440_;
 wire _2441_;
 wire _2442_;
 wire _2443_;
 wire _2444_;
 wire _2445_;
 wire _2446_;
 wire _2447_;
 wire _2448_;
 wire _2449_;
 wire _2450_;
 wire _2451_;
 wire _2452_;
 wire _2453_;
 wire _2454_;
 wire _2455_;
 wire _2456_;
 wire _2457_;
 wire _2458_;
 wire _2459_;
 wire _2460_;
 wire _2461_;
 wire _2462_;
 wire _2463_;
 wire _2464_;
 wire _2465_;
 wire _2466_;
 wire _2467_;
 wire _2468_;
 wire _2469_;
 wire _2470_;
 wire _2471_;
 wire _2472_;
 wire _2473_;
 wire _2474_;
 wire _2475_;
 wire _2476_;
 wire _2477_;
 wire _2478_;
 wire _2479_;
 wire _2480_;
 wire _2481_;
 wire _2482_;
 wire _2483_;
 wire _2484_;
 wire _2485_;
 wire _2486_;
 wire _2487_;
 wire _2488_;
 wire _2489_;
 wire _2490_;
 wire _2491_;
 wire _2492_;
 wire _2493_;
 wire _2494_;
 wire _2495_;
 wire _2496_;
 wire _2497_;
 wire _2498_;
 wire _2499_;
 wire _2500_;
 wire _2501_;
 wire _2502_;
 wire _2503_;
 wire _2504_;
 wire _2505_;
 wire _2506_;
 wire _2507_;
 wire _2508_;
 wire _2509_;
 wire _2510_;
 wire _2511_;
 wire _2512_;
 wire _2513_;
 wire _2514_;
 wire _2515_;
 wire _2516_;
 wire _2517_;
 wire _2518_;
 wire _2519_;
 wire _2520_;
 wire _2521_;
 wire _2522_;
 wire _2523_;
 wire _2524_;
 wire _2525_;
 wire _2526_;
 wire _2527_;
 wire _2528_;
 wire _2529_;
 wire _2530_;
 wire _2531_;
 wire _2532_;
 wire _2533_;
 wire _2534_;
 wire _2535_;
 wire _2536_;
 wire _2537_;
 wire _2538_;
 wire _2539_;
 wire _2540_;
 wire _2541_;
 wire _2542_;
 wire _2543_;
 wire _2544_;
 wire _2545_;
 wire _2546_;
 wire _2547_;
 wire _2548_;
 wire _2549_;
 wire _2550_;
 wire _2551_;
 wire _2552_;
 wire _2553_;
 wire _2554_;
 wire _2555_;
 wire _2556_;
 wire _2557_;
 wire _2558_;
 wire _2559_;
 wire _2560_;
 wire _2561_;
 wire _2562_;
 wire _2563_;
 wire _2564_;
 wire _2565_;
 wire _2566_;
 wire _2567_;
 wire _2568_;
 wire _2569_;
 wire _2570_;
 wire _2571_;
 wire _2572_;
 wire _2573_;
 wire _2574_;
 wire _2575_;
 wire _2576_;
 wire _2577_;
 wire _2578_;
 wire _2579_;
 wire _2580_;
 wire _2581_;
 wire _2582_;
 wire _2583_;
 wire _2584_;
 wire _2585_;
 wire _2586_;
 wire _2587_;
 wire _2588_;
 wire _2589_;
 wire _2590_;
 wire _2591_;
 wire _2592_;
 wire _2593_;
 wire _2594_;
 wire _2595_;
 wire _2596_;
 wire _2597_;
 wire _2598_;
 wire _2599_;
 wire _2600_;
 wire _2601_;
 wire _2602_;
 wire _2603_;
 wire _2604_;
 wire _2605_;
 wire _2606_;
 wire _2607_;
 wire _2608_;
 wire _2609_;
 wire _2610_;
 wire _2611_;
 wire _2612_;
 wire _2613_;
 wire _2614_;
 wire _2615_;
 wire _2616_;
 wire _2617_;
 wire _2618_;
 wire _2619_;
 wire _2620_;
 wire _2621_;
 wire _2622_;
 wire _2623_;
 wire _2624_;
 wire _2625_;
 wire _2626_;
 wire _2627_;
 wire _2628_;
 wire _2629_;
 wire _2630_;
 wire _2631_;
 wire _2632_;
 wire _2633_;
 wire _2634_;
 wire _2635_;
 wire _2636_;
 wire _2637_;
 wire _2638_;
 wire _2639_;
 wire _2640_;
 wire _2641_;
 wire _2642_;
 wire _2643_;
 wire _2644_;
 wire _2645_;
 wire _2646_;
 wire _2647_;
 wire _2648_;
 wire _2649_;
 wire _2650_;
 wire _2651_;
 wire _2652_;
 wire _2653_;
 wire _2654_;
 wire _2655_;
 wire _2656_;
 wire _2657_;
 wire _2658_;
 wire _2659_;
 wire _2660_;
 wire _2661_;
 wire _2662_;
 wire _2663_;
 wire _2664_;
 wire _2665_;
 wire _2666_;
 wire _2667_;
 wire _2668_;
 wire _2669_;
 wire _2670_;
 wire _2671_;
 wire _2672_;
 wire _2673_;
 wire _2674_;
 wire _2675_;
 wire _2676_;
 wire _2677_;
 wire _2678_;
 wire _2679_;
 wire _2680_;
 wire _2681_;
 wire _2682_;
 wire _2683_;
 wire _2684_;
 wire _2685_;
 wire _2686_;
 wire _2687_;
 wire _2688_;
 wire _2689_;
 wire _2690_;
 wire _2691_;
 wire _2692_;
 wire _2693_;
 wire _2694_;
 wire _2695_;
 wire _2696_;
 wire _2697_;
 wire _2698_;
 wire _2699_;
 wire _2700_;
 wire _2701_;
 wire _2702_;
 wire _2703_;
 wire _2704_;
 wire _2705_;
 wire _2706_;
 wire _2707_;
 wire _2708_;
 wire _2709_;
 wire _2710_;
 wire _2711_;
 wire _2712_;
 wire _2713_;
 wire _2714_;
 wire _2715_;
 wire _2716_;
 wire _2717_;
 wire _2718_;
 wire _2719_;
 wire _2720_;
 wire _2721_;
 wire _2722_;
 wire _2723_;
 wire _2724_;
 wire _2725_;
 wire _2726_;
 wire _2727_;
 wire _2728_;
 wire _2729_;
 wire _2730_;
 wire _2731_;
 wire _2732_;
 wire _2733_;
 wire _2734_;
 wire _2735_;
 wire _2736_;
 wire _2737_;
 wire _2738_;
 wire _2739_;
 wire _2740_;
 wire _2741_;
 wire _2742_;
 wire _2743_;
 wire _2744_;
 wire _2745_;
 wire _2746_;
 wire _2747_;
 wire _2748_;
 wire _2749_;
 wire _2750_;
 wire _2751_;
 wire _2752_;
 wire _2753_;
 wire _2754_;
 wire _2755_;
 wire _2756_;
 wire _2757_;
 wire _2758_;
 wire _2759_;
 wire _2760_;
 wire _2761_;
 wire _2762_;
 wire _2763_;
 wire _2764_;
 wire _2765_;
 wire _2766_;
 wire _2767_;
 wire _2768_;
 wire _2769_;
 wire _2770_;
 wire _2771_;
 wire _2772_;
 wire _2773_;
 wire _2774_;
 wire _2775_;
 wire _2776_;
 wire _2777_;
 wire _2778_;
 wire _2779_;
 wire _2780_;
 wire _2781_;
 wire _2782_;
 wire _2783_;
 wire _2784_;
 wire _2785_;
 wire _2786_;
 wire _2787_;
 wire _2788_;
 wire _2789_;
 wire _2790_;
 wire _2791_;
 wire _2792_;
 wire _2793_;
 wire _2794_;
 wire _2795_;
 wire _2796_;
 wire _2797_;
 wire _2798_;
 wire _2799_;
 wire _2800_;
 wire _2801_;
 wire _2802_;
 wire _2803_;
 wire _2804_;
 wire _2805_;
 wire _2806_;
 wire _2807_;
 wire _2808_;
 wire _2809_;
 wire _2810_;
 wire _2811_;
 wire _2812_;
 wire _2813_;
 wire _2814_;
 wire _2815_;
 wire _2816_;
 wire _2817_;
 wire _2818_;
 wire _2819_;
 wire _2820_;
 wire _2821_;
 wire _2822_;
 wire _2823_;
 wire _2824_;
 wire _2825_;
 wire _2826_;
 wire _2827_;
 wire _2828_;
 wire _2829_;
 wire _2830_;
 wire _2831_;
 wire _2832_;
 wire _2833_;
 wire _2834_;
 wire _2835_;
 wire _2836_;
 wire _2837_;
 wire _2838_;
 wire _2839_;
 wire _2840_;
 wire _2841_;
 wire _2842_;
 wire _2843_;
 wire _2844_;
 wire _2845_;
 wire _2846_;
 wire _2847_;
 wire _2848_;
 wire _2849_;
 wire _2850_;
 wire _2851_;
 wire _2852_;
 wire _2853_;
 wire _2854_;
 wire _2855_;
 wire _2856_;
 wire _2857_;
 wire _2858_;
 wire _2859_;
 wire _2860_;
 wire _2861_;
 wire _2862_;
 wire _2863_;
 wire _2864_;
 wire _2865_;
 wire _2866_;
 wire _2867_;
 wire _2868_;
 wire _2869_;
 wire _2870_;
 wire _2871_;
 wire _2872_;
 wire _2873_;
 wire _2874_;
 wire _2875_;
 wire _2876_;
 wire _2877_;
 wire _2878_;
 wire _2879_;
 wire _2880_;
 wire _2881_;
 wire _2882_;
 wire _2883_;
 wire _2884_;
 wire _2885_;
 wire _2886_;
 wire _2887_;
 wire _2888_;
 wire _2889_;
 wire _2890_;
 wire _2891_;
 wire _2892_;
 wire _2893_;
 wire _2894_;
 wire _2895_;
 wire _2896_;
 wire _2897_;
 wire _2898_;
 wire _2899_;
 wire _2900_;
 wire _2901_;
 wire _2902_;
 wire _2903_;
 wire _2904_;
 wire _2905_;
 wire _2906_;
 wire _2907_;
 wire _2908_;
 wire _2909_;
 wire _2910_;
 wire _2911_;
 wire _2912_;
 wire _2913_;
 wire _2914_;
 wire _2915_;
 wire _2916_;
 wire _2917_;
 wire _2918_;
 wire _2919_;
 wire _2920_;
 wire _2921_;
 wire _2922_;
 wire _2923_;
 wire _2924_;
 wire _2925_;
 wire _2926_;
 wire _2927_;
 wire _2928_;
 wire _2929_;
 wire _2930_;
 wire _2931_;
 wire _2932_;
 wire _2933_;
 wire _2934_;
 wire _2935_;
 wire _2936_;
 wire _2937_;
 wire _2938_;
 wire _2939_;
 wire _2940_;
 wire _2941_;
 wire _2942_;
 wire _2943_;
 wire _2944_;
 wire _2945_;
 wire _2946_;
 wire _2947_;
 wire _2948_;
 wire _2949_;
 wire _2950_;
 wire _2951_;
 wire _2952_;
 wire _2953_;
 wire _2954_;
 wire _2955_;
 wire _2956_;
 wire _2957_;
 wire _2958_;
 wire _2959_;
 wire _2960_;
 wire _2961_;
 wire _2962_;
 wire _2963_;
 wire _2964_;
 wire _2965_;
 wire _2966_;
 wire _2967_;
 wire _2968_;
 wire _2969_;
 wire _2970_;
 wire _2971_;
 wire _2972_;
 wire _2973_;
 wire _2974_;
 wire _2975_;
 wire _2976_;
 wire _2977_;
 wire _2978_;
 wire _2979_;
 wire _2980_;
 wire _2981_;
 wire _2982_;
 wire _2983_;
 wire _2984_;
 wire _2985_;
 wire _2986_;
 wire _2987_;
 wire _2988_;
 wire _2989_;
 wire _2990_;
 wire _2991_;
 wire _2992_;
 wire _2993_;
 wire _2994_;
 wire _2995_;
 wire _2996_;
 wire _2997_;
 wire _2998_;
 wire _2999_;
 wire _3000_;
 wire _3001_;
 wire _3002_;
 wire _3003_;
 wire _3004_;
 wire _3005_;
 wire _3006_;
 wire _3007_;
 wire _3008_;
 wire _3009_;
 wire _3010_;
 wire _3011_;
 wire _3012_;
 wire _3013_;
 wire _3014_;
 wire _3015_;
 wire _3016_;
 wire _3017_;
 wire _3018_;
 wire _3019_;
 wire _3020_;
 wire _3021_;
 wire _3022_;
 wire _3023_;
 wire _3024_;
 wire _3025_;
 wire _3026_;
 wire _3027_;
 wire _3028_;
 wire _3029_;
 wire _3030_;
 wire _3031_;
 wire _3032_;
 wire _3033_;
 wire _3034_;
 wire _3035_;
 wire _3036_;
 wire _3037_;
 wire _3038_;
 wire _3039_;
 wire _3040_;
 wire _3041_;
 wire _3042_;
 wire _3043_;
 wire _3044_;
 wire _3045_;
 wire _3046_;
 wire _3047_;
 wire _3048_;
 wire _3049_;
 wire _3050_;
 wire _3051_;
 wire _3052_;
 wire _3053_;
 wire _3054_;
 wire _3055_;
 wire _3056_;
 wire _3057_;
 wire _3058_;
 wire _3059_;
 wire _3060_;
 wire _3061_;
 wire _3062_;
 wire _3063_;
 wire _3064_;
 wire _3065_;
 wire _3066_;
 wire _3067_;
 wire _3068_;
 wire _3069_;
 wire _3070_;
 wire _3071_;
 wire _3072_;
 wire _3073_;
 wire _3074_;
 wire _3075_;
 wire _3076_;
 wire _3077_;
 wire _3078_;
 wire _3079_;
 wire _3080_;
 wire _3081_;
 wire _3082_;
 wire _3083_;
 wire _3084_;
 wire _3085_;
 wire _3086_;
 wire _3087_;
 wire _3088_;
 wire _3089_;
 wire _3090_;
 wire _3091_;
 wire _3092_;
 wire _3093_;
 wire _3094_;
 wire _3095_;
 wire _3096_;
 wire _3097_;
 wire _3098_;
 wire _3099_;
 wire _3100_;
 wire _3101_;
 wire _3102_;
 wire _3103_;
 wire _3104_;
 wire _3105_;
 wire _3106_;
 wire _3107_;
 wire _3108_;
 wire _3109_;
 wire _3110_;
 wire _3111_;
 wire _3112_;
 wire _3113_;
 wire _3114_;
 wire _3115_;
 wire _3116_;
 wire _3117_;
 wire _3118_;
 wire _3119_;
 wire _3120_;
 wire _3121_;
 wire _3122_;
 wire _3123_;
 wire _3124_;
 wire _3125_;
 wire _3126_;
 wire _3127_;
 wire _3128_;
 wire _3129_;
 wire _3130_;
 wire _3131_;
 wire _3132_;
 wire _3133_;
 wire _3134_;
 wire _3135_;
 wire _3136_;
 wire _3137_;
 wire _3138_;
 wire _3139_;
 wire _3140_;
 wire _3141_;
 wire _3142_;
 wire _3143_;
 wire _3144_;
 wire _3145_;
 wire _3146_;
 wire _3147_;
 wire _3148_;
 wire _3149_;
 wire _3150_;
 wire _3151_;
 wire _3152_;
 wire _3153_;
 wire _3154_;
 wire _3155_;
 wire _3156_;
 wire _3157_;
 wire _3158_;
 wire _3159_;
 wire _3160_;
 wire _3161_;
 wire _3162_;
 wire _3163_;
 wire _3164_;
 wire clknet_leaf_0_clk;
 wire net137;
 wire \btn.button_state[0] ;
 wire \btn.button_state[1] ;
 wire \btn.button_state[2] ;
 wire \btn.button_state[3] ;
 wire \btn.change_timer[0] ;
 wire \btn.change_timer[1] ;
 wire \btn.change_timer[2] ;
 wire \btn.change_timer[3] ;
 wire \btn.change_timer[4] ;
 wire \btn.change_timer[5] ;
 wire \btn.change_timer[6] ;
 wire \btn.current_event[0] ;
 wire \btn.current_event[1] ;
 wire \btn.current_event[2] ;
 wire \btn.current_event[3] ;
 wire \btn.gate_200hz ;
 wire \btn.input_event[0] ;
 wire \btn.input_event[1] ;
 wire \btn.input_event[2] ;
 wire \btn.input_event[3] ;
 wire \btn.input_event[4] ;
 wire \btn.long_press ;
 wire \btn.sample_10ms[0] ;
 wire \btn.sample_10ms[1] ;
 wire \btn.sample_10ms[2] ;
 wire \btn.sample_10ms[3] ;
 wire \btn.sample_15ms[0] ;
 wire \btn.sample_15ms[1] ;
 wire \btn.sample_15ms[2] ;
 wire \btn.sample_15ms[3] ;
 wire \btn.sample_5ms[0] ;
 wire \btn.sample_5ms[1] ;
 wire \btn.sample_5ms[2] ;
 wire \btn.sample_5ms[3] ;
 wire \clk_div_counter[0] ;
 wire \clk_div_counter[1] ;
 wire \clk_div_counter[2] ;
 wire \clk_div_counter[3] ;
 wire \clk_div_counter[4] ;
 wire \clk_div_counter[5] ;
 wire \clk_div_counter[6] ;
 wire \clk_div_counter[7] ;
 wire display_graphical;
 wire \display_value[0] ;
 wire \display_value[1] ;
 wire \display_value[2] ;
 wire \display_value[3] ;
 wire \display_value[4] ;
 wire \dsp.digit ;
 wire \dsp.digit_sel_raw[1] ;
 wire \dsp.segments_raw[0] ;
 wire \dsp.segments_raw[1] ;
 wire \dsp.segments_raw[2] ;
 wire \dsp.segments_raw[3] ;
 wire \dsp.segments_raw[4] ;
 wire \dsp.segments_raw[5] ;
 wire \dsp.segments_raw[6] ;
 wire \game.challenge_mode ;
 wire \game.challenge_num[0] ;
 wire \game.challenge_num[1] ;
 wire \game.challenge_num[2] ;
 wire \game.challenge_num[3] ;
 wire \game.counter[0] ;
 wire \game.counter[1] ;
 wire \game.counter[2] ;
 wire \game.counter[3] ;
 wire \game.counter[4] ;
 wire \game.counter[5] ;
 wire \game.counter[6] ;
 wire \game.counter[7] ;
 wire \game.current_level[0] ;
 wire \game.current_level[1] ;
 wire \game.current_level[2] ;
 wire \game.current_level[3] ;
 wire \game.current_level[4] ;
 wire \game.fsm.block_len[0][0] ;
 wire \game.fsm.block_len[0][1] ;
 wire \game.fsm.block_len[0][2] ;
 wire \game.fsm.block_len[1][0] ;
 wire \game.fsm.block_len[1][1] ;
 wire \game.fsm.block_len[1][2] ;
 wire \game.fsm.block_len[2][0] ;
 wire \game.fsm.block_len[2][1] ;
 wire \game.fsm.block_len[2][2] ;
 wire \game.fsm.block_len[3][0] ;
 wire \game.fsm.block_len[3][1] ;
 wire \game.fsm.block_len[3][2] ;
 wire \game.fsm.block_len[4][0] ;
 wire \game.fsm.block_len[4][1] ;
 wire \game.fsm.block_len[4][2] ;
 wire \game.fsm.block_len[5][0] ;
 wire \game.fsm.block_len[5][1] ;
 wire \game.fsm.block_len[5][2] ;
 wire \game.fsm.block_len[6][0] ;
 wire \game.fsm.block_len[6][1] ;
 wire \game.fsm.block_len[6][2] ;
 wire \game.fsm.block_len[7][0] ;
 wire \game.fsm.block_len[7][1] ;
 wire \game.fsm.block_len[7][2] ;
 wire \game.fsm.color_count[0][0] ;
 wire \game.fsm.color_count[0][1] ;
 wire \game.fsm.color_count[0][2] ;
 wire \game.fsm.color_count[1][0] ;
 wire \game.fsm.color_count[1][1] ;
 wire \game.fsm.color_count[1][2] ;
 wire \game.fsm.color_count[2][0] ;
 wire \game.fsm.color_count[2][1] ;
 wire \game.fsm.color_count[2][2] ;
 wire \game.fsm.color_count[3][0] ;
 wire \game.fsm.color_count[3][1] ;
 wire \game.fsm.color_count[3][2] ;
 wire \game.fsm.green_block_count[0] ;
 wire \game.fsm.green_block_count[1] ;
 wire \game.fsm.green_block_count[2] ;
 wire \game.fsm.len1_block_count[0] ;
 wire \game.fsm.len1_block_count[1] ;
 wire \game.fsm.len1_block_count[2] ;
 wire \game.fsm.len1_color_count[0][0] ;
 wire \game.fsm.len1_color_count[0][1] ;
 wire \game.fsm.len1_color_count[0][2] ;
 wire \game.fsm.len1_color_count[1][0] ;
 wire \game.fsm.len1_color_count[1][1] ;
 wire \game.fsm.len1_color_count[1][2] ;
 wire \game.fsm.len1_color_count[2][0] ;
 wire \game.fsm.len1_color_count[2][1] ;
 wire \game.fsm.len1_color_count[2][2] ;
 wire \game.fsm.len1_color_count[3][0] ;
 wire \game.fsm.len1_color_count[3][1] ;
 wire \game.fsm.len1_color_count[3][2] ;
 wire \game.fsm.len2_block_count[0] ;
 wire \game.fsm.len2_block_count[1] ;
 wire \game.fsm.len2_color_count[0][0] ;
 wire \game.fsm.len2_color_count[0][1] ;
 wire \game.fsm.len2_color_count[1][0] ;
 wire \game.fsm.len2_color_count[1][1] ;
 wire \game.fsm.len2_color_count[2][0] ;
 wire \game.fsm.len2_color_count[2][1] ;
 wire \game.fsm.len2_color_count[3][0] ;
 wire \game.fsm.len2_color_count[3][1] ;
 wire \game.fsm.len3_block_count[0] ;
 wire \game.fsm.len3_block_count[1] ;
 wire \game.fsm.len3_color_count[0][0] ;
 wire \game.fsm.len3_color_count[0][1] ;
 wire \game.fsm.len3_color_count[1][0] ;
 wire \game.fsm.len3_color_count[1][1] ;
 wire \game.fsm.len3_color_count[2][0] ;
 wire \game.fsm.len3_color_count[2][1] ;
 wire \game.fsm.len3_color_count[3][0] ;
 wire \game.fsm.len3_color_count[3][1] ;
 wire \game.fsm.length[0] ;
 wire \game.fsm.length[1] ;
 wire \game.fsm.length[2] ;
 wire \game.fsm.num_blocks[0] ;
 wire \game.fsm.num_blocks[1] ;
 wire \game.fsm.num_blocks[2] ;
 wire \game.fsm.read_pos[0] ;
 wire \game.fsm.read_pos[1] ;
 wire \game.fsm.read_pos[2] ;
 wire \game.fsm.seq[0][0] ;
 wire \game.fsm.seq[0][1] ;
 wire \game.fsm.seq[1][0] ;
 wire \game.fsm.seq[1][1] ;
 wire \game.fsm.seq[2][0] ;
 wire \game.fsm.seq[2][1] ;
 wire \game.fsm.seq[3][0] ;
 wire \game.fsm.seq[3][1] ;
 wire \game.fsm.seq[4][0] ;
 wire \game.fsm.seq[4][1] ;
 wire \game.fsm.seq[5][0] ;
 wire \game.fsm.seq[5][1] ;
 wire \game.fsm.seq[6][0] ;
 wire \game.fsm.seq[6][1] ;
 wire \game.fsm.seq[7][0] ;
 wire \game.fsm.seq[7][1] ;
 wire \game.input_color[0] ;
 wire \game.input_color[1] ;
 wire \game.input_erase ;
 wire \game.input_reset ;
 wire \game.input_update ;
 wire \game.next_state[0] ;
 wire \game.next_state[2] ;
 wire \game.slv.fsm_color[0] ;
 wire \game.slv.fsm_color[1] ;
 wire \game.slv.fsm_reset ;
 wire \game.slv.fsm_update ;
 wire \game.slv.length[0] ;
 wire \game.slv.length[1] ;
 wire \game.slv.length[2] ;
 wire \game.slv.lfsr[0] ;
 wire \game.slv.lfsr[10] ;
 wire \game.slv.lfsr[11] ;
 wire \game.slv.lfsr[12] ;
 wire \game.slv.lfsr[13] ;
 wire \game.slv.lfsr[14] ;
 wire \game.slv.lfsr[15] ;
 wire \game.slv.lfsr[16] ;
 wire \game.slv.lfsr[17] ;
 wire \game.slv.lfsr[18] ;
 wire \game.slv.lfsr[19] ;
 wire \game.slv.lfsr[1] ;
 wire \game.slv.lfsr[20] ;
 wire \game.slv.lfsr[2] ;
 wire \game.slv.lfsr[3] ;
 wire \game.slv.lfsr[4] ;
 wire \game.slv.lfsr[5] ;
 wire \game.slv.lfsr[6] ;
 wire \game.slv.lfsr[7] ;
 wire \game.slv.lfsr[8] ;
 wire \game.slv.lfsr[9] ;
 wire \game.slv.pos[0] ;
 wire \game.slv.pos[1] ;
 wire \game.slv.pos[2] ;
 wire \game.slv.ready ;
 wire \game.slv.retries[0] ;
 wire \game.slv.retries[1] ;
 wire \game.slv.retries[2] ;
 wire \game.slv.saved_target ;
 wire \game.slv.state[1] ;
 wire \game.slv.state[2] ;
 wire \game.slv.state[3] ;
 wire \game.slv.target[0] ;
 wire \game.slv.target[1] ;
 wire \game.slv.trigger ;
 wire \game.solver_active ;
 wire \game.solver_trigger_delayed ;
 wire \game.sound_mode[0] ;
 wire \game.sound_mode[1] ;
 wire \game.sound_mode[2] ;
 wire \game.sound_on ;
 wire \game.state[0] ;
 wire \game.state[1] ;
 wire \game.state[2] ;
 wire \game.state[3] ;
 wire \game.tune[0] ;
 wire \game.tune[1] ;
 wire \snd.active_tune[0] ;
 wire \snd.active_tune[1] ;
 wire \snd.chord[0][0] ;
 wire \snd.chord[0][1] ;
 wire \snd.chord[0][2] ;
 wire \snd.chord[0][3] ;
 wire \snd.chord[0][4] ;
 wire \snd.chord[0][5] ;
 wire \snd.chord[1][0] ;
 wire \snd.chord[1][5] ;
 wire \snd.chord[2][2] ;
 wire \snd.chord[3][0] ;
 wire \snd.counter[0] ;
 wire \snd.counter[1] ;
 wire \snd.counter[2] ;
 wire \snd.counter[3] ;
 wire \snd.counter[4] ;
 wire \snd.counter[5] ;
 wire \snd.counter[6] ;
 wire \snd.counter[7] ;
 wire \snd.counter[8] ;
 wire \snd.next_note_sel[0] ;
 wire \snd.next_note_sel[1] ;
 wire \snd.next_note_timing[0] ;
 wire \snd.next_note_timing[1] ;
 wire \snd.next_note_timing[2] ;
 wire \snd.next_note_timing[3] ;
 wire \snd.next_note_timing[4] ;
 wire \snd.next_note_timing[5] ;
 wire \snd.next_note_timing[6] ;
 wire \snd.next_note_timing[7] ;
 wire \snd.next_note_timing[8] ;
 wire \snd.note_sel[0] ;
 wire \snd.note_sel[1] ;
 wire \snd.note_timing[0] ;
 wire \snd.note_timing[1] ;
 wire \snd.note_timing[2] ;
 wire \snd.note_timing[3] ;
 wire \snd.note_timing[4] ;
 wire \snd.note_timing[5] ;
 wire \snd.note_timing[6] ;
 wire \snd.note_timing[7] ;
 wire \snd.note_timing[8] ;
 wire \snd.sequencer_state[0] ;
 wire \snd.sequencer_state[1] ;
 wire \snd.sound ;
 wire \snd.tune_counter[0] ;
 wire \snd.tune_counter[1] ;
 wire \snd.tune_counter[2] ;
 wire \snd.tune_counter[3] ;
 wire \snd.tune_counter[4] ;
 wire \snd.tune_counter[5] ;
 wire \snd.tune_counter[6] ;
 wire \snd.tune_pos[0] ;
 wire \snd.tune_pos[1] ;
 wire \snd.tune_pos[2] ;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net138;
 wire net139;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net180;
 wire net181;
 wire net182;
 wire net183;
 wire net184;
 wire net185;
 wire net186;
 wire net187;
 wire net188;
 wire net189;
 wire net190;
 wire net191;
 wire net192;
 wire net193;
 wire net194;
 wire net195;
 wire net196;
 wire net197;
 wire net198;
 wire net199;
 wire net200;
 wire net201;
 wire net202;
 wire net203;
 wire net204;
 wire net205;
 wire net206;
 wire net207;
 wire net208;
 wire net209;
 wire net210;
 wire net211;
 wire net212;
 wire net213;
 wire net214;
 wire net215;
 wire net216;
 wire net217;
 wire net218;
 wire net219;
 wire net220;
 wire net221;
 wire net222;
 wire net223;
 wire net224;
 wire net225;
 wire net226;
 wire net227;
 wire net228;
 wire net229;
 wire net230;
 wire net231;
 wire net232;
 wire net233;
 wire net234;
 wire net235;
 wire net236;
 wire net237;
 wire net238;
 wire net239;
 wire net240;
 wire net241;
 wire net242;
 wire net243;
 wire net244;
 wire net245;
 wire net246;
 wire net247;
 wire net248;
 wire net249;
 wire net250;
 wire net251;
 wire net252;
 wire net253;
 wire net254;
 wire net255;
 wire net256;
 wire net257;
 wire net258;
 wire net259;
 wire net260;
 wire net261;
 wire net262;
 wire net263;
 wire net264;
 wire net265;
 wire net266;
 wire net267;
 wire net268;
 wire net269;
 wire net270;
 wire net271;
 wire net272;
 wire net273;
 wire net274;
 wire net275;
 wire net276;
 wire net277;
 wire net278;
 wire net279;
 wire net280;
 wire net281;
 wire net282;
 wire net283;
 wire net284;
 wire net285;
 wire net286;
 wire net287;
 wire net288;
 wire net289;
 wire net290;
 wire net291;
 wire net292;
 wire net293;
 wire net294;
 wire net295;
 wire net296;
 wire net297;
 wire net298;
 wire net299;
 wire net300;
 wire net301;
 wire net302;
 wire net303;
 wire net304;
 wire net305;
 wire net306;
 wire net307;
 wire net308;
 wire net309;
 wire net310;
 wire net311;
 wire net312;
 wire net313;
 wire net314;
 wire net315;
 wire net316;
 wire net317;
 wire net318;
 wire net319;
 wire net320;
 wire net321;
 wire net322;
 wire net323;
 wire net324;
 wire net325;
 wire net326;
 wire net327;
 wire net328;
 wire net329;
 wire net330;
 wire net331;
 wire net332;
 wire net333;
 wire net334;
 wire net335;
 wire net336;
 wire net337;
 wire net338;
 wire net339;
 wire net340;
 wire net341;
 wire net342;
 wire net343;
 wire net344;
 wire net345;
 wire net346;
 wire net347;
 wire net348;
 wire net349;
 wire net350;
 wire net351;
 wire net352;
 wire net353;
 wire net354;
 wire net355;
 wire net356;
 wire net357;
 wire net358;
 wire net359;
 wire net360;
 wire net361;
 wire net362;
 wire net363;
 wire net364;
 wire net365;
 wire net366;
 wire net367;
 wire net368;
 wire net369;
 wire net370;
 wire net371;
 wire net372;
 wire net373;
 wire net374;
 wire net375;
 wire net376;
 wire net377;
 wire net378;
 wire net379;
 wire net380;
 wire net381;
 wire net382;
 wire net383;
 wire net384;
 wire net385;
 wire net386;
 wire net387;
 wire net388;
 wire net389;
 wire net390;
 wire net391;
 wire net392;
 wire net393;
 wire net394;
 wire net395;
 wire net396;
 wire net397;
 wire net398;
 wire net399;
 wire net400;
 wire net401;
 wire net402;
 wire net403;
 wire net404;
 wire net405;
 wire net406;
 wire net407;
 wire net408;
 wire net409;
 wire net410;
 wire net411;
 wire net412;
 wire net413;
 wire net414;
 wire net415;
 wire net416;
 wire net417;
 wire net418;
 wire net419;
 wire net420;
 wire net421;
 wire net422;
 wire net423;
 wire net424;
 wire net425;
 wire net426;
 wire net427;
 wire net428;
 wire net429;
 wire net430;
 wire net431;
 wire net432;
 wire net433;
 wire net434;
 wire net435;
 wire net436;
 wire net437;
 wire net438;
 wire net439;
 wire net440;
 wire net441;
 wire net442;
 wire net443;
 wire net444;
 wire net445;
 wire net446;
 wire net447;
 wire net448;
 wire net449;
 wire clknet_leaf_1_clk;
 wire clknet_leaf_2_clk;
 wire clknet_leaf_3_clk;
 wire clknet_leaf_4_clk;
 wire clknet_leaf_6_clk;
 wire clknet_leaf_7_clk;
 wire clknet_leaf_8_clk;
 wire clknet_leaf_9_clk;
 wire clknet_leaf_10_clk;
 wire clknet_leaf_11_clk;
 wire clknet_leaf_12_clk;
 wire clknet_leaf_13_clk;
 wire clknet_leaf_14_clk;
 wire clknet_leaf_15_clk;
 wire clknet_leaf_16_clk;
 wire clknet_leaf_17_clk;
 wire clknet_leaf_18_clk;
 wire clknet_leaf_19_clk;
 wire clknet_leaf_20_clk;
 wire clknet_leaf_21_clk;
 wire clknet_leaf_22_clk;
 wire clknet_leaf_23_clk;
 wire clknet_leaf_24_clk;
 wire clknet_leaf_25_clk;
 wire clknet_leaf_26_clk;
 wire clknet_leaf_27_clk;
 wire clknet_leaf_28_clk;
 wire clknet_leaf_29_clk;
 wire clknet_leaf_30_clk;
 wire clknet_leaf_31_clk;
 wire clknet_leaf_32_clk;
 wire clknet_leaf_34_clk;
 wire clknet_leaf_35_clk;
 wire clknet_leaf_36_clk;
 wire clknet_leaf_37_clk;
 wire clknet_leaf_38_clk;
 wire clknet_leaf_39_clk;
 wire clknet_leaf_40_clk;
 wire clknet_leaf_41_clk;
 wire clknet_leaf_42_clk;
 wire clknet_leaf_43_clk;
 wire clknet_leaf_44_clk;
 wire clknet_leaf_45_clk;
 wire clknet_0_clk;
 wire clknet_3_0__leaf_clk;
 wire clknet_3_1__leaf_clk;
 wire clknet_3_2__leaf_clk;
 wire clknet_3_3__leaf_clk;
 wire clknet_3_4__leaf_clk;
 wire clknet_3_5__leaf_clk;
 wire clknet_3_6__leaf_clk;
 wire clknet_3_7__leaf_clk;
 wire net450;

 sg13g2_inv_1 _3167_ (.Y(_2632_),
    .A(\game.slv.trigger ));
 sg13g2_buf_1 _3168_ (.A(\game.slv.lfsr[2] ),
    .X(_2633_));
 sg13g2_buf_1 _3169_ (.A(\game.slv.lfsr[1] ),
    .X(_2634_));
 sg13g2_buf_2 _3170_ (.A(\game.slv.lfsr[0] ),
    .X(_2635_));
 sg13g2_and3_1 _3171_ (.X(_2636_),
    .A(_2633_),
    .B(_2634_),
    .C(_2635_));
 sg13g2_nor3_1 _3172_ (.A(_2633_),
    .B(_2634_),
    .C(_2635_),
    .Y(_2637_));
 sg13g2_buf_2 _3173_ (.A(\game.slv.state[2] ),
    .X(_2638_));
 sg13g2_o21ai_1 _3174_ (.B1(_2638_),
    .Y(_2639_),
    .A1(_2636_),
    .A2(_2637_));
 sg13g2_buf_1 _3175_ (.A(rst_n),
    .X(_2640_));
 sg13g2_inv_2 _3176_ (.Y(_2641_),
    .A(_2640_));
 sg13g2_buf_1 _3177_ (.A(_2641_),
    .X(_2642_));
 sg13g2_buf_1 _3178_ (.A(net108),
    .X(_2643_));
 sg13g2_a21oi_1 _3179_ (.A1(_2632_),
    .A2(_2639_),
    .Y(_0012_),
    .B1(net73));
 sg13g2_buf_1 _3180_ (.A(_2640_),
    .X(_2644_));
 sg13g2_nand2_1 _3181_ (.Y(_2645_),
    .A(net134),
    .B(_2632_));
 sg13g2_buf_2 _3182_ (.A(\game.fsm.block_len[6][1] ),
    .X(_2646_));
 sg13g2_inv_1 _3183_ (.Y(_2647_),
    .A(_2646_));
 sg13g2_buf_1 _3184_ (.A(_0078_),
    .X(_2648_));
 sg13g2_buf_2 _3185_ (.A(_0077_),
    .X(_2649_));
 sg13g2_buf_8 _3186_ (.A(\game.fsm.block_len[4][0] ),
    .X(_2650_));
 sg13g2_inv_1 _3187_ (.Y(_2651_),
    .A(_2650_));
 sg13g2_buf_1 _3188_ (.A(\game.fsm.block_len[4][2] ),
    .X(_2652_));
 sg13g2_buf_8 _3189_ (.A(\game.fsm.block_len[5][2] ),
    .X(_2653_));
 sg13g2_nor2b_1 _3190_ (.A(net133),
    .B_N(_2653_),
    .Y(_2654_));
 sg13g2_buf_8 _3191_ (.A(\game.fsm.block_len[4][1] ),
    .X(_2655_));
 sg13g2_buf_8 _3192_ (.A(\game.fsm.block_len[5][1] ),
    .X(_2656_));
 sg13g2_nor2b_1 _3193_ (.A(_2655_),
    .B_N(_2656_),
    .Y(_2657_));
 sg13g2_or4_1 _3194_ (.A(_2651_),
    .B(\game.fsm.block_len[5][0] ),
    .C(_2654_),
    .D(_2657_),
    .X(_2658_));
 sg13g2_buf_1 _3195_ (.A(_2658_),
    .X(_2659_));
 sg13g2_nand2b_1 _3196_ (.Y(_2660_),
    .B(_2653_),
    .A_N(net133));
 sg13g2_nor2b_1 _3197_ (.A(_2656_),
    .B_N(_2655_),
    .Y(_2661_));
 sg13g2_nor2b_1 _3198_ (.A(_2653_),
    .B_N(net133),
    .Y(_2662_));
 sg13g2_a21oi_1 _3199_ (.A1(_2660_),
    .A2(_2661_),
    .Y(_2663_),
    .B1(_2662_));
 sg13g2_inv_1 _3200_ (.Y(_2664_),
    .A(\game.fsm.num_blocks[2] ));
 sg13g2_buf_2 _3201_ (.A(\game.fsm.num_blocks[1] ),
    .X(_2665_));
 sg13g2_inv_4 _3202_ (.A(_2665_),
    .Y(_2666_));
 sg13g2_nor2_2 _3203_ (.A(_2664_),
    .B(_2666_),
    .Y(_2667_));
 sg13g2_nand2b_1 _3204_ (.Y(_2668_),
    .B(net133),
    .A_N(_2653_));
 sg13g2_xnor2_1 _3205_ (.Y(_2669_),
    .A(_2650_),
    .B(\game.fsm.block_len[5][0] ));
 sg13g2_xnor2_1 _3206_ (.Y(_2670_),
    .A(_2655_),
    .B(_2656_));
 sg13g2_nand4_1 _3207_ (.B(_2668_),
    .C(_2669_),
    .A(_2660_),
    .Y(_2671_),
    .D(_2670_));
 sg13g2_and4_1 _3208_ (.A(_2659_),
    .B(_2663_),
    .C(_2667_),
    .D(_2671_),
    .X(_2672_));
 sg13g2_buf_8 _3209_ (.A(_2672_),
    .X(_2673_));
 sg13g2_mux2_1 _3210_ (.A0(_2648_),
    .A1(_2649_),
    .S(net42),
    .X(_2674_));
 sg13g2_buf_8 _3211_ (.A(_2674_),
    .X(_2675_));
 sg13g2_xnor2_1 _3212_ (.Y(_2676_),
    .A(_2647_),
    .B(_2675_));
 sg13g2_buf_1 _3213_ (.A(_0079_),
    .X(_2677_));
 sg13g2_buf_1 _3214_ (.A(_0081_),
    .X(_2678_));
 sg13g2_buf_1 _3215_ (.A(_0080_),
    .X(_2679_));
 sg13g2_mux2_1 _3216_ (.A0(_2678_),
    .A1(_2679_),
    .S(net42),
    .X(_2680_));
 sg13g2_buf_8 _3217_ (.A(_2680_),
    .X(_2681_));
 sg13g2_xnor2_1 _3218_ (.Y(_2682_),
    .A(_2677_),
    .B(_2681_));
 sg13g2_buf_2 _3219_ (.A(_2682_),
    .X(_2683_));
 sg13g2_mux2_1 _3220_ (.A0(_0076_),
    .A1(_0075_),
    .S(net42),
    .X(_2684_));
 sg13g2_buf_2 _3221_ (.A(_2684_),
    .X(_2685_));
 sg13g2_buf_1 _3222_ (.A(_0074_),
    .X(_2686_));
 sg13g2_buf_1 _3223_ (.A(\game.fsm.num_blocks[0] ),
    .X(_2687_));
 sg13g2_buf_2 _3224_ (.A(_2687_),
    .X(_2688_));
 sg13g2_nand2_2 _3225_ (.Y(_2689_),
    .A(_2688_),
    .B(_2667_));
 sg13g2_nor2_1 _3226_ (.A(net132),
    .B(_2689_),
    .Y(_2690_));
 sg13g2_and4_1 _3227_ (.A(_2676_),
    .B(_2683_),
    .C(_2685_),
    .D(_2690_),
    .X(_2691_));
 sg13g2_buf_2 _3228_ (.A(_2691_),
    .X(_2692_));
 sg13g2_nand2_1 _3229_ (.Y(_2693_),
    .A(_2649_),
    .B(net42));
 sg13g2_nand2b_1 _3230_ (.Y(_2694_),
    .B(_2648_),
    .A_N(net42));
 sg13g2_inv_1 _3231_ (.Y(_2695_),
    .A(_0076_));
 sg13g2_nand2_1 _3232_ (.Y(_2696_),
    .A(_2695_),
    .B(net132));
 sg13g2_inv_1 _3233_ (.Y(_2697_),
    .A(_0075_));
 sg13g2_nand2_1 _3234_ (.Y(_2698_),
    .A(_2697_),
    .B(net132));
 sg13g2_mux2_1 _3235_ (.A0(_2696_),
    .A1(_2698_),
    .S(net42),
    .X(_2699_));
 sg13g2_buf_1 _3236_ (.A(_0082_),
    .X(_2700_));
 sg13g2_inv_1 _3237_ (.Y(_2701_),
    .A(net131));
 sg13g2_and2_1 _3238_ (.A(_2687_),
    .B(_2667_),
    .X(_2702_));
 sg13g2_buf_1 _3239_ (.A(_2702_),
    .X(_2703_));
 sg13g2_nand2_1 _3240_ (.Y(_2704_),
    .A(_2701_),
    .B(_2703_));
 sg13g2_a221oi_1 _3241_ (.B2(_2647_),
    .C1(_2704_),
    .B1(_2699_),
    .A1(_2693_),
    .Y(_2705_),
    .A2(_2694_));
 sg13g2_a21oi_1 _3242_ (.A1(_2653_),
    .A2(_2667_),
    .Y(_2706_),
    .B1(_2652_));
 sg13g2_a21o_1 _3243_ (.A2(_2705_),
    .A1(_2683_),
    .B1(_2706_),
    .X(_2707_));
 sg13g2_buf_1 _3244_ (.A(_2707_),
    .X(_2708_));
 sg13g2_buf_2 _3245_ (.A(\game.fsm.block_len[1][2] ),
    .X(_2709_));
 sg13g2_nor2b_1 _3246_ (.A(_2709_),
    .B_N(\game.fsm.block_len[0][2] ),
    .Y(_2710_));
 sg13g2_inv_1 _3247_ (.Y(_2711_),
    .A(\game.fsm.block_len[0][2] ));
 sg13g2_buf_2 _3248_ (.A(\game.fsm.block_len[1][1] ),
    .X(_2712_));
 sg13g2_nand2b_1 _3249_ (.Y(_2713_),
    .B(\game.fsm.block_len[0][1] ),
    .A_N(_2712_));
 sg13g2_nor2b_1 _3250_ (.A(\game.fsm.block_len[0][0] ),
    .B_N(\game.fsm.block_len[1][0] ),
    .Y(_2714_));
 sg13g2_nor2b_1 _3251_ (.A(\game.fsm.block_len[0][1] ),
    .B_N(_2712_),
    .Y(_2715_));
 sg13g2_a221oi_1 _3252_ (.B2(_2714_),
    .C1(_2715_),
    .B1(_2713_),
    .A1(_2711_),
    .Y(_2716_),
    .A2(_2709_));
 sg13g2_nor2_1 _3253_ (.A(\game.fsm.num_blocks[2] ),
    .B(_2665_),
    .Y(_2717_));
 sg13g2_nor3_2 _3254_ (.A(_2710_),
    .B(_2716_),
    .C(_2717_),
    .Y(_2718_));
 sg13g2_mux2_1 _3255_ (.A0(_0089_),
    .A1(_0088_),
    .S(_2718_),
    .X(_2719_));
 sg13g2_buf_2 _3256_ (.A(_2719_),
    .X(_2720_));
 sg13g2_buf_2 _3257_ (.A(\game.fsm.block_len[3][2] ),
    .X(_2721_));
 sg13g2_buf_2 _3258_ (.A(_0085_),
    .X(_2722_));
 sg13g2_nand3_1 _3259_ (.B(_2665_),
    .C(_2722_),
    .A(_2687_),
    .Y(_2723_));
 sg13g2_buf_2 _3260_ (.A(\game.fsm.block_len[2][2] ),
    .X(_2724_));
 sg13g2_a21oi_1 _3261_ (.A1(_2721_),
    .A2(_2723_),
    .Y(_2725_),
    .B1(_2724_));
 sg13g2_buf_1 _3262_ (.A(_2665_),
    .X(_2726_));
 sg13g2_and2_1 _3263_ (.A(net107),
    .B(net106),
    .X(_2727_));
 sg13g2_buf_1 _3264_ (.A(\game.fsm.num_blocks[2] ),
    .X(_2728_));
 sg13g2_a21oi_1 _3265_ (.A1(_2724_),
    .A2(_2727_),
    .Y(_2729_),
    .B1(net130));
 sg13g2_or2_1 _3266_ (.X(_2730_),
    .B(_2729_),
    .A(_2725_));
 sg13g2_nand2_1 _3267_ (.Y(_2731_),
    .A(_2720_),
    .B(_2730_));
 sg13g2_buf_2 _3268_ (.A(_2731_),
    .X(_2732_));
 sg13g2_inv_1 _3269_ (.Y(_2733_),
    .A(_0023_));
 sg13g2_nor3_2 _3270_ (.A(\game.fsm.len1_color_count[1][1] ),
    .B(\game.fsm.len1_color_count[1][0] ),
    .C(_2733_),
    .Y(_2734_));
 sg13g2_inv_1 _3271_ (.Y(_2735_),
    .A(_0022_));
 sg13g2_nor3_2 _3272_ (.A(\game.fsm.len1_color_count[0][1] ),
    .B(\game.fsm.len1_color_count[0][0] ),
    .C(_2735_),
    .Y(_2736_));
 sg13g2_inv_1 _3273_ (.Y(_2737_),
    .A(_0024_));
 sg13g2_nor3_1 _3274_ (.A(\game.fsm.len1_color_count[3][1] ),
    .B(\game.fsm.len1_color_count[3][0] ),
    .C(_2737_),
    .Y(_2738_));
 sg13g2_xnor2_1 _3275_ (.Y(_2739_),
    .A(_2736_),
    .B(_2738_));
 sg13g2_xnor2_1 _3276_ (.Y(_2740_),
    .A(_2734_),
    .B(_2739_));
 sg13g2_buf_2 _3277_ (.A(_2740_),
    .X(_2741_));
 sg13g2_nor2_1 _3278_ (.A(\game.fsm.len3_color_count[1][1] ),
    .B(\game.fsm.len3_color_count[1][0] ),
    .Y(_2742_));
 sg13g2_nor2_1 _3279_ (.A(\game.fsm.len2_color_count[3][1] ),
    .B(\game.fsm.len2_color_count[3][0] ),
    .Y(_2743_));
 sg13g2_nor2_1 _3280_ (.A(\game.fsm.len2_color_count[1][1] ),
    .B(\game.fsm.len2_color_count[1][0] ),
    .Y(_2744_));
 sg13g2_xor2_1 _3281_ (.B(_2744_),
    .A(_2743_),
    .X(_2745_));
 sg13g2_xnor2_1 _3282_ (.Y(_2746_),
    .A(_2742_),
    .B(_2745_));
 sg13g2_nor2_1 _3283_ (.A(\game.fsm.len3_color_count[2][1] ),
    .B(\game.fsm.len3_color_count[2][0] ),
    .Y(_2747_));
 sg13g2_nor2_1 _3284_ (.A(\game.fsm.len3_color_count[0][1] ),
    .B(\game.fsm.len3_color_count[0][0] ),
    .Y(_2748_));
 sg13g2_xor2_1 _3285_ (.B(_2748_),
    .A(_2747_),
    .X(_2749_));
 sg13g2_xnor2_1 _3286_ (.Y(_2750_),
    .A(_2746_),
    .B(_2749_));
 sg13g2_xnor2_1 _3287_ (.Y(_2751_),
    .A(_2741_),
    .B(_2750_));
 sg13g2_nor2_2 _3288_ (.A(\game.fsm.len2_color_count[2][1] ),
    .B(\game.fsm.len2_color_count[2][0] ),
    .Y(_2752_));
 sg13g2_nor2_2 _3289_ (.A(\game.fsm.len3_color_count[3][1] ),
    .B(\game.fsm.len3_color_count[3][0] ),
    .Y(_2753_));
 sg13g2_xnor2_1 _3290_ (.Y(_2754_),
    .A(_2752_),
    .B(_2753_));
 sg13g2_nor3_1 _3291_ (.A(_2732_),
    .B(_2751_),
    .C(_2754_),
    .Y(_2755_));
 sg13g2_o21ai_1 _3292_ (.B1(_2755_),
    .Y(_2756_),
    .A1(_2692_),
    .A2(_2708_));
 sg13g2_nand2b_1 _3293_ (.Y(_2757_),
    .B(_0073_),
    .A_N(net107));
 sg13g2_and2_1 _3294_ (.A(net130),
    .B(_2757_),
    .X(_2758_));
 sg13g2_buf_1 _3295_ (.A(_2758_),
    .X(_2759_));
 sg13g2_xor2_1 _3296_ (.B(_2753_),
    .A(_2752_),
    .X(_2760_));
 sg13g2_nand3_1 _3297_ (.B(_2751_),
    .C(_2760_),
    .A(_2759_),
    .Y(_2761_));
 sg13g2_xnor2_1 _3298_ (.Y(_2762_),
    .A(net132),
    .B(_2685_));
 sg13g2_and3_1 _3299_ (.X(_2763_),
    .A(_2676_),
    .B(_2683_),
    .C(_2762_));
 sg13g2_buf_2 _3300_ (.A(\game.fsm.block_len[6][2] ),
    .X(_2764_));
 sg13g2_nand2_1 _3301_ (.Y(_2765_),
    .A(_2764_),
    .B(_2703_));
 sg13g2_and2_1 _3302_ (.A(_2681_),
    .B(_2699_),
    .X(_2766_));
 sg13g2_nand2_1 _3303_ (.Y(_2767_),
    .A(_2648_),
    .B(_2678_));
 sg13g2_nand2_1 _3304_ (.Y(_2768_),
    .A(_2649_),
    .B(_2679_));
 sg13g2_mux2_1 _3305_ (.A0(_2767_),
    .A1(_2768_),
    .S(_2673_),
    .X(_2769_));
 sg13g2_o21ai_1 _3306_ (.B1(_2677_),
    .Y(_2770_),
    .A1(_2700_),
    .A2(_2769_));
 sg13g2_a21oi_1 _3307_ (.A1(_2676_),
    .A2(_2766_),
    .Y(_2771_),
    .B1(_2770_));
 sg13g2_nor3_2 _3308_ (.A(_2763_),
    .B(_2765_),
    .C(_2771_),
    .Y(_2772_));
 sg13g2_mux2_1 _3309_ (.A0(_2756_),
    .A1(_2761_),
    .S(_2772_),
    .X(_2773_));
 sg13g2_xor2_1 _3310_ (.B(_2750_),
    .A(_2741_),
    .X(_2774_));
 sg13g2_nor3_1 _3311_ (.A(_2732_),
    .B(_2774_),
    .C(_2760_),
    .Y(_2775_));
 sg13g2_o21ai_1 _3312_ (.B1(_2775_),
    .Y(_2776_),
    .A1(_2692_),
    .A2(_2708_));
 sg13g2_nand3_1 _3313_ (.B(_2774_),
    .C(_2754_),
    .A(_2759_),
    .Y(_2777_));
 sg13g2_mux2_1 _3314_ (.A0(_2776_),
    .A1(_2777_),
    .S(_2772_),
    .X(_2778_));
 sg13g2_nor3_1 _3315_ (.A(_2692_),
    .B(_2708_),
    .C(_2761_),
    .Y(_2779_));
 sg13g2_nor3_1 _3316_ (.A(_2692_),
    .B(_2708_),
    .C(_2777_),
    .Y(_2780_));
 sg13g2_nand3_1 _3317_ (.B(_2751_),
    .C(_2760_),
    .A(_2732_),
    .Y(_2781_));
 sg13g2_nand2_1 _3318_ (.Y(_2782_),
    .A(_2728_),
    .B(_2757_));
 sg13g2_buf_2 _3319_ (.A(_2782_),
    .X(_2783_));
 sg13g2_and2_1 _3320_ (.A(_2720_),
    .B(_2730_),
    .X(_2784_));
 sg13g2_buf_1 _3321_ (.A(_2784_),
    .X(_2785_));
 sg13g2_nand4_1 _3322_ (.B(_2785_),
    .C(_2774_),
    .A(_2783_),
    .Y(_2786_),
    .D(_2760_));
 sg13g2_nand3_1 _3323_ (.B(_2774_),
    .C(_2754_),
    .A(_2732_),
    .Y(_2787_));
 sg13g2_nand4_1 _3324_ (.B(_2785_),
    .C(_2751_),
    .A(_2783_),
    .Y(_2788_),
    .D(_2754_));
 sg13g2_nand4_1 _3325_ (.B(_2786_),
    .C(_2787_),
    .A(_2781_),
    .Y(_2789_),
    .D(_2788_));
 sg13g2_nor3_1 _3326_ (.A(_2779_),
    .B(_2780_),
    .C(_2789_),
    .Y(_2790_));
 sg13g2_nand3_1 _3327_ (.B(_2778_),
    .C(_2790_),
    .A(_2773_),
    .Y(_2791_));
 sg13g2_nor2_1 _3328_ (.A(\game.fsm.len1_color_count[2][1] ),
    .B(\game.fsm.len1_color_count[2][0] ),
    .Y(_2792_));
 sg13g2_nand2_1 _3329_ (.Y(_2793_),
    .A(_0025_),
    .B(_2792_));
 sg13g2_inv_1 _3330_ (.Y(_2794_),
    .A(\game.current_level[0] ));
 sg13g2_buf_1 _3331_ (.A(_2794_),
    .X(_2795_));
 sg13g2_or3_1 _3332_ (.A(net105),
    .B(\game.fsm.len2_color_count[0][1] ),
    .C(\game.fsm.len2_color_count[0][0] ),
    .X(_2796_));
 sg13g2_nor3_1 _3333_ (.A(_2791_),
    .B(_2793_),
    .C(_2796_),
    .Y(_2797_));
 sg13g2_and2_1 _3334_ (.A(_0025_),
    .B(_2792_),
    .X(_2798_));
 sg13g2_nor2_1 _3335_ (.A(_2798_),
    .B(_2796_),
    .Y(_2799_));
 sg13g2_buf_1 _3336_ (.A(\game.current_level[0] ),
    .X(_2800_));
 sg13g2_o21ai_1 _3337_ (.B1(net129),
    .Y(_2801_),
    .A1(\game.fsm.len2_color_count[0][1] ),
    .A2(\game.fsm.len2_color_count[0][0] ));
 sg13g2_nor2_1 _3338_ (.A(_2793_),
    .B(_2801_),
    .Y(_2802_));
 sg13g2_o21ai_1 _3339_ (.B1(_2791_),
    .Y(_2803_),
    .A1(_2799_),
    .A2(_2802_));
 sg13g2_nor2b_1 _3340_ (.A(_2797_),
    .B_N(_2803_),
    .Y(_2804_));
 sg13g2_or3_1 _3341_ (.A(_2791_),
    .B(_2798_),
    .C(_2801_),
    .X(_2805_));
 sg13g2_nor3_1 _3342_ (.A(_2783_),
    .B(_2692_),
    .C(_2708_),
    .Y(_2806_));
 sg13g2_or3_1 _3343_ (.A(_2763_),
    .B(_2765_),
    .C(_2771_),
    .X(_2807_));
 sg13g2_buf_8 _3344_ (.A(_2807_),
    .X(_2808_));
 sg13g2_nand3b_1 _3345_ (.B(_2785_),
    .C(_2808_),
    .Y(_2809_),
    .A_N(_2806_));
 sg13g2_nor2_1 _3346_ (.A(_2747_),
    .B(_2748_),
    .Y(_2810_));
 sg13g2_nand2_1 _3347_ (.Y(_2811_),
    .A(_2747_),
    .B(_2748_));
 sg13g2_o21ai_1 _3348_ (.B1(_2811_),
    .Y(_2812_),
    .A1(_2746_),
    .A2(_2810_));
 sg13g2_nand2_1 _3349_ (.Y(_2813_),
    .A(_2746_),
    .B(_2810_));
 sg13g2_o21ai_1 _3350_ (.B1(_2813_),
    .Y(_2814_),
    .A1(_2741_),
    .A2(_2812_));
 sg13g2_nor2_1 _3351_ (.A(_2746_),
    .B(_2811_),
    .Y(_2815_));
 sg13g2_a21oi_1 _3352_ (.A1(_2741_),
    .A2(_2812_),
    .Y(_2816_),
    .B1(_2815_));
 sg13g2_nor2_1 _3353_ (.A(_2732_),
    .B(_2816_),
    .Y(_2817_));
 sg13g2_nor2_1 _3354_ (.A(_2772_),
    .B(_2806_),
    .Y(_2818_));
 sg13g2_nand2_1 _3355_ (.Y(_2819_),
    .A(_2741_),
    .B(_2815_));
 sg13g2_o21ai_1 _3356_ (.B1(_2819_),
    .Y(_2820_),
    .A1(_2741_),
    .A2(_2813_));
 sg13g2_a221oi_1 _3357_ (.B2(_2818_),
    .C1(_2820_),
    .B1(_2817_),
    .A1(_2809_),
    .Y(_2821_),
    .A2(_2814_));
 sg13g2_a21o_1 _3358_ (.A2(_2736_),
    .A1(_2734_),
    .B1(_2738_),
    .X(_2822_));
 sg13g2_o21ai_1 _3359_ (.B1(_2822_),
    .Y(_2823_),
    .A1(_2734_),
    .A2(_2736_));
 sg13g2_nor2_1 _3360_ (.A(_2742_),
    .B(_2743_),
    .Y(_2824_));
 sg13g2_a21oi_1 _3361_ (.A1(_2742_),
    .A2(_2743_),
    .Y(_2825_),
    .B1(_2744_));
 sg13g2_or2_1 _3362_ (.X(_2826_),
    .B(_2825_),
    .A(_2824_));
 sg13g2_xnor2_1 _3363_ (.Y(_2827_),
    .A(_2823_),
    .B(_2826_));
 sg13g2_xnor2_1 _3364_ (.Y(_2828_),
    .A(_2821_),
    .B(_2827_));
 sg13g2_nand2_1 _3365_ (.Y(_2829_),
    .A(_2752_),
    .B(_2753_));
 sg13g2_nand2_1 _3366_ (.Y(_2830_),
    .A(_2751_),
    .B(_2829_));
 sg13g2_nand2_1 _3367_ (.Y(_2831_),
    .A(_2774_),
    .B(_2829_));
 sg13g2_nor3_1 _3368_ (.A(_2732_),
    .B(_2772_),
    .C(_2806_),
    .Y(_2832_));
 sg13g2_mux2_1 _3369_ (.A0(_2830_),
    .A1(_2831_),
    .S(_2832_),
    .X(_2833_));
 sg13g2_o21ai_1 _3370_ (.B1(_2833_),
    .Y(_2834_),
    .A1(_2752_),
    .A2(_2753_));
 sg13g2_xnor2_1 _3371_ (.Y(_2835_),
    .A(_2828_),
    .B(_2834_));
 sg13g2_mux2_1 _3372_ (.A0(_2804_),
    .A1(_2805_),
    .S(_2835_),
    .X(_2836_));
 sg13g2_nand4_1 _3373_ (.B(_2683_),
    .C(_2685_),
    .A(_2676_),
    .Y(_2837_),
    .D(_2690_));
 sg13g2_a21oi_1 _3374_ (.A1(_2683_),
    .A2(_2705_),
    .Y(_2838_),
    .B1(_2706_));
 sg13g2_nand2_1 _3375_ (.Y(_2839_),
    .A(_2837_),
    .B(_2838_));
 sg13g2_a21oi_1 _3376_ (.A1(_2808_),
    .A2(_2839_),
    .Y(_2840_),
    .B1(_2732_));
 sg13g2_inv_2 _3377_ (.Y(_2841_),
    .A(_2677_));
 sg13g2_and2_1 _3378_ (.A(_2841_),
    .B(_2706_),
    .X(_2842_));
 sg13g2_buf_1 _3379_ (.A(_2842_),
    .X(_2843_));
 sg13g2_xnor2_1 _3380_ (.Y(_2844_),
    .A(_2646_),
    .B(_2675_));
 sg13g2_xnor2_1 _3381_ (.Y(_2845_),
    .A(_2841_),
    .B(_2681_));
 sg13g2_nand3_1 _3382_ (.B(net132),
    .C(net42),
    .A(_2697_),
    .Y(_2846_));
 sg13g2_o21ai_1 _3383_ (.B1(_2846_),
    .Y(_2847_),
    .A1(net42),
    .A2(_2696_));
 sg13g2_nor3_1 _3384_ (.A(_2844_),
    .B(_2845_),
    .C(_2847_),
    .Y(_2848_));
 sg13g2_nor3_1 _3385_ (.A(_2646_),
    .B(_2701_),
    .C(_2689_),
    .Y(_2849_));
 sg13g2_o21ai_1 _3386_ (.B1(_2849_),
    .Y(_2850_),
    .A1(_2843_),
    .A2(_2848_));
 sg13g2_or2_1 _3387_ (.X(_2851_),
    .B(_2706_),
    .A(_2677_));
 sg13g2_mux2_1 _3388_ (.A0(_2841_),
    .A1(_2851_),
    .S(_2681_),
    .X(_2852_));
 sg13g2_nand2b_1 _3389_ (.Y(_2853_),
    .B(_2852_),
    .A_N(_2704_));
 sg13g2_a221oi_1 _3390_ (.B2(_2701_),
    .C1(_2689_),
    .B1(_2852_),
    .A1(_2683_),
    .Y(_2854_),
    .A2(_2762_));
 sg13g2_nand2_1 _3391_ (.Y(_2855_),
    .A(_2646_),
    .B(_2699_));
 sg13g2_nor2_1 _3392_ (.A(_2675_),
    .B(_2843_),
    .Y(_2856_));
 sg13g2_o21ai_1 _3393_ (.B1(_2856_),
    .Y(_2857_),
    .A1(_2845_),
    .A2(_2855_));
 sg13g2_and4_1 _3394_ (.A(_2647_),
    .B(_2675_),
    .C(_2683_),
    .D(_2762_),
    .X(_2858_));
 sg13g2_a221oi_1 _3395_ (.B2(_2857_),
    .C1(_2858_),
    .B1(_2854_),
    .A1(_2675_),
    .Y(_2859_),
    .A2(_2853_));
 sg13g2_and2_1 _3396_ (.A(_2850_),
    .B(_2859_),
    .X(_2860_));
 sg13g2_buf_1 _3397_ (.A(_2860_),
    .X(_2861_));
 sg13g2_a21oi_1 _3398_ (.A1(_2837_),
    .A2(_2838_),
    .Y(_2862_),
    .B1(_2785_));
 sg13g2_a21oi_2 _3399_ (.B1(_2783_),
    .Y(_2863_),
    .A2(_2862_),
    .A1(_2808_));
 sg13g2_o21ai_1 _3400_ (.B1(_2863_),
    .Y(_2864_),
    .A1(_2840_),
    .A2(_2861_));
 sg13g2_and2_1 _3401_ (.A(net130),
    .B(_2723_),
    .X(_2865_));
 sg13g2_a21o_1 _3402_ (.A2(_2865_),
    .A1(_2721_),
    .B1(_2724_),
    .X(_2866_));
 sg13g2_buf_1 _3403_ (.A(_2866_),
    .X(_2867_));
 sg13g2_nand2_1 _3404_ (.Y(_2868_),
    .A(net107),
    .B(net106));
 sg13g2_nand2_1 _3405_ (.Y(_2869_),
    .A(_2664_),
    .B(_2868_));
 sg13g2_buf_2 _3406_ (.A(_2869_),
    .X(_2870_));
 sg13g2_o21ai_1 _3407_ (.B1(_2870_),
    .Y(_2871_),
    .A1(_2720_),
    .A2(_2867_));
 sg13g2_nor2b_1 _3408_ (.A(_2724_),
    .B_N(_2721_),
    .Y(_2872_));
 sg13g2_buf_1 _3409_ (.A(_2872_),
    .X(_2873_));
 sg13g2_inv_1 _3410_ (.Y(_2874_),
    .A(_2721_));
 sg13g2_buf_8 _3411_ (.A(\game.fsm.block_len[2][1] ),
    .X(_2875_));
 sg13g2_buf_2 _3412_ (.A(\game.fsm.block_len[3][1] ),
    .X(_2876_));
 sg13g2_nand2b_1 _3413_ (.Y(_2877_),
    .B(_2876_),
    .A_N(_2875_));
 sg13g2_buf_2 _3414_ (.A(\game.fsm.block_len[3][0] ),
    .X(_2878_));
 sg13g2_buf_2 _3415_ (.A(\game.fsm.block_len[2][0] ),
    .X(_2879_));
 sg13g2_nor2b_1 _3416_ (.A(_2878_),
    .B_N(_2879_),
    .Y(_2880_));
 sg13g2_nor2b_1 _3417_ (.A(_2876_),
    .B_N(_2875_),
    .Y(_2881_));
 sg13g2_a221oi_1 _3418_ (.B2(_2880_),
    .C1(_2881_),
    .B1(_2877_),
    .A1(_2724_),
    .Y(_2882_),
    .A2(_2874_));
 sg13g2_buf_1 _3419_ (.A(_2882_),
    .X(_2883_));
 sg13g2_or2_1 _3420_ (.X(_2884_),
    .B(_2883_),
    .A(_2873_));
 sg13g2_nor2b_1 _3421_ (.A(_2875_),
    .B_N(_2876_),
    .Y(_2885_));
 sg13g2_xor2_1 _3422_ (.B(_2878_),
    .A(_2879_),
    .X(_2886_));
 sg13g2_or4_1 _3423_ (.A(_2873_),
    .B(_2885_),
    .C(_2881_),
    .D(_2886_),
    .X(_2887_));
 sg13g2_nand4_1 _3424_ (.B(_2884_),
    .C(_2865_),
    .A(_0092_),
    .Y(_2888_),
    .D(_2887_));
 sg13g2_nor2_1 _3425_ (.A(_2873_),
    .B(_2883_),
    .Y(_2889_));
 sg13g2_nand2_1 _3426_ (.Y(_2890_),
    .A(_2865_),
    .B(_2887_));
 sg13g2_o21ai_1 _3427_ (.B1(_0093_),
    .Y(_2891_),
    .A1(_2889_),
    .A2(_2890_));
 sg13g2_mux2_1 _3428_ (.A0(_0091_),
    .A1(_0090_),
    .S(_2718_),
    .X(_2892_));
 sg13g2_buf_1 _3429_ (.A(_2892_),
    .X(_2893_));
 sg13g2_a221oi_1 _3430_ (.B2(_2891_),
    .C1(_2893_),
    .B1(_2888_),
    .A1(_2720_),
    .Y(_2894_),
    .A2(_2867_));
 sg13g2_mux2_1 _3431_ (.A0(_0087_),
    .A1(_0086_),
    .S(_2718_),
    .X(_2895_));
 sg13g2_o21ai_1 _3432_ (.B1(_2895_),
    .Y(_2896_),
    .A1(_2871_),
    .A2(_2894_));
 sg13g2_nand2_1 _3433_ (.Y(_2897_),
    .A(_2720_),
    .B(_2867_));
 sg13g2_nand3_1 _3434_ (.B(_2891_),
    .C(_2893_),
    .A(_2888_),
    .Y(_2898_));
 sg13g2_a21oi_1 _3435_ (.A1(_2897_),
    .A2(_2898_),
    .Y(_2899_),
    .B1(_2871_));
 sg13g2_inv_1 _3436_ (.Y(_2900_),
    .A(_0083_));
 sg13g2_nand2b_1 _3437_ (.Y(_2901_),
    .B(_2884_),
    .A_N(_2890_));
 sg13g2_nand2_1 _3438_ (.Y(_2902_),
    .A(_0084_),
    .B(_2901_));
 sg13g2_o21ai_1 _3439_ (.B1(_2902_),
    .Y(_2903_),
    .A1(_2900_),
    .A2(_2901_));
 sg13g2_o21ai_1 _3440_ (.B1(_2903_),
    .Y(_2904_),
    .A1(_2895_),
    .A2(_2899_));
 sg13g2_and2_1 _3441_ (.A(_2896_),
    .B(_2904_),
    .X(_2905_));
 sg13g2_buf_2 _3442_ (.A(_2905_),
    .X(_2906_));
 sg13g2_nand3_1 _3443_ (.B(_2720_),
    .C(_2867_),
    .A(_2870_),
    .Y(_2907_));
 sg13g2_nor2b_1 _3444_ (.A(_2893_),
    .B_N(_2907_),
    .Y(_2908_));
 sg13g2_nand2_1 _3445_ (.Y(_2909_),
    .A(_2888_),
    .B(_2891_));
 sg13g2_a21oi_1 _3446_ (.A1(_2871_),
    .A2(_2893_),
    .Y(_2910_),
    .B1(_2909_));
 sg13g2_nor2_1 _3447_ (.A(_2908_),
    .B(_2910_),
    .Y(_2911_));
 sg13g2_nor2_1 _3448_ (.A(_2906_),
    .B(_2911_),
    .Y(_2912_));
 sg13g2_a21oi_1 _3449_ (.A1(_2701_),
    .A2(_2675_),
    .Y(_2913_),
    .B1(_2843_));
 sg13g2_o21ai_1 _3450_ (.B1(_2913_),
    .Y(_2914_),
    .A1(_2844_),
    .A2(_2847_));
 sg13g2_and3_1 _3451_ (.X(_2915_),
    .A(_2703_),
    .B(_2852_),
    .C(_2914_));
 sg13g2_mux2_1 _3452_ (.A0(_2685_),
    .A1(_2686_),
    .S(_2915_),
    .X(_2916_));
 sg13g2_and3_1 _3453_ (.X(_2917_),
    .A(_2861_),
    .B(_2863_),
    .C(_2916_));
 sg13g2_a21o_1 _3454_ (.A2(_2839_),
    .A1(_2808_),
    .B1(_2732_),
    .X(_2918_));
 sg13g2_or2_1 _3455_ (.X(_2919_),
    .B(_2910_),
    .A(_2908_));
 sg13g2_buf_1 _3456_ (.A(_2919_),
    .X(_2920_));
 sg13g2_nand3_1 _3457_ (.B(_2906_),
    .C(_2920_),
    .A(_2918_),
    .Y(_2921_));
 sg13g2_a22oi_1 _3458_ (.Y(_2922_),
    .B1(_2917_),
    .B2(_2921_),
    .A2(_2912_),
    .A1(_2864_));
 sg13g2_buf_1 _3459_ (.A(\game.fsm.length[2] ),
    .X(_2923_));
 sg13g2_inv_1 _3460_ (.Y(_2924_),
    .A(net128));
 sg13g2_buf_1 _3461_ (.A(_2924_),
    .X(_2925_));
 sg13g2_buf_2 _3462_ (.A(\game.fsm.seq[1][1] ),
    .X(_2926_));
 sg13g2_buf_2 _3463_ (.A(\game.fsm.length[0] ),
    .X(_2927_));
 sg13g2_buf_2 _3464_ (.A(\game.fsm.length[1] ),
    .X(_2928_));
 sg13g2_nor2_1 _3465_ (.A(_2927_),
    .B(_2928_),
    .Y(_2929_));
 sg13g2_buf_1 _3466_ (.A(\game.fsm.seq[2][1] ),
    .X(_2930_));
 sg13g2_nor2_1 _3467_ (.A(net127),
    .B(_2924_),
    .Y(_2931_));
 sg13g2_buf_2 _3468_ (.A(\game.fsm.seq[3][1] ),
    .X(_2932_));
 sg13g2_nand2b_1 _3469_ (.Y(_2933_),
    .B(net128),
    .A_N(_2928_));
 sg13g2_nand2b_1 _3470_ (.Y(_2934_),
    .B(_2928_),
    .A_N(net128));
 sg13g2_o21ai_1 _3471_ (.B1(_2934_),
    .Y(_0387_),
    .A1(_2932_),
    .A2(_2933_));
 sg13g2_buf_1 _3472_ (.A(_2927_),
    .X(_0388_));
 sg13g2_buf_2 _3473_ (.A(\game.fsm.seq[0][1] ),
    .X(_0389_));
 sg13g2_nor2_1 _3474_ (.A(_0389_),
    .B(_2934_),
    .Y(_0390_));
 sg13g2_a221oi_1 _3475_ (.B2(net104),
    .C1(_0390_),
    .B1(_0387_),
    .A1(_2929_),
    .Y(_0391_),
    .A2(_2931_));
 sg13g2_or2_1 _3476_ (.X(_0392_),
    .B(_0391_),
    .A(_2926_));
 sg13g2_buf_2 _3477_ (.A(\game.fsm.seq[5][1] ),
    .X(_0393_));
 sg13g2_buf_1 _3478_ (.A(_2928_),
    .X(_0394_));
 sg13g2_nand2_1 _3479_ (.Y(_0395_),
    .A(_0394_),
    .B(net128));
 sg13g2_nor2_1 _3480_ (.A(_0393_),
    .B(_0395_),
    .Y(_0396_));
 sg13g2_buf_1 _3481_ (.A(net103),
    .X(_0397_));
 sg13g2_buf_1 _3482_ (.A(\game.fsm.seq[7][1] ),
    .X(_0398_));
 sg13g2_buf_1 _3483_ (.A(net128),
    .X(_0399_));
 sg13g2_nor3_1 _3484_ (.A(net71),
    .B(_0398_),
    .C(net102),
    .Y(_0400_));
 sg13g2_nor2_1 _3485_ (.A(_0396_),
    .B(_0400_),
    .Y(_0401_));
 sg13g2_buf_1 _3486_ (.A(net71),
    .X(_0402_));
 sg13g2_o21ai_1 _3487_ (.B1(_0401_),
    .Y(_0403_),
    .A1(_0402_),
    .A2(_0391_));
 sg13g2_buf_2 _3488_ (.A(\game.fsm.seq[4][1] ),
    .X(_0404_));
 sg13g2_nor2_1 _3489_ (.A(_0404_),
    .B(_0395_),
    .Y(_0405_));
 sg13g2_buf_2 _3490_ (.A(\game.fsm.seq[6][1] ),
    .X(_0406_));
 sg13g2_nor3_1 _3491_ (.A(net71),
    .B(_0406_),
    .C(net102),
    .Y(_0407_));
 sg13g2_nor2_1 _3492_ (.A(_0405_),
    .B(_0407_),
    .Y(_0408_));
 sg13g2_nand2_1 _3493_ (.Y(_0409_),
    .A(_0391_),
    .B(_0408_));
 sg13g2_inv_1 _3494_ (.Y(_0410_),
    .A(_2927_));
 sg13g2_buf_1 _3495_ (.A(_0410_),
    .X(_0411_));
 sg13g2_mux4_1 _3496_ (.S0(_2926_),
    .A0(_0401_),
    .A1(_0403_),
    .A2(_0408_),
    .A3(_0409_),
    .S1(net70),
    .X(_0412_));
 sg13g2_buf_1 _3497_ (.A(\game.fsm.seq[2][0] ),
    .X(_0413_));
 sg13g2_inv_1 _3498_ (.Y(_0414_),
    .A(net126));
 sg13g2_nor2_1 _3499_ (.A(net104),
    .B(_0414_),
    .Y(_0415_));
 sg13g2_buf_1 _3500_ (.A(\game.fsm.seq[3][0] ),
    .X(_0416_));
 sg13g2_inv_1 _3501_ (.Y(_0417_),
    .A(_0416_));
 sg13g2_nor2_1 _3502_ (.A(net71),
    .B(_2924_),
    .Y(_0418_));
 sg13g2_buf_1 _3503_ (.A(\game.fsm.seq[0][0] ),
    .X(_0419_));
 sg13g2_o21ai_1 _3504_ (.B1(_2933_),
    .Y(_0420_),
    .A1(_0419_),
    .A2(_2934_));
 sg13g2_nand2_2 _3505_ (.Y(_0421_),
    .A(_2927_),
    .B(net103));
 sg13g2_nor3_1 _3506_ (.A(net128),
    .B(\game.fsm.seq[1][0] ),
    .C(_0421_),
    .Y(_0422_));
 sg13g2_a221oi_1 _3507_ (.B2(_0410_),
    .C1(_0422_),
    .B1(_0420_),
    .A1(_0417_),
    .Y(_0423_),
    .A2(_0418_));
 sg13g2_buf_2 _3508_ (.A(\game.fsm.seq[6][0] ),
    .X(_0424_));
 sg13g2_buf_1 _3509_ (.A(\game.fsm.seq[7][0] ),
    .X(_0425_));
 sg13g2_buf_2 _3510_ (.A(\game.fsm.seq[4][0] ),
    .X(_0426_));
 sg13g2_buf_1 _3511_ (.A(\game.fsm.seq[5][0] ),
    .X(_0427_));
 sg13g2_mux4_1 _3512_ (.S0(net104),
    .A0(_0424_),
    .A1(_0425_),
    .A2(_0426_),
    .A3(_0427_),
    .S1(net103),
    .X(_0428_));
 sg13g2_inv_2 _3513_ (.Y(_0429_),
    .A(net103));
 sg13g2_nand3b_1 _3514_ (.B(_2925_),
    .C(_0429_),
    .Y(_0430_),
    .A_N(_0428_));
 sg13g2_o21ai_1 _3515_ (.B1(_0430_),
    .Y(_0431_),
    .A1(_0415_),
    .A2(_0423_));
 sg13g2_or2_1 _3516_ (.X(_0432_),
    .B(_0428_),
    .A(_2924_));
 sg13g2_a21oi_1 _3517_ (.A1(_0423_),
    .A2(_0432_),
    .Y(_0433_),
    .B1(_0429_));
 sg13g2_o21ai_1 _3518_ (.B1(_0065_),
    .Y(_0434_),
    .A1(_0431_),
    .A2(_0433_));
 sg13g2_or3_1 _3519_ (.A(_0065_),
    .B(_0431_),
    .C(_0433_),
    .X(_0435_));
 sg13g2_buf_2 _3520_ (.A(_0067_),
    .X(_0436_));
 sg13g2_buf_1 _3521_ (.A(_0436_),
    .X(_0437_));
 sg13g2_nand2_1 _3522_ (.Y(_0438_),
    .A(_0414_),
    .B(net101));
 sg13g2_inv_1 _3523_ (.Y(_0439_),
    .A(_0064_));
 sg13g2_mux2_1 _3524_ (.A0(_0426_),
    .A1(_0439_),
    .S(_0436_),
    .X(_0440_));
 sg13g2_or2_1 _3525_ (.X(_0441_),
    .B(_0427_),
    .A(_0436_));
 sg13g2_mux2_1 _3526_ (.A0(_0416_),
    .A1(_0425_),
    .S(_0436_),
    .X(_0442_));
 sg13g2_mux4_1 _3527_ (.S0(_0429_),
    .A0(_0438_),
    .A1(_0440_),
    .A2(_0441_),
    .A3(_0442_),
    .S1(_0410_),
    .X(_0443_));
 sg13g2_mux2_1 _3528_ (.A0(_0424_),
    .A1(net126),
    .S(_0436_),
    .X(_0444_));
 sg13g2_nand3b_1 _3529_ (.B(net101),
    .C(_0065_),
    .Y(_0445_),
    .A_N(net104));
 sg13g2_o21ai_1 _3530_ (.B1(_0445_),
    .Y(_0446_),
    .A1(_0410_),
    .A2(_0444_));
 sg13g2_nand2_1 _3531_ (.Y(_0447_),
    .A(net71),
    .B(_0446_));
 sg13g2_a21oi_1 _3532_ (.A1(_0443_),
    .A2(_0447_),
    .Y(_0448_),
    .B1(_0439_));
 sg13g2_and3_1 _3533_ (.X(_0449_),
    .A(_0439_),
    .B(_0443_),
    .C(_0447_));
 sg13g2_mux4_1 _3534_ (.S0(_2927_),
    .A0(_0398_),
    .A1(_0404_),
    .A2(_0393_),
    .A3(_0406_),
    .S1(net103),
    .X(_0450_));
 sg13g2_inv_1 _3535_ (.Y(_0451_),
    .A(_0450_));
 sg13g2_mux4_1 _3536_ (.S0(_2927_),
    .A0(_2932_),
    .A1(_0389_),
    .A2(_2926_),
    .A3(net127),
    .S1(_2928_),
    .X(_0452_));
 sg13g2_inv_1 _3537_ (.Y(_0453_),
    .A(_0452_));
 sg13g2_xor2_1 _3538_ (.B(_2929_),
    .A(_0436_),
    .X(_0454_));
 sg13g2_mux2_1 _3539_ (.A0(_0451_),
    .A1(_0453_),
    .S(_0454_),
    .X(_0455_));
 sg13g2_buf_2 _3540_ (.A(_0455_),
    .X(_0456_));
 sg13g2_xor2_1 _3541_ (.B(_0456_),
    .A(_0389_),
    .X(_0457_));
 sg13g2_o21ai_1 _3542_ (.B1(_0457_),
    .Y(_0458_),
    .A1(_0448_),
    .A2(_0449_));
 sg13g2_a221oi_1 _3543_ (.B2(_0435_),
    .C1(_0458_),
    .B1(_0434_),
    .A1(_0392_),
    .Y(_0459_),
    .A2(_0412_));
 sg13g2_nor3_1 _3544_ (.A(net72),
    .B(net129),
    .C(_0459_),
    .Y(_0460_));
 sg13g2_o21ai_1 _3545_ (.B1(net102),
    .Y(_0461_),
    .A1(_0429_),
    .A2(_0426_));
 sg13g2_o21ai_1 _3546_ (.B1(_2925_),
    .Y(_0462_),
    .A1(_0397_),
    .A2(_0424_));
 sg13g2_nand3b_1 _3547_ (.B(net103),
    .C(_0064_),
    .Y(_0463_),
    .A_N(_2923_));
 sg13g2_a21oi_1 _3548_ (.A1(_2933_),
    .A2(_0463_),
    .Y(_0464_),
    .B1(net70));
 sg13g2_a221oi_1 _3549_ (.B2(_0397_),
    .C1(net70),
    .B1(_0464_),
    .A1(_0461_),
    .Y(_0465_),
    .A2(_0462_));
 sg13g2_buf_1 _3550_ (.A(net104),
    .X(_0466_));
 sg13g2_mux2_1 _3551_ (.A0(_0427_),
    .A1(_0425_),
    .S(net103),
    .X(_0467_));
 sg13g2_nor2_1 _3552_ (.A(_0399_),
    .B(_0467_),
    .Y(_0468_));
 sg13g2_o21ai_1 _3553_ (.B1(net126),
    .Y(_0469_),
    .A1(_0466_),
    .A2(_0468_));
 sg13g2_or2_1 _3554_ (.X(_0470_),
    .B(_0469_),
    .A(_0465_));
 sg13g2_mux4_1 _3555_ (.S0(net71),
    .A0(_2926_),
    .A1(_2932_),
    .A2(net127),
    .A3(_0389_),
    .S1(net104),
    .X(_0471_));
 sg13g2_mux4_1 _3556_ (.S0(net71),
    .A0(_0393_),
    .A1(_0398_),
    .A2(_0406_),
    .A3(_0404_),
    .S1(net104),
    .X(_0472_));
 sg13g2_xnor2_1 _3557_ (.Y(_0473_),
    .A(_2924_),
    .B(_0421_));
 sg13g2_mux2_1 _3558_ (.A0(_0471_),
    .A1(_0472_),
    .S(_0473_),
    .X(_0474_));
 sg13g2_xnor2_1 _3559_ (.Y(_0475_),
    .A(net127),
    .B(_0474_));
 sg13g2_o21ai_1 _3560_ (.B1(net128),
    .Y(_0476_),
    .A1(_0065_),
    .A2(_0394_));
 sg13g2_nor2_1 _3561_ (.A(_0388_),
    .B(_0476_),
    .Y(_0477_));
 sg13g2_nand4_1 _3562_ (.B(_0417_),
    .C(net126),
    .A(_0411_),
    .Y(_0478_),
    .D(_0477_));
 sg13g2_nor2_1 _3563_ (.A(_0477_),
    .B(_0464_),
    .Y(_0479_));
 sg13g2_nor3_1 _3564_ (.A(net71),
    .B(_0424_),
    .C(_0399_),
    .Y(_0480_));
 sg13g2_nor3_1 _3565_ (.A(_0429_),
    .B(_0426_),
    .C(net72),
    .Y(_0481_));
 sg13g2_nor4_1 _3566_ (.A(_0411_),
    .B(net126),
    .C(_0480_),
    .D(_0481_),
    .Y(_0482_));
 sg13g2_o21ai_1 _3567_ (.B1(_0417_),
    .Y(_0483_),
    .A1(_0477_),
    .A2(_0464_));
 sg13g2_nor3_1 _3568_ (.A(_0388_),
    .B(net126),
    .C(_0468_),
    .Y(_0484_));
 sg13g2_nor4_1 _3569_ (.A(_0466_),
    .B(net50),
    .C(_0414_),
    .D(_0476_),
    .Y(_0485_));
 sg13g2_a221oi_1 _3570_ (.B2(_0484_),
    .C1(_0485_),
    .B1(_0483_),
    .A1(_0479_),
    .Y(_0486_),
    .A2(_0482_));
 sg13g2_nand4_1 _3571_ (.B(_0475_),
    .C(_0478_),
    .A(_0470_),
    .Y(_0487_),
    .D(_0486_));
 sg13g2_nor2_1 _3572_ (.A(net129),
    .B(_0395_),
    .Y(_0488_));
 sg13g2_nor2_1 _3573_ (.A(_0429_),
    .B(net129),
    .Y(_0489_));
 sg13g2_a22oi_1 _3574_ (.Y(_0490_),
    .B1(_0489_),
    .B2(_0458_),
    .A2(_0488_),
    .A1(_0487_));
 sg13g2_o21ai_1 _3575_ (.B1(_0490_),
    .Y(_0491_),
    .A1(_2795_),
    .A2(_0458_));
 sg13g2_buf_2 _3576_ (.A(\game.current_level[1] ),
    .X(_0492_));
 sg13g2_inv_2 _3577_ (.Y(_0493_),
    .A(_0492_));
 sg13g2_o21ai_1 _3578_ (.B1(_0493_),
    .Y(_0494_),
    .A1(_0460_),
    .A2(_0491_));
 sg13g2_buf_1 _3579_ (.A(\game.current_level[2] ),
    .X(_0495_));
 sg13g2_buf_1 _3580_ (.A(_0495_),
    .X(_0496_));
 sg13g2_buf_2 _3581_ (.A(\game.fsm.color_count[3][1] ),
    .X(_0497_));
 sg13g2_buf_1 _3582_ (.A(\game.fsm.color_count[3][0] ),
    .X(_0498_));
 sg13g2_nor2_1 _3583_ (.A(_0497_),
    .B(net125),
    .Y(_0499_));
 sg13g2_buf_1 _3584_ (.A(\game.fsm.color_count[0][0] ),
    .X(_0500_));
 sg13g2_buf_1 _3585_ (.A(_0500_),
    .X(_0501_));
 sg13g2_buf_1 _3586_ (.A(\game.fsm.color_count[0][1] ),
    .X(_0502_));
 sg13g2_buf_1 _3587_ (.A(\game.fsm.color_count[0][2] ),
    .X(_0503_));
 sg13g2_or2_1 _3588_ (.X(_0504_),
    .B(_0503_),
    .A(_0502_));
 sg13g2_buf_1 _3589_ (.A(_0504_),
    .X(_0505_));
 sg13g2_nor2_1 _3590_ (.A(net99),
    .B(_0505_),
    .Y(_0506_));
 sg13g2_a21oi_1 _3591_ (.A1(_0071_),
    .A2(_0499_),
    .Y(_0507_),
    .B1(_0506_));
 sg13g2_buf_2 _3592_ (.A(\game.fsm.color_count[1][1] ),
    .X(_0508_));
 sg13g2_inv_1 _3593_ (.Y(_0509_),
    .A(_0508_));
 sg13g2_inv_1 _3594_ (.Y(_0510_),
    .A(\game.fsm.color_count[1][0] ));
 sg13g2_nand3_1 _3595_ (.B(_0510_),
    .C(_0070_),
    .A(_0509_),
    .Y(_0511_));
 sg13g2_buf_1 _3596_ (.A(_0511_),
    .X(_0512_));
 sg13g2_nor2_1 _3597_ (.A(_2800_),
    .B(_0512_),
    .Y(_0513_));
 sg13g2_a21oi_1 _3598_ (.A1(_2800_),
    .A2(_0507_),
    .Y(_0514_),
    .B1(_0513_));
 sg13g2_nor2_1 _3599_ (.A(_0493_),
    .B(_0514_),
    .Y(_0515_));
 sg13g2_nor3_1 _3600_ (.A(net100),
    .B(\game.current_level[4] ),
    .C(_0515_),
    .Y(_0516_));
 sg13g2_xnor2_1 _3601_ (.Y(_0517_),
    .A(_2932_),
    .B(net127));
 sg13g2_nor4_1 _3602_ (.A(_0416_),
    .B(net126),
    .C(net72),
    .D(_0517_),
    .Y(_0518_));
 sg13g2_inv_1 _3603_ (.Y(_0519_),
    .A(net127));
 sg13g2_nand3b_1 _3604_ (.B(net103),
    .C(net101),
    .Y(_0520_),
    .A_N(net104));
 sg13g2_nand2b_1 _3605_ (.Y(_0521_),
    .B(_0066_),
    .A_N(net128));
 sg13g2_nand4_1 _3606_ (.B(_0519_),
    .C(_0520_),
    .A(_0414_),
    .Y(_0522_),
    .D(_0521_));
 sg13g2_o21ai_1 _3607_ (.B1(_2926_),
    .Y(_0523_),
    .A1(_0389_),
    .A2(_0419_));
 sg13g2_inv_1 _3608_ (.Y(_0524_),
    .A(_0523_));
 sg13g2_inv_1 _3609_ (.Y(_0525_),
    .A(_0419_));
 sg13g2_a21oi_1 _3610_ (.A1(_0389_),
    .A2(_0525_),
    .Y(_0526_),
    .B1(_2926_));
 sg13g2_nand4_1 _3611_ (.B(net127),
    .C(_0520_),
    .A(_0414_),
    .Y(_0527_),
    .D(_0521_));
 sg13g2_a221oi_1 _3612_ (.B2(_0527_),
    .C1(\game.fsm.seq[1][0] ),
    .B1(_0526_),
    .A1(_0522_),
    .Y(_0528_),
    .A2(_0524_));
 sg13g2_or2_1 _3613_ (.X(_0529_),
    .B(_0528_),
    .A(_0518_));
 sg13g2_nor2_1 _3614_ (.A(_0424_),
    .B(_0066_),
    .Y(_0530_));
 sg13g2_xor2_1 _3615_ (.B(_0406_),
    .A(_0393_),
    .X(_0531_));
 sg13g2_xor2_1 _3616_ (.B(_0404_),
    .A(_0393_),
    .X(_0532_));
 sg13g2_inv_1 _3617_ (.Y(_0533_),
    .A(_0426_));
 sg13g2_a22oi_1 _3618_ (.Y(_0534_),
    .B1(_0532_),
    .B2(_0533_),
    .A2(_0531_),
    .A1(_0530_));
 sg13g2_nor3_1 _3619_ (.A(_0427_),
    .B(net72),
    .C(_0534_),
    .Y(_0535_));
 sg13g2_o21ai_1 _3620_ (.B1(net50),
    .Y(_0536_),
    .A1(_0529_),
    .A2(_0535_));
 sg13g2_xnor2_1 _3621_ (.Y(_0537_),
    .A(_2932_),
    .B(_0404_));
 sg13g2_nor4_1 _3622_ (.A(_0416_),
    .B(net101),
    .C(_2929_),
    .D(_0537_),
    .Y(_0538_));
 sg13g2_a221oi_1 _3623_ (.B2(_0533_),
    .C1(_0493_),
    .B1(_0538_),
    .A1(net102),
    .Y(_0539_),
    .A2(_0529_));
 sg13g2_inv_1 _3624_ (.Y(_0540_),
    .A(_0502_));
 sg13g2_inv_1 _3625_ (.Y(_0541_),
    .A(net99));
 sg13g2_buf_1 _3626_ (.A(_0503_),
    .X(_0542_));
 sg13g2_nor4_1 _3627_ (.A(net98),
    .B(_0541_),
    .C(_0542_),
    .D(_0492_),
    .Y(_0543_));
 sg13g2_a21oi_1 _3628_ (.A1(_0536_),
    .A2(_0539_),
    .Y(_0544_),
    .B1(_0543_));
 sg13g2_buf_1 _3629_ (.A(\game.fsm.color_count[2][2] ),
    .X(_0545_));
 sg13g2_inv_1 _3630_ (.Y(_0546_),
    .A(net124));
 sg13g2_buf_1 _3631_ (.A(\game.fsm.color_count[3][2] ),
    .X(_0547_));
 sg13g2_inv_1 _3632_ (.Y(_0548_),
    .A(net123));
 sg13g2_buf_2 _3633_ (.A(\game.fsm.color_count[2][0] ),
    .X(_0549_));
 sg13g2_inv_1 _3634_ (.Y(_0550_),
    .A(_0549_));
 sg13g2_nand2_1 _3635_ (.Y(_0551_),
    .A(net125),
    .B(_0550_));
 sg13g2_buf_2 _3636_ (.A(\game.fsm.color_count[2][1] ),
    .X(_0552_));
 sg13g2_nor2_1 _3637_ (.A(_0552_),
    .B(_0549_),
    .Y(_0553_));
 sg13g2_a21oi_1 _3638_ (.A1(net125),
    .A2(_0553_),
    .Y(_0554_),
    .B1(_0497_));
 sg13g2_a221oi_1 _3639_ (.B2(_0552_),
    .C1(_0554_),
    .B1(_0551_),
    .A1(_0545_),
    .Y(_0555_),
    .A2(_0548_));
 sg13g2_a21oi_1 _3640_ (.A1(_0546_),
    .A2(_0547_),
    .Y(_0556_),
    .B1(_0555_));
 sg13g2_nand2_1 _3641_ (.Y(_0557_),
    .A(_0072_),
    .B(_0553_));
 sg13g2_nand2_1 _3642_ (.Y(_0558_),
    .A(_0071_),
    .B(_0499_));
 sg13g2_xnor2_1 _3643_ (.Y(_0559_),
    .A(_0558_),
    .B(_0506_));
 sg13g2_mux2_1 _3644_ (.A0(_0507_),
    .A1(_0559_),
    .S(_0512_),
    .X(_0560_));
 sg13g2_nor2b_1 _3645_ (.A(_0557_),
    .B_N(_0512_),
    .Y(_0561_));
 sg13g2_a221oi_1 _3646_ (.B2(_0507_),
    .C1(_0492_),
    .B1(_0561_),
    .A1(_0557_),
    .Y(_0562_),
    .A2(_0560_));
 sg13g2_a21o_1 _3647_ (.A2(_0556_),
    .A1(_0492_),
    .B1(_0562_),
    .X(_0563_));
 sg13g2_mux2_1 _3648_ (.A0(_0544_),
    .A1(_0563_),
    .S(_2795_),
    .X(_0564_));
 sg13g2_inv_1 _3649_ (.Y(_0565_),
    .A(\game.current_level[4] ));
 sg13g2_nand2_1 _3650_ (.Y(_0566_),
    .A(_0495_),
    .B(_0565_));
 sg13g2_buf_2 _3651_ (.A(\game.current_level[3] ),
    .X(_0567_));
 sg13g2_nand2_1 _3652_ (.Y(_0568_),
    .A(_0567_),
    .B(_0565_));
 sg13g2_o21ai_1 _3653_ (.B1(_0568_),
    .Y(_0569_),
    .A1(_0564_),
    .A2(_0566_));
 sg13g2_a21o_1 _3654_ (.A2(_0516_),
    .A1(_0494_),
    .B1(_0569_),
    .X(_0570_));
 sg13g2_buf_1 _3655_ (.A(\game.fsm.color_count[1][2] ),
    .X(_0571_));
 sg13g2_nand2b_1 _3656_ (.Y(_0572_),
    .B(net122),
    .A_N(_0502_));
 sg13g2_nand2_1 _3657_ (.Y(_0573_),
    .A(_0509_),
    .B(_0572_));
 sg13g2_nand3_1 _3658_ (.B(net97),
    .C(net122),
    .A(_0502_),
    .Y(_0574_));
 sg13g2_or2_1 _3659_ (.X(_0575_),
    .B(net122),
    .A(net97));
 sg13g2_nand3_1 _3660_ (.B(_0574_),
    .C(_0575_),
    .A(_0508_),
    .Y(_0576_));
 sg13g2_nand3_1 _3661_ (.B(_0573_),
    .C(_0576_),
    .A(_0510_),
    .Y(_0577_));
 sg13g2_a21oi_1 _3662_ (.A1(_0505_),
    .A2(_0577_),
    .Y(_0578_),
    .B1(net99));
 sg13g2_xor2_1 _3663_ (.B(net122),
    .A(net97),
    .X(_0579_));
 sg13g2_nor3_1 _3664_ (.A(_0509_),
    .B(net98),
    .C(_0579_),
    .Y(_0580_));
 sg13g2_inv_1 _3665_ (.Y(_0581_),
    .A(_0503_));
 sg13g2_nor3_1 _3666_ (.A(_0508_),
    .B(_0581_),
    .C(_0572_),
    .Y(_0582_));
 sg13g2_o21ai_1 _3667_ (.B1(net99),
    .Y(_0583_),
    .A1(_0580_),
    .A2(_0582_));
 sg13g2_or3_1 _3668_ (.A(_0508_),
    .B(net122),
    .C(_0505_),
    .X(_0584_));
 sg13g2_a21oi_1 _3669_ (.A1(_0583_),
    .A2(_0584_),
    .Y(_0585_),
    .B1(_0510_));
 sg13g2_xnor2_1 _3670_ (.Y(_0586_),
    .A(_0508_),
    .B(_0497_));
 sg13g2_xnor2_1 _3671_ (.Y(_0587_),
    .A(net123),
    .B(net122));
 sg13g2_xnor2_1 _3672_ (.Y(_0588_),
    .A(\game.fsm.color_count[1][0] ),
    .B(net125));
 sg13g2_nand3_1 _3673_ (.B(_0587_),
    .C(_0588_),
    .A(_0586_),
    .Y(_0589_));
 sg13g2_xnor2_1 _3674_ (.Y(_0590_),
    .A(_0508_),
    .B(_0552_));
 sg13g2_xnor2_1 _3675_ (.Y(_0591_),
    .A(net124),
    .B(net122));
 sg13g2_xnor2_1 _3676_ (.Y(_0592_),
    .A(\game.fsm.color_count[1][0] ),
    .B(_0549_));
 sg13g2_nand3_1 _3677_ (.B(_0591_),
    .C(_0592_),
    .A(_0590_),
    .Y(_0593_));
 sg13g2_a22oi_1 _3678_ (.Y(_0594_),
    .B1(_0593_),
    .B2(_0557_),
    .A2(_0589_),
    .A1(_0558_));
 sg13g2_o21ai_1 _3679_ (.B1(_0594_),
    .Y(_0595_),
    .A1(_0578_),
    .A2(_0585_));
 sg13g2_nand2_1 _3680_ (.Y(_0596_),
    .A(_0541_),
    .B(_0581_));
 sg13g2_nand3_1 _3681_ (.B(net97),
    .C(_0549_),
    .A(net99),
    .Y(_0597_));
 sg13g2_or2_1 _3682_ (.X(_0598_),
    .B(_0549_),
    .A(_0500_));
 sg13g2_a21oi_1 _3683_ (.A1(_0597_),
    .A2(_0598_),
    .Y(_0599_),
    .B1(_0546_));
 sg13g2_nor3_1 _3684_ (.A(net97),
    .B(_0550_),
    .C(net124),
    .Y(_0600_));
 sg13g2_inv_1 _3685_ (.Y(_0601_),
    .A(_0552_));
 sg13g2_o21ai_1 _3686_ (.B1(_0601_),
    .Y(_0602_),
    .A1(_0599_),
    .A2(_0600_));
 sg13g2_a21o_1 _3687_ (.A2(_0602_),
    .A1(_0596_),
    .B1(_0502_),
    .X(_0603_));
 sg13g2_xnor2_1 _3688_ (.Y(_0604_),
    .A(net97),
    .B(net124));
 sg13g2_nand3_1 _3689_ (.B(_0549_),
    .C(_0604_),
    .A(net99),
    .Y(_0605_));
 sg13g2_nor2b_1 _3690_ (.A(_0500_),
    .B_N(_0503_),
    .Y(_0606_));
 sg13g2_nand3_1 _3691_ (.B(net124),
    .C(_0606_),
    .A(_0550_),
    .Y(_0607_));
 sg13g2_a21oi_1 _3692_ (.A1(_0605_),
    .A2(_0607_),
    .Y(_0608_),
    .B1(net98));
 sg13g2_nor3_1 _3693_ (.A(_0549_),
    .B(net124),
    .C(_0596_),
    .Y(_0609_));
 sg13g2_o21ai_1 _3694_ (.B1(_0552_),
    .Y(_0610_),
    .A1(_0608_),
    .A2(_0609_));
 sg13g2_xnor2_1 _3695_ (.Y(_0611_),
    .A(net124),
    .B(net123));
 sg13g2_xnor2_1 _3696_ (.Y(_0612_),
    .A(_0497_),
    .B(_0552_));
 sg13g2_inv_1 _3697_ (.Y(_0613_),
    .A(net125));
 sg13g2_nand2_1 _3698_ (.Y(_0614_),
    .A(_0613_),
    .B(_0549_));
 sg13g2_and3_1 _3699_ (.X(_0615_),
    .A(_0551_),
    .B(_0612_),
    .C(_0614_));
 sg13g2_a22oi_1 _3700_ (.Y(_0616_),
    .B1(_0611_),
    .B2(_0615_),
    .A2(_0499_),
    .A1(_0071_));
 sg13g2_a21o_1 _3701_ (.A2(_0610_),
    .A1(_0603_),
    .B1(_0616_),
    .X(_0617_));
 sg13g2_xnor2_1 _3702_ (.Y(_0618_),
    .A(_0503_),
    .B(net123));
 sg13g2_nand3_1 _3703_ (.B(net125),
    .C(_0618_),
    .A(net99),
    .Y(_0619_));
 sg13g2_nand3_1 _3704_ (.B(net123),
    .C(_0606_),
    .A(_0613_),
    .Y(_0620_));
 sg13g2_a21oi_1 _3705_ (.A1(_0619_),
    .A2(_0620_),
    .Y(_0621_),
    .B1(net98));
 sg13g2_nor3_1 _3706_ (.A(net125),
    .B(net123),
    .C(_0596_),
    .Y(_0622_));
 sg13g2_o21ai_1 _3707_ (.B1(_0497_),
    .Y(_0623_),
    .A1(_0621_),
    .A2(_0622_));
 sg13g2_nand2b_1 _3708_ (.Y(_0624_),
    .B(_0606_),
    .A_N(_0499_));
 sg13g2_nand3_1 _3709_ (.B(_0581_),
    .C(net123),
    .A(_0501_),
    .Y(_0625_));
 sg13g2_inv_1 _3710_ (.Y(_0626_),
    .A(_0497_));
 sg13g2_nand2_1 _3711_ (.Y(_0627_),
    .A(_0626_),
    .B(_0498_));
 sg13g2_a22oi_1 _3712_ (.Y(_0628_),
    .B1(_0627_),
    .B2(_0501_),
    .A2(_0548_),
    .A1(_0542_));
 sg13g2_nand4_1 _3713_ (.B(_0624_),
    .C(_0625_),
    .A(net98),
    .Y(_0629_),
    .D(_0628_));
 sg13g2_and3_1 _3714_ (.X(_0630_),
    .A(_0558_),
    .B(_0623_),
    .C(_0629_));
 sg13g2_a221oi_1 _3715_ (.B2(_0557_),
    .C1(_0630_),
    .B1(_0617_),
    .A1(_0512_),
    .Y(_0631_),
    .A2(_0595_));
 sg13g2_nor2_1 _3716_ (.A(_2710_),
    .B(_2716_),
    .Y(_0632_));
 sg13g2_nand2b_1 _3717_ (.Y(_0633_),
    .B(_2655_),
    .A_N(_2656_));
 sg13g2_nor2b_1 _3718_ (.A(_2650_),
    .B_N(\game.fsm.block_len[5][0] ),
    .Y(_0634_));
 sg13g2_a21oi_1 _3719_ (.A1(_0633_),
    .A2(_0634_),
    .Y(_0635_),
    .B1(_2657_));
 sg13g2_nand2_1 _3720_ (.Y(_0636_),
    .A(_2726_),
    .B(_2668_));
 sg13g2_a21oi_1 _3721_ (.A1(_2660_),
    .A2(_0635_),
    .Y(_0637_),
    .B1(_0636_));
 sg13g2_o21ai_1 _3722_ (.B1(net130),
    .Y(_0638_),
    .A1(_0632_),
    .A2(_0637_));
 sg13g2_nand2b_1 _3723_ (.Y(_0639_),
    .B(_2709_),
    .A_N(_2724_));
 sg13g2_inv_1 _3724_ (.Y(_0640_),
    .A(_2712_));
 sg13g2_nor2_1 _3725_ (.A(_2875_),
    .B(_0640_),
    .Y(_0641_));
 sg13g2_inv_1 _3726_ (.Y(_0642_),
    .A(\game.fsm.block_len[1][0] ));
 sg13g2_a22oi_1 _3727_ (.Y(_0643_),
    .B1(_0640_),
    .B2(_2875_),
    .A2(_0642_),
    .A1(_2879_));
 sg13g2_nand2b_1 _3728_ (.Y(_0644_),
    .B(_2724_),
    .A_N(_2709_));
 sg13g2_o21ai_1 _3729_ (.B1(_0644_),
    .Y(_0645_),
    .A1(_0641_),
    .A2(_0643_));
 sg13g2_nand3_1 _3730_ (.B(_0639_),
    .C(_0645_),
    .A(_2870_),
    .Y(_0646_));
 sg13g2_nand2_1 _3731_ (.Y(_0647_),
    .A(net133),
    .B(_2874_));
 sg13g2_nor2b_1 _3732_ (.A(_2876_),
    .B_N(_2655_),
    .Y(_0648_));
 sg13g2_nand2b_1 _3733_ (.Y(_0649_),
    .B(_2878_),
    .A_N(_2650_));
 sg13g2_nand2b_1 _3734_ (.Y(_0650_),
    .B(_2876_),
    .A_N(_2655_));
 sg13g2_o21ai_1 _3735_ (.B1(_0650_),
    .Y(_0651_),
    .A1(_0648_),
    .A2(_0649_));
 sg13g2_nor2b_1 _3736_ (.A(net133),
    .B_N(_2721_),
    .Y(_0652_));
 sg13g2_a21oi_1 _3737_ (.A1(_0647_),
    .A2(_0651_),
    .Y(_0653_),
    .B1(_0652_));
 sg13g2_nor2b_1 _3738_ (.A(_0648_),
    .B_N(_0650_),
    .Y(_0654_));
 sg13g2_nor2b_1 _3739_ (.A(_2721_),
    .B_N(net133),
    .Y(_0655_));
 sg13g2_xor2_1 _3740_ (.B(_2878_),
    .A(_2650_),
    .X(_0656_));
 sg13g2_nor3_1 _3741_ (.A(_0655_),
    .B(_0652_),
    .C(_0656_),
    .Y(_0657_));
 sg13g2_a21oi_1 _3742_ (.A1(_0654_),
    .A2(_0657_),
    .Y(_0658_),
    .B1(_2783_));
 sg13g2_a22oi_1 _3743_ (.Y(_0659_),
    .B1(_0653_),
    .B2(_0658_),
    .A2(_0632_),
    .A1(net106));
 sg13g2_nand4_1 _3744_ (.B(_0638_),
    .C(_0646_),
    .A(_2901_),
    .Y(_0660_),
    .D(_0659_));
 sg13g2_nand2b_1 _3745_ (.Y(_0661_),
    .B(_2759_),
    .A_N(_0653_));
 sg13g2_xor2_1 _3746_ (.B(_2712_),
    .A(_2875_),
    .X(_0662_));
 sg13g2_xnor2_1 _3747_ (.Y(_0663_),
    .A(_2879_),
    .B(\game.fsm.block_len[1][0] ));
 sg13g2_nand3_1 _3748_ (.B(_0644_),
    .C(_0663_),
    .A(_0639_),
    .Y(_0664_));
 sg13g2_o21ai_1 _3749_ (.B1(_2870_),
    .Y(_0665_),
    .A1(_0662_),
    .A2(_0664_));
 sg13g2_a21o_1 _3750_ (.A2(_0645_),
    .A1(_0639_),
    .B1(_0665_),
    .X(_0666_));
 sg13g2_buf_1 _3751_ (.A(net106),
    .X(_0667_));
 sg13g2_nand2_1 _3752_ (.Y(_0668_),
    .A(_2711_),
    .B(_2709_));
 sg13g2_nand2b_1 _3753_ (.Y(_0669_),
    .B(\game.fsm.block_len[0][0] ),
    .A_N(\game.fsm.block_len[1][0] ));
 sg13g2_o21ai_1 _3754_ (.B1(_2713_),
    .Y(_0670_),
    .A1(_2715_),
    .A2(_0669_));
 sg13g2_a21o_1 _3755_ (.A2(_0670_),
    .A1(_0668_),
    .B1(_2710_),
    .X(_0671_));
 sg13g2_nand2_1 _3756_ (.Y(_0672_),
    .A(net130),
    .B(_2723_));
 sg13g2_nor3_2 _3757_ (.A(_2873_),
    .B(_2883_),
    .C(_0672_),
    .Y(_0673_));
 sg13g2_a21oi_1 _3758_ (.A1(_0667_),
    .A2(_0671_),
    .Y(_0674_),
    .B1(_0673_));
 sg13g2_a21oi_1 _3759_ (.A1(_2659_),
    .A2(_2663_),
    .Y(_0675_),
    .B1(_2666_));
 sg13g2_o21ai_1 _3760_ (.B1(_2728_),
    .Y(_0676_),
    .A1(_0671_),
    .A2(_0675_));
 sg13g2_nand4_1 _3761_ (.B(_0666_),
    .C(_0674_),
    .A(_0661_),
    .Y(_0677_),
    .D(_0676_));
 sg13g2_nand3_1 _3762_ (.B(_0660_),
    .C(_0677_),
    .A(_2794_),
    .Y(_0678_));
 sg13g2_o21ai_1 _3763_ (.B1(_0678_),
    .Y(_0679_),
    .A1(net105),
    .A2(_0631_));
 sg13g2_nand2_2 _3764_ (.Y(_0680_),
    .A(_2794_),
    .B(_0493_));
 sg13g2_buf_1 _3765_ (.A(\game.fsm.len2_block_count[0] ),
    .X(_0681_));
 sg13g2_nor2b_1 _3766_ (.A(_0681_),
    .B_N(\game.fsm.len2_block_count[1] ),
    .Y(_0682_));
 sg13g2_o21ai_1 _3767_ (.B1(_0495_),
    .Y(_0683_),
    .A1(_0680_),
    .A2(_0682_));
 sg13g2_a21oi_1 _3768_ (.A1(_0492_),
    .A2(_0679_),
    .Y(_0684_),
    .B1(_0683_));
 sg13g2_nand3_1 _3769_ (.B(_0684_),
    .C(_2832_),
    .A(_0570_),
    .Y(_0685_));
 sg13g2_nor2_1 _3770_ (.A(net98),
    .B(_0626_),
    .Y(_0686_));
 sg13g2_nor2_1 _3771_ (.A(_0497_),
    .B(_0618_),
    .Y(_0687_));
 sg13g2_a22oi_1 _3772_ (.Y(_0688_),
    .B1(_0687_),
    .B2(_0540_),
    .A2(_0686_),
    .A1(_0618_));
 sg13g2_xnor2_1 _3773_ (.Y(_0689_),
    .A(net99),
    .B(_0498_));
 sg13g2_nor3_1 _3774_ (.A(net129),
    .B(_0688_),
    .C(_0689_),
    .Y(_0690_));
 sg13g2_buf_1 _3775_ (.A(\game.fsm.len1_block_count[0] ),
    .X(_0691_));
 sg13g2_or2_1 _3776_ (.X(_0692_),
    .B(\game.fsm.len1_block_count[2] ),
    .A(\game.fsm.len1_block_count[1] ));
 sg13g2_nor2_1 _3777_ (.A(_0681_),
    .B(\game.fsm.len2_block_count[1] ),
    .Y(_0693_));
 sg13g2_nor4_1 _3778_ (.A(net105),
    .B(_0691_),
    .C(_0692_),
    .D(_0693_),
    .Y(_0694_));
 sg13g2_nor3_1 _3779_ (.A(_0492_),
    .B(_0690_),
    .C(_0694_),
    .Y(_0695_));
 sg13g2_nand2_1 _3780_ (.Y(_0696_),
    .A(net105),
    .B(_0492_));
 sg13g2_nor2_1 _3781_ (.A(_2664_),
    .B(_2757_),
    .Y(_0697_));
 sg13g2_nor2_1 _3782_ (.A(_2794_),
    .B(_0493_),
    .Y(_0698_));
 sg13g2_buf_1 _3783_ (.A(_0698_),
    .X(_0699_));
 sg13g2_buf_1 _3784_ (.A(\game.fsm.green_block_count[0] ),
    .X(_0700_));
 sg13g2_inv_1 _3785_ (.Y(_0701_),
    .A(\game.fsm.green_block_count[2] ));
 sg13g2_nand3b_1 _3786_ (.B(\game.fsm.green_block_count[1] ),
    .C(_0701_),
    .Y(_0702_),
    .A_N(_0700_));
 sg13g2_a21oi_1 _3787_ (.A1(net49),
    .A2(_0702_),
    .Y(_0703_),
    .B1(net100));
 sg13g2_o21ai_1 _3788_ (.B1(_0703_),
    .Y(_0704_),
    .A1(_0696_),
    .A2(_0697_));
 sg13g2_o21ai_1 _3789_ (.B1(_0567_),
    .Y(_0705_),
    .A1(_0695_),
    .A2(_0704_));
 sg13g2_nand2_1 _3790_ (.Y(_0706_),
    .A(net129),
    .B(_0493_));
 sg13g2_and2_1 _3791_ (.A(_0684_),
    .B(_0706_),
    .X(_0707_));
 sg13g2_o21ai_1 _3792_ (.B1(_0570_),
    .Y(_0708_),
    .A1(_0705_),
    .A2(_0707_));
 sg13g2_o21ai_1 _3793_ (.B1(_0708_),
    .Y(_0709_),
    .A1(_2922_),
    .A2(_0685_));
 sg13g2_buf_2 _3794_ (.A(_0709_),
    .X(_0710_));
 sg13g2_nor4_1 _3795_ (.A(_2840_),
    .B(_2861_),
    .C(_2906_),
    .D(_2911_),
    .Y(_0711_));
 sg13g2_nor2_1 _3796_ (.A(_2863_),
    .B(_2906_),
    .Y(_0712_));
 sg13g2_or3_1 _3797_ (.A(net129),
    .B(_0711_),
    .C(_0712_),
    .X(_0713_));
 sg13g2_and3_1 _3798_ (.X(_0714_),
    .A(_2850_),
    .B(_2859_),
    .C(_2911_));
 sg13g2_o21ai_1 _3799_ (.B1(_2863_),
    .Y(_0715_),
    .A1(_2840_),
    .A2(_0714_));
 sg13g2_inv_1 _3800_ (.Y(_0716_),
    .A(_2916_));
 sg13g2_a21oi_1 _3801_ (.A1(_2906_),
    .A2(_0715_),
    .Y(_0717_),
    .B1(_0716_));
 sg13g2_inv_1 _3802_ (.Y(_0718_),
    .A(_0691_));
 sg13g2_or2_1 _3803_ (.X(_0719_),
    .B(_0692_),
    .A(_0718_));
 sg13g2_o21ai_1 _3804_ (.B1(_2920_),
    .Y(_0720_),
    .A1(_2783_),
    .A2(_2918_));
 sg13g2_o21ai_1 _3805_ (.B1(_2861_),
    .Y(_0721_),
    .A1(_2863_),
    .A2(_2920_));
 sg13g2_and3_1 _3806_ (.X(_0722_),
    .A(_0719_),
    .B(_0720_),
    .C(_0721_));
 sg13g2_buf_2 _3807_ (.A(\game.fsm.len3_block_count[0] ),
    .X(_0723_));
 sg13g2_inv_1 _3808_ (.Y(_0724_),
    .A(\game.fsm.len3_block_count[1] ));
 sg13g2_a22oi_1 _3809_ (.Y(_0725_),
    .B1(_0720_),
    .B2(_0721_),
    .A2(_0724_),
    .A1(_0723_));
 sg13g2_nor4_2 _3810_ (.A(_0713_),
    .B(_0717_),
    .C(_0722_),
    .Y(_0726_),
    .D(_0725_));
 sg13g2_nor2b_1 _3811_ (.A(\game.fsm.len2_block_count[1] ),
    .B_N(_0681_),
    .Y(_0727_));
 sg13g2_nand2_1 _3812_ (.Y(_0728_),
    .A(net105),
    .B(_0727_));
 sg13g2_a21oi_1 _3813_ (.A1(net105),
    .A2(_2809_),
    .Y(_0729_),
    .B1(_0492_));
 sg13g2_o21ai_1 _3814_ (.B1(_0729_),
    .Y(_0730_),
    .A1(_2922_),
    .A2(_0728_));
 sg13g2_nor3_1 _3815_ (.A(_0710_),
    .B(_0726_),
    .C(_0730_),
    .Y(_0731_));
 sg13g2_nand2_1 _3816_ (.Y(_0732_),
    .A(_2648_),
    .B(net131));
 sg13g2_nand2_1 _3817_ (.Y(_0733_),
    .A(_2649_),
    .B(net131));
 sg13g2_nand2_1 _3818_ (.Y(_0734_),
    .A(net130),
    .B(_2726_));
 sg13g2_a21oi_1 _3819_ (.A1(_2659_),
    .A2(_2663_),
    .Y(_0735_),
    .B1(_0734_));
 sg13g2_buf_1 _3820_ (.A(_0735_),
    .X(_0736_));
 sg13g2_mux2_1 _3821_ (.A0(_0732_),
    .A1(_0733_),
    .S(net41),
    .X(_0737_));
 sg13g2_inv_1 _3822_ (.Y(_0738_),
    .A(_2648_));
 sg13g2_nand2_1 _3823_ (.Y(_0739_),
    .A(_0738_),
    .B(_2701_));
 sg13g2_inv_1 _3824_ (.Y(_0740_),
    .A(_2649_));
 sg13g2_nand2_1 _3825_ (.Y(_0741_),
    .A(_0740_),
    .B(_2701_));
 sg13g2_mux2_1 _3826_ (.A0(_0739_),
    .A1(_0741_),
    .S(net41),
    .X(_0742_));
 sg13g2_mux2_1 _3827_ (.A0(_2695_),
    .A1(_2697_),
    .S(net41),
    .X(_0743_));
 sg13g2_inv_1 _3828_ (.Y(_0744_),
    .A(_2764_));
 sg13g2_a221oi_1 _3829_ (.B2(net132),
    .C1(_0744_),
    .B1(_0743_),
    .A1(_0737_),
    .Y(_0745_),
    .A2(_0742_));
 sg13g2_mux2_1 _3830_ (.A0(_0738_),
    .A1(_0740_),
    .S(net41),
    .X(_0746_));
 sg13g2_buf_2 _3831_ (.A(_0746_),
    .X(_0747_));
 sg13g2_nand2_1 _3832_ (.Y(_0748_),
    .A(_2646_),
    .B(_2764_));
 sg13g2_nor2_1 _3833_ (.A(_2841_),
    .B(_2689_),
    .Y(_0749_));
 sg13g2_o21ai_1 _3834_ (.B1(_0749_),
    .Y(_0750_),
    .A1(_0747_),
    .A2(_0748_));
 sg13g2_inv_1 _3835_ (.Y(_0751_),
    .A(_2678_));
 sg13g2_inv_1 _3836_ (.Y(_0752_),
    .A(_2679_));
 sg13g2_mux2_1 _3837_ (.A0(_0751_),
    .A1(_0752_),
    .S(_0735_),
    .X(_0753_));
 sg13g2_buf_1 _3838_ (.A(_0753_),
    .X(_0754_));
 sg13g2_o21ai_1 _3839_ (.B1(_0754_),
    .Y(_0755_),
    .A1(_0745_),
    .A2(_0750_));
 sg13g2_a21oi_1 _3840_ (.A1(_2711_),
    .A2(_2709_),
    .Y(_0756_),
    .B1(_2717_));
 sg13g2_nor2b_1 _3841_ (.A(_2717_),
    .B_N(_2710_),
    .Y(_0757_));
 sg13g2_a21oi_2 _3842_ (.B1(_0757_),
    .Y(_0758_),
    .A2(_0756_),
    .A1(_0670_));
 sg13g2_mux2_1 _3843_ (.A0(_0027_),
    .A1(_0026_),
    .S(_0673_),
    .X(_0759_));
 sg13g2_buf_8 _3844_ (.A(_0759_),
    .X(_0760_));
 sg13g2_inv_1 _3845_ (.Y(_0761_),
    .A(_0088_));
 sg13g2_nor2_1 _3846_ (.A(_0761_),
    .B(_0758_),
    .Y(_0762_));
 sg13g2_a221oi_1 _3847_ (.B2(_2870_),
    .C1(_0762_),
    .B1(_0760_),
    .A1(_0089_),
    .Y(_0763_),
    .A2(_0758_));
 sg13g2_buf_1 _3848_ (.A(_0763_),
    .X(_0764_));
 sg13g2_and2_1 _3849_ (.A(_2759_),
    .B(_0764_),
    .X(_0765_));
 sg13g2_and2_1 _3850_ (.A(_0755_),
    .B(_0765_),
    .X(_0766_));
 sg13g2_or2_1 _3851_ (.X(_0767_),
    .B(_0750_),
    .A(_0745_));
 sg13g2_mux2_1 _3852_ (.A0(_2678_),
    .A1(_2679_),
    .S(net41),
    .X(_0768_));
 sg13g2_o21ai_1 _3853_ (.B1(_2759_),
    .Y(_0769_),
    .A1(_0764_),
    .A2(_0768_));
 sg13g2_nand2_1 _3854_ (.Y(_0770_),
    .A(_2678_),
    .B(_2841_));
 sg13g2_nand2_1 _3855_ (.Y(_0771_),
    .A(_2679_),
    .B(_2841_));
 sg13g2_mux2_1 _3856_ (.A0(_0770_),
    .A1(_0771_),
    .S(_0736_),
    .X(_0772_));
 sg13g2_and2_1 _3857_ (.A(_2703_),
    .B(_0772_),
    .X(_0773_));
 sg13g2_xnor2_1 _3858_ (.Y(_0774_),
    .A(_2764_),
    .B(_0754_));
 sg13g2_nor2_1 _3859_ (.A(_2647_),
    .B(_0747_),
    .Y(_0775_));
 sg13g2_a21oi_1 _3860_ (.A1(_2703_),
    .A2(_0772_),
    .Y(_0776_),
    .B1(_0747_));
 sg13g2_a221oi_1 _3861_ (.B2(_0775_),
    .C1(_0776_),
    .B1(_0774_),
    .A1(net131),
    .Y(_0777_),
    .A2(_0773_));
 sg13g2_inv_1 _3862_ (.Y(_0778_),
    .A(_0089_));
 sg13g2_mux2_1 _3863_ (.A0(_0761_),
    .A1(_0778_),
    .S(_0758_),
    .X(_0779_));
 sg13g2_buf_1 _3864_ (.A(_0779_),
    .X(_0780_));
 sg13g2_and2_1 _3865_ (.A(_0780_),
    .B(_0760_),
    .X(_0781_));
 sg13g2_mux2_1 _3866_ (.A0(_0093_),
    .A1(_0092_),
    .S(_0673_),
    .X(_0782_));
 sg13g2_buf_1 _3867_ (.A(_0782_),
    .X(_0783_));
 sg13g2_nor2b_1 _3868_ (.A(_0783_),
    .B_N(_2870_),
    .Y(_0784_));
 sg13g2_o21ai_1 _3869_ (.B1(_2870_),
    .Y(_0785_),
    .A1(_0780_),
    .A2(_0760_));
 sg13g2_inv_1 _3870_ (.Y(_0786_),
    .A(_0090_));
 sg13g2_inv_1 _3871_ (.Y(_0787_),
    .A(_0091_));
 sg13g2_mux2_1 _3872_ (.A0(_0786_),
    .A1(_0787_),
    .S(_0758_),
    .X(_0788_));
 sg13g2_buf_1 _3873_ (.A(_0788_),
    .X(_0789_));
 sg13g2_nor2b_1 _3874_ (.A(_0783_),
    .B_N(_0789_),
    .Y(_0790_));
 sg13g2_a221oi_1 _3875_ (.B2(_0789_),
    .C1(_0790_),
    .B1(_0785_),
    .A1(_0781_),
    .Y(_0791_),
    .A2(_0784_));
 sg13g2_buf_1 _3876_ (.A(_0791_),
    .X(_0792_));
 sg13g2_a22oi_1 _3877_ (.Y(_0793_),
    .B1(_0777_),
    .B2(_0792_),
    .A2(_0769_),
    .A1(_0767_));
 sg13g2_mux2_1 _3878_ (.A0(_2696_),
    .A1(_2698_),
    .S(net41),
    .X(_0794_));
 sg13g2_a21oi_1 _3879_ (.A1(net131),
    .A2(_0794_),
    .Y(_0795_),
    .B1(_2646_));
 sg13g2_or2_1 _3880_ (.X(_0796_),
    .B(_0795_),
    .A(_0747_));
 sg13g2_nor2_1 _3881_ (.A(_2648_),
    .B(net131),
    .Y(_0797_));
 sg13g2_nor2_1 _3882_ (.A(_2649_),
    .B(net131),
    .Y(_0798_));
 sg13g2_mux2_1 _3883_ (.A0(_0797_),
    .A1(_0798_),
    .S(_0736_),
    .X(_0799_));
 sg13g2_a221oi_1 _3884_ (.B2(_0794_),
    .C1(_2689_),
    .B1(_0799_),
    .A1(_2841_),
    .Y(_0800_),
    .A2(_0768_));
 sg13g2_nor2b_1 _3885_ (.A(net132),
    .B_N(_0800_),
    .Y(_0801_));
 sg13g2_xnor2_1 _3886_ (.Y(_0802_),
    .A(_0744_),
    .B(_0754_));
 sg13g2_nor2_1 _3887_ (.A(_2695_),
    .B(net41),
    .Y(_0803_));
 sg13g2_a221oi_1 _3888_ (.B2(_0802_),
    .C1(_0803_),
    .B1(_0773_),
    .A1(_0075_),
    .Y(_0804_),
    .A2(net41));
 sg13g2_o21ai_1 _3889_ (.B1(_0800_),
    .Y(_0805_),
    .A1(_0747_),
    .A2(_0795_));
 sg13g2_nand2_1 _3890_ (.Y(_0806_),
    .A(_2703_),
    .B(_0772_));
 sg13g2_nor3_1 _3891_ (.A(net132),
    .B(_0806_),
    .C(_0774_),
    .Y(_0807_));
 sg13g2_a221oi_1 _3892_ (.B2(_0805_),
    .C1(_0807_),
    .B1(_0804_),
    .A1(_0796_),
    .Y(_0808_),
    .A2(_0801_));
 sg13g2_o21ai_1 _3893_ (.B1(_0808_),
    .Y(_0809_),
    .A1(_0766_),
    .A2(_0793_));
 sg13g2_mux2_1 _3894_ (.A0(_0086_),
    .A1(_0087_),
    .S(_0758_),
    .X(_0810_));
 sg13g2_inv_1 _3895_ (.Y(_0811_),
    .A(_0810_));
 sg13g2_nand2_1 _3896_ (.Y(_0812_),
    .A(_0780_),
    .B(_0760_));
 sg13g2_nor2_1 _3897_ (.A(_0783_),
    .B(_0789_),
    .Y(_0813_));
 sg13g2_a21o_1 _3898_ (.A2(_0813_),
    .A1(_0812_),
    .B1(_0785_),
    .X(_0814_));
 sg13g2_a22oi_1 _3899_ (.Y(_0815_),
    .B1(_0783_),
    .B2(_0789_),
    .A2(_0760_),
    .A1(_0780_));
 sg13g2_or3_1 _3900_ (.A(_2873_),
    .B(_2883_),
    .C(_0672_),
    .X(_0816_));
 sg13g2_nor4_1 _3901_ (.A(_2900_),
    .B(_2873_),
    .C(_2883_),
    .D(_0672_),
    .Y(_0817_));
 sg13g2_a221oi_1 _3902_ (.B2(_0084_),
    .C1(_0817_),
    .B1(_0816_),
    .A1(_2664_),
    .Y(_0818_),
    .A2(_2868_));
 sg13g2_o21ai_1 _3903_ (.B1(_0818_),
    .Y(_0819_),
    .A1(_0780_),
    .A2(_0760_));
 sg13g2_and2_1 _3904_ (.A(_0084_),
    .B(_0816_),
    .X(_0820_));
 sg13g2_or3_1 _3905_ (.A(_0810_),
    .B(_0820_),
    .C(_0817_),
    .X(_0821_));
 sg13g2_o21ai_1 _3906_ (.B1(_0821_),
    .Y(_0822_),
    .A1(_0815_),
    .A2(_0819_));
 sg13g2_a21o_1 _3907_ (.A2(_0814_),
    .A1(_0811_),
    .B1(_0822_),
    .X(_0823_));
 sg13g2_a21oi_1 _3908_ (.A1(_0775_),
    .A2(_0774_),
    .Y(_0824_),
    .B1(_0776_));
 sg13g2_nand2_1 _3909_ (.Y(_0825_),
    .A(net131),
    .B(_0773_));
 sg13g2_a221oi_1 _3910_ (.B2(_0825_),
    .C1(_0792_),
    .B1(_0824_),
    .A1(_0767_),
    .Y(_0826_),
    .A2(_0769_));
 sg13g2_or3_1 _3911_ (.A(_0766_),
    .B(_0823_),
    .C(_0826_),
    .X(_0827_));
 sg13g2_nand2b_1 _3912_ (.Y(_0828_),
    .B(_0808_),
    .A_N(_0823_));
 sg13g2_nand3_1 _3913_ (.B(_0827_),
    .C(_0828_),
    .A(_0809_),
    .Y(_0829_));
 sg13g2_nor2_1 _3914_ (.A(_0745_),
    .B(_0750_),
    .Y(_0830_));
 sg13g2_nor2_1 _3915_ (.A(_2783_),
    .B(_0754_),
    .Y(_0831_));
 sg13g2_or4_1 _3916_ (.A(_0830_),
    .B(_0765_),
    .C(_0831_),
    .D(_0792_),
    .X(_0832_));
 sg13g2_nand3_1 _3917_ (.B(_0765_),
    .C(_0777_),
    .A(_0755_),
    .Y(_0833_));
 sg13g2_nand2b_1 _3918_ (.Y(_0834_),
    .B(_0777_),
    .A_N(_0792_));
 sg13g2_nand3_1 _3919_ (.B(_0833_),
    .C(_0834_),
    .A(_0832_),
    .Y(_0835_));
 sg13g2_or2_1 _3920_ (.X(_0836_),
    .B(_0719_),
    .A(_0835_));
 sg13g2_nand2_1 _3921_ (.Y(_0837_),
    .A(_2759_),
    .B(_0755_));
 sg13g2_nor2b_1 _3922_ (.A(\game.fsm.len3_block_count[1] ),
    .B_N(_0723_),
    .Y(_0838_));
 sg13g2_a221oi_1 _3923_ (.B2(_0838_),
    .C1(_0696_),
    .B1(_0835_),
    .A1(_0764_),
    .Y(_0839_),
    .A2(_0837_));
 sg13g2_nand3b_1 _3924_ (.B(_0836_),
    .C(_0839_),
    .Y(_0840_),
    .A_N(_0829_));
 sg13g2_nor4_1 _3925_ (.A(\game.fsm.len2_color_count[2][1] ),
    .B(\game.fsm.len3_color_count[3][1] ),
    .C(\game.fsm.len2_color_count[0][1] ),
    .D(\game.fsm.len1_color_count[3][2] ),
    .Y(_0841_));
 sg13g2_nor4_1 _3926_ (.A(\game.fsm.len1_color_count[2][1] ),
    .B(\game.fsm.len1_color_count[0][2] ),
    .C(\game.fsm.len1_color_count[1][2] ),
    .D(\game.fsm.len1_color_count[2][2] ),
    .Y(_0842_));
 sg13g2_nor4_1 _3927_ (.A(\game.fsm.len1_color_count[0][1] ),
    .B(\game.fsm.len1_color_count[1][1] ),
    .C(\game.fsm.len1_color_count[3][1] ),
    .D(\game.fsm.len3_color_count[2][1] ),
    .Y(_0843_));
 sg13g2_nor4_1 _3928_ (.A(\game.fsm.len2_color_count[1][1] ),
    .B(\game.fsm.len2_color_count[3][1] ),
    .C(\game.fsm.len3_color_count[1][1] ),
    .D(\game.fsm.len3_color_count[0][1] ),
    .Y(_0844_));
 sg13g2_nand4_1 _3929_ (.B(_0842_),
    .C(_0843_),
    .A(_0841_),
    .Y(_0845_),
    .D(_0844_));
 sg13g2_a221oi_1 _3930_ (.B2(_0727_),
    .C1(_0696_),
    .B1(_0835_),
    .A1(_0764_),
    .Y(_0846_),
    .A2(_0837_));
 sg13g2_nor2_1 _3931_ (.A(_0567_),
    .B(_0565_),
    .Y(_0847_));
 sg13g2_nand2b_1 _3932_ (.Y(_0848_),
    .B(_0847_),
    .A_N(net100));
 sg13g2_a221oi_1 _3933_ (.B2(_0846_),
    .C1(_0848_),
    .B1(_0829_),
    .A1(net49),
    .Y(_0849_),
    .A2(_0845_));
 sg13g2_nand2_1 _3934_ (.Y(_0850_),
    .A(_0840_),
    .B(_0849_));
 sg13g2_nor2b_1 _3935_ (.A(_0710_),
    .B_N(_0850_),
    .Y(_0851_));
 sg13g2_a21oi_1 _3936_ (.A1(_2836_),
    .A2(_0731_),
    .Y(_0852_),
    .B1(_0851_));
 sg13g2_buf_2 _3937_ (.A(_0852_),
    .X(_0853_));
 sg13g2_xor2_1 _3938_ (.B(_0853_),
    .A(\game.slv.saved_target ),
    .X(_0854_));
 sg13g2_buf_1 _3939_ (.A(\game.slv.pos[0] ),
    .X(_0855_));
 sg13g2_or3_1 _3940_ (.A(_0855_),
    .B(\game.slv.pos[1] ),
    .C(\game.slv.pos[2] ),
    .X(_0856_));
 sg13g2_buf_1 _3941_ (.A(_0856_),
    .X(_0857_));
 sg13g2_buf_1 _3942_ (.A(\game.slv.state[1] ),
    .X(_0858_));
 sg13g2_inv_2 _3943_ (.Y(_0859_),
    .A(_2638_));
 sg13g2_nor3_1 _3944_ (.A(_0859_),
    .B(_2636_),
    .C(_2637_),
    .Y(_0860_));
 sg13g2_a221oi_1 _3945_ (.B2(net121),
    .C1(_0860_),
    .B1(_0857_),
    .A1(\game.slv.state[3] ),
    .Y(_0861_),
    .A2(_0854_));
 sg13g2_nor2_1 _3946_ (.A(_2645_),
    .B(_0861_),
    .Y(_0011_));
 sg13g2_buf_1 _3947_ (.A(\game.state[1] ),
    .X(_0862_));
 sg13g2_buf_1 _3948_ (.A(\game.state[2] ),
    .X(_0863_));
 sg13g2_buf_1 _3949_ (.A(\game.challenge_num[1] ),
    .X(_0864_));
 sg13g2_buf_1 _3950_ (.A(\game.challenge_num[0] ),
    .X(_0865_));
 sg13g2_inv_1 _3951_ (.Y(_0866_),
    .A(_0865_));
 sg13g2_buf_2 _3952_ (.A(\game.challenge_num[2] ),
    .X(_0867_));
 sg13g2_buf_1 _3953_ (.A(\game.challenge_num[3] ),
    .X(_0868_));
 sg13g2_nand4_1 _3954_ (.B(_0866_),
    .C(_0867_),
    .A(_0864_),
    .Y(_0869_),
    .D(_0868_));
 sg13g2_nand2_1 _3955_ (.Y(_0870_),
    .A(net119),
    .B(_0869_));
 sg13g2_buf_2 _3956_ (.A(\game.state[0] ),
    .X(_0871_));
 sg13g2_buf_1 _3957_ (.A(\game.state[3] ),
    .X(_0872_));
 sg13g2_or2_1 _3958_ (.X(_0873_),
    .B(net118),
    .A(_0871_));
 sg13g2_buf_1 _3959_ (.A(_0873_),
    .X(_0874_));
 sg13g2_a21oi_1 _3960_ (.A1(net120),
    .A2(_0870_),
    .Y(_0875_),
    .B1(_0874_));
 sg13g2_buf_1 _3961_ (.A(_0875_),
    .X(_0876_));
 sg13g2_buf_1 _3962_ (.A(_0876_),
    .X(_0877_));
 sg13g2_nor2_1 _3963_ (.A(net120),
    .B(_0871_),
    .Y(_0878_));
 sg13g2_buf_1 _3964_ (.A(_0878_),
    .X(_0879_));
 sg13g2_nor2_1 _3965_ (.A(_0872_),
    .B(\game.state[2] ),
    .Y(_0880_));
 sg13g2_buf_2 _3966_ (.A(_0880_),
    .X(_0881_));
 sg13g2_and2_1 _3967_ (.A(_0879_),
    .B(_0881_),
    .X(_0882_));
 sg13g2_buf_1 _3968_ (.A(_0882_),
    .X(_0883_));
 sg13g2_buf_1 _3969_ (.A(\btn.input_event[4] ),
    .X(_0884_));
 sg13g2_buf_1 _3970_ (.A(\btn.input_event[0] ),
    .X(_0885_));
 sg13g2_buf_1 _3971_ (.A(\btn.input_event[1] ),
    .X(_0886_));
 sg13g2_inv_2 _3972_ (.Y(_0887_),
    .A(_0886_));
 sg13g2_nor2_2 _3973_ (.A(_0885_),
    .B(_0887_),
    .Y(_0888_));
 sg13g2_buf_1 _3974_ (.A(\btn.input_event[2] ),
    .X(_0889_));
 sg13g2_buf_2 _3975_ (.A(\btn.input_event[3] ),
    .X(_0890_));
 sg13g2_nor2_2 _3976_ (.A(_0889_),
    .B(_0890_),
    .Y(_0891_));
 sg13g2_nand3_1 _3977_ (.B(_0888_),
    .C(_0891_),
    .A(net117),
    .Y(_0892_));
 sg13g2_buf_1 _3978_ (.A(_0892_),
    .X(_0893_));
 sg13g2_and2_1 _3979_ (.A(_0883_),
    .B(_0893_),
    .X(_0894_));
 sg13g2_buf_1 _3980_ (.A(_0894_),
    .X(_0895_));
 sg13g2_inv_1 _3981_ (.Y(_0896_),
    .A(_0061_));
 sg13g2_nand3_1 _3982_ (.B(_0567_),
    .C(net49),
    .A(net100),
    .Y(_0897_));
 sg13g2_xnor2_1 _3983_ (.Y(_0898_),
    .A(_0896_),
    .B(_0897_));
 sg13g2_nand2_1 _3984_ (.Y(_0899_),
    .A(_0867_),
    .B(_0868_));
 sg13g2_nor3_1 _3985_ (.A(net120),
    .B(_0871_),
    .C(net118),
    .Y(_0900_));
 sg13g2_buf_2 _3986_ (.A(_0900_),
    .X(_0901_));
 sg13g2_nand2_1 _3987_ (.Y(_0902_),
    .A(_0864_),
    .B(_0865_));
 sg13g2_nor3_1 _3988_ (.A(_0899_),
    .B(_0901_),
    .C(_0902_),
    .Y(_0903_));
 sg13g2_a21oi_1 _3989_ (.A1(_0895_),
    .A2(_0898_),
    .Y(_0904_),
    .B1(_0903_));
 sg13g2_buf_1 _3990_ (.A(\display_value[4] ),
    .X(_0905_));
 sg13g2_nor2_1 _3991_ (.A(_0905_),
    .B(net30),
    .Y(_0906_));
 sg13g2_a21oi_2 _3992_ (.B1(_0906_),
    .Y(_0907_),
    .A2(_0904_),
    .A1(net30));
 sg13g2_inv_1 _3993_ (.Y(_0908_),
    .A(_0053_));
 sg13g2_xnor2_1 _3994_ (.Y(_0909_),
    .A(_0063_),
    .B(net49));
 sg13g2_nor2b_1 _3995_ (.A(net118),
    .B_N(net119),
    .Y(_0910_));
 sg13g2_buf_2 _3996_ (.A(_0910_),
    .X(_0911_));
 sg13g2_and2_1 _3997_ (.A(_0879_),
    .B(_0911_),
    .X(_0912_));
 sg13g2_buf_2 _3998_ (.A(_0912_),
    .X(_0913_));
 sg13g2_buf_1 _3999_ (.A(_0054_),
    .X(_0914_));
 sg13g2_inv_1 _4000_ (.Y(_0915_),
    .A(_0914_));
 sg13g2_xnor2_1 _4001_ (.Y(_0916_),
    .A(_0914_),
    .B(_0902_));
 sg13g2_nor2_1 _4002_ (.A(_0901_),
    .B(_0916_),
    .Y(_0917_));
 sg13g2_a221oi_1 _4003_ (.B2(_0915_),
    .C1(_0917_),
    .B1(_0913_),
    .A1(_0895_),
    .Y(_0918_),
    .A2(_0909_));
 sg13g2_nand2_1 _4004_ (.Y(_0919_),
    .A(_0876_),
    .B(_0918_));
 sg13g2_o21ai_1 _4005_ (.B1(_0919_),
    .Y(_0920_),
    .A1(_0908_),
    .A2(_0877_));
 sg13g2_buf_1 _4006_ (.A(_0920_),
    .X(_0921_));
 sg13g2_buf_1 _4007_ (.A(_0865_),
    .X(_0922_));
 sg13g2_nand3_1 _4008_ (.B(net96),
    .C(_0901_),
    .A(net119),
    .Y(_0923_));
 sg13g2_o21ai_1 _4009_ (.B1(_0923_),
    .Y(_0924_),
    .A1(net96),
    .A2(_0901_));
 sg13g2_a21o_1 _4010_ (.A2(_0895_),
    .A1(_0069_),
    .B1(_0924_),
    .X(_0925_));
 sg13g2_buf_1 _4011_ (.A(\display_value[0] ),
    .X(_0926_));
 sg13g2_nor2b_1 _4012_ (.A(_0876_),
    .B_N(_0926_),
    .Y(_0927_));
 sg13g2_a21o_1 _4013_ (.A2(_0925_),
    .A1(net30),
    .B1(_0927_),
    .X(_0928_));
 sg13g2_buf_1 _4014_ (.A(_0928_),
    .X(_0929_));
 sg13g2_nand2_1 _4015_ (.Y(_0930_),
    .A(_0879_),
    .B(_0881_));
 sg13g2_buf_2 _4016_ (.A(_0930_),
    .X(_0931_));
 sg13g2_nand2_1 _4017_ (.Y(_0932_),
    .A(_0879_),
    .B(_0911_));
 sg13g2_buf_1 _4018_ (.A(_0932_),
    .X(_0933_));
 sg13g2_xor2_1 _4019_ (.B(net96),
    .A(_0864_),
    .X(_0934_));
 sg13g2_nand2_1 _4020_ (.Y(_0935_),
    .A(net47),
    .B(_0934_));
 sg13g2_o21ai_1 _4021_ (.B1(_0935_),
    .Y(_0936_),
    .A1(_0052_),
    .A2(net47));
 sg13g2_nand2_1 _4022_ (.Y(_0937_),
    .A(_0696_),
    .B(_0706_));
 sg13g2_a22oi_1 _4023_ (.Y(_0938_),
    .B1(_0937_),
    .B2(_0895_),
    .A2(_0936_),
    .A1(_0931_));
 sg13g2_buf_2 _4024_ (.A(\display_value[1] ),
    .X(_0939_));
 sg13g2_nor2_1 _4025_ (.A(_0939_),
    .B(_0876_),
    .Y(_0940_));
 sg13g2_a21oi_2 _4026_ (.B1(_0940_),
    .Y(_0941_),
    .A2(_0938_),
    .A1(net30));
 sg13g2_nand2_1 _4027_ (.Y(_0942_),
    .A(_2640_),
    .B(_0941_));
 sg13g2_buf_2 _4028_ (.A(_0942_),
    .X(_0943_));
 sg13g2_inv_2 _4029_ (.Y(_0168_),
    .A(_0943_));
 sg13g2_nor2_1 _4030_ (.A(net24),
    .B(_0168_),
    .Y(_0944_));
 sg13g2_buf_1 _4031_ (.A(\display_value[3] ),
    .X(_0945_));
 sg13g2_inv_1 _4032_ (.Y(_0946_),
    .A(_0945_));
 sg13g2_buf_1 _4033_ (.A(_0055_),
    .X(_0947_));
 sg13g2_nor2_1 _4034_ (.A(_0947_),
    .B(net47),
    .Y(_0948_));
 sg13g2_buf_1 _4035_ (.A(_0883_),
    .X(_0949_));
 sg13g2_nand2_1 _4036_ (.Y(_0950_),
    .A(net40),
    .B(_0893_));
 sg13g2_nand2_1 _4037_ (.Y(_0951_),
    .A(net100),
    .B(net49));
 sg13g2_xnor2_1 _4038_ (.Y(_0952_),
    .A(_0062_),
    .B(_0951_));
 sg13g2_nand3_1 _4039_ (.B(_0865_),
    .C(_0867_),
    .A(_0864_),
    .Y(_0953_));
 sg13g2_xor2_1 _4040_ (.B(_0953_),
    .A(_0947_),
    .X(_0954_));
 sg13g2_nand2b_1 _4041_ (.Y(_0955_),
    .B(_0954_),
    .A_N(_0901_));
 sg13g2_o21ai_1 _4042_ (.B1(_0955_),
    .Y(_0956_),
    .A1(_0950_),
    .A2(_0952_));
 sg13g2_o21ai_1 _4043_ (.B1(_0876_),
    .Y(_0957_),
    .A1(_0948_),
    .A2(_0956_));
 sg13g2_o21ai_1 _4044_ (.B1(_0957_),
    .Y(_0958_),
    .A1(_0946_),
    .A2(_0876_));
 sg13g2_buf_2 _4045_ (.A(_0958_),
    .X(_0959_));
 sg13g2_inv_2 _4046_ (.Y(_0960_),
    .A(_0959_));
 sg13g2_o21ai_1 _4047_ (.B1(_0960_),
    .Y(_0961_),
    .A1(net21),
    .A2(_0944_));
 sg13g2_and2_1 _4048_ (.A(_0907_),
    .B(_0961_),
    .X(_0962_));
 sg13g2_a21oi_2 _4049_ (.B1(_0927_),
    .Y(_0963_),
    .A2(_0925_),
    .A1(net30));
 sg13g2_a21oi_1 _4050_ (.A1(_0921_),
    .A2(_0963_),
    .Y(_0964_),
    .B1(_0960_));
 sg13g2_nor2_1 _4051_ (.A(_0943_),
    .B(_0964_),
    .Y(_0965_));
 sg13g2_a21o_1 _4052_ (.A2(_0904_),
    .A1(net30),
    .B1(_0906_),
    .X(_0966_));
 sg13g2_buf_1 _4053_ (.A(_0966_),
    .X(_0967_));
 sg13g2_nand2b_1 _4054_ (.Y(_0968_),
    .B(net24),
    .A_N(net21));
 sg13g2_nand2_1 _4055_ (.Y(_0969_),
    .A(_0943_),
    .B(_0959_));
 sg13g2_nand3_1 _4056_ (.B(_0968_),
    .C(_0969_),
    .A(net23),
    .Y(_0970_));
 sg13g2_buf_1 _4057_ (.A(net134),
    .X(_0971_));
 sg13g2_o21ai_1 _4058_ (.B1(net95),
    .Y(_0972_),
    .A1(_0965_),
    .A2(_0970_));
 sg13g2_nor2_1 _4059_ (.A(_0962_),
    .B(_0972_),
    .Y(_0000_));
 sg13g2_buf_1 _4060_ (.A(net134),
    .X(_0973_));
 sg13g2_buf_1 _4061_ (.A(net94),
    .X(_0974_));
 sg13g2_nor2_1 _4062_ (.A(net21),
    .B(net24),
    .Y(_0975_));
 sg13g2_and2_1 _4063_ (.A(net21),
    .B(net24),
    .X(_0976_));
 sg13g2_nor3_1 _4064_ (.A(_0941_),
    .B(_0975_),
    .C(_0976_),
    .Y(_0977_));
 sg13g2_a21oi_1 _4065_ (.A1(_0941_),
    .A2(_0975_),
    .Y(_0978_),
    .B1(_0977_));
 sg13g2_nor2b_1 _4066_ (.A(_0921_),
    .B_N(_0941_),
    .Y(_0979_));
 sg13g2_o21ai_1 _4067_ (.B1(net23),
    .Y(_0980_),
    .A1(_0963_),
    .A2(_0960_));
 sg13g2_a22oi_1 _4068_ (.Y(_0981_),
    .B1(_0979_),
    .B2(_0980_),
    .A2(_0959_),
    .A1(_0907_));
 sg13g2_o21ai_1 _4069_ (.B1(_0981_),
    .Y(_0982_),
    .A1(_0959_),
    .A2(_0978_));
 sg13g2_nand2_1 _4070_ (.Y(_0001_),
    .A(_0974_),
    .B(_0982_));
 sg13g2_and2_1 _4071_ (.A(net21),
    .B(_0960_),
    .X(_0983_));
 sg13g2_buf_1 _4072_ (.A(_0983_),
    .X(_0984_));
 sg13g2_nor2_1 _4073_ (.A(net21),
    .B(_0960_),
    .Y(_0985_));
 sg13g2_a22oi_1 _4074_ (.Y(_0986_),
    .B1(_0985_),
    .B2(_0943_),
    .A2(_0984_),
    .A1(net23));
 sg13g2_nor2_1 _4075_ (.A(net24),
    .B(_0986_),
    .Y(_0987_));
 sg13g2_buf_1 _4076_ (.A(_0973_),
    .X(_0988_));
 sg13g2_o21ai_1 _4077_ (.B1(net66),
    .Y(_0002_),
    .A1(_0962_),
    .A2(_0987_));
 sg13g2_nand2_1 _4078_ (.Y(_0989_),
    .A(_0960_),
    .B(_0944_));
 sg13g2_nor3_1 _4079_ (.A(net24),
    .B(_0943_),
    .C(_0985_),
    .Y(_0990_));
 sg13g2_nor2_1 _4080_ (.A(_0943_),
    .B(_0959_),
    .Y(_0991_));
 sg13g2_o21ai_1 _4081_ (.B1(_0969_),
    .Y(_0992_),
    .A1(_0968_),
    .A2(_0991_));
 sg13g2_o21ai_1 _4082_ (.B1(net23),
    .Y(_0993_),
    .A1(_0990_),
    .A2(_0992_));
 sg13g2_o21ai_1 _4083_ (.B1(_0993_),
    .Y(_0994_),
    .A1(_0967_),
    .A2(_0989_));
 sg13g2_a22oi_1 _4084_ (.Y(_0995_),
    .B1(_0994_),
    .B2(net95),
    .A2(_0984_),
    .A1(_0168_));
 sg13g2_inv_1 _4085_ (.Y(_0003_),
    .A(_0995_));
 sg13g2_nor3_1 _4086_ (.A(net108),
    .B(net23),
    .C(_0960_),
    .Y(_0996_));
 sg13g2_nor2_1 _4087_ (.A(_2641_),
    .B(_0960_),
    .Y(_0170_));
 sg13g2_nor2_1 _4088_ (.A(_2641_),
    .B(net23),
    .Y(_0171_));
 sg13g2_nor2_1 _4089_ (.A(_0170_),
    .B(_0171_),
    .Y(_0997_));
 sg13g2_nor2_1 _4090_ (.A(net21),
    .B(_0943_),
    .Y(_0998_));
 sg13g2_nor2_1 _4091_ (.A(_0997_),
    .B(_0998_),
    .Y(_0999_));
 sg13g2_a21oi_1 _4092_ (.A1(_0168_),
    .A2(_0997_),
    .Y(_1000_),
    .B1(_0999_));
 sg13g2_nor3_1 _4093_ (.A(_0929_),
    .B(_0996_),
    .C(_1000_),
    .Y(_0004_));
 sg13g2_nor3_1 _4094_ (.A(net23),
    .B(_0959_),
    .C(_0998_),
    .Y(_1001_));
 sg13g2_nor3_1 _4095_ (.A(_0963_),
    .B(_0943_),
    .C(_0985_),
    .Y(_1002_));
 sg13g2_nor3_1 _4096_ (.A(_0907_),
    .B(_0984_),
    .C(_1002_),
    .Y(_1003_));
 sg13g2_nor2_1 _4097_ (.A(_1001_),
    .B(_1003_),
    .Y(_1004_));
 sg13g2_a21oi_1 _4098_ (.A1(_0907_),
    .A2(net24),
    .Y(_1005_),
    .B1(_0985_));
 sg13g2_o21ai_1 _4099_ (.B1(net95),
    .Y(_1006_),
    .A1(_0168_),
    .A2(_1005_));
 sg13g2_nor2_1 _4100_ (.A(_1004_),
    .B(_1006_),
    .Y(_0005_));
 sg13g2_nand2_1 _4101_ (.Y(_1007_),
    .A(net21),
    .B(_0959_));
 sg13g2_o21ai_1 _4102_ (.B1(_1007_),
    .Y(_1008_),
    .A1(_0968_),
    .A2(_0959_));
 sg13g2_nor2_1 _4103_ (.A(net23),
    .B(net24),
    .Y(_1009_));
 sg13g2_o21ai_1 _4104_ (.B1(_0984_),
    .Y(_1010_),
    .A1(_0168_),
    .A2(_1009_));
 sg13g2_nand2b_1 _4105_ (.Y(_1011_),
    .B(_0967_),
    .A_N(_0984_));
 sg13g2_buf_1 _4106_ (.A(net108),
    .X(_1012_));
 sg13g2_a221oi_1 _4107_ (.B2(_1011_),
    .C1(net65),
    .B1(_1010_),
    .A1(_0168_),
    .Y(_0006_),
    .A2(_1008_));
 sg13g2_inv_1 _4108_ (.Y(_1013_),
    .A(\game.slv.state[1] ));
 sg13g2_nor3_1 _4109_ (.A(_1013_),
    .B(_2645_),
    .C(_0857_),
    .Y(_0010_));
 sg13g2_nand2_1 _4110_ (.Y(_1014_),
    .A(_0443_),
    .B(_0447_));
 sg13g2_buf_1 _4111_ (.A(_1014_),
    .X(_1015_));
 sg13g2_buf_1 _4112_ (.A(\game.solver_active ),
    .X(_1016_));
 sg13g2_buf_1 _4113_ (.A(_1016_),
    .X(_1017_));
 sg13g2_nor2b_1 _4114_ (.A(net93),
    .B_N(\game.input_color[0] ),
    .Y(_1018_));
 sg13g2_a21oi_1 _4115_ (.A1(_1017_),
    .A2(\game.slv.fsm_color[0] ),
    .Y(_1019_),
    .B1(_1018_));
 sg13g2_buf_2 _4116_ (.A(_1019_),
    .X(_1020_));
 sg13g2_xnor2_1 _4117_ (.Y(_1021_),
    .A(_1015_),
    .B(_1020_));
 sg13g2_nor3_2 _4118_ (.A(net69),
    .B(net50),
    .C(net102),
    .Y(_1022_));
 sg13g2_inv_1 _4119_ (.Y(_1023_),
    .A(\game.input_color[1] ));
 sg13g2_nor2_1 _4120_ (.A(net93),
    .B(_1023_),
    .Y(_1024_));
 sg13g2_a21o_1 _4121_ (.A2(\game.slv.fsm_color[1] ),
    .A1(net93),
    .B1(_1024_),
    .X(_1025_));
 sg13g2_buf_1 _4122_ (.A(_1025_),
    .X(_1026_));
 sg13g2_xnor2_1 _4123_ (.Y(_1027_),
    .A(_0456_),
    .B(_1026_));
 sg13g2_nor2_1 _4124_ (.A(_1022_),
    .B(_1027_),
    .Y(_1028_));
 sg13g2_nand2_1 _4125_ (.Y(_1029_),
    .A(_1021_),
    .B(_1028_));
 sg13g2_buf_2 _4126_ (.A(_1029_),
    .X(_1030_));
 sg13g2_mux4_1 _4127_ (.S0(_2688_),
    .A0(_2697_),
    .A1(\game.fsm.block_len[6][0] ),
    .A2(_2900_),
    .A3(_2695_),
    .S1(_2666_),
    .X(_1031_));
 sg13g2_inv_1 _4128_ (.Y(_1032_),
    .A(\game.fsm.block_len[7][0] ));
 sg13g2_mux4_1 _4129_ (.S0(net106),
    .A0(_1032_),
    .A1(_0086_),
    .A2(_0087_),
    .A3(_0084_),
    .S1(net107),
    .X(_1033_));
 sg13g2_nand2_1 _4130_ (.Y(_1034_),
    .A(_2722_),
    .B(_1033_));
 sg13g2_o21ai_1 _4131_ (.B1(_1034_),
    .Y(_1035_),
    .A1(_2722_),
    .A2(_1031_));
 sg13g2_buf_1 _4132_ (.A(_1035_),
    .X(_1036_));
 sg13g2_nor2_1 _4133_ (.A(_0437_),
    .B(_0421_),
    .Y(_1037_));
 sg13g2_nor2b_1 _4134_ (.A(_1016_),
    .B_N(_0031_),
    .Y(_1038_));
 sg13g2_a21oi_1 _4135_ (.A1(_0032_),
    .A2(_1016_),
    .Y(_1039_),
    .B1(_1038_));
 sg13g2_buf_1 _4136_ (.A(_1039_),
    .X(_1040_));
 sg13g2_nor2b_1 _4137_ (.A(_1037_),
    .B_N(net48),
    .Y(_1041_));
 sg13g2_buf_2 _4138_ (.A(_1041_),
    .X(_1042_));
 sg13g2_buf_1 _4139_ (.A(_1042_),
    .X(_1043_));
 sg13g2_o21ai_1 _4140_ (.B1(net28),
    .Y(_1044_),
    .A1(_1030_),
    .A2(net39));
 sg13g2_inv_1 _4141_ (.Y(_1045_),
    .A(\game.input_erase ));
 sg13g2_nor3_1 _4142_ (.A(net93),
    .B(_1045_),
    .C(_1022_),
    .Y(_1046_));
 sg13g2_buf_2 _4143_ (.A(_1046_),
    .X(_1047_));
 sg13g2_nand2_1 _4144_ (.Y(_1048_),
    .A(net39),
    .B(_1047_));
 sg13g2_nor2b_1 _4145_ (.A(_1016_),
    .B_N(\game.input_reset ),
    .Y(_1049_));
 sg13g2_a21o_1 _4146_ (.A2(\game.slv.fsm_reset ),
    .A1(net93),
    .B1(_1049_),
    .X(_1050_));
 sg13g2_buf_1 _4147_ (.A(_1050_),
    .X(_1051_));
 sg13g2_buf_1 _4148_ (.A(_1051_),
    .X(_1052_));
 sg13g2_a21oi_1 _4149_ (.A1(_1044_),
    .A2(_1048_),
    .Y(_1053_),
    .B1(net46));
 sg13g2_buf_2 _4150_ (.A(_1053_),
    .X(_1054_));
 sg13g2_a21oi_1 _4151_ (.A1(net93),
    .A2(\game.slv.fsm_reset ),
    .Y(_1055_),
    .B1(_1049_));
 sg13g2_buf_2 _4152_ (.A(_1055_),
    .X(_1056_));
 sg13g2_buf_1 _4153_ (.A(_1056_),
    .X(_1057_));
 sg13g2_buf_1 _4154_ (.A(net45),
    .X(_1058_));
 sg13g2_and2_1 _4155_ (.A(\game.fsm.block_len[0][0] ),
    .B(net38),
    .X(_1059_));
 sg13g2_nand2b_1 _4156_ (.Y(_1060_),
    .B(net48),
    .A_N(_1037_));
 sg13g2_buf_1 _4157_ (.A(_1060_),
    .X(_1061_));
 sg13g2_nor2_1 _4158_ (.A(_1051_),
    .B(_1061_),
    .Y(_1062_));
 sg13g2_buf_2 _4159_ (.A(_1062_),
    .X(_1063_));
 sg13g2_nand2_1 _4160_ (.Y(_1064_),
    .A(_1030_),
    .B(_1063_));
 sg13g2_nor2_2 _4161_ (.A(net107),
    .B(net106),
    .Y(_1065_));
 sg13g2_nand2_2 _4162_ (.Y(_1066_),
    .A(net37),
    .B(_1047_));
 sg13g2_nand3_1 _4163_ (.B(_1021_),
    .C(_1028_),
    .A(_1042_),
    .Y(_1067_));
 sg13g2_buf_1 _4164_ (.A(_1067_),
    .X(_1068_));
 sg13g2_a21oi_2 _4165_ (.B1(_1051_),
    .Y(_1069_),
    .A2(_1068_),
    .A1(_1066_));
 sg13g2_o21ai_1 _4166_ (.B1(_1069_),
    .Y(_1070_),
    .A1(_2727_),
    .A2(_1065_));
 sg13g2_o21ai_1 _4167_ (.B1(_1070_),
    .Y(_1071_),
    .A1(_0073_),
    .A2(_1064_));
 sg13g2_buf_1 _4168_ (.A(_1071_),
    .X(_1072_));
 sg13g2_inv_2 _4169_ (.Y(_1073_),
    .A(_2722_));
 sg13g2_xnor2_1 _4170_ (.Y(_1074_),
    .A(_1073_),
    .B(_1065_));
 sg13g2_nand2_1 _4171_ (.Y(_1075_),
    .A(_1069_),
    .B(_1074_));
 sg13g2_o21ai_1 _4172_ (.B1(_1075_),
    .Y(_1076_),
    .A1(net130),
    .A2(_1064_));
 sg13g2_buf_1 _4173_ (.A(_1076_),
    .X(_1077_));
 sg13g2_nand2b_1 _4174_ (.Y(_1078_),
    .B(_1077_),
    .A_N(_1072_));
 sg13g2_buf_1 _4175_ (.A(net107),
    .X(_1079_));
 sg13g2_nand2_1 _4176_ (.Y(_1080_),
    .A(net64),
    .B(_1069_));
 sg13g2_o21ai_1 _4177_ (.B1(_1080_),
    .Y(_1081_),
    .A1(net64),
    .A2(_1064_));
 sg13g2_buf_1 _4178_ (.A(_1081_),
    .X(_1082_));
 sg13g2_nand2b_1 _4179_ (.Y(_1083_),
    .B(_1082_),
    .A_N(_1078_));
 sg13g2_buf_1 _4180_ (.A(_1083_),
    .X(_1084_));
 sg13g2_mux2_1 _4181_ (.A0(_1054_),
    .A1(_1059_),
    .S(_1084_),
    .X(_0172_));
 sg13g2_inv_1 _4182_ (.Y(_1085_),
    .A(\game.fsm.block_len[7][1] ));
 sg13g2_nand2_1 _4183_ (.Y(_1086_),
    .A(_1073_),
    .B(_2876_));
 sg13g2_nor2_1 _4184_ (.A(_2666_),
    .B(_2712_),
    .Y(_1087_));
 sg13g2_a22oi_1 _4185_ (.Y(_1088_),
    .B1(_1086_),
    .B2(_1087_),
    .A2(_1085_),
    .A1(_2666_));
 sg13g2_nand2_1 _4186_ (.Y(_1089_),
    .A(net68),
    .B(_2656_));
 sg13g2_o21ai_1 _4187_ (.B1(_1089_),
    .Y(_1090_),
    .A1(net68),
    .A2(_1086_));
 sg13g2_mux2_1 _4188_ (.A0(\game.fsm.block_len[0][1] ),
    .A1(_2875_),
    .S(net68),
    .X(_1091_));
 sg13g2_nor2_1 _4189_ (.A(net68),
    .B(_2655_),
    .Y(_1092_));
 sg13g2_a21oi_1 _4190_ (.A1(net68),
    .A2(_2647_),
    .Y(_1093_),
    .B1(_1092_));
 sg13g2_mux4_1 _4191_ (.S0(_1073_),
    .A0(_1088_),
    .A1(_1090_),
    .A2(_1091_),
    .A3(_1093_),
    .S1(net64),
    .X(_1094_));
 sg13g2_buf_1 _4192_ (.A(_1094_),
    .X(_1095_));
 sg13g2_nand2b_1 _4193_ (.Y(_1096_),
    .B(net39),
    .A_N(_1095_));
 sg13g2_inv_1 _4194_ (.Y(_1097_),
    .A(net39));
 sg13g2_nand2_1 _4195_ (.Y(_1098_),
    .A(_1097_),
    .B(_1095_));
 sg13g2_nand2_1 _4196_ (.Y(_1099_),
    .A(_1096_),
    .B(_1098_));
 sg13g2_or3_1 _4197_ (.A(net93),
    .B(_1045_),
    .C(_1022_),
    .X(_1100_));
 sg13g2_buf_1 _4198_ (.A(_1100_),
    .X(_1101_));
 sg13g2_nor2_1 _4199_ (.A(_1042_),
    .B(_1101_),
    .Y(_1102_));
 sg13g2_buf_2 _4200_ (.A(_1102_),
    .X(_1103_));
 sg13g2_nand2_1 _4201_ (.Y(_1104_),
    .A(_1103_),
    .B(_1099_));
 sg13g2_o21ai_1 _4202_ (.B1(_1104_),
    .Y(_1105_),
    .A1(_1068_),
    .A2(_1099_));
 sg13g2_nand2_2 _4203_ (.Y(_1106_),
    .A(net45),
    .B(_1105_));
 sg13g2_buf_1 _4204_ (.A(_1057_),
    .X(_1107_));
 sg13g2_nand3_1 _4205_ (.B(net36),
    .C(_1084_),
    .A(\game.fsm.block_len[0][1] ),
    .Y(_1108_));
 sg13g2_o21ai_1 _4206_ (.B1(_1108_),
    .Y(_0173_),
    .A1(_1084_),
    .A2(_1106_));
 sg13g2_nor2_1 _4207_ (.A(net106),
    .B(_2678_),
    .Y(_1109_));
 sg13g2_a21oi_1 _4208_ (.A1(_0667_),
    .A2(_2764_),
    .Y(_1110_),
    .B1(_1109_));
 sg13g2_nor2_1 _4209_ (.A(_2722_),
    .B(_1110_),
    .Y(_1111_));
 sg13g2_inv_1 _4210_ (.Y(_1112_),
    .A(_0026_));
 sg13g2_nand3_1 _4211_ (.B(_1112_),
    .C(_1065_),
    .A(_1073_),
    .Y(_1113_));
 sg13g2_o21ai_1 _4212_ (.B1(_1113_),
    .Y(_1114_),
    .A1(_1073_),
    .A2(_1065_));
 sg13g2_nor2_1 _4213_ (.A(net107),
    .B(_2666_),
    .Y(_1115_));
 sg13g2_nand2_1 _4214_ (.Y(_1116_),
    .A(net106),
    .B(_0027_));
 sg13g2_o21ai_1 _4215_ (.B1(_1116_),
    .Y(_1117_),
    .A1(net68),
    .A2(_0778_));
 sg13g2_a22oi_1 _4216_ (.Y(_1118_),
    .B1(_1117_),
    .B2(net107),
    .A2(_1115_),
    .A1(_0088_));
 sg13g2_nand3_1 _4217_ (.B(_2722_),
    .C(\game.fsm.block_len[7][2] ),
    .A(_2666_),
    .Y(_1119_));
 sg13g2_nand3_1 _4218_ (.B(_0752_),
    .C(_1073_),
    .A(net68),
    .Y(_1120_));
 sg13g2_a21oi_1 _4219_ (.A1(_1119_),
    .A2(_1120_),
    .Y(_1121_),
    .B1(net64));
 sg13g2_a221oi_1 _4220_ (.B2(_1118_),
    .C1(_1121_),
    .B1(_1114_),
    .A1(net64),
    .Y(_1122_),
    .A2(_1111_));
 sg13g2_buf_1 _4221_ (.A(_1122_),
    .X(_1123_));
 sg13g2_nor2_2 _4222_ (.A(net37),
    .B(_1030_),
    .Y(_1124_));
 sg13g2_inv_1 _4223_ (.Y(_1125_),
    .A(_1098_));
 sg13g2_nor2_1 _4224_ (.A(_1066_),
    .B(_1095_),
    .Y(_1126_));
 sg13g2_a22oi_1 _4225_ (.Y(_1127_),
    .B1(_1126_),
    .B2(net39),
    .A2(_1125_),
    .A1(_1124_));
 sg13g2_a221oi_1 _4226_ (.B2(_1124_),
    .C1(_1123_),
    .B1(_1098_),
    .A1(_1103_),
    .Y(_1128_),
    .A2(_1096_));
 sg13g2_a21oi_1 _4227_ (.A1(_1123_),
    .A2(_1127_),
    .Y(_1129_),
    .B1(_1128_));
 sg13g2_and2_1 _4228_ (.A(net45),
    .B(_1129_),
    .X(_1130_));
 sg13g2_buf_2 _4229_ (.A(_1130_),
    .X(_1131_));
 sg13g2_buf_1 _4230_ (.A(net46),
    .X(_1132_));
 sg13g2_nor2_1 _4231_ (.A(_2711_),
    .B(net35),
    .Y(_1133_));
 sg13g2_mux2_1 _4232_ (.A0(_1131_),
    .A1(_1133_),
    .S(_1084_),
    .X(_0174_));
 sg13g2_nor2_1 _4233_ (.A(_0642_),
    .B(net35),
    .Y(_1134_));
 sg13g2_a21o_1 _4234_ (.A2(_1068_),
    .A1(_1066_),
    .B1(net64),
    .X(_1135_));
 sg13g2_nand3_1 _4235_ (.B(_1042_),
    .C(_1030_),
    .A(_1079_),
    .Y(_1136_));
 sg13g2_nand3_1 _4236_ (.B(_1135_),
    .C(_1136_),
    .A(_1056_),
    .Y(_1137_));
 sg13g2_buf_1 _4237_ (.A(_1137_),
    .X(_1138_));
 sg13g2_nand2b_1 _4238_ (.Y(_1139_),
    .B(_1138_),
    .A_N(_1078_));
 sg13g2_buf_1 _4239_ (.A(_1139_),
    .X(_1140_));
 sg13g2_mux2_1 _4240_ (.A0(_1054_),
    .A1(_1134_),
    .S(_1140_),
    .X(_0175_));
 sg13g2_nand3_1 _4241_ (.B(net36),
    .C(_1140_),
    .A(_2712_),
    .Y(_1141_));
 sg13g2_o21ai_1 _4242_ (.B1(_1141_),
    .Y(_0176_),
    .A1(_1106_),
    .A2(_1140_));
 sg13g2_and2_1 _4243_ (.A(_2709_),
    .B(net38),
    .X(_1142_));
 sg13g2_mux2_1 _4244_ (.A0(_1131_),
    .A1(_1142_),
    .S(_1140_),
    .X(_0177_));
 sg13g2_and2_1 _4245_ (.A(_2879_),
    .B(net38),
    .X(_1143_));
 sg13g2_nand3_1 _4246_ (.B(_1077_),
    .C(_1072_),
    .A(_1082_),
    .Y(_1144_));
 sg13g2_buf_1 _4247_ (.A(_1144_),
    .X(_1145_));
 sg13g2_mux2_1 _4248_ (.A0(_1054_),
    .A1(_1143_),
    .S(_1145_),
    .X(_0178_));
 sg13g2_nand3_1 _4249_ (.B(net36),
    .C(_1145_),
    .A(_2875_),
    .Y(_1146_));
 sg13g2_o21ai_1 _4250_ (.B1(_1146_),
    .Y(_0179_),
    .A1(_1106_),
    .A2(_1145_));
 sg13g2_and2_1 _4251_ (.A(_2724_),
    .B(net38),
    .X(_1147_));
 sg13g2_mux2_1 _4252_ (.A0(_1131_),
    .A1(_1147_),
    .S(_1145_),
    .X(_0180_));
 sg13g2_buf_1 _4253_ (.A(net45),
    .X(_1148_));
 sg13g2_and2_1 _4254_ (.A(_2878_),
    .B(net34),
    .X(_1149_));
 sg13g2_nand3_1 _4255_ (.B(_1072_),
    .C(_1138_),
    .A(_1077_),
    .Y(_1150_));
 sg13g2_buf_1 _4256_ (.A(_1150_),
    .X(_1151_));
 sg13g2_mux2_1 _4257_ (.A0(_1054_),
    .A1(_1149_),
    .S(_1151_),
    .X(_0181_));
 sg13g2_nand3_1 _4258_ (.B(net36),
    .C(_1151_),
    .A(_2876_),
    .Y(_1152_));
 sg13g2_o21ai_1 _4259_ (.B1(_1152_),
    .Y(_0182_),
    .A1(_1106_),
    .A2(_1151_));
 sg13g2_nor2_1 _4260_ (.A(_2874_),
    .B(net35),
    .Y(_1153_));
 sg13g2_mux2_1 _4261_ (.A0(_1131_),
    .A1(_1153_),
    .S(_1151_),
    .X(_0183_));
 sg13g2_nor2_1 _4262_ (.A(_2651_),
    .B(net35),
    .Y(_1154_));
 sg13g2_nor2_1 _4263_ (.A(_1077_),
    .B(_1072_),
    .Y(_1155_));
 sg13g2_nand2_2 _4264_ (.Y(_1156_),
    .A(_1082_),
    .B(_1155_));
 sg13g2_mux2_1 _4265_ (.A0(_1054_),
    .A1(_1154_),
    .S(_1156_),
    .X(_0184_));
 sg13g2_nand3_1 _4266_ (.B(net36),
    .C(_1156_),
    .A(_2655_),
    .Y(_1157_));
 sg13g2_o21ai_1 _4267_ (.B1(_1157_),
    .Y(_0185_),
    .A1(_1106_),
    .A2(_1156_));
 sg13g2_and2_1 _4268_ (.A(net133),
    .B(net34),
    .X(_1158_));
 sg13g2_mux2_1 _4269_ (.A0(_1131_),
    .A1(_1158_),
    .S(_1156_),
    .X(_0186_));
 sg13g2_nand2_2 _4270_ (.Y(_1159_),
    .A(_1138_),
    .B(_1155_));
 sg13g2_mux2_1 _4271_ (.A0(_1054_),
    .A1(\game.fsm.block_len[5][0] ),
    .S(_1159_),
    .X(_0187_));
 sg13g2_and2_1 _4272_ (.A(net45),
    .B(_1105_),
    .X(_1160_));
 sg13g2_mux2_1 _4273_ (.A0(_1160_),
    .A1(_2656_),
    .S(_1159_),
    .X(_0188_));
 sg13g2_mux2_1 _4274_ (.A0(_1131_),
    .A1(_2653_),
    .S(_1159_),
    .X(_0189_));
 sg13g2_nand3b_1 _4275_ (.B(_1072_),
    .C(_1138_),
    .Y(_1161_),
    .A_N(_1077_));
 sg13g2_buf_1 _4276_ (.A(_1161_),
    .X(_1162_));
 sg13g2_mux2_1 _4277_ (.A0(_1054_),
    .A1(\game.fsm.block_len[7][0] ),
    .S(_1162_),
    .X(_0193_));
 sg13g2_mux2_1 _4278_ (.A0(_1160_),
    .A1(\game.fsm.block_len[7][1] ),
    .S(_1162_),
    .X(_0194_));
 sg13g2_mux2_1 _4279_ (.A0(_1131_),
    .A1(\game.fsm.block_len[7][2] ),
    .S(_1162_),
    .X(_0195_));
 sg13g2_nand2_1 _4280_ (.Y(_1163_),
    .A(_1056_),
    .B(_1042_));
 sg13g2_buf_2 _4281_ (.A(_1163_),
    .X(_1164_));
 sg13g2_nor2_1 _4282_ (.A(_1026_),
    .B(_1164_),
    .Y(_1165_));
 sg13g2_a21oi_1 _4283_ (.A1(_0456_),
    .A2(_1164_),
    .Y(_1166_),
    .B1(_1165_));
 sg13g2_buf_4 _4284_ (.X(_1167_),
    .A(_1166_));
 sg13g2_and2_1 _4285_ (.A(_1020_),
    .B(_1063_),
    .X(_1168_));
 sg13g2_a21oi_1 _4286_ (.A1(_1015_),
    .A2(_1164_),
    .Y(_1169_),
    .B1(_1168_));
 sg13g2_buf_4 _4287_ (.X(_1170_),
    .A(_1169_));
 sg13g2_mux4_1 _4288_ (.S0(_1167_),
    .A0(_0541_),
    .A1(_0550_),
    .A2(_0510_),
    .A3(_0613_),
    .S1(_1170_),
    .X(_1171_));
 sg13g2_buf_1 _4289_ (.A(_1171_),
    .X(_1172_));
 sg13g2_inv_1 _4290_ (.Y(_1173_),
    .A(_1172_));
 sg13g2_nor2_1 _4291_ (.A(_1043_),
    .B(_1047_),
    .Y(_1174_));
 sg13g2_nor3_2 _4292_ (.A(_1052_),
    .B(_1173_),
    .C(_1174_),
    .Y(_1175_));
 sg13g2_nor2_1 _4293_ (.A(_0541_),
    .B(net35),
    .Y(_1176_));
 sg13g2_nor2_1 _4294_ (.A(_1051_),
    .B(_1066_),
    .Y(_1177_));
 sg13g2_buf_1 _4295_ (.A(_1177_),
    .X(_1178_));
 sg13g2_a21oi_2 _4296_ (.B1(_1168_),
    .Y(_1179_),
    .A2(_1178_),
    .A1(net29));
 sg13g2_a21oi_2 _4297_ (.B1(_1024_),
    .Y(_1180_),
    .A2(\game.slv.fsm_color[1] ),
    .A1(net93));
 sg13g2_a22oi_1 _4298_ (.Y(_1181_),
    .B1(_1103_),
    .B2(_0456_),
    .A2(_1180_),
    .A1(_1042_));
 sg13g2_nor2_1 _4299_ (.A(_1051_),
    .B(_1181_),
    .Y(_1182_));
 sg13g2_nand2b_1 _4300_ (.Y(_1183_),
    .B(_1182_),
    .A_N(_1179_));
 sg13g2_buf_1 _4301_ (.A(_1183_),
    .X(_1184_));
 sg13g2_mux2_1 _4302_ (.A0(_1175_),
    .A1(_1176_),
    .S(_1184_),
    .X(_0196_));
 sg13g2_mux4_1 _4303_ (.S0(_1167_),
    .A0(net98),
    .A1(_0601_),
    .A2(_0509_),
    .A3(_0626_),
    .S1(_1170_),
    .X(_1185_));
 sg13g2_buf_1 _4304_ (.A(_1185_),
    .X(_1186_));
 sg13g2_xnor2_1 _4305_ (.Y(_1187_),
    .A(_1172_),
    .B(_1186_));
 sg13g2_nand2_1 _4306_ (.Y(_1188_),
    .A(net22),
    .B(_1187_));
 sg13g2_o21ai_1 _4307_ (.B1(_1188_),
    .Y(_1189_),
    .A1(_1164_),
    .A2(_1187_));
 sg13g2_nor2_1 _4308_ (.A(net98),
    .B(net46),
    .Y(_1190_));
 sg13g2_mux2_1 _4309_ (.A0(_1189_),
    .A1(_1190_),
    .S(_1184_),
    .X(_0197_));
 sg13g2_inv_1 _4310_ (.Y(_1191_),
    .A(_0072_));
 sg13g2_inv_1 _4311_ (.Y(_1192_),
    .A(_0071_));
 sg13g2_mux4_1 _4312_ (.S0(_1167_),
    .A0(net97),
    .A1(_1191_),
    .A2(net122),
    .A3(_1192_),
    .S1(_1170_),
    .X(_1193_));
 sg13g2_buf_1 _4313_ (.A(_1193_),
    .X(_1194_));
 sg13g2_nor3_1 _4314_ (.A(_1172_),
    .B(_1186_),
    .C(_1194_),
    .Y(_1195_));
 sg13g2_a21o_1 _4315_ (.A2(_1194_),
    .A1(_1186_),
    .B1(_1195_),
    .X(_1196_));
 sg13g2_nand2_1 _4316_ (.Y(_1197_),
    .A(net22),
    .B(_1186_));
 sg13g2_nand2_1 _4317_ (.Y(_1198_),
    .A(_1063_),
    .B(_1194_));
 sg13g2_o21ai_1 _4318_ (.B1(_1198_),
    .Y(_1199_),
    .A1(_1194_),
    .A2(_1197_));
 sg13g2_nand2_1 _4319_ (.Y(_1200_),
    .A(_1178_),
    .B(_1194_));
 sg13g2_a21oi_1 _4320_ (.A1(_1172_),
    .A2(_1186_),
    .Y(_1201_),
    .B1(_1200_));
 sg13g2_a221oi_1 _4321_ (.B2(_1172_),
    .C1(_1201_),
    .B1(_1199_),
    .A1(_1063_),
    .Y(_1202_),
    .A2(_1196_));
 sg13g2_buf_1 _4322_ (.A(_1202_),
    .X(_1203_));
 sg13g2_nand3_1 _4323_ (.B(net36),
    .C(_1184_),
    .A(net97),
    .Y(_1204_));
 sg13g2_o21ai_1 _4324_ (.B1(_1204_),
    .Y(_0198_),
    .A1(_1184_),
    .A2(_1203_));
 sg13g2_nor2_1 _4325_ (.A(_0510_),
    .B(net46),
    .Y(_1205_));
 sg13g2_nand2_2 _4326_ (.Y(_1206_),
    .A(_1179_),
    .B(_1182_));
 sg13g2_mux2_1 _4327_ (.A0(_1175_),
    .A1(_1205_),
    .S(_1206_),
    .X(_0199_));
 sg13g2_nor2_1 _4328_ (.A(_0509_),
    .B(net46),
    .Y(_1207_));
 sg13g2_mux2_1 _4329_ (.A0(_1189_),
    .A1(_1207_),
    .S(_1206_),
    .X(_0200_));
 sg13g2_nand3_1 _4330_ (.B(net36),
    .C(_1206_),
    .A(_0571_),
    .Y(_1208_));
 sg13g2_o21ai_1 _4331_ (.B1(_1208_),
    .Y(_0201_),
    .A1(_1203_),
    .A2(_1206_));
 sg13g2_nor2_1 _4332_ (.A(_0550_),
    .B(net46),
    .Y(_1209_));
 sg13g2_a21oi_1 _4333_ (.A1(_1056_),
    .A2(_1174_),
    .Y(_1210_),
    .B1(_1182_));
 sg13g2_nand2b_1 _4334_ (.Y(_1211_),
    .B(_1210_),
    .A_N(_1179_));
 sg13g2_buf_1 _4335_ (.A(_1211_),
    .X(_1212_));
 sg13g2_mux2_1 _4336_ (.A0(_1175_),
    .A1(_1209_),
    .S(_1212_),
    .X(_0202_));
 sg13g2_nor2_1 _4337_ (.A(_0601_),
    .B(net46),
    .Y(_1213_));
 sg13g2_mux2_1 _4338_ (.A0(_1189_),
    .A1(_1213_),
    .S(_1212_),
    .X(_0203_));
 sg13g2_buf_1 _4339_ (.A(_1057_),
    .X(_1214_));
 sg13g2_nand3_1 _4340_ (.B(_1214_),
    .C(_1212_),
    .A(net124),
    .Y(_1215_));
 sg13g2_o21ai_1 _4341_ (.B1(_1215_),
    .Y(_0204_),
    .A1(_1203_),
    .A2(_1212_));
 sg13g2_nand2_2 _4342_ (.Y(_1216_),
    .A(_1179_),
    .B(_1210_));
 sg13g2_mux2_1 _4343_ (.A0(_1175_),
    .A1(net125),
    .S(_1216_),
    .X(_0205_));
 sg13g2_nor2_1 _4344_ (.A(_1189_),
    .B(_1216_),
    .Y(_1217_));
 sg13g2_a21oi_1 _4345_ (.A1(_0626_),
    .A2(_1216_),
    .Y(_0206_),
    .B1(_1217_));
 sg13g2_nand2_1 _4346_ (.Y(_1218_),
    .A(net123),
    .B(_1216_));
 sg13g2_o21ai_1 _4347_ (.B1(_1218_),
    .Y(_0207_),
    .A1(_1203_),
    .A2(_1216_));
 sg13g2_nand2_1 _4348_ (.Y(_1219_),
    .A(_1097_),
    .B(_1123_));
 sg13g2_or2_1 _4349_ (.X(_1220_),
    .B(_1219_),
    .A(_1095_));
 sg13g2_buf_1 _4350_ (.A(_1220_),
    .X(_1221_));
 sg13g2_nand2b_1 _4351_ (.Y(_1222_),
    .B(_1221_),
    .A_N(_1030_));
 sg13g2_nor2b_1 _4352_ (.A(_1099_),
    .B_N(_1123_),
    .Y(_1223_));
 sg13g2_a22oi_1 _4353_ (.Y(_1224_),
    .B1(_1223_),
    .B2(_1103_),
    .A2(_1222_),
    .A1(_1042_));
 sg13g2_buf_1 _4354_ (.A(_1224_),
    .X(_1225_));
 sg13g2_mux4_1 _4355_ (.S0(_1170_),
    .A0(\game.fsm.len1_color_count[0][0] ),
    .A1(\game.fsm.len1_color_count[1][0] ),
    .A2(\game.fsm.len1_color_count[2][0] ),
    .A3(\game.fsm.len1_color_count[3][0] ),
    .S1(_1167_),
    .X(_1226_));
 sg13g2_nor3_2 _4356_ (.A(_1052_),
    .B(_1225_),
    .C(_1226_),
    .Y(_1227_));
 sg13g2_and2_1 _4357_ (.A(\game.fsm.len1_color_count[0][0] ),
    .B(net34),
    .X(_1228_));
 sg13g2_inv_1 _4358_ (.Y(_1229_),
    .A(net29));
 sg13g2_nand2_1 _4359_ (.Y(_1230_),
    .A(net22),
    .B(_1223_));
 sg13g2_and2_1 _4360_ (.A(_1063_),
    .B(_1222_),
    .X(_1231_));
 sg13g2_buf_1 _4361_ (.A(_1231_),
    .X(_1232_));
 sg13g2_nand2_1 _4362_ (.Y(_1233_),
    .A(_1020_),
    .B(_1232_));
 sg13g2_o21ai_1 _4363_ (.B1(_1233_),
    .Y(_1234_),
    .A1(_1229_),
    .A2(_1230_));
 sg13g2_buf_1 _4364_ (.A(_1234_),
    .X(_1235_));
 sg13g2_inv_2 _4365_ (.Y(_1236_),
    .A(_0456_));
 sg13g2_nand2_1 _4366_ (.Y(_1237_),
    .A(_1180_),
    .B(_1232_));
 sg13g2_o21ai_1 _4367_ (.B1(_1237_),
    .Y(_1238_),
    .A1(_1236_),
    .A2(_1230_));
 sg13g2_nand2_2 _4368_ (.Y(_1239_),
    .A(_1235_),
    .B(_1238_));
 sg13g2_mux2_1 _4369_ (.A0(_1227_),
    .A1(_1228_),
    .S(_1239_),
    .X(_0214_));
 sg13g2_mux4_1 _4370_ (.S0(_1167_),
    .A0(_0040_),
    .A1(_0042_),
    .A2(_0041_),
    .A3(_0043_),
    .S1(_1170_),
    .X(_1240_));
 sg13g2_nand2b_1 _4371_ (.Y(_1241_),
    .B(_1226_),
    .A_N(_1240_));
 sg13g2_nand2b_1 _4372_ (.Y(_1242_),
    .B(_1240_),
    .A_N(_1226_));
 sg13g2_nand2_1 _4373_ (.Y(_1243_),
    .A(_1241_),
    .B(_1242_));
 sg13g2_and2_1 _4374_ (.A(_1095_),
    .B(_1123_),
    .X(_1244_));
 sg13g2_buf_1 _4375_ (.A(_1244_),
    .X(_1245_));
 sg13g2_and2_1 _4376_ (.A(net39),
    .B(net26),
    .X(_1246_));
 sg13g2_buf_1 _4377_ (.A(_1246_),
    .X(_1247_));
 sg13g2_xnor2_1 _4378_ (.Y(_1248_),
    .A(_1243_),
    .B(_1247_));
 sg13g2_nor2_1 _4379_ (.A(_1030_),
    .B(_1221_),
    .Y(_1249_));
 sg13g2_mux2_1 _4380_ (.A0(_1030_),
    .A1(_1249_),
    .S(_1243_),
    .X(_1250_));
 sg13g2_nand2_1 _4381_ (.Y(_1251_),
    .A(_1063_),
    .B(_1250_));
 sg13g2_o21ai_1 _4382_ (.B1(_1251_),
    .Y(_1252_),
    .A1(_1230_),
    .A2(_1248_));
 sg13g2_buf_1 _4383_ (.A(_1252_),
    .X(_1253_));
 sg13g2_nand2b_1 _4384_ (.Y(_1254_),
    .B(_1253_),
    .A_N(_1239_));
 sg13g2_buf_1 _4385_ (.A(net45),
    .X(_1255_));
 sg13g2_nand3_1 _4386_ (.B(net32),
    .C(_1239_),
    .A(\game.fsm.len1_color_count[0][1] ),
    .Y(_1256_));
 sg13g2_nand2_1 _4387_ (.Y(_0215_),
    .A(_1254_),
    .B(_1256_));
 sg13g2_mux4_1 _4388_ (.S0(_1170_),
    .A0(_0022_),
    .A1(_0023_),
    .A2(_0025_),
    .A3(_0024_),
    .S1(_1167_),
    .X(_1257_));
 sg13g2_nand2_1 _4389_ (.Y(_1258_),
    .A(_1036_),
    .B(_1245_));
 sg13g2_mux2_1 _4390_ (.A0(_1241_),
    .A1(_1242_),
    .S(_1258_),
    .X(_1259_));
 sg13g2_xnor2_1 _4391_ (.Y(_1260_),
    .A(_1257_),
    .B(_1259_));
 sg13g2_nand2_1 _4392_ (.Y(_1261_),
    .A(_1056_),
    .B(_1124_));
 sg13g2_nor2_1 _4393_ (.A(_1221_),
    .B(_1261_),
    .Y(_1262_));
 sg13g2_mux2_1 _4394_ (.A0(_1241_),
    .A1(_1242_),
    .S(_1262_),
    .X(_1263_));
 sg13g2_xor2_1 _4395_ (.B(_1263_),
    .A(_1257_),
    .X(_1264_));
 sg13g2_nand2_1 _4396_ (.Y(_1265_),
    .A(_1232_),
    .B(_1264_));
 sg13g2_o21ai_1 _4397_ (.B1(_1265_),
    .Y(_1266_),
    .A1(_1230_),
    .A2(_1260_));
 sg13g2_buf_1 _4398_ (.A(_1266_),
    .X(_1267_));
 sg13g2_nand2b_1 _4399_ (.Y(_1268_),
    .B(_1267_),
    .A_N(_1239_));
 sg13g2_nand3_1 _4400_ (.B(net32),
    .C(_1239_),
    .A(\game.fsm.len1_color_count[0][2] ),
    .Y(_1269_));
 sg13g2_nand2_1 _4401_ (.Y(_0216_),
    .A(_1268_),
    .B(_1269_));
 sg13g2_and2_1 _4402_ (.A(\game.fsm.len1_color_count[1][0] ),
    .B(net34),
    .X(_1270_));
 sg13g2_nand2b_1 _4403_ (.Y(_1271_),
    .B(_1238_),
    .A_N(_1235_));
 sg13g2_buf_1 _4404_ (.A(_1271_),
    .X(_1272_));
 sg13g2_mux2_1 _4405_ (.A0(_1227_),
    .A1(_1270_),
    .S(_1272_),
    .X(_0217_));
 sg13g2_nand2b_1 _4406_ (.Y(_1273_),
    .B(_1253_),
    .A_N(_1272_));
 sg13g2_nand3_1 _4407_ (.B(net32),
    .C(_1272_),
    .A(\game.fsm.len1_color_count[1][1] ),
    .Y(_1274_));
 sg13g2_nand2_1 _4408_ (.Y(_0218_),
    .A(_1273_),
    .B(_1274_));
 sg13g2_nand2b_1 _4409_ (.Y(_1275_),
    .B(_1267_),
    .A_N(_1272_));
 sg13g2_nand3_1 _4410_ (.B(net32),
    .C(_1272_),
    .A(\game.fsm.len1_color_count[1][2] ),
    .Y(_1276_));
 sg13g2_nand2_1 _4411_ (.Y(_0219_),
    .A(_1275_),
    .B(_1276_));
 sg13g2_a21oi_1 _4412_ (.A1(_1056_),
    .A2(_1225_),
    .Y(_1277_),
    .B1(_1238_));
 sg13g2_and2_1 _4413_ (.A(_1235_),
    .B(_1277_),
    .X(_1278_));
 sg13g2_buf_1 _4414_ (.A(_1278_),
    .X(_1279_));
 sg13g2_nand2_1 _4415_ (.Y(_1280_),
    .A(\game.fsm.len1_color_count[2][0] ),
    .B(net38));
 sg13g2_nand2_1 _4416_ (.Y(_1281_),
    .A(_1227_),
    .B(_1279_));
 sg13g2_o21ai_1 _4417_ (.B1(_1281_),
    .Y(_0220_),
    .A1(_1279_),
    .A2(_1280_));
 sg13g2_nand2_1 _4418_ (.Y(_1282_),
    .A(\game.fsm.len1_color_count[2][1] ),
    .B(_1058_));
 sg13g2_nand2_1 _4419_ (.Y(_1283_),
    .A(_1253_),
    .B(_1279_));
 sg13g2_o21ai_1 _4420_ (.B1(_1283_),
    .Y(_0221_),
    .A1(_1279_),
    .A2(_1282_));
 sg13g2_nand2_1 _4421_ (.Y(_1284_),
    .A(\game.fsm.len1_color_count[2][2] ),
    .B(net38));
 sg13g2_nand2_1 _4422_ (.Y(_1285_),
    .A(_1267_),
    .B(_1279_));
 sg13g2_o21ai_1 _4423_ (.B1(_1285_),
    .Y(_0222_),
    .A1(_1279_),
    .A2(_1284_));
 sg13g2_nor2b_2 _4424_ (.A(_1235_),
    .B_N(_1277_),
    .Y(_1286_));
 sg13g2_mux2_1 _4425_ (.A0(\game.fsm.len1_color_count[3][0] ),
    .A1(_1227_),
    .S(_1286_),
    .X(_0223_));
 sg13g2_mux2_1 _4426_ (.A0(\game.fsm.len1_color_count[3][1] ),
    .A1(_1253_),
    .S(_1286_),
    .X(_0224_));
 sg13g2_mux2_1 _4427_ (.A0(\game.fsm.len1_color_count[3][2] ),
    .A1(_1267_),
    .S(_1286_),
    .X(_0225_));
 sg13g2_mux4_1 _4428_ (.S0(_1236_),
    .A0(\game.fsm.len2_color_count[1][0] ),
    .A1(\game.fsm.len2_color_count[3][0] ),
    .A2(\game.fsm.len2_color_count[0][0] ),
    .A3(\game.fsm.len2_color_count[2][0] ),
    .S1(net29),
    .X(_1287_));
 sg13g2_nor2_1 _4429_ (.A(_1051_),
    .B(_1068_),
    .Y(_1288_));
 sg13g2_and2_1 _4430_ (.A(_1223_),
    .B(_1288_),
    .X(_1289_));
 sg13g2_buf_1 _4431_ (.A(_1289_),
    .X(_1290_));
 sg13g2_and2_1 _4432_ (.A(net22),
    .B(net26),
    .X(_1291_));
 sg13g2_nor2_1 _4433_ (.A(_1290_),
    .B(_1291_),
    .Y(_1292_));
 sg13g2_nor2_1 _4434_ (.A(_1287_),
    .B(_1292_),
    .Y(_1293_));
 sg13g2_and2_1 _4435_ (.A(\game.fsm.len2_color_count[0][0] ),
    .B(net34),
    .X(_1294_));
 sg13g2_nand2_1 _4436_ (.Y(_1295_),
    .A(_1177_),
    .B(_1244_));
 sg13g2_nand2_1 _4437_ (.Y(_1296_),
    .A(_1180_),
    .B(_1290_));
 sg13g2_o21ai_1 _4438_ (.B1(_1296_),
    .Y(_1297_),
    .A1(_1236_),
    .A2(_1295_));
 sg13g2_buf_1 _4439_ (.A(_1297_),
    .X(_1298_));
 sg13g2_nand2_1 _4440_ (.Y(_1299_),
    .A(_1020_),
    .B(_1290_));
 sg13g2_o21ai_1 _4441_ (.B1(_1299_),
    .Y(_1300_),
    .A1(_1229_),
    .A2(_1295_));
 sg13g2_buf_1 _4442_ (.A(_1300_),
    .X(_1301_));
 sg13g2_nand2_1 _4443_ (.Y(_1302_),
    .A(_1298_),
    .B(_1301_));
 sg13g2_mux2_1 _4444_ (.A0(_1293_),
    .A1(_1294_),
    .S(_1302_),
    .X(_0228_));
 sg13g2_mux4_1 _4445_ (.S0(net29),
    .A0(_0045_),
    .A1(_0044_),
    .A2(_0047_),
    .A3(_0046_),
    .S1(_1236_),
    .X(_1303_));
 sg13g2_xor2_1 _4446_ (.B(_1303_),
    .A(_1287_),
    .X(_1304_));
 sg13g2_nor2_1 _4447_ (.A(net39),
    .B(_1304_),
    .Y(_1305_));
 sg13g2_o21ai_1 _4448_ (.B1(_1305_),
    .Y(_1306_),
    .A1(_1262_),
    .A2(_1291_));
 sg13g2_nand3_1 _4449_ (.B(_1247_),
    .C(_1304_),
    .A(_1069_),
    .Y(_1307_));
 sg13g2_nand2_1 _4450_ (.Y(_1308_),
    .A(_1306_),
    .B(_1307_));
 sg13g2_nand3_1 _4451_ (.B(_1301_),
    .C(_1308_),
    .A(_1298_),
    .Y(_1309_));
 sg13g2_nand3_1 _4452_ (.B(net32),
    .C(_1302_),
    .A(\game.fsm.len2_color_count[0][1] ),
    .Y(_1310_));
 sg13g2_nand2_1 _4453_ (.Y(_0229_),
    .A(_1309_),
    .B(_1310_));
 sg13g2_and2_1 _4454_ (.A(\game.fsm.len2_color_count[1][0] ),
    .B(net34),
    .X(_1311_));
 sg13g2_nand2b_1 _4455_ (.Y(_1312_),
    .B(_1298_),
    .A_N(_1301_));
 sg13g2_mux2_1 _4456_ (.A0(_1293_),
    .A1(_1311_),
    .S(_1312_),
    .X(_0230_));
 sg13g2_nand2b_1 _4457_ (.Y(_1313_),
    .B(_1308_),
    .A_N(_1312_));
 sg13g2_nand3_1 _4458_ (.B(net32),
    .C(_1312_),
    .A(\game.fsm.len2_color_count[1][1] ),
    .Y(_1314_));
 sg13g2_nand2_1 _4459_ (.Y(_0231_),
    .A(_1313_),
    .B(_1314_));
 sg13g2_and2_1 _4460_ (.A(\game.fsm.len2_color_count[2][0] ),
    .B(net34),
    .X(_1315_));
 sg13g2_a21oi_1 _4461_ (.A1(net45),
    .A2(_1292_),
    .Y(_1316_),
    .B1(_1298_));
 sg13g2_nand2_1 _4462_ (.Y(_1317_),
    .A(_1301_),
    .B(_1316_));
 sg13g2_mux2_1 _4463_ (.A0(_1293_),
    .A1(_1315_),
    .S(_1317_),
    .X(_0232_));
 sg13g2_nand3_1 _4464_ (.B(_1308_),
    .C(_1316_),
    .A(_1301_),
    .Y(_1318_));
 sg13g2_nand3_1 _4465_ (.B(net32),
    .C(_1317_),
    .A(\game.fsm.len2_color_count[2][1] ),
    .Y(_1319_));
 sg13g2_nand2_1 _4466_ (.Y(_0233_),
    .A(_1318_),
    .B(_1319_));
 sg13g2_nor2b_1 _4467_ (.A(_1301_),
    .B_N(_1316_),
    .Y(_1320_));
 sg13g2_mux2_1 _4468_ (.A0(\game.fsm.len2_color_count[3][0] ),
    .A1(_1293_),
    .S(_1320_),
    .X(_0234_));
 sg13g2_mux2_1 _4469_ (.A0(\game.fsm.len2_color_count[3][1] ),
    .A1(_1308_),
    .S(_1320_),
    .X(_0235_));
 sg13g2_nor2_1 _4470_ (.A(_1096_),
    .B(_1123_),
    .Y(_1321_));
 sg13g2_nand2_1 _4471_ (.Y(_1322_),
    .A(_1177_),
    .B(_1321_));
 sg13g2_o21ai_1 _4472_ (.B1(_1322_),
    .Y(_1323_),
    .A1(net39),
    .A2(_1295_));
 sg13g2_buf_1 _4473_ (.A(_1323_),
    .X(_1324_));
 sg13g2_inv_1 _4474_ (.Y(_1325_),
    .A(_1324_));
 sg13g2_nand2_1 _4475_ (.Y(_1326_),
    .A(net26),
    .B(_1288_));
 sg13g2_mux4_1 _4476_ (.S0(net29),
    .A0(\game.fsm.len3_color_count[1][0] ),
    .A1(\game.fsm.len3_color_count[0][0] ),
    .A2(\game.fsm.len3_color_count[3][0] ),
    .A3(\game.fsm.len3_color_count[2][0] ),
    .S1(_1236_),
    .X(_1327_));
 sg13g2_a21oi_2 _4477_ (.B1(_1327_),
    .Y(_1328_),
    .A2(_1326_),
    .A1(_1325_));
 sg13g2_and2_1 _4478_ (.A(\game.fsm.len3_color_count[0][0] ),
    .B(net34),
    .X(_1329_));
 sg13g2_nand2_1 _4479_ (.Y(_1330_),
    .A(_0456_),
    .B(_1324_));
 sg13g2_o21ai_1 _4480_ (.B1(_1330_),
    .Y(_1331_),
    .A1(_1026_),
    .A2(_1326_));
 sg13g2_and4_1 _4481_ (.A(_1056_),
    .B(_1020_),
    .C(_1124_),
    .D(net26),
    .X(_1332_));
 sg13g2_a21o_1 _4482_ (.A2(_1324_),
    .A1(net29),
    .B1(_1332_),
    .X(_1333_));
 sg13g2_nand2_1 _4483_ (.Y(_1334_),
    .A(_1331_),
    .B(_1333_));
 sg13g2_mux2_1 _4484_ (.A0(_1328_),
    .A1(_1329_),
    .S(_1334_),
    .X(_0238_));
 sg13g2_mux4_1 _4485_ (.S0(net29),
    .A0(_0049_),
    .A1(_0048_),
    .A2(_0051_),
    .A3(_0050_),
    .S1(_1236_),
    .X(_1335_));
 sg13g2_xor2_1 _4486_ (.B(_1335_),
    .A(_1327_),
    .X(_1336_));
 sg13g2_nor3_1 _4487_ (.A(_1097_),
    .B(_1261_),
    .C(_1336_),
    .Y(_1337_));
 sg13g2_and3_1 _4488_ (.X(_1338_),
    .A(_1097_),
    .B(_1069_),
    .C(_1336_));
 sg13g2_o21ai_1 _4489_ (.B1(net26),
    .Y(_1339_),
    .A1(_1337_),
    .A2(_1338_));
 sg13g2_o21ai_1 _4490_ (.B1(_1339_),
    .Y(_1340_),
    .A1(_1322_),
    .A2(_1336_));
 sg13g2_buf_1 _4491_ (.A(_1340_),
    .X(_1341_));
 sg13g2_nand2b_1 _4492_ (.Y(_1342_),
    .B(_1341_),
    .A_N(_1334_));
 sg13g2_nand3_1 _4493_ (.B(_1107_),
    .C(_1334_),
    .A(\game.fsm.len3_color_count[0][1] ),
    .Y(_1343_));
 sg13g2_nand2_1 _4494_ (.Y(_0239_),
    .A(_1342_),
    .B(_1343_));
 sg13g2_and2_1 _4495_ (.A(\game.fsm.len3_color_count[1][0] ),
    .B(_1148_),
    .X(_1344_));
 sg13g2_a21oi_1 _4496_ (.A1(net29),
    .A2(_1324_),
    .Y(_1345_),
    .B1(_1332_));
 sg13g2_nand2_1 _4497_ (.Y(_1346_),
    .A(_1331_),
    .B(_1345_));
 sg13g2_mux2_1 _4498_ (.A0(_1328_),
    .A1(_1344_),
    .S(_1346_),
    .X(_0240_));
 sg13g2_nand2b_1 _4499_ (.Y(_1347_),
    .B(_1341_),
    .A_N(_1346_));
 sg13g2_nand3_1 _4500_ (.B(net36),
    .C(_1346_),
    .A(\game.fsm.len3_color_count[1][1] ),
    .Y(_1348_));
 sg13g2_nand2_1 _4501_ (.Y(_0241_),
    .A(_1347_),
    .B(_1348_));
 sg13g2_and2_1 _4502_ (.A(\game.fsm.len3_color_count[2][0] ),
    .B(_1148_),
    .X(_1349_));
 sg13g2_nand2_1 _4503_ (.Y(_1350_),
    .A(_1124_),
    .B(net26));
 sg13g2_mux2_1 _4504_ (.A0(_1180_),
    .A1(_1325_),
    .S(_1350_),
    .X(_1351_));
 sg13g2_a22oi_1 _4505_ (.Y(_1352_),
    .B1(_1351_),
    .B2(net45),
    .A2(_1324_),
    .A1(_0456_));
 sg13g2_nand2_1 _4506_ (.Y(_1353_),
    .A(_1333_),
    .B(_1352_));
 sg13g2_mux2_1 _4507_ (.A0(_1328_),
    .A1(_1349_),
    .S(_1353_),
    .X(_0242_));
 sg13g2_nand2b_1 _4508_ (.Y(_1354_),
    .B(_1341_),
    .A_N(_1353_));
 sg13g2_nand3_1 _4509_ (.B(_1107_),
    .C(_1353_),
    .A(\game.fsm.len3_color_count[2][1] ),
    .Y(_1355_));
 sg13g2_nand2_1 _4510_ (.Y(_0243_),
    .A(_1354_),
    .B(_1355_));
 sg13g2_nand2_1 _4511_ (.Y(_1356_),
    .A(_1345_),
    .B(_1352_));
 sg13g2_mux2_1 _4512_ (.A0(_1328_),
    .A1(\game.fsm.len3_color_count[3][0] ),
    .S(_1356_),
    .X(_0244_));
 sg13g2_mux2_1 _4513_ (.A0(_1341_),
    .A1(\game.fsm.len3_color_count[3][1] ),
    .S(_1356_),
    .X(_0245_));
 sg13g2_nor2_1 _4514_ (.A(_1020_),
    .B(_1164_),
    .Y(_1357_));
 sg13g2_inv_2 _4515_ (.Y(_1358_),
    .A(_1357_));
 sg13g2_nand2_1 _4516_ (.Y(_1359_),
    .A(net69),
    .B(net22));
 sg13g2_o21ai_1 _4517_ (.B1(_1359_),
    .Y(_1360_),
    .A1(net69),
    .A2(_1164_));
 sg13g2_buf_1 _4518_ (.A(_1360_),
    .X(_1361_));
 sg13g2_inv_1 _4519_ (.Y(_1362_),
    .A(_0068_));
 sg13g2_nand2b_1 _4520_ (.Y(_1363_),
    .B(_0421_),
    .A_N(_2929_));
 sg13g2_a22oi_1 _4521_ (.Y(_1364_),
    .B1(net22),
    .B2(_1363_),
    .A2(_1063_),
    .A1(_1362_));
 sg13g2_buf_1 _4522_ (.A(_1364_),
    .X(_1365_));
 sg13g2_a22oi_1 _4523_ (.Y(_1366_),
    .B1(net22),
    .B2(_0454_),
    .A2(_1063_),
    .A1(net72));
 sg13g2_buf_1 _4524_ (.A(_1366_),
    .X(_1367_));
 sg13g2_inv_1 _4525_ (.Y(_1368_),
    .A(_1367_));
 sg13g2_nand3_1 _4526_ (.B(_1365_),
    .C(_1368_),
    .A(_1361_),
    .Y(_1369_));
 sg13g2_buf_1 _4527_ (.A(_1369_),
    .X(_1370_));
 sg13g2_nand3_1 _4528_ (.B(net33),
    .C(_1370_),
    .A(_0419_),
    .Y(_1371_));
 sg13g2_o21ai_1 _4529_ (.B1(_1371_),
    .Y(_0252_),
    .A1(_1358_),
    .A2(_1370_));
 sg13g2_nor2_1 _4530_ (.A(_1180_),
    .B(_1164_),
    .Y(_1372_));
 sg13g2_inv_2 _4531_ (.Y(_1373_),
    .A(_1372_));
 sg13g2_nand3_1 _4532_ (.B(net33),
    .C(_1370_),
    .A(_0389_),
    .Y(_1374_));
 sg13g2_o21ai_1 _4533_ (.B1(_1374_),
    .Y(_0253_),
    .A1(_1370_),
    .A2(_1373_));
 sg13g2_nand2b_1 _4534_ (.Y(_1375_),
    .B(_1047_),
    .A_N(net48));
 sg13g2_nand2_1 _4535_ (.Y(_1376_),
    .A(net70),
    .B(_1375_));
 sg13g2_o21ai_1 _4536_ (.B1(_1376_),
    .Y(_1377_),
    .A1(net70),
    .A2(_1043_));
 sg13g2_nand2_1 _4537_ (.Y(_1378_),
    .A(_1056_),
    .B(_1377_));
 sg13g2_nand3_1 _4538_ (.B(_1368_),
    .C(_1378_),
    .A(_1365_),
    .Y(_1379_));
 sg13g2_buf_1 _4539_ (.A(_1379_),
    .X(_1380_));
 sg13g2_nand3_1 _4540_ (.B(net33),
    .C(_1380_),
    .A(\game.fsm.seq[1][0] ),
    .Y(_1381_));
 sg13g2_o21ai_1 _4541_ (.B1(_1381_),
    .Y(_0254_),
    .A1(_1358_),
    .A2(_1380_));
 sg13g2_nand3_1 _4542_ (.B(net33),
    .C(_1380_),
    .A(_2926_),
    .Y(_1382_));
 sg13g2_o21ai_1 _4543_ (.B1(_1382_),
    .Y(_0255_),
    .A1(_1373_),
    .A2(_1380_));
 sg13g2_nor2_1 _4544_ (.A(_1365_),
    .B(_1367_),
    .Y(_1383_));
 sg13g2_nand2_1 _4545_ (.Y(_1384_),
    .A(_1361_),
    .B(_1383_));
 sg13g2_nand3_1 _4546_ (.B(net33),
    .C(_1384_),
    .A(net126),
    .Y(_1385_));
 sg13g2_o21ai_1 _4547_ (.B1(_1385_),
    .Y(_0256_),
    .A1(_1358_),
    .A2(_1384_));
 sg13g2_nand3_1 _4548_ (.B(net33),
    .C(_1384_),
    .A(net127),
    .Y(_1386_));
 sg13g2_o21ai_1 _4549_ (.B1(_1386_),
    .Y(_0257_),
    .A1(_1373_),
    .A2(_1384_));
 sg13g2_nand2_1 _4550_ (.Y(_1387_),
    .A(_1378_),
    .B(_1383_));
 sg13g2_nand3_1 _4551_ (.B(net33),
    .C(_1387_),
    .A(_0416_),
    .Y(_1388_));
 sg13g2_o21ai_1 _4552_ (.B1(_1388_),
    .Y(_0258_),
    .A1(_1358_),
    .A2(_1387_));
 sg13g2_nand3_1 _4553_ (.B(_1214_),
    .C(_1387_),
    .A(_2932_),
    .Y(_1389_));
 sg13g2_o21ai_1 _4554_ (.B1(_1389_),
    .Y(_0259_),
    .A1(_1373_),
    .A2(_1387_));
 sg13g2_nand3_1 _4555_ (.B(_1365_),
    .C(_1367_),
    .A(_1361_),
    .Y(_1390_));
 sg13g2_buf_1 _4556_ (.A(_1390_),
    .X(_1391_));
 sg13g2_nand3_1 _4557_ (.B(net33),
    .C(_1391_),
    .A(_0426_),
    .Y(_1392_));
 sg13g2_o21ai_1 _4558_ (.B1(_1392_),
    .Y(_0260_),
    .A1(_1358_),
    .A2(_1391_));
 sg13g2_nand3_1 _4559_ (.B(_1058_),
    .C(_1391_),
    .A(_0404_),
    .Y(_1393_));
 sg13g2_o21ai_1 _4560_ (.B1(_1393_),
    .Y(_0261_),
    .A1(_1373_),
    .A2(_1391_));
 sg13g2_nand3_1 _4561_ (.B(_1367_),
    .C(_1378_),
    .A(_1365_),
    .Y(_1394_));
 sg13g2_buf_1 _4562_ (.A(_1394_),
    .X(_1395_));
 sg13g2_nand2_1 _4563_ (.Y(_1396_),
    .A(_0427_),
    .B(_1395_));
 sg13g2_o21ai_1 _4564_ (.B1(_1396_),
    .Y(_0262_),
    .A1(_1358_),
    .A2(_1395_));
 sg13g2_nand2_1 _4565_ (.Y(_1397_),
    .A(_0393_),
    .B(_1395_));
 sg13g2_o21ai_1 _4566_ (.B1(_1397_),
    .Y(_0263_),
    .A1(_1373_),
    .A2(_1395_));
 sg13g2_nand2_1 _4567_ (.Y(_1398_),
    .A(net22),
    .B(_1363_));
 sg13g2_o21ai_1 _4568_ (.B1(_1398_),
    .Y(_1399_),
    .A1(_0068_),
    .A2(_1164_));
 sg13g2_nand3_1 _4569_ (.B(_1367_),
    .C(_1378_),
    .A(_1399_),
    .Y(_1400_));
 sg13g2_buf_1 _4570_ (.A(_1400_),
    .X(_1401_));
 sg13g2_nand2_1 _4571_ (.Y(_1402_),
    .A(_0425_),
    .B(_1401_));
 sg13g2_o21ai_1 _4572_ (.B1(_1402_),
    .Y(_0266_),
    .A1(_1358_),
    .A2(_1401_));
 sg13g2_nand2_1 _4573_ (.Y(_1403_),
    .A(_0398_),
    .B(_1401_));
 sg13g2_o21ai_1 _4574_ (.B1(_1403_),
    .Y(_0267_),
    .A1(_1373_),
    .A2(_1401_));
 sg13g2_inv_1 _4575_ (.Y(_1404_),
    .A(_0094_));
 sg13g2_buf_1 _4576_ (.A(\clk_div_counter[2] ),
    .X(_1405_));
 sg13g2_inv_1 _4577_ (.Y(_1406_),
    .A(\clk_div_counter[7] ));
 sg13g2_buf_1 _4578_ (.A(\clk_div_counter[3] ),
    .X(_1407_));
 sg13g2_buf_1 _4579_ (.A(\clk_div_counter[5] ),
    .X(_1408_));
 sg13g2_nand4_1 _4580_ (.B(_1408_),
    .C(\clk_div_counter[4] ),
    .A(_1407_),
    .Y(_1409_),
    .D(\clk_div_counter[6] ));
 sg13g2_buf_1 _4581_ (.A(\clk_div_counter[1] ),
    .X(_1410_));
 sg13g2_buf_1 _4582_ (.A(\clk_div_counter[0] ),
    .X(_1411_));
 sg13g2_nand2b_1 _4583_ (.Y(_1412_),
    .B(_1411_),
    .A_N(_1410_));
 sg13g2_nor4_1 _4584_ (.A(_1405_),
    .B(_1406_),
    .C(_1409_),
    .D(_1412_),
    .Y(_1413_));
 sg13g2_nand2b_1 _4585_ (.Y(_1414_),
    .B(net134),
    .A_N(_1413_));
 sg13g2_buf_2 _4586_ (.A(_1414_),
    .X(_1415_));
 sg13g2_nor2_1 _4587_ (.A(_1404_),
    .B(_1415_),
    .Y(_0131_));
 sg13g2_nand2b_1 _4588_ (.Y(_1416_),
    .B(_1410_),
    .A_N(_1411_));
 sg13g2_a21oi_1 _4589_ (.A1(_1412_),
    .A2(_1416_),
    .Y(_0132_),
    .B1(_1415_));
 sg13g2_buf_1 _4590_ (.A(_2641_),
    .X(_1417_));
 sg13g2_buf_1 _4591_ (.A(net92),
    .X(_1418_));
 sg13g2_nand2_1 _4592_ (.Y(_1419_),
    .A(_1411_),
    .B(_1410_));
 sg13g2_xor2_1 _4593_ (.B(_1419_),
    .A(_1405_),
    .X(_1420_));
 sg13g2_nor2_1 _4594_ (.A(net63),
    .B(_1420_),
    .Y(_0133_));
 sg13g2_nand3_1 _4595_ (.B(_1410_),
    .C(_1405_),
    .A(_1411_),
    .Y(_1421_));
 sg13g2_xor2_1 _4596_ (.B(_1421_),
    .A(_1407_),
    .X(_1422_));
 sg13g2_nor2_1 _4597_ (.A(_1415_),
    .B(_1422_),
    .Y(_0134_));
 sg13g2_nand4_1 _4598_ (.B(_1410_),
    .C(_1405_),
    .A(_1411_),
    .Y(_1423_),
    .D(_1407_));
 sg13g2_xor2_1 _4599_ (.B(_1423_),
    .A(\clk_div_counter[4] ),
    .X(_1424_));
 sg13g2_nor2_1 _4600_ (.A(_1415_),
    .B(_1424_),
    .Y(_0135_));
 sg13g2_nand2_1 _4601_ (.Y(_1425_),
    .A(_1407_),
    .B(\clk_div_counter[4] ));
 sg13g2_nor2_1 _4602_ (.A(_1425_),
    .B(_1421_),
    .Y(_1426_));
 sg13g2_xnor2_1 _4603_ (.Y(_1427_),
    .A(_1408_),
    .B(_1426_));
 sg13g2_nor2_1 _4604_ (.A(_1415_),
    .B(_1427_),
    .Y(_0136_));
 sg13g2_nand2_1 _4605_ (.Y(_1428_),
    .A(_1408_),
    .B(_1426_));
 sg13g2_xor2_1 _4606_ (.B(_1428_),
    .A(\clk_div_counter[6] ),
    .X(_1429_));
 sg13g2_nor2_1 _4607_ (.A(_1415_),
    .B(_1429_),
    .Y(_0137_));
 sg13g2_nand3_1 _4608_ (.B(\clk_div_counter[6] ),
    .C(_1426_),
    .A(_1408_),
    .Y(_1430_));
 sg13g2_xnor2_1 _4609_ (.Y(_1431_),
    .A(_1406_),
    .B(_1430_));
 sg13g2_nor2_1 _4610_ (.A(_1415_),
    .B(_1431_),
    .Y(_0138_));
 sg13g2_nand3b_1 _4611_ (.B(_1072_),
    .C(_1082_),
    .Y(_1432_),
    .A_N(_1077_));
 sg13g2_buf_1 _4612_ (.A(_1432_),
    .X(_1433_));
 sg13g2_mux2_1 _4613_ (.A0(_1054_),
    .A1(\game.fsm.block_len[6][0] ),
    .S(_1433_),
    .X(_1434_));
 sg13g2_and2_1 _4614_ (.A(net32),
    .B(_1434_),
    .X(_0190_));
 sg13g2_mux2_1 _4615_ (.A0(_1160_),
    .A1(_2646_),
    .S(_1433_),
    .X(_1435_));
 sg13g2_and2_1 _4616_ (.A(_1255_),
    .B(_1435_),
    .X(_0191_));
 sg13g2_mux2_1 _4617_ (.A0(_1131_),
    .A1(_2764_),
    .S(_1433_),
    .X(_1436_));
 sg13g2_and2_1 _4618_ (.A(_1255_),
    .B(_1436_),
    .X(_0192_));
 sg13g2_buf_1 _4619_ (.A(net46),
    .X(_1437_));
 sg13g2_nand3_1 _4620_ (.B(_1229_),
    .C(net37),
    .A(_0456_),
    .Y(_1438_));
 sg13g2_nor2_1 _4621_ (.A(_1020_),
    .B(_1026_),
    .Y(_1439_));
 sg13g2_nand2_1 _4622_ (.Y(_1440_),
    .A(net28),
    .B(_1439_));
 sg13g2_inv_1 _4623_ (.Y(_1441_),
    .A(_1221_));
 sg13g2_a22oi_1 _4624_ (.Y(_1442_),
    .B1(_1103_),
    .B2(_1441_),
    .A2(_1030_),
    .A1(net28));
 sg13g2_buf_2 _4625_ (.A(_1442_),
    .X(_1443_));
 sg13g2_a21oi_1 _4626_ (.A1(_1438_),
    .A2(_1440_),
    .Y(_1444_),
    .B1(_1443_));
 sg13g2_xnor2_1 _4627_ (.Y(_1445_),
    .A(_0700_),
    .B(_1444_));
 sg13g2_nor2_1 _4628_ (.A(net31),
    .B(_1445_),
    .Y(_0208_));
 sg13g2_nand3_1 _4629_ (.B(net28),
    .C(_1439_),
    .A(_0700_),
    .Y(_1446_));
 sg13g2_o21ai_1 _4630_ (.B1(_1446_),
    .Y(_1447_),
    .A1(_0700_),
    .A2(_1438_));
 sg13g2_nor2b_1 _4631_ (.A(_1443_),
    .B_N(_1447_),
    .Y(_1448_));
 sg13g2_xnor2_1 _4632_ (.Y(_1449_),
    .A(\game.fsm.green_block_count[1] ),
    .B(_1448_));
 sg13g2_nor2_1 _4633_ (.A(_1437_),
    .B(_1449_),
    .Y(_0209_));
 sg13g2_or3_1 _4634_ (.A(_0700_),
    .B(\game.fsm.green_block_count[1] ),
    .C(_1438_),
    .X(_1450_));
 sg13g2_nand4_1 _4635_ (.B(\game.fsm.green_block_count[1] ),
    .C(net28),
    .A(_0700_),
    .Y(_1451_),
    .D(_1439_));
 sg13g2_a21oi_1 _4636_ (.A1(_1450_),
    .A2(_1451_),
    .Y(_1452_),
    .B1(_1443_));
 sg13g2_xnor2_1 _4637_ (.Y(_1453_),
    .A(\game.fsm.green_block_count[2] ),
    .B(_1452_));
 sg13g2_nor2_1 _4638_ (.A(_1437_),
    .B(_1453_),
    .Y(_0210_));
 sg13g2_xnor2_1 _4639_ (.Y(_1454_),
    .A(_0718_),
    .B(_1225_));
 sg13g2_nor2_1 _4640_ (.A(net31),
    .B(_1454_),
    .Y(_0211_));
 sg13g2_o21ai_1 _4641_ (.B1(_1068_),
    .Y(_1455_),
    .A1(net28),
    .A2(_1221_));
 sg13g2_xnor2_1 _4642_ (.Y(_1456_),
    .A(_0691_),
    .B(_1455_));
 sg13g2_nor2_1 _4643_ (.A(_1225_),
    .B(_1456_),
    .Y(_1457_));
 sg13g2_xnor2_1 _4644_ (.Y(_1458_),
    .A(\game.fsm.len1_block_count[1] ),
    .B(_1457_));
 sg13g2_nor2_1 _4645_ (.A(net31),
    .B(_1458_),
    .Y(_0212_));
 sg13g2_nor2_1 _4646_ (.A(_0718_),
    .B(_1455_),
    .Y(_1459_));
 sg13g2_nor2_1 _4647_ (.A(\game.fsm.len1_block_count[1] ),
    .B(_0691_),
    .Y(_1460_));
 sg13g2_a22oi_1 _4648_ (.Y(_1461_),
    .B1(_1460_),
    .B2(_1455_),
    .A2(_1459_),
    .A1(\game.fsm.len1_block_count[1] ));
 sg13g2_nor2_1 _4649_ (.A(_1225_),
    .B(_1461_),
    .Y(_1462_));
 sg13g2_xnor2_1 _4650_ (.Y(_1463_),
    .A(\game.fsm.len1_block_count[2] ),
    .B(_1462_));
 sg13g2_nor2_1 _4651_ (.A(net31),
    .B(_1463_),
    .Y(_0213_));
 sg13g2_a22oi_1 _4652_ (.Y(_1464_),
    .B1(net26),
    .B2(_1103_),
    .A2(_1223_),
    .A1(_1124_));
 sg13g2_xor2_1 _4653_ (.B(_1464_),
    .A(_0681_),
    .X(_1465_));
 sg13g2_nor2_1 _4654_ (.A(net31),
    .B(_1465_),
    .Y(_0226_));
 sg13g2_o21ai_1 _4655_ (.B1(_1221_),
    .Y(_1466_),
    .A1(net28),
    .A2(_1247_));
 sg13g2_xor2_1 _4656_ (.B(_1466_),
    .A(_0681_),
    .X(_1467_));
 sg13g2_nor2_1 _4657_ (.A(_1464_),
    .B(_1467_),
    .Y(_1468_));
 sg13g2_xnor2_1 _4658_ (.Y(_1469_),
    .A(\game.fsm.len2_block_count[1] ),
    .B(_1468_));
 sg13g2_nor2_1 _4659_ (.A(net31),
    .B(_1469_),
    .Y(_0227_));
 sg13g2_a21oi_1 _4660_ (.A1(_1097_),
    .A2(net26),
    .Y(_1470_),
    .B1(_1321_));
 sg13g2_o21ai_1 _4661_ (.B1(_1350_),
    .Y(_1471_),
    .A1(_1066_),
    .A2(_1470_));
 sg13g2_xnor2_1 _4662_ (.Y(_1472_),
    .A(_0723_),
    .B(_1471_));
 sg13g2_nor2_1 _4663_ (.A(net31),
    .B(_1472_),
    .Y(_0236_));
 sg13g2_o21ai_1 _4664_ (.B1(_1258_),
    .Y(_1473_),
    .A1(net28),
    .A2(_1245_));
 sg13g2_xnor2_1 _4665_ (.Y(_1474_),
    .A(_0723_),
    .B(_1473_));
 sg13g2_nand2_1 _4666_ (.Y(_1475_),
    .A(_1471_),
    .B(_1474_));
 sg13g2_xnor2_1 _4667_ (.Y(_1476_),
    .A(_0724_),
    .B(_1475_));
 sg13g2_nor2_1 _4668_ (.A(net31),
    .B(_1476_),
    .Y(_0237_));
 sg13g2_o21ai_1 _4669_ (.B1(_1061_),
    .Y(_1477_),
    .A1(_0066_),
    .A2(_1101_));
 sg13g2_nor2_1 _4670_ (.A(net69),
    .B(net48),
    .Y(_1478_));
 sg13g2_nand2_1 _4671_ (.Y(_1479_),
    .A(_0066_),
    .B(_1047_));
 sg13g2_a221oi_1 _4672_ (.B2(_1479_),
    .C1(_1132_),
    .B1(_1478_),
    .A1(net69),
    .Y(_0246_),
    .A2(_1477_));
 sg13g2_xnor2_1 _4673_ (.Y(_1480_),
    .A(net50),
    .B(_1375_));
 sg13g2_nand3_1 _4674_ (.B(net101),
    .C(net48),
    .A(net50),
    .Y(_1481_));
 sg13g2_o21ai_1 _4675_ (.B1(_1481_),
    .Y(_1482_),
    .A1(_0402_),
    .A2(net48));
 sg13g2_nor2_1 _4676_ (.A(net70),
    .B(_1482_),
    .Y(_1483_));
 sg13g2_a21oi_1 _4677_ (.A1(net70),
    .A2(_1480_),
    .Y(_1484_),
    .B1(_1483_));
 sg13g2_nor2_1 _4678_ (.A(_1132_),
    .B(_1484_),
    .Y(_0247_));
 sg13g2_nand3_1 _4679_ (.B(net102),
    .C(net48),
    .A(net69),
    .Y(_1485_));
 sg13g2_nand2_1 _4680_ (.Y(_1486_),
    .A(_1375_),
    .B(_1485_));
 sg13g2_nand2_1 _4681_ (.Y(_1487_),
    .A(net102),
    .B(_1101_));
 sg13g2_nor2_1 _4682_ (.A(net70),
    .B(net48),
    .Y(_1488_));
 sg13g2_a22oi_1 _4683_ (.Y(_1489_),
    .B1(_1487_),
    .B2(_1488_),
    .A2(_1486_),
    .A1(net50));
 sg13g2_inv_1 _4684_ (.Y(_1490_),
    .A(_1489_));
 sg13g2_o21ai_1 _4685_ (.B1(_1376_),
    .Y(_1491_),
    .A1(net101),
    .A2(_1047_));
 sg13g2_nor3_1 _4686_ (.A(net69),
    .B(net101),
    .C(_1040_),
    .Y(_1492_));
 sg13g2_a22oi_1 _4687_ (.Y(_1493_),
    .B1(_1047_),
    .B2(_1492_),
    .A2(_1040_),
    .A1(net72));
 sg13g2_o21ai_1 _4688_ (.B1(net38),
    .Y(_1494_),
    .A1(net50),
    .A2(_1493_));
 sg13g2_a221oi_1 _4689_ (.B2(net72),
    .C1(_1494_),
    .B1(_1491_),
    .A1(net101),
    .Y(_0248_),
    .A2(_1490_));
 sg13g2_nor3_1 _4690_ (.A(_1079_),
    .B(net37),
    .C(_1443_),
    .Y(_1495_));
 sg13g2_a21oi_1 _4691_ (.A1(net64),
    .A2(_1443_),
    .Y(_1496_),
    .B1(_1495_));
 sg13g2_nand4_1 _4692_ (.B(net37),
    .C(_1103_),
    .A(_0033_),
    .Y(_1497_),
    .D(_1441_));
 sg13g2_a21oi_1 _4693_ (.A1(_1496_),
    .A2(_1497_),
    .Y(_0249_),
    .B1(net35));
 sg13g2_xnor2_1 _4694_ (.Y(_1498_),
    .A(net64),
    .B(net37));
 sg13g2_nor2_1 _4695_ (.A(_1443_),
    .B(_1498_),
    .Y(_1499_));
 sg13g2_xnor2_1 _4696_ (.Y(_1500_),
    .A(net68),
    .B(_1499_));
 sg13g2_nor2_1 _4697_ (.A(net35),
    .B(_1500_),
    .Y(_0250_));
 sg13g2_nand2_1 _4698_ (.Y(_1501_),
    .A(net37),
    .B(_1065_));
 sg13g2_o21ai_1 _4699_ (.B1(_1501_),
    .Y(_1502_),
    .A1(_2868_),
    .A2(net37));
 sg13g2_xnor2_1 _4700_ (.Y(_1503_),
    .A(_1073_),
    .B(_1502_));
 sg13g2_nor2_1 _4701_ (.A(_1443_),
    .B(_1503_),
    .Y(_1504_));
 sg13g2_a21oi_1 _4702_ (.A1(net130),
    .A2(_1443_),
    .Y(_1505_),
    .B1(_1504_));
 sg13g2_nor2_1 _4703_ (.A(net35),
    .B(_1505_),
    .Y(_0251_));
 sg13g2_inv_1 _4704_ (.Y(_1506_),
    .A(_0424_));
 sg13g2_nand3_1 _4705_ (.B(_1399_),
    .C(_1367_),
    .A(_1361_),
    .Y(_1507_));
 sg13g2_nand2_1 _4706_ (.Y(_1508_),
    .A(net38),
    .B(_1507_));
 sg13g2_a22oi_1 _4707_ (.Y(_0264_),
    .B1(_1508_),
    .B2(_1358_),
    .A2(_1507_),
    .A1(_1506_));
 sg13g2_inv_1 _4708_ (.Y(_1509_),
    .A(_0406_));
 sg13g2_a22oi_1 _4709_ (.Y(_0265_),
    .B1(_1508_),
    .B2(_1373_),
    .A2(_1507_),
    .A1(_1509_));
 sg13g2_buf_8 _4710_ (.A(_2638_),
    .X(_1510_));
 sg13g2_nand2_1 _4711_ (.Y(_1511_),
    .A(net121),
    .B(_0857_));
 sg13g2_nor3_1 _4712_ (.A(net91),
    .B(_2645_),
    .C(_1511_),
    .Y(_0282_));
 sg13g2_and2_1 _4713_ (.A(_2635_),
    .B(_0282_),
    .X(_0279_));
 sg13g2_and2_1 _4714_ (.A(_2634_),
    .B(_0282_),
    .X(_0280_));
 sg13g2_nand2b_1 _4715_ (.Y(_1512_),
    .B(\game.slv.state[3] ),
    .A_N(\game.slv.saved_target ));
 sg13g2_nor4_1 _4716_ (.A(_0710_),
    .B(_0726_),
    .C(_0730_),
    .D(_1512_),
    .Y(_1513_));
 sg13g2_and2_1 _4717_ (.A(\game.slv.saved_target ),
    .B(\game.slv.state[3] ),
    .X(_1514_));
 sg13g2_nor2b_1 _4718_ (.A(_0850_),
    .B_N(_1514_),
    .Y(_1515_));
 sg13g2_or2_1 _4719_ (.X(_1516_),
    .B(_0730_),
    .A(_0726_));
 sg13g2_a21oi_1 _4720_ (.A1(_0840_),
    .A2(_0849_),
    .Y(_1517_),
    .B1(_1512_));
 sg13g2_mux2_1 _4721_ (.A0(_1517_),
    .A1(_1514_),
    .S(_0710_),
    .X(_1518_));
 sg13g2_a221oi_1 _4722_ (.B2(_1516_),
    .C1(_1518_),
    .B1(_1515_),
    .A1(_2836_),
    .Y(_1519_),
    .A2(_1513_));
 sg13g2_nand2b_1 _4723_ (.Y(_1520_),
    .B(_1515_),
    .A_N(_2836_));
 sg13g2_nand2_1 _4724_ (.Y(_1521_),
    .A(_1013_),
    .B(_0859_));
 sg13g2_a21o_1 _4725_ (.A2(_1520_),
    .A1(_1519_),
    .B1(_1521_),
    .X(_1522_));
 sg13g2_buf_2 _4726_ (.A(_1522_),
    .X(_1523_));
 sg13g2_nor2_1 _4727_ (.A(_2645_),
    .B(_1523_),
    .Y(_0310_));
 sg13g2_buf_1 _4728_ (.A(net118),
    .X(_1524_));
 sg13g2_buf_1 _4729_ (.A(net119),
    .X(_1525_));
 sg13g2_nand2_2 _4730_ (.Y(_1526_),
    .A(net120),
    .B(_0871_));
 sg13g2_nor3_2 _4731_ (.A(net90),
    .B(net89),
    .C(_1526_),
    .Y(_1527_));
 sg13g2_and3_1 _4732_ (.X(_0318_),
    .A(net95),
    .B(\game.solver_trigger_delayed ),
    .C(_1527_));
 sg13g2_buf_1 _4733_ (.A(\snd.note_timing[8] ),
    .X(_1528_));
 sg13g2_inv_1 _4734_ (.Y(_1529_),
    .A(_1528_));
 sg13g2_buf_1 _4735_ (.A(\snd.counter[8] ),
    .X(_1530_));
 sg13g2_inv_1 _4736_ (.Y(_1531_),
    .A(_1530_));
 sg13g2_buf_1 _4737_ (.A(\snd.counter[7] ),
    .X(_1532_));
 sg13g2_buf_1 _4738_ (.A(\snd.note_timing[6] ),
    .X(_1533_));
 sg13g2_inv_1 _4739_ (.Y(_1534_),
    .A(\snd.counter[6] ));
 sg13g2_nor2b_1 _4740_ (.A(\snd.counter[6] ),
    .B_N(_1533_),
    .Y(_1535_));
 sg13g2_buf_2 _4741_ (.A(\snd.counter[5] ),
    .X(_1536_));
 sg13g2_buf_1 _4742_ (.A(\snd.note_timing[4] ),
    .X(_1537_));
 sg13g2_buf_2 _4743_ (.A(\snd.counter[4] ),
    .X(_1538_));
 sg13g2_inv_1 _4744_ (.Y(_1539_),
    .A(_1538_));
 sg13g2_nor2_1 _4745_ (.A(_1537_),
    .B(_1539_),
    .Y(_1540_));
 sg13g2_buf_1 _4746_ (.A(\snd.counter[3] ),
    .X(_1541_));
 sg13g2_buf_1 _4747_ (.A(\snd.counter[2] ),
    .X(_1542_));
 sg13g2_inv_1 _4748_ (.Y(_1543_),
    .A(_1542_));
 sg13g2_inv_1 _4749_ (.Y(_1544_),
    .A(\snd.note_timing[2] ));
 sg13g2_buf_2 _4750_ (.A(\snd.counter[0] ),
    .X(_1545_));
 sg13g2_nand2b_1 _4751_ (.Y(_1546_),
    .B(\snd.note_timing[0] ),
    .A_N(_1545_));
 sg13g2_buf_2 _4752_ (.A(\snd.counter[1] ),
    .X(_1547_));
 sg13g2_buf_1 _4753_ (.A(\snd.note_timing[1] ),
    .X(_1548_));
 sg13g2_nor2_1 _4754_ (.A(_1547_),
    .B(_1546_),
    .Y(_1549_));
 sg13g2_nor2_1 _4755_ (.A(_1548_),
    .B(_1549_),
    .Y(_1550_));
 sg13g2_a221oi_1 _4756_ (.B2(_1547_),
    .C1(_1550_),
    .B1(_1546_),
    .A1(_1544_),
    .Y(_1551_),
    .A2(_1542_));
 sg13g2_a21oi_1 _4757_ (.A1(\snd.note_timing[2] ),
    .A2(_1543_),
    .Y(_1552_),
    .B1(_1551_));
 sg13g2_nand2_1 _4758_ (.Y(_1553_),
    .A(_1541_),
    .B(_1552_));
 sg13g2_inv_1 _4759_ (.Y(_1554_),
    .A(\snd.note_timing[3] ));
 sg13g2_o21ai_1 _4760_ (.B1(_1554_),
    .Y(_1555_),
    .A1(_1541_),
    .A2(_1552_));
 sg13g2_a22oi_1 _4761_ (.Y(_1556_),
    .B1(_1553_),
    .B2(_1555_),
    .A2(_1539_),
    .A1(_1537_));
 sg13g2_or2_1 _4762_ (.X(_1557_),
    .B(_1556_),
    .A(_1540_));
 sg13g2_nor2_1 _4763_ (.A(_1536_),
    .B(_1557_),
    .Y(_1558_));
 sg13g2_inv_1 _4764_ (.Y(_1559_),
    .A(\snd.note_timing[5] ));
 sg13g2_a21oi_1 _4765_ (.A1(_1536_),
    .A2(_1557_),
    .Y(_1560_),
    .B1(_1559_));
 sg13g2_or3_1 _4766_ (.A(_1535_),
    .B(_1558_),
    .C(_1560_),
    .X(_1561_));
 sg13g2_o21ai_1 _4767_ (.B1(_1561_),
    .Y(_1562_),
    .A1(_1533_),
    .A2(_1534_));
 sg13g2_inv_1 _4768_ (.Y(_1563_),
    .A(\snd.note_timing[7] ));
 sg13g2_o21ai_1 _4769_ (.B1(_1563_),
    .Y(_1564_),
    .A1(_1532_),
    .A2(_1562_));
 sg13g2_nand2_1 _4770_ (.Y(_1565_),
    .A(_1532_),
    .B(_1562_));
 sg13g2_a22oi_1 _4771_ (.Y(_1566_),
    .B1(_1564_),
    .B2(_1565_),
    .A2(_1531_),
    .A1(_1528_));
 sg13g2_a21oi_1 _4772_ (.A1(_1529_),
    .A2(_1530_),
    .Y(_1567_),
    .B1(_1566_));
 sg13g2_buf_2 _4773_ (.A(_1567_),
    .X(_1568_));
 sg13g2_nand2_1 _4774_ (.Y(_1569_),
    .A(net134),
    .B(_1568_));
 sg13g2_buf_1 _4775_ (.A(_1569_),
    .X(_1570_));
 sg13g2_xnor2_1 _4776_ (.Y(_1571_),
    .A(_1545_),
    .B(_1547_));
 sg13g2_nor2_1 _4777_ (.A(net19),
    .B(_1571_),
    .Y(_0344_));
 sg13g2_nand2_1 _4778_ (.Y(_1572_),
    .A(_1545_),
    .B(_1547_));
 sg13g2_xnor2_1 _4779_ (.Y(_1573_),
    .A(_1543_),
    .B(_1572_));
 sg13g2_nor2_1 _4780_ (.A(net19),
    .B(_1573_),
    .Y(_0345_));
 sg13g2_inv_1 _4781_ (.Y(_1574_),
    .A(_1541_));
 sg13g2_nand3_1 _4782_ (.B(_1547_),
    .C(_1542_),
    .A(_1545_),
    .Y(_1575_));
 sg13g2_xnor2_1 _4783_ (.Y(_1576_),
    .A(_1574_),
    .B(_1575_));
 sg13g2_nor2_1 _4784_ (.A(net19),
    .B(_1576_),
    .Y(_0346_));
 sg13g2_nor2_1 _4785_ (.A(_1574_),
    .B(_1575_),
    .Y(_1577_));
 sg13g2_xnor2_1 _4786_ (.Y(_1578_),
    .A(_1538_),
    .B(_1577_));
 sg13g2_nor2_1 _4787_ (.A(net19),
    .B(_1578_),
    .Y(_0347_));
 sg13g2_nand2_1 _4788_ (.Y(_1579_),
    .A(_1538_),
    .B(_1577_));
 sg13g2_xor2_1 _4789_ (.B(_1579_),
    .A(_1536_),
    .X(_1580_));
 sg13g2_nor2_1 _4790_ (.A(_1570_),
    .B(_1580_),
    .Y(_0348_));
 sg13g2_nand3_1 _4791_ (.B(_1536_),
    .C(_1577_),
    .A(_1538_),
    .Y(_1581_));
 sg13g2_xnor2_1 _4792_ (.Y(_1582_),
    .A(_1534_),
    .B(_1581_));
 sg13g2_nor2_1 _4793_ (.A(net19),
    .B(_1582_),
    .Y(_0349_));
 sg13g2_inv_1 _4794_ (.Y(_1583_),
    .A(_1532_));
 sg13g2_or2_1 _4795_ (.X(_1584_),
    .B(_1581_),
    .A(_1534_));
 sg13g2_xnor2_1 _4796_ (.Y(_1585_),
    .A(_1583_),
    .B(_1584_));
 sg13g2_nor2_1 _4797_ (.A(net19),
    .B(_1585_),
    .Y(_0350_));
 sg13g2_nor2_1 _4798_ (.A(_1583_),
    .B(_1584_),
    .Y(_1586_));
 sg13g2_xnor2_1 _4799_ (.Y(_1587_),
    .A(_1530_),
    .B(_1586_));
 sg13g2_nor2_1 _4800_ (.A(net19),
    .B(_1587_),
    .Y(_0351_));
 sg13g2_nand2_1 _4801_ (.Y(_1588_),
    .A(\snd.note_timing[7] ),
    .B(_1534_));
 sg13g2_inv_1 _4802_ (.Y(_1589_),
    .A(_1545_));
 sg13g2_nor2_1 _4803_ (.A(_1544_),
    .B(_1547_),
    .Y(_1590_));
 sg13g2_nor3_1 _4804_ (.A(_1548_),
    .B(_1589_),
    .C(_1590_),
    .Y(_1591_));
 sg13g2_a221oi_1 _4805_ (.B2(_1542_),
    .C1(_1591_),
    .B1(_1554_),
    .A1(_1544_),
    .Y(_1592_),
    .A2(_1547_));
 sg13g2_a21oi_1 _4806_ (.A1(\snd.note_timing[3] ),
    .A2(_1543_),
    .Y(_1593_),
    .B1(_1592_));
 sg13g2_nor2_1 _4807_ (.A(_1541_),
    .B(_1593_),
    .Y(_1594_));
 sg13g2_nor2_1 _4808_ (.A(_1537_),
    .B(_1594_),
    .Y(_1595_));
 sg13g2_a221oi_1 _4809_ (.B2(_1541_),
    .C1(_1595_),
    .B1(_1593_),
    .A1(_1559_),
    .Y(_1596_),
    .A2(_1538_));
 sg13g2_a21oi_1 _4810_ (.A1(\snd.note_timing[5] ),
    .A2(_1539_),
    .Y(_1597_),
    .B1(_1596_));
 sg13g2_nor2_1 _4811_ (.A(_1536_),
    .B(_1597_),
    .Y(_1598_));
 sg13g2_nand2_1 _4812_ (.Y(_1599_),
    .A(_1536_),
    .B(_1597_));
 sg13g2_o21ai_1 _4813_ (.B1(_1599_),
    .Y(_1600_),
    .A1(_1533_),
    .A2(_1598_));
 sg13g2_xor2_1 _4814_ (.B(_1532_),
    .A(_1528_),
    .X(_1601_));
 sg13g2_a21oi_1 _4815_ (.A1(_1563_),
    .A2(\snd.counter[6] ),
    .Y(_1602_),
    .B1(_1601_));
 sg13g2_nand2_1 _4816_ (.Y(_1603_),
    .A(_0036_),
    .B(_1602_));
 sg13g2_a21oi_1 _4817_ (.A1(_1588_),
    .A2(_1600_),
    .Y(_1604_),
    .B1(_1603_));
 sg13g2_nor3_1 _4818_ (.A(_1529_),
    .B(_1532_),
    .C(_1530_),
    .Y(_1605_));
 sg13g2_nor2_1 _4819_ (.A(_1604_),
    .B(_1605_),
    .Y(_1606_));
 sg13g2_xnor2_1 _4820_ (.Y(_1607_),
    .A(\snd.note_timing[3] ),
    .B(_1542_));
 sg13g2_xnor2_1 _4821_ (.Y(_1608_),
    .A(_1537_),
    .B(_1541_));
 sg13g2_xnor2_1 _4822_ (.Y(_1609_),
    .A(_1548_),
    .B(_1545_));
 sg13g2_nand4_1 _4823_ (.B(_1607_),
    .C(_1608_),
    .A(_1588_),
    .Y(_1610_),
    .D(_1609_));
 sg13g2_xnor2_1 _4824_ (.Y(_1611_),
    .A(\snd.note_timing[5] ),
    .B(_1538_));
 sg13g2_xnor2_1 _4825_ (.Y(_1612_),
    .A(_1533_),
    .B(_1536_));
 sg13g2_xnor2_1 _4826_ (.Y(_1613_),
    .A(\snd.note_timing[2] ),
    .B(_1547_));
 sg13g2_nand3_1 _4827_ (.B(_1612_),
    .C(_1613_),
    .A(_1611_),
    .Y(_1614_));
 sg13g2_nor3_1 _4828_ (.A(_1603_),
    .B(_1610_),
    .C(_1614_),
    .Y(_1615_));
 sg13g2_nor3_1 _4829_ (.A(\snd.sound ),
    .B(_1606_),
    .C(_1615_),
    .Y(_1616_));
 sg13g2_nor2_1 _4830_ (.A(net19),
    .B(_1616_),
    .Y(_0376_));
 sg13g2_inv_1 _4831_ (.Y(_1617_),
    .A(_0871_));
 sg13g2_nor2_1 _4832_ (.A(net120),
    .B(_1617_),
    .Y(_1618_));
 sg13g2_and2_1 _4833_ (.A(_0881_),
    .B(_1618_),
    .X(_1619_));
 sg13g2_buf_1 _4834_ (.A(_1619_),
    .X(_1620_));
 sg13g2_nor2_1 _4835_ (.A(\game.fsm.read_pos[0] ),
    .B(net44),
    .Y(_1621_));
 sg13g2_buf_1 _4836_ (.A(\game.counter[6] ),
    .X(_1622_));
 sg13g2_buf_1 _4837_ (.A(\game.counter[5] ),
    .X(_1623_));
 sg13g2_and2_1 _4838_ (.A(_1622_),
    .B(_1623_),
    .X(_1624_));
 sg13g2_buf_1 _4839_ (.A(\game.counter[4] ),
    .X(_1625_));
 sg13g2_buf_2 _4840_ (.A(\game.counter[2] ),
    .X(_1626_));
 sg13g2_buf_1 _4841_ (.A(\game.counter[3] ),
    .X(_1627_));
 sg13g2_or3_1 _4842_ (.A(_1625_),
    .B(_1626_),
    .C(_1627_),
    .X(_1628_));
 sg13g2_buf_1 _4843_ (.A(\game.counter[7] ),
    .X(_1629_));
 sg13g2_a21oi_1 _4844_ (.A1(_1624_),
    .A2(_1628_),
    .Y(_1630_),
    .B1(_1629_));
 sg13g2_nand2_2 _4845_ (.Y(_1631_),
    .A(_0862_),
    .B(_1617_));
 sg13g2_nor3_2 _4846_ (.A(net118),
    .B(net119),
    .C(_1631_),
    .Y(_1632_));
 sg13g2_buf_1 _4847_ (.A(\game.fsm.read_pos[2] ),
    .X(_1633_));
 sg13g2_inv_1 _4848_ (.Y(_1634_),
    .A(_1633_));
 sg13g2_buf_1 _4849_ (.A(\game.fsm.read_pos[1] ),
    .X(_1635_));
 sg13g2_inv_1 _4850_ (.Y(_1636_),
    .A(\game.fsm.read_pos[0] ));
 sg13g2_inv_1 _4851_ (.Y(_1637_),
    .A(_1635_));
 sg13g2_a22oi_1 _4852_ (.Y(_1638_),
    .B1(_1637_),
    .B2(net50),
    .A2(_1636_),
    .A1(net69));
 sg13g2_a221oi_1 _4853_ (.B2(net72),
    .C1(_1638_),
    .B1(_1633_),
    .A1(_0429_),
    .Y(_1639_),
    .A2(_1635_));
 sg13g2_a21oi_2 _4854_ (.B1(_1639_),
    .Y(_1640_),
    .A2(_1634_),
    .A1(net102));
 sg13g2_a21o_1 _4855_ (.A2(_1640_),
    .A1(_1632_),
    .B1(_1630_),
    .X(_1641_));
 sg13g2_buf_1 _4856_ (.A(\btn.gate_200hz ),
    .X(_1642_));
 sg13g2_buf_1 _4857_ (.A(_0035_),
    .X(_1643_));
 sg13g2_inv_1 _4858_ (.Y(_1644_),
    .A(_1643_));
 sg13g2_o21ai_1 _4859_ (.B1(_1644_),
    .Y(_1645_),
    .A1(net44),
    .A2(_1632_));
 sg13g2_a221oi_1 _4860_ (.B2(_1642_),
    .C1(_1645_),
    .B1(_1641_),
    .A1(net44),
    .Y(_1646_),
    .A2(_1630_));
 sg13g2_buf_1 _4861_ (.A(_1646_),
    .X(_1647_));
 sg13g2_nand2_1 _4862_ (.Y(_1648_),
    .A(_1621_),
    .B(_1647_));
 sg13g2_inv_1 _4863_ (.Y(_1649_),
    .A(_1647_));
 sg13g2_nand2_1 _4864_ (.Y(_1650_),
    .A(\game.fsm.read_pos[0] ),
    .B(_1649_));
 sg13g2_a21oi_1 _4865_ (.A1(_1648_),
    .A2(_1650_),
    .Y(_0095_),
    .B1(_2643_));
 sg13g2_nand2b_1 _4866_ (.Y(_1651_),
    .B(_1647_),
    .A_N(_1621_));
 sg13g2_nor3_1 _4867_ (.A(_1636_),
    .B(_1635_),
    .C(net44),
    .Y(_1652_));
 sg13g2_a22oi_1 _4868_ (.Y(_1653_),
    .B1(_1652_),
    .B2(_1647_),
    .A2(_1651_),
    .A1(_1635_));
 sg13g2_nor2_1 _4869_ (.A(net63),
    .B(_1653_),
    .Y(_0096_));
 sg13g2_nand2_1 _4870_ (.Y(_1654_),
    .A(\game.fsm.read_pos[0] ),
    .B(_1635_));
 sg13g2_nor3_1 _4871_ (.A(_1633_),
    .B(_1649_),
    .C(_1654_),
    .Y(_1655_));
 sg13g2_a21oi_1 _4872_ (.A1(_1633_),
    .A2(_1654_),
    .Y(_1656_),
    .B1(_1655_));
 sg13g2_nand2_1 _4873_ (.Y(_1657_),
    .A(_1633_),
    .B(_1649_));
 sg13g2_o21ai_1 _4874_ (.B1(_1657_),
    .Y(_1658_),
    .A1(net44),
    .A2(_1656_));
 sg13g2_and2_1 _4875_ (.A(net66),
    .B(_1658_),
    .X(_0097_));
 sg13g2_buf_2 _4876_ (.A(\btn.button_state[0] ),
    .X(_1659_));
 sg13g2_inv_1 _4877_ (.Y(_1660_),
    .A(_1642_));
 sg13g2_nand3_1 _4878_ (.B(\btn.sample_10ms[0] ),
    .C(\btn.sample_15ms[0] ),
    .A(\btn.sample_5ms[0] ),
    .Y(_1661_));
 sg13g2_or2_1 _4879_ (.X(_1662_),
    .B(_1661_),
    .A(net88));
 sg13g2_mux2_1 _4880_ (.A0(net1),
    .A1(_1659_),
    .S(_1662_),
    .X(_1663_));
 sg13g2_and2_1 _4881_ (.A(net66),
    .B(_1663_),
    .X(_0098_));
 sg13g2_buf_2 _4882_ (.A(\btn.button_state[1] ),
    .X(_1664_));
 sg13g2_buf_1 _4883_ (.A(_1642_),
    .X(_1665_));
 sg13g2_buf_1 _4884_ (.A(_1665_),
    .X(_1666_));
 sg13g2_nor2_1 _4885_ (.A(_1664_),
    .B(net62),
    .Y(_1667_));
 sg13g2_buf_1 _4886_ (.A(_1660_),
    .X(_1668_));
 sg13g2_nand3_1 _4887_ (.B(\btn.sample_10ms[1] ),
    .C(\btn.sample_15ms[1] ),
    .A(\btn.sample_5ms[1] ),
    .Y(_1669_));
 sg13g2_mux2_1 _4888_ (.A0(net2),
    .A1(_1664_),
    .S(_1669_),
    .X(_1670_));
 sg13g2_nor2_1 _4889_ (.A(net61),
    .B(_1670_),
    .Y(_1671_));
 sg13g2_nor3_1 _4890_ (.A(net65),
    .B(_1667_),
    .C(_1671_),
    .Y(_0099_));
 sg13g2_buf_1 _4891_ (.A(_2642_),
    .X(_1672_));
 sg13g2_buf_2 _4892_ (.A(\btn.button_state[2] ),
    .X(_1673_));
 sg13g2_nor2_1 _4893_ (.A(_1673_),
    .B(net62),
    .Y(_1674_));
 sg13g2_nand3_1 _4894_ (.B(\btn.sample_10ms[2] ),
    .C(\btn.sample_15ms[2] ),
    .A(\btn.sample_5ms[2] ),
    .Y(_1675_));
 sg13g2_mux2_1 _4895_ (.A0(net3),
    .A1(_1673_),
    .S(_1675_),
    .X(_1676_));
 sg13g2_nor2_1 _4896_ (.A(net61),
    .B(_1676_),
    .Y(_1677_));
 sg13g2_nor3_1 _4897_ (.A(net60),
    .B(_1674_),
    .C(_1677_),
    .Y(_0100_));
 sg13g2_buf_2 _4898_ (.A(\btn.button_state[3] ),
    .X(_1678_));
 sg13g2_nor2_1 _4899_ (.A(_1678_),
    .B(net62),
    .Y(_1679_));
 sg13g2_nand3_1 _4900_ (.B(\btn.sample_10ms[3] ),
    .C(\btn.sample_15ms[3] ),
    .A(\btn.sample_5ms[3] ),
    .Y(_1680_));
 sg13g2_mux2_1 _4901_ (.A0(net4),
    .A1(_1678_),
    .S(_1680_),
    .X(_1681_));
 sg13g2_nor2_1 _4902_ (.A(net61),
    .B(_1681_),
    .Y(_1682_));
 sg13g2_nor3_1 _4903_ (.A(net60),
    .B(_1679_),
    .C(_1682_),
    .Y(_0101_));
 sg13g2_buf_1 _4904_ (.A(\btn.change_timer[0] ),
    .X(_1683_));
 sg13g2_xor2_1 _4905_ (.B(_1664_),
    .A(net2),
    .X(_1684_));
 sg13g2_nand2b_1 _4906_ (.Y(_1685_),
    .B(_1684_),
    .A_N(_1669_));
 sg13g2_xor2_1 _4907_ (.B(_1673_),
    .A(net3),
    .X(_1686_));
 sg13g2_nand2b_1 _4908_ (.Y(_1687_),
    .B(_1686_),
    .A_N(_1675_));
 sg13g2_xor2_1 _4909_ (.B(_1659_),
    .A(net1),
    .X(_1688_));
 sg13g2_nand2b_1 _4910_ (.Y(_1689_),
    .B(_1688_),
    .A_N(_1661_));
 sg13g2_xor2_1 _4911_ (.B(_1678_),
    .A(net4),
    .X(_1690_));
 sg13g2_nand2b_1 _4912_ (.Y(_1691_),
    .B(_1690_),
    .A_N(_1680_));
 sg13g2_and4_1 _4913_ (.A(_1685_),
    .B(_1687_),
    .C(_1689_),
    .D(_1691_),
    .X(_1692_));
 sg13g2_buf_1 _4914_ (.A(_1692_),
    .X(_1693_));
 sg13g2_nor4_2 _4915_ (.A(_1659_),
    .B(_1664_),
    .C(_1673_),
    .Y(_1694_),
    .D(_1678_));
 sg13g2_nand2_1 _4916_ (.Y(_1695_),
    .A(net43),
    .B(_1694_));
 sg13g2_buf_1 _4917_ (.A(\btn.change_timer[3] ),
    .X(_1696_));
 sg13g2_buf_1 _4918_ (.A(\btn.change_timer[4] ),
    .X(_1697_));
 sg13g2_and2_1 _4919_ (.A(\btn.change_timer[1] ),
    .B(_1683_),
    .X(_1698_));
 sg13g2_and2_1 _4920_ (.A(\btn.change_timer[2] ),
    .B(_1698_),
    .X(_1699_));
 sg13g2_buf_1 _4921_ (.A(_1699_),
    .X(_1700_));
 sg13g2_and4_1 _4922_ (.A(_1696_),
    .B(\btn.change_timer[5] ),
    .C(_1697_),
    .D(_1700_),
    .X(_1701_));
 sg13g2_nand2_1 _4923_ (.Y(_1702_),
    .A(\btn.change_timer[6] ),
    .B(_1701_));
 sg13g2_nand3_1 _4924_ (.B(_1695_),
    .C(_1702_),
    .A(_1642_),
    .Y(_1703_));
 sg13g2_buf_1 _4925_ (.A(_1703_),
    .X(_1704_));
 sg13g2_inv_1 _4926_ (.Y(_1705_),
    .A(\btn.change_timer[2] ));
 sg13g2_or2_1 _4927_ (.X(_1706_),
    .B(_1683_),
    .A(\btn.change_timer[1] ));
 sg13g2_nor4_1 _4928_ (.A(_1705_),
    .B(\btn.change_timer[6] ),
    .C(_1694_),
    .D(_1706_),
    .Y(_1707_));
 sg13g2_nand4_1 _4929_ (.B(\btn.change_timer[5] ),
    .C(_1697_),
    .A(_1696_),
    .Y(_1708_),
    .D(_1707_));
 sg13g2_a21o_1 _4930_ (.A2(_1708_),
    .A1(net43),
    .B1(net88),
    .X(_1709_));
 sg13g2_buf_1 _4931_ (.A(_1709_),
    .X(_1710_));
 sg13g2_nand2_1 _4932_ (.Y(_1711_),
    .A(_1704_),
    .B(_1710_));
 sg13g2_buf_2 _4933_ (.A(_1711_),
    .X(_1712_));
 sg13g2_and3_1 _4934_ (.X(_1713_),
    .A(_1642_),
    .B(_1695_),
    .C(_1702_));
 sg13g2_buf_1 _4935_ (.A(_1713_),
    .X(_1714_));
 sg13g2_o21ai_1 _4936_ (.B1(net134),
    .Y(_1715_),
    .A1(net88),
    .A2(net43));
 sg13g2_buf_2 _4937_ (.A(_1715_),
    .X(_1716_));
 sg13g2_a21oi_1 _4938_ (.A1(_1683_),
    .A2(_1714_),
    .Y(_1717_),
    .B1(_1716_));
 sg13g2_o21ai_1 _4939_ (.B1(_1717_),
    .Y(_1718_),
    .A1(_1683_),
    .A2(_1712_));
 sg13g2_inv_1 _4940_ (.Y(_0102_),
    .A(_1718_));
 sg13g2_nand2_1 _4941_ (.Y(_1719_),
    .A(_1683_),
    .B(_1714_));
 sg13g2_o21ai_1 _4942_ (.B1(_1712_),
    .Y(_1720_),
    .A1(_1683_),
    .A2(_1704_));
 sg13g2_nor2_1 _4943_ (.A(\btn.change_timer[1] ),
    .B(_1720_),
    .Y(_1721_));
 sg13g2_a21oi_1 _4944_ (.A1(\btn.change_timer[1] ),
    .A2(_1719_),
    .Y(_1722_),
    .B1(_1721_));
 sg13g2_nor2_1 _4945_ (.A(_1716_),
    .B(_1722_),
    .Y(_0103_));
 sg13g2_o21ai_1 _4946_ (.B1(_1712_),
    .Y(_1723_),
    .A1(_1698_),
    .A2(_1704_));
 sg13g2_a221oi_1 _4947_ (.B2(_1705_),
    .C1(_1716_),
    .B1(_1723_),
    .A1(_1700_),
    .Y(_0104_),
    .A2(_1714_));
 sg13g2_nand2b_1 _4948_ (.Y(_1724_),
    .B(_1714_),
    .A_N(_1700_));
 sg13g2_a21oi_1 _4949_ (.A1(_1712_),
    .A2(_1724_),
    .Y(_1725_),
    .B1(_1696_));
 sg13g2_and3_1 _4950_ (.X(_1726_),
    .A(_1696_),
    .B(_1700_),
    .C(_1714_));
 sg13g2_nor3_1 _4951_ (.A(_1716_),
    .B(_1725_),
    .C(_1726_),
    .Y(_0105_));
 sg13g2_a21o_1 _4952_ (.A2(_1700_),
    .A1(_1696_),
    .B1(_1704_),
    .X(_1727_));
 sg13g2_a21oi_1 _4953_ (.A1(_1712_),
    .A2(_1727_),
    .Y(_1728_),
    .B1(_1697_));
 sg13g2_and4_1 _4954_ (.A(_1696_),
    .B(_1697_),
    .C(_1700_),
    .D(_1714_),
    .X(_1729_));
 sg13g2_nor3_1 _4955_ (.A(_1716_),
    .B(_1728_),
    .C(_1729_),
    .Y(_0106_));
 sg13g2_inv_1 _4956_ (.Y(_1730_),
    .A(\btn.change_timer[5] ));
 sg13g2_nand4_1 _4957_ (.B(_1697_),
    .C(_1700_),
    .A(_1696_),
    .Y(_1731_),
    .D(_1712_));
 sg13g2_nor3_1 _4958_ (.A(_1730_),
    .B(\btn.change_timer[6] ),
    .C(_1731_),
    .Y(_1732_));
 sg13g2_and2_1 _4959_ (.A(_1730_),
    .B(_1731_),
    .X(_1733_));
 sg13g2_nor3_1 _4960_ (.A(_1716_),
    .B(_1732_),
    .C(_1733_),
    .Y(_0107_));
 sg13g2_a21oi_1 _4961_ (.A1(_1701_),
    .A2(_1712_),
    .Y(_1734_),
    .B1(\btn.change_timer[6] ));
 sg13g2_nor2_1 _4962_ (.A(_1716_),
    .B(_1734_),
    .Y(_0108_));
 sg13g2_mux2_1 _4963_ (.A0(net1),
    .A1(_1659_),
    .S(_1661_),
    .X(_1735_));
 sg13g2_or2_1 _4964_ (.X(_1736_),
    .B(_1735_),
    .A(_1693_));
 sg13g2_or4_1 _4965_ (.A(_1670_),
    .B(_1676_),
    .C(_1681_),
    .D(_1736_),
    .X(_1737_));
 sg13g2_buf_1 _4966_ (.A(_1737_),
    .X(_1738_));
 sg13g2_o21ai_1 _4967_ (.B1(_2644_),
    .Y(_1739_),
    .A1(_1710_),
    .A2(_1738_));
 sg13g2_buf_1 _4968_ (.A(_1739_),
    .X(_1740_));
 sg13g2_nor2_1 _4969_ (.A(\btn.long_press ),
    .B(_1694_),
    .Y(_1741_));
 sg13g2_a21oi_2 _4970_ (.B1(_1710_),
    .Y(_1742_),
    .A2(_1741_),
    .A1(net43));
 sg13g2_a21oi_1 _4971_ (.A1(_1736_),
    .A2(_1742_),
    .Y(_1743_),
    .B1(\btn.current_event[0] ));
 sg13g2_nor2_1 _4972_ (.A(_1740_),
    .B(_1743_),
    .Y(_0109_));
 sg13g2_inv_1 _4973_ (.Y(_1744_),
    .A(\btn.current_event[1] ));
 sg13g2_o21ai_1 _4974_ (.B1(_1742_),
    .Y(_1745_),
    .A1(_1670_),
    .A2(net43));
 sg13g2_a21oi_1 _4975_ (.A1(_1744_),
    .A2(_1745_),
    .Y(_0110_),
    .B1(_1740_));
 sg13g2_inv_1 _4976_ (.Y(_1746_),
    .A(\btn.current_event[2] ));
 sg13g2_o21ai_1 _4977_ (.B1(_1742_),
    .Y(_1747_),
    .A1(_1676_),
    .A2(net43));
 sg13g2_a21oi_1 _4978_ (.A1(_1746_),
    .A2(_1747_),
    .Y(_0111_),
    .B1(_1740_));
 sg13g2_inv_1 _4979_ (.Y(_1748_),
    .A(\btn.current_event[3] ));
 sg13g2_o21ai_1 _4980_ (.B1(_1742_),
    .Y(_1749_),
    .A1(_1681_),
    .A2(net43));
 sg13g2_a21oi_1 _4981_ (.A1(_1748_),
    .A2(_1749_),
    .Y(_0112_),
    .B1(_1740_));
 sg13g2_nand2_1 _4982_ (.Y(_1750_),
    .A(_2644_),
    .B(net87));
 sg13g2_nor2_1 _4983_ (.A(_1738_),
    .B(_1750_),
    .Y(_1751_));
 sg13g2_and2_1 _4984_ (.A(\btn.current_event[0] ),
    .B(_1751_),
    .X(_0113_));
 sg13g2_nor3_1 _4985_ (.A(_1744_),
    .B(_1738_),
    .C(_1750_),
    .Y(_0114_));
 sg13g2_nor3_1 _4986_ (.A(_1746_),
    .B(_1738_),
    .C(_1750_),
    .Y(_0115_));
 sg13g2_nor3_1 _4987_ (.A(_1748_),
    .B(_1738_),
    .C(_1750_),
    .Y(_0116_));
 sg13g2_and2_1 _4988_ (.A(\btn.long_press ),
    .B(_1751_),
    .X(_0117_));
 sg13g2_inv_1 _4989_ (.Y(_1752_),
    .A(_1710_));
 sg13g2_a21oi_1 _4990_ (.A1(net43),
    .A2(_1752_),
    .Y(_1753_),
    .B1(\btn.long_press ));
 sg13g2_nor2_1 _4991_ (.A(_1740_),
    .B(_1753_),
    .Y(_0118_));
 sg13g2_buf_1 _4992_ (.A(_1665_),
    .X(_1754_));
 sg13g2_nand2_1 _4993_ (.Y(_1755_),
    .A(\btn.sample_5ms[0] ),
    .B(net59));
 sg13g2_buf_1 _4994_ (.A(net88),
    .X(_1756_));
 sg13g2_nand2_1 _4995_ (.Y(_1757_),
    .A(\btn.sample_10ms[0] ),
    .B(net58));
 sg13g2_a21oi_1 _4996_ (.A1(_1755_),
    .A2(_1757_),
    .Y(_0119_),
    .B1(net73));
 sg13g2_nand2_1 _4997_ (.Y(_1758_),
    .A(\btn.sample_5ms[1] ),
    .B(net59));
 sg13g2_nand2_1 _4998_ (.Y(_1759_),
    .A(\btn.sample_10ms[1] ),
    .B(net58));
 sg13g2_a21oi_1 _4999_ (.A1(_1758_),
    .A2(_1759_),
    .Y(_0120_),
    .B1(net73));
 sg13g2_nand2_1 _5000_ (.Y(_1760_),
    .A(\btn.sample_5ms[2] ),
    .B(net59));
 sg13g2_nand2_1 _5001_ (.Y(_1761_),
    .A(\btn.sample_10ms[2] ),
    .B(net58));
 sg13g2_a21oi_1 _5002_ (.A1(_1760_),
    .A2(_1761_),
    .Y(_0121_),
    .B1(net73));
 sg13g2_nand2_1 _5003_ (.Y(_1762_),
    .A(\btn.sample_5ms[3] ),
    .B(net59));
 sg13g2_nand2_1 _5004_ (.Y(_1763_),
    .A(\btn.sample_10ms[3] ),
    .B(net58));
 sg13g2_a21oi_1 _5005_ (.A1(_1762_),
    .A2(_1763_),
    .Y(_0122_),
    .B1(net73));
 sg13g2_nand2_1 _5006_ (.Y(_1764_),
    .A(\btn.sample_10ms[0] ),
    .B(net59));
 sg13g2_nand2_1 _5007_ (.Y(_1765_),
    .A(\btn.sample_15ms[0] ),
    .B(_1756_));
 sg13g2_a21oi_1 _5008_ (.A1(_1764_),
    .A2(_1765_),
    .Y(_0123_),
    .B1(net73));
 sg13g2_nand2_1 _5009_ (.Y(_1766_),
    .A(\btn.sample_10ms[1] ),
    .B(_1754_));
 sg13g2_nand2_1 _5010_ (.Y(_1767_),
    .A(\btn.sample_15ms[1] ),
    .B(net58));
 sg13g2_a21oi_1 _5011_ (.A1(_1766_),
    .A2(_1767_),
    .Y(_0124_),
    .B1(net73));
 sg13g2_nand2_1 _5012_ (.Y(_1768_),
    .A(\btn.sample_10ms[2] ),
    .B(_1754_));
 sg13g2_nand2_1 _5013_ (.Y(_1769_),
    .A(\btn.sample_15ms[2] ),
    .B(_1756_));
 sg13g2_a21oi_1 _5014_ (.A1(_1768_),
    .A2(_1769_),
    .Y(_0125_),
    .B1(_2643_));
 sg13g2_nand2_1 _5015_ (.Y(_1770_),
    .A(\btn.sample_10ms[3] ),
    .B(net59));
 sg13g2_nand2_1 _5016_ (.Y(_1771_),
    .A(\btn.sample_15ms[3] ),
    .B(net58));
 sg13g2_a21oi_1 _5017_ (.A1(_1770_),
    .A2(_1771_),
    .Y(_0126_),
    .B1(net73));
 sg13g2_nor2_1 _5018_ (.A(\btn.sample_5ms[0] ),
    .B(net62),
    .Y(_1772_));
 sg13g2_nor2_1 _5019_ (.A(net61),
    .B(_1688_),
    .Y(_1773_));
 sg13g2_nor3_1 _5020_ (.A(net60),
    .B(_1772_),
    .C(_1773_),
    .Y(_0127_));
 sg13g2_nor2_1 _5021_ (.A(\btn.sample_5ms[1] ),
    .B(_1666_),
    .Y(_1774_));
 sg13g2_nor2_1 _5022_ (.A(net61),
    .B(_1684_),
    .Y(_1775_));
 sg13g2_nor3_1 _5023_ (.A(net60),
    .B(_1774_),
    .C(_1775_),
    .Y(_0128_));
 sg13g2_nor2_1 _5024_ (.A(\btn.sample_5ms[2] ),
    .B(_1666_),
    .Y(_1776_));
 sg13g2_nor2_1 _5025_ (.A(_1668_),
    .B(_1686_),
    .Y(_1777_));
 sg13g2_nor3_1 _5026_ (.A(net60),
    .B(_1776_),
    .C(_1777_),
    .Y(_0129_));
 sg13g2_nor2_1 _5027_ (.A(\btn.sample_5ms[3] ),
    .B(net62),
    .Y(_1778_));
 sg13g2_nor2_1 _5028_ (.A(_1668_),
    .B(_1690_),
    .Y(_1779_));
 sg13g2_nor3_1 _5029_ (.A(_1672_),
    .B(_1778_),
    .C(_1779_),
    .Y(_0130_));
 sg13g2_and2_1 _5030_ (.A(net66),
    .B(_0021_),
    .X(_0139_));
 sg13g2_buf_2 _5031_ (.A(\dsp.digit ),
    .X(_1780_));
 sg13g2_inv_1 _5032_ (.Y(_1781_),
    .A(_1780_));
 sg13g2_nor2_1 _5033_ (.A(_2641_),
    .B(net86),
    .Y(_0140_));
 sg13g2_buf_1 _5034_ (.A(display_graphical),
    .X(_1782_));
 sg13g2_buf_1 _5035_ (.A(_1782_),
    .X(_1783_));
 sg13g2_buf_2 _5036_ (.A(\display_value[2] ),
    .X(_1784_));
 sg13g2_inv_1 _5037_ (.Y(_1785_),
    .A(_1784_));
 sg13g2_nand2b_1 _5038_ (.Y(_1786_),
    .B(_0059_),
    .A_N(_0926_));
 sg13g2_o21ai_1 _5039_ (.B1(_0058_),
    .Y(_1787_),
    .A1(net116),
    .A2(_1786_));
 sg13g2_nand2_1 _5040_ (.Y(_1788_),
    .A(_0939_),
    .B(_1787_));
 sg13g2_nor2_1 _5041_ (.A(net116),
    .B(_0905_),
    .Y(_1789_));
 sg13g2_nand4_1 _5042_ (.B(_1782_),
    .C(_1788_),
    .A(_1785_),
    .Y(_1790_),
    .D(_1789_));
 sg13g2_o21ai_1 _5043_ (.B1(_1790_),
    .Y(_1791_),
    .A1(_0014_),
    .A2(net85));
 sg13g2_nor2_2 _5044_ (.A(_0939_),
    .B(_0926_),
    .Y(_1792_));
 sg13g2_nand2_1 _5045_ (.Y(_1793_),
    .A(_1784_),
    .B(_1792_));
 sg13g2_nor2_1 _5046_ (.A(net116),
    .B(_1793_),
    .Y(_1794_));
 sg13g2_buf_1 _5047_ (.A(_0905_),
    .X(_1795_));
 sg13g2_o21ai_1 _5048_ (.B1(net84),
    .Y(_1796_),
    .A1(_1782_),
    .A2(_1794_));
 sg13g2_nand3_1 _5049_ (.B(_1785_),
    .C(_1792_),
    .A(_0946_),
    .Y(_1797_));
 sg13g2_a21oi_1 _5050_ (.A1(_1783_),
    .A2(_1797_),
    .Y(_1798_),
    .B1(net86));
 sg13g2_a221oi_1 _5051_ (.B2(_1798_),
    .C1(net65),
    .B1(_1796_),
    .A1(net86),
    .Y(_0141_),
    .A2(_1791_));
 sg13g2_nor2_1 _5052_ (.A(net108),
    .B(_1780_),
    .Y(_1799_));
 sg13g2_o21ai_1 _5053_ (.B1(_1799_),
    .Y(_1800_),
    .A1(net85),
    .A2(_0015_));
 sg13g2_and2_1 _5054_ (.A(_1784_),
    .B(_0939_),
    .X(_1801_));
 sg13g2_buf_1 _5055_ (.A(_1801_),
    .X(_1802_));
 sg13g2_nand2_1 _5056_ (.Y(_1803_),
    .A(_1782_),
    .B(_1789_));
 sg13g2_a21oi_1 _5057_ (.A1(_1787_),
    .A2(_1802_),
    .Y(_1804_),
    .B1(_1803_));
 sg13g2_inv_2 _5058_ (.Y(_1805_),
    .A(_1782_));
 sg13g2_nand2_1 _5059_ (.Y(_1806_),
    .A(_0058_),
    .B(_1786_));
 sg13g2_a21oi_1 _5060_ (.A1(_0939_),
    .A2(_1806_),
    .Y(_1807_),
    .B1(_1784_));
 sg13g2_inv_1 _5061_ (.Y(_1808_),
    .A(_0905_));
 sg13g2_o21ai_1 _5062_ (.B1(_1808_),
    .Y(_1809_),
    .A1(_0946_),
    .A2(_1807_));
 sg13g2_nand3b_1 _5063_ (.B(_0058_),
    .C(_1784_),
    .Y(_1810_),
    .A_N(_0939_));
 sg13g2_nand2_1 _5064_ (.Y(_1811_),
    .A(_0908_),
    .B(_1810_));
 sg13g2_nand3_1 _5065_ (.B(_1793_),
    .C(_1811_),
    .A(_0946_),
    .Y(_1812_));
 sg13g2_nand2_1 _5066_ (.Y(_1813_),
    .A(net84),
    .B(_1812_));
 sg13g2_nand2_1 _5067_ (.Y(_1814_),
    .A(_1809_),
    .B(_1813_));
 sg13g2_nand2_1 _5068_ (.Y(_1815_),
    .A(net84),
    .B(_1794_));
 sg13g2_nand3_1 _5069_ (.B(_1814_),
    .C(_1815_),
    .A(_1805_),
    .Y(_1816_));
 sg13g2_nand2_1 _5070_ (.Y(_1817_),
    .A(_0908_),
    .B(_1793_));
 sg13g2_nand3_1 _5071_ (.B(_0059_),
    .C(_1792_),
    .A(_1784_),
    .Y(_1818_));
 sg13g2_nand4_1 _5072_ (.B(_1789_),
    .C(_1817_),
    .A(net85),
    .Y(_1819_),
    .D(_1818_));
 sg13g2_nand3_1 _5073_ (.B(_1816_),
    .C(_1819_),
    .A(_0140_),
    .Y(_1820_));
 sg13g2_o21ai_1 _5074_ (.B1(_1820_),
    .Y(_0142_),
    .A1(_1800_),
    .A2(_1804_));
 sg13g2_nand3_1 _5075_ (.B(_1805_),
    .C(_1812_),
    .A(net84),
    .Y(_1821_));
 sg13g2_nand3_1 _5076_ (.B(_1809_),
    .C(_1821_),
    .A(_1780_),
    .Y(_1822_));
 sg13g2_nor2_1 _5077_ (.A(_1782_),
    .B(_0016_),
    .Y(_1823_));
 sg13g2_a21oi_1 _5078_ (.A1(_1811_),
    .A2(_1818_),
    .Y(_1824_),
    .B1(_0946_));
 sg13g2_nor3_1 _5079_ (.A(net84),
    .B(_1805_),
    .C(_1824_),
    .Y(_1825_));
 sg13g2_or3_1 _5080_ (.A(_1780_),
    .B(_1823_),
    .C(_1825_),
    .X(_1826_));
 sg13g2_buf_1 _5081_ (.A(net108),
    .X(_1827_));
 sg13g2_a21oi_1 _5082_ (.A1(_1822_),
    .A2(_1826_),
    .Y(_0143_),
    .B1(_1827_));
 sg13g2_nand3_1 _5083_ (.B(_1806_),
    .C(_1802_),
    .A(net116),
    .Y(_1828_));
 sg13g2_nand3b_1 _5084_ (.B(_1783_),
    .C(_1828_),
    .Y(_1829_),
    .A_N(_1795_));
 sg13g2_o21ai_1 _5085_ (.B1(_1829_),
    .Y(_1830_),
    .A1(net85),
    .A2(_0017_));
 sg13g2_nor2_1 _5086_ (.A(_1785_),
    .B(_1792_),
    .Y(_1831_));
 sg13g2_nor2_1 _5087_ (.A(_0946_),
    .B(_1805_),
    .Y(_1832_));
 sg13g2_a21oi_1 _5088_ (.A1(_1831_),
    .A2(_1832_),
    .Y(_1833_),
    .B1(_1781_));
 sg13g2_a221oi_1 _5089_ (.B2(_1796_),
    .C1(_1012_),
    .B1(_1833_),
    .A1(net86),
    .Y(_0144_),
    .A2(_1830_));
 sg13g2_nand2_1 _5090_ (.Y(_1834_),
    .A(_1785_),
    .B(_1792_));
 sg13g2_a21oi_1 _5091_ (.A1(net116),
    .A2(_1834_),
    .Y(_1835_),
    .B1(net84));
 sg13g2_o21ai_1 _5092_ (.B1(_1815_),
    .Y(_1836_),
    .A1(_1805_),
    .A2(_1835_));
 sg13g2_nand2_1 _5093_ (.Y(_1837_),
    .A(_0939_),
    .B(_0926_));
 sg13g2_o21ai_1 _5094_ (.B1(_0053_),
    .Y(_1838_),
    .A1(_1784_),
    .A2(_1837_));
 sg13g2_a21oi_1 _5095_ (.A1(_0945_),
    .A2(_1838_),
    .Y(_1839_),
    .B1(net84));
 sg13g2_nor2_1 _5096_ (.A(_1805_),
    .B(_1839_),
    .Y(_1840_));
 sg13g2_a21oi_1 _5097_ (.A1(_1805_),
    .A2(_0018_),
    .Y(_1841_),
    .B1(_1840_));
 sg13g2_nor2_1 _5098_ (.A(_1780_),
    .B(_1841_),
    .Y(_1842_));
 sg13g2_a21oi_1 _5099_ (.A1(_1780_),
    .A2(_1836_),
    .Y(_1843_),
    .B1(_1842_));
 sg13g2_nor2_1 _5100_ (.A(net63),
    .B(_1843_),
    .Y(_0145_));
 sg13g2_a21oi_1 _5101_ (.A1(net86),
    .A2(_0019_),
    .Y(_1844_),
    .B1(net85));
 sg13g2_nor3_1 _5102_ (.A(_1780_),
    .B(_1803_),
    .C(_1831_),
    .Y(_1845_));
 sg13g2_nor4_1 _5103_ (.A(net116),
    .B(_1795_),
    .C(net86),
    .D(_1838_),
    .Y(_1846_));
 sg13g2_nor4_1 _5104_ (.A(net92),
    .B(_1844_),
    .C(_1845_),
    .D(_1846_),
    .Y(_0146_));
 sg13g2_o21ai_1 _5105_ (.B1(net116),
    .Y(_1847_),
    .A1(_0059_),
    .A2(_1834_));
 sg13g2_nand3b_1 _5106_ (.B(net85),
    .C(_1847_),
    .Y(_1848_),
    .A_N(net84));
 sg13g2_o21ai_1 _5107_ (.B1(_1848_),
    .Y(_1849_),
    .A1(net85),
    .A2(_0020_));
 sg13g2_a21oi_1 _5108_ (.A1(_0926_),
    .A2(_1802_),
    .Y(_1850_),
    .B1(net116));
 sg13g2_nor2_1 _5109_ (.A(_1805_),
    .B(_1850_),
    .Y(_1851_));
 sg13g2_nor2_1 _5110_ (.A(net86),
    .B(_1851_),
    .Y(_1852_));
 sg13g2_a221oi_1 _5111_ (.B2(_1796_),
    .C1(_1012_),
    .B1(_1852_),
    .A1(net86),
    .Y(_0147_),
    .A2(_1849_));
 sg13g2_nor2_1 _5112_ (.A(_0869_),
    .B(_1631_),
    .Y(_1853_));
 sg13g2_buf_1 _5113_ (.A(_0871_),
    .X(_1854_));
 sg13g2_nand2_1 _5114_ (.Y(_1855_),
    .A(_0885_),
    .B(_0887_));
 sg13g2_buf_1 _5115_ (.A(_0889_),
    .X(_1856_));
 sg13g2_buf_1 _5116_ (.A(_0034_),
    .X(_1857_));
 sg13g2_nand2_2 _5117_ (.Y(_1858_),
    .A(_0890_),
    .B(_1857_));
 sg13g2_nor2_1 _5118_ (.A(net82),
    .B(_1858_),
    .Y(_1859_));
 sg13g2_nor2b_1 _5119_ (.A(_1855_),
    .B_N(_1859_),
    .Y(_1860_));
 sg13g2_buf_1 _5120_ (.A(net120),
    .X(_1861_));
 sg13g2_inv_1 _5121_ (.Y(_1862_),
    .A(net81));
 sg13g2_o21ai_1 _5122_ (.B1(_1862_),
    .Y(_1863_),
    .A1(net83),
    .A2(_1860_));
 sg13g2_nand3b_1 _5123_ (.B(net89),
    .C(_1863_),
    .Y(_1864_),
    .A_N(_1853_));
 sg13g2_nand2b_1 _5124_ (.Y(_1865_),
    .B(_1864_),
    .A_N(net90));
 sg13g2_o21ai_1 _5125_ (.B1(_0973_),
    .Y(_1866_),
    .A1(_0881_),
    .A2(_1865_));
 sg13g2_nor4_1 _5126_ (.A(net81),
    .B(net83),
    .C(_0893_),
    .D(_1865_),
    .Y(_1867_));
 sg13g2_nor2_1 _5127_ (.A(\game.challenge_mode ),
    .B(_1867_),
    .Y(_1868_));
 sg13g2_nor2_1 _5128_ (.A(_1866_),
    .B(_1868_),
    .Y(_0148_));
 sg13g2_nand2b_1 _5129_ (.Y(_1869_),
    .B(_0893_),
    .A_N(net89));
 sg13g2_buf_1 _5130_ (.A(_0886_),
    .X(_1870_));
 sg13g2_nor2_2 _5131_ (.A(_0885_),
    .B(_1870_),
    .Y(_1871_));
 sg13g2_nand4_1 _5132_ (.B(_0890_),
    .C(_1857_),
    .A(_1856_),
    .Y(_1872_),
    .D(_1871_));
 sg13g2_buf_2 _5133_ (.A(_1872_),
    .X(_1873_));
 sg13g2_buf_1 _5134_ (.A(_0885_),
    .X(_1874_));
 sg13g2_nor2_1 _5135_ (.A(_0887_),
    .B(net117),
    .Y(_1875_));
 sg13g2_nand3_1 _5136_ (.B(_0891_),
    .C(_1875_),
    .A(net79),
    .Y(_1876_));
 sg13g2_nand3_1 _5137_ (.B(_1873_),
    .C(_1876_),
    .A(_0913_),
    .Y(_1877_));
 sg13g2_nand3_1 _5138_ (.B(_1869_),
    .C(_1877_),
    .A(_0877_),
    .Y(_1878_));
 sg13g2_buf_2 _5139_ (.A(_1878_),
    .X(_1879_));
 sg13g2_buf_1 _5140_ (.A(_0864_),
    .X(_1880_));
 sg13g2_inv_1 _5141_ (.Y(_1881_),
    .A(_0889_));
 sg13g2_nor4_1 _5142_ (.A(net79),
    .B(net80),
    .C(_1881_),
    .D(_1858_),
    .Y(_1882_));
 sg13g2_buf_2 _5143_ (.A(_1882_),
    .X(_1883_));
 sg13g2_nor2_1 _5144_ (.A(net78),
    .B(_1883_),
    .Y(_1884_));
 sg13g2_nor2_1 _5145_ (.A(_0867_),
    .B(_0868_),
    .Y(_1885_));
 sg13g2_and3_1 _5146_ (.X(_1886_),
    .A(_1880_),
    .B(_0867_),
    .C(_1883_));
 sg13g2_buf_1 _5147_ (.A(_1886_),
    .X(_1887_));
 sg13g2_a22oi_1 _5148_ (.Y(_1888_),
    .B1(_1887_),
    .B2(_0868_),
    .A2(_1885_),
    .A1(_1884_));
 sg13g2_o21ai_1 _5149_ (.B1(_0931_),
    .Y(_1889_),
    .A1(net47),
    .A2(_1888_));
 sg13g2_nor3_1 _5150_ (.A(net96),
    .B(_1889_),
    .C(_1879_),
    .Y(_1890_));
 sg13g2_a21oi_1 _5151_ (.A1(net96),
    .A2(_1879_),
    .Y(_1891_),
    .B1(_1890_));
 sg13g2_nor2_1 _5152_ (.A(net63),
    .B(_1891_),
    .Y(_0149_));
 sg13g2_inv_1 _5153_ (.Y(_1892_),
    .A(_1880_));
 sg13g2_nor3_1 _5154_ (.A(_1892_),
    .B(net96),
    .C(_0899_),
    .Y(_1893_));
 sg13g2_o21ai_1 _5155_ (.B1(_0913_),
    .Y(_1894_),
    .A1(_1893_),
    .A2(_1873_));
 sg13g2_nor3_1 _5156_ (.A(net47),
    .B(_0934_),
    .C(_1883_),
    .Y(_1895_));
 sg13g2_a21oi_1 _5157_ (.A1(_0934_),
    .A2(_1894_),
    .Y(_1896_),
    .B1(_1895_));
 sg13g2_nor3_1 _5158_ (.A(net40),
    .B(_1879_),
    .C(_1896_),
    .Y(_1897_));
 sg13g2_a21oi_1 _5159_ (.A1(net78),
    .A2(_1879_),
    .Y(_1898_),
    .B1(_1897_));
 sg13g2_nor2_1 _5160_ (.A(_1418_),
    .B(_1898_),
    .Y(_0150_));
 sg13g2_nand3_1 _5161_ (.B(_0914_),
    .C(_1883_),
    .A(net78),
    .Y(_1899_));
 sg13g2_o21ai_1 _5162_ (.B1(_1899_),
    .Y(_1900_),
    .A1(net78),
    .A2(_0914_));
 sg13g2_nor3_1 _5163_ (.A(net78),
    .B(net96),
    .C(_1883_),
    .Y(_1901_));
 sg13g2_a21oi_1 _5164_ (.A1(_0866_),
    .A2(_0899_),
    .Y(_1902_),
    .B1(_1873_));
 sg13g2_nor2_1 _5165_ (.A(net78),
    .B(_1885_),
    .Y(_1903_));
 sg13g2_a221oi_1 _5166_ (.B2(_1873_),
    .C1(_0914_),
    .B1(_1903_),
    .A1(net78),
    .Y(_1904_),
    .A2(_1902_));
 sg13g2_a221oi_1 _5167_ (.B2(_0914_),
    .C1(_1904_),
    .B1(_1901_),
    .A1(net96),
    .Y(_1905_),
    .A2(_1900_));
 sg13g2_nor2_1 _5168_ (.A(_0933_),
    .B(_1905_),
    .Y(_1906_));
 sg13g2_nor2_1 _5169_ (.A(_0917_),
    .B(_1906_),
    .Y(_1907_));
 sg13g2_nor2_1 _5170_ (.A(_1879_),
    .B(_1907_),
    .Y(_1908_));
 sg13g2_a21oi_1 _5171_ (.A1(_0867_),
    .A2(_1879_),
    .Y(_1909_),
    .B1(_1908_));
 sg13g2_nor2_1 _5172_ (.A(_1418_),
    .B(_1909_),
    .Y(_0151_));
 sg13g2_mux2_1 _5173_ (.A0(_1892_),
    .A1(_1887_),
    .S(_0947_),
    .X(_1910_));
 sg13g2_nor2b_1 _5174_ (.A(_0867_),
    .B_N(_0947_),
    .Y(_1911_));
 sg13g2_nor3_1 _5175_ (.A(net78),
    .B(_0867_),
    .C(_1883_),
    .Y(_1912_));
 sg13g2_or2_1 _5176_ (.X(_1913_),
    .B(_0868_),
    .A(_0922_));
 sg13g2_o21ai_1 _5177_ (.B1(_1913_),
    .Y(_1914_),
    .A1(_1887_),
    .A2(_1912_));
 sg13g2_nor2b_1 _5178_ (.A(_0947_),
    .B_N(_1914_),
    .Y(_1915_));
 sg13g2_a221oi_1 _5179_ (.B2(_1901_),
    .C1(_1915_),
    .B1(_1911_),
    .A1(_0922_),
    .Y(_1916_),
    .A2(_1910_));
 sg13g2_o21ai_1 _5180_ (.B1(_0955_),
    .Y(_1917_),
    .A1(net47),
    .A2(_1916_));
 sg13g2_nor2_1 _5181_ (.A(_1879_),
    .B(_1917_),
    .Y(_1918_));
 sg13g2_nor2b_1 _5182_ (.A(_0868_),
    .B_N(_1879_),
    .Y(_1919_));
 sg13g2_nor3_1 _5183_ (.A(_1672_),
    .B(_1918_),
    .C(_1919_),
    .Y(_0152_));
 sg13g2_buf_1 _5184_ (.A(\game.counter[0] ),
    .X(_1920_));
 sg13g2_nor2b_1 _5185_ (.A(\game.solver_trigger_delayed ),
    .B_N(\game.slv.ready ),
    .Y(_1921_));
 sg13g2_nand2_1 _5186_ (.Y(_1922_),
    .A(_1854_),
    .B(_1921_));
 sg13g2_o21ai_1 _5187_ (.B1(_1922_),
    .Y(_1923_),
    .A1(net83),
    .A2(net115));
 sg13g2_a22oi_1 _5188_ (.Y(_1924_),
    .B1(_1923_),
    .B2(_1861_),
    .A2(_1618_),
    .A1(_1644_));
 sg13g2_buf_1 _5189_ (.A(_0890_),
    .X(_1925_));
 sg13g2_nor2_1 _5190_ (.A(_1881_),
    .B(net77),
    .Y(_1926_));
 sg13g2_buf_1 _5191_ (.A(_1857_),
    .X(_1927_));
 sg13g2_nand2b_1 _5192_ (.Y(_1928_),
    .B(net76),
    .A_N(net119));
 sg13g2_nand4_1 _5193_ (.B(_1871_),
    .C(_1926_),
    .A(_0879_),
    .Y(_1929_),
    .D(_1928_));
 sg13g2_o21ai_1 _5194_ (.B1(_1929_),
    .Y(_1930_),
    .A1(net89),
    .A2(_1924_));
 sg13g2_nand2b_1 _5195_ (.Y(_1931_),
    .B(_1930_),
    .A_N(net90));
 sg13g2_buf_1 _5196_ (.A(_1931_),
    .X(_1932_));
 sg13g2_nor2_1 _5197_ (.A(net44),
    .B(_1632_),
    .Y(_1933_));
 sg13g2_inv_1 _5198_ (.Y(_1934_),
    .A(net44));
 sg13g2_a21oi_1 _5199_ (.A1(_1934_),
    .A2(_1640_),
    .Y(_1935_),
    .B1(_1630_));
 sg13g2_nor2_1 _5200_ (.A(_1933_),
    .B(_1935_),
    .Y(_1936_));
 sg13g2_buf_2 _5201_ (.A(_1936_),
    .X(_1937_));
 sg13g2_nand2b_1 _5202_ (.Y(_1938_),
    .B(_1937_),
    .A_N(_1931_));
 sg13g2_buf_1 _5203_ (.A(_1938_),
    .X(_1939_));
 sg13g2_nor2_1 _5204_ (.A(net114),
    .B(_1939_),
    .Y(_1940_));
 sg13g2_a21oi_1 _5205_ (.A1(net114),
    .A2(net27),
    .Y(_1941_),
    .B1(_1940_));
 sg13g2_nor2_1 _5206_ (.A(net63),
    .B(_1941_),
    .Y(_0153_));
 sg13g2_buf_2 _5207_ (.A(\game.counter[1] ),
    .X(_1942_));
 sg13g2_nand2b_1 _5208_ (.Y(_1943_),
    .B(net114),
    .A_N(_1942_));
 sg13g2_nand2b_1 _5209_ (.Y(_1944_),
    .B(_1942_),
    .A_N(net114));
 sg13g2_o21ai_1 _5210_ (.B1(_1944_),
    .Y(_1945_),
    .A1(net27),
    .A2(_1943_));
 sg13g2_a22oi_1 _5211_ (.Y(_1946_),
    .B1(_1937_),
    .B2(_1945_),
    .A2(net27),
    .A1(_1942_));
 sg13g2_nor2_1 _5212_ (.A(net63),
    .B(_1946_),
    .Y(_0154_));
 sg13g2_nand2_1 _5213_ (.Y(_1947_),
    .A(_1942_),
    .B(_1920_));
 sg13g2_nor3_1 _5214_ (.A(_1626_),
    .B(net27),
    .C(_1947_),
    .Y(_1948_));
 sg13g2_a21o_1 _5215_ (.A2(_1947_),
    .A1(_1626_),
    .B1(_1948_),
    .X(_1949_));
 sg13g2_a22oi_1 _5216_ (.Y(_1950_),
    .B1(_1937_),
    .B2(_1949_),
    .A2(net27),
    .A1(_1626_));
 sg13g2_nor2_1 _5217_ (.A(net63),
    .B(_1950_),
    .Y(_0155_));
 sg13g2_nand3_1 _5218_ (.B(_1942_),
    .C(net114),
    .A(_1626_),
    .Y(_1951_));
 sg13g2_buf_1 _5219_ (.A(_1951_),
    .X(_1952_));
 sg13g2_a21o_1 _5220_ (.A2(_1952_),
    .A1(_1937_),
    .B1(net27),
    .X(_1953_));
 sg13g2_nor3_1 _5221_ (.A(_1627_),
    .B(_1939_),
    .C(_1952_),
    .Y(_1954_));
 sg13g2_a21oi_1 _5222_ (.A1(_1627_),
    .A2(_1953_),
    .Y(_1955_),
    .B1(_1954_));
 sg13g2_nor2_1 _5223_ (.A(net63),
    .B(_1955_),
    .Y(_0156_));
 sg13g2_buf_1 _5224_ (.A(net92),
    .X(_1956_));
 sg13g2_nand4_1 _5225_ (.B(_1627_),
    .C(_1942_),
    .A(_1626_),
    .Y(_1957_),
    .D(net114));
 sg13g2_a21o_1 _5226_ (.A2(_1957_),
    .A1(_1937_),
    .B1(net27),
    .X(_1958_));
 sg13g2_nor3_1 _5227_ (.A(_1625_),
    .B(_1939_),
    .C(_1957_),
    .Y(_1959_));
 sg13g2_a21oi_1 _5228_ (.A1(_1625_),
    .A2(_1958_),
    .Y(_1960_),
    .B1(_1959_));
 sg13g2_nor2_1 _5229_ (.A(net56),
    .B(_1960_),
    .Y(_0157_));
 sg13g2_nand2_1 _5230_ (.Y(_1961_),
    .A(_1625_),
    .B(_1627_));
 sg13g2_nor2_1 _5231_ (.A(_1952_),
    .B(_1961_),
    .Y(_1962_));
 sg13g2_nor3_1 _5232_ (.A(_1933_),
    .B(_1935_),
    .C(_1962_),
    .Y(_1963_));
 sg13g2_o21ai_1 _5233_ (.B1(_1623_),
    .Y(_1964_),
    .A1(_1932_),
    .A2(_1963_));
 sg13g2_or4_1 _5234_ (.A(_1623_),
    .B(_1939_),
    .C(_1952_),
    .D(_1961_),
    .X(_1965_));
 sg13g2_a21oi_1 _5235_ (.A1(_1964_),
    .A2(_1965_),
    .Y(_0158_),
    .B1(net57));
 sg13g2_nand2_1 _5236_ (.Y(_1966_),
    .A(_1623_),
    .B(_1962_));
 sg13g2_a21o_1 _5237_ (.A2(_1966_),
    .A1(_1937_),
    .B1(net27),
    .X(_1967_));
 sg13g2_nor3_1 _5238_ (.A(_1622_),
    .B(_1939_),
    .C(_1966_),
    .Y(_1968_));
 sg13g2_a21oi_1 _5239_ (.A1(_1622_),
    .A2(_1967_),
    .Y(_1969_),
    .B1(_1968_));
 sg13g2_nor2_1 _5240_ (.A(_1956_),
    .B(_1969_),
    .Y(_0159_));
 sg13g2_nand3_1 _5241_ (.B(_1623_),
    .C(_1962_),
    .A(_1622_),
    .Y(_1970_));
 sg13g2_nor3_1 _5242_ (.A(_1629_),
    .B(_1931_),
    .C(_1970_),
    .Y(_1971_));
 sg13g2_a21o_1 _5243_ (.A2(_1970_),
    .A1(_1629_),
    .B1(_1971_),
    .X(_1972_));
 sg13g2_a22oi_1 _5244_ (.Y(_1973_),
    .B1(_1937_),
    .B2(_1972_),
    .A2(_1932_),
    .A1(_1629_));
 sg13g2_nor2_1 _5245_ (.A(_1956_),
    .B(_1973_),
    .Y(_0160_));
 sg13g2_nor2_1 _5246_ (.A(_0931_),
    .B(_1883_),
    .Y(_1974_));
 sg13g2_buf_2 _5247_ (.A(_1974_),
    .X(_1975_));
 sg13g2_nand3_1 _5248_ (.B(net89),
    .C(_1893_),
    .A(net81),
    .Y(_1976_));
 sg13g2_or2_1 _5249_ (.X(_1977_),
    .B(net119),
    .A(net120));
 sg13g2_buf_1 _5250_ (.A(_1977_),
    .X(_1978_));
 sg13g2_a221oi_1 _5251_ (.B2(_1978_),
    .C1(_0874_),
    .B1(_1976_),
    .A1(_1876_),
    .Y(_1979_),
    .A2(_1975_));
 sg13g2_buf_1 _5252_ (.A(_1979_),
    .X(_1980_));
 sg13g2_nand2b_1 _5253_ (.Y(_1981_),
    .B(net129),
    .A_N(net25));
 sg13g2_inv_1 _5254_ (.Y(_1982_),
    .A(_0069_));
 sg13g2_nor3_2 _5255_ (.A(net100),
    .B(_0567_),
    .C(_0680_),
    .Y(_1983_));
 sg13g2_nand3_1 _5256_ (.B(_1975_),
    .C(_1983_),
    .A(_0061_),
    .Y(_1984_));
 sg13g2_nor3_1 _5257_ (.A(net105),
    .B(_0493_),
    .C(_0848_),
    .Y(_1985_));
 sg13g2_nand2_2 _5258_ (.Y(_1986_),
    .A(_0949_),
    .B(_1873_));
 sg13g2_a22oi_1 _5259_ (.Y(_1987_),
    .B1(_1985_),
    .B2(_1986_),
    .A2(_1984_),
    .A1(_1982_));
 sg13g2_nand2_1 _5260_ (.Y(_1988_),
    .A(net25),
    .B(_1987_));
 sg13g2_a21oi_1 _5261_ (.A1(_1981_),
    .A2(_1988_),
    .Y(_0161_),
    .B1(net57));
 sg13g2_xnor2_1 _5262_ (.Y(_1989_),
    .A(net105),
    .B(_1975_));
 sg13g2_nand2_1 _5263_ (.Y(_1990_),
    .A(net25),
    .B(_1989_));
 sg13g2_xnor2_1 _5264_ (.Y(_1991_),
    .A(_0493_),
    .B(_1990_));
 sg13g2_nor2_1 _5265_ (.A(net56),
    .B(_1991_),
    .Y(_0162_));
 sg13g2_nor2_1 _5266_ (.A(net100),
    .B(_0680_),
    .Y(_1992_));
 sg13g2_o21ai_1 _5267_ (.B1(_1992_),
    .Y(_1993_),
    .A1(_0567_),
    .A2(_0896_));
 sg13g2_nand3_1 _5268_ (.B(net49),
    .C(_0848_),
    .A(_0063_),
    .Y(_1994_));
 sg13g2_o21ai_1 _5269_ (.B1(_1994_),
    .Y(_1995_),
    .A1(_0063_),
    .A2(net49));
 sg13g2_nand2_1 _5270_ (.Y(_1996_),
    .A(_1986_),
    .B(_1995_));
 sg13g2_o21ai_1 _5271_ (.B1(_1996_),
    .Y(_1997_),
    .A1(_1986_),
    .A2(_1993_));
 sg13g2_nand2_1 _5272_ (.Y(_1998_),
    .A(_0680_),
    .B(_1975_));
 sg13g2_nand2_1 _5273_ (.Y(_1999_),
    .A(net25),
    .B(_1998_));
 sg13g2_a22oi_1 _5274_ (.Y(_2000_),
    .B1(_1999_),
    .B2(net100),
    .A2(_1997_),
    .A1(net25));
 sg13g2_nor2_1 _5275_ (.A(net56),
    .B(_2000_),
    .Y(_0163_));
 sg13g2_o21ai_1 _5276_ (.B1(_0699_),
    .Y(_2001_),
    .A1(_0496_),
    .A2(_0847_));
 sg13g2_nand2_1 _5277_ (.Y(_2002_),
    .A(_0062_),
    .B(_0951_));
 sg13g2_o21ai_1 _5278_ (.B1(_2002_),
    .Y(_2003_),
    .A1(_0062_),
    .A2(_2001_));
 sg13g2_nand3_1 _5279_ (.B(_1975_),
    .C(_1983_),
    .A(_0896_),
    .Y(_2004_));
 sg13g2_o21ai_1 _5280_ (.B1(_2004_),
    .Y(_2005_),
    .A1(_1975_),
    .A2(_2003_));
 sg13g2_o21ai_1 _5281_ (.B1(net25),
    .Y(_2006_),
    .A1(_1986_),
    .A2(_1992_));
 sg13g2_a22oi_1 _5282_ (.Y(_2007_),
    .B1(_2006_),
    .B2(_0567_),
    .A2(_2005_),
    .A1(_1980_));
 sg13g2_nor2_1 _5283_ (.A(net56),
    .B(_2007_),
    .Y(_0164_));
 sg13g2_nand3_1 _5284_ (.B(_0896_),
    .C(_1983_),
    .A(\game.current_level[4] ),
    .Y(_2008_));
 sg13g2_nor2_1 _5285_ (.A(_0061_),
    .B(_0897_),
    .Y(_2009_));
 sg13g2_a21oi_1 _5286_ (.A1(net49),
    .A2(_0847_),
    .Y(_2010_),
    .B1(_0061_));
 sg13g2_o21ai_1 _5287_ (.B1(_1986_),
    .Y(_2011_),
    .A1(_0496_),
    .A2(_2010_));
 sg13g2_a21oi_1 _5288_ (.A1(_0567_),
    .A2(_0699_),
    .Y(_2012_),
    .B1(_0896_));
 sg13g2_nor3_1 _5289_ (.A(_2009_),
    .B(_2011_),
    .C(_2012_),
    .Y(_2013_));
 sg13g2_a21oi_1 _5290_ (.A1(_1975_),
    .A2(_2008_),
    .Y(_2014_),
    .B1(_2013_));
 sg13g2_o21ai_1 _5291_ (.B1(net25),
    .Y(_2015_),
    .A1(_1983_),
    .A2(_2013_));
 sg13g2_a221oi_1 _5292_ (.B2(_0565_),
    .C1(net65),
    .B1(_2015_),
    .A1(net25),
    .Y(_0165_),
    .A2(_2014_));
 sg13g2_o21ai_1 _5293_ (.B1(net95),
    .Y(_2016_),
    .A1(net85),
    .A2(_0901_));
 sg13g2_nor2_1 _5294_ (.A(_0895_),
    .B(_2016_),
    .Y(_0166_));
 sg13g2_nand2_1 _5295_ (.Y(_0167_),
    .A(net67),
    .B(_0963_));
 sg13g2_buf_1 _5296_ (.A(net134),
    .X(_2017_));
 sg13g2_o21ai_1 _5297_ (.B1(net75),
    .Y(_2018_),
    .A1(_1784_),
    .A2(net30));
 sg13g2_a21oi_1 _5298_ (.A1(net30),
    .A2(_0918_),
    .Y(_0169_),
    .B1(_2018_));
 sg13g2_nor2_1 _5299_ (.A(net82),
    .B(_1855_),
    .Y(_2019_));
 sg13g2_nor2_1 _5300_ (.A(_0890_),
    .B(_0884_),
    .Y(_2020_));
 sg13g2_nor2b_1 _5301_ (.A(_0885_),
    .B_N(_1857_),
    .Y(_2021_));
 sg13g2_xor2_1 _5302_ (.B(_0890_),
    .A(_0889_),
    .X(_2022_));
 sg13g2_mux2_1 _5303_ (.A0(_0891_),
    .A1(_2022_),
    .S(_0887_),
    .X(_2023_));
 sg13g2_a22oi_1 _5304_ (.Y(_2024_),
    .B1(_2021_),
    .B2(_2023_),
    .A2(_2020_),
    .A1(_2019_));
 sg13g2_nor2_1 _5305_ (.A(_0931_),
    .B(_1037_),
    .Y(_2025_));
 sg13g2_nor2b_1 _5306_ (.A(_2024_),
    .B_N(_2025_),
    .Y(_2026_));
 sg13g2_buf_1 _5307_ (.A(_2026_),
    .X(_2027_));
 sg13g2_nand2b_1 _5308_ (.Y(_2028_),
    .B(\game.input_color[0] ),
    .A_N(_2027_));
 sg13g2_nand2_1 _5309_ (.Y(_2029_),
    .A(_1881_),
    .B(net76));
 sg13g2_xnor2_1 _5310_ (.Y(_2030_),
    .A(net80),
    .B(net77));
 sg13g2_nor3_1 _5311_ (.A(net79),
    .B(_2029_),
    .C(_2030_),
    .Y(_2031_));
 sg13g2_nand2_1 _5312_ (.Y(_2032_),
    .A(_2027_),
    .B(_2031_));
 sg13g2_a21oi_1 _5313_ (.A1(_2028_),
    .A2(_2032_),
    .Y(_0268_),
    .B1(net57));
 sg13g2_buf_1 _5314_ (.A(net94),
    .X(_2033_));
 sg13g2_nand4_1 _5315_ (.B(_1871_),
    .C(_2022_),
    .A(net76),
    .Y(_2034_),
    .D(_2025_));
 sg13g2_o21ai_1 _5316_ (.B1(_2034_),
    .Y(_2035_),
    .A1(_1023_),
    .A2(_2027_));
 sg13g2_and2_1 _5317_ (.A(net55),
    .B(_2035_),
    .X(_0269_));
 sg13g2_and4_1 _5318_ (.A(_1881_),
    .B(net77),
    .C(net117),
    .D(_1871_),
    .X(_2036_));
 sg13g2_buf_1 _5319_ (.A(_2036_),
    .X(_2037_));
 sg13g2_inv_1 _5320_ (.Y(_2038_),
    .A(_2037_));
 sg13g2_nor2_1 _5321_ (.A(_0931_),
    .B(_1022_),
    .Y(_2039_));
 sg13g2_inv_1 _5322_ (.Y(_2040_),
    .A(_2039_));
 sg13g2_nor3_1 _5323_ (.A(net60),
    .B(_2038_),
    .C(_2040_),
    .Y(_0270_));
 sg13g2_xor2_1 _5324_ (.B(net117),
    .A(net80),
    .X(_2041_));
 sg13g2_nand3_1 _5325_ (.B(_0891_),
    .C(_2041_),
    .A(net79),
    .Y(_2042_));
 sg13g2_a21oi_1 _5326_ (.A1(_1873_),
    .A2(_2042_),
    .Y(_2043_),
    .B1(_0931_));
 sg13g2_or2_1 _5327_ (.X(_0271_),
    .B(_2043_),
    .A(_1866_));
 sg13g2_and2_1 _5328_ (.A(net55),
    .B(_2027_),
    .X(_0272_));
 sg13g2_nor2_1 _5329_ (.A(_0871_),
    .B(_1978_),
    .Y(_2044_));
 sg13g2_a21oi_1 _5330_ (.A1(net120),
    .A2(_0871_),
    .Y(_2045_),
    .B1(_0863_));
 sg13g2_a21oi_1 _5331_ (.A1(_0035_),
    .A2(_2045_),
    .Y(_2046_),
    .B1(net118));
 sg13g2_nor2_1 _5332_ (.A(_2044_),
    .B(_2046_),
    .Y(_2047_));
 sg13g2_buf_1 _5333_ (.A(_2047_),
    .X(_2048_));
 sg13g2_buf_2 _5334_ (.A(_0007_),
    .X(_2049_));
 sg13g2_buf_2 _5335_ (.A(_0008_),
    .X(_2050_));
 sg13g2_mux4_1 _5336_ (.S0(_2049_),
    .A0(_0419_),
    .A1(\game.fsm.seq[1][0] ),
    .A2(_0413_),
    .A3(_0416_),
    .S1(_2050_),
    .X(_2051_));
 sg13g2_mux4_1 _5337_ (.S0(_2050_),
    .A0(_0426_),
    .A1(_0424_),
    .A2(_0427_),
    .A3(_0425_),
    .S1(_2049_),
    .X(_2052_));
 sg13g2_mux2_1 _5338_ (.A0(_2051_),
    .A1(_2052_),
    .S(_0009_),
    .X(_2053_));
 sg13g2_buf_1 _5339_ (.A(_2053_),
    .X(_2054_));
 sg13g2_mux4_1 _5340_ (.S0(_2050_),
    .A0(_0389_),
    .A1(_2930_),
    .A2(_2926_),
    .A3(_2932_),
    .S1(_2049_),
    .X(_2055_));
 sg13g2_mux4_1 _5341_ (.S0(_2050_),
    .A0(_0404_),
    .A1(_0406_),
    .A2(_0393_),
    .A3(_0398_),
    .S1(_2049_),
    .X(_2056_));
 sg13g2_mux2_1 _5342_ (.A0(_2055_),
    .A1(_2056_),
    .S(_0009_),
    .X(_2057_));
 sg13g2_nor3_1 _5343_ (.A(_1626_),
    .B(_1942_),
    .C(net114),
    .Y(_2058_));
 sg13g2_nor3_1 _5344_ (.A(_1622_),
    .B(_1629_),
    .C(_1623_),
    .Y(_2059_));
 sg13g2_o21ai_1 _5345_ (.B1(_2059_),
    .Y(_2060_),
    .A1(_1961_),
    .A2(_2058_));
 sg13g2_nand2_1 _5346_ (.Y(_2061_),
    .A(_1632_),
    .B(_2060_));
 sg13g2_nor3_1 _5347_ (.A(_1640_),
    .B(_2057_),
    .C(_2061_),
    .Y(_2062_));
 sg13g2_nand2b_1 _5348_ (.Y(_2063_),
    .B(_2062_),
    .A_N(_2054_));
 sg13g2_o21ai_1 _5349_ (.B1(_2063_),
    .Y(_2064_),
    .A1(_0853_),
    .A2(_2040_));
 sg13g2_nand2b_1 _5350_ (.Y(_2065_),
    .B(_2048_),
    .A_N(net12));
 sg13g2_o21ai_1 _5351_ (.B1(_2065_),
    .Y(_2066_),
    .A1(_2048_),
    .A2(_2064_));
 sg13g2_nor2_1 _5352_ (.A(net56),
    .B(_2066_),
    .Y(_0273_));
 sg13g2_nor3_1 _5353_ (.A(net13),
    .B(_2044_),
    .C(_2046_),
    .Y(_2067_));
 sg13g2_a221oi_1 _5354_ (.B2(_2062_),
    .C1(_2048_),
    .B1(_2054_),
    .A1(_0853_),
    .Y(_2068_),
    .A2(_2039_));
 sg13g2_nor3_1 _5355_ (.A(net60),
    .B(_2067_),
    .C(_2068_),
    .Y(_0274_));
 sg13g2_nor2_1 _5356_ (.A(_1640_),
    .B(_2061_),
    .Y(_2069_));
 sg13g2_nand2_1 _5357_ (.Y(_2070_),
    .A(_2057_),
    .B(_2069_));
 sg13g2_nor2_1 _5358_ (.A(_2054_),
    .B(_2070_),
    .Y(_2071_));
 sg13g2_a21oi_1 _5359_ (.A1(net40),
    .A2(_1022_),
    .Y(_2072_),
    .B1(_2071_));
 sg13g2_nor2_1 _5360_ (.A(_2048_),
    .B(_2072_),
    .Y(_2073_));
 sg13g2_a21oi_1 _5361_ (.A1(net14),
    .A2(_2048_),
    .Y(_2074_),
    .B1(_2073_));
 sg13g2_nand2_1 _5362_ (.Y(_0275_),
    .A(_0974_),
    .B(_2074_));
 sg13g2_nor3_1 _5363_ (.A(net15),
    .B(_2044_),
    .C(_2046_),
    .Y(_2075_));
 sg13g2_inv_1 _5364_ (.Y(_2076_),
    .A(_2070_));
 sg13g2_a221oi_1 _5365_ (.B2(_2076_),
    .C1(_2048_),
    .B1(_2054_),
    .A1(net40),
    .Y(_2077_),
    .A2(_1037_));
 sg13g2_nor3_1 _5366_ (.A(net60),
    .B(_2075_),
    .C(_2077_),
    .Y(_0276_));
 sg13g2_inv_1 _5367_ (.Y(_2078_),
    .A(_1874_));
 sg13g2_nor2b_1 _5368_ (.A(net77),
    .B_N(_0884_),
    .Y(_2079_));
 sg13g2_a21oi_1 _5369_ (.A1(_1925_),
    .A2(net76),
    .Y(_2080_),
    .B1(_2079_));
 sg13g2_nand2_1 _5370_ (.Y(_2081_),
    .A(_2078_),
    .B(_2080_));
 sg13g2_or2_1 _5371_ (.X(_2082_),
    .B(net117),
    .A(_0890_));
 sg13g2_buf_1 _5372_ (.A(_2082_),
    .X(_2083_));
 sg13g2_xnor2_1 _5373_ (.Y(_2084_),
    .A(_1870_),
    .B(net82));
 sg13g2_a21oi_1 _5374_ (.A1(net79),
    .A2(_2083_),
    .Y(_2085_),
    .B1(_2084_));
 sg13g2_nand3b_1 _5375_ (.B(_1856_),
    .C(net80),
    .Y(_2086_),
    .A_N(net117));
 sg13g2_o21ai_1 _5376_ (.B1(_2086_),
    .Y(_2087_),
    .A1(net80),
    .A2(_2029_));
 sg13g2_a22oi_1 _5377_ (.Y(_2088_),
    .B1(_2087_),
    .B2(_2078_),
    .A2(_2019_),
    .A1(net117));
 sg13g2_nor2_1 _5378_ (.A(net77),
    .B(_2088_),
    .Y(_2089_));
 sg13g2_a21oi_1 _5379_ (.A1(_2081_),
    .A2(_2085_),
    .Y(_2090_),
    .B1(_2089_));
 sg13g2_nand2b_1 _5380_ (.Y(_2091_),
    .B(net40),
    .A_N(_2090_));
 sg13g2_o21ai_1 _5381_ (.B1(net82),
    .Y(_2092_),
    .A1(_1927_),
    .A2(_2079_));
 sg13g2_nand3b_1 _5382_ (.B(_1927_),
    .C(net80),
    .Y(_2093_),
    .A_N(_1925_));
 sg13g2_o21ai_1 _5383_ (.B1(_2093_),
    .Y(_2094_),
    .A1(net80),
    .A2(_2092_));
 sg13g2_and2_1 _5384_ (.A(_2078_),
    .B(_2094_),
    .X(_2095_));
 sg13g2_o21ai_1 _5385_ (.B1(_2083_),
    .Y(_2096_),
    .A1(net80),
    .A2(_1858_));
 sg13g2_a22oi_1 _5386_ (.Y(_2097_),
    .B1(_2096_),
    .B2(_1874_),
    .A2(_2020_),
    .A1(_0887_));
 sg13g2_nor2_1 _5387_ (.A(net82),
    .B(_2097_),
    .Y(_2098_));
 sg13g2_o21ai_1 _5388_ (.B1(_0913_),
    .Y(_2099_),
    .A1(_2095_),
    .A2(_2098_));
 sg13g2_a21oi_1 _5389_ (.A1(_2037_),
    .A2(_2039_),
    .Y(_2100_),
    .B1(_2027_));
 sg13g2_buf_2 _5390_ (.A(\game.sound_on ),
    .X(_2101_));
 sg13g2_nand3_1 _5391_ (.B(net83),
    .C(_2101_),
    .A(_1861_),
    .Y(_2102_));
 sg13g2_a21o_1 _5392_ (.A2(_2102_),
    .A1(_0911_),
    .B1(_0901_),
    .X(_2103_));
 sg13g2_nand4_1 _5393_ (.B(_2099_),
    .C(_2100_),
    .A(_2091_),
    .Y(_2104_),
    .D(_2103_));
 sg13g2_buf_1 _5394_ (.A(_2104_),
    .X(_2105_));
 sg13g2_nand2b_2 _5395_ (.Y(_2106_),
    .B(net119),
    .A_N(net118));
 sg13g2_nor3_1 _5396_ (.A(_1893_),
    .B(_2106_),
    .C(_1631_),
    .Y(_2107_));
 sg13g2_a21oi_1 _5397_ (.A1(\game.next_state[0] ),
    .A2(_2105_),
    .Y(_2108_),
    .B1(_2107_));
 sg13g2_nor2_1 _5398_ (.A(net56),
    .B(_2108_),
    .Y(_0277_));
 sg13g2_nor2_1 _5399_ (.A(_0933_),
    .B(_2105_),
    .Y(_2109_));
 sg13g2_a21oi_1 _5400_ (.A1(\game.next_state[2] ),
    .A2(_2105_),
    .Y(_2110_),
    .B1(_2109_));
 sg13g2_nor2_1 _5401_ (.A(net56),
    .B(_2110_),
    .Y(_0278_));
 sg13g2_inv_1 _5402_ (.Y(_2111_),
    .A(_0030_));
 sg13g2_nor3_1 _5403_ (.A(net91),
    .B(_0029_),
    .C(_2111_),
    .Y(_2112_));
 sg13g2_a21oi_1 _5404_ (.A1(_0854_),
    .A2(_2112_),
    .Y(_2113_),
    .B1(_0860_));
 sg13g2_o21ai_1 _5405_ (.B1(net66),
    .Y(_0281_),
    .A1(\game.slv.trigger ),
    .A2(_2113_));
 sg13g2_buf_1 _5406_ (.A(\game.slv.retries[0] ),
    .X(_2114_));
 sg13g2_nor3_1 _5407_ (.A(_2114_),
    .B(\game.slv.retries[1] ),
    .C(\game.slv.retries[2] ),
    .Y(_2115_));
 sg13g2_inv_1 _5408_ (.Y(_2116_),
    .A(_2115_));
 sg13g2_a21oi_1 _5409_ (.A1(\game.slv.length[2] ),
    .A2(\game.slv.length[1] ),
    .Y(_2117_),
    .B1(_2116_));
 sg13g2_xnor2_1 _5410_ (.Y(_2118_),
    .A(\game.slv.length[0] ),
    .B(_2117_));
 sg13g2_nand2_1 _5411_ (.Y(_2119_),
    .A(_2638_),
    .B(_2635_));
 sg13g2_o21ai_1 _5412_ (.B1(_2119_),
    .Y(_2120_),
    .A1(net91),
    .A2(_2118_));
 sg13g2_and2_1 _5413_ (.A(net94),
    .B(_2120_),
    .X(_2121_));
 sg13g2_and2_1 _5414_ (.A(net94),
    .B(\game.slv.length[0] ),
    .X(_2122_));
 sg13g2_nor2_1 _5415_ (.A(\game.slv.state[1] ),
    .B(_2638_),
    .Y(_2123_));
 sg13g2_nand2_1 _5416_ (.Y(_2124_),
    .A(_0029_),
    .B(_2123_));
 sg13g2_and3_1 _5417_ (.X(_2125_),
    .A(_0028_),
    .B(_2639_),
    .C(_2124_));
 sg13g2_buf_1 _5418_ (.A(_2125_),
    .X(_2126_));
 sg13g2_nand3_1 _5419_ (.B(_2639_),
    .C(_2124_),
    .A(_0028_),
    .Y(_2127_));
 sg13g2_buf_1 _5420_ (.A(_2127_),
    .X(_2128_));
 sg13g2_nor2_1 _5421_ (.A(net121),
    .B(_2128_),
    .Y(_2129_));
 sg13g2_and2_1 _5422_ (.A(_1519_),
    .B(_1520_),
    .X(_2130_));
 sg13g2_buf_8 _5423_ (.A(_2130_),
    .X(_2131_));
 sg13g2_a22oi_1 _5424_ (.Y(_2132_),
    .B1(_2129_),
    .B2(_2131_),
    .A2(_2126_),
    .A1(net91));
 sg13g2_buf_1 _5425_ (.A(_2132_),
    .X(_2133_));
 sg13g2_mux2_1 _5426_ (.A0(_2121_),
    .A1(_2122_),
    .S(_2133_),
    .X(_0283_));
 sg13g2_nand3_1 _5427_ (.B(\game.slv.length[0] ),
    .C(_2115_),
    .A(\game.slv.length[1] ),
    .Y(_2134_));
 sg13g2_a21o_1 _5428_ (.A2(_2115_),
    .A1(\game.slv.length[0] ),
    .B1(\game.slv.length[1] ),
    .X(_2135_));
 sg13g2_o21ai_1 _5429_ (.B1(_2135_),
    .Y(_2136_),
    .A1(\game.slv.length[2] ),
    .A2(_2134_));
 sg13g2_nand2_1 _5430_ (.Y(_2137_),
    .A(_2638_),
    .B(_2634_));
 sg13g2_o21ai_1 _5431_ (.B1(_2137_),
    .Y(_2138_),
    .A1(net91),
    .A2(_2136_));
 sg13g2_and2_1 _5432_ (.A(net94),
    .B(_2138_),
    .X(_2139_));
 sg13g2_and2_1 _5433_ (.A(net94),
    .B(\game.slv.length[1] ),
    .X(_2140_));
 sg13g2_mux2_1 _5434_ (.A0(_2139_),
    .A1(_2140_),
    .S(_2133_),
    .X(_0284_));
 sg13g2_inv_1 _5435_ (.Y(_2141_),
    .A(\game.slv.length[2] ));
 sg13g2_and2_1 _5436_ (.A(_2141_),
    .B(_2134_),
    .X(_2142_));
 sg13g2_nor2_1 _5437_ (.A(_2634_),
    .B(_2635_),
    .Y(_2143_));
 sg13g2_nand3b_1 _5438_ (.B(_0028_),
    .C(net91),
    .Y(_2144_),
    .A_N(_2633_));
 sg13g2_o21ai_1 _5439_ (.B1(net75),
    .Y(_2145_),
    .A1(_2143_),
    .A2(_2144_));
 sg13g2_a221oi_1 _5440_ (.B2(_0859_),
    .C1(_2145_),
    .B1(_2142_),
    .A1(_2141_),
    .Y(_0285_),
    .A2(_2133_));
 sg13g2_xnor2_1 _5441_ (.Y(_2146_),
    .A(\game.slv.lfsr[16] ),
    .B(\game.slv.lfsr[18] ));
 sg13g2_nand2_1 _5442_ (.Y(_0286_),
    .A(net67),
    .B(_2146_));
 sg13g2_nand2b_1 _5443_ (.Y(_0287_),
    .B(net67),
    .A_N(\game.slv.lfsr[7] ));
 sg13g2_nand2b_1 _5444_ (.Y(_0288_),
    .B(net67),
    .A_N(\game.slv.lfsr[8] ));
 sg13g2_nand2b_1 _5445_ (.Y(_0289_),
    .B(net67),
    .A_N(\game.slv.lfsr[9] ));
 sg13g2_nand2b_1 _5446_ (.Y(_0290_),
    .B(net67),
    .A_N(\game.slv.lfsr[10] ));
 sg13g2_buf_1 _5447_ (.A(net94),
    .X(_2147_));
 sg13g2_nand2b_1 _5448_ (.Y(_0291_),
    .B(net54),
    .A_N(\game.slv.lfsr[11] ));
 sg13g2_nand2b_1 _5449_ (.Y(_0292_),
    .B(net54),
    .A_N(\game.slv.lfsr[12] ));
 sg13g2_nand2b_1 _5450_ (.Y(_0293_),
    .B(net54),
    .A_N(\game.slv.lfsr[13] ));
 sg13g2_nand2b_1 _5451_ (.Y(_0294_),
    .B(net54),
    .A_N(\game.slv.lfsr[14] ));
 sg13g2_nand2b_1 _5452_ (.Y(_0295_),
    .B(_2147_),
    .A_N(\game.slv.lfsr[15] ));
 sg13g2_nand2b_1 _5453_ (.Y(_0296_),
    .B(_2147_),
    .A_N(\game.slv.lfsr[16] ));
 sg13g2_xnor2_1 _5454_ (.Y(_2148_),
    .A(\game.slv.lfsr[17] ),
    .B(\game.slv.lfsr[19] ));
 sg13g2_nand2_1 _5455_ (.Y(_0297_),
    .A(net67),
    .B(_2148_));
 sg13g2_nand2b_1 _5456_ (.Y(_0298_),
    .B(net54),
    .A_N(\game.slv.lfsr[17] ));
 sg13g2_xnor2_1 _5457_ (.Y(_2149_),
    .A(\game.slv.lfsr[18] ),
    .B(\game.slv.lfsr[20] ));
 sg13g2_nand2_1 _5458_ (.Y(_0299_),
    .A(net67),
    .B(_2149_));
 sg13g2_nand2b_1 _5459_ (.Y(_0300_),
    .B(net54),
    .A_N(_2635_));
 sg13g2_nand2b_1 _5460_ (.Y(_0301_),
    .B(net54),
    .A_N(_2634_));
 sg13g2_nand2b_1 _5461_ (.Y(_0302_),
    .B(net54),
    .A_N(_2633_));
 sg13g2_nand2b_1 _5462_ (.Y(_0303_),
    .B(net66),
    .A_N(\game.slv.lfsr[3] ));
 sg13g2_nand2b_1 _5463_ (.Y(_0304_),
    .B(_0988_),
    .A_N(\game.slv.lfsr[4] ));
 sg13g2_nand2b_1 _5464_ (.Y(_0305_),
    .B(net66),
    .A_N(\game.slv.lfsr[5] ));
 sg13g2_nand2b_1 _5465_ (.Y(_0306_),
    .B(_0988_),
    .A_N(\game.slv.lfsr[6] ));
 sg13g2_and2_1 _5466_ (.A(_1523_),
    .B(_2126_),
    .X(_2150_));
 sg13g2_nand2_1 _5467_ (.Y(_2151_),
    .A(_0855_),
    .B(net75));
 sg13g2_nor2_1 _5468_ (.A(net121),
    .B(_2118_),
    .Y(_2152_));
 sg13g2_a21oi_1 _5469_ (.A1(net121),
    .A2(_0056_),
    .Y(_2153_),
    .B1(_2152_));
 sg13g2_o21ai_1 _5470_ (.B1(_2119_),
    .Y(_2154_),
    .A1(net91),
    .A2(_2153_));
 sg13g2_nor3_1 _5471_ (.A(_2638_),
    .B(_0030_),
    .C(_0857_),
    .Y(_2155_));
 sg13g2_nor2_1 _5472_ (.A(_2128_),
    .B(_2155_),
    .Y(_2156_));
 sg13g2_nand4_1 _5473_ (.B(_1523_),
    .C(_2154_),
    .A(net75),
    .Y(_2157_),
    .D(_2156_));
 sg13g2_o21ai_1 _5474_ (.B1(_2157_),
    .Y(_0307_),
    .A1(_2150_),
    .A2(_2151_));
 sg13g2_nand2_1 _5475_ (.Y(_2158_),
    .A(\game.slv.pos[1] ),
    .B(net75));
 sg13g2_xnor2_1 _5476_ (.Y(_2159_),
    .A(_0855_),
    .B(\game.slv.pos[1] ));
 sg13g2_nor2_1 _5477_ (.A(net121),
    .B(_2136_),
    .Y(_2160_));
 sg13g2_a21oi_1 _5478_ (.A1(net121),
    .A2(_2159_),
    .Y(_2161_),
    .B1(_2160_));
 sg13g2_o21ai_1 _5479_ (.B1(_2137_),
    .Y(_2162_),
    .A1(_1510_),
    .A2(_2161_));
 sg13g2_nand4_1 _5480_ (.B(_1523_),
    .C(_2156_),
    .A(net75),
    .Y(_2163_),
    .D(_2162_));
 sg13g2_o21ai_1 _5481_ (.B1(_2163_),
    .Y(_0308_),
    .A1(_2150_),
    .A2(_2158_));
 sg13g2_nand2_1 _5482_ (.Y(_2164_),
    .A(_1013_),
    .B(_2142_));
 sg13g2_o21ai_1 _5483_ (.B1(\game.slv.pos[2] ),
    .Y(_2165_),
    .A1(_0855_),
    .A2(\game.slv.pos[1] ));
 sg13g2_nand3_1 _5484_ (.B(_0857_),
    .C(_2165_),
    .A(net121),
    .Y(_2166_));
 sg13g2_and3_1 _5485_ (.X(_2167_),
    .A(_0859_),
    .B(_2164_),
    .C(_2166_));
 sg13g2_a21oi_1 _5486_ (.A1(net91),
    .A2(_2633_),
    .Y(_2168_),
    .B1(_2167_));
 sg13g2_nor2_1 _5487_ (.A(net92),
    .B(_2168_),
    .Y(_2169_));
 sg13g2_and2_1 _5488_ (.A(\game.slv.pos[2] ),
    .B(net94),
    .X(_2170_));
 sg13g2_nand2_1 _5489_ (.Y(_2171_),
    .A(_1523_),
    .B(_2156_));
 sg13g2_mux2_1 _5490_ (.A0(_2169_),
    .A1(_2170_),
    .S(_2171_),
    .X(_0309_));
 sg13g2_inv_1 _5491_ (.Y(_2172_),
    .A(_2114_));
 sg13g2_nor3_1 _5492_ (.A(_2172_),
    .B(_1521_),
    .C(_2128_),
    .Y(_2173_));
 sg13g2_a221oi_1 _5493_ (.B2(_2131_),
    .C1(net65),
    .B1(_2173_),
    .A1(_2172_),
    .Y(_0311_),
    .A2(_2133_));
 sg13g2_nand4_1 _5494_ (.B(_2131_),
    .C(_2123_),
    .A(_2172_),
    .Y(_2174_),
    .D(_2126_));
 sg13g2_inv_1 _5495_ (.Y(_2175_),
    .A(\game.slv.retries[1] ));
 sg13g2_nor2_1 _5496_ (.A(net108),
    .B(_2175_),
    .Y(_2176_));
 sg13g2_nand2_1 _5497_ (.Y(_2177_),
    .A(_1519_),
    .B(_1520_));
 sg13g2_o21ai_1 _5498_ (.B1(_0859_),
    .Y(_2178_),
    .A1(_0858_),
    .A2(_2114_));
 sg13g2_nand4_1 _5499_ (.B(_2175_),
    .C(_2126_),
    .A(net134),
    .Y(_2179_),
    .D(_2178_));
 sg13g2_a21oi_1 _5500_ (.A1(_0859_),
    .A2(_2177_),
    .Y(_2180_),
    .B1(_2179_));
 sg13g2_a21o_1 _5501_ (.A2(_2176_),
    .A1(_2174_),
    .B1(_2180_),
    .X(_0312_));
 sg13g2_nor4_1 _5502_ (.A(_2114_),
    .B(\game.slv.retries[1] ),
    .C(_1521_),
    .D(_2128_),
    .Y(_2181_));
 sg13g2_a21oi_1 _5503_ (.A1(_2131_),
    .A2(_2181_),
    .Y(_2182_),
    .B1(net108));
 sg13g2_nor3_1 _5504_ (.A(_0858_),
    .B(_2114_),
    .C(\game.slv.retries[1] ),
    .Y(_2183_));
 sg13g2_nor2_1 _5505_ (.A(_1510_),
    .B(_2183_),
    .Y(_2184_));
 sg13g2_or4_1 _5506_ (.A(_2641_),
    .B(\game.slv.retries[2] ),
    .C(_2128_),
    .D(_2184_),
    .X(_2185_));
 sg13g2_a21oi_1 _5507_ (.A1(_0859_),
    .A2(_2177_),
    .Y(_2186_),
    .B1(_2185_));
 sg13g2_a21o_1 _5508_ (.A2(_2182_),
    .A1(\game.slv.retries[2] ),
    .B1(_2186_),
    .X(_0313_));
 sg13g2_mux2_1 _5509_ (.A0(\game.slv.target[0] ),
    .A1(_2635_),
    .S(\game.slv.target[1] ),
    .X(_2187_));
 sg13g2_nor2b_1 _5510_ (.A(\game.slv.trigger ),
    .B_N(\game.slv.saved_target ),
    .Y(_2188_));
 sg13g2_a21oi_1 _5511_ (.A1(\game.slv.trigger ),
    .A2(_2187_),
    .Y(_2189_),
    .B1(_2188_));
 sg13g2_nor2_1 _5512_ (.A(net56),
    .B(_2189_),
    .Y(_0314_));
 sg13g2_buf_1 _5513_ (.A(net92),
    .X(_2190_));
 sg13g2_nand2_1 _5514_ (.Y(_2191_),
    .A(\game.slv.ready ),
    .B(_1527_));
 sg13g2_a22oi_1 _5515_ (.Y(_2192_),
    .B1(_2191_),
    .B2(_1017_),
    .A2(_1527_),
    .A1(\game.solver_trigger_delayed ));
 sg13g2_nor2_1 _5516_ (.A(net53),
    .B(_2192_),
    .Y(_0315_));
 sg13g2_nor3_1 _5517_ (.A(_1881_),
    .B(_1855_),
    .C(_2083_),
    .Y(_2193_));
 sg13g2_a21o_1 _5518_ (.A2(_1859_),
    .A1(_0888_),
    .B1(_2193_),
    .X(_2194_));
 sg13g2_buf_1 _5519_ (.A(_2194_),
    .X(_2195_));
 sg13g2_nand3_1 _5520_ (.B(_1525_),
    .C(_0869_),
    .A(net81),
    .Y(_2196_));
 sg13g2_a21oi_1 _5521_ (.A1(_1978_),
    .A2(_2196_),
    .Y(_2197_),
    .B1(_0874_));
 sg13g2_o21ai_1 _5522_ (.B1(_2197_),
    .Y(_2198_),
    .A1(_0950_),
    .A2(_2195_));
 sg13g2_nand2_1 _5523_ (.Y(_2199_),
    .A(\game.slv.target[0] ),
    .B(_2198_));
 sg13g2_nand3_1 _5524_ (.B(_0888_),
    .C(_1859_),
    .A(_0949_),
    .Y(_2200_));
 sg13g2_a21oi_1 _5525_ (.A1(_2199_),
    .A2(_2200_),
    .Y(_0316_),
    .B1(net57));
 sg13g2_inv_1 _5526_ (.Y(_2201_),
    .A(\game.slv.target[1] ));
 sg13g2_a221oi_1 _5527_ (.B2(_2201_),
    .C1(net65),
    .B1(_2198_),
    .A1(net40),
    .Y(_0317_),
    .A2(_2195_));
 sg13g2_nor2_1 _5528_ (.A(_0950_),
    .B(_2195_),
    .Y(_2202_));
 sg13g2_nand2b_1 _5529_ (.Y(_2203_),
    .B(net83),
    .A_N(net89));
 sg13g2_o21ai_1 _5530_ (.B1(_2203_),
    .Y(_2204_),
    .A1(net83),
    .A2(_0870_));
 sg13g2_a21oi_1 _5531_ (.A1(net81),
    .A2(_2204_),
    .Y(_2205_),
    .B1(_2044_));
 sg13g2_nor3_1 _5532_ (.A(net90),
    .B(_2202_),
    .C(_2205_),
    .Y(_2206_));
 sg13g2_nor2_1 _5533_ (.A(\game.solver_trigger_delayed ),
    .B(_2206_),
    .Y(_2207_));
 sg13g2_nor3_1 _5534_ (.A(net92),
    .B(_1527_),
    .C(_2207_),
    .Y(_0319_));
 sg13g2_or2_1 _5535_ (.X(_2208_),
    .B(net89),
    .A(net83));
 sg13g2_o21ai_1 _5536_ (.B1(_2208_),
    .Y(_2209_),
    .A1(net90),
    .A2(net115));
 sg13g2_nor2_1 _5537_ (.A(_1524_),
    .B(_2045_),
    .Y(_2210_));
 sg13g2_a21oi_2 _5538_ (.B1(_2210_),
    .Y(_2211_),
    .A2(_2209_),
    .A1(_1862_));
 sg13g2_buf_1 _5539_ (.A(\game.sound_mode[0] ),
    .X(_2212_));
 sg13g2_buf_1 _5540_ (.A(\snd.sequencer_state[1] ),
    .X(_2213_));
 sg13g2_buf_1 _5541_ (.A(\snd.sequencer_state[0] ),
    .X(_2214_));
 sg13g2_or2_1 _5542_ (.X(_2215_),
    .B(_2214_),
    .A(net112));
 sg13g2_nor3_2 _5543_ (.A(_2106_),
    .B(_1526_),
    .C(_2215_),
    .Y(_2216_));
 sg13g2_nand2_1 _5544_ (.Y(_2217_),
    .A(\game.tune[0] ),
    .B(_2216_));
 sg13g2_a221oi_1 _5545_ (.B2(_2217_),
    .C1(_0013_),
    .B1(_2099_),
    .A1(_0881_),
    .Y(_2218_),
    .A2(_1631_));
 sg13g2_a221oi_1 _5546_ (.B2(_2212_),
    .C1(_2218_),
    .B1(_2211_),
    .A1(_2101_),
    .Y(_2219_),
    .A2(net40));
 sg13g2_nor2_1 _5547_ (.A(net53),
    .B(_2219_),
    .Y(_0320_));
 sg13g2_buf_1 _5548_ (.A(\game.sound_mode[1] ),
    .X(_2220_));
 sg13g2_inv_1 _5549_ (.Y(_2221_),
    .A(_2220_));
 sg13g2_nor4_1 _5550_ (.A(_0437_),
    .B(_0421_),
    .C(_2024_),
    .D(_2037_),
    .Y(_2222_));
 sg13g2_a21oi_1 _5551_ (.A1(_1022_),
    .A2(_2037_),
    .Y(_2223_),
    .B1(_2222_));
 sg13g2_nand4_1 _5552_ (.B(_2024_),
    .C(_2038_),
    .A(_2101_),
    .Y(_2224_),
    .D(_2090_));
 sg13g2_o21ai_1 _5553_ (.B1(_2224_),
    .Y(_2225_),
    .A1(_0013_),
    .A2(_2223_));
 sg13g2_a21oi_1 _5554_ (.A1(net40),
    .A2(_2225_),
    .Y(_2226_),
    .B1(_2211_));
 sg13g2_inv_1 _5555_ (.Y(_2227_),
    .A(\game.tune[1] ));
 sg13g2_nor2_1 _5556_ (.A(_0013_),
    .B(_2227_),
    .Y(_2228_));
 sg13g2_a22oi_1 _5557_ (.Y(_2229_),
    .B1(_2216_),
    .B2(_2228_),
    .A2(_1620_),
    .A1(_2101_));
 sg13g2_a221oi_1 _5558_ (.B2(_2229_),
    .C1(net65),
    .B1(_2226_),
    .A1(_2221_),
    .Y(_0321_),
    .A2(_2211_));
 sg13g2_inv_1 _5559_ (.Y(_2230_),
    .A(\game.sound_mode[2] ));
 sg13g2_nand2_1 _5560_ (.Y(_2231_),
    .A(_2101_),
    .B(_2216_));
 sg13g2_a221oi_1 _5561_ (.B2(_2231_),
    .C1(net65),
    .B1(_2226_),
    .A1(_2230_),
    .Y(_0322_),
    .A2(_2211_));
 sg13g2_nand4_1 _5562_ (.B(_0888_),
    .C(_0901_),
    .A(net76),
    .Y(_2232_),
    .D(_1926_));
 sg13g2_nor2_1 _5563_ (.A(_0013_),
    .B(_2232_),
    .Y(_2233_));
 sg13g2_nor2b_1 _5564_ (.A(_2101_),
    .B_N(_2232_),
    .Y(_2234_));
 sg13g2_o21ai_1 _5565_ (.B1(net66),
    .Y(_0323_),
    .A1(_2233_),
    .A2(_2234_));
 sg13g2_or2_1 _5566_ (.X(_2235_),
    .B(_1855_),
    .A(net117));
 sg13g2_nand3_1 _5567_ (.B(_0853_),
    .C(_0888_),
    .A(net76),
    .Y(_2236_));
 sg13g2_o21ai_1 _5568_ (.B1(_2236_),
    .Y(_2237_),
    .A1(_0853_),
    .A2(_2235_));
 sg13g2_and2_1 _5569_ (.A(_0891_),
    .B(_0913_),
    .X(_2238_));
 sg13g2_nand3_1 _5570_ (.B(_1627_),
    .C(_1624_),
    .A(_1625_),
    .Y(_2239_));
 sg13g2_o21ai_1 _5571_ (.B1(_1626_),
    .Y(_2240_),
    .A1(_1942_),
    .A2(net114));
 sg13g2_a21oi_1 _5572_ (.A1(_1862_),
    .A2(_0881_),
    .Y(_2241_),
    .B1(_1629_));
 sg13g2_o21ai_1 _5573_ (.B1(_2241_),
    .Y(_2242_),
    .A1(_2239_),
    .A2(_2240_));
 sg13g2_nand2_1 _5574_ (.Y(_2243_),
    .A(_1640_),
    .B(_2242_));
 sg13g2_nand3_1 _5575_ (.B(_1632_),
    .C(_2243_),
    .A(_1642_),
    .Y(_2244_));
 sg13g2_and3_1 _5576_ (.X(_2245_),
    .A(_1644_),
    .B(net44),
    .C(_1630_));
 sg13g2_nand2_1 _5577_ (.Y(_2246_),
    .A(_2021_),
    .B(_2084_));
 sg13g2_or3_1 _5578_ (.A(net77),
    .B(_0931_),
    .C(_2246_),
    .X(_2247_));
 sg13g2_nand3b_1 _5579_ (.B(_2231_),
    .C(_2247_),
    .Y(_2248_),
    .A_N(_2043_));
 sg13g2_nand3_1 _5580_ (.B(_0879_),
    .C(_2215_),
    .A(net90),
    .Y(_2249_));
 sg13g2_or3_1 _5581_ (.A(net118),
    .B(_1526_),
    .C(_1921_),
    .X(_2250_));
 sg13g2_a21oi_1 _5582_ (.A1(_2249_),
    .A2(_2250_),
    .Y(_2251_),
    .B1(_0863_));
 sg13g2_nor4_1 _5583_ (.A(_2048_),
    .B(_2245_),
    .C(_2248_),
    .D(_2251_),
    .Y(_2252_));
 sg13g2_nand3_1 _5584_ (.B(_1881_),
    .C(_1875_),
    .A(net79),
    .Y(_2253_));
 sg13g2_a21oi_1 _5585_ (.A1(_2246_),
    .A2(_2253_),
    .Y(_2254_),
    .B1(net77));
 sg13g2_o21ai_1 _5586_ (.B1(_0913_),
    .Y(_2255_),
    .A1(_1883_),
    .A2(_2254_));
 sg13g2_nand4_1 _5587_ (.B(_2244_),
    .C(_2252_),
    .A(_2100_),
    .Y(_2256_),
    .D(_2255_));
 sg13g2_buf_1 _5588_ (.A(_2256_),
    .X(_2257_));
 sg13g2_a21o_1 _5589_ (.A2(_0881_),
    .A1(net81),
    .B1(_2257_),
    .X(_2258_));
 sg13g2_nand2_1 _5590_ (.Y(_2259_),
    .A(_2101_),
    .B(_0911_));
 sg13g2_a221oi_1 _5591_ (.B2(\game.next_state[0] ),
    .C1(_0881_),
    .B1(_2259_),
    .A1(_0911_),
    .Y(_2260_),
    .A2(_1526_));
 sg13g2_nor4_1 _5592_ (.A(net82),
    .B(net47),
    .C(_1855_),
    .D(_1858_),
    .Y(_2261_));
 sg13g2_nor3_1 _5593_ (.A(_1620_),
    .B(_2260_),
    .C(_2261_),
    .Y(_2262_));
 sg13g2_o21ai_1 _5594_ (.B1(net75),
    .Y(_2263_),
    .A1(_2257_),
    .A2(_2262_));
 sg13g2_a221oi_1 _5595_ (.B2(_1617_),
    .C1(_2263_),
    .B1(_2258_),
    .A1(_2237_),
    .Y(_0324_),
    .A2(_2238_));
 sg13g2_nor2_1 _5596_ (.A(net79),
    .B(net77),
    .Y(_2264_));
 sg13g2_nand2_1 _5597_ (.Y(_2265_),
    .A(_0887_),
    .B(net82));
 sg13g2_o21ai_1 _5598_ (.B1(_2265_),
    .Y(_2266_),
    .A1(_0887_),
    .A2(_2029_));
 sg13g2_a21oi_1 _5599_ (.A1(_2264_),
    .A2(_2266_),
    .Y(_2267_),
    .B1(_1860_));
 sg13g2_a21oi_1 _5600_ (.A1(_1858_),
    .A2(_2083_),
    .Y(_2268_),
    .B1(net82));
 sg13g2_mux2_1 _5601_ (.A0(_1926_),
    .A1(_2268_),
    .S(net79),
    .X(_2269_));
 sg13g2_nand2_1 _5602_ (.Y(_2270_),
    .A(_0887_),
    .B(_2269_));
 sg13g2_mux2_1 _5603_ (.A0(_2267_),
    .A1(_2270_),
    .S(_0853_),
    .X(_2271_));
 sg13g2_nand2_1 _5604_ (.Y(_2272_),
    .A(_1871_),
    .B(_1926_));
 sg13g2_nor4_1 _5605_ (.A(net76),
    .B(_0950_),
    .C(_2272_),
    .D(_2195_),
    .Y(_2273_));
 sg13g2_nor4_1 _5606_ (.A(_2641_),
    .B(_2260_),
    .C(_2258_),
    .D(_2273_),
    .Y(_2274_));
 sg13g2_o21ai_1 _5607_ (.B1(_2274_),
    .Y(_2275_),
    .A1(net47),
    .A2(_2271_));
 sg13g2_nand3_1 _5608_ (.B(net81),
    .C(_2257_),
    .A(net75),
    .Y(_2276_));
 sg13g2_nand2_1 _5609_ (.Y(_0325_),
    .A(_2275_),
    .B(_2276_));
 sg13g2_o21ai_1 _5610_ (.B1(_2202_),
    .Y(_2277_),
    .A1(net76),
    .A2(_2272_));
 sg13g2_nand2b_1 _5611_ (.Y(_2278_),
    .B(_2272_),
    .A_N(_1860_));
 sg13g2_inv_1 _5612_ (.Y(_2279_),
    .A(\game.next_state[2] ));
 sg13g2_nand2b_1 _5613_ (.Y(_2280_),
    .B(_1526_),
    .A_N(net90));
 sg13g2_o21ai_1 _5614_ (.B1(_2280_),
    .Y(_2281_),
    .A1(_2101_),
    .A2(_2279_));
 sg13g2_a22oi_1 _5615_ (.Y(_2282_),
    .B1(_2281_),
    .B2(net89),
    .A2(\game.next_state[2] ),
    .A1(net90));
 sg13g2_a21oi_1 _5616_ (.A1(_0913_),
    .A2(_2278_),
    .Y(_2283_),
    .B1(_2282_));
 sg13g2_a21oi_1 _5617_ (.A1(\game.challenge_mode ),
    .A2(_1632_),
    .Y(_2284_),
    .B1(_2283_));
 sg13g2_a21o_1 _5618_ (.A2(_2284_),
    .A1(_2277_),
    .B1(_2257_),
    .X(_2285_));
 sg13g2_nand2_1 _5619_ (.Y(_2286_),
    .A(_1525_),
    .B(_2257_));
 sg13g2_a21oi_1 _5620_ (.A1(_2285_),
    .A2(_2286_),
    .Y(_0326_),
    .B1(net57));
 sg13g2_nand2_1 _5621_ (.Y(_2287_),
    .A(_1524_),
    .B(_2257_));
 sg13g2_or3_1 _5622_ (.A(_2106_),
    .B(_2102_),
    .C(_2257_),
    .X(_2288_));
 sg13g2_a21oi_1 _5623_ (.A1(_2287_),
    .A2(_2288_),
    .Y(_0327_),
    .B1(_1827_));
 sg13g2_o21ai_1 _5624_ (.B1(_0911_),
    .Y(_2289_),
    .A1(_1618_),
    .A2(_1853_));
 sg13g2_nand2_1 _5625_ (.Y(_2290_),
    .A(_0911_),
    .B(_1526_));
 sg13g2_a21oi_1 _5626_ (.A1(_0879_),
    .A2(_2105_),
    .Y(_2291_),
    .B1(_2290_));
 sg13g2_or2_1 _5627_ (.X(_2292_),
    .B(_2291_),
    .A(\game.tune[0] ));
 sg13g2_and3_1 _5628_ (.X(_0328_),
    .A(net95),
    .B(_2289_),
    .C(_2292_));
 sg13g2_o21ai_1 _5629_ (.B1(_2227_),
    .Y(_2293_),
    .A1(net83),
    .A2(_2106_));
 sg13g2_nand2_1 _5630_ (.Y(_2294_),
    .A(_2017_),
    .B(_2293_));
 sg13g2_a22oi_1 _5631_ (.Y(_2295_),
    .B1(_2105_),
    .B2(_2227_),
    .A2(_0911_),
    .A1(_1854_));
 sg13g2_nor2_1 _5632_ (.A(net81),
    .B(_2295_),
    .Y(_2296_));
 sg13g2_nor3_1 _5633_ (.A(_2107_),
    .B(_2294_),
    .C(_2296_),
    .Y(_0329_));
 sg13g2_and2_1 _5634_ (.A(net55),
    .B(_1413_),
    .X(_0330_));
 sg13g2_buf_1 _5635_ (.A(\snd.active_tune[0] ),
    .X(_2297_));
 sg13g2_nand2_1 _5636_ (.Y(_2298_),
    .A(_2220_),
    .B(net113));
 sg13g2_nor2_1 _5637_ (.A(\game.sound_mode[2] ),
    .B(_2298_),
    .Y(_2299_));
 sg13g2_a21oi_2 _5638_ (.B1(_2299_),
    .Y(_2300_),
    .A2(_2298_),
    .A1(_0038_));
 sg13g2_nor2b_1 _5639_ (.A(net112),
    .B_N(net113),
    .Y(_2301_));
 sg13g2_a22oi_1 _5640_ (.Y(_2302_),
    .B1(_2300_),
    .B2(_2301_),
    .A2(net111),
    .A1(net112));
 sg13g2_or2_1 _5641_ (.X(_2303_),
    .B(_2302_),
    .A(_2214_));
 sg13g2_inv_1 _5642_ (.Y(_2304_),
    .A(_2214_));
 sg13g2_nand2b_1 _5643_ (.Y(_2305_),
    .B(net111),
    .A_N(net112));
 sg13g2_a21o_1 _5644_ (.A2(_2300_),
    .A1(_2304_),
    .B1(_2305_),
    .X(_2306_));
 sg13g2_a21oi_1 _5645_ (.A1(_2303_),
    .A2(_2306_),
    .Y(_0331_),
    .B1(net57));
 sg13g2_nor2_1 _5646_ (.A(_2213_),
    .B(_2214_),
    .Y(_2307_));
 sg13g2_nand2b_1 _5647_ (.Y(_2308_),
    .B(net113),
    .A_N(\game.sound_mode[2] ));
 sg13g2_nand2b_1 _5648_ (.Y(_2309_),
    .B(_0038_),
    .A_N(net113));
 sg13g2_nand4_1 _5649_ (.B(_2307_),
    .C(_2308_),
    .A(_2220_),
    .Y(_2310_),
    .D(_2309_));
 sg13g2_buf_2 _5650_ (.A(\snd.active_tune[1] ),
    .X(_2311_));
 sg13g2_inv_1 _5651_ (.Y(_2312_),
    .A(_2311_));
 sg13g2_a21oi_1 _5652_ (.A1(_2213_),
    .A2(_2214_),
    .Y(_2313_),
    .B1(_2312_));
 sg13g2_nand2_1 _5653_ (.Y(_2314_),
    .A(_2307_),
    .B(_2300_));
 sg13g2_nand2_1 _5654_ (.Y(_2315_),
    .A(_2313_),
    .B(_2314_));
 sg13g2_a21oi_1 _5655_ (.A1(_2310_),
    .A2(_2315_),
    .Y(_0332_),
    .B1(net57));
 sg13g2_buf_1 _5656_ (.A(\snd.tune_pos[0] ),
    .X(_2316_));
 sg13g2_buf_2 _5657_ (.A(\snd.tune_pos[2] ),
    .X(_2317_));
 sg13g2_nor2_1 _5658_ (.A(\snd.tune_pos[1] ),
    .B(_2317_),
    .Y(_2318_));
 sg13g2_nand2_1 _5659_ (.Y(_2319_),
    .A(net110),
    .B(_2318_));
 sg13g2_a21oi_1 _5660_ (.A1(net111),
    .A2(_2319_),
    .Y(_2320_),
    .B1(_2311_));
 sg13g2_buf_1 _5661_ (.A(\snd.tune_pos[1] ),
    .X(_2321_));
 sg13g2_buf_2 _5662_ (.A(_0039_),
    .X(_2322_));
 sg13g2_xor2_1 _5663_ (.B(_2322_),
    .A(net109),
    .X(_2323_));
 sg13g2_nor3_1 _5664_ (.A(net111),
    .B(net110),
    .C(_2323_),
    .Y(_2324_));
 sg13g2_nor3_1 _5665_ (.A(_2311_),
    .B(net111),
    .C(_2319_),
    .Y(_2325_));
 sg13g2_buf_1 _5666_ (.A(\snd.tune_counter[2] ),
    .X(_2326_));
 sg13g2_buf_1 _5667_ (.A(\snd.tune_counter[5] ),
    .X(_2327_));
 sg13g2_buf_1 _5668_ (.A(\snd.tune_counter[1] ),
    .X(_2328_));
 sg13g2_buf_1 _5669_ (.A(\snd.tune_counter[4] ),
    .X(_2329_));
 sg13g2_nor2_1 _5670_ (.A(_2328_),
    .B(_2329_),
    .Y(_2330_));
 sg13g2_buf_2 _5671_ (.A(\snd.tune_counter[0] ),
    .X(_2331_));
 sg13g2_buf_1 _5672_ (.A(\snd.tune_counter[3] ),
    .X(_2332_));
 sg13g2_nor3_1 _5673_ (.A(_2331_),
    .B(_2332_),
    .C(_0037_),
    .Y(_2333_));
 sg13g2_nand4_1 _5674_ (.B(_2327_),
    .C(_2330_),
    .A(_2326_),
    .Y(_2334_),
    .D(_2333_));
 sg13g2_nor2b_1 _5675_ (.A(_2214_),
    .B_N(net112),
    .Y(_2335_));
 sg13g2_buf_2 _5676_ (.A(_2335_),
    .X(_2336_));
 sg13g2_and2_1 _5677_ (.A(_2334_),
    .B(_2336_),
    .X(_2337_));
 sg13g2_buf_1 _5678_ (.A(_2337_),
    .X(_2338_));
 sg13g2_nor4_1 _5679_ (.A(_2331_),
    .B(_2332_),
    .C(_2326_),
    .D(\snd.tune_counter[6] ),
    .Y(_2339_));
 sg13g2_nand3b_1 _5680_ (.B(_2330_),
    .C(_2339_),
    .Y(_2340_),
    .A_N(_2327_));
 sg13g2_buf_1 _5681_ (.A(_2340_),
    .X(_2341_));
 sg13g2_nand2_1 _5682_ (.Y(_2342_),
    .A(_2317_),
    .B(_2322_));
 sg13g2_inv_1 _5683_ (.Y(_2343_),
    .A(net110));
 sg13g2_nor2_1 _5684_ (.A(_2343_),
    .B(_2317_),
    .Y(_2344_));
 sg13g2_a21oi_1 _5685_ (.A1(_2343_),
    .A2(_2322_),
    .Y(_2345_),
    .B1(_2344_));
 sg13g2_nand2_1 _5686_ (.Y(_2346_),
    .A(net109),
    .B(_2345_));
 sg13g2_o21ai_1 _5687_ (.B1(_2346_),
    .Y(_2347_),
    .A1(net109),
    .A2(_2342_));
 sg13g2_nor3_1 _5688_ (.A(net115),
    .B(_2312_),
    .C(\snd.active_tune[0] ),
    .Y(_2348_));
 sg13g2_nor2_1 _5689_ (.A(_1660_),
    .B(_2318_),
    .Y(_2349_));
 sg13g2_a22oi_1 _5690_ (.Y(_2350_),
    .B1(_2349_),
    .B2(_2312_),
    .A2(_2348_),
    .A1(_2347_));
 sg13g2_and2_1 _5691_ (.A(_2311_),
    .B(\snd.active_tune[0] ),
    .X(_2351_));
 sg13g2_nand2_1 _5692_ (.Y(_2352_),
    .A(_2343_),
    .B(_2318_));
 sg13g2_a21oi_1 _5693_ (.A1(_2351_),
    .A2(_2352_),
    .Y(_2353_),
    .B1(_2341_));
 sg13g2_or2_1 _5694_ (.X(_2354_),
    .B(_2353_),
    .A(net115));
 sg13g2_o21ai_1 _5695_ (.B1(_2354_),
    .Y(_2355_),
    .A1(_2341_),
    .A2(_2350_));
 sg13g2_nor2_2 _5696_ (.A(net112),
    .B(_2304_),
    .Y(_2356_));
 sg13g2_a21oi_1 _5697_ (.A1(_2338_),
    .A2(_2355_),
    .Y(_2357_),
    .B1(_2356_));
 sg13g2_inv_1 _5698_ (.Y(_2358_),
    .A(_2338_));
 sg13g2_nor2_1 _5699_ (.A(net115),
    .B(_2358_),
    .Y(_2359_));
 sg13g2_and2_1 _5700_ (.A(_2357_),
    .B(_2359_),
    .X(_2360_));
 sg13g2_nor2b_1 _5701_ (.A(_2325_),
    .B_N(_2360_),
    .Y(_2361_));
 sg13g2_o21ai_1 _5702_ (.B1(_2361_),
    .Y(_2362_),
    .A1(_2320_),
    .A2(_2324_));
 sg13g2_nand2_1 _5703_ (.Y(_2363_),
    .A(net115),
    .B(_2336_));
 sg13g2_nand2_1 _5704_ (.Y(_2364_),
    .A(_2357_),
    .B(_2363_));
 sg13g2_buf_2 _5705_ (.A(_2364_),
    .X(_2365_));
 sg13g2_o21ai_1 _5706_ (.B1(_2307_),
    .Y(_2366_),
    .A1(_2220_),
    .A2(_2309_));
 sg13g2_buf_1 _5707_ (.A(_2366_),
    .X(_2367_));
 sg13g2_nor2_2 _5708_ (.A(_2221_),
    .B(\game.sound_mode[2] ),
    .Y(_2368_));
 sg13g2_a21o_1 _5709_ (.A2(_0038_),
    .A1(_2221_),
    .B1(_2368_),
    .X(_2369_));
 sg13g2_buf_1 _5710_ (.A(_2369_),
    .X(_2370_));
 sg13g2_a22oi_1 _5711_ (.Y(_2371_),
    .B1(_2370_),
    .B2(_1659_),
    .A2(_2368_),
    .A1(net12));
 sg13g2_inv_1 _5712_ (.Y(_2372_),
    .A(_2371_));
 sg13g2_nor2_2 _5713_ (.A(_2221_),
    .B(_2309_),
    .Y(_2373_));
 sg13g2_a22oi_1 _5714_ (.Y(_2374_),
    .B1(_2373_),
    .B2(net12),
    .A2(_2372_),
    .A1(net113));
 sg13g2_nor2_1 _5715_ (.A(_2367_),
    .B(_2374_),
    .Y(_2375_));
 sg13g2_a21oi_1 _5716_ (.A1(\snd.chord[0][0] ),
    .A2(_2365_),
    .Y(_2376_),
    .B1(_2375_));
 sg13g2_a21oi_1 _5717_ (.A1(_2362_),
    .A2(_2376_),
    .Y(_0333_),
    .B1(net57));
 sg13g2_nand2_1 _5718_ (.Y(_2377_),
    .A(_2316_),
    .B(_2321_));
 sg13g2_or3_1 _5719_ (.A(_2316_),
    .B(_2321_),
    .C(_2322_),
    .X(_2378_));
 sg13g2_o21ai_1 _5720_ (.B1(_2378_),
    .Y(_2379_),
    .A1(_2317_),
    .A2(_2377_));
 sg13g2_nor2b_1 _5721_ (.A(net111),
    .B_N(_2379_),
    .Y(_2380_));
 sg13g2_o21ai_1 _5722_ (.B1(_2338_),
    .Y(_2381_),
    .A1(_2312_),
    .A2(_2380_));
 sg13g2_nand2_1 _5723_ (.Y(_2382_),
    .A(\snd.chord[0][1] ),
    .B(_2365_));
 sg13g2_o21ai_1 _5724_ (.B1(_2382_),
    .Y(_2383_),
    .A1(_2365_),
    .A2(_2381_));
 sg13g2_o21ai_1 _5725_ (.B1(_0971_),
    .Y(_2384_),
    .A1(_2375_),
    .A2(_2383_));
 sg13g2_inv_1 _5726_ (.Y(_0334_),
    .A(_2384_));
 sg13g2_xnor2_1 _5727_ (.Y(_2385_),
    .A(net110),
    .B(_2317_));
 sg13g2_nor3_1 _5728_ (.A(net111),
    .B(net109),
    .C(_2385_),
    .Y(_2386_));
 sg13g2_o21ai_1 _5729_ (.B1(_2361_),
    .Y(_2387_),
    .A1(_2320_),
    .A2(_2386_));
 sg13g2_a21oi_1 _5730_ (.A1(\snd.chord[0][2] ),
    .A2(_2365_),
    .Y(_2388_),
    .B1(_2375_));
 sg13g2_buf_1 _5731_ (.A(net108),
    .X(_2389_));
 sg13g2_a21oi_1 _5732_ (.A1(_2387_),
    .A2(_2388_),
    .Y(_0335_),
    .B1(net52));
 sg13g2_buf_1 _5733_ (.A(\snd.chord[0][3] ),
    .X(_2390_));
 sg13g2_nand3_1 _5734_ (.B(net109),
    .C(_2322_),
    .A(_2311_),
    .Y(_2391_));
 sg13g2_nor3_1 _5735_ (.A(_2297_),
    .B(net110),
    .C(_2391_),
    .Y(_2392_));
 sg13g2_a22oi_1 _5736_ (.Y(_2393_),
    .B1(_2392_),
    .B2(_2360_),
    .A2(_2365_),
    .A1(_2390_));
 sg13g2_nor2_1 _5737_ (.A(net53),
    .B(_2393_),
    .Y(_0336_));
 sg13g2_xor2_1 _5738_ (.B(_2317_),
    .A(_2311_),
    .X(_2394_));
 sg13g2_nor4_1 _5739_ (.A(net111),
    .B(_2343_),
    .C(net109),
    .D(_2394_),
    .Y(_2395_));
 sg13g2_a221oi_1 _5740_ (.B2(_2360_),
    .C1(_2375_),
    .B1(_2395_),
    .A1(\snd.chord[0][4] ),
    .Y(_2396_),
    .A2(_2365_));
 sg13g2_nor2_1 _5741_ (.A(net53),
    .B(_2396_),
    .Y(_0337_));
 sg13g2_buf_1 _5742_ (.A(\snd.chord[0][5] ),
    .X(_2397_));
 sg13g2_buf_1 _5743_ (.A(_2397_),
    .X(_2398_));
 sg13g2_a21oi_1 _5744_ (.A1(net74),
    .A2(_2365_),
    .Y(_2399_),
    .B1(_2361_));
 sg13g2_nor2_1 _5745_ (.A(net53),
    .B(_2399_),
    .Y(_0338_));
 sg13g2_o21ai_1 _5746_ (.B1(_2354_),
    .Y(_2400_),
    .A1(_2341_),
    .A2(_2351_));
 sg13g2_a21oi_1 _5747_ (.A1(_2338_),
    .A2(_2400_),
    .Y(_2401_),
    .B1(_2356_));
 sg13g2_nand2_1 _5748_ (.Y(_2402_),
    .A(_2363_),
    .B(_2401_));
 sg13g2_a22oi_1 _5749_ (.Y(_2403_),
    .B1(_2402_),
    .B2(\snd.chord[1][0] ),
    .A2(_2401_),
    .A1(_2359_));
 sg13g2_nor2_1 _5750_ (.A(net53),
    .B(_2403_),
    .Y(_0339_));
 sg13g2_a22oi_1 _5751_ (.Y(_2404_),
    .B1(_2370_),
    .B2(_1664_),
    .A2(_2368_),
    .A1(net13));
 sg13g2_inv_1 _5752_ (.Y(_2405_),
    .A(_2404_));
 sg13g2_a22oi_1 _5753_ (.Y(_2406_),
    .B1(_2405_),
    .B2(net113),
    .A2(_2373_),
    .A1(net13));
 sg13g2_o21ai_1 _5754_ (.B1(_2358_),
    .Y(_2407_),
    .A1(_2367_),
    .A2(_2406_));
 sg13g2_mux2_1 _5755_ (.A0(_2407_),
    .A1(\snd.chord[1][5] ),
    .S(_2402_),
    .X(_2408_));
 sg13g2_and2_1 _5756_ (.A(net55),
    .B(_2408_),
    .X(_0340_));
 sg13g2_buf_2 _5757_ (.A(\snd.chord[2][2] ),
    .X(_2409_));
 sg13g2_o21ai_1 _5758_ (.B1(_2336_),
    .Y(_2410_),
    .A1(net115),
    .A2(_2334_));
 sg13g2_nand2b_1 _5759_ (.Y(_2411_),
    .B(_2410_),
    .A_N(_2356_));
 sg13g2_a22oi_1 _5760_ (.Y(_2412_),
    .B1(_2370_),
    .B2(_1673_),
    .A2(_2368_),
    .A1(net14));
 sg13g2_inv_1 _5761_ (.Y(_2413_),
    .A(_2412_));
 sg13g2_a22oi_1 _5762_ (.Y(_2414_),
    .B1(_2413_),
    .B2(net113),
    .A2(_2373_),
    .A1(net14));
 sg13g2_nor2_1 _5763_ (.A(_2367_),
    .B(_2414_),
    .Y(_2415_));
 sg13g2_a21oi_1 _5764_ (.A1(_2409_),
    .A2(_2411_),
    .Y(_2416_),
    .B1(_2415_));
 sg13g2_nor2_1 _5765_ (.A(net53),
    .B(_2416_),
    .Y(_0341_));
 sg13g2_buf_1 _5766_ (.A(\snd.chord[3][0] ),
    .X(_2417_));
 sg13g2_a22oi_1 _5767_ (.Y(_2418_),
    .B1(_2370_),
    .B2(_1678_),
    .A2(_2368_),
    .A1(net15));
 sg13g2_inv_1 _5768_ (.Y(_2419_),
    .A(_2418_));
 sg13g2_a22oi_1 _5769_ (.Y(_2420_),
    .B1(_2419_),
    .B2(net113),
    .A2(_2373_),
    .A1(net15));
 sg13g2_nor2_1 _5770_ (.A(_2367_),
    .B(_2420_),
    .Y(_2421_));
 sg13g2_a21oi_1 _5771_ (.A1(_2417_),
    .A2(_2411_),
    .Y(_2422_),
    .B1(_2421_));
 sg13g2_nor2_1 _5772_ (.A(net53),
    .B(_2422_),
    .Y(_0342_));
 sg13g2_buf_1 _5773_ (.A(_1568_),
    .X(_2423_));
 sg13g2_a21oi_1 _5774_ (.A1(_1545_),
    .A2(net20),
    .Y(_0343_),
    .B1(net52));
 sg13g2_buf_1 _5775_ (.A(\snd.note_sel[1] ),
    .X(_2424_));
 sg13g2_nor2_2 _5776_ (.A(\snd.chord[1][5] ),
    .B(\snd.chord[1][0] ),
    .Y(_2425_));
 sg13g2_buf_2 _5777_ (.A(\snd.note_sel[0] ),
    .X(_2426_));
 sg13g2_nand3b_1 _5778_ (.B(_2426_),
    .C(_2417_),
    .Y(_2427_),
    .A_N(_2409_));
 sg13g2_nor2_1 _5779_ (.A(_2390_),
    .B(\snd.chord[0][2] ),
    .Y(_2428_));
 sg13g2_nor4_2 _5780_ (.A(\snd.chord[0][1] ),
    .B(\snd.chord[0][0] ),
    .C(_2397_),
    .Y(_2429_),
    .D(\snd.chord[0][4] ));
 sg13g2_nand2_1 _5781_ (.Y(_2430_),
    .A(_2428_),
    .B(_2429_));
 sg13g2_a21oi_1 _5782_ (.A1(_2425_),
    .A2(_2427_),
    .Y(_2431_),
    .B1(_2430_));
 sg13g2_nor2_1 _5783_ (.A(_2426_),
    .B(_0060_),
    .Y(_2432_));
 sg13g2_nor2_1 _5784_ (.A(_2431_),
    .B(_2432_),
    .Y(_2433_));
 sg13g2_nand3b_1 _5785_ (.B(_2428_),
    .C(_2429_),
    .Y(_2434_),
    .A_N(_2425_));
 sg13g2_nand2b_1 _5786_ (.Y(_2435_),
    .B(_2426_),
    .A_N(_0060_));
 sg13g2_a21oi_1 _5787_ (.A1(_2434_),
    .A2(_2435_),
    .Y(_2436_),
    .B1(_2409_));
 sg13g2_nand2b_1 _5788_ (.Y(_2437_),
    .B(_2417_),
    .A_N(_2409_));
 sg13g2_a21oi_1 _5789_ (.A1(_2425_),
    .A2(_2437_),
    .Y(_2438_),
    .B1(_2426_));
 sg13g2_nor3_1 _5790_ (.A(_2424_),
    .B(_2436_),
    .C(_2438_),
    .Y(_2439_));
 sg13g2_a21oi_1 _5791_ (.A1(_2424_),
    .A2(_2433_),
    .Y(_2440_),
    .B1(_2439_));
 sg13g2_buf_2 _5792_ (.A(_2440_),
    .X(_2441_));
 sg13g2_nor2b_1 _5793_ (.A(net87),
    .B_N(\snd.next_note_sel[0] ),
    .Y(_2442_));
 sg13g2_a21oi_1 _5794_ (.A1(net59),
    .A2(_2441_),
    .Y(_2443_),
    .B1(_2442_));
 sg13g2_nor2_1 _5795_ (.A(_2190_),
    .B(_2443_),
    .Y(_0352_));
 sg13g2_nor2b_1 _5796_ (.A(_2426_),
    .B_N(_2424_),
    .Y(_2444_));
 sg13g2_nand2_1 _5797_ (.Y(_2445_),
    .A(_2409_),
    .B(_2425_));
 sg13g2_o21ai_1 _5798_ (.B1(_0060_),
    .Y(_2446_),
    .A1(_2430_),
    .A2(_2445_));
 sg13g2_or2_1 _5799_ (.X(_2447_),
    .B(_2409_),
    .A(_2417_));
 sg13g2_nor2_1 _5800_ (.A(_2426_),
    .B(_2425_),
    .Y(_2448_));
 sg13g2_nand4_1 _5801_ (.B(_2425_),
    .C(_2428_),
    .A(_2426_),
    .Y(_2449_),
    .D(_2429_));
 sg13g2_o21ai_1 _5802_ (.B1(_2449_),
    .Y(_2450_),
    .A1(_2424_),
    .A2(_2448_));
 sg13g2_a22oi_1 _5803_ (.Y(_2451_),
    .B1(_2447_),
    .B2(_2450_),
    .A2(_2446_),
    .A1(_2444_));
 sg13g2_buf_2 _5804_ (.A(_2451_),
    .X(_2452_));
 sg13g2_nand2_1 _5805_ (.Y(_2453_),
    .A(net87),
    .B(_2452_));
 sg13g2_o21ai_1 _5806_ (.B1(_2453_),
    .Y(_2454_),
    .A1(net62),
    .A2(\snd.next_note_sel[1] ));
 sg13g2_nor2_1 _5807_ (.A(_2190_),
    .B(_2454_),
    .Y(_0353_));
 sg13g2_mux4_1 _5808_ (.S0(_2452_),
    .A0(_2409_),
    .A1(_2397_),
    .A2(_2417_),
    .A3(\snd.chord[1][5] ),
    .S1(_2441_),
    .X(_2455_));
 sg13g2_nor2b_1 _5809_ (.A(_2441_),
    .B_N(_2452_),
    .Y(_2456_));
 sg13g2_buf_1 _5810_ (.A(_2456_),
    .X(_2457_));
 sg13g2_and2_1 _5811_ (.A(\snd.chord[0][4] ),
    .B(_2457_),
    .X(_2458_));
 sg13g2_buf_2 _5812_ (.A(_2458_),
    .X(_2459_));
 sg13g2_o21ai_1 _5813_ (.B1(net87),
    .Y(_2460_),
    .A1(_2455_),
    .A2(_2459_));
 sg13g2_nor2b_1 _5814_ (.A(_2452_),
    .B_N(_2417_),
    .Y(_2461_));
 sg13g2_a22oi_1 _5815_ (.Y(_2462_),
    .B1(_2457_),
    .B2(\snd.chord[0][1] ),
    .A2(_2461_),
    .A1(_2441_));
 sg13g2_buf_2 _5816_ (.A(_2462_),
    .X(_2463_));
 sg13g2_inv_1 _5817_ (.Y(_2464_),
    .A(_2463_));
 sg13g2_nand3_1 _5818_ (.B(_2457_),
    .C(_2464_),
    .A(_0057_),
    .Y(_2465_));
 sg13g2_buf_1 _5819_ (.A(_2465_),
    .X(_2466_));
 sg13g2_inv_1 _5820_ (.Y(_2467_),
    .A(_2466_));
 sg13g2_nand2b_1 _5821_ (.Y(_2468_),
    .B(\snd.chord[0][2] ),
    .A_N(_2390_));
 sg13g2_nor2_1 _5822_ (.A(_2409_),
    .B(_2452_),
    .Y(_2469_));
 sg13g2_a21oi_1 _5823_ (.A1(_2452_),
    .A2(_2468_),
    .Y(_2470_),
    .B1(_2469_));
 sg13g2_a21o_1 _5824_ (.A2(_2452_),
    .A1(\snd.chord[1][0] ),
    .B1(_2461_),
    .X(_2471_));
 sg13g2_mux2_1 _5825_ (.A0(_2470_),
    .A1(_2471_),
    .S(_2441_),
    .X(_2472_));
 sg13g2_buf_2 _5826_ (.A(_2472_),
    .X(_2473_));
 sg13g2_nand3b_1 _5827_ (.B(_2457_),
    .C(_2390_),
    .Y(_2474_),
    .A_N(\snd.chord[0][2] ));
 sg13g2_buf_1 _5828_ (.A(_2474_),
    .X(_2475_));
 sg13g2_inv_1 _5829_ (.Y(_2476_),
    .A(_2475_));
 sg13g2_inv_1 _5830_ (.Y(_2477_),
    .A(_0057_));
 sg13g2_a22oi_1 _5831_ (.Y(_2478_),
    .B1(_2471_),
    .B2(_2441_),
    .A2(_2457_),
    .A1(_2477_));
 sg13g2_buf_2 _5832_ (.A(_2478_),
    .X(_2479_));
 sg13g2_a21oi_1 _5833_ (.A1(_2428_),
    .A2(_2452_),
    .Y(_2480_),
    .B1(_2469_));
 sg13g2_mux2_1 _5834_ (.A0(_2480_),
    .A1(_2471_),
    .S(_2441_),
    .X(_2481_));
 sg13g2_buf_2 _5835_ (.A(_2481_),
    .X(_2482_));
 sg13g2_a21oi_1 _5836_ (.A1(_2463_),
    .A2(_2479_),
    .Y(_2483_),
    .B1(_2482_));
 sg13g2_nor2_1 _5837_ (.A(_2476_),
    .B(_2483_),
    .Y(_2484_));
 sg13g2_nor3_1 _5838_ (.A(_2467_),
    .B(_2473_),
    .C(_2484_),
    .Y(_2485_));
 sg13g2_nor2b_1 _5839_ (.A(_2485_),
    .B_N(net74),
    .Y(_2486_));
 sg13g2_nand2_1 _5840_ (.Y(_2487_),
    .A(\snd.chord[0][4] ),
    .B(_2457_));
 sg13g2_and2_1 _5841_ (.A(_2455_),
    .B(_2487_),
    .X(_2488_));
 sg13g2_buf_1 _5842_ (.A(_2488_),
    .X(_2489_));
 sg13g2_nand2_1 _5843_ (.Y(_2490_),
    .A(_2463_),
    .B(_2479_));
 sg13g2_nand2_1 _5844_ (.Y(_2491_),
    .A(_2482_),
    .B(_2490_));
 sg13g2_o21ai_1 _5845_ (.B1(_2491_),
    .Y(_2492_),
    .A1(_2476_),
    .A2(_2490_));
 sg13g2_o21ai_1 _5846_ (.B1(_2466_),
    .Y(_2493_),
    .A1(_2464_),
    .A2(_2479_));
 sg13g2_nand2_1 _5847_ (.Y(_2494_),
    .A(_2482_),
    .B(_2493_));
 sg13g2_o21ai_1 _5848_ (.B1(_2494_),
    .Y(_2495_),
    .A1(_2473_),
    .A2(_2483_));
 sg13g2_nand2_1 _5849_ (.Y(_2496_),
    .A(_2390_),
    .B(_2477_));
 sg13g2_nor2_2 _5850_ (.A(_2397_),
    .B(_2487_),
    .Y(_2497_));
 sg13g2_o21ai_1 _5851_ (.B1(_2497_),
    .Y(_2498_),
    .A1(_2463_),
    .A2(_2496_));
 sg13g2_a21oi_1 _5852_ (.A1(_2475_),
    .A2(_2495_),
    .Y(_2499_),
    .B1(_2498_));
 sg13g2_a221oi_1 _5853_ (.B2(_2492_),
    .C1(_2499_),
    .B1(_2489_),
    .A1(_2459_),
    .Y(_2500_),
    .A2(_2486_));
 sg13g2_nand2_1 _5854_ (.Y(_2501_),
    .A(net88),
    .B(\snd.next_note_timing[0] ));
 sg13g2_o21ai_1 _5855_ (.B1(_2501_),
    .Y(_2502_),
    .A1(_2460_),
    .A2(_2500_));
 sg13g2_and2_1 _5856_ (.A(net55),
    .B(_2502_),
    .X(_0354_));
 sg13g2_o21ai_1 _5857_ (.B1(_2463_),
    .Y(_2503_),
    .A1(_2397_),
    .A2(_2479_));
 sg13g2_nor2b_1 _5858_ (.A(_2482_),
    .B_N(_2503_),
    .Y(_2504_));
 sg13g2_a21oi_1 _5859_ (.A1(_2463_),
    .A2(_2482_),
    .Y(_2505_),
    .B1(_2479_));
 sg13g2_nand2b_1 _5860_ (.Y(_2506_),
    .B(net74),
    .A_N(_2505_));
 sg13g2_a21oi_1 _5861_ (.A1(_2490_),
    .A2(_2506_),
    .Y(_2507_),
    .B1(_2475_));
 sg13g2_nor3_1 _5862_ (.A(_2487_),
    .B(_2504_),
    .C(_2507_),
    .Y(_2508_));
 sg13g2_nor2b_1 _5863_ (.A(_2485_),
    .B_N(_2489_),
    .Y(_2509_));
 sg13g2_nor2_1 _5864_ (.A(_2508_),
    .B(_2509_),
    .Y(_2510_));
 sg13g2_o21ai_1 _5865_ (.B1(_2017_),
    .Y(_2511_),
    .A1(net87),
    .A2(\snd.next_note_timing[1] ));
 sg13g2_a21oi_1 _5866_ (.A1(net59),
    .A2(_2510_),
    .Y(_0355_),
    .B1(_2511_));
 sg13g2_nor2_1 _5867_ (.A(_2475_),
    .B(_2505_),
    .Y(_2512_));
 sg13g2_nor2_1 _5868_ (.A(_2463_),
    .B(_2482_),
    .Y(_2513_));
 sg13g2_nor2_1 _5869_ (.A(_2512_),
    .B(_2513_),
    .Y(_2514_));
 sg13g2_nand2_1 _5870_ (.Y(_2515_),
    .A(_2475_),
    .B(_2482_));
 sg13g2_mux2_1 _5871_ (.A0(_2473_),
    .A1(_2466_),
    .S(_2515_),
    .X(_2516_));
 sg13g2_inv_1 _5872_ (.Y(_2517_),
    .A(_2516_));
 sg13g2_nand2b_1 _5873_ (.Y(_2518_),
    .B(_2473_),
    .A_N(_2479_));
 sg13g2_o21ai_1 _5874_ (.B1(_2518_),
    .Y(_2519_),
    .A1(_2473_),
    .A2(_2490_));
 sg13g2_o21ai_1 _5875_ (.B1(_2398_),
    .Y(_2520_),
    .A1(_2517_),
    .A2(_2519_));
 sg13g2_o21ai_1 _5876_ (.B1(_2520_),
    .Y(_2521_),
    .A1(net74),
    .A2(_2485_));
 sg13g2_a22oi_1 _5877_ (.Y(_2522_),
    .B1(_2521_),
    .B2(_2459_),
    .A2(_2514_),
    .A1(_2489_));
 sg13g2_nand2_1 _5878_ (.Y(_2523_),
    .A(net88),
    .B(\snd.next_note_timing[2] ));
 sg13g2_o21ai_1 _5879_ (.B1(_2523_),
    .Y(_2524_),
    .A1(_2460_),
    .A2(_2522_));
 sg13g2_and2_1 _5880_ (.A(net55),
    .B(_2524_),
    .X(_0356_));
 sg13g2_nor2_1 _5881_ (.A(net62),
    .B(\snd.next_note_timing[3] ),
    .Y(_2525_));
 sg13g2_nor2_1 _5882_ (.A(_2517_),
    .B(_2519_),
    .Y(_2526_));
 sg13g2_inv_1 _5883_ (.Y(_2527_),
    .A(_2526_));
 sg13g2_nand2_1 _5884_ (.Y(_2528_),
    .A(_2463_),
    .B(_2482_));
 sg13g2_o21ai_1 _5885_ (.B1(_2466_),
    .Y(_2529_),
    .A1(_2479_),
    .A2(_2528_));
 sg13g2_a22oi_1 _5886_ (.Y(_2530_),
    .B1(_2529_),
    .B2(_2473_),
    .A2(_2515_),
    .A1(_2464_));
 sg13g2_mux2_1 _5887_ (.A0(_2514_),
    .A1(_2530_),
    .S(net74),
    .X(_2531_));
 sg13g2_a221oi_1 _5888_ (.B2(_2459_),
    .C1(net58),
    .B1(_2531_),
    .A1(_2489_),
    .Y(_2532_),
    .A2(_2527_));
 sg13g2_nor3_1 _5889_ (.A(net92),
    .B(_2525_),
    .C(_2532_),
    .Y(_0357_));
 sg13g2_nor2_1 _5890_ (.A(net62),
    .B(\snd.next_note_timing[4] ),
    .Y(_2533_));
 sg13g2_nand2b_1 _5891_ (.Y(_2534_),
    .B(_2464_),
    .A_N(_2518_));
 sg13g2_and2_1 _5892_ (.A(_2475_),
    .B(_2534_),
    .X(_2535_));
 sg13g2_buf_1 _5893_ (.A(_2535_),
    .X(_2536_));
 sg13g2_nand2_1 _5894_ (.Y(_2537_),
    .A(_2473_),
    .B(_2536_));
 sg13g2_nand2_1 _5895_ (.Y(_2538_),
    .A(net74),
    .B(_2537_));
 sg13g2_o21ai_1 _5896_ (.B1(_2538_),
    .Y(_2539_),
    .A1(net74),
    .A2(_2526_));
 sg13g2_a221oi_1 _5897_ (.B2(_2459_),
    .C1(net88),
    .B1(_2539_),
    .A1(_2489_),
    .Y(_2540_),
    .A2(_2530_));
 sg13g2_nor3_1 _5898_ (.A(_1417_),
    .B(_2533_),
    .C(_2540_),
    .Y(_0358_));
 sg13g2_buf_1 _5899_ (.A(_2642_),
    .X(_2541_));
 sg13g2_o21ai_1 _5900_ (.B1(_2536_),
    .Y(_2542_),
    .A1(_2459_),
    .A2(_2473_));
 sg13g2_a22oi_1 _5901_ (.Y(_2543_),
    .B1(_2542_),
    .B2(_2455_),
    .A2(_2530_),
    .A1(_2497_));
 sg13g2_nor2_1 _5902_ (.A(_2460_),
    .B(_2543_),
    .Y(_2544_));
 sg13g2_a21oi_1 _5903_ (.A1(net61),
    .A2(\snd.next_note_timing[5] ),
    .Y(_2545_),
    .B1(_2544_));
 sg13g2_nor2_1 _5904_ (.A(_2541_),
    .B(_2545_),
    .Y(_0359_));
 sg13g2_nand2_1 _5905_ (.Y(_2546_),
    .A(_2475_),
    .B(_2534_));
 sg13g2_a21oi_1 _5906_ (.A1(_2455_),
    .A2(_2546_),
    .Y(_2547_),
    .B1(_2459_));
 sg13g2_nand3_1 _5907_ (.B(_2459_),
    .C(_2546_),
    .A(net74),
    .Y(_2548_));
 sg13g2_o21ai_1 _5908_ (.B1(_2548_),
    .Y(_2549_),
    .A1(_2398_),
    .A2(_2537_));
 sg13g2_or3_1 _5909_ (.A(net88),
    .B(_2547_),
    .C(_2549_),
    .X(_2550_));
 sg13g2_nand2_1 _5910_ (.Y(_2551_),
    .A(net61),
    .B(\snd.next_note_timing[6] ));
 sg13g2_a21oi_1 _5911_ (.A1(_2550_),
    .A2(_2551_),
    .Y(_0360_),
    .B1(net52));
 sg13g2_nor2_1 _5912_ (.A(net87),
    .B(\snd.next_note_timing[7] ),
    .Y(_2552_));
 sg13g2_mux2_1 _5913_ (.A0(_2497_),
    .A1(_2489_),
    .S(_2536_),
    .X(_2553_));
 sg13g2_nor2_1 _5914_ (.A(net58),
    .B(_2553_),
    .Y(_2554_));
 sg13g2_nor3_1 _5915_ (.A(_1417_),
    .B(_2552_),
    .C(_2554_),
    .Y(_0361_));
 sg13g2_nand2_1 _5916_ (.Y(_2555_),
    .A(net61),
    .B(\snd.next_note_timing[8] ));
 sg13g2_nand3_1 _5917_ (.B(_2497_),
    .C(_2536_),
    .A(net87),
    .Y(_2556_));
 sg13g2_a21oi_1 _5918_ (.A1(_2555_),
    .A2(_2556_),
    .Y(_0362_),
    .B1(net52));
 sg13g2_nand2_1 _5919_ (.Y(_2557_),
    .A(_2426_),
    .B(net20));
 sg13g2_nand2b_1 _5920_ (.Y(_2558_),
    .B(\snd.next_note_sel[0] ),
    .A_N(net20));
 sg13g2_a21oi_1 _5921_ (.A1(_2557_),
    .A2(_2558_),
    .Y(_0363_),
    .B1(net52));
 sg13g2_mux2_1 _5922_ (.A0(\snd.next_note_sel[1] ),
    .A1(_2424_),
    .S(net20),
    .X(_2559_));
 sg13g2_and2_1 _5923_ (.A(_2033_),
    .B(_2559_),
    .X(_0364_));
 sg13g2_mux2_1 _5924_ (.A0(\snd.next_note_timing[0] ),
    .A1(\snd.note_timing[0] ),
    .S(_1568_),
    .X(_2560_));
 sg13g2_and2_1 _5925_ (.A(_2033_),
    .B(_2560_),
    .X(_0365_));
 sg13g2_nand2_1 _5926_ (.Y(_2561_),
    .A(_1548_),
    .B(net20));
 sg13g2_nand2b_1 _5927_ (.Y(_2562_),
    .B(\snd.next_note_timing[1] ),
    .A_N(net20));
 sg13g2_a21oi_1 _5928_ (.A1(_2561_),
    .A2(_2562_),
    .Y(_0366_),
    .B1(net52));
 sg13g2_mux2_1 _5929_ (.A0(\snd.next_note_timing[2] ),
    .A1(\snd.note_timing[2] ),
    .S(_1568_),
    .X(_2563_));
 sg13g2_and2_1 _5930_ (.A(net55),
    .B(_2563_),
    .X(_0367_));
 sg13g2_mux2_1 _5931_ (.A0(\snd.next_note_timing[3] ),
    .A1(\snd.note_timing[3] ),
    .S(_1568_),
    .X(_2564_));
 sg13g2_and2_1 _5932_ (.A(net55),
    .B(_2564_),
    .X(_0368_));
 sg13g2_mux2_1 _5933_ (.A0(\snd.next_note_timing[4] ),
    .A1(_1537_),
    .S(_1568_),
    .X(_2565_));
 sg13g2_and2_1 _5934_ (.A(net95),
    .B(_2565_),
    .X(_0369_));
 sg13g2_mux2_1 _5935_ (.A0(\snd.next_note_timing[5] ),
    .A1(\snd.note_timing[5] ),
    .S(_1568_),
    .X(_2566_));
 sg13g2_and2_1 _5936_ (.A(net95),
    .B(_2566_),
    .X(_0370_));
 sg13g2_nand2_1 _5937_ (.Y(_2567_),
    .A(_1533_),
    .B(net20));
 sg13g2_nand2b_1 _5938_ (.Y(_2568_),
    .B(\snd.next_note_timing[6] ),
    .A_N(_2423_));
 sg13g2_a21oi_1 _5939_ (.A1(_2567_),
    .A2(_2568_),
    .Y(_0371_),
    .B1(net52));
 sg13g2_nand2_1 _5940_ (.Y(_2569_),
    .A(\snd.note_timing[7] ),
    .B(_2423_));
 sg13g2_nand2b_1 _5941_ (.Y(_2570_),
    .B(\snd.next_note_timing[7] ),
    .A_N(net20));
 sg13g2_a21oi_1 _5942_ (.A1(_2569_),
    .A2(_2570_),
    .Y(_0372_),
    .B1(_2389_));
 sg13g2_o21ai_1 _5943_ (.B1(\snd.next_note_timing[8] ),
    .Y(_2571_),
    .A1(_1530_),
    .A2(_1566_));
 sg13g2_nand2b_1 _5944_ (.Y(_2572_),
    .B(_1528_),
    .A_N(_1566_));
 sg13g2_a21oi_1 _5945_ (.A1(_2571_),
    .A2(_2572_),
    .Y(_0373_),
    .B1(_2389_));
 sg13g2_o21ai_1 _5946_ (.B1(_1643_),
    .Y(_2573_),
    .A1(_2356_),
    .A2(_2336_));
 sg13g2_nand2b_1 _5947_ (.Y(_2574_),
    .B(_2307_),
    .A_N(_2300_));
 sg13g2_nand2_1 _5948_ (.Y(_2575_),
    .A(_2573_),
    .B(_2574_));
 sg13g2_buf_2 _5949_ (.A(_2575_),
    .X(_2576_));
 sg13g2_nand4_1 _5950_ (.B(_2329_),
    .C(_2327_),
    .A(_2328_),
    .Y(_2577_),
    .D(_2339_));
 sg13g2_and2_1 _5951_ (.A(_2356_),
    .B(_2577_),
    .X(_2578_));
 sg13g2_buf_1 _5952_ (.A(_2578_),
    .X(_2579_));
 sg13g2_nor3_1 _5953_ (.A(_2304_),
    .B(_2576_),
    .C(_2579_),
    .Y(_2580_));
 sg13g2_and2_1 _5954_ (.A(_2573_),
    .B(_2574_),
    .X(_2581_));
 sg13g2_buf_1 _5955_ (.A(_2581_),
    .X(_2582_));
 sg13g2_nand3_1 _5956_ (.B(_2297_),
    .C(_2343_),
    .A(_1644_),
    .Y(_2583_));
 sg13g2_nand2_1 _5957_ (.Y(_2584_),
    .A(_2311_),
    .B(_2583_));
 sg13g2_a21oi_1 _5958_ (.A1(_2318_),
    .A2(_2584_),
    .Y(_2585_),
    .B1(_2341_));
 sg13g2_nand2b_1 _5959_ (.Y(_2586_),
    .B(_2348_),
    .A_N(_2347_));
 sg13g2_o21ai_1 _5960_ (.B1(_2336_),
    .Y(_2587_),
    .A1(net87),
    .A2(_2334_));
 sg13g2_a21o_1 _5961_ (.A2(_2586_),
    .A1(_2585_),
    .B1(_2587_),
    .X(_2588_));
 sg13g2_a21oi_1 _5962_ (.A1(_2582_),
    .A2(_2588_),
    .Y(_2589_),
    .B1(_2214_));
 sg13g2_nor3_1 _5963_ (.A(net92),
    .B(_2580_),
    .C(_2589_),
    .Y(_0374_));
 sg13g2_nor4_1 _5964_ (.A(net115),
    .B(net112),
    .C(_2304_),
    .D(_2577_),
    .Y(_2590_));
 sg13g2_o21ai_1 _5965_ (.B1(_0971_),
    .Y(_2591_),
    .A1(_2336_),
    .A2(_2590_));
 sg13g2_inv_1 _5966_ (.Y(_0375_),
    .A(_2591_));
 sg13g2_nor2_2 _5967_ (.A(_2338_),
    .B(_2579_),
    .Y(_2592_));
 sg13g2_nor3_1 _5968_ (.A(_2331_),
    .B(_2576_),
    .C(_2592_),
    .Y(_2593_));
 sg13g2_a21oi_1 _5969_ (.A1(_2331_),
    .A2(_2576_),
    .Y(_2594_),
    .B1(_2593_));
 sg13g2_nor2_1 _5970_ (.A(net51),
    .B(_2594_),
    .Y(_0377_));
 sg13g2_nor2_1 _5971_ (.A(_2336_),
    .B(_2579_),
    .Y(_2595_));
 sg13g2_o21ai_1 _5972_ (.B1(_2582_),
    .Y(_2596_),
    .A1(_2331_),
    .A2(_2595_));
 sg13g2_inv_1 _5973_ (.Y(_2597_),
    .A(_2331_));
 sg13g2_nor3_1 _5974_ (.A(_2328_),
    .B(_2597_),
    .C(_2595_),
    .Y(_2598_));
 sg13g2_a22oi_1 _5975_ (.Y(_2599_),
    .B1(_2598_),
    .B2(_2582_),
    .A2(_2596_),
    .A1(_2328_));
 sg13g2_nor2_1 _5976_ (.A(_2541_),
    .B(_2599_),
    .Y(_0378_));
 sg13g2_nand2_1 _5977_ (.Y(_2600_),
    .A(_2328_),
    .B(_2331_));
 sg13g2_nor3_1 _5978_ (.A(_2326_),
    .B(_2576_),
    .C(_2600_),
    .Y(_2601_));
 sg13g2_a21oi_1 _5979_ (.A1(_2326_),
    .A2(_2600_),
    .Y(_2602_),
    .B1(_2601_));
 sg13g2_nor2_1 _5980_ (.A(_2592_),
    .B(_2602_),
    .Y(_2603_));
 sg13g2_a21oi_1 _5981_ (.A1(_2326_),
    .A2(_2576_),
    .Y(_2604_),
    .B1(_2603_));
 sg13g2_nor2_1 _5982_ (.A(net51),
    .B(_2604_),
    .Y(_0379_));
 sg13g2_and3_1 _5983_ (.X(_2605_),
    .A(_2328_),
    .B(_2331_),
    .C(_2326_));
 sg13g2_o21ai_1 _5984_ (.B1(_2582_),
    .Y(_2606_),
    .A1(_2592_),
    .A2(_2605_));
 sg13g2_nor2b_1 _5985_ (.A(_2332_),
    .B_N(_2605_),
    .Y(_2607_));
 sg13g2_nor2_2 _5986_ (.A(_2576_),
    .B(_2592_),
    .Y(_2608_));
 sg13g2_a22oi_1 _5987_ (.Y(_2609_),
    .B1(_2607_),
    .B2(_2608_),
    .A2(_2606_),
    .A1(_2332_));
 sg13g2_nor2_1 _5988_ (.A(net51),
    .B(_2609_),
    .Y(_0380_));
 sg13g2_and2_1 _5989_ (.A(_2332_),
    .B(_2605_),
    .X(_2610_));
 sg13g2_o21ai_1 _5990_ (.B1(_2582_),
    .Y(_2611_),
    .A1(_2592_),
    .A2(_2610_));
 sg13g2_nor2b_1 _5991_ (.A(_2329_),
    .B_N(_2610_),
    .Y(_2612_));
 sg13g2_a22oi_1 _5992_ (.Y(_2613_),
    .B1(_2612_),
    .B2(_2608_),
    .A2(_2611_),
    .A1(_2329_));
 sg13g2_nor2_1 _5993_ (.A(net51),
    .B(_2613_),
    .Y(_0381_));
 sg13g2_and2_1 _5994_ (.A(_2329_),
    .B(_2610_),
    .X(_2614_));
 sg13g2_nor2b_1 _5995_ (.A(_2327_),
    .B_N(_2614_),
    .Y(_2615_));
 sg13g2_o21ai_1 _5996_ (.B1(_2582_),
    .Y(_2616_),
    .A1(_2592_),
    .A2(_2614_));
 sg13g2_a22oi_1 _5997_ (.Y(_2617_),
    .B1(_2616_),
    .B2(_2327_),
    .A2(_2615_),
    .A1(_2608_));
 sg13g2_nor2_1 _5998_ (.A(net51),
    .B(_2617_),
    .Y(_0382_));
 sg13g2_nand2_1 _5999_ (.Y(_2618_),
    .A(_2327_),
    .B(_2614_));
 sg13g2_xor2_1 _6000_ (.B(_2618_),
    .A(_0037_),
    .X(_2619_));
 sg13g2_a22oi_1 _6001_ (.Y(_2620_),
    .B1(_2608_),
    .B2(_2619_),
    .A2(_2576_),
    .A1(\snd.tune_counter[6] ));
 sg13g2_nor2_1 _6002_ (.A(net51),
    .B(_2620_),
    .Y(_0383_));
 sg13g2_nand2b_1 _6003_ (.Y(_2621_),
    .B(_2574_),
    .A_N(_2411_));
 sg13g2_nand2_1 _6004_ (.Y(_2622_),
    .A(net112),
    .B(_2304_));
 sg13g2_nor2_1 _6005_ (.A(net110),
    .B(_2622_),
    .Y(_2623_));
 sg13g2_nor2b_1 _6006_ (.A(_2621_),
    .B_N(_2623_),
    .Y(_2624_));
 sg13g2_a21oi_1 _6007_ (.A1(net110),
    .A2(_2621_),
    .Y(_2625_),
    .B1(_2624_));
 sg13g2_nor2_1 _6008_ (.A(net51),
    .B(_2625_),
    .Y(_0384_));
 sg13g2_o21ai_1 _6009_ (.B1(net109),
    .Y(_2626_),
    .A1(_2621_),
    .A2(_2623_));
 sg13g2_nor2_1 _6010_ (.A(_2622_),
    .B(_2411_),
    .Y(_2627_));
 sg13g2_nand3b_1 _6011_ (.B(_2627_),
    .C(net110),
    .Y(_2628_),
    .A_N(net109));
 sg13g2_a21oi_1 _6012_ (.A1(_2626_),
    .A2(_2628_),
    .Y(_0385_),
    .B1(net52));
 sg13g2_xor2_1 _6013_ (.B(_2377_),
    .A(_2322_),
    .X(_2629_));
 sg13g2_a22oi_1 _6014_ (.Y(_2630_),
    .B1(_2627_),
    .B2(_2629_),
    .A2(_2621_),
    .A1(_2317_));
 sg13g2_nor2_1 _6015_ (.A(net51),
    .B(_2630_),
    .Y(_0386_));
 sg13g2_buf_4 _6016_ (.X(_2631_),
    .A(ui_in[4]));
 sg13g2_xor2_1 _6017_ (.B(net450),
    .A(\dsp.segments_raw[0] ),
    .X(net5));
 sg13g2_xor2_1 _6018_ (.B(\dsp.segments_raw[1] ),
    .A(net450),
    .X(net6));
 sg13g2_xor2_1 _6019_ (.B(\dsp.segments_raw[2] ),
    .A(_2631_),
    .X(net7));
 sg13g2_xor2_1 _6020_ (.B(\dsp.segments_raw[3] ),
    .A(net450),
    .X(net8));
 sg13g2_xor2_1 _6021_ (.B(\dsp.segments_raw[4] ),
    .A(net450),
    .X(net9));
 sg13g2_xor2_1 _6022_ (.B(\dsp.segments_raw[5] ),
    .A(net450),
    .X(net10));
 sg13g2_xor2_1 _6023_ (.B(\dsp.segments_raw[6] ),
    .A(net450),
    .X(net11));
 sg13g2_xor2_1 _6024_ (.B(net450),
    .A(_1780_),
    .X(net17));
 sg13g2_xor2_1 _6025_ (.B(\dsp.digit_sel_raw[1] ),
    .A(net450),
    .X(net18));
 sg13g2_dfrbp_1 _6026_ (.CLK(clknet_leaf_11_clk),
    .RESET_B(net137),
    .D(_0000_),
    .Q_N(_3157_),
    .Q(_0014_));
 sg13g2_dfrbp_1 _6027_ (.CLK(clknet_leaf_15_clk),
    .RESET_B(net138),
    .D(_0001_),
    .Q_N(_3158_),
    .Q(_0015_));
 sg13g2_dfrbp_1 _6028_ (.CLK(clknet_leaf_12_clk),
    .RESET_B(net139),
    .D(_0002_),
    .Q_N(_3159_),
    .Q(_0016_));
 sg13g2_dfrbp_1 _6029_ (.CLK(clknet_leaf_11_clk),
    .RESET_B(net140),
    .D(_0003_),
    .Q_N(_3160_),
    .Q(_0017_));
 sg13g2_dfrbp_1 _6030_ (.CLK(clknet_leaf_11_clk),
    .RESET_B(net141),
    .D(_0004_),
    .Q_N(_3161_),
    .Q(_0018_));
 sg13g2_dfrbp_1 _6031_ (.CLK(clknet_leaf_11_clk),
    .RESET_B(net142),
    .D(_0005_),
    .Q_N(_3162_),
    .Q(_0019_));
 sg13g2_dfrbp_1 _6032_ (.CLK(clknet_leaf_12_clk),
    .RESET_B(net143),
    .D(_0006_),
    .Q_N(_3156_),
    .Q(_0020_));
 sg13g2_dfrbp_1 _6033_ (.CLK(clknet_leaf_29_clk),
    .RESET_B(net144),
    .D(_0095_),
    .Q_N(_3155_),
    .Q(_0007_));
 sg13g2_dfrbp_1 _6034_ (.CLK(clknet_leaf_30_clk),
    .RESET_B(net145),
    .D(_0096_),
    .Q_N(_3154_),
    .Q(_0008_));
 sg13g2_dfrbp_1 _6035_ (.CLK(clknet_leaf_29_clk),
    .RESET_B(net146),
    .D(_0097_),
    .Q_N(_3153_),
    .Q(_0009_));
 sg13g2_buf_2 clkbuf_leaf_0_clk (.A(clknet_3_0__leaf_clk),
    .X(clknet_leaf_0_clk));
 sg13g2_tiehi _6026__137 (.L_HI(net137));
 sg13g2_buf_1 _6038_ (.A(net147),
    .X(uio_oe[0]));
 sg13g2_buf_1 _6039_ (.A(net148),
    .X(uio_oe[1]));
 sg13g2_buf_1 _6040_ (.A(net149),
    .X(uio_oe[2]));
 sg13g2_buf_1 _6041_ (.A(net150),
    .X(uio_oe[3]));
 sg13g2_buf_1 _6042_ (.A(net151),
    .X(uio_oe[4]));
 sg13g2_buf_1 _6043_ (.A(net152),
    .X(uio_oe[5]));
 sg13g2_buf_1 _6044_ (.A(net153),
    .X(uio_oe[6]));
 sg13g2_buf_1 _6045_ (.A(net154),
    .X(uio_oe[7]));
 sg13g2_buf_1 _6046_ (.A(net135),
    .X(uio_out[7]));
 sg13g2_buf_1 _6047_ (.A(\snd.sound ),
    .X(net16));
 sg13g2_buf_1 _6048_ (.A(net136),
    .X(uo_out[7]));
 sg13g2_dfrbp_1 \btn.button_state[0]$_SDFFE_PN0P_  (.CLK(clknet_leaf_20_clk),
    .RESET_B(net155),
    .D(_0098_),
    .Q_N(_3152_),
    .Q(\btn.button_state[0] ));
 sg13g2_dfrbp_1 \btn.button_state[1]$_SDFFE_PN0P_  (.CLK(clknet_leaf_19_clk),
    .RESET_B(net156),
    .D(_0099_),
    .Q_N(_3151_),
    .Q(\btn.button_state[1] ));
 sg13g2_dfrbp_1 \btn.button_state[2]$_SDFFE_PN0P_  (.CLK(clknet_leaf_21_clk),
    .RESET_B(net157),
    .D(_0100_),
    .Q_N(_3150_),
    .Q(\btn.button_state[2] ));
 sg13g2_dfrbp_1 \btn.button_state[3]$_SDFFE_PN0P_  (.CLK(clknet_leaf_22_clk),
    .RESET_B(net158),
    .D(_0101_),
    .Q_N(_3149_),
    .Q(\btn.button_state[3] ));
 sg13g2_dfrbp_1 \btn.change_timer[0]$_SDFFE_PN0P_  (.CLK(clknet_leaf_13_clk),
    .RESET_B(net159),
    .D(_0102_),
    .Q_N(_3148_),
    .Q(\btn.change_timer[0] ));
 sg13g2_dfrbp_1 \btn.change_timer[1]$_SDFFE_PN0P_  (.CLK(clknet_leaf_14_clk),
    .RESET_B(net160),
    .D(_0103_),
    .Q_N(_3147_),
    .Q(\btn.change_timer[1] ));
 sg13g2_dfrbp_1 \btn.change_timer[2]$_SDFFE_PN0P_  (.CLK(clknet_leaf_14_clk),
    .RESET_B(net161),
    .D(_0104_),
    .Q_N(_3146_),
    .Q(\btn.change_timer[2] ));
 sg13g2_dfrbp_1 \btn.change_timer[3]$_SDFFE_PN0P_  (.CLK(clknet_leaf_19_clk),
    .RESET_B(net162),
    .D(_0105_),
    .Q_N(_3145_),
    .Q(\btn.change_timer[3] ));
 sg13g2_dfrbp_1 \btn.change_timer[4]$_SDFFE_PN0P_  (.CLK(clknet_leaf_19_clk),
    .RESET_B(net163),
    .D(_0106_),
    .Q_N(_3144_),
    .Q(\btn.change_timer[4] ));
 sg13g2_dfrbp_1 \btn.change_timer[5]$_SDFFE_PN0P_  (.CLK(clknet_leaf_18_clk),
    .RESET_B(net164),
    .D(_0107_),
    .Q_N(_3143_),
    .Q(\btn.change_timer[5] ));
 sg13g2_dfrbp_1 \btn.change_timer[6]$_SDFFE_PN0P_  (.CLK(clknet_leaf_14_clk),
    .RESET_B(net165),
    .D(_0108_),
    .Q_N(_3142_),
    .Q(\btn.change_timer[6] ));
 sg13g2_dfrbp_1 \btn.current_event[0]$_SDFFE_PN0P_  (.CLK(clknet_leaf_19_clk),
    .RESET_B(net166),
    .D(_0109_),
    .Q_N(_3141_),
    .Q(\btn.current_event[0] ));
 sg13g2_dfrbp_1 \btn.current_event[1]$_SDFFE_PN0P_  (.CLK(clknet_leaf_19_clk),
    .RESET_B(net167),
    .D(_0110_),
    .Q_N(_3140_),
    .Q(\btn.current_event[1] ));
 sg13g2_dfrbp_1 \btn.current_event[2]$_SDFFE_PN0P_  (.CLK(clknet_leaf_19_clk),
    .RESET_B(net168),
    .D(_0111_),
    .Q_N(_3139_),
    .Q(\btn.current_event[2] ));
 sg13g2_dfrbp_1 \btn.current_event[3]$_SDFFE_PN0P_  (.CLK(clknet_leaf_19_clk),
    .RESET_B(net169),
    .D(_0112_),
    .Q_N(_3138_),
    .Q(\btn.current_event[3] ));
 sg13g2_dfrbp_1 \btn.input_event[0]$_SDFF_PN0_  (.CLK(clknet_leaf_17_clk),
    .RESET_B(net170),
    .D(_0113_),
    .Q_N(_3137_),
    .Q(\btn.input_event[0] ));
 sg13g2_dfrbp_1 \btn.input_event[1]$_SDFF_PN0_  (.CLK(clknet_leaf_20_clk),
    .RESET_B(net171),
    .D(_0114_),
    .Q_N(_3136_),
    .Q(\btn.input_event[1] ));
 sg13g2_dfrbp_1 \btn.input_event[2]$_SDFF_PN0_  (.CLK(clknet_leaf_18_clk),
    .RESET_B(net172),
    .D(_0115_),
    .Q_N(_3135_),
    .Q(\btn.input_event[2] ));
 sg13g2_dfrbp_1 \btn.input_event[3]$_SDFF_PN0_  (.CLK(clknet_leaf_20_clk),
    .RESET_B(net173),
    .D(_0116_),
    .Q_N(_3134_),
    .Q(\btn.input_event[3] ));
 sg13g2_dfrbp_1 \btn.input_event[4]$_SDFF_PN0_  (.CLK(clknet_leaf_18_clk),
    .RESET_B(net174),
    .D(_0117_),
    .Q_N(_0034_),
    .Q(\btn.input_event[4] ));
 sg13g2_dfrbp_1 \btn.long_press$_SDFFE_PN0P_  (.CLK(clknet_leaf_19_clk),
    .RESET_B(net175),
    .D(_0118_),
    .Q_N(_3133_),
    .Q(\btn.long_press ));
 sg13g2_dfrbp_1 \btn.sample_10ms[0]$_SDFFE_PN0P_  (.CLK(clknet_leaf_20_clk),
    .RESET_B(net176),
    .D(_0119_),
    .Q_N(_3132_),
    .Q(\btn.sample_10ms[0] ));
 sg13g2_dfrbp_1 \btn.sample_10ms[1]$_SDFFE_PN0P_  (.CLK(clknet_leaf_17_clk),
    .RESET_B(net177),
    .D(_0120_),
    .Q_N(_3131_),
    .Q(\btn.sample_10ms[1] ));
 sg13g2_dfrbp_1 \btn.sample_10ms[2]$_SDFFE_PN0P_  (.CLK(clknet_leaf_21_clk),
    .RESET_B(net178),
    .D(_0121_),
    .Q_N(_3130_),
    .Q(\btn.sample_10ms[2] ));
 sg13g2_dfrbp_1 \btn.sample_10ms[3]$_SDFFE_PN0P_  (.CLK(clknet_leaf_17_clk),
    .RESET_B(net179),
    .D(_0122_),
    .Q_N(_3129_),
    .Q(\btn.sample_10ms[3] ));
 sg13g2_dfrbp_1 \btn.sample_15ms[0]$_SDFFE_PN0P_  (.CLK(clknet_leaf_20_clk),
    .RESET_B(net180),
    .D(_0123_),
    .Q_N(_3128_),
    .Q(\btn.sample_15ms[0] ));
 sg13g2_dfrbp_1 \btn.sample_15ms[1]$_SDFFE_PN0P_  (.CLK(clknet_leaf_17_clk),
    .RESET_B(net181),
    .D(_0124_),
    .Q_N(_3127_),
    .Q(\btn.sample_15ms[1] ));
 sg13g2_dfrbp_1 \btn.sample_15ms[2]$_SDFFE_PN0P_  (.CLK(clknet_leaf_20_clk),
    .RESET_B(net182),
    .D(_0125_),
    .Q_N(_3126_),
    .Q(\btn.sample_15ms[2] ));
 sg13g2_dfrbp_1 \btn.sample_15ms[3]$_SDFFE_PN0P_  (.CLK(clknet_leaf_27_clk),
    .RESET_B(net183),
    .D(_0126_),
    .Q_N(_3125_),
    .Q(\btn.sample_15ms[3] ));
 sg13g2_dfrbp_1 \btn.sample_5ms[0]$_SDFFE_PN0P_  (.CLK(clknet_leaf_20_clk),
    .RESET_B(net184),
    .D(_0127_),
    .Q_N(_3124_),
    .Q(\btn.sample_5ms[0] ));
 sg13g2_dfrbp_1 \btn.sample_5ms[1]$_SDFFE_PN0P_  (.CLK(clknet_leaf_20_clk),
    .RESET_B(net185),
    .D(_0128_),
    .Q_N(_3123_),
    .Q(\btn.sample_5ms[1] ));
 sg13g2_dfrbp_1 \btn.sample_5ms[2]$_SDFFE_PN0P_  (.CLK(clknet_leaf_21_clk),
    .RESET_B(net186),
    .D(_0129_),
    .Q_N(_3122_),
    .Q(\btn.sample_5ms[2] ));
 sg13g2_dfrbp_1 \btn.sample_5ms[3]$_SDFFE_PN0P_  (.CLK(clknet_leaf_24_clk),
    .RESET_B(net187),
    .D(_0130_),
    .Q_N(_3121_),
    .Q(\btn.sample_5ms[3] ));
 sg13g2_dfrbp_1 \clk_div_counter[0]$_SDFF_PP0_  (.CLK(clknet_leaf_10_clk),
    .RESET_B(net188),
    .D(_0131_),
    .Q_N(_0094_),
    .Q(\clk_div_counter[0] ));
 sg13g2_dfrbp_1 \clk_div_counter[1]$_SDFF_PP0_  (.CLK(clknet_leaf_10_clk),
    .RESET_B(net189),
    .D(_0132_),
    .Q_N(_3120_),
    .Q(\clk_div_counter[1] ));
 sg13g2_dfrbp_1 \clk_div_counter[2]$_SDFF_PP0_  (.CLK(clknet_leaf_11_clk),
    .RESET_B(net190),
    .D(_0133_),
    .Q_N(_3119_),
    .Q(\clk_div_counter[2] ));
 sg13g2_dfrbp_1 \clk_div_counter[3]$_SDFF_PP0_  (.CLK(clknet_leaf_10_clk),
    .RESET_B(net191),
    .D(_0134_),
    .Q_N(_3118_),
    .Q(\clk_div_counter[3] ));
 sg13g2_dfrbp_1 \clk_div_counter[4]$_SDFF_PP0_  (.CLK(clknet_leaf_10_clk),
    .RESET_B(net192),
    .D(_0135_),
    .Q_N(_3117_),
    .Q(\clk_div_counter[4] ));
 sg13g2_dfrbp_1 \clk_div_counter[5]$_SDFF_PP0_  (.CLK(clknet_leaf_9_clk),
    .RESET_B(net193),
    .D(_0136_),
    .Q_N(_3116_),
    .Q(\clk_div_counter[5] ));
 sg13g2_dfrbp_1 \clk_div_counter[6]$_SDFF_PP0_  (.CLK(clknet_leaf_10_clk),
    .RESET_B(net194),
    .D(_0137_),
    .Q_N(_3115_),
    .Q(\clk_div_counter[6] ));
 sg13g2_dfrbp_1 \clk_div_counter[7]$_SDFF_PP0_  (.CLK(clknet_leaf_11_clk),
    .RESET_B(net195),
    .D(_0138_),
    .Q_N(_3114_),
    .Q(\clk_div_counter[7] ));
 sg13g2_dfrbp_1 \dsp.digit_sel_raw[0]$_SDFF_PN0_  (.CLK(clknet_leaf_11_clk),
    .RESET_B(net196),
    .D(_0139_),
    .Q_N(_0021_),
    .Q(\dsp.digit ));
 sg13g2_dfrbp_1 \dsp.digit_sel_raw[1]$_SDFF_PN0_  (.CLK(clknet_leaf_14_clk),
    .RESET_B(net197),
    .D(_0140_),
    .Q_N(_3113_),
    .Q(\dsp.digit_sel_raw[1] ));
 sg13g2_dfrbp_1 \dsp.segments_raw[0]$_SDFF_PN0_  (.CLK(clknet_leaf_13_clk),
    .RESET_B(net198),
    .D(_0141_),
    .Q_N(_3112_),
    .Q(\dsp.segments_raw[0] ));
 sg13g2_dfrbp_1 \dsp.segments_raw[1]$_SDFF_PN0_  (.CLK(clknet_leaf_13_clk),
    .RESET_B(net199),
    .D(_0142_),
    .Q_N(_3111_),
    .Q(\dsp.segments_raw[1] ));
 sg13g2_dfrbp_1 \dsp.segments_raw[2]$_SDFF_PN0_  (.CLK(clknet_leaf_13_clk),
    .RESET_B(net200),
    .D(_0143_),
    .Q_N(_3110_),
    .Q(\dsp.segments_raw[2] ));
 sg13g2_dfrbp_1 \dsp.segments_raw[3]$_SDFF_PN0_  (.CLK(clknet_leaf_13_clk),
    .RESET_B(net201),
    .D(_0144_),
    .Q_N(_3109_),
    .Q(\dsp.segments_raw[3] ));
 sg13g2_dfrbp_1 \dsp.segments_raw[4]$_SDFF_PN0_  (.CLK(clknet_leaf_13_clk),
    .RESET_B(net202),
    .D(_0145_),
    .Q_N(_3108_),
    .Q(\dsp.segments_raw[4] ));
 sg13g2_dfrbp_1 \dsp.segments_raw[5]$_SDFF_PN0_  (.CLK(clknet_leaf_13_clk),
    .RESET_B(net203),
    .D(_0146_),
    .Q_N(_3107_),
    .Q(\dsp.segments_raw[5] ));
 sg13g2_dfrbp_1 \dsp.segments_raw[6]$_SDFF_PN0_  (.CLK(clknet_leaf_13_clk),
    .RESET_B(net204),
    .D(_0147_),
    .Q_N(_3106_),
    .Q(\dsp.segments_raw[6] ));
 sg13g2_dfrbp_1 \game.challenge_mode$_SDFFE_PN0P_  (.CLK(clknet_leaf_16_clk),
    .RESET_B(net205),
    .D(_0148_),
    .Q_N(_3105_),
    .Q(\game.challenge_mode ));
 sg13g2_dfrbp_1 \game.challenge_num[0]$_SDFFE_PN0P_  (.CLK(clknet_leaf_15_clk),
    .RESET_B(net206),
    .D(_0149_),
    .Q_N(_3104_),
    .Q(\game.challenge_num[0] ));
 sg13g2_dfrbp_1 \game.challenge_num[1]$_SDFFE_PN0P_  (.CLK(clknet_leaf_15_clk),
    .RESET_B(net207),
    .D(_0150_),
    .Q_N(_0052_),
    .Q(\game.challenge_num[1] ));
 sg13g2_dfrbp_1 \game.challenge_num[2]$_SDFFE_PN0P_  (.CLK(clknet_leaf_14_clk),
    .RESET_B(net208),
    .D(_0151_),
    .Q_N(_0054_),
    .Q(\game.challenge_num[2] ));
 sg13g2_dfrbp_1 \game.challenge_num[3]$_SDFFE_PN0P_  (.CLK(clknet_leaf_14_clk),
    .RESET_B(net209),
    .D(_0152_),
    .Q_N(_0055_),
    .Q(\game.challenge_num[3] ));
 sg13g2_dfrbp_1 \game.counter[0]$_SDFFE_PN0P_  (.CLK(clknet_leaf_39_clk),
    .RESET_B(net210),
    .D(_0153_),
    .Q_N(_3103_),
    .Q(\game.counter[0] ));
 sg13g2_dfrbp_1 \game.counter[1]$_SDFFE_PN0P_  (.CLK(clknet_leaf_39_clk),
    .RESET_B(net211),
    .D(_0154_),
    .Q_N(_3102_),
    .Q(\game.counter[1] ));
 sg13g2_dfrbp_1 \game.counter[2]$_SDFFE_PN0P_  (.CLK(clknet_leaf_29_clk),
    .RESET_B(net212),
    .D(_0155_),
    .Q_N(_3101_),
    .Q(\game.counter[2] ));
 sg13g2_dfrbp_1 \game.counter[3]$_SDFFE_PN0P_  (.CLK(clknet_leaf_39_clk),
    .RESET_B(net213),
    .D(_0156_),
    .Q_N(_3100_),
    .Q(\game.counter[3] ));
 sg13g2_dfrbp_1 \game.counter[4]$_SDFFE_PN0P_  (.CLK(clknet_leaf_39_clk),
    .RESET_B(net214),
    .D(_0157_),
    .Q_N(_3099_),
    .Q(\game.counter[4] ));
 sg13g2_dfrbp_1 \game.counter[5]$_SDFFE_PN0P_  (.CLK(clknet_leaf_29_clk),
    .RESET_B(net215),
    .D(_0158_),
    .Q_N(_3098_),
    .Q(\game.counter[5] ));
 sg13g2_dfrbp_1 \game.counter[6]$_SDFFE_PN0P_  (.CLK(clknet_leaf_40_clk),
    .RESET_B(net216),
    .D(_0159_),
    .Q_N(_3097_),
    .Q(\game.counter[6] ));
 sg13g2_dfrbp_1 \game.counter[7]$_SDFFE_PN0P_  (.CLK(clknet_leaf_28_clk),
    .RESET_B(net217),
    .D(_0160_),
    .Q_N(_3096_),
    .Q(\game.counter[7] ));
 sg13g2_dfrbp_1 \game.current_level[0]$_SDFFE_PN0P_  (.CLK(clknet_leaf_3_clk),
    .RESET_B(net218),
    .D(_0161_),
    .Q_N(_0069_),
    .Q(\game.current_level[0] ));
 sg13g2_dfrbp_1 \game.current_level[1]$_SDFFE_PN0P_  (.CLK(clknet_leaf_3_clk),
    .RESET_B(net219),
    .D(_0162_),
    .Q_N(_3095_),
    .Q(\game.current_level[1] ));
 sg13g2_dfrbp_1 \game.current_level[2]$_SDFFE_PN0P_  (.CLK(clknet_leaf_3_clk),
    .RESET_B(net220),
    .D(_0163_),
    .Q_N(_0063_),
    .Q(\game.current_level[2] ));
 sg13g2_dfrbp_1 \game.current_level[3]$_SDFFE_PN0P_  (.CLK(clknet_leaf_3_clk),
    .RESET_B(net221),
    .D(_0164_),
    .Q_N(_0062_),
    .Q(\game.current_level[3] ));
 sg13g2_dfrbp_1 \game.current_level[4]$_SDFFE_PN0P_  (.CLK(clknet_leaf_3_clk),
    .RESET_B(net222),
    .D(_0165_),
    .Q_N(_0061_),
    .Q(\game.current_level[4] ));
 sg13g2_dfrbp_1 \game.display_graphical$_SDFFE_PN0P_  (.CLK(clknet_leaf_14_clk),
    .RESET_B(net223),
    .D(_0166_),
    .Q_N(_3094_),
    .Q(display_graphical));
 sg13g2_dfrbp_1 \game.display_value[0]$_SDFFE_PN1P_  (.CLK(clknet_leaf_12_clk),
    .RESET_B(net224),
    .D(_0167_),
    .Q_N(_0058_),
    .Q(\display_value[0] ));
 sg13g2_dfrbp_1 \game.display_value[1]$_SDFFE_PN0P_  (.CLK(clknet_leaf_11_clk),
    .RESET_B(net225),
    .D(_0168_),
    .Q_N(_3093_),
    .Q(\display_value[1] ));
 sg13g2_dfrbp_1 \game.display_value[2]$_SDFFE_PN0P_  (.CLK(clknet_leaf_15_clk),
    .RESET_B(net226),
    .D(_0169_),
    .Q_N(_0053_),
    .Q(\display_value[2] ));
 sg13g2_dfrbp_1 \game.display_value[3]$_SDFFE_PN0P_  (.CLK(clknet_leaf_12_clk),
    .RESET_B(net227),
    .D(_0170_),
    .Q_N(_3092_),
    .Q(\display_value[3] ));
 sg13g2_dfrbp_1 \game.display_value[4]$_SDFFE_PN0P_  (.CLK(clknet_leaf_12_clk),
    .RESET_B(net228),
    .D(_0171_),
    .Q_N(_0059_),
    .Q(\display_value[4] ));
 sg13g2_dfrbp_1 \game.fsm.block_len[0][0]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_45_clk),
    .RESET_B(net229),
    .D(_0172_),
    .Q_N(_0087_),
    .Q(\game.fsm.block_len[0][0] ));
 sg13g2_dfrbp_1 \game.fsm.block_len[0][1]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_45_clk),
    .RESET_B(net230),
    .D(_0173_),
    .Q_N(_0091_),
    .Q(\game.fsm.block_len[0][1] ));
 sg13g2_dfrbp_1 \game.fsm.block_len[0][2]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_45_clk),
    .RESET_B(net231),
    .D(_0174_),
    .Q_N(_0089_),
    .Q(\game.fsm.block_len[0][2] ));
 sg13g2_dfrbp_1 \game.fsm.block_len[1][0]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_45_clk),
    .RESET_B(net232),
    .D(_0175_),
    .Q_N(_0086_),
    .Q(\game.fsm.block_len[1][0] ));
 sg13g2_dfrbp_1 \game.fsm.block_len[1][1]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_45_clk),
    .RESET_B(net233),
    .D(_0176_),
    .Q_N(_0090_),
    .Q(\game.fsm.block_len[1][1] ));
 sg13g2_dfrbp_1 \game.fsm.block_len[1][2]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_45_clk),
    .RESET_B(net234),
    .D(_0177_),
    .Q_N(_0088_),
    .Q(\game.fsm.block_len[1][2] ));
 sg13g2_dfrbp_1 \game.fsm.block_len[2][0]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_45_clk),
    .RESET_B(net235),
    .D(_0178_),
    .Q_N(_0084_),
    .Q(\game.fsm.block_len[2][0] ));
 sg13g2_dfrbp_1 \game.fsm.block_len[2][1]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_0_clk),
    .RESET_B(net236),
    .D(_0179_),
    .Q_N(_0093_),
    .Q(\game.fsm.block_len[2][1] ));
 sg13g2_dfrbp_1 \game.fsm.block_len[2][2]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_0_clk),
    .RESET_B(net237),
    .D(_0180_),
    .Q_N(_0027_),
    .Q(\game.fsm.block_len[2][2] ));
 sg13g2_dfrbp_1 \game.fsm.block_len[3][0]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_0_clk),
    .RESET_B(net238),
    .D(_0181_),
    .Q_N(_0083_),
    .Q(\game.fsm.block_len[3][0] ));
 sg13g2_dfrbp_1 \game.fsm.block_len[3][1]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_0_clk),
    .RESET_B(net239),
    .D(_0182_),
    .Q_N(_0092_),
    .Q(\game.fsm.block_len[3][1] ));
 sg13g2_dfrbp_1 \game.fsm.block_len[3][2]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_0_clk),
    .RESET_B(net240),
    .D(_0183_),
    .Q_N(_0026_),
    .Q(\game.fsm.block_len[3][2] ));
 sg13g2_dfrbp_1 \game.fsm.block_len[4][0]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_1_clk),
    .RESET_B(net241),
    .D(_0184_),
    .Q_N(_0076_),
    .Q(\game.fsm.block_len[4][0] ));
 sg13g2_dfrbp_1 \game.fsm.block_len[4][1]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_1_clk),
    .RESET_B(net242),
    .D(_0185_),
    .Q_N(_0078_),
    .Q(\game.fsm.block_len[4][1] ));
 sg13g2_dfrbp_1 \game.fsm.block_len[4][2]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_6_clk),
    .RESET_B(net243),
    .D(_0186_),
    .Q_N(_0081_),
    .Q(\game.fsm.block_len[4][2] ));
 sg13g2_dfrbp_1 \game.fsm.block_len[5][0]$_DFFE_PP_  (.CLK(clknet_leaf_1_clk),
    .RESET_B(net244),
    .D(_0187_),
    .Q_N(_0075_),
    .Q(\game.fsm.block_len[5][0] ));
 sg13g2_dfrbp_1 \game.fsm.block_len[5][1]$_DFFE_PP_  (.CLK(clknet_leaf_6_clk),
    .RESET_B(net245),
    .D(_0188_),
    .Q_N(_0077_),
    .Q(\game.fsm.block_len[5][1] ));
 sg13g2_dfrbp_1 \game.fsm.block_len[5][2]$_DFFE_PP_  (.CLK(clknet_leaf_6_clk),
    .RESET_B(net246),
    .D(_0189_),
    .Q_N(_0080_),
    .Q(\game.fsm.block_len[5][2] ));
 sg13g2_dfrbp_1 \game.fsm.block_len[6][0]$_SDFFE_PP0P_  (.CLK(clknet_leaf_1_clk),
    .RESET_B(net247),
    .D(_0190_),
    .Q_N(_0074_),
    .Q(\game.fsm.block_len[6][0] ));
 sg13g2_dfrbp_1 \game.fsm.block_len[6][1]$_SDFFE_PP0P_  (.CLK(clknet_leaf_6_clk),
    .RESET_B(net248),
    .D(_0191_),
    .Q_N(_0082_),
    .Q(\game.fsm.block_len[6][1] ));
 sg13g2_dfrbp_1 \game.fsm.block_len[6][2]$_SDFFE_PP0P_  (.CLK(clknet_leaf_6_clk),
    .RESET_B(net249),
    .D(_0192_),
    .Q_N(_0079_),
    .Q(\game.fsm.block_len[6][2] ));
 sg13g2_dfrbp_1 \game.fsm.block_len[7][0]$_DFFE_PP_  (.CLK(clknet_leaf_45_clk),
    .RESET_B(net250),
    .D(_0193_),
    .Q_N(_3091_),
    .Q(\game.fsm.block_len[7][0] ));
 sg13g2_dfrbp_1 \game.fsm.block_len[7][1]$_DFFE_PP_  (.CLK(clknet_leaf_0_clk),
    .RESET_B(net251),
    .D(_0194_),
    .Q_N(_3090_),
    .Q(\game.fsm.block_len[7][1] ));
 sg13g2_dfrbp_1 \game.fsm.block_len[7][2]$_DFFE_PP_  (.CLK(clknet_leaf_0_clk),
    .RESET_B(net252),
    .D(_0195_),
    .Q_N(_3089_),
    .Q(\game.fsm.block_len[7][2] ));
 sg13g2_dfrbp_1 \game.fsm.color_count[0][0]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_36_clk),
    .RESET_B(net253),
    .D(_0196_),
    .Q_N(_3088_),
    .Q(\game.fsm.color_count[0][0] ));
 sg13g2_dfrbp_1 \game.fsm.color_count[0][1]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_37_clk),
    .RESET_B(net254),
    .D(_0197_),
    .Q_N(_3087_),
    .Q(\game.fsm.color_count[0][1] ));
 sg13g2_dfrbp_1 \game.fsm.color_count[0][2]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_37_clk),
    .RESET_B(net255),
    .D(_0198_),
    .Q_N(_3086_),
    .Q(\game.fsm.color_count[0][2] ));
 sg13g2_dfrbp_1 \game.fsm.color_count[1][0]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_37_clk),
    .RESET_B(net256),
    .D(_0199_),
    .Q_N(_3085_),
    .Q(\game.fsm.color_count[1][0] ));
 sg13g2_dfrbp_1 \game.fsm.color_count[1][1]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_37_clk),
    .RESET_B(net257),
    .D(_0200_),
    .Q_N(_3084_),
    .Q(\game.fsm.color_count[1][1] ));
 sg13g2_dfrbp_1 \game.fsm.color_count[1][2]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_38_clk),
    .RESET_B(net258),
    .D(_0201_),
    .Q_N(_0070_),
    .Q(\game.fsm.color_count[1][2] ));
 sg13g2_dfrbp_1 \game.fsm.color_count[2][0]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_36_clk),
    .RESET_B(net259),
    .D(_0202_),
    .Q_N(_3083_),
    .Q(\game.fsm.color_count[2][0] ));
 sg13g2_dfrbp_1 \game.fsm.color_count[2][1]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_36_clk),
    .RESET_B(net260),
    .D(_0203_),
    .Q_N(_3082_),
    .Q(\game.fsm.color_count[2][1] ));
 sg13g2_dfrbp_1 \game.fsm.color_count[2][2]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_36_clk),
    .RESET_B(net261),
    .D(_0204_),
    .Q_N(_0072_),
    .Q(\game.fsm.color_count[2][2] ));
 sg13g2_dfrbp_1 \game.fsm.color_count[3][0]$_DFFE_PP_  (.CLK(clknet_leaf_36_clk),
    .RESET_B(net262),
    .D(_0205_),
    .Q_N(_3081_),
    .Q(\game.fsm.color_count[3][0] ));
 sg13g2_dfrbp_1 \game.fsm.color_count[3][1]$_DFFE_PP_  (.CLK(clknet_leaf_36_clk),
    .RESET_B(net263),
    .D(_0206_),
    .Q_N(_3080_),
    .Q(\game.fsm.color_count[3][1] ));
 sg13g2_dfrbp_1 \game.fsm.color_count[3][2]$_DFFE_PP_  (.CLK(clknet_leaf_38_clk),
    .RESET_B(net264),
    .D(_0207_),
    .Q_N(_0071_),
    .Q(\game.fsm.color_count[3][2] ));
 sg13g2_dfrbp_1 \game.fsm.green_block_count[0]$_SDFFE_PP0P_  (.CLK(clknet_leaf_41_clk),
    .RESET_B(net265),
    .D(_0208_),
    .Q_N(_3079_),
    .Q(\game.fsm.green_block_count[0] ));
 sg13g2_dfrbp_1 \game.fsm.green_block_count[1]$_SDFFE_PP0P_  (.CLK(clknet_leaf_39_clk),
    .RESET_B(net266),
    .D(_0209_),
    .Q_N(_3078_),
    .Q(\game.fsm.green_block_count[1] ));
 sg13g2_dfrbp_1 \game.fsm.green_block_count[2]$_SDFFE_PP0P_  (.CLK(clknet_leaf_39_clk),
    .RESET_B(net267),
    .D(_0210_),
    .Q_N(_3077_),
    .Q(\game.fsm.green_block_count[2] ));
 sg13g2_dfrbp_1 \game.fsm.len1_block_count[0]$_SDFFE_PP0P_  (.CLK(clknet_leaf_40_clk),
    .RESET_B(net268),
    .D(_0211_),
    .Q_N(_3076_),
    .Q(\game.fsm.len1_block_count[0] ));
 sg13g2_dfrbp_1 \game.fsm.len1_block_count[1]$_SDFFE_PP0P_  (.CLK(clknet_leaf_40_clk),
    .RESET_B(net269),
    .D(_0212_),
    .Q_N(_3075_),
    .Q(\game.fsm.len1_block_count[1] ));
 sg13g2_dfrbp_1 \game.fsm.len1_block_count[2]$_SDFFE_PP0P_  (.CLK(clknet_leaf_40_clk),
    .RESET_B(net270),
    .D(_0213_),
    .Q_N(_3074_),
    .Q(\game.fsm.len1_block_count[2] ));
 sg13g2_dfrbp_1 \game.fsm.len1_color_count[0][0]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_42_clk),
    .RESET_B(net271),
    .D(_0214_),
    .Q_N(_3073_),
    .Q(\game.fsm.len1_color_count[0][0] ));
 sg13g2_dfrbp_1 \game.fsm.len1_color_count[0][1]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_38_clk),
    .RESET_B(net272),
    .D(_0215_),
    .Q_N(_0040_),
    .Q(\game.fsm.len1_color_count[0][1] ));
 sg13g2_dfrbp_1 \game.fsm.len1_color_count[0][2]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_42_clk),
    .RESET_B(net273),
    .D(_0216_),
    .Q_N(_0022_),
    .Q(\game.fsm.len1_color_count[0][2] ));
 sg13g2_dfrbp_1 \game.fsm.len1_color_count[1][0]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_37_clk),
    .RESET_B(net274),
    .D(_0217_),
    .Q_N(_3072_),
    .Q(\game.fsm.len1_color_count[1][0] ));
 sg13g2_dfrbp_1 \game.fsm.len1_color_count[1][1]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_38_clk),
    .RESET_B(net275),
    .D(_0218_),
    .Q_N(_0041_),
    .Q(\game.fsm.len1_color_count[1][1] ));
 sg13g2_dfrbp_1 \game.fsm.len1_color_count[1][2]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_37_clk),
    .RESET_B(net276),
    .D(_0219_),
    .Q_N(_0023_),
    .Q(\game.fsm.len1_color_count[1][2] ));
 sg13g2_dfrbp_1 \game.fsm.len1_color_count[2][0]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_39_clk),
    .RESET_B(net277),
    .D(_0220_),
    .Q_N(_3071_),
    .Q(\game.fsm.len1_color_count[2][0] ));
 sg13g2_dfrbp_1 \game.fsm.len1_color_count[2][1]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_38_clk),
    .RESET_B(net278),
    .D(_0221_),
    .Q_N(_0042_),
    .Q(\game.fsm.len1_color_count[2][1] ));
 sg13g2_dfrbp_1 \game.fsm.len1_color_count[2][2]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_38_clk),
    .RESET_B(net279),
    .D(_0222_),
    .Q_N(_0025_),
    .Q(\game.fsm.len1_color_count[2][2] ));
 sg13g2_dfrbp_1 \game.fsm.len1_color_count[3][0]$_DFFE_PP_  (.CLK(clknet_leaf_37_clk),
    .RESET_B(net280),
    .D(_0223_),
    .Q_N(_3070_),
    .Q(\game.fsm.len1_color_count[3][0] ));
 sg13g2_dfrbp_1 \game.fsm.len1_color_count[3][1]$_DFFE_PP_  (.CLK(clknet_leaf_38_clk),
    .RESET_B(net281),
    .D(_0224_),
    .Q_N(_0043_),
    .Q(\game.fsm.len1_color_count[3][1] ));
 sg13g2_dfrbp_1 \game.fsm.len1_color_count[3][2]$_DFFE_PP_  (.CLK(clknet_leaf_37_clk),
    .RESET_B(net282),
    .D(_0225_),
    .Q_N(_0024_),
    .Q(\game.fsm.len1_color_count[3][2] ));
 sg13g2_dfrbp_1 \game.fsm.len2_block_count[0]$_SDFFE_PP0P_  (.CLK(clknet_leaf_41_clk),
    .RESET_B(net283),
    .D(_0226_),
    .Q_N(_3069_),
    .Q(\game.fsm.len2_block_count[0] ));
 sg13g2_dfrbp_1 \game.fsm.len2_block_count[1]$_SDFFE_PP0P_  (.CLK(clknet_leaf_40_clk),
    .RESET_B(net284),
    .D(_0227_),
    .Q_N(_3068_),
    .Q(\game.fsm.len2_block_count[1] ));
 sg13g2_dfrbp_1 \game.fsm.len2_color_count[0][0]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_43_clk),
    .RESET_B(net285),
    .D(_0228_),
    .Q_N(_3067_),
    .Q(\game.fsm.len2_color_count[0][0] ));
 sg13g2_dfrbp_1 \game.fsm.len2_color_count[0][1]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_43_clk),
    .RESET_B(net286),
    .D(_0229_),
    .Q_N(_0044_),
    .Q(\game.fsm.len2_color_count[0][1] ));
 sg13g2_dfrbp_1 \game.fsm.len2_color_count[1][0]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_44_clk),
    .RESET_B(net287),
    .D(_0230_),
    .Q_N(_3066_),
    .Q(\game.fsm.len2_color_count[1][0] ));
 sg13g2_dfrbp_1 \game.fsm.len2_color_count[1][1]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_44_clk),
    .RESET_B(net288),
    .D(_0231_),
    .Q_N(_0045_),
    .Q(\game.fsm.len2_color_count[1][1] ));
 sg13g2_dfrbp_1 \game.fsm.len2_color_count[2][0]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_43_clk),
    .RESET_B(net289),
    .D(_0232_),
    .Q_N(_3065_),
    .Q(\game.fsm.len2_color_count[2][0] ));
 sg13g2_dfrbp_1 \game.fsm.len2_color_count[2][1]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_43_clk),
    .RESET_B(net290),
    .D(_0233_),
    .Q_N(_0046_),
    .Q(\game.fsm.len2_color_count[2][1] ));
 sg13g2_dfrbp_1 \game.fsm.len2_color_count[3][0]$_DFFE_PP_  (.CLK(clknet_leaf_44_clk),
    .RESET_B(net291),
    .D(_0234_),
    .Q_N(_3064_),
    .Q(\game.fsm.len2_color_count[3][0] ));
 sg13g2_dfrbp_1 \game.fsm.len2_color_count[3][1]$_DFFE_PP_  (.CLK(clknet_leaf_43_clk),
    .RESET_B(net292),
    .D(_0235_),
    .Q_N(_0047_),
    .Q(\game.fsm.len2_color_count[3][1] ));
 sg13g2_dfrbp_1 \game.fsm.len3_block_count[0]$_SDFFE_PP0P_  (.CLK(clknet_leaf_2_clk),
    .RESET_B(net293),
    .D(_0236_),
    .Q_N(_3063_),
    .Q(\game.fsm.len3_block_count[0] ));
 sg13g2_dfrbp_1 \game.fsm.len3_block_count[1]$_SDFFE_PP0P_  (.CLK(clknet_leaf_2_clk),
    .RESET_B(net294),
    .D(_0237_),
    .Q_N(_3062_),
    .Q(\game.fsm.len3_block_count[1] ));
 sg13g2_dfrbp_1 \game.fsm.len3_color_count[0][0]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_42_clk),
    .RESET_B(net295),
    .D(_0238_),
    .Q_N(_3061_),
    .Q(\game.fsm.len3_color_count[0][0] ));
 sg13g2_dfrbp_1 \game.fsm.len3_color_count[0][1]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_42_clk),
    .RESET_B(net296),
    .D(_0239_),
    .Q_N(_0048_),
    .Q(\game.fsm.len3_color_count[0][1] ));
 sg13g2_dfrbp_1 \game.fsm.len3_color_count[1][0]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_43_clk),
    .RESET_B(net297),
    .D(_0240_),
    .Q_N(_3060_),
    .Q(\game.fsm.len3_color_count[1][0] ));
 sg13g2_dfrbp_1 \game.fsm.len3_color_count[1][1]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_42_clk),
    .RESET_B(net298),
    .D(_0241_),
    .Q_N(_0049_),
    .Q(\game.fsm.len3_color_count[1][1] ));
 sg13g2_dfrbp_1 \game.fsm.len3_color_count[2][0]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_42_clk),
    .RESET_B(net299),
    .D(_0242_),
    .Q_N(_3059_),
    .Q(\game.fsm.len3_color_count[2][0] ));
 sg13g2_dfrbp_1 \game.fsm.len3_color_count[2][1]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_42_clk),
    .RESET_B(net300),
    .D(_0243_),
    .Q_N(_0050_),
    .Q(\game.fsm.len3_color_count[2][1] ));
 sg13g2_dfrbp_1 \game.fsm.len3_color_count[3][0]$_DFFE_PP_  (.CLK(clknet_leaf_42_clk),
    .RESET_B(net301),
    .D(_0244_),
    .Q_N(_3058_),
    .Q(\game.fsm.len3_color_count[3][0] ));
 sg13g2_dfrbp_1 \game.fsm.len3_color_count[3][1]$_DFFE_PP_  (.CLK(clknet_leaf_43_clk),
    .RESET_B(net302),
    .D(_0245_),
    .Q_N(_0051_),
    .Q(\game.fsm.len3_color_count[3][1] ));
 sg13g2_dfrbp_1 \game.fsm.length[0]$_SDFFE_PP0P_  (.CLK(clknet_3_2__leaf_clk),
    .RESET_B(net303),
    .D(_0246_),
    .Q_N(_0066_),
    .Q(\game.fsm.length[0] ));
 sg13g2_dfrbp_1 \game.fsm.length[1]$_SDFFE_PP0P_  (.CLK(clknet_leaf_36_clk),
    .RESET_B(net304),
    .D(_0247_),
    .Q_N(_0068_),
    .Q(\game.fsm.length[1] ));
 sg13g2_dfrbp_1 \game.fsm.length[2]$_SDFFE_PP0P_  (.CLK(clknet_leaf_29_clk),
    .RESET_B(net305),
    .D(_0248_),
    .Q_N(_0067_),
    .Q(\game.fsm.length[2] ));
 sg13g2_dfrbp_1 \game.fsm.num_blocks[0]$_SDFFE_PP0P_  (.CLK(clknet_leaf_41_clk),
    .RESET_B(net306),
    .D(_0249_),
    .Q_N(_0033_),
    .Q(\game.fsm.num_blocks[0] ));
 sg13g2_dfrbp_1 \game.fsm.num_blocks[1]$_SDFFE_PP0P_  (.CLK(clknet_leaf_2_clk),
    .RESET_B(net307),
    .D(_0250_),
    .Q_N(_0073_),
    .Q(\game.fsm.num_blocks[1] ));
 sg13g2_dfrbp_1 \game.fsm.num_blocks[2]$_SDFFE_PP0P_  (.CLK(clknet_leaf_44_clk),
    .RESET_B(net308),
    .D(_0251_),
    .Q_N(_0085_),
    .Q(\game.fsm.num_blocks[2] ));
 sg13g2_dfrbp_1 \game.fsm.seq[0][0]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_35_clk),
    .RESET_B(net309),
    .D(_0252_),
    .Q_N(_0064_),
    .Q(\game.fsm.seq[0][0] ));
 sg13g2_dfrbp_1 \game.fsm.seq[0][1]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_35_clk),
    .RESET_B(net310),
    .D(_0253_),
    .Q_N(_3057_),
    .Q(\game.fsm.seq[0][1] ));
 sg13g2_dfrbp_1 \game.fsm.seq[1][0]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_35_clk),
    .RESET_B(net311),
    .D(_0254_),
    .Q_N(_0065_),
    .Q(\game.fsm.seq[1][0] ));
 sg13g2_dfrbp_1 \game.fsm.seq[1][1]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_35_clk),
    .RESET_B(net312),
    .D(_0255_),
    .Q_N(_3056_),
    .Q(\game.fsm.seq[1][1] ));
 sg13g2_dfrbp_1 \game.fsm.seq[2][0]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_34_clk),
    .RESET_B(net313),
    .D(_0256_),
    .Q_N(_3055_),
    .Q(\game.fsm.seq[2][0] ));
 sg13g2_dfrbp_1 \game.fsm.seq[2][1]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_34_clk),
    .RESET_B(net314),
    .D(_0257_),
    .Q_N(_3054_),
    .Q(\game.fsm.seq[2][1] ));
 sg13g2_dfrbp_1 \game.fsm.seq[3][0]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_34_clk),
    .RESET_B(net315),
    .D(_0258_),
    .Q_N(_3053_),
    .Q(\game.fsm.seq[3][0] ));
 sg13g2_dfrbp_1 \game.fsm.seq[3][1]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_34_clk),
    .RESET_B(net316),
    .D(_0259_),
    .Q_N(_3052_),
    .Q(\game.fsm.seq[3][1] ));
 sg13g2_dfrbp_1 \game.fsm.seq[4][0]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_35_clk),
    .RESET_B(net317),
    .D(_0260_),
    .Q_N(_3051_),
    .Q(\game.fsm.seq[4][0] ));
 sg13g2_dfrbp_1 \game.fsm.seq[4][1]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_35_clk),
    .RESET_B(net318),
    .D(_0261_),
    .Q_N(_3050_),
    .Q(\game.fsm.seq[4][1] ));
 sg13g2_dfrbp_1 \game.fsm.seq[5][0]$_DFFE_PP_  (.CLK(clknet_leaf_34_clk),
    .RESET_B(net319),
    .D(_0262_),
    .Q_N(_3049_),
    .Q(\game.fsm.seq[5][0] ));
 sg13g2_dfrbp_1 \game.fsm.seq[5][1]$_DFFE_PP_  (.CLK(clknet_leaf_34_clk),
    .RESET_B(net320),
    .D(_0263_),
    .Q_N(_3048_),
    .Q(\game.fsm.seq[5][1] ));
 sg13g2_dfrbp_1 \game.fsm.seq[6][0]$_SDFFE_PP0P_  (.CLK(clknet_leaf_35_clk),
    .RESET_B(net321),
    .D(_0264_),
    .Q_N(_3047_),
    .Q(\game.fsm.seq[6][0] ));
 sg13g2_dfrbp_1 \game.fsm.seq[6][1]$_SDFFE_PP0P_  (.CLK(clknet_leaf_35_clk),
    .RESET_B(net322),
    .D(_0265_),
    .Q_N(_3046_),
    .Q(\game.fsm.seq[6][1] ));
 sg13g2_dfrbp_1 \game.fsm.seq[7][0]$_DFFE_PP_  (.CLK(clknet_leaf_34_clk),
    .RESET_B(net323),
    .D(_0266_),
    .Q_N(_3045_),
    .Q(\game.fsm.seq[7][0] ));
 sg13g2_dfrbp_1 \game.fsm.seq[7][1]$_DFFE_PP_  (.CLK(clknet_leaf_34_clk),
    .RESET_B(net324),
    .D(_0267_),
    .Q_N(_3044_),
    .Q(\game.fsm.seq[7][1] ));
 sg13g2_dfrbp_1 \game.fsm_read_pos[0]$_SDFFE_PN0P_  (.CLK(clknet_leaf_30_clk),
    .RESET_B(net325),
    .D(_0095_),
    .Q_N(_3043_),
    .Q(\game.fsm.read_pos[0] ));
 sg13g2_dfrbp_1 \game.fsm_read_pos[1]$_SDFFE_PN0P_  (.CLK(clknet_leaf_29_clk),
    .RESET_B(net326),
    .D(_0096_),
    .Q_N(_3042_),
    .Q(\game.fsm.read_pos[1] ));
 sg13g2_dfrbp_1 \game.fsm_read_pos[2]$_SDFFE_PN0P_  (.CLK(clknet_leaf_30_clk),
    .RESET_B(net327),
    .D(_0097_),
    .Q_N(_3041_),
    .Q(\game.fsm.read_pos[2] ));
 sg13g2_dfrbp_1 \game.input_color[0]$_SDFFE_PN0P_  (.CLK(clknet_leaf_3_clk),
    .RESET_B(net328),
    .D(_0268_),
    .Q_N(_3040_),
    .Q(\game.input_color[0] ));
 sg13g2_dfrbp_1 \game.input_color[1]$_SDFFE_PN0P_  (.CLK(clknet_leaf_28_clk),
    .RESET_B(net329),
    .D(_0269_),
    .Q_N(_3039_),
    .Q(\game.input_color[1] ));
 sg13g2_dfrbp_1 \game.input_erase$_SDFF_PN0_  (.CLK(clknet_leaf_39_clk),
    .RESET_B(net330),
    .D(_0270_),
    .Q_N(_3038_),
    .Q(\game.input_erase ));
 sg13g2_dfrbp_1 \game.input_reset$_SDFF_PN1_  (.CLK(clknet_leaf_40_clk),
    .RESET_B(net331),
    .D(_0271_),
    .Q_N(_3037_),
    .Q(\game.input_reset ));
 sg13g2_dfrbp_1 \game.input_update$_SDFF_PN0_  (.CLK(clknet_leaf_40_clk),
    .RESET_B(net332),
    .D(_0272_),
    .Q_N(_0031_),
    .Q(\game.input_update ));
 sg13g2_dfrbp_1 \game.leds[0]$_SDFFE_PN0P_  (.CLK(clknet_leaf_28_clk),
    .RESET_B(net333),
    .D(_0273_),
    .Q_N(_3036_),
    .Q(net12));
 sg13g2_dfrbp_1 \game.leds[1]$_SDFFE_PN0P_  (.CLK(clknet_leaf_28_clk),
    .RESET_B(net334),
    .D(_0274_),
    .Q_N(_3035_),
    .Q(net13));
 sg13g2_dfrbp_1 \game.leds[2]$_SDFFE_PN1P_  (.CLK(clknet_leaf_18_clk),
    .RESET_B(net335),
    .D(_0275_),
    .Q_N(_3034_),
    .Q(net14));
 sg13g2_dfrbp_1 \game.leds[3]$_SDFFE_PN0P_  (.CLK(clknet_leaf_28_clk),
    .RESET_B(net336),
    .D(_0276_),
    .Q_N(_3033_),
    .Q(net15));
 sg13g2_dfrbp_1 \game.next_state[1]$_SDFFE_PN0P_  (.CLK(clknet_leaf_16_clk),
    .RESET_B(net337),
    .D(_0277_),
    .Q_N(_3032_),
    .Q(\game.next_state[0] ));
 sg13g2_dfrbp_1 \game.next_state[2]$_SDFFE_PN0P_  (.CLK(clknet_leaf_16_clk),
    .RESET_B(net338),
    .D(_0278_),
    .Q_N(_3031_),
    .Q(\game.next_state[2] ));
 sg13g2_dfrbp_1 \game.slv.fsm_color[0]$_SDFF_PP0_  (.CLK(clknet_leaf_15_clk),
    .RESET_B(net339),
    .D(_0279_),
    .Q_N(_3030_),
    .Q(\game.slv.fsm_color[0] ));
 sg13g2_dfrbp_1 \game.slv.fsm_color[1]$_SDFF_PP0_  (.CLK(clknet_leaf_4_clk),
    .RESET_B(net340),
    .D(_0280_),
    .Q_N(_3029_),
    .Q(\game.slv.fsm_color[1] ));
 sg13g2_dfrbp_1 \game.slv.fsm_reset$_SDFF_PN1_  (.CLK(clknet_leaf_4_clk),
    .RESET_B(net341),
    .D(_0281_),
    .Q_N(_3028_),
    .Q(\game.slv.fsm_reset ));
 sg13g2_dfrbp_1 \game.slv.fsm_update$_SDFF_PP0_  (.CLK(clknet_leaf_15_clk),
    .RESET_B(net342),
    .D(_0282_),
    .Q_N(_0032_),
    .Q(\game.slv.fsm_update ));
 sg13g2_dfrbp_1 \game.slv.length[0]$_SDFFE_PN0P_  (.CLK(clknet_leaf_8_clk),
    .RESET_B(net343),
    .D(_0283_),
    .Q_N(_3027_),
    .Q(\game.slv.length[0] ));
 sg13g2_dfrbp_1 \game.slv.length[1]$_SDFFE_PN0P_  (.CLK(clknet_leaf_8_clk),
    .RESET_B(net344),
    .D(_0284_),
    .Q_N(_3026_),
    .Q(\game.slv.length[1] ));
 sg13g2_dfrbp_1 \game.slv.length[2]$_SDFFE_PN0P_  (.CLK(clknet_leaf_7_clk),
    .RESET_B(net345),
    .D(_0285_),
    .Q_N(_3025_),
    .Q(\game.slv.length[2] ));
 sg13g2_dfrbp_1 \game.slv.lfsr[0]$_SDFF_PN1_  (.CLK(clknet_leaf_9_clk),
    .RESET_B(net346),
    .D(_0286_),
    .Q_N(_3024_),
    .Q(\game.slv.lfsr[0] ));
 sg13g2_dfrbp_1 \game.slv.lfsr[10]$_SDFF_PN1_  (.CLK(clknet_leaf_8_clk),
    .RESET_B(net347),
    .D(_0287_),
    .Q_N(_3023_),
    .Q(\game.slv.lfsr[10] ));
 sg13g2_dfrbp_1 \game.slv.lfsr[11]$_SDFF_PN1_  (.CLK(clknet_leaf_7_clk),
    .RESET_B(net348),
    .D(_0288_),
    .Q_N(_3022_),
    .Q(\game.slv.lfsr[11] ));
 sg13g2_dfrbp_1 \game.slv.lfsr[12]$_SDFF_PN1_  (.CLK(clknet_leaf_9_clk),
    .RESET_B(net349),
    .D(_0289_),
    .Q_N(_3021_),
    .Q(\game.slv.lfsr[12] ));
 sg13g2_dfrbp_1 \game.slv.lfsr[13]$_SDFF_PN1_  (.CLK(clknet_leaf_9_clk),
    .RESET_B(net350),
    .D(_0290_),
    .Q_N(_3020_),
    .Q(\game.slv.lfsr[13] ));
 sg13g2_dfrbp_1 \game.slv.lfsr[14]$_SDFF_PN1_  (.CLK(clknet_leaf_7_clk),
    .RESET_B(net351),
    .D(_0291_),
    .Q_N(_3019_),
    .Q(\game.slv.lfsr[14] ));
 sg13g2_dfrbp_1 \game.slv.lfsr[15]$_SDFF_PN1_  (.CLK(clknet_leaf_9_clk),
    .RESET_B(net352),
    .D(_0292_),
    .Q_N(_3018_),
    .Q(\game.slv.lfsr[15] ));
 sg13g2_dfrbp_1 \game.slv.lfsr[16]$_SDFF_PN1_  (.CLK(clknet_leaf_9_clk),
    .RESET_B(net353),
    .D(_0293_),
    .Q_N(_3017_),
    .Q(\game.slv.lfsr[16] ));
 sg13g2_dfrbp_1 \game.slv.lfsr[17]$_SDFF_PN1_  (.CLK(clknet_leaf_7_clk),
    .RESET_B(net354),
    .D(_0294_),
    .Q_N(_3016_),
    .Q(\game.slv.lfsr[17] ));
 sg13g2_dfrbp_1 \game.slv.lfsr[18]$_SDFF_PN1_  (.CLK(clknet_leaf_9_clk),
    .RESET_B(net355),
    .D(_0295_),
    .Q_N(_3015_),
    .Q(\game.slv.lfsr[18] ));
 sg13g2_dfrbp_1 \game.slv.lfsr[19]$_SDFF_PN1_  (.CLK(clknet_leaf_8_clk),
    .RESET_B(net356),
    .D(_0296_),
    .Q_N(_3014_),
    .Q(\game.slv.lfsr[19] ));
 sg13g2_dfrbp_1 \game.slv.lfsr[1]$_SDFF_PN1_  (.CLK(clknet_leaf_9_clk),
    .RESET_B(net357),
    .D(_0297_),
    .Q_N(_3013_),
    .Q(\game.slv.lfsr[1] ));
 sg13g2_dfrbp_1 \game.slv.lfsr[20]$_SDFF_PN1_  (.CLK(clknet_leaf_7_clk),
    .RESET_B(net358),
    .D(_0298_),
    .Q_N(_3012_),
    .Q(\game.slv.lfsr[20] ));
 sg13g2_dfrbp_1 \game.slv.lfsr[2]$_SDFF_PN1_  (.CLK(clknet_leaf_7_clk),
    .RESET_B(net359),
    .D(_0299_),
    .Q_N(_3011_),
    .Q(\game.slv.lfsr[2] ));
 sg13g2_dfrbp_1 \game.slv.lfsr[3]$_SDFF_PN1_  (.CLK(clknet_leaf_10_clk),
    .RESET_B(net360),
    .D(_0300_),
    .Q_N(_3010_),
    .Q(\game.slv.lfsr[3] ));
 sg13g2_dfrbp_1 \game.slv.lfsr[4]$_SDFF_PN1_  (.CLK(clknet_leaf_8_clk),
    .RESET_B(net361),
    .D(_0301_),
    .Q_N(_3009_),
    .Q(\game.slv.lfsr[4] ));
 sg13g2_dfrbp_1 \game.slv.lfsr[5]$_SDFF_PN1_  (.CLK(clknet_leaf_7_clk),
    .RESET_B(net362),
    .D(_0302_),
    .Q_N(_3008_),
    .Q(\game.slv.lfsr[5] ));
 sg13g2_dfrbp_1 \game.slv.lfsr[6]$_SDFF_PN1_  (.CLK(clknet_leaf_10_clk),
    .RESET_B(net363),
    .D(_0303_),
    .Q_N(_3007_),
    .Q(\game.slv.lfsr[6] ));
 sg13g2_dfrbp_1 \game.slv.lfsr[7]$_SDFF_PN1_  (.CLK(clknet_leaf_8_clk),
    .RESET_B(net364),
    .D(_0304_),
    .Q_N(_3006_),
    .Q(\game.slv.lfsr[7] ));
 sg13g2_dfrbp_1 \game.slv.lfsr[8]$_SDFF_PN1_  (.CLK(clknet_leaf_7_clk),
    .RESET_B(net365),
    .D(_0305_),
    .Q_N(_3005_),
    .Q(\game.slv.lfsr[8] ));
 sg13g2_dfrbp_1 \game.slv.lfsr[9]$_SDFF_PN1_  (.CLK(clknet_leaf_10_clk),
    .RESET_B(net366),
    .D(_0306_),
    .Q_N(_3004_),
    .Q(\game.slv.lfsr[9] ));
 sg13g2_dfrbp_1 \game.slv.pos[0]$_SDFFE_PN0P_  (.CLK(clknet_leaf_6_clk),
    .RESET_B(net367),
    .D(_0307_),
    .Q_N(_0056_),
    .Q(\game.slv.pos[0] ));
 sg13g2_dfrbp_1 \game.slv.pos[1]$_SDFFE_PN0P_  (.CLK(clknet_leaf_6_clk),
    .RESET_B(net368),
    .D(_0308_),
    .Q_N(_3003_),
    .Q(\game.slv.pos[1] ));
 sg13g2_dfrbp_1 \game.slv.pos[2]$_SDFFE_PN0P_  (.CLK(clknet_leaf_6_clk),
    .RESET_B(net369),
    .D(_0309_),
    .Q_N(_3002_),
    .Q(\game.slv.pos[2] ));
 sg13g2_dfrbp_1 \game.slv.ready$_SDFF_PP0_  (.CLK(clknet_leaf_4_clk),
    .RESET_B(net370),
    .D(_0310_),
    .Q_N(_3001_),
    .Q(\game.slv.ready ));
 sg13g2_dfrbp_1 \game.slv.retries[0]$_SDFFE_PN0P_  (.CLK(clknet_leaf_4_clk),
    .RESET_B(net371),
    .D(_0311_),
    .Q_N(_3000_),
    .Q(\game.slv.retries[0] ));
 sg13g2_dfrbp_1 \game.slv.retries[1]$_SDFFE_PN0P_  (.CLK(clknet_leaf_8_clk),
    .RESET_B(net372),
    .D(_0312_),
    .Q_N(_2999_),
    .Q(\game.slv.retries[1] ));
 sg13g2_dfrbp_1 \game.slv.retries[2]$_SDFFE_PN0P_  (.CLK(clknet_leaf_8_clk),
    .RESET_B(net373),
    .D(_0313_),
    .Q_N(_2998_),
    .Q(\game.slv.retries[2] ));
 sg13g2_dfrbp_1 \game.slv.saved_target$_SDFFE_PN0P_  (.CLK(clknet_leaf_4_clk),
    .RESET_B(net374),
    .D(_0314_),
    .Q_N(_3163_),
    .Q(\game.slv.saved_target ));
 sg13g2_dfrbp_1 \game.slv.state[1]$_DFF_P_  (.CLK(clknet_leaf_4_clk),
    .RESET_B(net375),
    .D(_0011_),
    .Q_N(_0030_),
    .Q(\game.slv.state[1] ));
 sg13g2_dfrbp_1 \game.slv.state[2]$_DFF_P_  (.CLK(clknet_leaf_4_clk),
    .RESET_B(net376),
    .D(_0012_),
    .Q_N(_3164_),
    .Q(\game.slv.state[2] ));
 sg13g2_dfrbp_1 \game.slv.state[3]$_DFF_P_  (.CLK(clknet_leaf_4_clk),
    .RESET_B(net377),
    .D(_0010_),
    .Q_N(_0029_),
    .Q(\game.slv.state[3] ));
 sg13g2_dfrbp_1 \game.solver_active$_SDFFE_PN0P_  (.CLK(clknet_leaf_40_clk),
    .RESET_B(net378),
    .D(_0315_),
    .Q_N(_2997_),
    .Q(\game.solver_active ));
 sg13g2_dfrbp_1 \game.solver_target[0]$_SDFFE_PN0P_  (.CLK(clknet_leaf_15_clk),
    .RESET_B(net379),
    .D(_0316_),
    .Q_N(_2996_),
    .Q(\game.slv.target[0] ));
 sg13g2_dfrbp_1 \game.solver_target[1]$_SDFFE_PN0P_  (.CLK(clknet_leaf_15_clk),
    .RESET_B(net380),
    .D(_0317_),
    .Q_N(_2995_),
    .Q(\game.slv.target[1] ));
 sg13g2_dfrbp_1 \game.solver_trigger$_SDFF_PP0_  (.CLK(clknet_3_4__leaf_clk),
    .RESET_B(net381),
    .D(_0318_),
    .Q_N(_0028_),
    .Q(\game.slv.trigger ));
 sg13g2_dfrbp_1 \game.solver_trigger_delayed$_SDFFE_PN0P_  (.CLK(clknet_leaf_16_clk),
    .RESET_B(net382),
    .D(_0319_),
    .Q_N(_2994_),
    .Q(\game.solver_trigger_delayed ));
 sg13g2_dfrbp_1 \game.sound_mode[0]$_SDFFE_PN0P_  (.CLK(clknet_leaf_27_clk),
    .RESET_B(net383),
    .D(_0320_),
    .Q_N(_2993_),
    .Q(\game.sound_mode[0] ));
 sg13g2_dfrbp_1 \game.sound_mode[1]$_SDFFE_PN0P_  (.CLK(clknet_leaf_27_clk),
    .RESET_B(net384),
    .D(_0321_),
    .Q_N(_2992_),
    .Q(\game.sound_mode[1] ));
 sg13g2_dfrbp_1 \game.sound_mode[2]$_SDFFE_PN0P_  (.CLK(clknet_leaf_27_clk),
    .RESET_B(net385),
    .D(_0322_),
    .Q_N(_0038_),
    .Q(\game.sound_mode[2] ));
 sg13g2_dfrbp_1 \game.sound_on$_SDFFE_PN1P_  (.CLK(clknet_leaf_27_clk),
    .RESET_B(net386),
    .D(_0323_),
    .Q_N(_0013_),
    .Q(\game.sound_on ));
 sg13g2_dfrbp_1 \game.state[0]$_SDFFE_PN0P_  (.CLK(clknet_leaf_17_clk),
    .RESET_B(net387),
    .D(_0324_),
    .Q_N(_2991_),
    .Q(\game.state[0] ));
 sg13g2_dfrbp_1 \game.state[1]$_SDFFE_PN0P_  (.CLK(clknet_leaf_17_clk),
    .RESET_B(net388),
    .D(_0325_),
    .Q_N(_2990_),
    .Q(\game.state[1] ));
 sg13g2_dfrbp_1 \game.state[2]$_SDFFE_PN0P_  (.CLK(clknet_leaf_17_clk),
    .RESET_B(net389),
    .D(_0326_),
    .Q_N(_2989_),
    .Q(\game.state[2] ));
 sg13g2_dfrbp_1 \game.state[3]$_SDFFE_PN0P_  (.CLK(clknet_leaf_17_clk),
    .RESET_B(net390),
    .D(_0327_),
    .Q_N(_2988_),
    .Q(\game.state[3] ));
 sg13g2_dfrbp_1 \game.tune[0]$_SDFFE_PN0P_  (.CLK(clknet_leaf_27_clk),
    .RESET_B(net391),
    .D(_0328_),
    .Q_N(_2987_),
    .Q(\game.tune[0] ));
 sg13g2_dfrbp_1 \game.tune[1]$_SDFFE_PN0P_  (.CLK(clknet_leaf_27_clk),
    .RESET_B(net392),
    .D(_0329_),
    .Q_N(_2986_),
    .Q(\game.tune[1] ));
 sg13g2_dfrbp_1 \gate_200hz$_SDFF_PN0_  (.CLK(clknet_leaf_18_clk),
    .RESET_B(net393),
    .D(_0330_),
    .Q_N(_0035_),
    .Q(\btn.gate_200hz ));
 sg13g2_dfrbp_1 \snd.active_tune[0]$_SDFFE_PN0P_  (.CLK(clknet_leaf_30_clk),
    .RESET_B(net394),
    .D(_0331_),
    .Q_N(_2985_),
    .Q(\snd.active_tune[0] ));
 sg13g2_dfrbp_1 \snd.active_tune[1]$_SDFFE_PN0P_  (.CLK(clknet_leaf_26_clk),
    .RESET_B(net395),
    .D(_0332_),
    .Q_N(_2984_),
    .Q(\snd.active_tune[1] ));
 sg13g2_dfrbp_1 \snd.chord[0][0]$_SDFFE_PN0P_  (.CLK(clknet_leaf_26_clk),
    .RESET_B(net396),
    .D(_0333_),
    .Q_N(_0057_),
    .Q(\snd.chord[0][0] ));
 sg13g2_dfrbp_1 \snd.chord[0][1]$_SDFFE_PN0P_  (.CLK(clknet_leaf_26_clk),
    .RESET_B(net397),
    .D(_0334_),
    .Q_N(_2983_),
    .Q(\snd.chord[0][1] ));
 sg13g2_dfrbp_1 \snd.chord[0][2]$_SDFFE_PN0P_  (.CLK(clknet_leaf_25_clk),
    .RESET_B(net398),
    .D(_0335_),
    .Q_N(_2982_),
    .Q(\snd.chord[0][2] ));
 sg13g2_dfrbp_1 \snd.chord[0][3]$_SDFFE_PN0P_  (.CLK(clknet_leaf_25_clk),
    .RESET_B(net399),
    .D(_0336_),
    .Q_N(_2981_),
    .Q(\snd.chord[0][3] ));
 sg13g2_dfrbp_1 \snd.chord[0][4]$_SDFFE_PN0P_  (.CLK(clknet_leaf_25_clk),
    .RESET_B(net400),
    .D(_0337_),
    .Q_N(_2980_),
    .Q(\snd.chord[0][4] ));
 sg13g2_dfrbp_1 \snd.chord[0][5]$_SDFFE_PN0P_  (.CLK(clknet_leaf_26_clk),
    .RESET_B(net401),
    .D(_0338_),
    .Q_N(_2979_),
    .Q(\snd.chord[0][5] ));
 sg13g2_dfrbp_1 \snd.chord[1][2]$_SDFFE_PN0P_  (.CLK(clknet_leaf_26_clk),
    .RESET_B(net402),
    .D(_0339_),
    .Q_N(_2978_),
    .Q(\snd.chord[1][0] ));
 sg13g2_dfrbp_1 \snd.chord[1][5]$_SDFFE_PN0P_  (.CLK(clknet_leaf_26_clk),
    .RESET_B(net403),
    .D(_0340_),
    .Q_N(_2977_),
    .Q(\snd.chord[1][5] ));
 sg13g2_dfrbp_1 \snd.chord[2][2]$_SDFFE_PN0P_  (.CLK(clknet_leaf_26_clk),
    .RESET_B(net404),
    .D(_0341_),
    .Q_N(_2976_),
    .Q(\snd.chord[2][2] ));
 sg13g2_dfrbp_1 \snd.chord[3][2]$_SDFFE_PN0P_  (.CLK(clknet_leaf_25_clk),
    .RESET_B(net405),
    .D(_0342_),
    .Q_N(_0060_),
    .Q(\snd.chord[3][0] ));
 sg13g2_dfrbp_1 \snd.counter[0]$_SDFF_PN0_  (.CLK(clknet_leaf_23_clk),
    .RESET_B(net406),
    .D(_0343_),
    .Q_N(_2975_),
    .Q(\snd.counter[0] ));
 sg13g2_dfrbp_1 \snd.counter[1]$_SDFF_PP0_  (.CLK(clknet_leaf_23_clk),
    .RESET_B(net407),
    .D(_0344_),
    .Q_N(_2974_),
    .Q(\snd.counter[1] ));
 sg13g2_dfrbp_1 \snd.counter[2]$_SDFF_PP0_  (.CLK(clknet_leaf_23_clk),
    .RESET_B(net408),
    .D(_0345_),
    .Q_N(_2973_),
    .Q(\snd.counter[2] ));
 sg13g2_dfrbp_1 \snd.counter[3]$_SDFF_PP0_  (.CLK(clknet_leaf_22_clk),
    .RESET_B(net409),
    .D(_0346_),
    .Q_N(_2972_),
    .Q(\snd.counter[3] ));
 sg13g2_dfrbp_1 \snd.counter[4]$_SDFF_PP0_  (.CLK(clknet_leaf_22_clk),
    .RESET_B(net410),
    .D(_0347_),
    .Q_N(_2971_),
    .Q(\snd.counter[4] ));
 sg13g2_dfrbp_1 \snd.counter[5]$_SDFF_PP0_  (.CLK(clknet_leaf_22_clk),
    .RESET_B(net411),
    .D(_0348_),
    .Q_N(_2970_),
    .Q(\snd.counter[5] ));
 sg13g2_dfrbp_1 \snd.counter[6]$_SDFF_PP0_  (.CLK(clknet_leaf_22_clk),
    .RESET_B(net412),
    .D(_0349_),
    .Q_N(_2969_),
    .Q(\snd.counter[6] ));
 sg13g2_dfrbp_1 \snd.counter[7]$_SDFF_PP0_  (.CLK(clknet_leaf_22_clk),
    .RESET_B(net413),
    .D(_0350_),
    .Q_N(_2968_),
    .Q(\snd.counter[7] ));
 sg13g2_dfrbp_1 \snd.counter[8]$_SDFF_PP0_  (.CLK(clknet_leaf_22_clk),
    .RESET_B(net414),
    .D(_0351_),
    .Q_N(_0036_),
    .Q(\snd.counter[8] ));
 sg13g2_dfrbp_1 \snd.next_note_sel[0]$_SDFFE_PN0P_  (.CLK(clknet_leaf_27_clk),
    .RESET_B(net415),
    .D(_0352_),
    .Q_N(_2967_),
    .Q(\snd.next_note_sel[0] ));
 sg13g2_dfrbp_1 \snd.next_note_sel[1]$_SDFFE_PN0P_  (.CLK(clknet_leaf_26_clk),
    .RESET_B(net416),
    .D(_0353_),
    .Q_N(_2966_),
    .Q(\snd.next_note_sel[1] ));
 sg13g2_dfrbp_1 \snd.next_note_timing[0]$_SDFFE_PN0P_  (.CLK(clknet_leaf_23_clk),
    .RESET_B(net417),
    .D(_0354_),
    .Q_N(_2965_),
    .Q(\snd.next_note_timing[0] ));
 sg13g2_dfrbp_1 \snd.next_note_timing[1]$_SDFFE_PN0P_  (.CLK(clknet_leaf_24_clk),
    .RESET_B(net418),
    .D(_0355_),
    .Q_N(_2964_),
    .Q(\snd.next_note_timing[1] ));
 sg13g2_dfrbp_1 \snd.next_note_timing[2]$_SDFFE_PN0P_  (.CLK(clknet_leaf_24_clk),
    .RESET_B(net419),
    .D(_0356_),
    .Q_N(_2963_),
    .Q(\snd.next_note_timing[2] ));
 sg13g2_dfrbp_1 \snd.next_note_timing[3]$_SDFFE_PN0P_  (.CLK(clknet_leaf_24_clk),
    .RESET_B(net420),
    .D(_0357_),
    .Q_N(_2962_),
    .Q(\snd.next_note_timing[3] ));
 sg13g2_dfrbp_1 \snd.next_note_timing[4]$_SDFFE_PN0P_  (.CLK(clknet_leaf_21_clk),
    .RESET_B(net421),
    .D(_0358_),
    .Q_N(_2961_),
    .Q(\snd.next_note_timing[4] ));
 sg13g2_dfrbp_1 \snd.next_note_timing[5]$_SDFFE_PN0P_  (.CLK(clknet_leaf_24_clk),
    .RESET_B(net422),
    .D(_0359_),
    .Q_N(_2960_),
    .Q(\snd.next_note_timing[5] ));
 sg13g2_dfrbp_1 \snd.next_note_timing[6]$_SDFFE_PN0P_  (.CLK(clknet_leaf_24_clk),
    .RESET_B(net423),
    .D(_0360_),
    .Q_N(_2959_),
    .Q(\snd.next_note_timing[6] ));
 sg13g2_dfrbp_1 \snd.next_note_timing[7]$_SDFFE_PN0P_  (.CLK(clknet_leaf_21_clk),
    .RESET_B(net424),
    .D(_0361_),
    .Q_N(_2958_),
    .Q(\snd.next_note_timing[7] ));
 sg13g2_dfrbp_1 \snd.next_note_timing[8]$_SDFFE_PN0P_  (.CLK(clknet_leaf_21_clk),
    .RESET_B(net425),
    .D(_0362_),
    .Q_N(_2957_),
    .Q(\snd.next_note_timing[8] ));
 sg13g2_dfrbp_1 \snd.note_sel[0]$_SDFFE_PN0P_  (.CLK(clknet_leaf_25_clk),
    .RESET_B(net426),
    .D(_0363_),
    .Q_N(_2956_),
    .Q(\snd.note_sel[0] ));
 sg13g2_dfrbp_1 \snd.note_sel[1]$_SDFFE_PN0P_  (.CLK(clknet_leaf_25_clk),
    .RESET_B(net427),
    .D(_0364_),
    .Q_N(_2955_),
    .Q(\snd.note_sel[1] ));
 sg13g2_dfrbp_1 \snd.note_timing[0]$_SDFFE_PN0P_  (.CLK(clknet_leaf_24_clk),
    .RESET_B(net428),
    .D(_0365_),
    .Q_N(_2954_),
    .Q(\snd.note_timing[0] ));
 sg13g2_dfrbp_1 \snd.note_timing[1]$_SDFFE_PN0P_  (.CLK(clknet_leaf_25_clk),
    .RESET_B(net429),
    .D(_0366_),
    .Q_N(_2953_),
    .Q(\snd.note_timing[1] ));
 sg13g2_dfrbp_1 \snd.note_timing[2]$_SDFFE_PN0P_  (.CLK(clknet_leaf_23_clk),
    .RESET_B(net430),
    .D(_0367_),
    .Q_N(_2952_),
    .Q(\snd.note_timing[2] ));
 sg13g2_dfrbp_1 \snd.note_timing[3]$_SDFFE_PN0P_  (.CLK(clknet_leaf_23_clk),
    .RESET_B(net431),
    .D(_0368_),
    .Q_N(_2951_),
    .Q(\snd.note_timing[3] ));
 sg13g2_dfrbp_1 \snd.note_timing[4]$_SDFFE_PN0P_  (.CLK(clknet_leaf_23_clk),
    .RESET_B(net432),
    .D(_0369_),
    .Q_N(_2950_),
    .Q(\snd.note_timing[4] ));
 sg13g2_dfrbp_1 \snd.note_timing[5]$_SDFFE_PN0P_  (.CLK(clknet_leaf_24_clk),
    .RESET_B(net433),
    .D(_0370_),
    .Q_N(_2949_),
    .Q(\snd.note_timing[5] ));
 sg13g2_dfrbp_1 \snd.note_timing[6]$_SDFFE_PN0P_  (.CLK(clknet_leaf_23_clk),
    .RESET_B(net434),
    .D(_0371_),
    .Q_N(_2948_),
    .Q(\snd.note_timing[6] ));
 sg13g2_dfrbp_1 \snd.note_timing[7]$_SDFFE_PN0P_  (.CLK(clknet_leaf_21_clk),
    .RESET_B(net435),
    .D(_0372_),
    .Q_N(_2947_),
    .Q(\snd.note_timing[7] ));
 sg13g2_dfrbp_1 \snd.note_timing[8]$_SDFFE_PN0P_  (.CLK(clknet_leaf_21_clk),
    .RESET_B(net436),
    .D(_0373_),
    .Q_N(_2946_),
    .Q(\snd.note_timing[8] ));
 sg13g2_dfrbp_1 \snd.sequencer_state[0]$_SDFFE_PN0P_  (.CLK(clknet_leaf_29_clk),
    .RESET_B(net437),
    .D(_0374_),
    .Q_N(_2945_),
    .Q(\snd.sequencer_state[0] ));
 sg13g2_dfrbp_1 \snd.sequencer_state[1]$_SDFFE_PN0P_  (.CLK(clknet_leaf_29_clk),
    .RESET_B(net438),
    .D(_0375_),
    .Q_N(_2944_),
    .Q(\snd.sequencer_state[1] ));
 sg13g2_dfrbp_1 \snd.sound$_SDFFE_PP0P_  (.CLK(clknet_leaf_22_clk),
    .RESET_B(net439),
    .D(_0376_),
    .Q_N(_2943_),
    .Q(\snd.sound ));
 sg13g2_dfrbp_1 \snd.tune_counter[0]$_SDFFE_PN0P_  (.CLK(clknet_leaf_32_clk),
    .RESET_B(net440),
    .D(_0377_),
    .Q_N(_2942_),
    .Q(\snd.tune_counter[0] ));
 sg13g2_dfrbp_1 \snd.tune_counter[1]$_SDFFE_PN0P_  (.CLK(clknet_leaf_31_clk),
    .RESET_B(net441),
    .D(_0378_),
    .Q_N(_2941_),
    .Q(\snd.tune_counter[1] ));
 sg13g2_dfrbp_1 \snd.tune_counter[2]$_SDFFE_PN0P_  (.CLK(clknet_leaf_32_clk),
    .RESET_B(net442),
    .D(_0379_),
    .Q_N(_2940_),
    .Q(\snd.tune_counter[2] ));
 sg13g2_dfrbp_1 \snd.tune_counter[3]$_SDFFE_PN0P_  (.CLK(clknet_leaf_31_clk),
    .RESET_B(net443),
    .D(_0380_),
    .Q_N(_2939_),
    .Q(\snd.tune_counter[3] ));
 sg13g2_dfrbp_1 \snd.tune_counter[4]$_SDFFE_PN0P_  (.CLK(clknet_leaf_31_clk),
    .RESET_B(net444),
    .D(_0381_),
    .Q_N(_2938_),
    .Q(\snd.tune_counter[4] ));
 sg13g2_dfrbp_1 \snd.tune_counter[5]$_SDFFE_PN0P_  (.CLK(clknet_leaf_31_clk),
    .RESET_B(net445),
    .D(_0382_),
    .Q_N(_2937_),
    .Q(\snd.tune_counter[5] ));
 sg13g2_dfrbp_1 \snd.tune_counter[6]$_SDFFE_PN0P_  (.CLK(clknet_leaf_31_clk),
    .RESET_B(net446),
    .D(_0383_),
    .Q_N(_0037_),
    .Q(\snd.tune_counter[6] ));
 sg13g2_dfrbp_1 \snd.tune_pos[0]$_SDFFE_PN0P_  (.CLK(clknet_leaf_31_clk),
    .RESET_B(net447),
    .D(_0384_),
    .Q_N(_2936_),
    .Q(\snd.tune_pos[0] ));
 sg13g2_dfrbp_1 \snd.tune_pos[1]$_SDFFE_PN0P_  (.CLK(clknet_leaf_31_clk),
    .RESET_B(net448),
    .D(_0385_),
    .Q_N(_2935_),
    .Q(\snd.tune_pos[1] ));
 sg13g2_dfrbp_1 \snd.tune_pos[2]$_SDFFE_PN0P_  (.CLK(clknet_leaf_31_clk),
    .RESET_B(net449),
    .D(_0386_),
    .Q_N(_0039_),
    .Q(\snd.tune_pos[2] ));
 sg13g2_buf_1 input1 (.A(ui_in[0]),
    .X(net1));
 sg13g2_buf_1 input2 (.A(ui_in[1]),
    .X(net2));
 sg13g2_buf_1 input3 (.A(ui_in[2]),
    .X(net3));
 sg13g2_buf_1 input4 (.A(ui_in[3]),
    .X(net4));
 sg13g2_buf_1 output5 (.A(net5),
    .X(uio_out[0]));
 sg13g2_buf_1 output6 (.A(net6),
    .X(uio_out[1]));
 sg13g2_buf_1 output7 (.A(net7),
    .X(uio_out[2]));
 sg13g2_buf_1 output8 (.A(net8),
    .X(uio_out[3]));
 sg13g2_buf_1 output9 (.A(net9),
    .X(uio_out[4]));
 sg13g2_buf_1 output10 (.A(net10),
    .X(uio_out[5]));
 sg13g2_buf_1 output11 (.A(net11),
    .X(uio_out[6]));
 sg13g2_buf_1 output12 (.A(net12),
    .X(uo_out[0]));
 sg13g2_buf_1 output13 (.A(net13),
    .X(uo_out[1]));
 sg13g2_buf_1 output14 (.A(net14),
    .X(uo_out[2]));
 sg13g2_buf_1 output15 (.A(net15),
    .X(uo_out[3]));
 sg13g2_buf_1 output16 (.A(net16),
    .X(uo_out[4]));
 sg13g2_buf_1 output17 (.A(net17),
    .X(uo_out[5]));
 sg13g2_buf_1 output18 (.A(net18),
    .X(uo_out[6]));
 sg13g2_buf_2 fanout19 (.A(_1570_),
    .X(net19));
 sg13g2_buf_2 fanout20 (.A(_2423_),
    .X(net20));
 sg13g2_buf_2 fanout21 (.A(_0921_),
    .X(net21));
 sg13g2_buf_2 fanout22 (.A(_1178_),
    .X(net22));
 sg13g2_buf_2 fanout23 (.A(_0967_),
    .X(net23));
 sg13g2_buf_2 fanout24 (.A(_0929_),
    .X(net24));
 sg13g2_buf_2 fanout25 (.A(_1980_),
    .X(net25));
 sg13g2_buf_2 fanout26 (.A(_1245_),
    .X(net26));
 sg13g2_buf_2 fanout27 (.A(_1932_),
    .X(net27));
 sg13g2_buf_2 fanout28 (.A(_1043_),
    .X(net28));
 sg13g2_buf_4 fanout29 (.X(net29),
    .A(_1015_));
 sg13g2_buf_2 fanout30 (.A(_0877_),
    .X(net30));
 sg13g2_buf_2 fanout31 (.A(_1437_),
    .X(net31));
 sg13g2_buf_2 fanout32 (.A(_1255_),
    .X(net32));
 sg13g2_buf_2 fanout33 (.A(_1214_),
    .X(net33));
 sg13g2_buf_2 fanout34 (.A(_1148_),
    .X(net34));
 sg13g2_buf_2 fanout35 (.A(_1132_),
    .X(net35));
 sg13g2_buf_2 fanout36 (.A(_1107_),
    .X(net36));
 sg13g2_buf_2 fanout37 (.A(_1061_),
    .X(net37));
 sg13g2_buf_2 fanout38 (.A(_1058_),
    .X(net38));
 sg13g2_buf_2 fanout39 (.A(_1036_),
    .X(net39));
 sg13g2_buf_2 fanout40 (.A(_0949_),
    .X(net40));
 sg13g2_buf_2 fanout41 (.A(_0736_),
    .X(net41));
 sg13g2_buf_2 fanout42 (.A(_2673_),
    .X(net42));
 sg13g2_buf_2 fanout43 (.A(_1693_),
    .X(net43));
 sg13g2_buf_2 fanout44 (.A(_1620_),
    .X(net44));
 sg13g2_buf_2 fanout45 (.A(_1057_),
    .X(net45));
 sg13g2_buf_2 fanout46 (.A(_1052_),
    .X(net46));
 sg13g2_buf_2 fanout47 (.A(_0933_),
    .X(net47));
 sg13g2_buf_2 fanout48 (.A(_1040_),
    .X(net48));
 sg13g2_buf_2 fanout49 (.A(_0699_),
    .X(net49));
 sg13g2_buf_2 fanout50 (.A(_0402_),
    .X(net50));
 sg13g2_buf_2 fanout51 (.A(_2541_),
    .X(net51));
 sg13g2_buf_2 fanout52 (.A(_2389_),
    .X(net52));
 sg13g2_buf_2 fanout53 (.A(_2190_),
    .X(net53));
 sg13g2_buf_2 fanout54 (.A(_2147_),
    .X(net54));
 sg13g2_buf_2 fanout55 (.A(_2033_),
    .X(net55));
 sg13g2_buf_2 fanout56 (.A(_1956_),
    .X(net56));
 sg13g2_buf_2 fanout57 (.A(_1827_),
    .X(net57));
 sg13g2_buf_2 fanout58 (.A(_1756_),
    .X(net58));
 sg13g2_buf_2 fanout59 (.A(_1754_),
    .X(net59));
 sg13g2_buf_2 fanout60 (.A(_1672_),
    .X(net60));
 sg13g2_buf_2 fanout61 (.A(_1668_),
    .X(net61));
 sg13g2_buf_2 fanout62 (.A(_1666_),
    .X(net62));
 sg13g2_buf_2 fanout63 (.A(_1418_),
    .X(net63));
 sg13g2_buf_2 fanout64 (.A(_1079_),
    .X(net64));
 sg13g2_buf_2 fanout65 (.A(_1012_),
    .X(net65));
 sg13g2_buf_2 fanout66 (.A(_0988_),
    .X(net66));
 sg13g2_buf_2 fanout67 (.A(_0974_),
    .X(net67));
 sg13g2_buf_2 fanout68 (.A(_0667_),
    .X(net68));
 sg13g2_buf_2 fanout69 (.A(_0466_),
    .X(net69));
 sg13g2_buf_2 fanout70 (.A(_0411_),
    .X(net70));
 sg13g2_buf_2 fanout71 (.A(_0397_),
    .X(net71));
 sg13g2_buf_2 fanout72 (.A(_2925_),
    .X(net72));
 sg13g2_buf_2 fanout73 (.A(_2643_),
    .X(net73));
 sg13g2_buf_2 fanout74 (.A(_2398_),
    .X(net74));
 sg13g2_buf_2 fanout75 (.A(_2017_),
    .X(net75));
 sg13g2_buf_2 fanout76 (.A(_1927_),
    .X(net76));
 sg13g2_buf_2 fanout77 (.A(_1925_),
    .X(net77));
 sg13g2_buf_2 fanout78 (.A(_1880_),
    .X(net78));
 sg13g2_buf_2 fanout79 (.A(_1874_),
    .X(net79));
 sg13g2_buf_2 fanout80 (.A(_1870_),
    .X(net80));
 sg13g2_buf_2 fanout81 (.A(_1861_),
    .X(net81));
 sg13g2_buf_2 fanout82 (.A(_1856_),
    .X(net82));
 sg13g2_buf_2 fanout83 (.A(_1854_),
    .X(net83));
 sg13g2_buf_2 fanout84 (.A(_1795_),
    .X(net84));
 sg13g2_buf_2 fanout85 (.A(_1783_),
    .X(net85));
 sg13g2_buf_2 fanout86 (.A(_1781_),
    .X(net86));
 sg13g2_buf_2 fanout87 (.A(_1665_),
    .X(net87));
 sg13g2_buf_2 fanout88 (.A(_1660_),
    .X(net88));
 sg13g2_buf_2 fanout89 (.A(_1525_),
    .X(net89));
 sg13g2_buf_2 fanout90 (.A(_1524_),
    .X(net90));
 sg13g2_buf_2 fanout91 (.A(_1510_),
    .X(net91));
 sg13g2_buf_2 fanout92 (.A(_1417_),
    .X(net92));
 sg13g2_buf_2 fanout93 (.A(_1017_),
    .X(net93));
 sg13g2_buf_2 fanout94 (.A(_0973_),
    .X(net94));
 sg13g2_buf_2 fanout95 (.A(_0971_),
    .X(net95));
 sg13g2_buf_2 fanout96 (.A(_0922_),
    .X(net96));
 sg13g2_buf_2 fanout97 (.A(_0542_),
    .X(net97));
 sg13g2_buf_2 fanout98 (.A(_0540_),
    .X(net98));
 sg13g2_buf_2 fanout99 (.A(_0501_),
    .X(net99));
 sg13g2_buf_2 fanout100 (.A(_0496_),
    .X(net100));
 sg13g2_buf_2 fanout101 (.A(_0437_),
    .X(net101));
 sg13g2_buf_2 fanout102 (.A(_0399_),
    .X(net102));
 sg13g2_buf_2 fanout103 (.A(_0394_),
    .X(net103));
 sg13g2_buf_2 fanout104 (.A(_0388_),
    .X(net104));
 sg13g2_buf_2 fanout105 (.A(_2795_),
    .X(net105));
 sg13g2_buf_2 fanout106 (.A(_2726_),
    .X(net106));
 sg13g2_buf_2 fanout107 (.A(_2688_),
    .X(net107));
 sg13g2_buf_2 fanout108 (.A(_2642_),
    .X(net108));
 sg13g2_buf_2 fanout109 (.A(_2321_),
    .X(net109));
 sg13g2_buf_2 fanout110 (.A(_2316_),
    .X(net110));
 sg13g2_buf_2 fanout111 (.A(_2297_),
    .X(net111));
 sg13g2_buf_2 fanout112 (.A(_2213_),
    .X(net112));
 sg13g2_buf_2 fanout113 (.A(_2212_),
    .X(net113));
 sg13g2_buf_2 fanout114 (.A(_1920_),
    .X(net114));
 sg13g2_buf_2 fanout115 (.A(_1643_),
    .X(net115));
 sg13g2_buf_2 fanout116 (.A(_0945_),
    .X(net116));
 sg13g2_buf_2 fanout117 (.A(_0884_),
    .X(net117));
 sg13g2_buf_2 fanout118 (.A(_0872_),
    .X(net118));
 sg13g2_buf_2 fanout119 (.A(_0863_),
    .X(net119));
 sg13g2_buf_2 fanout120 (.A(_0862_),
    .X(net120));
 sg13g2_buf_2 fanout121 (.A(_0858_),
    .X(net121));
 sg13g2_buf_2 fanout122 (.A(_0571_),
    .X(net122));
 sg13g2_buf_2 fanout123 (.A(_0547_),
    .X(net123));
 sg13g2_buf_2 fanout124 (.A(_0545_),
    .X(net124));
 sg13g2_buf_2 fanout125 (.A(_0498_),
    .X(net125));
 sg13g2_buf_2 fanout126 (.A(_0413_),
    .X(net126));
 sg13g2_buf_2 fanout127 (.A(_2930_),
    .X(net127));
 sg13g2_buf_2 fanout128 (.A(_2923_),
    .X(net128));
 sg13g2_buf_2 fanout129 (.A(_2800_),
    .X(net129));
 sg13g2_buf_2 fanout130 (.A(_2728_),
    .X(net130));
 sg13g2_buf_2 fanout131 (.A(_2700_),
    .X(net131));
 sg13g2_buf_2 fanout132 (.A(_2686_),
    .X(net132));
 sg13g2_buf_2 fanout133 (.A(_2652_),
    .X(net133));
 sg13g2_buf_2 fanout134 (.A(_2644_),
    .X(net134));
 sg13g2_tielo _6046__135 (.L_LO(net135));
 sg13g2_tielo _6048__136 (.L_LO(net136));
 sg13g2_tiehi _6027__138 (.L_HI(net138));
 sg13g2_tiehi _6028__139 (.L_HI(net139));
 sg13g2_tiehi _6029__140 (.L_HI(net140));
 sg13g2_tiehi _6030__141 (.L_HI(net141));
 sg13g2_tiehi _6031__142 (.L_HI(net142));
 sg13g2_tiehi _6032__143 (.L_HI(net143));
 sg13g2_tiehi _6033__144 (.L_HI(net144));
 sg13g2_tiehi _6034__145 (.L_HI(net145));
 sg13g2_tiehi _6035__146 (.L_HI(net146));
 sg13g2_tiehi _6038__147 (.L_HI(net147));
 sg13g2_tiehi _6039__148 (.L_HI(net148));
 sg13g2_tiehi _6040__149 (.L_HI(net149));
 sg13g2_tiehi _6041__150 (.L_HI(net150));
 sg13g2_tiehi _6042__151 (.L_HI(net151));
 sg13g2_tiehi _6043__152 (.L_HI(net152));
 sg13g2_tiehi _6044__153 (.L_HI(net153));
 sg13g2_tiehi _6045__154 (.L_HI(net154));
 sg13g2_tiehi \btn.button_state[0]$_SDFFE_PN0P__155  (.L_HI(net155));
 sg13g2_tiehi \btn.button_state[1]$_SDFFE_PN0P__156  (.L_HI(net156));
 sg13g2_tiehi \btn.button_state[2]$_SDFFE_PN0P__157  (.L_HI(net157));
 sg13g2_tiehi \btn.button_state[3]$_SDFFE_PN0P__158  (.L_HI(net158));
 sg13g2_tiehi \btn.change_timer[0]$_SDFFE_PN0P__159  (.L_HI(net159));
 sg13g2_tiehi \btn.change_timer[1]$_SDFFE_PN0P__160  (.L_HI(net160));
 sg13g2_tiehi \btn.change_timer[2]$_SDFFE_PN0P__161  (.L_HI(net161));
 sg13g2_tiehi \btn.change_timer[3]$_SDFFE_PN0P__162  (.L_HI(net162));
 sg13g2_tiehi \btn.change_timer[4]$_SDFFE_PN0P__163  (.L_HI(net163));
 sg13g2_tiehi \btn.change_timer[5]$_SDFFE_PN0P__164  (.L_HI(net164));
 sg13g2_tiehi \btn.change_timer[6]$_SDFFE_PN0P__165  (.L_HI(net165));
 sg13g2_tiehi \btn.current_event[0]$_SDFFE_PN0P__166  (.L_HI(net166));
 sg13g2_tiehi \btn.current_event[1]$_SDFFE_PN0P__167  (.L_HI(net167));
 sg13g2_tiehi \btn.current_event[2]$_SDFFE_PN0P__168  (.L_HI(net168));
 sg13g2_tiehi \btn.current_event[3]$_SDFFE_PN0P__169  (.L_HI(net169));
 sg13g2_tiehi \btn.input_event[0]$_SDFF_PN0__170  (.L_HI(net170));
 sg13g2_tiehi \btn.input_event[1]$_SDFF_PN0__171  (.L_HI(net171));
 sg13g2_tiehi \btn.input_event[2]$_SDFF_PN0__172  (.L_HI(net172));
 sg13g2_tiehi \btn.input_event[3]$_SDFF_PN0__173  (.L_HI(net173));
 sg13g2_tiehi \btn.input_event[4]$_SDFF_PN0__174  (.L_HI(net174));
 sg13g2_tiehi \btn.long_press$_SDFFE_PN0P__175  (.L_HI(net175));
 sg13g2_tiehi \btn.sample_10ms[0]$_SDFFE_PN0P__176  (.L_HI(net176));
 sg13g2_tiehi \btn.sample_10ms[1]$_SDFFE_PN0P__177  (.L_HI(net177));
 sg13g2_tiehi \btn.sample_10ms[2]$_SDFFE_PN0P__178  (.L_HI(net178));
 sg13g2_tiehi \btn.sample_10ms[3]$_SDFFE_PN0P__179  (.L_HI(net179));
 sg13g2_tiehi \btn.sample_15ms[0]$_SDFFE_PN0P__180  (.L_HI(net180));
 sg13g2_tiehi \btn.sample_15ms[1]$_SDFFE_PN0P__181  (.L_HI(net181));
 sg13g2_tiehi \btn.sample_15ms[2]$_SDFFE_PN0P__182  (.L_HI(net182));
 sg13g2_tiehi \btn.sample_15ms[3]$_SDFFE_PN0P__183  (.L_HI(net183));
 sg13g2_tiehi \btn.sample_5ms[0]$_SDFFE_PN0P__184  (.L_HI(net184));
 sg13g2_tiehi \btn.sample_5ms[1]$_SDFFE_PN0P__185  (.L_HI(net185));
 sg13g2_tiehi \btn.sample_5ms[2]$_SDFFE_PN0P__186  (.L_HI(net186));
 sg13g2_tiehi \btn.sample_5ms[3]$_SDFFE_PN0P__187  (.L_HI(net187));
 sg13g2_tiehi \clk_div_counter[0]$_SDFF_PP0__188  (.L_HI(net188));
 sg13g2_tiehi \clk_div_counter[1]$_SDFF_PP0__189  (.L_HI(net189));
 sg13g2_tiehi \clk_div_counter[2]$_SDFF_PP0__190  (.L_HI(net190));
 sg13g2_tiehi \clk_div_counter[3]$_SDFF_PP0__191  (.L_HI(net191));
 sg13g2_tiehi \clk_div_counter[4]$_SDFF_PP0__192  (.L_HI(net192));
 sg13g2_tiehi \clk_div_counter[5]$_SDFF_PP0__193  (.L_HI(net193));
 sg13g2_tiehi \clk_div_counter[6]$_SDFF_PP0__194  (.L_HI(net194));
 sg13g2_tiehi \clk_div_counter[7]$_SDFF_PP0__195  (.L_HI(net195));
 sg13g2_tiehi \dsp.digit_sel_raw[0]$_SDFF_PN0__196  (.L_HI(net196));
 sg13g2_tiehi \dsp.digit_sel_raw[1]$_SDFF_PN0__197  (.L_HI(net197));
 sg13g2_tiehi \dsp.segments_raw[0]$_SDFF_PN0__198  (.L_HI(net198));
 sg13g2_tiehi \dsp.segments_raw[1]$_SDFF_PN0__199  (.L_HI(net199));
 sg13g2_tiehi \dsp.segments_raw[2]$_SDFF_PN0__200  (.L_HI(net200));
 sg13g2_tiehi \dsp.segments_raw[3]$_SDFF_PN0__201  (.L_HI(net201));
 sg13g2_tiehi \dsp.segments_raw[4]$_SDFF_PN0__202  (.L_HI(net202));
 sg13g2_tiehi \dsp.segments_raw[5]$_SDFF_PN0__203  (.L_HI(net203));
 sg13g2_tiehi \dsp.segments_raw[6]$_SDFF_PN0__204  (.L_HI(net204));
 sg13g2_tiehi \game.challenge_mode$_SDFFE_PN0P__205  (.L_HI(net205));
 sg13g2_tiehi \game.challenge_num[0]$_SDFFE_PN0P__206  (.L_HI(net206));
 sg13g2_tiehi \game.challenge_num[1]$_SDFFE_PN0P__207  (.L_HI(net207));
 sg13g2_tiehi \game.challenge_num[2]$_SDFFE_PN0P__208  (.L_HI(net208));
 sg13g2_tiehi \game.challenge_num[3]$_SDFFE_PN0P__209  (.L_HI(net209));
 sg13g2_tiehi \game.counter[0]$_SDFFE_PN0P__210  (.L_HI(net210));
 sg13g2_tiehi \game.counter[1]$_SDFFE_PN0P__211  (.L_HI(net211));
 sg13g2_tiehi \game.counter[2]$_SDFFE_PN0P__212  (.L_HI(net212));
 sg13g2_tiehi \game.counter[3]$_SDFFE_PN0P__213  (.L_HI(net213));
 sg13g2_tiehi \game.counter[4]$_SDFFE_PN0P__214  (.L_HI(net214));
 sg13g2_tiehi \game.counter[5]$_SDFFE_PN0P__215  (.L_HI(net215));
 sg13g2_tiehi \game.counter[6]$_SDFFE_PN0P__216  (.L_HI(net216));
 sg13g2_tiehi \game.counter[7]$_SDFFE_PN0P__217  (.L_HI(net217));
 sg13g2_tiehi \game.current_level[0]$_SDFFE_PN0P__218  (.L_HI(net218));
 sg13g2_tiehi \game.current_level[1]$_SDFFE_PN0P__219  (.L_HI(net219));
 sg13g2_tiehi \game.current_level[2]$_SDFFE_PN0P__220  (.L_HI(net220));
 sg13g2_tiehi \game.current_level[3]$_SDFFE_PN0P__221  (.L_HI(net221));
 sg13g2_tiehi \game.current_level[4]$_SDFFE_PN0P__222  (.L_HI(net222));
 sg13g2_tiehi \game.display_graphical$_SDFFE_PN0P__223  (.L_HI(net223));
 sg13g2_tiehi \game.display_value[0]$_SDFFE_PN1P__224  (.L_HI(net224));
 sg13g2_tiehi \game.display_value[1]$_SDFFE_PN0P__225  (.L_HI(net225));
 sg13g2_tiehi \game.display_value[2]$_SDFFE_PN0P__226  (.L_HI(net226));
 sg13g2_tiehi \game.display_value[3]$_SDFFE_PN0P__227  (.L_HI(net227));
 sg13g2_tiehi \game.display_value[4]$_SDFFE_PN0P__228  (.L_HI(net228));
 sg13g2_tiehi \game.fsm.block_len[0][0]$_SDFFCE_PN0P__229  (.L_HI(net229));
 sg13g2_tiehi \game.fsm.block_len[0][1]$_SDFFCE_PN0P__230  (.L_HI(net230));
 sg13g2_tiehi \game.fsm.block_len[0][2]$_SDFFCE_PN0P__231  (.L_HI(net231));
 sg13g2_tiehi \game.fsm.block_len[1][0]$_SDFFCE_PN0P__232  (.L_HI(net232));
 sg13g2_tiehi \game.fsm.block_len[1][1]$_SDFFCE_PN0P__233  (.L_HI(net233));
 sg13g2_tiehi \game.fsm.block_len[1][2]$_SDFFCE_PN0P__234  (.L_HI(net234));
 sg13g2_tiehi \game.fsm.block_len[2][0]$_SDFFCE_PN0P__235  (.L_HI(net235));
 sg13g2_tiehi \game.fsm.block_len[2][1]$_SDFFCE_PN0P__236  (.L_HI(net236));
 sg13g2_tiehi \game.fsm.block_len[2][2]$_SDFFCE_PN0P__237  (.L_HI(net237));
 sg13g2_tiehi \game.fsm.block_len[3][0]$_SDFFCE_PN0P__238  (.L_HI(net238));
 sg13g2_tiehi \game.fsm.block_len[3][1]$_SDFFCE_PN0P__239  (.L_HI(net239));
 sg13g2_tiehi \game.fsm.block_len[3][2]$_SDFFCE_PN0P__240  (.L_HI(net240));
 sg13g2_tiehi \game.fsm.block_len[4][0]$_SDFFCE_PN0P__241  (.L_HI(net241));
 sg13g2_tiehi \game.fsm.block_len[4][1]$_SDFFCE_PN0P__242  (.L_HI(net242));
 sg13g2_tiehi \game.fsm.block_len[4][2]$_SDFFCE_PN0P__243  (.L_HI(net243));
 sg13g2_tiehi \game.fsm.block_len[5][0]$_DFFE_PP__244  (.L_HI(net244));
 sg13g2_tiehi \game.fsm.block_len[5][1]$_DFFE_PP__245  (.L_HI(net245));
 sg13g2_tiehi \game.fsm.block_len[5][2]$_DFFE_PP__246  (.L_HI(net246));
 sg13g2_tiehi \game.fsm.block_len[6][0]$_SDFFE_PP0P__247  (.L_HI(net247));
 sg13g2_tiehi \game.fsm.block_len[6][1]$_SDFFE_PP0P__248  (.L_HI(net248));
 sg13g2_tiehi \game.fsm.block_len[6][2]$_SDFFE_PP0P__249  (.L_HI(net249));
 sg13g2_tiehi \game.fsm.block_len[7][0]$_DFFE_PP__250  (.L_HI(net250));
 sg13g2_tiehi \game.fsm.block_len[7][1]$_DFFE_PP__251  (.L_HI(net251));
 sg13g2_tiehi \game.fsm.block_len[7][2]$_DFFE_PP__252  (.L_HI(net252));
 sg13g2_tiehi \game.fsm.color_count[0][0]$_SDFFCE_PN0P__253  (.L_HI(net253));
 sg13g2_tiehi \game.fsm.color_count[0][1]$_SDFFCE_PN0P__254  (.L_HI(net254));
 sg13g2_tiehi \game.fsm.color_count[0][2]$_SDFFCE_PN0P__255  (.L_HI(net255));
 sg13g2_tiehi \game.fsm.color_count[1][0]$_SDFFCE_PN0P__256  (.L_HI(net256));
 sg13g2_tiehi \game.fsm.color_count[1][1]$_SDFFCE_PN0P__257  (.L_HI(net257));
 sg13g2_tiehi \game.fsm.color_count[1][2]$_SDFFCE_PN0P__258  (.L_HI(net258));
 sg13g2_tiehi \game.fsm.color_count[2][0]$_SDFFCE_PN0P__259  (.L_HI(net259));
 sg13g2_tiehi \game.fsm.color_count[2][1]$_SDFFCE_PN0P__260  (.L_HI(net260));
 sg13g2_tiehi \game.fsm.color_count[2][2]$_SDFFCE_PN0P__261  (.L_HI(net261));
 sg13g2_tiehi \game.fsm.color_count[3][0]$_DFFE_PP__262  (.L_HI(net262));
 sg13g2_tiehi \game.fsm.color_count[3][1]$_DFFE_PP__263  (.L_HI(net263));
 sg13g2_tiehi \game.fsm.color_count[3][2]$_DFFE_PP__264  (.L_HI(net264));
 sg13g2_tiehi \game.fsm.green_block_count[0]$_SDFFE_PP0P__265  (.L_HI(net265));
 sg13g2_tiehi \game.fsm.green_block_count[1]$_SDFFE_PP0P__266  (.L_HI(net266));
 sg13g2_tiehi \game.fsm.green_block_count[2]$_SDFFE_PP0P__267  (.L_HI(net267));
 sg13g2_tiehi \game.fsm.len1_block_count[0]$_SDFFE_PP0P__268  (.L_HI(net268));
 sg13g2_tiehi \game.fsm.len1_block_count[1]$_SDFFE_PP0P__269  (.L_HI(net269));
 sg13g2_tiehi \game.fsm.len1_block_count[2]$_SDFFE_PP0P__270  (.L_HI(net270));
 sg13g2_tiehi \game.fsm.len1_color_count[0][0]$_SDFFCE_PN0P__271  (.L_HI(net271));
 sg13g2_tiehi \game.fsm.len1_color_count[0][1]$_SDFFCE_PN0P__272  (.L_HI(net272));
 sg13g2_tiehi \game.fsm.len1_color_count[0][2]$_SDFFCE_PN0P__273  (.L_HI(net273));
 sg13g2_tiehi \game.fsm.len1_color_count[1][0]$_SDFFCE_PN0P__274  (.L_HI(net274));
 sg13g2_tiehi \game.fsm.len1_color_count[1][1]$_SDFFCE_PN0P__275  (.L_HI(net275));
 sg13g2_tiehi \game.fsm.len1_color_count[1][2]$_SDFFCE_PN0P__276  (.L_HI(net276));
 sg13g2_tiehi \game.fsm.len1_color_count[2][0]$_SDFFCE_PN0P__277  (.L_HI(net277));
 sg13g2_tiehi \game.fsm.len1_color_count[2][1]$_SDFFCE_PN0P__278  (.L_HI(net278));
 sg13g2_tiehi \game.fsm.len1_color_count[2][2]$_SDFFCE_PN0P__279  (.L_HI(net279));
 sg13g2_tiehi \game.fsm.len1_color_count[3][0]$_DFFE_PP__280  (.L_HI(net280));
 sg13g2_tiehi \game.fsm.len1_color_count[3][1]$_DFFE_PP__281  (.L_HI(net281));
 sg13g2_tiehi \game.fsm.len1_color_count[3][2]$_DFFE_PP__282  (.L_HI(net282));
 sg13g2_tiehi \game.fsm.len2_block_count[0]$_SDFFE_PP0P__283  (.L_HI(net283));
 sg13g2_tiehi \game.fsm.len2_block_count[1]$_SDFFE_PP0P__284  (.L_HI(net284));
 sg13g2_tiehi \game.fsm.len2_color_count[0][0]$_SDFFCE_PN0P__285  (.L_HI(net285));
 sg13g2_tiehi \game.fsm.len2_color_count[0][1]$_SDFFCE_PN0P__286  (.L_HI(net286));
 sg13g2_tiehi \game.fsm.len2_color_count[1][0]$_SDFFCE_PN0P__287  (.L_HI(net287));
 sg13g2_tiehi \game.fsm.len2_color_count[1][1]$_SDFFCE_PN0P__288  (.L_HI(net288));
 sg13g2_tiehi \game.fsm.len2_color_count[2][0]$_SDFFCE_PN0P__289  (.L_HI(net289));
 sg13g2_tiehi \game.fsm.len2_color_count[2][1]$_SDFFCE_PN0P__290  (.L_HI(net290));
 sg13g2_tiehi \game.fsm.len2_color_count[3][0]$_DFFE_PP__291  (.L_HI(net291));
 sg13g2_tiehi \game.fsm.len2_color_count[3][1]$_DFFE_PP__292  (.L_HI(net292));
 sg13g2_tiehi \game.fsm.len3_block_count[0]$_SDFFE_PP0P__293  (.L_HI(net293));
 sg13g2_tiehi \game.fsm.len3_block_count[1]$_SDFFE_PP0P__294  (.L_HI(net294));
 sg13g2_tiehi \game.fsm.len3_color_count[0][0]$_SDFFCE_PN0P__295  (.L_HI(net295));
 sg13g2_tiehi \game.fsm.len3_color_count[0][1]$_SDFFCE_PN0P__296  (.L_HI(net296));
 sg13g2_tiehi \game.fsm.len3_color_count[1][0]$_SDFFCE_PN0P__297  (.L_HI(net297));
 sg13g2_tiehi \game.fsm.len3_color_count[1][1]$_SDFFCE_PN0P__298  (.L_HI(net298));
 sg13g2_tiehi \game.fsm.len3_color_count[2][0]$_SDFFCE_PN0P__299  (.L_HI(net299));
 sg13g2_tiehi \game.fsm.len3_color_count[2][1]$_SDFFCE_PN0P__300  (.L_HI(net300));
 sg13g2_tiehi \game.fsm.len3_color_count[3][0]$_DFFE_PP__301  (.L_HI(net301));
 sg13g2_tiehi \game.fsm.len3_color_count[3][1]$_DFFE_PP__302  (.L_HI(net302));
 sg13g2_tiehi \game.fsm.length[0]$_SDFFE_PP0P__303  (.L_HI(net303));
 sg13g2_tiehi \game.fsm.length[1]$_SDFFE_PP0P__304  (.L_HI(net304));
 sg13g2_tiehi \game.fsm.length[2]$_SDFFE_PP0P__305  (.L_HI(net305));
 sg13g2_tiehi \game.fsm.num_blocks[0]$_SDFFE_PP0P__306  (.L_HI(net306));
 sg13g2_tiehi \game.fsm.num_blocks[1]$_SDFFE_PP0P__307  (.L_HI(net307));
 sg13g2_tiehi \game.fsm.num_blocks[2]$_SDFFE_PP0P__308  (.L_HI(net308));
 sg13g2_tiehi \game.fsm.seq[0][0]$_SDFFCE_PN0P__309  (.L_HI(net309));
 sg13g2_tiehi \game.fsm.seq[0][1]$_SDFFCE_PN0P__310  (.L_HI(net310));
 sg13g2_tiehi \game.fsm.seq[1][0]$_SDFFCE_PN0P__311  (.L_HI(net311));
 sg13g2_tiehi \game.fsm.seq[1][1]$_SDFFCE_PN0P__312  (.L_HI(net312));
 sg13g2_tiehi \game.fsm.seq[2][0]$_SDFFCE_PN0P__313  (.L_HI(net313));
 sg13g2_tiehi \game.fsm.seq[2][1]$_SDFFCE_PN0P__314  (.L_HI(net314));
 sg13g2_tiehi \game.fsm.seq[3][0]$_SDFFCE_PN0P__315  (.L_HI(net315));
 sg13g2_tiehi \game.fsm.seq[3][1]$_SDFFCE_PN0P__316  (.L_HI(net316));
 sg13g2_tiehi \game.fsm.seq[4][0]$_SDFFCE_PN0P__317  (.L_HI(net317));
 sg13g2_tiehi \game.fsm.seq[4][1]$_SDFFCE_PN0P__318  (.L_HI(net318));
 sg13g2_tiehi \game.fsm.seq[5][0]$_DFFE_PP__319  (.L_HI(net319));
 sg13g2_tiehi \game.fsm.seq[5][1]$_DFFE_PP__320  (.L_HI(net320));
 sg13g2_tiehi \game.fsm.seq[6][0]$_SDFFE_PP0P__321  (.L_HI(net321));
 sg13g2_tiehi \game.fsm.seq[6][1]$_SDFFE_PP0P__322  (.L_HI(net322));
 sg13g2_tiehi \game.fsm.seq[7][0]$_DFFE_PP__323  (.L_HI(net323));
 sg13g2_tiehi \game.fsm.seq[7][1]$_DFFE_PP__324  (.L_HI(net324));
 sg13g2_tiehi \game.fsm_read_pos[0]$_SDFFE_PN0P__325  (.L_HI(net325));
 sg13g2_tiehi \game.fsm_read_pos[1]$_SDFFE_PN0P__326  (.L_HI(net326));
 sg13g2_tiehi \game.fsm_read_pos[2]$_SDFFE_PN0P__327  (.L_HI(net327));
 sg13g2_tiehi \game.input_color[0]$_SDFFE_PN0P__328  (.L_HI(net328));
 sg13g2_tiehi \game.input_color[1]$_SDFFE_PN0P__329  (.L_HI(net329));
 sg13g2_tiehi \game.input_erase$_SDFF_PN0__330  (.L_HI(net330));
 sg13g2_tiehi \game.input_reset$_SDFF_PN1__331  (.L_HI(net331));
 sg13g2_tiehi \game.input_update$_SDFF_PN0__332  (.L_HI(net332));
 sg13g2_tiehi \game.leds[0]$_SDFFE_PN0P__333  (.L_HI(net333));
 sg13g2_tiehi \game.leds[1]$_SDFFE_PN0P__334  (.L_HI(net334));
 sg13g2_tiehi \game.leds[2]$_SDFFE_PN1P__335  (.L_HI(net335));
 sg13g2_tiehi \game.leds[3]$_SDFFE_PN0P__336  (.L_HI(net336));
 sg13g2_tiehi \game.next_state[1]$_SDFFE_PN0P__337  (.L_HI(net337));
 sg13g2_tiehi \game.next_state[2]$_SDFFE_PN0P__338  (.L_HI(net338));
 sg13g2_tiehi \game.slv.fsm_color[0]$_SDFF_PP0__339  (.L_HI(net339));
 sg13g2_tiehi \game.slv.fsm_color[1]$_SDFF_PP0__340  (.L_HI(net340));
 sg13g2_tiehi \game.slv.fsm_reset$_SDFF_PN1__341  (.L_HI(net341));
 sg13g2_tiehi \game.slv.fsm_update$_SDFF_PP0__342  (.L_HI(net342));
 sg13g2_tiehi \game.slv.length[0]$_SDFFE_PN0P__343  (.L_HI(net343));
 sg13g2_tiehi \game.slv.length[1]$_SDFFE_PN0P__344  (.L_HI(net344));
 sg13g2_tiehi \game.slv.length[2]$_SDFFE_PN0P__345  (.L_HI(net345));
 sg13g2_tiehi \game.slv.lfsr[0]$_SDFF_PN1__346  (.L_HI(net346));
 sg13g2_tiehi \game.slv.lfsr[10]$_SDFF_PN1__347  (.L_HI(net347));
 sg13g2_tiehi \game.slv.lfsr[11]$_SDFF_PN1__348  (.L_HI(net348));
 sg13g2_tiehi \game.slv.lfsr[12]$_SDFF_PN1__349  (.L_HI(net349));
 sg13g2_tiehi \game.slv.lfsr[13]$_SDFF_PN1__350  (.L_HI(net350));
 sg13g2_tiehi \game.slv.lfsr[14]$_SDFF_PN1__351  (.L_HI(net351));
 sg13g2_tiehi \game.slv.lfsr[15]$_SDFF_PN1__352  (.L_HI(net352));
 sg13g2_tiehi \game.slv.lfsr[16]$_SDFF_PN1__353  (.L_HI(net353));
 sg13g2_tiehi \game.slv.lfsr[17]$_SDFF_PN1__354  (.L_HI(net354));
 sg13g2_tiehi \game.slv.lfsr[18]$_SDFF_PN1__355  (.L_HI(net355));
 sg13g2_tiehi \game.slv.lfsr[19]$_SDFF_PN1__356  (.L_HI(net356));
 sg13g2_tiehi \game.slv.lfsr[1]$_SDFF_PN1__357  (.L_HI(net357));
 sg13g2_tiehi \game.slv.lfsr[20]$_SDFF_PN1__358  (.L_HI(net358));
 sg13g2_tiehi \game.slv.lfsr[2]$_SDFF_PN1__359  (.L_HI(net359));
 sg13g2_tiehi \game.slv.lfsr[3]$_SDFF_PN1__360  (.L_HI(net360));
 sg13g2_tiehi \game.slv.lfsr[4]$_SDFF_PN1__361  (.L_HI(net361));
 sg13g2_tiehi \game.slv.lfsr[5]$_SDFF_PN1__362  (.L_HI(net362));
 sg13g2_tiehi \game.slv.lfsr[6]$_SDFF_PN1__363  (.L_HI(net363));
 sg13g2_tiehi \game.slv.lfsr[7]$_SDFF_PN1__364  (.L_HI(net364));
 sg13g2_tiehi \game.slv.lfsr[8]$_SDFF_PN1__365  (.L_HI(net365));
 sg13g2_tiehi \game.slv.lfsr[9]$_SDFF_PN1__366  (.L_HI(net366));
 sg13g2_tiehi \game.slv.pos[0]$_SDFFE_PN0P__367  (.L_HI(net367));
 sg13g2_tiehi \game.slv.pos[1]$_SDFFE_PN0P__368  (.L_HI(net368));
 sg13g2_tiehi \game.slv.pos[2]$_SDFFE_PN0P__369  (.L_HI(net369));
 sg13g2_tiehi \game.slv.ready$_SDFF_PP0__370  (.L_HI(net370));
 sg13g2_tiehi \game.slv.retries[0]$_SDFFE_PN0P__371  (.L_HI(net371));
 sg13g2_tiehi \game.slv.retries[1]$_SDFFE_PN0P__372  (.L_HI(net372));
 sg13g2_tiehi \game.slv.retries[2]$_SDFFE_PN0P__373  (.L_HI(net373));
 sg13g2_tiehi \game.slv.saved_target$_SDFFE_PN0P__374  (.L_HI(net374));
 sg13g2_tiehi \game.slv.state[1]$_DFF_P__375  (.L_HI(net375));
 sg13g2_tiehi \game.slv.state[2]$_DFF_P__376  (.L_HI(net376));
 sg13g2_tiehi \game.slv.state[3]$_DFF_P__377  (.L_HI(net377));
 sg13g2_tiehi \game.solver_active$_SDFFE_PN0P__378  (.L_HI(net378));
 sg13g2_tiehi \game.solver_target[0]$_SDFFE_PN0P__379  (.L_HI(net379));
 sg13g2_tiehi \game.solver_target[1]$_SDFFE_PN0P__380  (.L_HI(net380));
 sg13g2_tiehi \game.solver_trigger$_SDFF_PP0__381  (.L_HI(net381));
 sg13g2_tiehi \game.solver_trigger_delayed$_SDFFE_PN0P__382  (.L_HI(net382));
 sg13g2_tiehi \game.sound_mode[0]$_SDFFE_PN0P__383  (.L_HI(net383));
 sg13g2_tiehi \game.sound_mode[1]$_SDFFE_PN0P__384  (.L_HI(net384));
 sg13g2_tiehi \game.sound_mode[2]$_SDFFE_PN0P__385  (.L_HI(net385));
 sg13g2_tiehi \game.sound_on$_SDFFE_PN1P__386  (.L_HI(net386));
 sg13g2_tiehi \game.state[0]$_SDFFE_PN0P__387  (.L_HI(net387));
 sg13g2_tiehi \game.state[1]$_SDFFE_PN0P__388  (.L_HI(net388));
 sg13g2_tiehi \game.state[2]$_SDFFE_PN0P__389  (.L_HI(net389));
 sg13g2_tiehi \game.state[3]$_SDFFE_PN0P__390  (.L_HI(net390));
 sg13g2_tiehi \game.tune[0]$_SDFFE_PN0P__391  (.L_HI(net391));
 sg13g2_tiehi \game.tune[1]$_SDFFE_PN0P__392  (.L_HI(net392));
 sg13g2_tiehi \gate_200hz$_SDFF_PN0__393  (.L_HI(net393));
 sg13g2_tiehi \snd.active_tune[0]$_SDFFE_PN0P__394  (.L_HI(net394));
 sg13g2_tiehi \snd.active_tune[1]$_SDFFE_PN0P__395  (.L_HI(net395));
 sg13g2_tiehi \snd.chord[0][0]$_SDFFE_PN0P__396  (.L_HI(net396));
 sg13g2_tiehi \snd.chord[0][1]$_SDFFE_PN0P__397  (.L_HI(net397));
 sg13g2_tiehi \snd.chord[0][2]$_SDFFE_PN0P__398  (.L_HI(net398));
 sg13g2_tiehi \snd.chord[0][3]$_SDFFE_PN0P__399  (.L_HI(net399));
 sg13g2_tiehi \snd.chord[0][4]$_SDFFE_PN0P__400  (.L_HI(net400));
 sg13g2_tiehi \snd.chord[0][5]$_SDFFE_PN0P__401  (.L_HI(net401));
 sg13g2_tiehi \snd.chord[1][2]$_SDFFE_PN0P__402  (.L_HI(net402));
 sg13g2_tiehi \snd.chord[1][5]$_SDFFE_PN0P__403  (.L_HI(net403));
 sg13g2_tiehi \snd.chord[2][2]$_SDFFE_PN0P__404  (.L_HI(net404));
 sg13g2_tiehi \snd.chord[3][2]$_SDFFE_PN0P__405  (.L_HI(net405));
 sg13g2_tiehi \snd.counter[0]$_SDFF_PN0__406  (.L_HI(net406));
 sg13g2_tiehi \snd.counter[1]$_SDFF_PP0__407  (.L_HI(net407));
 sg13g2_tiehi \snd.counter[2]$_SDFF_PP0__408  (.L_HI(net408));
 sg13g2_tiehi \snd.counter[3]$_SDFF_PP0__409  (.L_HI(net409));
 sg13g2_tiehi \snd.counter[4]$_SDFF_PP0__410  (.L_HI(net410));
 sg13g2_tiehi \snd.counter[5]$_SDFF_PP0__411  (.L_HI(net411));
 sg13g2_tiehi \snd.counter[6]$_SDFF_PP0__412  (.L_HI(net412));
 sg13g2_tiehi \snd.counter[7]$_SDFF_PP0__413  (.L_HI(net413));
 sg13g2_tiehi \snd.counter[8]$_SDFF_PP0__414  (.L_HI(net414));
 sg13g2_tiehi \snd.next_note_sel[0]$_SDFFE_PN0P__415  (.L_HI(net415));
 sg13g2_tiehi \snd.next_note_sel[1]$_SDFFE_PN0P__416  (.L_HI(net416));
 sg13g2_tiehi \snd.next_note_timing[0]$_SDFFE_PN0P__417  (.L_HI(net417));
 sg13g2_tiehi \snd.next_note_timing[1]$_SDFFE_PN0P__418  (.L_HI(net418));
 sg13g2_tiehi \snd.next_note_timing[2]$_SDFFE_PN0P__419  (.L_HI(net419));
 sg13g2_tiehi \snd.next_note_timing[3]$_SDFFE_PN0P__420  (.L_HI(net420));
 sg13g2_tiehi \snd.next_note_timing[4]$_SDFFE_PN0P__421  (.L_HI(net421));
 sg13g2_tiehi \snd.next_note_timing[5]$_SDFFE_PN0P__422  (.L_HI(net422));
 sg13g2_tiehi \snd.next_note_timing[6]$_SDFFE_PN0P__423  (.L_HI(net423));
 sg13g2_tiehi \snd.next_note_timing[7]$_SDFFE_PN0P__424  (.L_HI(net424));
 sg13g2_tiehi \snd.next_note_timing[8]$_SDFFE_PN0P__425  (.L_HI(net425));
 sg13g2_tiehi \snd.note_sel[0]$_SDFFE_PN0P__426  (.L_HI(net426));
 sg13g2_tiehi \snd.note_sel[1]$_SDFFE_PN0P__427  (.L_HI(net427));
 sg13g2_tiehi \snd.note_timing[0]$_SDFFE_PN0P__428  (.L_HI(net428));
 sg13g2_tiehi \snd.note_timing[1]$_SDFFE_PN0P__429  (.L_HI(net429));
 sg13g2_tiehi \snd.note_timing[2]$_SDFFE_PN0P__430  (.L_HI(net430));
 sg13g2_tiehi \snd.note_timing[3]$_SDFFE_PN0P__431  (.L_HI(net431));
 sg13g2_tiehi \snd.note_timing[4]$_SDFFE_PN0P__432  (.L_HI(net432));
 sg13g2_tiehi \snd.note_timing[5]$_SDFFE_PN0P__433  (.L_HI(net433));
 sg13g2_tiehi \snd.note_timing[6]$_SDFFE_PN0P__434  (.L_HI(net434));
 sg13g2_tiehi \snd.note_timing[7]$_SDFFE_PN0P__435  (.L_HI(net435));
 sg13g2_tiehi \snd.note_timing[8]$_SDFFE_PN0P__436  (.L_HI(net436));
 sg13g2_tiehi \snd.sequencer_state[0]$_SDFFE_PN0P__437  (.L_HI(net437));
 sg13g2_tiehi \snd.sequencer_state[1]$_SDFFE_PN0P__438  (.L_HI(net438));
 sg13g2_tiehi \snd.sound$_SDFFE_PP0P__439  (.L_HI(net439));
 sg13g2_tiehi \snd.tune_counter[0]$_SDFFE_PN0P__440  (.L_HI(net440));
 sg13g2_tiehi \snd.tune_counter[1]$_SDFFE_PN0P__441  (.L_HI(net441));
 sg13g2_tiehi \snd.tune_counter[2]$_SDFFE_PN0P__442  (.L_HI(net442));
 sg13g2_tiehi \snd.tune_counter[3]$_SDFFE_PN0P__443  (.L_HI(net443));
 sg13g2_tiehi \snd.tune_counter[4]$_SDFFE_PN0P__444  (.L_HI(net444));
 sg13g2_tiehi \snd.tune_counter[5]$_SDFFE_PN0P__445  (.L_HI(net445));
 sg13g2_tiehi \snd.tune_counter[6]$_SDFFE_PN0P__446  (.L_HI(net446));
 sg13g2_tiehi \snd.tune_pos[0]$_SDFFE_PN0P__447  (.L_HI(net447));
 sg13g2_tiehi \snd.tune_pos[1]$_SDFFE_PN0P__448  (.L_HI(net448));
 sg13g2_tiehi \snd.tune_pos[2]$_SDFFE_PN0P__449  (.L_HI(net449));
 sg13g2_buf_2 clkbuf_leaf_1_clk (.A(clknet_3_1__leaf_clk),
    .X(clknet_leaf_1_clk));
 sg13g2_buf_2 clkbuf_leaf_2_clk (.A(clknet_3_1__leaf_clk),
    .X(clknet_leaf_2_clk));
 sg13g2_buf_2 clkbuf_leaf_3_clk (.A(clknet_3_1__leaf_clk),
    .X(clknet_leaf_3_clk));
 sg13g2_buf_2 clkbuf_leaf_4_clk (.A(clknet_3_4__leaf_clk),
    .X(clknet_leaf_4_clk));
 sg13g2_buf_2 clkbuf_leaf_6_clk (.A(clknet_3_4__leaf_clk),
    .X(clknet_leaf_6_clk));
 sg13g2_buf_2 clkbuf_leaf_7_clk (.A(clknet_3_4__leaf_clk),
    .X(clknet_leaf_7_clk));
 sg13g2_buf_2 clkbuf_leaf_8_clk (.A(clknet_3_4__leaf_clk),
    .X(clknet_leaf_8_clk));
 sg13g2_buf_2 clkbuf_leaf_9_clk (.A(clknet_3_5__leaf_clk),
    .X(clknet_leaf_9_clk));
 sg13g2_buf_2 clkbuf_leaf_10_clk (.A(clknet_3_5__leaf_clk),
    .X(clknet_leaf_10_clk));
 sg13g2_buf_2 clkbuf_leaf_11_clk (.A(clknet_3_5__leaf_clk),
    .X(clknet_leaf_11_clk));
 sg13g2_buf_2 clkbuf_leaf_12_clk (.A(clknet_3_5__leaf_clk),
    .X(clknet_leaf_12_clk));
 sg13g2_buf_2 clkbuf_leaf_13_clk (.A(clknet_3_5__leaf_clk),
    .X(clknet_leaf_13_clk));
 sg13g2_buf_2 clkbuf_leaf_14_clk (.A(clknet_3_5__leaf_clk),
    .X(clknet_leaf_14_clk));
 sg13g2_buf_2 clkbuf_leaf_15_clk (.A(clknet_3_4__leaf_clk),
    .X(clknet_leaf_15_clk));
 sg13g2_buf_2 clkbuf_leaf_16_clk (.A(clknet_3_1__leaf_clk),
    .X(clknet_leaf_16_clk));
 sg13g2_buf_2 clkbuf_leaf_17_clk (.A(clknet_3_6__leaf_clk),
    .X(clknet_leaf_17_clk));
 sg13g2_buf_2 clkbuf_leaf_18_clk (.A(clknet_3_7__leaf_clk),
    .X(clknet_leaf_18_clk));
 sg13g2_buf_2 clkbuf_leaf_19_clk (.A(clknet_3_7__leaf_clk),
    .X(clknet_leaf_19_clk));
 sg13g2_buf_2 clkbuf_leaf_20_clk (.A(clknet_3_6__leaf_clk),
    .X(clknet_leaf_20_clk));
 sg13g2_buf_2 clkbuf_leaf_21_clk (.A(clknet_3_7__leaf_clk),
    .X(clknet_leaf_21_clk));
 sg13g2_buf_2 clkbuf_leaf_22_clk (.A(clknet_3_7__leaf_clk),
    .X(clknet_leaf_22_clk));
 sg13g2_buf_2 clkbuf_leaf_23_clk (.A(clknet_3_7__leaf_clk),
    .X(clknet_leaf_23_clk));
 sg13g2_buf_2 clkbuf_leaf_24_clk (.A(clknet_3_6__leaf_clk),
    .X(clknet_leaf_24_clk));
 sg13g2_buf_2 clkbuf_leaf_25_clk (.A(clknet_3_6__leaf_clk),
    .X(clknet_leaf_25_clk));
 sg13g2_buf_2 clkbuf_leaf_26_clk (.A(clknet_3_6__leaf_clk),
    .X(clknet_leaf_26_clk));
 sg13g2_buf_2 clkbuf_leaf_27_clk (.A(clknet_3_6__leaf_clk),
    .X(clknet_leaf_27_clk));
 sg13g2_buf_2 clkbuf_leaf_28_clk (.A(clknet_3_3__leaf_clk),
    .X(clknet_leaf_28_clk));
 sg13g2_buf_2 clkbuf_leaf_29_clk (.A(clknet_3_3__leaf_clk),
    .X(clknet_leaf_29_clk));
 sg13g2_buf_2 clkbuf_leaf_30_clk (.A(clknet_3_3__leaf_clk),
    .X(clknet_leaf_30_clk));
 sg13g2_buf_2 clkbuf_leaf_31_clk (.A(clknet_3_3__leaf_clk),
    .X(clknet_leaf_31_clk));
 sg13g2_buf_2 clkbuf_leaf_32_clk (.A(clknet_3_2__leaf_clk),
    .X(clknet_leaf_32_clk));
 sg13g2_buf_2 clkbuf_leaf_34_clk (.A(clknet_3_2__leaf_clk),
    .X(clknet_leaf_34_clk));
 sg13g2_buf_2 clkbuf_leaf_35_clk (.A(clknet_3_2__leaf_clk),
    .X(clknet_leaf_35_clk));
 sg13g2_buf_2 clkbuf_leaf_36_clk (.A(clknet_3_2__leaf_clk),
    .X(clknet_leaf_36_clk));
 sg13g2_buf_2 clkbuf_leaf_37_clk (.A(clknet_3_2__leaf_clk),
    .X(clknet_leaf_37_clk));
 sg13g2_buf_2 clkbuf_leaf_38_clk (.A(clknet_3_0__leaf_clk),
    .X(clknet_leaf_38_clk));
 sg13g2_buf_2 clkbuf_leaf_39_clk (.A(clknet_3_3__leaf_clk),
    .X(clknet_leaf_39_clk));
 sg13g2_buf_2 clkbuf_leaf_40_clk (.A(clknet_3_1__leaf_clk),
    .X(clknet_leaf_40_clk));
 sg13g2_buf_2 clkbuf_leaf_41_clk (.A(clknet_3_1__leaf_clk),
    .X(clknet_leaf_41_clk));
 sg13g2_buf_2 clkbuf_leaf_42_clk (.A(clknet_3_0__leaf_clk),
    .X(clknet_leaf_42_clk));
 sg13g2_buf_2 clkbuf_leaf_43_clk (.A(clknet_3_0__leaf_clk),
    .X(clknet_leaf_43_clk));
 sg13g2_buf_2 clkbuf_leaf_44_clk (.A(clknet_3_0__leaf_clk),
    .X(clknet_leaf_44_clk));
 sg13g2_buf_2 clkbuf_leaf_45_clk (.A(clknet_3_0__leaf_clk),
    .X(clknet_leaf_45_clk));
 sg13g2_buf_1 clkbuf_0_clk (.A(clk),
    .X(clknet_0_clk));
 sg13g2_buf_1 clkbuf_3_0__f_clk (.A(clknet_0_clk),
    .X(clknet_3_0__leaf_clk));
 sg13g2_buf_1 clkbuf_3_1__f_clk (.A(clknet_0_clk),
    .X(clknet_3_1__leaf_clk));
 sg13g2_buf_1 clkbuf_3_2__f_clk (.A(clknet_0_clk),
    .X(clknet_3_2__leaf_clk));
 sg13g2_buf_1 clkbuf_3_3__f_clk (.A(clknet_0_clk),
    .X(clknet_3_3__leaf_clk));
 sg13g2_buf_1 clkbuf_3_4__f_clk (.A(clknet_0_clk),
    .X(clknet_3_4__leaf_clk));
 sg13g2_buf_1 clkbuf_3_5__f_clk (.A(clknet_0_clk),
    .X(clknet_3_5__leaf_clk));
 sg13g2_buf_1 clkbuf_3_6__f_clk (.A(clknet_0_clk),
    .X(clknet_3_6__leaf_clk));
 sg13g2_buf_1 clkbuf_3_7__f_clk (.A(clknet_0_clk),
    .X(clknet_3_7__leaf_clk));
 sg13g2_buf_1 clkload0 (.A(clknet_3_0__leaf_clk));
 sg13g2_buf_1 clkload1 (.A(clknet_3_1__leaf_clk));
 sg13g2_inv_1 clkload2 (.A(clknet_3_3__leaf_clk));
 sg13g2_buf_1 clkload3 (.A(clknet_3_5__leaf_clk));
 sg13g2_buf_1 clkload4 (.A(clknet_3_6__leaf_clk));
 sg13g2_inv_1 clkload5 (.A(clknet_3_7__leaf_clk));
 sg13g2_inv_1 clkload6 (.A(clknet_leaf_0_clk));
 sg13g2_inv_1 clkload7 (.A(clknet_leaf_38_clk));
 sg13g2_inv_1 clkload8 (.A(clknet_leaf_43_clk));
 sg13g2_inv_4 clkload9 (.A(clknet_leaf_44_clk));
 sg13g2_inv_4 clkload10 (.A(clknet_leaf_1_clk));
 sg13g2_buf_16 clkload11 (.A(clknet_leaf_2_clk));
 sg13g2_inv_2 clkload12 (.A(clknet_leaf_3_clk));
 sg13g2_inv_4 clkload13 (.A(clknet_leaf_16_clk));
 sg13g2_buf_16 clkload14 (.A(clknet_leaf_41_clk));
 sg13g2_buf_16 clkload15 (.A(clknet_leaf_32_clk));
 sg13g2_inv_1 clkload16 (.A(clknet_leaf_36_clk));
 sg13g2_buf_8 clkload17 (.A(clknet_leaf_28_clk));
 sg13g2_inv_4 clkload18 (.A(clknet_leaf_30_clk));
 sg13g2_buf_8 clkload19 (.A(clknet_leaf_12_clk));
 sg13g2_inv_1 clkload20 (.A(clknet_leaf_14_clk));
 sg13g2_inv_1 clkload21 (.A(clknet_leaf_25_clk));
 sg13g2_buf_8 clkload22 (.A(clknet_leaf_18_clk));
 sg13g2_buf_1 fanout1 (.A(_2631_),
    .X(net450));
 sg13g2_antennanp ANTENNA_1 (.A(clk));
 sg13g2_antennanp ANTENNA_2 (.A(clk));
 sg13g2_antennanp ANTENNA_3 (.A(clk));
 sg13g2_antennanp ANTENNA_4 (.A(clk));
 sg13g2_antennanp ANTENNA_5 (.A(clk));
 sg13g2_decap_8 FILLER_0_0 ();
 sg13g2_decap_8 FILLER_0_7 ();
 sg13g2_decap_8 FILLER_0_14 ();
 sg13g2_decap_8 FILLER_0_21 ();
 sg13g2_decap_8 FILLER_0_32 ();
 sg13g2_decap_4 FILLER_0_39 ();
 sg13g2_fill_1 FILLER_0_43 ();
 sg13g2_decap_8 FILLER_0_49 ();
 sg13g2_decap_8 FILLER_0_56 ();
 sg13g2_decap_8 FILLER_0_63 ();
 sg13g2_decap_8 FILLER_0_70 ();
 sg13g2_decap_8 FILLER_0_77 ();
 sg13g2_decap_8 FILLER_0_84 ();
 sg13g2_decap_8 FILLER_0_91 ();
 sg13g2_decap_8 FILLER_0_98 ();
 sg13g2_decap_8 FILLER_0_105 ();
 sg13g2_decap_8 FILLER_0_112 ();
 sg13g2_decap_8 FILLER_0_119 ();
 sg13g2_decap_8 FILLER_0_126 ();
 sg13g2_decap_4 FILLER_0_133 ();
 sg13g2_fill_2 FILLER_0_137 ();
 sg13g2_decap_8 FILLER_0_143 ();
 sg13g2_decap_8 FILLER_0_150 ();
 sg13g2_decap_8 FILLER_0_157 ();
 sg13g2_decap_8 FILLER_0_164 ();
 sg13g2_decap_8 FILLER_0_171 ();
 sg13g2_decap_8 FILLER_0_178 ();
 sg13g2_decap_8 FILLER_0_185 ();
 sg13g2_decap_8 FILLER_0_192 ();
 sg13g2_decap_8 FILLER_0_199 ();
 sg13g2_decap_8 FILLER_0_210 ();
 sg13g2_decap_8 FILLER_0_217 ();
 sg13g2_decap_8 FILLER_0_224 ();
 sg13g2_decap_8 FILLER_0_231 ();
 sg13g2_decap_8 FILLER_0_238 ();
 sg13g2_decap_8 FILLER_0_245 ();
 sg13g2_decap_8 FILLER_0_252 ();
 sg13g2_decap_8 FILLER_0_259 ();
 sg13g2_decap_4 FILLER_0_266 ();
 sg13g2_decap_8 FILLER_0_274 ();
 sg13g2_decap_8 FILLER_0_281 ();
 sg13g2_decap_8 FILLER_0_288 ();
 sg13g2_decap_8 FILLER_0_295 ();
 sg13g2_fill_2 FILLER_0_302 ();
 sg13g2_decap_8 FILLER_0_309 ();
 sg13g2_decap_8 FILLER_0_316 ();
 sg13g2_decap_8 FILLER_0_323 ();
 sg13g2_decap_8 FILLER_0_330 ();
 sg13g2_decap_8 FILLER_0_337 ();
 sg13g2_decap_4 FILLER_0_344 ();
 sg13g2_decap_4 FILLER_0_352 ();
 sg13g2_decap_8 FILLER_0_360 ();
 sg13g2_decap_8 FILLER_0_367 ();
 sg13g2_decap_8 FILLER_0_374 ();
 sg13g2_decap_8 FILLER_0_381 ();
 sg13g2_decap_8 FILLER_0_388 ();
 sg13g2_decap_8 FILLER_0_395 ();
 sg13g2_decap_8 FILLER_0_402 ();
 sg13g2_decap_8 FILLER_0_409 ();
 sg13g2_decap_8 FILLER_0_416 ();
 sg13g2_decap_8 FILLER_0_423 ();
 sg13g2_decap_8 FILLER_1_0 ();
 sg13g2_decap_8 FILLER_1_7 ();
 sg13g2_decap_8 FILLER_1_14 ();
 sg13g2_decap_8 FILLER_1_82 ();
 sg13g2_decap_8 FILLER_1_89 ();
 sg13g2_decap_4 FILLER_1_96 ();
 sg13g2_fill_2 FILLER_1_100 ();
 sg13g2_fill_1 FILLER_1_158 ();
 sg13g2_decap_8 FILLER_1_169 ();
 sg13g2_fill_2 FILLER_1_217 ();
 sg13g2_fill_1 FILLER_1_219 ();
 sg13g2_decap_4 FILLER_1_246 ();
 sg13g2_fill_2 FILLER_1_250 ();
 sg13g2_decap_4 FILLER_1_256 ();
 sg13g2_fill_1 FILLER_1_260 ();
 sg13g2_decap_4 FILLER_1_330 ();
 sg13g2_fill_2 FILLER_1_334 ();
 sg13g2_fill_1 FILLER_1_372 ();
 sg13g2_fill_1 FILLER_1_378 ();
 sg13g2_fill_1 FILLER_1_405 ();
 sg13g2_decap_8 FILLER_1_410 ();
 sg13g2_decap_8 FILLER_1_417 ();
 sg13g2_decap_4 FILLER_1_424 ();
 sg13g2_fill_2 FILLER_1_428 ();
 sg13g2_decap_8 FILLER_2_0 ();
 sg13g2_decap_8 FILLER_2_7 ();
 sg13g2_decap_8 FILLER_2_14 ();
 sg13g2_fill_2 FILLER_2_21 ();
 sg13g2_decap_8 FILLER_2_80 ();
 sg13g2_decap_8 FILLER_2_87 ();
 sg13g2_fill_1 FILLER_2_94 ();
 sg13g2_decap_8 FILLER_2_125 ();
 sg13g2_decap_4 FILLER_2_163 ();
 sg13g2_fill_2 FILLER_2_243 ();
 sg13g2_fill_2 FILLER_2_271 ();
 sg13g2_fill_1 FILLER_2_273 ();
 sg13g2_decap_4 FILLER_2_341 ();
 sg13g2_fill_2 FILLER_2_375 ();
 sg13g2_fill_1 FILLER_2_377 ();
 sg13g2_decap_8 FILLER_2_409 ();
 sg13g2_decap_8 FILLER_2_416 ();
 sg13g2_decap_8 FILLER_2_423 ();
 sg13g2_decap_8 FILLER_3_0 ();
 sg13g2_decap_8 FILLER_3_7 ();
 sg13g2_decap_8 FILLER_3_14 ();
 sg13g2_decap_8 FILLER_3_21 ();
 sg13g2_fill_2 FILLER_3_28 ();
 sg13g2_fill_1 FILLER_3_30 ();
 sg13g2_decap_8 FILLER_3_35 ();
 sg13g2_fill_2 FILLER_3_42 ();
 sg13g2_fill_2 FILLER_3_54 ();
 sg13g2_decap_4 FILLER_3_60 ();
 sg13g2_fill_2 FILLER_3_77 ();
 sg13g2_decap_8 FILLER_3_83 ();
 sg13g2_decap_4 FILLER_3_90 ();
 sg13g2_fill_2 FILLER_3_94 ();
 sg13g2_decap_8 FILLER_3_121 ();
 sg13g2_decap_4 FILLER_3_133 ();
 sg13g2_fill_2 FILLER_3_137 ();
 sg13g2_fill_1 FILLER_3_143 ();
 sg13g2_fill_2 FILLER_3_232 ();
 sg13g2_decap_8 FILLER_3_238 ();
 sg13g2_decap_8 FILLER_3_245 ();
 sg13g2_fill_2 FILLER_3_252 ();
 sg13g2_fill_1 FILLER_3_254 ();
 sg13g2_fill_2 FILLER_3_285 ();
 sg13g2_fill_1 FILLER_3_287 ();
 sg13g2_fill_2 FILLER_3_304 ();
 sg13g2_fill_1 FILLER_3_332 ();
 sg13g2_fill_1 FILLER_3_369 ();
 sg13g2_fill_1 FILLER_3_375 ();
 sg13g2_fill_1 FILLER_3_381 ();
 sg13g2_fill_2 FILLER_3_387 ();
 sg13g2_fill_2 FILLER_3_393 ();
 sg13g2_fill_1 FILLER_3_395 ();
 sg13g2_decap_8 FILLER_3_401 ();
 sg13g2_decap_8 FILLER_3_408 ();
 sg13g2_decap_8 FILLER_3_415 ();
 sg13g2_decap_8 FILLER_3_422 ();
 sg13g2_fill_1 FILLER_3_429 ();
 sg13g2_decap_8 FILLER_4_0 ();
 sg13g2_decap_8 FILLER_4_7 ();
 sg13g2_fill_2 FILLER_4_14 ();
 sg13g2_fill_2 FILLER_4_36 ();
 sg13g2_fill_1 FILLER_4_38 ();
 sg13g2_fill_2 FILLER_4_49 ();
 sg13g2_decap_8 FILLER_4_56 ();
 sg13g2_fill_2 FILLER_4_63 ();
 sg13g2_fill_2 FILLER_4_86 ();
 sg13g2_decap_8 FILLER_4_114 ();
 sg13g2_decap_8 FILLER_4_121 ();
 sg13g2_fill_2 FILLER_4_140 ();
 sg13g2_decap_4 FILLER_4_147 ();
 sg13g2_decap_8 FILLER_4_155 ();
 sg13g2_decap_8 FILLER_4_162 ();
 sg13g2_fill_1 FILLER_4_174 ();
 sg13g2_fill_2 FILLER_4_185 ();
 sg13g2_decap_8 FILLER_4_192 ();
 sg13g2_decap_8 FILLER_4_199 ();
 sg13g2_decap_4 FILLER_4_206 ();
 sg13g2_fill_1 FILLER_4_210 ();
 sg13g2_fill_1 FILLER_4_221 ();
 sg13g2_decap_8 FILLER_4_226 ();
 sg13g2_fill_2 FILLER_4_233 ();
 sg13g2_fill_1 FILLER_4_235 ();
 sg13g2_decap_4 FILLER_4_241 ();
 sg13g2_fill_1 FILLER_4_245 ();
 sg13g2_fill_2 FILLER_4_264 ();
 sg13g2_decap_4 FILLER_4_275 ();
 sg13g2_fill_2 FILLER_4_279 ();
 sg13g2_fill_2 FILLER_4_287 ();
 sg13g2_fill_1 FILLER_4_289 ();
 sg13g2_decap_4 FILLER_4_324 ();
 sg13g2_fill_1 FILLER_4_328 ();
 sg13g2_fill_2 FILLER_4_334 ();
 sg13g2_decap_4 FILLER_4_341 ();
 sg13g2_fill_1 FILLER_4_345 ();
 sg13g2_decap_4 FILLER_4_356 ();
 sg13g2_fill_2 FILLER_4_360 ();
 sg13g2_decap_8 FILLER_4_371 ();
 sg13g2_decap_8 FILLER_4_391 ();
 sg13g2_decap_8 FILLER_4_398 ();
 sg13g2_decap_8 FILLER_4_405 ();
 sg13g2_decap_8 FILLER_4_412 ();
 sg13g2_decap_8 FILLER_4_419 ();
 sg13g2_decap_4 FILLER_4_426 ();
 sg13g2_decap_8 FILLER_5_0 ();
 sg13g2_decap_8 FILLER_5_7 ();
 sg13g2_decap_8 FILLER_5_14 ();
 sg13g2_decap_8 FILLER_5_21 ();
 sg13g2_decap_4 FILLER_5_28 ();
 sg13g2_fill_2 FILLER_5_32 ();
 sg13g2_fill_1 FILLER_5_58 ();
 sg13g2_fill_2 FILLER_5_63 ();
 sg13g2_fill_1 FILLER_5_78 ();
 sg13g2_fill_2 FILLER_5_84 ();
 sg13g2_fill_1 FILLER_5_90 ();
 sg13g2_fill_2 FILLER_5_95 ();
 sg13g2_fill_1 FILLER_5_117 ();
 sg13g2_fill_1 FILLER_5_122 ();
 sg13g2_fill_2 FILLER_5_127 ();
 sg13g2_fill_2 FILLER_5_139 ();
 sg13g2_fill_1 FILLER_5_141 ();
 sg13g2_decap_4 FILLER_5_150 ();
 sg13g2_fill_1 FILLER_5_154 ();
 sg13g2_fill_2 FILLER_5_169 ();
 sg13g2_fill_1 FILLER_5_171 ();
 sg13g2_fill_2 FILLER_5_177 ();
 sg13g2_decap_8 FILLER_5_184 ();
 sg13g2_decap_8 FILLER_5_191 ();
 sg13g2_fill_1 FILLER_5_198 ();
 sg13g2_fill_1 FILLER_5_214 ();
 sg13g2_fill_1 FILLER_5_241 ();
 sg13g2_fill_1 FILLER_5_268 ();
 sg13g2_fill_2 FILLER_5_273 ();
 sg13g2_fill_2 FILLER_5_279 ();
 sg13g2_fill_1 FILLER_5_281 ();
 sg13g2_fill_2 FILLER_5_287 ();
 sg13g2_fill_1 FILLER_5_289 ();
 sg13g2_decap_4 FILLER_5_298 ();
 sg13g2_fill_2 FILLER_5_314 ();
 sg13g2_fill_1 FILLER_5_316 ();
 sg13g2_decap_8 FILLER_5_320 ();
 sg13g2_decap_8 FILLER_5_327 ();
 sg13g2_fill_2 FILLER_5_334 ();
 sg13g2_fill_1 FILLER_5_336 ();
 sg13g2_decap_4 FILLER_5_341 ();
 sg13g2_fill_1 FILLER_5_345 ();
 sg13g2_decap_8 FILLER_5_356 ();
 sg13g2_fill_1 FILLER_5_366 ();
 sg13g2_decap_8 FILLER_5_402 ();
 sg13g2_decap_8 FILLER_5_409 ();
 sg13g2_decap_8 FILLER_5_416 ();
 sg13g2_decap_8 FILLER_5_423 ();
 sg13g2_decap_8 FILLER_6_0 ();
 sg13g2_decap_4 FILLER_6_7 ();
 sg13g2_decap_4 FILLER_6_47 ();
 sg13g2_fill_2 FILLER_6_83 ();
 sg13g2_decap_4 FILLER_6_137 ();
 sg13g2_fill_2 FILLER_6_202 ();
 sg13g2_fill_1 FILLER_6_204 ();
 sg13g2_fill_1 FILLER_6_209 ();
 sg13g2_fill_2 FILLER_6_236 ();
 sg13g2_fill_1 FILLER_6_238 ();
 sg13g2_fill_1 FILLER_6_243 ();
 sg13g2_fill_2 FILLER_6_254 ();
 sg13g2_fill_2 FILLER_6_260 ();
 sg13g2_fill_2 FILLER_6_285 ();
 sg13g2_decap_8 FILLER_6_312 ();
 sg13g2_decap_4 FILLER_6_326 ();
 sg13g2_fill_2 FILLER_6_330 ();
 sg13g2_fill_1 FILLER_6_362 ();
 sg13g2_fill_1 FILLER_6_366 ();
 sg13g2_fill_1 FILLER_6_393 ();
 sg13g2_decap_8 FILLER_6_420 ();
 sg13g2_fill_2 FILLER_6_427 ();
 sg13g2_fill_1 FILLER_6_429 ();
 sg13g2_decap_4 FILLER_7_0 ();
 sg13g2_fill_2 FILLER_7_4 ();
 sg13g2_fill_1 FILLER_7_67 ();
 sg13g2_decap_8 FILLER_7_78 ();
 sg13g2_decap_4 FILLER_7_85 ();
 sg13g2_fill_1 FILLER_7_89 ();
 sg13g2_decap_4 FILLER_7_94 ();
 sg13g2_fill_2 FILLER_7_98 ();
 sg13g2_fill_1 FILLER_7_109 ();
 sg13g2_fill_1 FILLER_7_115 ();
 sg13g2_fill_1 FILLER_7_141 ();
 sg13g2_decap_4 FILLER_7_152 ();
 sg13g2_fill_1 FILLER_7_156 ();
 sg13g2_decap_4 FILLER_7_186 ();
 sg13g2_fill_2 FILLER_7_190 ();
 sg13g2_fill_1 FILLER_7_201 ();
 sg13g2_fill_1 FILLER_7_210 ();
 sg13g2_fill_1 FILLER_7_216 ();
 sg13g2_fill_1 FILLER_7_220 ();
 sg13g2_decap_4 FILLER_7_225 ();
 sg13g2_fill_1 FILLER_7_235 ();
 sg13g2_fill_2 FILLER_7_266 ();
 sg13g2_fill_1 FILLER_7_325 ();
 sg13g2_fill_1 FILLER_7_330 ();
 sg13g2_fill_1 FILLER_7_336 ();
 sg13g2_fill_1 FILLER_7_342 ();
 sg13g2_decap_4 FILLER_7_350 ();
 sg13g2_fill_2 FILLER_7_383 ();
 sg13g2_fill_1 FILLER_7_385 ();
 sg13g2_decap_8 FILLER_7_421 ();
 sg13g2_fill_2 FILLER_7_428 ();
 sg13g2_decap_4 FILLER_8_0 ();
 sg13g2_fill_1 FILLER_8_4 ();
 sg13g2_fill_1 FILLER_8_15 ();
 sg13g2_fill_2 FILLER_8_24 ();
 sg13g2_fill_1 FILLER_8_30 ();
 sg13g2_decap_4 FILLER_8_35 ();
 sg13g2_decap_4 FILLER_8_46 ();
 sg13g2_fill_2 FILLER_8_50 ();
 sg13g2_decap_8 FILLER_8_56 ();
 sg13g2_decap_8 FILLER_8_63 ();
 sg13g2_fill_2 FILLER_8_91 ();
 sg13g2_fill_1 FILLER_8_98 ();
 sg13g2_decap_8 FILLER_8_110 ();
 sg13g2_decap_4 FILLER_8_117 ();
 sg13g2_fill_2 FILLER_8_121 ();
 sg13g2_decap_4 FILLER_8_131 ();
 sg13g2_fill_1 FILLER_8_135 ();
 sg13g2_fill_2 FILLER_8_154 ();
 sg13g2_fill_1 FILLER_8_177 ();
 sg13g2_fill_1 FILLER_8_182 ();
 sg13g2_decap_8 FILLER_8_236 ();
 sg13g2_fill_2 FILLER_8_243 ();
 sg13g2_fill_1 FILLER_8_245 ();
 sg13g2_decap_4 FILLER_8_260 ();
 sg13g2_decap_4 FILLER_8_292 ();
 sg13g2_fill_2 FILLER_8_296 ();
 sg13g2_decap_8 FILLER_8_335 ();
 sg13g2_decap_8 FILLER_8_342 ();
 sg13g2_decap_8 FILLER_8_349 ();
 sg13g2_decap_4 FILLER_8_369 ();
 sg13g2_fill_2 FILLER_8_373 ();
 sg13g2_fill_1 FILLER_8_379 ();
 sg13g2_fill_1 FILLER_8_384 ();
 sg13g2_fill_2 FILLER_8_400 ();
 sg13g2_fill_1 FILLER_8_407 ();
 sg13g2_fill_1 FILLER_8_417 ();
 sg13g2_fill_1 FILLER_8_422 ();
 sg13g2_fill_2 FILLER_8_427 ();
 sg13g2_fill_1 FILLER_8_429 ();
 sg13g2_decap_8 FILLER_9_0 ();
 sg13g2_fill_2 FILLER_9_7 ();
 sg13g2_decap_4 FILLER_9_35 ();
 sg13g2_fill_1 FILLER_9_39 ();
 sg13g2_decap_8 FILLER_9_58 ();
 sg13g2_decap_8 FILLER_9_65 ();
 sg13g2_fill_1 FILLER_9_72 ();
 sg13g2_fill_2 FILLER_9_89 ();
 sg13g2_decap_4 FILLER_9_101 ();
 sg13g2_decap_8 FILLER_9_114 ();
 sg13g2_fill_2 FILLER_9_121 ();
 sg13g2_fill_1 FILLER_9_127 ();
 sg13g2_decap_4 FILLER_9_134 ();
 sg13g2_fill_1 FILLER_9_138 ();
 sg13g2_fill_2 FILLER_9_171 ();
 sg13g2_decap_4 FILLER_9_181 ();
 sg13g2_fill_2 FILLER_9_185 ();
 sg13g2_fill_2 FILLER_9_192 ();
 sg13g2_fill_1 FILLER_9_194 ();
 sg13g2_fill_1 FILLER_9_208 ();
 sg13g2_fill_1 FILLER_9_218 ();
 sg13g2_decap_4 FILLER_9_240 ();
 sg13g2_fill_2 FILLER_9_244 ();
 sg13g2_fill_1 FILLER_9_290 ();
 sg13g2_fill_2 FILLER_9_304 ();
 sg13g2_fill_1 FILLER_9_306 ();
 sg13g2_fill_1 FILLER_9_312 ();
 sg13g2_fill_1 FILLER_9_318 ();
 sg13g2_fill_2 FILLER_9_329 ();
 sg13g2_fill_1 FILLER_9_331 ();
 sg13g2_fill_2 FILLER_9_336 ();
 sg13g2_fill_1 FILLER_9_342 ();
 sg13g2_decap_4 FILLER_9_375 ();
 sg13g2_fill_2 FILLER_9_379 ();
 sg13g2_fill_1 FILLER_9_385 ();
 sg13g2_fill_1 FILLER_9_391 ();
 sg13g2_fill_1 FILLER_9_402 ();
 sg13g2_fill_1 FILLER_9_429 ();
 sg13g2_decap_4 FILLER_10_0 ();
 sg13g2_fill_1 FILLER_10_4 ();
 sg13g2_decap_8 FILLER_10_15 ();
 sg13g2_decap_8 FILLER_10_22 ();
 sg13g2_fill_2 FILLER_10_29 ();
 sg13g2_fill_1 FILLER_10_31 ();
 sg13g2_fill_1 FILLER_10_35 ();
 sg13g2_decap_4 FILLER_10_40 ();
 sg13g2_fill_2 FILLER_10_57 ();
 sg13g2_fill_2 FILLER_10_64 ();
 sg13g2_fill_1 FILLER_10_66 ();
 sg13g2_decap_4 FILLER_10_72 ();
 sg13g2_fill_1 FILLER_10_85 ();
 sg13g2_fill_1 FILLER_10_92 ();
 sg13g2_fill_2 FILLER_10_106 ();
 sg13g2_fill_1 FILLER_10_108 ();
 sg13g2_fill_2 FILLER_10_113 ();
 sg13g2_fill_2 FILLER_10_141 ();
 sg13g2_fill_1 FILLER_10_143 ();
 sg13g2_fill_2 FILLER_10_172 ();
 sg13g2_fill_1 FILLER_10_182 ();
 sg13g2_decap_8 FILLER_10_189 ();
 sg13g2_decap_8 FILLER_10_196 ();
 sg13g2_fill_1 FILLER_10_203 ();
 sg13g2_decap_4 FILLER_10_208 ();
 sg13g2_fill_1 FILLER_10_212 ();
 sg13g2_decap_8 FILLER_10_240 ();
 sg13g2_decap_4 FILLER_10_247 ();
 sg13g2_fill_1 FILLER_10_251 ();
 sg13g2_decap_4 FILLER_10_257 ();
 sg13g2_decap_4 FILLER_10_324 ();
 sg13g2_fill_1 FILLER_10_336 ();
 sg13g2_fill_2 FILLER_10_341 ();
 sg13g2_decap_4 FILLER_10_348 ();
 sg13g2_decap_4 FILLER_10_367 ();
 sg13g2_decap_4 FILLER_10_384 ();
 sg13g2_fill_1 FILLER_10_388 ();
 sg13g2_decap_8 FILLER_10_394 ();
 sg13g2_fill_1 FILLER_10_401 ();
 sg13g2_fill_2 FILLER_10_428 ();
 sg13g2_decap_8 FILLER_11_26 ();
 sg13g2_fill_2 FILLER_11_45 ();
 sg13g2_fill_1 FILLER_11_84 ();
 sg13g2_fill_1 FILLER_11_97 ();
 sg13g2_fill_2 FILLER_11_102 ();
 sg13g2_decap_8 FILLER_11_114 ();
 sg13g2_fill_1 FILLER_11_121 ();
 sg13g2_decap_8 FILLER_11_143 ();
 sg13g2_decap_8 FILLER_11_150 ();
 sg13g2_decap_8 FILLER_11_157 ();
 sg13g2_fill_2 FILLER_11_164 ();
 sg13g2_fill_1 FILLER_11_166 ();
 sg13g2_fill_1 FILLER_11_178 ();
 sg13g2_fill_1 FILLER_11_196 ();
 sg13g2_fill_1 FILLER_11_202 ();
 sg13g2_decap_4 FILLER_11_208 ();
 sg13g2_fill_1 FILLER_11_212 ();
 sg13g2_decap_8 FILLER_11_222 ();
 sg13g2_decap_8 FILLER_11_229 ();
 sg13g2_decap_8 FILLER_11_236 ();
 sg13g2_decap_4 FILLER_11_243 ();
 sg13g2_fill_1 FILLER_11_247 ();
 sg13g2_fill_2 FILLER_11_252 ();
 sg13g2_decap_4 FILLER_11_259 ();
 sg13g2_fill_2 FILLER_11_263 ();
 sg13g2_decap_4 FILLER_11_269 ();
 sg13g2_fill_2 FILLER_11_273 ();
 sg13g2_decap_8 FILLER_11_305 ();
 sg13g2_fill_1 FILLER_11_312 ();
 sg13g2_fill_2 FILLER_11_320 ();
 sg13g2_fill_2 FILLER_11_326 ();
 sg13g2_fill_2 FILLER_11_340 ();
 sg13g2_decap_4 FILLER_11_359 ();
 sg13g2_decap_8 FILLER_11_370 ();
 sg13g2_fill_2 FILLER_11_377 ();
 sg13g2_decap_4 FILLER_11_386 ();
 sg13g2_decap_8 FILLER_11_399 ();
 sg13g2_fill_2 FILLER_11_427 ();
 sg13g2_fill_1 FILLER_11_429 ();
 sg13g2_decap_8 FILLER_12_0 ();
 sg13g2_decap_8 FILLER_12_11 ();
 sg13g2_fill_2 FILLER_12_18 ();
 sg13g2_fill_1 FILLER_12_20 ();
 sg13g2_fill_1 FILLER_12_31 ();
 sg13g2_decap_8 FILLER_12_63 ();
 sg13g2_decap_8 FILLER_12_93 ();
 sg13g2_decap_8 FILLER_12_100 ();
 sg13g2_decap_8 FILLER_12_120 ();
 sg13g2_fill_2 FILLER_12_127 ();
 sg13g2_decap_4 FILLER_12_134 ();
 sg13g2_fill_1 FILLER_12_138 ();
 sg13g2_decap_4 FILLER_12_151 ();
 sg13g2_fill_2 FILLER_12_155 ();
 sg13g2_fill_1 FILLER_12_169 ();
 sg13g2_fill_2 FILLER_12_174 ();
 sg13g2_fill_2 FILLER_12_186 ();
 sg13g2_fill_1 FILLER_12_188 ();
 sg13g2_fill_1 FILLER_12_200 ();
 sg13g2_fill_2 FILLER_12_205 ();
 sg13g2_decap_4 FILLER_12_233 ();
 sg13g2_fill_1 FILLER_12_237 ();
 sg13g2_decap_8 FILLER_12_273 ();
 sg13g2_decap_8 FILLER_12_280 ();
 sg13g2_fill_2 FILLER_12_287 ();
 sg13g2_fill_1 FILLER_12_289 ();
 sg13g2_fill_2 FILLER_12_306 ();
 sg13g2_fill_2 FILLER_12_339 ();
 sg13g2_fill_2 FILLER_12_362 ();
 sg13g2_fill_1 FILLER_12_364 ();
 sg13g2_decap_8 FILLER_12_390 ();
 sg13g2_fill_2 FILLER_12_397 ();
 sg13g2_decap_8 FILLER_13_0 ();
 sg13g2_decap_8 FILLER_13_7 ();
 sg13g2_decap_4 FILLER_13_14 ();
 sg13g2_fill_1 FILLER_13_18 ();
 sg13g2_decap_8 FILLER_13_29 ();
 sg13g2_fill_2 FILLER_13_79 ();
 sg13g2_decap_8 FILLER_13_88 ();
 sg13g2_decap_8 FILLER_13_95 ();
 sg13g2_fill_2 FILLER_13_102 ();
 sg13g2_fill_1 FILLER_13_104 ();
 sg13g2_fill_2 FILLER_13_140 ();
 sg13g2_fill_1 FILLER_13_142 ();
 sg13g2_decap_8 FILLER_13_175 ();
 sg13g2_fill_1 FILLER_13_182 ();
 sg13g2_fill_2 FILLER_13_201 ();
 sg13g2_fill_2 FILLER_13_226 ();
 sg13g2_fill_2 FILLER_13_245 ();
 sg13g2_fill_1 FILLER_13_247 ();
 sg13g2_fill_1 FILLER_13_258 ();
 sg13g2_decap_8 FILLER_13_265 ();
 sg13g2_fill_1 FILLER_13_272 ();
 sg13g2_decap_8 FILLER_13_277 ();
 sg13g2_decap_4 FILLER_13_284 ();
 sg13g2_decap_8 FILLER_13_313 ();
 sg13g2_decap_8 FILLER_13_320 ();
 sg13g2_fill_2 FILLER_13_327 ();
 sg13g2_fill_1 FILLER_13_329 ();
 sg13g2_decap_4 FILLER_13_339 ();
 sg13g2_fill_2 FILLER_13_343 ();
 sg13g2_decap_4 FILLER_13_350 ();
 sg13g2_fill_2 FILLER_13_354 ();
 sg13g2_fill_1 FILLER_13_361 ();
 sg13g2_fill_1 FILLER_13_366 ();
 sg13g2_fill_2 FILLER_13_372 ();
 sg13g2_fill_2 FILLER_13_395 ();
 sg13g2_fill_2 FILLER_13_401 ();
 sg13g2_fill_1 FILLER_13_403 ();
 sg13g2_decap_4 FILLER_14_0 ();
 sg13g2_fill_1 FILLER_14_4 ();
 sg13g2_fill_1 FILLER_14_15 ();
 sg13g2_fill_2 FILLER_14_42 ();
 sg13g2_fill_1 FILLER_14_44 ();
 sg13g2_fill_2 FILLER_14_76 ();
 sg13g2_decap_8 FILLER_14_86 ();
 sg13g2_decap_8 FILLER_14_93 ();
 sg13g2_decap_8 FILLER_14_100 ();
 sg13g2_fill_2 FILLER_14_107 ();
 sg13g2_fill_1 FILLER_14_139 ();
 sg13g2_fill_1 FILLER_14_174 ();
 sg13g2_fill_1 FILLER_14_194 ();
 sg13g2_fill_1 FILLER_14_200 ();
 sg13g2_fill_1 FILLER_14_208 ();
 sg13g2_fill_1 FILLER_14_214 ();
 sg13g2_fill_1 FILLER_14_241 ();
 sg13g2_fill_1 FILLER_14_250 ();
 sg13g2_fill_1 FILLER_14_257 ();
 sg13g2_fill_2 FILLER_14_279 ();
 sg13g2_fill_1 FILLER_14_281 ();
 sg13g2_decap_8 FILLER_14_285 ();
 sg13g2_decap_8 FILLER_14_316 ();
 sg13g2_decap_4 FILLER_14_323 ();
 sg13g2_fill_1 FILLER_14_340 ();
 sg13g2_decap_8 FILLER_14_346 ();
 sg13g2_fill_2 FILLER_14_353 ();
 sg13g2_fill_2 FILLER_14_403 ();
 sg13g2_fill_2 FILLER_14_409 ();
 sg13g2_fill_1 FILLER_14_419 ();
 sg13g2_decap_4 FILLER_14_425 ();
 sg13g2_fill_1 FILLER_14_429 ();
 sg13g2_fill_2 FILLER_15_4 ();
 sg13g2_fill_1 FILLER_15_6 ();
 sg13g2_fill_2 FILLER_15_43 ();
 sg13g2_fill_2 FILLER_15_50 ();
 sg13g2_fill_1 FILLER_15_52 ();
 sg13g2_fill_2 FILLER_15_57 ();
 sg13g2_fill_1 FILLER_15_59 ();
 sg13g2_fill_1 FILLER_15_85 ();
 sg13g2_decap_8 FILLER_15_94 ();
 sg13g2_decap_8 FILLER_15_101 ();
 sg13g2_fill_2 FILLER_15_108 ();
 sg13g2_fill_1 FILLER_15_110 ();
 sg13g2_fill_2 FILLER_15_121 ();
 sg13g2_fill_2 FILLER_15_136 ();
 sg13g2_fill_1 FILLER_15_142 ();
 sg13g2_fill_2 FILLER_15_147 ();
 sg13g2_fill_1 FILLER_15_157 ();
 sg13g2_fill_1 FILLER_15_163 ();
 sg13g2_fill_1 FILLER_15_199 ();
 sg13g2_fill_1 FILLER_15_205 ();
 sg13g2_fill_1 FILLER_15_210 ();
 sg13g2_fill_2 FILLER_15_237 ();
 sg13g2_fill_2 FILLER_15_247 ();
 sg13g2_fill_1 FILLER_15_258 ();
 sg13g2_fill_1 FILLER_15_280 ();
 sg13g2_fill_1 FILLER_15_289 ();
 sg13g2_fill_1 FILLER_15_294 ();
 sg13g2_fill_1 FILLER_15_300 ();
 sg13g2_fill_1 FILLER_15_315 ();
 sg13g2_fill_2 FILLER_15_332 ();
 sg13g2_fill_1 FILLER_15_340 ();
 sg13g2_fill_2 FILLER_15_349 ();
 sg13g2_decap_8 FILLER_15_382 ();
 sg13g2_decap_8 FILLER_15_407 ();
 sg13g2_decap_8 FILLER_15_414 ();
 sg13g2_decap_8 FILLER_15_421 ();
 sg13g2_fill_2 FILLER_15_428 ();
 sg13g2_fill_2 FILLER_16_0 ();
 sg13g2_fill_2 FILLER_16_30 ();
 sg13g2_fill_1 FILLER_16_32 ();
 sg13g2_decap_8 FILLER_16_36 ();
 sg13g2_fill_1 FILLER_16_43 ();
 sg13g2_decap_8 FILLER_16_54 ();
 sg13g2_fill_2 FILLER_16_84 ();
 sg13g2_fill_1 FILLER_16_86 ();
 sg13g2_decap_4 FILLER_16_97 ();
 sg13g2_fill_2 FILLER_16_105 ();
 sg13g2_decap_8 FILLER_16_111 ();
 sg13g2_decap_4 FILLER_16_118 ();
 sg13g2_decap_4 FILLER_16_126 ();
 sg13g2_fill_1 FILLER_16_130 ();
 sg13g2_fill_2 FILLER_16_165 ();
 sg13g2_decap_8 FILLER_16_171 ();
 sg13g2_fill_2 FILLER_16_221 ();
 sg13g2_fill_1 FILLER_16_223 ();
 sg13g2_fill_1 FILLER_16_245 ();
 sg13g2_fill_2 FILLER_16_259 ();
 sg13g2_fill_1 FILLER_16_261 ();
 sg13g2_fill_2 FILLER_16_266 ();
 sg13g2_fill_1 FILLER_16_268 ();
 sg13g2_decap_4 FILLER_16_276 ();
 sg13g2_fill_1 FILLER_16_315 ();
 sg13g2_fill_2 FILLER_16_324 ();
 sg13g2_decap_8 FILLER_16_334 ();
 sg13g2_fill_2 FILLER_16_341 ();
 sg13g2_fill_2 FILLER_16_356 ();
 sg13g2_fill_2 FILLER_16_363 ();
 sg13g2_fill_1 FILLER_16_368 ();
 sg13g2_fill_1 FILLER_16_390 ();
 sg13g2_fill_1 FILLER_16_395 ();
 sg13g2_fill_1 FILLER_16_401 ();
 sg13g2_fill_2 FILLER_16_407 ();
 sg13g2_decap_4 FILLER_16_413 ();
 sg13g2_fill_1 FILLER_16_417 ();
 sg13g2_decap_8 FILLER_16_422 ();
 sg13g2_fill_1 FILLER_16_429 ();
 sg13g2_fill_1 FILLER_17_0 ();
 sg13g2_decap_4 FILLER_17_12 ();
 sg13g2_decap_8 FILLER_17_35 ();
 sg13g2_fill_2 FILLER_17_42 ();
 sg13g2_fill_1 FILLER_17_44 ();
 sg13g2_fill_1 FILLER_17_51 ();
 sg13g2_decap_4 FILLER_17_61 ();
 sg13g2_fill_1 FILLER_17_88 ();
 sg13g2_fill_1 FILLER_17_92 ();
 sg13g2_fill_2 FILLER_17_119 ();
 sg13g2_fill_1 FILLER_17_121 ();
 sg13g2_fill_1 FILLER_17_132 ();
 sg13g2_fill_2 FILLER_17_151 ();
 sg13g2_fill_2 FILLER_17_163 ();
 sg13g2_fill_1 FILLER_17_165 ();
 sg13g2_decap_8 FILLER_17_171 ();
 sg13g2_fill_1 FILLER_17_178 ();
 sg13g2_fill_2 FILLER_17_187 ();
 sg13g2_fill_1 FILLER_17_189 ();
 sg13g2_decap_8 FILLER_17_198 ();
 sg13g2_decap_8 FILLER_17_209 ();
 sg13g2_decap_8 FILLER_17_216 ();
 sg13g2_decap_4 FILLER_17_223 ();
 sg13g2_decap_8 FILLER_17_253 ();
 sg13g2_decap_8 FILLER_17_260 ();
 sg13g2_fill_2 FILLER_17_267 ();
 sg13g2_fill_2 FILLER_17_273 ();
 sg13g2_fill_2 FILLER_17_279 ();
 sg13g2_fill_2 FILLER_17_296 ();
 sg13g2_decap_8 FILLER_17_311 ();
 sg13g2_decap_4 FILLER_17_318 ();
 sg13g2_fill_2 FILLER_17_322 ();
 sg13g2_decap_4 FILLER_17_329 ();
 sg13g2_fill_1 FILLER_17_333 ();
 sg13g2_fill_2 FILLER_17_346 ();
 sg13g2_decap_4 FILLER_17_390 ();
 sg13g2_decap_4 FILLER_18_0 ();
 sg13g2_decap_8 FILLER_18_8 ();
 sg13g2_fill_2 FILLER_18_15 ();
 sg13g2_fill_1 FILLER_18_17 ();
 sg13g2_decap_8 FILLER_18_22 ();
 sg13g2_decap_4 FILLER_18_29 ();
 sg13g2_fill_1 FILLER_18_33 ();
 sg13g2_decap_4 FILLER_18_38 ();
 sg13g2_fill_1 FILLER_18_42 ();
 sg13g2_fill_1 FILLER_18_103 ();
 sg13g2_fill_1 FILLER_18_112 ();
 sg13g2_decap_4 FILLER_18_117 ();
 sg13g2_decap_8 FILLER_18_125 ();
 sg13g2_fill_1 FILLER_18_136 ();
 sg13g2_decap_4 FILLER_18_145 ();
 sg13g2_fill_1 FILLER_18_149 ();
 sg13g2_fill_2 FILLER_18_160 ();
 sg13g2_decap_4 FILLER_18_174 ();
 sg13g2_fill_2 FILLER_18_217 ();
 sg13g2_fill_1 FILLER_18_219 ();
 sg13g2_decap_8 FILLER_18_224 ();
 sg13g2_decap_8 FILLER_18_231 ();
 sg13g2_fill_2 FILLER_18_247 ();
 sg13g2_fill_1 FILLER_18_267 ();
 sg13g2_decap_8 FILLER_18_273 ();
 sg13g2_decap_8 FILLER_18_280 ();
 sg13g2_fill_1 FILLER_18_287 ();
 sg13g2_fill_2 FILLER_18_301 ();
 sg13g2_decap_8 FILLER_18_308 ();
 sg13g2_decap_8 FILLER_18_315 ();
 sg13g2_decap_4 FILLER_18_322 ();
 sg13g2_fill_1 FILLER_18_326 ();
 sg13g2_fill_1 FILLER_18_335 ();
 sg13g2_fill_1 FILLER_18_342 ();
 sg13g2_decap_4 FILLER_18_353 ();
 sg13g2_fill_2 FILLER_18_357 ();
 sg13g2_fill_2 FILLER_18_364 ();
 sg13g2_fill_2 FILLER_18_391 ();
 sg13g2_fill_1 FILLER_18_393 ();
 sg13g2_fill_2 FILLER_18_397 ();
 sg13g2_fill_1 FILLER_18_399 ();
 sg13g2_fill_1 FILLER_19_0 ();
 sg13g2_fill_2 FILLER_19_24 ();
 sg13g2_fill_1 FILLER_19_26 ();
 sg13g2_decap_8 FILLER_19_57 ();
 sg13g2_fill_2 FILLER_19_64 ();
 sg13g2_fill_1 FILLER_19_66 ();
 sg13g2_fill_2 FILLER_19_76 ();
 sg13g2_fill_1 FILLER_19_78 ();
 sg13g2_fill_2 FILLER_19_85 ();
 sg13g2_fill_1 FILLER_19_87 ();
 sg13g2_decap_4 FILLER_19_114 ();
 sg13g2_decap_8 FILLER_19_122 ();
 sg13g2_decap_8 FILLER_19_129 ();
 sg13g2_decap_8 FILLER_19_136 ();
 sg13g2_fill_2 FILLER_19_143 ();
 sg13g2_fill_1 FILLER_19_145 ();
 sg13g2_decap_4 FILLER_19_163 ();
 sg13g2_fill_2 FILLER_19_167 ();
 sg13g2_fill_1 FILLER_19_192 ();
 sg13g2_fill_2 FILLER_19_205 ();
 sg13g2_fill_2 FILLER_19_233 ();
 sg13g2_fill_1 FILLER_19_235 ();
 sg13g2_fill_1 FILLER_19_242 ();
 sg13g2_fill_2 FILLER_19_247 ();
 sg13g2_fill_1 FILLER_19_280 ();
 sg13g2_fill_1 FILLER_19_299 ();
 sg13g2_decap_8 FILLER_19_309 ();
 sg13g2_decap_4 FILLER_19_316 ();
 sg13g2_fill_1 FILLER_19_320 ();
 sg13g2_decap_8 FILLER_19_344 ();
 sg13g2_decap_8 FILLER_19_351 ();
 sg13g2_fill_2 FILLER_19_358 ();
 sg13g2_fill_1 FILLER_19_363 ();
 sg13g2_decap_8 FILLER_19_381 ();
 sg13g2_fill_2 FILLER_19_388 ();
 sg13g2_fill_2 FILLER_19_394 ();
 sg13g2_fill_1 FILLER_19_396 ();
 sg13g2_decap_8 FILLER_19_402 ();
 sg13g2_fill_2 FILLER_19_409 ();
 sg13g2_decap_8 FILLER_19_415 ();
 sg13g2_decap_4 FILLER_19_426 ();
 sg13g2_fill_2 FILLER_20_0 ();
 sg13g2_fill_2 FILLER_20_13 ();
 sg13g2_decap_8 FILLER_20_51 ();
 sg13g2_decap_8 FILLER_20_58 ();
 sg13g2_decap_8 FILLER_20_65 ();
 sg13g2_fill_2 FILLER_20_72 ();
 sg13g2_fill_1 FILLER_20_74 ();
 sg13g2_fill_1 FILLER_20_79 ();
 sg13g2_fill_2 FILLER_20_91 ();
 sg13g2_decap_8 FILLER_20_112 ();
 sg13g2_fill_2 FILLER_20_119 ();
 sg13g2_decap_8 FILLER_20_131 ();
 sg13g2_decap_8 FILLER_20_143 ();
 sg13g2_fill_2 FILLER_20_155 ();
 sg13g2_decap_4 FILLER_20_162 ();
 sg13g2_decap_8 FILLER_20_172 ();
 sg13g2_fill_2 FILLER_20_183 ();
 sg13g2_decap_8 FILLER_20_190 ();
 sg13g2_fill_2 FILLER_20_197 ();
 sg13g2_fill_1 FILLER_20_199 ();
 sg13g2_decap_8 FILLER_20_244 ();
 sg13g2_fill_1 FILLER_20_264 ();
 sg13g2_decap_4 FILLER_20_270 ();
 sg13g2_decap_8 FILLER_20_278 ();
 sg13g2_decap_4 FILLER_20_303 ();
 sg13g2_fill_2 FILLER_20_307 ();
 sg13g2_decap_4 FILLER_20_344 ();
 sg13g2_fill_1 FILLER_20_348 ();
 sg13g2_fill_1 FILLER_20_359 ();
 sg13g2_fill_1 FILLER_20_391 ();
 sg13g2_decap_8 FILLER_20_400 ();
 sg13g2_fill_2 FILLER_20_407 ();
 sg13g2_decap_8 FILLER_20_414 ();
 sg13g2_decap_8 FILLER_20_421 ();
 sg13g2_fill_2 FILLER_20_428 ();
 sg13g2_fill_2 FILLER_21_0 ();
 sg13g2_decap_4 FILLER_21_14 ();
 sg13g2_fill_2 FILLER_21_41 ();
 sg13g2_fill_1 FILLER_21_53 ();
 sg13g2_decap_4 FILLER_21_58 ();
 sg13g2_fill_1 FILLER_21_96 ();
 sg13g2_decap_8 FILLER_21_102 ();
 sg13g2_fill_1 FILLER_21_109 ();
 sg13g2_fill_2 FILLER_21_159 ();
 sg13g2_fill_1 FILLER_21_161 ();
 sg13g2_fill_1 FILLER_21_168 ();
 sg13g2_decap_8 FILLER_21_175 ();
 sg13g2_decap_4 FILLER_21_197 ();
 sg13g2_fill_1 FILLER_21_201 ();
 sg13g2_fill_1 FILLER_21_206 ();
 sg13g2_fill_1 FILLER_21_212 ();
 sg13g2_fill_2 FILLER_21_217 ();
 sg13g2_fill_2 FILLER_21_223 ();
 sg13g2_fill_1 FILLER_21_225 ();
 sg13g2_decap_8 FILLER_21_230 ();
 sg13g2_decap_8 FILLER_21_246 ();
 sg13g2_fill_2 FILLER_21_253 ();
 sg13g2_fill_2 FILLER_21_259 ();
 sg13g2_fill_1 FILLER_21_261 ();
 sg13g2_fill_2 FILLER_21_316 ();
 sg13g2_decap_8 FILLER_21_322 ();
 sg13g2_fill_2 FILLER_21_329 ();
 sg13g2_decap_8 FILLER_22_0 ();
 sg13g2_decap_4 FILLER_22_17 ();
 sg13g2_fill_1 FILLER_22_21 ();
 sg13g2_fill_2 FILLER_22_75 ();
 sg13g2_decap_8 FILLER_22_95 ();
 sg13g2_decap_4 FILLER_22_102 ();
 sg13g2_fill_2 FILLER_22_106 ();
 sg13g2_fill_1 FILLER_22_130 ();
 sg13g2_fill_2 FILLER_22_148 ();
 sg13g2_fill_1 FILLER_22_172 ();
 sg13g2_fill_1 FILLER_22_178 ();
 sg13g2_fill_2 FILLER_22_184 ();
 sg13g2_fill_1 FILLER_22_186 ();
 sg13g2_fill_1 FILLER_22_210 ();
 sg13g2_decap_4 FILLER_22_237 ();
 sg13g2_fill_2 FILLER_22_241 ();
 sg13g2_fill_2 FILLER_22_247 ();
 sg13g2_decap_8 FILLER_22_254 ();
 sg13g2_decap_8 FILLER_22_261 ();
 sg13g2_decap_8 FILLER_22_272 ();
 sg13g2_decap_4 FILLER_22_279 ();
 sg13g2_fill_2 FILLER_22_283 ();
 sg13g2_decap_8 FILLER_22_290 ();
 sg13g2_decap_4 FILLER_22_301 ();
 sg13g2_decap_8 FILLER_22_317 ();
 sg13g2_decap_4 FILLER_22_324 ();
 sg13g2_fill_1 FILLER_22_358 ();
 sg13g2_fill_1 FILLER_22_373 ();
 sg13g2_fill_1 FILLER_22_379 ();
 sg13g2_fill_2 FILLER_22_401 ();
 sg13g2_fill_1 FILLER_22_403 ();
 sg13g2_decap_4 FILLER_23_0 ();
 sg13g2_fill_2 FILLER_23_4 ();
 sg13g2_fill_1 FILLER_23_16 ();
 sg13g2_decap_4 FILLER_23_22 ();
 sg13g2_fill_2 FILLER_23_26 ();
 sg13g2_fill_1 FILLER_23_33 ();
 sg13g2_fill_1 FILLER_23_37 ();
 sg13g2_fill_1 FILLER_23_47 ();
 sg13g2_fill_1 FILLER_23_53 ();
 sg13g2_decap_4 FILLER_23_81 ();
 sg13g2_fill_2 FILLER_23_85 ();
 sg13g2_decap_8 FILLER_23_121 ();
 sg13g2_decap_8 FILLER_23_128 ();
 sg13g2_fill_2 FILLER_23_135 ();
 sg13g2_fill_2 FILLER_23_146 ();
 sg13g2_fill_2 FILLER_23_153 ();
 sg13g2_fill_1 FILLER_23_155 ();
 sg13g2_fill_2 FILLER_23_165 ();
 sg13g2_fill_2 FILLER_23_172 ();
 sg13g2_fill_2 FILLER_23_196 ();
 sg13g2_fill_1 FILLER_23_198 ();
 sg13g2_decap_8 FILLER_23_203 ();
 sg13g2_fill_1 FILLER_23_210 ();
 sg13g2_fill_2 FILLER_23_220 ();
 sg13g2_decap_8 FILLER_23_243 ();
 sg13g2_decap_8 FILLER_23_264 ();
 sg13g2_decap_4 FILLER_23_271 ();
 sg13g2_fill_1 FILLER_23_275 ();
 sg13g2_decap_8 FILLER_23_280 ();
 sg13g2_fill_1 FILLER_23_287 ();
 sg13g2_decap_4 FILLER_23_298 ();
 sg13g2_fill_2 FILLER_23_329 ();
 sg13g2_fill_2 FILLER_23_344 ();
 sg13g2_fill_1 FILLER_23_346 ();
 sg13g2_fill_2 FILLER_23_363 ();
 sg13g2_fill_2 FILLER_23_370 ();
 sg13g2_fill_2 FILLER_23_377 ();
 sg13g2_fill_1 FILLER_23_379 ();
 sg13g2_fill_2 FILLER_23_394 ();
 sg13g2_fill_2 FILLER_24_0 ();
 sg13g2_fill_1 FILLER_24_2 ();
 sg13g2_fill_1 FILLER_24_29 ();
 sg13g2_decap_4 FILLER_24_49 ();
 sg13g2_fill_1 FILLER_24_58 ();
 sg13g2_fill_1 FILLER_24_64 ();
 sg13g2_fill_1 FILLER_24_74 ();
 sg13g2_decap_8 FILLER_24_102 ();
 sg13g2_decap_8 FILLER_24_109 ();
 sg13g2_decap_8 FILLER_24_116 ();
 sg13g2_fill_2 FILLER_24_123 ();
 sg13g2_fill_1 FILLER_24_125 ();
 sg13g2_decap_4 FILLER_24_149 ();
 sg13g2_fill_2 FILLER_24_153 ();
 sg13g2_fill_1 FILLER_24_159 ();
 sg13g2_fill_1 FILLER_24_165 ();
 sg13g2_fill_1 FILLER_24_194 ();
 sg13g2_decap_8 FILLER_24_209 ();
 sg13g2_decap_4 FILLER_24_216 ();
 sg13g2_fill_1 FILLER_24_220 ();
 sg13g2_decap_4 FILLER_24_230 ();
 sg13g2_decap_8 FILLER_24_238 ();
 sg13g2_decap_8 FILLER_24_245 ();
 sg13g2_fill_2 FILLER_24_252 ();
 sg13g2_fill_1 FILLER_24_254 ();
 sg13g2_decap_4 FILLER_24_259 ();
 sg13g2_decap_8 FILLER_24_267 ();
 sg13g2_decap_4 FILLER_24_274 ();
 sg13g2_fill_1 FILLER_24_278 ();
 sg13g2_decap_8 FILLER_24_284 ();
 sg13g2_decap_8 FILLER_24_291 ();
 sg13g2_fill_1 FILLER_24_312 ();
 sg13g2_decap_8 FILLER_24_318 ();
 sg13g2_decap_4 FILLER_24_330 ();
 sg13g2_decap_8 FILLER_24_339 ();
 sg13g2_decap_4 FILLER_24_346 ();
 sg13g2_decap_8 FILLER_24_360 ();
 sg13g2_decap_8 FILLER_24_367 ();
 sg13g2_fill_2 FILLER_24_374 ();
 sg13g2_fill_1 FILLER_24_376 ();
 sg13g2_fill_1 FILLER_24_385 ();
 sg13g2_decap_4 FILLER_24_396 ();
 sg13g2_fill_2 FILLER_24_404 ();
 sg13g2_fill_1 FILLER_24_429 ();
 sg13g2_decap_4 FILLER_25_0 ();
 sg13g2_fill_1 FILLER_25_4 ();
 sg13g2_fill_2 FILLER_25_25 ();
 sg13g2_fill_1 FILLER_25_27 ();
 sg13g2_fill_2 FILLER_25_31 ();
 sg13g2_fill_2 FILLER_25_53 ();
 sg13g2_fill_1 FILLER_25_55 ();
 sg13g2_fill_1 FILLER_25_62 ();
 sg13g2_fill_1 FILLER_25_68 ();
 sg13g2_fill_1 FILLER_25_73 ();
 sg13g2_fill_1 FILLER_25_97 ();
 sg13g2_decap_8 FILLER_25_107 ();
 sg13g2_fill_1 FILLER_25_114 ();
 sg13g2_decap_4 FILLER_25_123 ();
 sg13g2_fill_1 FILLER_25_127 ();
 sg13g2_fill_1 FILLER_25_133 ();
 sg13g2_fill_2 FILLER_25_191 ();
 sg13g2_fill_1 FILLER_25_193 ();
 sg13g2_decap_4 FILLER_25_224 ();
 sg13g2_fill_1 FILLER_25_228 ();
 sg13g2_fill_1 FILLER_25_239 ();
 sg13g2_decap_4 FILLER_25_251 ();
 sg13g2_fill_1 FILLER_25_255 ();
 sg13g2_fill_1 FILLER_25_286 ();
 sg13g2_decap_8 FILLER_25_291 ();
 sg13g2_decap_4 FILLER_25_298 ();
 sg13g2_fill_1 FILLER_25_321 ();
 sg13g2_decap_4 FILLER_25_332 ();
 sg13g2_fill_1 FILLER_25_342 ();
 sg13g2_fill_2 FILLER_25_351 ();
 sg13g2_fill_1 FILLER_25_353 ();
 sg13g2_decap_8 FILLER_25_388 ();
 sg13g2_decap_4 FILLER_25_395 ();
 sg13g2_fill_2 FILLER_25_399 ();
 sg13g2_decap_4 FILLER_25_405 ();
 sg13g2_fill_1 FILLER_25_409 ();
 sg13g2_fill_1 FILLER_25_414 ();
 sg13g2_decap_8 FILLER_25_423 ();
 sg13g2_decap_4 FILLER_26_0 ();
 sg13g2_fill_1 FILLER_26_4 ();
 sg13g2_fill_1 FILLER_26_19 ();
 sg13g2_decap_4 FILLER_26_32 ();
 sg13g2_fill_1 FILLER_26_41 ();
 sg13g2_fill_1 FILLER_26_47 ();
 sg13g2_fill_1 FILLER_26_53 ();
 sg13g2_fill_2 FILLER_26_60 ();
 sg13g2_decap_4 FILLER_26_73 ();
 sg13g2_fill_2 FILLER_26_77 ();
 sg13g2_fill_2 FILLER_26_84 ();
 sg13g2_fill_2 FILLER_26_91 ();
 sg13g2_fill_1 FILLER_26_93 ();
 sg13g2_decap_4 FILLER_26_99 ();
 sg13g2_fill_2 FILLER_26_107 ();
 sg13g2_fill_1 FILLER_26_109 ();
 sg13g2_fill_2 FILLER_26_132 ();
 sg13g2_fill_1 FILLER_26_142 ();
 sg13g2_fill_1 FILLER_26_152 ();
 sg13g2_fill_2 FILLER_26_158 ();
 sg13g2_fill_2 FILLER_26_164 ();
 sg13g2_decap_4 FILLER_26_170 ();
 sg13g2_fill_2 FILLER_26_174 ();
 sg13g2_fill_2 FILLER_26_188 ();
 sg13g2_fill_1 FILLER_26_190 ();
 sg13g2_fill_2 FILLER_26_196 ();
 sg13g2_decap_8 FILLER_26_229 ();
 sg13g2_fill_2 FILLER_26_236 ();
 sg13g2_fill_1 FILLER_26_298 ();
 sg13g2_fill_1 FILLER_26_348 ();
 sg13g2_fill_2 FILLER_26_379 ();
 sg13g2_fill_2 FILLER_26_386 ();
 sg13g2_fill_2 FILLER_26_395 ();
 sg13g2_fill_2 FILLER_26_401 ();
 sg13g2_fill_1 FILLER_26_403 ();
 sg13g2_decap_8 FILLER_27_0 ();
 sg13g2_decap_8 FILLER_27_7 ();
 sg13g2_decap_4 FILLER_27_14 ();
 sg13g2_fill_2 FILLER_27_18 ();
 sg13g2_decap_8 FILLER_27_23 ();
 sg13g2_decap_8 FILLER_27_30 ();
 sg13g2_decap_4 FILLER_27_37 ();
 sg13g2_fill_1 FILLER_27_41 ();
 sg13g2_decap_8 FILLER_27_46 ();
 sg13g2_decap_8 FILLER_27_53 ();
 sg13g2_decap_4 FILLER_27_60 ();
 sg13g2_decap_8 FILLER_27_73 ();
 sg13g2_decap_8 FILLER_27_80 ();
 sg13g2_decap_4 FILLER_27_87 ();
 sg13g2_decap_4 FILLER_27_96 ();
 sg13g2_fill_2 FILLER_27_100 ();
 sg13g2_decap_8 FILLER_27_107 ();
 sg13g2_fill_1 FILLER_27_114 ();
 sg13g2_fill_2 FILLER_27_139 ();
 sg13g2_fill_1 FILLER_27_150 ();
 sg13g2_fill_1 FILLER_27_159 ();
 sg13g2_fill_2 FILLER_27_191 ();
 sg13g2_fill_1 FILLER_27_193 ();
 sg13g2_fill_2 FILLER_27_257 ();
 sg13g2_fill_1 FILLER_27_274 ();
 sg13g2_fill_1 FILLER_27_285 ();
 sg13g2_fill_2 FILLER_27_291 ();
 sg13g2_fill_1 FILLER_27_293 ();
 sg13g2_fill_2 FILLER_27_299 ();
 sg13g2_fill_1 FILLER_27_301 ();
 sg13g2_fill_2 FILLER_27_311 ();
 sg13g2_fill_1 FILLER_27_316 ();
 sg13g2_fill_2 FILLER_27_322 ();
 sg13g2_decap_8 FILLER_27_328 ();
 sg13g2_fill_1 FILLER_27_339 ();
 sg13g2_fill_2 FILLER_27_344 ();
 sg13g2_fill_2 FILLER_27_350 ();
 sg13g2_fill_1 FILLER_27_352 ();
 sg13g2_fill_2 FILLER_27_357 ();
 sg13g2_fill_1 FILLER_27_359 ();
 sg13g2_fill_2 FILLER_27_365 ();
 sg13g2_fill_1 FILLER_27_367 ();
 sg13g2_decap_8 FILLER_27_373 ();
 sg13g2_decap_8 FILLER_27_380 ();
 sg13g2_fill_1 FILLER_27_387 ();
 sg13g2_decap_4 FILLER_27_418 ();
 sg13g2_fill_1 FILLER_27_422 ();
 sg13g2_fill_2 FILLER_27_427 ();
 sg13g2_fill_1 FILLER_27_429 ();
 sg13g2_decap_8 FILLER_28_0 ();
 sg13g2_fill_1 FILLER_28_7 ();
 sg13g2_fill_2 FILLER_28_13 ();
 sg13g2_fill_1 FILLER_28_15 ();
 sg13g2_decap_4 FILLER_28_29 ();
 sg13g2_fill_1 FILLER_28_33 ();
 sg13g2_fill_1 FILLER_28_39 ();
 sg13g2_fill_2 FILLER_28_49 ();
 sg13g2_fill_1 FILLER_28_51 ();
 sg13g2_fill_2 FILLER_28_65 ();
 sg13g2_fill_1 FILLER_28_72 ();
 sg13g2_decap_8 FILLER_28_78 ();
 sg13g2_decap_8 FILLER_28_85 ();
 sg13g2_decap_4 FILLER_28_92 ();
 sg13g2_fill_1 FILLER_28_96 ();
 sg13g2_decap_4 FILLER_28_106 ();
 sg13g2_fill_2 FILLER_28_110 ();
 sg13g2_fill_1 FILLER_28_123 ();
 sg13g2_decap_4 FILLER_28_129 ();
 sg13g2_fill_1 FILLER_28_133 ();
 sg13g2_fill_2 FILLER_28_142 ();
 sg13g2_decap_4 FILLER_28_149 ();
 sg13g2_fill_1 FILLER_28_171 ();
 sg13g2_fill_2 FILLER_28_176 ();
 sg13g2_fill_1 FILLER_28_178 ();
 sg13g2_fill_1 FILLER_28_183 ();
 sg13g2_fill_1 FILLER_28_214 ();
 sg13g2_decap_8 FILLER_28_219 ();
 sg13g2_fill_2 FILLER_28_233 ();
 sg13g2_fill_1 FILLER_28_235 ();
 sg13g2_decap_4 FILLER_28_249 ();
 sg13g2_fill_2 FILLER_28_266 ();
 sg13g2_fill_1 FILLER_28_273 ();
 sg13g2_fill_2 FILLER_28_279 ();
 sg13g2_fill_1 FILLER_28_281 ();
 sg13g2_decap_8 FILLER_28_291 ();
 sg13g2_decap_8 FILLER_28_298 ();
 sg13g2_decap_8 FILLER_28_324 ();
 sg13g2_decap_8 FILLER_28_331 ();
 sg13g2_decap_4 FILLER_28_338 ();
 sg13g2_decap_8 FILLER_28_347 ();
 sg13g2_fill_2 FILLER_28_354 ();
 sg13g2_decap_4 FILLER_28_368 ();
 sg13g2_fill_1 FILLER_28_372 ();
 sg13g2_decap_4 FILLER_29_45 ();
 sg13g2_decap_8 FILLER_29_54 ();
 sg13g2_fill_2 FILLER_29_65 ();
 sg13g2_fill_1 FILLER_29_72 ();
 sg13g2_fill_1 FILLER_29_78 ();
 sg13g2_fill_1 FILLER_29_89 ();
 sg13g2_decap_8 FILLER_29_103 ();
 sg13g2_decap_4 FILLER_29_110 ();
 sg13g2_fill_2 FILLER_29_126 ();
 sg13g2_fill_1 FILLER_29_128 ();
 sg13g2_fill_2 FILLER_29_139 ();
 sg13g2_decap_8 FILLER_29_158 ();
 sg13g2_fill_1 FILLER_29_173 ();
 sg13g2_decap_8 FILLER_29_178 ();
 sg13g2_decap_8 FILLER_29_185 ();
 sg13g2_decap_8 FILLER_29_196 ();
 sg13g2_decap_8 FILLER_29_203 ();
 sg13g2_decap_4 FILLER_29_210 ();
 sg13g2_decap_8 FILLER_29_233 ();
 sg13g2_decap_8 FILLER_29_240 ();
 sg13g2_decap_8 FILLER_29_247 ();
 sg13g2_fill_2 FILLER_29_254 ();
 sg13g2_decap_8 FILLER_29_289 ();
 sg13g2_decap_4 FILLER_29_296 ();
 sg13g2_fill_1 FILLER_29_300 ();
 sg13g2_fill_1 FILLER_29_306 ();
 sg13g2_decap_4 FILLER_29_316 ();
 sg13g2_fill_2 FILLER_29_320 ();
 sg13g2_decap_8 FILLER_29_356 ();
 sg13g2_decap_8 FILLER_29_373 ();
 sg13g2_decap_4 FILLER_29_380 ();
 sg13g2_fill_2 FILLER_29_384 ();
 sg13g2_fill_1 FILLER_29_414 ();
 sg13g2_decap_8 FILLER_29_419 ();
 sg13g2_decap_4 FILLER_29_426 ();
 sg13g2_fill_1 FILLER_30_0 ();
 sg13g2_decap_4 FILLER_30_36 ();
 sg13g2_fill_1 FILLER_30_45 ();
 sg13g2_fill_2 FILLER_30_72 ();
 sg13g2_fill_1 FILLER_30_74 ();
 sg13g2_decap_8 FILLER_30_80 ();
 sg13g2_decap_8 FILLER_30_87 ();
 sg13g2_fill_2 FILLER_30_103 ();
 sg13g2_fill_2 FILLER_30_150 ();
 sg13g2_fill_1 FILLER_30_152 ();
 sg13g2_fill_2 FILLER_30_161 ();
 sg13g2_decap_8 FILLER_30_205 ();
 sg13g2_decap_8 FILLER_30_212 ();
 sg13g2_fill_2 FILLER_30_219 ();
 sg13g2_decap_8 FILLER_30_226 ();
 sg13g2_decap_4 FILLER_30_233 ();
 sg13g2_fill_2 FILLER_30_237 ();
 sg13g2_decap_8 FILLER_30_243 ();
 sg13g2_decap_4 FILLER_30_250 ();
 sg13g2_fill_2 FILLER_30_276 ();
 sg13g2_fill_1 FILLER_30_315 ();
 sg13g2_decap_8 FILLER_30_342 ();
 sg13g2_decap_8 FILLER_30_349 ();
 sg13g2_decap_8 FILLER_30_356 ();
 sg13g2_fill_2 FILLER_30_363 ();
 sg13g2_fill_1 FILLER_30_403 ();
 sg13g2_decap_8 FILLER_31_0 ();
 sg13g2_fill_1 FILLER_31_16 ();
 sg13g2_fill_1 FILLER_31_26 ();
 sg13g2_decap_8 FILLER_31_45 ();
 sg13g2_fill_2 FILLER_31_52 ();
 sg13g2_fill_1 FILLER_31_54 ();
 sg13g2_decap_4 FILLER_31_68 ();
 sg13g2_fill_1 FILLER_31_72 ();
 sg13g2_decap_8 FILLER_31_83 ();
 sg13g2_decap_4 FILLER_31_90 ();
 sg13g2_fill_2 FILLER_31_94 ();
 sg13g2_decap_4 FILLER_31_100 ();
 sg13g2_fill_1 FILLER_31_104 ();
 sg13g2_fill_1 FILLER_31_125 ();
 sg13g2_fill_2 FILLER_31_136 ();
 sg13g2_fill_1 FILLER_31_138 ();
 sg13g2_fill_2 FILLER_31_165 ();
 sg13g2_fill_1 FILLER_31_171 ();
 sg13g2_fill_2 FILLER_31_176 ();
 sg13g2_fill_1 FILLER_31_178 ();
 sg13g2_fill_2 FILLER_31_197 ();
 sg13g2_fill_1 FILLER_31_269 ();
 sg13g2_fill_2 FILLER_31_277 ();
 sg13g2_fill_1 FILLER_31_279 ();
 sg13g2_decap_4 FILLER_31_285 ();
 sg13g2_fill_1 FILLER_31_289 ();
 sg13g2_fill_2 FILLER_31_294 ();
 sg13g2_fill_2 FILLER_31_353 ();
 sg13g2_decap_8 FILLER_31_360 ();
 sg13g2_decap_8 FILLER_31_367 ();
 sg13g2_fill_2 FILLER_31_374 ();
 sg13g2_fill_1 FILLER_31_397 ();
 sg13g2_fill_1 FILLER_31_402 ();
 sg13g2_fill_1 FILLER_31_407 ();
 sg13g2_fill_2 FILLER_31_413 ();
 sg13g2_decap_8 FILLER_31_419 ();
 sg13g2_decap_4 FILLER_31_426 ();
 sg13g2_decap_4 FILLER_32_0 ();
 sg13g2_fill_1 FILLER_32_4 ();
 sg13g2_decap_8 FILLER_32_15 ();
 sg13g2_decap_8 FILLER_32_22 ();
 sg13g2_decap_8 FILLER_32_29 ();
 sg13g2_fill_1 FILLER_32_36 ();
 sg13g2_fill_2 FILLER_32_42 ();
 sg13g2_fill_2 FILLER_32_47 ();
 sg13g2_decap_8 FILLER_32_53 ();
 sg13g2_fill_1 FILLER_32_60 ();
 sg13g2_fill_2 FILLER_32_64 ();
 sg13g2_fill_1 FILLER_32_66 ();
 sg13g2_decap_8 FILLER_32_71 ();
 sg13g2_decap_8 FILLER_32_78 ();
 sg13g2_decap_8 FILLER_32_85 ();
 sg13g2_decap_4 FILLER_32_92 ();
 sg13g2_fill_2 FILLER_32_96 ();
 sg13g2_decap_8 FILLER_32_103 ();
 sg13g2_decap_4 FILLER_32_110 ();
 sg13g2_fill_1 FILLER_32_119 ();
 sg13g2_fill_2 FILLER_32_167 ();
 sg13g2_fill_2 FILLER_32_195 ();
 sg13g2_fill_1 FILLER_32_205 ();
 sg13g2_fill_1 FILLER_32_232 ();
 sg13g2_fill_1 FILLER_32_241 ();
 sg13g2_fill_1 FILLER_32_247 ();
 sg13g2_fill_1 FILLER_32_252 ();
 sg13g2_fill_1 FILLER_32_258 ();
 sg13g2_fill_1 FILLER_32_264 ();
 sg13g2_fill_1 FILLER_32_279 ();
 sg13g2_decap_8 FILLER_32_285 ();
 sg13g2_fill_2 FILLER_32_292 ();
 sg13g2_fill_1 FILLER_32_294 ();
 sg13g2_fill_1 FILLER_32_299 ();
 sg13g2_fill_1 FILLER_32_304 ();
 sg13g2_decap_8 FILLER_32_343 ();
 sg13g2_decap_8 FILLER_32_350 ();
 sg13g2_decap_8 FILLER_32_357 ();
 sg13g2_decap_8 FILLER_32_364 ();
 sg13g2_fill_2 FILLER_32_371 ();
 sg13g2_decap_4 FILLER_32_388 ();
 sg13g2_decap_4 FILLER_32_398 ();
 sg13g2_decap_4 FILLER_32_407 ();
 sg13g2_decap_8 FILLER_32_415 ();
 sg13g2_decap_8 FILLER_32_422 ();
 sg13g2_fill_1 FILLER_32_429 ();
 sg13g2_decap_8 FILLER_33_0 ();
 sg13g2_fill_2 FILLER_33_12 ();
 sg13g2_fill_1 FILLER_33_14 ();
 sg13g2_decap_4 FILLER_33_41 ();
 sg13g2_fill_1 FILLER_33_45 ();
 sg13g2_decap_4 FILLER_33_51 ();
 sg13g2_fill_2 FILLER_33_55 ();
 sg13g2_fill_2 FILLER_33_67 ();
 sg13g2_fill_1 FILLER_33_69 ();
 sg13g2_fill_1 FILLER_33_99 ();
 sg13g2_fill_2 FILLER_33_105 ();
 sg13g2_fill_1 FILLER_33_111 ();
 sg13g2_fill_2 FILLER_33_121 ();
 sg13g2_decap_8 FILLER_33_157 ();
 sg13g2_decap_8 FILLER_33_164 ();
 sg13g2_decap_4 FILLER_33_171 ();
 sg13g2_fill_1 FILLER_33_175 ();
 sg13g2_fill_2 FILLER_33_180 ();
 sg13g2_fill_1 FILLER_33_206 ();
 sg13g2_fill_2 FILLER_33_211 ();
 sg13g2_fill_2 FILLER_33_217 ();
 sg13g2_fill_2 FILLER_33_223 ();
 sg13g2_fill_1 FILLER_33_225 ();
 sg13g2_fill_2 FILLER_33_252 ();
 sg13g2_fill_1 FILLER_33_254 ();
 sg13g2_fill_2 FILLER_33_309 ();
 sg13g2_decap_8 FILLER_33_315 ();
 sg13g2_decap_4 FILLER_33_322 ();
 sg13g2_fill_2 FILLER_33_360 ();
 sg13g2_fill_1 FILLER_33_362 ();
 sg13g2_decap_4 FILLER_33_381 ();
 sg13g2_fill_1 FILLER_33_388 ();
 sg13g2_fill_2 FILLER_34_0 ();
 sg13g2_fill_1 FILLER_34_2 ();
 sg13g2_fill_1 FILLER_34_34 ();
 sg13g2_fill_1 FILLER_34_59 ();
 sg13g2_fill_1 FILLER_34_68 ();
 sg13g2_fill_1 FILLER_34_74 ();
 sg13g2_fill_1 FILLER_34_79 ();
 sg13g2_fill_1 FILLER_34_96 ();
 sg13g2_fill_1 FILLER_34_102 ();
 sg13g2_fill_1 FILLER_34_108 ();
 sg13g2_fill_2 FILLER_34_114 ();
 sg13g2_decap_4 FILLER_34_121 ();
 sg13g2_fill_2 FILLER_34_125 ();
 sg13g2_fill_2 FILLER_34_132 ();
 sg13g2_fill_1 FILLER_34_134 ();
 sg13g2_decap_8 FILLER_34_151 ();
 sg13g2_decap_4 FILLER_34_158 ();
 sg13g2_fill_1 FILLER_34_167 ();
 sg13g2_fill_2 FILLER_34_173 ();
 sg13g2_decap_8 FILLER_34_199 ();
 sg13g2_decap_8 FILLER_34_216 ();
 sg13g2_decap_8 FILLER_34_223 ();
 sg13g2_decap_8 FILLER_34_230 ();
 sg13g2_decap_4 FILLER_34_237 ();
 sg13g2_fill_2 FILLER_34_241 ();
 sg13g2_fill_2 FILLER_34_247 ();
 sg13g2_fill_1 FILLER_34_249 ();
 sg13g2_fill_2 FILLER_34_254 ();
 sg13g2_fill_1 FILLER_34_256 ();
 sg13g2_fill_1 FILLER_34_272 ();
 sg13g2_fill_1 FILLER_34_292 ();
 sg13g2_decap_4 FILLER_34_297 ();
 sg13g2_fill_2 FILLER_34_315 ();
 sg13g2_fill_1 FILLER_34_317 ();
 sg13g2_fill_1 FILLER_34_322 ();
 sg13g2_decap_8 FILLER_34_328 ();
 sg13g2_fill_2 FILLER_34_335 ();
 sg13g2_fill_1 FILLER_34_337 ();
 sg13g2_fill_2 FILLER_34_377 ();
 sg13g2_fill_1 FILLER_34_379 ();
 sg13g2_fill_2 FILLER_34_398 ();
 sg13g2_fill_2 FILLER_35_0 ();
 sg13g2_fill_2 FILLER_35_26 ();
 sg13g2_decap_4 FILLER_35_32 ();
 sg13g2_fill_1 FILLER_35_36 ();
 sg13g2_fill_1 FILLER_35_47 ();
 sg13g2_fill_2 FILLER_35_63 ();
 sg13g2_fill_1 FILLER_35_70 ();
 sg13g2_fill_2 FILLER_35_84 ();
 sg13g2_fill_1 FILLER_35_86 ();
 sg13g2_decap_8 FILLER_35_113 ();
 sg13g2_decap_8 FILLER_35_120 ();
 sg13g2_fill_1 FILLER_35_134 ();
 sg13g2_decap_8 FILLER_35_143 ();
 sg13g2_fill_2 FILLER_35_150 ();
 sg13g2_fill_1 FILLER_35_152 ();
 sg13g2_fill_1 FILLER_35_171 ();
 sg13g2_decap_8 FILLER_35_177 ();
 sg13g2_fill_2 FILLER_35_184 ();
 sg13g2_decap_8 FILLER_35_191 ();
 sg13g2_decap_8 FILLER_35_198 ();
 sg13g2_decap_4 FILLER_35_205 ();
 sg13g2_decap_4 FILLER_35_213 ();
 sg13g2_fill_1 FILLER_35_217 ();
 sg13g2_decap_4 FILLER_35_222 ();
 sg13g2_decap_8 FILLER_35_231 ();
 sg13g2_decap_8 FILLER_35_238 ();
 sg13g2_fill_1 FILLER_35_245 ();
 sg13g2_fill_2 FILLER_35_250 ();
 sg13g2_decap_8 FILLER_35_292 ();
 sg13g2_fill_2 FILLER_35_299 ();
 sg13g2_fill_1 FILLER_35_301 ();
 sg13g2_decap_4 FILLER_35_306 ();
 sg13g2_fill_2 FILLER_35_310 ();
 sg13g2_fill_1 FILLER_35_357 ();
 sg13g2_fill_1 FILLER_35_367 ();
 sg13g2_fill_2 FILLER_35_373 ();
 sg13g2_fill_2 FILLER_35_379 ();
 sg13g2_decap_8 FILLER_35_386 ();
 sg13g2_decap_8 FILLER_35_403 ();
 sg13g2_fill_2 FILLER_35_414 ();
 sg13g2_fill_2 FILLER_35_420 ();
 sg13g2_fill_1 FILLER_35_422 ();
 sg13g2_fill_2 FILLER_35_427 ();
 sg13g2_fill_1 FILLER_35_429 ();
 sg13g2_decap_8 FILLER_36_0 ();
 sg13g2_decap_8 FILLER_36_11 ();
 sg13g2_decap_4 FILLER_36_31 ();
 sg13g2_fill_1 FILLER_36_35 ();
 sg13g2_fill_2 FILLER_36_59 ();
 sg13g2_fill_1 FILLER_36_70 ();
 sg13g2_fill_1 FILLER_36_83 ();
 sg13g2_decap_8 FILLER_36_89 ();
 sg13g2_decap_4 FILLER_36_96 ();
 sg13g2_fill_1 FILLER_36_100 ();
 sg13g2_decap_4 FILLER_36_106 ();
 sg13g2_fill_2 FILLER_36_110 ();
 sg13g2_decap_8 FILLER_36_119 ();
 sg13g2_decap_8 FILLER_36_126 ();
 sg13g2_fill_2 FILLER_36_133 ();
 sg13g2_fill_1 FILLER_36_177 ();
 sg13g2_decap_8 FILLER_36_190 ();
 sg13g2_decap_4 FILLER_36_197 ();
 sg13g2_fill_1 FILLER_36_201 ();
 sg13g2_fill_2 FILLER_36_232 ();
 sg13g2_fill_2 FILLER_36_244 ();
 sg13g2_decap_4 FILLER_36_250 ();
 sg13g2_fill_2 FILLER_36_254 ();
 sg13g2_decap_8 FILLER_36_260 ();
 sg13g2_fill_1 FILLER_36_267 ();
 sg13g2_fill_1 FILLER_36_281 ();
 sg13g2_decap_8 FILLER_36_286 ();
 sg13g2_decap_4 FILLER_36_293 ();
 sg13g2_fill_1 FILLER_36_297 ();
 sg13g2_fill_1 FILLER_36_311 ();
 sg13g2_fill_2 FILLER_36_342 ();
 sg13g2_fill_1 FILLER_36_349 ();
 sg13g2_fill_1 FILLER_36_354 ();
 sg13g2_fill_2 FILLER_36_361 ();
 sg13g2_fill_1 FILLER_36_368 ();
 sg13g2_decap_4 FILLER_36_374 ();
 sg13g2_fill_1 FILLER_36_378 ();
 sg13g2_fill_1 FILLER_36_388 ();
 sg13g2_decap_4 FILLER_36_393 ();
 sg13g2_fill_1 FILLER_36_402 ();
 sg13g2_decap_8 FILLER_36_408 ();
 sg13g2_decap_8 FILLER_36_415 ();
 sg13g2_decap_8 FILLER_36_422 ();
 sg13g2_fill_1 FILLER_36_429 ();
 sg13g2_fill_1 FILLER_37_26 ();
 sg13g2_fill_1 FILLER_37_31 ();
 sg13g2_fill_1 FILLER_37_46 ();
 sg13g2_fill_1 FILLER_37_66 ();
 sg13g2_fill_1 FILLER_37_77 ();
 sg13g2_decap_8 FILLER_37_83 ();
 sg13g2_decap_4 FILLER_37_90 ();
 sg13g2_fill_1 FILLER_37_94 ();
 sg13g2_fill_1 FILLER_37_99 ();
 sg13g2_fill_1 FILLER_37_117 ();
 sg13g2_fill_2 FILLER_37_132 ();
 sg13g2_decap_4 FILLER_37_143 ();
 sg13g2_fill_2 FILLER_37_152 ();
 sg13g2_fill_1 FILLER_37_154 ();
 sg13g2_fill_1 FILLER_37_183 ();
 sg13g2_fill_1 FILLER_37_210 ();
 sg13g2_fill_2 FILLER_37_237 ();
 sg13g2_fill_1 FILLER_37_269 ();
 sg13g2_fill_2 FILLER_37_278 ();
 sg13g2_decap_8 FILLER_37_292 ();
 sg13g2_fill_2 FILLER_37_316 ();
 sg13g2_fill_1 FILLER_37_318 ();
 sg13g2_decap_8 FILLER_37_323 ();
 sg13g2_decap_8 FILLER_37_335 ();
 sg13g2_fill_2 FILLER_37_342 ();
 sg13g2_fill_1 FILLER_37_344 ();
 sg13g2_fill_1 FILLER_37_383 ();
 sg13g2_fill_2 FILLER_37_417 ();
 sg13g2_decap_4 FILLER_37_424 ();
 sg13g2_fill_2 FILLER_37_428 ();
 sg13g2_decap_4 FILLER_38_0 ();
 sg13g2_fill_1 FILLER_38_4 ();
 sg13g2_fill_1 FILLER_38_15 ();
 sg13g2_decap_8 FILLER_38_26 ();
 sg13g2_fill_2 FILLER_38_37 ();
 sg13g2_fill_1 FILLER_38_43 ();
 sg13g2_fill_1 FILLER_38_54 ();
 sg13g2_fill_1 FILLER_38_59 ();
 sg13g2_fill_1 FILLER_38_73 ();
 sg13g2_fill_2 FILLER_38_78 ();
 sg13g2_fill_2 FILLER_38_85 ();
 sg13g2_fill_2 FILLER_38_99 ();
 sg13g2_fill_1 FILLER_38_101 ();
 sg13g2_fill_1 FILLER_38_121 ();
 sg13g2_fill_1 FILLER_38_127 ();
 sg13g2_decap_8 FILLER_38_141 ();
 sg13g2_decap_8 FILLER_38_148 ();
 sg13g2_fill_2 FILLER_38_155 ();
 sg13g2_fill_2 FILLER_38_170 ();
 sg13g2_decap_4 FILLER_38_197 ();
 sg13g2_fill_2 FILLER_38_201 ();
 sg13g2_fill_1 FILLER_38_234 ();
 sg13g2_decap_8 FILLER_38_243 ();
 sg13g2_decap_8 FILLER_38_250 ();
 sg13g2_decap_4 FILLER_38_257 ();
 sg13g2_fill_2 FILLER_38_266 ();
 sg13g2_fill_2 FILLER_38_290 ();
 sg13g2_fill_1 FILLER_38_292 ();
 sg13g2_decap_8 FILLER_38_297 ();
 sg13g2_fill_1 FILLER_38_304 ();
 sg13g2_decap_8 FILLER_38_310 ();
 sg13g2_decap_4 FILLER_38_322 ();
 sg13g2_fill_1 FILLER_38_326 ();
 sg13g2_decap_8 FILLER_38_353 ();
 sg13g2_fill_1 FILLER_38_360 ();
 sg13g2_fill_1 FILLER_38_376 ();
 sg13g2_fill_1 FILLER_38_381 ();
 sg13g2_fill_1 FILLER_38_387 ();
 sg13g2_fill_1 FILLER_38_397 ();
 sg13g2_fill_1 FILLER_38_403 ();
 sg13g2_decap_4 FILLER_39_0 ();
 sg13g2_fill_1 FILLER_39_4 ();
 sg13g2_decap_4 FILLER_39_20 ();
 sg13g2_fill_1 FILLER_39_24 ();
 sg13g2_decap_4 FILLER_39_30 ();
 sg13g2_fill_1 FILLER_39_38 ();
 sg13g2_fill_2 FILLER_39_67 ();
 sg13g2_fill_1 FILLER_39_78 ();
 sg13g2_decap_4 FILLER_39_83 ();
 sg13g2_fill_1 FILLER_39_87 ();
 sg13g2_fill_1 FILLER_39_102 ();
 sg13g2_fill_1 FILLER_39_108 ();
 sg13g2_fill_1 FILLER_39_120 ();
 sg13g2_decap_8 FILLER_39_137 ();
 sg13g2_fill_1 FILLER_39_144 ();
 sg13g2_fill_2 FILLER_39_150 ();
 sg13g2_decap_4 FILLER_39_161 ();
 sg13g2_fill_1 FILLER_39_168 ();
 sg13g2_decap_8 FILLER_39_181 ();
 sg13g2_fill_2 FILLER_39_188 ();
 sg13g2_decap_8 FILLER_39_193 ();
 sg13g2_decap_8 FILLER_39_200 ();
 sg13g2_fill_2 FILLER_39_207 ();
 sg13g2_fill_1 FILLER_39_223 ();
 sg13g2_decap_8 FILLER_39_253 ();
 sg13g2_decap_8 FILLER_39_260 ();
 sg13g2_fill_1 FILLER_39_267 ();
 sg13g2_decap_4 FILLER_39_290 ();
 sg13g2_decap_8 FILLER_39_306 ();
 sg13g2_decap_8 FILLER_39_313 ();
 sg13g2_decap_8 FILLER_39_320 ();
 sg13g2_fill_2 FILLER_39_327 ();
 sg13g2_decap_4 FILLER_39_338 ();
 sg13g2_fill_1 FILLER_39_342 ();
 sg13g2_decap_8 FILLER_40_0 ();
 sg13g2_decap_8 FILLER_40_17 ();
 sg13g2_decap_8 FILLER_40_24 ();
 sg13g2_decap_4 FILLER_40_31 ();
 sg13g2_fill_1 FILLER_40_38 ();
 sg13g2_fill_2 FILLER_40_64 ();
 sg13g2_decap_8 FILLER_40_69 ();
 sg13g2_fill_1 FILLER_40_76 ();
 sg13g2_fill_1 FILLER_40_85 ();
 sg13g2_decap_8 FILLER_40_96 ();
 sg13g2_fill_2 FILLER_40_103 ();
 sg13g2_fill_1 FILLER_40_105 ();
 sg13g2_fill_2 FILLER_40_109 ();
 sg13g2_fill_1 FILLER_40_111 ();
 sg13g2_decap_4 FILLER_40_119 ();
 sg13g2_decap_8 FILLER_40_130 ();
 sg13g2_decap_4 FILLER_40_137 ();
 sg13g2_fill_1 FILLER_40_141 ();
 sg13g2_decap_8 FILLER_40_173 ();
 sg13g2_decap_8 FILLER_40_180 ();
 sg13g2_decap_4 FILLER_40_187 ();
 sg13g2_fill_1 FILLER_40_191 ();
 sg13g2_fill_2 FILLER_40_229 ();
 sg13g2_decap_4 FILLER_40_239 ();
 sg13g2_decap_4 FILLER_40_248 ();
 sg13g2_fill_1 FILLER_40_252 ();
 sg13g2_fill_1 FILLER_40_256 ();
 sg13g2_fill_1 FILLER_40_262 ();
 sg13g2_fill_1 FILLER_40_268 ();
 sg13g2_decap_8 FILLER_40_313 ();
 sg13g2_decap_4 FILLER_40_320 ();
 sg13g2_fill_2 FILLER_40_324 ();
 sg13g2_fill_1 FILLER_40_342 ();
 sg13g2_fill_1 FILLER_40_348 ();
 sg13g2_fill_1 FILLER_40_366 ();
 sg13g2_fill_1 FILLER_40_372 ();
 sg13g2_fill_1 FILLER_40_377 ();
 sg13g2_fill_1 FILLER_40_425 ();
 sg13g2_fill_1 FILLER_41_36 ();
 sg13g2_fill_1 FILLER_41_48 ();
 sg13g2_decap_8 FILLER_41_59 ();
 sg13g2_fill_1 FILLER_41_70 ();
 sg13g2_fill_2 FILLER_41_78 ();
 sg13g2_fill_1 FILLER_41_80 ();
 sg13g2_decap_8 FILLER_41_85 ();
 sg13g2_decap_8 FILLER_41_92 ();
 sg13g2_fill_1 FILLER_41_99 ();
 sg13g2_decap_8 FILLER_41_111 ();
 sg13g2_decap_8 FILLER_41_118 ();
 sg13g2_fill_2 FILLER_41_125 ();
 sg13g2_fill_2 FILLER_41_147 ();
 sg13g2_fill_1 FILLER_41_153 ();
 sg13g2_fill_1 FILLER_41_176 ();
 sg13g2_decap_8 FILLER_41_184 ();
 sg13g2_decap_8 FILLER_41_191 ();
 sg13g2_fill_1 FILLER_41_198 ();
 sg13g2_fill_2 FILLER_41_212 ();
 sg13g2_fill_1 FILLER_41_214 ();
 sg13g2_decap_8 FILLER_41_230 ();
 sg13g2_fill_2 FILLER_41_237 ();
 sg13g2_fill_2 FILLER_41_256 ();
 sg13g2_fill_1 FILLER_41_263 ();
 sg13g2_fill_1 FILLER_41_286 ();
 sg13g2_decap_8 FILLER_41_313 ();
 sg13g2_fill_2 FILLER_41_320 ();
 sg13g2_fill_1 FILLER_41_322 ();
 sg13g2_fill_2 FILLER_41_349 ();
 sg13g2_fill_1 FILLER_41_351 ();
 sg13g2_decap_4 FILLER_41_357 ();
 sg13g2_fill_1 FILLER_41_361 ();
 sg13g2_decap_4 FILLER_41_374 ();
 sg13g2_fill_1 FILLER_41_397 ();
 sg13g2_fill_2 FILLER_41_403 ();
 sg13g2_fill_2 FILLER_41_410 ();
 sg13g2_fill_2 FILLER_41_416 ();
 sg13g2_fill_1 FILLER_41_418 ();
 sg13g2_decap_8 FILLER_41_423 ();
 sg13g2_decap_4 FILLER_42_0 ();
 sg13g2_fill_1 FILLER_42_8 ();
 sg13g2_fill_2 FILLER_42_42 ();
 sg13g2_fill_1 FILLER_42_44 ();
 sg13g2_fill_2 FILLER_42_59 ();
 sg13g2_fill_1 FILLER_42_61 ();
 sg13g2_fill_1 FILLER_42_70 ();
 sg13g2_fill_2 FILLER_42_76 ();
 sg13g2_fill_2 FILLER_42_86 ();
 sg13g2_fill_1 FILLER_42_88 ();
 sg13g2_fill_2 FILLER_42_96 ();
 sg13g2_fill_1 FILLER_42_98 ();
 sg13g2_decap_8 FILLER_42_112 ();
 sg13g2_fill_2 FILLER_42_119 ();
 sg13g2_fill_2 FILLER_42_154 ();
 sg13g2_fill_1 FILLER_42_156 ();
 sg13g2_decap_8 FILLER_42_197 ();
 sg13g2_fill_2 FILLER_42_204 ();
 sg13g2_decap_8 FILLER_42_210 ();
 sg13g2_decap_4 FILLER_42_217 ();
 sg13g2_fill_1 FILLER_42_221 ();
 sg13g2_decap_8 FILLER_42_226 ();
 sg13g2_decap_8 FILLER_42_233 ();
 sg13g2_fill_2 FILLER_42_240 ();
 sg13g2_fill_1 FILLER_42_242 ();
 sg13g2_decap_4 FILLER_42_248 ();
 sg13g2_fill_2 FILLER_42_252 ();
 sg13g2_decap_4 FILLER_42_278 ();
 sg13g2_decap_4 FILLER_42_308 ();
 sg13g2_fill_1 FILLER_42_312 ();
 sg13g2_decap_8 FILLER_42_317 ();
 sg13g2_fill_1 FILLER_42_324 ();
 sg13g2_fill_1 FILLER_42_330 ();
 sg13g2_decap_8 FILLER_42_343 ();
 sg13g2_fill_2 FILLER_42_350 ();
 sg13g2_decap_8 FILLER_42_369 ();
 sg13g2_decap_4 FILLER_42_376 ();
 sg13g2_decap_8 FILLER_42_395 ();
 sg13g2_decap_8 FILLER_42_402 ();
 sg13g2_decap_8 FILLER_42_409 ();
 sg13g2_decap_8 FILLER_42_416 ();
 sg13g2_decap_8 FILLER_42_423 ();
 sg13g2_decap_8 FILLER_43_0 ();
 sg13g2_decap_8 FILLER_43_7 ();
 sg13g2_fill_2 FILLER_43_14 ();
 sg13g2_fill_2 FILLER_43_20 ();
 sg13g2_decap_8 FILLER_43_35 ();
 sg13g2_fill_1 FILLER_43_46 ();
 sg13g2_fill_2 FILLER_43_55 ();
 sg13g2_fill_1 FILLER_43_57 ();
 sg13g2_fill_1 FILLER_43_102 ();
 sg13g2_decap_8 FILLER_43_108 ();
 sg13g2_decap_8 FILLER_43_115 ();
 sg13g2_decap_4 FILLER_43_122 ();
 sg13g2_fill_2 FILLER_43_126 ();
 sg13g2_fill_2 FILLER_43_133 ();
 sg13g2_decap_4 FILLER_43_140 ();
 sg13g2_fill_1 FILLER_43_149 ();
 sg13g2_fill_1 FILLER_43_159 ();
 sg13g2_decap_8 FILLER_43_197 ();
 sg13g2_fill_2 FILLER_43_204 ();
 sg13g2_fill_2 FILLER_43_212 ();
 sg13g2_fill_1 FILLER_43_214 ();
 sg13g2_decap_4 FILLER_43_241 ();
 sg13g2_fill_2 FILLER_43_249 ();
 sg13g2_decap_4 FILLER_43_254 ();
 sg13g2_fill_2 FILLER_43_262 ();
 sg13g2_fill_1 FILLER_43_274 ();
 sg13g2_decap_4 FILLER_43_285 ();
 sg13g2_fill_1 FILLER_43_289 ();
 sg13g2_decap_8 FILLER_43_298 ();
 sg13g2_fill_2 FILLER_43_305 ();
 sg13g2_fill_1 FILLER_43_307 ();
 sg13g2_decap_8 FILLER_43_331 ();
 sg13g2_decap_4 FILLER_43_338 ();
 sg13g2_fill_2 FILLER_43_342 ();
 sg13g2_decap_4 FILLER_43_348 ();
 sg13g2_decap_8 FILLER_43_358 ();
 sg13g2_fill_2 FILLER_43_365 ();
 sg13g2_fill_1 FILLER_43_367 ();
 sg13g2_decap_8 FILLER_43_373 ();
 sg13g2_fill_1 FILLER_43_380 ();
 sg13g2_decap_4 FILLER_43_425 ();
 sg13g2_fill_1 FILLER_43_429 ();
 sg13g2_fill_1 FILLER_44_0 ();
 sg13g2_fill_1 FILLER_44_27 ();
 sg13g2_fill_1 FILLER_44_33 ();
 sg13g2_fill_1 FILLER_44_38 ();
 sg13g2_fill_1 FILLER_44_54 ();
 sg13g2_fill_1 FILLER_44_77 ();
 sg13g2_decap_4 FILLER_44_91 ();
 sg13g2_decap_8 FILLER_44_102 ();
 sg13g2_decap_8 FILLER_44_109 ();
 sg13g2_decap_8 FILLER_44_116 ();
 sg13g2_decap_8 FILLER_44_123 ();
 sg13g2_decap_8 FILLER_44_130 ();
 sg13g2_fill_2 FILLER_44_137 ();
 sg13g2_decap_8 FILLER_44_143 ();
 sg13g2_fill_1 FILLER_44_155 ();
 sg13g2_fill_1 FILLER_44_160 ();
 sg13g2_fill_2 FILLER_44_167 ();
 sg13g2_fill_1 FILLER_44_184 ();
 sg13g2_fill_1 FILLER_44_211 ();
 sg13g2_fill_1 FILLER_44_216 ();
 sg13g2_fill_1 FILLER_44_243 ();
 sg13g2_fill_2 FILLER_44_250 ();
 sg13g2_fill_1 FILLER_44_258 ();
 sg13g2_decap_8 FILLER_44_267 ();
 sg13g2_decap_8 FILLER_44_274 ();
 sg13g2_decap_8 FILLER_44_281 ();
 sg13g2_fill_1 FILLER_44_288 ();
 sg13g2_fill_1 FILLER_44_320 ();
 sg13g2_decap_4 FILLER_44_326 ();
 sg13g2_fill_2 FILLER_44_339 ();
 sg13g2_fill_2 FILLER_44_379 ();
 sg13g2_fill_1 FILLER_44_381 ();
 sg13g2_fill_1 FILLER_44_386 ();
 sg13g2_fill_2 FILLER_44_417 ();
 sg13g2_decap_8 FILLER_44_423 ();
 sg13g2_decap_8 FILLER_45_0 ();
 sg13g2_decap_8 FILLER_45_11 ();
 sg13g2_decap_8 FILLER_45_18 ();
 sg13g2_decap_8 FILLER_45_25 ();
 sg13g2_decap_4 FILLER_45_32 ();
 sg13g2_fill_1 FILLER_45_36 ();
 sg13g2_decap_4 FILLER_45_71 ();
 sg13g2_fill_1 FILLER_45_75 ();
 sg13g2_decap_8 FILLER_45_85 ();
 sg13g2_fill_2 FILLER_45_92 ();
 sg13g2_fill_1 FILLER_45_94 ();
 sg13g2_fill_1 FILLER_45_126 ();
 sg13g2_fill_1 FILLER_45_132 ();
 sg13g2_fill_1 FILLER_45_159 ();
 sg13g2_fill_1 FILLER_45_165 ();
 sg13g2_fill_1 FILLER_45_171 ();
 sg13g2_fill_1 FILLER_45_177 ();
 sg13g2_fill_1 FILLER_45_183 ();
 sg13g2_fill_2 FILLER_45_203 ();
 sg13g2_fill_1 FILLER_45_221 ();
 sg13g2_fill_1 FILLER_45_227 ();
 sg13g2_fill_1 FILLER_45_232 ();
 sg13g2_fill_1 FILLER_45_238 ();
 sg13g2_fill_2 FILLER_45_244 ();
 sg13g2_decap_4 FILLER_45_250 ();
 sg13g2_decap_4 FILLER_45_265 ();
 sg13g2_fill_2 FILLER_45_269 ();
 sg13g2_decap_4 FILLER_45_324 ();
 sg13g2_fill_2 FILLER_45_328 ();
 sg13g2_fill_2 FILLER_45_396 ();
 sg13g2_fill_2 FILLER_45_402 ();
 sg13g2_fill_1 FILLER_46_0 ();
 sg13g2_fill_2 FILLER_46_27 ();
 sg13g2_fill_1 FILLER_46_29 ();
 sg13g2_decap_8 FILLER_46_79 ();
 sg13g2_decap_8 FILLER_46_86 ();
 sg13g2_decap_8 FILLER_46_93 ();
 sg13g2_fill_1 FILLER_46_100 ();
 sg13g2_decap_4 FILLER_46_105 ();
 sg13g2_fill_2 FILLER_46_135 ();
 sg13g2_decap_4 FILLER_46_145 ();
 sg13g2_fill_1 FILLER_46_149 ();
 sg13g2_fill_1 FILLER_46_158 ();
 sg13g2_fill_1 FILLER_46_180 ();
 sg13g2_decap_8 FILLER_46_186 ();
 sg13g2_decap_8 FILLER_46_193 ();
 sg13g2_fill_1 FILLER_46_200 ();
 sg13g2_fill_2 FILLER_46_215 ();
 sg13g2_fill_1 FILLER_46_221 ();
 sg13g2_fill_2 FILLER_46_226 ();
 sg13g2_fill_2 FILLER_46_231 ();
 sg13g2_fill_1 FILLER_46_237 ();
 sg13g2_fill_1 FILLER_46_278 ();
 sg13g2_decap_4 FILLER_46_287 ();
 sg13g2_decap_4 FILLER_46_302 ();
 sg13g2_fill_1 FILLER_46_317 ();
 sg13g2_decap_8 FILLER_46_324 ();
 sg13g2_fill_1 FILLER_46_331 ();
 sg13g2_decap_4 FILLER_46_359 ();
 sg13g2_fill_1 FILLER_46_363 ();
 sg13g2_fill_1 FILLER_46_378 ();
 sg13g2_fill_1 FILLER_46_389 ();
 sg13g2_decap_4 FILLER_46_424 ();
 sg13g2_fill_2 FILLER_46_428 ();
 sg13g2_decap_4 FILLER_47_43 ();
 sg13g2_decap_8 FILLER_47_60 ();
 sg13g2_decap_8 FILLER_47_67 ();
 sg13g2_decap_8 FILLER_47_74 ();
 sg13g2_decap_8 FILLER_47_81 ();
 sg13g2_decap_8 FILLER_47_88 ();
 sg13g2_decap_8 FILLER_47_95 ();
 sg13g2_decap_8 FILLER_47_102 ();
 sg13g2_decap_8 FILLER_47_109 ();
 sg13g2_fill_1 FILLER_47_116 ();
 sg13g2_decap_8 FILLER_47_121 ();
 sg13g2_decap_4 FILLER_47_128 ();
 sg13g2_fill_2 FILLER_47_132 ();
 sg13g2_decap_8 FILLER_47_144 ();
 sg13g2_fill_1 FILLER_47_151 ();
 sg13g2_fill_1 FILLER_47_171 ();
 sg13g2_decap_8 FILLER_47_182 ();
 sg13g2_decap_8 FILLER_47_189 ();
 sg13g2_fill_2 FILLER_47_214 ();
 sg13g2_fill_1 FILLER_47_220 ();
 sg13g2_fill_1 FILLER_47_242 ();
 sg13g2_decap_4 FILLER_47_265 ();
 sg13g2_fill_1 FILLER_47_273 ();
 sg13g2_decap_8 FILLER_47_284 ();
 sg13g2_decap_8 FILLER_47_291 ();
 sg13g2_fill_1 FILLER_47_298 ();
 sg13g2_fill_2 FILLER_47_304 ();
 sg13g2_decap_8 FILLER_47_325 ();
 sg13g2_fill_2 FILLER_47_340 ();
 sg13g2_fill_2 FILLER_47_352 ();
 sg13g2_fill_1 FILLER_47_354 ();
 sg13g2_decap_8 FILLER_47_389 ();
 sg13g2_decap_8 FILLER_47_396 ();
 sg13g2_fill_1 FILLER_47_403 ();
 sg13g2_decap_4 FILLER_47_408 ();
 sg13g2_fill_1 FILLER_47_412 ();
 sg13g2_fill_2 FILLER_47_417 ();
 sg13g2_decap_8 FILLER_47_423 ();
 sg13g2_decap_8 FILLER_48_0 ();
 sg13g2_fill_2 FILLER_48_7 ();
 sg13g2_fill_1 FILLER_48_9 ();
 sg13g2_decap_4 FILLER_48_14 ();
 sg13g2_fill_2 FILLER_48_18 ();
 sg13g2_fill_2 FILLER_48_25 ();
 sg13g2_fill_1 FILLER_48_27 ();
 sg13g2_decap_8 FILLER_48_36 ();
 sg13g2_decap_8 FILLER_48_43 ();
 sg13g2_decap_8 FILLER_48_50 ();
 sg13g2_decap_8 FILLER_48_57 ();
 sg13g2_decap_8 FILLER_48_64 ();
 sg13g2_decap_8 FILLER_48_71 ();
 sg13g2_decap_8 FILLER_48_78 ();
 sg13g2_decap_4 FILLER_48_85 ();
 sg13g2_decap_4 FILLER_48_115 ();
 sg13g2_fill_2 FILLER_48_119 ();
 sg13g2_decap_4 FILLER_48_129 ();
 sg13g2_decap_8 FILLER_48_137 ();
 sg13g2_decap_8 FILLER_48_144 ();
 sg13g2_fill_1 FILLER_48_181 ();
 sg13g2_decap_4 FILLER_48_191 ();
 sg13g2_fill_2 FILLER_48_195 ();
 sg13g2_decap_8 FILLER_48_201 ();
 sg13g2_decap_4 FILLER_48_208 ();
 sg13g2_fill_1 FILLER_48_234 ();
 sg13g2_decap_4 FILLER_48_277 ();
 sg13g2_fill_2 FILLER_48_281 ();
 sg13g2_decap_8 FILLER_48_295 ();
 sg13g2_decap_4 FILLER_48_302 ();
 sg13g2_fill_2 FILLER_48_306 ();
 sg13g2_decap_8 FILLER_48_325 ();
 sg13g2_fill_1 FILLER_48_332 ();
 sg13g2_fill_1 FILLER_48_337 ();
 sg13g2_fill_1 FILLER_48_364 ();
 sg13g2_fill_1 FILLER_48_369 ();
 sg13g2_fill_1 FILLER_48_376 ();
 sg13g2_fill_2 FILLER_48_381 ();
 sg13g2_fill_1 FILLER_48_395 ();
 sg13g2_decap_4 FILLER_48_426 ();
 sg13g2_decap_8 FILLER_49_0 ();
 sg13g2_decap_8 FILLER_49_7 ();
 sg13g2_decap_8 FILLER_49_14 ();
 sg13g2_decap_8 FILLER_49_21 ();
 sg13g2_decap_8 FILLER_49_28 ();
 sg13g2_decap_8 FILLER_49_35 ();
 sg13g2_decap_8 FILLER_49_42 ();
 sg13g2_decap_8 FILLER_49_49 ();
 sg13g2_decap_8 FILLER_49_56 ();
 sg13g2_fill_2 FILLER_49_63 ();
 sg13g2_fill_1 FILLER_49_73 ();
 sg13g2_fill_1 FILLER_49_100 ();
 sg13g2_fill_1 FILLER_49_114 ();
 sg13g2_fill_1 FILLER_49_125 ();
 sg13g2_decap_8 FILLER_49_152 ();
 sg13g2_fill_1 FILLER_49_163 ();
 sg13g2_decap_4 FILLER_49_168 ();
 sg13g2_fill_2 FILLER_49_185 ();
 sg13g2_fill_1 FILLER_49_187 ();
 sg13g2_decap_8 FILLER_49_214 ();
 sg13g2_decap_4 FILLER_49_221 ();
 sg13g2_fill_1 FILLER_49_225 ();
 sg13g2_fill_2 FILLER_49_236 ();
 sg13g2_fill_2 FILLER_49_242 ();
 sg13g2_fill_1 FILLER_49_259 ();
 sg13g2_fill_2 FILLER_49_286 ();
 sg13g2_fill_1 FILLER_49_288 ();
 sg13g2_fill_1 FILLER_49_292 ();
 sg13g2_decap_8 FILLER_49_297 ();
 sg13g2_fill_2 FILLER_49_304 ();
 sg13g2_fill_2 FILLER_49_318 ();
 sg13g2_fill_1 FILLER_49_323 ();
 sg13g2_fill_1 FILLER_49_350 ();
 sg13g2_fill_1 FILLER_49_356 ();
 sg13g2_fill_2 FILLER_49_362 ();
 sg13g2_fill_1 FILLER_49_364 ();
 sg13g2_fill_2 FILLER_49_369 ();
 sg13g2_fill_1 FILLER_49_371 ();
 sg13g2_decap_4 FILLER_49_377 ();
 sg13g2_fill_1 FILLER_49_381 ();
 sg13g2_fill_2 FILLER_49_387 ();
 sg13g2_fill_1 FILLER_49_394 ();
 sg13g2_fill_2 FILLER_49_407 ();
 sg13g2_fill_1 FILLER_49_425 ();
 sg13g2_decap_8 FILLER_50_0 ();
 sg13g2_decap_8 FILLER_50_7 ();
 sg13g2_decap_8 FILLER_50_14 ();
 sg13g2_decap_8 FILLER_50_21 ();
 sg13g2_fill_2 FILLER_50_28 ();
 sg13g2_fill_1 FILLER_50_70 ();
 sg13g2_fill_1 FILLER_50_84 ();
 sg13g2_fill_2 FILLER_50_102 ();
 sg13g2_fill_2 FILLER_50_116 ();
 sg13g2_fill_2 FILLER_50_122 ();
 sg13g2_fill_1 FILLER_50_124 ();
 sg13g2_decap_4 FILLER_50_151 ();
 sg13g2_fill_2 FILLER_50_181 ();
 sg13g2_fill_1 FILLER_50_183 ();
 sg13g2_fill_2 FILLER_50_225 ();
 sg13g2_fill_1 FILLER_50_240 ();
 sg13g2_fill_1 FILLER_50_246 ();
 sg13g2_fill_1 FILLER_50_298 ();
 sg13g2_fill_2 FILLER_50_304 ();
 sg13g2_decap_4 FILLER_50_324 ();
 sg13g2_decap_8 FILLER_50_336 ();
 sg13g2_fill_2 FILLER_50_343 ();
 sg13g2_fill_2 FILLER_50_383 ();
 sg13g2_fill_1 FILLER_50_420 ();
 sg13g2_decap_4 FILLER_50_426 ();
 sg13g2_fill_1 FILLER_51_63 ();
 sg13g2_fill_1 FILLER_51_88 ();
 sg13g2_fill_1 FILLER_51_102 ();
 sg13g2_fill_2 FILLER_51_112 ();
 sg13g2_fill_1 FILLER_51_114 ();
 sg13g2_fill_1 FILLER_51_120 ();
 sg13g2_fill_2 FILLER_51_155 ();
 sg13g2_fill_1 FILLER_51_157 ();
 sg13g2_fill_2 FILLER_51_184 ();
 sg13g2_fill_1 FILLER_51_186 ();
 sg13g2_fill_1 FILLER_51_197 ();
 sg13g2_fill_2 FILLER_51_202 ();
 sg13g2_fill_1 FILLER_51_209 ();
 sg13g2_fill_2 FILLER_51_215 ();
 sg13g2_fill_2 FILLER_51_222 ();
 sg13g2_fill_2 FILLER_51_228 ();
 sg13g2_fill_2 FILLER_51_235 ();
 sg13g2_fill_1 FILLER_51_237 ();
 sg13g2_fill_1 FILLER_51_296 ();
 sg13g2_decap_8 FILLER_51_327 ();
 sg13g2_decap_8 FILLER_51_334 ();
 sg13g2_decap_4 FILLER_51_341 ();
 sg13g2_decap_8 FILLER_51_349 ();
 sg13g2_decap_8 FILLER_51_356 ();
 sg13g2_decap_4 FILLER_51_363 ();
 sg13g2_fill_1 FILLER_51_367 ();
 sg13g2_fill_2 FILLER_51_396 ();
 sg13g2_fill_1 FILLER_51_402 ();
 sg13g2_fill_2 FILLER_51_420 ();
 sg13g2_fill_2 FILLER_51_427 ();
 sg13g2_fill_1 FILLER_51_429 ();
 sg13g2_decap_4 FILLER_52_31 ();
 sg13g2_fill_2 FILLER_52_39 ();
 sg13g2_fill_2 FILLER_52_45 ();
 sg13g2_fill_1 FILLER_52_47 ();
 sg13g2_fill_2 FILLER_52_73 ();
 sg13g2_fill_1 FILLER_52_126 ();
 sg13g2_fill_2 FILLER_52_132 ();
 sg13g2_decap_8 FILLER_52_142 ();
 sg13g2_fill_1 FILLER_52_149 ();
 sg13g2_fill_2 FILLER_52_155 ();
 sg13g2_fill_1 FILLER_52_157 ();
 sg13g2_fill_2 FILLER_52_162 ();
 sg13g2_fill_1 FILLER_52_164 ();
 sg13g2_decap_8 FILLER_52_174 ();
 sg13g2_fill_1 FILLER_52_181 ();
 sg13g2_fill_2 FILLER_52_200 ();
 sg13g2_fill_1 FILLER_52_216 ();
 sg13g2_fill_1 FILLER_52_222 ();
 sg13g2_decap_8 FILLER_52_233 ();
 sg13g2_decap_8 FILLER_52_240 ();
 sg13g2_fill_1 FILLER_52_247 ();
 sg13g2_decap_4 FILLER_52_269 ();
 sg13g2_decap_8 FILLER_52_282 ();
 sg13g2_decap_8 FILLER_52_289 ();
 sg13g2_fill_2 FILLER_52_301 ();
 sg13g2_decap_8 FILLER_52_307 ();
 sg13g2_decap_8 FILLER_52_314 ();
 sg13g2_fill_1 FILLER_52_347 ();
 sg13g2_fill_2 FILLER_52_354 ();
 sg13g2_fill_2 FILLER_52_361 ();
 sg13g2_fill_2 FILLER_52_373 ();
 sg13g2_fill_1 FILLER_52_383 ();
 sg13g2_fill_2 FILLER_52_392 ();
 sg13g2_decap_8 FILLER_52_399 ();
 sg13g2_fill_2 FILLER_52_406 ();
 sg13g2_fill_1 FILLER_52_408 ();
 sg13g2_fill_2 FILLER_52_428 ();
 sg13g2_fill_1 FILLER_53_0 ();
 sg13g2_fill_2 FILLER_53_5 ();
 sg13g2_fill_1 FILLER_53_11 ();
 sg13g2_fill_2 FILLER_53_17 ();
 sg13g2_fill_2 FILLER_53_24 ();
 sg13g2_fill_2 FILLER_53_74 ();
 sg13g2_fill_2 FILLER_53_85 ();
 sg13g2_fill_1 FILLER_53_87 ();
 sg13g2_fill_2 FILLER_53_100 ();
 sg13g2_fill_1 FILLER_53_107 ();
 sg13g2_fill_2 FILLER_53_112 ();
 sg13g2_decap_4 FILLER_53_140 ();
 sg13g2_fill_2 FILLER_53_144 ();
 sg13g2_fill_2 FILLER_53_161 ();
 sg13g2_decap_4 FILLER_53_166 ();
 sg13g2_fill_2 FILLER_53_180 ();
 sg13g2_decap_8 FILLER_53_187 ();
 sg13g2_fill_1 FILLER_53_194 ();
 sg13g2_fill_2 FILLER_53_199 ();
 sg13g2_fill_2 FILLER_53_220 ();
 sg13g2_decap_4 FILLER_53_238 ();
 sg13g2_fill_2 FILLER_53_242 ();
 sg13g2_fill_1 FILLER_53_269 ();
 sg13g2_fill_2 FILLER_53_279 ();
 sg13g2_fill_1 FILLER_53_281 ();
 sg13g2_decap_8 FILLER_53_290 ();
 sg13g2_fill_2 FILLER_53_297 ();
 sg13g2_fill_1 FILLER_53_299 ();
 sg13g2_decap_8 FILLER_53_308 ();
 sg13g2_fill_1 FILLER_53_350 ();
 sg13g2_fill_1 FILLER_53_371 ();
 sg13g2_fill_1 FILLER_53_376 ();
 sg13g2_fill_2 FILLER_53_397 ();
 sg13g2_decap_8 FILLER_53_403 ();
 sg13g2_decap_4 FILLER_53_410 ();
 sg13g2_fill_2 FILLER_53_419 ();
 sg13g2_fill_1 FILLER_53_421 ();
 sg13g2_decap_4 FILLER_53_426 ();
 sg13g2_decap_4 FILLER_54_31 ();
 sg13g2_fill_1 FILLER_54_35 ();
 sg13g2_fill_2 FILLER_54_40 ();
 sg13g2_fill_1 FILLER_54_42 ();
 sg13g2_fill_1 FILLER_54_47 ();
 sg13g2_fill_2 FILLER_54_72 ();
 sg13g2_fill_1 FILLER_54_74 ();
 sg13g2_decap_8 FILLER_54_90 ();
 sg13g2_fill_1 FILLER_54_97 ();
 sg13g2_decap_8 FILLER_54_113 ();
 sg13g2_decap_8 FILLER_54_120 ();
 sg13g2_decap_4 FILLER_54_127 ();
 sg13g2_fill_2 FILLER_54_161 ();
 sg13g2_decap_4 FILLER_54_175 ();
 sg13g2_fill_1 FILLER_54_179 ();
 sg13g2_decap_8 FILLER_54_185 ();
 sg13g2_fill_1 FILLER_54_192 ();
 sg13g2_fill_2 FILLER_54_214 ();
 sg13g2_fill_1 FILLER_54_222 ();
 sg13g2_fill_1 FILLER_54_233 ();
 sg13g2_fill_2 FILLER_54_248 ();
 sg13g2_fill_1 FILLER_54_250 ();
 sg13g2_decap_8 FILLER_54_262 ();
 sg13g2_fill_2 FILLER_54_269 ();
 sg13g2_decap_4 FILLER_54_306 ();
 sg13g2_fill_1 FILLER_54_315 ();
 sg13g2_fill_2 FILLER_54_328 ();
 sg13g2_fill_2 FILLER_54_334 ();
 sg13g2_decap_8 FILLER_54_346 ();
 sg13g2_fill_2 FILLER_54_353 ();
 sg13g2_fill_2 FILLER_54_384 ();
 sg13g2_fill_2 FILLER_54_396 ();
 sg13g2_fill_1 FILLER_54_403 ();
 sg13g2_fill_1 FILLER_55_0 ();
 sg13g2_fill_2 FILLER_55_14 ();
 sg13g2_fill_1 FILLER_55_21 ();
 sg13g2_fill_2 FILLER_55_48 ();
 sg13g2_fill_2 FILLER_55_54 ();
 sg13g2_fill_1 FILLER_55_56 ();
 sg13g2_fill_2 FILLER_55_61 ();
 sg13g2_fill_1 FILLER_55_63 ();
 sg13g2_fill_2 FILLER_55_68 ();
 sg13g2_decap_8 FILLER_55_79 ();
 sg13g2_fill_2 FILLER_55_86 ();
 sg13g2_fill_1 FILLER_55_88 ();
 sg13g2_decap_8 FILLER_55_93 ();
 sg13g2_decap_4 FILLER_55_103 ();
 sg13g2_fill_1 FILLER_55_107 ();
 sg13g2_decap_8 FILLER_55_117 ();
 sg13g2_fill_2 FILLER_55_124 ();
 sg13g2_decap_4 FILLER_55_161 ();
 sg13g2_fill_1 FILLER_55_165 ();
 sg13g2_fill_1 FILLER_55_185 ();
 sg13g2_fill_1 FILLER_55_190 ();
 sg13g2_decap_8 FILLER_55_205 ();
 sg13g2_fill_1 FILLER_55_212 ();
 sg13g2_decap_8 FILLER_55_217 ();
 sg13g2_decap_4 FILLER_55_228 ();
 sg13g2_fill_2 FILLER_55_245 ();
 sg13g2_fill_1 FILLER_55_247 ();
 sg13g2_fill_1 FILLER_55_279 ();
 sg13g2_decap_8 FILLER_55_310 ();
 sg13g2_decap_8 FILLER_55_317 ();
 sg13g2_decap_8 FILLER_55_324 ();
 sg13g2_decap_8 FILLER_55_331 ();
 sg13g2_decap_8 FILLER_55_338 ();
 sg13g2_decap_8 FILLER_55_345 ();
 sg13g2_fill_2 FILLER_55_352 ();
 sg13g2_decap_8 FILLER_55_358 ();
 sg13g2_decap_4 FILLER_55_365 ();
 sg13g2_decap_4 FILLER_55_386 ();
 sg13g2_decap_4 FILLER_55_425 ();
 sg13g2_fill_1 FILLER_55_429 ();
 sg13g2_fill_1 FILLER_56_26 ();
 sg13g2_decap_4 FILLER_56_31 ();
 sg13g2_decap_8 FILLER_56_39 ();
 sg13g2_decap_4 FILLER_56_46 ();
 sg13g2_fill_1 FILLER_56_50 ();
 sg13g2_fill_1 FILLER_56_56 ();
 sg13g2_fill_1 FILLER_56_62 ();
 sg13g2_fill_1 FILLER_56_66 ();
 sg13g2_fill_1 FILLER_56_75 ();
 sg13g2_fill_1 FILLER_56_104 ();
 sg13g2_decap_4 FILLER_56_110 ();
 sg13g2_fill_2 FILLER_56_131 ();
 sg13g2_fill_1 FILLER_56_133 ();
 sg13g2_decap_8 FILLER_56_142 ();
 sg13g2_decap_8 FILLER_56_149 ();
 sg13g2_fill_1 FILLER_56_156 ();
 sg13g2_fill_2 FILLER_56_164 ();
 sg13g2_fill_1 FILLER_56_166 ();
 sg13g2_fill_1 FILLER_56_172 ();
 sg13g2_fill_1 FILLER_56_183 ();
 sg13g2_fill_2 FILLER_56_199 ();
 sg13g2_fill_2 FILLER_56_215 ();
 sg13g2_decap_4 FILLER_56_227 ();
 sg13g2_fill_2 FILLER_56_231 ();
 sg13g2_fill_1 FILLER_56_254 ();
 sg13g2_fill_1 FILLER_56_267 ();
 sg13g2_fill_1 FILLER_56_286 ();
 sg13g2_fill_2 FILLER_56_291 ();
 sg13g2_fill_2 FILLER_56_324 ();
 sg13g2_decap_8 FILLER_56_331 ();
 sg13g2_decap_8 FILLER_56_338 ();
 sg13g2_fill_1 FILLER_56_345 ();
 sg13g2_decap_4 FILLER_56_397 ();
 sg13g2_decap_8 FILLER_56_405 ();
 sg13g2_decap_8 FILLER_56_412 ();
 sg13g2_decap_8 FILLER_56_419 ();
 sg13g2_decap_4 FILLER_56_426 ();
 sg13g2_fill_2 FILLER_57_0 ();
 sg13g2_fill_1 FILLER_57_2 ();
 sg13g2_decap_8 FILLER_57_7 ();
 sg13g2_decap_4 FILLER_57_14 ();
 sg13g2_fill_1 FILLER_57_18 ();
 sg13g2_decap_4 FILLER_57_24 ();
 sg13g2_fill_1 FILLER_57_54 ();
 sg13g2_fill_1 FILLER_57_60 ();
 sg13g2_fill_1 FILLER_57_69 ();
 sg13g2_fill_1 FILLER_57_75 ();
 sg13g2_decap_4 FILLER_57_112 ();
 sg13g2_decap_8 FILLER_57_120 ();
 sg13g2_decap_4 FILLER_57_127 ();
 sg13g2_fill_2 FILLER_57_131 ();
 sg13g2_fill_1 FILLER_57_137 ();
 sg13g2_fill_2 FILLER_57_173 ();
 sg13g2_fill_1 FILLER_57_175 ();
 sg13g2_fill_2 FILLER_57_193 ();
 sg13g2_decap_8 FILLER_57_200 ();
 sg13g2_fill_1 FILLER_57_212 ();
 sg13g2_fill_1 FILLER_57_220 ();
 sg13g2_decap_8 FILLER_57_226 ();
 sg13g2_fill_2 FILLER_57_233 ();
 sg13g2_fill_2 FILLER_57_240 ();
 sg13g2_fill_1 FILLER_57_242 ();
 sg13g2_fill_2 FILLER_57_261 ();
 sg13g2_decap_4 FILLER_57_268 ();
 sg13g2_fill_1 FILLER_57_272 ();
 sg13g2_decap_4 FILLER_57_278 ();
 sg13g2_fill_1 FILLER_57_282 ();
 sg13g2_fill_2 FILLER_57_317 ();
 sg13g2_fill_1 FILLER_57_350 ();
 sg13g2_fill_1 FILLER_57_396 ();
 sg13g2_decap_4 FILLER_57_406 ();
 sg13g2_fill_1 FILLER_57_410 ();
 sg13g2_decap_4 FILLER_57_415 ();
 sg13g2_decap_8 FILLER_57_423 ();
 sg13g2_fill_1 FILLER_58_26 ();
 sg13g2_fill_2 FILLER_58_35 ();
 sg13g2_fill_1 FILLER_58_37 ();
 sg13g2_decap_8 FILLER_58_73 ();
 sg13g2_fill_2 FILLER_58_100 ();
 sg13g2_decap_8 FILLER_58_128 ();
 sg13g2_decap_8 FILLER_58_135 ();
 sg13g2_fill_2 FILLER_58_142 ();
 sg13g2_fill_2 FILLER_58_148 ();
 sg13g2_decap_4 FILLER_58_154 ();
 sg13g2_fill_2 FILLER_58_158 ();
 sg13g2_decap_4 FILLER_58_166 ();
 sg13g2_fill_2 FILLER_58_174 ();
 sg13g2_fill_2 FILLER_58_185 ();
 sg13g2_decap_4 FILLER_58_196 ();
 sg13g2_fill_1 FILLER_58_200 ();
 sg13g2_fill_2 FILLER_58_234 ();
 sg13g2_fill_2 FILLER_58_256 ();
 sg13g2_decap_8 FILLER_58_284 ();
 sg13g2_fill_2 FILLER_58_291 ();
 sg13g2_fill_1 FILLER_58_293 ();
 sg13g2_fill_2 FILLER_58_298 ();
 sg13g2_fill_1 FILLER_58_305 ();
 sg13g2_fill_2 FILLER_58_315 ();
 sg13g2_fill_1 FILLER_58_322 ();
 sg13g2_fill_2 FILLER_58_327 ();
 sg13g2_fill_1 FILLER_58_333 ();
 sg13g2_fill_1 FILLER_58_388 ();
 sg13g2_fill_2 FILLER_58_392 ();
 sg13g2_fill_2 FILLER_59_0 ();
 sg13g2_fill_1 FILLER_59_2 ();
 sg13g2_decap_4 FILLER_59_33 ();
 sg13g2_fill_1 FILLER_59_37 ();
 sg13g2_fill_1 FILLER_59_58 ();
 sg13g2_decap_8 FILLER_59_113 ();
 sg13g2_decap_8 FILLER_59_120 ();
 sg13g2_decap_4 FILLER_59_127 ();
 sg13g2_fill_1 FILLER_59_131 ();
 sg13g2_fill_1 FILLER_59_137 ();
 sg13g2_fill_1 FILLER_59_147 ();
 sg13g2_fill_1 FILLER_59_152 ();
 sg13g2_fill_1 FILLER_59_158 ();
 sg13g2_fill_1 FILLER_59_167 ();
 sg13g2_fill_1 FILLER_59_173 ();
 sg13g2_fill_2 FILLER_59_179 ();
 sg13g2_decap_8 FILLER_59_191 ();
 sg13g2_decap_4 FILLER_59_198 ();
 sg13g2_fill_1 FILLER_59_202 ();
 sg13g2_fill_2 FILLER_59_208 ();
 sg13g2_fill_1 FILLER_59_218 ();
 sg13g2_fill_1 FILLER_59_233 ();
 sg13g2_fill_2 FILLER_59_240 ();
 sg13g2_decap_8 FILLER_59_248 ();
 sg13g2_decap_4 FILLER_59_286 ();
 sg13g2_fill_2 FILLER_59_308 ();
 sg13g2_decap_8 FILLER_59_326 ();
 sg13g2_fill_2 FILLER_59_354 ();
 sg13g2_fill_2 FILLER_59_361 ();
 sg13g2_fill_1 FILLER_59_363 ();
 sg13g2_fill_2 FILLER_59_368 ();
 sg13g2_decap_8 FILLER_59_380 ();
 sg13g2_decap_4 FILLER_59_387 ();
 sg13g2_fill_2 FILLER_59_391 ();
 sg13g2_fill_2 FILLER_59_397 ();
 sg13g2_decap_8 FILLER_60_0 ();
 sg13g2_decap_4 FILLER_60_7 ();
 sg13g2_fill_1 FILLER_60_20 ();
 sg13g2_fill_2 FILLER_60_47 ();
 sg13g2_fill_1 FILLER_60_49 ();
 sg13g2_fill_2 FILLER_60_80 ();
 sg13g2_fill_2 FILLER_60_108 ();
 sg13g2_fill_2 FILLER_60_136 ();
 sg13g2_fill_1 FILLER_60_138 ();
 sg13g2_fill_1 FILLER_60_165 ();
 sg13g2_fill_2 FILLER_60_170 ();
 sg13g2_fill_1 FILLER_60_172 ();
 sg13g2_fill_1 FILLER_60_178 ();
 sg13g2_fill_1 FILLER_60_182 ();
 sg13g2_decap_8 FILLER_60_193 ();
 sg13g2_decap_8 FILLER_60_200 ();
 sg13g2_fill_2 FILLER_60_212 ();
 sg13g2_fill_1 FILLER_60_214 ();
 sg13g2_decap_8 FILLER_60_224 ();
 sg13g2_decap_4 FILLER_60_231 ();
 sg13g2_fill_1 FILLER_60_235 ();
 sg13g2_decap_8 FILLER_60_251 ();
 sg13g2_decap_4 FILLER_60_258 ();
 sg13g2_fill_2 FILLER_60_270 ();
 sg13g2_fill_2 FILLER_60_298 ();
 sg13g2_fill_2 FILLER_60_305 ();
 sg13g2_fill_1 FILLER_60_307 ();
 sg13g2_decap_4 FILLER_60_338 ();
 sg13g2_fill_1 FILLER_60_350 ();
 sg13g2_fill_1 FILLER_60_356 ();
 sg13g2_fill_2 FILLER_60_369 ();
 sg13g2_fill_1 FILLER_60_371 ();
 sg13g2_decap_8 FILLER_60_416 ();
 sg13g2_decap_8 FILLER_60_423 ();
 sg13g2_decap_8 FILLER_61_0 ();
 sg13g2_fill_2 FILLER_61_7 ();
 sg13g2_fill_1 FILLER_61_9 ();
 sg13g2_decap_8 FILLER_61_22 ();
 sg13g2_decap_8 FILLER_61_29 ();
 sg13g2_decap_8 FILLER_61_36 ();
 sg13g2_fill_1 FILLER_61_43 ();
 sg13g2_fill_2 FILLER_61_48 ();
 sg13g2_fill_1 FILLER_61_50 ();
 sg13g2_decap_8 FILLER_61_77 ();
 sg13g2_decap_4 FILLER_61_84 ();
 sg13g2_fill_2 FILLER_61_88 ();
 sg13g2_decap_8 FILLER_61_94 ();
 sg13g2_decap_8 FILLER_61_101 ();
 sg13g2_decap_8 FILLER_61_108 ();
 sg13g2_fill_2 FILLER_61_115 ();
 sg13g2_fill_2 FILLER_61_121 ();
 sg13g2_fill_1 FILLER_61_123 ();
 sg13g2_fill_2 FILLER_61_134 ();
 sg13g2_decap_8 FILLER_61_140 ();
 sg13g2_fill_1 FILLER_61_147 ();
 sg13g2_fill_1 FILLER_61_155 ();
 sg13g2_fill_2 FILLER_61_169 ();
 sg13g2_fill_1 FILLER_61_171 ();
 sg13g2_fill_2 FILLER_61_177 ();
 sg13g2_fill_1 FILLER_61_179 ();
 sg13g2_fill_2 FILLER_61_198 ();
 sg13g2_fill_1 FILLER_61_200 ();
 sg13g2_fill_1 FILLER_61_209 ();
 sg13g2_fill_2 FILLER_61_225 ();
 sg13g2_fill_1 FILLER_61_227 ();
 sg13g2_fill_1 FILLER_61_237 ();
 sg13g2_fill_2 FILLER_61_249 ();
 sg13g2_decap_8 FILLER_61_259 ();
 sg13g2_decap_4 FILLER_61_266 ();
 sg13g2_fill_2 FILLER_61_274 ();
 sg13g2_decap_4 FILLER_61_310 ();
 sg13g2_fill_2 FILLER_61_314 ();
 sg13g2_decap_8 FILLER_61_325 ();
 sg13g2_decap_4 FILLER_61_341 ();
 sg13g2_fill_1 FILLER_61_359 ();
 sg13g2_fill_2 FILLER_61_365 ();
 sg13g2_fill_1 FILLER_61_367 ();
 sg13g2_decap_8 FILLER_61_373 ();
 sg13g2_fill_2 FILLER_61_380 ();
 sg13g2_fill_1 FILLER_61_386 ();
 sg13g2_decap_8 FILLER_61_391 ();
 sg13g2_fill_2 FILLER_61_398 ();
 sg13g2_fill_1 FILLER_61_400 ();
 sg13g2_decap_8 FILLER_61_411 ();
 sg13g2_decap_8 FILLER_61_418 ();
 sg13g2_decap_4 FILLER_61_425 ();
 sg13g2_fill_1 FILLER_61_429 ();
 sg13g2_fill_2 FILLER_62_26 ();
 sg13g2_fill_1 FILLER_62_28 ();
 sg13g2_decap_8 FILLER_62_33 ();
 sg13g2_decap_8 FILLER_62_40 ();
 sg13g2_decap_8 FILLER_62_47 ();
 sg13g2_decap_8 FILLER_62_62 ();
 sg13g2_decap_8 FILLER_62_69 ();
 sg13g2_decap_8 FILLER_62_76 ();
 sg13g2_decap_8 FILLER_62_83 ();
 sg13g2_decap_8 FILLER_62_90 ();
 sg13g2_decap_8 FILLER_62_97 ();
 sg13g2_fill_2 FILLER_62_120 ();
 sg13g2_fill_1 FILLER_62_131 ();
 sg13g2_decap_8 FILLER_62_140 ();
 sg13g2_decap_8 FILLER_62_147 ();
 sg13g2_fill_1 FILLER_62_154 ();
 sg13g2_fill_2 FILLER_62_172 ();
 sg13g2_fill_2 FILLER_62_190 ();
 sg13g2_decap_4 FILLER_62_198 ();
 sg13g2_fill_1 FILLER_62_217 ();
 sg13g2_fill_2 FILLER_62_222 ();
 sg13g2_fill_1 FILLER_62_224 ();
 sg13g2_fill_1 FILLER_62_245 ();
 sg13g2_decap_4 FILLER_62_262 ();
 sg13g2_decap_8 FILLER_62_274 ();
 sg13g2_decap_8 FILLER_62_281 ();
 sg13g2_fill_1 FILLER_62_288 ();
 sg13g2_fill_2 FILLER_62_293 ();
 sg13g2_decap_8 FILLER_62_304 ();
 sg13g2_decap_8 FILLER_62_311 ();
 sg13g2_fill_2 FILLER_62_318 ();
 sg13g2_fill_1 FILLER_62_324 ();
 sg13g2_decap_4 FILLER_62_365 ();
 sg13g2_fill_1 FILLER_62_369 ();
 sg13g2_fill_2 FILLER_62_401 ();
 sg13g2_fill_1 FILLER_62_403 ();
 sg13g2_decap_8 FILLER_63_0 ();
 sg13g2_fill_1 FILLER_63_7 ();
 sg13g2_decap_8 FILLER_63_12 ();
 sg13g2_fill_2 FILLER_63_19 ();
 sg13g2_fill_1 FILLER_63_21 ();
 sg13g2_decap_4 FILLER_63_27 ();
 sg13g2_fill_1 FILLER_63_31 ();
 sg13g2_decap_8 FILLER_63_36 ();
 sg13g2_decap_8 FILLER_63_43 ();
 sg13g2_fill_2 FILLER_63_50 ();
 sg13g2_fill_1 FILLER_63_52 ();
 sg13g2_decap_8 FILLER_63_58 ();
 sg13g2_decap_8 FILLER_63_65 ();
 sg13g2_fill_1 FILLER_63_72 ();
 sg13g2_fill_2 FILLER_63_77 ();
 sg13g2_decap_8 FILLER_63_83 ();
 sg13g2_decap_4 FILLER_63_90 ();
 sg13g2_fill_2 FILLER_63_94 ();
 sg13g2_decap_8 FILLER_63_141 ();
 sg13g2_decap_8 FILLER_63_148 ();
 sg13g2_decap_8 FILLER_63_155 ();
 sg13g2_decap_8 FILLER_63_162 ();
 sg13g2_fill_1 FILLER_63_213 ();
 sg13g2_fill_1 FILLER_63_249 ();
 sg13g2_fill_2 FILLER_63_256 ();
 sg13g2_decap_4 FILLER_63_288 ();
 sg13g2_fill_2 FILLER_63_292 ();
 sg13g2_decap_4 FILLER_63_298 ();
 sg13g2_fill_1 FILLER_63_302 ();
 sg13g2_decap_8 FILLER_63_307 ();
 sg13g2_fill_2 FILLER_63_344 ();
 sg13g2_fill_2 FILLER_63_351 ();
 sg13g2_fill_1 FILLER_63_353 ();
 sg13g2_fill_1 FILLER_63_380 ();
 sg13g2_fill_1 FILLER_63_385 ();
 sg13g2_fill_1 FILLER_63_396 ();
 sg13g2_fill_2 FILLER_63_402 ();
 sg13g2_decap_8 FILLER_64_0 ();
 sg13g2_decap_4 FILLER_64_16 ();
 sg13g2_decap_8 FILLER_64_51 ();
 sg13g2_decap_8 FILLER_64_58 ();
 sg13g2_fill_1 FILLER_64_92 ();
 sg13g2_fill_1 FILLER_64_107 ();
 sg13g2_fill_1 FILLER_64_120 ();
 sg13g2_fill_2 FILLER_64_155 ();
 sg13g2_fill_1 FILLER_64_161 ();
 sg13g2_fill_1 FILLER_64_167 ();
 sg13g2_fill_1 FILLER_64_173 ();
 sg13g2_fill_1 FILLER_64_186 ();
 sg13g2_fill_2 FILLER_64_200 ();
 sg13g2_fill_2 FILLER_64_249 ();
 sg13g2_fill_1 FILLER_64_255 ();
 sg13g2_fill_2 FILLER_64_282 ();
 sg13g2_fill_1 FILLER_64_284 ();
 sg13g2_fill_1 FILLER_64_307 ();
 sg13g2_fill_2 FILLER_64_334 ();
 sg13g2_fill_1 FILLER_64_362 ();
 sg13g2_fill_2 FILLER_64_367 ();
 sg13g2_decap_8 FILLER_64_423 ();
 sg13g2_fill_2 FILLER_65_26 ();
 sg13g2_fill_1 FILLER_65_28 ();
 sg13g2_fill_1 FILLER_65_89 ();
 sg13g2_fill_2 FILLER_65_99 ();
 sg13g2_fill_1 FILLER_65_125 ();
 sg13g2_fill_2 FILLER_65_130 ();
 sg13g2_fill_1 FILLER_65_140 ();
 sg13g2_fill_1 FILLER_65_145 ();
 sg13g2_fill_2 FILLER_65_205 ();
 sg13g2_fill_1 FILLER_65_217 ();
 sg13g2_fill_2 FILLER_65_259 ();
 sg13g2_fill_1 FILLER_65_261 ();
 sg13g2_decap_4 FILLER_65_266 ();
 sg13g2_fill_1 FILLER_65_270 ();
 sg13g2_decap_4 FILLER_65_275 ();
 sg13g2_fill_1 FILLER_65_310 ();
 sg13g2_fill_1 FILLER_65_319 ();
 sg13g2_decap_8 FILLER_65_328 ();
 sg13g2_decap_8 FILLER_65_335 ();
 sg13g2_decap_4 FILLER_65_346 ();
 sg13g2_fill_2 FILLER_65_350 ();
 sg13g2_decap_4 FILLER_65_356 ();
 sg13g2_fill_2 FILLER_65_360 ();
 sg13g2_decap_4 FILLER_65_372 ();
 sg13g2_fill_2 FILLER_65_376 ();
 sg13g2_decap_8 FILLER_65_382 ();
 sg13g2_decap_8 FILLER_65_389 ();
 sg13g2_decap_8 FILLER_65_396 ();
 sg13g2_decap_8 FILLER_65_403 ();
 sg13g2_decap_8 FILLER_65_410 ();
 sg13g2_fill_2 FILLER_65_417 ();
 sg13g2_decap_4 FILLER_65_424 ();
 sg13g2_fill_2 FILLER_65_428 ();
 sg13g2_fill_1 FILLER_66_71 ();
 sg13g2_fill_2 FILLER_66_98 ();
 sg13g2_fill_1 FILLER_66_100 ();
 sg13g2_fill_1 FILLER_66_106 ();
 sg13g2_fill_1 FILLER_66_112 ();
 sg13g2_fill_1 FILLER_66_118 ();
 sg13g2_fill_2 FILLER_66_130 ();
 sg13g2_fill_2 FILLER_66_137 ();
 sg13g2_fill_1 FILLER_66_139 ();
 sg13g2_decap_8 FILLER_66_145 ();
 sg13g2_fill_2 FILLER_66_156 ();
 sg13g2_fill_2 FILLER_66_162 ();
 sg13g2_fill_2 FILLER_66_168 ();
 sg13g2_fill_2 FILLER_66_175 ();
 sg13g2_fill_2 FILLER_66_182 ();
 sg13g2_fill_1 FILLER_66_189 ();
 sg13g2_decap_8 FILLER_66_195 ();
 sg13g2_decap_4 FILLER_66_202 ();
 sg13g2_decap_8 FILLER_66_215 ();
 sg13g2_decap_8 FILLER_66_222 ();
 sg13g2_decap_4 FILLER_66_234 ();
 sg13g2_fill_1 FILLER_66_238 ();
 sg13g2_fill_2 FILLER_66_243 ();
 sg13g2_fill_1 FILLER_66_245 ();
 sg13g2_decap_8 FILLER_66_254 ();
 sg13g2_fill_2 FILLER_66_261 ();
 sg13g2_fill_1 FILLER_66_263 ();
 sg13g2_fill_2 FILLER_66_273 ();
 sg13g2_fill_1 FILLER_66_275 ();
 sg13g2_decap_4 FILLER_66_306 ();
 sg13g2_fill_2 FILLER_66_323 ();
 sg13g2_fill_1 FILLER_66_325 ();
 sg13g2_fill_1 FILLER_66_341 ();
 sg13g2_fill_2 FILLER_66_346 ();
 sg13g2_fill_1 FILLER_66_353 ();
 sg13g2_fill_2 FILLER_66_359 ();
 sg13g2_fill_2 FILLER_66_370 ();
 sg13g2_decap_8 FILLER_66_376 ();
 sg13g2_decap_8 FILLER_66_383 ();
 sg13g2_decap_8 FILLER_66_390 ();
 sg13g2_fill_2 FILLER_66_397 ();
 sg13g2_fill_2 FILLER_67_39 ();
 sg13g2_fill_1 FILLER_67_41 ();
 sg13g2_fill_2 FILLER_67_50 ();
 sg13g2_fill_2 FILLER_67_57 ();
 sg13g2_fill_1 FILLER_67_59 ();
 sg13g2_fill_1 FILLER_67_64 ();
 sg13g2_decap_4 FILLER_67_92 ();
 sg13g2_fill_1 FILLER_67_96 ();
 sg13g2_decap_8 FILLER_67_101 ();
 sg13g2_fill_1 FILLER_67_108 ();
 sg13g2_fill_2 FILLER_67_113 ();
 sg13g2_decap_4 FILLER_67_120 ();
 sg13g2_fill_1 FILLER_67_127 ();
 sg13g2_decap_8 FILLER_67_140 ();
 sg13g2_decap_8 FILLER_67_147 ();
 sg13g2_fill_1 FILLER_67_154 ();
 sg13g2_decap_4 FILLER_67_164 ();
 sg13g2_decap_4 FILLER_67_173 ();
 sg13g2_decap_4 FILLER_67_181 ();
 sg13g2_fill_2 FILLER_67_194 ();
 sg13g2_fill_1 FILLER_67_196 ();
 sg13g2_decap_8 FILLER_67_201 ();
 sg13g2_fill_2 FILLER_67_208 ();
 sg13g2_fill_1 FILLER_67_210 ();
 sg13g2_decap_4 FILLER_67_215 ();
 sg13g2_decap_4 FILLER_67_223 ();
 sg13g2_decap_4 FILLER_67_253 ();
 sg13g2_fill_1 FILLER_67_287 ();
 sg13g2_fill_1 FILLER_67_292 ();
 sg13g2_decap_8 FILLER_67_301 ();
 sg13g2_decap_8 FILLER_67_308 ();
 sg13g2_decap_8 FILLER_67_315 ();
 sg13g2_decap_8 FILLER_67_322 ();
 sg13g2_fill_1 FILLER_67_329 ();
 sg13g2_fill_1 FILLER_67_356 ();
 sg13g2_fill_1 FILLER_67_396 ();
 sg13g2_decap_8 FILLER_67_402 ();
 sg13g2_fill_2 FILLER_67_409 ();
 sg13g2_fill_1 FILLER_67_415 ();
 sg13g2_fill_1 FILLER_67_424 ();
 sg13g2_fill_1 FILLER_67_429 ();
 sg13g2_decap_4 FILLER_68_0 ();
 sg13g2_fill_1 FILLER_68_4 ();
 sg13g2_decap_4 FILLER_68_14 ();
 sg13g2_fill_1 FILLER_68_57 ();
 sg13g2_fill_1 FILLER_68_71 ();
 sg13g2_fill_1 FILLER_68_76 ();
 sg13g2_fill_1 FILLER_68_82 ();
 sg13g2_fill_1 FILLER_68_87 ();
 sg13g2_decap_8 FILLER_68_159 ();
 sg13g2_decap_8 FILLER_68_166 ();
 sg13g2_decap_4 FILLER_68_208 ();
 sg13g2_fill_1 FILLER_68_212 ();
 sg13g2_fill_2 FILLER_68_309 ();
 sg13g2_fill_1 FILLER_68_311 ();
 sg13g2_fill_2 FILLER_68_325 ();
 sg13g2_fill_1 FILLER_68_331 ();
 sg13g2_decap_8 FILLER_68_358 ();
 sg13g2_decap_8 FILLER_68_391 ();
 sg13g2_fill_1 FILLER_68_398 ();
 sg13g2_fill_2 FILLER_68_407 ();
 sg13g2_fill_2 FILLER_69_31 ();
 sg13g2_fill_1 FILLER_69_33 ();
 sg13g2_decap_4 FILLER_69_60 ();
 sg13g2_decap_4 FILLER_69_68 ();
 sg13g2_fill_1 FILLER_69_82 ();
 sg13g2_fill_2 FILLER_69_106 ();
 sg13g2_fill_2 FILLER_69_121 ();
 sg13g2_fill_2 FILLER_69_149 ();
 sg13g2_fill_2 FILLER_69_156 ();
 sg13g2_decap_8 FILLER_69_188 ();
 sg13g2_decap_8 FILLER_69_195 ();
 sg13g2_decap_8 FILLER_69_202 ();
 sg13g2_decap_8 FILLER_69_209 ();
 sg13g2_decap_8 FILLER_69_216 ();
 sg13g2_decap_8 FILLER_69_250 ();
 sg13g2_decap_4 FILLER_69_257 ();
 sg13g2_fill_1 FILLER_69_261 ();
 sg13g2_fill_2 FILLER_69_306 ();
 sg13g2_fill_1 FILLER_69_346 ();
 sg13g2_fill_1 FILLER_69_351 ();
 sg13g2_fill_2 FILLER_69_367 ();
 sg13g2_fill_1 FILLER_69_369 ();
 sg13g2_decap_8 FILLER_69_374 ();
 sg13g2_decap_8 FILLER_69_381 ();
 sg13g2_decap_8 FILLER_69_392 ();
 sg13g2_fill_2 FILLER_69_399 ();
 sg13g2_fill_1 FILLER_69_401 ();
 sg13g2_fill_1 FILLER_69_429 ();
 sg13g2_decap_4 FILLER_70_0 ();
 sg13g2_decap_4 FILLER_70_12 ();
 sg13g2_fill_2 FILLER_70_16 ();
 sg13g2_decap_8 FILLER_70_23 ();
 sg13g2_decap_8 FILLER_70_30 ();
 sg13g2_decap_4 FILLER_70_37 ();
 sg13g2_decap_8 FILLER_70_45 ();
 sg13g2_fill_2 FILLER_70_52 ();
 sg13g2_decap_4 FILLER_70_59 ();
 sg13g2_fill_1 FILLER_70_63 ();
 sg13g2_fill_1 FILLER_70_69 ();
 sg13g2_fill_2 FILLER_70_75 ();
 sg13g2_fill_2 FILLER_70_117 ();
 sg13g2_fill_1 FILLER_70_129 ();
 sg13g2_fill_1 FILLER_70_166 ();
 sg13g2_fill_2 FILLER_70_171 ();
 sg13g2_decap_8 FILLER_70_184 ();
 sg13g2_decap_8 FILLER_70_191 ();
 sg13g2_fill_2 FILLER_70_198 ();
 sg13g2_decap_4 FILLER_70_230 ();
 sg13g2_decap_8 FILLER_70_238 ();
 sg13g2_decap_8 FILLER_70_245 ();
 sg13g2_fill_2 FILLER_70_252 ();
 sg13g2_fill_1 FILLER_70_254 ();
 sg13g2_fill_1 FILLER_70_270 ();
 sg13g2_decap_8 FILLER_70_323 ();
 sg13g2_decap_4 FILLER_70_335 ();
 sg13g2_fill_2 FILLER_70_339 ();
 sg13g2_decap_8 FILLER_70_367 ();
 sg13g2_decap_8 FILLER_70_374 ();
 sg13g2_fill_2 FILLER_70_381 ();
 sg13g2_fill_1 FILLER_70_383 ();
 sg13g2_fill_2 FILLER_70_396 ();
 sg13g2_fill_1 FILLER_70_419 ();
 sg13g2_decap_4 FILLER_70_425 ();
 sg13g2_fill_1 FILLER_70_429 ();
 sg13g2_decap_8 FILLER_71_26 ();
 sg13g2_decap_4 FILLER_71_33 ();
 sg13g2_fill_1 FILLER_71_37 ();
 sg13g2_fill_1 FILLER_71_42 ();
 sg13g2_decap_8 FILLER_71_48 ();
 sg13g2_decap_4 FILLER_71_55 ();
 sg13g2_fill_1 FILLER_71_80 ();
 sg13g2_fill_1 FILLER_71_138 ();
 sg13g2_fill_1 FILLER_71_143 ();
 sg13g2_fill_2 FILLER_71_190 ();
 sg13g2_fill_2 FILLER_71_218 ();
 sg13g2_fill_2 FILLER_71_223 ();
 sg13g2_fill_1 FILLER_71_225 ();
 sg13g2_decap_8 FILLER_71_230 ();
 sg13g2_decap_4 FILLER_71_237 ();
 sg13g2_decap_8 FILLER_71_246 ();
 sg13g2_decap_8 FILLER_71_253 ();
 sg13g2_decap_4 FILLER_71_260 ();
 sg13g2_fill_2 FILLER_71_264 ();
 sg13g2_decap_4 FILLER_71_274 ();
 sg13g2_decap_8 FILLER_71_282 ();
 sg13g2_decap_8 FILLER_71_289 ();
 sg13g2_fill_1 FILLER_71_300 ();
 sg13g2_fill_2 FILLER_71_306 ();
 sg13g2_fill_1 FILLER_71_308 ();
 sg13g2_decap_8 FILLER_71_325 ();
 sg13g2_decap_8 FILLER_71_332 ();
 sg13g2_decap_8 FILLER_71_339 ();
 sg13g2_decap_8 FILLER_71_363 ();
 sg13g2_fill_1 FILLER_71_370 ();
 sg13g2_decap_4 FILLER_71_378 ();
 sg13g2_decap_8 FILLER_71_422 ();
 sg13g2_fill_1 FILLER_71_429 ();
 sg13g2_fill_1 FILLER_72_31 ();
 sg13g2_fill_2 FILLER_72_62 ();
 sg13g2_fill_1 FILLER_72_90 ();
 sg13g2_fill_2 FILLER_72_95 ();
 sg13g2_fill_2 FILLER_72_101 ();
 sg13g2_fill_1 FILLER_72_124 ();
 sg13g2_fill_2 FILLER_72_147 ();
 sg13g2_fill_2 FILLER_72_153 ();
 sg13g2_decap_4 FILLER_72_159 ();
 sg13g2_fill_1 FILLER_72_163 ();
 sg13g2_decap_4 FILLER_72_168 ();
 sg13g2_fill_1 FILLER_72_172 ();
 sg13g2_decap_8 FILLER_72_203 ();
 sg13g2_fill_1 FILLER_72_210 ();
 sg13g2_fill_2 FILLER_72_226 ();
 sg13g2_fill_1 FILLER_72_228 ();
 sg13g2_fill_1 FILLER_72_255 ();
 sg13g2_decap_8 FILLER_72_286 ();
 sg13g2_decap_4 FILLER_72_293 ();
 sg13g2_fill_1 FILLER_72_297 ();
 sg13g2_fill_2 FILLER_72_311 ();
 sg13g2_decap_4 FILLER_72_323 ();
 sg13g2_fill_1 FILLER_72_385 ();
 sg13g2_fill_2 FILLER_72_411 ();
 sg13g2_fill_2 FILLER_72_417 ();
 sg13g2_fill_1 FILLER_72_419 ();
 sg13g2_decap_4 FILLER_72_424 ();
 sg13g2_fill_2 FILLER_72_428 ();
 sg13g2_decap_4 FILLER_73_0 ();
 sg13g2_fill_2 FILLER_73_4 ();
 sg13g2_decap_4 FILLER_73_15 ();
 sg13g2_decap_8 FILLER_73_61 ();
 sg13g2_fill_2 FILLER_73_68 ();
 sg13g2_fill_1 FILLER_73_70 ();
 sg13g2_decap_8 FILLER_73_101 ();
 sg13g2_decap_4 FILLER_73_108 ();
 sg13g2_fill_1 FILLER_73_152 ();
 sg13g2_decap_8 FILLER_73_157 ();
 sg13g2_decap_8 FILLER_73_164 ();
 sg13g2_decap_8 FILLER_73_171 ();
 sg13g2_fill_2 FILLER_73_178 ();
 sg13g2_fill_1 FILLER_73_180 ();
 sg13g2_decap_8 FILLER_73_185 ();
 sg13g2_decap_8 FILLER_73_192 ();
 sg13g2_decap_8 FILLER_73_199 ();
 sg13g2_fill_2 FILLER_73_206 ();
 sg13g2_fill_2 FILLER_73_231 ();
 sg13g2_fill_2 FILLER_73_276 ();
 sg13g2_fill_1 FILLER_73_278 ();
 sg13g2_fill_1 FILLER_73_293 ();
 sg13g2_fill_2 FILLER_73_330 ();
 sg13g2_fill_2 FILLER_73_363 ();
 sg13g2_fill_1 FILLER_73_371 ();
 sg13g2_fill_2 FILLER_73_389 ();
 sg13g2_fill_1 FILLER_73_391 ();
 sg13g2_fill_1 FILLER_74_26 ();
 sg13g2_decap_4 FILLER_74_69 ();
 sg13g2_decap_8 FILLER_74_76 ();
 sg13g2_fill_1 FILLER_74_83 ();
 sg13g2_fill_1 FILLER_74_110 ();
 sg13g2_decap_4 FILLER_74_127 ();
 sg13g2_fill_2 FILLER_74_153 ();
 sg13g2_fill_1 FILLER_74_181 ();
 sg13g2_fill_1 FILLER_74_247 ();
 sg13g2_fill_1 FILLER_74_252 ();
 sg13g2_fill_1 FILLER_74_258 ();
 sg13g2_fill_1 FILLER_74_271 ();
 sg13g2_fill_2 FILLER_74_285 ();
 sg13g2_fill_1 FILLER_74_336 ();
 sg13g2_fill_1 FILLER_74_349 ();
 sg13g2_fill_1 FILLER_74_355 ();
 sg13g2_fill_1 FILLER_74_360 ();
 sg13g2_fill_1 FILLER_74_369 ();
 sg13g2_fill_1 FILLER_74_380 ();
 sg13g2_fill_2 FILLER_74_423 ();
 sg13g2_decap_8 FILLER_75_0 ();
 sg13g2_decap_8 FILLER_75_15 ();
 sg13g2_decap_8 FILLER_75_22 ();
 sg13g2_decap_4 FILLER_75_29 ();
 sg13g2_fill_2 FILLER_75_33 ();
 sg13g2_fill_2 FILLER_75_52 ();
 sg13g2_fill_1 FILLER_75_54 ();
 sg13g2_decap_4 FILLER_75_62 ();
 sg13g2_fill_2 FILLER_75_66 ();
 sg13g2_decap_8 FILLER_75_98 ();
 sg13g2_fill_2 FILLER_75_105 ();
 sg13g2_fill_1 FILLER_75_119 ();
 sg13g2_fill_1 FILLER_75_155 ();
 sg13g2_fill_2 FILLER_75_182 ();
 sg13g2_fill_1 FILLER_75_241 ();
 sg13g2_fill_1 FILLER_75_246 ();
 sg13g2_decap_8 FILLER_75_251 ();
 sg13g2_decap_4 FILLER_75_258 ();
 sg13g2_fill_2 FILLER_75_262 ();
 sg13g2_fill_2 FILLER_75_279 ();
 sg13g2_fill_1 FILLER_75_281 ();
 sg13g2_decap_4 FILLER_75_291 ();
 sg13g2_decap_4 FILLER_75_299 ();
 sg13g2_fill_2 FILLER_75_324 ();
 sg13g2_fill_1 FILLER_75_326 ();
 sg13g2_decap_8 FILLER_75_332 ();
 sg13g2_decap_4 FILLER_75_339 ();
 sg13g2_decap_8 FILLER_75_347 ();
 sg13g2_decap_8 FILLER_75_363 ();
 sg13g2_decap_8 FILLER_75_374 ();
 sg13g2_decap_8 FILLER_75_381 ();
 sg13g2_decap_8 FILLER_75_388 ();
 sg13g2_decap_4 FILLER_75_395 ();
 sg13g2_fill_1 FILLER_75_399 ();
 sg13g2_decap_8 FILLER_76_0 ();
 sg13g2_decap_8 FILLER_76_7 ();
 sg13g2_fill_1 FILLER_76_14 ();
 sg13g2_fill_1 FILLER_76_23 ();
 sg13g2_fill_2 FILLER_76_46 ();
 sg13g2_fill_1 FILLER_76_48 ();
 sg13g2_decap_8 FILLER_76_55 ();
 sg13g2_decap_8 FILLER_76_62 ();
 sg13g2_fill_2 FILLER_76_69 ();
 sg13g2_fill_1 FILLER_76_71 ();
 sg13g2_fill_2 FILLER_76_81 ();
 sg13g2_fill_2 FILLER_76_118 ();
 sg13g2_fill_2 FILLER_76_130 ();
 sg13g2_fill_1 FILLER_76_132 ();
 sg13g2_decap_8 FILLER_76_138 ();
 sg13g2_fill_2 FILLER_76_145 ();
 sg13g2_fill_1 FILLER_76_147 ();
 sg13g2_fill_2 FILLER_76_151 ();
 sg13g2_fill_1 FILLER_76_153 ();
 sg13g2_fill_2 FILLER_76_163 ();
 sg13g2_fill_1 FILLER_76_165 ();
 sg13g2_decap_8 FILLER_76_170 ();
 sg13g2_decap_8 FILLER_76_177 ();
 sg13g2_decap_4 FILLER_76_184 ();
 sg13g2_fill_1 FILLER_76_188 ();
 sg13g2_fill_1 FILLER_76_197 ();
 sg13g2_fill_2 FILLER_76_202 ();
 sg13g2_fill_1 FILLER_76_209 ();
 sg13g2_fill_1 FILLER_76_215 ();
 sg13g2_decap_8 FILLER_76_232 ();
 sg13g2_decap_8 FILLER_76_239 ();
 sg13g2_decap_8 FILLER_76_246 ();
 sg13g2_decap_8 FILLER_76_253 ();
 sg13g2_fill_2 FILLER_76_270 ();
 sg13g2_decap_4 FILLER_76_280 ();
 sg13g2_fill_1 FILLER_76_287 ();
 sg13g2_decap_8 FILLER_76_298 ();
 sg13g2_fill_1 FILLER_76_310 ();
 sg13g2_decap_8 FILLER_76_337 ();
 sg13g2_fill_1 FILLER_76_357 ();
 sg13g2_decap_4 FILLER_76_361 ();
 sg13g2_fill_2 FILLER_76_365 ();
 sg13g2_decap_4 FILLER_76_371 ();
 sg13g2_decap_8 FILLER_76_382 ();
 sg13g2_decap_8 FILLER_76_389 ();
 sg13g2_decap_8 FILLER_76_396 ();
 sg13g2_fill_2 FILLER_76_403 ();
 sg13g2_decap_8 FILLER_76_412 ();
 sg13g2_decap_8 FILLER_76_419 ();
 sg13g2_decap_4 FILLER_76_426 ();
 sg13g2_fill_1 FILLER_77_0 ();
 sg13g2_fill_2 FILLER_77_35 ();
 sg13g2_fill_1 FILLER_77_61 ();
 sg13g2_fill_1 FILLER_77_66 ();
 sg13g2_fill_2 FILLER_77_71 ();
 sg13g2_decap_4 FILLER_77_77 ();
 sg13g2_decap_4 FILLER_77_85 ();
 sg13g2_fill_2 FILLER_77_115 ();
 sg13g2_fill_1 FILLER_77_117 ();
 sg13g2_decap_8 FILLER_77_183 ();
 sg13g2_decap_8 FILLER_77_190 ();
 sg13g2_decap_8 FILLER_77_197 ();
 sg13g2_decap_8 FILLER_77_244 ();
 sg13g2_decap_4 FILLER_77_251 ();
 sg13g2_fill_1 FILLER_77_255 ();
 sg13g2_fill_2 FILLER_77_292 ();
 sg13g2_decap_4 FILLER_77_298 ();
 sg13g2_fill_2 FILLER_77_302 ();
 sg13g2_fill_1 FILLER_77_309 ();
 sg13g2_fill_1 FILLER_77_315 ();
 sg13g2_fill_1 FILLER_77_376 ();
 sg13g2_fill_1 FILLER_77_419 ();
 sg13g2_decap_4 FILLER_77_425 ();
 sg13g2_fill_1 FILLER_77_429 ();
 sg13g2_decap_4 FILLER_78_0 ();
 sg13g2_fill_1 FILLER_78_12 ();
 sg13g2_fill_1 FILLER_78_83 ();
 sg13g2_decap_8 FILLER_78_88 ();
 sg13g2_decap_8 FILLER_78_95 ();
 sg13g2_decap_8 FILLER_78_102 ();
 sg13g2_decap_8 FILLER_78_109 ();
 sg13g2_decap_4 FILLER_78_116 ();
 sg13g2_decap_8 FILLER_78_124 ();
 sg13g2_decap_4 FILLER_78_178 ();
 sg13g2_fill_2 FILLER_78_182 ();
 sg13g2_fill_1 FILLER_78_256 ();
 sg13g2_fill_2 FILLER_78_361 ();
 sg13g2_fill_2 FILLER_78_402 ();
 sg13g2_fill_1 FILLER_79_0 ();
 sg13g2_fill_1 FILLER_79_27 ();
 sg13g2_fill_1 FILLER_79_32 ();
 sg13g2_fill_2 FILLER_79_41 ();
 sg13g2_fill_2 FILLER_79_69 ();
 sg13g2_fill_1 FILLER_79_76 ();
 sg13g2_fill_1 FILLER_79_107 ();
 sg13g2_fill_1 FILLER_79_113 ();
 sg13g2_fill_2 FILLER_79_118 ();
 sg13g2_fill_1 FILLER_79_150 ();
 sg13g2_fill_2 FILLER_79_155 ();
 sg13g2_fill_1 FILLER_79_161 ();
 sg13g2_fill_2 FILLER_79_166 ();
 sg13g2_fill_2 FILLER_79_176 ();
 sg13g2_fill_1 FILLER_79_206 ();
 sg13g2_decap_8 FILLER_79_215 ();
 sg13g2_fill_2 FILLER_79_253 ();
 sg13g2_fill_1 FILLER_79_255 ();
 sg13g2_fill_1 FILLER_79_282 ();
 sg13g2_fill_2 FILLER_79_286 ();
 sg13g2_fill_1 FILLER_79_288 ();
 sg13g2_fill_1 FILLER_79_315 ();
 sg13g2_fill_2 FILLER_79_320 ();
 sg13g2_fill_1 FILLER_79_327 ();
 sg13g2_fill_2 FILLER_79_332 ();
 sg13g2_fill_2 FILLER_79_338 ();
 sg13g2_fill_2 FILLER_79_345 ();
 sg13g2_fill_1 FILLER_79_347 ();
 sg13g2_fill_2 FILLER_79_369 ();
 sg13g2_fill_1 FILLER_79_371 ();
 sg13g2_fill_2 FILLER_79_385 ();
 sg13g2_decap_8 FILLER_80_0 ();
 sg13g2_decap_8 FILLER_80_11 ();
 sg13g2_decap_8 FILLER_80_18 ();
 sg13g2_fill_2 FILLER_80_25 ();
 sg13g2_fill_1 FILLER_80_27 ();
 sg13g2_decap_8 FILLER_80_32 ();
 sg13g2_decap_8 FILLER_80_39 ();
 sg13g2_fill_2 FILLER_80_46 ();
 sg13g2_decap_8 FILLER_80_56 ();
 sg13g2_decap_8 FILLER_80_63 ();
 sg13g2_fill_2 FILLER_80_70 ();
 sg13g2_fill_1 FILLER_80_72 ();
 sg13g2_fill_2 FILLER_80_81 ();
 sg13g2_fill_1 FILLER_80_83 ();
 sg13g2_decap_4 FILLER_80_96 ();
 sg13g2_fill_2 FILLER_80_116 ();
 sg13g2_fill_2 FILLER_80_126 ();
 sg13g2_fill_1 FILLER_80_152 ();
 sg13g2_fill_2 FILLER_80_165 ();
 sg13g2_fill_1 FILLER_80_167 ();
 sg13g2_fill_2 FILLER_80_192 ();
 sg13g2_fill_1 FILLER_80_198 ();
 sg13g2_fill_1 FILLER_80_207 ();
 sg13g2_fill_2 FILLER_80_216 ();
 sg13g2_fill_2 FILLER_80_222 ();
 sg13g2_fill_1 FILLER_80_224 ();
 sg13g2_fill_1 FILLER_80_233 ();
 sg13g2_fill_1 FILLER_80_238 ();
 sg13g2_fill_1 FILLER_80_243 ();
 sg13g2_fill_1 FILLER_80_252 ();
 sg13g2_fill_2 FILLER_80_273 ();
 sg13g2_decap_8 FILLER_80_279 ();
 sg13g2_decap_8 FILLER_80_286 ();
 sg13g2_fill_2 FILLER_80_293 ();
 sg13g2_decap_8 FILLER_80_299 ();
 sg13g2_decap_8 FILLER_80_306 ();
 sg13g2_decap_8 FILLER_80_313 ();
 sg13g2_decap_8 FILLER_80_320 ();
 sg13g2_decap_8 FILLER_80_327 ();
 sg13g2_decap_4 FILLER_80_334 ();
 sg13g2_fill_1 FILLER_80_338 ();
 sg13g2_fill_2 FILLER_80_347 ();
 sg13g2_fill_2 FILLER_80_353 ();
 sg13g2_fill_1 FILLER_80_367 ();
 sg13g2_fill_2 FILLER_80_380 ();
 sg13g2_decap_4 FILLER_80_390 ();
 sg13g2_fill_1 FILLER_80_394 ();
 sg13g2_decap_4 FILLER_80_399 ();
 sg13g2_fill_1 FILLER_80_403 ();
 sg13g2_fill_2 FILLER_80_408 ();
 sg13g2_fill_1 FILLER_80_410 ();
 sg13g2_decap_8 FILLER_80_419 ();
 sg13g2_decap_4 FILLER_80_426 ();
endmodule
