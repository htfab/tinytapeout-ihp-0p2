module tt_um_htfab_bouncy_capsule (clk,
    ena,
    rst_n,
    ui_in,
    uio_in,
    uio_oe,
    uio_out,
    uo_out);
 input clk;
 input ena;
 input rst_n;
 input [7:0] ui_in;
 input [7:0] uio_in;
 output [7:0] uio_oe;
 output [7:0] uio_out;
 output [7:0] uo_out;

 wire _0000_;
 wire _0001_;
 wire _0002_;
 wire _0003_;
 wire _0004_;
 wire _0005_;
 wire _0006_;
 wire _0007_;
 wire _0008_;
 wire _0009_;
 wire _0010_;
 wire _0011_;
 wire _0012_;
 wire _0013_;
 wire _0014_;
 wire _0015_;
 wire _0016_;
 wire _0017_;
 wire _0018_;
 wire _0019_;
 wire _0020_;
 wire _0021_;
 wire _0022_;
 wire _0023_;
 wire _0024_;
 wire _0025_;
 wire _0026_;
 wire _0027_;
 wire _0028_;
 wire _0029_;
 wire _0030_;
 wire _0031_;
 wire _0032_;
 wire _0033_;
 wire _0034_;
 wire _0035_;
 wire _0036_;
 wire _0037_;
 wire _0038_;
 wire _0039_;
 wire _0040_;
 wire _0041_;
 wire _0042_;
 wire _0043_;
 wire _0044_;
 wire _0045_;
 wire _0046_;
 wire _0047_;
 wire _0048_;
 wire _0049_;
 wire _0050_;
 wire _0051_;
 wire _0052_;
 wire _0053_;
 wire _0054_;
 wire _0055_;
 wire _0056_;
 wire _0057_;
 wire _0058_;
 wire _0059_;
 wire _0060_;
 wire _0061_;
 wire _0062_;
 wire _0063_;
 wire _0064_;
 wire _0065_;
 wire _0066_;
 wire _0067_;
 wire _0068_;
 wire _0069_;
 wire _0070_;
 wire _0071_;
 wire _0072_;
 wire _0073_;
 wire _0074_;
 wire _0075_;
 wire _0076_;
 wire _0077_;
 wire _0078_;
 wire _0079_;
 wire _0080_;
 wire _0081_;
 wire _0082_;
 wire _0083_;
 wire _0084_;
 wire _0085_;
 wire _0086_;
 wire _0087_;
 wire _0088_;
 wire _0089_;
 wire _0090_;
 wire _0091_;
 wire _0092_;
 wire _0093_;
 wire _0094_;
 wire _0095_;
 wire _0096_;
 wire _0097_;
 wire _0098_;
 wire _0099_;
 wire _0100_;
 wire _0101_;
 wire _0102_;
 wire _0103_;
 wire _0104_;
 wire _0105_;
 wire _0106_;
 wire _0107_;
 wire _0108_;
 wire _0109_;
 wire _0110_;
 wire _0111_;
 wire _0112_;
 wire _0113_;
 wire _0114_;
 wire _0115_;
 wire _0116_;
 wire _0117_;
 wire _0118_;
 wire _0119_;
 wire _0120_;
 wire _0121_;
 wire _0122_;
 wire _0123_;
 wire _0124_;
 wire _0125_;
 wire _0126_;
 wire _0127_;
 wire _0128_;
 wire _0129_;
 wire _0130_;
 wire _0131_;
 wire _0132_;
 wire _0133_;
 wire _0134_;
 wire _0135_;
 wire _0136_;
 wire _0137_;
 wire _0138_;
 wire _0139_;
 wire _0140_;
 wire _0141_;
 wire _0142_;
 wire _0143_;
 wire _0144_;
 wire _0145_;
 wire _0146_;
 wire _0147_;
 wire _0148_;
 wire _0149_;
 wire _0150_;
 wire _0151_;
 wire _0152_;
 wire _0153_;
 wire _0154_;
 wire _0155_;
 wire _0156_;
 wire _0157_;
 wire _0158_;
 wire _0159_;
 wire _0160_;
 wire _0161_;
 wire _0162_;
 wire _0163_;
 wire _0164_;
 wire _0165_;
 wire _0166_;
 wire _0167_;
 wire _0168_;
 wire _0169_;
 wire _0170_;
 wire _0171_;
 wire _0172_;
 wire _0173_;
 wire _0174_;
 wire _0175_;
 wire _0176_;
 wire _0177_;
 wire _0178_;
 wire _0179_;
 wire _0180_;
 wire _0181_;
 wire _0182_;
 wire _0183_;
 wire _0184_;
 wire _0185_;
 wire _0186_;
 wire _0187_;
 wire _0188_;
 wire _0189_;
 wire _0190_;
 wire _0191_;
 wire _0192_;
 wire _0193_;
 wire _0194_;
 wire _0195_;
 wire _0196_;
 wire _0197_;
 wire _0198_;
 wire _0199_;
 wire _0200_;
 wire _0201_;
 wire _0202_;
 wire _0203_;
 wire _0204_;
 wire _0205_;
 wire _0206_;
 wire _0207_;
 wire _0208_;
 wire _0209_;
 wire _0210_;
 wire _0211_;
 wire _0212_;
 wire _0213_;
 wire _0214_;
 wire _0215_;
 wire _0216_;
 wire _0217_;
 wire _0218_;
 wire _0219_;
 wire _0220_;
 wire _0221_;
 wire _0222_;
 wire _0223_;
 wire _0224_;
 wire _0225_;
 wire _0226_;
 wire _0227_;
 wire _0228_;
 wire _0229_;
 wire _0230_;
 wire _0231_;
 wire _0232_;
 wire _0233_;
 wire _0234_;
 wire _0235_;
 wire _0236_;
 wire _0237_;
 wire _0238_;
 wire _0239_;
 wire _0240_;
 wire _0241_;
 wire _0242_;
 wire _0243_;
 wire _0244_;
 wire _0245_;
 wire _0246_;
 wire _0247_;
 wire _0248_;
 wire _0249_;
 wire _0250_;
 wire _0251_;
 wire _0252_;
 wire _0253_;
 wire _0254_;
 wire _0255_;
 wire _0256_;
 wire _0257_;
 wire _0258_;
 wire _0259_;
 wire _0260_;
 wire _0261_;
 wire _0262_;
 wire _0263_;
 wire _0264_;
 wire _0265_;
 wire _0266_;
 wire _0267_;
 wire _0268_;
 wire _0269_;
 wire _0270_;
 wire _0271_;
 wire _0272_;
 wire _0273_;
 wire _0274_;
 wire _0275_;
 wire _0276_;
 wire _0277_;
 wire _0278_;
 wire _0279_;
 wire _0280_;
 wire _0281_;
 wire _0282_;
 wire _0283_;
 wire _0284_;
 wire _0285_;
 wire _0286_;
 wire _0287_;
 wire _0288_;
 wire _0289_;
 wire _0290_;
 wire _0291_;
 wire _0292_;
 wire _0293_;
 wire _0294_;
 wire _0295_;
 wire _0296_;
 wire _0297_;
 wire _0298_;
 wire _0299_;
 wire _0300_;
 wire _0301_;
 wire _0302_;
 wire _0303_;
 wire _0304_;
 wire _0305_;
 wire _0306_;
 wire _0307_;
 wire _0308_;
 wire _0309_;
 wire _0310_;
 wire _0311_;
 wire _0312_;
 wire _0313_;
 wire _0314_;
 wire _0315_;
 wire _0316_;
 wire _0317_;
 wire _0318_;
 wire _0319_;
 wire _0320_;
 wire _0321_;
 wire _0322_;
 wire _0323_;
 wire _0324_;
 wire _0325_;
 wire _0326_;
 wire _0327_;
 wire _0328_;
 wire _0329_;
 wire _0330_;
 wire _0331_;
 wire _0332_;
 wire _0333_;
 wire _0334_;
 wire _0335_;
 wire _0336_;
 wire _0337_;
 wire _0338_;
 wire _0339_;
 wire _0340_;
 wire _0341_;
 wire _0342_;
 wire _0343_;
 wire _0344_;
 wire _0345_;
 wire _0346_;
 wire _0347_;
 wire _0348_;
 wire _0349_;
 wire _0350_;
 wire _0351_;
 wire _0352_;
 wire _0353_;
 wire _0354_;
 wire _0355_;
 wire _0356_;
 wire _0357_;
 wire _0358_;
 wire _0359_;
 wire _0360_;
 wire _0361_;
 wire _0362_;
 wire _0363_;
 wire _0364_;
 wire _0365_;
 wire _0366_;
 wire _0367_;
 wire _0368_;
 wire _0369_;
 wire _0370_;
 wire _0371_;
 wire _0372_;
 wire _0373_;
 wire _0374_;
 wire _0375_;
 wire _0376_;
 wire _0377_;
 wire _0378_;
 wire _0379_;
 wire _0380_;
 wire _0381_;
 wire _0382_;
 wire _0383_;
 wire _0384_;
 wire _0385_;
 wire _0386_;
 wire _0387_;
 wire _0388_;
 wire _0389_;
 wire _0390_;
 wire _0391_;
 wire _0392_;
 wire _0393_;
 wire _0394_;
 wire _0395_;
 wire _0396_;
 wire _0397_;
 wire _0398_;
 wire _0399_;
 wire _0400_;
 wire _0401_;
 wire _0402_;
 wire _0403_;
 wire _0404_;
 wire _0405_;
 wire _0406_;
 wire _0407_;
 wire _0408_;
 wire _0409_;
 wire _0410_;
 wire _0411_;
 wire _0412_;
 wire _0413_;
 wire _0414_;
 wire _0415_;
 wire _0416_;
 wire _0417_;
 wire _0418_;
 wire _0419_;
 wire _0420_;
 wire _0421_;
 wire _0422_;
 wire _0423_;
 wire _0424_;
 wire _0425_;
 wire _0426_;
 wire _0427_;
 wire _0428_;
 wire _0429_;
 wire _0430_;
 wire _0431_;
 wire _0432_;
 wire _0433_;
 wire _0434_;
 wire _0435_;
 wire _0436_;
 wire _0437_;
 wire _0438_;
 wire _0439_;
 wire _0440_;
 wire _0441_;
 wire _0442_;
 wire _0443_;
 wire _0444_;
 wire _0445_;
 wire _0446_;
 wire _0447_;
 wire _0448_;
 wire _0449_;
 wire _0450_;
 wire _0451_;
 wire _0452_;
 wire _0453_;
 wire _0454_;
 wire _0455_;
 wire _0456_;
 wire _0457_;
 wire _0458_;
 wire _0459_;
 wire _0460_;
 wire _0461_;
 wire _0462_;
 wire _0463_;
 wire _0464_;
 wire _0465_;
 wire _0466_;
 wire _0467_;
 wire _0468_;
 wire _0469_;
 wire _0470_;
 wire _0471_;
 wire _0472_;
 wire _0473_;
 wire _0474_;
 wire _0475_;
 wire _0476_;
 wire _0477_;
 wire _0478_;
 wire _0479_;
 wire _0480_;
 wire _0481_;
 wire _0482_;
 wire _0483_;
 wire _0484_;
 wire _0485_;
 wire _0486_;
 wire _0487_;
 wire _0488_;
 wire _0489_;
 wire _0490_;
 wire _0491_;
 wire _0492_;
 wire _0493_;
 wire _0494_;
 wire _0495_;
 wire _0496_;
 wire _0497_;
 wire _0498_;
 wire _0499_;
 wire _0500_;
 wire _0501_;
 wire _0502_;
 wire _0503_;
 wire _0504_;
 wire _0505_;
 wire _0506_;
 wire _0507_;
 wire _0508_;
 wire _0509_;
 wire _0510_;
 wire _0511_;
 wire _0512_;
 wire _0513_;
 wire _0514_;
 wire _0515_;
 wire _0516_;
 wire _0517_;
 wire _0518_;
 wire _0519_;
 wire _0520_;
 wire _0521_;
 wire _0522_;
 wire _0523_;
 wire _0524_;
 wire _0525_;
 wire _0526_;
 wire _0527_;
 wire _0528_;
 wire _0529_;
 wire _0530_;
 wire _0531_;
 wire _0532_;
 wire _0533_;
 wire _0534_;
 wire _0535_;
 wire _0536_;
 wire _0537_;
 wire _0538_;
 wire _0539_;
 wire _0540_;
 wire _0541_;
 wire _0542_;
 wire _0543_;
 wire _0544_;
 wire _0545_;
 wire _0546_;
 wire _0547_;
 wire _0548_;
 wire _0549_;
 wire _0550_;
 wire _0551_;
 wire _0552_;
 wire _0553_;
 wire _0554_;
 wire _0555_;
 wire _0556_;
 wire _0557_;
 wire _0558_;
 wire _0559_;
 wire _0560_;
 wire _0561_;
 wire _0562_;
 wire _0563_;
 wire _0564_;
 wire _0565_;
 wire _0566_;
 wire _0567_;
 wire _0568_;
 wire _0569_;
 wire _0570_;
 wire _0571_;
 wire _0572_;
 wire _0573_;
 wire _0574_;
 wire _0575_;
 wire _0576_;
 wire _0577_;
 wire _0578_;
 wire _0579_;
 wire _0580_;
 wire _0581_;
 wire _0582_;
 wire _0583_;
 wire _0584_;
 wire _0585_;
 wire _0586_;
 wire _0587_;
 wire _0588_;
 wire _0589_;
 wire _0590_;
 wire _0591_;
 wire _0592_;
 wire _0593_;
 wire _0594_;
 wire _0595_;
 wire _0596_;
 wire _0597_;
 wire _0598_;
 wire _0599_;
 wire _0600_;
 wire _0601_;
 wire _0602_;
 wire _0603_;
 wire _0604_;
 wire _0605_;
 wire _0606_;
 wire _0607_;
 wire _0608_;
 wire _0609_;
 wire _0610_;
 wire _0611_;
 wire _0612_;
 wire _0613_;
 wire _0614_;
 wire _0615_;
 wire _0616_;
 wire _0617_;
 wire _0618_;
 wire _0619_;
 wire _0620_;
 wire _0621_;
 wire _0622_;
 wire _0623_;
 wire _0624_;
 wire _0625_;
 wire _0626_;
 wire _0627_;
 wire _0628_;
 wire _0629_;
 wire _0630_;
 wire _0631_;
 wire _0632_;
 wire _0633_;
 wire _0634_;
 wire _0635_;
 wire _0636_;
 wire _0637_;
 wire _0638_;
 wire _0639_;
 wire _0640_;
 wire _0641_;
 wire _0642_;
 wire _0643_;
 wire _0644_;
 wire _0645_;
 wire _0646_;
 wire _0647_;
 wire _0648_;
 wire _0649_;
 wire _0650_;
 wire _0651_;
 wire _0652_;
 wire _0653_;
 wire _0654_;
 wire _0655_;
 wire _0656_;
 wire _0657_;
 wire _0658_;
 wire _0659_;
 wire _0660_;
 wire _0661_;
 wire _0662_;
 wire _0663_;
 wire _0664_;
 wire _0665_;
 wire _0666_;
 wire _0667_;
 wire _0668_;
 wire _0669_;
 wire _0670_;
 wire _0671_;
 wire _0672_;
 wire _0673_;
 wire _0674_;
 wire _0675_;
 wire _0676_;
 wire _0677_;
 wire _0678_;
 wire _0679_;
 wire _0680_;
 wire _0681_;
 wire _0682_;
 wire _0683_;
 wire _0684_;
 wire _0685_;
 wire _0686_;
 wire _0687_;
 wire _0688_;
 wire _0689_;
 wire _0690_;
 wire _0691_;
 wire _0692_;
 wire _0693_;
 wire _0694_;
 wire _0695_;
 wire _0696_;
 wire _0697_;
 wire _0698_;
 wire _0699_;
 wire _0700_;
 wire _0701_;
 wire _0702_;
 wire _0703_;
 wire _0704_;
 wire _0705_;
 wire _0706_;
 wire _0707_;
 wire _0708_;
 wire _0709_;
 wire _0710_;
 wire _0711_;
 wire _0712_;
 wire _0713_;
 wire _0714_;
 wire _0715_;
 wire _0716_;
 wire _0717_;
 wire _0718_;
 wire _0719_;
 wire _0720_;
 wire _0721_;
 wire _0722_;
 wire _0723_;
 wire _0724_;
 wire _0725_;
 wire _0726_;
 wire _0727_;
 wire _0728_;
 wire _0729_;
 wire _0730_;
 wire _0731_;
 wire _0732_;
 wire _0733_;
 wire _0734_;
 wire _0735_;
 wire _0736_;
 wire _0737_;
 wire _0738_;
 wire _0739_;
 wire _0740_;
 wire _0741_;
 wire _0742_;
 wire _0743_;
 wire _0744_;
 wire _0745_;
 wire _0746_;
 wire _0747_;
 wire _0748_;
 wire _0749_;
 wire _0750_;
 wire _0751_;
 wire _0752_;
 wire _0753_;
 wire _0754_;
 wire _0755_;
 wire _0756_;
 wire _0757_;
 wire _0758_;
 wire _0759_;
 wire _0760_;
 wire _0761_;
 wire _0762_;
 wire _0763_;
 wire _0764_;
 wire _0765_;
 wire _0766_;
 wire _0767_;
 wire _0768_;
 wire _0769_;
 wire _0770_;
 wire _0771_;
 wire _0772_;
 wire _0773_;
 wire _0774_;
 wire _0775_;
 wire _0776_;
 wire _0777_;
 wire _0778_;
 wire _0779_;
 wire _0780_;
 wire _0781_;
 wire _0782_;
 wire _0783_;
 wire _0784_;
 wire _0785_;
 wire _0786_;
 wire _0787_;
 wire _0788_;
 wire _0789_;
 wire _0790_;
 wire _0791_;
 wire _0792_;
 wire _0793_;
 wire _0794_;
 wire _0795_;
 wire _0796_;
 wire _0797_;
 wire _0798_;
 wire _0799_;
 wire _0800_;
 wire _0801_;
 wire _0802_;
 wire _0803_;
 wire _0804_;
 wire _0805_;
 wire _0806_;
 wire _0807_;
 wire _0808_;
 wire _0809_;
 wire _0810_;
 wire _0811_;
 wire _0812_;
 wire _0813_;
 wire _0814_;
 wire _0815_;
 wire _0816_;
 wire _0817_;
 wire _0818_;
 wire _0819_;
 wire _0820_;
 wire _0821_;
 wire _0822_;
 wire _0823_;
 wire _0824_;
 wire _0825_;
 wire _0826_;
 wire _0827_;
 wire _0828_;
 wire _0829_;
 wire _0830_;
 wire _0831_;
 wire _0832_;
 wire _0833_;
 wire _0834_;
 wire _0835_;
 wire _0836_;
 wire _0837_;
 wire _0838_;
 wire _0839_;
 wire _0840_;
 wire _0841_;
 wire _0842_;
 wire _0843_;
 wire _0844_;
 wire _0845_;
 wire _0846_;
 wire _0847_;
 wire _0848_;
 wire _0849_;
 wire _0850_;
 wire _0851_;
 wire _0852_;
 wire _0853_;
 wire _0854_;
 wire _0855_;
 wire _0856_;
 wire _0857_;
 wire _0858_;
 wire _0859_;
 wire _0860_;
 wire _0861_;
 wire _0862_;
 wire _0863_;
 wire _0864_;
 wire _0865_;
 wire _0866_;
 wire _0867_;
 wire _0868_;
 wire _0869_;
 wire _0870_;
 wire _0871_;
 wire _0872_;
 wire _0873_;
 wire _0874_;
 wire _0875_;
 wire _0876_;
 wire _0877_;
 wire _0878_;
 wire _0879_;
 wire _0880_;
 wire _0881_;
 wire _0882_;
 wire _0883_;
 wire _0884_;
 wire _0885_;
 wire _0886_;
 wire _0887_;
 wire _0888_;
 wire _0889_;
 wire _0890_;
 wire _0891_;
 wire _0892_;
 wire _0893_;
 wire _0894_;
 wire _0895_;
 wire _0896_;
 wire _0897_;
 wire _0898_;
 wire _0899_;
 wire _0900_;
 wire _0901_;
 wire _0902_;
 wire _0903_;
 wire _0904_;
 wire _0905_;
 wire _0906_;
 wire _0907_;
 wire _0908_;
 wire _0909_;
 wire _0910_;
 wire _0911_;
 wire _0912_;
 wire _0913_;
 wire _0914_;
 wire _0915_;
 wire _0916_;
 wire _0917_;
 wire _0918_;
 wire _0919_;
 wire _0920_;
 wire _0921_;
 wire _0922_;
 wire _0923_;
 wire _0924_;
 wire _0925_;
 wire _0926_;
 wire _0927_;
 wire _0928_;
 wire _0929_;
 wire _0930_;
 wire _0931_;
 wire _0932_;
 wire _0933_;
 wire _0934_;
 wire _0935_;
 wire _0936_;
 wire _0937_;
 wire _0938_;
 wire _0939_;
 wire _0940_;
 wire _0941_;
 wire _0942_;
 wire _0943_;
 wire _0944_;
 wire _0945_;
 wire _0946_;
 wire _0947_;
 wire _0948_;
 wire _0949_;
 wire _0950_;
 wire _0951_;
 wire _0952_;
 wire _0953_;
 wire _0954_;
 wire _0955_;
 wire _0956_;
 wire _0957_;
 wire _0958_;
 wire _0959_;
 wire _0960_;
 wire _0961_;
 wire _0962_;
 wire _0963_;
 wire _0964_;
 wire _0965_;
 wire _0966_;
 wire _0967_;
 wire _0968_;
 wire _0969_;
 wire _0970_;
 wire _0971_;
 wire _0972_;
 wire _0973_;
 wire _0974_;
 wire _0975_;
 wire _0976_;
 wire _0977_;
 wire _0978_;
 wire _0979_;
 wire _0980_;
 wire _0981_;
 wire _0982_;
 wire _0983_;
 wire _0984_;
 wire _0985_;
 wire _0986_;
 wire _0987_;
 wire _0988_;
 wire _0989_;
 wire _0990_;
 wire _0991_;
 wire _0992_;
 wire _0993_;
 wire _0994_;
 wire _0995_;
 wire _0996_;
 wire _0997_;
 wire _0998_;
 wire _0999_;
 wire _1000_;
 wire _1001_;
 wire _1002_;
 wire _1003_;
 wire _1004_;
 wire _1005_;
 wire _1006_;
 wire _1007_;
 wire _1008_;
 wire _1009_;
 wire _1010_;
 wire _1011_;
 wire _1012_;
 wire _1013_;
 wire _1014_;
 wire _1015_;
 wire _1016_;
 wire _1017_;
 wire _1018_;
 wire _1019_;
 wire _1020_;
 wire _1021_;
 wire _1022_;
 wire _1023_;
 wire _1024_;
 wire _1025_;
 wire _1026_;
 wire _1027_;
 wire _1028_;
 wire _1029_;
 wire _1030_;
 wire _1031_;
 wire _1032_;
 wire _1033_;
 wire _1034_;
 wire _1035_;
 wire _1036_;
 wire _1037_;
 wire _1038_;
 wire _1039_;
 wire _1040_;
 wire _1041_;
 wire _1042_;
 wire _1043_;
 wire _1044_;
 wire _1045_;
 wire _1046_;
 wire _1047_;
 wire _1048_;
 wire _1049_;
 wire _1050_;
 wire _1051_;
 wire _1052_;
 wire _1053_;
 wire _1054_;
 wire _1055_;
 wire _1056_;
 wire _1057_;
 wire _1058_;
 wire _1059_;
 wire _1060_;
 wire _1061_;
 wire _1062_;
 wire _1063_;
 wire _1064_;
 wire _1065_;
 wire _1066_;
 wire _1067_;
 wire _1068_;
 wire _1069_;
 wire _1070_;
 wire _1071_;
 wire _1072_;
 wire _1073_;
 wire _1074_;
 wire _1075_;
 wire _1076_;
 wire _1077_;
 wire _1078_;
 wire _1079_;
 wire _1080_;
 wire _1081_;
 wire _1082_;
 wire _1083_;
 wire _1084_;
 wire _1085_;
 wire _1086_;
 wire _1087_;
 wire _1088_;
 wire _1089_;
 wire _1090_;
 wire _1091_;
 wire _1092_;
 wire _1093_;
 wire _1094_;
 wire _1095_;
 wire _1096_;
 wire _1097_;
 wire _1098_;
 wire _1099_;
 wire _1100_;
 wire _1101_;
 wire _1102_;
 wire _1103_;
 wire _1104_;
 wire _1105_;
 wire _1106_;
 wire _1107_;
 wire _1108_;
 wire _1109_;
 wire _1110_;
 wire _1111_;
 wire _1112_;
 wire _1113_;
 wire _1114_;
 wire _1115_;
 wire _1116_;
 wire _1117_;
 wire _1118_;
 wire _1119_;
 wire _1120_;
 wire _1121_;
 wire _1122_;
 wire _1123_;
 wire _1124_;
 wire _1125_;
 wire _1126_;
 wire _1127_;
 wire _1128_;
 wire _1129_;
 wire _1130_;
 wire _1131_;
 wire _1132_;
 wire _1133_;
 wire _1134_;
 wire _1135_;
 wire _1136_;
 wire _1137_;
 wire _1138_;
 wire _1139_;
 wire _1140_;
 wire _1141_;
 wire _1142_;
 wire _1143_;
 wire _1144_;
 wire _1145_;
 wire _1146_;
 wire _1147_;
 wire _1148_;
 wire _1149_;
 wire _1150_;
 wire _1151_;
 wire _1152_;
 wire _1153_;
 wire _1154_;
 wire _1155_;
 wire _1156_;
 wire _1157_;
 wire _1158_;
 wire _1159_;
 wire _1160_;
 wire _1161_;
 wire _1162_;
 wire _1163_;
 wire _1164_;
 wire _1165_;
 wire _1166_;
 wire _1167_;
 wire _1168_;
 wire _1169_;
 wire _1170_;
 wire _1171_;
 wire _1172_;
 wire _1173_;
 wire _1174_;
 wire _1175_;
 wire _1176_;
 wire _1177_;
 wire _1178_;
 wire _1179_;
 wire _1180_;
 wire _1181_;
 wire _1182_;
 wire _1183_;
 wire _1184_;
 wire _1185_;
 wire _1186_;
 wire _1187_;
 wire _1188_;
 wire _1189_;
 wire _1190_;
 wire _1191_;
 wire _1192_;
 wire _1193_;
 wire _1194_;
 wire _1195_;
 wire _1196_;
 wire _1197_;
 wire _1198_;
 wire _1199_;
 wire _1200_;
 wire _1201_;
 wire _1202_;
 wire _1203_;
 wire _1204_;
 wire _1205_;
 wire _1206_;
 wire _1207_;
 wire _1208_;
 wire _1209_;
 wire _1210_;
 wire _1211_;
 wire _1212_;
 wire _1213_;
 wire _1214_;
 wire _1215_;
 wire _1216_;
 wire _1217_;
 wire _1218_;
 wire _1219_;
 wire _1220_;
 wire _1221_;
 wire _1222_;
 wire _1223_;
 wire _1224_;
 wire _1225_;
 wire _1226_;
 wire _1227_;
 wire _1228_;
 wire _1229_;
 wire _1230_;
 wire _1231_;
 wire _1232_;
 wire _1233_;
 wire _1234_;
 wire _1235_;
 wire _1236_;
 wire _1237_;
 wire _1238_;
 wire _1239_;
 wire _1240_;
 wire _1241_;
 wire _1242_;
 wire _1243_;
 wire _1244_;
 wire _1245_;
 wire _1246_;
 wire _1247_;
 wire _1248_;
 wire _1249_;
 wire _1250_;
 wire _1251_;
 wire _1252_;
 wire _1253_;
 wire _1254_;
 wire _1255_;
 wire _1256_;
 wire _1257_;
 wire _1258_;
 wire _1259_;
 wire _1260_;
 wire _1261_;
 wire _1262_;
 wire _1263_;
 wire _1264_;
 wire _1265_;
 wire _1266_;
 wire _1267_;
 wire _1268_;
 wire _1269_;
 wire _1270_;
 wire _1271_;
 wire _1272_;
 wire _1273_;
 wire _1274_;
 wire _1275_;
 wire _1276_;
 wire _1277_;
 wire _1278_;
 wire _1279_;
 wire _1280_;
 wire _1281_;
 wire _1282_;
 wire _1283_;
 wire _1284_;
 wire _1285_;
 wire _1286_;
 wire _1287_;
 wire _1288_;
 wire _1289_;
 wire _1290_;
 wire _1291_;
 wire _1292_;
 wire _1293_;
 wire _1294_;
 wire _1295_;
 wire _1296_;
 wire _1297_;
 wire _1298_;
 wire _1299_;
 wire _1300_;
 wire _1301_;
 wire _1302_;
 wire _1303_;
 wire _1304_;
 wire _1305_;
 wire _1306_;
 wire _1307_;
 wire _1308_;
 wire _1309_;
 wire _1310_;
 wire _1311_;
 wire _1312_;
 wire _1313_;
 wire _1314_;
 wire _1315_;
 wire _1316_;
 wire _1317_;
 wire _1318_;
 wire _1319_;
 wire _1320_;
 wire _1321_;
 wire _1322_;
 wire _1323_;
 wire _1324_;
 wire _1325_;
 wire _1326_;
 wire _1327_;
 wire _1328_;
 wire _1329_;
 wire _1330_;
 wire _1331_;
 wire _1332_;
 wire _1333_;
 wire _1334_;
 wire _1335_;
 wire _1336_;
 wire _1337_;
 wire _1338_;
 wire _1339_;
 wire _1340_;
 wire _1341_;
 wire _1342_;
 wire _1343_;
 wire _1344_;
 wire _1345_;
 wire _1346_;
 wire _1347_;
 wire _1348_;
 wire _1349_;
 wire _1350_;
 wire _1351_;
 wire _1352_;
 wire _1353_;
 wire _1354_;
 wire _1355_;
 wire _1356_;
 wire _1357_;
 wire _1358_;
 wire _1359_;
 wire _1360_;
 wire _1361_;
 wire _1362_;
 wire _1363_;
 wire _1364_;
 wire _1365_;
 wire _1366_;
 wire _1367_;
 wire _1368_;
 wire _1369_;
 wire _1370_;
 wire _1371_;
 wire _1372_;
 wire _1373_;
 wire _1374_;
 wire _1375_;
 wire _1376_;
 wire _1377_;
 wire _1378_;
 wire _1379_;
 wire _1380_;
 wire _1381_;
 wire _1382_;
 wire _1383_;
 wire _1384_;
 wire _1385_;
 wire _1386_;
 wire _1387_;
 wire _1388_;
 wire _1389_;
 wire _1390_;
 wire _1391_;
 wire _1392_;
 wire _1393_;
 wire _1394_;
 wire _1395_;
 wire _1396_;
 wire _1397_;
 wire _1398_;
 wire _1399_;
 wire _1400_;
 wire _1401_;
 wire _1402_;
 wire _1403_;
 wire _1404_;
 wire _1405_;
 wire _1406_;
 wire _1407_;
 wire _1408_;
 wire _1409_;
 wire _1410_;
 wire _1411_;
 wire _1412_;
 wire _1413_;
 wire _1414_;
 wire _1415_;
 wire _1416_;
 wire _1417_;
 wire _1418_;
 wire _1419_;
 wire _1420_;
 wire _1421_;
 wire _1422_;
 wire _1423_;
 wire _1424_;
 wire _1425_;
 wire _1426_;
 wire _1427_;
 wire _1428_;
 wire _1429_;
 wire _1430_;
 wire _1431_;
 wire _1432_;
 wire _1433_;
 wire _1434_;
 wire _1435_;
 wire _1436_;
 wire _1437_;
 wire _1438_;
 wire _1439_;
 wire _1440_;
 wire _1441_;
 wire _1442_;
 wire _1443_;
 wire _1444_;
 wire _1445_;
 wire _1446_;
 wire _1447_;
 wire _1448_;
 wire _1449_;
 wire _1450_;
 wire _1451_;
 wire _1452_;
 wire _1453_;
 wire _1454_;
 wire _1455_;
 wire _1456_;
 wire _1457_;
 wire _1458_;
 wire _1459_;
 wire _1460_;
 wire _1461_;
 wire _1462_;
 wire _1463_;
 wire _1464_;
 wire _1465_;
 wire _1466_;
 wire _1467_;
 wire _1468_;
 wire _1469_;
 wire _1470_;
 wire _1471_;
 wire _1472_;
 wire _1473_;
 wire _1474_;
 wire _1475_;
 wire _1476_;
 wire _1477_;
 wire _1478_;
 wire _1479_;
 wire _1480_;
 wire _1481_;
 wire _1482_;
 wire _1483_;
 wire _1484_;
 wire _1485_;
 wire _1486_;
 wire _1487_;
 wire _1488_;
 wire _1489_;
 wire _1490_;
 wire _1491_;
 wire _1492_;
 wire _1493_;
 wire _1494_;
 wire _1495_;
 wire _1496_;
 wire _1497_;
 wire _1498_;
 wire _1499_;
 wire _1500_;
 wire _1501_;
 wire _1502_;
 wire _1503_;
 wire _1504_;
 wire _1505_;
 wire _1506_;
 wire _1507_;
 wire _1508_;
 wire _1509_;
 wire _1510_;
 wire _1511_;
 wire _1512_;
 wire _1513_;
 wire _1514_;
 wire _1515_;
 wire _1516_;
 wire _1517_;
 wire _1518_;
 wire _1519_;
 wire _1520_;
 wire _1521_;
 wire _1522_;
 wire _1523_;
 wire _1524_;
 wire _1525_;
 wire _1526_;
 wire _1527_;
 wire _1528_;
 wire _1529_;
 wire _1530_;
 wire _1531_;
 wire _1532_;
 wire _1533_;
 wire _1534_;
 wire _1535_;
 wire _1536_;
 wire _1537_;
 wire _1538_;
 wire _1539_;
 wire _1540_;
 wire _1541_;
 wire _1542_;
 wire _1543_;
 wire _1544_;
 wire _1545_;
 wire _1546_;
 wire _1547_;
 wire _1548_;
 wire _1549_;
 wire _1550_;
 wire _1551_;
 wire _1552_;
 wire _1553_;
 wire _1554_;
 wire _1555_;
 wire _1556_;
 wire _1557_;
 wire _1558_;
 wire _1559_;
 wire _1560_;
 wire _1561_;
 wire _1562_;
 wire _1563_;
 wire _1564_;
 wire _1565_;
 wire _1566_;
 wire _1567_;
 wire _1568_;
 wire _1569_;
 wire _1570_;
 wire _1571_;
 wire _1572_;
 wire _1573_;
 wire _1574_;
 wire _1575_;
 wire _1576_;
 wire _1577_;
 wire _1578_;
 wire _1579_;
 wire _1580_;
 wire _1581_;
 wire _1582_;
 wire _1583_;
 wire _1584_;
 wire _1585_;
 wire _1586_;
 wire _1587_;
 wire _1588_;
 wire _1589_;
 wire _1590_;
 wire _1591_;
 wire _1592_;
 wire _1593_;
 wire _1594_;
 wire _1595_;
 wire _1596_;
 wire _1597_;
 wire _1598_;
 wire _1599_;
 wire _1600_;
 wire _1601_;
 wire _1602_;
 wire _1603_;
 wire _1604_;
 wire _1605_;
 wire _1606_;
 wire _1607_;
 wire _1608_;
 wire _1609_;
 wire _1610_;
 wire _1611_;
 wire _1612_;
 wire _1613_;
 wire _1614_;
 wire _1615_;
 wire _1616_;
 wire _1617_;
 wire _1618_;
 wire _1619_;
 wire _1620_;
 wire _1621_;
 wire _1622_;
 wire _1623_;
 wire _1624_;
 wire _1625_;
 wire _1626_;
 wire _1627_;
 wire _1628_;
 wire _1629_;
 wire _1630_;
 wire _1631_;
 wire _1632_;
 wire _1633_;
 wire _1634_;
 wire _1635_;
 wire _1636_;
 wire _1637_;
 wire _1638_;
 wire _1639_;
 wire _1640_;
 wire _1641_;
 wire _1642_;
 wire _1643_;
 wire _1644_;
 wire _1645_;
 wire _1646_;
 wire _1647_;
 wire _1648_;
 wire _1649_;
 wire _1650_;
 wire _1651_;
 wire _1652_;
 wire _1653_;
 wire _1654_;
 wire _1655_;
 wire _1656_;
 wire _1657_;
 wire _1658_;
 wire _1659_;
 wire _1660_;
 wire _1661_;
 wire _1662_;
 wire _1663_;
 wire _1664_;
 wire _1665_;
 wire _1666_;
 wire _1667_;
 wire _1668_;
 wire _1669_;
 wire _1670_;
 wire _1671_;
 wire _1672_;
 wire _1673_;
 wire _1674_;
 wire _1675_;
 wire _1676_;
 wire _1677_;
 wire _1678_;
 wire _1679_;
 wire _1680_;
 wire _1681_;
 wire _1682_;
 wire _1683_;
 wire _1684_;
 wire _1685_;
 wire _1686_;
 wire _1687_;
 wire _1688_;
 wire _1689_;
 wire _1690_;
 wire _1691_;
 wire _1692_;
 wire _1693_;
 wire _1694_;
 wire _1695_;
 wire _1696_;
 wire _1697_;
 wire _1698_;
 wire _1699_;
 wire _1700_;
 wire _1701_;
 wire _1702_;
 wire _1703_;
 wire _1704_;
 wire _1705_;
 wire _1706_;
 wire _1707_;
 wire _1708_;
 wire _1709_;
 wire _1710_;
 wire _1711_;
 wire _1712_;
 wire _1713_;
 wire _1714_;
 wire _1715_;
 wire _1716_;
 wire _1717_;
 wire _1718_;
 wire _1719_;
 wire _1720_;
 wire _1721_;
 wire _1722_;
 wire _1723_;
 wire _1724_;
 wire _1725_;
 wire _1726_;
 wire _1727_;
 wire _1728_;
 wire _1729_;
 wire _1730_;
 wire _1731_;
 wire _1732_;
 wire _1733_;
 wire _1734_;
 wire _1735_;
 wire _1736_;
 wire _1737_;
 wire _1738_;
 wire _1739_;
 wire _1740_;
 wire _1741_;
 wire _1742_;
 wire _1743_;
 wire _1744_;
 wire _1745_;
 wire _1746_;
 wire _1747_;
 wire _1748_;
 wire _1749_;
 wire _1750_;
 wire _1751_;
 wire _1752_;
 wire _1753_;
 wire _1754_;
 wire _1755_;
 wire _1756_;
 wire _1757_;
 wire _1758_;
 wire _1759_;
 wire _1760_;
 wire _1761_;
 wire _1762_;
 wire _1763_;
 wire _1764_;
 wire _1765_;
 wire _1766_;
 wire _1767_;
 wire _1768_;
 wire _1769_;
 wire _1770_;
 wire _1771_;
 wire _1772_;
 wire _1773_;
 wire _1774_;
 wire _1775_;
 wire _1776_;
 wire _1777_;
 wire _1778_;
 wire _1779_;
 wire _1780_;
 wire _1781_;
 wire _1782_;
 wire _1783_;
 wire _1784_;
 wire _1785_;
 wire _1786_;
 wire _1787_;
 wire _1788_;
 wire _1789_;
 wire _1790_;
 wire _1791_;
 wire _1792_;
 wire _1793_;
 wire _1794_;
 wire _1795_;
 wire _1796_;
 wire _1797_;
 wire _1798_;
 wire _1799_;
 wire _1800_;
 wire _1801_;
 wire _1802_;
 wire _1803_;
 wire _1804_;
 wire _1805_;
 wire _1806_;
 wire _1807_;
 wire _1808_;
 wire _1809_;
 wire _1810_;
 wire _1811_;
 wire _1812_;
 wire _1813_;
 wire _1814_;
 wire _1815_;
 wire _1816_;
 wire _1817_;
 wire _1818_;
 wire _1819_;
 wire _1820_;
 wire _1821_;
 wire _1822_;
 wire _1823_;
 wire _1824_;
 wire _1825_;
 wire _1826_;
 wire _1827_;
 wire _1828_;
 wire _1829_;
 wire _1830_;
 wire _1831_;
 wire _1832_;
 wire _1833_;
 wire _1834_;
 wire _1835_;
 wire _1836_;
 wire _1837_;
 wire _1838_;
 wire _1839_;
 wire _1840_;
 wire _1841_;
 wire _1842_;
 wire _1843_;
 wire _1844_;
 wire _1845_;
 wire _1846_;
 wire _1847_;
 wire _1848_;
 wire _1849_;
 wire _1850_;
 wire _1851_;
 wire _1852_;
 wire _1853_;
 wire _1854_;
 wire _1855_;
 wire _1856_;
 wire _1857_;
 wire _1858_;
 wire _1859_;
 wire _1860_;
 wire _1861_;
 wire _1862_;
 wire _1863_;
 wire _1864_;
 wire _1865_;
 wire _1866_;
 wire _1867_;
 wire _1868_;
 wire _1869_;
 wire _1870_;
 wire _1871_;
 wire _1872_;
 wire _1873_;
 wire _1874_;
 wire _1875_;
 wire _1876_;
 wire _1877_;
 wire _1878_;
 wire _1879_;
 wire _1880_;
 wire _1881_;
 wire _1882_;
 wire _1883_;
 wire _1884_;
 wire _1885_;
 wire _1886_;
 wire _1887_;
 wire _1888_;
 wire _1889_;
 wire _1890_;
 wire _1891_;
 wire _1892_;
 wire _1893_;
 wire _1894_;
 wire _1895_;
 wire _1896_;
 wire _1897_;
 wire _1898_;
 wire _1899_;
 wire _1900_;
 wire _1901_;
 wire _1902_;
 wire _1903_;
 wire _1904_;
 wire _1905_;
 wire _1906_;
 wire _1907_;
 wire _1908_;
 wire _1909_;
 wire _1910_;
 wire _1911_;
 wire _1912_;
 wire _1913_;
 wire _1914_;
 wire _1915_;
 wire _1916_;
 wire _1917_;
 wire _1918_;
 wire _1919_;
 wire _1920_;
 wire _1921_;
 wire _1922_;
 wire _1923_;
 wire _1924_;
 wire _1925_;
 wire _1926_;
 wire _1927_;
 wire _1928_;
 wire _1929_;
 wire _1930_;
 wire _1931_;
 wire _1932_;
 wire _1933_;
 wire _1934_;
 wire _1935_;
 wire _1936_;
 wire _1937_;
 wire _1938_;
 wire _1939_;
 wire _1940_;
 wire _1941_;
 wire _1942_;
 wire _1943_;
 wire _1944_;
 wire _1945_;
 wire _1946_;
 wire _1947_;
 wire _1948_;
 wire _1949_;
 wire _1950_;
 wire _1951_;
 wire _1952_;
 wire _1953_;
 wire _1954_;
 wire _1955_;
 wire _1956_;
 wire _1957_;
 wire _1958_;
 wire _1959_;
 wire _1960_;
 wire _1961_;
 wire _1962_;
 wire _1963_;
 wire _1964_;
 wire _1965_;
 wire _1966_;
 wire _1967_;
 wire _1968_;
 wire _1969_;
 wire _1970_;
 wire _1971_;
 wire _1972_;
 wire _1973_;
 wire _1974_;
 wire _1975_;
 wire _1976_;
 wire _1977_;
 wire _1978_;
 wire _1979_;
 wire _1980_;
 wire _1981_;
 wire _1982_;
 wire _1983_;
 wire _1984_;
 wire _1985_;
 wire _1986_;
 wire _1987_;
 wire _1988_;
 wire _1989_;
 wire _1990_;
 wire _1991_;
 wire _1992_;
 wire _1993_;
 wire _1994_;
 wire _1995_;
 wire _1996_;
 wire _1997_;
 wire _1998_;
 wire _1999_;
 wire _2000_;
 wire _2001_;
 wire _2002_;
 wire _2003_;
 wire _2004_;
 wire _2005_;
 wire _2006_;
 wire _2007_;
 wire _2008_;
 wire _2009_;
 wire _2010_;
 wire _2011_;
 wire _2012_;
 wire _2013_;
 wire _2014_;
 wire _2015_;
 wire _2016_;
 wire _2017_;
 wire _2018_;
 wire _2019_;
 wire _2020_;
 wire _2021_;
 wire _2022_;
 wire _2023_;
 wire _2024_;
 wire _2025_;
 wire _2026_;
 wire _2027_;
 wire _2028_;
 wire _2029_;
 wire _2030_;
 wire _2031_;
 wire _2032_;
 wire _2033_;
 wire _2034_;
 wire _2035_;
 wire _2036_;
 wire _2037_;
 wire _2038_;
 wire _2039_;
 wire _2040_;
 wire _2041_;
 wire _2042_;
 wire _2043_;
 wire _2044_;
 wire _2045_;
 wire _2046_;
 wire _2047_;
 wire _2048_;
 wire _2049_;
 wire _2050_;
 wire _2051_;
 wire _2052_;
 wire _2053_;
 wire _2054_;
 wire _2055_;
 wire _2056_;
 wire _2057_;
 wire _2058_;
 wire _2059_;
 wire _2060_;
 wire _2061_;
 wire _2062_;
 wire _2063_;
 wire _2064_;
 wire _2065_;
 wire _2066_;
 wire _2067_;
 wire _2068_;
 wire _2069_;
 wire _2070_;
 wire _2071_;
 wire _2072_;
 wire _2073_;
 wire _2074_;
 wire _2075_;
 wire _2076_;
 wire _2077_;
 wire _2078_;
 wire _2079_;
 wire _2080_;
 wire _2081_;
 wire _2082_;
 wire _2083_;
 wire _2084_;
 wire _2085_;
 wire _2086_;
 wire _2087_;
 wire _2088_;
 wire _2089_;
 wire _2090_;
 wire _2091_;
 wire _2092_;
 wire _2093_;
 wire _2094_;
 wire _2095_;
 wire _2096_;
 wire _2097_;
 wire _2098_;
 wire _2099_;
 wire _2100_;
 wire _2101_;
 wire _2102_;
 wire _2103_;
 wire _2104_;
 wire _2105_;
 wire _2106_;
 wire _2107_;
 wire _2108_;
 wire _2109_;
 wire _2110_;
 wire _2111_;
 wire _2112_;
 wire _2113_;
 wire _2114_;
 wire _2115_;
 wire _2116_;
 wire _2117_;
 wire _2118_;
 wire _2119_;
 wire _2120_;
 wire _2121_;
 wire _2122_;
 wire _2123_;
 wire _2124_;
 wire _2125_;
 wire _2126_;
 wire _2127_;
 wire _2128_;
 wire _2129_;
 wire _2130_;
 wire _2131_;
 wire _2132_;
 wire _2133_;
 wire _2134_;
 wire _2135_;
 wire _2136_;
 wire _2137_;
 wire _2138_;
 wire _2139_;
 wire _2140_;
 wire _2141_;
 wire _2142_;
 wire _2143_;
 wire _2144_;
 wire _2145_;
 wire _2146_;
 wire _2147_;
 wire _2148_;
 wire _2149_;
 wire _2150_;
 wire _2151_;
 wire _2152_;
 wire _2153_;
 wire _2154_;
 wire _2155_;
 wire _2156_;
 wire _2157_;
 wire _2158_;
 wire _2159_;
 wire _2160_;
 wire _2161_;
 wire _2162_;
 wire _2163_;
 wire _2164_;
 wire _2165_;
 wire _2166_;
 wire _2167_;
 wire _2168_;
 wire _2169_;
 wire _2170_;
 wire _2171_;
 wire _2172_;
 wire _2173_;
 wire _2174_;
 wire _2175_;
 wire _2176_;
 wire _2177_;
 wire _2178_;
 wire _2179_;
 wire _2180_;
 wire _2181_;
 wire _2182_;
 wire _2183_;
 wire _2184_;
 wire _2185_;
 wire _2186_;
 wire _2187_;
 wire _2188_;
 wire _2189_;
 wire _2190_;
 wire _2191_;
 wire _2192_;
 wire _2193_;
 wire _2194_;
 wire _2195_;
 wire _2196_;
 wire _2197_;
 wire _2198_;
 wire _2199_;
 wire _2200_;
 wire _2201_;
 wire _2202_;
 wire _2203_;
 wire _2204_;
 wire _2205_;
 wire _2206_;
 wire _2207_;
 wire _2208_;
 wire _2209_;
 wire _2210_;
 wire _2211_;
 wire _2212_;
 wire _2213_;
 wire _2214_;
 wire _2215_;
 wire _2216_;
 wire _2217_;
 wire _2218_;
 wire _2219_;
 wire _2220_;
 wire _2221_;
 wire _2222_;
 wire _2223_;
 wire _2224_;
 wire _2225_;
 wire _2226_;
 wire _2227_;
 wire _2228_;
 wire _2229_;
 wire _2230_;
 wire _2231_;
 wire _2232_;
 wire _2233_;
 wire _2234_;
 wire _2235_;
 wire _2236_;
 wire _2237_;
 wire _2238_;
 wire _2239_;
 wire _2240_;
 wire _2241_;
 wire _2242_;
 wire _2243_;
 wire _2244_;
 wire _2245_;
 wire _2246_;
 wire _2247_;
 wire _2248_;
 wire _2249_;
 wire _2250_;
 wire _2251_;
 wire _2252_;
 wire _2253_;
 wire _2254_;
 wire _2255_;
 wire _2256_;
 wire _2257_;
 wire _2258_;
 wire _2259_;
 wire _2260_;
 wire _2261_;
 wire _2262_;
 wire _2263_;
 wire _2264_;
 wire _2265_;
 wire _2266_;
 wire _2267_;
 wire _2268_;
 wire _2269_;
 wire _2270_;
 wire _2271_;
 wire _2272_;
 wire _2273_;
 wire _2274_;
 wire _2275_;
 wire _2276_;
 wire _2277_;
 wire _2278_;
 wire _2279_;
 wire _2280_;
 wire _2281_;
 wire _2282_;
 wire _2283_;
 wire _2284_;
 wire _2285_;
 wire _2286_;
 wire _2287_;
 wire _2288_;
 wire _2289_;
 wire _2290_;
 wire _2291_;
 wire _2292_;
 wire _2293_;
 wire _2294_;
 wire _2295_;
 wire _2296_;
 wire _2297_;
 wire _2298_;
 wire _2299_;
 wire _2300_;
 wire _2301_;
 wire _2302_;
 wire _2303_;
 wire _2304_;
 wire _2305_;
 wire _2306_;
 wire _2307_;
 wire _2308_;
 wire _2309_;
 wire _2310_;
 wire _2311_;
 wire _2312_;
 wire _2313_;
 wire _2314_;
 wire _2315_;
 wire _2316_;
 wire _2317_;
 wire _2318_;
 wire _2319_;
 wire _2320_;
 wire _2321_;
 wire _2322_;
 wire _2323_;
 wire _2324_;
 wire _2325_;
 wire _2326_;
 wire _2327_;
 wire _2328_;
 wire _2329_;
 wire _2330_;
 wire _2331_;
 wire _2332_;
 wire _2333_;
 wire _2334_;
 wire _2335_;
 wire _2336_;
 wire _2337_;
 wire _2338_;
 wire _2339_;
 wire _2340_;
 wire _2341_;
 wire _2342_;
 wire _2343_;
 wire _2344_;
 wire _2345_;
 wire _2346_;
 wire _2347_;
 wire _2348_;
 wire _2349_;
 wire _2350_;
 wire _2351_;
 wire _2352_;
 wire _2353_;
 wire _2354_;
 wire _2355_;
 wire _2356_;
 wire _2357_;
 wire _2358_;
 wire _2359_;
 wire _2360_;
 wire _2361_;
 wire _2362_;
 wire _2363_;
 wire _2364_;
 wire _2365_;
 wire _2366_;
 wire _2367_;
 wire _2368_;
 wire _2369_;
 wire _2370_;
 wire _2371_;
 wire _2372_;
 wire _2373_;
 wire _2374_;
 wire _2375_;
 wire _2376_;
 wire _2377_;
 wire _2378_;
 wire _2379_;
 wire _2380_;
 wire _2381_;
 wire _2382_;
 wire _2383_;
 wire _2384_;
 wire _2385_;
 wire _2386_;
 wire _2387_;
 wire _2388_;
 wire _2389_;
 wire _2390_;
 wire _2391_;
 wire _2392_;
 wire _2393_;
 wire _2394_;
 wire _2395_;
 wire _2396_;
 wire _2397_;
 wire _2398_;
 wire _2399_;
 wire _2400_;
 wire _2401_;
 wire _2402_;
 wire _2403_;
 wire _2404_;
 wire _2405_;
 wire _2406_;
 wire _2407_;
 wire _2408_;
 wire _2409_;
 wire _2410_;
 wire _2411_;
 wire _2412_;
 wire _2413_;
 wire _2414_;
 wire _2415_;
 wire _2416_;
 wire _2417_;
 wire _2418_;
 wire _2419_;
 wire _2420_;
 wire _2421_;
 wire _2422_;
 wire _2423_;
 wire _2424_;
 wire _2425_;
 wire _2426_;
 wire _2427_;
 wire _2428_;
 wire _2429_;
 wire _2430_;
 wire _2431_;
 wire _2432_;
 wire _2433_;
 wire _2434_;
 wire _2435_;
 wire _2436_;
 wire _2437_;
 wire _2438_;
 wire _2439_;
 wire _2440_;
 wire _2441_;
 wire _2442_;
 wire _2443_;
 wire _2444_;
 wire _2445_;
 wire _2446_;
 wire _2447_;
 wire _2448_;
 wire _2449_;
 wire _2450_;
 wire _2451_;
 wire _2452_;
 wire _2453_;
 wire _2454_;
 wire _2455_;
 wire _2456_;
 wire _2457_;
 wire _2458_;
 wire _2459_;
 wire _2460_;
 wire _2461_;
 wire _2462_;
 wire _2463_;
 wire _2464_;
 wire _2465_;
 wire _2466_;
 wire _2467_;
 wire _2468_;
 wire _2469_;
 wire _2470_;
 wire _2471_;
 wire _2472_;
 wire _2473_;
 wire _2474_;
 wire _2475_;
 wire _2476_;
 wire _2477_;
 wire _2478_;
 wire _2479_;
 wire _2480_;
 wire _2481_;
 wire _2482_;
 wire _2483_;
 wire _2484_;
 wire _2485_;
 wire _2486_;
 wire _2487_;
 wire _2488_;
 wire _2489_;
 wire _2490_;
 wire _2491_;
 wire _2492_;
 wire _2493_;
 wire _2494_;
 wire _2495_;
 wire _2496_;
 wire _2497_;
 wire _2498_;
 wire _2499_;
 wire _2500_;
 wire _2501_;
 wire _2502_;
 wire _2503_;
 wire _2504_;
 wire _2505_;
 wire _2506_;
 wire _2507_;
 wire _2508_;
 wire _2509_;
 wire _2510_;
 wire _2511_;
 wire _2512_;
 wire _2513_;
 wire _2514_;
 wire _2515_;
 wire _2516_;
 wire _2517_;
 wire _2518_;
 wire _2519_;
 wire _2520_;
 wire _2521_;
 wire _2522_;
 wire _2523_;
 wire _2524_;
 wire _2525_;
 wire _2526_;
 wire _2527_;
 wire _2528_;
 wire _2529_;
 wire _2530_;
 wire _2531_;
 wire _2532_;
 wire _2533_;
 wire _2534_;
 wire _2535_;
 wire _2536_;
 wire _2537_;
 wire _2538_;
 wire _2539_;
 wire _2540_;
 wire _2541_;
 wire _2542_;
 wire _2543_;
 wire _2544_;
 wire _2545_;
 wire _2546_;
 wire _2547_;
 wire _2548_;
 wire _2549_;
 wire _2550_;
 wire _2551_;
 wire _2552_;
 wire _2553_;
 wire _2554_;
 wire _2555_;
 wire _2556_;
 wire _2557_;
 wire _2558_;
 wire _2559_;
 wire _2560_;
 wire _2561_;
 wire _2562_;
 wire _2563_;
 wire _2564_;
 wire _2565_;
 wire _2566_;
 wire _2567_;
 wire _2568_;
 wire _2569_;
 wire _2570_;
 wire _2571_;
 wire _2572_;
 wire _2573_;
 wire _2574_;
 wire _2575_;
 wire _2576_;
 wire _2577_;
 wire _2578_;
 wire _2579_;
 wire _2580_;
 wire _2581_;
 wire _2582_;
 wire _2583_;
 wire _2584_;
 wire _2585_;
 wire _2586_;
 wire _2587_;
 wire _2588_;
 wire _2589_;
 wire _2590_;
 wire _2591_;
 wire _2592_;
 wire _2593_;
 wire _2594_;
 wire _2595_;
 wire _2596_;
 wire _2597_;
 wire _2598_;
 wire _2599_;
 wire _2600_;
 wire _2601_;
 wire _2602_;
 wire _2603_;
 wire _2604_;
 wire _2605_;
 wire _2606_;
 wire _2607_;
 wire _2608_;
 wire _2609_;
 wire _2610_;
 wire _2611_;
 wire _2612_;
 wire _2613_;
 wire _2614_;
 wire _2615_;
 wire _2616_;
 wire _2617_;
 wire _2618_;
 wire _2619_;
 wire _2620_;
 wire _2621_;
 wire _2622_;
 wire _2623_;
 wire _2624_;
 wire _2625_;
 wire _2626_;
 wire _2627_;
 wire _2628_;
 wire _2629_;
 wire _2630_;
 wire _2631_;
 wire _2632_;
 wire _2633_;
 wire _2634_;
 wire _2635_;
 wire _2636_;
 wire _2637_;
 wire _2638_;
 wire _2639_;
 wire _2640_;
 wire _2641_;
 wire _2642_;
 wire _2643_;
 wire _2644_;
 wire _2645_;
 wire _2646_;
 wire _2647_;
 wire _2648_;
 wire _2649_;
 wire _2650_;
 wire _2651_;
 wire _2652_;
 wire _2653_;
 wire _2654_;
 wire _2655_;
 wire _2656_;
 wire _2657_;
 wire _2658_;
 wire _2659_;
 wire _2660_;
 wire _2661_;
 wire _2662_;
 wire _2663_;
 wire _2664_;
 wire _2665_;
 wire _2666_;
 wire _2667_;
 wire _2668_;
 wire _2669_;
 wire _2670_;
 wire _2671_;
 wire _2672_;
 wire _2673_;
 wire _2674_;
 wire _2675_;
 wire _2676_;
 wire _2677_;
 wire _2678_;
 wire _2679_;
 wire _2680_;
 wire _2681_;
 wire _2682_;
 wire _2683_;
 wire _2684_;
 wire _2685_;
 wire _2686_;
 wire _2687_;
 wire _2688_;
 wire _2689_;
 wire _2690_;
 wire _2691_;
 wire _2692_;
 wire _2693_;
 wire _2694_;
 wire _2695_;
 wire _2696_;
 wire _2697_;
 wire _2698_;
 wire _2699_;
 wire _2700_;
 wire _2701_;
 wire _2702_;
 wire _2703_;
 wire _2704_;
 wire _2705_;
 wire _2706_;
 wire _2707_;
 wire _2708_;
 wire _2709_;
 wire _2710_;
 wire _2711_;
 wire _2712_;
 wire _2713_;
 wire _2714_;
 wire _2715_;
 wire _2716_;
 wire _2717_;
 wire _2718_;
 wire _2719_;
 wire _2720_;
 wire _2721_;
 wire _2722_;
 wire _2723_;
 wire _2724_;
 wire _2725_;
 wire _2726_;
 wire _2727_;
 wire _2728_;
 wire _2729_;
 wire _2730_;
 wire _2731_;
 wire _2732_;
 wire _2733_;
 wire _2734_;
 wire _2735_;
 wire _2736_;
 wire _2737_;
 wire _2738_;
 wire _2739_;
 wire _2740_;
 wire _2741_;
 wire _2742_;
 wire _2743_;
 wire _2744_;
 wire _2745_;
 wire _2746_;
 wire _2747_;
 wire _2748_;
 wire _2749_;
 wire _2750_;
 wire _2751_;
 wire _2752_;
 wire _2753_;
 wire _2754_;
 wire _2755_;
 wire _2756_;
 wire _2757_;
 wire _2758_;
 wire _2759_;
 wire _2760_;
 wire _2761_;
 wire _2762_;
 wire _2763_;
 wire _2764_;
 wire _2765_;
 wire _2766_;
 wire _2767_;
 wire _2768_;
 wire _2769_;
 wire _2770_;
 wire _2771_;
 wire _2772_;
 wire _2773_;
 wire _2774_;
 wire _2775_;
 wire _2776_;
 wire _2777_;
 wire _2778_;
 wire _2779_;
 wire _2780_;
 wire _2781_;
 wire _2782_;
 wire _2783_;
 wire _2784_;
 wire _2785_;
 wire _2786_;
 wire _2787_;
 wire _2788_;
 wire _2789_;
 wire _2790_;
 wire _2791_;
 wire _2792_;
 wire _2793_;
 wire _2794_;
 wire _2795_;
 wire _2796_;
 wire _2797_;
 wire _2798_;
 wire _2799_;
 wire _2800_;
 wire _2801_;
 wire _2802_;
 wire _2803_;
 wire _2804_;
 wire _2805_;
 wire _2806_;
 wire _2807_;
 wire _2808_;
 wire _2809_;
 wire _2810_;
 wire _2811_;
 wire _2812_;
 wire _2813_;
 wire _2814_;
 wire _2815_;
 wire _2816_;
 wire _2817_;
 wire _2818_;
 wire _2819_;
 wire _2820_;
 wire _2821_;
 wire _2822_;
 wire _2823_;
 wire _2824_;
 wire _2825_;
 wire _2826_;
 wire _2827_;
 wire _2828_;
 wire _2829_;
 wire _2830_;
 wire _2831_;
 wire _2832_;
 wire _2833_;
 wire _2834_;
 wire _2835_;
 wire _2836_;
 wire _2837_;
 wire _2838_;
 wire _2839_;
 wire _2840_;
 wire _2841_;
 wire _2842_;
 wire _2843_;
 wire _2844_;
 wire _2845_;
 wire _2846_;
 wire _2847_;
 wire _2848_;
 wire _2849_;
 wire _2850_;
 wire _2851_;
 wire _2852_;
 wire _2853_;
 wire _2854_;
 wire _2855_;
 wire _2856_;
 wire _2857_;
 wire _2858_;
 wire _2859_;
 wire _2860_;
 wire _2861_;
 wire _2862_;
 wire _2863_;
 wire _2864_;
 wire _2865_;
 wire _2866_;
 wire _2867_;
 wire _2868_;
 wire _2869_;
 wire _2870_;
 wire _2871_;
 wire _2872_;
 wire _2873_;
 wire _2874_;
 wire _2875_;
 wire _2876_;
 wire _2877_;
 wire _2878_;
 wire _2879_;
 wire _2880_;
 wire _2881_;
 wire _2882_;
 wire _2883_;
 wire _2884_;
 wire _2885_;
 wire _2886_;
 wire _2887_;
 wire _2888_;
 wire _2889_;
 wire _2890_;
 wire _2891_;
 wire _2892_;
 wire _2893_;
 wire _2894_;
 wire _2895_;
 wire _2896_;
 wire _2897_;
 wire _2898_;
 wire _2899_;
 wire _2900_;
 wire _2901_;
 wire _2902_;
 wire _2903_;
 wire _2904_;
 wire _2905_;
 wire _2906_;
 wire _2907_;
 wire _2908_;
 wire _2909_;
 wire _2910_;
 wire _2911_;
 wire _2912_;
 wire _2913_;
 wire _2914_;
 wire _2915_;
 wire _2916_;
 wire _2917_;
 wire _2918_;
 wire _2919_;
 wire _2920_;
 wire _2921_;
 wire _2922_;
 wire _2923_;
 wire _2924_;
 wire _2925_;
 wire _2926_;
 wire _2927_;
 wire _2928_;
 wire _2929_;
 wire _2930_;
 wire _2931_;
 wire _2932_;
 wire _2933_;
 wire _2934_;
 wire _2935_;
 wire _2936_;
 wire _2937_;
 wire _2938_;
 wire _2939_;
 wire _2940_;
 wire _2941_;
 wire _2942_;
 wire _2943_;
 wire _2944_;
 wire _2945_;
 wire _2946_;
 wire _2947_;
 wire _2948_;
 wire _2949_;
 wire _2950_;
 wire _2951_;
 wire _2952_;
 wire _2953_;
 wire _2954_;
 wire _2955_;
 wire _2956_;
 wire _2957_;
 wire _2958_;
 wire _2959_;
 wire _2960_;
 wire _2961_;
 wire _2962_;
 wire _2963_;
 wire _2964_;
 wire _2965_;
 wire _2966_;
 wire _2967_;
 wire _2968_;
 wire _2969_;
 wire _2970_;
 wire _2971_;
 wire _2972_;
 wire _2973_;
 wire _2974_;
 wire _2975_;
 wire _2976_;
 wire _2977_;
 wire _2978_;
 wire _2979_;
 wire _2980_;
 wire _2981_;
 wire _2982_;
 wire _2983_;
 wire _2984_;
 wire _2985_;
 wire _2986_;
 wire _2987_;
 wire _2988_;
 wire _2989_;
 wire _2990_;
 wire _2991_;
 wire _2992_;
 wire _2993_;
 wire _2994_;
 wire _2995_;
 wire _2996_;
 wire _2997_;
 wire _2998_;
 wire _2999_;
 wire _3000_;
 wire _3001_;
 wire _3002_;
 wire _3003_;
 wire _3004_;
 wire _3005_;
 wire _3006_;
 wire _3007_;
 wire _3008_;
 wire _3009_;
 wire _3010_;
 wire _3011_;
 wire _3012_;
 wire _3013_;
 wire _3014_;
 wire _3015_;
 wire _3016_;
 wire _3017_;
 wire _3018_;
 wire _3019_;
 wire _3020_;
 wire _3021_;
 wire _3022_;
 wire _3023_;
 wire _3024_;
 wire _3025_;
 wire _3026_;
 wire _3027_;
 wire _3028_;
 wire _3029_;
 wire _3030_;
 wire _3031_;
 wire _3032_;
 wire _3033_;
 wire _3034_;
 wire _3035_;
 wire _3036_;
 wire _3037_;
 wire _3038_;
 wire _3039_;
 wire _3040_;
 wire _3041_;
 wire _3042_;
 wire _3043_;
 wire _3044_;
 wire _3045_;
 wire _3046_;
 wire _3047_;
 wire _3048_;
 wire _3049_;
 wire _3050_;
 wire _3051_;
 wire _3052_;
 wire _3053_;
 wire _3054_;
 wire _3055_;
 wire _3056_;
 wire _3057_;
 wire _3058_;
 wire _3059_;
 wire _3060_;
 wire _3061_;
 wire _3062_;
 wire _3063_;
 wire _3064_;
 wire _3065_;
 wire _3066_;
 wire _3067_;
 wire _3068_;
 wire _3069_;
 wire _3070_;
 wire _3071_;
 wire _3072_;
 wire _3073_;
 wire _3074_;
 wire _3075_;
 wire _3076_;
 wire _3077_;
 wire _3078_;
 wire _3079_;
 wire _3080_;
 wire _3081_;
 wire _3082_;
 wire _3083_;
 wire _3084_;
 wire _3085_;
 wire _3086_;
 wire _3087_;
 wire _3088_;
 wire _3089_;
 wire _3090_;
 wire _3091_;
 wire _3092_;
 wire _3093_;
 wire _3094_;
 wire _3095_;
 wire _3096_;
 wire _3097_;
 wire _3098_;
 wire _3099_;
 wire _3100_;
 wire _3101_;
 wire _3102_;
 wire _3103_;
 wire _3104_;
 wire _3105_;
 wire _3106_;
 wire _3107_;
 wire _3108_;
 wire _3109_;
 wire _3110_;
 wire _3111_;
 wire _3112_;
 wire _3113_;
 wire _3114_;
 wire _3115_;
 wire _3116_;
 wire _3117_;
 wire _3118_;
 wire _3119_;
 wire _3120_;
 wire _3121_;
 wire _3122_;
 wire _3123_;
 wire _3124_;
 wire _3125_;
 wire _3126_;
 wire _3127_;
 wire _3128_;
 wire _3129_;
 wire _3130_;
 wire _3131_;
 wire _3132_;
 wire _3133_;
 wire _3134_;
 wire _3135_;
 wire _3136_;
 wire _3137_;
 wire _3138_;
 wire _3139_;
 wire _3140_;
 wire _3141_;
 wire _3142_;
 wire _3143_;
 wire _3144_;
 wire _3145_;
 wire _3146_;
 wire _3147_;
 wire _3148_;
 wire _3149_;
 wire _3150_;
 wire _3151_;
 wire _3152_;
 wire _3153_;
 wire _3154_;
 wire _3155_;
 wire _3156_;
 wire _3157_;
 wire _3158_;
 wire _3159_;
 wire _3160_;
 wire _3161_;
 wire _3162_;
 wire _3163_;
 wire _3164_;
 wire _3165_;
 wire _3166_;
 wire _3167_;
 wire _3168_;
 wire _3169_;
 wire _3170_;
 wire _3171_;
 wire _3172_;
 wire _3173_;
 wire _3174_;
 wire _3175_;
 wire _3176_;
 wire _3177_;
 wire _3178_;
 wire _3179_;
 wire _3180_;
 wire _3181_;
 wire _3182_;
 wire _3183_;
 wire _3184_;
 wire _3185_;
 wire _3186_;
 wire _3187_;
 wire _3188_;
 wire _3189_;
 wire _3190_;
 wire _3191_;
 wire _3192_;
 wire _3193_;
 wire _3194_;
 wire _3195_;
 wire _3196_;
 wire _3197_;
 wire _3198_;
 wire _3199_;
 wire _3200_;
 wire _3201_;
 wire _3202_;
 wire _3203_;
 wire _3204_;
 wire _3205_;
 wire _3206_;
 wire _3207_;
 wire _3208_;
 wire _3209_;
 wire _3210_;
 wire _3211_;
 wire _3212_;
 wire _3213_;
 wire _3214_;
 wire _3215_;
 wire _3216_;
 wire _3217_;
 wire _3218_;
 wire _3219_;
 wire _3220_;
 wire _3221_;
 wire _3222_;
 wire _3223_;
 wire _3224_;
 wire _3225_;
 wire _3226_;
 wire _3227_;
 wire _3228_;
 wire _3229_;
 wire _3230_;
 wire _3231_;
 wire _3232_;
 wire _3233_;
 wire _3234_;
 wire _3235_;
 wire _3236_;
 wire _3237_;
 wire _3238_;
 wire _3239_;
 wire _3240_;
 wire _3241_;
 wire _3242_;
 wire _3243_;
 wire _3244_;
 wire _3245_;
 wire _3246_;
 wire _3247_;
 wire _3248_;
 wire _3249_;
 wire _3250_;
 wire _3251_;
 wire _3252_;
 wire _3253_;
 wire _3254_;
 wire _3255_;
 wire _3256_;
 wire _3257_;
 wire _3258_;
 wire _3259_;
 wire _3260_;
 wire _3261_;
 wire _3262_;
 wire _3263_;
 wire _3264_;
 wire _3265_;
 wire _3266_;
 wire _3267_;
 wire _3268_;
 wire _3269_;
 wire _3270_;
 wire _3271_;
 wire _3272_;
 wire _3273_;
 wire _3274_;
 wire _3275_;
 wire _3276_;
 wire _3277_;
 wire _3278_;
 wire _3279_;
 wire _3280_;
 wire _3281_;
 wire _3282_;
 wire _3283_;
 wire _3284_;
 wire _3285_;
 wire _3286_;
 wire _3287_;
 wire _3288_;
 wire _3289_;
 wire _3290_;
 wire _3291_;
 wire _3292_;
 wire _3293_;
 wire _3294_;
 wire _3295_;
 wire _3296_;
 wire _3297_;
 wire _3298_;
 wire _3299_;
 wire _3300_;
 wire _3301_;
 wire _3302_;
 wire _3303_;
 wire _3304_;
 wire _3305_;
 wire _3306_;
 wire _3307_;
 wire _3308_;
 wire _3309_;
 wire _3310_;
 wire _3311_;
 wire _3312_;
 wire _3313_;
 wire _3314_;
 wire _3315_;
 wire _3316_;
 wire _3317_;
 wire _3318_;
 wire _3319_;
 wire _3320_;
 wire _3321_;
 wire _3322_;
 wire _3323_;
 wire _3324_;
 wire _3325_;
 wire _3326_;
 wire _3327_;
 wire _3328_;
 wire _3329_;
 wire _3330_;
 wire _3331_;
 wire _3332_;
 wire _3333_;
 wire _3334_;
 wire _3335_;
 wire _3336_;
 wire _3337_;
 wire _3338_;
 wire _3339_;
 wire _3340_;
 wire _3341_;
 wire _3342_;
 wire _3343_;
 wire _3344_;
 wire _3345_;
 wire _3346_;
 wire _3347_;
 wire _3348_;
 wire _3349_;
 wire _3350_;
 wire _3351_;
 wire _3352_;
 wire _3353_;
 wire _3354_;
 wire _3355_;
 wire _3356_;
 wire _3357_;
 wire _3358_;
 wire _3359_;
 wire _3360_;
 wire _3361_;
 wire _3362_;
 wire _3363_;
 wire _3364_;
 wire _3365_;
 wire _3366_;
 wire _3367_;
 wire _3368_;
 wire _3369_;
 wire _3370_;
 wire _3371_;
 wire _3372_;
 wire _3373_;
 wire _3374_;
 wire _3375_;
 wire _3376_;
 wire _3377_;
 wire _3378_;
 wire _3379_;
 wire _3380_;
 wire _3381_;
 wire _3382_;
 wire _3383_;
 wire _3384_;
 wire _3385_;
 wire _3386_;
 wire _3387_;
 wire _3388_;
 wire _3389_;
 wire _3390_;
 wire _3391_;
 wire _3392_;
 wire _3393_;
 wire _3394_;
 wire _3395_;
 wire _3396_;
 wire _3397_;
 wire _3398_;
 wire _3399_;
 wire _3400_;
 wire _3401_;
 wire _3402_;
 wire _3403_;
 wire _3404_;
 wire _3405_;
 wire _3406_;
 wire _3407_;
 wire _3408_;
 wire _3409_;
 wire _3410_;
 wire _3411_;
 wire _3412_;
 wire _3413_;
 wire _3414_;
 wire _3415_;
 wire _3416_;
 wire _3417_;
 wire _3418_;
 wire _3419_;
 wire _3420_;
 wire _3421_;
 wire _3422_;
 wire _3423_;
 wire _3424_;
 wire _3425_;
 wire _3426_;
 wire _3427_;
 wire _3428_;
 wire _3429_;
 wire _3430_;
 wire _3431_;
 wire _3432_;
 wire _3433_;
 wire _3434_;
 wire _3435_;
 wire _3436_;
 wire _3437_;
 wire _3438_;
 wire _3439_;
 wire _3440_;
 wire _3441_;
 wire _3442_;
 wire _3443_;
 wire _3444_;
 wire _3445_;
 wire _3446_;
 wire _3447_;
 wire _3448_;
 wire _3449_;
 wire _3450_;
 wire _3451_;
 wire _3452_;
 wire _3453_;
 wire _3454_;
 wire _3455_;
 wire _3456_;
 wire _3457_;
 wire _3458_;
 wire _3459_;
 wire _3460_;
 wire _3461_;
 wire _3462_;
 wire _3463_;
 wire _3464_;
 wire _3465_;
 wire _3466_;
 wire _3467_;
 wire _3468_;
 wire _3469_;
 wire _3470_;
 wire _3471_;
 wire _3472_;
 wire _3473_;
 wire _3474_;
 wire _3475_;
 wire _3476_;
 wire _3477_;
 wire _3478_;
 wire _3479_;
 wire _3480_;
 wire _3481_;
 wire _3482_;
 wire _3483_;
 wire _3484_;
 wire _3485_;
 wire _3486_;
 wire _3487_;
 wire _3488_;
 wire _3489_;
 wire _3490_;
 wire _3491_;
 wire _3492_;
 wire _3493_;
 wire _3494_;
 wire _3495_;
 wire _3496_;
 wire _3497_;
 wire _3498_;
 wire _3499_;
 wire _3500_;
 wire _3501_;
 wire _3502_;
 wire _3503_;
 wire _3504_;
 wire _3505_;
 wire _3506_;
 wire _3507_;
 wire _3508_;
 wire _3509_;
 wire _3510_;
 wire _3511_;
 wire _3512_;
 wire _3513_;
 wire _3514_;
 wire _3515_;
 wire _3516_;
 wire _3517_;
 wire _3518_;
 wire _3519_;
 wire _3520_;
 wire _3521_;
 wire _3522_;
 wire _3523_;
 wire _3524_;
 wire _3525_;
 wire _3526_;
 wire _3527_;
 wire _3528_;
 wire _3529_;
 wire _3530_;
 wire _3531_;
 wire _3532_;
 wire _3533_;
 wire _3534_;
 wire _3535_;
 wire _3536_;
 wire _3537_;
 wire _3538_;
 wire _3539_;
 wire _3540_;
 wire _3541_;
 wire _3542_;
 wire _3543_;
 wire _3544_;
 wire _3545_;
 wire _3546_;
 wire _3547_;
 wire _3548_;
 wire _3549_;
 wire _3550_;
 wire _3551_;
 wire _3552_;
 wire _3553_;
 wire _3554_;
 wire _3555_;
 wire _3556_;
 wire _3557_;
 wire _3558_;
 wire _3559_;
 wire _3560_;
 wire _3561_;
 wire _3562_;
 wire _3563_;
 wire _3564_;
 wire _3565_;
 wire _3566_;
 wire _3567_;
 wire _3568_;
 wire _3569_;
 wire _3570_;
 wire _3571_;
 wire _3572_;
 wire _3573_;
 wire _3574_;
 wire _3575_;
 wire _3576_;
 wire _3577_;
 wire _3578_;
 wire _3579_;
 wire _3580_;
 wire _3581_;
 wire _3582_;
 wire _3583_;
 wire _3584_;
 wire _3585_;
 wire _3586_;
 wire _3587_;
 wire _3588_;
 wire _3589_;
 wire _3590_;
 wire _3591_;
 wire _3592_;
 wire _3593_;
 wire _3594_;
 wire _3595_;
 wire _3596_;
 wire _3597_;
 wire _3598_;
 wire _3599_;
 wire _3600_;
 wire _3601_;
 wire _3602_;
 wire _3603_;
 wire _3604_;
 wire _3605_;
 wire _3606_;
 wire _3607_;
 wire _3608_;
 wire _3609_;
 wire _3610_;
 wire _3611_;
 wire _3612_;
 wire _3613_;
 wire _3614_;
 wire _3615_;
 wire _3616_;
 wire _3617_;
 wire _3618_;
 wire _3619_;
 wire _3620_;
 wire _3621_;
 wire _3622_;
 wire _3623_;
 wire _3624_;
 wire _3625_;
 wire _3626_;
 wire _3627_;
 wire _3628_;
 wire _3629_;
 wire _3630_;
 wire _3631_;
 wire _3632_;
 wire _3633_;
 wire _3634_;
 wire _3635_;
 wire _3636_;
 wire _3637_;
 wire _3638_;
 wire _3639_;
 wire _3640_;
 wire _3641_;
 wire _3642_;
 wire _3643_;
 wire _3644_;
 wire _3645_;
 wire _3646_;
 wire _3647_;
 wire _3648_;
 wire _3649_;
 wire _3650_;
 wire _3651_;
 wire _3652_;
 wire _3653_;
 wire _3654_;
 wire _3655_;
 wire _3656_;
 wire _3657_;
 wire _3658_;
 wire _3659_;
 wire _3660_;
 wire _3661_;
 wire _3662_;
 wire _3663_;
 wire _3664_;
 wire _3665_;
 wire _3666_;
 wire _3667_;
 wire _3668_;
 wire _3669_;
 wire _3670_;
 wire _3671_;
 wire _3672_;
 wire _3673_;
 wire _3674_;
 wire _3675_;
 wire _3676_;
 wire _3677_;
 wire _3678_;
 wire _3679_;
 wire _3680_;
 wire _3681_;
 wire _3682_;
 wire _3683_;
 wire _3684_;
 wire _3685_;
 wire _3686_;
 wire _3687_;
 wire _3688_;
 wire _3689_;
 wire _3690_;
 wire _3691_;
 wire _3692_;
 wire _3693_;
 wire _3694_;
 wire _3695_;
 wire _3696_;
 wire _3697_;
 wire _3698_;
 wire _3699_;
 wire _3700_;
 wire _3701_;
 wire _3702_;
 wire _3703_;
 wire _3704_;
 wire _3705_;
 wire _3706_;
 wire _3707_;
 wire _3708_;
 wire _3709_;
 wire _3710_;
 wire _3711_;
 wire _3712_;
 wire _3713_;
 wire _3714_;
 wire _3715_;
 wire _3716_;
 wire _3717_;
 wire _3718_;
 wire _3719_;
 wire _3720_;
 wire _3721_;
 wire _3722_;
 wire _3723_;
 wire _3724_;
 wire _3725_;
 wire _3726_;
 wire _3727_;
 wire _3728_;
 wire _3729_;
 wire _3730_;
 wire _3731_;
 wire _3732_;
 wire _3733_;
 wire _3734_;
 wire _3735_;
 wire _3736_;
 wire _3737_;
 wire _3738_;
 wire _3739_;
 wire _3740_;
 wire _3741_;
 wire _3742_;
 wire _3743_;
 wire _3744_;
 wire _3745_;
 wire _3746_;
 wire _3747_;
 wire _3748_;
 wire _3749_;
 wire _3750_;
 wire _3751_;
 wire _3752_;
 wire _3753_;
 wire _3754_;
 wire _3755_;
 wire _3756_;
 wire _3757_;
 wire _3758_;
 wire _3759_;
 wire _3760_;
 wire _3761_;
 wire _3762_;
 wire _3763_;
 wire _3764_;
 wire _3765_;
 wire _3766_;
 wire _3767_;
 wire _3768_;
 wire _3769_;
 wire _3770_;
 wire _3771_;
 wire _3772_;
 wire _3773_;
 wire _3774_;
 wire _3775_;
 wire _3776_;
 wire _3777_;
 wire _3778_;
 wire _3779_;
 wire _3780_;
 wire _3781_;
 wire _3782_;
 wire _3783_;
 wire _3784_;
 wire _3785_;
 wire _3786_;
 wire _3787_;
 wire _3788_;
 wire _3789_;
 wire _3790_;
 wire _3791_;
 wire _3792_;
 wire _3793_;
 wire _3794_;
 wire _3795_;
 wire _3796_;
 wire _3797_;
 wire _3798_;
 wire _3799_;
 wire _3800_;
 wire _3801_;
 wire _3802_;
 wire _3803_;
 wire _3804_;
 wire _3805_;
 wire _3806_;
 wire _3807_;
 wire _3808_;
 wire _3809_;
 wire _3810_;
 wire _3811_;
 wire _3812_;
 wire _3813_;
 wire _3814_;
 wire _3815_;
 wire _3816_;
 wire _3817_;
 wire _3818_;
 wire _3819_;
 wire _3820_;
 wire _3821_;
 wire _3822_;
 wire _3823_;
 wire _3824_;
 wire _3825_;
 wire _3826_;
 wire _3827_;
 wire _3828_;
 wire _3829_;
 wire _3830_;
 wire _3831_;
 wire _3832_;
 wire _3833_;
 wire _3834_;
 wire _3835_;
 wire _3836_;
 wire _3837_;
 wire _3838_;
 wire _3839_;
 wire _3840_;
 wire _3841_;
 wire _3842_;
 wire _3843_;
 wire _3844_;
 wire _3845_;
 wire _3846_;
 wire _3847_;
 wire _3848_;
 wire _3849_;
 wire _3850_;
 wire _3851_;
 wire _3852_;
 wire _3853_;
 wire _3854_;
 wire _3855_;
 wire _3856_;
 wire _3857_;
 wire _3858_;
 wire _3859_;
 wire _3860_;
 wire _3861_;
 wire _3862_;
 wire _3863_;
 wire _3864_;
 wire _3865_;
 wire _3866_;
 wire _3867_;
 wire _3868_;
 wire _3869_;
 wire _3870_;
 wire _3871_;
 wire _3872_;
 wire _3873_;
 wire _3874_;
 wire _3875_;
 wire _3876_;
 wire _3877_;
 wire _3878_;
 wire _3879_;
 wire _3880_;
 wire _3881_;
 wire _3882_;
 wire _3883_;
 wire _3884_;
 wire _3885_;
 wire _3886_;
 wire _3887_;
 wire _3888_;
 wire _3889_;
 wire _3890_;
 wire _3891_;
 wire _3892_;
 wire _3893_;
 wire _3894_;
 wire _3895_;
 wire _3896_;
 wire _3897_;
 wire _3898_;
 wire _3899_;
 wire _3900_;
 wire _3901_;
 wire _3902_;
 wire _3903_;
 wire _3904_;
 wire _3905_;
 wire _3906_;
 wire _3907_;
 wire _3908_;
 wire _3909_;
 wire _3910_;
 wire _3911_;
 wire _3912_;
 wire _3913_;
 wire _3914_;
 wire _3915_;
 wire _3916_;
 wire _3917_;
 wire _3918_;
 wire _3919_;
 wire _3920_;
 wire _3921_;
 wire _3922_;
 wire _3923_;
 wire _3924_;
 wire _3925_;
 wire _3926_;
 wire _3927_;
 wire _3928_;
 wire _3929_;
 wire _3930_;
 wire _3931_;
 wire _3932_;
 wire _3933_;
 wire _3934_;
 wire _3935_;
 wire _3936_;
 wire _3937_;
 wire _3938_;
 wire _3939_;
 wire _3940_;
 wire _3941_;
 wire _3942_;
 wire _3943_;
 wire _3944_;
 wire _3945_;
 wire _3946_;
 wire _3947_;
 wire _3948_;
 wire _3949_;
 wire _3950_;
 wire _3951_;
 wire _3952_;
 wire _3953_;
 wire _3954_;
 wire _3955_;
 wire _3956_;
 wire _3957_;
 wire _3958_;
 wire _3959_;
 wire _3960_;
 wire _3961_;
 wire _3962_;
 wire _3963_;
 wire _3964_;
 wire _3965_;
 wire _3966_;
 wire _3967_;
 wire _3968_;
 wire _3969_;
 wire _3970_;
 wire _3971_;
 wire _3972_;
 wire _3973_;
 wire _3974_;
 wire _3975_;
 wire _3976_;
 wire _3977_;
 wire _3978_;
 wire _3979_;
 wire _3980_;
 wire _3981_;
 wire _3982_;
 wire _3983_;
 wire _3984_;
 wire _3985_;
 wire _3986_;
 wire _3987_;
 wire _3988_;
 wire _3989_;
 wire _3990_;
 wire _3991_;
 wire _3992_;
 wire _3993_;
 wire _3994_;
 wire _3995_;
 wire _3996_;
 wire _3997_;
 wire _3998_;
 wire _3999_;
 wire _4000_;
 wire _4001_;
 wire _4002_;
 wire _4003_;
 wire _4004_;
 wire _4005_;
 wire _4006_;
 wire _4007_;
 wire _4008_;
 wire _4009_;
 wire _4010_;
 wire _4011_;
 wire _4012_;
 wire _4013_;
 wire _4014_;
 wire _4015_;
 wire _4016_;
 wire _4017_;
 wire _4018_;
 wire _4019_;
 wire _4020_;
 wire _4021_;
 wire _4022_;
 wire _4023_;
 wire _4024_;
 wire _4025_;
 wire _4026_;
 wire _4027_;
 wire _4028_;
 wire _4029_;
 wire _4030_;
 wire _4031_;
 wire _4032_;
 wire _4033_;
 wire _4034_;
 wire _4035_;
 wire _4036_;
 wire _4037_;
 wire _4038_;
 wire _4039_;
 wire _4040_;
 wire _4041_;
 wire _4042_;
 wire _4043_;
 wire _4044_;
 wire _4045_;
 wire _4046_;
 wire _4047_;
 wire _4048_;
 wire _4049_;
 wire _4050_;
 wire _4051_;
 wire _4052_;
 wire _4053_;
 wire _4054_;
 wire _4055_;
 wire _4056_;
 wire _4057_;
 wire _4058_;
 wire _4059_;
 wire _4060_;
 wire _4061_;
 wire _4062_;
 wire _4063_;
 wire _4064_;
 wire _4065_;
 wire _4066_;
 wire _4067_;
 wire _4068_;
 wire _4069_;
 wire _4070_;
 wire _4071_;
 wire _4072_;
 wire _4073_;
 wire _4074_;
 wire _4075_;
 wire _4076_;
 wire _4077_;
 wire _4078_;
 wire _4079_;
 wire _4080_;
 wire _4081_;
 wire _4082_;
 wire _4083_;
 wire _4084_;
 wire _4085_;
 wire _4086_;
 wire _4087_;
 wire _4088_;
 wire _4089_;
 wire _4090_;
 wire _4091_;
 wire _4092_;
 wire _4093_;
 wire _4094_;
 wire _4095_;
 wire _4096_;
 wire _4097_;
 wire _4098_;
 wire _4099_;
 wire _4100_;
 wire _4101_;
 wire _4102_;
 wire _4103_;
 wire _4104_;
 wire _4105_;
 wire _4106_;
 wire _4107_;
 wire _4108_;
 wire _4109_;
 wire _4110_;
 wire _4111_;
 wire _4112_;
 wire _4113_;
 wire _4114_;
 wire _4115_;
 wire _4116_;
 wire _4117_;
 wire _4118_;
 wire _4119_;
 wire _4120_;
 wire _4121_;
 wire clknet_leaf_0_clk;
 wire bitmap_pixel;
 wire \capsule_color[0] ;
 wire \capsule_color[1] ;
 wire \capsule_color[2] ;
 wire \capsule_color[3] ;
 wire \capsule_color[4] ;
 wire \capsule_color[5] ;
 wire \center_x[0] ;
 wire \center_x[1] ;
 wire \center_x[2] ;
 wire \center_x[3] ;
 wire \center_x[4] ;
 wire \center_x[5] ;
 wire \center_x[6] ;
 wire \center_x[7] ;
 wire \center_x[8] ;
 wire \center_x[9] ;
 wire \center_y[0] ;
 wire \center_y[1] ;
 wire \center_y[2] ;
 wire \center_y[3] ;
 wire \center_y[4] ;
 wire \center_y[5] ;
 wire \center_y[6] ;
 wire \center_y[7] ;
 wire \center_y[8] ;
 wire \center_y[9] ;
 wire \collision_impact[0] ;
 wire \collision_impact[1] ;
 wire \color_entropy[0] ;
 wire \color_entropy[1] ;
 wire handle_impact;
 wire hsync;
 wire \i_bitmap.in[0] ;
 wire \i_bitmap.in[10] ;
 wire \i_bitmap.in[11] ;
 wire \i_bitmap.in[12] ;
 wire \i_bitmap.in[1] ;
 wire \i_bitmap.in[2] ;
 wire \i_bitmap.in[3] ;
 wire \i_bitmap.in[4] ;
 wire \i_bitmap.in[5] ;
 wire \i_bitmap.in[6] ;
 wire \i_bitmap.in[7] ;
 wire \i_bitmap.in[8] ;
 wire \i_bitmap.in[9] ;
 wire \i_capsule.tf_x[0] ;
 wire \i_capsule.tf_x[8] ;
 wire \i_capsule.tf_x[9] ;
 wire \i_capsule.tf_y[0] ;
 wire \i_capsule.tf_y[7] ;
 wire \i_capsule.tf_y[8] ;
 wire \i_capsule.tf_y[9] ;
 wire \i_collision.i_coll_table.in[0] ;
 wire \i_collision.i_coll_table.in[1] ;
 wire \i_collision.i_coll_table.in[3] ;
 wire \i_collision.i_coll_table.in[4] ;
 wire \i_collision.i_coll_table.in[5] ;
 wire \i_collision.mirror ;
 wire \i_collision.phi[1] ;
 wire \i_collision.rotate ;
 wire \i_collision.update ;
 wire \i_collision.vx[0] ;
 wire \i_collision.vx[1] ;
 wire \i_collision.vx[2] ;
 wire \i_collision.vy[0] ;
 wire \i_collision.vy[1] ;
 wire \i_collision.vy[2] ;
 wire \i_colors.channel[0] ;
 wire \i_colors.channel[1] ;
 wire \i_colors.channel[2] ;
 wire \i_delta_sigma.acc[0] ;
 wire \i_delta_sigma.acc[10] ;
 wire \i_delta_sigma.acc[11] ;
 wire \i_delta_sigma.acc[12] ;
 wire \i_delta_sigma.acc[13] ;
 wire \i_delta_sigma.acc[1] ;
 wire \i_delta_sigma.acc[2] ;
 wire \i_delta_sigma.acc[3] ;
 wire \i_delta_sigma.acc[4] ;
 wire \i_delta_sigma.acc[5] ;
 wire \i_delta_sigma.acc[6] ;
 wire \i_delta_sigma.acc[7] ;
 wire \i_delta_sigma.acc[8] ;
 wire \i_delta_sigma.acc[9] ;
 wire \i_delta_sigma.sample[0] ;
 wire \i_delta_sigma.sample[10] ;
 wire \i_delta_sigma.sample[11] ;
 wire \i_delta_sigma.sample[1] ;
 wire \i_delta_sigma.sample[2] ;
 wire \i_delta_sigma.sample[3] ;
 wire \i_delta_sigma.sample[4] ;
 wire \i_delta_sigma.sample[5] ;
 wire \i_delta_sigma.sample[6] ;
 wire \i_delta_sigma.sample[7] ;
 wire \i_delta_sigma.sample[8] ;
 wire \i_delta_sigma.sample[9] ;
 wire \i_kinematics.center_x_lo[0] ;
 wire \i_kinematics.center_x_lo[1] ;
 wire \i_kinematics.center_y_lo[0] ;
 wire \i_kinematics.center_y_lo[1] ;
 wire \i_kinematics.phi[0] ;
 wire \i_kinematics.phi[10] ;
 wire \i_kinematics.phi[1] ;
 wire \i_kinematics.phi[2] ;
 wire \i_kinematics.phi[3] ;
 wire \i_kinematics.phi[4] ;
 wire \i_kinematics.phi[5] ;
 wire \i_kinematics.phi[6] ;
 wire \i_kinematics.phi[7] ;
 wire \i_kinematics.update ;
 wire \i_orchestrator.hit_bottom ;
 wire \i_orchestrator.hit_left ;
 wire \i_orchestrator.hit_priority[0] ;
 wire \i_orchestrator.hit_priority[1] ;
 wire \i_orchestrator.hit_right ;
 wire \i_orchestrator.hit_top ;
 wire \i_orchestrator.lfsr[1] ;
 wire \i_orchestrator.lfsr[2] ;
 wire \i_orchestrator.lfsr[3] ;
 wire \i_orchestrator.lfsr[4] ;
 wire \i_orchestrator.lfsr[5] ;
 wire \i_orchestrator.lfsr[6] ;
 wire \i_orchestrator.lfsr[7] ;
 wire \i_orchestrator.sample_counter[0] ;
 wire \i_orchestrator.sample_counter[1] ;
 wire \i_orchestrator.sample_counter[2] ;
 wire \i_orchestrator.sample_counter[3] ;
 wire \i_orchestrator.sample_counter[4] ;
 wire \i_orchestrator.sample_counter[5] ;
 wire \i_orchestrator.sample_counter[6] ;
 wire \i_orchestrator.sample_counter[7] ;
 wire \i_orchestrator.sample_counter[8] ;
 wire \i_orchestrator.sample_counter[9] ;
 wire \i_orchestrator.tension[1] ;
 wire \i_orchestrator.tension[2] ;
 wire \i_orchestrator.tension[3] ;
 wire \i_orchestrator.trigger_debounce ;
 wire \i_orchestrator.trigger_resonator[0] ;
 wire \i_orchestrator.trigger_resonator[1] ;
 wire \i_orchestrator.update_resonator ;
 wire \i_orchestrator.update_transform ;
 wire \i_orchestrator.vga_x[0] ;
 wire \i_orchestrator.vga_x[1] ;
 wire \i_orchestrator.vga_x[2] ;
 wire \i_orchestrator.vga_x[3] ;
 wire \i_orchestrator.vga_x[4] ;
 wire \i_orchestrator.vga_x[5] ;
 wire \i_orchestrator.vga_x[6] ;
 wire \i_orchestrator.vga_x[7] ;
 wire \i_orchestrator.vga_x[8] ;
 wire \i_orchestrator.vga_x[9] ;
 wire \i_orchestrator.vga_y[0] ;
 wire \i_orchestrator.vga_y[1] ;
 wire \i_orchestrator.vga_y[2] ;
 wire \i_orchestrator.vga_y[3] ;
 wire \i_orchestrator.vga_y[4] ;
 wire \i_orchestrator.vga_y[5] ;
 wire \i_orchestrator.vga_y[6] ;
 wire \i_orchestrator.vga_y[7] ;
 wire \i_orchestrator.vga_y[8] ;
 wire \i_orchestrator.vga_y[9] ;
 wire \i_resonator.counter[0] ;
 wire \i_resonator.counter[1] ;
 wire \i_resonator.counter[2] ;
 wire \i_resonator.counter[3] ;
 wire \i_resonator.v[0] ;
 wire \i_resonator.v[10] ;
 wire \i_resonator.v[11] ;
 wire \i_resonator.v[12] ;
 wire \i_resonator.v[13] ;
 wire \i_resonator.v[14] ;
 wire \i_resonator.v[15] ;
 wire \i_resonator.v[1] ;
 wire \i_resonator.v[2] ;
 wire \i_resonator.v[3] ;
 wire \i_resonator.v[4] ;
 wire \i_resonator.v[5] ;
 wire \i_resonator.v[6] ;
 wire \i_resonator.v[7] ;
 wire \i_resonator.v[8] ;
 wire \i_resonator.v[9] ;
 wire \i_transform.image_x[0] ;
 wire \i_transform.image_x[1] ;
 wire \i_transform.image_x[2] ;
 wire \i_transform.image_x[3] ;
 wire \i_transform.image_x[4] ;
 wire \i_transform.image_x[5] ;
 wire \i_transform.image_y[0] ;
 wire \i_transform.image_y[1] ;
 wire \i_transform.image_y[2] ;
 wire \i_transform.image_y[3] ;
 wire \i_transform.image_y[4] ;
 wire \i_transform.image_y[5] ;
 wire \i_transform.track_x[0] ;
 wire \i_transform.track_x[1] ;
 wire \i_transform.track_x[2] ;
 wire \i_transform.track_x[3] ;
 wire \i_transform.track_x[4] ;
 wire \i_transform.track_x[5] ;
 wire \i_transform.track_x[6] ;
 wire \i_transform.track_x[7] ;
 wire \i_transform.track_x[8] ;
 wire \i_transform.track_x[9] ;
 wire \i_transform.track_y[0] ;
 wire \i_transform.track_y[1] ;
 wire \i_transform.track_y[2] ;
 wire \i_transform.track_y[3] ;
 wire \i_transform.track_y[4] ;
 wire \i_transform.track_y[5] ;
 wire \i_transform.track_y[6] ;
 wire \i_transform.track_y[7] ;
 wire \i_transform.track_y[8] ;
 wire \i_transform.track_y[9] ;
 wire \i_vga_beam.vsync ;
 wire orient;
 wire pdm_out;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net180;
 wire net181;
 wire net182;
 wire net183;
 wire net184;
 wire net185;
 wire net186;
 wire net187;
 wire net188;
 wire net189;
 wire net190;
 wire net191;
 wire net192;
 wire net193;
 wire net194;
 wire net195;
 wire net196;
 wire net197;
 wire net198;
 wire net199;
 wire net200;
 wire net201;
 wire net202;
 wire net203;
 wire net204;
 wire net205;
 wire net206;
 wire net207;
 wire net208;
 wire net209;
 wire net210;
 wire net211;
 wire net212;
 wire net213;
 wire net214;
 wire net215;
 wire net216;
 wire net217;
 wire net218;
 wire net219;
 wire net220;
 wire net221;
 wire net222;
 wire net223;
 wire net224;
 wire net225;
 wire net226;
 wire net227;
 wire net228;
 wire net229;
 wire net230;
 wire net231;
 wire net232;
 wire net233;
 wire net234;
 wire net235;
 wire net236;
 wire net237;
 wire net238;
 wire net239;
 wire net240;
 wire net241;
 wire net242;
 wire net243;
 wire net244;
 wire net245;
 wire net246;
 wire net247;
 wire net248;
 wire net249;
 wire net250;
 wire net251;
 wire net252;
 wire net253;
 wire net254;
 wire net255;
 wire net256;
 wire net257;
 wire net258;
 wire net259;
 wire net260;
 wire net261;
 wire net262;
 wire net263;
 wire net264;
 wire net265;
 wire net266;
 wire net267;
 wire net268;
 wire net269;
 wire net270;
 wire net271;
 wire net272;
 wire net273;
 wire net274;
 wire net275;
 wire net276;
 wire net277;
 wire net278;
 wire net279;
 wire net280;
 wire net281;
 wire net282;
 wire net283;
 wire net284;
 wire net285;
 wire net286;
 wire net287;
 wire net288;
 wire net289;
 wire net290;
 wire net291;
 wire net292;
 wire net293;
 wire net294;
 wire net295;
 wire net296;
 wire net297;
 wire net298;
 wire net299;
 wire net300;
 wire net301;
 wire net302;
 wire net303;
 wire net304;
 wire net305;
 wire net306;
 wire net307;
 wire net308;
 wire net309;
 wire net310;
 wire net311;
 wire net312;
 wire net313;
 wire net314;
 wire net315;
 wire net316;
 wire net317;
 wire net318;
 wire net319;
 wire net320;
 wire net321;
 wire net322;
 wire net323;
 wire net324;
 wire net325;
 wire net326;
 wire net327;
 wire net328;
 wire net329;
 wire net330;
 wire net331;
 wire net332;
 wire net333;
 wire net334;
 wire net335;
 wire net336;
 wire net337;
 wire net338;
 wire net339;
 wire net340;
 wire net341;
 wire net342;
 wire net343;
 wire net344;
 wire net345;
 wire net346;
 wire net347;
 wire net348;
 wire net349;
 wire net350;
 wire net351;
 wire net352;
 wire net353;
 wire net354;
 wire net355;
 wire net356;
 wire net357;
 wire net358;
 wire net359;
 wire net360;
 wire net361;
 wire net362;
 wire net363;
 wire net364;
 wire net365;
 wire net366;
 wire net367;
 wire net368;
 wire net369;
 wire net370;
 wire net371;
 wire net372;
 wire net373;
 wire net374;
 wire net375;
 wire net376;
 wire net377;
 wire net378;
 wire net379;
 wire net380;
 wire net381;
 wire net382;
 wire net383;
 wire net384;
 wire net385;
 wire net386;
 wire net387;
 wire net388;
 wire net389;
 wire net390;
 wire net391;
 wire net392;
 wire net393;
 wire net394;
 wire net395;
 wire net396;
 wire net397;
 wire net398;
 wire net399;
 wire net400;
 wire net401;
 wire net402;
 wire net403;
 wire net404;
 wire net405;
 wire net406;
 wire net407;
 wire net408;
 wire net409;
 wire net410;
 wire net411;
 wire net412;
 wire net413;
 wire clknet_leaf_1_clk;
 wire clknet_leaf_2_clk;
 wire clknet_leaf_3_clk;
 wire clknet_leaf_4_clk;
 wire clknet_leaf_5_clk;
 wire clknet_leaf_6_clk;
 wire clknet_leaf_7_clk;
 wire clknet_leaf_8_clk;
 wire clknet_leaf_9_clk;
 wire clknet_leaf_10_clk;
 wire clknet_leaf_11_clk;
 wire clknet_leaf_12_clk;
 wire clknet_leaf_13_clk;
 wire clknet_leaf_14_clk;
 wire clknet_leaf_15_clk;
 wire clknet_leaf_16_clk;
 wire clknet_leaf_17_clk;
 wire clknet_leaf_18_clk;
 wire clknet_leaf_19_clk;
 wire clknet_leaf_20_clk;
 wire clknet_leaf_21_clk;
 wire clknet_leaf_22_clk;
 wire clknet_leaf_23_clk;
 wire clknet_leaf_24_clk;
 wire clknet_leaf_25_clk;
 wire clknet_leaf_26_clk;
 wire clknet_leaf_27_clk;
 wire clknet_leaf_28_clk;
 wire clknet_leaf_29_clk;
 wire clknet_leaf_30_clk;
 wire clknet_leaf_31_clk;
 wire clknet_leaf_32_clk;
 wire clknet_leaf_33_clk;
 wire clknet_leaf_34_clk;
 wire clknet_leaf_35_clk;
 wire clknet_leaf_36_clk;
 wire clknet_0_clk;
 wire clknet_3_0__leaf_clk;
 wire clknet_3_1__leaf_clk;
 wire clknet_3_2__leaf_clk;
 wire clknet_3_3__leaf_clk;
 wire clknet_3_4__leaf_clk;
 wire clknet_3_5__leaf_clk;
 wire clknet_3_6__leaf_clk;
 wire clknet_3_7__leaf_clk;

 sg13g2_dfrbp_1 \B_reg[0]$_SDFF_PP0_  (.CLK(clknet_leaf_6_clk),
    .RESET_B(net184),
    .D(_0070_),
    .Q_N(_4116_),
    .Q(net23));
 sg13g2_dfrbp_1 \B_reg[1]$_SDFF_PP0_  (.CLK(clknet_leaf_11_clk),
    .RESET_B(net185),
    .D(_0071_),
    .Q_N(_4115_),
    .Q(net19));
 sg13g2_dfrbp_1 \G_reg[0]$_SDFF_PP0_  (.CLK(clknet_leaf_6_clk),
    .RESET_B(net186),
    .D(_0072_),
    .Q_N(_4114_),
    .Q(net22));
 sg13g2_dfrbp_1 \G_reg[1]$_SDFF_PP0_  (.CLK(clknet_leaf_11_clk),
    .RESET_B(net187),
    .D(_0073_),
    .Q_N(_4113_),
    .Q(net18));
 sg13g2_dfrbp_1 \R_reg[0]$_SDFF_PP0_  (.CLK(clknet_leaf_11_clk),
    .RESET_B(net188),
    .D(_0074_),
    .Q_N(_4112_),
    .Q(net21));
 sg13g2_dfrbp_1 \R_reg[1]$_SDFF_PP0_  (.CLK(clknet_leaf_11_clk),
    .RESET_B(net189),
    .D(_0075_),
    .Q_N(_4117_),
    .Q(net17));
 sg13g2_inv_1 _4123_ (.Y(_3478_),
    .A(handle_impact));
 sg13g2_nor2_1 _4124_ (.A(net7),
    .B(_3478_),
    .Y(_3479_));
 sg13g2_buf_2 _4125_ (.A(_3479_),
    .X(_3480_));
 sg13g2_buf_1 _4126_ (.A(rst_n),
    .X(_3481_));
 sg13g2_buf_1 _4127_ (.A(_3481_),
    .X(_3482_));
 sg13g2_buf_1 _4128_ (.A(net183),
    .X(_3483_));
 sg13g2_buf_1 _4129_ (.A(\color_entropy[1] ),
    .X(_3484_));
 sg13g2_buf_2 _4130_ (.A(\i_colors.channel[2] ),
    .X(_3485_));
 sg13g2_nand4_1 _4131_ (.B(net169),
    .C(_3484_),
    .A(_3480_),
    .Y(_3486_),
    .D(_3485_));
 sg13g2_inv_1 _4132_ (.Y(_3487_),
    .A(_3484_));
 sg13g2_buf_1 _4133_ (.A(\i_colors.channel[1] ),
    .X(_3488_));
 sg13g2_nand4_1 _4134_ (.B(net183),
    .C(_3487_),
    .A(_3480_),
    .Y(_3489_),
    .D(_3488_));
 sg13g2_inv_1 _4135_ (.Y(_3490_),
    .A(_3480_));
 sg13g2_buf_1 _4136_ (.A(\i_colors.channel[0] ),
    .X(_3491_));
 sg13g2_inv_2 _4137_ (.Y(_3492_),
    .A(_3481_));
 sg13g2_buf_1 _4138_ (.A(_3492_),
    .X(_3493_));
 sg13g2_a21oi_1 _4139_ (.A1(_3490_),
    .A2(_3491_),
    .Y(_3494_),
    .B1(_3493_));
 sg13g2_nand3_1 _4140_ (.B(_3489_),
    .C(_3494_),
    .A(_3486_),
    .Y(_0001_));
 sg13g2_nand4_1 _4141_ (.B(net183),
    .C(_3491_),
    .A(_3480_),
    .Y(_3495_),
    .D(_3484_));
 sg13g2_nand4_1 _4142_ (.B(net183),
    .C(_3487_),
    .A(_3480_),
    .Y(_3496_),
    .D(_3485_));
 sg13g2_nand3_1 _4143_ (.B(net169),
    .C(_3488_),
    .A(_3490_),
    .Y(_3497_));
 sg13g2_nand3_1 _4144_ (.B(_3496_),
    .C(_3497_),
    .A(_3495_),
    .Y(_0002_));
 sg13g2_nand4_1 _4145_ (.B(_3482_),
    .C(_3484_),
    .A(_3480_),
    .Y(_3498_),
    .D(_3488_));
 sg13g2_nand4_1 _4146_ (.B(_3482_),
    .C(_3491_),
    .A(_3480_),
    .Y(_3499_),
    .D(_3487_));
 sg13g2_nand3_1 _4147_ (.B(net169),
    .C(_3485_),
    .A(_3490_),
    .Y(_3500_));
 sg13g2_nand3_1 _4148_ (.B(_3499_),
    .C(_3500_),
    .A(_3498_),
    .Y(_0003_));
 sg13g2_buf_2 _4149_ (.A(\i_orchestrator.vga_y[5] ),
    .X(_3501_));
 sg13g2_inv_1 _4150_ (.Y(_3502_),
    .A(_3501_));
 sg13g2_buf_2 _4151_ (.A(\i_orchestrator.vga_y[8] ),
    .X(_3503_));
 sg13g2_inv_2 _4152_ (.Y(_3504_),
    .A(_3503_));
 sg13g2_buf_2 _4153_ (.A(\i_orchestrator.vga_y[7] ),
    .X(_3505_));
 sg13g2_buf_2 _4154_ (.A(\i_orchestrator.vga_y[6] ),
    .X(_3506_));
 sg13g2_nand2_1 _4155_ (.Y(_3507_),
    .A(_3505_),
    .B(_3506_));
 sg13g2_nor3_1 _4156_ (.A(_3502_),
    .B(_3504_),
    .C(_3507_),
    .Y(_3508_));
 sg13g2_buf_2 _4157_ (.A(\i_orchestrator.vga_y[1] ),
    .X(_3509_));
 sg13g2_buf_2 _4158_ (.A(\i_orchestrator.vga_y[0] ),
    .X(_3510_));
 sg13g2_nand2_1 _4159_ (.Y(_3511_),
    .A(_3509_),
    .B(_3510_));
 sg13g2_buf_1 _4160_ (.A(\i_orchestrator.vga_y[2] ),
    .X(_3512_));
 sg13g2_inv_1 _4161_ (.Y(_3513_),
    .A(_3512_));
 sg13g2_buf_1 _4162_ (.A(\i_orchestrator.vga_y[3] ),
    .X(_3514_));
 sg13g2_inv_1 _4163_ (.Y(_3515_),
    .A(net182));
 sg13g2_a21oi_1 _4164_ (.A1(_3511_),
    .A2(_3513_),
    .Y(_3516_),
    .B1(_3515_));
 sg13g2_inv_1 _4165_ (.Y(_3517_),
    .A(_3509_));
 sg13g2_nor2_1 _4166_ (.A(_3510_),
    .B(_3517_),
    .Y(_3518_));
 sg13g2_nand3_1 _4167_ (.B(_3513_),
    .C(net182),
    .A(_3518_),
    .Y(_3519_));
 sg13g2_inv_1 _4168_ (.Y(_3520_),
    .A(_3519_));
 sg13g2_buf_2 _4169_ (.A(\i_orchestrator.vga_y[9] ),
    .X(_3521_));
 sg13g2_nor2_1 _4170_ (.A(_3521_),
    .B(_3504_),
    .Y(_3522_));
 sg13g2_inv_1 _4171_ (.Y(_3523_),
    .A(_3522_));
 sg13g2_inv_1 _4172_ (.Y(_3524_),
    .A(_3507_));
 sg13g2_buf_1 _4173_ (.A(\i_orchestrator.vga_y[4] ),
    .X(_3525_));
 sg13g2_inv_1 _4174_ (.Y(_3526_),
    .A(_3525_));
 sg13g2_nand3_1 _4175_ (.B(_3526_),
    .C(_3501_),
    .A(_3524_),
    .Y(_3527_));
 sg13g2_nor2_1 _4176_ (.A(_3523_),
    .B(_3527_),
    .Y(_3528_));
 sg13g2_a22oi_1 _4177_ (.Y(_3529_),
    .B1(_3520_),
    .B2(_3528_),
    .A2(_3516_),
    .A1(_3508_));
 sg13g2_nand2_1 _4178_ (.Y(_3530_),
    .A(_3512_),
    .B(net182));
 sg13g2_a21oi_1 _4179_ (.A1(_3530_),
    .A2(_3526_),
    .Y(_3531_),
    .B1(_3502_));
 sg13g2_nor2_1 _4180_ (.A(_3504_),
    .B(_3507_),
    .Y(_3532_));
 sg13g2_a21oi_1 _4181_ (.A1(_3531_),
    .A2(_3532_),
    .Y(_3533_),
    .B1(_3521_));
 sg13g2_nor2b_1 _4182_ (.A(_3529_),
    .B_N(_3533_),
    .Y(_0007_));
 sg13g2_buf_2 _4183_ (.A(\i_orchestrator.vga_x[8] ),
    .X(_3534_));
 sg13g2_nand2_1 _4184_ (.Y(_3535_),
    .A(\i_orchestrator.vga_x[9] ),
    .B(_3534_));
 sg13g2_buf_1 _4185_ (.A(\i_orchestrator.vga_x[6] ),
    .X(_3536_));
 sg13g2_inv_1 _4186_ (.Y(_3537_),
    .A(_3536_));
 sg13g2_buf_2 _4187_ (.A(\i_orchestrator.vga_x[5] ),
    .X(_3538_));
 sg13g2_inv_1 _4188_ (.Y(_3539_),
    .A(_3538_));
 sg13g2_buf_2 _4189_ (.A(\i_orchestrator.vga_x[4] ),
    .X(_3540_));
 sg13g2_inv_1 _4190_ (.Y(_3541_),
    .A(_3540_));
 sg13g2_nand3_1 _4191_ (.B(_3539_),
    .C(_3541_),
    .A(_3537_),
    .Y(_3542_));
 sg13g2_inv_1 _4192_ (.Y(_3543_),
    .A(\i_orchestrator.vga_x[9] ));
 sg13g2_nor2_1 _4193_ (.A(_3534_),
    .B(\i_orchestrator.vga_x[7] ),
    .Y(_3544_));
 sg13g2_nor2_1 _4194_ (.A(_3543_),
    .B(_3544_),
    .Y(_3545_));
 sg13g2_nand3_1 _4195_ (.B(_3538_),
    .C(_3540_),
    .A(_3536_),
    .Y(_3546_));
 sg13g2_and4_1 _4196_ (.A(_3535_),
    .B(_3542_),
    .C(_3545_),
    .D(_3546_),
    .X(_0006_));
 sg13g2_a21oi_2 _4197_ (.B1(_3521_),
    .Y(_3547_),
    .A2(_3501_),
    .A1(_3532_));
 sg13g2_buf_1 _4198_ (.A(_3547_),
    .X(_3548_));
 sg13g2_a21o_1 _4199_ (.A2(net182),
    .A1(net127),
    .B1(_0058_),
    .X(_3549_));
 sg13g2_inv_4 _4200_ (.A(_3547_),
    .Y(_3550_));
 sg13g2_o21ai_1 _4201_ (.B1(\i_transform.track_y[2] ),
    .Y(_3551_),
    .A1(_3513_),
    .A2(_3550_));
 sg13g2_nand3_1 _4202_ (.B(net182),
    .C(_0058_),
    .A(net127),
    .Y(_3552_));
 sg13g2_inv_1 _4203_ (.Y(_3553_),
    .A(\i_transform.track_y[2] ));
 sg13g2_nand3_1 _4204_ (.B(_3512_),
    .C(_3553_),
    .A(net127),
    .Y(_3554_));
 sg13g2_nand4_1 _4205_ (.B(_3551_),
    .C(_3552_),
    .A(_3549_),
    .Y(_3555_),
    .D(_3554_));
 sg13g2_buf_2 _4206_ (.A(\i_transform.track_y[8] ),
    .X(_3556_));
 sg13g2_inv_1 _4207_ (.Y(_3557_),
    .A(_3556_));
 sg13g2_a21oi_1 _4208_ (.A1(net127),
    .A2(_3503_),
    .Y(_3558_),
    .B1(_3557_));
 sg13g2_nor3_1 _4209_ (.A(_3504_),
    .B(_3556_),
    .C(_3550_),
    .Y(_3559_));
 sg13g2_nor3_1 _4210_ (.A(\i_transform.track_y[9] ),
    .B(_3558_),
    .C(_3559_),
    .Y(_3560_));
 sg13g2_inv_1 _4211_ (.Y(_3561_),
    .A(_3560_));
 sg13g2_nand2_1 _4212_ (.Y(_3562_),
    .A(_3547_),
    .B(_3505_));
 sg13g2_xnor2_1 _4213_ (.Y(_3563_),
    .A(_0059_),
    .B(_3562_));
 sg13g2_inv_1 _4214_ (.Y(_3564_),
    .A(_3506_));
 sg13g2_buf_1 _4215_ (.A(\i_transform.track_y[6] ),
    .X(_3565_));
 sg13g2_o21ai_1 _4216_ (.B1(_3565_),
    .Y(_3566_),
    .A1(_3564_),
    .A2(_3550_));
 sg13g2_inv_1 _4217_ (.Y(_3567_),
    .A(_3565_));
 sg13g2_nand3_1 _4218_ (.B(_3506_),
    .C(_3567_),
    .A(_3548_),
    .Y(_3568_));
 sg13g2_nand3_1 _4219_ (.B(_3566_),
    .C(_3568_),
    .A(_3563_),
    .Y(_3569_));
 sg13g2_nor2_1 _4220_ (.A(_3561_),
    .B(_3569_),
    .Y(_3570_));
 sg13g2_inv_1 _4221_ (.Y(_3571_),
    .A(\i_transform.track_y[4] ));
 sg13g2_a21oi_1 _4222_ (.A1(net127),
    .A2(_3525_),
    .Y(_3572_),
    .B1(_3571_));
 sg13g2_inv_1 _4223_ (.Y(_3573_),
    .A(_0060_));
 sg13g2_nand2_1 _4224_ (.Y(_3574_),
    .A(net127),
    .B(_3501_));
 sg13g2_nor2_1 _4225_ (.A(_3573_),
    .B(_3574_),
    .Y(_3575_));
 sg13g2_nor3_1 _4226_ (.A(_3526_),
    .B(\i_transform.track_y[4] ),
    .C(_3550_),
    .Y(_3576_));
 sg13g2_nand2_1 _4227_ (.Y(_3577_),
    .A(_3574_),
    .B(_3573_));
 sg13g2_inv_1 _4228_ (.Y(_3578_),
    .A(_3577_));
 sg13g2_nor4_1 _4229_ (.A(_3572_),
    .B(_3575_),
    .C(_3576_),
    .D(_3578_),
    .Y(_3579_));
 sg13g2_nand3b_1 _4230_ (.B(_3570_),
    .C(_3579_),
    .Y(_3580_),
    .A_N(_3555_));
 sg13g2_buf_1 _4231_ (.A(\i_transform.track_y[1] ),
    .X(_3581_));
 sg13g2_nor3_1 _4232_ (.A(_3517_),
    .B(_3581_),
    .C(_3550_),
    .Y(_3582_));
 sg13g2_buf_1 _4233_ (.A(\i_transform.track_y[0] ),
    .X(_3583_));
 sg13g2_nand2_1 _4234_ (.Y(_3584_),
    .A(net127),
    .B(_3510_));
 sg13g2_nor2_1 _4235_ (.A(_3583_),
    .B(_3584_),
    .Y(_3585_));
 sg13g2_nand2_1 _4236_ (.Y(_3586_),
    .A(_3548_),
    .B(_3509_));
 sg13g2_a22oi_1 _4237_ (.Y(_3587_),
    .B1(_3583_),
    .B2(_3584_),
    .A2(_3581_),
    .A1(_3586_));
 sg13g2_inv_1 _4238_ (.Y(_3588_),
    .A(_3587_));
 sg13g2_nor3_1 _4239_ (.A(_3582_),
    .B(_3585_),
    .C(_3588_),
    .Y(_3589_));
 sg13g2_nor2b_1 _4240_ (.A(_3580_),
    .B_N(_3589_),
    .Y(_3590_));
 sg13g2_buf_2 _4241_ (.A(_3590_),
    .X(_3591_));
 sg13g2_inv_2 _4242_ (.Y(_3592_),
    .A(_3591_));
 sg13g2_nor2_1 _4243_ (.A(_3545_),
    .B(_3550_),
    .Y(_3593_));
 sg13g2_inv_2 _4244_ (.Y(_3594_),
    .A(_3593_));
 sg13g2_nor3_1 _4245_ (.A(_3541_),
    .B(\i_transform.track_x[4] ),
    .C(_3594_),
    .Y(_3595_));
 sg13g2_buf_1 _4246_ (.A(_3593_),
    .X(_3596_));
 sg13g2_inv_1 _4247_ (.Y(_3597_),
    .A(\i_transform.track_x[4] ));
 sg13g2_a21oi_1 _4248_ (.A1(_3596_),
    .A2(_3540_),
    .Y(_3598_),
    .B1(_3597_));
 sg13g2_buf_1 _4249_ (.A(\i_transform.track_x[5] ),
    .X(_3599_));
 sg13g2_nand2_1 _4250_ (.Y(_3600_),
    .A(_3593_),
    .B(_3538_));
 sg13g2_nor2_1 _4251_ (.A(_3599_),
    .B(_3600_),
    .Y(_3601_));
 sg13g2_nand2_1 _4252_ (.Y(_3602_),
    .A(_3600_),
    .B(_3599_));
 sg13g2_nand2b_1 _4253_ (.Y(_3603_),
    .B(_3602_),
    .A_N(_3601_));
 sg13g2_nor3_1 _4254_ (.A(_3595_),
    .B(_3598_),
    .C(_3603_),
    .Y(_3604_));
 sg13g2_inv_1 _4255_ (.Y(_3605_),
    .A(\i_orchestrator.vga_x[2] ));
 sg13g2_nor3_1 _4256_ (.A(_3605_),
    .B(\i_transform.track_x[2] ),
    .C(net103),
    .Y(_3606_));
 sg13g2_inv_1 _4257_ (.Y(_3607_),
    .A(_3606_));
 sg13g2_buf_2 _4258_ (.A(\i_orchestrator.vga_x[3] ),
    .X(_3608_));
 sg13g2_inv_1 _4259_ (.Y(_3609_),
    .A(\i_transform.track_x[3] ));
 sg13g2_a21oi_1 _4260_ (.A1(net102),
    .A2(_3608_),
    .Y(_3610_),
    .B1(_3609_));
 sg13g2_nand3_1 _4261_ (.B(_3608_),
    .C(_3609_),
    .A(net102),
    .Y(_3611_));
 sg13g2_nor2b_1 _4262_ (.A(_3610_),
    .B_N(_3611_),
    .Y(_3612_));
 sg13g2_o21ai_1 _4263_ (.B1(\i_transform.track_x[2] ),
    .Y(_3613_),
    .A1(_3605_),
    .A2(net103));
 sg13g2_nand4_1 _4264_ (.B(_3607_),
    .C(_3612_),
    .A(_3604_),
    .Y(_3614_),
    .D(_3613_));
 sg13g2_buf_1 _4265_ (.A(\i_transform.track_x[8] ),
    .X(_3615_));
 sg13g2_inv_1 _4266_ (.Y(_3616_),
    .A(_3615_));
 sg13g2_a21oi_1 _4267_ (.A1(net102),
    .A2(_3534_),
    .Y(_3617_),
    .B1(_3616_));
 sg13g2_and3_1 _4268_ (.X(_3618_),
    .A(_3593_),
    .B(_3534_),
    .C(_3616_));
 sg13g2_buf_1 _4269_ (.A(\i_transform.track_x[9] ),
    .X(_3619_));
 sg13g2_nor2_1 _4270_ (.A(_3543_),
    .B(net103),
    .Y(_3620_));
 sg13g2_inv_1 _4271_ (.Y(_3621_),
    .A(_3620_));
 sg13g2_nor2_1 _4272_ (.A(_3619_),
    .B(_3621_),
    .Y(_3622_));
 sg13g2_nand2_1 _4273_ (.Y(_3623_),
    .A(_3621_),
    .B(_3619_));
 sg13g2_inv_1 _4274_ (.Y(_3624_),
    .A(_3623_));
 sg13g2_nor4_1 _4275_ (.A(_3617_),
    .B(_3618_),
    .C(_3622_),
    .D(_3624_),
    .Y(_3625_));
 sg13g2_buf_1 _4276_ (.A(\i_transform.track_x[7] ),
    .X(_3626_));
 sg13g2_nand2_1 _4277_ (.Y(_3627_),
    .A(net102),
    .B(\i_orchestrator.vga_x[7] ));
 sg13g2_nor2_1 _4278_ (.A(_3626_),
    .B(_3627_),
    .Y(_3628_));
 sg13g2_inv_1 _4279_ (.Y(_3629_),
    .A(_3628_));
 sg13g2_nand2_1 _4280_ (.Y(_3630_),
    .A(_3627_),
    .B(_3626_));
 sg13g2_buf_2 _4281_ (.A(\i_transform.track_x[6] ),
    .X(_3631_));
 sg13g2_inv_1 _4282_ (.Y(_3632_),
    .A(_3631_));
 sg13g2_a21oi_1 _4283_ (.A1(net102),
    .A2(_3536_),
    .Y(_3633_),
    .B1(_3632_));
 sg13g2_nor3_1 _4284_ (.A(_3537_),
    .B(_3631_),
    .C(net103),
    .Y(_3634_));
 sg13g2_nor2_1 _4285_ (.A(_3633_),
    .B(_3634_),
    .Y(_3635_));
 sg13g2_nand4_1 _4286_ (.B(_3629_),
    .C(_3630_),
    .A(_3625_),
    .Y(_3636_),
    .D(_3635_));
 sg13g2_nor2_1 _4287_ (.A(_3614_),
    .B(_3636_),
    .Y(_3637_));
 sg13g2_buf_1 _4288_ (.A(\i_transform.track_x[1] ),
    .X(_3638_));
 sg13g2_inv_1 _4289_ (.Y(_3639_),
    .A(_3638_));
 sg13g2_a21oi_1 _4290_ (.A1(net102),
    .A2(\i_orchestrator.vga_x[1] ),
    .Y(_3640_),
    .B1(_3639_));
 sg13g2_buf_1 _4291_ (.A(\i_transform.track_x[0] ),
    .X(_3641_));
 sg13g2_inv_1 _4292_ (.Y(_3642_),
    .A(_3641_));
 sg13g2_a21oi_1 _4293_ (.A1(net102),
    .A2(\i_orchestrator.vga_x[0] ),
    .Y(_3643_),
    .B1(_3642_));
 sg13g2_inv_1 _4294_ (.Y(_3644_),
    .A(\i_orchestrator.vga_x[1] ));
 sg13g2_nor3_1 _4295_ (.A(_3644_),
    .B(_3638_),
    .C(net103),
    .Y(_3645_));
 sg13g2_nor3_1 _4296_ (.A(_3640_),
    .B(_3643_),
    .C(_3645_),
    .Y(_3646_));
 sg13g2_nand3_1 _4297_ (.B(\i_orchestrator.vga_x[0] ),
    .C(_3642_),
    .A(net102),
    .Y(_3647_));
 sg13g2_and2_1 _4298_ (.A(_3646_),
    .B(_3647_),
    .X(_3648_));
 sg13g2_nand2_1 _4299_ (.Y(_3649_),
    .A(_3637_),
    .B(_3648_));
 sg13g2_inv_1 _4300_ (.Y(_3650_),
    .A(_3649_));
 sg13g2_nor2_1 _4301_ (.A(net84),
    .B(_3650_),
    .Y(_3651_));
 sg13g2_buf_2 _4302_ (.A(_3651_),
    .X(_3652_));
 sg13g2_inv_4 _4303_ (.A(_3652_),
    .Y(_3653_));
 sg13g2_o21ai_1 _4304_ (.B1(_3637_),
    .Y(_3654_),
    .A1(_3645_),
    .A2(_3646_));
 sg13g2_o21ai_1 _4305_ (.B1(_3630_),
    .Y(_3655_),
    .A1(_3628_),
    .A2(_3634_));
 sg13g2_nand2b_1 _4306_ (.Y(_3656_),
    .B(_3625_),
    .A_N(_3655_));
 sg13g2_nor2_1 _4307_ (.A(_3631_),
    .B(_3599_),
    .Y(_3657_));
 sg13g2_inv_1 _4308_ (.Y(_3658_),
    .A(_3626_));
 sg13g2_nand2_1 _4309_ (.Y(_3659_),
    .A(_3657_),
    .B(_3658_));
 sg13g2_nor2_1 _4310_ (.A(_3615_),
    .B(_3659_),
    .Y(_3660_));
 sg13g2_nand2b_1 _4311_ (.Y(_3661_),
    .B(_3660_),
    .A_N(_3619_));
 sg13g2_o21ai_1 _4312_ (.B1(_3623_),
    .Y(_3662_),
    .A1(_3618_),
    .A2(_3622_));
 sg13g2_nand4_1 _4313_ (.B(_3656_),
    .C(_3661_),
    .A(_3654_),
    .Y(_3663_),
    .D(_3662_));
 sg13g2_a21oi_1 _4314_ (.A1(_3607_),
    .A2(_3611_),
    .Y(_3664_),
    .B1(_3610_));
 sg13g2_nand2_1 _4315_ (.Y(_3665_),
    .A(_3604_),
    .B(_3664_));
 sg13g2_a21oi_1 _4316_ (.A1(_3595_),
    .A2(_3602_),
    .Y(_3666_),
    .B1(_3601_));
 sg13g2_a21o_1 _4317_ (.A2(_3666_),
    .A1(_3665_),
    .B1(_3636_),
    .X(_3667_));
 sg13g2_nor2b_1 _4318_ (.A(_3663_),
    .B_N(_3667_),
    .Y(_3668_));
 sg13g2_buf_1 _4319_ (.A(_3668_),
    .X(_3669_));
 sg13g2_nor2_1 _4320_ (.A(net63),
    .B(_3669_),
    .Y(_3670_));
 sg13g2_buf_2 _4321_ (.A(_3670_),
    .X(_3671_));
 sg13g2_inv_1 _4322_ (.Y(_3672_),
    .A(_0027_));
 sg13g2_buf_8 _4323_ (.A(\i_collision.i_coll_table.in[1] ),
    .X(_3673_));
 sg13g2_buf_8 _4324_ (.A(\i_kinematics.phi[3] ),
    .X(_3674_));
 sg13g2_xor2_1 _4325_ (.B(_3674_),
    .A(net181),
    .X(_3675_));
 sg13g2_buf_8 _4326_ (.A(\i_kinematics.phi[4] ),
    .X(_3676_));
 sg13g2_xor2_1 _4327_ (.B(_3676_),
    .A(net181),
    .X(_3677_));
 sg13g2_buf_2 _4328_ (.A(_3677_),
    .X(_3678_));
 sg13g2_nand2_1 _4329_ (.Y(_3679_),
    .A(_3675_),
    .B(_3678_));
 sg13g2_xnor2_1 _4330_ (.Y(_3680_),
    .A(net181),
    .B(_3674_));
 sg13g2_xnor2_1 _4331_ (.Y(_3681_),
    .A(net181),
    .B(_3676_));
 sg13g2_nand2_2 _4332_ (.Y(_3682_),
    .A(_3680_),
    .B(_3681_));
 sg13g2_buf_2 _4333_ (.A(\i_kinematics.phi[5] ),
    .X(_3683_));
 sg13g2_xnor2_1 _4334_ (.Y(_3684_),
    .A(net181),
    .B(_3683_));
 sg13g2_buf_8 _4335_ (.A(_3684_),
    .X(_3685_));
 sg13g2_inv_2 _4336_ (.Y(_3686_),
    .A(net149));
 sg13g2_nand3_1 _4337_ (.B(_3682_),
    .C(_3686_),
    .A(_3679_),
    .Y(_3687_));
 sg13g2_xnor2_1 _4338_ (.Y(_3688_),
    .A(_3673_),
    .B(\i_kinematics.phi[6] ));
 sg13g2_buf_2 _4339_ (.A(_3688_),
    .X(_3689_));
 sg13g2_buf_1 _4340_ (.A(_3689_),
    .X(_3690_));
 sg13g2_nand2_1 _4341_ (.Y(_3691_),
    .A(_3681_),
    .B(net149));
 sg13g2_nand3_1 _4342_ (.B(_3690_),
    .C(_3691_),
    .A(_3687_),
    .Y(_3692_));
 sg13g2_a21oi_1 _4343_ (.A1(_3675_),
    .A2(net149),
    .Y(_3693_),
    .B1(net134));
 sg13g2_nand2_1 _4344_ (.Y(_3694_),
    .A(_3678_),
    .B(_3680_));
 sg13g2_buf_2 _4345_ (.A(\i_kinematics.phi[7] ),
    .X(_3695_));
 sg13g2_xnor2_1 _4346_ (.Y(_3696_),
    .A(net181),
    .B(_3695_));
 sg13g2_buf_1 _4347_ (.A(_3696_),
    .X(_3697_));
 sg13g2_a21oi_1 _4348_ (.A1(_3693_),
    .A2(_3694_),
    .Y(_3698_),
    .B1(net148));
 sg13g2_nand2_1 _4349_ (.Y(_3699_),
    .A(_3692_),
    .B(_3698_));
 sg13g2_buf_2 _4350_ (.A(\i_collision.phi[1] ),
    .X(_3700_));
 sg13g2_nor2_1 _4351_ (.A(net181),
    .B(_3700_),
    .Y(_3701_));
 sg13g2_nand2_1 _4352_ (.Y(_3702_),
    .A(_3673_),
    .B(_3700_));
 sg13g2_inv_1 _4353_ (.Y(_3703_),
    .A(_3702_));
 sg13g2_nor2_1 _4354_ (.A(_3701_),
    .B(_3703_),
    .Y(_3704_));
 sg13g2_buf_2 _4355_ (.A(_3704_),
    .X(_3705_));
 sg13g2_a21oi_1 _4356_ (.A1(_3681_),
    .A2(net149),
    .Y(_3706_),
    .B1(_3689_));
 sg13g2_nor2_1 _4357_ (.A(_3681_),
    .B(net149),
    .Y(_3707_));
 sg13g2_nand2_1 _4358_ (.Y(_3708_),
    .A(_3707_),
    .B(_3675_));
 sg13g2_inv_2 _4359_ (.Y(_3709_),
    .A(net148));
 sg13g2_a21oi_1 _4360_ (.A1(_3706_),
    .A2(_3708_),
    .Y(_3710_),
    .B1(_3709_));
 sg13g2_inv_1 _4361_ (.Y(_3711_),
    .A(_3710_));
 sg13g2_nand3_1 _4362_ (.B(_3705_),
    .C(_3711_),
    .A(_3699_),
    .Y(_3712_));
 sg13g2_a21oi_1 _4363_ (.A1(_3678_),
    .A2(_3680_),
    .Y(_3713_),
    .B1(net134));
 sg13g2_nor2_1 _4364_ (.A(_3680_),
    .B(_3678_),
    .Y(_3714_));
 sg13g2_nand2_1 _4365_ (.Y(_3715_),
    .A(_3714_),
    .B(_3686_));
 sg13g2_a21oi_1 _4366_ (.A1(_3713_),
    .A2(_3715_),
    .Y(_3716_),
    .B1(net148));
 sg13g2_inv_1 _4367_ (.Y(_3717_),
    .A(_3689_));
 sg13g2_nand2_1 _4368_ (.Y(_3718_),
    .A(_3675_),
    .B(net149));
 sg13g2_nor2_1 _4369_ (.A(_3678_),
    .B(_3718_),
    .Y(_3719_));
 sg13g2_nor2_1 _4370_ (.A(_3717_),
    .B(_3719_),
    .Y(_3720_));
 sg13g2_nand2_1 _4371_ (.Y(_3721_),
    .A(_3679_),
    .B(_3682_));
 sg13g2_nand2_1 _4372_ (.Y(_3722_),
    .A(_3721_),
    .B(_3686_));
 sg13g2_nand2_1 _4373_ (.Y(_3723_),
    .A(_3720_),
    .B(_3722_));
 sg13g2_nand2_1 _4374_ (.Y(_3724_),
    .A(_3716_),
    .B(_3723_));
 sg13g2_inv_2 _4375_ (.Y(_3725_),
    .A(_3705_));
 sg13g2_nor2_1 _4376_ (.A(net149),
    .B(_3675_),
    .Y(_3726_));
 sg13g2_a21oi_1 _4377_ (.A1(_3678_),
    .A2(net134),
    .Y(_3727_),
    .B1(_3718_));
 sg13g2_o21ai_1 _4378_ (.B1(net148),
    .Y(_3728_),
    .A1(_3726_),
    .A2(_3727_));
 sg13g2_nand3_1 _4379_ (.B(_3725_),
    .C(_3728_),
    .A(_3724_),
    .Y(_3729_));
 sg13g2_nand2_1 _4380_ (.Y(_3730_),
    .A(_3712_),
    .B(_3729_));
 sg13g2_a21oi_1 _4381_ (.A1(_3708_),
    .A2(net134),
    .Y(_3731_),
    .B1(_3709_));
 sg13g2_nand2_1 _4382_ (.Y(_3732_),
    .A(_3687_),
    .B(_3706_));
 sg13g2_nand2_1 _4383_ (.Y(_3733_),
    .A(_3731_),
    .B(_3732_));
 sg13g2_nand2_1 _4384_ (.Y(_3734_),
    .A(_3726_),
    .B(_3690_));
 sg13g2_nand2_1 _4385_ (.Y(_3735_),
    .A(_3714_),
    .B(_3717_));
 sg13g2_nand2_1 _4386_ (.Y(_3736_),
    .A(_3694_),
    .B(net149));
 sg13g2_nand3_1 _4387_ (.B(_3735_),
    .C(_3736_),
    .A(_3734_),
    .Y(_3737_));
 sg13g2_nor2_1 _4388_ (.A(_3689_),
    .B(_3686_),
    .Y(_3738_));
 sg13g2_a21oi_1 _4389_ (.A1(_3738_),
    .A2(_3714_),
    .Y(_3739_),
    .B1(net148));
 sg13g2_nand2_1 _4390_ (.Y(_3740_),
    .A(_3737_),
    .B(_3739_));
 sg13g2_buf_1 _4391_ (.A(_3705_),
    .X(_3741_));
 sg13g2_nand3_1 _4392_ (.B(_3740_),
    .C(net116),
    .A(_3733_),
    .Y(_3742_));
 sg13g2_nand2_1 _4393_ (.Y(_3743_),
    .A(_3685_),
    .B(_3689_));
 sg13g2_nor2_1 _4394_ (.A(_3681_),
    .B(_3709_),
    .Y(_3744_));
 sg13g2_nor2_1 _4395_ (.A(_3743_),
    .B(_3721_),
    .Y(_3745_));
 sg13g2_a21oi_1 _4396_ (.A1(_3743_),
    .A2(_3744_),
    .Y(_3746_),
    .B1(_3745_));
 sg13g2_nand2_1 _4397_ (.Y(_3747_),
    .A(_3714_),
    .B(_3689_));
 sg13g2_o21ai_1 _4398_ (.B1(_3747_),
    .Y(_3748_),
    .A1(net134),
    .A2(_3726_));
 sg13g2_nor2_1 _4399_ (.A(net148),
    .B(_3719_),
    .Y(_3749_));
 sg13g2_nand2_1 _4400_ (.Y(_3750_),
    .A(_3748_),
    .B(_3749_));
 sg13g2_buf_1 _4401_ (.A(_3725_),
    .X(_3751_));
 sg13g2_nand3_1 _4402_ (.B(_3750_),
    .C(_3751_),
    .A(_3746_),
    .Y(_3752_));
 sg13g2_nand2_2 _4403_ (.Y(_3753_),
    .A(_3742_),
    .B(_3752_));
 sg13g2_buf_1 _4404_ (.A(\i_kinematics.phi[10] ),
    .X(_3754_));
 sg13g2_inv_1 _4405_ (.Y(_3755_),
    .A(orient));
 sg13g2_nand2b_1 _4406_ (.Y(_3756_),
    .B(_3755_),
    .A_N(_3754_));
 sg13g2_nand2_1 _4407_ (.Y(_3757_),
    .A(orient),
    .B(_3754_));
 sg13g2_nand2_1 _4408_ (.Y(_3758_),
    .A(_3756_),
    .B(_3757_));
 sg13g2_inv_1 _4409_ (.Y(_3759_),
    .A(_3758_));
 sg13g2_buf_1 _4410_ (.A(_3759_),
    .X(_3760_));
 sg13g2_nand2_1 _4411_ (.Y(_3761_),
    .A(_3753_),
    .B(net126));
 sg13g2_xnor2_1 _4412_ (.Y(_3762_),
    .A(_3730_),
    .B(_3761_));
 sg13g2_buf_2 _4413_ (.A(_3762_),
    .X(_3763_));
 sg13g2_buf_1 _4414_ (.A(_0028_),
    .X(_3764_));
 sg13g2_inv_1 _4415_ (.Y(_3765_),
    .A(_3764_));
 sg13g2_nand2_1 _4416_ (.Y(_3766_),
    .A(_3733_),
    .B(_3740_));
 sg13g2_nand2_1 _4417_ (.Y(_3767_),
    .A(_3766_),
    .B(_3705_));
 sg13g2_nand2_1 _4418_ (.Y(_3768_),
    .A(_3746_),
    .B(_3750_));
 sg13g2_nand2_1 _4419_ (.Y(_3769_),
    .A(_3768_),
    .B(_3725_));
 sg13g2_nand2_1 _4420_ (.Y(_3770_),
    .A(_3767_),
    .B(_3769_));
 sg13g2_buf_2 _4421_ (.A(_3770_),
    .X(_3771_));
 sg13g2_nor2_1 _4422_ (.A(_3765_),
    .B(_3771_),
    .Y(_3772_));
 sg13g2_buf_2 _4423_ (.A(\i_capsule.tf_y[0] ),
    .X(_3773_));
 sg13g2_xnor2_1 _4424_ (.Y(_3774_),
    .A(_3773_),
    .B(_3763_));
 sg13g2_nor2_1 _4425_ (.A(_3772_),
    .B(_3774_),
    .Y(_3775_));
 sg13g2_a21oi_1 _4426_ (.A1(_3672_),
    .A2(_3763_),
    .Y(_3776_),
    .B1(_3775_));
 sg13g2_buf_2 _4427_ (.A(_0026_),
    .X(_3777_));
 sg13g2_nand2_1 _4428_ (.Y(_3778_),
    .A(_3678_),
    .B(_3685_));
 sg13g2_nand3_1 _4429_ (.B(_3717_),
    .C(_3778_),
    .A(_3722_),
    .Y(_3779_));
 sg13g2_nand3_1 _4430_ (.B(_3692_),
    .C(_3697_),
    .A(_3779_),
    .Y(_3780_));
 sg13g2_nand2_1 _4431_ (.Y(_3781_),
    .A(_3682_),
    .B(_3686_));
 sg13g2_nand3_1 _4432_ (.B(net134),
    .C(_3691_),
    .A(_3781_),
    .Y(_3782_));
 sg13g2_a21oi_1 _4433_ (.A1(_3738_),
    .A2(_3679_),
    .Y(_3783_),
    .B1(net148));
 sg13g2_nand2_1 _4434_ (.Y(_3784_),
    .A(_3707_),
    .B(_3717_));
 sg13g2_inv_1 _4435_ (.Y(_3785_),
    .A(_3784_));
 sg13g2_nand2_1 _4436_ (.Y(_3786_),
    .A(_3785_),
    .B(_3675_));
 sg13g2_nand3_1 _4437_ (.B(_3783_),
    .C(_3786_),
    .A(_3782_),
    .Y(_3787_));
 sg13g2_a21oi_1 _4438_ (.A1(_3780_),
    .A2(_3787_),
    .Y(_3788_),
    .B1(net116));
 sg13g2_o21ai_1 _4439_ (.B1(_3717_),
    .Y(_3789_),
    .A1(_3686_),
    .A2(_3682_));
 sg13g2_nand2_1 _4440_ (.Y(_3790_),
    .A(_3781_),
    .B(net134));
 sg13g2_nand2_2 _4441_ (.Y(_3791_),
    .A(_3790_),
    .B(_3709_));
 sg13g2_inv_1 _4442_ (.Y(_3792_),
    .A(_3791_));
 sg13g2_o21ai_1 _4443_ (.B1(_3792_),
    .Y(_3793_),
    .A1(_3707_),
    .A2(_3789_));
 sg13g2_nand2_1 _4444_ (.Y(_3794_),
    .A(_3786_),
    .B(net148));
 sg13g2_nand3_1 _4445_ (.B(net116),
    .C(_3794_),
    .A(_3793_),
    .Y(_3795_));
 sg13g2_nor2b_1 _4446_ (.A(_3788_),
    .B_N(_3795_),
    .Y(_3796_));
 sg13g2_nand2_1 _4447_ (.Y(_3797_),
    .A(_3730_),
    .B(_3771_));
 sg13g2_nand3_1 _4448_ (.B(_3797_),
    .C(net126),
    .A(_3796_),
    .Y(_3798_));
 sg13g2_nand2_1 _4449_ (.Y(_3799_),
    .A(_3797_),
    .B(_3759_));
 sg13g2_nand2_1 _4450_ (.Y(_3800_),
    .A(_3779_),
    .B(_3692_));
 sg13g2_nand2_1 _4451_ (.Y(_3801_),
    .A(_3800_),
    .B(_3697_));
 sg13g2_nand2_1 _4452_ (.Y(_3802_),
    .A(_3738_),
    .B(_3679_));
 sg13g2_nand3_1 _4453_ (.B(_3802_),
    .C(_3786_),
    .A(_3782_),
    .Y(_3803_));
 sg13g2_nand2_1 _4454_ (.Y(_3804_),
    .A(_3803_),
    .B(_3709_));
 sg13g2_nand3_1 _4455_ (.B(net101),
    .C(_3804_),
    .A(_3801_),
    .Y(_3805_));
 sg13g2_nand2_1 _4456_ (.Y(_3806_),
    .A(_3805_),
    .B(_3795_));
 sg13g2_nand2_1 _4457_ (.Y(_3807_),
    .A(_3799_),
    .B(_3806_));
 sg13g2_nand2_1 _4458_ (.Y(_3808_),
    .A(_3798_),
    .B(_3807_));
 sg13g2_buf_8 _4459_ (.A(_3808_),
    .X(_3809_));
 sg13g2_xnor2_1 _4460_ (.Y(_3810_),
    .A(_3777_),
    .B(_3809_));
 sg13g2_nor2b_1 _4461_ (.A(_3776_),
    .B_N(_3810_),
    .Y(_3811_));
 sg13g2_nor2b_1 _4462_ (.A(_3810_),
    .B_N(_3776_),
    .Y(_3812_));
 sg13g2_nor3_1 _4463_ (.A(net63),
    .B(_3811_),
    .C(_3812_),
    .Y(_3813_));
 sg13g2_buf_1 _4464_ (.A(_3758_),
    .X(_3814_));
 sg13g2_buf_1 _4465_ (.A(_3814_),
    .X(_3815_));
 sg13g2_xnor2_1 _4466_ (.Y(_3816_),
    .A(_3777_),
    .B(net125));
 sg13g2_nor2_1 _4467_ (.A(_0031_),
    .B(_3809_),
    .Y(_3817_));
 sg13g2_inv_1 _4468_ (.Y(_3818_),
    .A(\i_transform.image_y[2] ));
 sg13g2_xnor2_1 _4469_ (.Y(_3819_),
    .A(_3818_),
    .B(_3809_));
 sg13g2_inv_1 _4470_ (.Y(_3820_),
    .A(_3763_));
 sg13g2_inv_1 _4471_ (.Y(_3821_),
    .A(\i_transform.image_y[0] ));
 sg13g2_nor2_1 _4472_ (.A(_3821_),
    .B(_3771_),
    .Y(_3822_));
 sg13g2_xnor2_1 _4473_ (.Y(_3823_),
    .A(_0032_),
    .B(_3763_));
 sg13g2_inv_1 _4474_ (.Y(_3824_),
    .A(_3823_));
 sg13g2_a22oi_1 _4475_ (.Y(_3825_),
    .B1(_3822_),
    .B2(_3824_),
    .A2(_3820_),
    .A1(\i_transform.image_y[1] ));
 sg13g2_nor2_1 _4476_ (.A(_3819_),
    .B(_3825_),
    .Y(_3826_));
 sg13g2_nor2_1 _4477_ (.A(_3817_),
    .B(_3826_),
    .Y(_3827_));
 sg13g2_nand2_1 _4478_ (.Y(_3828_),
    .A(_3699_),
    .B(_3711_));
 sg13g2_nand2_1 _4479_ (.Y(_3829_),
    .A(_3828_),
    .B(_3741_));
 sg13g2_nand2_1 _4480_ (.Y(_3830_),
    .A(_3724_),
    .B(_3728_));
 sg13g2_nand2_1 _4481_ (.Y(_3831_),
    .A(_3830_),
    .B(net101));
 sg13g2_nand2_1 _4482_ (.Y(_3832_),
    .A(_3829_),
    .B(_3831_));
 sg13g2_nor2_1 _4483_ (.A(_3753_),
    .B(_3832_),
    .Y(_3833_));
 sg13g2_nand2_1 _4484_ (.Y(_3834_),
    .A(_3710_),
    .B(_3790_));
 sg13g2_nand3_1 _4485_ (.B(_3686_),
    .C(net134),
    .A(_3682_),
    .Y(_3835_));
 sg13g2_nand2_1 _4486_ (.Y(_3836_),
    .A(_3783_),
    .B(_3835_));
 sg13g2_nand3_1 _4487_ (.B(net101),
    .C(_3836_),
    .A(_3834_),
    .Y(_3837_));
 sg13g2_nor2_1 _4488_ (.A(_3785_),
    .B(_3791_),
    .Y(_3838_));
 sg13g2_nand2_1 _4489_ (.Y(_3839_),
    .A(_3838_),
    .B(net116));
 sg13g2_nand2_1 _4490_ (.Y(_3840_),
    .A(_3837_),
    .B(_3839_));
 sg13g2_nand3_1 _4491_ (.B(_3806_),
    .C(_3840_),
    .A(_3833_),
    .Y(_3841_));
 sg13g2_nand2_1 _4492_ (.Y(_3842_),
    .A(_3841_),
    .B(net126));
 sg13g2_nor2_1 _4493_ (.A(_3709_),
    .B(_3706_),
    .Y(_3843_));
 sg13g2_nand2_1 _4494_ (.Y(_3844_),
    .A(_3791_),
    .B(net101));
 sg13g2_nand2_1 _4495_ (.Y(_3845_),
    .A(_3785_),
    .B(_3709_));
 sg13g2_nand2_1 _4496_ (.Y(_3846_),
    .A(_3845_),
    .B(net116));
 sg13g2_o21ai_1 _4497_ (.B1(_3846_),
    .Y(_3847_),
    .A1(_3843_),
    .A2(_3844_));
 sg13g2_inv_1 _4498_ (.Y(_3848_),
    .A(_3847_));
 sg13g2_nand2_1 _4499_ (.Y(_3849_),
    .A(_3842_),
    .B(_3848_));
 sg13g2_nand3_1 _4500_ (.B(net126),
    .C(_3847_),
    .A(_3841_),
    .Y(_3850_));
 sg13g2_nand2_1 _4501_ (.Y(_3851_),
    .A(_3849_),
    .B(_3850_));
 sg13g2_buf_8 _4502_ (.A(_3851_),
    .X(_3852_));
 sg13g2_xor2_1 _4503_ (.B(_3852_),
    .A(\i_transform.image_y[4] ),
    .X(_3853_));
 sg13g2_xnor2_1 _4504_ (.Y(_3854_),
    .A(_0027_),
    .B(net125));
 sg13g2_buf_1 _4505_ (.A(\i_transform.image_y[5] ),
    .X(_3855_));
 sg13g2_a21oi_1 _4506_ (.A1(_3837_),
    .A2(_3839_),
    .Y(_3856_),
    .B1(_3847_));
 sg13g2_nand4_1 _4507_ (.B(_3771_),
    .C(_3730_),
    .A(_3806_),
    .Y(_3857_),
    .D(_3856_));
 sg13g2_nand3_1 _4508_ (.B(net126),
    .C(_3844_),
    .A(_3857_),
    .Y(_3858_));
 sg13g2_nand3_1 _4509_ (.B(_3751_),
    .C(_3814_),
    .A(_3791_),
    .Y(_3859_));
 sg13g2_nand2_1 _4510_ (.Y(_3860_),
    .A(_3858_),
    .B(_3859_));
 sg13g2_buf_1 _4511_ (.A(_3860_),
    .X(_3861_));
 sg13g2_xnor2_1 _4512_ (.Y(_3862_),
    .A(_3855_),
    .B(net79));
 sg13g2_inv_1 _4513_ (.Y(_3863_),
    .A(_3862_));
 sg13g2_nor2_1 _4514_ (.A(_3854_),
    .B(_3863_),
    .Y(_3864_));
 sg13g2_nand2_1 _4515_ (.Y(_3865_),
    .A(_3833_),
    .B(_3806_));
 sg13g2_nand2_1 _4516_ (.Y(_3866_),
    .A(_3865_),
    .B(net126));
 sg13g2_nand2_1 _4517_ (.Y(_3867_),
    .A(_3866_),
    .B(_3840_));
 sg13g2_inv_1 _4518_ (.Y(_3868_),
    .A(_3840_));
 sg13g2_nand3_1 _4519_ (.B(net126),
    .C(_3868_),
    .A(_3865_),
    .Y(_3869_));
 sg13g2_nand2_1 _4520_ (.Y(_3870_),
    .A(_3867_),
    .B(_3869_));
 sg13g2_buf_8 _4521_ (.A(_3870_),
    .X(_3871_));
 sg13g2_xnor2_1 _4522_ (.Y(_3872_),
    .A(\i_transform.image_y[3] ),
    .B(_3871_));
 sg13g2_nand3b_1 _4523_ (.B(_3864_),
    .C(_3872_),
    .Y(_3873_),
    .A_N(_3853_));
 sg13g2_nor2_1 _4524_ (.A(_0029_),
    .B(net72),
    .Y(_3874_));
 sg13g2_nor2_1 _4525_ (.A(_0030_),
    .B(_3871_),
    .Y(_3875_));
 sg13g2_nand2b_1 _4526_ (.Y(_3876_),
    .B(_3875_),
    .A_N(_3853_));
 sg13g2_nand2b_1 _4527_ (.Y(_3877_),
    .B(_3876_),
    .A_N(_3874_));
 sg13g2_nor2_1 _4528_ (.A(_3764_),
    .B(net79),
    .Y(_3878_));
 sg13g2_inv_1 _4529_ (.Y(_3879_),
    .A(_3854_));
 sg13g2_inv_1 _4530_ (.Y(_3880_),
    .A(_3773_));
 sg13g2_nor2_1 _4531_ (.A(_3880_),
    .B(net125),
    .Y(_3881_));
 sg13g2_a21o_1 _4532_ (.A2(_3879_),
    .A1(_3878_),
    .B1(_3881_),
    .X(_3882_));
 sg13g2_a21oi_1 _4533_ (.A1(_3877_),
    .A2(_3864_),
    .Y(_3883_),
    .B1(_3882_));
 sg13g2_o21ai_1 _4534_ (.B1(_3883_),
    .Y(_3884_),
    .A1(_3827_),
    .A2(_3873_));
 sg13g2_buf_1 _4535_ (.A(net68),
    .X(_3885_));
 sg13g2_a21oi_1 _4536_ (.A1(_3884_),
    .A2(_3816_),
    .Y(_3886_),
    .B1(net62));
 sg13g2_o21ai_1 _4537_ (.B1(_3886_),
    .Y(_3887_),
    .A1(_3816_),
    .A2(_3884_));
 sg13g2_o21ai_1 _4538_ (.B1(_3887_),
    .Y(_3888_),
    .A1(_3671_),
    .A2(_3813_));
 sg13g2_buf_2 _4539_ (.A(\i_bitmap.in[7] ),
    .X(_3889_));
 sg13g2_inv_1 _4540_ (.Y(_3890_),
    .A(_3889_));
 sg13g2_xnor2_1 _4541_ (.Y(_3891_),
    .A(_3754_),
    .B(_3700_));
 sg13g2_nand2b_1 _4542_ (.Y(_3892_),
    .B(orient),
    .A_N(_3891_));
 sg13g2_nand2_1 _4543_ (.Y(_3893_),
    .A(_3891_),
    .B(_3755_));
 sg13g2_nand2_1 _4544_ (.Y(_3894_),
    .A(_3892_),
    .B(_3893_));
 sg13g2_buf_1 _4545_ (.A(_3894_),
    .X(_3895_));
 sg13g2_buf_1 _4546_ (.A(net124),
    .X(_3896_));
 sg13g2_buf_1 _4547_ (.A(net115),
    .X(_3897_));
 sg13g2_xnor2_1 _4548_ (.Y(_3898_),
    .A(_3890_),
    .B(net100));
 sg13g2_a21oi_1 _4549_ (.A1(_3780_),
    .A2(_3787_),
    .Y(_3899_),
    .B1(net101));
 sg13g2_nand3_1 _4550_ (.B(net101),
    .C(_3794_),
    .A(_3793_),
    .Y(_3900_));
 sg13g2_nor2b_1 _4551_ (.A(_3899_),
    .B_N(_3900_),
    .Y(_3901_));
 sg13g2_nand3_1 _4552_ (.B(_3725_),
    .C(_3711_),
    .A(_3699_),
    .Y(_3902_));
 sg13g2_nand3_1 _4553_ (.B(_3705_),
    .C(_3728_),
    .A(_3724_),
    .Y(_3903_));
 sg13g2_nand2_1 _4554_ (.Y(_3904_),
    .A(_3902_),
    .B(_3903_));
 sg13g2_nand2_1 _4555_ (.Y(_3905_),
    .A(_3766_),
    .B(_3725_));
 sg13g2_nand2_1 _4556_ (.Y(_3906_),
    .A(_3768_),
    .B(_3705_));
 sg13g2_nand2_2 _4557_ (.Y(_3907_),
    .A(_3905_),
    .B(_3906_));
 sg13g2_nand2_1 _4558_ (.Y(_3908_),
    .A(_3904_),
    .B(_3907_));
 sg13g2_inv_2 _4559_ (.Y(_3909_),
    .A(net124));
 sg13g2_nand3_1 _4560_ (.B(_3908_),
    .C(_3909_),
    .A(_3901_),
    .Y(_3910_));
 sg13g2_nand2_1 _4561_ (.Y(_3911_),
    .A(_3908_),
    .B(_3909_));
 sg13g2_nand3_1 _4562_ (.B(net116),
    .C(_3804_),
    .A(_3801_),
    .Y(_3912_));
 sg13g2_nand2_1 _4563_ (.Y(_3913_),
    .A(_3912_),
    .B(_3900_));
 sg13g2_nand2_1 _4564_ (.Y(_3914_),
    .A(_3911_),
    .B(_3913_));
 sg13g2_nand2_1 _4565_ (.Y(_3915_),
    .A(_3910_),
    .B(_3914_));
 sg13g2_buf_8 _4566_ (.A(_3915_),
    .X(_3916_));
 sg13g2_inv_1 _4567_ (.Y(_3917_),
    .A(_3916_));
 sg13g2_nand3_1 _4568_ (.B(_3740_),
    .C(_3725_),
    .A(_3733_),
    .Y(_3918_));
 sg13g2_nand3_1 _4569_ (.B(_3750_),
    .C(_3705_),
    .A(_3746_),
    .Y(_3919_));
 sg13g2_nand2_2 _4570_ (.Y(_3920_),
    .A(_3918_),
    .B(_3919_));
 sg13g2_nand4_1 _4571_ (.B(_3902_),
    .C(_3909_),
    .A(_3920_),
    .Y(_3921_),
    .D(_3903_));
 sg13g2_o21ai_1 _4572_ (.B1(_3904_),
    .Y(_3922_),
    .A1(_3895_),
    .A2(_3907_));
 sg13g2_nand2_1 _4573_ (.Y(_3923_),
    .A(_3921_),
    .B(_3922_));
 sg13g2_buf_8 _4574_ (.A(_3923_),
    .X(_3924_));
 sg13g2_inv_1 _4575_ (.Y(_3925_),
    .A(_3924_));
 sg13g2_xor2_1 _4576_ (.B(_3924_),
    .A(\i_transform.image_y[1] ),
    .X(_3926_));
 sg13g2_nand2_1 _4577_ (.Y(_3927_),
    .A(_3920_),
    .B(_0033_));
 sg13g2_nand2_1 _4578_ (.Y(_3928_),
    .A(_3926_),
    .B(_3927_));
 sg13g2_o21ai_1 _4579_ (.B1(_3928_),
    .Y(_3929_),
    .A1(_0032_),
    .A2(_3925_));
 sg13g2_xnor2_1 _4580_ (.Y(_3930_),
    .A(_0031_),
    .B(_3916_));
 sg13g2_nand2_1 _4581_ (.Y(_3931_),
    .A(_3929_),
    .B(_3930_));
 sg13g2_o21ai_1 _4582_ (.B1(_3931_),
    .Y(_3932_),
    .A1(_3818_),
    .A2(_3917_));
 sg13g2_nand3_1 _4583_ (.B(net116),
    .C(_3836_),
    .A(_3834_),
    .Y(_3933_));
 sg13g2_nand2_1 _4584_ (.Y(_3934_),
    .A(_3838_),
    .B(net101));
 sg13g2_nand2_1 _4585_ (.Y(_3935_),
    .A(_3933_),
    .B(_3934_));
 sg13g2_a21oi_1 _4586_ (.A1(_3902_),
    .A2(_3903_),
    .Y(_3936_),
    .B1(_3920_));
 sg13g2_nand2_1 _4587_ (.Y(_3937_),
    .A(_3936_),
    .B(_3913_));
 sg13g2_nand2_1 _4588_ (.Y(_3938_),
    .A(_3937_),
    .B(_3909_));
 sg13g2_xnor2_1 _4589_ (.Y(_3939_),
    .A(_3935_),
    .B(_3938_));
 sg13g2_buf_1 _4590_ (.A(_3939_),
    .X(_3940_));
 sg13g2_xnor2_1 _4591_ (.Y(_3941_),
    .A(_0030_),
    .B(net78));
 sg13g2_xnor2_1 _4592_ (.Y(_3942_),
    .A(_3773_),
    .B(net115));
 sg13g2_nand2_1 _4593_ (.Y(_3943_),
    .A(_3791_),
    .B(net116));
 sg13g2_nand2_1 _4594_ (.Y(_3944_),
    .A(_3845_),
    .B(net101));
 sg13g2_o21ai_1 _4595_ (.B1(_3944_),
    .Y(_3945_),
    .A1(_3843_),
    .A2(_3943_));
 sg13g2_buf_1 _4596_ (.A(_3945_),
    .X(_3946_));
 sg13g2_inv_1 _4597_ (.Y(_3947_),
    .A(_3935_));
 sg13g2_nor2_1 _4598_ (.A(_3946_),
    .B(_3947_),
    .Y(_3948_));
 sg13g2_nand3_1 _4599_ (.B(_3913_),
    .C(_3948_),
    .A(_3936_),
    .Y(_3949_));
 sg13g2_buf_1 _4600_ (.A(_3909_),
    .X(_3950_));
 sg13g2_nand3_1 _4601_ (.B(net99),
    .C(_3943_),
    .A(_3949_),
    .Y(_3951_));
 sg13g2_nand3_1 _4602_ (.B(_3895_),
    .C(_3741_),
    .A(_3791_),
    .Y(_3952_));
 sg13g2_nand2_1 _4603_ (.Y(_3953_),
    .A(_3951_),
    .B(_3952_));
 sg13g2_buf_2 _4604_ (.A(_3953_),
    .X(_3954_));
 sg13g2_xnor2_1 _4605_ (.Y(_3955_),
    .A(_3764_),
    .B(net75));
 sg13g2_nand2b_1 _4606_ (.Y(_3956_),
    .B(_3955_),
    .A_N(_3942_));
 sg13g2_inv_1 _4607_ (.Y(_3957_),
    .A(_3956_));
 sg13g2_nand2_1 _4608_ (.Y(_3958_),
    .A(_3947_),
    .B(net99));
 sg13g2_nand3_1 _4609_ (.B(_3946_),
    .C(_3958_),
    .A(_3938_),
    .Y(_3959_));
 sg13g2_nand3_1 _4610_ (.B(_3913_),
    .C(_3935_),
    .A(_3936_),
    .Y(_3960_));
 sg13g2_inv_1 _4611_ (.Y(_3961_),
    .A(_3946_));
 sg13g2_nand3_1 _4612_ (.B(net99),
    .C(_3961_),
    .A(_3960_),
    .Y(_3962_));
 sg13g2_nand2_1 _4613_ (.Y(_0285_),
    .A(_3959_),
    .B(_3962_));
 sg13g2_buf_8 _4614_ (.A(_0285_),
    .X(_0286_));
 sg13g2_xnor2_1 _4615_ (.Y(_0287_),
    .A(_0029_),
    .B(_0286_));
 sg13g2_inv_1 _4616_ (.Y(_0288_),
    .A(_0287_));
 sg13g2_nand4_1 _4617_ (.B(_3941_),
    .C(_3957_),
    .A(_3932_),
    .Y(_0289_),
    .D(_0288_));
 sg13g2_nand2_1 _4618_ (.Y(_0290_),
    .A(net78),
    .B(\i_transform.image_y[3] ));
 sg13g2_inv_1 _4619_ (.Y(_0291_),
    .A(_0286_));
 sg13g2_nand2_1 _4620_ (.Y(_0292_),
    .A(_0291_),
    .B(\i_transform.image_y[4] ));
 sg13g2_o21ai_1 _4621_ (.B1(_0292_),
    .Y(_0293_),
    .A1(_0290_),
    .A2(_0287_));
 sg13g2_nand2_1 _4622_ (.Y(_0294_),
    .A(net75),
    .B(_3855_));
 sg13g2_nand2_1 _4623_ (.Y(_0295_),
    .A(net115),
    .B(_3672_));
 sg13g2_o21ai_1 _4624_ (.B1(_0295_),
    .Y(_0296_),
    .A1(_3942_),
    .A2(_0294_));
 sg13g2_a21oi_1 _4625_ (.A1(_0293_),
    .A2(_3957_),
    .Y(_0297_),
    .B1(_0296_));
 sg13g2_nand2_1 _4626_ (.Y(_0298_),
    .A(_0289_),
    .B(_0297_));
 sg13g2_xnor2_1 _4627_ (.Y(_0299_),
    .A(_3898_),
    .B(_0298_));
 sg13g2_inv_1 _4628_ (.Y(_0300_),
    .A(_3563_));
 sg13g2_nand3_1 _4629_ (.B(_3505_),
    .C(_0059_),
    .A(net127),
    .Y(_0301_));
 sg13g2_o21ai_1 _4630_ (.B1(_0301_),
    .Y(_0302_),
    .A1(_3568_),
    .A2(_0300_));
 sg13g2_nand2_1 _4631_ (.Y(_0303_),
    .A(_3552_),
    .B(_3554_));
 sg13g2_nand2_1 _4632_ (.Y(_0304_),
    .A(_0303_),
    .B(_3549_));
 sg13g2_inv_1 _4633_ (.Y(_0305_),
    .A(_3579_));
 sg13g2_o21ai_1 _4634_ (.B1(_3577_),
    .Y(_0306_),
    .A1(_3575_),
    .A2(_3576_));
 sg13g2_o21ai_1 _4635_ (.B1(_0306_),
    .Y(_0307_),
    .A1(_0304_),
    .A2(_0305_));
 sg13g2_buf_1 _4636_ (.A(\i_transform.track_y[5] ),
    .X(_0308_));
 sg13g2_nor2_1 _4637_ (.A(_3565_),
    .B(_0308_),
    .Y(_0309_));
 sg13g2_inv_1 _4638_ (.Y(_0310_),
    .A(\i_transform.track_y[7] ));
 sg13g2_nand2_1 _4639_ (.Y(_0311_),
    .A(_0309_),
    .B(_0310_));
 sg13g2_nor2_1 _4640_ (.A(_3556_),
    .B(_0311_),
    .Y(_0312_));
 sg13g2_nor2_1 _4641_ (.A(_0312_),
    .B(_3559_),
    .Y(_0313_));
 sg13g2_nor2_1 _4642_ (.A(\i_transform.track_y[9] ),
    .B(_0313_),
    .Y(_0314_));
 sg13g2_a221oi_1 _4643_ (.B2(_3570_),
    .C1(_0314_),
    .B1(_0307_),
    .A1(_3560_),
    .Y(_0315_),
    .A2(_0302_));
 sg13g2_inv_1 _4644_ (.Y(_0316_),
    .A(_3582_));
 sg13g2_a21o_1 _4645_ (.A2(_3588_),
    .A1(_0316_),
    .B1(_3580_),
    .X(_0317_));
 sg13g2_nand2_1 _4646_ (.Y(_0318_),
    .A(_0315_),
    .B(_0317_));
 sg13g2_buf_1 _4647_ (.A(_0318_),
    .X(_0319_));
 sg13g2_buf_1 _4648_ (.A(net80),
    .X(_0320_));
 sg13g2_nand2_1 _4649_ (.Y(_0321_),
    .A(_0299_),
    .B(net77));
 sg13g2_xnor2_1 _4650_ (.Y(_0322_),
    .A(_3672_),
    .B(_3924_));
 sg13g2_nor2b_1 _4651_ (.A(_3907_),
    .B_N(_3855_),
    .Y(_0323_));
 sg13g2_nand2_1 _4652_ (.Y(_0324_),
    .A(_0322_),
    .B(_0323_));
 sg13g2_nor2b_1 _4653_ (.A(net77),
    .B_N(_0324_),
    .Y(_0325_));
 sg13g2_xnor2_1 _4654_ (.Y(_0326_),
    .A(_3889_),
    .B(_3916_));
 sg13g2_inv_1 _4655_ (.Y(_0327_),
    .A(_0326_));
 sg13g2_nor2_1 _4656_ (.A(_3880_),
    .B(_3924_),
    .Y(_0328_));
 sg13g2_inv_1 _4657_ (.Y(_0329_),
    .A(_0328_));
 sg13g2_nand3_1 _4658_ (.B(_0327_),
    .C(_0329_),
    .A(_0325_),
    .Y(_0330_));
 sg13g2_a21oi_1 _4659_ (.A1(_0324_),
    .A2(_0329_),
    .Y(_0331_),
    .B1(_0327_));
 sg13g2_inv_2 _4660_ (.Y(_0332_),
    .A(_0319_));
 sg13g2_buf_1 _4661_ (.A(_3591_),
    .X(_0333_));
 sg13g2_a21oi_1 _4662_ (.A1(_0331_),
    .A2(net76),
    .Y(_0334_),
    .B1(_0333_));
 sg13g2_nand3_1 _4663_ (.B(_0330_),
    .C(_0334_),
    .A(_0321_),
    .Y(_0335_));
 sg13g2_nor2_1 _4664_ (.A(net84),
    .B(_3649_),
    .Y(_0336_));
 sg13g2_buf_1 _4665_ (.A(_0336_),
    .X(_0337_));
 sg13g2_inv_1 _4666_ (.Y(_0338_),
    .A(_3777_));
 sg13g2_nand2_1 _4667_ (.Y(_0339_),
    .A(net71),
    .B(_0338_));
 sg13g2_nand3_1 _4668_ (.B(_0335_),
    .C(_0339_),
    .A(_3888_),
    .Y(_0340_));
 sg13g2_buf_2 _4669_ (.A(_0340_),
    .X(_0341_));
 sg13g2_nor2_2 _4670_ (.A(\i_orchestrator.update_transform ),
    .B(_3492_),
    .Y(_0342_));
 sg13g2_buf_1 _4671_ (.A(_0342_),
    .X(_0343_));
 sg13g2_nand2_2 _4672_ (.Y(_0344_),
    .A(_0341_),
    .B(_0343_));
 sg13g2_inv_1 _4673_ (.Y(_0345_),
    .A(_0344_));
 sg13g2_buf_1 _4674_ (.A(_0345_),
    .X(_0346_));
 sg13g2_buf_2 _4675_ (.A(_0013_),
    .X(_0347_));
 sg13g2_xnor2_1 _4676_ (.Y(_0348_),
    .A(_0347_),
    .B(net133));
 sg13g2_buf_2 _4677_ (.A(\i_bitmap.in[0] ),
    .X(_0349_));
 sg13g2_xnor2_1 _4678_ (.Y(_0350_),
    .A(_0349_),
    .B(net133));
 sg13g2_inv_1 _4679_ (.Y(_0351_),
    .A(_0350_));
 sg13g2_nor2_1 _4680_ (.A(_0348_),
    .B(_0351_),
    .Y(_0352_));
 sg13g2_inv_1 _4681_ (.Y(_0353_),
    .A(_0352_));
 sg13g2_inv_1 _4682_ (.Y(_0354_),
    .A(\i_transform.image_x[5] ));
 sg13g2_nand2_1 _4683_ (.Y(_0355_),
    .A(net79),
    .B(_0354_));
 sg13g2_nand3_1 _4684_ (.B(\i_transform.image_x[5] ),
    .C(_3859_),
    .A(_3858_),
    .Y(_0356_));
 sg13g2_buf_1 _4685_ (.A(\i_capsule.tf_x[0] ),
    .X(_0357_));
 sg13g2_inv_1 _4686_ (.Y(_0358_),
    .A(_0357_));
 sg13g2_nor2_1 _4687_ (.A(_0358_),
    .B(net133),
    .Y(_0359_));
 sg13g2_nor2_1 _4688_ (.A(_0357_),
    .B(_3760_),
    .Y(_0360_));
 sg13g2_nor2_1 _4689_ (.A(_0359_),
    .B(_0360_),
    .Y(_0361_));
 sg13g2_nand3_1 _4690_ (.B(_0356_),
    .C(_0361_),
    .A(_0355_),
    .Y(_0362_));
 sg13g2_nor2_1 _4691_ (.A(_0353_),
    .B(_0362_),
    .Y(_0363_));
 sg13g2_nor2_1 _4692_ (.A(_0018_),
    .B(_3771_),
    .Y(_0364_));
 sg13g2_inv_1 _4693_ (.Y(_0365_),
    .A(\i_transform.image_x[2] ));
 sg13g2_nand2_1 _4694_ (.Y(_0366_),
    .A(_3809_),
    .B(_0365_));
 sg13g2_nand3_1 _4695_ (.B(_3807_),
    .C(\i_transform.image_x[2] ),
    .A(_3798_),
    .Y(_0367_));
 sg13g2_and2_1 _4696_ (.A(_0366_),
    .B(_0367_),
    .X(_0368_));
 sg13g2_buf_1 _4697_ (.A(_0368_),
    .X(_0369_));
 sg13g2_inv_1 _4698_ (.Y(_0370_),
    .A(\i_transform.image_x[1] ));
 sg13g2_nor2_1 _4699_ (.A(_0370_),
    .B(_3763_),
    .Y(_0371_));
 sg13g2_nand2_1 _4700_ (.Y(_0372_),
    .A(_3763_),
    .B(_0370_));
 sg13g2_nor2b_1 _4701_ (.A(_0371_),
    .B_N(_0372_),
    .Y(_0373_));
 sg13g2_nand2_1 _4702_ (.Y(_0374_),
    .A(_0369_),
    .B(_0373_));
 sg13g2_buf_1 _4703_ (.A(\i_transform.image_x[3] ),
    .X(_0375_));
 sg13g2_xnor2_1 _4704_ (.Y(_0376_),
    .A(_0375_),
    .B(_3871_));
 sg13g2_inv_4 _4705_ (.A(_0376_),
    .Y(_0377_));
 sg13g2_buf_1 _4706_ (.A(\i_transform.image_x[4] ),
    .X(_0378_));
 sg13g2_inv_1 _4707_ (.Y(_0379_),
    .A(_0378_));
 sg13g2_nand2_1 _4708_ (.Y(_0380_),
    .A(net72),
    .B(_0379_));
 sg13g2_nand3_1 _4709_ (.B(_3850_),
    .C(_0378_),
    .A(_3849_),
    .Y(_0381_));
 sg13g2_nand2_2 _4710_ (.Y(_0382_),
    .A(_0380_),
    .B(_0381_));
 sg13g2_nor3_1 _4711_ (.A(_0374_),
    .B(_0377_),
    .C(_0382_),
    .Y(_0383_));
 sg13g2_nand3_1 _4712_ (.B(_0364_),
    .C(_0383_),
    .A(_0363_),
    .Y(_0384_));
 sg13g2_nand2_1 _4713_ (.Y(_0385_),
    .A(net72),
    .B(_0378_));
 sg13g2_nand3_1 _4714_ (.B(_3850_),
    .C(_0379_),
    .A(_3849_),
    .Y(_0386_));
 sg13g2_nand2_1 _4715_ (.Y(_0387_),
    .A(_0385_),
    .B(_0386_));
 sg13g2_nor2_1 _4716_ (.A(_0016_),
    .B(_3871_),
    .Y(_0388_));
 sg13g2_nor2_1 _4717_ (.A(_0015_),
    .B(net72),
    .Y(_0389_));
 sg13g2_a21oi_1 _4718_ (.A1(_0387_),
    .A2(_0388_),
    .Y(_0390_),
    .B1(_0389_));
 sg13g2_nand3_1 _4719_ (.B(_0367_),
    .C(_0371_),
    .A(_0366_),
    .Y(_0391_));
 sg13g2_nor2_1 _4720_ (.A(_0017_),
    .B(_3809_),
    .Y(_0392_));
 sg13g2_inv_1 _4721_ (.Y(_0393_),
    .A(_0392_));
 sg13g2_nand2_1 _4722_ (.Y(_0394_),
    .A(_0391_),
    .B(_0393_));
 sg13g2_nand3_1 _4723_ (.B(_0394_),
    .C(_0376_),
    .A(_0387_),
    .Y(_0395_));
 sg13g2_nand2_1 _4724_ (.Y(_0396_),
    .A(_0390_),
    .B(_0395_));
 sg13g2_nand2_1 _4725_ (.Y(_0397_),
    .A(_0396_),
    .B(_0363_));
 sg13g2_inv_1 _4726_ (.Y(_0398_),
    .A(_0014_));
 sg13g2_inv_1 _4727_ (.Y(_0399_),
    .A(_0360_));
 sg13g2_nand4_1 _4728_ (.B(_0398_),
    .C(_3859_),
    .A(_3858_),
    .Y(_0400_),
    .D(_0399_));
 sg13g2_nand2b_1 _4729_ (.Y(_0401_),
    .B(_0400_),
    .A_N(_0359_));
 sg13g2_nand2_1 _4730_ (.Y(_0402_),
    .A(_0401_),
    .B(_0352_));
 sg13g2_buf_2 _4731_ (.A(\i_bitmap.in[1] ),
    .X(_0403_));
 sg13g2_nor2b_1 _4732_ (.A(net133),
    .B_N(_0349_),
    .Y(_0404_));
 sg13g2_a22oi_1 _4733_ (.Y(_0405_),
    .B1(_0347_),
    .B2(_0404_),
    .A2(_0403_),
    .A1(_3760_));
 sg13g2_nand2_1 _4734_ (.Y(_0406_),
    .A(_0402_),
    .B(_0405_));
 sg13g2_inv_1 _4735_ (.Y(_0407_),
    .A(_0406_));
 sg13g2_nand3_1 _4736_ (.B(_0397_),
    .C(_0407_),
    .A(_0384_),
    .Y(_0408_));
 sg13g2_buf_1 _4737_ (.A(_0021_),
    .X(_0409_));
 sg13g2_xnor2_1 _4738_ (.Y(_0410_),
    .A(_0409_),
    .B(net133));
 sg13g2_inv_1 _4739_ (.Y(_0411_),
    .A(_0410_));
 sg13g2_nand2_1 _4740_ (.Y(_0412_),
    .A(_0408_),
    .B(_0411_));
 sg13g2_a21oi_1 _4741_ (.A1(_0396_),
    .A2(_0363_),
    .Y(_0413_),
    .B1(_0406_));
 sg13g2_nand3_1 _4742_ (.B(_0410_),
    .C(_0384_),
    .A(_0413_),
    .Y(_0414_));
 sg13g2_nand2_1 _4743_ (.Y(_0415_),
    .A(_0412_),
    .B(_0414_));
 sg13g2_nand2_1 _4744_ (.Y(_0416_),
    .A(_0415_),
    .B(net80));
 sg13g2_inv_1 _4745_ (.Y(_0417_),
    .A(_0347_));
 sg13g2_xnor2_1 _4746_ (.Y(_0418_),
    .A(_0417_),
    .B(_3871_));
 sg13g2_nor2_1 _4747_ (.A(_0398_),
    .B(_3771_),
    .Y(_0419_));
 sg13g2_xnor2_1 _4748_ (.Y(_0420_),
    .A(_0358_),
    .B(_3763_));
 sg13g2_nand2b_1 _4749_ (.Y(_0421_),
    .B(_0420_),
    .A_N(_0419_));
 sg13g2_inv_1 _4750_ (.Y(_0422_),
    .A(_0020_));
 sg13g2_nand2_1 _4751_ (.Y(_0423_),
    .A(_3763_),
    .B(_0422_));
 sg13g2_nand2_1 _4752_ (.Y(_0424_),
    .A(_0421_),
    .B(_0423_));
 sg13g2_xnor2_1 _4753_ (.Y(_0425_),
    .A(_0019_),
    .B(_3809_));
 sg13g2_nand2_1 _4754_ (.Y(_0426_),
    .A(_0424_),
    .B(_0425_));
 sg13g2_nand2_1 _4755_ (.Y(_0427_),
    .A(_3809_),
    .B(_0349_));
 sg13g2_nand2_1 _4756_ (.Y(_0428_),
    .A(_0426_),
    .B(_0427_));
 sg13g2_nand2b_1 _4757_ (.Y(_0429_),
    .B(_0428_),
    .A_N(_0418_));
 sg13g2_inv_1 _4758_ (.Y(_0430_),
    .A(_0403_));
 sg13g2_inv_1 _4759_ (.Y(_0431_),
    .A(_3871_));
 sg13g2_nor2_1 _4760_ (.A(_0430_),
    .B(_0431_),
    .Y(_0432_));
 sg13g2_inv_1 _4761_ (.Y(_0433_),
    .A(_0432_));
 sg13g2_nand2_1 _4762_ (.Y(_0434_),
    .A(_0429_),
    .B(_0433_));
 sg13g2_inv_1 _4763_ (.Y(_0435_),
    .A(_0409_));
 sg13g2_xnor2_1 _4764_ (.Y(_0436_),
    .A(_0435_),
    .B(net72));
 sg13g2_inv_1 _4765_ (.Y(_0437_),
    .A(_0436_));
 sg13g2_nand2_1 _4766_ (.Y(_0438_),
    .A(_0434_),
    .B(_0437_));
 sg13g2_nand3_1 _4767_ (.B(_0433_),
    .C(_0436_),
    .A(_0429_),
    .Y(_0439_));
 sg13g2_nand2_1 _4768_ (.Y(_0440_),
    .A(_0438_),
    .B(_0439_));
 sg13g2_a21oi_1 _4769_ (.A1(_0440_),
    .A2(net76),
    .Y(_0441_),
    .B1(_3591_));
 sg13g2_nand2_1 _4770_ (.Y(_0442_),
    .A(_0416_),
    .B(_0441_));
 sg13g2_xnor2_1 _4771_ (.Y(_0443_),
    .A(_0409_),
    .B(net124));
 sg13g2_nand3_1 _4772_ (.B(_3962_),
    .C(_0378_),
    .A(_3959_),
    .Y(_0444_));
 sg13g2_nand3_1 _4773_ (.B(_3961_),
    .C(_3958_),
    .A(_3938_),
    .Y(_0445_));
 sg13g2_nand3_1 _4774_ (.B(net99),
    .C(_3946_),
    .A(_3960_),
    .Y(_0446_));
 sg13g2_nand3_1 _4775_ (.B(_0446_),
    .C(_0379_),
    .A(_0445_),
    .Y(_0447_));
 sg13g2_nand2_1 _4776_ (.Y(_0448_),
    .A(_0444_),
    .B(_0447_));
 sg13g2_nor2_1 _4777_ (.A(_0016_),
    .B(net78),
    .Y(_0449_));
 sg13g2_nand2b_1 _4778_ (.Y(_0450_),
    .B(_0286_),
    .A_N(_0015_));
 sg13g2_inv_2 _4779_ (.Y(_0451_),
    .A(_0450_));
 sg13g2_a21oi_1 _4780_ (.A1(_0448_),
    .A2(_0449_),
    .Y(_0452_),
    .B1(_0451_));
 sg13g2_nand2_1 _4781_ (.Y(_0453_),
    .A(_3916_),
    .B(_0365_));
 sg13g2_nand3_1 _4782_ (.B(_3914_),
    .C(\i_transform.image_x[2] ),
    .A(_3910_),
    .Y(_0454_));
 sg13g2_nor2_1 _4783_ (.A(_0370_),
    .B(_3924_),
    .Y(_0455_));
 sg13g2_nand3_1 _4784_ (.B(_0454_),
    .C(_0455_),
    .A(_0453_),
    .Y(_0456_));
 sg13g2_nor2_1 _4785_ (.A(_0017_),
    .B(_3916_),
    .Y(_0457_));
 sg13g2_inv_1 _4786_ (.Y(_0458_),
    .A(_0457_));
 sg13g2_nand2_1 _4787_ (.Y(_0459_),
    .A(_0456_),
    .B(_0458_));
 sg13g2_xnor2_1 _4788_ (.Y(_0460_),
    .A(_0375_),
    .B(net78));
 sg13g2_nand3_1 _4789_ (.B(_0459_),
    .C(_0460_),
    .A(_0448_),
    .Y(_0461_));
 sg13g2_nand2_1 _4790_ (.Y(_0462_),
    .A(_0452_),
    .B(_0461_));
 sg13g2_nand2_1 _4791_ (.Y(_0463_),
    .A(net75),
    .B(_0354_));
 sg13g2_nand3_1 _4792_ (.B(\i_transform.image_x[5] ),
    .C(_3952_),
    .A(_3951_),
    .Y(_0464_));
 sg13g2_nor2_1 _4793_ (.A(_0358_),
    .B(net124),
    .Y(_0465_));
 sg13g2_nor2_1 _4794_ (.A(_0357_),
    .B(net99),
    .Y(_0466_));
 sg13g2_nor2_1 _4795_ (.A(_0465_),
    .B(_0466_),
    .Y(_0467_));
 sg13g2_nand3_1 _4796_ (.B(_0464_),
    .C(_0467_),
    .A(_0463_),
    .Y(_0468_));
 sg13g2_xnor2_1 _4797_ (.Y(_0469_),
    .A(_0347_),
    .B(net124));
 sg13g2_xnor2_1 _4798_ (.Y(_0470_),
    .A(_0349_),
    .B(net124));
 sg13g2_inv_1 _4799_ (.Y(_0471_),
    .A(_0470_));
 sg13g2_nor2_1 _4800_ (.A(_0469_),
    .B(_0471_),
    .Y(_0472_));
 sg13g2_nor2b_1 _4801_ (.A(_0468_),
    .B_N(_0472_),
    .Y(_0473_));
 sg13g2_nand2_1 _4802_ (.Y(_0474_),
    .A(_0462_),
    .B(_0473_));
 sg13g2_inv_1 _4803_ (.Y(_0475_),
    .A(_0375_));
 sg13g2_xnor2_1 _4804_ (.Y(_0476_),
    .A(_0475_),
    .B(net78));
 sg13g2_nand2_2 _4805_ (.Y(_0477_),
    .A(_0453_),
    .B(_0454_));
 sg13g2_inv_4 _4806_ (.A(_0477_),
    .Y(_0478_));
 sg13g2_nand2_1 _4807_ (.Y(_0479_),
    .A(_3924_),
    .B(_0370_));
 sg13g2_nor2b_1 _4808_ (.A(_0455_),
    .B_N(_0479_),
    .Y(_0480_));
 sg13g2_nand2_1 _4809_ (.Y(_0481_),
    .A(_0478_),
    .B(_0480_));
 sg13g2_nand3_1 _4810_ (.B(_3962_),
    .C(_0379_),
    .A(_3959_),
    .Y(_0482_));
 sg13g2_nand3_1 _4811_ (.B(_0446_),
    .C(_0378_),
    .A(_0445_),
    .Y(_0483_));
 sg13g2_nand2_2 _4812_ (.Y(_0484_),
    .A(_0482_),
    .B(_0483_));
 sg13g2_nor3_1 _4813_ (.A(_0476_),
    .B(_0481_),
    .C(_0484_),
    .Y(_0485_));
 sg13g2_nor2_1 _4814_ (.A(_0018_),
    .B(_3907_),
    .Y(_0486_));
 sg13g2_nand3_1 _4815_ (.B(_0473_),
    .C(_0486_),
    .A(_0485_),
    .Y(_0487_));
 sg13g2_nor2_1 _4816_ (.A(_0014_),
    .B(net75),
    .Y(_0488_));
 sg13g2_inv_1 _4817_ (.Y(_0489_),
    .A(_0488_));
 sg13g2_inv_1 _4818_ (.Y(_0490_),
    .A(_0465_));
 sg13g2_a21oi_1 _4819_ (.A1(_0489_),
    .A2(_0490_),
    .Y(_0491_),
    .B1(_0466_));
 sg13g2_nand2_1 _4820_ (.Y(_0492_),
    .A(net99),
    .B(_0349_));
 sg13g2_nand2_1 _4821_ (.Y(_0493_),
    .A(net99),
    .B(_0403_));
 sg13g2_o21ai_1 _4822_ (.B1(_0493_),
    .Y(_0494_),
    .A1(_0492_),
    .A2(_0469_));
 sg13g2_a21oi_1 _4823_ (.A1(_0491_),
    .A2(_0472_),
    .Y(_0495_),
    .B1(_0494_));
 sg13g2_nand3_1 _4824_ (.B(_0487_),
    .C(_0495_),
    .A(_0474_),
    .Y(_0496_));
 sg13g2_nand2b_1 _4825_ (.Y(_0497_),
    .B(_0496_),
    .A_N(_0443_));
 sg13g2_nand4_1 _4826_ (.B(_0487_),
    .C(_0443_),
    .A(_0474_),
    .Y(_0498_),
    .D(_0495_));
 sg13g2_nand2_1 _4827_ (.Y(_0499_),
    .A(_0497_),
    .B(_0498_));
 sg13g2_inv_1 _4828_ (.Y(_0500_),
    .A(net68));
 sg13g2_buf_1 _4829_ (.A(_0500_),
    .X(_0501_));
 sg13g2_nand2_1 _4830_ (.Y(_0502_),
    .A(_0499_),
    .B(net60));
 sg13g2_nor2_1 _4831_ (.A(_0398_),
    .B(_3907_),
    .Y(_0503_));
 sg13g2_xnor2_1 _4832_ (.Y(_0504_),
    .A(_0358_),
    .B(_3924_));
 sg13g2_nand2b_1 _4833_ (.Y(_0505_),
    .B(_0504_),
    .A_N(_0503_));
 sg13g2_nand2_1 _4834_ (.Y(_0506_),
    .A(_3924_),
    .B(_0422_));
 sg13g2_nand2_1 _4835_ (.Y(_0507_),
    .A(_0505_),
    .B(_0506_));
 sg13g2_xnor2_1 _4836_ (.Y(_0508_),
    .A(_0019_),
    .B(_3916_));
 sg13g2_nand2_1 _4837_ (.Y(_0509_),
    .A(_0507_),
    .B(_0508_));
 sg13g2_nand2_1 _4838_ (.Y(_0510_),
    .A(_3916_),
    .B(_0349_));
 sg13g2_nand2_1 _4839_ (.Y(_0511_),
    .A(_0509_),
    .B(_0510_));
 sg13g2_xnor2_1 _4840_ (.Y(_0512_),
    .A(_0417_),
    .B(_3940_));
 sg13g2_inv_1 _4841_ (.Y(_0513_),
    .A(_0512_));
 sg13g2_nand2_1 _4842_ (.Y(_0514_),
    .A(_0511_),
    .B(_0513_));
 sg13g2_nand2_1 _4843_ (.Y(_0515_),
    .A(net78),
    .B(_0403_));
 sg13g2_xnor2_1 _4844_ (.Y(_0516_),
    .A(_0435_),
    .B(_0286_));
 sg13g2_inv_2 _4845_ (.Y(_0517_),
    .A(_0516_));
 sg13g2_nand3_1 _4846_ (.B(_0515_),
    .C(_0517_),
    .A(_0514_),
    .Y(_0518_));
 sg13g2_nand2b_1 _4847_ (.Y(_0519_),
    .B(_0516_),
    .A_N(_0515_));
 sg13g2_nand3_1 _4848_ (.B(_0513_),
    .C(_0516_),
    .A(_0511_),
    .Y(_0520_));
 sg13g2_nand3_1 _4849_ (.B(_0519_),
    .C(_0520_),
    .A(_0518_),
    .Y(_0521_));
 sg13g2_a21oi_1 _4850_ (.A1(_0521_),
    .A2(net68),
    .Y(_0522_),
    .B1(net63));
 sg13g2_nand2_1 _4851_ (.Y(_0523_),
    .A(_0502_),
    .B(_0522_));
 sg13g2_nand2_1 _4852_ (.Y(_0524_),
    .A(_0442_),
    .B(_0523_));
 sg13g2_nand2_1 _4853_ (.Y(_0525_),
    .A(net71),
    .B(_0435_));
 sg13g2_nor2b_1 _4854_ (.A(_0524_),
    .B_N(_0525_),
    .Y(_0526_));
 sg13g2_nand3_1 _4855_ (.B(_0356_),
    .C(_0389_),
    .A(_0355_),
    .Y(_0527_));
 sg13g2_nor2_1 _4856_ (.A(_0014_),
    .B(net79),
    .Y(_0528_));
 sg13g2_inv_1 _4857_ (.Y(_0529_),
    .A(_0528_));
 sg13g2_nand2_1 _4858_ (.Y(_0530_),
    .A(_0527_),
    .B(_0529_));
 sg13g2_inv_1 _4859_ (.Y(_0531_),
    .A(_0361_));
 sg13g2_nor2_1 _4860_ (.A(_0351_),
    .B(_0531_),
    .Y(_0532_));
 sg13g2_nor2_1 _4861_ (.A(_0404_),
    .B(_0359_),
    .Y(_0533_));
 sg13g2_inv_1 _4862_ (.Y(_0534_),
    .A(_0533_));
 sg13g2_a21oi_1 _4863_ (.A1(_0530_),
    .A2(_0532_),
    .Y(_0535_),
    .B1(_0534_));
 sg13g2_a21oi_1 _4864_ (.A1(_0372_),
    .A2(_0364_),
    .Y(_0536_),
    .B1(_0371_));
 sg13g2_inv_1 _4865_ (.Y(_0537_),
    .A(_0536_));
 sg13g2_nand2_1 _4866_ (.Y(_0538_),
    .A(_0369_),
    .B(_0537_));
 sg13g2_nand2_2 _4867_ (.Y(_0539_),
    .A(_0538_),
    .B(_0393_));
 sg13g2_nand2_1 _4868_ (.Y(_0540_),
    .A(_0539_),
    .B(_0376_));
 sg13g2_inv_1 _4869_ (.Y(_0541_),
    .A(_0388_));
 sg13g2_nand2_1 _4870_ (.Y(_0542_),
    .A(_0540_),
    .B(_0541_));
 sg13g2_inv_1 _4871_ (.Y(_0543_),
    .A(_0532_));
 sg13g2_nand2_2 _4872_ (.Y(_0544_),
    .A(_0355_),
    .B(_0356_));
 sg13g2_nor3_1 _4873_ (.A(_0543_),
    .B(_0382_),
    .C(_0544_),
    .Y(_0545_));
 sg13g2_nand2_1 _4874_ (.Y(_0546_),
    .A(_0542_),
    .B(_0545_));
 sg13g2_nand2_1 _4875_ (.Y(_0547_),
    .A(_0535_),
    .B(_0546_));
 sg13g2_inv_1 _4876_ (.Y(_0548_),
    .A(_0348_));
 sg13g2_nand2_1 _4877_ (.Y(_0549_),
    .A(_0547_),
    .B(_0548_));
 sg13g2_nand3_1 _4878_ (.B(_0348_),
    .C(_0546_),
    .A(_0535_),
    .Y(_0550_));
 sg13g2_nand2_1 _4879_ (.Y(_0551_),
    .A(_0549_),
    .B(_0550_));
 sg13g2_nand2_1 _4880_ (.Y(_0552_),
    .A(_0551_),
    .B(net80));
 sg13g2_nand3_1 _4881_ (.B(_0418_),
    .C(_0427_),
    .A(_0426_),
    .Y(_0553_));
 sg13g2_a21oi_1 _4882_ (.A1(_0429_),
    .A2(_0553_),
    .Y(_0554_),
    .B1(net80));
 sg13g2_nand2b_1 _4883_ (.Y(_0555_),
    .B(net84),
    .A_N(_0554_));
 sg13g2_inv_1 _4884_ (.Y(_0556_),
    .A(_0555_));
 sg13g2_nand2_1 _4885_ (.Y(_0557_),
    .A(_0552_),
    .B(_0556_));
 sg13g2_nand2_1 _4886_ (.Y(_0558_),
    .A(_0490_),
    .B(_0492_));
 sg13g2_nand2_1 _4887_ (.Y(_0559_),
    .A(_0463_),
    .B(_0464_));
 sg13g2_inv_1 _4888_ (.Y(_0560_),
    .A(_0559_));
 sg13g2_nand2_1 _4889_ (.Y(_0561_),
    .A(_0560_),
    .B(_0451_));
 sg13g2_inv_1 _4890_ (.Y(_0562_),
    .A(_0467_));
 sg13g2_nor2_1 _4891_ (.A(_0471_),
    .B(_0562_),
    .Y(_0563_));
 sg13g2_inv_1 _4892_ (.Y(_0564_),
    .A(_0563_));
 sg13g2_a21oi_1 _4893_ (.A1(_0561_),
    .A2(_0489_),
    .Y(_0565_),
    .B1(_0564_));
 sg13g2_nor2_1 _4894_ (.A(_0558_),
    .B(_0565_),
    .Y(_0566_));
 sg13g2_nor2_1 _4895_ (.A(_0559_),
    .B(_0484_),
    .Y(_0567_));
 sg13g2_inv_2 _4896_ (.Y(_0568_),
    .A(_0567_));
 sg13g2_nor2_1 _4897_ (.A(_0564_),
    .B(_0568_),
    .Y(_0569_));
 sg13g2_a21oi_1 _4898_ (.A1(_0479_),
    .A2(_0486_),
    .Y(_0570_),
    .B1(_0455_));
 sg13g2_inv_1 _4899_ (.Y(_0571_),
    .A(_0570_));
 sg13g2_nand2_1 _4900_ (.Y(_0572_),
    .A(_0571_),
    .B(_0478_));
 sg13g2_nand2_1 _4901_ (.Y(_0573_),
    .A(_0572_),
    .B(_0458_));
 sg13g2_nand2_1 _4902_ (.Y(_0574_),
    .A(_0573_),
    .B(_0460_));
 sg13g2_inv_1 _4903_ (.Y(_0575_),
    .A(_0449_));
 sg13g2_nand2_1 _4904_ (.Y(_0576_),
    .A(_0574_),
    .B(_0575_));
 sg13g2_nand2_1 _4905_ (.Y(_0577_),
    .A(_0569_),
    .B(_0576_));
 sg13g2_nand2_1 _4906_ (.Y(_0578_),
    .A(_0566_),
    .B(_0577_));
 sg13g2_nand2_1 _4907_ (.Y(_0579_),
    .A(_0578_),
    .B(_0469_));
 sg13g2_inv_1 _4908_ (.Y(_0580_),
    .A(_0469_));
 sg13g2_nand3_1 _4909_ (.B(_0580_),
    .C(_0577_),
    .A(_0566_),
    .Y(_0581_));
 sg13g2_nand3_1 _4910_ (.B(_0581_),
    .C(_0500_),
    .A(_0579_),
    .Y(_0582_));
 sg13g2_xnor2_1 _4911_ (.Y(_0583_),
    .A(_0513_),
    .B(_0511_));
 sg13g2_a21oi_1 _4912_ (.A1(_0583_),
    .A2(net68),
    .Y(_0584_),
    .B1(net63));
 sg13g2_nand2_1 _4913_ (.Y(_0585_),
    .A(_0582_),
    .B(_0584_));
 sg13g2_inv_1 _4914_ (.Y(_0586_),
    .A(net71));
 sg13g2_nor2_1 _4915_ (.A(_0347_),
    .B(_0586_),
    .Y(_0587_));
 sg13g2_inv_1 _4916_ (.Y(_0588_),
    .A(_0587_));
 sg13g2_nand3_1 _4917_ (.B(_0585_),
    .C(_0588_),
    .A(_0557_),
    .Y(_0589_));
 sg13g2_buf_8 _4918_ (.A(_0589_),
    .X(_0590_));
 sg13g2_nand2_2 _4919_ (.Y(_0591_),
    .A(_0590_),
    .B(_0342_));
 sg13g2_buf_8 _4920_ (.A(_0591_),
    .X(_0592_));
 sg13g2_nor2_1 _4921_ (.A(_0526_),
    .B(net38),
    .Y(_0593_));
 sg13g2_buf_1 _4922_ (.A(_0022_),
    .X(_0594_));
 sg13g2_nor2_1 _4923_ (.A(_0594_),
    .B(_0586_),
    .Y(_0595_));
 sg13g2_o21ai_1 _4924_ (.B1(_0541_),
    .Y(_0596_),
    .A1(_0393_),
    .A2(_0377_));
 sg13g2_nor2_1 _4925_ (.A(_0382_),
    .B(_0544_),
    .Y(_0597_));
 sg13g2_nand2_1 _4926_ (.Y(_0598_),
    .A(_0596_),
    .B(_0597_));
 sg13g2_inv_1 _4927_ (.Y(_0599_),
    .A(_0530_));
 sg13g2_nand2_1 _4928_ (.Y(_0600_),
    .A(_0598_),
    .B(_0599_));
 sg13g2_nor2_1 _4929_ (.A(_0410_),
    .B(_0348_),
    .Y(_0601_));
 sg13g2_inv_1 _4930_ (.Y(_0602_),
    .A(_0601_));
 sg13g2_nor2_1 _4931_ (.A(_0602_),
    .B(_0543_),
    .Y(_0603_));
 sg13g2_nand2_1 _4932_ (.Y(_0604_),
    .A(_0600_),
    .B(_0603_));
 sg13g2_buf_1 _4933_ (.A(net126),
    .X(_0605_));
 sg13g2_nand3_1 _4934_ (.B(_0403_),
    .C(_0409_),
    .A(net114),
    .Y(_0606_));
 sg13g2_buf_2 _4935_ (.A(\i_bitmap.in[2] ),
    .X(_0607_));
 sg13g2_nand2_1 _4936_ (.Y(_0608_),
    .A(net114),
    .B(_0607_));
 sg13g2_nand2_1 _4937_ (.Y(_0609_),
    .A(_0606_),
    .B(_0608_));
 sg13g2_a21oi_1 _4938_ (.A1(_0601_),
    .A2(_0534_),
    .Y(_0610_),
    .B1(_0609_));
 sg13g2_nor2b_1 _4939_ (.A(_0377_),
    .B_N(_0369_),
    .Y(_0611_));
 sg13g2_nand4_1 _4940_ (.B(_0537_),
    .C(_0611_),
    .A(_0597_),
    .Y(_0612_),
    .D(_0603_));
 sg13g2_nand3_1 _4941_ (.B(_0610_),
    .C(_0612_),
    .A(_0604_),
    .Y(_0613_));
 sg13g2_xnor2_1 _4942_ (.Y(_0614_),
    .A(_0594_),
    .B(net133));
 sg13g2_nand2_1 _4943_ (.Y(_0615_),
    .A(_0613_),
    .B(_0614_));
 sg13g2_inv_1 _4944_ (.Y(_0616_),
    .A(_0614_));
 sg13g2_nand4_1 _4945_ (.B(_0616_),
    .C(_0610_),
    .A(_0604_),
    .Y(_0617_),
    .D(_0612_));
 sg13g2_nand3_1 _4946_ (.B(_0617_),
    .C(net80),
    .A(_0615_),
    .Y(_0618_));
 sg13g2_inv_1 _4947_ (.Y(_0619_),
    .A(_0594_));
 sg13g2_xnor2_1 _4948_ (.Y(_0620_),
    .A(_0619_),
    .B(net79));
 sg13g2_nand2_1 _4949_ (.Y(_0621_),
    .A(net72),
    .B(_0607_));
 sg13g2_nand2_1 _4950_ (.Y(_0622_),
    .A(_0438_),
    .B(_0621_));
 sg13g2_xor2_1 _4951_ (.B(_0622_),
    .A(_0620_),
    .X(_0623_));
 sg13g2_a21oi_1 _4952_ (.A1(_0623_),
    .A2(net76),
    .Y(_0624_),
    .B1(_3591_));
 sg13g2_nand2_1 _4953_ (.Y(_0625_),
    .A(_0618_),
    .B(_0624_));
 sg13g2_o21ai_1 _4954_ (.B1(_0489_),
    .Y(_0626_),
    .A1(_0450_),
    .A2(_0559_));
 sg13g2_a21oi_1 _4955_ (.A1(_0460_),
    .A2(_0457_),
    .Y(_0627_),
    .B1(_0449_));
 sg13g2_nor2_1 _4956_ (.A(_0568_),
    .B(_0627_),
    .Y(_0628_));
 sg13g2_nor2_1 _4957_ (.A(_0443_),
    .B(_0469_),
    .Y(_0629_));
 sg13g2_inv_1 _4958_ (.Y(_0630_),
    .A(_0629_));
 sg13g2_nor2_1 _4959_ (.A(_0630_),
    .B(_0564_),
    .Y(_0631_));
 sg13g2_o21ai_1 _4960_ (.B1(_0631_),
    .Y(_0632_),
    .A1(_0626_),
    .A2(_0628_));
 sg13g2_nand2_1 _4961_ (.Y(_0633_),
    .A(net99),
    .B(_0607_));
 sg13g2_o21ai_1 _4962_ (.B1(_0633_),
    .Y(_0634_),
    .A1(_0493_),
    .A2(_0443_));
 sg13g2_a21oi_1 _4963_ (.A1(_0629_),
    .A2(_0558_),
    .Y(_0635_),
    .B1(_0634_));
 sg13g2_nor2_1 _4964_ (.A(_0477_),
    .B(_0476_),
    .Y(_0636_));
 sg13g2_nand4_1 _4965_ (.B(_0636_),
    .C(_0571_),
    .A(_0567_),
    .Y(_0637_),
    .D(_0631_));
 sg13g2_nand3_1 _4966_ (.B(_0635_),
    .C(_0637_),
    .A(_0632_),
    .Y(_0638_));
 sg13g2_xnor2_1 _4967_ (.Y(_0639_),
    .A(_0594_),
    .B(net124));
 sg13g2_nand2_1 _4968_ (.Y(_0640_),
    .A(_0638_),
    .B(_0639_));
 sg13g2_inv_1 _4969_ (.Y(_0641_),
    .A(_0639_));
 sg13g2_nand4_1 _4970_ (.B(_0641_),
    .C(_0635_),
    .A(_0632_),
    .Y(_0642_),
    .D(_0637_));
 sg13g2_nand3_1 _4971_ (.B(_0642_),
    .C(net60),
    .A(_0640_),
    .Y(_0643_));
 sg13g2_nand2_1 _4972_ (.Y(_0644_),
    .A(_0291_),
    .B(_0607_));
 sg13g2_nand3_1 _4973_ (.B(_0644_),
    .C(_0519_),
    .A(_0520_),
    .Y(_0645_));
 sg13g2_xnor2_1 _4974_ (.Y(_0646_),
    .A(_0619_),
    .B(net75));
 sg13g2_nor2b_1 _4975_ (.A(_0645_),
    .B_N(_0646_),
    .Y(_0647_));
 sg13g2_nand2b_1 _4976_ (.Y(_0648_),
    .B(_0645_),
    .A_N(_0646_));
 sg13g2_nand2_1 _4977_ (.Y(_0649_),
    .A(_0648_),
    .B(_3652_));
 sg13g2_inv_1 _4978_ (.Y(_0650_),
    .A(_3671_));
 sg13g2_o21ai_1 _4979_ (.B1(_0650_),
    .Y(_0651_),
    .A1(_0647_),
    .A2(_0649_));
 sg13g2_nand2_1 _4980_ (.Y(_0652_),
    .A(_0643_),
    .B(_0651_));
 sg13g2_nand3b_1 _4981_ (.B(_0625_),
    .C(_0652_),
    .Y(_0653_),
    .A_N(_0595_));
 sg13g2_buf_2 _4982_ (.A(_0653_),
    .X(_0654_));
 sg13g2_nand2_1 _4983_ (.Y(_0655_),
    .A(_0654_),
    .B(net147));
 sg13g2_buf_8 _4984_ (.A(_0655_),
    .X(_0656_));
 sg13g2_nand3_1 _4985_ (.B(_0381_),
    .C(_0388_),
    .A(_0380_),
    .Y(_0657_));
 sg13g2_inv_1 _4986_ (.Y(_0658_),
    .A(_0389_));
 sg13g2_nand2_1 _4987_ (.Y(_0659_),
    .A(_0657_),
    .B(_0658_));
 sg13g2_nor2_1 _4988_ (.A(_0531_),
    .B(_0544_),
    .Y(_0660_));
 sg13g2_a21oi_1 _4989_ (.A1(_0659_),
    .A2(_0660_),
    .Y(_0661_),
    .B1(_0401_));
 sg13g2_nor2_1 _4990_ (.A(_0377_),
    .B(_0382_),
    .Y(_0662_));
 sg13g2_nand3_1 _4991_ (.B(_0539_),
    .C(_0662_),
    .A(_0660_),
    .Y(_0663_));
 sg13g2_nand2_1 _4992_ (.Y(_0664_),
    .A(_0661_),
    .B(_0663_));
 sg13g2_nand2_1 _4993_ (.Y(_0665_),
    .A(_0664_),
    .B(_0351_));
 sg13g2_nand3_1 _4994_ (.B(_0350_),
    .C(_0663_),
    .A(_0661_),
    .Y(_0666_));
 sg13g2_nand3_1 _4995_ (.B(_0666_),
    .C(net80),
    .A(_0665_),
    .Y(_0667_));
 sg13g2_nor2_1 _4996_ (.A(_0425_),
    .B(_0424_),
    .Y(_0668_));
 sg13g2_inv_1 _4997_ (.Y(_0669_),
    .A(_0668_));
 sg13g2_a21oi_1 _4998_ (.A1(_0669_),
    .A2(_0426_),
    .Y(_0670_),
    .B1(net80));
 sg13g2_inv_1 _4999_ (.Y(_0671_),
    .A(_0670_));
 sg13g2_nand3_1 _5000_ (.B(net84),
    .C(_0671_),
    .A(_0667_),
    .Y(_0672_));
 sg13g2_nor2_1 _5001_ (.A(_0468_),
    .B(_0452_),
    .Y(_0673_));
 sg13g2_nor2_1 _5002_ (.A(_0491_),
    .B(_0673_),
    .Y(_0674_));
 sg13g2_nor3_1 _5003_ (.A(_0476_),
    .B(_0484_),
    .C(_0468_),
    .Y(_0675_));
 sg13g2_nand2_1 _5004_ (.Y(_0676_),
    .A(_0675_),
    .B(_0573_));
 sg13g2_a21oi_1 _5005_ (.A1(_0674_),
    .A2(_0676_),
    .Y(_0677_),
    .B1(_0470_));
 sg13g2_nand3_1 _5006_ (.B(_0470_),
    .C(_0676_),
    .A(_0674_),
    .Y(_0678_));
 sg13g2_nand2_1 _5007_ (.Y(_0679_),
    .A(_0678_),
    .B(_0500_));
 sg13g2_inv_1 _5008_ (.Y(_0680_),
    .A(_0507_));
 sg13g2_nand2b_1 _5009_ (.Y(_0681_),
    .B(_0680_),
    .A_N(_0508_));
 sg13g2_nand2_1 _5010_ (.Y(_0682_),
    .A(_0681_),
    .B(_0509_));
 sg13g2_nor2_1 _5011_ (.A(_3582_),
    .B(_3588_),
    .Y(_0683_));
 sg13g2_inv_1 _5012_ (.Y(_0684_),
    .A(_0683_));
 sg13g2_nor3_1 _5013_ (.A(_0684_),
    .B(_3585_),
    .C(_3580_),
    .Y(_0685_));
 sg13g2_buf_2 _5014_ (.A(_0685_),
    .X(_0686_));
 sg13g2_inv_2 _5015_ (.Y(_0687_),
    .A(_0686_));
 sg13g2_nor2_1 _5016_ (.A(net82),
    .B(_3650_),
    .Y(_0688_));
 sg13g2_buf_2 _5017_ (.A(_0688_),
    .X(_0689_));
 sg13g2_inv_1 _5018_ (.Y(_0690_),
    .A(_0689_));
 sg13g2_a21oi_1 _5019_ (.A1(net68),
    .A2(_0682_),
    .Y(_0691_),
    .B1(_0690_));
 sg13g2_o21ai_1 _5020_ (.B1(_0691_),
    .Y(_0692_),
    .A1(_0677_),
    .A2(_0679_));
 sg13g2_nand2b_1 _5021_ (.Y(_0693_),
    .B(net71),
    .A_N(_0019_));
 sg13g2_nand3_1 _5022_ (.B(_0692_),
    .C(_0693_),
    .A(_0672_),
    .Y(_0694_));
 sg13g2_buf_1 _5023_ (.A(_0694_),
    .X(_0695_));
 sg13g2_nand3_1 _5024_ (.B(_0590_),
    .C(_0342_),
    .A(_0695_),
    .Y(_0696_));
 sg13g2_buf_2 _5025_ (.A(_0696_),
    .X(_0697_));
 sg13g2_nand3_1 _5026_ (.B(_0523_),
    .C(_0525_),
    .A(_0442_),
    .Y(_0698_));
 sg13g2_buf_1 _5027_ (.A(_0698_),
    .X(_0699_));
 sg13g2_nand2_1 _5028_ (.Y(_0700_),
    .A(_0699_),
    .B(net147));
 sg13g2_buf_8 _5029_ (.A(_0700_),
    .X(_0701_));
 sg13g2_nand2_2 _5030_ (.Y(_0702_),
    .A(_0697_),
    .B(net52));
 sg13g2_inv_2 _5031_ (.Y(_0703_),
    .A(_0702_));
 sg13g2_nor2_1 _5032_ (.A(net53),
    .B(_0703_),
    .Y(_0704_));
 sg13g2_nand2b_1 _5033_ (.Y(_0705_),
    .B(_0704_),
    .A_N(_0593_));
 sg13g2_nand2_2 _5034_ (.Y(_0706_),
    .A(_0700_),
    .B(net38));
 sg13g2_inv_2 _5035_ (.Y(_0707_),
    .A(_0706_));
 sg13g2_nand2_1 _5036_ (.Y(_0708_),
    .A(_0707_),
    .B(net53));
 sg13g2_nand2_1 _5037_ (.Y(_0709_),
    .A(_0705_),
    .B(_0708_));
 sg13g2_buf_1 _5038_ (.A(_0024_),
    .X(_0710_));
 sg13g2_nor2_1 _5039_ (.A(_0710_),
    .B(_0586_),
    .Y(_0711_));
 sg13g2_xnor2_1 _5040_ (.Y(_0712_),
    .A(_0710_),
    .B(net125));
 sg13g2_inv_1 _5041_ (.Y(_0713_),
    .A(_0712_));
 sg13g2_buf_1 _5042_ (.A(_0023_),
    .X(_0714_));
 sg13g2_xnor2_1 _5043_ (.Y(_0715_),
    .A(_0714_),
    .B(net133));
 sg13g2_nor2_1 _5044_ (.A(_0715_),
    .B(_0614_),
    .Y(_0716_));
 sg13g2_nor2b_1 _5045_ (.A(_0602_),
    .B_N(_0716_),
    .Y(_0717_));
 sg13g2_nand2b_1 _5046_ (.Y(_0718_),
    .B(_0717_),
    .A_N(_0535_));
 sg13g2_inv_1 _5047_ (.Y(_0719_),
    .A(_0714_));
 sg13g2_buf_2 _5048_ (.A(\i_bitmap.in[3] ),
    .X(_0720_));
 sg13g2_nand2_1 _5049_ (.Y(_0721_),
    .A(net114),
    .B(_0720_));
 sg13g2_buf_2 _5050_ (.A(\i_bitmap.in[4] ),
    .X(_0722_));
 sg13g2_nand2_1 _5051_ (.Y(_0723_),
    .A(net114),
    .B(_0722_));
 sg13g2_o21ai_1 _5052_ (.B1(_0723_),
    .Y(_0724_),
    .A1(_0719_),
    .A2(_0721_));
 sg13g2_a21oi_1 _5053_ (.A1(_0716_),
    .A2(_0609_),
    .Y(_0725_),
    .B1(_0724_));
 sg13g2_nand3_1 _5054_ (.B(_0545_),
    .C(_0717_),
    .A(_0542_),
    .Y(_0726_));
 sg13g2_nand3_1 _5055_ (.B(_0725_),
    .C(_0726_),
    .A(_0718_),
    .Y(_0727_));
 sg13g2_xnor2_1 _5056_ (.Y(_0728_),
    .A(_0713_),
    .B(_0727_));
 sg13g2_nand2_1 _5057_ (.Y(_0729_),
    .A(_0728_),
    .B(net77));
 sg13g2_buf_2 _5058_ (.A(\i_bitmap.in[5] ),
    .X(_0730_));
 sg13g2_xnor2_1 _5059_ (.Y(_0731_),
    .A(_0730_),
    .B(net125));
 sg13g2_o21ai_1 _5060_ (.B1(_0621_),
    .Y(_0732_),
    .A1(_0433_),
    .A2(_0436_));
 sg13g2_xnor2_1 _5061_ (.Y(_0733_),
    .A(_0722_),
    .B(net133));
 sg13g2_nor2_1 _5062_ (.A(_0733_),
    .B(_0620_),
    .Y(_0734_));
 sg13g2_inv_1 _5063_ (.Y(_0735_),
    .A(_0733_));
 sg13g2_nand3_1 _5064_ (.B(_0720_),
    .C(_0735_),
    .A(net79),
    .Y(_0736_));
 sg13g2_o21ai_1 _5065_ (.B1(_0736_),
    .Y(_0737_),
    .A1(_0714_),
    .A2(net114));
 sg13g2_a21oi_1 _5066_ (.A1(_0732_),
    .A2(_0734_),
    .Y(_0738_),
    .B1(_0737_));
 sg13g2_nor2_1 _5067_ (.A(_0418_),
    .B(_0436_),
    .Y(_0739_));
 sg13g2_nand3_1 _5068_ (.B(_0428_),
    .C(_0739_),
    .A(_0734_),
    .Y(_0740_));
 sg13g2_nand2_1 _5069_ (.Y(_0741_),
    .A(_0738_),
    .B(_0740_));
 sg13g2_xor2_1 _5070_ (.B(_0741_),
    .A(_0731_),
    .X(_0742_));
 sg13g2_a21oi_1 _5071_ (.A1(_0742_),
    .A2(net76),
    .Y(_0743_),
    .B1(_3591_));
 sg13g2_nand2_1 _5072_ (.Y(_0744_),
    .A(_0729_),
    .B(_0743_));
 sg13g2_xnor2_1 _5073_ (.Y(_0745_),
    .A(_0710_),
    .B(net115));
 sg13g2_xnor2_1 _5074_ (.Y(_0746_),
    .A(_0714_),
    .B(net124));
 sg13g2_nor2_1 _5075_ (.A(_0746_),
    .B(_0639_),
    .Y(_0747_));
 sg13g2_nor2b_1 _5076_ (.A(_0630_),
    .B_N(_0747_),
    .Y(_0748_));
 sg13g2_o21ai_1 _5077_ (.B1(_0748_),
    .Y(_0749_),
    .A1(_0558_),
    .A2(_0565_));
 sg13g2_buf_1 _5078_ (.A(_3950_),
    .X(_0750_));
 sg13g2_nand2_1 _5079_ (.Y(_0751_),
    .A(_3950_),
    .B(_0720_));
 sg13g2_nor2_1 _5080_ (.A(_0751_),
    .B(_0746_),
    .Y(_0752_));
 sg13g2_a221oi_1 _5081_ (.B2(_0747_),
    .C1(_0752_),
    .B1(_0634_),
    .A1(_0722_),
    .Y(_0753_),
    .A2(net92));
 sg13g2_nand3_1 _5082_ (.B(_0576_),
    .C(_0748_),
    .A(_0569_),
    .Y(_0754_));
 sg13g2_nand3_1 _5083_ (.B(_0753_),
    .C(_0754_),
    .A(_0749_),
    .Y(_0755_));
 sg13g2_xnor2_1 _5084_ (.Y(_0756_),
    .A(_0745_),
    .B(_0755_));
 sg13g2_xnor2_1 _5085_ (.Y(_0757_),
    .A(_0730_),
    .B(net115));
 sg13g2_nand2_1 _5086_ (.Y(_0758_),
    .A(_0519_),
    .B(_0644_));
 sg13g2_xnor2_1 _5087_ (.Y(_0759_),
    .A(_0722_),
    .B(net115));
 sg13g2_nor2_1 _5088_ (.A(_0759_),
    .B(_0646_),
    .Y(_0760_));
 sg13g2_nand2_1 _5089_ (.Y(_0761_),
    .A(net75),
    .B(_0720_));
 sg13g2_nand2_1 _5090_ (.Y(_0762_),
    .A(net115),
    .B(_0719_));
 sg13g2_o21ai_1 _5091_ (.B1(_0762_),
    .Y(_0763_),
    .A1(_0759_),
    .A2(_0761_));
 sg13g2_a21oi_1 _5092_ (.A1(_0758_),
    .A2(_0760_),
    .Y(_0764_),
    .B1(_0763_));
 sg13g2_nand4_1 _5093_ (.B(_0760_),
    .C(_0513_),
    .A(_0511_),
    .Y(_0765_),
    .D(_0516_));
 sg13g2_nand2_1 _5094_ (.Y(_0766_),
    .A(_0764_),
    .B(_0765_));
 sg13g2_xor2_1 _5095_ (.B(_0766_),
    .A(_0757_),
    .X(_0767_));
 sg13g2_a21oi_1 _5096_ (.A1(_0767_),
    .A2(net68),
    .Y(_0768_),
    .B1(_0690_));
 sg13g2_o21ai_1 _5097_ (.B1(_0768_),
    .Y(_0769_),
    .A1(net62),
    .A2(_0756_));
 sg13g2_nand3b_1 _5098_ (.B(_0744_),
    .C(_0769_),
    .Y(_0770_),
    .A_N(_0711_));
 sg13g2_buf_2 _5099_ (.A(_0770_),
    .X(_0771_));
 sg13g2_nor2_1 _5100_ (.A(_0614_),
    .B(_0410_),
    .Y(_0772_));
 sg13g2_inv_1 _5101_ (.Y(_0773_),
    .A(_0772_));
 sg13g2_nor2_1 _5102_ (.A(_0773_),
    .B(_0353_),
    .Y(_0774_));
 sg13g2_nand2b_1 _5103_ (.Y(_0775_),
    .B(_0774_),
    .A_N(_0661_));
 sg13g2_inv_1 _5104_ (.Y(_0776_),
    .A(_0405_));
 sg13g2_o21ai_1 _5105_ (.B1(_0721_),
    .Y(_0777_),
    .A1(_0619_),
    .A2(_0608_));
 sg13g2_a21oi_1 _5106_ (.A1(_0776_),
    .A2(_0772_),
    .Y(_0778_),
    .B1(_0777_));
 sg13g2_nand4_1 _5107_ (.B(_0539_),
    .C(_0662_),
    .A(_0660_),
    .Y(_0779_),
    .D(_0774_));
 sg13g2_nand3_1 _5108_ (.B(_0778_),
    .C(_0779_),
    .A(_0775_),
    .Y(_0780_));
 sg13g2_xor2_1 _5109_ (.B(_0780_),
    .A(_0715_),
    .X(_0781_));
 sg13g2_nand2_1 _5110_ (.Y(_0782_),
    .A(_0781_),
    .B(net80));
 sg13g2_o21ai_1 _5111_ (.B1(_0433_),
    .Y(_0783_),
    .A1(_0427_),
    .A2(_0418_));
 sg13g2_nor2_1 _5112_ (.A(_0436_),
    .B(_0620_),
    .Y(_0784_));
 sg13g2_nand2_1 _5113_ (.Y(_0785_),
    .A(net79),
    .B(_0720_));
 sg13g2_o21ai_1 _5114_ (.B1(_0785_),
    .Y(_0786_),
    .A1(_0621_),
    .A2(_0620_));
 sg13g2_a21oi_1 _5115_ (.A1(_0783_),
    .A2(_0784_),
    .Y(_0787_),
    .B1(_0786_));
 sg13g2_nor2b_1 _5116_ (.A(_0418_),
    .B_N(_0425_),
    .Y(_0788_));
 sg13g2_nand3_1 _5117_ (.B(_0424_),
    .C(_0788_),
    .A(_0784_),
    .Y(_0789_));
 sg13g2_nand2_1 _5118_ (.Y(_0790_),
    .A(_0787_),
    .B(_0789_));
 sg13g2_xnor2_1 _5119_ (.Y(_0791_),
    .A(_0735_),
    .B(_0790_));
 sg13g2_a21oi_1 _5120_ (.A1(_0791_),
    .A2(net76),
    .Y(_0792_),
    .B1(_3591_));
 sg13g2_nand2_1 _5121_ (.Y(_0793_),
    .A(_0782_),
    .B(_0792_));
 sg13g2_nor2_1 _5122_ (.A(_0646_),
    .B(_0517_),
    .Y(_0794_));
 sg13g2_nand3_1 _5123_ (.B(_0513_),
    .C(_0508_),
    .A(_0794_),
    .Y(_0795_));
 sg13g2_o21ai_1 _5124_ (.B1(_0515_),
    .Y(_0796_),
    .A1(_0510_),
    .A2(_0512_));
 sg13g2_o21ai_1 _5125_ (.B1(_0761_),
    .Y(_0797_),
    .A1(_0644_),
    .A2(_0646_));
 sg13g2_a21oi_1 _5126_ (.A1(_0796_),
    .A2(_0794_),
    .Y(_0798_),
    .B1(_0797_));
 sg13g2_o21ai_1 _5127_ (.B1(_0798_),
    .Y(_0799_),
    .A1(_0680_),
    .A2(_0795_));
 sg13g2_xor2_1 _5128_ (.B(_0799_),
    .A(_0759_),
    .X(_0800_));
 sg13g2_a21oi_1 _5129_ (.A1(_0800_),
    .A2(net68),
    .Y(_0801_),
    .B1(net63));
 sg13g2_nor2_1 _5130_ (.A(_0639_),
    .B(_0443_),
    .Y(_0802_));
 sg13g2_and2_1 _5131_ (.A(_0472_),
    .B(_0802_),
    .X(_0803_));
 sg13g2_o21ai_1 _5132_ (.B1(_0803_),
    .Y(_0804_),
    .A1(_0491_),
    .A2(_0673_));
 sg13g2_o21ai_1 _5133_ (.B1(_0751_),
    .Y(_0805_),
    .A1(_0633_),
    .A2(_0639_));
 sg13g2_a21oi_1 _5134_ (.A1(_0494_),
    .A2(_0802_),
    .Y(_0806_),
    .B1(_0805_));
 sg13g2_nand3_1 _5135_ (.B(_0573_),
    .C(_0803_),
    .A(_0675_),
    .Y(_0807_));
 sg13g2_nand3_1 _5136_ (.B(_0806_),
    .C(_0807_),
    .A(_0804_),
    .Y(_0808_));
 sg13g2_nand2_1 _5137_ (.Y(_0809_),
    .A(_0808_),
    .B(_0746_));
 sg13g2_inv_1 _5138_ (.Y(_0810_),
    .A(_0746_));
 sg13g2_nand4_1 _5139_ (.B(_0810_),
    .C(_0806_),
    .A(_0804_),
    .Y(_0811_),
    .D(_0807_));
 sg13g2_nand3_1 _5140_ (.B(_0811_),
    .C(net60),
    .A(_0809_),
    .Y(_0812_));
 sg13g2_nand2_1 _5141_ (.Y(_0813_),
    .A(_0801_),
    .B(_0812_));
 sg13g2_nand2_1 _5142_ (.Y(_0814_),
    .A(net71),
    .B(_0719_));
 sg13g2_nand3_1 _5143_ (.B(_0813_),
    .C(_0814_),
    .A(_0793_),
    .Y(_0815_));
 sg13g2_buf_2 _5144_ (.A(_0815_),
    .X(_0816_));
 sg13g2_nand2_1 _5145_ (.Y(_0817_),
    .A(_0816_),
    .B(net147));
 sg13g2_buf_8 _5146_ (.A(_0817_),
    .X(_0818_));
 sg13g2_buf_8 _5147_ (.A(_0818_),
    .X(_0819_));
 sg13g2_nor2_2 _5148_ (.A(_0771_),
    .B(net51),
    .Y(_0820_));
 sg13g2_nand2_1 _5149_ (.Y(_0821_),
    .A(_0709_),
    .B(_0820_));
 sg13g2_nor2_1 _5150_ (.A(net54),
    .B(_0821_),
    .Y(_0822_));
 sg13g2_nand2_2 _5151_ (.Y(_0823_),
    .A(_0695_),
    .B(_0342_));
 sg13g2_nand2_1 _5152_ (.Y(_0824_),
    .A(_0823_),
    .B(_0591_));
 sg13g2_buf_8 _5153_ (.A(_0824_),
    .X(_0825_));
 sg13g2_nand2_2 _5154_ (.Y(_0826_),
    .A(_0825_),
    .B(_0697_));
 sg13g2_nand2_1 _5155_ (.Y(_0827_),
    .A(_0625_),
    .B(_0652_));
 sg13g2_nor2_2 _5156_ (.A(_0595_),
    .B(_0827_),
    .Y(_0828_));
 sg13g2_nor2_2 _5157_ (.A(_0592_),
    .B(_0828_),
    .Y(_0829_));
 sg13g2_a21oi_1 _5158_ (.A1(_0826_),
    .A2(net53),
    .Y(_0830_),
    .B1(_0829_));
 sg13g2_nand2_1 _5159_ (.Y(_0831_),
    .A(_0771_),
    .B(net147));
 sg13g2_buf_8 _5160_ (.A(_0831_),
    .X(_0832_));
 sg13g2_inv_4 _5161_ (.A(net48),
    .Y(_0833_));
 sg13g2_buf_1 _5162_ (.A(_0833_),
    .X(_0834_));
 sg13g2_inv_8 _5163_ (.Y(_0835_),
    .A(_0818_));
 sg13g2_buf_8 _5164_ (.A(_0835_),
    .X(_0836_));
 sg13g2_nand3_1 _5165_ (.B(_0834_),
    .C(_0836_),
    .A(_0830_),
    .Y(_0837_));
 sg13g2_inv_2 _5166_ (.Y(_0838_),
    .A(_0343_));
 sg13g2_buf_1 _5167_ (.A(_0034_),
    .X(_0839_));
 sg13g2_nor2_1 _5168_ (.A(_0839_),
    .B(_0586_),
    .Y(_0840_));
 sg13g2_nor2_1 _5169_ (.A(net83),
    .B(_0332_),
    .Y(_0841_));
 sg13g2_inv_1 _5170_ (.Y(_0842_),
    .A(_0841_));
 sg13g2_buf_2 _5171_ (.A(\i_bitmap.in[8] ),
    .X(_0843_));
 sg13g2_xnor2_1 _5172_ (.Y(_0844_),
    .A(_0843_),
    .B(net78));
 sg13g2_inv_1 _5173_ (.Y(_0845_),
    .A(_0844_));
 sg13g2_a21oi_1 _5174_ (.A1(_0338_),
    .A2(_3917_),
    .Y(_0846_),
    .B1(_0331_));
 sg13g2_nor2_1 _5175_ (.A(_0845_),
    .B(_0846_),
    .Y(_0847_));
 sg13g2_a21oi_1 _5176_ (.A1(_0846_),
    .A2(_0845_),
    .Y(_0848_),
    .B1(_0686_));
 sg13g2_nand2b_1 _5177_ (.Y(_0849_),
    .B(_0848_),
    .A_N(_0847_));
 sg13g2_xnor2_1 _5178_ (.Y(_0850_),
    .A(_0843_),
    .B(net100));
 sg13g2_inv_1 _5179_ (.Y(_0851_),
    .A(_0850_));
 sg13g2_nand2_1 _5180_ (.Y(_0852_),
    .A(_0298_),
    .B(_3898_));
 sg13g2_o21ai_1 _5181_ (.B1(_0852_),
    .Y(_0853_),
    .A1(_3777_),
    .A2(net92));
 sg13g2_xnor2_1 _5182_ (.Y(_0854_),
    .A(_0851_),
    .B(_0853_));
 sg13g2_a22oi_1 _5183_ (.Y(_0855_),
    .B1(net77),
    .B2(_0854_),
    .A2(_0849_),
    .A1(_0842_));
 sg13g2_buf_1 _5184_ (.A(net125),
    .X(_0856_));
 sg13g2_xnor2_1 _5185_ (.Y(_0857_),
    .A(_0839_),
    .B(net113));
 sg13g2_inv_1 _5186_ (.Y(_0858_),
    .A(_0857_));
 sg13g2_nor2_1 _5187_ (.A(_3816_),
    .B(_3854_),
    .Y(_0859_));
 sg13g2_inv_1 _5188_ (.Y(_0860_),
    .A(_0859_));
 sg13g2_inv_1 _5189_ (.Y(_0861_),
    .A(_3872_));
 sg13g2_nor2_1 _5190_ (.A(_0861_),
    .B(_3827_),
    .Y(_0862_));
 sg13g2_nor2_1 _5191_ (.A(_3875_),
    .B(_0862_),
    .Y(_0863_));
 sg13g2_nor2_1 _5192_ (.A(_3853_),
    .B(_0863_),
    .Y(_0864_));
 sg13g2_nor2_1 _5193_ (.A(_3874_),
    .B(_0864_),
    .Y(_0865_));
 sg13g2_inv_1 _5194_ (.Y(_0866_),
    .A(_0865_));
 sg13g2_a21oi_1 _5195_ (.A1(_0866_),
    .A2(_3862_),
    .Y(_0867_),
    .B1(_3878_));
 sg13g2_nor2_1 _5196_ (.A(_3890_),
    .B(net113),
    .Y(_0868_));
 sg13g2_a21oi_1 _5197_ (.A1(_3881_),
    .A2(_3777_),
    .Y(_0869_),
    .B1(_0868_));
 sg13g2_o21ai_1 _5198_ (.B1(_0869_),
    .Y(_0870_),
    .A1(_0860_),
    .A2(_0867_));
 sg13g2_xnor2_1 _5199_ (.Y(_0871_),
    .A(_0858_),
    .B(_0870_));
 sg13g2_a21oi_1 _5200_ (.A1(_3889_),
    .A2(_3809_),
    .Y(_0872_),
    .B1(_3811_));
 sg13g2_xnor2_1 _5201_ (.Y(_0873_),
    .A(_0839_),
    .B(_3871_));
 sg13g2_inv_1 _5202_ (.Y(_0874_),
    .A(_0873_));
 sg13g2_a21oi_1 _5203_ (.A1(_0872_),
    .A2(_0874_),
    .Y(_0875_),
    .B1(_0690_));
 sg13g2_nor2_1 _5204_ (.A(_0874_),
    .B(_0872_),
    .Y(_0876_));
 sg13g2_inv_1 _5205_ (.Y(_0877_),
    .A(_0876_));
 sg13g2_nor2_1 _5206_ (.A(_0690_),
    .B(net68),
    .Y(_0878_));
 sg13g2_a21oi_1 _5207_ (.A1(_0875_),
    .A2(_0877_),
    .Y(_0879_),
    .B1(_0878_));
 sg13g2_a21oi_1 _5208_ (.A1(_0871_),
    .A2(net60),
    .Y(_0880_),
    .B1(_0879_));
 sg13g2_nor3_1 _5209_ (.A(_0840_),
    .B(_0855_),
    .C(_0880_),
    .Y(_0881_));
 sg13g2_nor2_1 _5210_ (.A(_0838_),
    .B(_0881_),
    .Y(_0882_));
 sg13g2_buf_2 _5211_ (.A(_0882_),
    .X(_0883_));
 sg13g2_buf_8 _5212_ (.A(net48),
    .X(_0884_));
 sg13g2_inv_2 _5213_ (.Y(_0885_),
    .A(_0816_));
 sg13g2_nor2_1 _5214_ (.A(net38),
    .B(_0823_),
    .Y(_0886_));
 sg13g2_buf_8 _5215_ (.A(_0886_),
    .X(_0887_));
 sg13g2_nor2_2 _5216_ (.A(_0701_),
    .B(_0828_),
    .Y(_0888_));
 sg13g2_nand4_1 _5217_ (.B(_0885_),
    .C(_0887_),
    .A(net37),
    .Y(_0889_),
    .D(_0888_));
 sg13g2_nand3_1 _5218_ (.B(_0883_),
    .C(_0889_),
    .A(_0837_),
    .Y(_0890_));
 sg13g2_nor2_1 _5219_ (.A(_0822_),
    .B(_0890_),
    .Y(_0891_));
 sg13g2_nor2b_1 _5220_ (.A(_0526_),
    .B_N(net147),
    .Y(_0892_));
 sg13g2_buf_2 _5221_ (.A(_0892_),
    .X(_0893_));
 sg13g2_nor2_1 _5222_ (.A(_0893_),
    .B(_0825_),
    .Y(_0894_));
 sg13g2_inv_1 _5223_ (.Y(_0895_),
    .A(_0894_));
 sg13g2_nand2_1 _5224_ (.Y(_0896_),
    .A(_0825_),
    .B(_0893_));
 sg13g2_buf_8 _5225_ (.A(_0896_),
    .X(_0897_));
 sg13g2_nand2_1 _5226_ (.Y(_0898_),
    .A(_0895_),
    .B(_0897_));
 sg13g2_nand2_1 _5227_ (.Y(_0899_),
    .A(_0898_),
    .B(net53));
 sg13g2_nand2_1 _5228_ (.Y(_0900_),
    .A(_0899_),
    .B(_0705_));
 sg13g2_nand2_1 _5229_ (.Y(_0901_),
    .A(_0900_),
    .B(_0820_));
 sg13g2_nand3_1 _5230_ (.B(_0702_),
    .C(_0656_),
    .A(_0897_),
    .Y(_0902_));
 sg13g2_nand2_1 _5231_ (.Y(_0903_),
    .A(_0829_),
    .B(_0885_));
 sg13g2_nand2_1 _5232_ (.Y(_0904_),
    .A(_0902_),
    .B(_0903_));
 sg13g2_nor2_1 _5233_ (.A(_0816_),
    .B(_0832_),
    .Y(_0905_));
 sg13g2_nand2_1 _5234_ (.Y(_0906_),
    .A(_0904_),
    .B(_0905_));
 sg13g2_nand2_1 _5235_ (.Y(_0907_),
    .A(_0901_),
    .B(_0906_));
 sg13g2_nand2_1 _5236_ (.Y(_0908_),
    .A(_0907_),
    .B(_0346_));
 sg13g2_nand3_1 _5237_ (.B(_0656_),
    .C(_0706_),
    .A(_0897_),
    .Y(_0909_));
 sg13g2_nand2_1 _5238_ (.Y(_0910_),
    .A(_0909_),
    .B(_0903_));
 sg13g2_buf_1 _5239_ (.A(net32),
    .X(_0911_));
 sg13g2_nand2_2 _5240_ (.Y(_0912_),
    .A(_0344_),
    .B(_0819_));
 sg13g2_inv_2 _5241_ (.Y(_0913_),
    .A(_0912_));
 sg13g2_nand3_1 _5242_ (.B(net27),
    .C(_0913_),
    .A(_0910_),
    .Y(_0914_));
 sg13g2_nand3_1 _5243_ (.B(_0908_),
    .C(_0914_),
    .A(_0891_),
    .Y(_0915_));
 sg13g2_nor2_1 _5244_ (.A(_0838_),
    .B(_0828_),
    .Y(_0916_));
 sg13g2_buf_2 _5245_ (.A(_0916_),
    .X(_0917_));
 sg13g2_nor2_1 _5246_ (.A(net50),
    .B(_0702_),
    .Y(_0918_));
 sg13g2_inv_1 _5247_ (.Y(_0919_),
    .A(_0918_));
 sg13g2_nand2_1 _5248_ (.Y(_0920_),
    .A(_0705_),
    .B(_0919_));
 sg13g2_a21oi_1 _5249_ (.A1(_0920_),
    .A2(_0820_),
    .Y(_0921_),
    .B1(_0345_));
 sg13g2_nor2_1 _5250_ (.A(_0818_),
    .B(_0830_),
    .Y(_0922_));
 sg13g2_nor2_1 _5251_ (.A(net48),
    .B(_0922_),
    .Y(_0923_));
 sg13g2_nand2_2 _5252_ (.Y(_0924_),
    .A(_0825_),
    .B(net52));
 sg13g2_nor2_1 _5253_ (.A(_0917_),
    .B(_0924_),
    .Y(_0925_));
 sg13g2_nor2_1 _5254_ (.A(_0835_),
    .B(_0925_),
    .Y(_0926_));
 sg13g2_nor2_1 _5255_ (.A(_0699_),
    .B(_0591_),
    .Y(_0927_));
 sg13g2_buf_2 _5256_ (.A(_0927_),
    .X(_0928_));
 sg13g2_nand2_1 _5257_ (.Y(_0929_),
    .A(_0928_),
    .B(_0654_));
 sg13g2_nand2_1 _5258_ (.Y(_0930_),
    .A(_0926_),
    .B(_0929_));
 sg13g2_nand2_1 _5259_ (.Y(_0931_),
    .A(_0923_),
    .B(_0930_));
 sg13g2_nand2_1 _5260_ (.Y(_0932_),
    .A(_0921_),
    .B(_0931_));
 sg13g2_inv_1 _5261_ (.Y(_0933_),
    .A(_0928_));
 sg13g2_nor2_1 _5262_ (.A(_0816_),
    .B(_0933_),
    .Y(_0934_));
 sg13g2_buf_1 _5263_ (.A(_0344_),
    .X(_0935_));
 sg13g2_a21oi_1 _5264_ (.A1(_0834_),
    .A2(_0934_),
    .Y(_0936_),
    .B1(net55));
 sg13g2_nand3_1 _5265_ (.B(_0837_),
    .C(_0936_),
    .A(_0821_),
    .Y(_0937_));
 sg13g2_nand2_1 _5266_ (.Y(_0938_),
    .A(_0932_),
    .B(_0937_));
 sg13g2_inv_4 _5267_ (.A(_0883_),
    .Y(_0939_));
 sg13g2_nand2_1 _5268_ (.Y(_0940_),
    .A(_0938_),
    .B(net46));
 sg13g2_nand2_1 _5269_ (.Y(_0941_),
    .A(_0915_),
    .B(_0940_));
 sg13g2_buf_1 _5270_ (.A(_0025_),
    .X(_0942_));
 sg13g2_xnor2_1 _5271_ (.Y(_0943_),
    .A(_0942_),
    .B(net115));
 sg13g2_inv_1 _5272_ (.Y(_0944_),
    .A(_0745_));
 sg13g2_nand2_1 _5273_ (.Y(_0945_),
    .A(_0755_),
    .B(_0944_));
 sg13g2_nand2_1 _5274_ (.Y(_0946_),
    .A(net92),
    .B(_0730_));
 sg13g2_nand3b_1 _5275_ (.B(_0945_),
    .C(_0946_),
    .Y(_0947_),
    .A_N(_0943_));
 sg13g2_nand2_1 _5276_ (.Y(_0948_),
    .A(_0945_),
    .B(_0946_));
 sg13g2_nand2_1 _5277_ (.Y(_0949_),
    .A(_0948_),
    .B(_0943_));
 sg13g2_nand3_1 _5278_ (.B(_0949_),
    .C(_0501_),
    .A(_0947_),
    .Y(_0950_));
 sg13g2_nand2b_1 _5279_ (.Y(_0951_),
    .B(_0766_),
    .A_N(_0757_));
 sg13g2_inv_1 _5280_ (.Y(_0952_),
    .A(_0710_));
 sg13g2_nand2_1 _5281_ (.Y(_0953_),
    .A(_3896_),
    .B(_0952_));
 sg13g2_buf_2 _5282_ (.A(\i_bitmap.in[6] ),
    .X(_0954_));
 sg13g2_xnor2_1 _5283_ (.Y(_0955_),
    .A(_0954_),
    .B(_3896_));
 sg13g2_a21o_1 _5284_ (.A2(_0953_),
    .A1(_0951_),
    .B1(_0955_),
    .X(_0956_));
 sg13g2_nand3_1 _5285_ (.B(_0953_),
    .C(_0955_),
    .A(_0951_),
    .Y(_0957_));
 sg13g2_nand3_1 _5286_ (.B(_0689_),
    .C(_0957_),
    .A(_0956_),
    .Y(_0958_));
 sg13g2_inv_1 _5287_ (.Y(_0959_),
    .A(_0878_));
 sg13g2_nand2_1 _5288_ (.Y(_0960_),
    .A(_0958_),
    .B(_0959_));
 sg13g2_nand2_1 _5289_ (.Y(_0961_),
    .A(_0950_),
    .B(_0960_));
 sg13g2_nand2b_1 _5290_ (.Y(_0962_),
    .B(_0741_),
    .A_N(_0731_));
 sg13g2_nand2_1 _5291_ (.Y(_0963_),
    .A(net125),
    .B(_0952_));
 sg13g2_xnor2_1 _5292_ (.Y(_0964_),
    .A(_0954_),
    .B(net125));
 sg13g2_a21oi_1 _5293_ (.A1(_0962_),
    .A2(_0963_),
    .Y(_0965_),
    .B1(_0964_));
 sg13g2_inv_1 _5294_ (.Y(_0966_),
    .A(_0965_));
 sg13g2_nand3_1 _5295_ (.B(_0963_),
    .C(_0964_),
    .A(_0962_),
    .Y(_0967_));
 sg13g2_nand2_1 _5296_ (.Y(_0968_),
    .A(_0966_),
    .B(_0967_));
 sg13g2_a21oi_1 _5297_ (.A1(_0968_),
    .A2(net76),
    .Y(_0969_),
    .B1(_3591_));
 sg13g2_xnor2_1 _5298_ (.Y(_0970_),
    .A(_0942_),
    .B(_3815_));
 sg13g2_inv_1 _5299_ (.Y(_0971_),
    .A(_0970_));
 sg13g2_nor2_1 _5300_ (.A(_0712_),
    .B(_0715_),
    .Y(_0972_));
 sg13g2_nor2b_1 _5301_ (.A(_0773_),
    .B_N(_0972_),
    .Y(_0973_));
 sg13g2_inv_1 _5302_ (.Y(_0974_),
    .A(_0730_));
 sg13g2_nor2_1 _5303_ (.A(_0974_),
    .B(_3815_),
    .Y(_0975_));
 sg13g2_inv_1 _5304_ (.Y(_0976_),
    .A(_0975_));
 sg13g2_o21ai_1 _5305_ (.B1(_0976_),
    .Y(_0977_),
    .A1(_0952_),
    .A2(_0723_));
 sg13g2_a221oi_1 _5306_ (.B2(_0973_),
    .C1(_0977_),
    .B1(_0406_),
    .A1(_0777_),
    .Y(_0978_),
    .A2(_0972_));
 sg13g2_nand2_1 _5307_ (.Y(_0979_),
    .A(_0542_),
    .B(_0387_));
 sg13g2_nand2_1 _5308_ (.Y(_0980_),
    .A(_0979_),
    .B(_0658_));
 sg13g2_nand3_1 _5309_ (.B(_0363_),
    .C(_0973_),
    .A(_0980_),
    .Y(_0981_));
 sg13g2_nand2_1 _5310_ (.Y(_0982_),
    .A(_0978_),
    .B(_0981_));
 sg13g2_xnor2_1 _5311_ (.Y(_0983_),
    .A(_0971_),
    .B(_0982_));
 sg13g2_nand2_1 _5312_ (.Y(_0984_),
    .A(_0983_),
    .B(net77));
 sg13g2_nand2_1 _5313_ (.Y(_0985_),
    .A(_0969_),
    .B(_0984_));
 sg13g2_inv_1 _5314_ (.Y(_0986_),
    .A(_0942_));
 sg13g2_nand3_1 _5315_ (.B(_0986_),
    .C(_0686_),
    .A(_3650_),
    .Y(_0987_));
 sg13g2_nand3_1 _5316_ (.B(_0985_),
    .C(_0987_),
    .A(_0961_),
    .Y(_0988_));
 sg13g2_buf_2 _5317_ (.A(_0988_),
    .X(_0989_));
 sg13g2_nand2_1 _5318_ (.Y(_0990_),
    .A(_0989_),
    .B(net147));
 sg13g2_buf_1 _5319_ (.A(_0990_),
    .X(_0991_));
 sg13g2_inv_4 _5320_ (.A(net31),
    .Y(_0992_));
 sg13g2_buf_8 _5321_ (.A(_0992_),
    .X(_0993_));
 sg13g2_nand2_1 _5322_ (.Y(_0994_),
    .A(_0941_),
    .B(net25));
 sg13g2_nand2_1 _5323_ (.Y(_0995_),
    .A(_0887_),
    .B(_0893_));
 sg13g2_buf_8 _5324_ (.A(_0995_),
    .X(_0996_));
 sg13g2_buf_8 _5325_ (.A(net50),
    .X(_0997_));
 sg13g2_nand3_1 _5326_ (.B(_0997_),
    .C(_0706_),
    .A(_0996_),
    .Y(_0998_));
 sg13g2_nor2_1 _5327_ (.A(_0695_),
    .B(net38),
    .Y(_0999_));
 sg13g2_buf_2 _5328_ (.A(_0999_),
    .X(_1000_));
 sg13g2_nand2_1 _5329_ (.Y(_1001_),
    .A(_1000_),
    .B(net52));
 sg13g2_buf_8 _5330_ (.A(net53),
    .X(_1002_));
 sg13g2_nand2_1 _5331_ (.Y(_1003_),
    .A(_1001_),
    .B(_1002_));
 sg13g2_a21oi_1 _5332_ (.A1(_0998_),
    .A2(_1003_),
    .Y(_1004_),
    .B1(_0912_));
 sg13g2_nor2_2 _5333_ (.A(_0590_),
    .B(_0823_),
    .Y(_1005_));
 sg13g2_nand2_1 _5334_ (.Y(_1006_),
    .A(_1005_),
    .B(net52));
 sg13g2_buf_1 _5335_ (.A(net50),
    .X(_1007_));
 sg13g2_nand3_1 _5336_ (.B(_1006_),
    .C(net43),
    .A(_0996_),
    .Y(_1008_));
 sg13g2_nor2_1 _5337_ (.A(_0835_),
    .B(_0344_),
    .Y(_1009_));
 sg13g2_inv_1 _5338_ (.Y(_1010_),
    .A(_1009_));
 sg13g2_a21oi_1 _5339_ (.A1(_1008_),
    .A2(_1003_),
    .Y(_1011_),
    .B1(_1010_));
 sg13g2_o21ai_1 _5340_ (.B1(net46),
    .Y(_1012_),
    .A1(_1004_),
    .A2(_1011_));
 sg13g2_buf_8 _5341_ (.A(_0818_),
    .X(_1013_));
 sg13g2_buf_8 _5342_ (.A(_0893_),
    .X(_1014_));
 sg13g2_nand2_1 _5343_ (.Y(_1015_),
    .A(_0826_),
    .B(_1014_));
 sg13g2_nor2_1 _5344_ (.A(_0928_),
    .B(net53),
    .Y(_1016_));
 sg13g2_inv_1 _5345_ (.Y(_1017_),
    .A(_0902_));
 sg13g2_a21oi_1 _5346_ (.A1(_1015_),
    .A2(_1016_),
    .Y(_1018_),
    .B1(_1017_));
 sg13g2_nor2_1 _5347_ (.A(net49),
    .B(_1018_),
    .Y(_1019_));
 sg13g2_inv_1 _5348_ (.Y(_1020_),
    .A(_1019_));
 sg13g2_buf_8 _5349_ (.A(net53),
    .X(_1021_));
 sg13g2_buf_1 _5350_ (.A(net41),
    .X(_1022_));
 sg13g2_o21ai_1 _5351_ (.B1(net52),
    .Y(_1023_),
    .A1(_0590_),
    .A2(_0823_));
 sg13g2_nand3_1 _5352_ (.B(_0697_),
    .C(net42),
    .A(_0825_),
    .Y(_1024_));
 sg13g2_nor3_1 _5353_ (.A(_0695_),
    .B(_0699_),
    .C(net38),
    .Y(_1025_));
 sg13g2_nor2_1 _5354_ (.A(net50),
    .B(_1025_),
    .Y(_1026_));
 sg13g2_nand2_1 _5355_ (.Y(_1027_),
    .A(_1024_),
    .B(_1026_));
 sg13g2_o21ai_1 _5356_ (.B1(_1027_),
    .Y(_1028_),
    .A1(net36),
    .A2(_1023_));
 sg13g2_buf_1 _5357_ (.A(net49),
    .X(_1029_));
 sg13g2_nand3_1 _5358_ (.B(_1028_),
    .C(_1029_),
    .A(_0883_),
    .Y(_1030_));
 sg13g2_nand3_1 _5359_ (.B(_1020_),
    .C(_1030_),
    .A(_1012_),
    .Y(_1031_));
 sg13g2_buf_1 _5360_ (.A(net37),
    .X(_1032_));
 sg13g2_nand2_1 _5361_ (.Y(_1033_),
    .A(_1031_),
    .B(net30));
 sg13g2_nand3_1 _5362_ (.B(_0697_),
    .C(_0526_),
    .A(_0825_),
    .Y(_1034_));
 sg13g2_buf_1 _5363_ (.A(_1034_),
    .X(_1035_));
 sg13g2_nand2_1 _5364_ (.Y(_1036_),
    .A(net42),
    .B(net38));
 sg13g2_buf_2 _5365_ (.A(_1036_),
    .X(_1037_));
 sg13g2_a21oi_1 _5366_ (.A1(_1035_),
    .A2(_1037_),
    .Y(_1038_),
    .B1(net41));
 sg13g2_buf_1 _5367_ (.A(_0819_),
    .X(_1039_));
 sg13g2_nand3_1 _5368_ (.B(net41),
    .C(_0706_),
    .A(_1015_),
    .Y(_1040_));
 sg13g2_nand3b_1 _5369_ (.B(net39),
    .C(_1040_),
    .Y(_1041_),
    .A_N(_1038_));
 sg13g2_nand2_1 _5370_ (.Y(_1042_),
    .A(_0708_),
    .B(net47));
 sg13g2_inv_1 _5371_ (.Y(_1043_),
    .A(_1042_));
 sg13g2_nor2_1 _5372_ (.A(net37),
    .B(_1043_),
    .Y(_1044_));
 sg13g2_a21oi_1 _5373_ (.A1(_1041_),
    .A2(_1044_),
    .Y(_1045_),
    .B1(net25));
 sg13g2_nand2_1 _5374_ (.Y(_1046_),
    .A(_1033_),
    .B(_1045_));
 sg13g2_nand2_1 _5375_ (.Y(_1047_),
    .A(_0994_),
    .B(_1046_));
 sg13g2_buf_2 _5376_ (.A(_0035_),
    .X(_1048_));
 sg13g2_inv_1 _5377_ (.Y(_1049_),
    .A(_1048_));
 sg13g2_xnor2_1 _5378_ (.Y(_1050_),
    .A(_1048_),
    .B(net113));
 sg13g2_nor2_1 _5379_ (.A(_0857_),
    .B(_3816_),
    .Y(_1051_));
 sg13g2_inv_1 _5380_ (.Y(_1052_),
    .A(_0843_));
 sg13g2_nor2_1 _5381_ (.A(_1052_),
    .B(net113),
    .Y(_1053_));
 sg13g2_a21oi_1 _5382_ (.A1(_0868_),
    .A2(_0839_),
    .Y(_1054_),
    .B1(_1053_));
 sg13g2_inv_1 _5383_ (.Y(_1055_),
    .A(_1054_));
 sg13g2_a21oi_1 _5384_ (.A1(_3884_),
    .A2(_1051_),
    .Y(_1056_),
    .B1(_1055_));
 sg13g2_inv_1 _5385_ (.Y(_1057_),
    .A(_1056_));
 sg13g2_o21ai_1 _5386_ (.B1(net60),
    .Y(_1058_),
    .A1(_1050_),
    .A2(_1057_));
 sg13g2_a21oi_1 _5387_ (.A1(_1050_),
    .A2(_1057_),
    .Y(_1059_),
    .B1(_1058_));
 sg13g2_xnor2_1 _5388_ (.Y(_1060_),
    .A(_1049_),
    .B(net72));
 sg13g2_a21oi_1 _5389_ (.A1(_0843_),
    .A2(_3871_),
    .Y(_1061_),
    .B1(_0876_));
 sg13g2_or2_1 _5390_ (.X(_1062_),
    .B(_1061_),
    .A(_1060_));
 sg13g2_nand2_1 _5391_ (.Y(_1063_),
    .A(_1062_),
    .B(_3652_));
 sg13g2_a21oi_1 _5392_ (.A1(_1060_),
    .A2(_1061_),
    .Y(_1064_),
    .B1(_1063_));
 sg13g2_nor2_1 _5393_ (.A(_3671_),
    .B(_1064_),
    .Y(_1065_));
 sg13g2_buf_1 _5394_ (.A(net76),
    .X(_1066_));
 sg13g2_buf_2 _5395_ (.A(\i_bitmap.in[9] ),
    .X(_1067_));
 sg13g2_xnor2_1 _5396_ (.Y(_1068_),
    .A(_1067_),
    .B(net100));
 sg13g2_inv_1 _5397_ (.Y(_1069_),
    .A(_0839_));
 sg13g2_a22oi_1 _5398_ (.Y(_1070_),
    .B1(_0851_),
    .B2(_0853_),
    .A2(_3897_),
    .A1(_1069_));
 sg13g2_xor2_1 _5399_ (.B(_1070_),
    .A(_1068_),
    .X(_1071_));
 sg13g2_xnor2_1 _5400_ (.Y(_1072_),
    .A(_1067_),
    .B(_0286_));
 sg13g2_inv_1 _5401_ (.Y(_1073_),
    .A(net78));
 sg13g2_a21oi_1 _5402_ (.A1(_1069_),
    .A2(_1073_),
    .Y(_1074_),
    .B1(_0847_));
 sg13g2_xnor2_1 _5403_ (.Y(_1075_),
    .A(_1072_),
    .B(_1074_));
 sg13g2_a21oi_1 _5404_ (.A1(_1075_),
    .A2(net76),
    .Y(_1076_),
    .B1(_0686_));
 sg13g2_o21ai_1 _5405_ (.B1(_1076_),
    .Y(_1077_),
    .A1(net74),
    .A2(_1071_));
 sg13g2_o21ai_1 _5406_ (.B1(_1077_),
    .Y(_1078_),
    .A1(_1059_),
    .A2(_1065_));
 sg13g2_a21oi_1 _5407_ (.A1(_1049_),
    .A2(net71),
    .Y(_1079_),
    .B1(_1078_));
 sg13g2_nor2_1 _5408_ (.A(_0838_),
    .B(_1079_),
    .Y(_1080_));
 sg13g2_inv_1 _5409_ (.Y(_1081_),
    .A(_1080_));
 sg13g2_nand2_1 _5410_ (.Y(_1082_),
    .A(_1047_),
    .B(_1081_));
 sg13g2_nand2_1 _5411_ (.Y(_1083_),
    .A(_0697_),
    .B(_0893_));
 sg13g2_nand2_1 _5412_ (.Y(_1084_),
    .A(_0924_),
    .B(_1083_));
 sg13g2_nor2_1 _5413_ (.A(_0997_),
    .B(_1084_),
    .Y(_1085_));
 sg13g2_nor2_1 _5414_ (.A(_1013_),
    .B(_1085_),
    .Y(_1086_));
 sg13g2_nor2_1 _5415_ (.A(_0593_),
    .B(net50),
    .Y(_1087_));
 sg13g2_nand2_1 _5416_ (.Y(_1088_),
    .A(_1087_),
    .B(_0702_));
 sg13g2_nand2_2 _5417_ (.Y(_1089_),
    .A(_0706_),
    .B(_0654_));
 sg13g2_buf_8 _5418_ (.A(net47),
    .X(_1090_));
 sg13g2_a21oi_1 _5419_ (.A1(_1088_),
    .A2(_1089_),
    .Y(_1091_),
    .B1(_1090_));
 sg13g2_o21ai_1 _5420_ (.B1(net27),
    .Y(_1092_),
    .A1(_1086_),
    .A2(_1091_));
 sg13g2_buf_1 _5421_ (.A(_0884_),
    .X(_1093_));
 sg13g2_nand2_1 _5422_ (.Y(_1094_),
    .A(_0593_),
    .B(_0654_));
 sg13g2_nor2_1 _5423_ (.A(_1094_),
    .B(_0835_),
    .Y(_1095_));
 sg13g2_a22oi_1 _5424_ (.Y(_1096_),
    .B1(_0820_),
    .B2(_0900_),
    .A2(_1095_),
    .A1(net29));
 sg13g2_nor2_1 _5425_ (.A(_0345_),
    .B(net31),
    .Y(_1097_));
 sg13g2_inv_1 _5426_ (.Y(_1098_),
    .A(_1097_));
 sg13g2_a21oi_1 _5427_ (.A1(_1092_),
    .A2(_1096_),
    .Y(_1099_),
    .B1(_1098_));
 sg13g2_a21oi_1 _5428_ (.A1(_1006_),
    .A2(net43),
    .Y(_1100_),
    .B1(_1026_));
 sg13g2_nor2_1 _5429_ (.A(net35),
    .B(_1100_),
    .Y(_1101_));
 sg13g2_nor2_1 _5430_ (.A(_1002_),
    .B(_1001_),
    .Y(_1102_));
 sg13g2_nor3_1 _5431_ (.A(net51),
    .B(_1102_),
    .C(_1085_),
    .Y(_1103_));
 sg13g2_o21ai_1 _5432_ (.B1(net29),
    .Y(_1104_),
    .A1(_1101_),
    .A2(_1103_));
 sg13g2_nor2_1 _5433_ (.A(_0823_),
    .B(_0929_),
    .Y(_1105_));
 sg13g2_inv_2 _5434_ (.Y(_1106_),
    .A(_0897_));
 sg13g2_nand2_1 _5435_ (.Y(_1107_),
    .A(_1023_),
    .B(net44));
 sg13g2_nor2_1 _5436_ (.A(_1106_),
    .B(_1107_),
    .Y(_1108_));
 sg13g2_o21ai_1 _5437_ (.B1(net39),
    .Y(_1109_),
    .A1(_1105_),
    .A2(_1108_));
 sg13g2_nand2_1 _5438_ (.Y(_1110_),
    .A(_1109_),
    .B(_1044_));
 sg13g2_nor2_1 _5439_ (.A(_0345_),
    .B(_0992_),
    .Y(_1111_));
 sg13g2_inv_2 _5440_ (.Y(_1112_),
    .A(_1111_));
 sg13g2_a21oi_1 _5441_ (.A1(_1104_),
    .A2(_1110_),
    .Y(_1113_),
    .B1(_1112_));
 sg13g2_nor2_1 _5442_ (.A(_1099_),
    .B(_1113_),
    .Y(_1114_));
 sg13g2_nand3_1 _5443_ (.B(_0702_),
    .C(net45),
    .A(_0996_),
    .Y(_1115_));
 sg13g2_nand3_1 _5444_ (.B(_0828_),
    .C(net38),
    .A(net42),
    .Y(_1116_));
 sg13g2_buf_2 _5445_ (.A(_1116_),
    .X(_1117_));
 sg13g2_a21oi_1 _5446_ (.A1(_1115_),
    .A2(_1117_),
    .Y(_1118_),
    .B1(net35));
 sg13g2_buf_1 _5447_ (.A(_0833_),
    .X(_1119_));
 sg13g2_nor2_1 _5448_ (.A(_0928_),
    .B(net50),
    .Y(_1120_));
 sg13g2_nand2_1 _5449_ (.Y(_1121_),
    .A(_1120_),
    .B(_1037_));
 sg13g2_nand2_1 _5450_ (.Y(_1122_),
    .A(_0894_),
    .B(net45));
 sg13g2_nand3_1 _5451_ (.B(net35),
    .C(_1122_),
    .A(_1121_),
    .Y(_1123_));
 sg13g2_nand3b_1 _5452_ (.B(net28),
    .C(_1123_),
    .Y(_1124_),
    .A_N(_1118_));
 sg13g2_nor2_1 _5453_ (.A(net49),
    .B(_0705_),
    .Y(_1125_));
 sg13g2_nor2_1 _5454_ (.A(_0833_),
    .B(_1095_),
    .Y(_1126_));
 sg13g2_nand3_1 _5455_ (.B(_1106_),
    .C(net44),
    .A(net47),
    .Y(_1127_));
 sg13g2_nand2_1 _5456_ (.Y(_1128_),
    .A(_1126_),
    .B(_1127_));
 sg13g2_nor2_1 _5457_ (.A(_1125_),
    .B(_1128_),
    .Y(_1129_));
 sg13g2_nor2_1 _5458_ (.A(net31),
    .B(_1129_),
    .Y(_1130_));
 sg13g2_nand2_1 _5459_ (.Y(_1131_),
    .A(_1124_),
    .B(_1130_));
 sg13g2_nor3_1 _5460_ (.A(_1007_),
    .B(net51),
    .C(_0895_),
    .Y(_1132_));
 sg13g2_nand2_1 _5461_ (.Y(_1133_),
    .A(net51),
    .B(_0929_));
 sg13g2_a21oi_1 _5462_ (.A1(_1087_),
    .A2(_1023_),
    .Y(_1134_),
    .B1(_1133_));
 sg13g2_nor3_1 _5463_ (.A(net37),
    .B(_1132_),
    .C(_1134_),
    .Y(_1135_));
 sg13g2_nor2_1 _5464_ (.A(net25),
    .B(_1135_),
    .Y(_1136_));
 sg13g2_inv_1 _5465_ (.Y(_1137_),
    .A(_1006_));
 sg13g2_nor3_1 _5466_ (.A(_1137_),
    .B(net47),
    .C(_1003_),
    .Y(_1138_));
 sg13g2_o21ai_1 _5467_ (.B1(_0832_),
    .Y(_1139_),
    .A1(_1089_),
    .A2(net47));
 sg13g2_nor2_1 _5468_ (.A(_1138_),
    .B(_1139_),
    .Y(_1140_));
 sg13g2_nand2b_1 _5469_ (.Y(_1141_),
    .B(_1140_),
    .A_N(_1103_));
 sg13g2_nand2_1 _5470_ (.Y(_1142_),
    .A(_1136_),
    .B(_1141_));
 sg13g2_nand2_1 _5471_ (.Y(_1143_),
    .A(_1131_),
    .B(_1142_));
 sg13g2_nand2_1 _5472_ (.Y(_1144_),
    .A(_1143_),
    .B(_0346_));
 sg13g2_nand2_1 _5473_ (.Y(_1145_),
    .A(_1114_),
    .B(_1144_));
 sg13g2_nand2_1 _5474_ (.Y(_1146_),
    .A(_1145_),
    .B(net46));
 sg13g2_inv_1 _5475_ (.Y(_1147_),
    .A(_0771_));
 sg13g2_nand2_1 _5476_ (.Y(_1148_),
    .A(net44),
    .B(_0592_));
 sg13g2_buf_1 _5477_ (.A(_0836_),
    .X(_1149_));
 sg13g2_nor2_1 _5478_ (.A(_1148_),
    .B(net34),
    .Y(_1150_));
 sg13g2_nor2_1 _5479_ (.A(_1147_),
    .B(_1150_),
    .Y(_1151_));
 sg13g2_nand2_1 _5480_ (.Y(_1152_),
    .A(net49),
    .B(_1094_));
 sg13g2_nand2_1 _5481_ (.Y(_1153_),
    .A(_0897_),
    .B(net36));
 sg13g2_a21oi_1 _5482_ (.A1(_1152_),
    .A2(_1153_),
    .Y(_1154_),
    .B1(net27));
 sg13g2_nor3_1 _5483_ (.A(net31),
    .B(_1151_),
    .C(_1154_),
    .Y(_1155_));
 sg13g2_a21oi_1 _5484_ (.A1(_1155_),
    .A2(_0883_),
    .Y(_1156_),
    .B1(_1081_));
 sg13g2_nand2_1 _5485_ (.Y(_1157_),
    .A(_1146_),
    .B(_1156_));
 sg13g2_nand2_1 _5486_ (.Y(_1158_),
    .A(_1082_),
    .B(_1157_));
 sg13g2_buf_1 _5487_ (.A(_0036_),
    .X(_1159_));
 sg13g2_inv_1 _5488_ (.Y(_1160_),
    .A(_1159_));
 sg13g2_buf_2 _5489_ (.A(\i_bitmap.in[10] ),
    .X(_1161_));
 sg13g2_xnor2_1 _5490_ (.Y(_1162_),
    .A(_1161_),
    .B(net75));
 sg13g2_nand2_1 _5491_ (.Y(_1163_),
    .A(_0286_),
    .B(_1049_));
 sg13g2_o21ai_1 _5492_ (.B1(_1163_),
    .Y(_1164_),
    .A1(_1072_),
    .A2(_1074_));
 sg13g2_xor2_1 _5493_ (.B(_1164_),
    .A(_1162_),
    .X(_1165_));
 sg13g2_xnor2_1 _5494_ (.Y(_1166_),
    .A(_1161_),
    .B(net100));
 sg13g2_nor2_1 _5495_ (.A(_1068_),
    .B(_0850_),
    .Y(_1167_));
 sg13g2_nand3b_1 _5496_ (.B(_3897_),
    .C(_1069_),
    .Y(_1168_),
    .A_N(_1067_));
 sg13g2_o21ai_1 _5497_ (.B1(_1168_),
    .Y(_1169_),
    .A1(_1048_),
    .A2(_0750_));
 sg13g2_a21o_1 _5498_ (.A2(_1167_),
    .A1(_0853_),
    .B1(_1169_),
    .X(_1170_));
 sg13g2_a21oi_1 _5499_ (.A1(_1170_),
    .A2(_1166_),
    .Y(_1171_),
    .B1(net74));
 sg13g2_o21ai_1 _5500_ (.B1(_1171_),
    .Y(_1172_),
    .A1(_1166_),
    .A2(_1170_));
 sg13g2_o21ai_1 _5501_ (.B1(_1172_),
    .Y(_1173_),
    .A1(net77),
    .A2(_1165_));
 sg13g2_xnor2_1 _5502_ (.Y(_1174_),
    .A(_1159_),
    .B(net113));
 sg13g2_inv_1 _5503_ (.Y(_1175_),
    .A(_1174_));
 sg13g2_nor2_1 _5504_ (.A(_1050_),
    .B(_0857_),
    .Y(_1176_));
 sg13g2_nand2_1 _5505_ (.Y(_1177_),
    .A(net114),
    .B(_1067_));
 sg13g2_inv_1 _5506_ (.Y(_1178_),
    .A(_1177_));
 sg13g2_a21oi_1 _5507_ (.A1(_1048_),
    .A2(_1053_),
    .Y(_1179_),
    .B1(_1178_));
 sg13g2_inv_1 _5508_ (.Y(_1180_),
    .A(_1179_));
 sg13g2_a21oi_1 _5509_ (.A1(_0870_),
    .A2(_1176_),
    .Y(_1181_),
    .B1(_1180_));
 sg13g2_xnor2_1 _5510_ (.Y(_1182_),
    .A(_1175_),
    .B(_1181_));
 sg13g2_xnor2_1 _5511_ (.Y(_1183_),
    .A(_1159_),
    .B(net79));
 sg13g2_nand2_1 _5512_ (.Y(_1184_),
    .A(net72),
    .B(_1067_));
 sg13g2_nand2_1 _5513_ (.Y(_1185_),
    .A(_1062_),
    .B(_1184_));
 sg13g2_xnor2_1 _5514_ (.Y(_1186_),
    .A(_1183_),
    .B(_1185_));
 sg13g2_a21oi_1 _5515_ (.A1(_1186_),
    .A2(net62),
    .Y(_1187_),
    .B1(net63));
 sg13g2_o21ai_1 _5516_ (.B1(_1187_),
    .Y(_1188_),
    .A1(net62),
    .A2(_1182_));
 sg13g2_o21ai_1 _5517_ (.B1(_1188_),
    .Y(_1189_),
    .A1(_0686_),
    .A2(_1173_));
 sg13g2_a21oi_1 _5518_ (.A1(_1160_),
    .A2(net71),
    .Y(_1190_),
    .B1(_1189_));
 sg13g2_nor2_1 _5519_ (.A(_0838_),
    .B(_1190_),
    .Y(_1191_));
 sg13g2_inv_1 _5520_ (.Y(_1192_),
    .A(_1191_));
 sg13g2_nand2_1 _5521_ (.Y(_1193_),
    .A(_1158_),
    .B(_1192_));
 sg13g2_inv_1 _5522_ (.Y(_1194_),
    .A(_0925_));
 sg13g2_nand2_1 _5523_ (.Y(_1195_),
    .A(net43),
    .B(net38));
 sg13g2_nand3_1 _5524_ (.B(_1117_),
    .C(_1195_),
    .A(_1194_),
    .Y(_1196_));
 sg13g2_nand2_1 _5525_ (.Y(_1197_),
    .A(_1196_),
    .B(_1149_));
 sg13g2_a21oi_1 _5526_ (.A1(_0925_),
    .A2(_0885_),
    .Y(_1198_),
    .B1(net29));
 sg13g2_nand3_1 _5527_ (.B(_0903_),
    .C(_1198_),
    .A(_1197_),
    .Y(_1199_));
 sg13g2_o21ai_1 _5528_ (.B1(_1032_),
    .Y(_1200_),
    .A1(_1029_),
    .A2(_0919_));
 sg13g2_nand2_1 _5529_ (.Y(_1201_),
    .A(_1199_),
    .B(_1200_));
 sg13g2_nor2_1 _5530_ (.A(_0935_),
    .B(_0991_),
    .Y(_1202_));
 sg13g2_inv_1 _5531_ (.Y(_1203_),
    .A(_0903_));
 sg13g2_nor3_1 _5532_ (.A(_0934_),
    .B(net37),
    .C(_1203_),
    .Y(_1204_));
 sg13g2_inv_1 _5533_ (.Y(_1205_),
    .A(_0888_));
 sg13g2_a21oi_1 _5534_ (.A1(_1149_),
    .A2(_1205_),
    .Y(_1206_),
    .B1(net28));
 sg13g2_a21oi_1 _5535_ (.A1(_1197_),
    .A2(_1204_),
    .Y(_1207_),
    .B1(_1206_));
 sg13g2_nor2_1 _5536_ (.A(_1098_),
    .B(_1207_),
    .Y(_1208_));
 sg13g2_a21oi_1 _5537_ (.A1(_1201_),
    .A2(_1202_),
    .Y(_1209_),
    .B1(_1208_));
 sg13g2_nand2_1 _5538_ (.Y(_1210_),
    .A(_1008_),
    .B(_1027_));
 sg13g2_nand2_1 _5539_ (.Y(_1211_),
    .A(_1210_),
    .B(_1009_));
 sg13g2_buf_1 _5540_ (.A(net45),
    .X(_1212_));
 sg13g2_nand2_1 _5541_ (.Y(_1213_),
    .A(_1035_),
    .B(net33));
 sg13g2_nand2_1 _5542_ (.Y(_1214_),
    .A(_1027_),
    .B(_1213_));
 sg13g2_nand2_1 _5543_ (.Y(_1215_),
    .A(_1214_),
    .B(_0913_));
 sg13g2_nand2_1 _5544_ (.Y(_1216_),
    .A(_0826_),
    .B(net43));
 sg13g2_a21o_1 _5545_ (.A2(_1035_),
    .A1(_1216_),
    .B1(net39),
    .X(_1217_));
 sg13g2_nand3_1 _5546_ (.B(_1215_),
    .C(_1217_),
    .A(_1211_),
    .Y(_1218_));
 sg13g2_nand2_1 _5547_ (.Y(_1219_),
    .A(_1218_),
    .B(net30));
 sg13g2_a21oi_1 _5548_ (.A1(_1000_),
    .A2(net52),
    .Y(_1220_),
    .B1(_1005_));
 sg13g2_inv_1 _5549_ (.Y(_1221_),
    .A(_1220_));
 sg13g2_a21oi_2 _5550_ (.B1(net35),
    .Y(_1222_),
    .A2(_1022_),
    .A1(_1221_));
 sg13g2_nand2_1 _5551_ (.Y(_1223_),
    .A(_1222_),
    .B(net28));
 sg13g2_nor2_1 _5552_ (.A(_0704_),
    .B(_1223_),
    .Y(_1224_));
 sg13g2_nor2_1 _5553_ (.A(net25),
    .B(_1224_),
    .Y(_1225_));
 sg13g2_a21oi_1 _5554_ (.A1(_1219_),
    .A2(_1225_),
    .Y(_1226_),
    .B1(net46));
 sg13g2_nand2_1 _5555_ (.Y(_1227_),
    .A(_1209_),
    .B(_1226_));
 sg13g2_inv_1 _5556_ (.Y(_1228_),
    .A(_0829_));
 sg13g2_o21ai_1 _5557_ (.B1(_1228_),
    .Y(_1229_),
    .A1(_1137_),
    .A2(_1003_));
 sg13g2_nor2_1 _5558_ (.A(_0885_),
    .B(_1229_),
    .Y(_1230_));
 sg13g2_nor2_1 _5559_ (.A(net29),
    .B(_1230_),
    .Y(_1231_));
 sg13g2_nand2_1 _5560_ (.Y(_1232_),
    .A(_0904_),
    .B(_0913_));
 sg13g2_nand2_1 _5561_ (.Y(_1233_),
    .A(_0909_),
    .B(_1228_));
 sg13g2_nand3_1 _5562_ (.B(net40),
    .C(net54),
    .A(_1233_),
    .Y(_1234_));
 sg13g2_nand3_1 _5563_ (.B(_1232_),
    .C(_1234_),
    .A(_1231_),
    .Y(_1235_));
 sg13g2_nand3_1 _5564_ (.B(_0887_),
    .C(_0888_),
    .A(net40),
    .Y(_1236_));
 sg13g2_a21oi_1 _5565_ (.A1(_1206_),
    .A2(_1236_),
    .Y(_1237_),
    .B1(net31));
 sg13g2_nand2_1 _5566_ (.Y(_1238_),
    .A(_1235_),
    .B(_1237_));
 sg13g2_nand3_1 _5567_ (.B(_1037_),
    .C(net43),
    .A(_0924_),
    .Y(_1239_));
 sg13g2_nand2_1 _5568_ (.Y(_1240_),
    .A(_1027_),
    .B(_1239_));
 sg13g2_nand2_1 _5569_ (.Y(_1241_),
    .A(_1240_),
    .B(net49));
 sg13g2_nand2_1 _5570_ (.Y(_1242_),
    .A(_0826_),
    .B(net41));
 sg13g2_nand3_1 _5571_ (.B(net47),
    .C(_1242_),
    .A(_0998_),
    .Y(_1243_));
 sg13g2_nand2_1 _5572_ (.Y(_1244_),
    .A(_1241_),
    .B(_1243_));
 sg13g2_nand2_1 _5573_ (.Y(_1245_),
    .A(_1244_),
    .B(_1093_));
 sg13g2_nand4_1 _5574_ (.B(_1220_),
    .C(_1039_),
    .A(_1119_),
    .Y(_1246_),
    .D(_1022_));
 sg13g2_nand2_1 _5575_ (.Y(_1247_),
    .A(_1245_),
    .B(_1246_));
 sg13g2_buf_1 _5576_ (.A(net31),
    .X(_1248_));
 sg13g2_nand2_1 _5577_ (.Y(_1249_),
    .A(_1247_),
    .B(net26));
 sg13g2_nand2_1 _5578_ (.Y(_1250_),
    .A(_1238_),
    .B(_1249_));
 sg13g2_nand2_1 _5579_ (.Y(_1251_),
    .A(_1250_),
    .B(_0939_));
 sg13g2_nand2_1 _5580_ (.Y(_1252_),
    .A(_1227_),
    .B(_1251_));
 sg13g2_nand2_1 _5581_ (.Y(_1253_),
    .A(_1252_),
    .B(_1080_));
 sg13g2_nand3_1 _5582_ (.B(_1083_),
    .C(net44),
    .A(_0924_),
    .Y(_1254_));
 sg13g2_nand2_1 _5583_ (.Y(_1255_),
    .A(_0888_),
    .B(_1000_));
 sg13g2_nand2_1 _5584_ (.Y(_1256_),
    .A(_1254_),
    .B(_1255_));
 sg13g2_nand2_1 _5585_ (.Y(_1257_),
    .A(_1256_),
    .B(net34));
 sg13g2_nand2_1 _5586_ (.Y(_1258_),
    .A(_1100_),
    .B(net40));
 sg13g2_nor2_1 _5587_ (.A(_0989_),
    .B(net55),
    .Y(_1259_));
 sg13g2_nand4_1 _5588_ (.B(_1258_),
    .C(net30),
    .A(_1257_),
    .Y(_1260_),
    .D(_1259_));
 sg13g2_nand2_1 _5589_ (.Y(_1261_),
    .A(_1260_),
    .B(_0883_));
 sg13g2_a21oi_1 _5590_ (.A1(_1089_),
    .A2(_1088_),
    .Y(_1262_),
    .B1(_1010_));
 sg13g2_a21oi_1 _5591_ (.A1(_0998_),
    .A2(_1117_),
    .Y(_1263_),
    .B1(_0912_));
 sg13g2_nand3_1 _5592_ (.B(_0816_),
    .C(_1228_),
    .A(_1254_),
    .Y(_1264_));
 sg13g2_nand2_1 _5593_ (.Y(_1265_),
    .A(_1264_),
    .B(net25));
 sg13g2_nor3_1 _5594_ (.A(_1262_),
    .B(_1263_),
    .C(_1265_),
    .Y(_1266_));
 sg13g2_nand3_1 _5595_ (.B(net28),
    .C(_1205_),
    .A(_1222_),
    .Y(_1267_));
 sg13g2_nand2_1 _5596_ (.Y(_1268_),
    .A(net27),
    .B(_0989_));
 sg13g2_nand2_1 _5597_ (.Y(_1269_),
    .A(_1267_),
    .B(_1268_));
 sg13g2_nor2b_1 _5598_ (.A(_1266_),
    .B_N(_1269_),
    .Y(_1270_));
 sg13g2_nor2_1 _5599_ (.A(_1261_),
    .B(_1270_),
    .Y(_1271_));
 sg13g2_nor2_1 _5600_ (.A(net52),
    .B(_0887_),
    .Y(_1272_));
 sg13g2_nand2_1 _5601_ (.Y(_1273_),
    .A(_1272_),
    .B(net50));
 sg13g2_nand2_1 _5602_ (.Y(_1274_),
    .A(_1273_),
    .B(_0929_));
 sg13g2_nand2_1 _5603_ (.Y(_1275_),
    .A(_1274_),
    .B(net40));
 sg13g2_a21oi_2 _5604_ (.B1(net51),
    .Y(_1276_),
    .A2(_1000_),
    .A1(_0888_));
 sg13g2_nand2_1 _5605_ (.Y(_1277_),
    .A(_1276_),
    .B(_1121_));
 sg13g2_nand2_1 _5606_ (.Y(_1278_),
    .A(_1120_),
    .B(net40));
 sg13g2_nand3_1 _5607_ (.B(_1277_),
    .C(_1278_),
    .A(_1275_),
    .Y(_1279_));
 sg13g2_nand2_1 _5608_ (.Y(_1280_),
    .A(_1095_),
    .B(net55));
 sg13g2_a21oi_1 _5609_ (.A1(_1280_),
    .A2(_1127_),
    .Y(_1281_),
    .B1(net26));
 sg13g2_a21oi_1 _5610_ (.A1(_1279_),
    .A2(_1111_),
    .Y(_1282_),
    .B1(_1281_));
 sg13g2_nand2b_1 _5611_ (.Y(_1283_),
    .B(_1032_),
    .A_N(_1282_));
 sg13g2_nand2_1 _5612_ (.Y(_1284_),
    .A(_1271_),
    .B(_1283_));
 sg13g2_a21oi_1 _5613_ (.A1(_1155_),
    .A2(_0935_),
    .Y(_1285_),
    .B1(_0883_));
 sg13g2_o21ai_1 _5614_ (.B1(_0911_),
    .Y(_1286_),
    .A1(_0816_),
    .A2(_1117_));
 sg13g2_nand3_1 _5615_ (.B(_1202_),
    .C(_1286_),
    .A(_1128_),
    .Y(_1287_));
 sg13g2_a21oi_1 _5616_ (.A1(_1285_),
    .A2(_1287_),
    .Y(_1288_),
    .B1(_1080_));
 sg13g2_a21oi_1 _5617_ (.A1(_1284_),
    .A2(_1288_),
    .Y(_1289_),
    .B1(_1192_));
 sg13g2_inv_1 _5618_ (.Y(_1290_),
    .A(_0037_));
 sg13g2_buf_2 _5619_ (.A(\i_bitmap.in[11] ),
    .X(_1291_));
 sg13g2_xnor2_1 _5620_ (.Y(_1292_),
    .A(_1291_),
    .B(net113));
 sg13g2_a22oi_1 _5621_ (.Y(_1293_),
    .B1(_1183_),
    .B2(_1185_),
    .A2(_3861_),
    .A1(_1161_));
 sg13g2_nor2_1 _5622_ (.A(_1292_),
    .B(_1293_),
    .Y(_1294_));
 sg13g2_inv_1 _5623_ (.Y(_1295_),
    .A(_1294_));
 sg13g2_nand2_1 _5624_ (.Y(_1296_),
    .A(_1293_),
    .B(_1292_));
 sg13g2_a21oi_1 _5625_ (.A1(_1295_),
    .A2(_1296_),
    .Y(_1297_),
    .B1(net60));
 sg13g2_nor2_1 _5626_ (.A(_1174_),
    .B(_1050_),
    .Y(_1298_));
 sg13g2_inv_1 _5627_ (.Y(_1299_),
    .A(_1161_));
 sg13g2_nor2_1 _5628_ (.A(_1299_),
    .B(_0856_),
    .Y(_1300_));
 sg13g2_a221oi_1 _5629_ (.B2(_1298_),
    .C1(_1300_),
    .B1(_1057_),
    .A1(_1159_),
    .Y(_1301_),
    .A2(_1178_));
 sg13g2_xnor2_1 _5630_ (.Y(_1302_),
    .A(_0037_),
    .B(net113));
 sg13g2_nand2b_1 _5631_ (.Y(_1303_),
    .B(_1302_),
    .A_N(_1301_));
 sg13g2_inv_1 _5632_ (.Y(_1304_),
    .A(_1302_));
 sg13g2_nand2_1 _5633_ (.Y(_1305_),
    .A(_1301_),
    .B(_1304_));
 sg13g2_nand3_1 _5634_ (.B(net60),
    .C(_1305_),
    .A(_1303_),
    .Y(_1306_));
 sg13g2_nand3b_1 _5635_ (.B(_1306_),
    .C(_0689_),
    .Y(_1307_),
    .A_N(_1297_));
 sg13g2_xnor2_1 _5636_ (.Y(_1308_),
    .A(_1291_),
    .B(net100));
 sg13g2_inv_1 _5637_ (.Y(_1309_),
    .A(_1308_));
 sg13g2_inv_1 _5638_ (.Y(_1310_),
    .A(_1166_));
 sg13g2_a22oi_1 _5639_ (.Y(_1311_),
    .B1(_1310_),
    .B2(_1170_),
    .A2(net100),
    .A1(_1160_));
 sg13g2_xnor2_1 _5640_ (.Y(_1312_),
    .A(_1309_),
    .B(_1311_));
 sg13g2_xnor2_1 _5641_ (.Y(_1313_),
    .A(_1290_),
    .B(net100));
 sg13g2_nand2_1 _5642_ (.Y(_1314_),
    .A(_1164_),
    .B(_1162_));
 sg13g2_o21ai_1 _5643_ (.B1(_1314_),
    .Y(_1315_),
    .A1(_1159_),
    .A2(_3954_));
 sg13g2_xnor2_1 _5644_ (.Y(_1316_),
    .A(_1313_),
    .B(_1315_));
 sg13g2_a21oi_1 _5645_ (.A1(_1316_),
    .A2(_1066_),
    .Y(_1317_),
    .B1(_0686_));
 sg13g2_o21ai_1 _5646_ (.B1(_1317_),
    .Y(_1318_),
    .A1(_1066_),
    .A2(_1312_));
 sg13g2_nand2_1 _5647_ (.Y(_1319_),
    .A(_1307_),
    .B(_1318_));
 sg13g2_a21oi_1 _5648_ (.A1(_1290_),
    .A2(_0337_),
    .Y(_1320_),
    .B1(_1319_));
 sg13g2_nor2_1 _5649_ (.A(_0838_),
    .B(_1320_),
    .Y(_1321_));
 sg13g2_a21oi_1 _5650_ (.A1(_1253_),
    .A2(_1289_),
    .Y(_1322_),
    .B1(_1321_));
 sg13g2_nand2_1 _5651_ (.Y(_1323_),
    .A(_0996_),
    .B(_1212_));
 sg13g2_a21oi_1 _5652_ (.A1(_0899_),
    .A2(_1323_),
    .Y(_1324_),
    .B1(net54));
 sg13g2_nand2_1 _5653_ (.Y(_1325_),
    .A(_0655_),
    .B(_0933_));
 sg13g2_nor2_1 _5654_ (.A(_1272_),
    .B(_1325_),
    .Y(_1326_));
 sg13g2_nor2_1 _5655_ (.A(_0818_),
    .B(_1326_),
    .Y(_1327_));
 sg13g2_nand2_1 _5656_ (.Y(_1328_),
    .A(_0897_),
    .B(net33));
 sg13g2_nor2_1 _5657_ (.A(_0341_),
    .B(net39),
    .Y(_1329_));
 sg13g2_a21oi_1 _5658_ (.A1(_1327_),
    .A2(_1328_),
    .Y(_1330_),
    .B1(_1329_));
 sg13g2_nor3_1 _5659_ (.A(_0771_),
    .B(_1324_),
    .C(_1330_),
    .Y(_1331_));
 sg13g2_nand2_1 _5660_ (.Y(_1332_),
    .A(_1229_),
    .B(net34));
 sg13g2_nand2_1 _5661_ (.Y(_1333_),
    .A(_0708_),
    .B(net51));
 sg13g2_nor2_1 _5662_ (.A(_0829_),
    .B(_1333_),
    .Y(_1334_));
 sg13g2_nand2_1 _5663_ (.Y(_1335_),
    .A(_1334_),
    .B(net54));
 sg13g2_nor3_1 _5664_ (.A(_0829_),
    .B(_1090_),
    .C(_0918_),
    .Y(_1336_));
 sg13g2_nand2_1 _5665_ (.Y(_1337_),
    .A(_1336_),
    .B(net55));
 sg13g2_nand4_1 _5666_ (.B(_1335_),
    .C(_1337_),
    .A(_1332_),
    .Y(_1338_),
    .D(_0911_));
 sg13g2_nand3b_1 _5667_ (.B(_0993_),
    .C(_1338_),
    .Y(_1339_),
    .A_N(_1331_));
 sg13g2_nand2_1 _5668_ (.Y(_1340_),
    .A(_1028_),
    .B(net40));
 sg13g2_nand2_1 _5669_ (.Y(_1341_),
    .A(_1340_),
    .B(_1243_));
 sg13g2_nand2_1 _5670_ (.Y(_1342_),
    .A(_1341_),
    .B(net30));
 sg13g2_nand3_1 _5671_ (.B(net26),
    .C(_1246_),
    .A(_1342_),
    .Y(_1343_));
 sg13g2_a21oi_1 _5672_ (.A1(_1339_),
    .A2(_1343_),
    .Y(_1344_),
    .B1(_0883_));
 sg13g2_nand2_1 _5673_ (.Y(_1345_),
    .A(_1086_),
    .B(_1122_));
 sg13g2_nand3_1 _5674_ (.B(net27),
    .C(_1275_),
    .A(_1345_),
    .Y(_1346_));
 sg13g2_nor2b_1 _5675_ (.A(_1087_),
    .B_N(_1094_),
    .Y(_1347_));
 sg13g2_a21oi_1 _5676_ (.A1(_1347_),
    .A2(net47),
    .Y(_1348_),
    .B1(net32));
 sg13g2_nor2_1 _5677_ (.A(_1248_),
    .B(_1348_),
    .Y(_1349_));
 sg13g2_a21oi_1 _5678_ (.A1(_1346_),
    .A2(_1349_),
    .Y(_1350_),
    .B1(net55));
 sg13g2_nand2_1 _5679_ (.Y(_1351_),
    .A(_0703_),
    .B(net45));
 sg13g2_a22oi_1 _5680_ (.Y(_1352_),
    .B1(_1351_),
    .B2(_0926_),
    .A2(_1121_),
    .A1(_1276_));
 sg13g2_nor2_1 _5681_ (.A(_0888_),
    .B(net34),
    .Y(_1353_));
 sg13g2_a21oi_1 _5682_ (.A1(_1353_),
    .A2(_1117_),
    .Y(_1354_),
    .B1(net29));
 sg13g2_a21oi_1 _5683_ (.A1(_1352_),
    .A2(net30),
    .Y(_1355_),
    .B1(_1354_));
 sg13g2_nand2_1 _5684_ (.Y(_1356_),
    .A(_1355_),
    .B(net26));
 sg13g2_nand2_1 _5685_ (.Y(_1357_),
    .A(_1350_),
    .B(_1356_));
 sg13g2_nand3_1 _5686_ (.B(net30),
    .C(_1258_),
    .A(_1257_),
    .Y(_1358_));
 sg13g2_nand3_1 _5687_ (.B(_1005_),
    .C(net42),
    .A(net44),
    .Y(_1359_));
 sg13g2_nand3_1 _5688_ (.B(net27),
    .C(_1359_),
    .A(_1353_),
    .Y(_1360_));
 sg13g2_nor2b_1 _5689_ (.A(_1112_),
    .B_N(_1360_),
    .Y(_1361_));
 sg13g2_nor2_1 _5690_ (.A(net29),
    .B(_1086_),
    .Y(_1362_));
 sg13g2_nand2_1 _5691_ (.Y(_1363_),
    .A(_1362_),
    .B(_1089_));
 sg13g2_nor2_1 _5692_ (.A(_0699_),
    .B(net50),
    .Y(_1364_));
 sg13g2_o21ai_1 _5693_ (.B1(net48),
    .Y(_1365_),
    .A1(_0818_),
    .A2(_1364_));
 sg13g2_nand2_1 _5694_ (.Y(_1366_),
    .A(_1363_),
    .B(_1365_));
 sg13g2_a22oi_1 _5695_ (.Y(_1367_),
    .B1(_1097_),
    .B2(_1366_),
    .A2(_1361_),
    .A1(_1358_));
 sg13g2_a21o_1 _5696_ (.A2(_1367_),
    .A1(_1357_),
    .B1(net46),
    .X(_1368_));
 sg13g2_and3_1 _5697_ (.X(_1369_),
    .A(_1321_),
    .B(_1190_),
    .C(_1079_));
 sg13g2_nand3b_1 _5698_ (.B(_1368_),
    .C(_1369_),
    .Y(_1370_),
    .A_N(_1344_));
 sg13g2_buf_1 _5699_ (.A(_0686_),
    .X(_1371_));
 sg13g2_nand2_1 _5700_ (.Y(_1372_),
    .A(_3650_),
    .B(_1371_));
 sg13g2_nor2_1 _5701_ (.A(_0038_),
    .B(_1372_),
    .Y(_1373_));
 sg13g2_nand2b_1 _5702_ (.Y(_1374_),
    .B(_1309_),
    .A_N(_1311_));
 sg13g2_buf_2 _5703_ (.A(\i_bitmap.in[12] ),
    .X(_1375_));
 sg13g2_buf_1 _5704_ (.A(net100),
    .X(_1376_));
 sg13g2_xnor2_1 _5705_ (.Y(_1377_),
    .A(_1375_),
    .B(net91));
 sg13g2_nand2_1 _5706_ (.Y(_1378_),
    .A(net91),
    .B(_1290_));
 sg13g2_and2_1 _5707_ (.A(_1377_),
    .B(_1378_),
    .X(_1379_));
 sg13g2_a21oi_1 _5708_ (.A1(_1374_),
    .A2(_1378_),
    .Y(_1380_),
    .B1(_1377_));
 sg13g2_a21oi_1 _5709_ (.A1(_1374_),
    .A2(_1379_),
    .Y(_1381_),
    .B1(_1380_));
 sg13g2_nand2_1 _5710_ (.Y(_1382_),
    .A(_1315_),
    .B(_1313_));
 sg13g2_nand2_1 _5711_ (.Y(_1383_),
    .A(net92),
    .B(_1291_));
 sg13g2_xnor2_1 _5712_ (.Y(_1384_),
    .A(_0038_),
    .B(_1376_));
 sg13g2_a21o_1 _5713_ (.A2(_1383_),
    .A1(_1382_),
    .B1(_1384_),
    .X(_1385_));
 sg13g2_nand3_1 _5714_ (.B(_1383_),
    .C(_1384_),
    .A(_1382_),
    .Y(_1386_));
 sg13g2_a21o_1 _5715_ (.A2(_1386_),
    .A1(_1385_),
    .B1(_0320_),
    .X(_1387_));
 sg13g2_o21ai_1 _5716_ (.B1(_1387_),
    .Y(_1388_),
    .A1(net74),
    .A2(_1381_));
 sg13g2_inv_1 _5717_ (.Y(_1389_),
    .A(_0038_));
 sg13g2_buf_1 _5718_ (.A(_0856_),
    .X(_1390_));
 sg13g2_xnor2_1 _5719_ (.Y(_1391_),
    .A(_1389_),
    .B(net98));
 sg13g2_nand2_1 _5720_ (.Y(_1392_),
    .A(_1304_),
    .B(_1175_));
 sg13g2_a22oi_1 _5721_ (.Y(_1393_),
    .B1(_0037_),
    .B2(_1300_),
    .A2(_1291_),
    .A1(_0605_));
 sg13g2_o21ai_1 _5722_ (.B1(_1393_),
    .Y(_1394_),
    .A1(_1392_),
    .A2(_1181_));
 sg13g2_xor2_1 _5723_ (.B(_1394_),
    .A(_1391_),
    .X(_1395_));
 sg13g2_nand2_1 _5724_ (.Y(_1396_),
    .A(net98),
    .B(_1290_));
 sg13g2_xnor2_1 _5725_ (.Y(_1397_),
    .A(_1375_),
    .B(net113));
 sg13g2_a21oi_1 _5726_ (.A1(_1295_),
    .A2(_1396_),
    .Y(_1398_),
    .B1(_1397_));
 sg13g2_nand3_1 _5727_ (.B(_1396_),
    .C(_1397_),
    .A(_1295_),
    .Y(_1399_));
 sg13g2_nand3b_1 _5728_ (.B(_1399_),
    .C(_0689_),
    .Y(_1400_),
    .A_N(_1398_));
 sg13g2_nand2_1 _5729_ (.Y(_1401_),
    .A(_1400_),
    .B(_0959_));
 sg13g2_o21ai_1 _5730_ (.B1(_1401_),
    .Y(_1402_),
    .A1(net62),
    .A2(_1395_));
 sg13g2_o21ai_1 _5731_ (.B1(_1402_),
    .Y(_1403_),
    .A1(_1371_),
    .A2(_1388_));
 sg13g2_o21ai_1 _5732_ (.B1(net147),
    .Y(_1404_),
    .A1(_1373_),
    .A2(_1403_));
 sg13g2_nand2_1 _5733_ (.Y(_1405_),
    .A(_1370_),
    .B(_1404_));
 sg13g2_a21oi_1 _5734_ (.A1(_1193_),
    .A2(_1322_),
    .Y(_1406_),
    .B1(_1405_));
 sg13g2_a21oi_1 _5735_ (.A1(_0706_),
    .A2(_0654_),
    .Y(_1407_),
    .B1(_0816_));
 sg13g2_a21oi_1 _5736_ (.A1(_1407_),
    .A2(_1107_),
    .Y(_1408_),
    .B1(net29));
 sg13g2_inv_1 _5737_ (.Y(_1409_),
    .A(_0825_));
 sg13g2_a21oi_1 _5738_ (.A1(_1409_),
    .A2(net42),
    .Y(_1410_),
    .B1(_0887_));
 sg13g2_a21oi_1 _5739_ (.A1(_1410_),
    .A2(net33),
    .Y(_1411_),
    .B1(net39));
 sg13g2_nand3_1 _5740_ (.B(net36),
    .C(_1037_),
    .A(_1035_),
    .Y(_1412_));
 sg13g2_nand2_1 _5741_ (.Y(_1413_),
    .A(_1411_),
    .B(_1412_));
 sg13g2_nand3_1 _5742_ (.B(net43),
    .C(_0933_),
    .A(_1024_),
    .Y(_1414_));
 sg13g2_nand2_1 _5743_ (.Y(_1415_),
    .A(_1222_),
    .B(_1414_));
 sg13g2_nand3_1 _5744_ (.B(_1415_),
    .C(net29),
    .A(_1413_),
    .Y(_1416_));
 sg13g2_nand2b_1 _5745_ (.Y(_1417_),
    .B(_1416_),
    .A_N(_1408_));
 sg13g2_inv_1 _5746_ (.Y(_1418_),
    .A(_1079_));
 sg13g2_a21oi_1 _5747_ (.A1(_1417_),
    .A2(net26),
    .Y(_1419_),
    .B1(_1418_));
 sg13g2_nand3_1 _5748_ (.B(_0933_),
    .C(net44),
    .A(_0897_),
    .Y(_1420_));
 sg13g2_a21oi_1 _5749_ (.A1(_1115_),
    .A2(_1420_),
    .Y(_1421_),
    .B1(_0341_));
 sg13g2_nand2_1 _5750_ (.Y(_1422_),
    .A(_1035_),
    .B(_0996_));
 sg13g2_nand2_1 _5751_ (.Y(_1423_),
    .A(_1422_),
    .B(net33));
 sg13g2_nand3_1 _5752_ (.B(_1040_),
    .C(net54),
    .A(_1423_),
    .Y(_1424_));
 sg13g2_nand2b_1 _5753_ (.Y(_1425_),
    .B(_1424_),
    .A_N(_1421_));
 sg13g2_nand2_1 _5754_ (.Y(_1426_),
    .A(_1425_),
    .B(net34));
 sg13g2_nand2_1 _5755_ (.Y(_1427_),
    .A(_1221_),
    .B(net45));
 sg13g2_o21ai_1 _5756_ (.B1(net53),
    .Y(_1428_),
    .A1(_0928_),
    .A2(_1000_));
 sg13g2_nand2_1 _5757_ (.Y(_1429_),
    .A(_1427_),
    .B(_1428_));
 sg13g2_a21oi_1 _5758_ (.A1(_1429_),
    .A2(net49),
    .Y(_1430_),
    .B1(net37));
 sg13g2_nand2_1 _5759_ (.Y(_1431_),
    .A(_1426_),
    .B(_1430_));
 sg13g2_nand3_1 _5760_ (.B(_1216_),
    .C(_1148_),
    .A(_0820_),
    .Y(_1432_));
 sg13g2_nor2b_1 _5761_ (.A(net26),
    .B_N(_1432_),
    .Y(_1433_));
 sg13g2_nand2_1 _5762_ (.Y(_1434_),
    .A(_1431_),
    .B(_1433_));
 sg13g2_nand2_1 _5763_ (.Y(_1435_),
    .A(_1419_),
    .B(_1434_));
 sg13g2_nand2_1 _5764_ (.Y(_1436_),
    .A(_1435_),
    .B(_0883_));
 sg13g2_nand3_1 _5765_ (.B(_1273_),
    .C(net39),
    .A(_1428_),
    .Y(_1437_));
 sg13g2_nand2_1 _5766_ (.Y(_1438_),
    .A(_1437_),
    .B(net28));
 sg13g2_nand2b_1 _5767_ (.Y(_1439_),
    .B(net36),
    .A_N(_1410_));
 sg13g2_nand3_1 _5768_ (.B(net34),
    .C(_1213_),
    .A(_1439_),
    .Y(_1440_));
 sg13g2_nand2b_1 _5769_ (.Y(_1441_),
    .B(_1440_),
    .A_N(_1438_));
 sg13g2_nand2_1 _5770_ (.Y(_1442_),
    .A(_1016_),
    .B(_1037_));
 sg13g2_a21oi_1 _5771_ (.A1(_1327_),
    .A2(_1442_),
    .Y(_1443_),
    .B1(net32));
 sg13g2_nor2_1 _5772_ (.A(net55),
    .B(_1443_),
    .Y(_1444_));
 sg13g2_a21oi_1 _5773_ (.A1(_1441_),
    .A2(_1444_),
    .Y(_1445_),
    .B1(net26));
 sg13g2_nand3_1 _5774_ (.B(_1014_),
    .C(_1005_),
    .A(net33),
    .Y(_1446_));
 sg13g2_nand2_1 _5775_ (.Y(_1447_),
    .A(_1446_),
    .B(_1428_));
 sg13g2_a21oi_1 _5776_ (.A1(_1015_),
    .A2(net36),
    .Y(_1448_),
    .B1(net39));
 sg13g2_a22oi_1 _5777_ (.Y(_1449_),
    .B1(_1423_),
    .B2(_1448_),
    .A2(net40),
    .A1(_1447_));
 sg13g2_nor2_1 _5778_ (.A(_1021_),
    .B(_1084_),
    .Y(_1450_));
 sg13g2_o21ai_1 _5779_ (.B1(_0884_),
    .Y(_1451_),
    .A1(_1042_),
    .A2(_1450_));
 sg13g2_nor2b_1 _5780_ (.A(net54),
    .B_N(_1451_),
    .Y(_1452_));
 sg13g2_o21ai_1 _5781_ (.B1(_1452_),
    .Y(_1453_),
    .A1(net30),
    .A2(_1449_));
 sg13g2_nand2_1 _5782_ (.Y(_1454_),
    .A(_1445_),
    .B(_1453_));
 sg13g2_nand3_1 _5783_ (.B(_1409_),
    .C(net42),
    .A(net43),
    .Y(_1455_));
 sg13g2_nand2_1 _5784_ (.Y(_1456_),
    .A(_1272_),
    .B(net41));
 sg13g2_and2_1 _5785_ (.A(_1455_),
    .B(_1456_),
    .X(_1457_));
 sg13g2_nor2_1 _5786_ (.A(net35),
    .B(_1105_),
    .Y(_1458_));
 sg13g2_a21oi_1 _5787_ (.A1(_1457_),
    .A2(_1458_),
    .Y(_1459_),
    .B1(net55));
 sg13g2_a21oi_1 _5788_ (.A1(_1005_),
    .A2(net42),
    .Y(_1460_),
    .B1(_1000_));
 sg13g2_nor2_1 _5789_ (.A(net44),
    .B(_1460_),
    .Y(_1461_));
 sg13g2_nor2b_1 _5790_ (.A(_1461_),
    .B_N(_0909_),
    .Y(_1462_));
 sg13g2_nand2_1 _5791_ (.Y(_1463_),
    .A(_1462_),
    .B(net34));
 sg13g2_nand2_1 _5792_ (.Y(_1464_),
    .A(_1459_),
    .B(_1463_));
 sg13g2_nand2_1 _5793_ (.Y(_1465_),
    .A(_1364_),
    .B(_0887_));
 sg13g2_o21ai_1 _5794_ (.B1(_1465_),
    .Y(_1466_),
    .A1(net36),
    .A2(_1460_));
 sg13g2_a21oi_1 _5795_ (.A1(_1466_),
    .A2(_1329_),
    .Y(_1467_),
    .B1(net27));
 sg13g2_a21o_1 _5796_ (.A2(_1455_),
    .A1(_1359_),
    .B1(_0912_),
    .X(_1468_));
 sg13g2_nand3_1 _5797_ (.B(_1467_),
    .C(_1468_),
    .A(_1464_),
    .Y(_1469_));
 sg13g2_inv_1 _5798_ (.Y(_1470_),
    .A(_1107_));
 sg13g2_nor3_1 _5799_ (.A(net30),
    .B(_1152_),
    .C(_1470_),
    .Y(_1471_));
 sg13g2_nor2_1 _5800_ (.A(net25),
    .B(_1471_),
    .Y(_1472_));
 sg13g2_nand2_1 _5801_ (.Y(_1473_),
    .A(_1469_),
    .B(_1472_));
 sg13g2_nand2_1 _5802_ (.Y(_1474_),
    .A(_1454_),
    .B(_1473_));
 sg13g2_nand2_1 _5803_ (.Y(_1475_),
    .A(_1474_),
    .B(_1080_));
 sg13g2_a21oi_1 _5804_ (.A1(_1436_),
    .A2(_1475_),
    .Y(_1476_),
    .B1(_1191_));
 sg13g2_o21ai_1 _5805_ (.B1(_0826_),
    .Y(_1477_),
    .A1(net42),
    .A2(net45));
 sg13g2_nand2_1 _5806_ (.Y(_1478_),
    .A(_0926_),
    .B(_1477_));
 sg13g2_a21oi_1 _5807_ (.A1(_0894_),
    .A2(net45),
    .Y(_1479_),
    .B1(net51));
 sg13g2_nand2_1 _5808_ (.Y(_1480_),
    .A(_0887_),
    .B(_0701_));
 sg13g2_nand3_1 _5809_ (.B(_1083_),
    .C(net44),
    .A(_1480_),
    .Y(_1481_));
 sg13g2_nand2_1 _5810_ (.Y(_1482_),
    .A(_1479_),
    .B(_1481_));
 sg13g2_nand2_1 _5811_ (.Y(_1483_),
    .A(_1478_),
    .B(_1482_));
 sg13g2_a21oi_1 _5812_ (.A1(_1483_),
    .A2(net28),
    .Y(_1484_),
    .B1(_1443_));
 sg13g2_nor2_1 _5813_ (.A(_1098_),
    .B(_1484_),
    .Y(_1485_));
 sg13g2_nand3_1 _5814_ (.B(net49),
    .C(_1359_),
    .A(_1414_),
    .Y(_1486_));
 sg13g2_nand2_1 _5815_ (.Y(_1487_),
    .A(net48),
    .B(_1025_));
 sg13g2_nand2_1 _5816_ (.Y(_1488_),
    .A(_1365_),
    .B(_1487_));
 sg13g2_nand2_1 _5817_ (.Y(_1489_),
    .A(_1486_),
    .B(_1488_));
 sg13g2_a21oi_1 _5818_ (.A1(_0996_),
    .A2(_1006_),
    .Y(_1490_),
    .B1(net33));
 sg13g2_o21ai_1 _5819_ (.B1(net28),
    .Y(_1491_),
    .A1(_1152_),
    .A2(_1490_));
 sg13g2_inv_1 _5820_ (.Y(_1492_),
    .A(_1259_));
 sg13g2_a21oi_1 _5821_ (.A1(_1489_),
    .A2(_1491_),
    .Y(_1493_),
    .B1(_1492_));
 sg13g2_nor2_1 _5822_ (.A(_1485_),
    .B(_1493_),
    .Y(_1494_));
 sg13g2_inv_1 _5823_ (.Y(_1495_),
    .A(_1000_));
 sg13g2_nor2_1 _5824_ (.A(net52),
    .B(_1495_),
    .Y(_1496_));
 sg13g2_a21oi_1 _5825_ (.A1(_1496_),
    .A2(_1021_),
    .Y(_1497_),
    .B1(net47));
 sg13g2_nand2_1 _5826_ (.Y(_1498_),
    .A(_1497_),
    .B(_1427_));
 sg13g2_a21oi_1 _5827_ (.A1(_1272_),
    .A2(net41),
    .Y(_1499_),
    .B1(net51));
 sg13g2_nand2_1 _5828_ (.Y(_1500_),
    .A(_1084_),
    .B(net43));
 sg13g2_nand2_1 _5829_ (.Y(_1501_),
    .A(_1499_),
    .B(_1500_));
 sg13g2_nand3_1 _5830_ (.B(_1501_),
    .C(net32),
    .A(_1498_),
    .Y(_1502_));
 sg13g2_inv_1 _5831_ (.Y(_1503_),
    .A(_1202_));
 sg13g2_a21oi_1 _5832_ (.A1(_1502_),
    .A2(_1451_),
    .Y(_1504_),
    .B1(_1503_));
 sg13g2_nand3_1 _5833_ (.B(net49),
    .C(_1117_),
    .A(_1414_),
    .Y(_1505_));
 sg13g2_nand2b_1 _5834_ (.Y(_1506_),
    .B(net48),
    .A_N(_0924_));
 sg13g2_nand2_1 _5835_ (.Y(_1507_),
    .A(_1365_),
    .B(_1506_));
 sg13g2_nand2_1 _5836_ (.Y(_1508_),
    .A(_1505_),
    .B(_1507_));
 sg13g2_o21ai_1 _5837_ (.B1(net28),
    .Y(_1509_),
    .A1(_1152_),
    .A2(_1326_));
 sg13g2_a21oi_1 _5838_ (.A1(_1508_),
    .A2(_1509_),
    .Y(_1510_),
    .B1(_1112_));
 sg13g2_nor2_1 _5839_ (.A(_1504_),
    .B(_1510_),
    .Y(_1511_));
 sg13g2_nand2_1 _5840_ (.Y(_1512_),
    .A(_1494_),
    .B(_1511_));
 sg13g2_inv_1 _5841_ (.Y(_1513_),
    .A(_1321_));
 sg13g2_nand2_1 _5842_ (.Y(_1514_),
    .A(_1512_),
    .B(_1513_));
 sg13g2_o21ai_1 _5843_ (.B1(net32),
    .Y(_1515_),
    .A1(_1087_),
    .A2(_1274_));
 sg13g2_nand2_1 _5844_ (.Y(_1516_),
    .A(_1480_),
    .B(net41));
 sg13g2_nand3_1 _5845_ (.B(_1216_),
    .C(_1516_),
    .A(net31),
    .Y(_1517_));
 sg13g2_nand2_1 _5846_ (.Y(_1518_),
    .A(_1515_),
    .B(_1517_));
 sg13g2_nand2_1 _5847_ (.Y(_1519_),
    .A(_1518_),
    .B(net54));
 sg13g2_nor2_1 _5848_ (.A(_1462_),
    .B(_1112_),
    .Y(_1520_));
 sg13g2_nand3b_1 _5849_ (.B(_1122_),
    .C(_0996_),
    .Y(_1521_),
    .A_N(_0341_));
 sg13g2_a21oi_1 _5850_ (.A1(_1521_),
    .A2(_0989_),
    .Y(_1522_),
    .B1(net37));
 sg13g2_nor2_1 _5851_ (.A(_1520_),
    .B(_1522_),
    .Y(_1523_));
 sg13g2_nand2_1 _5852_ (.Y(_1524_),
    .A(_1519_),
    .B(_1523_));
 sg13g2_nand2_1 _5853_ (.Y(_1525_),
    .A(_1524_),
    .B(net34));
 sg13g2_nor2_1 _5854_ (.A(net31),
    .B(_1430_),
    .Y(_1526_));
 sg13g2_nand2_1 _5855_ (.Y(_1527_),
    .A(_1327_),
    .B(_1216_));
 sg13g2_o21ai_1 _5856_ (.B1(net33),
    .Y(_1528_),
    .A1(_0928_),
    .A2(_1106_));
 sg13g2_nand3_1 _5857_ (.B(_1037_),
    .C(net41),
    .A(_0924_),
    .Y(_1529_));
 sg13g2_nand4_1 _5858_ (.B(net37),
    .C(net39),
    .A(_1528_),
    .Y(_1530_),
    .D(_1529_));
 sg13g2_nor2_1 _5859_ (.A(net48),
    .B(_0989_),
    .Y(_1531_));
 sg13g2_o21ai_1 _5860_ (.B1(_1531_),
    .Y(_1532_),
    .A1(_1106_),
    .A2(_1470_));
 sg13g2_nand2_1 _5861_ (.Y(_1533_),
    .A(_1530_),
    .B(_1532_));
 sg13g2_a21oi_1 _5862_ (.A1(_1526_),
    .A2(_1527_),
    .Y(_1534_),
    .B1(_1533_));
 sg13g2_nand2_1 _5863_ (.Y(_1535_),
    .A(_1525_),
    .B(_1534_));
 sg13g2_nand2_1 _5864_ (.Y(_1536_),
    .A(_1535_),
    .B(_1081_));
 sg13g2_nand2_1 _5865_ (.Y(_1537_),
    .A(_1514_),
    .B(_1536_));
 sg13g2_nand2_1 _5866_ (.Y(_1538_),
    .A(_1537_),
    .B(net46));
 sg13g2_a22oi_1 _5867_ (.Y(_1539_),
    .B1(net33),
    .B2(_1084_),
    .A2(_0996_),
    .A1(_1120_));
 sg13g2_o21ai_1 _5868_ (.B1(_1430_),
    .Y(_1540_),
    .A1(net40),
    .A2(_1539_));
 sg13g2_a21oi_1 _5869_ (.A1(_1540_),
    .A2(_1432_),
    .Y(_1541_),
    .B1(net26));
 sg13g2_o21ai_1 _5870_ (.B1(_1222_),
    .Y(_1542_),
    .A1(net36),
    .A2(_1015_));
 sg13g2_nor2_1 _5871_ (.A(net36),
    .B(_0885_),
    .Y(_1543_));
 sg13g2_a21oi_1 _5872_ (.A1(_1460_),
    .A2(_1543_),
    .Y(_1544_),
    .B1(net27));
 sg13g2_nand2_1 _5873_ (.Y(_1545_),
    .A(_1542_),
    .B(_1544_));
 sg13g2_nor2_1 _5874_ (.A(net25),
    .B(_1408_),
    .Y(_1546_));
 sg13g2_a21oi_1 _5875_ (.A1(_1545_),
    .A2(_1546_),
    .Y(_1547_),
    .B1(_0881_));
 sg13g2_nor2b_1 _5876_ (.A(_1541_),
    .B_N(_1547_),
    .Y(_1548_));
 sg13g2_o21ai_1 _5877_ (.B1(_1320_),
    .Y(_1549_),
    .A1(_1192_),
    .A2(_1548_));
 sg13g2_nand2_1 _5878_ (.Y(_1550_),
    .A(_1538_),
    .B(_1549_));
 sg13g2_nor2_1 _5879_ (.A(_1476_),
    .B(_1550_),
    .Y(_1551_));
 sg13g2_nand2b_1 _5880_ (.Y(_1552_),
    .B(_0923_),
    .A_N(_1334_));
 sg13g2_nand2_1 _5881_ (.Y(_1553_),
    .A(_1351_),
    .B(_1147_));
 sg13g2_nor2b_1 _5882_ (.A(_1553_),
    .B_N(_1276_),
    .Y(_1554_));
 sg13g2_nand2b_1 _5883_ (.Y(_1555_),
    .B(_1554_),
    .A_N(_1326_));
 sg13g2_a21oi_1 _5884_ (.A1(_1552_),
    .A2(_1555_),
    .Y(_1556_),
    .B1(_1098_));
 sg13g2_nand2b_1 _5885_ (.Y(_1557_),
    .B(_0923_),
    .A_N(_1336_));
 sg13g2_nand2_1 _5886_ (.Y(_1558_),
    .A(_1554_),
    .B(_0899_));
 sg13g2_a21oi_1 _5887_ (.A1(_1557_),
    .A2(_1558_),
    .Y(_1559_),
    .B1(_1503_));
 sg13g2_nor3_1 _5888_ (.A(net46),
    .B(_1556_),
    .C(_1559_),
    .Y(_1560_));
 sg13g2_a21oi_1 _5889_ (.A1(_0897_),
    .A2(_1495_),
    .Y(_1561_),
    .B1(net45));
 sg13g2_nor3_1 _5890_ (.A(net35),
    .B(_1016_),
    .C(_1561_),
    .Y(_1562_));
 sg13g2_o21ai_1 _5891_ (.B1(_1093_),
    .Y(_1563_),
    .A1(_1562_),
    .A2(_1019_));
 sg13g2_nand2_1 _5892_ (.Y(_1564_),
    .A(_1041_),
    .B(_1044_));
 sg13g2_nand2_1 _5893_ (.Y(_1565_),
    .A(_1563_),
    .B(_1564_));
 sg13g2_nand2_1 _5894_ (.Y(_1566_),
    .A(_1565_),
    .B(_1248_));
 sg13g2_nand2_1 _5895_ (.Y(_1567_),
    .A(_1560_),
    .B(_1566_));
 sg13g2_o21ai_1 _5896_ (.B1(net32),
    .Y(_1568_),
    .A1(_1089_),
    .A2(net35));
 sg13g2_a21oi_1 _5897_ (.A1(net48),
    .A2(_1364_),
    .Y(_1569_),
    .B1(net55));
 sg13g2_o21ai_1 _5898_ (.B1(_1569_),
    .Y(_1570_),
    .A1(net32),
    .A2(_1276_));
 sg13g2_nand2_1 _5899_ (.Y(_1571_),
    .A(_1570_),
    .B(net25));
 sg13g2_o21ai_1 _5900_ (.B1(_1571_),
    .Y(_1572_),
    .A1(_1568_),
    .A2(_1265_));
 sg13g2_nor2b_1 _5901_ (.A(net35),
    .B_N(_1115_),
    .Y(_1573_));
 sg13g2_a21oi_1 _5902_ (.A1(_1121_),
    .A2(_1228_),
    .Y(_1574_),
    .B1(_1013_));
 sg13g2_o21ai_1 _5903_ (.B1(_1119_),
    .Y(_1575_),
    .A1(_1573_),
    .A2(_1574_));
 sg13g2_nor2_1 _5904_ (.A(net54),
    .B(_1348_),
    .Y(_1576_));
 sg13g2_nand2_1 _5905_ (.Y(_1577_),
    .A(_1575_),
    .B(_1576_));
 sg13g2_nand2_1 _5906_ (.Y(_1578_),
    .A(_1572_),
    .B(_1577_));
 sg13g2_a21oi_1 _5907_ (.A1(_1212_),
    .A2(_0707_),
    .Y(_1579_),
    .B1(_1561_));
 sg13g2_nand2_1 _5908_ (.Y(_1580_),
    .A(_1579_),
    .B(_1039_));
 sg13g2_nor2_1 _5909_ (.A(net32),
    .B(_0993_),
    .Y(_1581_));
 sg13g2_nand2_1 _5910_ (.Y(_1582_),
    .A(_1580_),
    .B(_1581_));
 sg13g2_nor2_1 _5911_ (.A(_1019_),
    .B(_1582_),
    .Y(_1583_));
 sg13g2_a21oi_1 _5912_ (.A1(_1228_),
    .A2(_1148_),
    .Y(_1584_),
    .B1(_0912_));
 sg13g2_nand3_1 _5913_ (.B(_1037_),
    .C(_1007_),
    .A(_0702_),
    .Y(_1585_));
 sg13g2_a21oi_1 _5914_ (.A1(_1420_),
    .A2(_1585_),
    .Y(_1586_),
    .B1(_1010_));
 sg13g2_nor3_1 _5915_ (.A(_1043_),
    .B(_1584_),
    .C(_1586_),
    .Y(_1587_));
 sg13g2_nor2b_1 _5916_ (.A(_1587_),
    .B_N(_1531_),
    .Y(_1588_));
 sg13g2_nor2_1 _5917_ (.A(_1583_),
    .B(_1588_),
    .Y(_1589_));
 sg13g2_nand2_1 _5918_ (.Y(_1590_),
    .A(_1578_),
    .B(_1589_));
 sg13g2_nand2_1 _5919_ (.Y(_1591_),
    .A(_1590_),
    .B(net46));
 sg13g2_nand2_1 _5920_ (.Y(_1592_),
    .A(_1567_),
    .B(_1591_));
 sg13g2_inv_1 _5921_ (.Y(_1593_),
    .A(_1320_));
 sg13g2_nand2_1 _5922_ (.Y(_1594_),
    .A(_1592_),
    .B(_1593_));
 sg13g2_nand2_1 _5923_ (.Y(_1595_),
    .A(_1594_),
    .B(_1418_));
 sg13g2_nand2_1 _5924_ (.Y(_1596_),
    .A(_1595_),
    .B(_1191_));
 sg13g2_a21oi_1 _5925_ (.A1(_1551_),
    .A2(_1596_),
    .Y(_1597_),
    .B1(_1404_));
 sg13g2_nor2_1 _5926_ (.A(_1406_),
    .B(_1597_),
    .Y(_0000_));
 sg13g2_inv_1 _5927_ (.Y(_1598_),
    .A(\center_x[0] ));
 sg13g2_buf_1 _5928_ (.A(_0838_),
    .X(_1599_));
 sg13g2_buf_1 _5929_ (.A(net123),
    .X(_1600_));
 sg13g2_nor2_2 _5930_ (.A(net123),
    .B(_3671_),
    .Y(_1601_));
 sg13g2_nor3_1 _5931_ (.A(_0047_),
    .B(net123),
    .C(_0650_),
    .Y(_1602_));
 sg13g2_a221oi_1 _5932_ (.B2(_3642_),
    .C1(_1602_),
    .B1(_1601_),
    .A1(_1598_),
    .Y(_0244_),
    .A2(net112));
 sg13g2_xnor2_1 _5933_ (.Y(_1603_),
    .A(_3641_),
    .B(_3638_));
 sg13g2_buf_1 _5934_ (.A(net147),
    .X(_1604_));
 sg13g2_nor2_1 _5935_ (.A(\center_x[1] ),
    .B(net132),
    .Y(_1605_));
 sg13g2_a21oi_1 _5936_ (.A1(_1603_),
    .A2(net132),
    .Y(_1606_),
    .B1(_1605_));
 sg13g2_nor2_1 _5937_ (.A(_1606_),
    .B(_1601_),
    .Y(_1607_));
 sg13g2_a21oi_1 _5938_ (.A1(_3639_),
    .A2(_1601_),
    .Y(_0245_),
    .B1(_1607_));
 sg13g2_inv_1 _5939_ (.Y(_1608_),
    .A(\center_x[2] ));
 sg13g2_nand2_1 _5940_ (.Y(_1609_),
    .A(_3641_),
    .B(_3638_));
 sg13g2_inv_1 _5941_ (.Y(_1610_),
    .A(\i_transform.track_x[2] ));
 sg13g2_o21ai_1 _5942_ (.B1(_1610_),
    .Y(_1611_),
    .A1(_1609_),
    .A2(_0650_));
 sg13g2_nand4_1 _5943_ (.B(_3641_),
    .C(_3638_),
    .A(_3671_),
    .Y(_1612_),
    .D(\i_transform.track_x[2] ));
 sg13g2_a21oi_1 _5944_ (.A1(_1611_),
    .A2(_1612_),
    .Y(_1613_),
    .B1(net112));
 sg13g2_a21oi_1 _5945_ (.A1(_1608_),
    .A2(net112),
    .Y(_0246_),
    .B1(_1613_));
 sg13g2_nor2_1 _5946_ (.A(_1610_),
    .B(_1609_),
    .Y(_1614_));
 sg13g2_inv_1 _5947_ (.Y(_1615_),
    .A(_1614_));
 sg13g2_nor2_1 _5948_ (.A(_3609_),
    .B(_1615_),
    .Y(_1616_));
 sg13g2_inv_1 _5949_ (.Y(_1617_),
    .A(_1616_));
 sg13g2_nand2_1 _5950_ (.Y(_1618_),
    .A(_1615_),
    .B(_3609_));
 sg13g2_nand3_1 _5951_ (.B(net132),
    .C(_1618_),
    .A(_1617_),
    .Y(_1619_));
 sg13g2_buf_1 _5952_ (.A(\center_x[3] ),
    .X(_1620_));
 sg13g2_a22oi_1 _5953_ (.Y(_1621_),
    .B1(\i_transform.track_x[3] ),
    .B2(_1601_),
    .A2(net112),
    .A1(_1620_));
 sg13g2_o21ai_1 _5954_ (.B1(_1621_),
    .Y(_0247_),
    .A1(_0959_),
    .A2(_1619_));
 sg13g2_nor2_1 _5955_ (.A(_3597_),
    .B(_1617_),
    .Y(_1622_));
 sg13g2_inv_1 _5956_ (.Y(_1623_),
    .A(_1622_));
 sg13g2_nand2_1 _5957_ (.Y(_1624_),
    .A(_1617_),
    .B(_3597_));
 sg13g2_nand3_1 _5958_ (.B(net132),
    .C(_1624_),
    .A(_1623_),
    .Y(_1625_));
 sg13g2_buf_1 _5959_ (.A(\center_x[4] ),
    .X(_1626_));
 sg13g2_a22oi_1 _5960_ (.Y(_1627_),
    .B1(\i_transform.track_x[4] ),
    .B2(_1601_),
    .A2(net112),
    .A1(_1626_));
 sg13g2_o21ai_1 _5961_ (.B1(_1627_),
    .Y(_0248_),
    .A1(_0959_),
    .A2(_1625_));
 sg13g2_buf_1 _5962_ (.A(net60),
    .X(_1628_));
 sg13g2_nor2_1 _5963_ (.A(_0044_),
    .B(net58),
    .Y(_1629_));
 sg13g2_inv_1 _5964_ (.Y(_1630_),
    .A(_3599_));
 sg13g2_nor2_1 _5965_ (.A(_1630_),
    .B(_1623_),
    .Y(_1631_));
 sg13g2_nor2_1 _5966_ (.A(_3599_),
    .B(_1622_),
    .Y(_1632_));
 sg13g2_o21ai_1 _5967_ (.B1(net58),
    .Y(_1633_),
    .A1(_1631_),
    .A2(_1632_));
 sg13g2_nand3_1 _5968_ (.B(net132),
    .C(_3652_),
    .A(_1633_),
    .Y(_1634_));
 sg13g2_buf_1 _5969_ (.A(\center_x[5] ),
    .X(_1635_));
 sg13g2_buf_1 _5970_ (.A(net123),
    .X(_1636_));
 sg13g2_nor2_2 _5971_ (.A(_0838_),
    .B(_0689_),
    .Y(_1637_));
 sg13g2_a22oi_1 _5972_ (.Y(_1638_),
    .B1(_3599_),
    .B2(_1637_),
    .A2(net111),
    .A1(_1635_));
 sg13g2_o21ai_1 _5973_ (.B1(_1638_),
    .Y(_0249_),
    .A1(_1629_),
    .A2(_1634_));
 sg13g2_nand2_2 _5974_ (.Y(_1639_),
    .A(_0689_),
    .B(net132));
 sg13g2_buf_1 _5975_ (.A(_3885_),
    .X(_1640_));
 sg13g2_nor2b_1 _5976_ (.A(_3885_),
    .B_N(_1631_),
    .Y(_1641_));
 sg13g2_a21oi_1 _5977_ (.A1(_1630_),
    .A2(net59),
    .Y(_1642_),
    .B1(_1641_));
 sg13g2_xnor2_1 _5978_ (.Y(_1643_),
    .A(_3632_),
    .B(_1642_));
 sg13g2_buf_1 _5979_ (.A(\center_x[6] ),
    .X(_1644_));
 sg13g2_a22oi_1 _5980_ (.Y(_1645_),
    .B1(_3631_),
    .B2(_1637_),
    .A2(net111),
    .A1(_1644_));
 sg13g2_o21ai_1 _5981_ (.B1(_1645_),
    .Y(_0250_),
    .A1(_1639_),
    .A2(_1643_));
 sg13g2_a22oi_1 _5982_ (.Y(_1646_),
    .B1(_3631_),
    .B2(_1641_),
    .A2(net59),
    .A1(_3657_));
 sg13g2_xnor2_1 _5983_ (.Y(_1647_),
    .A(_3658_),
    .B(_1646_));
 sg13g2_buf_2 _5984_ (.A(\center_x[7] ),
    .X(_1648_));
 sg13g2_a22oi_1 _5985_ (.Y(_1649_),
    .B1(_3626_),
    .B2(_1637_),
    .A2(net111),
    .A1(_1648_));
 sg13g2_o21ai_1 _5986_ (.B1(_1649_),
    .Y(_0251_),
    .A1(_1639_),
    .A2(_1647_));
 sg13g2_nand2_1 _5987_ (.Y(_1650_),
    .A(_1641_),
    .B(_3631_));
 sg13g2_a22oi_1 _5988_ (.Y(_1651_),
    .B1(_3659_),
    .B2(_1650_),
    .A2(net58),
    .A1(_3658_));
 sg13g2_xnor2_1 _5989_ (.Y(_1652_),
    .A(_3615_),
    .B(_1651_));
 sg13g2_buf_1 _5990_ (.A(\center_x[8] ),
    .X(_1653_));
 sg13g2_a22oi_1 _5991_ (.Y(_1654_),
    .B1(_3615_),
    .B2(_1637_),
    .A2(_1636_),
    .A1(_1653_));
 sg13g2_o21ai_1 _5992_ (.B1(_1654_),
    .Y(_0252_),
    .A1(_1639_),
    .A2(_1652_));
 sg13g2_nand2_1 _5993_ (.Y(_1655_),
    .A(net59),
    .B(_3660_));
 sg13g2_nor3_1 _5994_ (.A(_3658_),
    .B(_3616_),
    .C(_1650_),
    .Y(_1656_));
 sg13g2_a21oi_1 _5995_ (.A1(_3619_),
    .A2(_1655_),
    .Y(_1657_),
    .B1(_1656_));
 sg13g2_a22oi_1 _5996_ (.Y(_1658_),
    .B1(_3619_),
    .B2(_1637_),
    .A2(_1636_),
    .A1(\center_x[9] ));
 sg13g2_o21ai_1 _5997_ (.B1(_1658_),
    .Y(_0253_),
    .A1(_1639_),
    .A2(_1657_));
 sg13g2_inv_1 _5998_ (.Y(_1659_),
    .A(\center_y[0] ));
 sg13g2_nor2_2 _5999_ (.A(net123),
    .B(_0841_),
    .Y(_1660_));
 sg13g2_inv_1 _6000_ (.Y(_1661_),
    .A(_3583_));
 sg13g2_nor2_1 _6001_ (.A(_0838_),
    .B(net83),
    .Y(_1662_));
 sg13g2_inv_1 _6002_ (.Y(_1663_),
    .A(_1662_));
 sg13g2_buf_8 _6003_ (.A(net74),
    .X(_1664_));
 sg13g2_nor3_1 _6004_ (.A(_0045_),
    .B(_1663_),
    .C(_1664_),
    .Y(_1665_));
 sg13g2_a221oi_1 _6005_ (.B2(_1661_),
    .C1(_1665_),
    .B1(_1660_),
    .A1(_1659_),
    .Y(_0254_),
    .A2(net112));
 sg13g2_inv_1 _6006_ (.Y(_1666_),
    .A(\center_y[1] ));
 sg13g2_inv_1 _6007_ (.Y(_1667_),
    .A(_3581_));
 sg13g2_xor2_1 _6008_ (.B(_3581_),
    .A(_3583_),
    .X(_1668_));
 sg13g2_nor3_1 _6009_ (.A(net123),
    .B(_1668_),
    .C(_0842_),
    .Y(_1669_));
 sg13g2_a221oi_1 _6010_ (.B2(_1667_),
    .C1(_1669_),
    .B1(_1660_),
    .A1(_1666_),
    .Y(_0255_),
    .A2(_1600_));
 sg13g2_inv_1 _6011_ (.Y(_1670_),
    .A(\center_y[2] ));
 sg13g2_nand2_1 _6012_ (.Y(_1671_),
    .A(_3583_),
    .B(_3581_));
 sg13g2_nand2_1 _6013_ (.Y(_1672_),
    .A(_1671_),
    .B(_3553_));
 sg13g2_nor2_1 _6014_ (.A(_3553_),
    .B(_1671_),
    .Y(_1673_));
 sg13g2_inv_1 _6015_ (.Y(_1674_),
    .A(_1673_));
 sg13g2_a221oi_1 _6016_ (.B2(_0317_),
    .C1(_1663_),
    .B1(_0315_),
    .A1(_1672_),
    .Y(_1675_),
    .A2(_1674_));
 sg13g2_a221oi_1 _6017_ (.B2(_3553_),
    .C1(_1675_),
    .B1(_1660_),
    .A1(_1670_),
    .Y(_0256_),
    .A2(_1600_));
 sg13g2_inv_1 _6018_ (.Y(_1676_),
    .A(\i_transform.track_y[3] ));
 sg13g2_nor2_1 _6019_ (.A(_1676_),
    .B(_1674_),
    .Y(_1677_));
 sg13g2_inv_1 _6020_ (.Y(_1678_),
    .A(_1677_));
 sg13g2_nand2_1 _6021_ (.Y(_1679_),
    .A(_1674_),
    .B(_1676_));
 sg13g2_nand3_1 _6022_ (.B(_1604_),
    .C(_1679_),
    .A(_1678_),
    .Y(_1680_));
 sg13g2_a22oi_1 _6023_ (.Y(_1681_),
    .B1(\i_transform.track_y[3] ),
    .B2(_1660_),
    .A2(net111),
    .A1(\center_y[3] ));
 sg13g2_o21ai_1 _6024_ (.B1(_1681_),
    .Y(_0257_),
    .A1(_0842_),
    .A2(_1680_));
 sg13g2_nor2_1 _6025_ (.A(_3571_),
    .B(_1678_),
    .Y(_1682_));
 sg13g2_inv_1 _6026_ (.Y(_1683_),
    .A(_1682_));
 sg13g2_nand2_1 _6027_ (.Y(_1684_),
    .A(_1678_),
    .B(_3571_));
 sg13g2_nand3_1 _6028_ (.B(_1604_),
    .C(_1684_),
    .A(_1683_),
    .Y(_1685_));
 sg13g2_buf_1 _6029_ (.A(\center_y[4] ),
    .X(_1686_));
 sg13g2_a22oi_1 _6030_ (.Y(_1687_),
    .B1(\i_transform.track_y[4] ),
    .B2(_1660_),
    .A2(net111),
    .A1(_1686_));
 sg13g2_o21ai_1 _6031_ (.B1(_1687_),
    .Y(_0258_),
    .A1(_0842_),
    .A2(_1685_));
 sg13g2_buf_1 _6032_ (.A(net77),
    .X(_1688_));
 sg13g2_nor2_1 _6033_ (.A(_0060_),
    .B(net73),
    .Y(_1689_));
 sg13g2_nor2b_1 _6034_ (.A(_1683_),
    .B_N(_0308_),
    .Y(_1690_));
 sg13g2_nor2_1 _6035_ (.A(_0308_),
    .B(_1682_),
    .Y(_1691_));
 sg13g2_o21ai_1 _6036_ (.B1(net73),
    .Y(_1692_),
    .A1(_1690_),
    .A2(_1691_));
 sg13g2_nand2_1 _6037_ (.Y(_1693_),
    .A(_1692_),
    .B(_1662_));
 sg13g2_buf_1 _6038_ (.A(\center_y[5] ),
    .X(_1694_));
 sg13g2_nor2_2 _6039_ (.A(_1599_),
    .B(_3592_),
    .Y(_1695_));
 sg13g2_a22oi_1 _6040_ (.Y(_1696_),
    .B1(_0308_),
    .B2(_1695_),
    .A2(net111),
    .A1(_1694_));
 sg13g2_o21ai_1 _6041_ (.B1(_1696_),
    .Y(_0259_),
    .A1(_1689_),
    .A2(_1693_));
 sg13g2_nor2_1 _6042_ (.A(_0308_),
    .B(net73),
    .Y(_1697_));
 sg13g2_a21oi_1 _6043_ (.A1(_1688_),
    .A2(_1690_),
    .Y(_1698_),
    .B1(_1697_));
 sg13g2_xnor2_1 _6044_ (.Y(_1699_),
    .A(_3567_),
    .B(_1698_));
 sg13g2_buf_1 _6045_ (.A(\center_y[6] ),
    .X(_1700_));
 sg13g2_a22oi_1 _6046_ (.Y(_1701_),
    .B1(_3565_),
    .B2(_1695_),
    .A2(net111),
    .A1(_1700_));
 sg13g2_o21ai_1 _6047_ (.B1(_1701_),
    .Y(_0260_),
    .A1(_1663_),
    .A2(_1699_));
 sg13g2_nand3_1 _6048_ (.B(_3565_),
    .C(_1690_),
    .A(_0320_),
    .Y(_1702_));
 sg13g2_inv_1 _6049_ (.Y(_1703_),
    .A(_1702_));
 sg13g2_a21oi_1 _6050_ (.A1(_0309_),
    .A2(net70),
    .Y(_1704_),
    .B1(_1703_));
 sg13g2_xnor2_1 _6051_ (.Y(_1705_),
    .A(_0310_),
    .B(_1704_));
 sg13g2_buf_2 _6052_ (.A(\center_y[7] ),
    .X(_1706_));
 sg13g2_a22oi_1 _6053_ (.Y(_1707_),
    .B1(\i_transform.track_y[7] ),
    .B2(_1695_),
    .A2(net111),
    .A1(_1706_));
 sg13g2_o21ai_1 _6054_ (.B1(_1707_),
    .Y(_0261_),
    .A1(_1663_),
    .A2(_1705_));
 sg13g2_a22oi_1 _6055_ (.Y(_1708_),
    .B1(_0311_),
    .B2(_1702_),
    .A2(_1688_),
    .A1(_0310_));
 sg13g2_xnor2_1 _6056_ (.Y(_1709_),
    .A(_3556_),
    .B(_1708_));
 sg13g2_buf_1 _6057_ (.A(\center_y[8] ),
    .X(_1710_));
 sg13g2_a22oi_1 _6058_ (.Y(_1711_),
    .B1(_3556_),
    .B2(_1695_),
    .A2(_1599_),
    .A1(_1710_));
 sg13g2_o21ai_1 _6059_ (.B1(_1711_),
    .Y(_0262_),
    .A1(_1663_),
    .A2(_1709_));
 sg13g2_inv_1 _6060_ (.Y(_1712_),
    .A(\center_y[9] ));
 sg13g2_buf_1 _6061_ (.A(net132),
    .X(_1713_));
 sg13g2_inv_1 _6062_ (.Y(_1714_),
    .A(\i_transform.track_y[9] ));
 sg13g2_nand3_1 _6063_ (.B(_3556_),
    .C(\i_transform.track_y[7] ),
    .A(_1703_),
    .Y(_1715_));
 sg13g2_a22oi_1 _6064_ (.Y(_1716_),
    .B1(_1714_),
    .B2(_1715_),
    .A2(_1664_),
    .A1(_0312_));
 sg13g2_nand2_1 _6065_ (.Y(_1717_),
    .A(_1716_),
    .B(_1662_));
 sg13g2_o21ai_1 _6066_ (.B1(_1717_),
    .Y(_0263_),
    .A1(_1712_),
    .A2(net122));
 sg13g2_inv_1 _6067_ (.Y(_1718_),
    .A(_3510_));
 sg13g2_inv_1 _6068_ (.Y(_1719_),
    .A(\i_orchestrator.vga_x[7] ));
 sg13g2_nand2_1 _6069_ (.Y(_1720_),
    .A(_1719_),
    .B(_3537_));
 sg13g2_nor4_1 _6070_ (.A(_3538_),
    .B(_3541_),
    .C(_3535_),
    .D(_1720_),
    .Y(_1721_));
 sg13g2_nand2_1 _6071_ (.Y(_1722_),
    .A(\i_orchestrator.vga_x[0] ),
    .B(\i_orchestrator.vga_x[1] ));
 sg13g2_nor2_1 _6072_ (.A(_3605_),
    .B(_1722_),
    .Y(_1723_));
 sg13g2_nand2_1 _6073_ (.Y(_1724_),
    .A(_1723_),
    .B(_3608_));
 sg13g2_inv_1 _6074_ (.Y(_1725_),
    .A(_1724_));
 sg13g2_nand2_1 _6075_ (.Y(_1726_),
    .A(_1721_),
    .B(_1725_));
 sg13g2_nand2_1 _6076_ (.Y(_1727_),
    .A(_1726_),
    .B(_3481_));
 sg13g2_buf_1 _6077_ (.A(_1727_),
    .X(_1728_));
 sg13g2_nor4_1 _6078_ (.A(_3505_),
    .B(_3506_),
    .C(_3525_),
    .D(_3501_),
    .Y(_1729_));
 sg13g2_nor3_1 _6079_ (.A(_3509_),
    .B(_3510_),
    .C(_3530_),
    .Y(_1730_));
 sg13g2_nand4_1 _6080_ (.B(_3521_),
    .C(_3504_),
    .A(_1729_),
    .Y(_1731_),
    .D(_1730_));
 sg13g2_nand2_1 _6081_ (.Y(_1732_),
    .A(_1731_),
    .B(_3481_));
 sg13g2_nor2_1 _6082_ (.A(_1726_),
    .B(_1732_),
    .Y(_1733_));
 sg13g2_nand2_1 _6083_ (.Y(_1734_),
    .A(_1733_),
    .B(_0064_));
 sg13g2_o21ai_1 _6084_ (.B1(_1734_),
    .Y(_0274_),
    .A1(_1718_),
    .A2(net97));
 sg13g2_xnor2_1 _6085_ (.Y(_1735_),
    .A(_3509_),
    .B(_3510_));
 sg13g2_inv_1 _6086_ (.Y(_1736_),
    .A(_1733_));
 sg13g2_inv_1 _6087_ (.Y(_1737_),
    .A(_1727_));
 sg13g2_nand2_1 _6088_ (.Y(_1738_),
    .A(net96),
    .B(_3509_));
 sg13g2_o21ai_1 _6089_ (.B1(_1738_),
    .Y(_0275_),
    .A1(_1735_),
    .A2(_1736_));
 sg13g2_nand2b_1 _6090_ (.Y(_1739_),
    .B(net97),
    .A_N(_3511_));
 sg13g2_nor2_1 _6091_ (.A(_3513_),
    .B(_3511_),
    .Y(_1740_));
 sg13g2_o21ai_1 _6092_ (.B1(_1727_),
    .Y(_1741_),
    .A1(_1740_),
    .A2(_1732_));
 sg13g2_inv_1 _6093_ (.Y(_1742_),
    .A(_1741_));
 sg13g2_a21oi_1 _6094_ (.A1(_3513_),
    .A2(_1739_),
    .Y(_0276_),
    .B1(_1742_));
 sg13g2_nand2_1 _6095_ (.Y(_1743_),
    .A(_1740_),
    .B(_3515_));
 sg13g2_nand2_1 _6096_ (.Y(_1744_),
    .A(_1741_),
    .B(net182));
 sg13g2_o21ai_1 _6097_ (.B1(_1744_),
    .Y(_0277_),
    .A1(_1736_),
    .A2(_1743_));
 sg13g2_nor2_1 _6098_ (.A(_3511_),
    .B(_3530_),
    .Y(_1745_));
 sg13g2_inv_1 _6099_ (.Y(_1746_),
    .A(_1745_));
 sg13g2_nor2_1 _6100_ (.A(_3526_),
    .B(_1746_),
    .Y(_1747_));
 sg13g2_inv_1 _6101_ (.Y(_1748_),
    .A(_1747_));
 sg13g2_nor2_1 _6102_ (.A(_1748_),
    .B(net96),
    .Y(_1749_));
 sg13g2_a21oi_1 _6103_ (.A1(net97),
    .A2(_1745_),
    .Y(_1750_),
    .B1(_3525_));
 sg13g2_inv_1 _6104_ (.Y(_1751_),
    .A(_1732_));
 sg13g2_nor2_1 _6105_ (.A(_1737_),
    .B(_1751_),
    .Y(_1752_));
 sg13g2_nor3_1 _6106_ (.A(_1749_),
    .B(_1750_),
    .C(_1752_),
    .Y(_0278_));
 sg13g2_nor2_1 _6107_ (.A(_3502_),
    .B(_1748_),
    .Y(_1753_));
 sg13g2_inv_1 _6108_ (.Y(_1754_),
    .A(_1753_));
 sg13g2_nor2_1 _6109_ (.A(_1754_),
    .B(net96),
    .Y(_1755_));
 sg13g2_nor2_1 _6110_ (.A(_3501_),
    .B(_1749_),
    .Y(_1756_));
 sg13g2_nor3_1 _6111_ (.A(_1755_),
    .B(_1756_),
    .C(_1752_),
    .Y(_0279_));
 sg13g2_nor3_1 _6112_ (.A(_3564_),
    .B(_1754_),
    .C(net96),
    .Y(_1757_));
 sg13g2_nor2_1 _6113_ (.A(_3506_),
    .B(_1755_),
    .Y(_1758_));
 sg13g2_nor3_1 _6114_ (.A(_1757_),
    .B(_1758_),
    .C(_1752_),
    .Y(_0280_));
 sg13g2_nor2_1 _6115_ (.A(_3505_),
    .B(_1757_),
    .Y(_1759_));
 sg13g2_nor2_1 _6116_ (.A(_3507_),
    .B(_1754_),
    .Y(_1760_));
 sg13g2_inv_1 _6117_ (.Y(_1761_),
    .A(_1760_));
 sg13g2_a21oi_1 _6118_ (.A1(_1751_),
    .A2(_1761_),
    .Y(_1762_),
    .B1(net96));
 sg13g2_nor2_1 _6119_ (.A(_1759_),
    .B(_1762_),
    .Y(_0281_));
 sg13g2_nor2_1 _6120_ (.A(_3504_),
    .B(_1761_),
    .Y(_1763_));
 sg13g2_o21ai_1 _6121_ (.B1(_1733_),
    .Y(_1764_),
    .A1(_3503_),
    .A2(_1760_));
 sg13g2_nand2_1 _6122_ (.Y(_1765_),
    .A(net96),
    .B(_3503_));
 sg13g2_o21ai_1 _6123_ (.B1(_1765_),
    .Y(_0282_),
    .A1(_1763_),
    .A2(_1764_));
 sg13g2_xnor2_1 _6124_ (.Y(_1766_),
    .A(_3521_),
    .B(_1763_));
 sg13g2_nand2_1 _6125_ (.Y(_1767_),
    .A(net96),
    .B(_3521_));
 sg13g2_o21ai_1 _6126_ (.B1(_1767_),
    .Y(_0283_),
    .A1(_1736_),
    .A2(_1766_));
 sg13g2_buf_1 _6127_ (.A(\i_capsule.tf_x[9] ),
    .X(_1768_));
 sg13g2_xnor2_1 _6128_ (.Y(_1769_),
    .A(net180),
    .B(_0607_));
 sg13g2_inv_1 _6129_ (.Y(_1770_),
    .A(\i_capsule.tf_x[9] ));
 sg13g2_nor2_1 _6130_ (.A(_0730_),
    .B(_1770_),
    .Y(_1771_));
 sg13g2_nor2_1 _6131_ (.A(_1768_),
    .B(_0974_),
    .Y(_1772_));
 sg13g2_nor2_2 _6132_ (.A(_1771_),
    .B(_1772_),
    .Y(_1773_));
 sg13g2_nor2_1 _6133_ (.A(_1769_),
    .B(_1773_),
    .Y(_1774_));
 sg13g2_buf_1 _6134_ (.A(_1774_),
    .X(_1775_));
 sg13g2_inv_1 _6135_ (.Y(_1776_),
    .A(net110));
 sg13g2_xnor2_1 _6136_ (.Y(_1777_),
    .A(net180),
    .B(_0403_));
 sg13g2_nor2_2 _6137_ (.A(_1777_),
    .B(_1773_),
    .Y(_1778_));
 sg13g2_inv_1 _6138_ (.Y(_1779_),
    .A(_1773_));
 sg13g2_xor2_1 _6139_ (.B(_0349_),
    .A(net180),
    .X(_1780_));
 sg13g2_nand2_1 _6140_ (.Y(_1781_),
    .A(_1779_),
    .B(_1780_));
 sg13g2_inv_1 _6141_ (.Y(_1782_),
    .A(_1781_));
 sg13g2_nor2_1 _6142_ (.A(_1778_),
    .B(_1782_),
    .Y(_1783_));
 sg13g2_nor2_1 _6143_ (.A(_1776_),
    .B(_1783_),
    .Y(_1784_));
 sg13g2_inv_1 _6144_ (.Y(_1785_),
    .A(_1784_));
 sg13g2_xnor2_1 _6145_ (.Y(_1786_),
    .A(net180),
    .B(_0720_));
 sg13g2_nor2_1 _6146_ (.A(_1786_),
    .B(_1773_),
    .Y(_1787_));
 sg13g2_buf_2 _6147_ (.A(_1787_),
    .X(_1788_));
 sg13g2_inv_1 _6148_ (.Y(_1789_),
    .A(_1788_));
 sg13g2_inv_1 _6149_ (.Y(_1790_),
    .A(_1772_));
 sg13g2_nor2_1 _6150_ (.A(_0722_),
    .B(_1771_),
    .Y(_1791_));
 sg13g2_a21oi_2 _6151_ (.B1(_1791_),
    .Y(_1792_),
    .A2(_1790_),
    .A1(_0722_));
 sg13g2_inv_1 _6152_ (.Y(_1793_),
    .A(_1792_));
 sg13g2_a21oi_1 _6153_ (.A1(_1785_),
    .A2(net95),
    .Y(_1794_),
    .B1(_1793_));
 sg13g2_nor2_1 _6154_ (.A(_1777_),
    .B(_1781_),
    .Y(_1795_));
 sg13g2_nor2_1 _6155_ (.A(_1776_),
    .B(_1795_),
    .Y(_1796_));
 sg13g2_nand2_1 _6156_ (.Y(_1797_),
    .A(_1796_),
    .B(_1788_));
 sg13g2_buf_1 _6157_ (.A(\i_capsule.tf_y[9] ),
    .X(_1798_));
 sg13g2_xnor2_1 _6158_ (.Y(_1799_),
    .A(net179),
    .B(_1161_));
 sg13g2_inv_1 _6159_ (.Y(_1800_),
    .A(_1799_));
 sg13g2_a21oi_1 _6160_ (.A1(_1794_),
    .A2(_1797_),
    .Y(_1801_),
    .B1(_1800_));
 sg13g2_nor3_1 _6161_ (.A(net95),
    .B(_1776_),
    .C(_1793_),
    .Y(_1802_));
 sg13g2_xor2_1 _6162_ (.B(_1291_),
    .A(net179),
    .X(_1803_));
 sg13g2_nand2_1 _6163_ (.Y(_1804_),
    .A(_1802_),
    .B(_1803_));
 sg13g2_nand3_1 _6164_ (.B(_1797_),
    .C(_1800_),
    .A(_1794_),
    .Y(_1805_));
 sg13g2_nand3b_1 _6165_ (.B(_1804_),
    .C(_1805_),
    .Y(_1806_),
    .A_N(_1801_));
 sg13g2_xnor2_1 _6166_ (.Y(_1807_),
    .A(_1768_),
    .B(_0357_));
 sg13g2_nor2_1 _6167_ (.A(_1807_),
    .B(_1773_),
    .Y(_1808_));
 sg13g2_inv_1 _6168_ (.Y(_1809_),
    .A(_1808_));
 sg13g2_nand2_1 _6169_ (.Y(_1810_),
    .A(_1809_),
    .B(_1781_));
 sg13g2_nand2_1 _6170_ (.Y(_1811_),
    .A(_1810_),
    .B(_1778_));
 sg13g2_inv_1 _6171_ (.Y(_1812_),
    .A(_1783_));
 sg13g2_a21oi_1 _6172_ (.A1(_1811_),
    .A2(_1812_),
    .Y(_1813_),
    .B1(net110));
 sg13g2_nand2_1 _6173_ (.Y(_1814_),
    .A(net110),
    .B(_1780_));
 sg13g2_nand2b_1 _6174_ (.Y(_1815_),
    .B(_1814_),
    .A_N(_1813_));
 sg13g2_nand2_1 _6175_ (.Y(_1816_),
    .A(_1815_),
    .B(net95));
 sg13g2_inv_1 _6176_ (.Y(_1817_),
    .A(_1778_));
 sg13g2_nor2_1 _6177_ (.A(_1808_),
    .B(_1817_),
    .Y(_1818_));
 sg13g2_nor3_1 _6178_ (.A(_1795_),
    .B(_1818_),
    .C(_1783_),
    .Y(_1819_));
 sg13g2_nor2_1 _6179_ (.A(net110),
    .B(_1819_),
    .Y(_1820_));
 sg13g2_inv_1 _6180_ (.Y(_1821_),
    .A(_1820_));
 sg13g2_nor2_1 _6181_ (.A(_1778_),
    .B(_1809_),
    .Y(_1822_));
 sg13g2_nor2_1 _6182_ (.A(_1817_),
    .B(_1810_),
    .Y(_1823_));
 sg13g2_o21ai_1 _6183_ (.B1(net110),
    .Y(_1824_),
    .A1(_1822_),
    .A2(_1823_));
 sg13g2_nand3_1 _6184_ (.B(_1788_),
    .C(_1824_),
    .A(_1821_),
    .Y(_1825_));
 sg13g2_nand3_1 _6185_ (.B(_1825_),
    .C(_1792_),
    .A(_1816_),
    .Y(_1826_));
 sg13g2_nand2_1 _6186_ (.Y(_1827_),
    .A(_1808_),
    .B(_1780_));
 sg13g2_nor2_1 _6187_ (.A(_1817_),
    .B(_1827_),
    .Y(_1828_));
 sg13g2_nand2_1 _6188_ (.Y(_1829_),
    .A(_1811_),
    .B(_1776_));
 sg13g2_o21ai_1 _6189_ (.B1(_1829_),
    .Y(_1830_),
    .A1(_1828_),
    .A2(_1785_));
 sg13g2_nand2_1 _6190_ (.Y(_1831_),
    .A(_1795_),
    .B(net110));
 sg13g2_a21oi_1 _6191_ (.A1(_1831_),
    .A2(net95),
    .Y(_1832_),
    .B1(_1792_));
 sg13g2_o21ai_1 _6192_ (.B1(_1832_),
    .Y(_1833_),
    .A1(net95),
    .A2(_1830_));
 sg13g2_xnor2_1 _6193_ (.Y(_1834_),
    .A(_1798_),
    .B(_3889_));
 sg13g2_a21oi_1 _6194_ (.A1(_1826_),
    .A2(_1833_),
    .Y(_1835_),
    .B1(_1834_));
 sg13g2_xnor2_1 _6195_ (.Y(_1836_),
    .A(_1798_),
    .B(_3773_));
 sg13g2_o21ai_1 _6196_ (.B1(net110),
    .Y(_1837_),
    .A1(_1822_),
    .A2(_1828_));
 sg13g2_a21oi_1 _6197_ (.A1(_1821_),
    .A2(_1837_),
    .Y(_1838_),
    .B1(_1788_));
 sg13g2_nand2_1 _6198_ (.Y(_1839_),
    .A(_1810_),
    .B(_1827_));
 sg13g2_nand2_1 _6199_ (.Y(_1840_),
    .A(_1839_),
    .B(_1778_));
 sg13g2_nor2_1 _6200_ (.A(net110),
    .B(_1822_),
    .Y(_1841_));
 sg13g2_a221oi_1 _6201_ (.B2(_1841_),
    .C1(_1789_),
    .B1(_1840_),
    .A1(_1775_),
    .Y(_1842_),
    .A2(_1818_));
 sg13g2_nor3_1 _6202_ (.A(_1793_),
    .B(_1838_),
    .C(_1842_),
    .Y(_1843_));
 sg13g2_nor2_1 _6203_ (.A(net95),
    .B(_1813_),
    .Y(_1844_));
 sg13g2_o21ai_1 _6204_ (.B1(_1784_),
    .Y(_1845_),
    .A1(_1817_),
    .A2(_1839_));
 sg13g2_a221oi_1 _6205_ (.B2(_1845_),
    .C1(_1792_),
    .B1(_1844_),
    .A1(net95),
    .Y(_1846_),
    .A2(_1796_));
 sg13g2_nor3_1 _6206_ (.A(_1836_),
    .B(_1843_),
    .C(_1846_),
    .Y(_1847_));
 sg13g2_xnor2_1 _6207_ (.Y(_1848_),
    .A(\i_capsule.tf_y[9] ),
    .B(_0843_));
 sg13g2_inv_1 _6208_ (.Y(_1849_),
    .A(_1848_));
 sg13g2_o21ai_1 _6209_ (.B1(_1829_),
    .Y(_1850_),
    .A1(_1795_),
    .A2(_1785_));
 sg13g2_a21oi_1 _6210_ (.A1(_1850_),
    .A2(net95),
    .Y(_1851_),
    .B1(_1793_));
 sg13g2_o21ai_1 _6211_ (.B1(_1844_),
    .Y(_1852_),
    .A1(_1785_),
    .A2(_1818_));
 sg13g2_nand2_1 _6212_ (.Y(_1853_),
    .A(_1851_),
    .B(_1852_));
 sg13g2_nor3_1 _6213_ (.A(_1776_),
    .B(_1817_),
    .C(_1827_),
    .Y(_1854_));
 sg13g2_nor2_1 _6214_ (.A(_1792_),
    .B(_1854_),
    .Y(_1855_));
 sg13g2_nand3_1 _6215_ (.B(_1788_),
    .C(_1829_),
    .A(_1855_),
    .Y(_1856_));
 sg13g2_nand2_1 _6216_ (.Y(_1857_),
    .A(_1853_),
    .B(_1856_));
 sg13g2_nor2_1 _6217_ (.A(_1849_),
    .B(_1857_),
    .Y(_1858_));
 sg13g2_nand3_1 _6218_ (.B(_1834_),
    .C(_1833_),
    .A(_1826_),
    .Y(_1859_));
 sg13g2_nor2b_1 _6219_ (.A(_1858_),
    .B_N(_1859_),
    .Y(_1860_));
 sg13g2_o21ai_1 _6220_ (.B1(_1860_),
    .Y(_1861_),
    .A1(_1835_),
    .A2(_1847_));
 sg13g2_nand2_1 _6221_ (.Y(_1862_),
    .A(_1854_),
    .B(_1788_));
 sg13g2_nand3_1 _6222_ (.B(_1788_),
    .C(_1814_),
    .A(_1812_),
    .Y(_1863_));
 sg13g2_a22oi_1 _6223_ (.Y(_1864_),
    .B1(_1863_),
    .B2(_1794_),
    .A2(_1793_),
    .A1(_1862_));
 sg13g2_xor2_1 _6224_ (.B(_1067_),
    .A(net179),
    .X(_1865_));
 sg13g2_a22oi_1 _6225_ (.Y(_1866_),
    .B1(_1849_),
    .B2(_1857_),
    .A2(_1865_),
    .A1(_1864_));
 sg13g2_nor2_1 _6226_ (.A(_1865_),
    .B(_1864_),
    .Y(_1867_));
 sg13g2_a21oi_1 _6227_ (.A1(_1861_),
    .A2(_1866_),
    .Y(_1868_),
    .B1(_1867_));
 sg13g2_nor2_1 _6228_ (.A(_1803_),
    .B(_1802_),
    .Y(_1869_));
 sg13g2_a21oi_1 _6229_ (.A1(_1801_),
    .A2(_1804_),
    .Y(_1870_),
    .B1(_1869_));
 sg13g2_o21ai_1 _6230_ (.B1(_1870_),
    .Y(_1871_),
    .A1(_1806_),
    .A2(_1868_));
 sg13g2_buf_2 _6231_ (.A(\i_capsule.tf_x[8] ),
    .X(_1872_));
 sg13g2_inv_1 _6232_ (.Y(_1873_),
    .A(_1872_));
 sg13g2_a21oi_1 _6233_ (.A1(_0954_),
    .A2(net180),
    .Y(_1874_),
    .B1(_1873_));
 sg13g2_inv_1 _6234_ (.Y(_1875_),
    .A(_0954_));
 sg13g2_a21oi_1 _6235_ (.A1(_1875_),
    .A2(_1770_),
    .Y(_1876_),
    .B1(_1872_));
 sg13g2_buf_2 _6236_ (.A(\i_capsule.tf_y[7] ),
    .X(_1877_));
 sg13g2_inv_1 _6237_ (.Y(_1878_),
    .A(_1877_));
 sg13g2_buf_2 _6238_ (.A(\i_capsule.tf_y[8] ),
    .X(_1879_));
 sg13g2_inv_1 _6239_ (.Y(_1880_),
    .A(_1879_));
 sg13g2_a22oi_1 _6240_ (.Y(_1881_),
    .B1(_1878_),
    .B2(_1880_),
    .A2(net179),
    .A1(_1375_));
 sg13g2_inv_1 _6241_ (.Y(_1882_),
    .A(_1375_));
 sg13g2_inv_1 _6242_ (.Y(_1883_),
    .A(net179));
 sg13g2_a22oi_1 _6243_ (.Y(_1884_),
    .B1(_1882_),
    .B2(_1883_),
    .A2(_1879_),
    .A1(_1877_));
 sg13g2_nor4_1 _6244_ (.A(_1874_),
    .B(_1876_),
    .C(_1881_),
    .D(_1884_),
    .Y(_1885_));
 sg13g2_nand2_2 _6245_ (.Y(_1886_),
    .A(_1871_),
    .B(_1885_));
 sg13g2_inv_2 _6246_ (.Y(_1887_),
    .A(_1886_));
 sg13g2_buf_1 _6247_ (.A(\capsule_color[0] ),
    .X(_1888_));
 sg13g2_nor2b_1 _6248_ (.A(net6),
    .B_N(bitmap_pixel),
    .Y(_1889_));
 sg13g2_inv_1 _6249_ (.Y(_1890_),
    .A(_1889_));
 sg13g2_inv_1 _6250_ (.Y(_1891_),
    .A(\capsule_color[1] ));
 sg13g2_inv_1 _6251_ (.Y(_1892_),
    .A(_1888_));
 sg13g2_buf_2 _6252_ (.A(\capsule_color[2] ),
    .X(_1893_));
 sg13g2_nand2_1 _6253_ (.Y(_1894_),
    .A(\capsule_color[3] ),
    .B(_1893_));
 sg13g2_nor2_1 _6254_ (.A(_1892_),
    .B(_1894_),
    .Y(_1895_));
 sg13g2_nor3_1 _6255_ (.A(_1891_),
    .B(net167),
    .C(_1895_),
    .Y(_1896_));
 sg13g2_a21oi_1 _6256_ (.A1(_1888_),
    .A2(net167),
    .Y(_1897_),
    .B1(_1896_));
 sg13g2_a21oi_1 _6257_ (.A1(_3514_),
    .A2(_3608_),
    .Y(_1898_),
    .B1(net5));
 sg13g2_o21ai_1 _6258_ (.B1(_1898_),
    .Y(_1899_),
    .A1(_3514_),
    .A2(_3608_));
 sg13g2_a21o_1 _6259_ (.A2(_1899_),
    .A1(_1886_),
    .B1(net103),
    .X(_1900_));
 sg13g2_a21oi_1 _6260_ (.A1(_1887_),
    .A2(_1897_),
    .Y(_0070_),
    .B1(_1900_));
 sg13g2_o21ai_1 _6261_ (.B1(\capsule_color[1] ),
    .Y(_1901_),
    .A1(_1888_),
    .A2(net167));
 sg13g2_nand2_1 _6262_ (.Y(_1902_),
    .A(_1889_),
    .B(_1894_));
 sg13g2_nand2_1 _6263_ (.Y(_1903_),
    .A(_1887_),
    .B(_3596_));
 sg13g2_a21oi_1 _6264_ (.A1(_1901_),
    .A2(_1902_),
    .Y(_0071_),
    .B1(_1903_));
 sg13g2_inv_1 _6265_ (.Y(_1904_),
    .A(\capsule_color[3] ));
 sg13g2_nor3_1 _6266_ (.A(_1904_),
    .B(_1893_),
    .C(net167),
    .Y(_1905_));
 sg13g2_a21oi_1 _6267_ (.A1(_1893_),
    .A2(net167),
    .Y(_1906_),
    .B1(_1905_));
 sg13g2_a21oi_1 _6268_ (.A1(_3525_),
    .A2(_3540_),
    .Y(_1907_),
    .B1(net5));
 sg13g2_o21ai_1 _6269_ (.B1(_1907_),
    .Y(_1908_),
    .A1(_3525_),
    .A2(_3540_));
 sg13g2_a21o_1 _6270_ (.A2(_1908_),
    .A1(_1886_),
    .B1(net103),
    .X(_1909_));
 sg13g2_a21oi_1 _6271_ (.A1(_1887_),
    .A2(_1906_),
    .Y(_0072_),
    .B1(_1909_));
 sg13g2_a21oi_1 _6272_ (.A1(_1904_),
    .A2(net167),
    .Y(_0073_),
    .B1(_1903_));
 sg13g2_buf_1 _6273_ (.A(\capsule_color[4] ),
    .X(_1910_));
 sg13g2_inv_1 _6274_ (.Y(_1911_),
    .A(\capsule_color[5] ));
 sg13g2_inv_1 _6275_ (.Y(_1912_),
    .A(_1910_));
 sg13g2_nor2_1 _6276_ (.A(_1912_),
    .B(_1894_),
    .Y(_1913_));
 sg13g2_nor3_1 _6277_ (.A(_1911_),
    .B(net167),
    .C(_1913_),
    .Y(_1914_));
 sg13g2_a21oi_1 _6278_ (.A1(_1910_),
    .A2(_1890_),
    .Y(_1915_),
    .B1(_1914_));
 sg13g2_a21oi_1 _6279_ (.A1(_3501_),
    .A2(_3538_),
    .Y(_1916_),
    .B1(net5));
 sg13g2_o21ai_1 _6280_ (.B1(_1916_),
    .Y(_1917_),
    .A1(_3501_),
    .A2(_3538_));
 sg13g2_a21o_1 _6281_ (.A2(_1917_),
    .A1(_1886_),
    .B1(net103),
    .X(_1918_));
 sg13g2_a21oi_1 _6282_ (.A1(_1887_),
    .A2(_1915_),
    .Y(_0074_),
    .B1(_1918_));
 sg13g2_o21ai_1 _6283_ (.B1(\capsule_color[5] ),
    .Y(_1919_),
    .A1(_1910_),
    .A2(net167));
 sg13g2_a21oi_1 _6284_ (.A1(_1902_),
    .A2(_1919_),
    .Y(_0075_),
    .B1(_1903_));
 sg13g2_buf_1 _6285_ (.A(\i_collision.vx[2] ),
    .X(_1920_));
 sg13g2_inv_1 _6286_ (.Y(_1921_),
    .A(net178));
 sg13g2_buf_1 _6287_ (.A(\i_collision.vx[0] ),
    .X(_1922_));
 sg13g2_buf_1 _6288_ (.A(\i_collision.vx[1] ),
    .X(_1923_));
 sg13g2_inv_1 _6289_ (.Y(_1924_),
    .A(_1923_));
 sg13g2_o21ai_1 _6290_ (.B1(net178),
    .Y(_1925_),
    .A1(_1922_),
    .A2(_1924_));
 sg13g2_inv_1 _6291_ (.Y(_1926_),
    .A(_1925_));
 sg13g2_a21oi_1 _6292_ (.A1(_1921_),
    .A2(_0009_),
    .Y(_1927_),
    .B1(_1926_));
 sg13g2_nor2_1 _6293_ (.A(\center_x[0] ),
    .B(_1927_),
    .Y(_1928_));
 sg13g2_nor2b_1 _6294_ (.A(_1598_),
    .B_N(_1927_),
    .Y(_1929_));
 sg13g2_nor2_1 _6295_ (.A(_1928_),
    .B(_1929_),
    .Y(_1930_));
 sg13g2_nor2_1 _6296_ (.A(net178),
    .B(_1924_),
    .Y(_1931_));
 sg13g2_nand2_1 _6297_ (.Y(_1932_),
    .A(_1931_),
    .B(_1922_));
 sg13g2_o21ai_1 _6298_ (.B1(_1932_),
    .Y(_1933_),
    .A1(_1923_),
    .A2(_1922_));
 sg13g2_xnor2_1 _6299_ (.Y(_1934_),
    .A(\i_kinematics.center_x_lo[1] ),
    .B(_1933_));
 sg13g2_inv_1 _6300_ (.Y(_1935_),
    .A(\i_kinematics.center_x_lo[0] ));
 sg13g2_nand2_1 _6301_ (.Y(_1936_),
    .A(_1923_),
    .B(_1922_));
 sg13g2_nor2_1 _6302_ (.A(_1935_),
    .B(_1936_),
    .Y(_1937_));
 sg13g2_nor2b_1 _6303_ (.A(_1933_),
    .B_N(\i_kinematics.center_x_lo[1] ),
    .Y(_1938_));
 sg13g2_a21oi_1 _6304_ (.A1(_1934_),
    .A2(_1937_),
    .Y(_1939_),
    .B1(_1938_));
 sg13g2_xor2_1 _6305_ (.B(_1939_),
    .A(_1930_),
    .X(_1940_));
 sg13g2_buf_1 _6306_ (.A(\i_kinematics.update ),
    .X(_1941_));
 sg13g2_buf_1 _6307_ (.A(net177),
    .X(_1942_));
 sg13g2_buf_1 _6308_ (.A(net177),
    .X(_1943_));
 sg13g2_nor2_2 _6309_ (.A(net2),
    .B(_3492_),
    .Y(_1944_));
 sg13g2_buf_1 _6310_ (.A(_1944_),
    .X(_1945_));
 sg13g2_o21ai_1 _6311_ (.B1(net146),
    .Y(_1946_),
    .A1(\center_x[0] ),
    .A2(net165));
 sg13g2_a21oi_1 _6312_ (.A1(_1940_),
    .A2(net166),
    .Y(_0106_),
    .B1(_1946_));
 sg13g2_inv_1 _6313_ (.Y(_1947_),
    .A(\center_x[1] ));
 sg13g2_inv_1 _6314_ (.Y(_1948_),
    .A(_1922_));
 sg13g2_nor2_1 _6315_ (.A(_1923_),
    .B(_1921_),
    .Y(_1949_));
 sg13g2_nor2_1 _6316_ (.A(_1931_),
    .B(_1949_),
    .Y(_1950_));
 sg13g2_a21oi_1 _6317_ (.A1(_1924_),
    .A2(_1948_),
    .Y(_1951_),
    .B1(_1950_));
 sg13g2_nor2_1 _6318_ (.A(_1947_),
    .B(_1951_),
    .Y(_1952_));
 sg13g2_inv_1 _6319_ (.Y(_1953_),
    .A(_1952_));
 sg13g2_nand2_1 _6320_ (.Y(_1954_),
    .A(_1951_),
    .B(_1947_));
 sg13g2_nand2_1 _6321_ (.Y(_1955_),
    .A(_1953_),
    .B(_1954_));
 sg13g2_inv_1 _6322_ (.Y(_1956_),
    .A(_1929_));
 sg13g2_a21oi_1 _6323_ (.A1(_1939_),
    .A2(_1956_),
    .Y(_1957_),
    .B1(_1928_));
 sg13g2_xor2_1 _6324_ (.B(_1957_),
    .A(_1955_),
    .X(_1958_));
 sg13g2_o21ai_1 _6325_ (.B1(net146),
    .Y(_1959_),
    .A1(\center_x[1] ),
    .A2(net165));
 sg13g2_a21oi_1 _6326_ (.A1(_1958_),
    .A2(net166),
    .Y(_0107_),
    .B1(_1959_));
 sg13g2_nor3_1 _6327_ (.A(\center_x[2] ),
    .B(_1931_),
    .C(_1949_),
    .Y(_1960_));
 sg13g2_nor2_1 _6328_ (.A(_1608_),
    .B(_1950_),
    .Y(_1961_));
 sg13g2_nor2_1 _6329_ (.A(_1960_),
    .B(_1961_),
    .Y(_1962_));
 sg13g2_a21oi_1 _6330_ (.A1(_1957_),
    .A2(_1954_),
    .Y(_1963_),
    .B1(_1952_));
 sg13g2_xor2_1 _6331_ (.B(_1963_),
    .A(_1962_),
    .X(_1964_));
 sg13g2_o21ai_1 _6332_ (.B1(net146),
    .Y(_1965_),
    .A1(\center_x[2] ),
    .A2(net165));
 sg13g2_a21oi_1 _6333_ (.A1(_1964_),
    .A2(net166),
    .Y(_0108_),
    .B1(_1965_));
 sg13g2_xor2_1 _6334_ (.B(_1620_),
    .A(net178),
    .X(_1966_));
 sg13g2_inv_1 _6335_ (.Y(_1967_),
    .A(_1961_));
 sg13g2_o21ai_1 _6336_ (.B1(_1967_),
    .Y(_1968_),
    .A1(_1960_),
    .A2(_1963_));
 sg13g2_xnor2_1 _6337_ (.Y(_1969_),
    .A(_1966_),
    .B(_1968_));
 sg13g2_buf_1 _6338_ (.A(_1941_),
    .X(_1970_));
 sg13g2_buf_1 _6339_ (.A(_1944_),
    .X(_1971_));
 sg13g2_o21ai_1 _6340_ (.B1(net145),
    .Y(_1972_),
    .A1(_1620_),
    .A2(net164));
 sg13g2_a21oi_1 _6341_ (.A1(_1969_),
    .A2(net166),
    .Y(_0109_),
    .B1(_1972_));
 sg13g2_xor2_1 _6342_ (.B(_1626_),
    .A(net178),
    .X(_1973_));
 sg13g2_inv_1 _6343_ (.Y(_1974_),
    .A(_1620_));
 sg13g2_buf_1 _6344_ (.A(net178),
    .X(_1975_));
 sg13g2_a21oi_1 _6345_ (.A1(net163),
    .A2(_1620_),
    .Y(_1976_),
    .B1(_1961_));
 sg13g2_nand2b_1 _6346_ (.Y(_1977_),
    .B(_1962_),
    .A_N(_1963_));
 sg13g2_a22oi_1 _6347_ (.Y(_1978_),
    .B1(_1976_),
    .B2(_1977_),
    .A2(_1974_),
    .A1(_1921_));
 sg13g2_xnor2_1 _6348_ (.Y(_1979_),
    .A(_1973_),
    .B(_1978_));
 sg13g2_o21ai_1 _6349_ (.B1(net145),
    .Y(_1980_),
    .A1(_1626_),
    .A2(net164));
 sg13g2_a21oi_1 _6350_ (.A1(_1979_),
    .A2(net166),
    .Y(_0110_),
    .B1(_1980_));
 sg13g2_xor2_1 _6351_ (.B(_1635_),
    .A(net178),
    .X(_1981_));
 sg13g2_nand3_1 _6352_ (.B(_1966_),
    .C(_1973_),
    .A(_1968_),
    .Y(_1982_));
 sg13g2_o21ai_1 _6353_ (.B1(_1982_),
    .Y(_1983_),
    .A1(_1921_),
    .A2(_1974_));
 sg13g2_a21o_1 _6354_ (.A2(_1626_),
    .A1(_1975_),
    .B1(_1983_),
    .X(_1984_));
 sg13g2_xnor2_1 _6355_ (.Y(_1985_),
    .A(_1981_),
    .B(_1984_));
 sg13g2_o21ai_1 _6356_ (.B1(_1971_),
    .Y(_1986_),
    .A1(_1635_),
    .A2(_1970_));
 sg13g2_a21oi_1 _6357_ (.A1(_1985_),
    .A2(_1942_),
    .Y(_0111_),
    .B1(_1986_));
 sg13g2_inv_1 _6358_ (.Y(_1987_),
    .A(_1981_));
 sg13g2_nand2_1 _6359_ (.Y(_1988_),
    .A(_1978_),
    .B(_1973_));
 sg13g2_nor2_1 _6360_ (.A(_1987_),
    .B(_1988_),
    .Y(_1989_));
 sg13g2_inv_1 _6361_ (.Y(_1990_),
    .A(_1989_));
 sg13g2_o21ai_1 _6362_ (.B1(net163),
    .Y(_1991_),
    .A1(_1635_),
    .A2(_1626_));
 sg13g2_xor2_1 _6363_ (.B(_1644_),
    .A(_1920_),
    .X(_1992_));
 sg13g2_inv_1 _6364_ (.Y(_1993_),
    .A(_1992_));
 sg13g2_a21oi_1 _6365_ (.A1(_1990_),
    .A2(_1991_),
    .Y(_1994_),
    .B1(_1993_));
 sg13g2_nand3_1 _6366_ (.B(_1991_),
    .C(_1993_),
    .A(_1990_),
    .Y(_1995_));
 sg13g2_nand3b_1 _6367_ (.B(_1943_),
    .C(_1995_),
    .Y(_1996_),
    .A_N(_1994_));
 sg13g2_inv_1 _6368_ (.Y(_1997_),
    .A(net177));
 sg13g2_buf_1 _6369_ (.A(_1997_),
    .X(_1998_));
 sg13g2_nand2_1 _6370_ (.Y(_1999_),
    .A(_1998_),
    .B(_1644_));
 sg13g2_nand3_1 _6371_ (.B(_1945_),
    .C(_1999_),
    .A(_1996_),
    .Y(_0112_));
 sg13g2_xor2_1 _6372_ (.B(_1648_),
    .A(net163),
    .X(_2000_));
 sg13g2_inv_1 _6373_ (.Y(_2001_),
    .A(_2000_));
 sg13g2_nand3_1 _6374_ (.B(_1981_),
    .C(_1992_),
    .A(_1984_),
    .Y(_2002_));
 sg13g2_o21ai_1 _6375_ (.B1(net163),
    .Y(_2003_),
    .A1(_1635_),
    .A2(_1644_));
 sg13g2_and2_1 _6376_ (.A(_2002_),
    .B(_2003_),
    .X(_2004_));
 sg13g2_buf_1 _6377_ (.A(_2004_),
    .X(_2005_));
 sg13g2_xnor2_1 _6378_ (.Y(_2006_),
    .A(_2001_),
    .B(_2005_));
 sg13g2_o21ai_1 _6379_ (.B1(_1971_),
    .Y(_2007_),
    .A1(_1648_),
    .A2(_1970_));
 sg13g2_a21oi_1 _6380_ (.A1(_2006_),
    .A2(_1942_),
    .Y(_0113_),
    .B1(_2007_));
 sg13g2_nor2_1 _6381_ (.A(_1993_),
    .B(_2001_),
    .Y(_2008_));
 sg13g2_inv_1 _6382_ (.Y(_2009_),
    .A(_2008_));
 sg13g2_o21ai_1 _6383_ (.B1(net163),
    .Y(_2010_),
    .A1(_1644_),
    .A2(_1648_));
 sg13g2_o21ai_1 _6384_ (.B1(_2010_),
    .Y(_2011_),
    .A1(_1991_),
    .A2(_2009_));
 sg13g2_a21oi_1 _6385_ (.A1(_1989_),
    .A2(_2008_),
    .Y(_2012_),
    .B1(_2011_));
 sg13g2_xor2_1 _6386_ (.B(_1653_),
    .A(net163),
    .X(_2013_));
 sg13g2_nand2b_1 _6387_ (.Y(_2014_),
    .B(_2013_),
    .A_N(_2012_));
 sg13g2_nand2b_1 _6388_ (.Y(_2015_),
    .B(_2012_),
    .A_N(_2013_));
 sg13g2_nand3_1 _6389_ (.B(_2015_),
    .C(_1943_),
    .A(_2014_),
    .Y(_2016_));
 sg13g2_nand2_1 _6390_ (.Y(_2017_),
    .A(_1998_),
    .B(_1653_));
 sg13g2_nand3_1 _6391_ (.B(_1945_),
    .C(_2017_),
    .A(_2016_),
    .Y(_0114_));
 sg13g2_nand2b_1 _6392_ (.Y(_2018_),
    .B(_1648_),
    .A_N(_2005_));
 sg13g2_a21o_1 _6393_ (.A2(_1648_),
    .A1(net163),
    .B1(_1997_),
    .X(_2019_));
 sg13g2_a21oi_1 _6394_ (.A1(net163),
    .A2(_1653_),
    .Y(_2020_),
    .B1(_2019_));
 sg13g2_o21ai_1 _6395_ (.B1(_2020_),
    .Y(_2021_),
    .A1(_1653_),
    .A2(_2005_));
 sg13g2_a21oi_1 _6396_ (.A1(_1921_),
    .A2(_2018_),
    .Y(_2022_),
    .B1(_2021_));
 sg13g2_nor2_1 _6397_ (.A(\center_x[9] ),
    .B(_2022_),
    .Y(_2023_));
 sg13g2_inv_1 _6398_ (.Y(_2024_),
    .A(_1944_));
 sg13g2_a21oi_1 _6399_ (.A1(_2022_),
    .A2(\center_x[9] ),
    .Y(_2025_),
    .B1(_2024_));
 sg13g2_nor2b_1 _6400_ (.A(_2023_),
    .B_N(_2025_),
    .Y(_0115_));
 sg13g2_nor3_1 _6401_ (.A(_1935_),
    .B(net144),
    .C(_1936_),
    .Y(_2026_));
 sg13g2_inv_1 _6402_ (.Y(_2027_),
    .A(_1936_));
 sg13g2_buf_1 _6403_ (.A(net177),
    .X(_2028_));
 sg13g2_a21oi_1 _6404_ (.A1(_2027_),
    .A2(net162),
    .Y(_2029_),
    .B1(\i_kinematics.center_x_lo[0] ));
 sg13g2_nor3_1 _6405_ (.A(_2024_),
    .B(_2026_),
    .C(_2029_),
    .Y(_0116_));
 sg13g2_xnor2_1 _6406_ (.Y(_2030_),
    .A(_1937_),
    .B(_1934_));
 sg13g2_o21ai_1 _6407_ (.B1(net145),
    .Y(_2031_),
    .A1(\i_kinematics.center_x_lo[1] ),
    .A2(net164));
 sg13g2_a21oi_1 _6408_ (.A1(_2030_),
    .A2(net166),
    .Y(_0117_),
    .B1(_2031_));
 sg13g2_buf_1 _6409_ (.A(\i_collision.vy[2] ),
    .X(_2032_));
 sg13g2_inv_1 _6410_ (.Y(_2033_),
    .A(_0008_));
 sg13g2_buf_1 _6411_ (.A(\i_collision.vy[0] ),
    .X(_2034_));
 sg13g2_buf_1 _6412_ (.A(\i_collision.vy[1] ),
    .X(_2035_));
 sg13g2_inv_1 _6413_ (.Y(_2036_),
    .A(_2035_));
 sg13g2_o21ai_1 _6414_ (.B1(net176),
    .Y(_2037_),
    .A1(_2034_),
    .A2(_2036_));
 sg13g2_o21ai_1 _6415_ (.B1(_2037_),
    .Y(_2038_),
    .A1(net176),
    .A2(_2033_));
 sg13g2_nor2_1 _6416_ (.A(_1659_),
    .B(_2038_),
    .Y(_2039_));
 sg13g2_inv_1 _6417_ (.Y(_2040_),
    .A(_2039_));
 sg13g2_nand2_1 _6418_ (.Y(_2041_),
    .A(_2038_),
    .B(_1659_));
 sg13g2_nand2_1 _6419_ (.Y(_2042_),
    .A(_2040_),
    .B(_2041_));
 sg13g2_nor2_1 _6420_ (.A(net176),
    .B(_2036_),
    .Y(_2043_));
 sg13g2_nand2_1 _6421_ (.Y(_2044_),
    .A(_2043_),
    .B(_2034_));
 sg13g2_o21ai_1 _6422_ (.B1(_2044_),
    .Y(_2045_),
    .A1(_2035_),
    .A2(_2034_));
 sg13g2_xnor2_1 _6423_ (.Y(_2046_),
    .A(\i_kinematics.center_y_lo[1] ),
    .B(_2045_));
 sg13g2_inv_1 _6424_ (.Y(_2047_),
    .A(\i_kinematics.center_y_lo[0] ));
 sg13g2_nand2_1 _6425_ (.Y(_2048_),
    .A(_2035_),
    .B(_2034_));
 sg13g2_nor2_1 _6426_ (.A(_2047_),
    .B(_2048_),
    .Y(_2049_));
 sg13g2_nor2b_1 _6427_ (.A(_2045_),
    .B_N(\i_kinematics.center_y_lo[1] ),
    .Y(_2050_));
 sg13g2_a21oi_1 _6428_ (.A1(_2046_),
    .A2(_2049_),
    .Y(_2051_),
    .B1(_2050_));
 sg13g2_xnor2_1 _6429_ (.Y(_2052_),
    .A(_2042_),
    .B(_2051_));
 sg13g2_o21ai_1 _6430_ (.B1(net145),
    .Y(_2053_),
    .A1(\center_y[0] ),
    .A2(net164));
 sg13g2_a21oi_1 _6431_ (.A1(_2052_),
    .A2(net166),
    .Y(_0118_),
    .B1(_2053_));
 sg13g2_inv_1 _6432_ (.Y(_2054_),
    .A(_2034_));
 sg13g2_inv_1 _6433_ (.Y(_2055_),
    .A(net176));
 sg13g2_nor2_1 _6434_ (.A(_2035_),
    .B(_2055_),
    .Y(_2056_));
 sg13g2_nor2_1 _6435_ (.A(_2043_),
    .B(_2056_),
    .Y(_2057_));
 sg13g2_a21o_1 _6436_ (.A2(_2054_),
    .A1(_2036_),
    .B1(_2057_),
    .X(_2058_));
 sg13g2_inv_1 _6437_ (.Y(_2059_),
    .A(_2058_));
 sg13g2_nor2_1 _6438_ (.A(_1666_),
    .B(_2059_),
    .Y(_2060_));
 sg13g2_nand2_1 _6439_ (.Y(_2061_),
    .A(_2059_),
    .B(_1666_));
 sg13g2_nand2b_1 _6440_ (.Y(_2062_),
    .B(_2061_),
    .A_N(_2060_));
 sg13g2_inv_1 _6441_ (.Y(_2063_),
    .A(_2041_));
 sg13g2_a21oi_1 _6442_ (.A1(_2051_),
    .A2(_2040_),
    .Y(_2064_),
    .B1(_2063_));
 sg13g2_xor2_1 _6443_ (.B(_2064_),
    .A(_2062_),
    .X(_2065_));
 sg13g2_o21ai_1 _6444_ (.B1(net145),
    .Y(_2066_),
    .A1(\center_y[1] ),
    .A2(net164));
 sg13g2_a21oi_1 _6445_ (.A1(_2065_),
    .A2(net166),
    .Y(_0119_),
    .B1(_2066_));
 sg13g2_nor2_1 _6446_ (.A(_1670_),
    .B(_2057_),
    .Y(_2067_));
 sg13g2_inv_1 _6447_ (.Y(_2068_),
    .A(_2067_));
 sg13g2_nand2_1 _6448_ (.Y(_2069_),
    .A(_2057_),
    .B(_1670_));
 sg13g2_nand2_1 _6449_ (.Y(_2070_),
    .A(_2068_),
    .B(_2069_));
 sg13g2_inv_1 _6450_ (.Y(_2071_),
    .A(_2070_));
 sg13g2_a21o_1 _6451_ (.A2(_2061_),
    .A1(_2064_),
    .B1(_2060_),
    .X(_2072_));
 sg13g2_xnor2_1 _6452_ (.Y(_2073_),
    .A(_2071_),
    .B(_2072_));
 sg13g2_buf_1 _6453_ (.A(net177),
    .X(_2074_));
 sg13g2_o21ai_1 _6454_ (.B1(net145),
    .Y(_2075_),
    .A1(\center_y[2] ),
    .A2(net164));
 sg13g2_a21oi_1 _6455_ (.A1(_2073_),
    .A2(net161),
    .Y(_0120_),
    .B1(_2075_));
 sg13g2_nor2_1 _6456_ (.A(net176),
    .B(\center_y[3] ),
    .Y(_2076_));
 sg13g2_nand2_1 _6457_ (.Y(_2077_),
    .A(net176),
    .B(\center_y[3] ));
 sg13g2_inv_1 _6458_ (.Y(_2078_),
    .A(_2077_));
 sg13g2_nor2_1 _6459_ (.A(_2076_),
    .B(_2078_),
    .Y(_2079_));
 sg13g2_nand2b_1 _6460_ (.Y(_2080_),
    .B(_2064_),
    .A_N(_2062_));
 sg13g2_a21oi_1 _6461_ (.A1(_2060_),
    .A2(_2069_),
    .Y(_2081_),
    .B1(_2067_));
 sg13g2_o21ai_1 _6462_ (.B1(_2081_),
    .Y(_2082_),
    .A1(_2070_),
    .A2(_2080_));
 sg13g2_xnor2_1 _6463_ (.Y(_2083_),
    .A(_2079_),
    .B(_2082_));
 sg13g2_o21ai_1 _6464_ (.B1(net145),
    .Y(_2084_),
    .A1(\center_y[3] ),
    .A2(net164));
 sg13g2_a21oi_1 _6465_ (.A1(_2083_),
    .A2(net161),
    .Y(_0121_),
    .B1(_2084_));
 sg13g2_nor2_1 _6466_ (.A(net176),
    .B(_1686_),
    .Y(_2085_));
 sg13g2_inv_1 _6467_ (.Y(_2086_),
    .A(_2085_));
 sg13g2_nand2_1 _6468_ (.Y(_2087_),
    .A(net176),
    .B(_1686_));
 sg13g2_nand2_1 _6469_ (.Y(_2088_),
    .A(_2086_),
    .B(_2087_));
 sg13g2_nand2_1 _6470_ (.Y(_2089_),
    .A(_2072_),
    .B(_2071_));
 sg13g2_nor2_1 _6471_ (.A(_2078_),
    .B(_2067_),
    .Y(_2090_));
 sg13g2_a21oi_1 _6472_ (.A1(_2089_),
    .A2(_2090_),
    .Y(_2091_),
    .B1(_2076_));
 sg13g2_nor2b_1 _6473_ (.A(_2088_),
    .B_N(_2091_),
    .Y(_2092_));
 sg13g2_inv_1 _6474_ (.Y(_2093_),
    .A(_2092_));
 sg13g2_nand2b_1 _6475_ (.Y(_2094_),
    .B(_2088_),
    .A_N(_2091_));
 sg13g2_nand3_1 _6476_ (.B(net165),
    .C(_2094_),
    .A(_2093_),
    .Y(_2095_));
 sg13g2_nand2_1 _6477_ (.Y(_2096_),
    .A(net144),
    .B(_1686_));
 sg13g2_nand3_1 _6478_ (.B(net146),
    .C(_2096_),
    .A(_2095_),
    .Y(_0122_));
 sg13g2_buf_1 _6479_ (.A(_2032_),
    .X(_2097_));
 sg13g2_xor2_1 _6480_ (.B(_1694_),
    .A(_2097_),
    .X(_2098_));
 sg13g2_inv_1 _6481_ (.Y(_2099_),
    .A(_2098_));
 sg13g2_nand2_1 _6482_ (.Y(_2100_),
    .A(_2082_),
    .B(_2079_));
 sg13g2_o21ai_1 _6483_ (.B1(_2077_),
    .Y(_2101_),
    .A1(_2088_),
    .A2(_2100_));
 sg13g2_nor2b_1 _6484_ (.A(_2101_),
    .B_N(_2087_),
    .Y(_2102_));
 sg13g2_nor2_1 _6485_ (.A(_2099_),
    .B(_2102_),
    .Y(_2103_));
 sg13g2_inv_1 _6486_ (.Y(_2104_),
    .A(_2103_));
 sg13g2_a21oi_1 _6487_ (.A1(_2102_),
    .A2(_2099_),
    .Y(_2105_),
    .B1(_1997_));
 sg13g2_a22oi_1 _6488_ (.Y(_2106_),
    .B1(_2104_),
    .B2(_2105_),
    .A2(net144),
    .A1(_1694_));
 sg13g2_nand2_1 _6489_ (.Y(_0123_),
    .A(_2106_),
    .B(net146));
 sg13g2_nor2_1 _6490_ (.A(_2099_),
    .B(_2093_),
    .Y(_2107_));
 sg13g2_inv_1 _6491_ (.Y(_2108_),
    .A(_2107_));
 sg13g2_o21ai_1 _6492_ (.B1(net160),
    .Y(_2109_),
    .A1(_1686_),
    .A2(_1694_));
 sg13g2_xor2_1 _6493_ (.B(_1700_),
    .A(net160),
    .X(_2110_));
 sg13g2_inv_1 _6494_ (.Y(_2111_),
    .A(_2110_));
 sg13g2_a21oi_1 _6495_ (.A1(_2108_),
    .A2(_2109_),
    .Y(_2112_),
    .B1(_2111_));
 sg13g2_nand3_1 _6496_ (.B(_2109_),
    .C(_2111_),
    .A(_2108_),
    .Y(_2113_));
 sg13g2_nand3b_1 _6497_ (.B(net165),
    .C(_2113_),
    .Y(_2114_),
    .A_N(_2112_));
 sg13g2_nand2_1 _6498_ (.Y(_2115_),
    .A(net144),
    .B(_1700_));
 sg13g2_nand3_1 _6499_ (.B(net146),
    .C(_2115_),
    .A(_2114_),
    .Y(_0124_));
 sg13g2_nor2_1 _6500_ (.A(_2111_),
    .B(_2104_),
    .Y(_2116_));
 sg13g2_o21ai_1 _6501_ (.B1(net160),
    .Y(_2117_),
    .A1(_1694_),
    .A2(_1700_));
 sg13g2_nor2b_1 _6502_ (.A(_2116_),
    .B_N(_2117_),
    .Y(_2118_));
 sg13g2_xor2_1 _6503_ (.B(_1706_),
    .A(net160),
    .X(_2119_));
 sg13g2_nand2b_1 _6504_ (.Y(_2120_),
    .B(_2119_),
    .A_N(_2118_));
 sg13g2_nand2b_1 _6505_ (.Y(_2121_),
    .B(_2118_),
    .A_N(_2119_));
 sg13g2_nand3_1 _6506_ (.B(net165),
    .C(_2121_),
    .A(_2120_),
    .Y(_2122_));
 sg13g2_nand2_1 _6507_ (.Y(_2123_),
    .A(net144),
    .B(_1706_));
 sg13g2_nand3_1 _6508_ (.B(net146),
    .C(_2123_),
    .A(_2122_),
    .Y(_0125_));
 sg13g2_xor2_1 _6509_ (.B(_1710_),
    .A(net160),
    .X(_2124_));
 sg13g2_nand2_1 _6510_ (.Y(_2125_),
    .A(_2110_),
    .B(_2119_));
 sg13g2_nor2_1 _6511_ (.A(_2109_),
    .B(_2125_),
    .Y(_2126_));
 sg13g2_o21ai_1 _6512_ (.B1(net160),
    .Y(_2127_),
    .A1(_1700_),
    .A2(_1706_));
 sg13g2_nor2b_1 _6513_ (.A(_2126_),
    .B_N(_2127_),
    .Y(_2128_));
 sg13g2_o21ai_1 _6514_ (.B1(_2128_),
    .Y(_2129_),
    .A1(_2125_),
    .A2(_2108_));
 sg13g2_xnor2_1 _6515_ (.Y(_2130_),
    .A(_2124_),
    .B(_2129_));
 sg13g2_o21ai_1 _6516_ (.B1(net145),
    .Y(_2131_),
    .A1(_1710_),
    .A2(net164));
 sg13g2_a21oi_1 _6517_ (.A1(_2130_),
    .A2(_2074_),
    .Y(_0126_),
    .B1(_2131_));
 sg13g2_inv_1 _6518_ (.Y(_2132_),
    .A(_1710_));
 sg13g2_a21oi_1 _6519_ (.A1(net160),
    .A2(_1706_),
    .Y(_2133_),
    .B1(_1997_));
 sg13g2_o21ai_1 _6520_ (.B1(_2133_),
    .Y(_2134_),
    .A1(_2055_),
    .A2(_2132_));
 sg13g2_a21oi_1 _6521_ (.A1(_2116_),
    .A2(_1706_),
    .Y(_2135_),
    .B1(net160));
 sg13g2_nor2_1 _6522_ (.A(_1710_),
    .B(_2118_),
    .Y(_2136_));
 sg13g2_nor3_1 _6523_ (.A(_2134_),
    .B(_2135_),
    .C(_2136_),
    .Y(_2137_));
 sg13g2_buf_1 _6524_ (.A(_1944_),
    .X(_2138_));
 sg13g2_o21ai_1 _6525_ (.B1(_2138_),
    .Y(_2139_),
    .A1(\center_y[9] ),
    .A2(_2137_));
 sg13g2_a21oi_1 _6526_ (.A1(\center_y[9] ),
    .A2(_2137_),
    .Y(_0127_),
    .B1(_2139_));
 sg13g2_nor3_1 _6527_ (.A(_2047_),
    .B(net144),
    .C(_2048_),
    .Y(_2140_));
 sg13g2_inv_1 _6528_ (.Y(_2141_),
    .A(_2048_));
 sg13g2_a21oi_1 _6529_ (.A1(_2141_),
    .A2(_2028_),
    .Y(_2142_),
    .B1(\i_kinematics.center_y_lo[0] ));
 sg13g2_nor3_1 _6530_ (.A(_2024_),
    .B(_2140_),
    .C(_2142_),
    .Y(_0128_));
 sg13g2_xnor2_1 _6531_ (.Y(_2143_),
    .A(_2049_),
    .B(_2046_));
 sg13g2_o21ai_1 _6532_ (.B1(net143),
    .Y(_2144_),
    .A1(\i_kinematics.center_y_lo[1] ),
    .A2(_2028_));
 sg13g2_a21oi_1 _6533_ (.A1(_2143_),
    .A2(_2074_),
    .Y(_0129_),
    .B1(_2144_));
 sg13g2_inv_1 _6534_ (.Y(_2145_),
    .A(\i_kinematics.phi[0] ));
 sg13g2_buf_2 _6535_ (.A(\i_collision.i_coll_table.in[3] ),
    .X(_2146_));
 sg13g2_buf_2 _6536_ (.A(\i_collision.i_coll_table.in[4] ),
    .X(_2147_));
 sg13g2_nand2_1 _6537_ (.Y(_2148_),
    .A(_2146_),
    .B(_2147_));
 sg13g2_nor3_1 _6538_ (.A(_2145_),
    .B(net144),
    .C(_2148_),
    .Y(_2149_));
 sg13g2_inv_1 _6539_ (.Y(_2150_),
    .A(_2148_));
 sg13g2_a21oi_1 _6540_ (.A1(_2150_),
    .A2(net177),
    .Y(_2151_),
    .B1(\i_kinematics.phi[0] ));
 sg13g2_nor3_1 _6541_ (.A(_2024_),
    .B(_2149_),
    .C(_2151_),
    .Y(_0130_));
 sg13g2_buf_1 _6542_ (.A(\i_collision.i_coll_table.in[5] ),
    .X(_2152_));
 sg13g2_buf_1 _6543_ (.A(_2152_),
    .X(_2153_));
 sg13g2_buf_1 _6544_ (.A(net159),
    .X(_2154_));
 sg13g2_buf_1 _6545_ (.A(net142),
    .X(_2155_));
 sg13g2_inv_1 _6546_ (.Y(_2156_),
    .A(_3695_));
 sg13g2_inv_2 _6547_ (.Y(_2157_),
    .A(net142));
 sg13g2_nor2_1 _6548_ (.A(_3683_),
    .B(net159),
    .Y(_2158_));
 sg13g2_inv_2 _6549_ (.Y(_2159_),
    .A(_2147_));
 sg13g2_nor2_1 _6550_ (.A(_2146_),
    .B(_2159_),
    .Y(_2160_));
 sg13g2_nor2_1 _6551_ (.A(_2152_),
    .B(_0052_),
    .Y(_2161_));
 sg13g2_a21o_1 _6552_ (.A2(net159),
    .A1(_2160_),
    .B1(_2161_),
    .X(_2162_));
 sg13g2_nor2_1 _6553_ (.A(\i_kinematics.phi[2] ),
    .B(_2162_),
    .Y(_2163_));
 sg13g2_inv_1 _6554_ (.Y(_2164_),
    .A(_2146_));
 sg13g2_nor2_2 _6555_ (.A(_2147_),
    .B(net158),
    .Y(_2165_));
 sg13g2_nand2_1 _6556_ (.Y(_2166_),
    .A(_2147_),
    .B(_2152_));
 sg13g2_inv_1 _6557_ (.Y(_2167_),
    .A(_2166_));
 sg13g2_nor3_1 _6558_ (.A(_2165_),
    .B(_2167_),
    .C(_2160_),
    .Y(_2168_));
 sg13g2_xnor2_1 _6559_ (.Y(_2169_),
    .A(\i_kinematics.phi[1] ),
    .B(_2168_));
 sg13g2_nor2_1 _6560_ (.A(_2145_),
    .B(_2148_),
    .Y(_2170_));
 sg13g2_nor2b_1 _6561_ (.A(_2168_),
    .B_N(\i_kinematics.phi[1] ),
    .Y(_2171_));
 sg13g2_a21oi_1 _6562_ (.A1(_2169_),
    .A2(_2170_),
    .Y(_2172_),
    .B1(_2171_));
 sg13g2_nand2_1 _6563_ (.Y(_2173_),
    .A(_2162_),
    .B(\i_kinematics.phi[2] ));
 sg13g2_o21ai_1 _6564_ (.B1(_2173_),
    .Y(_2174_),
    .A1(_2163_),
    .A2(_2172_));
 sg13g2_nor2_2 _6565_ (.A(_2146_),
    .B(_2147_),
    .Y(_2175_));
 sg13g2_xor2_1 _6566_ (.B(net159),
    .A(_2147_),
    .X(_2176_));
 sg13g2_inv_1 _6567_ (.Y(_2177_),
    .A(_2176_));
 sg13g2_nor2_1 _6568_ (.A(_2175_),
    .B(_2177_),
    .Y(_2178_));
 sg13g2_inv_1 _6569_ (.Y(_2179_),
    .A(_3674_));
 sg13g2_nand2_1 _6570_ (.Y(_2180_),
    .A(_2178_),
    .B(_2179_));
 sg13g2_nor2_1 _6571_ (.A(_2179_),
    .B(_2178_),
    .Y(_2181_));
 sg13g2_a21oi_1 _6572_ (.A1(_2174_),
    .A2(_2180_),
    .Y(_2182_),
    .B1(_2181_));
 sg13g2_inv_1 _6573_ (.Y(_2183_),
    .A(_2182_));
 sg13g2_inv_1 _6574_ (.Y(_2184_),
    .A(_3676_));
 sg13g2_nand2_1 _6575_ (.Y(_2185_),
    .A(_2177_),
    .B(_2184_));
 sg13g2_nor2_1 _6576_ (.A(_2184_),
    .B(_2177_),
    .Y(_2186_));
 sg13g2_a221oi_1 _6577_ (.B2(_2185_),
    .C1(_2186_),
    .B1(_2183_),
    .A1(_3683_),
    .Y(_2187_),
    .A2(net159));
 sg13g2_nor2_1 _6578_ (.A(_2158_),
    .B(_2187_),
    .Y(_2188_));
 sg13g2_nor2_1 _6579_ (.A(\i_kinematics.phi[6] ),
    .B(net159),
    .Y(_2189_));
 sg13g2_inv_1 _6580_ (.Y(_2190_),
    .A(_2189_));
 sg13g2_nand2_1 _6581_ (.Y(_2191_),
    .A(\i_kinematics.phi[6] ),
    .B(net159));
 sg13g2_inv_1 _6582_ (.Y(_2192_),
    .A(_2191_));
 sg13g2_a21oi_2 _6583_ (.B1(_2192_),
    .Y(_2193_),
    .A2(_2190_),
    .A1(_2188_));
 sg13g2_a21oi_1 _6584_ (.A1(_2156_),
    .A2(_2157_),
    .Y(_2194_),
    .B1(_2193_));
 sg13g2_a21oi_1 _6585_ (.A1(_3695_),
    .A2(net131),
    .Y(_2195_),
    .B1(_2194_));
 sg13g2_nand3_1 _6586_ (.B(net131),
    .C(_3701_),
    .A(_2195_),
    .Y(_2196_));
 sg13g2_buf_1 _6587_ (.A(_2157_),
    .X(_2197_));
 sg13g2_nand3_1 _6588_ (.B(net121),
    .C(_3703_),
    .A(_2194_),
    .Y(_2198_));
 sg13g2_a21oi_1 _6589_ (.A1(_2196_),
    .A2(_2198_),
    .Y(_2199_),
    .B1(_1997_));
 sg13g2_o21ai_1 _6590_ (.B1(_2138_),
    .Y(_2200_),
    .A1(_3754_),
    .A2(_2199_));
 sg13g2_a21oi_1 _6591_ (.A1(_3754_),
    .A2(_2199_),
    .Y(_0131_),
    .B1(_2200_));
 sg13g2_xnor2_1 _6592_ (.Y(_2201_),
    .A(_2170_),
    .B(_2169_));
 sg13g2_o21ai_1 _6593_ (.B1(net143),
    .Y(_2202_),
    .A1(\i_kinematics.phi[1] ),
    .A2(net162));
 sg13g2_a21oi_1 _6594_ (.A1(_2201_),
    .A2(net161),
    .Y(_0132_),
    .B1(_2202_));
 sg13g2_nand2b_1 _6595_ (.Y(_2203_),
    .B(_2173_),
    .A_N(_2163_));
 sg13g2_xnor2_1 _6596_ (.Y(_2204_),
    .A(_2203_),
    .B(_2172_));
 sg13g2_o21ai_1 _6597_ (.B1(net143),
    .Y(_2205_),
    .A1(\i_kinematics.phi[2] ),
    .A2(net162));
 sg13g2_a21oi_1 _6598_ (.A1(_2204_),
    .A2(net161),
    .Y(_0133_),
    .B1(_2205_));
 sg13g2_nor2b_1 _6599_ (.A(_2181_),
    .B_N(_2180_),
    .Y(_2206_));
 sg13g2_xnor2_1 _6600_ (.Y(_2207_),
    .A(_2206_),
    .B(_2174_));
 sg13g2_o21ai_1 _6601_ (.B1(net143),
    .Y(_2208_),
    .A1(_3674_),
    .A2(net162));
 sg13g2_a21oi_1 _6602_ (.A1(_2207_),
    .A2(net161),
    .Y(_0134_),
    .B1(_2208_));
 sg13g2_inv_1 _6603_ (.Y(_2209_),
    .A(_2186_));
 sg13g2_nand2_1 _6604_ (.Y(_2210_),
    .A(_2209_),
    .B(_2185_));
 sg13g2_xnor2_1 _6605_ (.Y(_2211_),
    .A(_2210_),
    .B(_2182_));
 sg13g2_o21ai_1 _6606_ (.B1(net143),
    .Y(_2212_),
    .A1(_3676_),
    .A2(net162));
 sg13g2_a21oi_1 _6607_ (.A1(_2211_),
    .A2(net161),
    .Y(_0135_),
    .B1(_2212_));
 sg13g2_nand2_1 _6608_ (.Y(_2213_),
    .A(_3683_),
    .B(net131));
 sg13g2_nor2b_1 _6609_ (.A(_2158_),
    .B_N(_2213_),
    .Y(_2214_));
 sg13g2_nand2_1 _6610_ (.Y(_2215_),
    .A(_2174_),
    .B(_2206_));
 sg13g2_a21oi_1 _6611_ (.A1(_2181_),
    .A2(_2185_),
    .Y(_2216_),
    .B1(_2186_));
 sg13g2_o21ai_1 _6612_ (.B1(_2216_),
    .Y(_2217_),
    .A1(_2210_),
    .A2(_2215_));
 sg13g2_xnor2_1 _6613_ (.Y(_2218_),
    .A(_2214_),
    .B(_2217_));
 sg13g2_o21ai_1 _6614_ (.B1(net143),
    .Y(_2219_),
    .A1(_3683_),
    .A2(net162));
 sg13g2_a21oi_1 _6615_ (.A1(_2218_),
    .A2(net161),
    .Y(_0136_),
    .B1(_2219_));
 sg13g2_nor2_1 _6616_ (.A(_2189_),
    .B(_2192_),
    .Y(_2220_));
 sg13g2_xnor2_1 _6617_ (.Y(_2221_),
    .A(_2220_),
    .B(_2188_));
 sg13g2_o21ai_1 _6618_ (.B1(net143),
    .Y(_2222_),
    .A1(\i_kinematics.phi[6] ),
    .A2(net162));
 sg13g2_a21oi_1 _6619_ (.A1(_2221_),
    .A2(net161),
    .Y(_0137_),
    .B1(_2222_));
 sg13g2_xnor2_1 _6620_ (.Y(_2223_),
    .A(_3695_),
    .B(_2155_));
 sg13g2_xnor2_1 _6621_ (.Y(_2224_),
    .A(_2223_),
    .B(_2193_));
 sg13g2_o21ai_1 _6622_ (.B1(net143),
    .Y(_2225_),
    .A1(_3695_),
    .A2(net162));
 sg13g2_a21oi_1 _6623_ (.A1(_2224_),
    .A2(net165),
    .Y(_0138_),
    .B1(_2225_));
 sg13g2_buf_1 _6624_ (.A(net181),
    .X(_2226_));
 sg13g2_nor2_2 _6625_ (.A(net157),
    .B(net142),
    .Y(_2227_));
 sg13g2_nand2_1 _6626_ (.Y(_2228_),
    .A(net157),
    .B(net159));
 sg13g2_inv_1 _6627_ (.Y(_2229_),
    .A(_2228_));
 sg13g2_nor2_1 _6628_ (.A(_2227_),
    .B(_2229_),
    .Y(_2230_));
 sg13g2_xnor2_1 _6629_ (.Y(_2231_),
    .A(_2230_),
    .B(_2195_));
 sg13g2_nand2_1 _6630_ (.Y(_2232_),
    .A(_2231_),
    .B(net165));
 sg13g2_nand2_1 _6631_ (.Y(_2233_),
    .A(net144),
    .B(net157));
 sg13g2_nand3_1 _6632_ (.B(net146),
    .C(_2233_),
    .A(_2232_),
    .Y(_0139_));
 sg13g2_nand3_1 _6633_ (.B(_2226_),
    .C(_3695_),
    .A(net121),
    .Y(_2234_));
 sg13g2_inv_1 _6634_ (.Y(_2235_),
    .A(_2226_));
 sg13g2_nand4_1 _6635_ (.B(_2235_),
    .C(_2156_),
    .A(_2193_),
    .Y(_2236_),
    .D(_2155_));
 sg13g2_o21ai_1 _6636_ (.B1(_2236_),
    .Y(_2237_),
    .A1(_2193_),
    .A2(_2234_));
 sg13g2_a21oi_1 _6637_ (.A1(_2237_),
    .A2(net177),
    .Y(_2238_),
    .B1(_3700_));
 sg13g2_and3_1 _6638_ (.X(_2239_),
    .A(_2237_),
    .B(_3700_),
    .C(net177));
 sg13g2_nor3_1 _6639_ (.A(_2024_),
    .B(_2238_),
    .C(_2239_),
    .Y(_0140_));
 sg13g2_inv_1 _6640_ (.Y(_2240_),
    .A(_0004_));
 sg13g2_buf_1 _6641_ (.A(\i_orchestrator.hit_left ),
    .X(_2241_));
 sg13g2_nor2_1 _6642_ (.A(\i_orchestrator.hit_bottom ),
    .B(_2241_),
    .Y(_2242_));
 sg13g2_and3_1 _6643_ (.X(_2243_),
    .A(_2242_),
    .B(_0057_),
    .C(_0056_));
 sg13g2_inv_1 _6644_ (.Y(_2244_),
    .A(_2243_));
 sg13g2_inv_1 _6645_ (.Y(_2245_),
    .A(\collision_impact[1] ));
 sg13g2_inv_1 _6646_ (.Y(_2246_),
    .A(\collision_impact[0] ));
 sg13g2_nand2_1 _6647_ (.Y(_2247_),
    .A(_2245_),
    .B(_2246_));
 sg13g2_nand2_1 _6648_ (.Y(_2248_),
    .A(_2244_),
    .B(_2247_));
 sg13g2_nor4_1 _6649_ (.A(net182),
    .B(_3509_),
    .C(_3513_),
    .D(_1718_),
    .Y(_2249_));
 sg13g2_inv_1 _6650_ (.Y(_2250_),
    .A(_2249_));
 sg13g2_inv_1 _6651_ (.Y(_2251_),
    .A(_3528_));
 sg13g2_nor3_1 _6652_ (.A(_3608_),
    .B(_3538_),
    .C(_3540_),
    .Y(_2252_));
 sg13g2_nor2_1 _6653_ (.A(\i_orchestrator.vga_x[0] ),
    .B(\i_orchestrator.vga_x[1] ),
    .Y(_2253_));
 sg13g2_nand3_1 _6654_ (.B(_3605_),
    .C(_2253_),
    .A(_2252_),
    .Y(_2254_));
 sg13g2_nor4_2 _6655_ (.A(\i_orchestrator.vga_x[9] ),
    .B(_3534_),
    .C(_1720_),
    .Y(_2255_),
    .D(_2254_));
 sg13g2_inv_1 _6656_ (.Y(_2256_),
    .A(_2255_));
 sg13g2_nor2_1 _6657_ (.A(_2251_),
    .B(_2256_),
    .Y(_2257_));
 sg13g2_inv_1 _6658_ (.Y(_2258_),
    .A(_2257_));
 sg13g2_nor2_2 _6659_ (.A(_2250_),
    .B(_2258_),
    .Y(_2259_));
 sg13g2_inv_1 _6660_ (.Y(_2260_),
    .A(_2259_));
 sg13g2_nor3_1 _6661_ (.A(_3492_),
    .B(_2248_),
    .C(_2260_),
    .Y(_2261_));
 sg13g2_nor2b_1 _6662_ (.A(_2240_),
    .B_N(_2261_),
    .Y(_0141_));
 sg13g2_nor2_1 _6663_ (.A(net3),
    .B(\i_orchestrator.trigger_debounce ),
    .Y(_2262_));
 sg13g2_nand2_1 _6664_ (.Y(_2263_),
    .A(_2261_),
    .B(_2262_));
 sg13g2_nor2_1 _6665_ (.A(_2246_),
    .B(_2263_),
    .Y(_0174_));
 sg13g2_nor2_1 _6666_ (.A(_2245_),
    .B(_2263_),
    .Y(_0175_));
 sg13g2_buf_1 _6667_ (.A(net168),
    .X(_2264_));
 sg13g2_nor4_1 _6668_ (.A(net141),
    .B(net1),
    .C(_3519_),
    .D(_2258_),
    .Y(_0177_));
 sg13g2_buf_1 _6669_ (.A(net168),
    .X(_2265_));
 sg13g2_nor2_1 _6670_ (.A(_1746_),
    .B(_2258_),
    .Y(_2266_));
 sg13g2_inv_1 _6671_ (.Y(_2267_),
    .A(_2266_));
 sg13g2_nor3_1 _6672_ (.A(net140),
    .B(_3520_),
    .C(_2267_),
    .Y(_0179_));
 sg13g2_buf_1 _6673_ (.A(\i_orchestrator.trigger_resonator[0] ),
    .X(_2268_));
 sg13g2_nor2_1 _6674_ (.A(\i_orchestrator.trigger_resonator[1] ),
    .B(_2268_),
    .Y(_2269_));
 sg13g2_inv_1 _6675_ (.Y(_2270_),
    .A(_2269_));
 sg13g2_nor2_1 _6676_ (.A(net4),
    .B(_3492_),
    .Y(_2271_));
 sg13g2_inv_1 _6677_ (.Y(_2272_),
    .A(_2271_));
 sg13g2_nor2_1 _6678_ (.A(_2270_),
    .B(_2272_),
    .Y(_2273_));
 sg13g2_inv_1 _6679_ (.Y(_2274_),
    .A(_2273_));
 sg13g2_buf_1 _6680_ (.A(_2274_),
    .X(_2275_));
 sg13g2_buf_1 _6681_ (.A(\i_resonator.counter[0] ),
    .X(_2276_));
 sg13g2_nor2_1 _6682_ (.A(\i_resonator.counter[2] ),
    .B(\i_resonator.counter[3] ),
    .Y(_2277_));
 sg13g2_nand2_1 _6683_ (.Y(_2278_),
    .A(_2277_),
    .B(_0062_));
 sg13g2_inv_1 _6684_ (.Y(_2279_),
    .A(_2278_));
 sg13g2_nor2_1 _6685_ (.A(_2276_),
    .B(_2279_),
    .Y(_2280_));
 sg13g2_nand2_1 _6686_ (.Y(_2281_),
    .A(_2279_),
    .B(_0061_));
 sg13g2_buf_2 _6687_ (.A(_2281_),
    .X(_2282_));
 sg13g2_inv_1 _6688_ (.Y(_2283_),
    .A(_2282_));
 sg13g2_nand3b_1 _6689_ (.B(_2277_),
    .C(_2276_),
    .Y(_2284_),
    .A_N(\i_resonator.counter[1] ));
 sg13g2_buf_1 _6690_ (.A(_2284_),
    .X(_2285_));
 sg13g2_nand2_1 _6691_ (.Y(_2286_),
    .A(_2283_),
    .B(_2285_));
 sg13g2_inv_1 _6692_ (.Y(_2287_),
    .A(_2286_));
 sg13g2_a22oi_1 _6693_ (.Y(_2288_),
    .B1(_2276_),
    .B2(_2287_),
    .A2(_2280_),
    .A1(_0061_));
 sg13g2_nor2_1 _6694_ (.A(net109),
    .B(_2288_),
    .Y(_0180_));
 sg13g2_nor2_1 _6695_ (.A(\i_resonator.counter[1] ),
    .B(_2276_),
    .Y(_2289_));
 sg13g2_nand2_1 _6696_ (.Y(_2290_),
    .A(\i_resonator.counter[1] ),
    .B(_2276_));
 sg13g2_inv_1 _6697_ (.Y(_2291_),
    .A(_2290_));
 sg13g2_buf_1 _6698_ (.A(\i_orchestrator.update_resonator ),
    .X(_2292_));
 sg13g2_nor2_1 _6699_ (.A(_2292_),
    .B(_2279_),
    .Y(_2293_));
 sg13g2_o21ai_1 _6700_ (.B1(_2293_),
    .Y(_2294_),
    .A1(_2289_),
    .A2(_2291_));
 sg13g2_buf_1 _6701_ (.A(_2292_),
    .X(_2295_));
 sg13g2_nand2_1 _6702_ (.Y(_2296_),
    .A(_2295_),
    .B(\i_orchestrator.tension[1] ));
 sg13g2_a21o_1 _6703_ (.A2(_2296_),
    .A1(_2294_),
    .B1(_2287_),
    .X(_2297_));
 sg13g2_buf_1 _6704_ (.A(_2283_),
    .X(_2298_));
 sg13g2_buf_1 _6705_ (.A(_2298_),
    .X(_2299_));
 sg13g2_nand2_1 _6706_ (.Y(_2300_),
    .A(_2299_),
    .B(\i_resonator.counter[1] ));
 sg13g2_a21oi_1 _6707_ (.A1(_2297_),
    .A2(_2300_),
    .Y(_0181_),
    .B1(_2275_));
 sg13g2_buf_1 _6708_ (.A(_2295_),
    .X(_2301_));
 sg13g2_inv_1 _6709_ (.Y(_2302_),
    .A(\i_resonator.counter[2] ));
 sg13g2_xnor2_1 _6710_ (.Y(_2303_),
    .A(_2302_),
    .B(_2289_));
 sg13g2_a22oi_1 _6711_ (.Y(_2304_),
    .B1(_2303_),
    .B2(_2293_),
    .A2(\i_orchestrator.tension[2] ),
    .A1(_2301_));
 sg13g2_nor3_1 _6712_ (.A(_2275_),
    .B(_2287_),
    .C(_2304_),
    .Y(_0182_));
 sg13g2_nand2_1 _6713_ (.Y(_2305_),
    .A(_2289_),
    .B(_2302_));
 sg13g2_xnor2_1 _6714_ (.Y(_2306_),
    .A(\i_resonator.counter[3] ),
    .B(_2305_));
 sg13g2_a22oi_1 _6715_ (.Y(_2307_),
    .B1(_2293_),
    .B2(_2306_),
    .A2(\i_orchestrator.tension[3] ),
    .A1(_2301_));
 sg13g2_nor3_1 _6716_ (.A(_2274_),
    .B(_2287_),
    .C(_2307_),
    .Y(_0183_));
 sg13g2_inv_1 _6717_ (.Y(_2308_),
    .A(_0039_));
 sg13g2_buf_1 _6718_ (.A(\i_resonator.v[15] ),
    .X(_2309_));
 sg13g2_buf_2 _6719_ (.A(\i_resonator.v[14] ),
    .X(_2310_));
 sg13g2_xor2_1 _6720_ (.B(_2310_),
    .A(net175),
    .X(_2311_));
 sg13g2_buf_2 _6721_ (.A(\i_resonator.v[13] ),
    .X(_2312_));
 sg13g2_xnor2_1 _6722_ (.Y(_2313_),
    .A(net175),
    .B(_2312_));
 sg13g2_nor2b_1 _6723_ (.A(_2311_),
    .B_N(_2313_),
    .Y(_2314_));
 sg13g2_buf_1 _6724_ (.A(\i_delta_sigma.sample[11] ),
    .X(_2315_));
 sg13g2_buf_2 _6725_ (.A(\i_delta_sigma.sample[10] ),
    .X(_2316_));
 sg13g2_inv_1 _6726_ (.Y(_2317_),
    .A(_2316_));
 sg13g2_buf_2 _6727_ (.A(\i_delta_sigma.sample[9] ),
    .X(_2318_));
 sg13g2_inv_1 _6728_ (.Y(_2319_),
    .A(_2318_));
 sg13g2_nand2_1 _6729_ (.Y(_2320_),
    .A(_2317_),
    .B(_2319_));
 sg13g2_nand3_1 _6730_ (.B(_2316_),
    .C(_2318_),
    .A(_2315_),
    .Y(_2321_));
 sg13g2_o21ai_1 _6731_ (.B1(_2321_),
    .Y(_2322_),
    .A1(_2315_),
    .A2(_2320_));
 sg13g2_nand2_1 _6732_ (.Y(_2323_),
    .A(_2314_),
    .B(_2322_));
 sg13g2_buf_2 _6733_ (.A(_2323_),
    .X(_2324_));
 sg13g2_mux2_1 _6734_ (.A0(_0041_),
    .A1(_0040_),
    .S(_2324_),
    .X(_2325_));
 sg13g2_nor2_1 _6735_ (.A(_2308_),
    .B(_2325_),
    .Y(_2326_));
 sg13g2_inv_1 _6736_ (.Y(_2327_),
    .A(_2292_));
 sg13g2_a21o_1 _6737_ (.A2(_2308_),
    .A1(_2325_),
    .B1(_2327_),
    .X(_2328_));
 sg13g2_buf_2 _6738_ (.A(\i_delta_sigma.sample[4] ),
    .X(_2329_));
 sg13g2_xnor2_1 _6739_ (.Y(_2330_),
    .A(_2329_),
    .B(\i_resonator.v[0] ));
 sg13g2_buf_1 _6740_ (.A(net174),
    .X(_2331_));
 sg13g2_buf_1 _6741_ (.A(net175),
    .X(_2332_));
 sg13g2_inv_2 _6742_ (.Y(_2333_),
    .A(net154));
 sg13g2_buf_1 _6743_ (.A(_2333_),
    .X(_2334_));
 sg13g2_inv_1 _6744_ (.Y(_2335_),
    .A(net174));
 sg13g2_buf_1 _6745_ (.A(_2335_),
    .X(_2336_));
 sg13g2_inv_1 _6746_ (.Y(_2337_),
    .A(_2310_));
 sg13g2_inv_1 _6747_ (.Y(_2338_),
    .A(_2312_));
 sg13g2_nand2_1 _6748_ (.Y(_2339_),
    .A(_2337_),
    .B(_2338_));
 sg13g2_xnor2_1 _6749_ (.Y(_2340_),
    .A(net155),
    .B(_2310_));
 sg13g2_o21ai_1 _6750_ (.B1(_2340_),
    .Y(_2341_),
    .A1(net138),
    .A2(_2312_));
 sg13g2_inv_1 _6751_ (.Y(_2342_),
    .A(_2341_));
 sg13g2_inv_1 _6752_ (.Y(_2343_),
    .A(\i_resonator.v[5] ));
 sg13g2_nor2_1 _6753_ (.A(_2318_),
    .B(_2343_),
    .Y(_2344_));
 sg13g2_buf_2 _6754_ (.A(\i_delta_sigma.sample[6] ),
    .X(_2345_));
 sg13g2_nor2b_1 _6755_ (.A(\i_resonator.v[2] ),
    .B_N(_2345_),
    .Y(_2346_));
 sg13g2_buf_2 _6756_ (.A(\i_delta_sigma.sample[5] ),
    .X(_2347_));
 sg13g2_xnor2_1 _6757_ (.Y(_2348_),
    .A(_2347_),
    .B(\i_resonator.v[1] ));
 sg13g2_nor2b_1 _6758_ (.A(\i_resonator.v[0] ),
    .B_N(_2329_),
    .Y(_2349_));
 sg13g2_inv_1 _6759_ (.Y(_2350_),
    .A(_2349_));
 sg13g2_inv_1 _6760_ (.Y(_2351_),
    .A(\i_resonator.v[1] ));
 sg13g2_nor2_1 _6761_ (.A(_2347_),
    .B(_2351_),
    .Y(_2352_));
 sg13g2_a21oi_1 _6762_ (.A1(_2348_),
    .A2(_2350_),
    .Y(_2353_),
    .B1(_2352_));
 sg13g2_inv_1 _6763_ (.Y(_2354_),
    .A(\i_resonator.v[2] ));
 sg13g2_nor2_1 _6764_ (.A(_2345_),
    .B(_2354_),
    .Y(_2355_));
 sg13g2_inv_1 _6765_ (.Y(_2356_),
    .A(_2355_));
 sg13g2_o21ai_1 _6766_ (.B1(_2356_),
    .Y(_2357_),
    .A1(_2346_),
    .A2(_2353_));
 sg13g2_buf_2 _6767_ (.A(\i_delta_sigma.sample[7] ),
    .X(_2358_));
 sg13g2_inv_1 _6768_ (.Y(_2359_),
    .A(_2358_));
 sg13g2_nor2_1 _6769_ (.A(\i_resonator.v[3] ),
    .B(_2359_),
    .Y(_2360_));
 sg13g2_inv_1 _6770_ (.Y(_2361_),
    .A(_2360_));
 sg13g2_inv_1 _6771_ (.Y(_2362_),
    .A(\i_resonator.v[3] ));
 sg13g2_nor2_1 _6772_ (.A(_2358_),
    .B(_2362_),
    .Y(_2363_));
 sg13g2_a21oi_1 _6773_ (.A1(_2357_),
    .A2(_2361_),
    .Y(_2364_),
    .B1(_2363_));
 sg13g2_buf_2 _6774_ (.A(\i_delta_sigma.sample[8] ),
    .X(_2365_));
 sg13g2_inv_1 _6775_ (.Y(_2366_),
    .A(\i_resonator.v[4] ));
 sg13g2_nor2_1 _6776_ (.A(_2365_),
    .B(_2366_),
    .Y(_2367_));
 sg13g2_inv_1 _6777_ (.Y(_2368_),
    .A(_2367_));
 sg13g2_inv_1 _6778_ (.Y(_2369_),
    .A(_2365_));
 sg13g2_nor2_1 _6779_ (.A(\i_resonator.v[4] ),
    .B(_2369_),
    .Y(_2370_));
 sg13g2_a21oi_1 _6780_ (.A1(_2364_),
    .A2(_2368_),
    .Y(_2371_),
    .B1(_2370_));
 sg13g2_nor2_1 _6781_ (.A(\i_resonator.v[5] ),
    .B(_2319_),
    .Y(_2372_));
 sg13g2_inv_1 _6782_ (.Y(_2373_),
    .A(_2372_));
 sg13g2_o21ai_1 _6783_ (.B1(_2373_),
    .Y(_2374_),
    .A1(_2344_),
    .A2(_2371_));
 sg13g2_buf_2 _6784_ (.A(\i_resonator.v[6] ),
    .X(_2375_));
 sg13g2_inv_1 _6785_ (.Y(_2376_),
    .A(_2375_));
 sg13g2_nor2_1 _6786_ (.A(_2316_),
    .B(_2376_),
    .Y(_2377_));
 sg13g2_inv_1 _6787_ (.Y(_2378_),
    .A(_2377_));
 sg13g2_nor2_1 _6788_ (.A(_2375_),
    .B(_2317_),
    .Y(_2379_));
 sg13g2_a21oi_1 _6789_ (.A1(_2374_),
    .A2(_2378_),
    .Y(_2380_),
    .B1(_2379_));
 sg13g2_buf_2 _6790_ (.A(\i_resonator.v[7] ),
    .X(_2381_));
 sg13g2_nor2_1 _6791_ (.A(_2381_),
    .B(_2335_),
    .Y(_2382_));
 sg13g2_inv_1 _6792_ (.Y(_2383_),
    .A(_2381_));
 sg13g2_nor2_1 _6793_ (.A(net174),
    .B(_2383_),
    .Y(_2384_));
 sg13g2_nor2_1 _6794_ (.A(_2382_),
    .B(_2384_),
    .Y(_2385_));
 sg13g2_buf_2 _6795_ (.A(\i_resonator.v[8] ),
    .X(_2386_));
 sg13g2_xnor2_1 _6796_ (.Y(_2387_),
    .A(net174),
    .B(_2386_));
 sg13g2_nand3_1 _6797_ (.B(_2385_),
    .C(_2387_),
    .A(_2380_),
    .Y(_2388_));
 sg13g2_o21ai_1 _6798_ (.B1(_2335_),
    .Y(_2389_),
    .A1(_2386_),
    .A2(_2381_));
 sg13g2_nand2_1 _6799_ (.Y(_2390_),
    .A(_2388_),
    .B(_2389_));
 sg13g2_buf_1 _6800_ (.A(\i_resonator.v[10] ),
    .X(_2391_));
 sg13g2_xnor2_1 _6801_ (.Y(_2392_),
    .A(net174),
    .B(net173));
 sg13g2_buf_2 _6802_ (.A(\i_resonator.v[9] ),
    .X(_2393_));
 sg13g2_xnor2_1 _6803_ (.Y(_2394_),
    .A(net174),
    .B(_2393_));
 sg13g2_nand3_1 _6804_ (.B(_2392_),
    .C(_2394_),
    .A(_2390_),
    .Y(_2395_));
 sg13g2_o21ai_1 _6805_ (.B1(_2335_),
    .Y(_2396_),
    .A1(net173),
    .A2(_2393_));
 sg13g2_nand2_1 _6806_ (.Y(_2397_),
    .A(_2395_),
    .B(_2396_));
 sg13g2_buf_1 _6807_ (.A(\i_resonator.v[12] ),
    .X(_2398_));
 sg13g2_xnor2_1 _6808_ (.Y(_2399_),
    .A(net174),
    .B(net172));
 sg13g2_buf_1 _6809_ (.A(\i_resonator.v[11] ),
    .X(_2400_));
 sg13g2_xnor2_1 _6810_ (.Y(_2401_),
    .A(net174),
    .B(net171));
 sg13g2_nand3_1 _6811_ (.B(_2399_),
    .C(_2401_),
    .A(_2397_),
    .Y(_2402_));
 sg13g2_o21ai_1 _6812_ (.B1(_2335_),
    .Y(_2403_),
    .A1(net172),
    .A2(net171));
 sg13g2_nand2_1 _6813_ (.Y(_2404_),
    .A(_2402_),
    .B(_2403_));
 sg13g2_a22oi_1 _6814_ (.Y(_2405_),
    .B1(_2342_),
    .B2(_2404_),
    .A2(_2339_),
    .A1(net138));
 sg13g2_inv_1 _6815_ (.Y(_2406_),
    .A(_2405_));
 sg13g2_nor3_1 _6816_ (.A(net155),
    .B(_2334_),
    .C(_2406_),
    .Y(_2407_));
 sg13g2_buf_1 _6817_ (.A(_2407_),
    .X(_2408_));
 sg13g2_buf_1 _6818_ (.A(net154),
    .X(_2409_));
 sg13g2_nor3_1 _6819_ (.A(net138),
    .B(net137),
    .C(_2405_),
    .Y(_2410_));
 sg13g2_nor2_2 _6820_ (.A(net156),
    .B(_2410_),
    .Y(_2411_));
 sg13g2_o21ai_1 _6821_ (.B1(_2411_),
    .Y(_2412_),
    .A1(_2330_),
    .A2(net61));
 sg13g2_o21ai_1 _6822_ (.B1(_2412_),
    .Y(_2413_),
    .A1(_2326_),
    .A2(_2328_));
 sg13g2_buf_1 _6823_ (.A(_2282_),
    .X(_2414_));
 sg13g2_buf_1 _6824_ (.A(_2273_),
    .X(_2415_));
 sg13g2_o21ai_1 _6825_ (.B1(net120),
    .Y(_2416_),
    .A1(\i_resonator.v[0] ),
    .A2(net108));
 sg13g2_a21oi_1 _6826_ (.A1(_2413_),
    .A2(net108),
    .Y(_0184_),
    .B1(_2416_));
 sg13g2_o21ai_1 _6827_ (.B1(net120),
    .Y(_2417_),
    .A1(net173),
    .A2(net108));
 sg13g2_nor2_1 _6828_ (.A(_2381_),
    .B(_2333_),
    .Y(_2418_));
 sg13g2_inv_1 _6829_ (.Y(_2419_),
    .A(_0042_));
 sg13g2_nor2_1 _6830_ (.A(_2419_),
    .B(_2324_),
    .Y(_2420_));
 sg13g2_a21oi_1 _6831_ (.A1(_0043_),
    .A2(_2324_),
    .Y(_2421_),
    .B1(_2420_));
 sg13g2_xnor2_1 _6832_ (.Y(_2422_),
    .A(_2366_),
    .B(_2421_));
 sg13g2_nor2_1 _6833_ (.A(net172),
    .B(_2324_),
    .Y(_2423_));
 sg13g2_a21o_1 _6834_ (.A2(_2324_),
    .A1(_2337_),
    .B1(_2423_),
    .X(_2424_));
 sg13g2_nor2_1 _6835_ (.A(\i_resonator.v[3] ),
    .B(_2424_),
    .Y(_2425_));
 sg13g2_nand2_1 _6836_ (.Y(_2426_),
    .A(_2324_),
    .B(_2419_));
 sg13g2_o21ai_1 _6837_ (.B1(_2426_),
    .Y(_2427_),
    .A1(_0040_),
    .A2(_2324_));
 sg13g2_nor2_1 _6838_ (.A(_2354_),
    .B(_2427_),
    .Y(_2428_));
 sg13g2_xnor2_1 _6839_ (.Y(_2429_),
    .A(\i_resonator.v[2] ),
    .B(_2427_));
 sg13g2_inv_1 _6840_ (.Y(_2430_),
    .A(_2429_));
 sg13g2_mux2_1 _6841_ (.A0(_2391_),
    .A1(_2398_),
    .S(_2324_),
    .X(_2431_));
 sg13g2_nor2_1 _6842_ (.A(_2351_),
    .B(_2431_),
    .Y(_2432_));
 sg13g2_xnor2_1 _6843_ (.Y(_2433_),
    .A(_2351_),
    .B(_2431_));
 sg13g2_nor2_1 _6844_ (.A(_2326_),
    .B(_2433_),
    .Y(_2434_));
 sg13g2_nor2_1 _6845_ (.A(_2432_),
    .B(_2434_),
    .Y(_2435_));
 sg13g2_nor2_1 _6846_ (.A(_2430_),
    .B(_2435_),
    .Y(_2436_));
 sg13g2_nor2_1 _6847_ (.A(_2428_),
    .B(_2436_),
    .Y(_2437_));
 sg13g2_inv_1 _6848_ (.Y(_2438_),
    .A(_2424_));
 sg13g2_nor2_1 _6849_ (.A(_2362_),
    .B(_2438_),
    .Y(_2439_));
 sg13g2_inv_1 _6850_ (.Y(_2440_),
    .A(_2439_));
 sg13g2_o21ai_1 _6851_ (.B1(_2440_),
    .Y(_2441_),
    .A1(_2425_),
    .A2(_2437_));
 sg13g2_nand2b_1 _6852_ (.Y(_2442_),
    .B(_2441_),
    .A_N(_2422_));
 sg13g2_nor2_1 _6853_ (.A(net175),
    .B(_2343_),
    .Y(_2443_));
 sg13g2_nor2_1 _6854_ (.A(_2366_),
    .B(_2421_),
    .Y(_2444_));
 sg13g2_nor2_1 _6855_ (.A(_2443_),
    .B(_2444_),
    .Y(_2445_));
 sg13g2_nor2_1 _6856_ (.A(\i_resonator.v[5] ),
    .B(_2333_),
    .Y(_2446_));
 sg13g2_a21oi_1 _6857_ (.A1(_2442_),
    .A2(_2445_),
    .Y(_2447_),
    .B1(_2446_));
 sg13g2_xnor2_1 _6858_ (.Y(_2448_),
    .A(net154),
    .B(_2375_));
 sg13g2_nand2_1 _6859_ (.Y(_2449_),
    .A(_2447_),
    .B(_2448_));
 sg13g2_o21ai_1 _6860_ (.B1(_2333_),
    .Y(_2450_),
    .A1(_2381_),
    .A2(_2375_));
 sg13g2_o21ai_1 _6861_ (.B1(_2450_),
    .Y(_2451_),
    .A1(_2418_),
    .A2(_2449_));
 sg13g2_xnor2_1 _6862_ (.Y(_2452_),
    .A(net154),
    .B(_2393_));
 sg13g2_xnor2_1 _6863_ (.Y(_2453_),
    .A(net154),
    .B(_2386_));
 sg13g2_nand3_1 _6864_ (.B(_2452_),
    .C(_2453_),
    .A(_2451_),
    .Y(_2454_));
 sg13g2_o21ai_1 _6865_ (.B1(net130),
    .Y(_2455_),
    .A1(_2393_),
    .A2(_2386_));
 sg13g2_nand2_1 _6866_ (.Y(_2456_),
    .A(_2454_),
    .B(_2455_));
 sg13g2_xnor2_1 _6867_ (.Y(_2457_),
    .A(net173),
    .B(net154));
 sg13g2_o21ai_1 _6868_ (.B1(net156),
    .Y(_2458_),
    .A1(_2457_),
    .A2(_2456_));
 sg13g2_a21oi_1 _6869_ (.A1(_2456_),
    .A2(_2457_),
    .Y(_2459_),
    .B1(_2458_));
 sg13g2_inv_1 _6870_ (.Y(_2460_),
    .A(net61));
 sg13g2_nand2_1 _6871_ (.Y(_2461_),
    .A(_2394_),
    .B(_2387_));
 sg13g2_a21oi_1 _6872_ (.A1(_2385_),
    .A2(_2377_),
    .Y(_2462_),
    .B1(_2384_));
 sg13g2_o21ai_1 _6873_ (.B1(net138),
    .Y(_2463_),
    .A1(_2393_),
    .A2(_2386_));
 sg13g2_o21ai_1 _6874_ (.B1(_2463_),
    .Y(_2464_),
    .A1(_2461_),
    .A2(_2462_));
 sg13g2_nor2_1 _6875_ (.A(_2377_),
    .B(_2379_),
    .Y(_2465_));
 sg13g2_inv_1 _6876_ (.Y(_2466_),
    .A(_2465_));
 sg13g2_nor4_1 _6877_ (.A(_2382_),
    .B(_2384_),
    .C(_2466_),
    .D(_2374_),
    .Y(_2467_));
 sg13g2_nand2b_1 _6878_ (.Y(_2468_),
    .B(_2467_),
    .A_N(_2461_));
 sg13g2_nand2b_1 _6879_ (.Y(_2469_),
    .B(_2468_),
    .A_N(_2464_));
 sg13g2_xor2_1 _6880_ (.B(_2469_),
    .A(_2392_),
    .X(_2470_));
 sg13g2_nand2_1 _6881_ (.Y(_2471_),
    .A(_2460_),
    .B(_2470_));
 sg13g2_inv_1 _6882_ (.Y(_2472_),
    .A(_2410_));
 sg13g2_a21oi_1 _6883_ (.A1(_2471_),
    .A2(net67),
    .Y(_2473_),
    .B1(net156));
 sg13g2_nor3_1 _6884_ (.A(net90),
    .B(_2459_),
    .C(_2473_),
    .Y(_2474_));
 sg13g2_nor2_1 _6885_ (.A(_2417_),
    .B(_2474_),
    .Y(_0185_));
 sg13g2_o21ai_1 _6886_ (.B1(net120),
    .Y(_2475_),
    .A1(_2400_),
    .A2(net108));
 sg13g2_inv_1 _6887_ (.Y(_2476_),
    .A(_2437_));
 sg13g2_nor3_1 _6888_ (.A(_2425_),
    .B(_2422_),
    .C(_2439_),
    .Y(_2477_));
 sg13g2_inv_1 _6889_ (.Y(_2478_),
    .A(_2444_));
 sg13g2_o21ai_1 _6890_ (.B1(_2478_),
    .Y(_2479_),
    .A1(_2422_),
    .A2(_2440_));
 sg13g2_a21oi_1 _6891_ (.A1(_2476_),
    .A2(_2477_),
    .Y(_2480_),
    .B1(_2479_));
 sg13g2_inv_1 _6892_ (.Y(_2481_),
    .A(_2480_));
 sg13g2_nor2_1 _6893_ (.A(_2446_),
    .B(_2443_),
    .Y(_2482_));
 sg13g2_nand3_1 _6894_ (.B(_2448_),
    .C(_2482_),
    .A(_2481_),
    .Y(_2483_));
 sg13g2_o21ai_1 _6895_ (.B1(_2333_),
    .Y(_2484_),
    .A1(_2375_),
    .A2(\i_resonator.v[5] ));
 sg13g2_nand2_1 _6896_ (.Y(_2485_),
    .A(_2483_),
    .B(_2484_));
 sg13g2_xnor2_1 _6897_ (.Y(_2486_),
    .A(net154),
    .B(_2381_));
 sg13g2_nand2_1 _6898_ (.Y(_2487_),
    .A(_2486_),
    .B(_2453_));
 sg13g2_inv_1 _6899_ (.Y(_2488_),
    .A(_2452_));
 sg13g2_inv_1 _6900_ (.Y(_2489_),
    .A(_2457_));
 sg13g2_nor2_1 _6901_ (.A(_2488_),
    .B(_2489_),
    .Y(_2490_));
 sg13g2_inv_1 _6902_ (.Y(_2491_),
    .A(_2490_));
 sg13g2_nor2_1 _6903_ (.A(_2487_),
    .B(_2491_),
    .Y(_2492_));
 sg13g2_o21ai_1 _6904_ (.B1(_2333_),
    .Y(_2493_),
    .A1(_2386_),
    .A2(_2381_));
 sg13g2_inv_1 _6905_ (.Y(_2494_),
    .A(_2493_));
 sg13g2_o21ai_1 _6906_ (.B1(_2333_),
    .Y(_2495_),
    .A1(net173),
    .A2(_2393_));
 sg13g2_inv_1 _6907_ (.Y(_2496_),
    .A(_2495_));
 sg13g2_a21oi_1 _6908_ (.A1(_2490_),
    .A2(_2494_),
    .Y(_2497_),
    .B1(_2496_));
 sg13g2_inv_1 _6909_ (.Y(_2498_),
    .A(_2497_));
 sg13g2_a21oi_1 _6910_ (.A1(_2485_),
    .A2(_2492_),
    .Y(_2499_),
    .B1(_2498_));
 sg13g2_xnor2_1 _6911_ (.Y(_2500_),
    .A(net137),
    .B(net171));
 sg13g2_inv_1 _6912_ (.Y(_2501_),
    .A(_2500_));
 sg13g2_o21ai_1 _6913_ (.B1(net156),
    .Y(_2502_),
    .A1(_2501_),
    .A2(_2499_));
 sg13g2_a21oi_1 _6914_ (.A1(_2499_),
    .A2(_2501_),
    .Y(_2503_),
    .B1(_2502_));
 sg13g2_xor2_1 _6915_ (.B(_2397_),
    .A(_2401_),
    .X(_2504_));
 sg13g2_nand2_1 _6916_ (.Y(_2505_),
    .A(_2460_),
    .B(_2504_));
 sg13g2_a21oi_1 _6917_ (.A1(_2505_),
    .A2(net67),
    .Y(_2506_),
    .B1(net156));
 sg13g2_nor3_1 _6918_ (.A(net94),
    .B(_2503_),
    .C(_2506_),
    .Y(_2507_));
 sg13g2_nor2_1 _6919_ (.A(_2475_),
    .B(_2507_),
    .Y(_0186_));
 sg13g2_xnor2_1 _6920_ (.Y(_2508_),
    .A(net137),
    .B(net172));
 sg13g2_inv_1 _6921_ (.Y(_2509_),
    .A(_2508_));
 sg13g2_nand3_1 _6922_ (.B(_2457_),
    .C(_2500_),
    .A(_2456_),
    .Y(_2510_));
 sg13g2_o21ai_1 _6923_ (.B1(net130),
    .Y(_2511_),
    .A1(net173),
    .A2(net171));
 sg13g2_nand2_1 _6924_ (.Y(_2512_),
    .A(_2510_),
    .B(_2511_));
 sg13g2_xnor2_1 _6925_ (.Y(_2513_),
    .A(_2509_),
    .B(_2512_));
 sg13g2_a21oi_1 _6926_ (.A1(_2513_),
    .A2(net139),
    .Y(_2514_),
    .B1(net90));
 sg13g2_nor2b_1 _6927_ (.A(_2467_),
    .B_N(_2462_),
    .Y(_2515_));
 sg13g2_inv_1 _6928_ (.Y(_2516_),
    .A(_2515_));
 sg13g2_nand2_1 _6929_ (.Y(_2517_),
    .A(_2401_),
    .B(_2392_));
 sg13g2_nor2_1 _6930_ (.A(_2517_),
    .B(_2461_),
    .Y(_2518_));
 sg13g2_o21ai_1 _6931_ (.B1(net138),
    .Y(_2519_),
    .A1(net173),
    .A2(net171));
 sg13g2_o21ai_1 _6932_ (.B1(_2519_),
    .Y(_2520_),
    .A1(_2463_),
    .A2(_2517_));
 sg13g2_a21oi_1 _6933_ (.A1(_2516_),
    .A2(_2518_),
    .Y(_2521_),
    .B1(_2520_));
 sg13g2_xnor2_1 _6934_ (.Y(_2522_),
    .A(_2399_),
    .B(_2521_));
 sg13g2_nand2_1 _6935_ (.Y(_2523_),
    .A(_2460_),
    .B(_2522_));
 sg13g2_a21o_1 _6936_ (.A2(net67),
    .A1(_2523_),
    .B1(net139),
    .X(_2524_));
 sg13g2_o21ai_1 _6937_ (.B1(net120),
    .Y(_2525_),
    .A1(net172),
    .A2(_2414_));
 sg13g2_a21oi_1 _6938_ (.A1(_2514_),
    .A2(_2524_),
    .Y(_0187_),
    .B1(_2525_));
 sg13g2_xnor2_1 _6939_ (.Y(_2526_),
    .A(net155),
    .B(_2312_));
 sg13g2_xnor2_1 _6940_ (.Y(_2527_),
    .A(_2526_),
    .B(_2404_));
 sg13g2_o21ai_1 _6941_ (.B1(_2411_),
    .Y(_2528_),
    .A1(_2527_),
    .A2(net61));
 sg13g2_nor2_1 _6942_ (.A(_2501_),
    .B(_2509_),
    .Y(_2529_));
 sg13g2_o21ai_1 _6943_ (.B1(_2493_),
    .Y(_2530_),
    .A1(_2484_),
    .A2(_2487_));
 sg13g2_nor2_1 _6944_ (.A(_2487_),
    .B(_2483_),
    .Y(_2531_));
 sg13g2_nor2_1 _6945_ (.A(_2530_),
    .B(_2531_),
    .Y(_2532_));
 sg13g2_inv_1 _6946_ (.Y(_2533_),
    .A(_2532_));
 sg13g2_inv_1 _6947_ (.Y(_2534_),
    .A(_2529_));
 sg13g2_nor2_1 _6948_ (.A(_2491_),
    .B(_2534_),
    .Y(_2535_));
 sg13g2_o21ai_1 _6949_ (.B1(net130),
    .Y(_2536_),
    .A1(net172),
    .A2(net171));
 sg13g2_inv_1 _6950_ (.Y(_2537_),
    .A(_2536_));
 sg13g2_a221oi_1 _6951_ (.B2(_2535_),
    .C1(_2537_),
    .B1(_2533_),
    .A1(_2496_),
    .Y(_2538_),
    .A2(_2529_));
 sg13g2_a21oi_1 _6952_ (.A1(_2538_),
    .A2(_2313_),
    .Y(_2539_),
    .B1(_2327_));
 sg13g2_o21ai_1 _6953_ (.B1(_2539_),
    .Y(_2540_),
    .A1(_2313_),
    .A2(_2538_));
 sg13g2_nand3_1 _6954_ (.B(_2540_),
    .C(_2282_),
    .A(_2528_),
    .Y(_2541_));
 sg13g2_nand2_1 _6955_ (.Y(_2542_),
    .A(net90),
    .B(_2312_));
 sg13g2_a21oi_1 _6956_ (.A1(_2541_),
    .A2(_2542_),
    .Y(_0188_),
    .B1(net109));
 sg13g2_nand2_1 _6957_ (.Y(_2543_),
    .A(_2313_),
    .B(_2508_));
 sg13g2_nor2_1 _6958_ (.A(net137),
    .B(_2338_),
    .Y(_2544_));
 sg13g2_inv_1 _6959_ (.Y(_2545_),
    .A(_2544_));
 sg13g2_o21ai_1 _6960_ (.B1(_2545_),
    .Y(_2546_),
    .A1(_2511_),
    .A2(_2543_));
 sg13g2_a21oi_1 _6961_ (.A1(net130),
    .A2(net172),
    .Y(_2547_),
    .B1(_2546_));
 sg13g2_o21ai_1 _6962_ (.B1(_2547_),
    .Y(_2548_),
    .A1(_2543_),
    .A2(_2510_));
 sg13g2_xnor2_1 _6963_ (.Y(_2549_),
    .A(_2311_),
    .B(_2548_));
 sg13g2_a21oi_1 _6964_ (.A1(_2549_),
    .A2(net139),
    .Y(_2550_),
    .B1(_2298_));
 sg13g2_nand2_1 _6965_ (.Y(_2551_),
    .A(_2526_),
    .B(_2399_));
 sg13g2_o21ai_1 _6966_ (.B1(net138),
    .Y(_2552_),
    .A1(_2312_),
    .A2(net172));
 sg13g2_o21ai_1 _6967_ (.B1(_2552_),
    .Y(_2553_),
    .A1(_2551_),
    .A2(_2521_));
 sg13g2_xor2_1 _6968_ (.B(_2553_),
    .A(_2340_),
    .X(_2554_));
 sg13g2_nand2_1 _6969_ (.Y(_2555_),
    .A(_2460_),
    .B(_2554_));
 sg13g2_a21o_1 _6970_ (.A2(_2472_),
    .A1(_2555_),
    .B1(net139),
    .X(_2556_));
 sg13g2_a221oi_1 _6971_ (.B2(_2556_),
    .C1(net109),
    .B1(_2550_),
    .A1(_2337_),
    .Y(_0189_),
    .A2(_2299_));
 sg13g2_xnor2_1 _6972_ (.Y(_2557_),
    .A(net155),
    .B(net137));
 sg13g2_nor2_1 _6973_ (.A(_2409_),
    .B(net138),
    .Y(_2558_));
 sg13g2_a21oi_1 _6974_ (.A1(_2406_),
    .A2(_2557_),
    .Y(_2559_),
    .B1(_2558_));
 sg13g2_buf_1 _6975_ (.A(_2327_),
    .X(_2560_));
 sg13g2_nand2_1 _6976_ (.Y(_2561_),
    .A(_2559_),
    .B(net136));
 sg13g2_inv_1 _6977_ (.Y(_2562_),
    .A(_2499_));
 sg13g2_nor2b_1 _6978_ (.A(_2534_),
    .B_N(_2314_),
    .Y(_2563_));
 sg13g2_nand2_1 _6979_ (.Y(_2564_),
    .A(net130),
    .B(_2310_));
 sg13g2_nand3_1 _6980_ (.B(net156),
    .C(_2564_),
    .A(_2545_),
    .Y(_2565_));
 sg13g2_a221oi_1 _6981_ (.B2(_2563_),
    .C1(_2565_),
    .B1(_2562_),
    .A1(_2314_),
    .Y(_2566_),
    .A2(_2537_));
 sg13g2_nor2_1 _6982_ (.A(net94),
    .B(_2566_),
    .Y(_2567_));
 sg13g2_a221oi_1 _6983_ (.B2(_2567_),
    .C1(net109),
    .B1(_2561_),
    .A1(net130),
    .Y(_0190_),
    .A2(net90));
 sg13g2_xor2_1 _6984_ (.B(_2433_),
    .A(_2326_),
    .X(_2568_));
 sg13g2_xnor2_1 _6985_ (.Y(_2569_),
    .A(_2350_),
    .B(_2348_));
 sg13g2_o21ai_1 _6986_ (.B1(_2411_),
    .Y(_2570_),
    .A1(_2569_),
    .A2(_2408_));
 sg13g2_o21ai_1 _6987_ (.B1(_2570_),
    .Y(_2571_),
    .A1(_2560_),
    .A2(_2568_));
 sg13g2_o21ai_1 _6988_ (.B1(_2415_),
    .Y(_2572_),
    .A1(\i_resonator.v[1] ),
    .A2(_2414_));
 sg13g2_a21oi_1 _6989_ (.A1(_2571_),
    .A2(net108),
    .Y(_0191_),
    .B1(_2572_));
 sg13g2_nor2_1 _6990_ (.A(_2355_),
    .B(_2346_),
    .Y(_2573_));
 sg13g2_xor2_1 _6991_ (.B(_2353_),
    .A(_2573_),
    .X(_2574_));
 sg13g2_o21ai_1 _6992_ (.B1(net67),
    .Y(_2575_),
    .A1(_2574_),
    .A2(_2408_));
 sg13g2_nand2_1 _6993_ (.Y(_2576_),
    .A(_2575_),
    .B(_2560_));
 sg13g2_nor2_1 _6994_ (.A(net136),
    .B(_2436_),
    .Y(_2577_));
 sg13g2_nand2_1 _6995_ (.Y(_2578_),
    .A(_2435_),
    .B(_2430_));
 sg13g2_a21oi_1 _6996_ (.A1(_2577_),
    .A2(_2578_),
    .Y(_2579_),
    .B1(net94));
 sg13g2_a221oi_1 _6997_ (.B2(_2579_),
    .C1(net109),
    .B1(_2576_),
    .A1(_2354_),
    .Y(_0192_),
    .A2(net90));
 sg13g2_nor2_1 _6998_ (.A(_2363_),
    .B(_2360_),
    .Y(_2580_));
 sg13g2_xnor2_1 _6999_ (.Y(_2581_),
    .A(_2580_),
    .B(_2357_));
 sg13g2_o21ai_1 _7000_ (.B1(_2472_),
    .Y(_2582_),
    .A1(_2581_),
    .A2(net61));
 sg13g2_nand2_1 _7001_ (.Y(_2583_),
    .A(_2582_),
    .B(net136));
 sg13g2_nor2_1 _7002_ (.A(_2425_),
    .B(_2439_),
    .Y(_2584_));
 sg13g2_xnor2_1 _7003_ (.Y(_2585_),
    .A(_2584_),
    .B(_2437_));
 sg13g2_a21oi_1 _7004_ (.A1(_2585_),
    .A2(net139),
    .Y(_2586_),
    .B1(net94));
 sg13g2_a221oi_1 _7005_ (.B2(_2586_),
    .C1(net109),
    .B1(_2583_),
    .A1(_2362_),
    .Y(_0193_),
    .A2(net90));
 sg13g2_xnor2_1 _7006_ (.Y(_2587_),
    .A(_2422_),
    .B(_2441_));
 sg13g2_nor2_1 _7007_ (.A(_2370_),
    .B(_2367_),
    .Y(_2588_));
 sg13g2_xor2_1 _7008_ (.B(_2364_),
    .A(_2588_),
    .X(_2589_));
 sg13g2_o21ai_1 _7009_ (.B1(_2411_),
    .Y(_2590_),
    .A1(_2589_),
    .A2(net61));
 sg13g2_o21ai_1 _7010_ (.B1(_2590_),
    .Y(_2591_),
    .A1(net136),
    .A2(_2587_));
 sg13g2_o21ai_1 _7011_ (.B1(net120),
    .Y(_2592_),
    .A1(\i_resonator.v[4] ),
    .A2(_2282_));
 sg13g2_a21oi_1 _7012_ (.A1(_2591_),
    .A2(net108),
    .Y(_0194_),
    .B1(_2592_));
 sg13g2_nor2_1 _7013_ (.A(_2372_),
    .B(_2344_),
    .Y(_2593_));
 sg13g2_xnor2_1 _7014_ (.Y(_2594_),
    .A(_2593_),
    .B(_2371_));
 sg13g2_o21ai_1 _7015_ (.B1(net67),
    .Y(_2595_),
    .A1(_2594_),
    .A2(net61));
 sg13g2_nand2_1 _7016_ (.Y(_2596_),
    .A(_2595_),
    .B(net136));
 sg13g2_a21oi_1 _7017_ (.A1(_2481_),
    .A2(_2482_),
    .Y(_2597_),
    .B1(net136));
 sg13g2_nand2b_1 _7018_ (.Y(_2598_),
    .B(_2480_),
    .A_N(_2482_));
 sg13g2_a21oi_1 _7019_ (.A1(_2597_),
    .A2(_2598_),
    .Y(_2599_),
    .B1(net94));
 sg13g2_a221oi_1 _7020_ (.B2(_2599_),
    .C1(net109),
    .B1(_2596_),
    .A1(_2343_),
    .Y(_0195_),
    .A2(net90));
 sg13g2_xor2_1 _7021_ (.B(_2447_),
    .A(_2448_),
    .X(_2600_));
 sg13g2_xnor2_1 _7022_ (.Y(_2601_),
    .A(_2466_),
    .B(_2374_));
 sg13g2_o21ai_1 _7023_ (.B1(_2411_),
    .Y(_2602_),
    .A1(_2601_),
    .A2(net61));
 sg13g2_o21ai_1 _7024_ (.B1(_2602_),
    .Y(_2603_),
    .A1(net136),
    .A2(_2600_));
 sg13g2_o21ai_1 _7025_ (.B1(net120),
    .Y(_2604_),
    .A1(_2375_),
    .A2(_2282_));
 sg13g2_a21oi_1 _7026_ (.A1(_2603_),
    .A2(net108),
    .Y(_0196_),
    .B1(_2604_));
 sg13g2_xnor2_1 _7027_ (.Y(_2605_),
    .A(_2385_),
    .B(_2380_));
 sg13g2_o21ai_1 _7028_ (.B1(net67),
    .Y(_2606_),
    .A1(_2605_),
    .A2(net61));
 sg13g2_nand2_1 _7029_ (.Y(_2607_),
    .A(_2606_),
    .B(net136));
 sg13g2_xor2_1 _7030_ (.B(_2485_),
    .A(_2486_),
    .X(_2608_));
 sg13g2_a21oi_1 _7031_ (.A1(_2608_),
    .A2(net139),
    .Y(_2609_),
    .B1(net94));
 sg13g2_a221oi_1 _7032_ (.B2(_2609_),
    .C1(net109),
    .B1(_2607_),
    .A1(_2383_),
    .Y(_0197_),
    .A2(net90));
 sg13g2_xnor2_1 _7033_ (.Y(_2610_),
    .A(_2387_),
    .B(_2515_));
 sg13g2_nand2_1 _7034_ (.Y(_2611_),
    .A(_2460_),
    .B(_2610_));
 sg13g2_a21o_1 _7035_ (.A2(net67),
    .A1(_2611_),
    .B1(net139),
    .X(_2612_));
 sg13g2_xor2_1 _7036_ (.B(_2451_),
    .A(_2453_),
    .X(_2613_));
 sg13g2_a21oi_1 _7037_ (.A1(_2613_),
    .A2(net139),
    .Y(_2614_),
    .B1(net94));
 sg13g2_o21ai_1 _7038_ (.B1(net120),
    .Y(_2615_),
    .A1(_2386_),
    .A2(_2282_));
 sg13g2_a21oi_1 _7039_ (.A1(_2612_),
    .A2(_2614_),
    .Y(_0198_),
    .B1(_2615_));
 sg13g2_o21ai_1 _7040_ (.B1(net120),
    .Y(_2616_),
    .A1(_2393_),
    .A2(net108));
 sg13g2_o21ai_1 _7041_ (.B1(net156),
    .Y(_2617_),
    .A1(_2488_),
    .A2(_2532_));
 sg13g2_a21oi_1 _7042_ (.A1(_2488_),
    .A2(_2532_),
    .Y(_2618_),
    .B1(_2617_));
 sg13g2_xor2_1 _7043_ (.B(_2390_),
    .A(_2394_),
    .X(_2619_));
 sg13g2_nand2_1 _7044_ (.Y(_2620_),
    .A(_2460_),
    .B(_2619_));
 sg13g2_a21oi_1 _7045_ (.A1(_2620_),
    .A2(net67),
    .Y(_2621_),
    .B1(net156));
 sg13g2_nor3_1 _7046_ (.A(net94),
    .B(_2618_),
    .C(_2621_),
    .Y(_2622_));
 sg13g2_nor2_1 _7047_ (.A(_2616_),
    .B(_2622_),
    .Y(_0199_));
 sg13g2_buf_1 _7048_ (.A(\i_delta_sigma.sample[0] ),
    .X(_2623_));
 sg13g2_inv_1 _7049_ (.Y(_2624_),
    .A(_2623_));
 sg13g2_inv_1 _7050_ (.Y(_2625_),
    .A(_2285_));
 sg13g2_a21oi_1 _7051_ (.A1(_2283_),
    .A2(_2625_),
    .Y(_2626_),
    .B1(_2270_));
 sg13g2_buf_1 _7052_ (.A(_2626_),
    .X(_2627_));
 sg13g2_xnor2_1 _7053_ (.Y(_2628_),
    .A(_2623_),
    .B(_2391_));
 sg13g2_xor2_1 _7054_ (.B(net154),
    .A(_2318_),
    .X(_2629_));
 sg13g2_nor2_1 _7055_ (.A(_2345_),
    .B(net175),
    .Y(_2630_));
 sg13g2_nand2_1 _7056_ (.Y(_2631_),
    .A(_2623_),
    .B(net173));
 sg13g2_buf_2 _7057_ (.A(\i_delta_sigma.sample[1] ),
    .X(_2632_));
 sg13g2_xor2_1 _7058_ (.B(net171),
    .A(_2632_),
    .X(_2633_));
 sg13g2_inv_1 _7059_ (.Y(_2634_),
    .A(_2633_));
 sg13g2_nand2_1 _7060_ (.Y(_2635_),
    .A(_2632_),
    .B(net171));
 sg13g2_o21ai_1 _7061_ (.B1(_2635_),
    .Y(_2636_),
    .A1(_2631_),
    .A2(_2634_));
 sg13g2_buf_1 _7062_ (.A(\i_delta_sigma.sample[2] ),
    .X(_2637_));
 sg13g2_nor2_1 _7063_ (.A(_2637_),
    .B(\i_resonator.v[12] ),
    .Y(_2638_));
 sg13g2_inv_1 _7064_ (.Y(_2639_),
    .A(_2638_));
 sg13g2_nand2_1 _7065_ (.Y(_2640_),
    .A(_2637_),
    .B(_2398_));
 sg13g2_inv_1 _7066_ (.Y(_2641_),
    .A(_2640_));
 sg13g2_a21oi_1 _7067_ (.A1(_2636_),
    .A2(_2639_),
    .Y(_2642_),
    .B1(_2641_));
 sg13g2_buf_1 _7068_ (.A(\i_delta_sigma.sample[3] ),
    .X(_2643_));
 sg13g2_nand2_1 _7069_ (.Y(_2644_),
    .A(_2643_),
    .B(_2312_));
 sg13g2_nor2_1 _7070_ (.A(_2643_),
    .B(_2312_),
    .Y(_2645_));
 sg13g2_a21oi_1 _7071_ (.A1(_2642_),
    .A2(_2644_),
    .Y(_2646_),
    .B1(_2645_));
 sg13g2_nor2_1 _7072_ (.A(_2329_),
    .B(_2310_),
    .Y(_2647_));
 sg13g2_inv_1 _7073_ (.Y(_2648_),
    .A(_2647_));
 sg13g2_nand2_1 _7074_ (.Y(_2649_),
    .A(_2329_),
    .B(_2310_));
 sg13g2_inv_1 _7075_ (.Y(_2650_),
    .A(_2649_));
 sg13g2_a21oi_1 _7076_ (.A1(_2646_),
    .A2(_2648_),
    .Y(_2651_),
    .B1(_2650_));
 sg13g2_nand2_1 _7077_ (.Y(_2652_),
    .A(_2347_),
    .B(net175));
 sg13g2_nor2_1 _7078_ (.A(_2347_),
    .B(net175),
    .Y(_2653_));
 sg13g2_a21oi_1 _7079_ (.A1(_2651_),
    .A2(_2652_),
    .Y(_2654_),
    .B1(_2653_));
 sg13g2_inv_1 _7080_ (.Y(_2655_),
    .A(_2654_));
 sg13g2_nand2_1 _7081_ (.Y(_2656_),
    .A(_2345_),
    .B(net175));
 sg13g2_o21ai_1 _7082_ (.B1(_2656_),
    .Y(_2657_),
    .A1(_2630_),
    .A2(_2655_));
 sg13g2_nor2_1 _7083_ (.A(_2365_),
    .B(_2309_),
    .Y(_2658_));
 sg13g2_inv_1 _7084_ (.Y(_2659_),
    .A(_2658_));
 sg13g2_xor2_1 _7085_ (.B(_2309_),
    .A(_2358_),
    .X(_2660_));
 sg13g2_nand3_1 _7086_ (.B(_2659_),
    .C(_2660_),
    .A(_2657_),
    .Y(_2661_));
 sg13g2_o21ai_1 _7087_ (.B1(_2332_),
    .Y(_2662_),
    .A1(_2365_),
    .A2(_2358_));
 sg13g2_nand2_1 _7088_ (.Y(_2663_),
    .A(_2661_),
    .B(_2662_));
 sg13g2_xor2_1 _7089_ (.B(_2332_),
    .A(_2316_),
    .X(_2664_));
 sg13g2_and2_1 _7090_ (.A(_2663_),
    .B(_2664_),
    .X(_2665_));
 sg13g2_a22oi_1 _7091_ (.Y(_2666_),
    .B1(_2629_),
    .B2(_2665_),
    .A2(_2320_),
    .A1(net137));
 sg13g2_nand3b_1 _7092_ (.B(_2336_),
    .C(_2334_),
    .Y(_2667_),
    .A_N(_2666_));
 sg13g2_buf_1 _7093_ (.A(_2667_),
    .X(_2668_));
 sg13g2_nand3_1 _7094_ (.B(net155),
    .C(net137),
    .A(_2666_),
    .Y(_2669_));
 sg13g2_nand2_1 _7095_ (.Y(_2670_),
    .A(_2668_),
    .B(_2669_));
 sg13g2_buf_1 _7096_ (.A(_2670_),
    .X(_2671_));
 sg13g2_buf_1 _7097_ (.A(_2668_),
    .X(_2672_));
 sg13g2_o21ai_1 _7098_ (.B1(net69),
    .Y(_2673_),
    .A1(_2628_),
    .A2(net66));
 sg13g2_inv_2 _7099_ (.Y(_2674_),
    .A(_2268_));
 sg13g2_nand2_1 _7100_ (.Y(_2675_),
    .A(_2673_),
    .B(_2674_));
 sg13g2_nor2_1 _7101_ (.A(\i_orchestrator.trigger_resonator[1] ),
    .B(_2626_),
    .Y(_2676_));
 sg13g2_buf_2 _7102_ (.A(_2676_),
    .X(_2677_));
 sg13g2_buf_1 _7103_ (.A(_2272_),
    .X(_2678_));
 sg13g2_a221oi_1 _7104_ (.B2(_2677_),
    .C1(net129),
    .B1(_2675_),
    .A1(_2624_),
    .Y(_0200_),
    .A2(net89));
 sg13g2_nor3_2 _7105_ (.A(_2268_),
    .B(_2285_),
    .C(_2282_),
    .Y(_2679_));
 sg13g2_nand2_1 _7106_ (.Y(_2680_),
    .A(_2365_),
    .B(_2409_));
 sg13g2_nand2_1 _7107_ (.Y(_2681_),
    .A(_2659_),
    .B(_2680_));
 sg13g2_inv_1 _7108_ (.Y(_2682_),
    .A(_2681_));
 sg13g2_nand2_1 _7109_ (.Y(_2683_),
    .A(_2682_),
    .B(_2629_));
 sg13g2_nor2b_1 _7110_ (.A(_2630_),
    .B_N(_2656_),
    .Y(_2684_));
 sg13g2_nand3_1 _7111_ (.B(_2660_),
    .C(_2684_),
    .A(_2654_),
    .Y(_2685_));
 sg13g2_a21oi_1 _7112_ (.A1(_2319_),
    .A2(_2369_),
    .Y(_2686_),
    .B1(net130));
 sg13g2_o21ai_1 _7113_ (.B1(net137),
    .Y(_2687_),
    .A1(_2358_),
    .A2(_2345_));
 sg13g2_nor2_1 _7114_ (.A(_2687_),
    .B(_2683_),
    .Y(_2688_));
 sg13g2_nor2_1 _7115_ (.A(_2686_),
    .B(_2688_),
    .Y(_2689_));
 sg13g2_o21ai_1 _7116_ (.B1(_2689_),
    .Y(_2690_),
    .A1(_2683_),
    .A2(_2685_));
 sg13g2_xnor2_1 _7117_ (.Y(_2691_),
    .A(_2664_),
    .B(_2690_));
 sg13g2_o21ai_1 _7118_ (.B1(net69),
    .Y(_2692_),
    .A1(_2691_),
    .A2(net66));
 sg13g2_a22oi_1 _7119_ (.Y(_2693_),
    .B1(_2679_),
    .B2(_2692_),
    .A2(net89),
    .A1(_2316_));
 sg13g2_inv_1 _7120_ (.Y(_2694_),
    .A(\i_orchestrator.trigger_resonator[1] ));
 sg13g2_a21oi_1 _7121_ (.A1(_2693_),
    .A2(_2694_),
    .Y(_0201_),
    .B1(_2678_));
 sg13g2_nand2_1 _7122_ (.Y(_2695_),
    .A(net138),
    .B(net130));
 sg13g2_o21ai_1 _7123_ (.B1(_2695_),
    .Y(_2696_),
    .A1(_2557_),
    .A2(_2666_));
 sg13g2_and3_1 _7124_ (.X(_2697_),
    .A(_2279_),
    .B(_2276_),
    .C(_2327_));
 sg13g2_o21ai_1 _7125_ (.B1(_2415_),
    .Y(_2698_),
    .A1(net155),
    .A2(_2697_));
 sg13g2_a21oi_1 _7126_ (.A1(_2696_),
    .A2(_2697_),
    .Y(_0202_),
    .B1(_2698_));
 sg13g2_xor2_1 _7127_ (.B(_2633_),
    .A(_2631_),
    .X(_2699_));
 sg13g2_o21ai_1 _7128_ (.B1(net69),
    .Y(_2700_),
    .A1(_2699_),
    .A2(net66));
 sg13g2_a22oi_1 _7129_ (.Y(_2701_),
    .B1(_2677_),
    .B2(_2700_),
    .A2(net89),
    .A1(_2632_));
 sg13g2_a21oi_1 _7130_ (.A1(_2701_),
    .A2(_2674_),
    .Y(_0203_),
    .B1(net129));
 sg13g2_inv_1 _7131_ (.Y(_2702_),
    .A(_2637_));
 sg13g2_nor2_1 _7132_ (.A(_2638_),
    .B(_2641_),
    .Y(_2703_));
 sg13g2_xnor2_1 _7133_ (.Y(_2704_),
    .A(_2703_),
    .B(_2636_));
 sg13g2_o21ai_1 _7134_ (.B1(_2668_),
    .Y(_2705_),
    .A1(_2704_),
    .A2(_2670_));
 sg13g2_nand2_1 _7135_ (.Y(_2706_),
    .A(_2705_),
    .B(_2674_));
 sg13g2_a221oi_1 _7136_ (.B2(_2677_),
    .C1(_2272_),
    .B1(_2706_),
    .A1(_2702_),
    .Y(_0204_),
    .A2(_2627_));
 sg13g2_nand2b_1 _7137_ (.Y(_2707_),
    .B(_2644_),
    .A_N(_2645_));
 sg13g2_xnor2_1 _7138_ (.Y(_2708_),
    .A(_2707_),
    .B(_2642_));
 sg13g2_o21ai_1 _7139_ (.B1(_2672_),
    .Y(_2709_),
    .A1(_2708_),
    .A2(_2671_));
 sg13g2_a22oi_1 _7140_ (.Y(_2710_),
    .B1(_2677_),
    .B2(_2709_),
    .A2(_2627_),
    .A1(_2643_));
 sg13g2_a21oi_1 _7141_ (.A1(_2710_),
    .A2(_2674_),
    .Y(_0205_),
    .B1(_2678_));
 sg13g2_nor2_1 _7142_ (.A(_2647_),
    .B(_2650_),
    .Y(_2711_));
 sg13g2_xnor2_1 _7143_ (.Y(_2712_),
    .A(_2711_),
    .B(_2646_));
 sg13g2_o21ai_1 _7144_ (.B1(net69),
    .Y(_2713_),
    .A1(_2712_),
    .A2(net66));
 sg13g2_a22oi_1 _7145_ (.Y(_2714_),
    .B1(_2679_),
    .B2(_2713_),
    .A2(net89),
    .A1(_2329_));
 sg13g2_a21oi_1 _7146_ (.A1(_2714_),
    .A2(_2694_),
    .Y(_0206_),
    .B1(net129));
 sg13g2_nand2b_1 _7147_ (.Y(_2715_),
    .B(_2652_),
    .A_N(_2653_));
 sg13g2_xnor2_1 _7148_ (.Y(_2716_),
    .A(_2715_),
    .B(_2651_));
 sg13g2_o21ai_1 _7149_ (.B1(_2672_),
    .Y(_2717_),
    .A1(_2716_),
    .A2(_2671_));
 sg13g2_a22oi_1 _7150_ (.Y(_2718_),
    .B1(_2677_),
    .B2(_2717_),
    .A2(net89),
    .A1(_2347_));
 sg13g2_a21oi_1 _7151_ (.A1(_2718_),
    .A2(_2674_),
    .Y(_0207_),
    .B1(net129));
 sg13g2_xnor2_1 _7152_ (.Y(_2719_),
    .A(_2684_),
    .B(_2654_));
 sg13g2_o21ai_1 _7153_ (.B1(net69),
    .Y(_2720_),
    .A1(_2719_),
    .A2(net66));
 sg13g2_a22oi_1 _7154_ (.Y(_2721_),
    .B1(_2679_),
    .B2(_2720_),
    .A2(net89),
    .A1(_2345_));
 sg13g2_a21oi_1 _7155_ (.A1(_2721_),
    .A2(_2694_),
    .Y(_0208_),
    .B1(net129));
 sg13g2_xnor2_1 _7156_ (.Y(_2722_),
    .A(_2660_),
    .B(_2657_));
 sg13g2_o21ai_1 _7157_ (.B1(net69),
    .Y(_2723_),
    .A1(_2722_),
    .A2(net66));
 sg13g2_a22oi_1 _7158_ (.Y(_2724_),
    .B1(_2677_),
    .B2(_2723_),
    .A2(net89),
    .A1(_2358_));
 sg13g2_a21oi_1 _7159_ (.A1(_2724_),
    .A2(_2674_),
    .Y(_0209_),
    .B1(net129));
 sg13g2_nand2_1 _7160_ (.Y(_2725_),
    .A(_2685_),
    .B(_2687_));
 sg13g2_xnor2_1 _7161_ (.Y(_2726_),
    .A(_2682_),
    .B(_2725_));
 sg13g2_o21ai_1 _7162_ (.B1(net69),
    .Y(_2727_),
    .A1(_2726_),
    .A2(net66));
 sg13g2_a22oi_1 _7163_ (.Y(_2728_),
    .B1(_2679_),
    .B2(_2727_),
    .A2(net89),
    .A1(_2365_));
 sg13g2_a21oi_1 _7164_ (.A1(_2728_),
    .A2(_2694_),
    .Y(_0210_),
    .B1(net129));
 sg13g2_xnor2_1 _7165_ (.Y(_2729_),
    .A(_2629_),
    .B(_2663_));
 sg13g2_o21ai_1 _7166_ (.B1(net69),
    .Y(_2730_),
    .A1(_2729_),
    .A2(net66));
 sg13g2_a22oi_1 _7167_ (.Y(_2731_),
    .B1(_2677_),
    .B2(_2730_),
    .A2(_2626_),
    .A1(_2318_));
 sg13g2_a21oi_1 _7168_ (.A1(_2731_),
    .A2(_2674_),
    .Y(_0211_),
    .B1(net129));
 sg13g2_nor2b_1 _7169_ (.A(net97),
    .B_N(_0067_),
    .Y(_0264_));
 sg13g2_inv_1 _7170_ (.Y(_2732_),
    .A(_1722_));
 sg13g2_nor3_1 _7171_ (.A(_2732_),
    .B(_2253_),
    .C(net97),
    .Y(_0265_));
 sg13g2_nor2_1 _7172_ (.A(\i_orchestrator.vga_x[2] ),
    .B(_2732_),
    .Y(_2733_));
 sg13g2_nor3_1 _7173_ (.A(_1723_),
    .B(_2733_),
    .C(_1728_),
    .Y(_0266_));
 sg13g2_nor2_1 _7174_ (.A(_3608_),
    .B(_1723_),
    .Y(_2734_));
 sg13g2_nor3_1 _7175_ (.A(net140),
    .B(_2734_),
    .C(_1725_),
    .Y(_0267_));
 sg13g2_buf_1 _7176_ (.A(net168),
    .X(_2735_));
 sg13g2_nor2_1 _7177_ (.A(_3541_),
    .B(_1724_),
    .Y(_2736_));
 sg13g2_nor2_1 _7178_ (.A(_3540_),
    .B(_1725_),
    .Y(_2737_));
 sg13g2_nor3_1 _7179_ (.A(net135),
    .B(_2736_),
    .C(_2737_),
    .Y(_0268_));
 sg13g2_nor2_1 _7180_ (.A(_3538_),
    .B(_2736_),
    .Y(_2738_));
 sg13g2_nor3_1 _7181_ (.A(_3539_),
    .B(_3541_),
    .C(_1724_),
    .Y(_2739_));
 sg13g2_nor3_1 _7182_ (.A(_2738_),
    .B(_2739_),
    .C(_1728_),
    .Y(_0269_));
 sg13g2_nor2_1 _7183_ (.A(_3536_),
    .B(_2739_),
    .Y(_2740_));
 sg13g2_nand2_1 _7184_ (.Y(_2741_),
    .A(_2739_),
    .B(_3536_));
 sg13g2_inv_1 _7185_ (.Y(_2742_),
    .A(_2741_));
 sg13g2_nor3_1 _7186_ (.A(_2740_),
    .B(net97),
    .C(_2742_),
    .Y(_0270_));
 sg13g2_nor2_1 _7187_ (.A(_1719_),
    .B(_2741_),
    .Y(_2743_));
 sg13g2_nor2_1 _7188_ (.A(\i_orchestrator.vga_x[7] ),
    .B(_2742_),
    .Y(_2744_));
 sg13g2_nor3_1 _7189_ (.A(net97),
    .B(_2743_),
    .C(_2744_),
    .Y(_0271_));
 sg13g2_nor2_1 _7190_ (.A(_3534_),
    .B(_2743_),
    .Y(_2745_));
 sg13g2_nand2_1 _7191_ (.Y(_2746_),
    .A(_2743_),
    .B(_3534_));
 sg13g2_inv_1 _7192_ (.Y(_2747_),
    .A(_2746_));
 sg13g2_nor3_1 _7193_ (.A(net97),
    .B(_2745_),
    .C(_2747_),
    .Y(_0272_));
 sg13g2_o21ai_1 _7194_ (.B1(net96),
    .Y(_2748_),
    .A1(_3543_),
    .A2(_2746_));
 sg13g2_a21oi_1 _7195_ (.A1(_3543_),
    .A2(_2746_),
    .Y(_0273_),
    .B1(_2748_));
 sg13g2_buf_1 _7196_ (.A(\i_collision.rotate ),
    .X(_2749_));
 sg13g2_inv_1 _7197_ (.Y(_2750_),
    .A(net170));
 sg13g2_nand2_1 _7198_ (.Y(_2751_),
    .A(net170),
    .B(_1923_));
 sg13g2_inv_1 _7199_ (.Y(_2752_),
    .A(_2751_));
 sg13g2_a21oi_1 _7200_ (.A1(_2750_),
    .A2(_2035_),
    .Y(_2753_),
    .B1(_2752_));
 sg13g2_buf_1 _7201_ (.A(_2753_),
    .X(_2754_));
 sg13g2_nand2b_1 _7202_ (.Y(_2755_),
    .B(_2750_),
    .A_N(_3700_));
 sg13g2_nand2_1 _7203_ (.Y(_2756_),
    .A(net170),
    .B(_3700_));
 sg13g2_nand2_1 _7204_ (.Y(_2757_),
    .A(_2755_),
    .B(_2756_));
 sg13g2_buf_2 _7205_ (.A(_2757_),
    .X(_2758_));
 sg13g2_inv_2 _7206_ (.Y(_2759_),
    .A(_2758_));
 sg13g2_buf_1 _7207_ (.A(_2759_),
    .X(_2760_));
 sg13g2_buf_2 _7208_ (.A(\i_collision.i_coll_table.in[0] ),
    .X(_2761_));
 sg13g2_nor2_1 _7209_ (.A(net157),
    .B(_2761_),
    .Y(_2762_));
 sg13g2_a21oi_1 _7210_ (.A1(_2153_),
    .A2(_2761_),
    .Y(_2763_),
    .B1(_2762_));
 sg13g2_nand2_1 _7211_ (.Y(_2764_),
    .A(net170),
    .B(_0009_));
 sg13g2_o21ai_1 _7212_ (.B1(_2764_),
    .Y(_2765_),
    .A1(net170),
    .A2(_2033_));
 sg13g2_buf_1 _7213_ (.A(_2765_),
    .X(_2766_));
 sg13g2_inv_1 _7214_ (.Y(_2767_),
    .A(net128));
 sg13g2_o21ai_1 _7215_ (.B1(_2767_),
    .Y(_2768_),
    .A1(_2763_),
    .A2(net93));
 sg13g2_a21oi_1 _7216_ (.A1(net93),
    .A2(_2763_),
    .Y(_2769_),
    .B1(_2768_));
 sg13g2_buf_1 _7217_ (.A(_2767_),
    .X(_2770_));
 sg13g2_nand2_2 _7218_ (.Y(_2771_),
    .A(net157),
    .B(_2761_));
 sg13g2_inv_1 _7219_ (.Y(_2772_),
    .A(_2771_));
 sg13g2_buf_1 _7220_ (.A(_2146_),
    .X(_2773_));
 sg13g2_o21ai_1 _7221_ (.B1(net153),
    .Y(_2774_),
    .A1(_2772_),
    .A2(_2758_));
 sg13g2_nor2_1 _7222_ (.A(_2761_),
    .B(_2235_),
    .Y(_2775_));
 sg13g2_inv_1 _7223_ (.Y(_2776_),
    .A(_2775_));
 sg13g2_nor2_1 _7224_ (.A(_2146_),
    .B(_2776_),
    .Y(_2777_));
 sg13g2_nor2_1 _7225_ (.A(_2157_),
    .B(_2777_),
    .Y(_2778_));
 sg13g2_a21oi_1 _7226_ (.A1(_2762_),
    .A2(net158),
    .Y(_2779_),
    .B1(net142));
 sg13g2_inv_2 _7227_ (.Y(_2780_),
    .A(_2761_));
 sg13g2_nor2_1 _7228_ (.A(net157),
    .B(_2780_),
    .Y(_2781_));
 sg13g2_nor2_1 _7229_ (.A(_2781_),
    .B(_2759_),
    .Y(_2782_));
 sg13g2_inv_1 _7230_ (.Y(_2783_),
    .A(_2782_));
 sg13g2_nand2_1 _7231_ (.Y(_2784_),
    .A(_2783_),
    .B(net153));
 sg13g2_a22oi_1 _7232_ (.Y(_2785_),
    .B1(_2779_),
    .B2(_2784_),
    .A2(_2778_),
    .A1(_2774_));
 sg13g2_nor2_1 _7233_ (.A(net107),
    .B(_2785_),
    .Y(_2786_));
 sg13g2_nor2_1 _7234_ (.A(_2769_),
    .B(_2786_),
    .Y(_2787_));
 sg13g2_nor2_1 _7235_ (.A(net119),
    .B(_2787_),
    .Y(_2788_));
 sg13g2_buf_1 _7236_ (.A(net128),
    .X(_2789_));
 sg13g2_nor2_1 _7237_ (.A(_2159_),
    .B(net93),
    .Y(_2790_));
 sg13g2_buf_1 _7238_ (.A(_2147_),
    .X(_2791_));
 sg13g2_nand2_1 _7239_ (.Y(_2792_),
    .A(_2759_),
    .B(_2146_));
 sg13g2_nor2_1 _7240_ (.A(net152),
    .B(_2792_),
    .Y(_2793_));
 sg13g2_a21oi_1 _7241_ (.A1(_2790_),
    .A2(_2772_),
    .Y(_2794_),
    .B1(_2793_));
 sg13g2_inv_1 _7242_ (.Y(_2795_),
    .A(_2781_));
 sg13g2_buf_1 _7243_ (.A(_2758_),
    .X(_2796_));
 sg13g2_nor3_1 _7244_ (.A(_2159_),
    .B(_2795_),
    .C(net106),
    .Y(_2797_));
 sg13g2_nor3_1 _7245_ (.A(net152),
    .B(_0052_),
    .C(net93),
    .Y(_2798_));
 sg13g2_o21ai_1 _7246_ (.B1(net131),
    .Y(_2799_),
    .A1(_2797_),
    .A2(_2798_));
 sg13g2_o21ai_1 _7247_ (.B1(_2799_),
    .Y(_2800_),
    .A1(net131),
    .A2(_2794_));
 sg13g2_a21oi_1 _7248_ (.A1(_2759_),
    .A2(_2771_),
    .Y(_2801_),
    .B1(_2146_));
 sg13g2_nor2_1 _7249_ (.A(_2762_),
    .B(_2759_),
    .Y(_2802_));
 sg13g2_nor2_1 _7250_ (.A(_2802_),
    .B(_2774_),
    .Y(_2803_));
 sg13g2_nor4_1 _7251_ (.A(net152),
    .B(net121),
    .C(_2801_),
    .D(_2803_),
    .Y(_2804_));
 sg13g2_nor2_1 _7252_ (.A(net153),
    .B(_2782_),
    .Y(_2805_));
 sg13g2_nor2_1 _7253_ (.A(_2775_),
    .B(_2758_),
    .Y(_2806_));
 sg13g2_nor2_1 _7254_ (.A(_2806_),
    .B(_2784_),
    .Y(_2807_));
 sg13g2_nor4_1 _7255_ (.A(net152),
    .B(net142),
    .C(_2805_),
    .D(_2807_),
    .Y(_2808_));
 sg13g2_nor2_1 _7256_ (.A(_2804_),
    .B(_2808_),
    .Y(_2809_));
 sg13g2_nor2_1 _7257_ (.A(_2153_),
    .B(_2806_),
    .Y(_2810_));
 sg13g2_nor2_1 _7258_ (.A(net128),
    .B(_2810_),
    .Y(_2811_));
 sg13g2_o21ai_1 _7259_ (.B1(_2811_),
    .Y(_2812_),
    .A1(_2157_),
    .A2(_2802_));
 sg13g2_o21ai_1 _7260_ (.B1(_2812_),
    .Y(_2813_),
    .A1(net152),
    .A2(net128));
 sg13g2_inv_1 _7261_ (.Y(_2814_),
    .A(_2753_));
 sg13g2_a221oi_1 _7262_ (.B2(_2813_),
    .C1(net117),
    .B1(_2809_),
    .A1(net118),
    .Y(_2815_),
    .A2(_2800_));
 sg13g2_inv_1 _7263_ (.Y(_2816_),
    .A(\i_collision.mirror ));
 sg13g2_nand2_1 _7264_ (.Y(_2817_),
    .A(net170),
    .B(net178));
 sg13g2_o21ai_1 _7265_ (.B1(_2817_),
    .Y(_2818_),
    .A1(net170),
    .A2(_2055_));
 sg13g2_xnor2_1 _7266_ (.Y(_2819_),
    .A(_2816_),
    .B(_2818_));
 sg13g2_buf_2 _7267_ (.A(_2819_),
    .X(_2820_));
 sg13g2_inv_1 _7268_ (.Y(_2821_),
    .A(_2820_));
 sg13g2_o21ai_1 _7269_ (.B1(_2821_),
    .Y(_2822_),
    .A1(_2788_),
    .A2(_2815_));
 sg13g2_buf_2 _7270_ (.A(\i_collision.update ),
    .X(_2823_));
 sg13g2_nor2_1 _7271_ (.A(_2771_),
    .B(_2758_),
    .Y(_2824_));
 sg13g2_nor2_1 _7272_ (.A(_2776_),
    .B(_2758_),
    .Y(_2825_));
 sg13g2_inv_1 _7273_ (.Y(_2826_),
    .A(_2825_));
 sg13g2_nand2_1 _7274_ (.Y(_2827_),
    .A(_2826_),
    .B(_2165_));
 sg13g2_o21ai_1 _7275_ (.B1(_2827_),
    .Y(_2828_),
    .A1(_2148_),
    .A2(_2824_));
 sg13g2_a21o_1 _7276_ (.A2(_2824_),
    .A1(_2160_),
    .B1(_2828_),
    .X(_2829_));
 sg13g2_nor2_1 _7277_ (.A(_2795_),
    .B(_2759_),
    .Y(_2830_));
 sg13g2_inv_1 _7278_ (.Y(_2831_),
    .A(_2830_));
 sg13g2_inv_1 _7279_ (.Y(_2832_),
    .A(_2762_));
 sg13g2_nor2_1 _7280_ (.A(_2832_),
    .B(_2759_),
    .Y(_2833_));
 sg13g2_inv_1 _7281_ (.Y(_2834_),
    .A(_2833_));
 sg13g2_a22oi_1 _7282_ (.Y(_2835_),
    .B1(_2165_),
    .B2(_2834_),
    .A2(_2150_),
    .A1(_2831_));
 sg13g2_nand2_1 _7283_ (.Y(_2836_),
    .A(_2830_),
    .B(_2160_));
 sg13g2_a21oi_1 _7284_ (.A1(_2835_),
    .A2(_2836_),
    .Y(_2837_),
    .B1(net142));
 sg13g2_a21oi_1 _7285_ (.A1(_2829_),
    .A2(net131),
    .Y(_2838_),
    .B1(_2837_));
 sg13g2_nand2_1 _7286_ (.Y(_2839_),
    .A(_2838_),
    .B(net118));
 sg13g2_o21ai_1 _7287_ (.B1(_2767_),
    .Y(_2840_),
    .A1(_2780_),
    .A2(_2165_));
 sg13g2_a21o_1 _7288_ (.A2(_2165_),
    .A1(_2780_),
    .B1(_2840_),
    .X(_2841_));
 sg13g2_nand3_1 _7289_ (.B(net119),
    .C(_2841_),
    .A(_2839_),
    .Y(_2842_));
 sg13g2_nand2_1 _7290_ (.Y(_2843_),
    .A(_2773_),
    .B(_2761_));
 sg13g2_inv_1 _7291_ (.Y(_2844_),
    .A(_2843_));
 sg13g2_nand3_1 _7292_ (.B(net118),
    .C(_2844_),
    .A(net117),
    .Y(_2845_));
 sg13g2_nand3_1 _7293_ (.B(_2820_),
    .C(_2845_),
    .A(_2842_),
    .Y(_2846_));
 sg13g2_nor2_2 _7294_ (.A(_2157_),
    .B(_2796_),
    .Y(_2847_));
 sg13g2_a21oi_1 _7295_ (.A1(_0068_),
    .A2(net106),
    .Y(_2848_),
    .B1(_2847_));
 sg13g2_buf_1 _7296_ (.A(_0053_),
    .X(_2849_));
 sg13g2_inv_1 _7297_ (.Y(_2850_),
    .A(_2849_));
 sg13g2_nor2_2 _7298_ (.A(_2767_),
    .B(net117),
    .Y(_2851_));
 sg13g2_nand4_1 _7299_ (.B(_2848_),
    .C(_2850_),
    .A(_2821_),
    .Y(_2852_),
    .D(_2851_));
 sg13g2_nand4_1 _7300_ (.B(_2823_),
    .C(_2846_),
    .A(_2822_),
    .Y(_2853_),
    .D(_2852_));
 sg13g2_a21o_1 _7301_ (.A2(_2823_),
    .A1(_2852_),
    .B1(net158),
    .X(_2854_));
 sg13g2_a21oi_1 _7302_ (.A1(_2853_),
    .A2(_2854_),
    .Y(_0069_),
    .B1(net140));
 sg13g2_nor2_1 _7303_ (.A(_2235_),
    .B(net106),
    .Y(_2855_));
 sg13g2_inv_1 _7304_ (.Y(_2856_),
    .A(_2855_));
 sg13g2_nand2b_1 _7305_ (.Y(_2857_),
    .B(_2856_),
    .A_N(_2227_));
 sg13g2_inv_1 _7306_ (.Y(_2858_),
    .A(_2175_));
 sg13g2_nor2_2 _7307_ (.A(_2154_),
    .B(_2758_),
    .Y(_2859_));
 sg13g2_inv_1 _7308_ (.Y(_2860_),
    .A(_2859_));
 sg13g2_nand4_1 _7309_ (.B(_2851_),
    .C(_2858_),
    .A(_2857_),
    .Y(_2861_),
    .D(_2860_));
 sg13g2_o21ai_1 _7310_ (.B1(net128),
    .Y(_2862_),
    .A1(_2227_),
    .A2(_2796_));
 sg13g2_a21o_1 _7311_ (.A2(net106),
    .A1(_2228_),
    .B1(_2862_),
    .X(_2863_));
 sg13g2_nor2_1 _7312_ (.A(net157),
    .B(_2759_),
    .Y(_2864_));
 sg13g2_inv_1 _7313_ (.Y(_2865_),
    .A(_2864_));
 sg13g2_a21oi_2 _7314_ (.B1(_2227_),
    .Y(_2866_),
    .A2(_2860_),
    .A1(_2865_));
 sg13g2_a21oi_1 _7315_ (.A1(_2866_),
    .A2(net107),
    .Y(_2867_),
    .B1(net119));
 sg13g2_inv_1 _7316_ (.Y(_2868_),
    .A(_2866_));
 sg13g2_nor2_1 _7317_ (.A(_2858_),
    .B(_2766_),
    .Y(_2869_));
 sg13g2_a21oi_1 _7318_ (.A1(_2868_),
    .A2(_2869_),
    .Y(_2870_),
    .B1(net117));
 sg13g2_nor3_1 _7319_ (.A(_2235_),
    .B(net152),
    .C(net93),
    .Y(_2871_));
 sg13g2_buf_1 _7320_ (.A(_0051_),
    .X(_2872_));
 sg13g2_a22oi_1 _7321_ (.Y(_2873_),
    .B1(_2872_),
    .B2(_2859_),
    .A2(_2175_),
    .A1(net121));
 sg13g2_o21ai_1 _7322_ (.B1(_2858_),
    .Y(_2874_),
    .A1(_2872_),
    .A2(net93));
 sg13g2_a21oi_1 _7323_ (.A1(_2760_),
    .A2(_2235_),
    .Y(_2875_),
    .B1(net121));
 sg13g2_a21oi_1 _7324_ (.A1(_2874_),
    .A2(_2875_),
    .Y(_2876_),
    .B1(net107));
 sg13g2_o21ai_1 _7325_ (.B1(_2876_),
    .Y(_2877_),
    .A1(_2871_),
    .A2(_2873_));
 sg13g2_a22oi_1 _7326_ (.Y(_2878_),
    .B1(_2870_),
    .B2(_2877_),
    .A2(_2867_),
    .A1(_2863_));
 sg13g2_mux2_1 _7327_ (.A0(_2861_),
    .A1(_2878_),
    .S(_2821_),
    .X(_2879_));
 sg13g2_buf_1 _7328_ (.A(net183),
    .X(_2880_));
 sg13g2_o21ai_1 _7329_ (.B1(net151),
    .Y(_2881_),
    .A1(_2823_),
    .A2(\collision_impact[0] ));
 sg13g2_a21oi_1 _7330_ (.A1(_2879_),
    .A2(_2823_),
    .Y(_0076_),
    .B1(_2881_));
 sg13g2_nor2_1 _7331_ (.A(_2157_),
    .B(net93),
    .Y(_2882_));
 sg13g2_nor2_1 _7332_ (.A(_2859_),
    .B(_2882_),
    .Y(_2883_));
 sg13g2_nor2_1 _7333_ (.A(_2175_),
    .B(_2883_),
    .Y(_2884_));
 sg13g2_nand2b_1 _7334_ (.Y(_2885_),
    .B(_2868_),
    .A_N(_2884_));
 sg13g2_a21o_1 _7335_ (.A2(_2872_),
    .A1(_2175_),
    .B1(net131),
    .X(_2886_));
 sg13g2_o21ai_1 _7336_ (.B1(_2847_),
    .Y(_2887_),
    .A1(_2872_),
    .A2(_2858_));
 sg13g2_o21ai_1 _7337_ (.B1(_2887_),
    .Y(_2888_),
    .A1(net93),
    .A2(_2886_));
 sg13g2_a21oi_1 _7338_ (.A1(_2888_),
    .A2(_2789_),
    .Y(_2889_),
    .B1(_2814_));
 sg13g2_o21ai_1 _7339_ (.B1(_2889_),
    .Y(_2890_),
    .A1(net118),
    .A2(_2885_));
 sg13g2_nand3_1 _7340_ (.B(_2789_),
    .C(_2814_),
    .A(_2866_),
    .Y(_2891_));
 sg13g2_inv_2 _7341_ (.Y(_2892_),
    .A(_2823_));
 sg13g2_nor2_1 _7342_ (.A(_2892_),
    .B(_2820_),
    .Y(_2893_));
 sg13g2_nand3_1 _7343_ (.B(_2891_),
    .C(_2893_),
    .A(_2890_),
    .Y(_2894_));
 sg13g2_nand2_1 _7344_ (.Y(_2895_),
    .A(_2892_),
    .B(\collision_impact[1] ));
 sg13g2_a21oi_1 _7345_ (.A1(_2894_),
    .A2(_2895_),
    .Y(_0077_),
    .B1(net140));
 sg13g2_nand2_1 _7346_ (.Y(_2896_),
    .A(_2749_),
    .B(_2823_));
 sg13g2_inv_1 _7347_ (.Y(_2897_),
    .A(_2896_));
 sg13g2_o21ai_1 _7348_ (.B1(net151),
    .Y(_2898_),
    .A1(_1922_),
    .A2(_2897_));
 sg13g2_nand3_1 _7349_ (.B(net158),
    .C(_2772_),
    .A(net106),
    .Y(_2899_));
 sg13g2_nand3_1 _7350_ (.B(net153),
    .C(_2771_),
    .A(net106),
    .Y(_2900_));
 sg13g2_a21oi_1 _7351_ (.A1(_2899_),
    .A2(_2900_),
    .Y(_2901_),
    .B1(_2159_));
 sg13g2_o21ai_1 _7352_ (.B1(net121),
    .Y(_2902_),
    .A1(_2798_),
    .A2(_2901_));
 sg13g2_o21ai_1 _7353_ (.B1(net158),
    .Y(_2903_),
    .A1(_2159_),
    .A2(_2795_));
 sg13g2_nand3_1 _7354_ (.B(net153),
    .C(_2791_),
    .A(_2781_),
    .Y(_2904_));
 sg13g2_nand3_1 _7355_ (.B(_2847_),
    .C(_2904_),
    .A(_2903_),
    .Y(_2905_));
 sg13g2_nand3_1 _7356_ (.B(net128),
    .C(_2905_),
    .A(_2902_),
    .Y(_2906_));
 sg13g2_nor2_1 _7357_ (.A(_2772_),
    .B(_2792_),
    .Y(_2907_));
 sg13g2_nor4_1 _7358_ (.A(_2157_),
    .B(_2802_),
    .C(_2801_),
    .D(_2907_),
    .Y(_2908_));
 sg13g2_nor2_1 _7359_ (.A(net158),
    .B(_2783_),
    .Y(_2909_));
 sg13g2_nor4_1 _7360_ (.A(net142),
    .B(_2806_),
    .C(_2805_),
    .D(_2909_),
    .Y(_2910_));
 sg13g2_nor2_1 _7361_ (.A(_2908_),
    .B(_2910_),
    .Y(_2911_));
 sg13g2_nand2_1 _7362_ (.Y(_2912_),
    .A(_2911_),
    .B(_2813_));
 sg13g2_a21oi_1 _7363_ (.A1(_2906_),
    .A2(_2912_),
    .Y(_2913_),
    .B1(net117));
 sg13g2_o21ai_1 _7364_ (.B1(_2779_),
    .Y(_2914_),
    .A1(net158),
    .A2(_2783_));
 sg13g2_o21ai_1 _7365_ (.B1(_2778_),
    .Y(_2915_),
    .A1(_2772_),
    .A2(_2792_));
 sg13g2_nand3_1 _7366_ (.B(net128),
    .C(_2915_),
    .A(_2914_),
    .Y(_2916_));
 sg13g2_nor2_1 _7367_ (.A(net119),
    .B(_2769_),
    .Y(_2917_));
 sg13g2_a21o_1 _7368_ (.A2(_2917_),
    .A1(_2916_),
    .B1(_2820_),
    .X(_2918_));
 sg13g2_a221oi_1 _7369_ (.B2(_2833_),
    .C1(_2154_),
    .B1(_2165_),
    .A1(_2830_),
    .Y(_2919_),
    .A2(net152));
 sg13g2_a221oi_1 _7370_ (.B2(_2775_),
    .C1(_2157_),
    .B1(_2793_),
    .A1(_2791_),
    .Y(_2920_),
    .A2(_2824_));
 sg13g2_nor3_1 _7371_ (.A(_2767_),
    .B(_2919_),
    .C(_2920_),
    .Y(_2921_));
 sg13g2_a21oi_1 _7372_ (.A1(_0054_),
    .A2(net107),
    .Y(_2922_),
    .B1(_2921_));
 sg13g2_nand2_1 _7373_ (.Y(_2923_),
    .A(_2922_),
    .B(net119));
 sg13g2_nand2_1 _7374_ (.Y(_2924_),
    .A(_2780_),
    .B(net153));
 sg13g2_nand3_1 _7375_ (.B(net118),
    .C(_2924_),
    .A(net117),
    .Y(_2925_));
 sg13g2_nand3_1 _7376_ (.B(_2820_),
    .C(_2925_),
    .A(_2923_),
    .Y(_2926_));
 sg13g2_o21ai_1 _7377_ (.B1(_2926_),
    .Y(_2927_),
    .A1(_2913_),
    .A2(_2918_));
 sg13g2_nor2_1 _7378_ (.A(_2896_),
    .B(_2927_),
    .Y(_2928_));
 sg13g2_nor2_1 _7379_ (.A(_2898_),
    .B(_2928_),
    .Y(_0078_));
 sg13g2_nor2_1 _7380_ (.A(_2849_),
    .B(_2197_),
    .Y(_2929_));
 sg13g2_nor2_1 _7381_ (.A(net142),
    .B(_2849_),
    .Y(_2930_));
 sg13g2_a22oi_1 _7382_ (.Y(_2931_),
    .B1(_2930_),
    .B2(_2833_),
    .A2(_2929_),
    .A1(_2825_));
 sg13g2_o21ai_1 _7383_ (.B1(net119),
    .Y(_2932_),
    .A1(net107),
    .A2(_2931_));
 sg13g2_nor4_1 _7384_ (.A(_2773_),
    .B(_2780_),
    .C(_2227_),
    .D(_2229_),
    .Y(_2933_));
 sg13g2_o21ai_1 _7385_ (.B1(net118),
    .Y(_2934_),
    .A1(_2849_),
    .A2(_2933_));
 sg13g2_inv_1 _7386_ (.Y(_2935_),
    .A(_0052_));
 sg13g2_o21ai_1 _7387_ (.B1(_2935_),
    .Y(_2936_),
    .A1(_2780_),
    .A2(_2230_));
 sg13g2_nand3_1 _7388_ (.B(_2159_),
    .C(net107),
    .A(_2936_),
    .Y(_2937_));
 sg13g2_nand4_1 _7389_ (.B(_2937_),
    .C(_2754_),
    .A(_2934_),
    .Y(_2938_),
    .D(_2883_));
 sg13g2_a22oi_1 _7390_ (.Y(_2939_),
    .B1(net121),
    .B2(_2782_),
    .A2(_2771_),
    .A1(_2847_));
 sg13g2_a21oi_1 _7391_ (.A1(_2939_),
    .A2(net107),
    .Y(_2940_),
    .B1(net119));
 sg13g2_a21oi_1 _7392_ (.A1(_2872_),
    .A2(net158),
    .Y(_2941_),
    .B1(_2760_));
 sg13g2_nand2_1 _7393_ (.Y(_2942_),
    .A(_2941_),
    .B(_2197_));
 sg13g2_o21ai_1 _7394_ (.B1(_2847_),
    .Y(_2943_),
    .A1(_2872_),
    .A2(net153));
 sg13g2_nand3_1 _7395_ (.B(_2943_),
    .C(net128),
    .A(_2942_),
    .Y(_2944_));
 sg13g2_nand2_1 _7396_ (.Y(_2945_),
    .A(_2940_),
    .B(_2944_));
 sg13g2_nand3_1 _7397_ (.B(_2945_),
    .C(_2821_),
    .A(_2938_),
    .Y(_2946_));
 sg13g2_o21ai_1 _7398_ (.B1(_2946_),
    .Y(_2947_),
    .A1(_2821_),
    .A2(_2932_));
 sg13g2_a21oi_1 _7399_ (.A1(_2896_),
    .A2(_1923_),
    .Y(_2948_),
    .B1(net141));
 sg13g2_o21ai_1 _7400_ (.B1(_2948_),
    .Y(_0079_),
    .A1(_2896_),
    .A2(_2947_));
 sg13g2_a21oi_1 _7401_ (.A1(_2884_),
    .A2(_2851_),
    .Y(_2949_),
    .B1(_2866_));
 sg13g2_nor2b_1 _7402_ (.A(_2949_),
    .B_N(_2818_),
    .Y(_2950_));
 sg13g2_a21oi_1 _7403_ (.A1(_2816_),
    .A2(_2949_),
    .Y(_2951_),
    .B1(_2950_));
 sg13g2_buf_1 _7404_ (.A(net183),
    .X(_2952_));
 sg13g2_o21ai_1 _7405_ (.B1(net150),
    .Y(_2953_),
    .A1(_1975_),
    .A2(_2897_));
 sg13g2_a21oi_1 _7406_ (.A1(_2951_),
    .A2(_2897_),
    .Y(_0080_),
    .B1(_2953_));
 sg13g2_nor2_2 _7407_ (.A(net170),
    .B(_2892_),
    .Y(_2954_));
 sg13g2_a21oi_1 _7408_ (.A1(_2927_),
    .A2(_2954_),
    .Y(_2955_),
    .B1(net141));
 sg13g2_o21ai_1 _7409_ (.B1(_2955_),
    .Y(_0081_),
    .A1(_2054_),
    .A2(_2954_));
 sg13g2_o21ai_1 _7410_ (.B1(net150),
    .Y(_2956_),
    .A1(_2035_),
    .A2(_2954_));
 sg13g2_a21oi_1 _7411_ (.A1(_2947_),
    .A2(_2954_),
    .Y(_0082_),
    .B1(_2956_));
 sg13g2_o21ai_1 _7412_ (.B1(net150),
    .Y(_2957_),
    .A1(_2097_),
    .A2(_2954_));
 sg13g2_a21oi_1 _7413_ (.A1(_2951_),
    .A2(_2954_),
    .Y(_0083_),
    .B1(_2957_));
 sg13g2_a21oi_1 _7414_ (.A1(_2802_),
    .A2(_2935_),
    .Y(_2958_),
    .B1(_2790_));
 sg13g2_nor2_1 _7415_ (.A(net121),
    .B(_2958_),
    .Y(_2959_));
 sg13g2_o21ai_1 _7416_ (.B1(_2811_),
    .Y(_2960_),
    .A1(_2161_),
    .A2(_2959_));
 sg13g2_nand2_1 _7417_ (.Y(_2961_),
    .A(_2859_),
    .B(net152));
 sg13g2_nand3_1 _7418_ (.B(_2850_),
    .C(net118),
    .A(_2882_),
    .Y(_2962_));
 sg13g2_nand3_1 _7419_ (.B(_2961_),
    .C(_2962_),
    .A(_2960_),
    .Y(_2963_));
 sg13g2_nand3b_1 _7420_ (.B(_2875_),
    .C(_2792_),
    .Y(_2964_),
    .A_N(_2777_));
 sg13g2_o21ai_1 _7421_ (.B1(net106),
    .Y(_2965_),
    .A1(net157),
    .A2(net153));
 sg13g2_nand2_1 _7422_ (.Y(_2966_),
    .A(_2965_),
    .B(_2779_));
 sg13g2_a21o_1 _7423_ (.A2(_2966_),
    .A1(_2964_),
    .B1(net107),
    .X(_2967_));
 sg13g2_a21oi_1 _7424_ (.A1(_2967_),
    .A2(_2940_),
    .Y(_2968_),
    .B1(_2820_));
 sg13g2_o21ai_1 _7425_ (.B1(_2968_),
    .Y(_2969_),
    .A1(net117),
    .A2(_2963_));
 sg13g2_o21ai_1 _7426_ (.B1(_2930_),
    .Y(_2970_),
    .A1(_2844_),
    .A2(_2865_));
 sg13g2_o21ai_1 _7427_ (.B1(_2929_),
    .Y(_2971_),
    .A1(_2844_),
    .A2(_2856_));
 sg13g2_nand3_1 _7428_ (.B(net118),
    .C(_2971_),
    .A(_2970_),
    .Y(_2972_));
 sg13g2_nand3_1 _7429_ (.B(_2849_),
    .C(_2843_),
    .A(_2770_),
    .Y(_2973_));
 sg13g2_nand4_1 _7430_ (.B(net119),
    .C(_2820_),
    .A(_2972_),
    .Y(_2974_),
    .D(_2973_));
 sg13g2_nor2b_1 _7431_ (.A(_2892_),
    .B_N(_2974_),
    .Y(_2975_));
 sg13g2_a221oi_1 _7432_ (.B2(_2975_),
    .C1(net140),
    .B1(_2969_),
    .A1(_2892_),
    .Y(_0084_),
    .A2(_2159_));
 sg13g2_o21ai_1 _7433_ (.B1(net117),
    .Y(_2976_),
    .A1(_2164_),
    .A2(_2770_));
 sg13g2_nand3b_1 _7434_ (.B(_2976_),
    .C(_2865_),
    .Y(_2977_),
    .A_N(_2869_));
 sg13g2_a21oi_1 _7435_ (.A1(_2977_),
    .A2(_2893_),
    .Y(_2978_),
    .B1(net131));
 sg13g2_a21oi_1 _7436_ (.A1(_2864_),
    .A2(_2754_),
    .Y(_2979_),
    .B1(_2851_));
 sg13g2_nand3_1 _7437_ (.B(_2235_),
    .C(_2858_),
    .A(_2976_),
    .Y(_2980_));
 sg13g2_a22oi_1 _7438_ (.Y(_2981_),
    .B1(_2979_),
    .B2(_2980_),
    .A2(_2851_),
    .A1(_2229_));
 sg13g2_nor4_1 _7439_ (.A(_2892_),
    .B(net106),
    .C(_2820_),
    .D(_2981_),
    .Y(_2982_));
 sg13g2_nor3_1 _7440_ (.A(net135),
    .B(_2978_),
    .C(_2982_),
    .Y(_0085_));
 sg13g2_inv_1 _7441_ (.Y(_2983_),
    .A(_3491_));
 sg13g2_nor3_1 _7442_ (.A(_3485_),
    .B(_3488_),
    .C(_3490_),
    .Y(_2984_));
 sg13g2_o21ai_1 _7443_ (.B1(_2984_),
    .Y(_2985_),
    .A1(_2983_),
    .A2(_1892_));
 sg13g2_nand2b_1 _7444_ (.Y(_2986_),
    .B(_1888_),
    .A_N(_2984_));
 sg13g2_nand3_1 _7445_ (.B(_2986_),
    .C(net151),
    .A(_2985_),
    .Y(_0086_));
 sg13g2_nand2_1 _7446_ (.Y(_2987_),
    .A(_1888_),
    .B(_0011_));
 sg13g2_inv_1 _7447_ (.Y(_2988_),
    .A(_2987_));
 sg13g2_a21oi_1 _7448_ (.A1(_2984_),
    .A2(_2988_),
    .Y(_2989_),
    .B1(\capsule_color[1] ));
 sg13g2_inv_1 _7449_ (.Y(_2990_),
    .A(_1893_));
 sg13g2_nand3_1 _7450_ (.B(_2990_),
    .C(_1911_),
    .A(_1904_),
    .Y(_2991_));
 sg13g2_buf_1 _7451_ (.A(\color_entropy[0] ),
    .X(_2992_));
 sg13g2_a21oi_1 _7452_ (.A1(_2991_),
    .A2(_2992_),
    .Y(_2993_),
    .B1(_2983_));
 sg13g2_nor2_1 _7453_ (.A(_2993_),
    .B(_2985_),
    .Y(_2994_));
 sg13g2_nor3_1 _7454_ (.A(net135),
    .B(_2989_),
    .C(_2994_),
    .Y(_0087_));
 sg13g2_nand3b_1 _7455_ (.B(_3480_),
    .C(_2983_),
    .Y(_2995_),
    .A_N(_3488_));
 sg13g2_buf_1 _7456_ (.A(_2995_),
    .X(_2996_));
 sg13g2_a21oi_1 _7457_ (.A1(_3485_),
    .A2(_1893_),
    .Y(_2997_),
    .B1(_2996_));
 sg13g2_a21oi_1 _7458_ (.A1(_1893_),
    .A2(_2996_),
    .Y(_2998_),
    .B1(_2997_));
 sg13g2_nand2_1 _7459_ (.Y(_0088_),
    .A(_2998_),
    .B(net151));
 sg13g2_o21ai_1 _7460_ (.B1(_1911_),
    .Y(_2999_),
    .A1(_1893_),
    .A2(_1891_));
 sg13g2_nand3_1 _7461_ (.B(_2992_),
    .C(_1894_),
    .A(_2999_),
    .Y(_3000_));
 sg13g2_a21oi_1 _7462_ (.A1(_3000_),
    .A2(_3485_),
    .Y(_3001_),
    .B1(_2996_));
 sg13g2_o21ai_1 _7463_ (.B1(_1904_),
    .Y(_3002_),
    .A1(_2990_),
    .A2(_2996_));
 sg13g2_nand2_1 _7464_ (.Y(_3003_),
    .A(_3002_),
    .B(net151));
 sg13g2_nor2_1 _7465_ (.A(_3001_),
    .B(_3003_),
    .Y(_0089_));
 sg13g2_nor3_1 _7466_ (.A(_3491_),
    .B(_3485_),
    .C(_3490_),
    .Y(_3004_));
 sg13g2_inv_1 _7467_ (.Y(_3005_),
    .A(_3004_));
 sg13g2_o21ai_1 _7468_ (.B1(_1910_),
    .Y(_3006_),
    .A1(_0010_),
    .A2(_3005_));
 sg13g2_nand2_1 _7469_ (.Y(_3007_),
    .A(_3004_),
    .B(_1912_));
 sg13g2_nand3_1 _7470_ (.B(net151),
    .C(_3007_),
    .A(_3006_),
    .Y(_0090_));
 sg13g2_o21ai_1 _7471_ (.B1(_1904_),
    .Y(_3008_),
    .A1(_2990_),
    .A2(_1891_));
 sg13g2_nand2_1 _7472_ (.Y(_3009_),
    .A(_3008_),
    .B(_2992_));
 sg13g2_o21ai_1 _7473_ (.B1(\capsule_color[5] ),
    .Y(_3010_),
    .A1(_3009_),
    .A2(_3007_));
 sg13g2_a21oi_1 _7474_ (.A1(_1910_),
    .A2(_0011_),
    .Y(_3011_),
    .B1(_0010_));
 sg13g2_nand2b_1 _7475_ (.Y(_3012_),
    .B(_3004_),
    .A_N(_3011_));
 sg13g2_nand3_1 _7476_ (.B(net151),
    .C(_3012_),
    .A(_3010_),
    .Y(_0091_));
 sg13g2_nor2_1 _7477_ (.A(\i_delta_sigma.acc[0] ),
    .B(_2623_),
    .Y(_3013_));
 sg13g2_nand2_1 _7478_ (.Y(_3014_),
    .A(\i_delta_sigma.acc[0] ),
    .B(_2623_));
 sg13g2_inv_1 _7479_ (.Y(_3015_),
    .A(_3014_));
 sg13g2_nor3_1 _7480_ (.A(net135),
    .B(_3013_),
    .C(_3015_),
    .Y(_0092_));
 sg13g2_nor2_1 _7481_ (.A(\i_delta_sigma.acc[10] ),
    .B(_2316_),
    .Y(_3016_));
 sg13g2_nand2_1 _7482_ (.Y(_3017_),
    .A(\i_delta_sigma.acc[10] ),
    .B(_2316_));
 sg13g2_inv_1 _7483_ (.Y(_3018_),
    .A(_3017_));
 sg13g2_nor2_1 _7484_ (.A(_3016_),
    .B(_3018_),
    .Y(_3019_));
 sg13g2_inv_1 _7485_ (.Y(_3020_),
    .A(_3019_));
 sg13g2_nor2_1 _7486_ (.A(\i_delta_sigma.acc[5] ),
    .B(_2347_),
    .Y(_3021_));
 sg13g2_nor2_1 _7487_ (.A(\i_delta_sigma.acc[4] ),
    .B(_2329_),
    .Y(_3022_));
 sg13g2_xor2_1 _7488_ (.B(_2632_),
    .A(\i_delta_sigma.acc[1] ),
    .X(_3023_));
 sg13g2_nand2_1 _7489_ (.Y(_3024_),
    .A(_3023_),
    .B(_3015_));
 sg13g2_inv_1 _7490_ (.Y(_3025_),
    .A(_3024_));
 sg13g2_a21oi_1 _7491_ (.A1(\i_delta_sigma.acc[1] ),
    .A2(_2632_),
    .Y(_3026_),
    .B1(_3025_));
 sg13g2_inv_1 _7492_ (.Y(_3027_),
    .A(_3026_));
 sg13g2_xor2_1 _7493_ (.B(_2637_),
    .A(\i_delta_sigma.acc[2] ),
    .X(_3028_));
 sg13g2_nand2_1 _7494_ (.Y(_3029_),
    .A(_3027_),
    .B(_3028_));
 sg13g2_inv_1 _7495_ (.Y(_3030_),
    .A(_3029_));
 sg13g2_a21oi_1 _7496_ (.A1(\i_delta_sigma.acc[2] ),
    .A2(_2637_),
    .Y(_3031_),
    .B1(_3030_));
 sg13g2_nand2_1 _7497_ (.Y(_3032_),
    .A(\i_delta_sigma.acc[3] ),
    .B(_2643_));
 sg13g2_nor2_1 _7498_ (.A(\i_delta_sigma.acc[3] ),
    .B(_2643_),
    .Y(_3033_));
 sg13g2_a21oi_1 _7499_ (.A1(_3031_),
    .A2(_3032_),
    .Y(_3034_),
    .B1(_3033_));
 sg13g2_inv_1 _7500_ (.Y(_3035_),
    .A(_3034_));
 sg13g2_nand2_1 _7501_ (.Y(_3036_),
    .A(\i_delta_sigma.acc[4] ),
    .B(_2329_));
 sg13g2_o21ai_1 _7502_ (.B1(_3036_),
    .Y(_3037_),
    .A1(_3022_),
    .A2(_3035_));
 sg13g2_inv_1 _7503_ (.Y(_3038_),
    .A(_3037_));
 sg13g2_nand2_1 _7504_ (.Y(_3039_),
    .A(\i_delta_sigma.acc[5] ),
    .B(_2347_));
 sg13g2_o21ai_1 _7505_ (.B1(_3039_),
    .Y(_3040_),
    .A1(_3021_),
    .A2(_3038_));
 sg13g2_buf_1 _7506_ (.A(_3040_),
    .X(_3041_));
 sg13g2_nor2_1 _7507_ (.A(\i_delta_sigma.acc[7] ),
    .B(_2358_),
    .Y(_3042_));
 sg13g2_nand2_1 _7508_ (.Y(_3043_),
    .A(\i_delta_sigma.acc[7] ),
    .B(_2358_));
 sg13g2_inv_1 _7509_ (.Y(_3044_),
    .A(_3043_));
 sg13g2_nor2_1 _7510_ (.A(_3042_),
    .B(_3044_),
    .Y(_3045_));
 sg13g2_inv_1 _7511_ (.Y(_3046_),
    .A(_3045_));
 sg13g2_nor2_1 _7512_ (.A(\i_delta_sigma.acc[6] ),
    .B(_2345_),
    .Y(_3047_));
 sg13g2_nand2_1 _7513_ (.Y(_3048_),
    .A(\i_delta_sigma.acc[6] ),
    .B(_2345_));
 sg13g2_inv_1 _7514_ (.Y(_3049_),
    .A(_3048_));
 sg13g2_nor2_1 _7515_ (.A(_3047_),
    .B(_3049_),
    .Y(_3050_));
 sg13g2_nor2b_1 _7516_ (.A(_3046_),
    .B_N(_3050_),
    .Y(_3051_));
 sg13g2_a21oi_1 _7517_ (.A1(_3043_),
    .A2(_3048_),
    .Y(_3052_),
    .B1(_3042_));
 sg13g2_a21oi_1 _7518_ (.A1(_3041_),
    .A2(_3051_),
    .Y(_3053_),
    .B1(_3052_));
 sg13g2_inv_1 _7519_ (.Y(_3054_),
    .A(_3053_));
 sg13g2_nor2_1 _7520_ (.A(\i_delta_sigma.acc[9] ),
    .B(_2318_),
    .Y(_3055_));
 sg13g2_nand2_1 _7521_ (.Y(_3056_),
    .A(\i_delta_sigma.acc[9] ),
    .B(_2318_));
 sg13g2_inv_1 _7522_ (.Y(_3057_),
    .A(_3056_));
 sg13g2_nor2_1 _7523_ (.A(_3055_),
    .B(_3057_),
    .Y(_3058_));
 sg13g2_inv_1 _7524_ (.Y(_3059_),
    .A(_3058_));
 sg13g2_nor2_1 _7525_ (.A(\i_delta_sigma.acc[8] ),
    .B(_2365_),
    .Y(_3060_));
 sg13g2_nand2_1 _7526_ (.Y(_3061_),
    .A(\i_delta_sigma.acc[8] ),
    .B(_2365_));
 sg13g2_nor2b_1 _7527_ (.A(_3060_),
    .B_N(_3061_),
    .Y(_3062_));
 sg13g2_inv_1 _7528_ (.Y(_3063_),
    .A(_3062_));
 sg13g2_nor2_1 _7529_ (.A(_3059_),
    .B(_3063_),
    .Y(_3064_));
 sg13g2_a21oi_1 _7530_ (.A1(_3056_),
    .A2(_3061_),
    .Y(_3065_),
    .B1(_3055_));
 sg13g2_a21oi_1 _7531_ (.A1(_3054_),
    .A2(_3064_),
    .Y(_3066_),
    .B1(_3065_));
 sg13g2_nor2_1 _7532_ (.A(_3020_),
    .B(_3066_),
    .Y(_3067_));
 sg13g2_nor2b_1 _7533_ (.A(_3019_),
    .B_N(_3066_),
    .Y(_3068_));
 sg13g2_nor3_1 _7534_ (.A(_2735_),
    .B(_3067_),
    .C(_3068_),
    .Y(_0093_));
 sg13g2_nor2_1 _7535_ (.A(\i_delta_sigma.acc[11] ),
    .B(net155),
    .Y(_3069_));
 sg13g2_nand2_1 _7536_ (.Y(_3070_),
    .A(\i_delta_sigma.acc[11] ),
    .B(net155));
 sg13g2_inv_1 _7537_ (.Y(_3071_),
    .A(_3070_));
 sg13g2_nor2_1 _7538_ (.A(_3069_),
    .B(_3071_),
    .Y(_3072_));
 sg13g2_inv_1 _7539_ (.Y(_3073_),
    .A(_3041_));
 sg13g2_o21ai_1 _7540_ (.B1(_3048_),
    .Y(_3074_),
    .A1(_3047_),
    .A2(_3073_));
 sg13g2_nor2_1 _7541_ (.A(_3046_),
    .B(_3063_),
    .Y(_3075_));
 sg13g2_a21oi_1 _7542_ (.A1(_3061_),
    .A2(_3043_),
    .Y(_3076_),
    .B1(_3060_));
 sg13g2_a21oi_1 _7543_ (.A1(_3074_),
    .A2(_3075_),
    .Y(_3077_),
    .B1(_3076_));
 sg13g2_nor2_1 _7544_ (.A(_3059_),
    .B(_3077_),
    .Y(_3078_));
 sg13g2_nor3_1 _7545_ (.A(_3018_),
    .B(_3057_),
    .C(_3078_),
    .Y(_3079_));
 sg13g2_nor2_1 _7546_ (.A(_3016_),
    .B(_3079_),
    .Y(_3080_));
 sg13g2_xor2_1 _7547_ (.B(_3080_),
    .A(_3072_),
    .X(_3081_));
 sg13g2_nor2_1 _7548_ (.A(net140),
    .B(_3081_),
    .Y(_0094_));
 sg13g2_xor2_1 _7549_ (.B(\i_delta_sigma.acc[12] ),
    .A(_2331_),
    .X(_3082_));
 sg13g2_nor3_1 _7550_ (.A(_3018_),
    .B(_3071_),
    .C(_3067_),
    .Y(_3083_));
 sg13g2_nor2_1 _7551_ (.A(_3069_),
    .B(_3083_),
    .Y(_3084_));
 sg13g2_xnor2_1 _7552_ (.Y(_3085_),
    .A(_3082_),
    .B(_3084_));
 sg13g2_xnor2_1 _7553_ (.Y(_3086_),
    .A(_0055_),
    .B(_3085_));
 sg13g2_and2_1 _7554_ (.A(_3086_),
    .B(_3081_),
    .X(_3087_));
 sg13g2_o21ai_1 _7555_ (.B1(net151),
    .Y(_3088_),
    .A1(_3081_),
    .A2(_3086_));
 sg13g2_nor2_1 _7556_ (.A(_3087_),
    .B(_3088_),
    .Y(_0095_));
 sg13g2_xnor2_1 _7557_ (.Y(_3089_),
    .A(_0055_),
    .B(\i_delta_sigma.acc[13] ));
 sg13g2_xnor2_1 _7558_ (.Y(_3090_),
    .A(_2336_),
    .B(_3089_));
 sg13g2_nand3_1 _7559_ (.B(_3072_),
    .C(_3082_),
    .A(_3080_),
    .Y(_3091_));
 sg13g2_o21ai_1 _7560_ (.B1(_2331_),
    .Y(_3092_),
    .A1(\i_delta_sigma.acc[11] ),
    .A2(\i_delta_sigma.acc[12] ));
 sg13g2_nand2_1 _7561_ (.Y(_3093_),
    .A(_3091_),
    .B(_3092_));
 sg13g2_xnor2_1 _7562_ (.Y(_3094_),
    .A(_3090_),
    .B(_3093_));
 sg13g2_nor2_1 _7563_ (.A(\i_delta_sigma.acc[13] ),
    .B(_3085_),
    .Y(_3095_));
 sg13g2_nor2_1 _7564_ (.A(_3095_),
    .B(_3087_),
    .Y(_3096_));
 sg13g2_xor2_1 _7565_ (.B(_3096_),
    .A(_3094_),
    .X(_3097_));
 sg13g2_nor2_1 _7566_ (.A(net140),
    .B(_3097_),
    .Y(_0096_));
 sg13g2_nor2_1 _7567_ (.A(_3015_),
    .B(_3023_),
    .Y(_3098_));
 sg13g2_nor3_1 _7568_ (.A(net135),
    .B(_3098_),
    .C(_3025_),
    .Y(_0097_));
 sg13g2_nor2_1 _7569_ (.A(_3028_),
    .B(_3027_),
    .Y(_3099_));
 sg13g2_nor3_1 _7570_ (.A(net135),
    .B(_3099_),
    .C(_3030_),
    .Y(_0098_));
 sg13g2_nor2b_1 _7571_ (.A(_3033_),
    .B_N(_3032_),
    .Y(_3100_));
 sg13g2_nor2b_1 _7572_ (.A(_3031_),
    .B_N(_3100_),
    .Y(_3101_));
 sg13g2_nor2b_1 _7573_ (.A(_3100_),
    .B_N(_3031_),
    .Y(_3102_));
 sg13g2_nor3_1 _7574_ (.A(_2735_),
    .B(_3101_),
    .C(_3102_),
    .Y(_0099_));
 sg13g2_nor2b_1 _7575_ (.A(_3022_),
    .B_N(_3036_),
    .Y(_3103_));
 sg13g2_o21ai_1 _7576_ (.B1(net150),
    .Y(_3104_),
    .A1(_3103_),
    .A2(_3034_));
 sg13g2_a21oi_1 _7577_ (.A1(_3034_),
    .A2(_3103_),
    .Y(_0100_),
    .B1(_3104_));
 sg13g2_nor2b_1 _7578_ (.A(_3021_),
    .B_N(_3039_),
    .Y(_3105_));
 sg13g2_o21ai_1 _7579_ (.B1(net150),
    .Y(_3106_),
    .A1(_3105_),
    .A2(_3037_));
 sg13g2_a21oi_1 _7580_ (.A1(_3037_),
    .A2(_3105_),
    .Y(_0101_),
    .B1(_3106_));
 sg13g2_o21ai_1 _7581_ (.B1(net150),
    .Y(_3107_),
    .A1(_3050_),
    .A2(_3041_));
 sg13g2_a21oi_1 _7582_ (.A1(_3050_),
    .A2(_3041_),
    .Y(_0102_),
    .B1(_3107_));
 sg13g2_xnor2_1 _7583_ (.Y(_3108_),
    .A(_3045_),
    .B(_3074_));
 sg13g2_nor2_1 _7584_ (.A(net140),
    .B(_3108_),
    .Y(_0103_));
 sg13g2_o21ai_1 _7585_ (.B1(net150),
    .Y(_3109_),
    .A1(_3063_),
    .A2(_3053_));
 sg13g2_a21oi_1 _7586_ (.A1(_3063_),
    .A2(_3053_),
    .Y(_0104_),
    .B1(_3109_));
 sg13g2_nor2b_1 _7587_ (.A(_3058_),
    .B_N(_3077_),
    .Y(_3110_));
 sg13g2_nor3_1 _7588_ (.A(net135),
    .B(_3078_),
    .C(_3110_),
    .Y(_0105_));
 sg13g2_nor2_1 _7589_ (.A(_3550_),
    .B(_2256_),
    .Y(_3111_));
 sg13g2_nor2_1 _7590_ (.A(_2741_),
    .B(_3621_),
    .Y(_3112_));
 sg13g2_nor4_1 _7591_ (.A(_2266_),
    .B(_3111_),
    .C(_3112_),
    .D(_1887_),
    .Y(_3113_));
 sg13g2_nand3_1 _7592_ (.B(_3522_),
    .C(_3502_),
    .A(_3524_),
    .Y(_3114_));
 sg13g2_nor3_1 _7593_ (.A(_3545_),
    .B(_3114_),
    .C(_1748_),
    .Y(_3115_));
 sg13g2_nor4_1 _7594_ (.A(_3512_),
    .B(net182),
    .C(_3509_),
    .D(_3510_),
    .Y(_3116_));
 sg13g2_nor2b_1 _7595_ (.A(_2251_),
    .B_N(_3116_),
    .Y(_3117_));
 sg13g2_a221oi_1 _7596_ (.B2(_2257_),
    .C1(_2259_),
    .B1(_3520_),
    .A1(_3117_),
    .Y(_3118_),
    .A2(_2255_));
 sg13g2_nor2_1 _7597_ (.A(_3111_),
    .B(_3112_),
    .Y(_3119_));
 sg13g2_nand2_1 _7598_ (.Y(_3120_),
    .A(_3118_),
    .B(_3119_));
 sg13g2_inv_1 _7599_ (.Y(_3121_),
    .A(_3120_));
 sg13g2_a21oi_1 _7600_ (.A1(_3121_),
    .A2(_3115_),
    .Y(_3122_),
    .B1(_2266_));
 sg13g2_a21o_1 _7601_ (.A2(_3115_),
    .A1(_3113_),
    .B1(_3122_),
    .X(_3123_));
 sg13g2_inv_1 _7602_ (.Y(_3124_),
    .A(\i_orchestrator.hit_bottom ));
 sg13g2_nand2_1 _7603_ (.Y(_3125_),
    .A(_2267_),
    .B(net183));
 sg13g2_a21oi_1 _7604_ (.A1(_3123_),
    .A2(_3124_),
    .Y(_0142_),
    .B1(_3125_));
 sg13g2_nand2_1 _7605_ (.Y(_3126_),
    .A(_1887_),
    .B(_3111_));
 sg13g2_inv_1 _7606_ (.Y(_3127_),
    .A(_2241_));
 sg13g2_a21oi_1 _7607_ (.A1(_3126_),
    .A2(_3127_),
    .Y(_0143_),
    .B1(_3125_));
 sg13g2_buf_1 _7608_ (.A(\i_orchestrator.hit_priority[0] ),
    .X(_3128_));
 sg13g2_inv_1 _7609_ (.Y(_3129_),
    .A(_3128_));
 sg13g2_nand2_1 _7610_ (.Y(_3130_),
    .A(_2255_),
    .B(_3117_));
 sg13g2_buf_1 _7611_ (.A(_3130_),
    .X(_3131_));
 sg13g2_o21ai_1 _7612_ (.B1(_2952_),
    .Y(_3132_),
    .A1(_0066_),
    .A2(net87));
 sg13g2_a21oi_1 _7613_ (.A1(_3129_),
    .A2(net87),
    .Y(_0144_),
    .B1(_3132_));
 sg13g2_inv_1 _7614_ (.Y(_3133_),
    .A(\i_orchestrator.hit_priority[1] ));
 sg13g2_xor2_1 _7615_ (.B(\i_orchestrator.hit_priority[1] ),
    .A(_3128_),
    .X(_3134_));
 sg13g2_o21ai_1 _7616_ (.B1(_2952_),
    .Y(_3135_),
    .A1(_3134_),
    .A2(net87));
 sg13g2_a21oi_1 _7617_ (.A1(_3133_),
    .A2(net87),
    .Y(_0145_),
    .B1(_3135_));
 sg13g2_a22oi_1 _7618_ (.Y(_3136_),
    .B1(_3112_),
    .B2(_1887_),
    .A2(_2267_),
    .A1(\i_orchestrator.hit_right ));
 sg13g2_nor2_1 _7619_ (.A(_2265_),
    .B(_3136_),
    .Y(_0146_));
 sg13g2_nand2_1 _7620_ (.Y(_3137_),
    .A(_3116_),
    .B(_1729_));
 sg13g2_nor4_1 _7621_ (.A(_3521_),
    .B(_3503_),
    .C(_3545_),
    .D(_3137_),
    .Y(_3138_));
 sg13g2_a21oi_1 _7622_ (.A1(_3121_),
    .A2(_3138_),
    .Y(_3139_),
    .B1(_2266_));
 sg13g2_a21o_1 _7623_ (.A2(_3138_),
    .A1(_3113_),
    .B1(_3139_),
    .X(_3140_));
 sg13g2_inv_1 _7624_ (.Y(_3141_),
    .A(\i_orchestrator.hit_top ));
 sg13g2_a21oi_1 _7625_ (.A1(_3140_),
    .A2(_3141_),
    .Y(_0147_),
    .B1(_3125_));
 sg13g2_inv_1 _7626_ (.Y(_3142_),
    .A(_3130_));
 sg13g2_buf_1 _7627_ (.A(_3142_),
    .X(_3143_));
 sg13g2_xor2_1 _7628_ (.B(\i_orchestrator.lfsr[6] ),
    .A(_3484_),
    .X(_3144_));
 sg13g2_a21oi_1 _7629_ (.A1(net85),
    .A2(_3144_),
    .Y(_3145_),
    .B1(net168));
 sg13g2_o21ai_1 _7630_ (.B1(_3145_),
    .Y(_0148_),
    .A1(_2780_),
    .A2(net85));
 sg13g2_o21ai_1 _7631_ (.B1(net169),
    .Y(_3146_),
    .A1(_2780_),
    .A2(net87));
 sg13g2_a21o_1 _7632_ (.A2(net87),
    .A1(\i_orchestrator.lfsr[1] ),
    .B1(_3146_),
    .X(_0149_));
 sg13g2_inv_1 _7633_ (.Y(_3147_),
    .A(\i_orchestrator.lfsr[2] ));
 sg13g2_a21oi_1 _7634_ (.A1(net85),
    .A2(\i_orchestrator.lfsr[1] ),
    .Y(_3148_),
    .B1(net168));
 sg13g2_o21ai_1 _7635_ (.B1(_3148_),
    .Y(_0150_),
    .A1(_3147_),
    .A2(net85));
 sg13g2_o21ai_1 _7636_ (.B1(net169),
    .Y(_3149_),
    .A1(_3147_),
    .A2(net87));
 sg13g2_a21o_1 _7637_ (.A2(net87),
    .A1(\i_orchestrator.lfsr[3] ),
    .B1(_3149_),
    .X(_0151_));
 sg13g2_inv_1 _7638_ (.Y(_3150_),
    .A(\i_orchestrator.lfsr[4] ));
 sg13g2_a21oi_1 _7639_ (.A1(net85),
    .A2(\i_orchestrator.lfsr[3] ),
    .Y(_3151_),
    .B1(_3493_));
 sg13g2_o21ai_1 _7640_ (.B1(_3151_),
    .Y(_0152_),
    .A1(_3150_),
    .A2(net85));
 sg13g2_o21ai_1 _7641_ (.B1(_3483_),
    .Y(_3152_),
    .A1(_3150_),
    .A2(_3130_));
 sg13g2_a21o_1 _7642_ (.A2(_3131_),
    .A1(\i_orchestrator.lfsr[5] ),
    .B1(_3152_),
    .X(_0153_));
 sg13g2_inv_1 _7643_ (.Y(_3153_),
    .A(\i_orchestrator.lfsr[6] ));
 sg13g2_a21oi_1 _7644_ (.A1(net85),
    .A2(\i_orchestrator.lfsr[5] ),
    .Y(_3154_),
    .B1(net168));
 sg13g2_o21ai_1 _7645_ (.B1(_3154_),
    .Y(_0154_),
    .A1(_3153_),
    .A2(net85));
 sg13g2_o21ai_1 _7646_ (.B1(_3483_),
    .Y(_3155_),
    .A1(_3153_),
    .A2(_3130_));
 sg13g2_a21o_1 _7647_ (.A2(_3131_),
    .A1(\i_orchestrator.lfsr[7] ),
    .B1(_3155_),
    .X(_0155_));
 sg13g2_inv_1 _7648_ (.Y(_3156_),
    .A(_2992_));
 sg13g2_a21oi_1 _7649_ (.A1(_3142_),
    .A2(\i_orchestrator.lfsr[7] ),
    .Y(_3157_),
    .B1(net168));
 sg13g2_o21ai_1 _7650_ (.B1(_3157_),
    .Y(_0156_),
    .A1(_3156_),
    .A2(_3143_));
 sg13g2_a21oi_1 _7651_ (.A1(_3142_),
    .A2(_2992_),
    .Y(_3158_),
    .B1(net168));
 sg13g2_o21ai_1 _7652_ (.B1(_3158_),
    .Y(_0157_),
    .A1(_3487_),
    .A2(_3143_));
 sg13g2_nand2_1 _7653_ (.Y(_3159_),
    .A(_3124_),
    .B(\i_orchestrator.hit_top ));
 sg13g2_nand3_1 _7654_ (.B(_0057_),
    .C(_3128_),
    .A(_3133_),
    .Y(_3160_));
 sg13g2_a21oi_1 _7655_ (.A1(_0012_),
    .A2(_3159_),
    .Y(_3161_),
    .B1(_3160_));
 sg13g2_inv_1 _7656_ (.Y(_3162_),
    .A(\i_orchestrator.hit_right ));
 sg13g2_nand2_1 _7657_ (.Y(_3163_),
    .A(_3162_),
    .B(_2241_));
 sg13g2_nand3_1 _7658_ (.B(_3133_),
    .C(_0005_),
    .A(_3129_),
    .Y(_3164_));
 sg13g2_a21oi_1 _7659_ (.A1(_0056_),
    .A2(_3163_),
    .Y(_3165_),
    .B1(_3164_));
 sg13g2_nand2_1 _7660_ (.Y(_3166_),
    .A(_3129_),
    .B(\i_orchestrator.hit_priority[1] ));
 sg13g2_a21oi_1 _7661_ (.A1(_3124_),
    .A2(_2241_),
    .Y(_3167_),
    .B1(\i_orchestrator.hit_top ));
 sg13g2_o21ai_1 _7662_ (.B1(_0012_),
    .Y(_3168_),
    .A1(\i_orchestrator.hit_right ),
    .A2(_3141_));
 sg13g2_nand3_1 _7663_ (.B(_3128_),
    .C(\i_orchestrator.hit_priority[1] ),
    .A(_3168_),
    .Y(_3169_));
 sg13g2_o21ai_1 _7664_ (.B1(_3169_),
    .Y(_3170_),
    .A1(_3166_),
    .A2(_3167_));
 sg13g2_nor3_1 _7665_ (.A(_3161_),
    .B(_3165_),
    .C(_3170_),
    .Y(_3171_));
 sg13g2_nand2_1 _7666_ (.Y(_3172_),
    .A(_3142_),
    .B(net183));
 sg13g2_nor2_1 _7667_ (.A(_3171_),
    .B(_3172_),
    .Y(_0158_));
 sg13g2_nand2_1 _7668_ (.Y(_3173_),
    .A(_3124_),
    .B(_3141_));
 sg13g2_a221oi_1 _7669_ (.B2(_3173_),
    .C1(_3172_),
    .B1(_3129_),
    .A1(_3127_),
    .Y(_0159_),
    .A2(_3162_));
 sg13g2_nand2_1 _7670_ (.Y(_3174_),
    .A(_2880_),
    .B(_0065_));
 sg13g2_inv_1 _7671_ (.Y(_0160_),
    .A(_3174_));
 sg13g2_nor2_1 _7672_ (.A(\i_orchestrator.sample_counter[1] ),
    .B(\i_orchestrator.sample_counter[0] ),
    .Y(_3175_));
 sg13g2_nand2_1 _7673_ (.Y(_3176_),
    .A(\i_orchestrator.sample_counter[1] ),
    .B(\i_orchestrator.sample_counter[0] ));
 sg13g2_inv_1 _7674_ (.Y(_3177_),
    .A(_3176_));
 sg13g2_nor3_1 _7675_ (.A(net135),
    .B(_3175_),
    .C(_3177_),
    .Y(_0161_));
 sg13g2_nor2b_1 _7676_ (.A(_3176_),
    .B_N(\i_orchestrator.sample_counter[2] ),
    .Y(_3178_));
 sg13g2_nor2_1 _7677_ (.A(\i_orchestrator.sample_counter[2] ),
    .B(_3177_),
    .Y(_3179_));
 sg13g2_nor3_1 _7678_ (.A(_2264_),
    .B(_3178_),
    .C(_3179_),
    .Y(_0162_));
 sg13g2_nor2_1 _7679_ (.A(\i_orchestrator.sample_counter[3] ),
    .B(_3178_),
    .Y(_3180_));
 sg13g2_nand2_1 _7680_ (.Y(_3181_),
    .A(_3178_),
    .B(\i_orchestrator.sample_counter[3] ));
 sg13g2_inv_1 _7681_ (.Y(_3182_),
    .A(_3181_));
 sg13g2_nor3_1 _7682_ (.A(_2264_),
    .B(_3180_),
    .C(_3182_),
    .Y(_0163_));
 sg13g2_inv_1 _7683_ (.Y(_3183_),
    .A(\i_orchestrator.sample_counter[4] ));
 sg13g2_nor2_1 _7684_ (.A(_3183_),
    .B(_3181_),
    .Y(_3184_));
 sg13g2_nor2_1 _7685_ (.A(\i_orchestrator.sample_counter[4] ),
    .B(_3182_),
    .Y(_3185_));
 sg13g2_nor3_1 _7686_ (.A(net141),
    .B(_3184_),
    .C(_3185_),
    .Y(_0164_));
 sg13g2_nor2_1 _7687_ (.A(\i_orchestrator.sample_counter[5] ),
    .B(_3184_),
    .Y(_3186_));
 sg13g2_and2_1 _7688_ (.A(_3184_),
    .B(\i_orchestrator.sample_counter[5] ),
    .X(_3187_));
 sg13g2_nor3_1 _7689_ (.A(net141),
    .B(_3186_),
    .C(_3187_),
    .Y(_0165_));
 sg13g2_nor2_1 _7690_ (.A(\i_orchestrator.sample_counter[6] ),
    .B(_3187_),
    .Y(_3188_));
 sg13g2_nand2_1 _7691_ (.Y(_3189_),
    .A(_3187_),
    .B(\i_orchestrator.sample_counter[6] ));
 sg13g2_inv_1 _7692_ (.Y(_3190_),
    .A(_3189_));
 sg13g2_nor3_1 _7693_ (.A(net141),
    .B(_3188_),
    .C(_3190_),
    .Y(_0166_));
 sg13g2_nor2b_1 _7694_ (.A(_3189_),
    .B_N(\i_orchestrator.sample_counter[7] ),
    .Y(_3191_));
 sg13g2_nor2_1 _7695_ (.A(\i_orchestrator.sample_counter[7] ),
    .B(_3190_),
    .Y(_3192_));
 sg13g2_nor3_1 _7696_ (.A(net141),
    .B(_3191_),
    .C(_3192_),
    .Y(_0167_));
 sg13g2_nor2_1 _7697_ (.A(\i_orchestrator.sample_counter[8] ),
    .B(_3191_),
    .Y(_3193_));
 sg13g2_nand2_1 _7698_ (.Y(_3194_),
    .A(_3191_),
    .B(\i_orchestrator.sample_counter[8] ));
 sg13g2_inv_1 _7699_ (.Y(_3195_),
    .A(_3194_));
 sg13g2_nor3_1 _7700_ (.A(net141),
    .B(_3193_),
    .C(_3195_),
    .Y(_0168_));
 sg13g2_o21ai_1 _7701_ (.B1(net150),
    .Y(_3196_),
    .A1(\i_orchestrator.sample_counter[9] ),
    .A2(_3195_));
 sg13g2_a21oi_1 _7702_ (.A1(\i_orchestrator.sample_counter[9] ),
    .A2(_3195_),
    .Y(_0169_),
    .B1(_3196_));
 sg13g2_inv_1 _7703_ (.Y(_3197_),
    .A(\i_orchestrator.tension[1] ));
 sg13g2_nor3_1 _7704_ (.A(_2241_),
    .B(\i_orchestrator.hit_right ),
    .C(_3173_),
    .Y(_3198_));
 sg13g2_nor3_1 _7705_ (.A(_2240_),
    .B(_3198_),
    .C(_2248_),
    .Y(_3199_));
 sg13g2_nand2_1 _7706_ (.Y(_3200_),
    .A(_2259_),
    .B(_3199_));
 sg13g2_o21ai_1 _7707_ (.B1(net169),
    .Y(_3201_),
    .A1(_0005_),
    .A2(_3200_));
 sg13g2_a21oi_1 _7708_ (.A1(_3197_),
    .A2(_3200_),
    .Y(_0170_),
    .B1(_3201_));
 sg13g2_inv_1 _7709_ (.Y(_3202_),
    .A(\i_orchestrator.tension[2] ));
 sg13g2_nand3_1 _7710_ (.B(_2242_),
    .C(_3199_),
    .A(_2259_),
    .Y(_3203_));
 sg13g2_o21ai_1 _7711_ (.B1(net169),
    .Y(_3204_),
    .A1(_3162_),
    .A2(_3203_));
 sg13g2_a21oi_1 _7712_ (.A1(_3202_),
    .A2(_3200_),
    .Y(_0171_),
    .B1(_3204_));
 sg13g2_nand2_1 _7713_ (.Y(_3205_),
    .A(_3200_),
    .B(\i_orchestrator.tension[3] ));
 sg13g2_a21oi_1 _7714_ (.A1(_3205_),
    .A2(_3203_),
    .Y(_0172_),
    .B1(_2265_));
 sg13g2_a21oi_1 _7715_ (.A1(_2259_),
    .A2(_2247_),
    .Y(_3206_),
    .B1(\i_orchestrator.trigger_debounce ));
 sg13g2_o21ai_1 _7716_ (.B1(_2880_),
    .Y(_3207_),
    .A1(_2244_),
    .A2(_2260_));
 sg13g2_nor2_1 _7717_ (.A(_3206_),
    .B(_3207_),
    .Y(_0173_));
 sg13g2_nor2_1 _7718_ (.A(_3198_),
    .B(_3172_),
    .Y(_0176_));
 sg13g2_nor4_1 _7719_ (.A(\i_orchestrator.sample_counter[2] ),
    .B(\i_orchestrator.sample_counter[5] ),
    .C(\i_orchestrator.sample_counter[4] ),
    .D(\i_orchestrator.sample_counter[7] ),
    .Y(_3208_));
 sg13g2_nor4_1 _7720_ (.A(\i_orchestrator.sample_counter[1] ),
    .B(\i_orchestrator.sample_counter[0] ),
    .C(_3492_),
    .D(\i_orchestrator.sample_counter[3] ),
    .Y(_3209_));
 sg13g2_nand2_1 _7721_ (.Y(_3210_),
    .A(_3208_),
    .B(_3209_));
 sg13g2_nor4_1 _7722_ (.A(\i_orchestrator.sample_counter[6] ),
    .B(\i_orchestrator.sample_counter[9] ),
    .C(\i_orchestrator.sample_counter[8] ),
    .D(_3210_),
    .Y(_0178_));
 sg13g2_nor2_1 _7723_ (.A(_0841_),
    .B(_3671_),
    .Y(_3211_));
 sg13g2_inv_1 _7724_ (.Y(_3212_),
    .A(_3211_));
 sg13g2_buf_1 _7725_ (.A(net57),
    .X(_3213_));
 sg13g2_nand2_1 _7726_ (.Y(_3214_),
    .A(net83),
    .B(_3907_));
 sg13g2_o21ai_1 _7727_ (.B1(_3214_),
    .Y(_3215_),
    .A1(net83),
    .A2(_3753_));
 sg13g2_xnor2_1 _7728_ (.Y(_3216_),
    .A(_0018_),
    .B(_3215_));
 sg13g2_o21ai_1 _7729_ (.B1(net122),
    .Y(_3217_),
    .A1(\i_transform.image_x[0] ),
    .A2(net56));
 sg13g2_a21oi_1 _7730_ (.A1(net56),
    .A2(_3216_),
    .Y(_0212_),
    .B1(_3217_));
 sg13g2_buf_1 _7731_ (.A(net123),
    .X(_3218_));
 sg13g2_nand2b_1 _7732_ (.Y(_3219_),
    .B(_3589_),
    .A_N(_3555_));
 sg13g2_nor4_2 _7733_ (.A(_3561_),
    .B(_3569_),
    .C(_0305_),
    .Y(_3220_),
    .D(_3219_));
 sg13g2_nand2_1 _7734_ (.Y(_3221_),
    .A(_3650_),
    .B(_3220_));
 sg13g2_inv_1 _7735_ (.Y(_3222_),
    .A(_3221_));
 sg13g2_a21oi_1 _7736_ (.A1(_0720_),
    .A2(net65),
    .Y(_3223_),
    .B1(_0827_));
 sg13g2_nor2_1 _7737_ (.A(net105),
    .B(_3223_),
    .Y(_0213_));
 sg13g2_nand2_1 _7738_ (.Y(_3224_),
    .A(_0793_),
    .B(_0813_));
 sg13g2_inv_1 _7739_ (.Y(_3225_),
    .A(_3224_));
 sg13g2_buf_1 _7740_ (.A(net71),
    .X(_3226_));
 sg13g2_nand2_1 _7741_ (.Y(_3227_),
    .A(net64),
    .B(_0722_));
 sg13g2_buf_1 _7742_ (.A(net123),
    .X(_3228_));
 sg13g2_a21oi_1 _7743_ (.A1(_3225_),
    .A2(_3227_),
    .Y(_0214_),
    .B1(net104));
 sg13g2_nand2_1 _7744_ (.Y(_3229_),
    .A(_0744_),
    .B(_0769_));
 sg13g2_a21oi_1 _7745_ (.A1(_0730_),
    .A2(net65),
    .Y(_3230_),
    .B1(_3229_));
 sg13g2_nor2_1 _7746_ (.A(net105),
    .B(_3230_),
    .Y(_0215_));
 sg13g2_nand2_1 _7747_ (.Y(_3231_),
    .A(_0961_),
    .B(_0985_));
 sg13g2_a21oi_1 _7748_ (.A1(_0954_),
    .A2(net65),
    .Y(_3232_),
    .B1(_3231_));
 sg13g2_nor2_1 _7749_ (.A(net105),
    .B(_3232_),
    .Y(_0216_));
 sg13g2_xnor2_1 _7750_ (.Y(_3233_),
    .A(_1872_),
    .B(net91));
 sg13g2_o21ai_1 _7751_ (.B1(_0956_),
    .Y(_3234_),
    .A1(_0942_),
    .A2(net92));
 sg13g2_inv_1 _7752_ (.Y(_3235_),
    .A(_3234_));
 sg13g2_nor2_1 _7753_ (.A(_3233_),
    .B(_3235_),
    .Y(_3236_));
 sg13g2_a21o_1 _7754_ (.A2(_3233_),
    .A1(_3235_),
    .B1(net58),
    .X(_3237_));
 sg13g2_inv_1 _7755_ (.Y(_3238_),
    .A(_0943_));
 sg13g2_a22oi_1 _7756_ (.Y(_3239_),
    .B1(_3238_),
    .B2(_0948_),
    .A2(_0750_),
    .A1(_0954_));
 sg13g2_buf_1 _7757_ (.A(_0046_),
    .X(_3240_));
 sg13g2_buf_1 _7758_ (.A(net91),
    .X(_3241_));
 sg13g2_xnor2_1 _7759_ (.Y(_3242_),
    .A(_3240_),
    .B(net86));
 sg13g2_a21oi_1 _7760_ (.A1(_3239_),
    .A2(_3242_),
    .Y(_3243_),
    .B1(net62));
 sg13g2_o21ai_1 _7761_ (.B1(_3243_),
    .Y(_3244_),
    .A1(_3239_),
    .A2(_3242_));
 sg13g2_o21ai_1 _7762_ (.B1(_3244_),
    .Y(_3245_),
    .A1(_3236_),
    .A2(_3237_));
 sg13g2_nand2_1 _7763_ (.Y(_3246_),
    .A(_0713_),
    .B(_0971_));
 sg13g2_inv_1 _7764_ (.Y(_3247_),
    .A(_0727_));
 sg13g2_buf_1 _7765_ (.A(_1390_),
    .X(_3248_));
 sg13g2_nor2_1 _7766_ (.A(_1875_),
    .B(net88),
    .Y(_3249_));
 sg13g2_a21oi_1 _7767_ (.A1(_0975_),
    .A2(_0942_),
    .Y(_3250_),
    .B1(_3249_));
 sg13g2_o21ai_1 _7768_ (.B1(_3250_),
    .Y(_3251_),
    .A1(_3246_),
    .A2(_3247_));
 sg13g2_xnor2_1 _7769_ (.Y(_3252_),
    .A(_3240_),
    .B(net98));
 sg13g2_inv_1 _7770_ (.Y(_3253_),
    .A(_3252_));
 sg13g2_a21oi_1 _7771_ (.A1(_3251_),
    .A2(_3253_),
    .Y(_3254_),
    .B1(net74));
 sg13g2_o21ai_1 _7772_ (.B1(_3254_),
    .Y(_3255_),
    .A1(_3251_),
    .A2(_3253_));
 sg13g2_xnor2_1 _7773_ (.Y(_3256_),
    .A(_1872_),
    .B(net98));
 sg13g2_a21oi_1 _7774_ (.A1(_0986_),
    .A2(net88),
    .Y(_3257_),
    .B1(_0965_));
 sg13g2_nor2_1 _7775_ (.A(_3256_),
    .B(_3257_),
    .Y(_3258_));
 sg13g2_a21oi_1 _7776_ (.A1(_3257_),
    .A2(_3256_),
    .Y(_3259_),
    .B1(net73));
 sg13g2_nand2b_1 _7777_ (.Y(_3260_),
    .B(_3259_),
    .A_N(_3258_));
 sg13g2_a21oi_1 _7778_ (.A1(_3255_),
    .A2(_3260_),
    .Y(_3261_),
    .B1(_0333_));
 sg13g2_a221oi_1 _7779_ (.B2(_3652_),
    .C1(_3261_),
    .B1(_3245_),
    .A1(_1872_),
    .Y(_3262_),
    .A2(_0337_));
 sg13g2_nor2_1 _7780_ (.A(net105),
    .B(_3262_),
    .Y(_0217_));
 sg13g2_inv_1 _7781_ (.Y(_3263_),
    .A(_3240_));
 sg13g2_a21oi_1 _7782_ (.A1(_3263_),
    .A2(net88),
    .Y(_3264_),
    .B1(_3258_));
 sg13g2_xnor2_1 _7783_ (.Y(_3265_),
    .A(net180),
    .B(net88));
 sg13g2_o21ai_1 _7784_ (.B1(net74),
    .Y(_3266_),
    .A1(_3265_),
    .A2(_3264_));
 sg13g2_a21oi_1 _7785_ (.A1(_3264_),
    .A2(_3265_),
    .Y(_3267_),
    .B1(_3266_));
 sg13g2_nand2_1 _7786_ (.Y(_3268_),
    .A(_0971_),
    .B(_3253_));
 sg13g2_inv_1 _7787_ (.Y(_3269_),
    .A(_0982_));
 sg13g2_a22oi_1 _7788_ (.Y(_3270_),
    .B1(_3240_),
    .B2(_3249_),
    .A2(_1872_),
    .A1(net114));
 sg13g2_o21ai_1 _7789_ (.B1(_3270_),
    .Y(_3271_),
    .A1(_3268_),
    .A2(_3269_));
 sg13g2_inv_1 _7790_ (.Y(_3272_),
    .A(_0063_));
 sg13g2_xnor2_1 _7791_ (.Y(_3273_),
    .A(_3272_),
    .B(net88));
 sg13g2_a21oi_1 _7792_ (.A1(_3271_),
    .A2(_3273_),
    .Y(_3274_),
    .B1(net74));
 sg13g2_o21ai_1 _7793_ (.B1(_3274_),
    .Y(_3275_),
    .A1(_3271_),
    .A2(_3273_));
 sg13g2_nand2b_1 _7794_ (.Y(_3276_),
    .B(_3275_),
    .A_N(_3267_));
 sg13g2_a22oi_1 _7795_ (.Y(_3277_),
    .B1(_0687_),
    .B2(_3276_),
    .A2(net64),
    .A1(net180));
 sg13g2_xnor2_1 _7796_ (.Y(_3278_),
    .A(_3272_),
    .B(net86));
 sg13g2_nor2_1 _7797_ (.A(_0943_),
    .B(_3242_),
    .Y(_3279_));
 sg13g2_nor3_1 _7798_ (.A(_1875_),
    .B(_3263_),
    .C(net86),
    .Y(_3280_));
 sg13g2_a221oi_1 _7799_ (.B2(_3279_),
    .C1(_3280_),
    .B1(_0948_),
    .A1(_1872_),
    .Y(_3281_),
    .A2(net92));
 sg13g2_xor2_1 _7800_ (.B(_3281_),
    .A(_3278_),
    .X(_3282_));
 sg13g2_a21oi_1 _7801_ (.A1(_3263_),
    .A2(net86),
    .Y(_3283_),
    .B1(_3236_));
 sg13g2_xnor2_1 _7802_ (.Y(_3284_),
    .A(net180),
    .B(net86));
 sg13g2_a21oi_1 _7803_ (.A1(_3283_),
    .A2(_3284_),
    .Y(_3285_),
    .B1(_0501_));
 sg13g2_o21ai_1 _7804_ (.B1(_3285_),
    .Y(_3286_),
    .A1(_3283_),
    .A2(_3284_));
 sg13g2_o21ai_1 _7805_ (.B1(_3286_),
    .Y(_3287_),
    .A1(net59),
    .A2(_3282_));
 sg13g2_nand2_1 _7806_ (.Y(_3288_),
    .A(_3287_),
    .B(_0689_));
 sg13g2_a21oi_1 _7807_ (.A1(_3277_),
    .A2(_3288_),
    .Y(_0218_),
    .B1(net104));
 sg13g2_o21ai_1 _7808_ (.B1(net82),
    .Y(_3289_),
    .A1(_0364_),
    .A2(_0373_));
 sg13g2_a21oi_1 _7809_ (.A1(_0364_),
    .A2(_0373_),
    .Y(_3290_),
    .B1(_3289_));
 sg13g2_nor2_1 _7810_ (.A(_3290_),
    .B(_3211_),
    .Y(_3291_));
 sg13g2_a21oi_1 _7811_ (.A1(_0480_),
    .A2(_0486_),
    .Y(_3292_),
    .B1(net84));
 sg13g2_o21ai_1 _7812_ (.B1(_3292_),
    .Y(_3293_),
    .A1(_0486_),
    .A2(_0480_));
 sg13g2_a221oi_1 _7813_ (.B2(_3293_),
    .C1(net112),
    .B1(_3291_),
    .A1(_0370_),
    .Y(_0219_),
    .A2(_3211_));
 sg13g2_xor2_1 _7814_ (.B(_0570_),
    .A(_0477_),
    .X(_3294_));
 sg13g2_nor2_1 _7815_ (.A(_0537_),
    .B(_0369_),
    .Y(_3295_));
 sg13g2_nor2_1 _7816_ (.A(net81),
    .B(_3295_),
    .Y(_3296_));
 sg13g2_a22oi_1 _7817_ (.Y(_3297_),
    .B1(_0538_),
    .B2(_3296_),
    .A2(_3220_),
    .A1(_3294_));
 sg13g2_o21ai_1 _7818_ (.B1(net122),
    .Y(_3298_),
    .A1(\i_transform.image_x[2] ),
    .A2(net57));
 sg13g2_a21oi_1 _7819_ (.A1(_3297_),
    .A2(net56),
    .Y(_0220_),
    .B1(_3298_));
 sg13g2_xnor2_1 _7820_ (.Y(_3299_),
    .A(_0377_),
    .B(_0539_));
 sg13g2_inv_1 _7821_ (.Y(_3300_),
    .A(_0573_));
 sg13g2_a21oi_1 _7822_ (.A1(_3300_),
    .A2(_0476_),
    .Y(_3301_),
    .B1(net82));
 sg13g2_a22oi_1 _7823_ (.Y(_3302_),
    .B1(_0574_),
    .B2(_3301_),
    .A2(net82),
    .A1(_3299_));
 sg13g2_o21ai_1 _7824_ (.B1(net122),
    .Y(_3303_),
    .A1(_0375_),
    .A2(net57));
 sg13g2_a21oi_1 _7825_ (.A1(_3302_),
    .A2(net56),
    .Y(_0221_),
    .B1(_3303_));
 sg13g2_xnor2_1 _7826_ (.Y(_3304_),
    .A(_0382_),
    .B(_0542_));
 sg13g2_inv_1 _7827_ (.Y(_3305_),
    .A(_0576_));
 sg13g2_nor2_1 _7828_ (.A(_0484_),
    .B(_3305_),
    .Y(_3306_));
 sg13g2_inv_1 _7829_ (.Y(_3307_),
    .A(_3306_));
 sg13g2_a21oi_1 _7830_ (.A1(_3305_),
    .A2(_0484_),
    .Y(_3308_),
    .B1(net82));
 sg13g2_a22oi_1 _7831_ (.Y(_3309_),
    .B1(_3307_),
    .B2(_3308_),
    .A2(net82),
    .A1(_3304_));
 sg13g2_o21ai_1 _7832_ (.B1(net122),
    .Y(_3310_),
    .A1(_0378_),
    .A2(net57));
 sg13g2_a21oi_1 _7833_ (.A1(_3309_),
    .A2(net56),
    .Y(_0222_),
    .B1(_3310_));
 sg13g2_xnor2_1 _7834_ (.Y(_3311_),
    .A(_0398_),
    .B(_3753_));
 sg13g2_a21oi_1 _7835_ (.A1(net70),
    .A2(_3311_),
    .Y(_3312_),
    .B1(net83));
 sg13g2_a21oi_1 _7836_ (.A1(_0980_),
    .A2(_0544_),
    .Y(_3313_),
    .B1(net70));
 sg13g2_o21ai_1 _7837_ (.B1(_3313_),
    .Y(_3314_),
    .A1(_0544_),
    .A2(_0980_));
 sg13g2_a22oi_1 _7838_ (.Y(_3315_),
    .B1(_3312_),
    .B2(_3314_),
    .A2(net64),
    .A1(\i_transform.image_x[5] ));
 sg13g2_o21ai_1 _7839_ (.B1(_0559_),
    .Y(_3316_),
    .A1(_0451_),
    .A2(_3306_));
 sg13g2_nand3_1 _7840_ (.B(_0560_),
    .C(_0450_),
    .A(_3307_),
    .Y(_3317_));
 sg13g2_nand3_1 _7841_ (.B(_3317_),
    .C(net58),
    .A(_3316_),
    .Y(_3318_));
 sg13g2_xnor2_1 _7842_ (.Y(_3319_),
    .A(_0398_),
    .B(_3920_));
 sg13g2_a21oi_1 _7843_ (.A1(net59),
    .A2(_3319_),
    .Y(_3320_),
    .B1(net63));
 sg13g2_nand2_1 _7844_ (.Y(_3321_),
    .A(_3318_),
    .B(_3320_));
 sg13g2_a21oi_1 _7845_ (.A1(_3315_),
    .A2(_3321_),
    .Y(_0223_),
    .B1(net104));
 sg13g2_o21ai_1 _7846_ (.B1(_0599_),
    .Y(_3322_),
    .A1(_0544_),
    .A2(_0979_));
 sg13g2_a21oi_1 _7847_ (.A1(_3322_),
    .A2(_0361_),
    .Y(_3323_),
    .B1(net70));
 sg13g2_o21ai_1 _7848_ (.B1(_3323_),
    .Y(_3324_),
    .A1(_0361_),
    .A2(_3322_));
 sg13g2_nand2b_1 _7849_ (.Y(_3325_),
    .B(_0419_),
    .A_N(_0420_));
 sg13g2_nand3_1 _7850_ (.B(_0421_),
    .C(_3325_),
    .A(net70),
    .Y(_3326_));
 sg13g2_a21o_1 _7851_ (.A2(_3326_),
    .A1(_3324_),
    .B1(net83),
    .X(_3327_));
 sg13g2_a21oi_1 _7852_ (.A1(_0576_),
    .A2(_0567_),
    .Y(_3328_),
    .B1(_0626_));
 sg13g2_xnor2_1 _7853_ (.Y(_3329_),
    .A(_0562_),
    .B(_3328_));
 sg13g2_nand2b_1 _7854_ (.Y(_3330_),
    .B(_0503_),
    .A_N(_0504_));
 sg13g2_nand3_1 _7855_ (.B(_0505_),
    .C(_3330_),
    .A(net59),
    .Y(_3331_));
 sg13g2_o21ai_1 _7856_ (.B1(_3331_),
    .Y(_3332_),
    .A1(net59),
    .A2(_3329_));
 sg13g2_a22oi_1 _7857_ (.Y(_3333_),
    .B1(_3652_),
    .B2(_3332_),
    .A2(net64),
    .A1(_0357_));
 sg13g2_a21oi_1 _7858_ (.A1(_3327_),
    .A2(_3333_),
    .Y(_0224_),
    .B1(net104));
 sg13g2_nand2_1 _7859_ (.Y(_3334_),
    .A(_0672_),
    .B(_0692_));
 sg13g2_inv_1 _7860_ (.Y(_3335_),
    .A(_3334_));
 sg13g2_nand2_1 _7861_ (.Y(_3336_),
    .A(net64),
    .B(_0349_));
 sg13g2_a21oi_1 _7862_ (.A1(_3335_),
    .A2(_3336_),
    .Y(_0225_),
    .B1(net104));
 sg13g2_nand2_1 _7863_ (.Y(_3337_),
    .A(_0557_),
    .B(_0585_));
 sg13g2_a21oi_1 _7864_ (.A1(_0403_),
    .A2(net65),
    .Y(_3338_),
    .B1(_3337_));
 sg13g2_nor2_1 _7865_ (.A(net105),
    .B(_3338_),
    .Y(_0226_));
 sg13g2_inv_1 _7866_ (.Y(_3339_),
    .A(_0524_));
 sg13g2_nand2_1 _7867_ (.Y(_3340_),
    .A(net64),
    .B(_0607_));
 sg13g2_a21oi_1 _7868_ (.A1(_3339_),
    .A2(_3340_),
    .Y(_0227_),
    .B1(net104));
 sg13g2_nand2_1 _7869_ (.Y(_3341_),
    .A(net83),
    .B(_3771_));
 sg13g2_o21ai_1 _7870_ (.B1(_3341_),
    .Y(_3342_),
    .A1(_3920_),
    .A2(net83));
 sg13g2_xnor2_1 _7871_ (.Y(_3343_),
    .A(_0033_),
    .B(_3342_));
 sg13g2_o21ai_1 _7872_ (.B1(net122),
    .Y(_3344_),
    .A1(\i_transform.image_y[0] ),
    .A2(_3212_));
 sg13g2_a21oi_1 _7873_ (.A1(_3213_),
    .A2(_3343_),
    .Y(_0228_),
    .B1(_3344_));
 sg13g2_a21oi_1 _7874_ (.A1(_1161_),
    .A2(net65),
    .Y(_3345_),
    .B1(_1189_));
 sg13g2_nor2_1 _7875_ (.A(net105),
    .B(_3345_),
    .Y(_0229_));
 sg13g2_a21oi_1 _7876_ (.A1(_1291_),
    .A2(net65),
    .Y(_3346_),
    .B1(_1319_));
 sg13g2_nor2_1 _7877_ (.A(_3218_),
    .B(_3346_),
    .Y(_0230_));
 sg13g2_a21oi_1 _7878_ (.A1(_1375_),
    .A2(net65),
    .Y(_3347_),
    .B1(_1403_));
 sg13g2_nor2_1 _7879_ (.A(_3218_),
    .B(_3347_),
    .Y(_0231_));
 sg13g2_xnor2_1 _7880_ (.Y(_3348_),
    .A(_0048_),
    .B(net91));
 sg13g2_inv_1 _7881_ (.Y(_3349_),
    .A(_3348_));
 sg13g2_o21ai_1 _7882_ (.B1(_1385_),
    .Y(_3350_),
    .A1(_1882_),
    .A2(net91));
 sg13g2_xnor2_1 _7883_ (.Y(_3351_),
    .A(_3349_),
    .B(_3350_));
 sg13g2_nand2_1 _7884_ (.Y(_3352_),
    .A(net91),
    .B(_1389_));
 sg13g2_nand2b_1 _7885_ (.Y(_3353_),
    .B(_3352_),
    .A_N(_1380_));
 sg13g2_inv_1 _7886_ (.Y(_3354_),
    .A(_3353_));
 sg13g2_xnor2_1 _7887_ (.Y(_3355_),
    .A(_1877_),
    .B(net91));
 sg13g2_a21oi_1 _7888_ (.A1(_3354_),
    .A2(_3355_),
    .Y(_3356_),
    .B1(net70));
 sg13g2_nor2_1 _7889_ (.A(_3355_),
    .B(_3354_),
    .Y(_3357_));
 sg13g2_inv_1 _7890_ (.Y(_3358_),
    .A(_3357_));
 sg13g2_nand2_1 _7891_ (.Y(_3359_),
    .A(_3356_),
    .B(_3358_));
 sg13g2_o21ai_1 _7892_ (.B1(_3359_),
    .Y(_3360_),
    .A1(net73),
    .A2(_3351_));
 sg13g2_nand2_1 _7893_ (.Y(_3361_),
    .A(_3360_),
    .B(net84));
 sg13g2_xnor2_1 _7894_ (.Y(_3362_),
    .A(_1877_),
    .B(net98));
 sg13g2_a21oi_1 _7895_ (.A1(_1389_),
    .A2(net98),
    .Y(_3363_),
    .B1(_1398_));
 sg13g2_xnor2_1 _7896_ (.Y(_3364_),
    .A(_3362_),
    .B(_3363_));
 sg13g2_a21oi_1 _7897_ (.A1(_3364_),
    .A2(_1640_),
    .Y(_3365_),
    .B1(_3653_));
 sg13g2_xnor2_1 _7898_ (.Y(_3366_),
    .A(_0048_),
    .B(net98));
 sg13g2_a22oi_1 _7899_ (.Y(_3367_),
    .B1(_1391_),
    .B2(_1394_),
    .A2(_0605_),
    .A1(_1375_));
 sg13g2_nor2_1 _7900_ (.A(_3366_),
    .B(_3367_),
    .Y(_3368_));
 sg13g2_and2_1 _7901_ (.A(_3367_),
    .B(_3366_),
    .X(_3369_));
 sg13g2_o21ai_1 _7902_ (.B1(_1628_),
    .Y(_3370_),
    .A1(_3368_),
    .A2(_3369_));
 sg13g2_a22oi_1 _7903_ (.Y(_3371_),
    .B1(_3365_),
    .B2(_3370_),
    .A2(net64),
    .A1(_1877_));
 sg13g2_a21oi_1 _7904_ (.A1(_3361_),
    .A2(_3371_),
    .Y(_0232_),
    .B1(net104));
 sg13g2_buf_1 _7905_ (.A(_0049_),
    .X(_3372_));
 sg13g2_xnor2_1 _7906_ (.Y(_3373_),
    .A(_3372_),
    .B(net86));
 sg13g2_a22oi_1 _7907_ (.Y(_3374_),
    .B1(_3349_),
    .B2(_3350_),
    .A2(net92),
    .A1(_1877_));
 sg13g2_nor2_1 _7908_ (.A(_3373_),
    .B(_3374_),
    .Y(_3375_));
 sg13g2_a21o_1 _7909_ (.A2(_3373_),
    .A1(_3374_),
    .B1(net73),
    .X(_3376_));
 sg13g2_inv_1 _7910_ (.Y(_3377_),
    .A(_0048_));
 sg13g2_nand2_1 _7911_ (.Y(_3378_),
    .A(net86),
    .B(_3377_));
 sg13g2_xnor2_1 _7912_ (.Y(_3379_),
    .A(_1879_),
    .B(_1376_));
 sg13g2_nand3_1 _7913_ (.B(_3378_),
    .C(_3379_),
    .A(_3358_),
    .Y(_3380_));
 sg13g2_inv_1 _7914_ (.Y(_3381_),
    .A(_3379_));
 sg13g2_nand2_1 _7915_ (.Y(_3382_),
    .A(_3357_),
    .B(_3381_));
 sg13g2_nor2_1 _7916_ (.A(_3378_),
    .B(_3379_),
    .Y(_3383_));
 sg13g2_nor2_1 _7917_ (.A(_3383_),
    .B(net74),
    .Y(_3384_));
 sg13g2_nand3_1 _7918_ (.B(_3382_),
    .C(_3384_),
    .A(_3380_),
    .Y(_3385_));
 sg13g2_o21ai_1 _7919_ (.B1(_3385_),
    .Y(_3386_),
    .A1(_3375_),
    .A2(_3376_));
 sg13g2_a22oi_1 _7920_ (.Y(_3387_),
    .B1(_0687_),
    .B2(_3386_),
    .A2(_3226_),
    .A1(_1879_));
 sg13g2_xnor2_1 _7921_ (.Y(_3388_),
    .A(_1879_),
    .B(_1390_));
 sg13g2_nor2_1 _7922_ (.A(_3362_),
    .B(_3363_),
    .Y(_3389_));
 sg13g2_a21oi_1 _7923_ (.A1(_3377_),
    .A2(net98),
    .Y(_3390_),
    .B1(_3389_));
 sg13g2_nor2_1 _7924_ (.A(_3388_),
    .B(_3390_),
    .Y(_3391_));
 sg13g2_a21oi_1 _7925_ (.A1(_3390_),
    .A2(_3388_),
    .Y(_3392_),
    .B1(_1628_));
 sg13g2_nor2b_1 _7926_ (.A(_3391_),
    .B_N(_3392_),
    .Y(_3393_));
 sg13g2_nor2_1 _7927_ (.A(_1878_),
    .B(net88),
    .Y(_3394_));
 sg13g2_xnor2_1 _7928_ (.Y(_3395_),
    .A(_3372_),
    .B(net88));
 sg13g2_o21ai_1 _7929_ (.B1(_3395_),
    .Y(_3396_),
    .A1(_3394_),
    .A2(_3368_));
 sg13g2_inv_1 _7930_ (.Y(_3397_),
    .A(_3368_));
 sg13g2_inv_1 _7931_ (.Y(_3398_),
    .A(_3394_));
 sg13g2_nand3b_1 _7932_ (.B(_3397_),
    .C(_3398_),
    .Y(_3399_),
    .A_N(_3395_));
 sg13g2_a21oi_1 _7933_ (.A1(_3396_),
    .A2(_3399_),
    .Y(_3400_),
    .B1(_1640_));
 sg13g2_o21ai_1 _7934_ (.B1(_0689_),
    .Y(_3401_),
    .A1(_3393_),
    .A2(_3400_));
 sg13g2_a21oi_1 _7935_ (.A1(_3387_),
    .A2(_3401_),
    .Y(_0233_),
    .B1(net104));
 sg13g2_a21oi_1 _7936_ (.A1(_1879_),
    .A2(net92),
    .Y(_3402_),
    .B1(_3375_));
 sg13g2_xnor2_1 _7937_ (.Y(_3403_),
    .A(_0050_),
    .B(_3241_));
 sg13g2_o21ai_1 _7938_ (.B1(net70),
    .Y(_3404_),
    .A1(_3403_),
    .A2(_3402_));
 sg13g2_a21oi_1 _7939_ (.A1(_3402_),
    .A2(_3403_),
    .Y(_3405_),
    .B1(_3404_));
 sg13g2_inv_1 _7940_ (.Y(_3406_),
    .A(_3372_));
 sg13g2_a21oi_1 _7941_ (.A1(_3406_),
    .A2(_3241_),
    .Y(_3407_),
    .B1(_3383_));
 sg13g2_xnor2_1 _7942_ (.Y(_3408_),
    .A(net179),
    .B(net86));
 sg13g2_a21oi_1 _7943_ (.A1(_3382_),
    .A2(_3407_),
    .Y(_3409_),
    .B1(_3408_));
 sg13g2_nand3_1 _7944_ (.B(_3407_),
    .C(_3408_),
    .A(_3382_),
    .Y(_3410_));
 sg13g2_nand2b_1 _7945_ (.Y(_3411_),
    .B(_3410_),
    .A_N(_3409_));
 sg13g2_nor2_1 _7946_ (.A(net70),
    .B(_3411_),
    .Y(_3412_));
 sg13g2_o21ai_1 _7947_ (.B1(net84),
    .Y(_3413_),
    .A1(_3405_),
    .A2(_3412_));
 sg13g2_a21oi_1 _7948_ (.A1(_3406_),
    .A2(net88),
    .Y(_3414_),
    .B1(_3391_));
 sg13g2_xnor2_1 _7949_ (.Y(_3415_),
    .A(net179),
    .B(_3248_));
 sg13g2_o21ai_1 _7950_ (.B1(net62),
    .Y(_3416_),
    .A1(_3415_),
    .A2(_3414_));
 sg13g2_a21oi_1 _7951_ (.A1(_3414_),
    .A2(_3415_),
    .Y(_3417_),
    .B1(_3416_));
 sg13g2_a22oi_1 _7952_ (.Y(_3418_),
    .B1(_3372_),
    .B2(_3394_),
    .A2(_1879_),
    .A1(net114));
 sg13g2_o21ai_1 _7953_ (.B1(_3418_),
    .Y(_3419_),
    .A1(_3395_),
    .A2(_3397_));
 sg13g2_xor2_1 _7954_ (.B(_3248_),
    .A(_0050_),
    .X(_3420_));
 sg13g2_a21oi_1 _7955_ (.A1(_3419_),
    .A2(_3420_),
    .Y(_3421_),
    .B1(net62));
 sg13g2_o21ai_1 _7956_ (.B1(_3421_),
    .Y(_3422_),
    .A1(_3419_),
    .A2(_3420_));
 sg13g2_nand2b_1 _7957_ (.Y(_3423_),
    .B(_3422_),
    .A_N(_3417_));
 sg13g2_a22oi_1 _7958_ (.Y(_3424_),
    .B1(_3652_),
    .B2(_3423_),
    .A2(_3226_),
    .A1(net179));
 sg13g2_a21oi_1 _7959_ (.A1(_3413_),
    .A2(_3424_),
    .Y(_0234_),
    .B1(_3228_));
 sg13g2_xnor2_1 _7960_ (.Y(_3425_),
    .A(_3822_),
    .B(_3823_));
 sg13g2_nor2_1 _7961_ (.A(_3927_),
    .B(_3926_),
    .Y(_3426_));
 sg13g2_nor2_1 _7962_ (.A(net81),
    .B(_3426_),
    .Y(_3427_));
 sg13g2_a22oi_1 _7963_ (.Y(_3428_),
    .B1(_3928_),
    .B2(_3427_),
    .A2(net81),
    .A1(_3425_));
 sg13g2_o21ai_1 _7964_ (.B1(net122),
    .Y(_3429_),
    .A1(\i_transform.image_y[1] ),
    .A2(net57));
 sg13g2_a21oi_1 _7965_ (.A1(_3428_),
    .A2(net56),
    .Y(_0235_),
    .B1(_3429_));
 sg13g2_xor2_1 _7966_ (.B(_3825_),
    .A(_3819_),
    .X(_3430_));
 sg13g2_nor2_1 _7967_ (.A(_3930_),
    .B(_3929_),
    .Y(_3431_));
 sg13g2_nor2_1 _7968_ (.A(net81),
    .B(_3431_),
    .Y(_3432_));
 sg13g2_a22oi_1 _7969_ (.Y(_3433_),
    .B1(_3931_),
    .B2(_3432_),
    .A2(net81),
    .A1(_3430_));
 sg13g2_o21ai_1 _7970_ (.B1(_1713_),
    .Y(_3434_),
    .A1(\i_transform.image_y[2] ),
    .A2(net57));
 sg13g2_a21oi_1 _7971_ (.A1(_3433_),
    .A2(net56),
    .Y(_0236_),
    .B1(_3434_));
 sg13g2_nor2_1 _7972_ (.A(net82),
    .B(_0862_),
    .Y(_3435_));
 sg13g2_nand2_1 _7973_ (.Y(_3436_),
    .A(_3827_),
    .B(_0861_));
 sg13g2_nand2_1 _7974_ (.Y(_3437_),
    .A(_3932_),
    .B(_3941_));
 sg13g2_nor2_1 _7975_ (.A(_3941_),
    .B(_3932_),
    .Y(_3438_));
 sg13g2_nor2_1 _7976_ (.A(net81),
    .B(_3438_),
    .Y(_3439_));
 sg13g2_a22oi_1 _7977_ (.Y(_3440_),
    .B1(_3437_),
    .B2(_3439_),
    .A2(_3436_),
    .A1(_3435_));
 sg13g2_o21ai_1 _7978_ (.B1(net122),
    .Y(_3441_),
    .A1(\i_transform.image_y[3] ),
    .A2(net57));
 sg13g2_a21oi_1 _7979_ (.A1(_3440_),
    .A2(_3213_),
    .Y(_0237_),
    .B1(_3441_));
 sg13g2_nor2_1 _7980_ (.A(net82),
    .B(_0864_),
    .Y(_3442_));
 sg13g2_nand2_1 _7981_ (.Y(_3443_),
    .A(_0863_),
    .B(_3853_));
 sg13g2_nand2_1 _7982_ (.Y(_3444_),
    .A(_3437_),
    .B(_0290_));
 sg13g2_nand2_1 _7983_ (.Y(_3445_),
    .A(_3444_),
    .B(_0288_));
 sg13g2_inv_1 _7984_ (.Y(_3446_),
    .A(_3444_));
 sg13g2_a21oi_1 _7985_ (.A1(_3446_),
    .A2(_0287_),
    .Y(_3447_),
    .B1(net81));
 sg13g2_a22oi_1 _7986_ (.Y(_3448_),
    .B1(_3445_),
    .B2(_3447_),
    .A2(_3443_),
    .A1(_3442_));
 sg13g2_o21ai_1 _7987_ (.B1(_1713_),
    .Y(_3449_),
    .A1(\i_transform.image_y[4] ),
    .A2(net57));
 sg13g2_a21oi_1 _7988_ (.A1(_3448_),
    .A2(net56),
    .Y(_0238_),
    .B1(_3449_));
 sg13g2_nand2_1 _7989_ (.Y(_3450_),
    .A(_3445_),
    .B(_0292_));
 sg13g2_xnor2_1 _7990_ (.Y(_3451_),
    .A(_3955_),
    .B(_3450_));
 sg13g2_xnor2_1 _7991_ (.Y(_3452_),
    .A(_3764_),
    .B(_3920_));
 sg13g2_o21ai_1 _7992_ (.B1(net84),
    .Y(_3453_),
    .A1(_3452_),
    .A2(net73));
 sg13g2_a21o_1 _7993_ (.A2(net73),
    .A1(_3451_),
    .B1(_3453_),
    .X(_3454_));
 sg13g2_xnor2_1 _7994_ (.Y(_3455_),
    .A(_3765_),
    .B(_3753_));
 sg13g2_a21oi_1 _7995_ (.A1(net59),
    .A2(_3455_),
    .Y(_3456_),
    .B1(net63));
 sg13g2_xnor2_1 _7996_ (.Y(_3457_),
    .A(_3863_),
    .B(_0865_));
 sg13g2_nand2_1 _7997_ (.Y(_3458_),
    .A(_3457_),
    .B(net58));
 sg13g2_a22oi_1 _7998_ (.Y(_3459_),
    .B1(_3456_),
    .B2(_3458_),
    .A2(net64),
    .A1(_3855_));
 sg13g2_a21oi_1 _7999_ (.A1(_3454_),
    .A2(_3459_),
    .Y(_0239_),
    .B1(net112));
 sg13g2_nor2_1 _8000_ (.A(_3775_),
    .B(net58),
    .Y(_3460_));
 sg13g2_nand2_1 _8001_ (.Y(_3461_),
    .A(_3774_),
    .B(_3772_));
 sg13g2_xnor2_1 _8002_ (.Y(_3462_),
    .A(_3879_),
    .B(_0867_));
 sg13g2_a22oi_1 _8003_ (.Y(_3463_),
    .B1(net58),
    .B2(_3462_),
    .A2(_3461_),
    .A1(_3460_));
 sg13g2_nor2_1 _8004_ (.A(_3880_),
    .B(_1372_),
    .Y(_3464_));
 sg13g2_a22oi_1 _8005_ (.Y(_3465_),
    .B1(_3955_),
    .B2(_3450_),
    .A2(net75),
    .A1(_3855_));
 sg13g2_o21ai_1 _8006_ (.B1(net77),
    .Y(_3466_),
    .A1(_3942_),
    .A2(_3465_));
 sg13g2_a21o_1 _8007_ (.A2(_3465_),
    .A1(_3942_),
    .B1(_3466_),
    .X(_3467_));
 sg13g2_o21ai_1 _8008_ (.B1(_0325_),
    .Y(_3468_),
    .A1(_0323_),
    .A2(_0322_));
 sg13g2_a21oi_1 _8009_ (.A1(_3467_),
    .A2(_3468_),
    .Y(_3469_),
    .B1(net81));
 sg13g2_o21ai_1 _8010_ (.B1(net132),
    .Y(_3470_),
    .A1(_3464_),
    .A2(_3469_));
 sg13g2_o21ai_1 _8011_ (.B1(_3470_),
    .Y(_0240_),
    .A1(_1639_),
    .A2(_3463_));
 sg13g2_nand2_1 _8012_ (.Y(_3471_),
    .A(_3888_),
    .B(_0335_));
 sg13g2_a21oi_1 _8013_ (.A1(_3889_),
    .A2(net65),
    .Y(_3472_),
    .B1(_3471_));
 sg13g2_nor2_1 _8014_ (.A(net105),
    .B(_3472_),
    .Y(_0241_));
 sg13g2_nor2_1 _8015_ (.A(_1052_),
    .B(_0586_),
    .Y(_3473_));
 sg13g2_nor3_1 _8016_ (.A(_0855_),
    .B(_3473_),
    .C(_0880_),
    .Y(_3474_));
 sg13g2_nor2_1 _8017_ (.A(net105),
    .B(_3474_),
    .Y(_0242_));
 sg13g2_a21oi_1 _8018_ (.A1(_1067_),
    .A2(_3222_),
    .Y(_3475_),
    .B1(_1078_));
 sg13g2_nor2_1 _8019_ (.A(_3228_),
    .B(_3475_),
    .Y(_0243_));
 sg13g2_nor2_1 _8020_ (.A(net8),
    .B(_3478_),
    .Y(_3476_));
 sg13g2_o21ai_1 _8021_ (.B1(net169),
    .Y(_3477_),
    .A1(orient),
    .A2(_3476_));
 sg13g2_a21oi_1 _8022_ (.A1(_3891_),
    .A2(_3476_),
    .Y(_0284_),
    .B1(_3477_));
 sg13g2_nor2_2 _8023_ (.A(\i_delta_sigma.acc[13] ),
    .B(net4),
    .Y(pdm_out));
 sg13g2_dfrbp_1 _8024_ (.CLK(clknet_leaf_28_clk),
    .RESET_B(net190),
    .D(_0069_),
    .Q_N(_0052_),
    .Q(\i_collision.i_coll_table.in[3] ));
 sg13g2_buf_2 clkbuf_leaf_0_clk (.A(clknet_3_1__leaf_clk),
    .X(clknet_leaf_0_clk));
 sg13g2_buf_1 _8026_ (.A(net191),
    .X(uio_oe[0]));
 sg13g2_buf_1 _8027_ (.A(net192),
    .X(uio_oe[1]));
 sg13g2_buf_1 _8028_ (.A(net193),
    .X(uio_oe[2]));
 sg13g2_buf_1 _8029_ (.A(net194),
    .X(uio_oe[3]));
 sg13g2_buf_1 _8030_ (.A(net195),
    .X(uio_oe[4]));
 sg13g2_buf_1 _8031_ (.A(net196),
    .X(uio_oe[5]));
 sg13g2_buf_1 _8032_ (.A(net197),
    .X(uio_oe[6]));
 sg13g2_buf_1 _8033_ (.A(net198),
    .X(uio_oe[7]));
 sg13g2_buf_1 _8034_ (.A(pdm_out),
    .X(net9));
 sg13g2_buf_1 _8035_ (.A(pdm_out),
    .X(net10));
 sg13g2_buf_1 _8036_ (.A(pdm_out),
    .X(net11));
 sg13g2_buf_1 _8037_ (.A(pdm_out),
    .X(net12));
 sg13g2_buf_1 _8038_ (.A(pdm_out),
    .X(net13));
 sg13g2_buf_1 _8039_ (.A(pdm_out),
    .X(net14));
 sg13g2_buf_1 _8040_ (.A(pdm_out),
    .X(net15));
 sg13g2_buf_1 _8041_ (.A(pdm_out),
    .X(net16));
 sg13g2_buf_1 _8042_ (.A(\i_vga_beam.vsync ),
    .X(net20));
 sg13g2_buf_1 _8043_ (.A(hsync),
    .X(net24));
 sg13g2_dfrbp_1 \bitmap_pixel$_DFF_P_  (.CLK(clknet_leaf_5_clk),
    .RESET_B(net199),
    .D(_0000_),
    .Q_N(_4111_),
    .Q(bitmap_pixel));
 sg13g2_dfrbp_1 \i_collision.imp[0]$_SDFFE_PN0P_  (.CLK(clknet_leaf_20_clk),
    .RESET_B(net200),
    .D(_0076_),
    .Q_N(_4110_),
    .Q(\collision_impact[0] ));
 sg13g2_dfrbp_1 \i_collision.imp[1]$_SDFFE_PN0P_  (.CLK(clknet_leaf_23_clk),
    .RESET_B(net201),
    .D(_0077_),
    .Q_N(_4109_),
    .Q(\collision_impact[1] ));
 sg13g2_dfrbp_1 \i_collision.vx[0]$_SDFFE_PN0P_  (.CLK(clknet_leaf_22_clk),
    .RESET_B(net202),
    .D(_0078_),
    .Q_N(_0009_),
    .Q(\i_collision.vx[0] ));
 sg13g2_dfrbp_1 \i_collision.vx[1]$_SDFFE_PN1P_  (.CLK(clknet_leaf_23_clk),
    .RESET_B(net203),
    .D(_0079_),
    .Q_N(_4108_),
    .Q(\i_collision.vx[1] ));
 sg13g2_dfrbp_1 \i_collision.vx[2]$_SDFFE_PN0P_  (.CLK(clknet_leaf_22_clk),
    .RESET_B(net204),
    .D(_0080_),
    .Q_N(_4107_),
    .Q(\i_collision.vx[2] ));
 sg13g2_dfrbp_1 \i_collision.vy[0]$_SDFFE_PN1P_  (.CLK(clknet_leaf_22_clk),
    .RESET_B(net205),
    .D(_0081_),
    .Q_N(_0008_),
    .Q(\i_collision.vy[0] ));
 sg13g2_dfrbp_1 \i_collision.vy[1]$_SDFFE_PN0P_  (.CLK(clknet_leaf_23_clk),
    .RESET_B(net206),
    .D(_0082_),
    .Q_N(_4106_),
    .Q(\i_collision.vy[1] ));
 sg13g2_dfrbp_1 \i_collision.vy[2]$_SDFFE_PN0P_  (.CLK(clknet_leaf_22_clk),
    .RESET_B(net207),
    .D(_0083_),
    .Q_N(_4105_),
    .Q(\i_collision.vy[2] ));
 sg13g2_dfrbp_1 \i_collision.w[1]$_SDFFE_PN0P_  (.CLK(clknet_leaf_28_clk),
    .RESET_B(net208),
    .D(_0084_),
    .Q_N(_0053_),
    .Q(\i_collision.i_coll_table.in[4] ));
 sg13g2_dfrbp_1 \i_collision.w[2]$_SDFFE_PN0P_  (.CLK(clknet_leaf_30_clk),
    .RESET_B(net209),
    .D(_0085_),
    .Q_N(_0068_),
    .Q(\i_collision.i_coll_table.in[5] ));
 sg13g2_dfrbp_1 \i_colors.blue[0]$_SDFFE_PN1P_  (.CLK(clknet_leaf_12_clk),
    .RESET_B(net210),
    .D(_0086_),
    .Q_N(_4104_),
    .Q(\capsule_color[0] ));
 sg13g2_dfrbp_1 \i_colors.blue[1]$_SDFFE_PN0P_  (.CLK(clknet_leaf_10_clk),
    .RESET_B(net211),
    .D(_0087_),
    .Q_N(_4118_),
    .Q(\capsule_color[1] ));
 sg13g2_dfrbp_1 \i_colors.channel[0]$_DFF_P_  (.CLK(clknet_leaf_13_clk),
    .RESET_B(net212),
    .D(_0001_),
    .Q_N(_4119_),
    .Q(\i_colors.channel[0] ));
 sg13g2_dfrbp_1 \i_colors.channel[1]$_DFF_P_  (.CLK(clknet_leaf_12_clk),
    .RESET_B(net213),
    .D(_0002_),
    .Q_N(_0010_),
    .Q(\i_colors.channel[1] ));
 sg13g2_dfrbp_1 \i_colors.channel[2]$_DFF_P_  (.CLK(clknet_leaf_12_clk),
    .RESET_B(net214),
    .D(_0003_),
    .Q_N(_4103_),
    .Q(\i_colors.channel[2] ));
 sg13g2_dfrbp_1 \i_colors.green[0]$_SDFFE_PN1P_  (.CLK(clknet_leaf_12_clk),
    .RESET_B(net215),
    .D(_0088_),
    .Q_N(_4102_),
    .Q(\capsule_color[2] ));
 sg13g2_dfrbp_1 \i_colors.green[1]$_SDFFE_PN0P_  (.CLK(clknet_leaf_11_clk),
    .RESET_B(net216),
    .D(_0089_),
    .Q_N(_4101_),
    .Q(\capsule_color[3] ));
 sg13g2_dfrbp_1 \i_colors.red[0]$_SDFFE_PN1P_  (.CLK(clknet_leaf_12_clk),
    .RESET_B(net217),
    .D(_0090_),
    .Q_N(_4100_),
    .Q(\capsule_color[4] ));
 sg13g2_dfrbp_1 \i_colors.red[1]$_SDFFE_PN1P_  (.CLK(clknet_leaf_12_clk),
    .RESET_B(net218),
    .D(_0091_),
    .Q_N(_4099_),
    .Q(\capsule_color[5] ));
 sg13g2_dfrbp_1 \i_delta_sigma.acc[0]$_SDFF_PN0_  (.CLK(clknet_leaf_15_clk),
    .RESET_B(net219),
    .D(_0092_),
    .Q_N(_4098_),
    .Q(\i_delta_sigma.acc[0] ));
 sg13g2_dfrbp_1 \i_delta_sigma.acc[10]$_SDFF_PN0_  (.CLK(clknet_leaf_19_clk),
    .RESET_B(net220),
    .D(_0093_),
    .Q_N(_4097_),
    .Q(\i_delta_sigma.acc[10] ));
 sg13g2_dfrbp_1 \i_delta_sigma.acc[11]$_SDFF_PN0_  (.CLK(clknet_leaf_19_clk),
    .RESET_B(net221),
    .D(_0094_),
    .Q_N(_4096_),
    .Q(\i_delta_sigma.acc[11] ));
 sg13g2_dfrbp_1 \i_delta_sigma.acc[12]$_SDFF_PN0_  (.CLK(clknet_leaf_19_clk),
    .RESET_B(net222),
    .D(_0095_),
    .Q_N(_4095_),
    .Q(\i_delta_sigma.acc[12] ));
 sg13g2_dfrbp_1 \i_delta_sigma.acc[13]$_SDFF_PN0_  (.CLK(clknet_leaf_17_clk),
    .RESET_B(net223),
    .D(_0096_),
    .Q_N(_0055_),
    .Q(\i_delta_sigma.acc[13] ));
 sg13g2_dfrbp_1 \i_delta_sigma.acc[1]$_SDFF_PN0_  (.CLK(clknet_leaf_16_clk),
    .RESET_B(net224),
    .D(_0097_),
    .Q_N(_4094_),
    .Q(\i_delta_sigma.acc[1] ));
 sg13g2_dfrbp_1 \i_delta_sigma.acc[2]$_SDFF_PN0_  (.CLK(clknet_leaf_16_clk),
    .RESET_B(net225),
    .D(_0098_),
    .Q_N(_4093_),
    .Q(\i_delta_sigma.acc[2] ));
 sg13g2_dfrbp_1 \i_delta_sigma.acc[3]$_SDFF_PN0_  (.CLK(clknet_leaf_17_clk),
    .RESET_B(net226),
    .D(_0099_),
    .Q_N(_4092_),
    .Q(\i_delta_sigma.acc[3] ));
 sg13g2_dfrbp_1 \i_delta_sigma.acc[4]$_SDFF_PN0_  (.CLK(clknet_leaf_16_clk),
    .RESET_B(net227),
    .D(_0100_),
    .Q_N(_4091_),
    .Q(\i_delta_sigma.acc[4] ));
 sg13g2_dfrbp_1 \i_delta_sigma.acc[5]$_SDFF_PN0_  (.CLK(clknet_leaf_18_clk),
    .RESET_B(net228),
    .D(_0101_),
    .Q_N(_4090_),
    .Q(\i_delta_sigma.acc[5] ));
 sg13g2_dfrbp_1 \i_delta_sigma.acc[6]$_SDFF_PN0_  (.CLK(clknet_leaf_23_clk),
    .RESET_B(net229),
    .D(_0102_),
    .Q_N(_4089_),
    .Q(\i_delta_sigma.acc[6] ));
 sg13g2_dfrbp_1 \i_delta_sigma.acc[7]$_SDFF_PN0_  (.CLK(clknet_leaf_23_clk),
    .RESET_B(net230),
    .D(_0103_),
    .Q_N(_4088_),
    .Q(\i_delta_sigma.acc[7] ));
 sg13g2_dfrbp_1 \i_delta_sigma.acc[8]$_SDFF_PN0_  (.CLK(clknet_leaf_19_clk),
    .RESET_B(net231),
    .D(_0104_),
    .Q_N(_4087_),
    .Q(\i_delta_sigma.acc[8] ));
 sg13g2_dfrbp_1 \i_delta_sigma.acc[9]$_SDFF_PN0_  (.CLK(clknet_leaf_19_clk),
    .RESET_B(net232),
    .D(_0105_),
    .Q_N(_4086_),
    .Q(\i_delta_sigma.acc[9] ));
 sg13g2_dfrbp_1 \i_kinematics.center_x[0]$_SDFFE_PP0P_  (.CLK(clknet_leaf_21_clk),
    .RESET_B(net233),
    .D(_0106_),
    .Q_N(_4085_),
    .Q(\center_x[0] ));
 sg13g2_dfrbp_1 \i_kinematics.center_x[1]$_SDFFE_PP0P_  (.CLK(clknet_leaf_21_clk),
    .RESET_B(net234),
    .D(_0107_),
    .Q_N(_4084_),
    .Q(\center_x[1] ));
 sg13g2_dfrbp_1 \i_kinematics.center_x[2]$_SDFFE_PP0P_  (.CLK(clknet_leaf_21_clk),
    .RESET_B(net235),
    .D(_0108_),
    .Q_N(_4083_),
    .Q(\center_x[2] ));
 sg13g2_dfrbp_1 \i_kinematics.center_x[3]$_SDFFE_PP0P_  (.CLK(clknet_leaf_20_clk),
    .RESET_B(net236),
    .D(_0109_),
    .Q_N(_4082_),
    .Q(\center_x[3] ));
 sg13g2_dfrbp_1 \i_kinematics.center_x[4]$_SDFFE_PP0P_  (.CLK(clknet_leaf_20_clk),
    .RESET_B(net237),
    .D(_0110_),
    .Q_N(_4081_),
    .Q(\center_x[4] ));
 sg13g2_dfrbp_1 \i_kinematics.center_x[5]$_SDFFE_PP0P_  (.CLK(clknet_leaf_20_clk),
    .RESET_B(net238),
    .D(_0111_),
    .Q_N(_4080_),
    .Q(\center_x[5] ));
 sg13g2_dfrbp_1 \i_kinematics.center_x[6]$_SDFFE_PP1P_  (.CLK(clknet_leaf_21_clk),
    .RESET_B(net239),
    .D(_0112_),
    .Q_N(_4079_),
    .Q(\center_x[6] ));
 sg13g2_dfrbp_1 \i_kinematics.center_x[7]$_SDFFE_PP0P_  (.CLK(clknet_leaf_9_clk),
    .RESET_B(net240),
    .D(_0113_),
    .Q_N(_4078_),
    .Q(\center_x[7] ));
 sg13g2_dfrbp_1 \i_kinematics.center_x[8]$_SDFFE_PP1P_  (.CLK(clknet_leaf_21_clk),
    .RESET_B(net241),
    .D(_0114_),
    .Q_N(_4077_),
    .Q(\center_x[8] ));
 sg13g2_dfrbp_1 \i_kinematics.center_x[9]$_SDFFE_PP0P_  (.CLK(clknet_leaf_9_clk),
    .RESET_B(net242),
    .D(_0115_),
    .Q_N(_4076_),
    .Q(\center_x[9] ));
 sg13g2_dfrbp_1 \i_kinematics.center_x_lo[0]$_SDFFE_PP0P_  (.CLK(clknet_leaf_22_clk),
    .RESET_B(net243),
    .D(_0116_),
    .Q_N(_4075_),
    .Q(\i_kinematics.center_x_lo[0] ));
 sg13g2_dfrbp_1 \i_kinematics.center_x_lo[1]$_SDFFE_PP0P_  (.CLK(clknet_leaf_24_clk),
    .RESET_B(net244),
    .D(_0117_),
    .Q_N(_4074_),
    .Q(\i_kinematics.center_x_lo[1] ));
 sg13g2_dfrbp_1 \i_kinematics.center_y[0]$_SDFFE_PP0P_  (.CLK(clknet_leaf_23_clk),
    .RESET_B(net245),
    .D(_0118_),
    .Q_N(_4073_),
    .Q(\center_y[0] ));
 sg13g2_dfrbp_1 \i_kinematics.center_y[1]$_SDFFE_PP0P_  (.CLK(clknet_leaf_22_clk),
    .RESET_B(net246),
    .D(_0119_),
    .Q_N(_4072_),
    .Q(\center_y[1] ));
 sg13g2_dfrbp_1 \i_kinematics.center_y[2]$_SDFFE_PP0P_  (.CLK(clknet_leaf_22_clk),
    .RESET_B(net247),
    .D(_0120_),
    .Q_N(_4071_),
    .Q(\center_y[2] ));
 sg13g2_dfrbp_1 \i_kinematics.center_y[3]$_SDFFE_PP0P_  (.CLK(clknet_leaf_31_clk),
    .RESET_B(net248),
    .D(_0121_),
    .Q_N(_4070_),
    .Q(\center_y[3] ));
 sg13g2_dfrbp_1 \i_kinematics.center_y[4]$_SDFFE_PP1P_  (.CLK(clknet_leaf_31_clk),
    .RESET_B(net249),
    .D(_0122_),
    .Q_N(_4069_),
    .Q(\center_y[4] ));
 sg13g2_dfrbp_1 \i_kinematics.center_y[5]$_SDFFE_PP1P_  (.CLK(clknet_leaf_32_clk),
    .RESET_B(net250),
    .D(_0123_),
    .Q_N(_4068_),
    .Q(\center_y[5] ));
 sg13g2_dfrbp_1 \i_kinematics.center_y[6]$_SDFFE_PP1P_  (.CLK(clknet_leaf_31_clk),
    .RESET_B(net251),
    .D(_0124_),
    .Q_N(_4067_),
    .Q(\center_y[6] ));
 sg13g2_dfrbp_1 \i_kinematics.center_y[7]$_SDFFE_PP1P_  (.CLK(clknet_leaf_32_clk),
    .RESET_B(net252),
    .D(_0125_),
    .Q_N(_4066_),
    .Q(\center_y[7] ));
 sg13g2_dfrbp_1 \i_kinematics.center_y[8]$_SDFFE_PP0P_  (.CLK(clknet_leaf_31_clk),
    .RESET_B(net253),
    .D(_0126_),
    .Q_N(_4065_),
    .Q(\center_y[8] ));
 sg13g2_dfrbp_1 \i_kinematics.center_y[9]$_SDFFE_PP0P_  (.CLK(clknet_leaf_32_clk),
    .RESET_B(net254),
    .D(_0127_),
    .Q_N(_4064_),
    .Q(\center_y[9] ));
 sg13g2_dfrbp_1 \i_kinematics.center_y_lo[0]$_SDFFE_PP0P_  (.CLK(clknet_leaf_31_clk),
    .RESET_B(net255),
    .D(_0128_),
    .Q_N(_4063_),
    .Q(\i_kinematics.center_y_lo[0] ));
 sg13g2_dfrbp_1 \i_kinematics.center_y_lo[1]$_SDFFE_PP0P_  (.CLK(clknet_leaf_31_clk),
    .RESET_B(net256),
    .D(_0129_),
    .Q_N(_4062_),
    .Q(\i_kinematics.center_y_lo[1] ));
 sg13g2_dfrbp_1 \i_kinematics.phi[0]$_SDFFE_PP0P_  (.CLK(clknet_leaf_30_clk),
    .RESET_B(net257),
    .D(_0130_),
    .Q_N(_4061_),
    .Q(\i_kinematics.phi[0] ));
 sg13g2_dfrbp_1 \i_kinematics.phi[10]$_SDFFE_PP0P_  (.CLK(clknet_leaf_30_clk),
    .RESET_B(net258),
    .D(_0131_),
    .Q_N(_4060_),
    .Q(\i_kinematics.phi[10] ));
 sg13g2_dfrbp_1 \i_kinematics.phi[1]$_SDFFE_PP0P_  (.CLK(clknet_leaf_28_clk),
    .RESET_B(net259),
    .D(_0132_),
    .Q_N(_4059_),
    .Q(\i_kinematics.phi[1] ));
 sg13g2_dfrbp_1 \i_kinematics.phi[2]$_SDFFE_PP0P_  (.CLK(clknet_leaf_28_clk),
    .RESET_B(net260),
    .D(_0133_),
    .Q_N(_4058_),
    .Q(\i_kinematics.phi[2] ));
 sg13g2_dfrbp_1 \i_kinematics.phi[3]$_SDFFE_PP0P_  (.CLK(clknet_leaf_29_clk),
    .RESET_B(net261),
    .D(_0134_),
    .Q_N(_4057_),
    .Q(\i_kinematics.phi[3] ));
 sg13g2_dfrbp_1 \i_kinematics.phi[4]$_SDFFE_PP0P_  (.CLK(clknet_leaf_29_clk),
    .RESET_B(net262),
    .D(_0135_),
    .Q_N(_4056_),
    .Q(\i_kinematics.phi[4] ));
 sg13g2_dfrbp_1 \i_kinematics.phi[5]$_SDFFE_PP0P_  (.CLK(clknet_leaf_29_clk),
    .RESET_B(net263),
    .D(_0136_),
    .Q_N(_4055_),
    .Q(\i_kinematics.phi[5] ));
 sg13g2_dfrbp_1 \i_kinematics.phi[6]$_SDFFE_PP0P_  (.CLK(clknet_leaf_29_clk),
    .RESET_B(net264),
    .D(_0137_),
    .Q_N(_4054_),
    .Q(\i_kinematics.phi[6] ));
 sg13g2_dfrbp_1 \i_kinematics.phi[7]$_SDFFE_PP0P_  (.CLK(clknet_leaf_29_clk),
    .RESET_B(net265),
    .D(_0138_),
    .Q_N(_4053_),
    .Q(\i_kinematics.phi[7] ));
 sg13g2_dfrbp_1 \i_kinematics.phi[8]$_SDFFE_PP1P_  (.CLK(clknet_leaf_30_clk),
    .RESET_B(net266),
    .D(_0139_),
    .Q_N(_0051_),
    .Q(\i_collision.i_coll_table.in[1] ));
 sg13g2_dfrbp_1 \i_kinematics.phi[9]$_SDFFE_PP0P_  (.CLK(clknet_leaf_30_clk),
    .RESET_B(net267),
    .D(_0140_),
    .Q_N(_4052_),
    .Q(\i_collision.phi[1] ));
 sg13g2_dfrbp_1 \i_orchestrator.handle_impact$_SDFF_PP0_  (.CLK(clknet_leaf_14_clk),
    .RESET_B(net268),
    .D(_0141_),
    .Q_N(_4051_),
    .Q(handle_impact));
 sg13g2_dfrbp_1 \i_orchestrator.hit_bottom$_SDFFE_PN0P_  (.CLK(clknet_leaf_9_clk),
    .RESET_B(net269),
    .D(_0142_),
    .Q_N(_0005_),
    .Q(\i_orchestrator.hit_bottom ));
 sg13g2_dfrbp_1 \i_orchestrator.hit_left$_SDFFE_PN0P_  (.CLK(clknet_leaf_10_clk),
    .RESET_B(net270),
    .D(_0143_),
    .Q_N(_0012_),
    .Q(\i_orchestrator.hit_left ));
 sg13g2_dfrbp_1 \i_orchestrator.hit_priority[0]$_SDFFE_PN0P_  (.CLK(clknet_leaf_13_clk),
    .RESET_B(net271),
    .D(_0144_),
    .Q_N(_0066_),
    .Q(\i_orchestrator.hit_priority[0] ));
 sg13g2_dfrbp_1 \i_orchestrator.hit_priority[1]$_SDFFE_PN0P_  (.CLK(clknet_leaf_13_clk),
    .RESET_B(net272),
    .D(_0145_),
    .Q_N(_4050_),
    .Q(\i_orchestrator.hit_priority[1] ));
 sg13g2_dfrbp_1 \i_orchestrator.hit_right$_SDFFE_PN0P_  (.CLK(clknet_leaf_12_clk),
    .RESET_B(net273),
    .D(_0146_),
    .Q_N(_0057_),
    .Q(\i_orchestrator.hit_right ));
 sg13g2_dfrbp_1 \i_orchestrator.hit_top$_SDFFE_PN0P_  (.CLK(clknet_leaf_10_clk),
    .RESET_B(net274),
    .D(_0147_),
    .Q_N(_0056_),
    .Q(\i_orchestrator.hit_top ));
 sg13g2_dfrbp_1 \i_orchestrator.lfsr[0]$_SDFFE_PN1P_  (.CLK(clknet_leaf_28_clk),
    .RESET_B(net275),
    .D(_0148_),
    .Q_N(_0054_),
    .Q(\i_collision.i_coll_table.in[0] ));
 sg13g2_dfrbp_1 \i_orchestrator.lfsr[1]$_SDFFE_PN1P_  (.CLK(clknet_leaf_13_clk),
    .RESET_B(net276),
    .D(_0149_),
    .Q_N(_4049_),
    .Q(\i_orchestrator.lfsr[1] ));
 sg13g2_dfrbp_1 \i_orchestrator.lfsr[2]$_SDFFE_PN1P_  (.CLK(clknet_leaf_13_clk),
    .RESET_B(net277),
    .D(_0150_),
    .Q_N(_4048_),
    .Q(\i_orchestrator.lfsr[2] ));
 sg13g2_dfrbp_1 \i_orchestrator.lfsr[3]$_SDFFE_PN1P_  (.CLK(clknet_leaf_15_clk),
    .RESET_B(net278),
    .D(_0151_),
    .Q_N(_4047_),
    .Q(\i_orchestrator.lfsr[3] ));
 sg13g2_dfrbp_1 \i_orchestrator.lfsr[4]$_SDFFE_PN1P_  (.CLK(clknet_leaf_14_clk),
    .RESET_B(net279),
    .D(_0152_),
    .Q_N(_4046_),
    .Q(\i_orchestrator.lfsr[4] ));
 sg13g2_dfrbp_1 \i_orchestrator.lfsr[5]$_SDFFE_PN1P_  (.CLK(clknet_leaf_14_clk),
    .RESET_B(net280),
    .D(_0153_),
    .Q_N(_4045_),
    .Q(\i_orchestrator.lfsr[5] ));
 sg13g2_dfrbp_1 \i_orchestrator.lfsr[6]$_SDFFE_PN1P_  (.CLK(clknet_leaf_14_clk),
    .RESET_B(net281),
    .D(_0154_),
    .Q_N(_4044_),
    .Q(\i_orchestrator.lfsr[6] ));
 sg13g2_dfrbp_1 \i_orchestrator.lfsr[7]$_SDFFE_PN1P_  (.CLK(clknet_leaf_13_clk),
    .RESET_B(net282),
    .D(_0155_),
    .Q_N(_4043_),
    .Q(\i_orchestrator.lfsr[7] ));
 sg13g2_dfrbp_1 \i_orchestrator.lfsr[8]$_SDFFE_PN1P_  (.CLK(clknet_leaf_12_clk),
    .RESET_B(net283),
    .D(_0156_),
    .Q_N(_0011_),
    .Q(\color_entropy[0] ));
 sg13g2_dfrbp_1 \i_orchestrator.lfsr[9]$_SDFFE_PN1P_  (.CLK(clknet_leaf_13_clk),
    .RESET_B(net284),
    .D(_0157_),
    .Q_N(_4042_),
    .Q(\color_entropy[1] ));
 sg13g2_dfrbp_1 \i_orchestrator.mirror_collision$_SDFF_PN0_  (.CLK(clknet_leaf_20_clk),
    .RESET_B(net285),
    .D(_0158_),
    .Q_N(_4041_),
    .Q(\i_collision.mirror ));
 sg13g2_dfrbp_1 \i_orchestrator.rotate_collision$_SDFF_PN0_  (.CLK(clknet_leaf_20_clk),
    .RESET_B(net286),
    .D(_0159_),
    .Q_N(_4040_),
    .Q(\i_collision.rotate ));
 sg13g2_dfrbp_1 \i_orchestrator.sample_counter[0]$_SDFF_PN0_  (.CLK(clknet_leaf_14_clk),
    .RESET_B(net287),
    .D(_0160_),
    .Q_N(_0065_),
    .Q(\i_orchestrator.sample_counter[0] ));
 sg13g2_dfrbp_1 \i_orchestrator.sample_counter[1]$_SDFF_PN0_  (.CLK(clknet_leaf_14_clk),
    .RESET_B(net288),
    .D(_0161_),
    .Q_N(_4039_),
    .Q(\i_orchestrator.sample_counter[1] ));
 sg13g2_dfrbp_1 \i_orchestrator.sample_counter[2]$_SDFF_PN0_  (.CLK(clknet_leaf_14_clk),
    .RESET_B(net289),
    .D(_0162_),
    .Q_N(_4038_),
    .Q(\i_orchestrator.sample_counter[2] ));
 sg13g2_dfrbp_1 \i_orchestrator.sample_counter[3]$_SDFF_PN0_  (.CLK(clknet_leaf_15_clk),
    .RESET_B(net290),
    .D(_0163_),
    .Q_N(_4037_),
    .Q(\i_orchestrator.sample_counter[3] ));
 sg13g2_dfrbp_1 \i_orchestrator.sample_counter[4]$_SDFF_PN0_  (.CLK(clknet_leaf_15_clk),
    .RESET_B(net291),
    .D(_0164_),
    .Q_N(_4036_),
    .Q(\i_orchestrator.sample_counter[4] ));
 sg13g2_dfrbp_1 \i_orchestrator.sample_counter[5]$_SDFF_PN0_  (.CLK(clknet_leaf_15_clk),
    .RESET_B(net292),
    .D(_0165_),
    .Q_N(_4035_),
    .Q(\i_orchestrator.sample_counter[5] ));
 sg13g2_dfrbp_1 \i_orchestrator.sample_counter[6]$_SDFF_PN0_  (.CLK(clknet_leaf_15_clk),
    .RESET_B(net293),
    .D(_0166_),
    .Q_N(_4034_),
    .Q(\i_orchestrator.sample_counter[6] ));
 sg13g2_dfrbp_1 \i_orchestrator.sample_counter[7]$_SDFF_PN0_  (.CLK(clknet_leaf_15_clk),
    .RESET_B(net294),
    .D(_0167_),
    .Q_N(_4033_),
    .Q(\i_orchestrator.sample_counter[7] ));
 sg13g2_dfrbp_1 \i_orchestrator.sample_counter[8]$_SDFF_PN0_  (.CLK(clknet_leaf_14_clk),
    .RESET_B(net295),
    .D(_0168_),
    .Q_N(_4032_),
    .Q(\i_orchestrator.sample_counter[8] ));
 sg13g2_dfrbp_1 \i_orchestrator.sample_counter[9]$_SDFF_PN0_  (.CLK(clknet_leaf_15_clk),
    .RESET_B(net296),
    .D(_0169_),
    .Q_N(_4031_),
    .Q(\i_orchestrator.sample_counter[9] ));
 sg13g2_dfrbp_1 \i_orchestrator.tension[1]$_SDFFE_PN0P_  (.CLK(clknet_leaf_17_clk),
    .RESET_B(net297),
    .D(_0170_),
    .Q_N(_4030_),
    .Q(\i_orchestrator.tension[1] ));
 sg13g2_dfrbp_1 \i_orchestrator.tension[2]$_SDFFE_PN0P_  (.CLK(clknet_leaf_17_clk),
    .RESET_B(net298),
    .D(_0171_),
    .Q_N(_4029_),
    .Q(\i_orchestrator.tension[2] ));
 sg13g2_dfrbp_1 \i_orchestrator.tension[3]$_SDFFE_PN0P_  (.CLK(clknet_leaf_16_clk),
    .RESET_B(net299),
    .D(_0172_),
    .Q_N(_4028_),
    .Q(\i_orchestrator.tension[3] ));
 sg13g2_dfrbp_1 \i_orchestrator.trigger_debounce$_SDFFE_PN0P_  (.CLK(clknet_leaf_9_clk),
    .RESET_B(net300),
    .D(_0173_),
    .Q_N(_0004_),
    .Q(\i_orchestrator.trigger_debounce ));
 sg13g2_dfrbp_1 \i_orchestrator.trigger_resonator[0]$_SDFF_PP0_  (.CLK(clknet_leaf_17_clk),
    .RESET_B(net301),
    .D(_0174_),
    .Q_N(_4027_),
    .Q(\i_orchestrator.trigger_resonator[0] ));
 sg13g2_dfrbp_1 \i_orchestrator.trigger_resonator[1]$_SDFF_PP0_  (.CLK(clknet_leaf_17_clk),
    .RESET_B(net302),
    .D(_0175_),
    .Q_N(_4026_),
    .Q(\i_orchestrator.trigger_resonator[1] ));
 sg13g2_dfrbp_1 \i_orchestrator.update_collision$_SDFF_PN0_  (.CLK(clknet_leaf_20_clk),
    .RESET_B(net303),
    .D(_0176_),
    .Q_N(_4025_),
    .Q(\i_collision.update ));
 sg13g2_dfrbp_1 \i_orchestrator.update_kinematics$_SDFF_PP0_  (.CLK(clknet_leaf_9_clk),
    .RESET_B(net304),
    .D(_0177_),
    .Q_N(_4024_),
    .Q(\i_kinematics.update ));
 sg13g2_dfrbp_1 \i_orchestrator.update_resonator$_SDFF_PN0_  (.CLK(clknet_leaf_16_clk),
    .RESET_B(net305),
    .D(_0178_),
    .Q_N(_0061_),
    .Q(\i_orchestrator.update_resonator ));
 sg13g2_dfrbp_1 \i_orchestrator.update_transform$_SDFF_PP0_  (.CLK(clknet_leaf_10_clk),
    .RESET_B(net306),
    .D(_0179_),
    .Q_N(_4023_),
    .Q(\i_orchestrator.update_transform ));
 sg13g2_dfrbp_1 \i_resonator.counter[0]$_SDFFE_PP0P_  (.CLK(clknet_leaf_16_clk),
    .RESET_B(net307),
    .D(_0180_),
    .Q_N(_4022_),
    .Q(\i_resonator.counter[0] ));
 sg13g2_dfrbp_1 \i_resonator.counter[1]$_SDFFE_PP0P_  (.CLK(clknet_leaf_17_clk),
    .RESET_B(net308),
    .D(_0181_),
    .Q_N(_0062_),
    .Q(\i_resonator.counter[1] ));
 sg13g2_dfrbp_1 \i_resonator.counter[2]$_SDFFE_PP0P_  (.CLK(clknet_leaf_16_clk),
    .RESET_B(net309),
    .D(_0182_),
    .Q_N(_4021_),
    .Q(\i_resonator.counter[2] ));
 sg13g2_dfrbp_1 \i_resonator.counter[3]$_SDFFE_PP0P_  (.CLK(clknet_leaf_16_clk),
    .RESET_B(net310),
    .D(_0183_),
    .Q_N(_4020_),
    .Q(\i_resonator.counter[3] ));
 sg13g2_dfrbp_1 \i_resonator.v[0]$_SDFFE_PP0P_  (.CLK(clknet_leaf_25_clk),
    .RESET_B(net311),
    .D(_0184_),
    .Q_N(_0039_),
    .Q(\i_resonator.v[0] ));
 sg13g2_dfrbp_1 \i_resonator.v[10]$_SDFFE_PP0P_  (.CLK(clknet_leaf_27_clk),
    .RESET_B(net312),
    .D(_0185_),
    .Q_N(_4019_),
    .Q(\i_resonator.v[10] ));
 sg13g2_dfrbp_1 \i_resonator.v[11]$_SDFFE_PP0P_  (.CLK(clknet_leaf_25_clk),
    .RESET_B(net313),
    .D(_0186_),
    .Q_N(_0040_),
    .Q(\i_resonator.v[11] ));
 sg13g2_dfrbp_1 \i_resonator.v[12]$_SDFFE_PP0P_  (.CLK(clknet_leaf_24_clk),
    .RESET_B(net314),
    .D(_0187_),
    .Q_N(_4018_),
    .Q(\i_resonator.v[12] ));
 sg13g2_dfrbp_1 \i_resonator.v[13]$_SDFFE_PP0P_  (.CLK(clknet_leaf_25_clk),
    .RESET_B(net315),
    .D(_0188_),
    .Q_N(_0042_),
    .Q(\i_resonator.v[13] ));
 sg13g2_dfrbp_1 \i_resonator.v[14]$_SDFFE_PP0P_  (.CLK(clknet_leaf_25_clk),
    .RESET_B(net316),
    .D(_0189_),
    .Q_N(_4017_),
    .Q(\i_resonator.v[14] ));
 sg13g2_dfrbp_1 \i_resonator.v[15]$_SDFFE_PP0P_  (.CLK(clknet_leaf_25_clk),
    .RESET_B(net317),
    .D(_0190_),
    .Q_N(_0043_),
    .Q(\i_resonator.v[15] ));
 sg13g2_dfrbp_1 \i_resonator.v[1]$_SDFFE_PP0P_  (.CLK(clknet_leaf_24_clk),
    .RESET_B(net318),
    .D(_0191_),
    .Q_N(_4016_),
    .Q(\i_resonator.v[1] ));
 sg13g2_dfrbp_1 \i_resonator.v[2]$_SDFFE_PP0P_  (.CLK(clknet_leaf_23_clk),
    .RESET_B(net319),
    .D(_0192_),
    .Q_N(_4015_),
    .Q(\i_resonator.v[2] ));
 sg13g2_dfrbp_1 \i_resonator.v[3]$_SDFFE_PP0P_  (.CLK(clknet_leaf_23_clk),
    .RESET_B(net320),
    .D(_0193_),
    .Q_N(_4014_),
    .Q(\i_resonator.v[3] ));
 sg13g2_dfrbp_1 \i_resonator.v[4]$_SDFFE_PP0P_  (.CLK(clknet_leaf_26_clk),
    .RESET_B(net321),
    .D(_0194_),
    .Q_N(_4013_),
    .Q(\i_resonator.v[4] ));
 sg13g2_dfrbp_1 \i_resonator.v[5]$_SDFFE_PP0P_  (.CLK(clknet_leaf_26_clk),
    .RESET_B(net322),
    .D(_0195_),
    .Q_N(_4012_),
    .Q(\i_resonator.v[5] ));
 sg13g2_dfrbp_1 \i_resonator.v[6]$_SDFFE_PP0P_  (.CLK(clknet_leaf_27_clk),
    .RESET_B(net323),
    .D(_0196_),
    .Q_N(_4011_),
    .Q(\i_resonator.v[6] ));
 sg13g2_dfrbp_1 \i_resonator.v[7]$_SDFFE_PP0P_  (.CLK(clknet_leaf_27_clk),
    .RESET_B(net324),
    .D(_0197_),
    .Q_N(_4010_),
    .Q(\i_resonator.v[7] ));
 sg13g2_dfrbp_1 \i_resonator.v[8]$_SDFFE_PP0P_  (.CLK(clknet_leaf_27_clk),
    .RESET_B(net325),
    .D(_0198_),
    .Q_N(_4009_),
    .Q(\i_resonator.v[8] ));
 sg13g2_dfrbp_1 \i_resonator.v[9]$_SDFFE_PP0P_  (.CLK(clknet_leaf_27_clk),
    .RESET_B(net326),
    .D(_0199_),
    .Q_N(_0041_),
    .Q(\i_resonator.v[9] ));
 sg13g2_dfrbp_1 \i_resonator.x[0]$_SDFFE_PP0P_  (.CLK(clknet_leaf_18_clk),
    .RESET_B(net327),
    .D(_0200_),
    .Q_N(_4008_),
    .Q(\i_delta_sigma.sample[0] ));
 sg13g2_dfrbp_1 \i_resonator.x[10]$_SDFFE_PP0P_  (.CLK(clknet_leaf_18_clk),
    .RESET_B(net328),
    .D(_0201_),
    .Q_N(_4007_),
    .Q(\i_delta_sigma.sample[10] ));
 sg13g2_dfrbp_1 \i_resonator.x[11]$_SDFFE_PP0P_  (.CLK(clknet_leaf_25_clk),
    .RESET_B(net329),
    .D(_0202_),
    .Q_N(_4006_),
    .Q(\i_delta_sigma.sample[11] ));
 sg13g2_dfrbp_1 \i_resonator.x[1]$_SDFFE_PP0P_  (.CLK(clknet_leaf_18_clk),
    .RESET_B(net330),
    .D(_0203_),
    .Q_N(_4005_),
    .Q(\i_delta_sigma.sample[1] ));
 sg13g2_dfrbp_1 \i_resonator.x[2]$_SDFFE_PP0P_  (.CLK(clknet_leaf_18_clk),
    .RESET_B(net331),
    .D(_0204_),
    .Q_N(_4004_),
    .Q(\i_delta_sigma.sample[2] ));
 sg13g2_dfrbp_1 \i_resonator.x[3]$_SDFFE_PP0P_  (.CLK(clknet_leaf_18_clk),
    .RESET_B(net332),
    .D(_0205_),
    .Q_N(_4003_),
    .Q(\i_delta_sigma.sample[3] ));
 sg13g2_dfrbp_1 \i_resonator.x[4]$_SDFFE_PP0P_  (.CLK(clknet_leaf_18_clk),
    .RESET_B(net333),
    .D(_0206_),
    .Q_N(_4002_),
    .Q(\i_delta_sigma.sample[4] ));
 sg13g2_dfrbp_1 \i_resonator.x[5]$_SDFFE_PP0P_  (.CLK(clknet_leaf_18_clk),
    .RESET_B(net334),
    .D(_0207_),
    .Q_N(_4001_),
    .Q(\i_delta_sigma.sample[5] ));
 sg13g2_dfrbp_1 \i_resonator.x[6]$_SDFFE_PP0P_  (.CLK(clknet_leaf_19_clk),
    .RESET_B(net335),
    .D(_0208_),
    .Q_N(_4000_),
    .Q(\i_delta_sigma.sample[6] ));
 sg13g2_dfrbp_1 \i_resonator.x[7]$_SDFFE_PP0P_  (.CLK(clknet_leaf_19_clk),
    .RESET_B(net336),
    .D(_0209_),
    .Q_N(_3999_),
    .Q(\i_delta_sigma.sample[7] ));
 sg13g2_dfrbp_1 \i_resonator.x[8]$_SDFFE_PP0P_  (.CLK(clknet_leaf_19_clk),
    .RESET_B(net337),
    .D(_0210_),
    .Q_N(_3998_),
    .Q(\i_delta_sigma.sample[8] ));
 sg13g2_dfrbp_1 \i_resonator.x[9]$_SDFFE_PP0P_  (.CLK(clknet_leaf_17_clk),
    .RESET_B(net338),
    .D(_0211_),
    .Q_N(_3997_),
    .Q(\i_delta_sigma.sample[9] ));
 sg13g2_dfrbp_1 \i_transform.image_x[0]$_SDFFE_PN0P_  (.CLK(clknet_leaf_34_clk),
    .RESET_B(net339),
    .D(_0212_),
    .Q_N(_0018_),
    .Q(\i_transform.image_x[0] ));
 sg13g2_dfrbp_1 \i_transform.image_x[10]$_SDFFE_PN0N_  (.CLK(clknet_leaf_0_clk),
    .RESET_B(net340),
    .D(_0213_),
    .Q_N(_0022_),
    .Q(\i_bitmap.in[3] ));
 sg13g2_dfrbp_1 \i_transform.image_x[11]$_SDFFE_PN0N_  (.CLK(clknet_leaf_36_clk),
    .RESET_B(net341),
    .D(_0214_),
    .Q_N(_0023_),
    .Q(\i_bitmap.in[4] ));
 sg13g2_dfrbp_1 \i_transform.image_x[12]$_SDFFE_PN0N_  (.CLK(clknet_leaf_0_clk),
    .RESET_B(net342),
    .D(_0215_),
    .Q_N(_0024_),
    .Q(\i_bitmap.in[5] ));
 sg13g2_dfrbp_1 \i_transform.image_x[13]$_SDFFE_PN0N_  (.CLK(clknet_leaf_4_clk),
    .RESET_B(net343),
    .D(_0216_),
    .Q_N(_0025_),
    .Q(\i_bitmap.in[6] ));
 sg13g2_dfrbp_1 \i_transform.image_x[14]$_SDFFE_PN0N_  (.CLK(clknet_leaf_4_clk),
    .RESET_B(net344),
    .D(_0217_),
    .Q_N(_0046_),
    .Q(\i_capsule.tf_x[8] ));
 sg13g2_dfrbp_1 \i_transform.image_x[15]$_SDFFE_PN0N_  (.CLK(clknet_leaf_4_clk),
    .RESET_B(net345),
    .D(_0218_),
    .Q_N(_0063_),
    .Q(\i_capsule.tf_x[9] ));
 sg13g2_dfrbp_1 \i_transform.image_x[1]$_SDFFE_PN0P_  (.CLK(clknet_leaf_34_clk),
    .RESET_B(net346),
    .D(_0219_),
    .Q_N(_3996_),
    .Q(\i_transform.image_x[1] ));
 sg13g2_dfrbp_1 \i_transform.image_x[2]$_SDFFE_PN0P_  (.CLK(clknet_leaf_34_clk),
    .RESET_B(net347),
    .D(_0220_),
    .Q_N(_0017_),
    .Q(\i_transform.image_x[2] ));
 sg13g2_dfrbp_1 \i_transform.image_x[3]$_SDFFE_PN0P_  (.CLK(clknet_leaf_35_clk),
    .RESET_B(net348),
    .D(_0221_),
    .Q_N(_0016_),
    .Q(\i_transform.image_x[3] ));
 sg13g2_dfrbp_1 \i_transform.image_x[4]$_SDFFE_PN0P_  (.CLK(clknet_leaf_35_clk),
    .RESET_B(net349),
    .D(_0222_),
    .Q_N(_0015_),
    .Q(\i_transform.image_x[4] ));
 sg13g2_dfrbp_1 \i_transform.image_x[5]$_SDFFE_PN0N_  (.CLK(clknet_leaf_34_clk),
    .RESET_B(net350),
    .D(_0223_),
    .Q_N(_0014_),
    .Q(\i_transform.image_x[5] ));
 sg13g2_dfrbp_1 \i_transform.image_x[6]$_SDFFE_PN0N_  (.CLK(clknet_leaf_36_clk),
    .RESET_B(net351),
    .D(_0224_),
    .Q_N(_0020_),
    .Q(\i_capsule.tf_x[0] ));
 sg13g2_dfrbp_1 \i_transform.image_x[7]$_SDFFE_PN0N_  (.CLK(clknet_leaf_36_clk),
    .RESET_B(net352),
    .D(_0225_),
    .Q_N(_0019_),
    .Q(\i_bitmap.in[0] ));
 sg13g2_dfrbp_1 \i_transform.image_x[8]$_SDFFE_PN0N_  (.CLK(clknet_leaf_0_clk),
    .RESET_B(net353),
    .D(_0226_),
    .Q_N(_0013_),
    .Q(\i_bitmap.in[1] ));
 sg13g2_dfrbp_1 \i_transform.image_x[9]$_SDFFE_PN0N_  (.CLK(clknet_leaf_0_clk),
    .RESET_B(net354),
    .D(_0227_),
    .Q_N(_0021_),
    .Q(\i_bitmap.in[2] ));
 sg13g2_dfrbp_1 \i_transform.image_y[0]$_SDFFE_PN0P_  (.CLK(clknet_leaf_29_clk),
    .RESET_B(net355),
    .D(_0228_),
    .Q_N(_0033_),
    .Q(\i_transform.image_y[0] ));
 sg13g2_dfrbp_1 \i_transform.image_y[10]$_SDFFE_PN0N_  (.CLK(clknet_leaf_1_clk),
    .RESET_B(net356),
    .D(_0229_),
    .Q_N(_0036_),
    .Q(\i_bitmap.in[10] ));
 sg13g2_dfrbp_1 \i_transform.image_y[11]$_SDFFE_PN0N_  (.CLK(clknet_leaf_1_clk),
    .RESET_B(net357),
    .D(_0230_),
    .Q_N(_0037_),
    .Q(\i_bitmap.in[11] ));
 sg13g2_dfrbp_1 \i_transform.image_y[12]$_SDFFE_PN0N_  (.CLK(clknet_leaf_2_clk),
    .RESET_B(net358),
    .D(_0231_),
    .Q_N(_0038_),
    .Q(\i_bitmap.in[12] ));
 sg13g2_dfrbp_1 \i_transform.image_y[13]$_SDFFE_PN0N_  (.CLK(clknet_leaf_3_clk),
    .RESET_B(net359),
    .D(_0232_),
    .Q_N(_0048_),
    .Q(\i_capsule.tf_y[7] ));
 sg13g2_dfrbp_1 \i_transform.image_y[14]$_SDFFE_PN0N_  (.CLK(clknet_leaf_3_clk),
    .RESET_B(net360),
    .D(_0233_),
    .Q_N(_0049_),
    .Q(\i_capsule.tf_y[8] ));
 sg13g2_dfrbp_1 \i_transform.image_y[15]$_SDFFE_PN0N_  (.CLK(clknet_leaf_2_clk),
    .RESET_B(net361),
    .D(_0234_),
    .Q_N(_0050_),
    .Q(\i_capsule.tf_y[9] ));
 sg13g2_dfrbp_1 \i_transform.image_y[1]$_SDFFE_PN0P_  (.CLK(clknet_leaf_30_clk),
    .RESET_B(net362),
    .D(_0235_),
    .Q_N(_0032_),
    .Q(\i_transform.image_y[1] ));
 sg13g2_dfrbp_1 \i_transform.image_y[2]$_SDFFE_PN0P_  (.CLK(clknet_leaf_30_clk),
    .RESET_B(net363),
    .D(_0236_),
    .Q_N(_0031_),
    .Q(\i_transform.image_y[2] ));
 sg13g2_dfrbp_1 \i_transform.image_y[3]$_SDFFE_PN0P_  (.CLK(clknet_leaf_33_clk),
    .RESET_B(net364),
    .D(_0237_),
    .Q_N(_0030_),
    .Q(\i_transform.image_y[3] ));
 sg13g2_dfrbp_1 \i_transform.image_y[4]$_SDFFE_PN0P_  (.CLK(clknet_leaf_34_clk),
    .RESET_B(net365),
    .D(_0238_),
    .Q_N(_0029_),
    .Q(\i_transform.image_y[4] ));
 sg13g2_dfrbp_1 \i_transform.image_y[5]$_SDFFE_PN0N_  (.CLK(clknet_leaf_33_clk),
    .RESET_B(net366),
    .D(_0239_),
    .Q_N(_0028_),
    .Q(\i_transform.image_y[5] ));
 sg13g2_dfrbp_1 \i_transform.image_y[6]$_SDFFE_PN0N_  (.CLK(clknet_leaf_33_clk),
    .RESET_B(net367),
    .D(_0240_),
    .Q_N(_0027_),
    .Q(\i_capsule.tf_y[0] ));
 sg13g2_dfrbp_1 \i_transform.image_y[7]$_SDFFE_PN0N_  (.CLK(clknet_leaf_32_clk),
    .RESET_B(net368),
    .D(_0241_),
    .Q_N(_0026_),
    .Q(\i_bitmap.in[7] ));
 sg13g2_dfrbp_1 \i_transform.image_y[8]$_SDFFE_PN0N_  (.CLK(clknet_leaf_1_clk),
    .RESET_B(net369),
    .D(_0242_),
    .Q_N(_0034_),
    .Q(\i_bitmap.in[8] ));
 sg13g2_dfrbp_1 \i_transform.image_y[9]$_SDFFE_PN0N_  (.CLK(clknet_leaf_2_clk),
    .RESET_B(net370),
    .D(_0243_),
    .Q_N(_0035_),
    .Q(\i_bitmap.in[9] ));
 sg13g2_dfrbp_1 \i_transform.track_x[0]$_DFFE_PP_  (.CLK(clknet_leaf_2_clk),
    .RESET_B(net371),
    .D(_0244_),
    .Q_N(_0047_),
    .Q(\i_transform.track_x[0] ));
 sg13g2_dfrbp_1 \i_transform.track_x[1]$_DFFE_PP_  (.CLK(clknet_leaf_7_clk),
    .RESET_B(net372),
    .D(_0245_),
    .Q_N(_3995_),
    .Q(\i_transform.track_x[1] ));
 sg13g2_dfrbp_1 \i_transform.track_x[2]$_DFFE_PP_  (.CLK(clknet_leaf_2_clk),
    .RESET_B(net373),
    .D(_0246_),
    .Q_N(_3994_),
    .Q(\i_transform.track_x[2] ));
 sg13g2_dfrbp_1 \i_transform.track_x[3]$_DFFE_PP_  (.CLK(clknet_leaf_7_clk),
    .RESET_B(net374),
    .D(_0247_),
    .Q_N(_3993_),
    .Q(\i_transform.track_x[3] ));
 sg13g2_dfrbp_1 \i_transform.track_x[4]$_DFFE_PP_  (.CLK(clknet_leaf_7_clk),
    .RESET_B(net375),
    .D(_0248_),
    .Q_N(_3992_),
    .Q(\i_transform.track_x[4] ));
 sg13g2_dfrbp_1 \i_transform.track_x[5]$_DFFE_PP_  (.CLK(clknet_leaf_7_clk),
    .RESET_B(net376),
    .D(_0249_),
    .Q_N(_0044_),
    .Q(\i_transform.track_x[5] ));
 sg13g2_dfrbp_1 \i_transform.track_x[6]$_DFFE_PP_  (.CLK(clknet_leaf_7_clk),
    .RESET_B(net377),
    .D(_0250_),
    .Q_N(_3991_),
    .Q(\i_transform.track_x[6] ));
 sg13g2_dfrbp_1 \i_transform.track_x[7]$_DFFE_PP_  (.CLK(clknet_leaf_7_clk),
    .RESET_B(net378),
    .D(_0251_),
    .Q_N(_3990_),
    .Q(\i_transform.track_x[7] ));
 sg13g2_dfrbp_1 \i_transform.track_x[8]$_DFFE_PP_  (.CLK(clknet_leaf_7_clk),
    .RESET_B(net379),
    .D(_0252_),
    .Q_N(_3989_),
    .Q(\i_transform.track_x[8] ));
 sg13g2_dfrbp_1 \i_transform.track_x[9]$_DFFE_PP_  (.CLK(clknet_leaf_7_clk),
    .RESET_B(net380),
    .D(_0253_),
    .Q_N(_3988_),
    .Q(\i_transform.track_x[9] ));
 sg13g2_dfrbp_1 \i_transform.track_y[0]$_DFFE_PP_  (.CLK(clknet_leaf_32_clk),
    .RESET_B(net381),
    .D(_0254_),
    .Q_N(_0045_),
    .Q(\i_transform.track_y[0] ));
 sg13g2_dfrbp_1 \i_transform.track_y[1]$_DFFE_PP_  (.CLK(clknet_leaf_21_clk),
    .RESET_B(net382),
    .D(_0255_),
    .Q_N(_3987_),
    .Q(\i_transform.track_y[1] ));
 sg13g2_dfrbp_1 \i_transform.track_y[2]$_DFFE_PP_  (.CLK(clknet_leaf_21_clk),
    .RESET_B(net383),
    .D(_0256_),
    .Q_N(_3986_),
    .Q(\i_transform.track_y[2] ));
 sg13g2_dfrbp_1 \i_transform.track_y[3]$_DFFE_PP_  (.CLK(clknet_leaf_8_clk),
    .RESET_B(net384),
    .D(_0257_),
    .Q_N(_0058_),
    .Q(\i_transform.track_y[3] ));
 sg13g2_dfrbp_1 \i_transform.track_y[4]$_DFFE_PP_  (.CLK(clknet_leaf_21_clk),
    .RESET_B(net385),
    .D(_0258_),
    .Q_N(_3985_),
    .Q(\i_transform.track_y[4] ));
 sg13g2_dfrbp_1 \i_transform.track_y[5]$_DFFE_PP_  (.CLK(clknet_leaf_8_clk),
    .RESET_B(net386),
    .D(_0259_),
    .Q_N(_0060_),
    .Q(\i_transform.track_y[5] ));
 sg13g2_dfrbp_1 \i_transform.track_y[6]$_DFFE_PP_  (.CLK(clknet_leaf_31_clk),
    .RESET_B(net387),
    .D(_0260_),
    .Q_N(_3984_),
    .Q(\i_transform.track_y[6] ));
 sg13g2_dfrbp_1 \i_transform.track_y[7]$_DFFE_PP_  (.CLK(clknet_leaf_32_clk),
    .RESET_B(net388),
    .D(_0261_),
    .Q_N(_0059_),
    .Q(\i_transform.track_y[7] ));
 sg13g2_dfrbp_1 \i_transform.track_y[8]$_DFFE_PP_  (.CLK(clknet_leaf_32_clk),
    .RESET_B(net389),
    .D(_0262_),
    .Q_N(_3983_),
    .Q(\i_transform.track_y[8] ));
 sg13g2_dfrbp_1 \i_transform.track_y[9]$_DFFE_PP_  (.CLK(clknet_leaf_32_clk),
    .RESET_B(net390),
    .D(_0263_),
    .Q_N(_4120_),
    .Q(\i_transform.track_y[9] ));
 sg13g2_dfrbp_1 \i_vga_beam.hsync$_DFF_P_  (.CLK(clknet_leaf_6_clk),
    .RESET_B(net391),
    .D(_0006_),
    .Q_N(_4121_),
    .Q(hsync));
 sg13g2_dfrbp_1 \i_vga_beam.vsync$_DFF_P_  (.CLK(clknet_leaf_11_clk),
    .RESET_B(net392),
    .D(_0007_),
    .Q_N(_3982_),
    .Q(\i_vga_beam.vsync ));
 sg13g2_dfrbp_1 \i_vga_beam.x[0]$_SDFF_PP0_  (.CLK(clknet_leaf_5_clk),
    .RESET_B(net393),
    .D(_0264_),
    .Q_N(_0067_),
    .Q(\i_orchestrator.vga_x[0] ));
 sg13g2_dfrbp_1 \i_vga_beam.x[1]$_SDFF_PP0_  (.CLK(clknet_leaf_5_clk),
    .RESET_B(net394),
    .D(_0265_),
    .Q_N(_3981_),
    .Q(\i_orchestrator.vga_x[1] ));
 sg13g2_dfrbp_1 \i_vga_beam.x[2]$_SDFF_PP0_  (.CLK(clknet_leaf_5_clk),
    .RESET_B(net395),
    .D(_0266_),
    .Q_N(_3980_),
    .Q(\i_orchestrator.vga_x[2] ));
 sg13g2_dfrbp_1 \i_vga_beam.x[3]$_SDFF_PP0_  (.CLK(clknet_leaf_6_clk),
    .RESET_B(net396),
    .D(_0267_),
    .Q_N(_3979_),
    .Q(\i_orchestrator.vga_x[3] ));
 sg13g2_dfrbp_1 \i_vga_beam.x[4]$_SDFF_PP0_  (.CLK(clknet_leaf_6_clk),
    .RESET_B(net397),
    .D(_0268_),
    .Q_N(_3978_),
    .Q(\i_orchestrator.vga_x[4] ));
 sg13g2_dfrbp_1 \i_vga_beam.x[5]$_SDFF_PP0_  (.CLK(clknet_leaf_6_clk),
    .RESET_B(net398),
    .D(_0269_),
    .Q_N(_3977_),
    .Q(\i_orchestrator.vga_x[5] ));
 sg13g2_dfrbp_1 \i_vga_beam.x[6]$_SDFF_PP0_  (.CLK(clknet_leaf_5_clk),
    .RESET_B(net399),
    .D(_0270_),
    .Q_N(_3976_),
    .Q(\i_orchestrator.vga_x[6] ));
 sg13g2_dfrbp_1 \i_vga_beam.x[7]$_SDFF_PP0_  (.CLK(clknet_leaf_5_clk),
    .RESET_B(net400),
    .D(_0271_),
    .Q_N(_3975_),
    .Q(\i_orchestrator.vga_x[7] ));
 sg13g2_dfrbp_1 \i_vga_beam.x[8]$_SDFF_PP0_  (.CLK(clknet_leaf_5_clk),
    .RESET_B(net401),
    .D(_0272_),
    .Q_N(_3974_),
    .Q(\i_orchestrator.vga_x[8] ));
 sg13g2_dfrbp_1 \i_vga_beam.x[9]$_SDFF_PP0_  (.CLK(clknet_leaf_5_clk),
    .RESET_B(net402),
    .D(_0273_),
    .Q_N(_3973_),
    .Q(\i_orchestrator.vga_x[9] ));
 sg13g2_dfrbp_1 \i_vga_beam.y[0]$_SDFFCE_PP0P_  (.CLK(clknet_leaf_9_clk),
    .RESET_B(net403),
    .D(_0274_),
    .Q_N(_0064_),
    .Q(\i_orchestrator.vga_y[0] ));
 sg13g2_dfrbp_1 \i_vga_beam.y[1]$_SDFFCE_PP0P_  (.CLK(clknet_leaf_9_clk),
    .RESET_B(net404),
    .D(_0275_),
    .Q_N(_3972_),
    .Q(\i_orchestrator.vga_y[1] ));
 sg13g2_dfrbp_1 \i_vga_beam.y[2]$_SDFFCE_PP0P_  (.CLK(clknet_leaf_10_clk),
    .RESET_B(net405),
    .D(_0276_),
    .Q_N(_3971_),
    .Q(\i_orchestrator.vga_y[2] ));
 sg13g2_dfrbp_1 \i_vga_beam.y[3]$_SDFFCE_PP0P_  (.CLK(clknet_leaf_10_clk),
    .RESET_B(net406),
    .D(_0277_),
    .Q_N(_3970_),
    .Q(\i_orchestrator.vga_y[3] ));
 sg13g2_dfrbp_1 \i_vga_beam.y[4]$_SDFFCE_PP0P_  (.CLK(clknet_leaf_11_clk),
    .RESET_B(net407),
    .D(_0278_),
    .Q_N(_3969_),
    .Q(\i_orchestrator.vga_y[4] ));
 sg13g2_dfrbp_1 \i_vga_beam.y[5]$_SDFFCE_PP0P_  (.CLK(clknet_leaf_11_clk),
    .RESET_B(net408),
    .D(_0279_),
    .Q_N(_3968_),
    .Q(\i_orchestrator.vga_y[5] ));
 sg13g2_dfrbp_1 \i_vga_beam.y[6]$_SDFFCE_PP0P_  (.CLK(clknet_leaf_6_clk),
    .RESET_B(net409),
    .D(_0280_),
    .Q_N(_3967_),
    .Q(\i_orchestrator.vga_y[6] ));
 sg13g2_dfrbp_1 \i_vga_beam.y[7]$_SDFFCE_PP0P_  (.CLK(clknet_leaf_6_clk),
    .RESET_B(net410),
    .D(_0281_),
    .Q_N(_3966_),
    .Q(\i_orchestrator.vga_y[7] ));
 sg13g2_dfrbp_1 \i_vga_beam.y[8]$_SDFFCE_PP0P_  (.CLK(clknet_leaf_8_clk),
    .RESET_B(net411),
    .D(_0282_),
    .Q_N(_3965_),
    .Q(\i_orchestrator.vga_y[8] ));
 sg13g2_dfrbp_1 \i_vga_beam.y[9]$_SDFFCE_PP0P_  (.CLK(clknet_leaf_9_clk),
    .RESET_B(net412),
    .D(_0283_),
    .Q_N(_3964_),
    .Q(\i_orchestrator.vga_y[9] ));
 sg13g2_dfrbp_1 \orient$_SDFFE_PN0P_  (.CLK(clknet_leaf_20_clk),
    .RESET_B(net413),
    .D(_0284_),
    .Q_N(_3963_),
    .Q(orient));
 sg13g2_buf_1 input1 (.A(ui_in[0]),
    .X(net1));
 sg13g2_buf_1 input2 (.A(ui_in[1]),
    .X(net2));
 sg13g2_buf_1 input3 (.A(ui_in[2]),
    .X(net3));
 sg13g2_buf_1 input4 (.A(ui_in[3]),
    .X(net4));
 sg13g2_buf_1 input5 (.A(ui_in[4]),
    .X(net5));
 sg13g2_buf_1 input6 (.A(ui_in[5]),
    .X(net6));
 sg13g2_buf_1 input7 (.A(ui_in[6]),
    .X(net7));
 sg13g2_buf_1 input8 (.A(ui_in[7]),
    .X(net8));
 sg13g2_buf_1 output9 (.A(net9),
    .X(uio_out[0]));
 sg13g2_buf_1 output10 (.A(net10),
    .X(uio_out[1]));
 sg13g2_buf_1 output11 (.A(net11),
    .X(uio_out[2]));
 sg13g2_buf_1 output12 (.A(net12),
    .X(uio_out[3]));
 sg13g2_buf_1 output13 (.A(net13),
    .X(uio_out[4]));
 sg13g2_buf_1 output14 (.A(net14),
    .X(uio_out[5]));
 sg13g2_buf_1 output15 (.A(net15),
    .X(uio_out[6]));
 sg13g2_buf_1 output16 (.A(net16),
    .X(uio_out[7]));
 sg13g2_buf_1 output17 (.A(net17),
    .X(uo_out[0]));
 sg13g2_buf_1 output18 (.A(net18),
    .X(uo_out[1]));
 sg13g2_buf_1 output19 (.A(net19),
    .X(uo_out[2]));
 sg13g2_buf_1 output20 (.A(net20),
    .X(uo_out[3]));
 sg13g2_buf_1 output21 (.A(net21),
    .X(uo_out[4]));
 sg13g2_buf_1 output22 (.A(net22),
    .X(uo_out[5]));
 sg13g2_buf_1 output23 (.A(net23),
    .X(uo_out[6]));
 sg13g2_buf_1 output24 (.A(net24),
    .X(uo_out[7]));
 sg13g2_buf_2 fanout25 (.A(_0993_),
    .X(net25));
 sg13g2_buf_2 fanout26 (.A(_1248_),
    .X(net26));
 sg13g2_buf_2 fanout27 (.A(_0911_),
    .X(net27));
 sg13g2_buf_2 fanout28 (.A(_1119_),
    .X(net28));
 sg13g2_buf_2 fanout29 (.A(_1093_),
    .X(net29));
 sg13g2_buf_2 fanout30 (.A(_1032_),
    .X(net30));
 sg13g2_buf_2 fanout31 (.A(_0991_),
    .X(net31));
 sg13g2_buf_2 fanout32 (.A(_0834_),
    .X(net32));
 sg13g2_buf_2 fanout33 (.A(_1212_),
    .X(net33));
 sg13g2_buf_2 fanout34 (.A(_1149_),
    .X(net34));
 sg13g2_buf_2 fanout35 (.A(_1090_),
    .X(net35));
 sg13g2_buf_2 fanout36 (.A(_1022_),
    .X(net36));
 sg13g2_buf_2 fanout37 (.A(_0884_),
    .X(net37));
 sg13g2_buf_2 fanout38 (.A(_0592_),
    .X(net38));
 sg13g2_buf_2 fanout39 (.A(_1039_),
    .X(net39));
 sg13g2_buf_2 fanout40 (.A(_1029_),
    .X(net40));
 sg13g2_buf_2 fanout41 (.A(_1021_),
    .X(net41));
 sg13g2_buf_2 fanout42 (.A(_1014_),
    .X(net42));
 sg13g2_buf_2 fanout43 (.A(_1007_),
    .X(net43));
 sg13g2_buf_2 fanout44 (.A(_1002_),
    .X(net44));
 sg13g2_buf_2 fanout45 (.A(_0997_),
    .X(net45));
 sg13g2_buf_2 fanout46 (.A(_0939_),
    .X(net46));
 sg13g2_buf_2 fanout47 (.A(_0836_),
    .X(net47));
 sg13g2_buf_4 fanout48 (.X(net48),
    .A(_0832_));
 sg13g2_buf_2 fanout49 (.A(_1013_),
    .X(net49));
 sg13g2_buf_2 fanout50 (.A(_0917_),
    .X(net50));
 sg13g2_buf_2 fanout51 (.A(_0819_),
    .X(net51));
 sg13g2_buf_2 fanout52 (.A(_0701_),
    .X(net52));
 sg13g2_buf_2 fanout53 (.A(_0656_),
    .X(net53));
 sg13g2_buf_2 fanout54 (.A(_0346_),
    .X(net54));
 sg13g2_buf_2 fanout55 (.A(_0935_),
    .X(net55));
 sg13g2_buf_2 fanout56 (.A(_3213_),
    .X(net56));
 sg13g2_buf_2 fanout57 (.A(_3212_),
    .X(net57));
 sg13g2_buf_2 fanout58 (.A(_1628_),
    .X(net58));
 sg13g2_buf_2 fanout59 (.A(_1640_),
    .X(net59));
 sg13g2_buf_2 fanout60 (.A(_0501_),
    .X(net60));
 sg13g2_buf_2 fanout61 (.A(_2408_),
    .X(net61));
 sg13g2_buf_2 fanout62 (.A(_3885_),
    .X(net62));
 sg13g2_buf_2 fanout63 (.A(_3653_),
    .X(net63));
 sg13g2_buf_2 fanout64 (.A(_3226_),
    .X(net64));
 sg13g2_buf_2 fanout65 (.A(_3222_),
    .X(net65));
 sg13g2_buf_2 fanout66 (.A(_2671_),
    .X(net66));
 sg13g2_buf_2 fanout67 (.A(_2472_),
    .X(net67));
 sg13g2_buf_2 fanout68 (.A(_3669_),
    .X(net68));
 sg13g2_buf_2 fanout69 (.A(_2672_),
    .X(net69));
 sg13g2_buf_2 fanout70 (.A(_1664_),
    .X(net70));
 sg13g2_buf_2 fanout71 (.A(_0337_),
    .X(net71));
 sg13g2_buf_2 fanout72 (.A(_3852_),
    .X(net72));
 sg13g2_buf_2 fanout73 (.A(_1688_),
    .X(net73));
 sg13g2_buf_2 fanout74 (.A(_1066_),
    .X(net74));
 sg13g2_buf_2 fanout75 (.A(_3954_),
    .X(net75));
 sg13g2_buf_2 fanout76 (.A(_0332_),
    .X(net76));
 sg13g2_buf_2 fanout77 (.A(_0320_),
    .X(net77));
 sg13g2_buf_2 fanout78 (.A(_3940_),
    .X(net78));
 sg13g2_buf_2 fanout79 (.A(_3861_),
    .X(net79));
 sg13g2_buf_2 fanout80 (.A(_0319_),
    .X(net80));
 sg13g2_buf_2 fanout81 (.A(_1371_),
    .X(net81));
 sg13g2_buf_2 fanout82 (.A(_0687_),
    .X(net82));
 sg13g2_buf_2 fanout83 (.A(_0333_),
    .X(net83));
 sg13g2_buf_2 fanout84 (.A(_3592_),
    .X(net84));
 sg13g2_buf_2 fanout85 (.A(_3143_),
    .X(net85));
 sg13g2_buf_2 fanout86 (.A(_3241_),
    .X(net86));
 sg13g2_buf_2 fanout87 (.A(_3131_),
    .X(net87));
 sg13g2_buf_2 fanout88 (.A(_3248_),
    .X(net88));
 sg13g2_buf_2 fanout89 (.A(_2627_),
    .X(net89));
 sg13g2_buf_2 fanout90 (.A(_2299_),
    .X(net90));
 sg13g2_buf_2 fanout91 (.A(_1376_),
    .X(net91));
 sg13g2_buf_2 fanout92 (.A(_0750_),
    .X(net92));
 sg13g2_buf_2 fanout93 (.A(_2760_),
    .X(net93));
 sg13g2_buf_2 fanout94 (.A(_2298_),
    .X(net94));
 sg13g2_buf_2 fanout95 (.A(_1789_),
    .X(net95));
 sg13g2_buf_2 fanout96 (.A(_1737_),
    .X(net96));
 sg13g2_buf_2 fanout97 (.A(_1728_),
    .X(net97));
 sg13g2_buf_2 fanout98 (.A(_1390_),
    .X(net98));
 sg13g2_buf_2 fanout99 (.A(_3950_),
    .X(net99));
 sg13g2_buf_2 fanout100 (.A(_3897_),
    .X(net100));
 sg13g2_buf_2 fanout101 (.A(_3751_),
    .X(net101));
 sg13g2_buf_2 fanout102 (.A(_3596_),
    .X(net102));
 sg13g2_buf_2 fanout103 (.A(_3594_),
    .X(net103));
 sg13g2_buf_2 fanout104 (.A(_3228_),
    .X(net104));
 sg13g2_buf_2 fanout105 (.A(_3218_),
    .X(net105));
 sg13g2_buf_2 fanout106 (.A(_2796_),
    .X(net106));
 sg13g2_buf_2 fanout107 (.A(_2770_),
    .X(net107));
 sg13g2_buf_2 fanout108 (.A(_2414_),
    .X(net108));
 sg13g2_buf_2 fanout109 (.A(_2275_),
    .X(net109));
 sg13g2_buf_2 fanout110 (.A(_1775_),
    .X(net110));
 sg13g2_buf_2 fanout111 (.A(_1636_),
    .X(net111));
 sg13g2_buf_2 fanout112 (.A(_1600_),
    .X(net112));
 sg13g2_buf_2 fanout113 (.A(_0856_),
    .X(net113));
 sg13g2_buf_2 fanout114 (.A(_0605_),
    .X(net114));
 sg13g2_buf_2 fanout115 (.A(_3896_),
    .X(net115));
 sg13g2_buf_2 fanout116 (.A(_3741_),
    .X(net116));
 sg13g2_buf_2 fanout117 (.A(_2814_),
    .X(net117));
 sg13g2_buf_2 fanout118 (.A(_2789_),
    .X(net118));
 sg13g2_buf_2 fanout119 (.A(_2754_),
    .X(net119));
 sg13g2_buf_2 fanout120 (.A(_2415_),
    .X(net120));
 sg13g2_buf_2 fanout121 (.A(_2197_),
    .X(net121));
 sg13g2_buf_2 fanout122 (.A(_1713_),
    .X(net122));
 sg13g2_buf_2 fanout123 (.A(_1599_),
    .X(net123));
 sg13g2_buf_2 fanout124 (.A(_3895_),
    .X(net124));
 sg13g2_buf_2 fanout125 (.A(_3815_),
    .X(net125));
 sg13g2_buf_2 fanout126 (.A(_3760_),
    .X(net126));
 sg13g2_buf_2 fanout127 (.A(_3548_),
    .X(net127));
 sg13g2_buf_2 fanout128 (.A(_2766_),
    .X(net128));
 sg13g2_buf_2 fanout129 (.A(_2678_),
    .X(net129));
 sg13g2_buf_2 fanout130 (.A(_2334_),
    .X(net130));
 sg13g2_buf_2 fanout131 (.A(_2155_),
    .X(net131));
 sg13g2_buf_2 fanout132 (.A(_1604_),
    .X(net132));
 sg13g2_buf_2 fanout133 (.A(_3814_),
    .X(net133));
 sg13g2_buf_2 fanout134 (.A(_3690_),
    .X(net134));
 sg13g2_buf_2 fanout135 (.A(_2735_),
    .X(net135));
 sg13g2_buf_2 fanout136 (.A(_2560_),
    .X(net136));
 sg13g2_buf_2 fanout137 (.A(_2409_),
    .X(net137));
 sg13g2_buf_2 fanout138 (.A(_2336_),
    .X(net138));
 sg13g2_buf_2 fanout139 (.A(_2301_),
    .X(net139));
 sg13g2_buf_2 fanout140 (.A(_2265_),
    .X(net140));
 sg13g2_buf_2 fanout141 (.A(_2264_),
    .X(net141));
 sg13g2_buf_2 fanout142 (.A(_2154_),
    .X(net142));
 sg13g2_buf_2 fanout143 (.A(_2138_),
    .X(net143));
 sg13g2_buf_2 fanout144 (.A(_1998_),
    .X(net144));
 sg13g2_buf_2 fanout145 (.A(_1971_),
    .X(net145));
 sg13g2_buf_2 fanout146 (.A(_1945_),
    .X(net146));
 sg13g2_buf_2 fanout147 (.A(_0343_),
    .X(net147));
 sg13g2_buf_2 fanout148 (.A(_3697_),
    .X(net148));
 sg13g2_buf_2 fanout149 (.A(_3685_),
    .X(net149));
 sg13g2_buf_2 fanout150 (.A(_2952_),
    .X(net150));
 sg13g2_buf_2 fanout151 (.A(_2880_),
    .X(net151));
 sg13g2_buf_2 fanout152 (.A(_2791_),
    .X(net152));
 sg13g2_buf_2 fanout153 (.A(_2773_),
    .X(net153));
 sg13g2_buf_4 fanout154 (.X(net154),
    .A(_2332_));
 sg13g2_buf_2 fanout155 (.A(_2331_),
    .X(net155));
 sg13g2_buf_2 fanout156 (.A(_2295_),
    .X(net156));
 sg13g2_buf_2 fanout157 (.A(_2226_),
    .X(net157));
 sg13g2_buf_2 fanout158 (.A(_2164_),
    .X(net158));
 sg13g2_buf_2 fanout159 (.A(_2153_),
    .X(net159));
 sg13g2_buf_2 fanout160 (.A(_2097_),
    .X(net160));
 sg13g2_buf_2 fanout161 (.A(_2074_),
    .X(net161));
 sg13g2_buf_2 fanout162 (.A(_2028_),
    .X(net162));
 sg13g2_buf_2 fanout163 (.A(_1975_),
    .X(net163));
 sg13g2_buf_2 fanout164 (.A(_1970_),
    .X(net164));
 sg13g2_buf_2 fanout165 (.A(_1943_),
    .X(net165));
 sg13g2_buf_2 fanout166 (.A(_1942_),
    .X(net166));
 sg13g2_buf_2 fanout167 (.A(_1890_),
    .X(net167));
 sg13g2_buf_2 fanout168 (.A(_3493_),
    .X(net168));
 sg13g2_buf_2 fanout169 (.A(_3483_),
    .X(net169));
 sg13g2_buf_2 fanout170 (.A(_2749_),
    .X(net170));
 sg13g2_buf_2 fanout171 (.A(_2400_),
    .X(net171));
 sg13g2_buf_2 fanout172 (.A(_2398_),
    .X(net172));
 sg13g2_buf_2 fanout173 (.A(_2391_),
    .X(net173));
 sg13g2_buf_2 fanout174 (.A(_2315_),
    .X(net174));
 sg13g2_buf_2 fanout175 (.A(_2309_),
    .X(net175));
 sg13g2_buf_2 fanout176 (.A(_2032_),
    .X(net176));
 sg13g2_buf_2 fanout177 (.A(_1941_),
    .X(net177));
 sg13g2_buf_2 fanout178 (.A(_1920_),
    .X(net178));
 sg13g2_buf_2 fanout179 (.A(_1798_),
    .X(net179));
 sg13g2_buf_4 fanout180 (.X(net180),
    .A(_1768_));
 sg13g2_buf_4 fanout181 (.X(net181),
    .A(_3673_));
 sg13g2_buf_2 fanout182 (.A(_3514_),
    .X(net182));
 sg13g2_buf_2 fanout183 (.A(_3482_),
    .X(net183));
 sg13g2_tiehi \B_reg[0]$_SDFF_PP0__184  (.L_HI(net184));
 sg13g2_tiehi \B_reg[1]$_SDFF_PP0__185  (.L_HI(net185));
 sg13g2_tiehi \G_reg[0]$_SDFF_PP0__186  (.L_HI(net186));
 sg13g2_tiehi \G_reg[1]$_SDFF_PP0__187  (.L_HI(net187));
 sg13g2_tiehi \R_reg[0]$_SDFF_PP0__188  (.L_HI(net188));
 sg13g2_tiehi \R_reg[1]$_SDFF_PP0__189  (.L_HI(net189));
 sg13g2_tiehi _8024__190 (.L_HI(net190));
 sg13g2_tiehi _8026__191 (.L_HI(net191));
 sg13g2_tiehi _8027__192 (.L_HI(net192));
 sg13g2_tiehi _8028__193 (.L_HI(net193));
 sg13g2_tiehi _8029__194 (.L_HI(net194));
 sg13g2_tiehi _8030__195 (.L_HI(net195));
 sg13g2_tiehi _8031__196 (.L_HI(net196));
 sg13g2_tiehi _8032__197 (.L_HI(net197));
 sg13g2_tiehi _8033__198 (.L_HI(net198));
 sg13g2_tiehi \bitmap_pixel$_DFF_P__199  (.L_HI(net199));
 sg13g2_tiehi \i_collision.imp[0]$_SDFFE_PN0P__200  (.L_HI(net200));
 sg13g2_tiehi \i_collision.imp[1]$_SDFFE_PN0P__201  (.L_HI(net201));
 sg13g2_tiehi \i_collision.vx[0]$_SDFFE_PN0P__202  (.L_HI(net202));
 sg13g2_tiehi \i_collision.vx[1]$_SDFFE_PN1P__203  (.L_HI(net203));
 sg13g2_tiehi \i_collision.vx[2]$_SDFFE_PN0P__204  (.L_HI(net204));
 sg13g2_tiehi \i_collision.vy[0]$_SDFFE_PN1P__205  (.L_HI(net205));
 sg13g2_tiehi \i_collision.vy[1]$_SDFFE_PN0P__206  (.L_HI(net206));
 sg13g2_tiehi \i_collision.vy[2]$_SDFFE_PN0P__207  (.L_HI(net207));
 sg13g2_tiehi \i_collision.w[1]$_SDFFE_PN0P__208  (.L_HI(net208));
 sg13g2_tiehi \i_collision.w[2]$_SDFFE_PN0P__209  (.L_HI(net209));
 sg13g2_tiehi \i_colors.blue[0]$_SDFFE_PN1P__210  (.L_HI(net210));
 sg13g2_tiehi \i_colors.blue[1]$_SDFFE_PN0P__211  (.L_HI(net211));
 sg13g2_tiehi \i_colors.channel[0]$_DFF_P__212  (.L_HI(net212));
 sg13g2_tiehi \i_colors.channel[1]$_DFF_P__213  (.L_HI(net213));
 sg13g2_tiehi \i_colors.channel[2]$_DFF_P__214  (.L_HI(net214));
 sg13g2_tiehi \i_colors.green[0]$_SDFFE_PN1P__215  (.L_HI(net215));
 sg13g2_tiehi \i_colors.green[1]$_SDFFE_PN0P__216  (.L_HI(net216));
 sg13g2_tiehi \i_colors.red[0]$_SDFFE_PN1P__217  (.L_HI(net217));
 sg13g2_tiehi \i_colors.red[1]$_SDFFE_PN1P__218  (.L_HI(net218));
 sg13g2_tiehi \i_delta_sigma.acc[0]$_SDFF_PN0__219  (.L_HI(net219));
 sg13g2_tiehi \i_delta_sigma.acc[10]$_SDFF_PN0__220  (.L_HI(net220));
 sg13g2_tiehi \i_delta_sigma.acc[11]$_SDFF_PN0__221  (.L_HI(net221));
 sg13g2_tiehi \i_delta_sigma.acc[12]$_SDFF_PN0__222  (.L_HI(net222));
 sg13g2_tiehi \i_delta_sigma.acc[13]$_SDFF_PN0__223  (.L_HI(net223));
 sg13g2_tiehi \i_delta_sigma.acc[1]$_SDFF_PN0__224  (.L_HI(net224));
 sg13g2_tiehi \i_delta_sigma.acc[2]$_SDFF_PN0__225  (.L_HI(net225));
 sg13g2_tiehi \i_delta_sigma.acc[3]$_SDFF_PN0__226  (.L_HI(net226));
 sg13g2_tiehi \i_delta_sigma.acc[4]$_SDFF_PN0__227  (.L_HI(net227));
 sg13g2_tiehi \i_delta_sigma.acc[5]$_SDFF_PN0__228  (.L_HI(net228));
 sg13g2_tiehi \i_delta_sigma.acc[6]$_SDFF_PN0__229  (.L_HI(net229));
 sg13g2_tiehi \i_delta_sigma.acc[7]$_SDFF_PN0__230  (.L_HI(net230));
 sg13g2_tiehi \i_delta_sigma.acc[8]$_SDFF_PN0__231  (.L_HI(net231));
 sg13g2_tiehi \i_delta_sigma.acc[9]$_SDFF_PN0__232  (.L_HI(net232));
 sg13g2_tiehi \i_kinematics.center_x[0]$_SDFFE_PP0P__233  (.L_HI(net233));
 sg13g2_tiehi \i_kinematics.center_x[1]$_SDFFE_PP0P__234  (.L_HI(net234));
 sg13g2_tiehi \i_kinematics.center_x[2]$_SDFFE_PP0P__235  (.L_HI(net235));
 sg13g2_tiehi \i_kinematics.center_x[3]$_SDFFE_PP0P__236  (.L_HI(net236));
 sg13g2_tiehi \i_kinematics.center_x[4]$_SDFFE_PP0P__237  (.L_HI(net237));
 sg13g2_tiehi \i_kinematics.center_x[5]$_SDFFE_PP0P__238  (.L_HI(net238));
 sg13g2_tiehi \i_kinematics.center_x[6]$_SDFFE_PP1P__239  (.L_HI(net239));
 sg13g2_tiehi \i_kinematics.center_x[7]$_SDFFE_PP0P__240  (.L_HI(net240));
 sg13g2_tiehi \i_kinematics.center_x[8]$_SDFFE_PP1P__241  (.L_HI(net241));
 sg13g2_tiehi \i_kinematics.center_x[9]$_SDFFE_PP0P__242  (.L_HI(net242));
 sg13g2_tiehi \i_kinematics.center_x_lo[0]$_SDFFE_PP0P__243  (.L_HI(net243));
 sg13g2_tiehi \i_kinematics.center_x_lo[1]$_SDFFE_PP0P__244  (.L_HI(net244));
 sg13g2_tiehi \i_kinematics.center_y[0]$_SDFFE_PP0P__245  (.L_HI(net245));
 sg13g2_tiehi \i_kinematics.center_y[1]$_SDFFE_PP0P__246  (.L_HI(net246));
 sg13g2_tiehi \i_kinematics.center_y[2]$_SDFFE_PP0P__247  (.L_HI(net247));
 sg13g2_tiehi \i_kinematics.center_y[3]$_SDFFE_PP0P__248  (.L_HI(net248));
 sg13g2_tiehi \i_kinematics.center_y[4]$_SDFFE_PP1P__249  (.L_HI(net249));
 sg13g2_tiehi \i_kinematics.center_y[5]$_SDFFE_PP1P__250  (.L_HI(net250));
 sg13g2_tiehi \i_kinematics.center_y[6]$_SDFFE_PP1P__251  (.L_HI(net251));
 sg13g2_tiehi \i_kinematics.center_y[7]$_SDFFE_PP1P__252  (.L_HI(net252));
 sg13g2_tiehi \i_kinematics.center_y[8]$_SDFFE_PP0P__253  (.L_HI(net253));
 sg13g2_tiehi \i_kinematics.center_y[9]$_SDFFE_PP0P__254  (.L_HI(net254));
 sg13g2_tiehi \i_kinematics.center_y_lo[0]$_SDFFE_PP0P__255  (.L_HI(net255));
 sg13g2_tiehi \i_kinematics.center_y_lo[1]$_SDFFE_PP0P__256  (.L_HI(net256));
 sg13g2_tiehi \i_kinematics.phi[0]$_SDFFE_PP0P__257  (.L_HI(net257));
 sg13g2_tiehi \i_kinematics.phi[10]$_SDFFE_PP0P__258  (.L_HI(net258));
 sg13g2_tiehi \i_kinematics.phi[1]$_SDFFE_PP0P__259  (.L_HI(net259));
 sg13g2_tiehi \i_kinematics.phi[2]$_SDFFE_PP0P__260  (.L_HI(net260));
 sg13g2_tiehi \i_kinematics.phi[3]$_SDFFE_PP0P__261  (.L_HI(net261));
 sg13g2_tiehi \i_kinematics.phi[4]$_SDFFE_PP0P__262  (.L_HI(net262));
 sg13g2_tiehi \i_kinematics.phi[5]$_SDFFE_PP0P__263  (.L_HI(net263));
 sg13g2_tiehi \i_kinematics.phi[6]$_SDFFE_PP0P__264  (.L_HI(net264));
 sg13g2_tiehi \i_kinematics.phi[7]$_SDFFE_PP0P__265  (.L_HI(net265));
 sg13g2_tiehi \i_kinematics.phi[8]$_SDFFE_PP1P__266  (.L_HI(net266));
 sg13g2_tiehi \i_kinematics.phi[9]$_SDFFE_PP0P__267  (.L_HI(net267));
 sg13g2_tiehi \i_orchestrator.handle_impact$_SDFF_PP0__268  (.L_HI(net268));
 sg13g2_tiehi \i_orchestrator.hit_bottom$_SDFFE_PN0P__269  (.L_HI(net269));
 sg13g2_tiehi \i_orchestrator.hit_left$_SDFFE_PN0P__270  (.L_HI(net270));
 sg13g2_tiehi \i_orchestrator.hit_priority[0]$_SDFFE_PN0P__271  (.L_HI(net271));
 sg13g2_tiehi \i_orchestrator.hit_priority[1]$_SDFFE_PN0P__272  (.L_HI(net272));
 sg13g2_tiehi \i_orchestrator.hit_right$_SDFFE_PN0P__273  (.L_HI(net273));
 sg13g2_tiehi \i_orchestrator.hit_top$_SDFFE_PN0P__274  (.L_HI(net274));
 sg13g2_tiehi \i_orchestrator.lfsr[0]$_SDFFE_PN1P__275  (.L_HI(net275));
 sg13g2_tiehi \i_orchestrator.lfsr[1]$_SDFFE_PN1P__276  (.L_HI(net276));
 sg13g2_tiehi \i_orchestrator.lfsr[2]$_SDFFE_PN1P__277  (.L_HI(net277));
 sg13g2_tiehi \i_orchestrator.lfsr[3]$_SDFFE_PN1P__278  (.L_HI(net278));
 sg13g2_tiehi \i_orchestrator.lfsr[4]$_SDFFE_PN1P__279  (.L_HI(net279));
 sg13g2_tiehi \i_orchestrator.lfsr[5]$_SDFFE_PN1P__280  (.L_HI(net280));
 sg13g2_tiehi \i_orchestrator.lfsr[6]$_SDFFE_PN1P__281  (.L_HI(net281));
 sg13g2_tiehi \i_orchestrator.lfsr[7]$_SDFFE_PN1P__282  (.L_HI(net282));
 sg13g2_tiehi \i_orchestrator.lfsr[8]$_SDFFE_PN1P__283  (.L_HI(net283));
 sg13g2_tiehi \i_orchestrator.lfsr[9]$_SDFFE_PN1P__284  (.L_HI(net284));
 sg13g2_tiehi \i_orchestrator.mirror_collision$_SDFF_PN0__285  (.L_HI(net285));
 sg13g2_tiehi \i_orchestrator.rotate_collision$_SDFF_PN0__286  (.L_HI(net286));
 sg13g2_tiehi \i_orchestrator.sample_counter[0]$_SDFF_PN0__287  (.L_HI(net287));
 sg13g2_tiehi \i_orchestrator.sample_counter[1]$_SDFF_PN0__288  (.L_HI(net288));
 sg13g2_tiehi \i_orchestrator.sample_counter[2]$_SDFF_PN0__289  (.L_HI(net289));
 sg13g2_tiehi \i_orchestrator.sample_counter[3]$_SDFF_PN0__290  (.L_HI(net290));
 sg13g2_tiehi \i_orchestrator.sample_counter[4]$_SDFF_PN0__291  (.L_HI(net291));
 sg13g2_tiehi \i_orchestrator.sample_counter[5]$_SDFF_PN0__292  (.L_HI(net292));
 sg13g2_tiehi \i_orchestrator.sample_counter[6]$_SDFF_PN0__293  (.L_HI(net293));
 sg13g2_tiehi \i_orchestrator.sample_counter[7]$_SDFF_PN0__294  (.L_HI(net294));
 sg13g2_tiehi \i_orchestrator.sample_counter[8]$_SDFF_PN0__295  (.L_HI(net295));
 sg13g2_tiehi \i_orchestrator.sample_counter[9]$_SDFF_PN0__296  (.L_HI(net296));
 sg13g2_tiehi \i_orchestrator.tension[1]$_SDFFE_PN0P__297  (.L_HI(net297));
 sg13g2_tiehi \i_orchestrator.tension[2]$_SDFFE_PN0P__298  (.L_HI(net298));
 sg13g2_tiehi \i_orchestrator.tension[3]$_SDFFE_PN0P__299  (.L_HI(net299));
 sg13g2_tiehi \i_orchestrator.trigger_debounce$_SDFFE_PN0P__300  (.L_HI(net300));
 sg13g2_tiehi \i_orchestrator.trigger_resonator[0]$_SDFF_PP0__301  (.L_HI(net301));
 sg13g2_tiehi \i_orchestrator.trigger_resonator[1]$_SDFF_PP0__302  (.L_HI(net302));
 sg13g2_tiehi \i_orchestrator.update_collision$_SDFF_PN0__303  (.L_HI(net303));
 sg13g2_tiehi \i_orchestrator.update_kinematics$_SDFF_PP0__304  (.L_HI(net304));
 sg13g2_tiehi \i_orchestrator.update_resonator$_SDFF_PN0__305  (.L_HI(net305));
 sg13g2_tiehi \i_orchestrator.update_transform$_SDFF_PP0__306  (.L_HI(net306));
 sg13g2_tiehi \i_resonator.counter[0]$_SDFFE_PP0P__307  (.L_HI(net307));
 sg13g2_tiehi \i_resonator.counter[1]$_SDFFE_PP0P__308  (.L_HI(net308));
 sg13g2_tiehi \i_resonator.counter[2]$_SDFFE_PP0P__309  (.L_HI(net309));
 sg13g2_tiehi \i_resonator.counter[3]$_SDFFE_PP0P__310  (.L_HI(net310));
 sg13g2_tiehi \i_resonator.v[0]$_SDFFE_PP0P__311  (.L_HI(net311));
 sg13g2_tiehi \i_resonator.v[10]$_SDFFE_PP0P__312  (.L_HI(net312));
 sg13g2_tiehi \i_resonator.v[11]$_SDFFE_PP0P__313  (.L_HI(net313));
 sg13g2_tiehi \i_resonator.v[12]$_SDFFE_PP0P__314  (.L_HI(net314));
 sg13g2_tiehi \i_resonator.v[13]$_SDFFE_PP0P__315  (.L_HI(net315));
 sg13g2_tiehi \i_resonator.v[14]$_SDFFE_PP0P__316  (.L_HI(net316));
 sg13g2_tiehi \i_resonator.v[15]$_SDFFE_PP0P__317  (.L_HI(net317));
 sg13g2_tiehi \i_resonator.v[1]$_SDFFE_PP0P__318  (.L_HI(net318));
 sg13g2_tiehi \i_resonator.v[2]$_SDFFE_PP0P__319  (.L_HI(net319));
 sg13g2_tiehi \i_resonator.v[3]$_SDFFE_PP0P__320  (.L_HI(net320));
 sg13g2_tiehi \i_resonator.v[4]$_SDFFE_PP0P__321  (.L_HI(net321));
 sg13g2_tiehi \i_resonator.v[5]$_SDFFE_PP0P__322  (.L_HI(net322));
 sg13g2_tiehi \i_resonator.v[6]$_SDFFE_PP0P__323  (.L_HI(net323));
 sg13g2_tiehi \i_resonator.v[7]$_SDFFE_PP0P__324  (.L_HI(net324));
 sg13g2_tiehi \i_resonator.v[8]$_SDFFE_PP0P__325  (.L_HI(net325));
 sg13g2_tiehi \i_resonator.v[9]$_SDFFE_PP0P__326  (.L_HI(net326));
 sg13g2_tiehi \i_resonator.x[0]$_SDFFE_PP0P__327  (.L_HI(net327));
 sg13g2_tiehi \i_resonator.x[10]$_SDFFE_PP0P__328  (.L_HI(net328));
 sg13g2_tiehi \i_resonator.x[11]$_SDFFE_PP0P__329  (.L_HI(net329));
 sg13g2_tiehi \i_resonator.x[1]$_SDFFE_PP0P__330  (.L_HI(net330));
 sg13g2_tiehi \i_resonator.x[2]$_SDFFE_PP0P__331  (.L_HI(net331));
 sg13g2_tiehi \i_resonator.x[3]$_SDFFE_PP0P__332  (.L_HI(net332));
 sg13g2_tiehi \i_resonator.x[4]$_SDFFE_PP0P__333  (.L_HI(net333));
 sg13g2_tiehi \i_resonator.x[5]$_SDFFE_PP0P__334  (.L_HI(net334));
 sg13g2_tiehi \i_resonator.x[6]$_SDFFE_PP0P__335  (.L_HI(net335));
 sg13g2_tiehi \i_resonator.x[7]$_SDFFE_PP0P__336  (.L_HI(net336));
 sg13g2_tiehi \i_resonator.x[8]$_SDFFE_PP0P__337  (.L_HI(net337));
 sg13g2_tiehi \i_resonator.x[9]$_SDFFE_PP0P__338  (.L_HI(net338));
 sg13g2_tiehi \i_transform.image_x[0]$_SDFFE_PN0P__339  (.L_HI(net339));
 sg13g2_tiehi \i_transform.image_x[10]$_SDFFE_PN0N__340  (.L_HI(net340));
 sg13g2_tiehi \i_transform.image_x[11]$_SDFFE_PN0N__341  (.L_HI(net341));
 sg13g2_tiehi \i_transform.image_x[12]$_SDFFE_PN0N__342  (.L_HI(net342));
 sg13g2_tiehi \i_transform.image_x[13]$_SDFFE_PN0N__343  (.L_HI(net343));
 sg13g2_tiehi \i_transform.image_x[14]$_SDFFE_PN0N__344  (.L_HI(net344));
 sg13g2_tiehi \i_transform.image_x[15]$_SDFFE_PN0N__345  (.L_HI(net345));
 sg13g2_tiehi \i_transform.image_x[1]$_SDFFE_PN0P__346  (.L_HI(net346));
 sg13g2_tiehi \i_transform.image_x[2]$_SDFFE_PN0P__347  (.L_HI(net347));
 sg13g2_tiehi \i_transform.image_x[3]$_SDFFE_PN0P__348  (.L_HI(net348));
 sg13g2_tiehi \i_transform.image_x[4]$_SDFFE_PN0P__349  (.L_HI(net349));
 sg13g2_tiehi \i_transform.image_x[5]$_SDFFE_PN0N__350  (.L_HI(net350));
 sg13g2_tiehi \i_transform.image_x[6]$_SDFFE_PN0N__351  (.L_HI(net351));
 sg13g2_tiehi \i_transform.image_x[7]$_SDFFE_PN0N__352  (.L_HI(net352));
 sg13g2_tiehi \i_transform.image_x[8]$_SDFFE_PN0N__353  (.L_HI(net353));
 sg13g2_tiehi \i_transform.image_x[9]$_SDFFE_PN0N__354  (.L_HI(net354));
 sg13g2_tiehi \i_transform.image_y[0]$_SDFFE_PN0P__355  (.L_HI(net355));
 sg13g2_tiehi \i_transform.image_y[10]$_SDFFE_PN0N__356  (.L_HI(net356));
 sg13g2_tiehi \i_transform.image_y[11]$_SDFFE_PN0N__357  (.L_HI(net357));
 sg13g2_tiehi \i_transform.image_y[12]$_SDFFE_PN0N__358  (.L_HI(net358));
 sg13g2_tiehi \i_transform.image_y[13]$_SDFFE_PN0N__359  (.L_HI(net359));
 sg13g2_tiehi \i_transform.image_y[14]$_SDFFE_PN0N__360  (.L_HI(net360));
 sg13g2_tiehi \i_transform.image_y[15]$_SDFFE_PN0N__361  (.L_HI(net361));
 sg13g2_tiehi \i_transform.image_y[1]$_SDFFE_PN0P__362  (.L_HI(net362));
 sg13g2_tiehi \i_transform.image_y[2]$_SDFFE_PN0P__363  (.L_HI(net363));
 sg13g2_tiehi \i_transform.image_y[3]$_SDFFE_PN0P__364  (.L_HI(net364));
 sg13g2_tiehi \i_transform.image_y[4]$_SDFFE_PN0P__365  (.L_HI(net365));
 sg13g2_tiehi \i_transform.image_y[5]$_SDFFE_PN0N__366  (.L_HI(net366));
 sg13g2_tiehi \i_transform.image_y[6]$_SDFFE_PN0N__367  (.L_HI(net367));
 sg13g2_tiehi \i_transform.image_y[7]$_SDFFE_PN0N__368  (.L_HI(net368));
 sg13g2_tiehi \i_transform.image_y[8]$_SDFFE_PN0N__369  (.L_HI(net369));
 sg13g2_tiehi \i_transform.image_y[9]$_SDFFE_PN0N__370  (.L_HI(net370));
 sg13g2_tiehi \i_transform.track_x[0]$_DFFE_PP__371  (.L_HI(net371));
 sg13g2_tiehi \i_transform.track_x[1]$_DFFE_PP__372  (.L_HI(net372));
 sg13g2_tiehi \i_transform.track_x[2]$_DFFE_PP__373  (.L_HI(net373));
 sg13g2_tiehi \i_transform.track_x[3]$_DFFE_PP__374  (.L_HI(net374));
 sg13g2_tiehi \i_transform.track_x[4]$_DFFE_PP__375  (.L_HI(net375));
 sg13g2_tiehi \i_transform.track_x[5]$_DFFE_PP__376  (.L_HI(net376));
 sg13g2_tiehi \i_transform.track_x[6]$_DFFE_PP__377  (.L_HI(net377));
 sg13g2_tiehi \i_transform.track_x[7]$_DFFE_PP__378  (.L_HI(net378));
 sg13g2_tiehi \i_transform.track_x[8]$_DFFE_PP__379  (.L_HI(net379));
 sg13g2_tiehi \i_transform.track_x[9]$_DFFE_PP__380  (.L_HI(net380));
 sg13g2_tiehi \i_transform.track_y[0]$_DFFE_PP__381  (.L_HI(net381));
 sg13g2_tiehi \i_transform.track_y[1]$_DFFE_PP__382  (.L_HI(net382));
 sg13g2_tiehi \i_transform.track_y[2]$_DFFE_PP__383  (.L_HI(net383));
 sg13g2_tiehi \i_transform.track_y[3]$_DFFE_PP__384  (.L_HI(net384));
 sg13g2_tiehi \i_transform.track_y[4]$_DFFE_PP__385  (.L_HI(net385));
 sg13g2_tiehi \i_transform.track_y[5]$_DFFE_PP__386  (.L_HI(net386));
 sg13g2_tiehi \i_transform.track_y[6]$_DFFE_PP__387  (.L_HI(net387));
 sg13g2_tiehi \i_transform.track_y[7]$_DFFE_PP__388  (.L_HI(net388));
 sg13g2_tiehi \i_transform.track_y[8]$_DFFE_PP__389  (.L_HI(net389));
 sg13g2_tiehi \i_transform.track_y[9]$_DFFE_PP__390  (.L_HI(net390));
 sg13g2_tiehi \i_vga_beam.hsync$_DFF_P__391  (.L_HI(net391));
 sg13g2_tiehi \i_vga_beam.vsync$_DFF_P__392  (.L_HI(net392));
 sg13g2_tiehi \i_vga_beam.x[0]$_SDFF_PP0__393  (.L_HI(net393));
 sg13g2_tiehi \i_vga_beam.x[1]$_SDFF_PP0__394  (.L_HI(net394));
 sg13g2_tiehi \i_vga_beam.x[2]$_SDFF_PP0__395  (.L_HI(net395));
 sg13g2_tiehi \i_vga_beam.x[3]$_SDFF_PP0__396  (.L_HI(net396));
 sg13g2_tiehi \i_vga_beam.x[4]$_SDFF_PP0__397  (.L_HI(net397));
 sg13g2_tiehi \i_vga_beam.x[5]$_SDFF_PP0__398  (.L_HI(net398));
 sg13g2_tiehi \i_vga_beam.x[6]$_SDFF_PP0__399  (.L_HI(net399));
 sg13g2_tiehi \i_vga_beam.x[7]$_SDFF_PP0__400  (.L_HI(net400));
 sg13g2_tiehi \i_vga_beam.x[8]$_SDFF_PP0__401  (.L_HI(net401));
 sg13g2_tiehi \i_vga_beam.x[9]$_SDFF_PP0__402  (.L_HI(net402));
 sg13g2_tiehi \i_vga_beam.y[0]$_SDFFCE_PP0P__403  (.L_HI(net403));
 sg13g2_tiehi \i_vga_beam.y[1]$_SDFFCE_PP0P__404  (.L_HI(net404));
 sg13g2_tiehi \i_vga_beam.y[2]$_SDFFCE_PP0P__405  (.L_HI(net405));
 sg13g2_tiehi \i_vga_beam.y[3]$_SDFFCE_PP0P__406  (.L_HI(net406));
 sg13g2_tiehi \i_vga_beam.y[4]$_SDFFCE_PP0P__407  (.L_HI(net407));
 sg13g2_tiehi \i_vga_beam.y[5]$_SDFFCE_PP0P__408  (.L_HI(net408));
 sg13g2_tiehi \i_vga_beam.y[6]$_SDFFCE_PP0P__409  (.L_HI(net409));
 sg13g2_tiehi \i_vga_beam.y[7]$_SDFFCE_PP0P__410  (.L_HI(net410));
 sg13g2_tiehi \i_vga_beam.y[8]$_SDFFCE_PP0P__411  (.L_HI(net411));
 sg13g2_tiehi \i_vga_beam.y[9]$_SDFFCE_PP0P__412  (.L_HI(net412));
 sg13g2_tiehi \orient$_SDFFE_PN0P__413  (.L_HI(net413));
 sg13g2_buf_2 clkbuf_leaf_1_clk (.A(clknet_3_1__leaf_clk),
    .X(clknet_leaf_1_clk));
 sg13g2_buf_2 clkbuf_leaf_2_clk (.A(clknet_3_4__leaf_clk),
    .X(clknet_leaf_2_clk));
 sg13g2_buf_2 clkbuf_leaf_3_clk (.A(clknet_3_4__leaf_clk),
    .X(clknet_leaf_3_clk));
 sg13g2_buf_2 clkbuf_leaf_4_clk (.A(clknet_3_4__leaf_clk),
    .X(clknet_leaf_4_clk));
 sg13g2_buf_2 clkbuf_leaf_5_clk (.A(clknet_3_5__leaf_clk),
    .X(clknet_leaf_5_clk));
 sg13g2_buf_2 clkbuf_leaf_6_clk (.A(clknet_3_5__leaf_clk),
    .X(clknet_leaf_6_clk));
 sg13g2_buf_2 clkbuf_leaf_7_clk (.A(clknet_3_4__leaf_clk),
    .X(clknet_leaf_7_clk));
 sg13g2_buf_2 clkbuf_leaf_8_clk (.A(clknet_3_1__leaf_clk),
    .X(clknet_leaf_8_clk));
 sg13g2_buf_2 clkbuf_leaf_9_clk (.A(clknet_3_4__leaf_clk),
    .X(clknet_leaf_9_clk));
 sg13g2_buf_2 clkbuf_leaf_10_clk (.A(clknet_3_5__leaf_clk),
    .X(clknet_leaf_10_clk));
 sg13g2_buf_2 clkbuf_leaf_11_clk (.A(clknet_3_5__leaf_clk),
    .X(clknet_leaf_11_clk));
 sg13g2_buf_2 clkbuf_leaf_12_clk (.A(clknet_3_7__leaf_clk),
    .X(clknet_leaf_12_clk));
 sg13g2_buf_2 clkbuf_leaf_13_clk (.A(clknet_3_7__leaf_clk),
    .X(clknet_leaf_13_clk));
 sg13g2_buf_2 clkbuf_leaf_14_clk (.A(clknet_3_7__leaf_clk),
    .X(clknet_leaf_14_clk));
 sg13g2_buf_2 clkbuf_leaf_15_clk (.A(clknet_3_7__leaf_clk),
    .X(clknet_leaf_15_clk));
 sg13g2_buf_2 clkbuf_leaf_16_clk (.A(clknet_3_6__leaf_clk),
    .X(clknet_leaf_16_clk));
 sg13g2_buf_2 clkbuf_leaf_17_clk (.A(clknet_3_6__leaf_clk),
    .X(clknet_leaf_17_clk));
 sg13g2_buf_2 clkbuf_leaf_18_clk (.A(clknet_3_6__leaf_clk),
    .X(clknet_leaf_18_clk));
 sg13g2_buf_2 clkbuf_leaf_19_clk (.A(clknet_3_6__leaf_clk),
    .X(clknet_leaf_19_clk));
 sg13g2_buf_2 clkbuf_leaf_20_clk (.A(clknet_3_6__leaf_clk),
    .X(clknet_leaf_20_clk));
 sg13g2_buf_2 clkbuf_leaf_21_clk (.A(clknet_3_3__leaf_clk),
    .X(clknet_leaf_21_clk));
 sg13g2_buf_2 clkbuf_leaf_22_clk (.A(clknet_3_3__leaf_clk),
    .X(clknet_leaf_22_clk));
 sg13g2_buf_2 clkbuf_leaf_23_clk (.A(clknet_3_2__leaf_clk),
    .X(clknet_leaf_23_clk));
 sg13g2_buf_2 clkbuf_leaf_24_clk (.A(clknet_3_3__leaf_clk),
    .X(clknet_leaf_24_clk));
 sg13g2_buf_2 clkbuf_leaf_25_clk (.A(clknet_3_3__leaf_clk),
    .X(clknet_leaf_25_clk));
 sg13g2_buf_2 clkbuf_leaf_26_clk (.A(clknet_3_2__leaf_clk),
    .X(clknet_leaf_26_clk));
 sg13g2_buf_2 clkbuf_leaf_27_clk (.A(clknet_3_2__leaf_clk),
    .X(clknet_leaf_27_clk));
 sg13g2_buf_2 clkbuf_leaf_28_clk (.A(clknet_3_2__leaf_clk),
    .X(clknet_leaf_28_clk));
 sg13g2_buf_2 clkbuf_leaf_29_clk (.A(clknet_3_2__leaf_clk),
    .X(clknet_leaf_29_clk));
 sg13g2_buf_2 clkbuf_leaf_30_clk (.A(clknet_3_0__leaf_clk),
    .X(clknet_leaf_30_clk));
 sg13g2_buf_2 clkbuf_leaf_31_clk (.A(clknet_3_1__leaf_clk),
    .X(clknet_leaf_31_clk));
 sg13g2_buf_2 clkbuf_leaf_32_clk (.A(clknet_3_1__leaf_clk),
    .X(clknet_leaf_32_clk));
 sg13g2_buf_2 clkbuf_leaf_33_clk (.A(clknet_3_0__leaf_clk),
    .X(clknet_leaf_33_clk));
 sg13g2_buf_2 clkbuf_leaf_34_clk (.A(clknet_3_0__leaf_clk),
    .X(clknet_leaf_34_clk));
 sg13g2_buf_2 clkbuf_leaf_35_clk (.A(clknet_3_0__leaf_clk),
    .X(clknet_leaf_35_clk));
 sg13g2_buf_2 clkbuf_leaf_36_clk (.A(clknet_3_0__leaf_clk),
    .X(clknet_leaf_36_clk));
 sg13g2_buf_1 clkbuf_0_clk (.A(clk),
    .X(clknet_0_clk));
 sg13g2_buf_1 clkbuf_3_0__f_clk (.A(clknet_0_clk),
    .X(clknet_3_0__leaf_clk));
 sg13g2_buf_1 clkbuf_3_1__f_clk (.A(clknet_0_clk),
    .X(clknet_3_1__leaf_clk));
 sg13g2_buf_1 clkbuf_3_2__f_clk (.A(clknet_0_clk),
    .X(clknet_3_2__leaf_clk));
 sg13g2_buf_1 clkbuf_3_3__f_clk (.A(clknet_0_clk),
    .X(clknet_3_3__leaf_clk));
 sg13g2_buf_1 clkbuf_3_4__f_clk (.A(clknet_0_clk),
    .X(clknet_3_4__leaf_clk));
 sg13g2_buf_1 clkbuf_3_5__f_clk (.A(clknet_0_clk),
    .X(clknet_3_5__leaf_clk));
 sg13g2_buf_1 clkbuf_3_6__f_clk (.A(clknet_0_clk),
    .X(clknet_3_6__leaf_clk));
 sg13g2_buf_1 clkbuf_3_7__f_clk (.A(clknet_0_clk),
    .X(clknet_3_7__leaf_clk));
 sg13g2_buf_2 clkload0 (.A(clknet_3_3__leaf_clk));
 sg13g2_buf_2 clkload1 (.A(clknet_3_5__leaf_clk));
 sg13g2_buf_2 clkload2 (.A(clknet_3_7__leaf_clk));
 sg13g2_inv_4 clkload3 (.A(clknet_leaf_33_clk));
 sg13g2_inv_2 clkload4 (.A(clknet_leaf_34_clk));
 sg13g2_buf_16 clkload5 (.A(clknet_leaf_35_clk));
 sg13g2_inv_4 clkload6 (.A(clknet_leaf_36_clk));
 sg13g2_inv_4 clkload7 (.A(clknet_leaf_0_clk));
 sg13g2_buf_16 clkload8 (.A(clknet_leaf_1_clk));
 sg13g2_buf_16 clkload9 (.A(clknet_leaf_8_clk));
 sg13g2_inv_1 clkload10 (.A(clknet_leaf_31_clk));
 sg13g2_buf_16 clkload11 (.A(clknet_leaf_26_clk));
 sg13g2_buf_8 clkload12 (.A(clknet_leaf_27_clk));
 sg13g2_buf_8 clkload13 (.A(clknet_leaf_28_clk));
 sg13g2_inv_2 clkload14 (.A(clknet_leaf_29_clk));
 sg13g2_inv_1 clkload15 (.A(clknet_leaf_22_clk));
 sg13g2_buf_16 clkload16 (.A(clknet_leaf_24_clk));
 sg13g2_inv_2 clkload17 (.A(clknet_leaf_25_clk));
 sg13g2_buf_8 clkload18 (.A(clknet_leaf_2_clk));
 sg13g2_buf_16 clkload19 (.A(clknet_leaf_3_clk));
 sg13g2_buf_16 clkload20 (.A(clknet_leaf_4_clk));
 sg13g2_inv_2 clkload21 (.A(clknet_leaf_10_clk));
 sg13g2_inv_1 clkload22 (.A(clknet_leaf_13_clk));
 sg13g2_antennanp ANTENNA_1 (.A(_0148_));
 sg13g2_antennanp ANTENNA_2 (.A(clk));
 sg13g2_antennanp ANTENNA_3 (.A(clk));
 sg13g2_antennanp ANTENNA_4 (.A(clk));
 sg13g2_antennanp ANTENNA_5 (.A(_0148_));
 sg13g2_antennanp ANTENNA_6 (.A(_0148_));
 sg13g2_antennanp ANTENNA_7 (.A(_0148_));
 sg13g2_antennanp ANTENNA_8 (.A(_0148_));
 sg13g2_decap_8 FILLER_0_0 ();
 sg13g2_decap_8 FILLER_0_7 ();
 sg13g2_decap_8 FILLER_0_14 ();
 sg13g2_decap_8 FILLER_0_21 ();
 sg13g2_decap_8 FILLER_0_28 ();
 sg13g2_fill_2 FILLER_0_35 ();
 sg13g2_decap_8 FILLER_0_58 ();
 sg13g2_fill_1 FILLER_0_65 ();
 sg13g2_fill_1 FILLER_0_75 ();
 sg13g2_fill_2 FILLER_0_98 ();
 sg13g2_fill_2 FILLER_0_113 ();
 sg13g2_fill_2 FILLER_0_119 ();
 sg13g2_fill_1 FILLER_0_121 ();
 sg13g2_fill_2 FILLER_0_129 ();
 sg13g2_fill_1 FILLER_0_131 ();
 sg13g2_fill_1 FILLER_0_153 ();
 sg13g2_fill_2 FILLER_0_162 ();
 sg13g2_fill_1 FILLER_0_164 ();
 sg13g2_fill_1 FILLER_0_178 ();
 sg13g2_decap_4 FILLER_0_183 ();
 sg13g2_decap_8 FILLER_0_211 ();
 sg13g2_fill_2 FILLER_0_218 ();
 sg13g2_decap_8 FILLER_0_223 ();
 sg13g2_decap_4 FILLER_0_230 ();
 sg13g2_fill_1 FILLER_0_234 ();
 sg13g2_decap_8 FILLER_0_261 ();
 sg13g2_decap_4 FILLER_0_268 ();
 sg13g2_decap_8 FILLER_0_298 ();
 sg13g2_fill_2 FILLER_0_309 ();
 sg13g2_fill_1 FILLER_0_315 ();
 sg13g2_decap_4 FILLER_0_324 ();
 sg13g2_fill_1 FILLER_0_328 ();
 sg13g2_decap_8 FILLER_0_355 ();
 sg13g2_decap_8 FILLER_0_362 ();
 sg13g2_decap_8 FILLER_0_369 ();
 sg13g2_fill_1 FILLER_0_376 ();
 sg13g2_decap_8 FILLER_0_381 ();
 sg13g2_fill_1 FILLER_0_388 ();
 sg13g2_decap_8 FILLER_0_394 ();
 sg13g2_fill_2 FILLER_0_401 ();
 sg13g2_fill_1 FILLER_0_403 ();
 sg13g2_decap_8 FILLER_0_408 ();
 sg13g2_decap_8 FILLER_0_415 ();
 sg13g2_decap_8 FILLER_0_422 ();
 sg13g2_fill_1 FILLER_0_429 ();
 sg13g2_decap_8 FILLER_1_0 ();
 sg13g2_decap_8 FILLER_1_7 ();
 sg13g2_fill_2 FILLER_1_14 ();
 sg13g2_fill_2 FILLER_1_42 ();
 sg13g2_fill_1 FILLER_1_44 ();
 sg13g2_fill_1 FILLER_1_49 ();
 sg13g2_fill_1 FILLER_1_64 ();
 sg13g2_fill_1 FILLER_1_72 ();
 sg13g2_fill_1 FILLER_1_90 ();
 sg13g2_decap_4 FILLER_1_96 ();
 sg13g2_fill_2 FILLER_1_100 ();
 sg13g2_fill_1 FILLER_1_107 ();
 sg13g2_decap_8 FILLER_1_113 ();
 sg13g2_fill_2 FILLER_1_125 ();
 sg13g2_fill_2 FILLER_1_132 ();
 sg13g2_fill_1 FILLER_1_134 ();
 sg13g2_fill_2 FILLER_1_139 ();
 sg13g2_fill_2 FILLER_1_159 ();
 sg13g2_fill_1 FILLER_1_171 ();
 sg13g2_fill_2 FILLER_1_176 ();
 sg13g2_fill_1 FILLER_1_197 ();
 sg13g2_decap_4 FILLER_1_220 ();
 sg13g2_fill_1 FILLER_1_224 ();
 sg13g2_decap_8 FILLER_1_234 ();
 sg13g2_fill_2 FILLER_1_241 ();
 sg13g2_fill_1 FILLER_1_243 ();
 sg13g2_fill_2 FILLER_1_248 ();
 sg13g2_fill_2 FILLER_1_280 ();
 sg13g2_fill_2 FILLER_1_286 ();
 sg13g2_decap_4 FILLER_1_292 ();
 sg13g2_fill_2 FILLER_1_330 ();
 sg13g2_fill_1 FILLER_1_332 ();
 sg13g2_decap_8 FILLER_1_349 ();
 sg13g2_decap_8 FILLER_1_356 ();
 sg13g2_decap_8 FILLER_1_363 ();
 sg13g2_fill_2 FILLER_1_427 ();
 sg13g2_fill_1 FILLER_1_429 ();
 sg13g2_decap_8 FILLER_2_0 ();
 sg13g2_decap_8 FILLER_2_7 ();
 sg13g2_decap_8 FILLER_2_14 ();
 sg13g2_fill_2 FILLER_2_47 ();
 sg13g2_decap_4 FILLER_2_62 ();
 sg13g2_fill_2 FILLER_2_66 ();
 sg13g2_decap_8 FILLER_2_73 ();
 sg13g2_decap_8 FILLER_2_80 ();
 sg13g2_decap_4 FILLER_2_87 ();
 sg13g2_decap_8 FILLER_2_102 ();
 sg13g2_fill_2 FILLER_2_109 ();
 sg13g2_fill_1 FILLER_2_111 ();
 sg13g2_decap_4 FILLER_2_129 ();
 sg13g2_fill_1 FILLER_2_147 ();
 sg13g2_fill_2 FILLER_2_152 ();
 sg13g2_decap_8 FILLER_2_158 ();
 sg13g2_fill_2 FILLER_2_165 ();
 sg13g2_fill_1 FILLER_2_167 ();
 sg13g2_decap_8 FILLER_2_178 ();
 sg13g2_fill_1 FILLER_2_185 ();
 sg13g2_fill_1 FILLER_2_190 ();
 sg13g2_fill_2 FILLER_2_195 ();
 sg13g2_decap_8 FILLER_2_202 ();
 sg13g2_fill_1 FILLER_2_209 ();
 sg13g2_fill_2 FILLER_2_221 ();
 sg13g2_fill_2 FILLER_2_227 ();
 sg13g2_fill_1 FILLER_2_229 ();
 sg13g2_decap_8 FILLER_2_251 ();
 sg13g2_fill_1 FILLER_2_271 ();
 sg13g2_decap_4 FILLER_2_277 ();
 sg13g2_fill_1 FILLER_2_315 ();
 sg13g2_fill_1 FILLER_2_321 ();
 sg13g2_decap_4 FILLER_2_356 ();
 sg13g2_decap_8 FILLER_2_422 ();
 sg13g2_fill_1 FILLER_2_429 ();
 sg13g2_decap_4 FILLER_3_0 ();
 sg13g2_fill_2 FILLER_3_4 ();
 sg13g2_decap_4 FILLER_3_40 ();
 sg13g2_decap_4 FILLER_3_50 ();
 sg13g2_fill_2 FILLER_3_64 ();
 sg13g2_fill_1 FILLER_3_66 ();
 sg13g2_fill_2 FILLER_3_70 ();
 sg13g2_decap_8 FILLER_3_80 ();
 sg13g2_fill_1 FILLER_3_118 ();
 sg13g2_decap_8 FILLER_3_151 ();
 sg13g2_decap_4 FILLER_3_158 ();
 sg13g2_fill_2 FILLER_3_162 ();
 sg13g2_decap_4 FILLER_3_168 ();
 sg13g2_fill_1 FILLER_3_172 ();
 sg13g2_decap_4 FILLER_3_178 ();
 sg13g2_fill_2 FILLER_3_182 ();
 sg13g2_fill_2 FILLER_3_188 ();
 sg13g2_fill_1 FILLER_3_204 ();
 sg13g2_fill_2 FILLER_3_214 ();
 sg13g2_fill_1 FILLER_3_221 ();
 sg13g2_fill_1 FILLER_3_226 ();
 sg13g2_fill_2 FILLER_3_237 ();
 sg13g2_decap_8 FILLER_3_257 ();
 sg13g2_fill_1 FILLER_3_264 ();
 sg13g2_fill_2 FILLER_3_274 ();
 sg13g2_fill_1 FILLER_3_276 ();
 sg13g2_decap_4 FILLER_3_287 ();
 sg13g2_fill_1 FILLER_3_291 ();
 sg13g2_fill_1 FILLER_3_296 ();
 sg13g2_fill_2 FILLER_3_333 ();
 sg13g2_fill_1 FILLER_3_335 ();
 sg13g2_decap_8 FILLER_3_355 ();
 sg13g2_fill_2 FILLER_3_362 ();
 sg13g2_fill_2 FILLER_3_383 ();
 sg13g2_fill_1 FILLER_3_385 ();
 sg13g2_decap_4 FILLER_4_0 ();
 sg13g2_fill_1 FILLER_4_34 ();
 sg13g2_fill_2 FILLER_4_43 ();
 sg13g2_fill_2 FILLER_4_49 ();
 sg13g2_fill_2 FILLER_4_55 ();
 sg13g2_fill_1 FILLER_4_73 ();
 sg13g2_fill_1 FILLER_4_78 ();
 sg13g2_decap_8 FILLER_4_89 ();
 sg13g2_fill_1 FILLER_4_96 ();
 sg13g2_decap_8 FILLER_4_111 ();
 sg13g2_decap_4 FILLER_4_118 ();
 sg13g2_decap_8 FILLER_4_126 ();
 sg13g2_decap_8 FILLER_4_133 ();
 sg13g2_decap_8 FILLER_4_140 ();
 sg13g2_fill_2 FILLER_4_151 ();
 sg13g2_fill_1 FILLER_4_153 ();
 sg13g2_fill_1 FILLER_4_163 ();
 sg13g2_fill_1 FILLER_4_173 ();
 sg13g2_decap_8 FILLER_4_184 ();
 sg13g2_decap_8 FILLER_4_191 ();
 sg13g2_fill_2 FILLER_4_198 ();
 sg13g2_decap_4 FILLER_4_204 ();
 sg13g2_fill_2 FILLER_4_208 ();
 sg13g2_fill_1 FILLER_4_231 ();
 sg13g2_fill_1 FILLER_4_240 ();
 sg13g2_fill_1 FILLER_4_262 ();
 sg13g2_decap_4 FILLER_4_271 ();
 sg13g2_fill_1 FILLER_4_275 ();
 sg13g2_fill_2 FILLER_4_286 ();
 sg13g2_fill_1 FILLER_4_297 ();
 sg13g2_fill_2 FILLER_4_302 ();
 sg13g2_fill_1 FILLER_4_304 ();
 sg13g2_fill_2 FILLER_4_310 ();
 sg13g2_fill_1 FILLER_4_348 ();
 sg13g2_decap_8 FILLER_4_359 ();
 sg13g2_fill_2 FILLER_4_366 ();
 sg13g2_fill_1 FILLER_4_381 ();
 sg13g2_fill_1 FILLER_4_390 ();
 sg13g2_fill_1 FILLER_4_396 ();
 sg13g2_fill_2 FILLER_4_402 ();
 sg13g2_decap_8 FILLER_5_0 ();
 sg13g2_decap_8 FILLER_5_7 ();
 sg13g2_decap_8 FILLER_5_14 ();
 sg13g2_fill_1 FILLER_5_31 ();
 sg13g2_fill_1 FILLER_5_56 ();
 sg13g2_fill_1 FILLER_5_61 ();
 sg13g2_fill_1 FILLER_5_68 ();
 sg13g2_fill_1 FILLER_5_73 ();
 sg13g2_fill_1 FILLER_5_91 ();
 sg13g2_fill_1 FILLER_5_96 ();
 sg13g2_fill_1 FILLER_5_102 ();
 sg13g2_fill_1 FILLER_5_107 ();
 sg13g2_decap_8 FILLER_5_115 ();
 sg13g2_fill_1 FILLER_5_122 ();
 sg13g2_decap_4 FILLER_5_141 ();
 sg13g2_fill_2 FILLER_5_154 ();
 sg13g2_fill_2 FILLER_5_160 ();
 sg13g2_fill_1 FILLER_5_162 ();
 sg13g2_fill_2 FILLER_5_171 ();
 sg13g2_decap_4 FILLER_5_186 ();
 sg13g2_decap_4 FILLER_5_203 ();
 sg13g2_fill_1 FILLER_5_216 ();
 sg13g2_fill_2 FILLER_5_221 ();
 sg13g2_fill_1 FILLER_5_228 ();
 sg13g2_fill_2 FILLER_5_233 ();
 sg13g2_decap_4 FILLER_5_239 ();
 sg13g2_fill_2 FILLER_5_243 ();
 sg13g2_fill_1 FILLER_5_265 ();
 sg13g2_fill_2 FILLER_5_274 ();
 sg13g2_fill_1 FILLER_5_276 ();
 sg13g2_fill_2 FILLER_5_329 ();
 sg13g2_fill_2 FILLER_5_336 ();
 sg13g2_fill_1 FILLER_5_338 ();
 sg13g2_fill_1 FILLER_5_352 ();
 sg13g2_fill_2 FILLER_5_358 ();
 sg13g2_fill_1 FILLER_5_360 ();
 sg13g2_decap_4 FILLER_5_375 ();
 sg13g2_fill_2 FILLER_5_392 ();
 sg13g2_fill_2 FILLER_5_398 ();
 sg13g2_decap_4 FILLER_5_409 ();
 sg13g2_decap_4 FILLER_5_417 ();
 sg13g2_fill_2 FILLER_5_421 ();
 sg13g2_fill_2 FILLER_5_428 ();
 sg13g2_decap_8 FILLER_6_0 ();
 sg13g2_decap_8 FILLER_6_7 ();
 sg13g2_fill_2 FILLER_6_14 ();
 sg13g2_fill_2 FILLER_6_25 ();
 sg13g2_decap_4 FILLER_6_31 ();
 sg13g2_fill_1 FILLER_6_35 ();
 sg13g2_fill_2 FILLER_6_45 ();
 sg13g2_fill_1 FILLER_6_47 ();
 sg13g2_decap_8 FILLER_6_54 ();
 sg13g2_fill_1 FILLER_6_61 ();
 sg13g2_decap_8 FILLER_6_66 ();
 sg13g2_decap_8 FILLER_6_76 ();
 sg13g2_fill_2 FILLER_6_83 ();
 sg13g2_decap_4 FILLER_6_93 ();
 sg13g2_fill_1 FILLER_6_103 ();
 sg13g2_fill_1 FILLER_6_108 ();
 sg13g2_fill_1 FILLER_6_119 ();
 sg13g2_fill_1 FILLER_6_129 ();
 sg13g2_decap_4 FILLER_6_153 ();
 sg13g2_fill_1 FILLER_6_157 ();
 sg13g2_fill_1 FILLER_6_171 ();
 sg13g2_fill_1 FILLER_6_176 ();
 sg13g2_fill_2 FILLER_6_181 ();
 sg13g2_fill_1 FILLER_6_196 ();
 sg13g2_fill_1 FILLER_6_201 ();
 sg13g2_fill_1 FILLER_6_211 ();
 sg13g2_fill_2 FILLER_6_225 ();
 sg13g2_fill_1 FILLER_6_227 ();
 sg13g2_fill_2 FILLER_6_232 ();
 sg13g2_decap_8 FILLER_6_242 ();
 sg13g2_fill_2 FILLER_6_249 ();
 sg13g2_fill_2 FILLER_6_271 ();
 sg13g2_decap_8 FILLER_6_286 ();
 sg13g2_fill_2 FILLER_6_293 ();
 sg13g2_fill_2 FILLER_6_299 ();
 sg13g2_fill_2 FILLER_6_311 ();
 sg13g2_fill_1 FILLER_6_313 ();
 sg13g2_fill_1 FILLER_6_319 ();
 sg13g2_decap_8 FILLER_6_333 ();
 sg13g2_fill_2 FILLER_6_362 ();
 sg13g2_decap_8 FILLER_6_368 ();
 sg13g2_fill_1 FILLER_6_375 ();
 sg13g2_fill_1 FILLER_6_380 ();
 sg13g2_fill_1 FILLER_6_386 ();
 sg13g2_fill_2 FILLER_6_390 ();
 sg13g2_decap_8 FILLER_6_413 ();
 sg13g2_fill_1 FILLER_6_420 ();
 sg13g2_fill_1 FILLER_6_429 ();
 sg13g2_decap_8 FILLER_7_0 ();
 sg13g2_fill_2 FILLER_7_7 ();
 sg13g2_fill_1 FILLER_7_9 ();
 sg13g2_fill_1 FILLER_7_21 ();
 sg13g2_decap_4 FILLER_7_27 ();
 sg13g2_fill_2 FILLER_7_31 ();
 sg13g2_fill_2 FILLER_7_51 ();
 sg13g2_fill_1 FILLER_7_53 ();
 sg13g2_decap_4 FILLER_7_76 ();
 sg13g2_decap_8 FILLER_7_106 ();
 sg13g2_decap_8 FILLER_7_113 ();
 sg13g2_fill_2 FILLER_7_120 ();
 sg13g2_fill_1 FILLER_7_122 ();
 sg13g2_decap_4 FILLER_7_128 ();
 sg13g2_fill_1 FILLER_7_132 ();
 sg13g2_decap_8 FILLER_7_145 ();
 sg13g2_decap_8 FILLER_7_152 ();
 sg13g2_fill_2 FILLER_7_159 ();
 sg13g2_fill_1 FILLER_7_161 ();
 sg13g2_fill_2 FILLER_7_186 ();
 sg13g2_fill_2 FILLER_7_220 ();
 sg13g2_fill_1 FILLER_7_222 ();
 sg13g2_fill_2 FILLER_7_232 ();
 sg13g2_fill_1 FILLER_7_234 ();
 sg13g2_fill_2 FILLER_7_243 ();
 sg13g2_fill_1 FILLER_7_245 ();
 sg13g2_decap_4 FILLER_7_275 ();
 sg13g2_fill_1 FILLER_7_279 ();
 sg13g2_fill_1 FILLER_7_298 ();
 sg13g2_fill_1 FILLER_7_303 ();
 sg13g2_fill_1 FILLER_7_314 ();
 sg13g2_fill_2 FILLER_7_333 ();
 sg13g2_fill_2 FILLER_7_339 ();
 sg13g2_fill_2 FILLER_7_362 ();
 sg13g2_fill_1 FILLER_7_364 ();
 sg13g2_fill_1 FILLER_7_382 ();
 sg13g2_fill_1 FILLER_7_399 ();
 sg13g2_fill_2 FILLER_7_405 ();
 sg13g2_fill_2 FILLER_7_411 ();
 sg13g2_decap_8 FILLER_8_0 ();
 sg13g2_decap_4 FILLER_8_7 ();
 sg13g2_fill_1 FILLER_8_11 ();
 sg13g2_decap_8 FILLER_8_20 ();
 sg13g2_fill_2 FILLER_8_27 ();
 sg13g2_decap_4 FILLER_8_35 ();
 sg13g2_decap_8 FILLER_8_44 ();
 sg13g2_decap_8 FILLER_8_51 ();
 sg13g2_decap_4 FILLER_8_58 ();
 sg13g2_fill_2 FILLER_8_62 ();
 sg13g2_fill_1 FILLER_8_67 ();
 sg13g2_fill_1 FILLER_8_80 ();
 sg13g2_fill_2 FILLER_8_90 ();
 sg13g2_fill_2 FILLER_8_95 ();
 sg13g2_fill_1 FILLER_8_97 ();
 sg13g2_decap_8 FILLER_8_130 ();
 sg13g2_fill_2 FILLER_8_137 ();
 sg13g2_fill_1 FILLER_8_139 ();
 sg13g2_fill_1 FILLER_8_145 ();
 sg13g2_fill_2 FILLER_8_155 ();
 sg13g2_decap_4 FILLER_8_167 ();
 sg13g2_fill_1 FILLER_8_180 ();
 sg13g2_decap_4 FILLER_8_192 ();
 sg13g2_fill_2 FILLER_8_196 ();
 sg13g2_decap_4 FILLER_8_203 ();
 sg13g2_fill_1 FILLER_8_207 ();
 sg13g2_fill_1 FILLER_8_229 ();
 sg13g2_fill_1 FILLER_8_235 ();
 sg13g2_fill_2 FILLER_8_255 ();
 sg13g2_fill_2 FILLER_8_265 ();
 sg13g2_fill_1 FILLER_8_267 ();
 sg13g2_fill_1 FILLER_8_272 ();
 sg13g2_fill_2 FILLER_8_276 ();
 sg13g2_fill_1 FILLER_8_278 ();
 sg13g2_fill_2 FILLER_8_292 ();
 sg13g2_decap_4 FILLER_8_299 ();
 sg13g2_fill_2 FILLER_8_321 ();
 sg13g2_fill_1 FILLER_8_334 ();
 sg13g2_fill_1 FILLER_8_340 ();
 sg13g2_fill_1 FILLER_8_367 ();
 sg13g2_fill_1 FILLER_8_373 ();
 sg13g2_fill_1 FILLER_8_378 ();
 sg13g2_fill_2 FILLER_8_387 ();
 sg13g2_fill_1 FILLER_8_411 ();
 sg13g2_decap_4 FILLER_8_420 ();
 sg13g2_fill_2 FILLER_8_424 ();
 sg13g2_decap_8 FILLER_9_0 ();
 sg13g2_fill_2 FILLER_9_7 ();
 sg13g2_fill_1 FILLER_9_13 ();
 sg13g2_fill_2 FILLER_9_19 ();
 sg13g2_fill_1 FILLER_9_21 ();
 sg13g2_decap_4 FILLER_9_27 ();
 sg13g2_decap_8 FILLER_9_42 ();
 sg13g2_fill_1 FILLER_9_49 ();
 sg13g2_decap_8 FILLER_9_55 ();
 sg13g2_fill_2 FILLER_9_62 ();
 sg13g2_fill_1 FILLER_9_64 ();
 sg13g2_decap_4 FILLER_9_75 ();
 sg13g2_fill_2 FILLER_9_84 ();
 sg13g2_fill_1 FILLER_9_86 ();
 sg13g2_decap_8 FILLER_9_96 ();
 sg13g2_decap_8 FILLER_9_103 ();
 sg13g2_fill_2 FILLER_9_110 ();
 sg13g2_fill_2 FILLER_9_125 ();
 sg13g2_fill_1 FILLER_9_127 ();
 sg13g2_fill_1 FILLER_9_132 ();
 sg13g2_decap_8 FILLER_9_140 ();
 sg13g2_decap_8 FILLER_9_147 ();
 sg13g2_decap_4 FILLER_9_154 ();
 sg13g2_fill_1 FILLER_9_167 ();
 sg13g2_fill_1 FILLER_9_178 ();
 sg13g2_fill_2 FILLER_9_187 ();
 sg13g2_fill_2 FILLER_9_198 ();
 sg13g2_decap_8 FILLER_9_206 ();
 sg13g2_decap_4 FILLER_9_213 ();
 sg13g2_fill_1 FILLER_9_217 ();
 sg13g2_fill_1 FILLER_9_222 ();
 sg13g2_decap_8 FILLER_9_266 ();
 sg13g2_decap_4 FILLER_9_273 ();
 sg13g2_fill_2 FILLER_9_277 ();
 sg13g2_decap_4 FILLER_9_287 ();
 sg13g2_fill_1 FILLER_9_291 ();
 sg13g2_fill_1 FILLER_9_307 ();
 sg13g2_fill_1 FILLER_9_344 ();
 sg13g2_fill_2 FILLER_9_349 ();
 sg13g2_fill_2 FILLER_9_356 ();
 sg13g2_fill_2 FILLER_9_363 ();
 sg13g2_fill_1 FILLER_9_365 ();
 sg13g2_fill_1 FILLER_9_378 ();
 sg13g2_fill_2 FILLER_9_386 ();
 sg13g2_fill_1 FILLER_9_388 ();
 sg13g2_fill_1 FILLER_9_397 ();
 sg13g2_fill_1 FILLER_9_403 ();
 sg13g2_fill_1 FILLER_9_412 ();
 sg13g2_fill_1 FILLER_9_421 ();
 sg13g2_decap_8 FILLER_10_0 ();
 sg13g2_decap_4 FILLER_10_7 ();
 sg13g2_fill_2 FILLER_10_19 ();
 sg13g2_fill_1 FILLER_10_25 ();
 sg13g2_decap_4 FILLER_10_30 ();
 sg13g2_decap_4 FILLER_10_42 ();
 sg13g2_fill_2 FILLER_10_46 ();
 sg13g2_fill_2 FILLER_10_70 ();
 sg13g2_decap_4 FILLER_10_77 ();
 sg13g2_fill_2 FILLER_10_81 ();
 sg13g2_decap_4 FILLER_10_91 ();
 sg13g2_fill_1 FILLER_10_95 ();
 sg13g2_decap_8 FILLER_10_123 ();
 sg13g2_fill_2 FILLER_10_130 ();
 sg13g2_fill_2 FILLER_10_141 ();
 sg13g2_decap_8 FILLER_10_156 ();
 sg13g2_decap_8 FILLER_10_167 ();
 sg13g2_decap_8 FILLER_10_174 ();
 sg13g2_fill_2 FILLER_10_181 ();
 sg13g2_fill_2 FILLER_10_212 ();
 sg13g2_decap_8 FILLER_10_218 ();
 sg13g2_decap_4 FILLER_10_225 ();
 sg13g2_fill_1 FILLER_10_229 ();
 sg13g2_fill_2 FILLER_10_235 ();
 sg13g2_fill_2 FILLER_10_245 ();
 sg13g2_fill_1 FILLER_10_247 ();
 sg13g2_fill_2 FILLER_10_253 ();
 sg13g2_fill_1 FILLER_10_255 ();
 sg13g2_fill_2 FILLER_10_260 ();
 sg13g2_fill_1 FILLER_10_281 ();
 sg13g2_decap_4 FILLER_10_286 ();
 sg13g2_decap_8 FILLER_10_297 ();
 sg13g2_fill_2 FILLER_10_304 ();
 sg13g2_fill_2 FILLER_10_327 ();
 sg13g2_fill_1 FILLER_10_329 ();
 sg13g2_decap_4 FILLER_10_361 ();
 sg13g2_fill_2 FILLER_10_365 ();
 sg13g2_fill_2 FILLER_10_377 ();
 sg13g2_fill_1 FILLER_10_379 ();
 sg13g2_decap_4 FILLER_10_385 ();
 sg13g2_fill_1 FILLER_10_389 ();
 sg13g2_fill_2 FILLER_10_398 ();
 sg13g2_fill_1 FILLER_10_405 ();
 sg13g2_decap_4 FILLER_10_410 ();
 sg13g2_fill_1 FILLER_10_414 ();
 sg13g2_fill_2 FILLER_10_419 ();
 sg13g2_fill_1 FILLER_10_421 ();
 sg13g2_fill_2 FILLER_10_427 ();
 sg13g2_fill_1 FILLER_10_429 ();
 sg13g2_fill_2 FILLER_11_0 ();
 sg13g2_fill_1 FILLER_11_14 ();
 sg13g2_fill_1 FILLER_11_20 ();
 sg13g2_fill_2 FILLER_11_29 ();
 sg13g2_fill_1 FILLER_11_38 ();
 sg13g2_fill_1 FILLER_11_48 ();
 sg13g2_decap_4 FILLER_11_54 ();
 sg13g2_fill_2 FILLER_11_58 ();
 sg13g2_fill_2 FILLER_11_73 ();
 sg13g2_decap_8 FILLER_11_79 ();
 sg13g2_fill_2 FILLER_11_95 ();
 sg13g2_decap_8 FILLER_11_100 ();
 sg13g2_decap_4 FILLER_11_107 ();
 sg13g2_fill_2 FILLER_11_120 ();
 sg13g2_fill_1 FILLER_11_126 ();
 sg13g2_fill_1 FILLER_11_131 ();
 sg13g2_fill_1 FILLER_11_176 ();
 sg13g2_fill_2 FILLER_11_187 ();
 sg13g2_decap_4 FILLER_11_193 ();
 sg13g2_fill_2 FILLER_11_197 ();
 sg13g2_fill_2 FILLER_11_204 ();
 sg13g2_fill_1 FILLER_11_206 ();
 sg13g2_decap_4 FILLER_11_233 ();
 sg13g2_decap_8 FILLER_11_278 ();
 sg13g2_fill_2 FILLER_11_285 ();
 sg13g2_fill_1 FILLER_11_287 ();
 sg13g2_fill_2 FILLER_11_300 ();
 sg13g2_fill_2 FILLER_11_313 ();
 sg13g2_decap_4 FILLER_11_319 ();
 sg13g2_fill_2 FILLER_11_323 ();
 sg13g2_fill_2 FILLER_11_332 ();
 sg13g2_fill_2 FILLER_11_347 ();
 sg13g2_decap_8 FILLER_11_353 ();
 sg13g2_fill_2 FILLER_11_368 ();
 sg13g2_fill_1 FILLER_11_370 ();
 sg13g2_decap_8 FILLER_11_379 ();
 sg13g2_fill_2 FILLER_11_386 ();
 sg13g2_fill_1 FILLER_11_388 ();
 sg13g2_fill_1 FILLER_11_404 ();
 sg13g2_decap_4 FILLER_11_410 ();
 sg13g2_fill_2 FILLER_11_419 ();
 sg13g2_fill_2 FILLER_12_0 ();
 sg13g2_fill_1 FILLER_12_2 ();
 sg13g2_fill_1 FILLER_12_15 ();
 sg13g2_fill_2 FILLER_12_21 ();
 sg13g2_fill_1 FILLER_12_23 ();
 sg13g2_decap_8 FILLER_12_47 ();
 sg13g2_decap_4 FILLER_12_54 ();
 sg13g2_fill_2 FILLER_12_58 ();
 sg13g2_fill_2 FILLER_12_68 ();
 sg13g2_fill_1 FILLER_12_70 ();
 sg13g2_fill_1 FILLER_12_76 ();
 sg13g2_fill_2 FILLER_12_89 ();
 sg13g2_fill_1 FILLER_12_91 ();
 sg13g2_decap_4 FILLER_12_97 ();
 sg13g2_fill_2 FILLER_12_111 ();
 sg13g2_fill_1 FILLER_12_113 ();
 sg13g2_decap_8 FILLER_12_141 ();
 sg13g2_decap_4 FILLER_12_148 ();
 sg13g2_decap_4 FILLER_12_157 ();
 sg13g2_decap_8 FILLER_12_166 ();
 sg13g2_fill_1 FILLER_12_173 ();
 sg13g2_decap_4 FILLER_12_178 ();
 sg13g2_decap_4 FILLER_12_191 ();
 sg13g2_fill_1 FILLER_12_195 ();
 sg13g2_fill_2 FILLER_12_204 ();
 sg13g2_fill_1 FILLER_12_206 ();
 sg13g2_decap_8 FILLER_12_219 ();
 sg13g2_fill_1 FILLER_12_226 ();
 sg13g2_decap_8 FILLER_12_253 ();
 sg13g2_decap_8 FILLER_12_260 ();
 sg13g2_fill_1 FILLER_12_267 ();
 sg13g2_fill_2 FILLER_12_272 ();
 sg13g2_fill_2 FILLER_12_279 ();
 sg13g2_decap_4 FILLER_12_286 ();
 sg13g2_fill_2 FILLER_12_290 ();
 sg13g2_fill_1 FILLER_12_318 ();
 sg13g2_fill_1 FILLER_12_324 ();
 sg13g2_fill_2 FILLER_12_335 ();
 sg13g2_fill_1 FILLER_12_337 ();
 sg13g2_fill_1 FILLER_12_346 ();
 sg13g2_decap_8 FILLER_12_352 ();
 sg13g2_decap_4 FILLER_12_359 ();
 sg13g2_fill_1 FILLER_12_363 ();
 sg13g2_decap_4 FILLER_12_372 ();
 sg13g2_fill_2 FILLER_12_376 ();
 sg13g2_fill_2 FILLER_12_389 ();
 sg13g2_fill_1 FILLER_12_391 ();
 sg13g2_fill_1 FILLER_12_398 ();
 sg13g2_decap_4 FILLER_12_404 ();
 sg13g2_fill_1 FILLER_12_408 ();
 sg13g2_fill_1 FILLER_12_429 ();
 sg13g2_fill_1 FILLER_13_0 ();
 sg13g2_fill_1 FILLER_13_9 ();
 sg13g2_decap_4 FILLER_13_14 ();
 sg13g2_fill_2 FILLER_13_18 ();
 sg13g2_fill_2 FILLER_13_28 ();
 sg13g2_decap_8 FILLER_13_37 ();
 sg13g2_fill_2 FILLER_13_44 ();
 sg13g2_fill_1 FILLER_13_46 ();
 sg13g2_decap_4 FILLER_13_66 ();
 sg13g2_decap_8 FILLER_13_77 ();
 sg13g2_decap_4 FILLER_13_84 ();
 sg13g2_fill_1 FILLER_13_118 ();
 sg13g2_decap_4 FILLER_13_148 ();
 sg13g2_fill_1 FILLER_13_152 ();
 sg13g2_decap_4 FILLER_13_184 ();
 sg13g2_fill_1 FILLER_13_188 ();
 sg13g2_fill_2 FILLER_13_192 ();
 sg13g2_fill_1 FILLER_13_216 ();
 sg13g2_decap_8 FILLER_13_225 ();
 sg13g2_decap_4 FILLER_13_232 ();
 sg13g2_fill_2 FILLER_13_236 ();
 sg13g2_decap_4 FILLER_13_242 ();
 sg13g2_fill_1 FILLER_13_246 ();
 sg13g2_fill_1 FILLER_13_257 ();
 sg13g2_decap_8 FILLER_13_293 ();
 sg13g2_fill_1 FILLER_13_300 ();
 sg13g2_fill_1 FILLER_13_305 ();
 sg13g2_fill_1 FILLER_13_311 ();
 sg13g2_fill_1 FILLER_13_316 ();
 sg13g2_fill_1 FILLER_13_321 ();
 sg13g2_fill_1 FILLER_13_327 ();
 sg13g2_fill_1 FILLER_13_332 ();
 sg13g2_fill_1 FILLER_13_339 ();
 sg13g2_fill_1 FILLER_13_345 ();
 sg13g2_decap_4 FILLER_13_358 ();
 sg13g2_fill_2 FILLER_13_370 ();
 sg13g2_fill_1 FILLER_13_413 ();
 sg13g2_fill_1 FILLER_13_417 ();
 sg13g2_decap_8 FILLER_13_422 ();
 sg13g2_fill_1 FILLER_13_429 ();
 sg13g2_decap_4 FILLER_14_0 ();
 sg13g2_fill_1 FILLER_14_4 ();
 sg13g2_fill_2 FILLER_14_12 ();
 sg13g2_fill_1 FILLER_14_37 ();
 sg13g2_fill_1 FILLER_14_46 ();
 sg13g2_fill_2 FILLER_14_61 ();
 sg13g2_fill_1 FILLER_14_63 ();
 sg13g2_fill_1 FILLER_14_87 ();
 sg13g2_fill_2 FILLER_14_103 ();
 sg13g2_fill_1 FILLER_14_105 ();
 sg13g2_fill_1 FILLER_14_109 ();
 sg13g2_fill_2 FILLER_14_119 ();
 sg13g2_fill_1 FILLER_14_121 ();
 sg13g2_fill_1 FILLER_14_134 ();
 sg13g2_fill_2 FILLER_14_139 ();
 sg13g2_decap_8 FILLER_14_157 ();
 sg13g2_fill_1 FILLER_14_164 ();
 sg13g2_fill_2 FILLER_14_185 ();
 sg13g2_fill_1 FILLER_14_214 ();
 sg13g2_decap_8 FILLER_14_220 ();
 sg13g2_decap_4 FILLER_14_227 ();
 sg13g2_fill_1 FILLER_14_231 ();
 sg13g2_fill_2 FILLER_14_269 ();
 sg13g2_fill_1 FILLER_14_271 ();
 sg13g2_fill_2 FILLER_14_297 ();
 sg13g2_fill_1 FILLER_14_299 ();
 sg13g2_fill_2 FILLER_14_345 ();
 sg13g2_decap_8 FILLER_14_352 ();
 sg13g2_decap_4 FILLER_14_359 ();
 sg13g2_decap_8 FILLER_14_368 ();
 sg13g2_fill_1 FILLER_14_375 ();
 sg13g2_fill_2 FILLER_14_385 ();
 sg13g2_decap_4 FILLER_14_391 ();
 sg13g2_decap_4 FILLER_14_425 ();
 sg13g2_fill_1 FILLER_14_429 ();
 sg13g2_fill_2 FILLER_15_0 ();
 sg13g2_decap_4 FILLER_15_15 ();
 sg13g2_fill_1 FILLER_15_26 ();
 sg13g2_fill_1 FILLER_15_32 ();
 sg13g2_fill_1 FILLER_15_37 ();
 sg13g2_fill_2 FILLER_15_43 ();
 sg13g2_fill_2 FILLER_15_55 ();
 sg13g2_fill_2 FILLER_15_75 ();
 sg13g2_fill_1 FILLER_15_77 ();
 sg13g2_fill_1 FILLER_15_88 ();
 sg13g2_fill_1 FILLER_15_93 ();
 sg13g2_decap_8 FILLER_15_100 ();
 sg13g2_fill_2 FILLER_15_107 ();
 sg13g2_decap_8 FILLER_15_113 ();
 sg13g2_fill_1 FILLER_15_120 ();
 sg13g2_decap_4 FILLER_15_126 ();
 sg13g2_fill_1 FILLER_15_130 ();
 sg13g2_fill_2 FILLER_15_162 ();
 sg13g2_fill_2 FILLER_15_170 ();
 sg13g2_fill_1 FILLER_15_172 ();
 sg13g2_decap_4 FILLER_15_181 ();
 sg13g2_fill_2 FILLER_15_185 ();
 sg13g2_decap_4 FILLER_15_230 ();
 sg13g2_fill_2 FILLER_15_234 ();
 sg13g2_fill_1 FILLER_15_246 ();
 sg13g2_fill_1 FILLER_15_255 ();
 sg13g2_fill_1 FILLER_15_264 ();
 sg13g2_fill_2 FILLER_15_270 ();
 sg13g2_fill_1 FILLER_15_272 ();
 sg13g2_fill_2 FILLER_15_290 ();
 sg13g2_fill_2 FILLER_15_338 ();
 sg13g2_decap_8 FILLER_15_350 ();
 sg13g2_fill_1 FILLER_15_357 ();
 sg13g2_fill_1 FILLER_15_366 ();
 sg13g2_fill_1 FILLER_15_372 ();
 sg13g2_fill_1 FILLER_15_385 ();
 sg13g2_fill_1 FILLER_15_402 ();
 sg13g2_decap_4 FILLER_15_411 ();
 sg13g2_fill_1 FILLER_15_420 ();
 sg13g2_fill_1 FILLER_15_429 ();
 sg13g2_decap_8 FILLER_16_0 ();
 sg13g2_fill_2 FILLER_16_7 ();
 sg13g2_fill_1 FILLER_16_9 ();
 sg13g2_fill_1 FILLER_16_15 ();
 sg13g2_fill_1 FILLER_16_26 ();
 sg13g2_fill_1 FILLER_16_36 ();
 sg13g2_fill_1 FILLER_16_40 ();
 sg13g2_fill_1 FILLER_16_52 ();
 sg13g2_fill_2 FILLER_16_57 ();
 sg13g2_fill_1 FILLER_16_59 ();
 sg13g2_fill_1 FILLER_16_67 ();
 sg13g2_decap_4 FILLER_16_72 ();
 sg13g2_fill_2 FILLER_16_102 ();
 sg13g2_fill_1 FILLER_16_104 ();
 sg13g2_decap_8 FILLER_16_122 ();
 sg13g2_decap_8 FILLER_16_129 ();
 sg13g2_decap_8 FILLER_16_136 ();
 sg13g2_fill_1 FILLER_16_143 ();
 sg13g2_fill_1 FILLER_16_165 ();
 sg13g2_decap_4 FILLER_16_173 ();
 sg13g2_fill_2 FILLER_16_201 ();
 sg13g2_fill_2 FILLER_16_211 ();
 sg13g2_fill_1 FILLER_16_213 ();
 sg13g2_decap_8 FILLER_16_217 ();
 sg13g2_fill_1 FILLER_16_224 ();
 sg13g2_fill_2 FILLER_16_229 ();
 sg13g2_decap_4 FILLER_16_236 ();
 sg13g2_fill_2 FILLER_16_254 ();
 sg13g2_fill_2 FILLER_16_266 ();
 sg13g2_fill_1 FILLER_16_268 ();
 sg13g2_fill_1 FILLER_16_302 ();
 sg13g2_fill_1 FILLER_16_313 ();
 sg13g2_decap_4 FILLER_16_354 ();
 sg13g2_fill_1 FILLER_16_358 ();
 sg13g2_fill_2 FILLER_16_383 ();
 sg13g2_fill_2 FILLER_16_388 ();
 sg13g2_fill_1 FILLER_16_390 ();
 sg13g2_fill_1 FILLER_16_394 ();
 sg13g2_fill_2 FILLER_16_410 ();
 sg13g2_fill_1 FILLER_16_412 ();
 sg13g2_fill_1 FILLER_16_420 ();
 sg13g2_fill_1 FILLER_16_429 ();
 sg13g2_decap_4 FILLER_17_4 ();
 sg13g2_fill_1 FILLER_17_8 ();
 sg13g2_fill_2 FILLER_17_17 ();
 sg13g2_fill_1 FILLER_17_23 ();
 sg13g2_fill_2 FILLER_17_27 ();
 sg13g2_fill_1 FILLER_17_29 ();
 sg13g2_fill_1 FILLER_17_35 ();
 sg13g2_fill_2 FILLER_17_41 ();
 sg13g2_fill_1 FILLER_17_59 ();
 sg13g2_fill_1 FILLER_17_69 ();
 sg13g2_fill_1 FILLER_17_75 ();
 sg13g2_decap_4 FILLER_17_81 ();
 sg13g2_fill_1 FILLER_17_91 ();
 sg13g2_decap_8 FILLER_17_96 ();
 sg13g2_fill_1 FILLER_17_103 ();
 sg13g2_decap_8 FILLER_17_122 ();
 sg13g2_fill_1 FILLER_17_129 ();
 sg13g2_fill_1 FILLER_17_144 ();
 sg13g2_fill_1 FILLER_17_150 ();
 sg13g2_fill_1 FILLER_17_161 ();
 sg13g2_fill_1 FILLER_17_167 ();
 sg13g2_fill_1 FILLER_17_175 ();
 sg13g2_fill_2 FILLER_17_193 ();
 sg13g2_fill_2 FILLER_17_201 ();
 sg13g2_fill_2 FILLER_17_207 ();
 sg13g2_fill_2 FILLER_17_217 ();
 sg13g2_fill_1 FILLER_17_219 ();
 sg13g2_decap_8 FILLER_17_274 ();
 sg13g2_decap_8 FILLER_17_281 ();
 sg13g2_fill_2 FILLER_17_288 ();
 sg13g2_fill_1 FILLER_17_290 ();
 sg13g2_decap_4 FILLER_17_296 ();
 sg13g2_fill_1 FILLER_17_300 ();
 sg13g2_fill_1 FILLER_17_307 ();
 sg13g2_fill_1 FILLER_17_324 ();
 sg13g2_decap_8 FILLER_17_348 ();
 sg13g2_fill_2 FILLER_17_355 ();
 sg13g2_decap_4 FILLER_17_373 ();
 sg13g2_fill_1 FILLER_17_395 ();
 sg13g2_decap_8 FILLER_17_407 ();
 sg13g2_fill_1 FILLER_17_414 ();
 sg13g2_decap_4 FILLER_17_420 ();
 sg13g2_fill_1 FILLER_17_429 ();
 sg13g2_decap_8 FILLER_18_0 ();
 sg13g2_decap_8 FILLER_18_7 ();
 sg13g2_fill_2 FILLER_18_14 ();
 sg13g2_fill_1 FILLER_18_16 ();
 sg13g2_fill_1 FILLER_18_33 ();
 sg13g2_fill_2 FILLER_18_42 ();
 sg13g2_decap_4 FILLER_18_52 ();
 sg13g2_fill_1 FILLER_18_60 ();
 sg13g2_fill_2 FILLER_18_73 ();
 sg13g2_fill_1 FILLER_18_75 ();
 sg13g2_fill_2 FILLER_18_85 ();
 sg13g2_fill_1 FILLER_18_87 ();
 sg13g2_decap_8 FILLER_18_101 ();
 sg13g2_fill_2 FILLER_18_141 ();
 sg13g2_fill_1 FILLER_18_152 ();
 sg13g2_decap_8 FILLER_18_161 ();
 sg13g2_fill_2 FILLER_18_173 ();
 sg13g2_fill_1 FILLER_18_180 ();
 sg13g2_fill_2 FILLER_18_188 ();
 sg13g2_decap_4 FILLER_18_226 ();
 sg13g2_fill_1 FILLER_18_230 ();
 sg13g2_decap_4 FILLER_18_236 ();
 sg13g2_fill_2 FILLER_18_240 ();
 sg13g2_fill_1 FILLER_18_250 ();
 sg13g2_fill_2 FILLER_18_273 ();
 sg13g2_decap_4 FILLER_18_288 ();
 sg13g2_fill_2 FILLER_18_292 ();
 sg13g2_fill_1 FILLER_18_311 ();
 sg13g2_decap_4 FILLER_18_317 ();
 sg13g2_fill_2 FILLER_18_321 ();
 sg13g2_fill_1 FILLER_18_328 ();
 sg13g2_fill_1 FILLER_18_334 ();
 sg13g2_fill_1 FILLER_18_339 ();
 sg13g2_decap_4 FILLER_18_387 ();
 sg13g2_fill_1 FILLER_18_391 ();
 sg13g2_fill_1 FILLER_18_401 ();
 sg13g2_fill_2 FILLER_18_427 ();
 sg13g2_fill_1 FILLER_18_429 ();
 sg13g2_fill_2 FILLER_19_0 ();
 sg13g2_fill_1 FILLER_19_5 ();
 sg13g2_fill_2 FILLER_19_10 ();
 sg13g2_fill_2 FILLER_19_17 ();
 sg13g2_fill_1 FILLER_19_19 ();
 sg13g2_fill_1 FILLER_19_37 ();
 sg13g2_fill_2 FILLER_19_42 ();
 sg13g2_decap_8 FILLER_19_52 ();
 sg13g2_fill_2 FILLER_19_59 ();
 sg13g2_fill_1 FILLER_19_72 ();
 sg13g2_decap_8 FILLER_19_87 ();
 sg13g2_fill_1 FILLER_19_94 ();
 sg13g2_fill_1 FILLER_19_101 ();
 sg13g2_decap_4 FILLER_19_126 ();
 sg13g2_fill_2 FILLER_19_130 ();
 sg13g2_fill_2 FILLER_19_136 ();
 sg13g2_fill_1 FILLER_19_138 ();
 sg13g2_fill_2 FILLER_19_154 ();
 sg13g2_fill_2 FILLER_19_173 ();
 sg13g2_fill_2 FILLER_19_179 ();
 sg13g2_fill_1 FILLER_19_181 ();
 sg13g2_decap_4 FILLER_19_188 ();
 sg13g2_decap_8 FILLER_19_197 ();
 sg13g2_fill_2 FILLER_19_204 ();
 sg13g2_fill_1 FILLER_19_206 ();
 sg13g2_decap_8 FILLER_19_211 ();
 sg13g2_decap_4 FILLER_19_218 ();
 sg13g2_fill_1 FILLER_19_222 ();
 sg13g2_decap_8 FILLER_19_240 ();
 sg13g2_decap_4 FILLER_19_255 ();
 sg13g2_fill_2 FILLER_19_293 ();
 sg13g2_fill_2 FILLER_19_302 ();
 sg13g2_decap_4 FILLER_19_309 ();
 sg13g2_fill_1 FILLER_19_323 ();
 sg13g2_fill_2 FILLER_19_335 ();
 sg13g2_fill_1 FILLER_19_346 ();
 sg13g2_fill_1 FILLER_19_356 ();
 sg13g2_fill_1 FILLER_19_365 ();
 sg13g2_fill_2 FILLER_19_370 ();
 sg13g2_fill_1 FILLER_19_379 ();
 sg13g2_decap_4 FILLER_19_384 ();
 sg13g2_fill_1 FILLER_19_388 ();
 sg13g2_decap_4 FILLER_19_394 ();
 sg13g2_fill_2 FILLER_19_402 ();
 sg13g2_fill_1 FILLER_19_404 ();
 sg13g2_fill_1 FILLER_19_429 ();
 sg13g2_fill_1 FILLER_20_30 ();
 sg13g2_decap_8 FILLER_20_39 ();
 sg13g2_decap_8 FILLER_20_46 ();
 sg13g2_fill_2 FILLER_20_53 ();
 sg13g2_fill_2 FILLER_20_60 ();
 sg13g2_fill_1 FILLER_20_62 ();
 sg13g2_fill_2 FILLER_20_68 ();
 sg13g2_fill_1 FILLER_20_70 ();
 sg13g2_fill_2 FILLER_20_76 ();
 sg13g2_fill_1 FILLER_20_78 ();
 sg13g2_decap_4 FILLER_20_89 ();
 sg13g2_decap_4 FILLER_20_98 ();
 sg13g2_fill_1 FILLER_20_102 ();
 sg13g2_fill_2 FILLER_20_107 ();
 sg13g2_fill_1 FILLER_20_109 ();
 sg13g2_fill_2 FILLER_20_113 ();
 sg13g2_fill_2 FILLER_20_119 ();
 sg13g2_fill_1 FILLER_20_121 ();
 sg13g2_fill_2 FILLER_20_130 ();
 sg13g2_fill_1 FILLER_20_132 ();
 sg13g2_fill_1 FILLER_20_152 ();
 sg13g2_fill_1 FILLER_20_200 ();
 sg13g2_decap_8 FILLER_20_218 ();
 sg13g2_fill_2 FILLER_20_225 ();
 sg13g2_fill_1 FILLER_20_227 ();
 sg13g2_fill_2 FILLER_20_232 ();
 sg13g2_fill_1 FILLER_20_234 ();
 sg13g2_fill_1 FILLER_20_247 ();
 sg13g2_decap_8 FILLER_20_257 ();
 sg13g2_decap_4 FILLER_20_264 ();
 sg13g2_fill_2 FILLER_20_268 ();
 sg13g2_decap_4 FILLER_20_282 ();
 sg13g2_decap_8 FILLER_20_290 ();
 sg13g2_decap_4 FILLER_20_297 ();
 sg13g2_fill_1 FILLER_20_301 ();
 sg13g2_decap_8 FILLER_20_306 ();
 sg13g2_decap_4 FILLER_20_313 ();
 sg13g2_fill_1 FILLER_20_317 ();
 sg13g2_fill_2 FILLER_20_332 ();
 sg13g2_fill_2 FILLER_20_341 ();
 sg13g2_fill_2 FILLER_20_378 ();
 sg13g2_fill_2 FILLER_20_384 ();
 sg13g2_fill_2 FILLER_20_391 ();
 sg13g2_decap_8 FILLER_20_408 ();
 sg13g2_decap_4 FILLER_20_415 ();
 sg13g2_fill_2 FILLER_20_419 ();
 sg13g2_fill_2 FILLER_21_0 ();
 sg13g2_fill_1 FILLER_21_10 ();
 sg13g2_fill_2 FILLER_21_18 ();
 sg13g2_decap_4 FILLER_21_25 ();
 sg13g2_fill_1 FILLER_21_29 ();
 sg13g2_fill_2 FILLER_21_43 ();
 sg13g2_fill_1 FILLER_21_45 ();
 sg13g2_fill_1 FILLER_21_54 ();
 sg13g2_fill_2 FILLER_21_86 ();
 sg13g2_fill_1 FILLER_21_119 ();
 sg13g2_fill_1 FILLER_21_124 ();
 sg13g2_fill_1 FILLER_21_129 ();
 sg13g2_fill_1 FILLER_21_139 ();
 sg13g2_decap_4 FILLER_21_152 ();
 sg13g2_fill_1 FILLER_21_156 ();
 sg13g2_decap_8 FILLER_21_162 ();
 sg13g2_fill_1 FILLER_21_169 ();
 sg13g2_decap_4 FILLER_21_174 ();
 sg13g2_fill_2 FILLER_21_178 ();
 sg13g2_decap_8 FILLER_21_188 ();
 sg13g2_fill_1 FILLER_21_245 ();
 sg13g2_fill_2 FILLER_21_276 ();
 sg13g2_fill_1 FILLER_21_311 ();
 sg13g2_fill_1 FILLER_21_340 ();
 sg13g2_fill_2 FILLER_21_382 ();
 sg13g2_fill_1 FILLER_21_408 ();
 sg13g2_decap_4 FILLER_21_413 ();
 sg13g2_fill_1 FILLER_21_417 ();
 sg13g2_decap_4 FILLER_21_426 ();
 sg13g2_fill_2 FILLER_22_0 ();
 sg13g2_fill_1 FILLER_22_2 ();
 sg13g2_fill_1 FILLER_22_14 ();
 sg13g2_fill_1 FILLER_22_18 ();
 sg13g2_decap_8 FILLER_22_27 ();
 sg13g2_fill_1 FILLER_22_38 ();
 sg13g2_fill_1 FILLER_22_47 ();
 sg13g2_decap_8 FILLER_22_51 ();
 sg13g2_fill_1 FILLER_22_71 ();
 sg13g2_fill_1 FILLER_22_75 ();
 sg13g2_fill_1 FILLER_22_80 ();
 sg13g2_decap_4 FILLER_22_90 ();
 sg13g2_fill_1 FILLER_22_108 ();
 sg13g2_fill_1 FILLER_22_112 ();
 sg13g2_fill_1 FILLER_22_117 ();
 sg13g2_decap_8 FILLER_22_127 ();
 sg13g2_fill_2 FILLER_22_134 ();
 sg13g2_fill_1 FILLER_22_141 ();
 sg13g2_fill_1 FILLER_22_157 ();
 sg13g2_fill_1 FILLER_22_162 ();
 sg13g2_fill_2 FILLER_22_167 ();
 sg13g2_fill_2 FILLER_22_177 ();
 sg13g2_fill_1 FILLER_22_179 ();
 sg13g2_fill_1 FILLER_22_187 ();
 sg13g2_fill_2 FILLER_22_223 ();
 sg13g2_decap_8 FILLER_22_230 ();
 sg13g2_fill_2 FILLER_22_237 ();
 sg13g2_fill_2 FILLER_22_251 ();
 sg13g2_fill_1 FILLER_22_262 ();
 sg13g2_fill_2 FILLER_22_267 ();
 sg13g2_fill_1 FILLER_22_269 ();
 sg13g2_decap_4 FILLER_22_278 ();
 sg13g2_fill_1 FILLER_22_282 ();
 sg13g2_decap_8 FILLER_22_288 ();
 sg13g2_fill_1 FILLER_22_295 ();
 sg13g2_fill_2 FILLER_22_301 ();
 sg13g2_fill_2 FILLER_22_341 ();
 sg13g2_decap_8 FILLER_22_346 ();
 sg13g2_fill_1 FILLER_22_353 ();
 sg13g2_decap_8 FILLER_22_365 ();
 sg13g2_decap_4 FILLER_22_380 ();
 sg13g2_fill_1 FILLER_22_392 ();
 sg13g2_fill_1 FILLER_22_405 ();
 sg13g2_fill_2 FILLER_22_413 ();
 sg13g2_decap_4 FILLER_22_425 ();
 sg13g2_fill_1 FILLER_22_429 ();
 sg13g2_decap_8 FILLER_23_0 ();
 sg13g2_fill_1 FILLER_23_7 ();
 sg13g2_fill_1 FILLER_23_13 ();
 sg13g2_fill_2 FILLER_23_19 ();
 sg13g2_fill_1 FILLER_23_50 ();
 sg13g2_fill_1 FILLER_23_62 ();
 sg13g2_fill_2 FILLER_23_68 ();
 sg13g2_fill_1 FILLER_23_70 ();
 sg13g2_fill_2 FILLER_23_76 ();
 sg13g2_fill_1 FILLER_23_78 ();
 sg13g2_fill_1 FILLER_23_82 ();
 sg13g2_decap_4 FILLER_23_91 ();
 sg13g2_fill_2 FILLER_23_99 ();
 sg13g2_fill_1 FILLER_23_105 ();
 sg13g2_decap_8 FILLER_23_140 ();
 sg13g2_decap_4 FILLER_23_147 ();
 sg13g2_fill_2 FILLER_23_151 ();
 sg13g2_decap_4 FILLER_23_218 ();
 sg13g2_fill_2 FILLER_23_222 ();
 sg13g2_decap_4 FILLER_23_232 ();
 sg13g2_fill_2 FILLER_23_246 ();
 sg13g2_fill_2 FILLER_23_251 ();
 sg13g2_fill_1 FILLER_23_253 ();
 sg13g2_fill_1 FILLER_23_258 ();
 sg13g2_fill_2 FILLER_23_293 ();
 sg13g2_fill_1 FILLER_23_316 ();
 sg13g2_fill_1 FILLER_23_339 ();
 sg13g2_fill_2 FILLER_23_344 ();
 sg13g2_fill_1 FILLER_23_346 ();
 sg13g2_fill_2 FILLER_23_381 ();
 sg13g2_fill_2 FILLER_23_386 ();
 sg13g2_fill_2 FILLER_23_396 ();
 sg13g2_fill_1 FILLER_23_398 ();
 sg13g2_fill_2 FILLER_23_407 ();
 sg13g2_fill_1 FILLER_23_409 ();
 sg13g2_fill_2 FILLER_23_419 ();
 sg13g2_fill_1 FILLER_23_429 ();
 sg13g2_decap_4 FILLER_24_0 ();
 sg13g2_fill_2 FILLER_24_4 ();
 sg13g2_fill_1 FILLER_24_21 ();
 sg13g2_fill_2 FILLER_24_38 ();
 sg13g2_fill_1 FILLER_24_52 ();
 sg13g2_decap_8 FILLER_24_57 ();
 sg13g2_decap_4 FILLER_24_64 ();
 sg13g2_fill_1 FILLER_24_68 ();
 sg13g2_fill_1 FILLER_24_77 ();
 sg13g2_fill_1 FILLER_24_87 ();
 sg13g2_decap_4 FILLER_24_101 ();
 sg13g2_decap_4 FILLER_24_113 ();
 sg13g2_fill_1 FILLER_24_117 ();
 sg13g2_decap_8 FILLER_24_122 ();
 sg13g2_decap_8 FILLER_24_138 ();
 sg13g2_fill_1 FILLER_24_149 ();
 sg13g2_fill_1 FILLER_24_158 ();
 sg13g2_fill_1 FILLER_24_176 ();
 sg13g2_fill_1 FILLER_24_181 ();
 sg13g2_fill_2 FILLER_24_192 ();
 sg13g2_fill_1 FILLER_24_197 ();
 sg13g2_fill_1 FILLER_24_202 ();
 sg13g2_fill_1 FILLER_24_233 ();
 sg13g2_fill_2 FILLER_24_258 ();
 sg13g2_decap_4 FILLER_24_265 ();
 sg13g2_fill_2 FILLER_24_274 ();
 sg13g2_decap_4 FILLER_24_280 ();
 sg13g2_fill_2 FILLER_24_292 ();
 sg13g2_fill_1 FILLER_24_294 ();
 sg13g2_fill_1 FILLER_24_299 ();
 sg13g2_decap_4 FILLER_24_309 ();
 sg13g2_fill_1 FILLER_24_337 ();
 sg13g2_decap_8 FILLER_24_343 ();
 sg13g2_decap_4 FILLER_24_350 ();
 sg13g2_fill_2 FILLER_24_380 ();
 sg13g2_fill_2 FILLER_24_396 ();
 sg13g2_fill_1 FILLER_24_398 ();
 sg13g2_fill_2 FILLER_24_428 ();
 sg13g2_decap_8 FILLER_25_0 ();
 sg13g2_fill_2 FILLER_25_7 ();
 sg13g2_fill_1 FILLER_25_23 ();
 sg13g2_fill_2 FILLER_25_28 ();
 sg13g2_fill_1 FILLER_25_30 ();
 sg13g2_fill_2 FILLER_25_46 ();
 sg13g2_decap_8 FILLER_25_57 ();
 sg13g2_fill_2 FILLER_25_64 ();
 sg13g2_fill_1 FILLER_25_75 ();
 sg13g2_fill_1 FILLER_25_84 ();
 sg13g2_fill_1 FILLER_25_94 ();
 sg13g2_fill_1 FILLER_25_107 ();
 sg13g2_fill_1 FILLER_25_127 ();
 sg13g2_fill_1 FILLER_25_131 ();
 sg13g2_fill_2 FILLER_25_137 ();
 sg13g2_decap_4 FILLER_25_151 ();
 sg13g2_fill_2 FILLER_25_155 ();
 sg13g2_fill_1 FILLER_25_170 ();
 sg13g2_fill_1 FILLER_25_200 ();
 sg13g2_decap_8 FILLER_25_206 ();
 sg13g2_decap_8 FILLER_25_213 ();
 sg13g2_fill_1 FILLER_25_220 ();
 sg13g2_decap_8 FILLER_25_226 ();
 sg13g2_fill_2 FILLER_25_233 ();
 sg13g2_fill_2 FILLER_25_246 ();
 sg13g2_fill_1 FILLER_25_248 ();
 sg13g2_decap_4 FILLER_25_261 ();
 sg13g2_decap_8 FILLER_25_294 ();
 sg13g2_decap_8 FILLER_25_301 ();
 sg13g2_decap_8 FILLER_25_308 ();
 sg13g2_fill_2 FILLER_25_315 ();
 sg13g2_fill_2 FILLER_25_325 ();
 sg13g2_fill_2 FILLER_25_332 ();
 sg13g2_fill_2 FILLER_25_338 ();
 sg13g2_fill_1 FILLER_25_340 ();
 sg13g2_fill_2 FILLER_25_360 ();
 sg13g2_fill_1 FILLER_25_362 ();
 sg13g2_fill_1 FILLER_25_372 ();
 sg13g2_fill_2 FILLER_25_376 ();
 sg13g2_decap_4 FILLER_25_383 ();
 sg13g2_decap_4 FILLER_25_413 ();
 sg13g2_fill_1 FILLER_25_417 ();
 sg13g2_decap_8 FILLER_25_423 ();
 sg13g2_decap_4 FILLER_26_0 ();
 sg13g2_fill_2 FILLER_26_8 ();
 sg13g2_fill_2 FILLER_26_14 ();
 sg13g2_decap_4 FILLER_26_35 ();
 sg13g2_fill_2 FILLER_26_39 ();
 sg13g2_decap_8 FILLER_26_48 ();
 sg13g2_fill_1 FILLER_26_65 ();
 sg13g2_fill_1 FILLER_26_100 ();
 sg13g2_fill_2 FILLER_26_115 ();
 sg13g2_fill_1 FILLER_26_117 ();
 sg13g2_fill_1 FILLER_26_130 ();
 sg13g2_fill_1 FILLER_26_140 ();
 sg13g2_fill_2 FILLER_26_154 ();
 sg13g2_decap_4 FILLER_26_169 ();
 sg13g2_fill_1 FILLER_26_173 ();
 sg13g2_decap_4 FILLER_26_195 ();
 sg13g2_fill_1 FILLER_26_199 ();
 sg13g2_decap_4 FILLER_26_249 ();
 sg13g2_fill_1 FILLER_26_271 ();
 sg13g2_fill_2 FILLER_26_277 ();
 sg13g2_fill_1 FILLER_26_295 ();
 sg13g2_fill_1 FILLER_26_322 ();
 sg13g2_fill_1 FILLER_26_349 ();
 sg13g2_fill_1 FILLER_26_361 ();
 sg13g2_fill_2 FILLER_26_370 ();
 sg13g2_fill_1 FILLER_26_372 ();
 sg13g2_decap_4 FILLER_26_386 ();
 sg13g2_decap_4 FILLER_26_395 ();
 sg13g2_fill_1 FILLER_26_399 ();
 sg13g2_fill_2 FILLER_27_0 ();
 sg13g2_fill_1 FILLER_27_12 ();
 sg13g2_fill_1 FILLER_27_18 ();
 sg13g2_fill_2 FILLER_27_23 ();
 sg13g2_fill_1 FILLER_27_25 ();
 sg13g2_fill_1 FILLER_27_30 ();
 sg13g2_fill_1 FILLER_27_39 ();
 sg13g2_fill_1 FILLER_27_71 ();
 sg13g2_fill_1 FILLER_27_77 ();
 sg13g2_fill_1 FILLER_27_82 ();
 sg13g2_fill_1 FILLER_27_88 ();
 sg13g2_decap_8 FILLER_27_93 ();
 sg13g2_fill_2 FILLER_27_117 ();
 sg13g2_fill_1 FILLER_27_131 ();
 sg13g2_decap_8 FILLER_27_137 ();
 sg13g2_fill_1 FILLER_27_144 ();
 sg13g2_fill_2 FILLER_27_155 ();
 sg13g2_fill_1 FILLER_27_182 ();
 sg13g2_fill_2 FILLER_27_186 ();
 sg13g2_fill_2 FILLER_27_193 ();
 sg13g2_decap_8 FILLER_27_199 ();
 sg13g2_decap_8 FILLER_27_214 ();
 sg13g2_decap_8 FILLER_27_221 ();
 sg13g2_decap_4 FILLER_27_228 ();
 sg13g2_fill_1 FILLER_27_255 ();
 sg13g2_fill_2 FILLER_27_274 ();
 sg13g2_fill_2 FILLER_27_279 ();
 sg13g2_fill_1 FILLER_27_281 ();
 sg13g2_fill_2 FILLER_27_287 ();
 sg13g2_fill_1 FILLER_27_289 ();
 sg13g2_decap_8 FILLER_27_295 ();
 sg13g2_fill_1 FILLER_27_302 ();
 sg13g2_fill_2 FILLER_27_307 ();
 sg13g2_fill_1 FILLER_27_309 ();
 sg13g2_decap_4 FILLER_27_318 ();
 sg13g2_fill_1 FILLER_27_322 ();
 sg13g2_fill_2 FILLER_27_333 ();
 sg13g2_fill_2 FILLER_27_339 ();
 sg13g2_fill_1 FILLER_27_341 ();
 sg13g2_decap_8 FILLER_27_346 ();
 sg13g2_decap_4 FILLER_27_353 ();
 sg13g2_fill_1 FILLER_27_357 ();
 sg13g2_decap_8 FILLER_27_367 ();
 sg13g2_decap_8 FILLER_27_404 ();
 sg13g2_fill_2 FILLER_27_411 ();
 sg13g2_fill_1 FILLER_27_422 ();
 sg13g2_fill_2 FILLER_27_428 ();
 sg13g2_fill_2 FILLER_28_0 ();
 sg13g2_fill_1 FILLER_28_12 ();
 sg13g2_fill_1 FILLER_28_18 ();
 sg13g2_decap_8 FILLER_28_31 ();
 sg13g2_decap_8 FILLER_28_38 ();
 sg13g2_fill_2 FILLER_28_45 ();
 sg13g2_fill_1 FILLER_28_47 ();
 sg13g2_decap_8 FILLER_28_57 ();
 sg13g2_fill_2 FILLER_28_64 ();
 sg13g2_fill_1 FILLER_28_66 ();
 sg13g2_fill_2 FILLER_28_75 ();
 sg13g2_decap_4 FILLER_28_82 ();
 sg13g2_decap_8 FILLER_28_94 ();
 sg13g2_decap_8 FILLER_28_101 ();
 sg13g2_decap_4 FILLER_28_136 ();
 sg13g2_decap_8 FILLER_28_148 ();
 sg13g2_fill_2 FILLER_28_155 ();
 sg13g2_fill_1 FILLER_28_157 ();
 sg13g2_decap_4 FILLER_28_167 ();
 sg13g2_fill_1 FILLER_28_181 ();
 sg13g2_fill_2 FILLER_28_187 ();
 sg13g2_fill_1 FILLER_28_189 ();
 sg13g2_fill_1 FILLER_28_195 ();
 sg13g2_decap_4 FILLER_28_222 ();
 sg13g2_fill_1 FILLER_28_226 ();
 sg13g2_fill_1 FILLER_28_237 ();
 sg13g2_decap_4 FILLER_28_280 ();
 sg13g2_fill_1 FILLER_28_284 ();
 sg13g2_decap_8 FILLER_28_302 ();
 sg13g2_fill_1 FILLER_28_313 ();
 sg13g2_fill_1 FILLER_28_319 ();
 sg13g2_fill_1 FILLER_28_360 ();
 sg13g2_fill_1 FILLER_28_377 ();
 sg13g2_fill_2 FILLER_28_386 ();
 sg13g2_fill_2 FILLER_28_397 ();
 sg13g2_decap_4 FILLER_29_0 ();
 sg13g2_fill_1 FILLER_29_10 ();
 sg13g2_fill_2 FILLER_29_19 ();
 sg13g2_fill_1 FILLER_29_21 ();
 sg13g2_fill_1 FILLER_29_26 ();
 sg13g2_fill_1 FILLER_29_36 ();
 sg13g2_decap_8 FILLER_29_48 ();
 sg13g2_fill_2 FILLER_29_55 ();
 sg13g2_decap_8 FILLER_29_61 ();
 sg13g2_fill_2 FILLER_29_68 ();
 sg13g2_fill_2 FILLER_29_82 ();
 sg13g2_fill_2 FILLER_29_102 ();
 sg13g2_fill_2 FILLER_29_117 ();
 sg13g2_fill_1 FILLER_29_119 ();
 sg13g2_fill_1 FILLER_29_125 ();
 sg13g2_decap_4 FILLER_29_137 ();
 sg13g2_fill_2 FILLER_29_159 ();
 sg13g2_decap_4 FILLER_29_170 ();
 sg13g2_decap_4 FILLER_29_200 ();
 sg13g2_decap_4 FILLER_29_208 ();
 sg13g2_fill_1 FILLER_29_225 ();
 sg13g2_fill_2 FILLER_29_257 ();
 sg13g2_fill_1 FILLER_29_271 ();
 sg13g2_fill_1 FILLER_29_279 ();
 sg13g2_fill_1 FILLER_29_295 ();
 sg13g2_fill_1 FILLER_29_321 ();
 sg13g2_decap_8 FILLER_29_352 ();
 sg13g2_decap_4 FILLER_29_359 ();
 sg13g2_fill_2 FILLER_29_363 ();
 sg13g2_decap_4 FILLER_29_383 ();
 sg13g2_fill_1 FILLER_29_404 ();
 sg13g2_fill_1 FILLER_29_409 ();
 sg13g2_fill_2 FILLER_29_428 ();
 sg13g2_decap_4 FILLER_30_4 ();
 sg13g2_fill_1 FILLER_30_8 ();
 sg13g2_fill_1 FILLER_30_18 ();
 sg13g2_fill_1 FILLER_30_23 ();
 sg13g2_fill_1 FILLER_30_29 ();
 sg13g2_fill_1 FILLER_30_34 ();
 sg13g2_fill_2 FILLER_30_39 ();
 sg13g2_decap_8 FILLER_30_49 ();
 sg13g2_fill_2 FILLER_30_56 ();
 sg13g2_decap_8 FILLER_30_63 ();
 sg13g2_fill_1 FILLER_30_83 ();
 sg13g2_fill_2 FILLER_30_103 ();
 sg13g2_fill_1 FILLER_30_105 ();
 sg13g2_fill_2 FILLER_30_140 ();
 sg13g2_fill_1 FILLER_30_161 ();
 sg13g2_fill_1 FILLER_30_176 ();
 sg13g2_fill_1 FILLER_30_180 ();
 sg13g2_decap_4 FILLER_30_190 ();
 sg13g2_fill_2 FILLER_30_199 ();
 sg13g2_decap_8 FILLER_30_215 ();
 sg13g2_decap_4 FILLER_30_222 ();
 sg13g2_fill_2 FILLER_30_226 ();
 sg13g2_decap_8 FILLER_30_232 ();
 sg13g2_decap_4 FILLER_30_239 ();
 sg13g2_fill_2 FILLER_30_243 ();
 sg13g2_decap_8 FILLER_30_253 ();
 sg13g2_fill_2 FILLER_30_264 ();
 sg13g2_fill_1 FILLER_30_266 ();
 sg13g2_fill_1 FILLER_30_304 ();
 sg13g2_decap_4 FILLER_30_310 ();
 sg13g2_fill_1 FILLER_30_318 ();
 sg13g2_fill_2 FILLER_30_331 ();
 sg13g2_fill_2 FILLER_30_337 ();
 sg13g2_fill_1 FILLER_30_339 ();
 sg13g2_decap_8 FILLER_30_344 ();
 sg13g2_fill_2 FILLER_30_351 ();
 sg13g2_fill_1 FILLER_30_353 ();
 sg13g2_fill_1 FILLER_30_376 ();
 sg13g2_fill_2 FILLER_30_381 ();
 sg13g2_fill_1 FILLER_30_388 ();
 sg13g2_fill_1 FILLER_30_400 ();
 sg13g2_fill_2 FILLER_30_414 ();
 sg13g2_fill_1 FILLER_30_416 ();
 sg13g2_fill_2 FILLER_31_26 ();
 sg13g2_fill_1 FILLER_31_28 ();
 sg13g2_fill_2 FILLER_31_52 ();
 sg13g2_fill_1 FILLER_31_54 ();
 sg13g2_fill_1 FILLER_31_59 ();
 sg13g2_fill_2 FILLER_31_71 ();
 sg13g2_fill_1 FILLER_31_73 ();
 sg13g2_fill_1 FILLER_31_82 ();
 sg13g2_fill_2 FILLER_31_93 ();
 sg13g2_fill_1 FILLER_31_95 ();
 sg13g2_fill_2 FILLER_31_108 ();
 sg13g2_fill_2 FILLER_31_123 ();
 sg13g2_fill_1 FILLER_31_133 ();
 sg13g2_fill_2 FILLER_31_139 ();
 sg13g2_decap_4 FILLER_31_151 ();
 sg13g2_fill_2 FILLER_31_173 ();
 sg13g2_decap_8 FILLER_31_189 ();
 sg13g2_fill_2 FILLER_31_196 ();
 sg13g2_fill_2 FILLER_31_224 ();
 sg13g2_fill_2 FILLER_31_264 ();
 sg13g2_fill_1 FILLER_31_266 ();
 sg13g2_fill_1 FILLER_31_271 ();
 sg13g2_fill_2 FILLER_31_275 ();
 sg13g2_decap_4 FILLER_31_282 ();
 sg13g2_fill_1 FILLER_31_286 ();
 sg13g2_fill_1 FILLER_31_295 ();
 sg13g2_fill_1 FILLER_31_363 ();
 sg13g2_fill_2 FILLER_31_372 ();
 sg13g2_fill_1 FILLER_31_374 ();
 sg13g2_fill_2 FILLER_31_383 ();
 sg13g2_fill_1 FILLER_31_385 ();
 sg13g2_decap_4 FILLER_32_20 ();
 sg13g2_fill_2 FILLER_32_24 ();
 sg13g2_decap_8 FILLER_32_31 ();
 sg13g2_decap_8 FILLER_32_38 ();
 sg13g2_decap_8 FILLER_32_45 ();
 sg13g2_decap_4 FILLER_32_60 ();
 sg13g2_fill_1 FILLER_32_83 ();
 sg13g2_fill_1 FILLER_32_129 ();
 sg13g2_fill_2 FILLER_32_138 ();
 sg13g2_fill_1 FILLER_32_140 ();
 sg13g2_decap_4 FILLER_32_158 ();
 sg13g2_fill_1 FILLER_32_162 ();
 sg13g2_fill_2 FILLER_32_176 ();
 sg13g2_fill_2 FILLER_32_192 ();
 sg13g2_fill_2 FILLER_32_229 ();
 sg13g2_fill_1 FILLER_32_231 ();
 sg13g2_fill_1 FILLER_32_263 ();
 sg13g2_fill_2 FILLER_32_272 ();
 sg13g2_decap_8 FILLER_32_282 ();
 sg13g2_fill_1 FILLER_32_289 ();
 sg13g2_fill_2 FILLER_32_298 ();
 sg13g2_decap_4 FILLER_32_308 ();
 sg13g2_fill_2 FILLER_32_312 ();
 sg13g2_fill_2 FILLER_32_331 ();
 sg13g2_decap_4 FILLER_32_342 ();
 sg13g2_fill_1 FILLER_32_346 ();
 sg13g2_fill_2 FILLER_32_351 ();
 sg13g2_fill_1 FILLER_32_353 ();
 sg13g2_fill_2 FILLER_32_360 ();
 sg13g2_fill_1 FILLER_32_369 ();
 sg13g2_fill_2 FILLER_32_379 ();
 sg13g2_fill_1 FILLER_32_381 ();
 sg13g2_fill_2 FILLER_32_399 ();
 sg13g2_fill_1 FILLER_32_401 ();
 sg13g2_decap_4 FILLER_32_415 ();
 sg13g2_fill_2 FILLER_32_427 ();
 sg13g2_fill_1 FILLER_32_429 ();
 sg13g2_fill_2 FILLER_33_0 ();
 sg13g2_fill_1 FILLER_33_2 ();
 sg13g2_fill_1 FILLER_33_7 ();
 sg13g2_fill_1 FILLER_33_12 ();
 sg13g2_fill_1 FILLER_33_18 ();
 sg13g2_fill_2 FILLER_33_24 ();
 sg13g2_fill_2 FILLER_33_34 ();
 sg13g2_decap_8 FILLER_33_44 ();
 sg13g2_fill_1 FILLER_33_70 ();
 sg13g2_fill_2 FILLER_33_79 ();
 sg13g2_decap_4 FILLER_33_127 ();
 sg13g2_decap_8 FILLER_33_136 ();
 sg13g2_decap_4 FILLER_33_143 ();
 sg13g2_fill_1 FILLER_33_147 ();
 sg13g2_fill_1 FILLER_33_193 ();
 sg13g2_fill_2 FILLER_33_198 ();
 sg13g2_fill_2 FILLER_33_205 ();
 sg13g2_fill_2 FILLER_33_213 ();
 sg13g2_fill_2 FILLER_33_219 ();
 sg13g2_fill_1 FILLER_33_221 ();
 sg13g2_fill_2 FILLER_33_227 ();
 sg13g2_fill_1 FILLER_33_229 ();
 sg13g2_fill_1 FILLER_33_241 ();
 sg13g2_decap_4 FILLER_33_246 ();
 sg13g2_fill_2 FILLER_33_250 ();
 sg13g2_fill_1 FILLER_33_257 ();
 sg13g2_fill_1 FILLER_33_263 ();
 sg13g2_fill_1 FILLER_33_284 ();
 sg13g2_fill_1 FILLER_33_296 ();
 sg13g2_fill_2 FILLER_33_302 ();
 sg13g2_fill_2 FILLER_33_309 ();
 sg13g2_decap_4 FILLER_33_315 ();
 sg13g2_fill_2 FILLER_33_350 ();
 sg13g2_fill_1 FILLER_33_352 ();
 sg13g2_fill_2 FILLER_33_379 ();
 sg13g2_fill_1 FILLER_33_389 ();
 sg13g2_fill_2 FILLER_33_395 ();
 sg13g2_fill_1 FILLER_33_402 ();
 sg13g2_fill_2 FILLER_33_408 ();
 sg13g2_fill_2 FILLER_33_415 ();
 sg13g2_decap_4 FILLER_33_424 ();
 sg13g2_fill_2 FILLER_33_428 ();
 sg13g2_fill_2 FILLER_34_39 ();
 sg13g2_fill_1 FILLER_34_54 ();
 sg13g2_decap_4 FILLER_34_60 ();
 sg13g2_fill_1 FILLER_34_81 ();
 sg13g2_fill_2 FILLER_34_100 ();
 sg13g2_fill_2 FILLER_34_127 ();
 sg13g2_fill_1 FILLER_34_134 ();
 sg13g2_fill_1 FILLER_34_148 ();
 sg13g2_fill_1 FILLER_34_163 ();
 sg13g2_fill_1 FILLER_34_179 ();
 sg13g2_fill_1 FILLER_34_188 ();
 sg13g2_fill_1 FILLER_34_192 ();
 sg13g2_fill_1 FILLER_34_199 ();
 sg13g2_decap_4 FILLER_34_240 ();
 sg13g2_fill_1 FILLER_34_244 ();
 sg13g2_decap_4 FILLER_34_271 ();
 sg13g2_fill_2 FILLER_34_283 ();
 sg13g2_fill_1 FILLER_34_299 ();
 sg13g2_fill_1 FILLER_34_326 ();
 sg13g2_fill_2 FILLER_34_332 ();
 sg13g2_fill_1 FILLER_34_360 ();
 sg13g2_fill_1 FILLER_34_370 ();
 sg13g2_decap_4 FILLER_34_384 ();
 sg13g2_decap_4 FILLER_35_0 ();
 sg13g2_fill_2 FILLER_35_4 ();
 sg13g2_decap_4 FILLER_35_10 ();
 sg13g2_fill_2 FILLER_35_18 ();
 sg13g2_fill_1 FILLER_35_20 ();
 sg13g2_fill_1 FILLER_35_30 ();
 sg13g2_fill_2 FILLER_35_38 ();
 sg13g2_decap_8 FILLER_35_45 ();
 sg13g2_fill_1 FILLER_35_52 ();
 sg13g2_fill_2 FILLER_35_60 ();
 sg13g2_fill_1 FILLER_35_62 ();
 sg13g2_fill_2 FILLER_35_67 ();
 sg13g2_fill_1 FILLER_35_80 ();
 sg13g2_decap_4 FILLER_35_84 ();
 sg13g2_fill_2 FILLER_35_97 ();
 sg13g2_fill_1 FILLER_35_99 ();
 sg13g2_fill_1 FILLER_35_108 ();
 sg13g2_fill_1 FILLER_35_146 ();
 sg13g2_fill_2 FILLER_35_161 ();
 sg13g2_fill_1 FILLER_35_175 ();
 sg13g2_decap_8 FILLER_35_188 ();
 sg13g2_decap_4 FILLER_35_195 ();
 sg13g2_fill_1 FILLER_35_199 ();
 sg13g2_fill_1 FILLER_35_213 ();
 sg13g2_fill_2 FILLER_35_220 ();
 sg13g2_fill_2 FILLER_35_228 ();
 sg13g2_fill_1 FILLER_35_230 ();
 sg13g2_decap_8 FILLER_35_239 ();
 sg13g2_decap_4 FILLER_35_246 ();
 sg13g2_fill_1 FILLER_35_250 ();
 sg13g2_decap_8 FILLER_35_260 ();
 sg13g2_decap_8 FILLER_35_267 ();
 sg13g2_fill_1 FILLER_35_274 ();
 sg13g2_fill_1 FILLER_35_283 ();
 sg13g2_fill_1 FILLER_35_295 ();
 sg13g2_fill_1 FILLER_35_313 ();
 sg13g2_fill_2 FILLER_35_318 ();
 sg13g2_fill_1 FILLER_35_320 ();
 sg13g2_fill_2 FILLER_35_325 ();
 sg13g2_fill_1 FILLER_35_332 ();
 sg13g2_fill_1 FILLER_35_337 ();
 sg13g2_fill_2 FILLER_35_350 ();
 sg13g2_fill_1 FILLER_35_403 ();
 sg13g2_fill_2 FILLER_35_416 ();
 sg13g2_fill_2 FILLER_36_11 ();
 sg13g2_fill_1 FILLER_36_13 ();
 sg13g2_decap_4 FILLER_36_25 ();
 sg13g2_fill_2 FILLER_36_29 ();
 sg13g2_fill_2 FILLER_36_46 ();
 sg13g2_fill_2 FILLER_36_51 ();
 sg13g2_decap_4 FILLER_36_58 ();
 sg13g2_fill_1 FILLER_36_62 ();
 sg13g2_decap_4 FILLER_36_74 ();
 sg13g2_decap_8 FILLER_36_83 ();
 sg13g2_decap_4 FILLER_36_90 ();
 sg13g2_fill_1 FILLER_36_94 ();
 sg13g2_fill_2 FILLER_36_99 ();
 sg13g2_fill_1 FILLER_36_104 ();
 sg13g2_fill_1 FILLER_36_108 ();
 sg13g2_decap_4 FILLER_36_114 ();
 sg13g2_fill_1 FILLER_36_118 ();
 sg13g2_decap_4 FILLER_36_142 ();
 sg13g2_fill_1 FILLER_36_159 ();
 sg13g2_fill_2 FILLER_36_164 ();
 sg13g2_fill_2 FILLER_36_170 ();
 sg13g2_fill_2 FILLER_36_176 ();
 sg13g2_decap_4 FILLER_36_183 ();
 sg13g2_fill_1 FILLER_36_187 ();
 sg13g2_fill_1 FILLER_36_218 ();
 sg13g2_fill_1 FILLER_36_251 ();
 sg13g2_fill_2 FILLER_36_288 ();
 sg13g2_fill_1 FILLER_36_290 ();
 sg13g2_fill_2 FILLER_36_295 ();
 sg13g2_fill_1 FILLER_36_327 ();
 sg13g2_fill_1 FILLER_36_332 ();
 sg13g2_fill_2 FILLER_36_337 ();
 sg13g2_fill_1 FILLER_36_342 ();
 sg13g2_fill_2 FILLER_36_358 ();
 sg13g2_fill_1 FILLER_36_360 ();
 sg13g2_fill_2 FILLER_36_365 ();
 sg13g2_fill_2 FILLER_36_375 ();
 sg13g2_fill_1 FILLER_36_383 ();
 sg13g2_fill_2 FILLER_36_388 ();
 sg13g2_fill_1 FILLER_36_398 ();
 sg13g2_fill_1 FILLER_37_31 ();
 sg13g2_fill_1 FILLER_37_37 ();
 sg13g2_decap_8 FILLER_37_55 ();
 sg13g2_fill_2 FILLER_37_62 ();
 sg13g2_fill_1 FILLER_37_64 ();
 sg13g2_fill_1 FILLER_37_69 ();
 sg13g2_decap_8 FILLER_37_75 ();
 sg13g2_fill_1 FILLER_37_86 ();
 sg13g2_fill_1 FILLER_37_113 ();
 sg13g2_fill_2 FILLER_37_118 ();
 sg13g2_fill_2 FILLER_37_125 ();
 sg13g2_fill_1 FILLER_37_131 ();
 sg13g2_fill_2 FILLER_37_156 ();
 sg13g2_fill_1 FILLER_37_158 ();
 sg13g2_decap_8 FILLER_37_189 ();
 sg13g2_fill_2 FILLER_37_196 ();
 sg13g2_decap_8 FILLER_37_202 ();
 sg13g2_fill_2 FILLER_37_212 ();
 sg13g2_fill_1 FILLER_37_248 ();
 sg13g2_decap_4 FILLER_37_253 ();
 sg13g2_fill_1 FILLER_37_257 ();
 sg13g2_decap_8 FILLER_37_262 ();
 sg13g2_fill_2 FILLER_37_269 ();
 sg13g2_fill_1 FILLER_37_271 ();
 sg13g2_decap_4 FILLER_37_297 ();
 sg13g2_fill_1 FILLER_37_301 ();
 sg13g2_decap_8 FILLER_37_318 ();
 sg13g2_fill_2 FILLER_37_325 ();
 sg13g2_fill_1 FILLER_37_327 ();
 sg13g2_fill_2 FILLER_37_354 ();
 sg13g2_fill_2 FILLER_37_385 ();
 sg13g2_fill_1 FILLER_37_396 ();
 sg13g2_decap_4 FILLER_37_407 ();
 sg13g2_fill_1 FILLER_37_411 ();
 sg13g2_decap_4 FILLER_37_416 ();
 sg13g2_decap_4 FILLER_37_424 ();
 sg13g2_fill_2 FILLER_37_428 ();
 sg13g2_fill_2 FILLER_38_0 ();
 sg13g2_fill_1 FILLER_38_2 ();
 sg13g2_fill_1 FILLER_38_11 ();
 sg13g2_fill_1 FILLER_38_18 ();
 sg13g2_fill_2 FILLER_38_23 ();
 sg13g2_fill_2 FILLER_38_33 ();
 sg13g2_fill_2 FILLER_38_38 ();
 sg13g2_fill_1 FILLER_38_49 ();
 sg13g2_decap_4 FILLER_38_66 ();
 sg13g2_fill_2 FILLER_38_70 ();
 sg13g2_decap_4 FILLER_38_81 ();
 sg13g2_fill_2 FILLER_38_85 ();
 sg13g2_fill_2 FILLER_38_92 ();
 sg13g2_decap_8 FILLER_38_98 ();
 sg13g2_fill_2 FILLER_38_113 ();
 sg13g2_fill_1 FILLER_38_115 ();
 sg13g2_fill_2 FILLER_38_124 ();
 sg13g2_fill_1 FILLER_38_126 ();
 sg13g2_fill_2 FILLER_38_132 ();
 sg13g2_fill_1 FILLER_38_134 ();
 sg13g2_fill_2 FILLER_38_143 ();
 sg13g2_fill_1 FILLER_38_145 ();
 sg13g2_decap_4 FILLER_38_155 ();
 sg13g2_fill_1 FILLER_38_159 ();
 sg13g2_fill_2 FILLER_38_164 ();
 sg13g2_fill_1 FILLER_38_166 ();
 sg13g2_decap_4 FILLER_38_172 ();
 sg13g2_fill_2 FILLER_38_176 ();
 sg13g2_decap_8 FILLER_38_183 ();
 sg13g2_decap_4 FILLER_38_190 ();
 sg13g2_fill_1 FILLER_38_194 ();
 sg13g2_fill_2 FILLER_38_207 ();
 sg13g2_fill_2 FILLER_38_215 ();
 sg13g2_decap_8 FILLER_38_230 ();
 sg13g2_fill_2 FILLER_38_237 ();
 sg13g2_fill_1 FILLER_38_239 ();
 sg13g2_fill_2 FILLER_38_295 ();
 sg13g2_fill_1 FILLER_38_328 ();
 sg13g2_decap_4 FILLER_38_338 ();
 sg13g2_decap_4 FILLER_39_31 ();
 sg13g2_fill_2 FILLER_39_35 ();
 sg13g2_fill_2 FILLER_39_57 ();
 sg13g2_fill_1 FILLER_39_59 ();
 sg13g2_fill_2 FILLER_39_74 ();
 sg13g2_fill_2 FILLER_39_87 ();
 sg13g2_decap_4 FILLER_39_99 ();
 sg13g2_fill_2 FILLER_39_148 ();
 sg13g2_fill_2 FILLER_39_159 ();
 sg13g2_decap_8 FILLER_39_177 ();
 sg13g2_decap_8 FILLER_39_184 ();
 sg13g2_fill_2 FILLER_39_208 ();
 sg13g2_fill_1 FILLER_39_210 ();
 sg13g2_decap_4 FILLER_39_220 ();
 sg13g2_decap_8 FILLER_39_229 ();
 sg13g2_fill_1 FILLER_39_236 ();
 sg13g2_fill_2 FILLER_39_243 ();
 sg13g2_fill_1 FILLER_39_245 ();
 sg13g2_decap_8 FILLER_39_254 ();
 sg13g2_decap_8 FILLER_39_261 ();
 sg13g2_decap_4 FILLER_39_268 ();
 sg13g2_fill_2 FILLER_39_272 ();
 sg13g2_fill_2 FILLER_39_290 ();
 sg13g2_fill_1 FILLER_39_292 ();
 sg13g2_decap_4 FILLER_39_303 ();
 sg13g2_fill_1 FILLER_39_307 ();
 sg13g2_fill_1 FILLER_39_312 ();
 sg13g2_decap_8 FILLER_39_317 ();
 sg13g2_fill_2 FILLER_39_324 ();
 sg13g2_fill_1 FILLER_39_357 ();
 sg13g2_fill_2 FILLER_39_375 ();
 sg13g2_decap_4 FILLER_39_386 ();
 sg13g2_decap_8 FILLER_39_403 ();
 sg13g2_fill_2 FILLER_39_410 ();
 sg13g2_fill_1 FILLER_39_412 ();
 sg13g2_fill_2 FILLER_39_417 ();
 sg13g2_fill_1 FILLER_39_423 ();
 sg13g2_fill_2 FILLER_39_428 ();
 sg13g2_decap_8 FILLER_40_0 ();
 sg13g2_fill_1 FILLER_40_7 ();
 sg13g2_decap_4 FILLER_40_12 ();
 sg13g2_fill_2 FILLER_40_16 ();
 sg13g2_decap_4 FILLER_40_23 ();
 sg13g2_fill_1 FILLER_40_27 ();
 sg13g2_decap_4 FILLER_40_32 ();
 sg13g2_fill_2 FILLER_40_36 ();
 sg13g2_fill_1 FILLER_40_61 ();
 sg13g2_fill_2 FILLER_40_71 ();
 sg13g2_fill_1 FILLER_40_73 ();
 sg13g2_fill_1 FILLER_40_79 ();
 sg13g2_fill_1 FILLER_40_85 ();
 sg13g2_fill_1 FILLER_40_90 ();
 sg13g2_fill_2 FILLER_40_96 ();
 sg13g2_fill_2 FILLER_40_111 ();
 sg13g2_decap_4 FILLER_40_117 ();
 sg13g2_decap_4 FILLER_40_126 ();
 sg13g2_fill_1 FILLER_40_159 ();
 sg13g2_decap_4 FILLER_40_168 ();
 sg13g2_fill_1 FILLER_40_172 ();
 sg13g2_fill_2 FILLER_40_176 ();
 sg13g2_fill_1 FILLER_40_178 ();
 sg13g2_decap_4 FILLER_40_185 ();
 sg13g2_fill_1 FILLER_40_189 ();
 sg13g2_fill_1 FILLER_40_217 ();
 sg13g2_fill_1 FILLER_40_222 ();
 sg13g2_fill_1 FILLER_40_226 ();
 sg13g2_fill_1 FILLER_40_231 ();
 sg13g2_fill_1 FILLER_40_237 ();
 sg13g2_decap_8 FILLER_40_264 ();
 sg13g2_fill_2 FILLER_40_276 ();
 sg13g2_fill_2 FILLER_40_291 ();
 sg13g2_fill_1 FILLER_40_301 ();
 sg13g2_decap_8 FILLER_40_328 ();
 sg13g2_fill_1 FILLER_40_335 ();
 sg13g2_decap_8 FILLER_40_343 ();
 sg13g2_fill_2 FILLER_40_350 ();
 sg13g2_fill_1 FILLER_40_352 ();
 sg13g2_fill_1 FILLER_40_364 ();
 sg13g2_decap_8 FILLER_40_382 ();
 sg13g2_fill_1 FILLER_40_389 ();
 sg13g2_fill_2 FILLER_40_400 ();
 sg13g2_fill_2 FILLER_40_427 ();
 sg13g2_fill_1 FILLER_40_429 ();
 sg13g2_fill_1 FILLER_41_0 ();
 sg13g2_fill_1 FILLER_41_5 ();
 sg13g2_fill_1 FILLER_41_36 ();
 sg13g2_decap_8 FILLER_41_46 ();
 sg13g2_decap_4 FILLER_41_60 ();
 sg13g2_fill_1 FILLER_41_74 ();
 sg13g2_fill_1 FILLER_41_83 ();
 sg13g2_fill_1 FILLER_41_88 ();
 sg13g2_fill_2 FILLER_41_102 ();
 sg13g2_fill_1 FILLER_41_104 ();
 sg13g2_decap_8 FILLER_41_121 ();
 sg13g2_fill_1 FILLER_41_137 ();
 sg13g2_fill_2 FILLER_41_141 ();
 sg13g2_fill_2 FILLER_41_148 ();
 sg13g2_fill_2 FILLER_41_153 ();
 sg13g2_decap_4 FILLER_41_164 ();
 sg13g2_fill_1 FILLER_41_168 ();
 sg13g2_fill_2 FILLER_41_173 ();
 sg13g2_fill_1 FILLER_41_175 ();
 sg13g2_fill_2 FILLER_41_184 ();
 sg13g2_fill_1 FILLER_41_186 ();
 sg13g2_decap_4 FILLER_41_193 ();
 sg13g2_fill_1 FILLER_41_197 ();
 sg13g2_fill_1 FILLER_41_214 ();
 sg13g2_fill_2 FILLER_41_222 ();
 sg13g2_fill_1 FILLER_41_224 ();
 sg13g2_fill_2 FILLER_41_234 ();
 sg13g2_fill_1 FILLER_41_236 ();
 sg13g2_fill_2 FILLER_41_246 ();
 sg13g2_fill_1 FILLER_41_248 ();
 sg13g2_fill_2 FILLER_41_292 ();
 sg13g2_fill_1 FILLER_41_294 ();
 sg13g2_fill_2 FILLER_41_300 ();
 sg13g2_fill_1 FILLER_41_312 ();
 sg13g2_decap_4 FILLER_41_317 ();
 sg13g2_fill_2 FILLER_41_321 ();
 sg13g2_decap_4 FILLER_41_328 ();
 sg13g2_decap_8 FILLER_41_350 ();
 sg13g2_decap_4 FILLER_41_357 ();
 sg13g2_fill_1 FILLER_41_361 ();
 sg13g2_decap_4 FILLER_41_383 ();
 sg13g2_fill_1 FILLER_41_387 ();
 sg13g2_decap_4 FILLER_41_405 ();
 sg13g2_fill_1 FILLER_41_409 ();
 sg13g2_decap_4 FILLER_42_0 ();
 sg13g2_fill_1 FILLER_42_4 ();
 sg13g2_decap_8 FILLER_42_18 ();
 sg13g2_decap_4 FILLER_42_25 ();
 sg13g2_fill_2 FILLER_42_29 ();
 sg13g2_decap_4 FILLER_42_35 ();
 sg13g2_fill_2 FILLER_42_50 ();
 sg13g2_decap_4 FILLER_42_92 ();
 sg13g2_fill_2 FILLER_42_108 ();
 sg13g2_fill_1 FILLER_42_110 ();
 sg13g2_fill_2 FILLER_42_117 ();
 sg13g2_fill_1 FILLER_42_119 ();
 sg13g2_fill_2 FILLER_42_128 ();
 sg13g2_decap_4 FILLER_42_139 ();
 sg13g2_fill_2 FILLER_42_143 ();
 sg13g2_fill_1 FILLER_42_161 ();
 sg13g2_fill_2 FILLER_42_167 ();
 sg13g2_fill_1 FILLER_42_214 ();
 sg13g2_fill_2 FILLER_42_224 ();
 sg13g2_fill_1 FILLER_42_238 ();
 sg13g2_fill_2 FILLER_42_243 ();
 sg13g2_fill_1 FILLER_42_253 ();
 sg13g2_fill_2 FILLER_42_258 ();
 sg13g2_decap_8 FILLER_42_264 ();
 sg13g2_fill_1 FILLER_42_271 ();
 sg13g2_fill_1 FILLER_42_275 ();
 sg13g2_fill_1 FILLER_42_281 ();
 sg13g2_fill_2 FILLER_42_290 ();
 sg13g2_fill_2 FILLER_42_300 ();
 sg13g2_fill_2 FILLER_42_307 ();
 sg13g2_fill_1 FILLER_42_309 ();
 sg13g2_fill_2 FILLER_42_318 ();
 sg13g2_fill_1 FILLER_42_320 ();
 sg13g2_fill_2 FILLER_42_359 ();
 sg13g2_fill_1 FILLER_42_361 ();
 sg13g2_decap_8 FILLER_42_370 ();
 sg13g2_decap_4 FILLER_42_377 ();
 sg13g2_decap_4 FILLER_42_394 ();
 sg13g2_decap_8 FILLER_42_411 ();
 sg13g2_fill_2 FILLER_42_418 ();
 sg13g2_fill_2 FILLER_42_428 ();
 sg13g2_decap_8 FILLER_43_0 ();
 sg13g2_decap_8 FILLER_43_7 ();
 sg13g2_fill_2 FILLER_43_14 ();
 sg13g2_fill_1 FILLER_43_16 ();
 sg13g2_fill_2 FILLER_43_47 ();
 sg13g2_decap_4 FILLER_43_53 ();
 sg13g2_fill_2 FILLER_43_78 ();
 sg13g2_fill_1 FILLER_43_80 ();
 sg13g2_decap_8 FILLER_43_86 ();
 sg13g2_fill_2 FILLER_43_97 ();
 sg13g2_fill_1 FILLER_43_99 ();
 sg13g2_fill_2 FILLER_43_127 ();
 sg13g2_decap_4 FILLER_43_133 ();
 sg13g2_fill_2 FILLER_43_140 ();
 sg13g2_fill_2 FILLER_43_191 ();
 sg13g2_fill_1 FILLER_43_193 ();
 sg13g2_fill_1 FILLER_43_233 ();
 sg13g2_fill_1 FILLER_43_269 ();
 sg13g2_fill_2 FILLER_43_278 ();
 sg13g2_fill_1 FILLER_43_292 ();
 sg13g2_fill_2 FILLER_43_300 ();
 sg13g2_fill_1 FILLER_43_302 ();
 sg13g2_fill_2 FILLER_43_311 ();
 sg13g2_decap_4 FILLER_43_319 ();
 sg13g2_fill_1 FILLER_43_328 ();
 sg13g2_fill_1 FILLER_43_333 ();
 sg13g2_fill_1 FILLER_43_337 ();
 sg13g2_fill_1 FILLER_43_369 ();
 sg13g2_fill_1 FILLER_43_375 ();
 sg13g2_decap_4 FILLER_43_391 ();
 sg13g2_fill_2 FILLER_43_418 ();
 sg13g2_fill_2 FILLER_43_428 ();
 sg13g2_decap_8 FILLER_44_0 ();
 sg13g2_decap_8 FILLER_44_7 ();
 sg13g2_fill_2 FILLER_44_14 ();
 sg13g2_fill_2 FILLER_44_33 ();
 sg13g2_fill_1 FILLER_44_59 ();
 sg13g2_decap_8 FILLER_44_73 ();
 sg13g2_decap_4 FILLER_44_80 ();
 sg13g2_fill_2 FILLER_44_98 ();
 sg13g2_fill_1 FILLER_44_113 ();
 sg13g2_fill_2 FILLER_44_117 ();
 sg13g2_fill_2 FILLER_44_125 ();
 sg13g2_fill_2 FILLER_44_181 ();
 sg13g2_fill_1 FILLER_44_183 ();
 sg13g2_decap_4 FILLER_44_214 ();
 sg13g2_fill_2 FILLER_44_218 ();
 sg13g2_decap_8 FILLER_44_243 ();
 sg13g2_fill_2 FILLER_44_276 ();
 sg13g2_fill_1 FILLER_44_290 ();
 sg13g2_fill_2 FILLER_44_303 ();
 sg13g2_fill_1 FILLER_44_310 ();
 sg13g2_decap_8 FILLER_44_320 ();
 sg13g2_decap_4 FILLER_44_327 ();
 sg13g2_fill_1 FILLER_44_331 ();
 sg13g2_fill_1 FILLER_44_340 ();
 sg13g2_fill_1 FILLER_44_345 ();
 sg13g2_fill_2 FILLER_44_349 ();
 sg13g2_decap_4 FILLER_44_359 ();
 sg13g2_fill_2 FILLER_44_363 ();
 sg13g2_decap_8 FILLER_44_383 ();
 sg13g2_fill_1 FILLER_44_390 ();
 sg13g2_fill_1 FILLER_44_396 ();
 sg13g2_decap_4 FILLER_44_407 ();
 sg13g2_fill_2 FILLER_44_416 ();
 sg13g2_fill_1 FILLER_44_418 ();
 sg13g2_fill_2 FILLER_44_427 ();
 sg13g2_fill_1 FILLER_44_429 ();
 sg13g2_fill_1 FILLER_45_18 ();
 sg13g2_decap_4 FILLER_45_49 ();
 sg13g2_fill_1 FILLER_45_58 ();
 sg13g2_decap_4 FILLER_45_67 ();
 sg13g2_fill_2 FILLER_45_71 ();
 sg13g2_fill_2 FILLER_45_91 ();
 sg13g2_fill_1 FILLER_45_93 ();
 sg13g2_fill_2 FILLER_45_99 ();
 sg13g2_fill_1 FILLER_45_111 ();
 sg13g2_decap_4 FILLER_45_124 ();
 sg13g2_fill_1 FILLER_45_136 ();
 sg13g2_fill_2 FILLER_45_141 ();
 sg13g2_fill_2 FILLER_45_148 ();
 sg13g2_fill_1 FILLER_45_160 ();
 sg13g2_fill_1 FILLER_45_174 ();
 sg13g2_fill_1 FILLER_45_184 ();
 sg13g2_fill_1 FILLER_45_190 ();
 sg13g2_decap_4 FILLER_45_217 ();
 sg13g2_fill_1 FILLER_45_221 ();
 sg13g2_fill_1 FILLER_45_227 ();
 sg13g2_fill_2 FILLER_45_258 ();
 sg13g2_decap_4 FILLER_45_279 ();
 sg13g2_fill_1 FILLER_45_287 ();
 sg13g2_decap_8 FILLER_45_301 ();
 sg13g2_decap_8 FILLER_45_316 ();
 sg13g2_fill_2 FILLER_45_328 ();
 sg13g2_decap_8 FILLER_45_339 ();
 sg13g2_decap_8 FILLER_45_346 ();
 sg13g2_decap_8 FILLER_45_353 ();
 sg13g2_fill_2 FILLER_45_364 ();
 sg13g2_fill_1 FILLER_45_377 ();
 sg13g2_fill_2 FILLER_45_384 ();
 sg13g2_decap_4 FILLER_45_395 ();
 sg13g2_decap_4 FILLER_46_0 ();
 sg13g2_fill_1 FILLER_46_4 ();
 sg13g2_decap_8 FILLER_46_35 ();
 sg13g2_decap_4 FILLER_46_42 ();
 sg13g2_fill_1 FILLER_46_46 ();
 sg13g2_fill_1 FILLER_46_77 ();
 sg13g2_fill_2 FILLER_46_91 ();
 sg13g2_fill_1 FILLER_46_93 ();
 sg13g2_decap_4 FILLER_46_106 ();
 sg13g2_fill_2 FILLER_46_110 ();
 sg13g2_fill_1 FILLER_46_134 ();
 sg13g2_fill_2 FILLER_46_145 ();
 sg13g2_fill_1 FILLER_46_147 ();
 sg13g2_fill_2 FILLER_46_156 ();
 sg13g2_fill_1 FILLER_46_158 ();
 sg13g2_fill_1 FILLER_46_164 ();
 sg13g2_fill_2 FILLER_46_170 ();
 sg13g2_fill_1 FILLER_46_172 ();
 sg13g2_fill_1 FILLER_46_185 ();
 sg13g2_decap_8 FILLER_46_212 ();
 sg13g2_fill_2 FILLER_46_219 ();
 sg13g2_fill_1 FILLER_46_221 ();
 sg13g2_decap_8 FILLER_46_239 ();
 sg13g2_fill_2 FILLER_46_249 ();
 sg13g2_fill_1 FILLER_46_251 ();
 sg13g2_decap_8 FILLER_46_282 ();
 sg13g2_fill_2 FILLER_46_289 ();
 sg13g2_fill_2 FILLER_46_413 ();
 sg13g2_decap_4 FILLER_46_424 ();
 sg13g2_fill_2 FILLER_46_428 ();
 sg13g2_decap_4 FILLER_47_0 ();
 sg13g2_fill_2 FILLER_47_4 ();
 sg13g2_fill_2 FILLER_47_24 ();
 sg13g2_fill_1 FILLER_47_26 ();
 sg13g2_decap_4 FILLER_47_33 ();
 sg13g2_fill_1 FILLER_47_42 ();
 sg13g2_fill_2 FILLER_47_47 ();
 sg13g2_fill_1 FILLER_47_49 ();
 sg13g2_fill_2 FILLER_47_53 ();
 sg13g2_fill_2 FILLER_47_60 ();
 sg13g2_fill_1 FILLER_47_62 ();
 sg13g2_fill_2 FILLER_47_68 ();
 sg13g2_fill_1 FILLER_47_70 ();
 sg13g2_fill_2 FILLER_47_75 ();
 sg13g2_fill_1 FILLER_47_114 ();
 sg13g2_decap_4 FILLER_47_135 ();
 sg13g2_fill_1 FILLER_47_139 ();
 sg13g2_fill_1 FILLER_47_151 ();
 sg13g2_fill_1 FILLER_47_157 ();
 sg13g2_fill_1 FILLER_47_167 ();
 sg13g2_decap_4 FILLER_47_172 ();
 sg13g2_decap_4 FILLER_47_180 ();
 sg13g2_fill_1 FILLER_47_184 ();
 sg13g2_fill_2 FILLER_47_190 ();
 sg13g2_fill_1 FILLER_47_192 ();
 sg13g2_fill_1 FILLER_47_197 ();
 sg13g2_fill_2 FILLER_47_204 ();
 sg13g2_fill_1 FILLER_47_206 ();
 sg13g2_fill_2 FILLER_47_211 ();
 sg13g2_decap_4 FILLER_47_217 ();
 sg13g2_fill_1 FILLER_47_221 ();
 sg13g2_fill_2 FILLER_47_247 ();
 sg13g2_fill_2 FILLER_47_294 ();
 sg13g2_fill_2 FILLER_47_301 ();
 sg13g2_fill_2 FILLER_47_308 ();
 sg13g2_fill_1 FILLER_47_310 ();
 sg13g2_decap_8 FILLER_47_315 ();
 sg13g2_decap_8 FILLER_47_322 ();
 sg13g2_fill_2 FILLER_47_329 ();
 sg13g2_decap_8 FILLER_47_335 ();
 sg13g2_fill_1 FILLER_47_378 ();
 sg13g2_fill_1 FILLER_47_384 ();
 sg13g2_fill_1 FILLER_47_390 ();
 sg13g2_fill_1 FILLER_47_397 ();
 sg13g2_fill_2 FILLER_47_402 ();
 sg13g2_decap_4 FILLER_48_0 ();
 sg13g2_fill_2 FILLER_48_4 ();
 sg13g2_decap_4 FILLER_48_15 ();
 sg13g2_decap_4 FILLER_48_29 ();
 sg13g2_fill_1 FILLER_48_62 ();
 sg13g2_decap_4 FILLER_48_81 ();
 sg13g2_fill_1 FILLER_48_85 ();
 sg13g2_fill_1 FILLER_48_90 ();
 sg13g2_fill_2 FILLER_48_99 ();
 sg13g2_fill_1 FILLER_48_101 ();
 sg13g2_fill_1 FILLER_48_110 ();
 sg13g2_decap_4 FILLER_48_116 ();
 sg13g2_fill_2 FILLER_48_120 ();
 sg13g2_fill_2 FILLER_48_129 ();
 sg13g2_fill_1 FILLER_48_131 ();
 sg13g2_decap_4 FILLER_48_135 ();
 sg13g2_fill_1 FILLER_48_139 ();
 sg13g2_fill_2 FILLER_48_148 ();
 sg13g2_fill_2 FILLER_48_158 ();
 sg13g2_fill_1 FILLER_48_160 ();
 sg13g2_decap_8 FILLER_48_169 ();
 sg13g2_fill_1 FILLER_48_176 ();
 sg13g2_fill_1 FILLER_48_180 ();
 sg13g2_fill_2 FILLER_48_212 ();
 sg13g2_fill_2 FILLER_48_253 ();
 sg13g2_decap_8 FILLER_48_272 ();
 sg13g2_decap_4 FILLER_48_279 ();
 sg13g2_fill_1 FILLER_48_295 ();
 sg13g2_fill_1 FILLER_48_330 ();
 sg13g2_decap_8 FILLER_48_360 ();
 sg13g2_fill_1 FILLER_48_378 ();
 sg13g2_fill_1 FILLER_48_405 ();
 sg13g2_fill_1 FILLER_48_411 ();
 sg13g2_fill_1 FILLER_48_418 ();
 sg13g2_fill_2 FILLER_48_428 ();
 sg13g2_fill_2 FILLER_49_5 ();
 sg13g2_fill_1 FILLER_49_7 ();
 sg13g2_fill_1 FILLER_49_13 ();
 sg13g2_fill_1 FILLER_49_29 ();
 sg13g2_fill_2 FILLER_49_36 ();
 sg13g2_fill_1 FILLER_49_38 ();
 sg13g2_decap_8 FILLER_49_43 ();
 sg13g2_decap_8 FILLER_49_50 ();
 sg13g2_decap_8 FILLER_49_77 ();
 sg13g2_fill_2 FILLER_49_84 ();
 sg13g2_fill_1 FILLER_49_86 ();
 sg13g2_fill_2 FILLER_49_104 ();
 sg13g2_fill_1 FILLER_49_115 ();
 sg13g2_fill_1 FILLER_49_139 ();
 sg13g2_fill_1 FILLER_49_145 ();
 sg13g2_fill_1 FILLER_49_151 ();
 sg13g2_fill_1 FILLER_49_160 ();
 sg13g2_fill_2 FILLER_49_165 ();
 sg13g2_fill_1 FILLER_49_167 ();
 sg13g2_fill_2 FILLER_49_199 ();
 sg13g2_decap_8 FILLER_49_204 ();
 sg13g2_fill_1 FILLER_49_211 ();
 sg13g2_fill_2 FILLER_49_219 ();
 sg13g2_fill_1 FILLER_49_242 ();
 sg13g2_fill_1 FILLER_49_251 ();
 sg13g2_fill_1 FILLER_49_267 ();
 sg13g2_decap_4 FILLER_49_275 ();
 sg13g2_fill_2 FILLER_49_279 ();
 sg13g2_fill_1 FILLER_49_289 ();
 sg13g2_fill_1 FILLER_49_295 ();
 sg13g2_decap_4 FILLER_49_309 ();
 sg13g2_decap_8 FILLER_49_317 ();
 sg13g2_decap_8 FILLER_49_324 ();
 sg13g2_fill_2 FILLER_49_331 ();
 sg13g2_fill_2 FILLER_49_338 ();
 sg13g2_fill_1 FILLER_49_340 ();
 sg13g2_fill_2 FILLER_49_348 ();
 sg13g2_fill_1 FILLER_49_362 ();
 sg13g2_fill_2 FILLER_49_367 ();
 sg13g2_fill_1 FILLER_49_369 ();
 sg13g2_fill_2 FILLER_49_375 ();
 sg13g2_fill_1 FILLER_49_381 ();
 sg13g2_fill_2 FILLER_49_388 ();
 sg13g2_fill_2 FILLER_49_395 ();
 sg13g2_fill_2 FILLER_49_402 ();
 sg13g2_decap_4 FILLER_50_0 ();
 sg13g2_fill_2 FILLER_50_4 ();
 sg13g2_decap_8 FILLER_50_14 ();
 sg13g2_decap_8 FILLER_50_21 ();
 sg13g2_fill_1 FILLER_50_28 ();
 sg13g2_fill_2 FILLER_50_34 ();
 sg13g2_fill_2 FILLER_50_40 ();
 sg13g2_fill_1 FILLER_50_42 ();
 sg13g2_decap_4 FILLER_50_47 ();
 sg13g2_fill_1 FILLER_50_51 ();
 sg13g2_fill_2 FILLER_50_65 ();
 sg13g2_fill_1 FILLER_50_73 ();
 sg13g2_decap_4 FILLER_50_78 ();
 sg13g2_fill_1 FILLER_50_82 ();
 sg13g2_fill_1 FILLER_50_133 ();
 sg13g2_fill_2 FILLER_50_147 ();
 sg13g2_fill_1 FILLER_50_149 ();
 sg13g2_decap_4 FILLER_50_176 ();
 sg13g2_decap_8 FILLER_50_190 ();
 sg13g2_decap_8 FILLER_50_197 ();
 sg13g2_decap_8 FILLER_50_204 ();
 sg13g2_decap_4 FILLER_50_211 ();
 sg13g2_fill_2 FILLER_50_215 ();
 sg13g2_decap_8 FILLER_50_256 ();
 sg13g2_decap_4 FILLER_50_263 ();
 sg13g2_fill_1 FILLER_50_280 ();
 sg13g2_decap_8 FILLER_50_308 ();
 sg13g2_fill_2 FILLER_50_315 ();
 sg13g2_fill_2 FILLER_50_343 ();
 sg13g2_fill_1 FILLER_50_345 ();
 sg13g2_decap_4 FILLER_50_350 ();
 sg13g2_fill_2 FILLER_50_354 ();
 sg13g2_fill_1 FILLER_50_364 ();
 sg13g2_decap_8 FILLER_50_416 ();
 sg13g2_fill_2 FILLER_50_427 ();
 sg13g2_fill_1 FILLER_50_429 ();
 sg13g2_fill_1 FILLER_51_0 ();
 sg13g2_fill_1 FILLER_51_14 ();
 sg13g2_fill_2 FILLER_51_31 ();
 sg13g2_fill_1 FILLER_51_33 ();
 sg13g2_decap_4 FILLER_51_42 ();
 sg13g2_fill_1 FILLER_51_46 ();
 sg13g2_decap_4 FILLER_51_51 ();
 sg13g2_fill_2 FILLER_51_68 ();
 sg13g2_fill_1 FILLER_51_70 ();
 sg13g2_decap_8 FILLER_51_84 ();
 sg13g2_fill_1 FILLER_51_91 ();
 sg13g2_decap_4 FILLER_51_100 ();
 sg13g2_fill_2 FILLER_51_109 ();
 sg13g2_fill_1 FILLER_51_111 ();
 sg13g2_decap_4 FILLER_51_134 ();
 sg13g2_fill_2 FILLER_51_138 ();
 sg13g2_fill_2 FILLER_51_150 ();
 sg13g2_decap_4 FILLER_51_157 ();
 sg13g2_fill_1 FILLER_51_165 ();
 sg13g2_fill_1 FILLER_51_174 ();
 sg13g2_fill_1 FILLER_51_183 ();
 sg13g2_fill_1 FILLER_51_214 ();
 sg13g2_fill_1 FILLER_51_223 ();
 sg13g2_fill_1 FILLER_51_228 ();
 sg13g2_fill_1 FILLER_51_234 ();
 sg13g2_fill_1 FILLER_51_254 ();
 sg13g2_fill_2 FILLER_51_260 ();
 sg13g2_fill_1 FILLER_51_262 ();
 sg13g2_fill_2 FILLER_51_272 ();
 sg13g2_fill_1 FILLER_51_290 ();
 sg13g2_fill_1 FILLER_51_298 ();
 sg13g2_fill_1 FILLER_51_325 ();
 sg13g2_decap_4 FILLER_51_330 ();
 sg13g2_fill_1 FILLER_51_334 ();
 sg13g2_decap_4 FILLER_51_339 ();
 sg13g2_decap_4 FILLER_51_351 ();
 sg13g2_fill_2 FILLER_51_355 ();
 sg13g2_decap_4 FILLER_51_378 ();
 sg13g2_fill_2 FILLER_51_392 ();
 sg13g2_decap_8 FILLER_52_0 ();
 sg13g2_fill_1 FILLER_52_7 ();
 sg13g2_fill_1 FILLER_52_19 ();
 sg13g2_fill_1 FILLER_52_34 ();
 sg13g2_fill_2 FILLER_52_40 ();
 sg13g2_fill_1 FILLER_52_42 ();
 sg13g2_fill_1 FILLER_52_48 ();
 sg13g2_fill_1 FILLER_52_54 ();
 sg13g2_fill_2 FILLER_52_59 ();
 sg13g2_fill_1 FILLER_52_65 ();
 sg13g2_fill_2 FILLER_52_74 ();
 sg13g2_decap_8 FILLER_52_80 ();
 sg13g2_fill_2 FILLER_52_87 ();
 sg13g2_decap_4 FILLER_52_93 ();
 sg13g2_fill_1 FILLER_52_97 ();
 sg13g2_fill_1 FILLER_52_102 ();
 sg13g2_decap_4 FILLER_52_107 ();
 sg13g2_fill_2 FILLER_52_137 ();
 sg13g2_fill_1 FILLER_52_139 ();
 sg13g2_fill_2 FILLER_52_148 ();
 sg13g2_fill_1 FILLER_52_150 ();
 sg13g2_decap_4 FILLER_52_167 ();
 sg13g2_fill_2 FILLER_52_183 ();
 sg13g2_decap_4 FILLER_52_190 ();
 sg13g2_decap_4 FILLER_52_200 ();
 sg13g2_fill_2 FILLER_52_210 ();
 sg13g2_fill_1 FILLER_52_212 ();
 sg13g2_fill_2 FILLER_52_218 ();
 sg13g2_fill_1 FILLER_52_220 ();
 sg13g2_fill_2 FILLER_52_224 ();
 sg13g2_decap_4 FILLER_52_238 ();
 sg13g2_fill_1 FILLER_52_247 ();
 sg13g2_fill_2 FILLER_52_254 ();
 sg13g2_fill_2 FILLER_52_269 ();
 sg13g2_fill_1 FILLER_52_271 ();
 sg13g2_fill_1 FILLER_52_303 ();
 sg13g2_decap_8 FILLER_52_312 ();
 sg13g2_decap_4 FILLER_52_319 ();
 sg13g2_fill_1 FILLER_52_323 ();
 sg13g2_fill_1 FILLER_52_372 ();
 sg13g2_fill_2 FILLER_52_377 ();
 sg13g2_fill_1 FILLER_52_422 ();
 sg13g2_fill_2 FILLER_52_427 ();
 sg13g2_fill_1 FILLER_52_429 ();
 sg13g2_fill_1 FILLER_53_13 ();
 sg13g2_fill_2 FILLER_53_19 ();
 sg13g2_fill_2 FILLER_53_29 ();
 sg13g2_fill_2 FILLER_53_42 ();
 sg13g2_fill_1 FILLER_53_49 ();
 sg13g2_fill_1 FILLER_53_55 ();
 sg13g2_fill_1 FILLER_53_66 ();
 sg13g2_decap_4 FILLER_53_94 ();
 sg13g2_fill_1 FILLER_53_98 ();
 sg13g2_fill_2 FILLER_53_104 ();
 sg13g2_fill_1 FILLER_53_106 ();
 sg13g2_fill_2 FILLER_53_111 ();
 sg13g2_fill_1 FILLER_53_113 ();
 sg13g2_decap_8 FILLER_53_122 ();
 sg13g2_fill_1 FILLER_53_129 ();
 sg13g2_decap_8 FILLER_53_134 ();
 sg13g2_fill_2 FILLER_53_141 ();
 sg13g2_fill_1 FILLER_53_143 ();
 sg13g2_decap_8 FILLER_53_147 ();
 sg13g2_decap_4 FILLER_53_154 ();
 sg13g2_fill_1 FILLER_53_170 ();
 sg13g2_fill_1 FILLER_53_174 ();
 sg13g2_fill_1 FILLER_53_180 ();
 sg13g2_fill_1 FILLER_53_185 ();
 sg13g2_fill_1 FILLER_53_216 ();
 sg13g2_fill_2 FILLER_53_227 ();
 sg13g2_fill_1 FILLER_53_248 ();
 sg13g2_decap_4 FILLER_53_253 ();
 sg13g2_fill_1 FILLER_53_282 ();
 sg13g2_fill_1 FILLER_53_288 ();
 sg13g2_fill_2 FILLER_53_299 ();
 sg13g2_fill_1 FILLER_53_305 ();
 sg13g2_decap_4 FILLER_53_336 ();
 sg13g2_fill_1 FILLER_53_340 ();
 sg13g2_decap_4 FILLER_53_345 ();
 sg13g2_fill_1 FILLER_53_349 ();
 sg13g2_decap_8 FILLER_53_354 ();
 sg13g2_decap_4 FILLER_53_365 ();
 sg13g2_fill_1 FILLER_53_380 ();
 sg13g2_fill_1 FILLER_53_385 ();
 sg13g2_fill_1 FILLER_53_390 ();
 sg13g2_fill_1 FILLER_53_395 ();
 sg13g2_decap_8 FILLER_54_0 ();
 sg13g2_fill_1 FILLER_54_7 ();
 sg13g2_fill_2 FILLER_54_13 ();
 sg13g2_fill_1 FILLER_54_15 ();
 sg13g2_fill_1 FILLER_54_19 ();
 sg13g2_fill_1 FILLER_54_30 ();
 sg13g2_fill_1 FILLER_54_52 ();
 sg13g2_fill_2 FILLER_54_67 ();
 sg13g2_fill_1 FILLER_54_69 ();
 sg13g2_fill_1 FILLER_54_79 ();
 sg13g2_fill_1 FILLER_54_93 ();
 sg13g2_decap_4 FILLER_54_108 ();
 sg13g2_fill_1 FILLER_54_115 ();
 sg13g2_fill_2 FILLER_54_120 ();
 sg13g2_fill_1 FILLER_54_125 ();
 sg13g2_fill_1 FILLER_54_131 ();
 sg13g2_fill_2 FILLER_54_137 ();
 sg13g2_fill_1 FILLER_54_139 ();
 sg13g2_fill_1 FILLER_54_154 ();
 sg13g2_fill_1 FILLER_54_162 ();
 sg13g2_fill_1 FILLER_54_168 ();
 sg13g2_fill_2 FILLER_54_174 ();
 sg13g2_fill_1 FILLER_54_180 ();
 sg13g2_fill_2 FILLER_54_184 ();
 sg13g2_fill_1 FILLER_54_191 ();
 sg13g2_fill_2 FILLER_54_197 ();
 sg13g2_fill_2 FILLER_54_205 ();
 sg13g2_fill_1 FILLER_54_230 ();
 sg13g2_decap_4 FILLER_54_234 ();
 sg13g2_fill_1 FILLER_54_238 ();
 sg13g2_decap_8 FILLER_54_242 ();
 sg13g2_fill_1 FILLER_54_249 ();
 sg13g2_decap_8 FILLER_54_255 ();
 sg13g2_fill_2 FILLER_54_262 ();
 sg13g2_fill_1 FILLER_54_289 ();
 sg13g2_decap_8 FILLER_54_325 ();
 sg13g2_fill_1 FILLER_54_332 ();
 sg13g2_fill_2 FILLER_54_408 ();
 sg13g2_fill_1 FILLER_54_410 ();
 sg13g2_decap_8 FILLER_54_415 ();
 sg13g2_decap_8 FILLER_54_422 ();
 sg13g2_fill_1 FILLER_54_429 ();
 sg13g2_decap_8 FILLER_55_0 ();
 sg13g2_fill_2 FILLER_55_7 ();
 sg13g2_fill_2 FILLER_55_22 ();
 sg13g2_fill_1 FILLER_55_24 ();
 sg13g2_fill_2 FILLER_55_29 ();
 sg13g2_fill_1 FILLER_55_31 ();
 sg13g2_decap_8 FILLER_55_35 ();
 sg13g2_decap_4 FILLER_55_42 ();
 sg13g2_fill_2 FILLER_55_46 ();
 sg13g2_fill_1 FILLER_55_52 ();
 sg13g2_fill_2 FILLER_55_60 ();
 sg13g2_fill_1 FILLER_55_62 ();
 sg13g2_fill_2 FILLER_55_68 ();
 sg13g2_fill_1 FILLER_55_70 ();
 sg13g2_fill_1 FILLER_55_79 ();
 sg13g2_decap_4 FILLER_55_85 ();
 sg13g2_fill_1 FILLER_55_89 ();
 sg13g2_decap_4 FILLER_55_98 ();
 sg13g2_fill_2 FILLER_55_106 ();
 sg13g2_fill_1 FILLER_55_108 ();
 sg13g2_decap_4 FILLER_55_144 ();
 sg13g2_decap_4 FILLER_55_156 ();
 sg13g2_fill_2 FILLER_55_215 ();
 sg13g2_decap_4 FILLER_55_222 ();
 sg13g2_decap_8 FILLER_55_261 ();
 sg13g2_decap_4 FILLER_55_268 ();
 sg13g2_fill_1 FILLER_55_277 ();
 sg13g2_fill_1 FILLER_55_288 ();
 sg13g2_fill_2 FILLER_55_293 ();
 sg13g2_fill_1 FILLER_55_295 ();
 sg13g2_fill_2 FILLER_55_322 ();
 sg13g2_fill_1 FILLER_55_328 ();
 sg13g2_fill_2 FILLER_55_338 ();
 sg13g2_fill_1 FILLER_55_340 ();
 sg13g2_fill_1 FILLER_55_349 ();
 sg13g2_fill_1 FILLER_55_358 ();
 sg13g2_fill_2 FILLER_55_380 ();
 sg13g2_decap_4 FILLER_55_400 ();
 sg13g2_decap_8 FILLER_56_0 ();
 sg13g2_fill_1 FILLER_56_7 ();
 sg13g2_fill_1 FILLER_56_31 ();
 sg13g2_fill_2 FILLER_56_36 ();
 sg13g2_fill_1 FILLER_56_47 ();
 sg13g2_fill_2 FILLER_56_74 ();
 sg13g2_fill_1 FILLER_56_76 ();
 sg13g2_fill_1 FILLER_56_82 ();
 sg13g2_decap_4 FILLER_56_88 ();
 sg13g2_fill_2 FILLER_56_102 ();
 sg13g2_decap_8 FILLER_56_109 ();
 sg13g2_decap_4 FILLER_56_126 ();
 sg13g2_fill_1 FILLER_56_139 ();
 sg13g2_fill_1 FILLER_56_145 ();
 sg13g2_fill_1 FILLER_56_151 ();
 sg13g2_fill_2 FILLER_56_157 ();
 sg13g2_fill_2 FILLER_56_168 ();
 sg13g2_fill_1 FILLER_56_170 ();
 sg13g2_fill_2 FILLER_56_185 ();
 sg13g2_decap_4 FILLER_56_191 ();
 sg13g2_decap_4 FILLER_56_199 ();
 sg13g2_decap_4 FILLER_56_209 ();
 sg13g2_fill_2 FILLER_56_225 ();
 sg13g2_fill_2 FILLER_56_231 ();
 sg13g2_fill_1 FILLER_56_233 ();
 sg13g2_fill_2 FILLER_56_248 ();
 sg13g2_fill_1 FILLER_56_250 ();
 sg13g2_decap_8 FILLER_56_255 ();
 sg13g2_decap_4 FILLER_56_297 ();
 sg13g2_fill_2 FILLER_56_301 ();
 sg13g2_fill_2 FILLER_56_307 ();
 sg13g2_fill_1 FILLER_56_335 ();
 sg13g2_fill_2 FILLER_56_340 ();
 sg13g2_fill_1 FILLER_56_342 ();
 sg13g2_fill_2 FILLER_56_351 ();
 sg13g2_fill_2 FILLER_56_392 ();
 sg13g2_decap_8 FILLER_57_0 ();
 sg13g2_decap_8 FILLER_57_7 ();
 sg13g2_fill_1 FILLER_57_14 ();
 sg13g2_fill_2 FILLER_57_24 ();
 sg13g2_decap_4 FILLER_57_31 ();
 sg13g2_fill_2 FILLER_57_40 ();
 sg13g2_fill_2 FILLER_57_57 ();
 sg13g2_fill_1 FILLER_57_59 ();
 sg13g2_fill_1 FILLER_57_83 ();
 sg13g2_fill_1 FILLER_57_97 ();
 sg13g2_fill_1 FILLER_57_107 ();
 sg13g2_fill_2 FILLER_57_141 ();
 sg13g2_decap_8 FILLER_57_190 ();
 sg13g2_fill_1 FILLER_57_197 ();
 sg13g2_decap_8 FILLER_57_210 ();
 sg13g2_decap_4 FILLER_57_217 ();
 sg13g2_decap_4 FILLER_57_231 ();
 sg13g2_fill_1 FILLER_57_243 ();
 sg13g2_fill_2 FILLER_57_270 ();
 sg13g2_fill_1 FILLER_57_272 ();
 sg13g2_fill_1 FILLER_57_276 ();
 sg13g2_fill_2 FILLER_57_287 ();
 sg13g2_fill_1 FILLER_57_289 ();
 sg13g2_decap_4 FILLER_57_294 ();
 sg13g2_fill_1 FILLER_57_298 ();
 sg13g2_fill_2 FILLER_57_304 ();
 sg13g2_fill_1 FILLER_57_306 ();
 sg13g2_decap_8 FILLER_57_363 ();
 sg13g2_fill_1 FILLER_57_373 ();
 sg13g2_fill_1 FILLER_57_382 ();
 sg13g2_decap_8 FILLER_57_394 ();
 sg13g2_decap_4 FILLER_57_401 ();
 sg13g2_fill_1 FILLER_57_405 ();
 sg13g2_fill_2 FILLER_57_410 ();
 sg13g2_fill_1 FILLER_57_412 ();
 sg13g2_fill_2 FILLER_57_417 ();
 sg13g2_fill_2 FILLER_57_427 ();
 sg13g2_fill_1 FILLER_57_429 ();
 sg13g2_fill_2 FILLER_58_0 ();
 sg13g2_fill_1 FILLER_58_6 ();
 sg13g2_fill_1 FILLER_58_25 ();
 sg13g2_fill_1 FILLER_58_40 ();
 sg13g2_fill_1 FILLER_58_45 ();
 sg13g2_fill_1 FILLER_58_50 ();
 sg13g2_fill_1 FILLER_58_55 ();
 sg13g2_fill_1 FILLER_58_62 ();
 sg13g2_fill_2 FILLER_58_67 ();
 sg13g2_fill_2 FILLER_58_73 ();
 sg13g2_fill_2 FILLER_58_79 ();
 sg13g2_fill_1 FILLER_58_81 ();
 sg13g2_fill_1 FILLER_58_87 ();
 sg13g2_fill_2 FILLER_58_92 ();
 sg13g2_fill_1 FILLER_58_94 ();
 sg13g2_decap_8 FILLER_58_105 ();
 sg13g2_decap_8 FILLER_58_112 ();
 sg13g2_fill_1 FILLER_58_119 ();
 sg13g2_fill_1 FILLER_58_131 ();
 sg13g2_fill_1 FILLER_58_135 ();
 sg13g2_fill_1 FILLER_58_144 ();
 sg13g2_decap_4 FILLER_58_151 ();
 sg13g2_decap_8 FILLER_58_160 ();
 sg13g2_decap_8 FILLER_58_167 ();
 sg13g2_fill_2 FILLER_58_177 ();
 sg13g2_decap_8 FILLER_58_220 ();
 sg13g2_decap_8 FILLER_58_227 ();
 sg13g2_decap_4 FILLER_58_234 ();
 sg13g2_fill_1 FILLER_58_242 ();
 sg13g2_fill_1 FILLER_58_273 ();
 sg13g2_decap_4 FILLER_58_326 ();
 sg13g2_fill_2 FILLER_58_330 ();
 sg13g2_fill_2 FILLER_58_335 ();
 sg13g2_fill_2 FILLER_58_374 ();
 sg13g2_decap_4 FILLER_58_381 ();
 sg13g2_fill_2 FILLER_58_385 ();
 sg13g2_fill_1 FILLER_58_394 ();
 sg13g2_fill_1 FILLER_58_408 ();
 sg13g2_fill_1 FILLER_58_419 ();
 sg13g2_decap_4 FILLER_58_425 ();
 sg13g2_fill_1 FILLER_58_429 ();
 sg13g2_fill_2 FILLER_59_22 ();
 sg13g2_fill_2 FILLER_59_43 ();
 sg13g2_decap_4 FILLER_59_54 ();
 sg13g2_fill_2 FILLER_59_58 ();
 sg13g2_fill_1 FILLER_59_76 ();
 sg13g2_decap_4 FILLER_59_86 ();
 sg13g2_fill_1 FILLER_59_102 ();
 sg13g2_decap_8 FILLER_59_107 ();
 sg13g2_decap_8 FILLER_59_114 ();
 sg13g2_fill_2 FILLER_59_125 ();
 sg13g2_fill_1 FILLER_59_127 ();
 sg13g2_fill_1 FILLER_59_131 ();
 sg13g2_fill_2 FILLER_59_141 ();
 sg13g2_fill_1 FILLER_59_151 ();
 sg13g2_decap_4 FILLER_59_157 ();
 sg13g2_decap_4 FILLER_59_182 ();
 sg13g2_decap_8 FILLER_59_191 ();
 sg13g2_decap_8 FILLER_59_202 ();
 sg13g2_decap_4 FILLER_59_209 ();
 sg13g2_fill_2 FILLER_59_213 ();
 sg13g2_fill_1 FILLER_59_219 ();
 sg13g2_fill_1 FILLER_59_240 ();
 sg13g2_fill_2 FILLER_59_246 ();
 sg13g2_decap_4 FILLER_59_254 ();
 sg13g2_fill_1 FILLER_59_258 ();
 sg13g2_fill_2 FILLER_59_264 ();
 sg13g2_fill_2 FILLER_59_271 ();
 sg13g2_decap_8 FILLER_59_291 ();
 sg13g2_fill_2 FILLER_59_298 ();
 sg13g2_decap_4 FILLER_59_305 ();
 sg13g2_fill_1 FILLER_59_313 ();
 sg13g2_decap_8 FILLER_59_318 ();
 sg13g2_decap_8 FILLER_59_325 ();
 sg13g2_fill_2 FILLER_59_332 ();
 sg13g2_fill_1 FILLER_59_338 ();
 sg13g2_fill_2 FILLER_59_343 ();
 sg13g2_fill_1 FILLER_59_371 ();
 sg13g2_fill_1 FILLER_59_401 ();
 sg13g2_fill_2 FILLER_59_407 ();
 sg13g2_fill_2 FILLER_59_412 ();
 sg13g2_fill_2 FILLER_59_419 ();
 sg13g2_decap_4 FILLER_59_426 ();
 sg13g2_decap_8 FILLER_60_0 ();
 sg13g2_fill_2 FILLER_60_7 ();
 sg13g2_fill_1 FILLER_60_9 ();
 sg13g2_fill_1 FILLER_60_30 ();
 sg13g2_fill_2 FILLER_60_52 ();
 sg13g2_fill_1 FILLER_60_63 ();
 sg13g2_fill_2 FILLER_60_68 ();
 sg13g2_fill_1 FILLER_60_70 ();
 sg13g2_fill_1 FILLER_60_75 ();
 sg13g2_fill_1 FILLER_60_81 ();
 sg13g2_fill_1 FILLER_60_91 ();
 sg13g2_decap_8 FILLER_60_96 ();
 sg13g2_fill_2 FILLER_60_107 ();
 sg13g2_decap_4 FILLER_60_114 ();
 sg13g2_fill_2 FILLER_60_118 ();
 sg13g2_fill_1 FILLER_60_132 ();
 sg13g2_fill_1 FILLER_60_138 ();
 sg13g2_fill_1 FILLER_60_142 ();
 sg13g2_decap_8 FILLER_60_158 ();
 sg13g2_decap_4 FILLER_60_165 ();
 sg13g2_fill_2 FILLER_60_169 ();
 sg13g2_fill_2 FILLER_60_174 ();
 sg13g2_fill_1 FILLER_60_176 ();
 sg13g2_fill_2 FILLER_60_185 ();
 sg13g2_decap_4 FILLER_60_213 ();
 sg13g2_fill_1 FILLER_60_217 ();
 sg13g2_fill_2 FILLER_60_270 ();
 sg13g2_decap_8 FILLER_60_298 ();
 sg13g2_decap_8 FILLER_60_305 ();
 sg13g2_decap_4 FILLER_60_338 ();
 sg13g2_fill_1 FILLER_60_342 ();
 sg13g2_fill_2 FILLER_60_361 ();
 sg13g2_decap_4 FILLER_60_375 ();
 sg13g2_fill_1 FILLER_60_379 ();
 sg13g2_fill_2 FILLER_60_409 ();
 sg13g2_decap_8 FILLER_60_415 ();
 sg13g2_decap_8 FILLER_60_422 ();
 sg13g2_fill_1 FILLER_60_429 ();
 sg13g2_decap_8 FILLER_61_0 ();
 sg13g2_fill_1 FILLER_61_11 ();
 sg13g2_fill_1 FILLER_61_17 ();
 sg13g2_fill_1 FILLER_61_24 ();
 sg13g2_fill_2 FILLER_61_29 ();
 sg13g2_fill_2 FILLER_61_35 ();
 sg13g2_fill_1 FILLER_61_37 ();
 sg13g2_fill_1 FILLER_61_42 ();
 sg13g2_fill_2 FILLER_61_47 ();
 sg13g2_fill_2 FILLER_61_53 ();
 sg13g2_fill_2 FILLER_61_60 ();
 sg13g2_fill_1 FILLER_61_62 ();
 sg13g2_decap_4 FILLER_61_77 ();
 sg13g2_fill_2 FILLER_61_81 ();
 sg13g2_fill_1 FILLER_61_96 ();
 sg13g2_fill_1 FILLER_61_101 ();
 sg13g2_fill_1 FILLER_61_105 ();
 sg13g2_fill_1 FILLER_61_110 ();
 sg13g2_decap_8 FILLER_61_115 ();
 sg13g2_fill_1 FILLER_61_122 ();
 sg13g2_fill_1 FILLER_61_137 ();
 sg13g2_fill_2 FILLER_61_143 ();
 sg13g2_fill_2 FILLER_61_155 ();
 sg13g2_fill_1 FILLER_61_157 ();
 sg13g2_decap_4 FILLER_61_176 ();
 sg13g2_decap_8 FILLER_61_210 ();
 sg13g2_fill_2 FILLER_61_217 ();
 sg13g2_fill_1 FILLER_61_226 ();
 sg13g2_decap_4 FILLER_61_231 ();
 sg13g2_fill_2 FILLER_61_235 ();
 sg13g2_fill_1 FILLER_61_240 ();
 sg13g2_fill_1 FILLER_61_246 ();
 sg13g2_fill_1 FILLER_61_250 ();
 sg13g2_fill_2 FILLER_61_255 ();
 sg13g2_fill_2 FILLER_61_260 ();
 sg13g2_fill_2 FILLER_61_268 ();
 sg13g2_fill_2 FILLER_61_276 ();
 sg13g2_fill_1 FILLER_61_278 ();
 sg13g2_fill_2 FILLER_61_317 ();
 sg13g2_fill_1 FILLER_61_327 ();
 sg13g2_fill_1 FILLER_61_333 ();
 sg13g2_decap_8 FILLER_61_341 ();
 sg13g2_fill_2 FILLER_61_348 ();
 sg13g2_fill_1 FILLER_61_376 ();
 sg13g2_fill_1 FILLER_61_384 ();
 sg13g2_fill_1 FILLER_61_388 ();
 sg13g2_fill_1 FILLER_61_393 ();
 sg13g2_fill_1 FILLER_61_398 ();
 sg13g2_fill_2 FILLER_61_402 ();
 sg13g2_fill_2 FILLER_62_0 ();
 sg13g2_fill_1 FILLER_62_2 ();
 sg13g2_fill_2 FILLER_62_11 ();
 sg13g2_fill_2 FILLER_62_27 ();
 sg13g2_decap_4 FILLER_62_37 ();
 sg13g2_fill_2 FILLER_62_55 ();
 sg13g2_fill_2 FILLER_62_61 ();
 sg13g2_fill_1 FILLER_62_63 ();
 sg13g2_fill_1 FILLER_62_68 ();
 sg13g2_fill_1 FILLER_62_74 ();
 sg13g2_fill_1 FILLER_62_80 ();
 sg13g2_fill_1 FILLER_62_86 ();
 sg13g2_fill_1 FILLER_62_91 ();
 sg13g2_fill_2 FILLER_62_111 ();
 sg13g2_fill_2 FILLER_62_122 ();
 sg13g2_fill_1 FILLER_62_128 ();
 sg13g2_decap_4 FILLER_62_134 ();
 sg13g2_fill_1 FILLER_62_142 ();
 sg13g2_fill_2 FILLER_62_150 ();
 sg13g2_fill_1 FILLER_62_152 ();
 sg13g2_fill_1 FILLER_62_176 ();
 sg13g2_fill_2 FILLER_62_182 ();
 sg13g2_decap_4 FILLER_62_197 ();
 sg13g2_decap_4 FILLER_62_206 ();
 sg13g2_fill_2 FILLER_62_210 ();
 sg13g2_decap_8 FILLER_62_217 ();
 sg13g2_fill_2 FILLER_62_224 ();
 sg13g2_decap_4 FILLER_62_244 ();
 sg13g2_fill_1 FILLER_62_248 ();
 sg13g2_decap_4 FILLER_62_279 ();
 sg13g2_fill_1 FILLER_62_283 ();
 sg13g2_fill_1 FILLER_62_288 ();
 sg13g2_decap_8 FILLER_62_293 ();
 sg13g2_decap_4 FILLER_62_300 ();
 sg13g2_decap_4 FILLER_62_321 ();
 sg13g2_fill_1 FILLER_62_325 ();
 sg13g2_decap_4 FILLER_62_343 ();
 sg13g2_decap_4 FILLER_62_352 ();
 sg13g2_decap_8 FILLER_62_360 ();
 sg13g2_decap_8 FILLER_62_367 ();
 sg13g2_decap_8 FILLER_62_374 ();
 sg13g2_fill_2 FILLER_62_381 ();
 sg13g2_fill_1 FILLER_62_388 ();
 sg13g2_fill_1 FILLER_62_393 ();
 sg13g2_fill_1 FILLER_62_399 ();
 sg13g2_fill_1 FILLER_62_407 ();
 sg13g2_fill_2 FILLER_62_428 ();
 sg13g2_decap_4 FILLER_63_0 ();
 sg13g2_fill_1 FILLER_63_16 ();
 sg13g2_fill_1 FILLER_63_21 ();
 sg13g2_decap_4 FILLER_63_37 ();
 sg13g2_decap_8 FILLER_63_45 ();
 sg13g2_decap_4 FILLER_63_52 ();
 sg13g2_fill_1 FILLER_63_56 ();
 sg13g2_fill_2 FILLER_63_61 ();
 sg13g2_fill_1 FILLER_63_63 ();
 sg13g2_fill_2 FILLER_63_72 ();
 sg13g2_fill_1 FILLER_63_74 ();
 sg13g2_decap_8 FILLER_63_79 ();
 sg13g2_fill_2 FILLER_63_86 ();
 sg13g2_decap_8 FILLER_63_100 ();
 sg13g2_fill_2 FILLER_63_107 ();
 sg13g2_fill_1 FILLER_63_109 ();
 sg13g2_decap_8 FILLER_63_128 ();
 sg13g2_fill_1 FILLER_63_135 ();
 sg13g2_decap_8 FILLER_63_139 ();
 sg13g2_fill_2 FILLER_63_146 ();
 sg13g2_fill_1 FILLER_63_153 ();
 sg13g2_decap_8 FILLER_63_158 ();
 sg13g2_decap_8 FILLER_63_165 ();
 sg13g2_decap_8 FILLER_63_172 ();
 sg13g2_fill_2 FILLER_63_179 ();
 sg13g2_fill_1 FILLER_63_181 ();
 sg13g2_fill_2 FILLER_63_190 ();
 sg13g2_fill_1 FILLER_63_192 ();
 sg13g2_fill_2 FILLER_63_230 ();
 sg13g2_fill_2 FILLER_63_242 ();
 sg13g2_fill_1 FILLER_63_252 ();
 sg13g2_fill_1 FILLER_63_259 ();
 sg13g2_decap_8 FILLER_63_267 ();
 sg13g2_fill_2 FILLER_63_274 ();
 sg13g2_fill_1 FILLER_63_276 ();
 sg13g2_fill_2 FILLER_63_307 ();
 sg13g2_fill_2 FILLER_63_344 ();
 sg13g2_fill_1 FILLER_63_378 ();
 sg13g2_fill_2 FILLER_63_387 ();
 sg13g2_fill_1 FILLER_63_389 ();
 sg13g2_fill_2 FILLER_63_394 ();
 sg13g2_fill_1 FILLER_63_400 ();
 sg13g2_decap_8 FILLER_63_405 ();
 sg13g2_decap_4 FILLER_63_412 ();
 sg13g2_fill_2 FILLER_63_428 ();
 sg13g2_decap_4 FILLER_64_0 ();
 sg13g2_fill_2 FILLER_64_4 ();
 sg13g2_fill_1 FILLER_64_15 ();
 sg13g2_fill_1 FILLER_64_41 ();
 sg13g2_fill_1 FILLER_64_47 ();
 sg13g2_fill_1 FILLER_64_56 ();
 sg13g2_fill_2 FILLER_64_63 ();
 sg13g2_fill_1 FILLER_64_65 ();
 sg13g2_fill_2 FILLER_64_98 ();
 sg13g2_fill_1 FILLER_64_100 ();
 sg13g2_decap_4 FILLER_64_114 ();
 sg13g2_fill_1 FILLER_64_118 ();
 sg13g2_fill_2 FILLER_64_132 ();
 sg13g2_decap_8 FILLER_64_146 ();
 sg13g2_decap_8 FILLER_64_153 ();
 sg13g2_fill_1 FILLER_64_160 ();
 sg13g2_decap_4 FILLER_64_195 ();
 sg13g2_decap_8 FILLER_64_203 ();
 sg13g2_fill_1 FILLER_64_210 ();
 sg13g2_decap_4 FILLER_64_219 ();
 sg13g2_fill_1 FILLER_64_237 ();
 sg13g2_fill_1 FILLER_64_248 ();
 sg13g2_decap_4 FILLER_64_289 ();
 sg13g2_fill_1 FILLER_64_293 ();
 sg13g2_fill_2 FILLER_64_300 ();
 sg13g2_fill_1 FILLER_64_307 ();
 sg13g2_decap_4 FILLER_64_316 ();
 sg13g2_fill_2 FILLER_64_335 ();
 sg13g2_fill_1 FILLER_64_342 ();
 sg13g2_fill_2 FILLER_64_347 ();
 sg13g2_fill_2 FILLER_64_353 ();
 sg13g2_decap_4 FILLER_64_359 ();
 sg13g2_fill_1 FILLER_64_363 ();
 sg13g2_fill_1 FILLER_64_377 ();
 sg13g2_fill_1 FILLER_64_384 ();
 sg13g2_fill_2 FILLER_64_397 ();
 sg13g2_fill_1 FILLER_64_399 ();
 sg13g2_decap_4 FILLER_65_0 ();
 sg13g2_decap_8 FILLER_65_8 ();
 sg13g2_fill_1 FILLER_65_15 ();
 sg13g2_fill_1 FILLER_65_24 ();
 sg13g2_fill_1 FILLER_65_30 ();
 sg13g2_fill_1 FILLER_65_36 ();
 sg13g2_fill_1 FILLER_65_42 ();
 sg13g2_fill_1 FILLER_65_48 ();
 sg13g2_decap_8 FILLER_65_53 ();
 sg13g2_fill_1 FILLER_65_60 ();
 sg13g2_decap_4 FILLER_65_81 ();
 sg13g2_fill_2 FILLER_65_85 ();
 sg13g2_decap_8 FILLER_65_93 ();
 sg13g2_decap_4 FILLER_65_105 ();
 sg13g2_fill_1 FILLER_65_109 ();
 sg13g2_decap_8 FILLER_65_117 ();
 sg13g2_fill_2 FILLER_65_124 ();
 sg13g2_decap_8 FILLER_65_144 ();
 sg13g2_decap_8 FILLER_65_151 ();
 sg13g2_fill_1 FILLER_65_158 ();
 sg13g2_fill_1 FILLER_65_172 ();
 sg13g2_decap_4 FILLER_65_190 ();
 sg13g2_decap_4 FILLER_65_206 ();
 sg13g2_fill_1 FILLER_65_210 ();
 sg13g2_fill_1 FILLER_65_263 ();
 sg13g2_fill_1 FILLER_65_302 ();
 sg13g2_fill_1 FILLER_65_322 ();
 sg13g2_fill_2 FILLER_65_335 ();
 sg13g2_fill_2 FILLER_65_368 ();
 sg13g2_fill_2 FILLER_65_375 ();
 sg13g2_fill_1 FILLER_65_381 ();
 sg13g2_fill_2 FILLER_65_394 ();
 sg13g2_fill_2 FILLER_65_406 ();
 sg13g2_fill_1 FILLER_65_412 ();
 sg13g2_fill_2 FILLER_65_417 ();
 sg13g2_decap_4 FILLER_65_426 ();
 sg13g2_fill_2 FILLER_66_0 ();
 sg13g2_fill_1 FILLER_66_2 ();
 sg13g2_fill_2 FILLER_66_16 ();
 sg13g2_decap_4 FILLER_66_21 ();
 sg13g2_fill_2 FILLER_66_25 ();
 sg13g2_fill_2 FILLER_66_37 ();
 sg13g2_fill_1 FILLER_66_39 ();
 sg13g2_fill_1 FILLER_66_60 ();
 sg13g2_fill_1 FILLER_66_66 ();
 sg13g2_fill_1 FILLER_66_72 ();
 sg13g2_fill_1 FILLER_66_88 ();
 sg13g2_fill_1 FILLER_66_98 ();
 sg13g2_decap_8 FILLER_66_103 ();
 sg13g2_decap_4 FILLER_66_110 ();
 sg13g2_fill_2 FILLER_66_114 ();
 sg13g2_decap_8 FILLER_66_145 ();
 sg13g2_decap_8 FILLER_66_152 ();
 sg13g2_fill_2 FILLER_66_159 ();
 sg13g2_fill_1 FILLER_66_161 ();
 sg13g2_fill_2 FILLER_66_165 ();
 sg13g2_fill_2 FILLER_66_181 ();
 sg13g2_decap_4 FILLER_66_205 ();
 sg13g2_fill_1 FILLER_66_217 ();
 sg13g2_decap_8 FILLER_66_227 ();
 sg13g2_fill_2 FILLER_66_234 ();
 sg13g2_fill_2 FILLER_66_243 ();
 sg13g2_fill_1 FILLER_66_245 ();
 sg13g2_decap_8 FILLER_66_273 ();
 sg13g2_fill_2 FILLER_66_280 ();
 sg13g2_fill_1 FILLER_66_282 ();
 sg13g2_decap_4 FILLER_66_293 ();
 sg13g2_fill_2 FILLER_66_297 ();
 sg13g2_fill_2 FILLER_66_303 ();
 sg13g2_fill_2 FILLER_66_310 ();
 sg13g2_fill_2 FILLER_66_317 ();
 sg13g2_fill_1 FILLER_66_353 ();
 sg13g2_decap_8 FILLER_66_361 ();
 sg13g2_fill_2 FILLER_66_368 ();
 sg13g2_fill_2 FILLER_66_427 ();
 sg13g2_fill_1 FILLER_66_429 ();
 sg13g2_decap_4 FILLER_67_0 ();
 sg13g2_fill_1 FILLER_67_9 ();
 sg13g2_fill_1 FILLER_67_14 ();
 sg13g2_decap_4 FILLER_67_19 ();
 sg13g2_fill_1 FILLER_67_37 ();
 sg13g2_fill_1 FILLER_67_43 ();
 sg13g2_fill_1 FILLER_67_49 ();
 sg13g2_fill_2 FILLER_67_90 ();
 sg13g2_decap_8 FILLER_67_109 ();
 sg13g2_decap_8 FILLER_67_116 ();
 sg13g2_fill_2 FILLER_67_123 ();
 sg13g2_fill_1 FILLER_67_130 ();
 sg13g2_fill_1 FILLER_67_135 ();
 sg13g2_fill_2 FILLER_67_140 ();
 sg13g2_fill_2 FILLER_67_168 ();
 sg13g2_fill_2 FILLER_67_175 ();
 sg13g2_fill_1 FILLER_67_177 ();
 sg13g2_fill_2 FILLER_67_188 ();
 sg13g2_fill_2 FILLER_67_200 ();
 sg13g2_fill_2 FILLER_67_211 ();
 sg13g2_fill_1 FILLER_67_233 ();
 sg13g2_decap_4 FILLER_67_251 ();
 sg13g2_fill_1 FILLER_67_255 ();
 sg13g2_fill_1 FILLER_67_264 ();
 sg13g2_decap_4 FILLER_67_268 ();
 sg13g2_fill_1 FILLER_67_272 ();
 sg13g2_fill_1 FILLER_67_279 ();
 sg13g2_fill_1 FILLER_67_284 ();
 sg13g2_fill_1 FILLER_67_311 ();
 sg13g2_fill_1 FILLER_67_316 ();
 sg13g2_fill_1 FILLER_67_321 ();
 sg13g2_fill_1 FILLER_67_371 ();
 sg13g2_fill_2 FILLER_67_398 ();
 sg13g2_decap_4 FILLER_67_426 ();
 sg13g2_fill_2 FILLER_68_0 ();
 sg13g2_fill_1 FILLER_68_2 ();
 sg13g2_fill_1 FILLER_68_11 ();
 sg13g2_fill_2 FILLER_68_32 ();
 sg13g2_fill_1 FILLER_68_34 ();
 sg13g2_fill_2 FILLER_68_40 ();
 sg13g2_decap_4 FILLER_68_55 ();
 sg13g2_fill_2 FILLER_68_59 ();
 sg13g2_fill_2 FILLER_68_71 ();
 sg13g2_decap_4 FILLER_68_77 ();
 sg13g2_fill_2 FILLER_68_85 ();
 sg13g2_decap_4 FILLER_68_96 ();
 sg13g2_decap_8 FILLER_68_118 ();
 sg13g2_fill_1 FILLER_68_125 ();
 sg13g2_fill_1 FILLER_68_136 ();
 sg13g2_decap_4 FILLER_68_145 ();
 sg13g2_fill_1 FILLER_68_149 ();
 sg13g2_fill_2 FILLER_68_154 ();
 sg13g2_fill_2 FILLER_68_161 ();
 sg13g2_decap_4 FILLER_68_167 ();
 sg13g2_fill_1 FILLER_68_182 ();
 sg13g2_fill_1 FILLER_68_187 ();
 sg13g2_decap_8 FILLER_68_229 ();
 sg13g2_fill_1 FILLER_68_236 ();
 sg13g2_fill_1 FILLER_68_249 ();
 sg13g2_decap_4 FILLER_68_255 ();
 sg13g2_fill_1 FILLER_68_259 ();
 sg13g2_decap_8 FILLER_68_282 ();
 sg13g2_decap_4 FILLER_68_329 ();
 sg13g2_fill_2 FILLER_68_333 ();
 sg13g2_fill_2 FILLER_68_339 ();
 sg13g2_fill_1 FILLER_68_355 ();
 sg13g2_fill_1 FILLER_68_361 ();
 sg13g2_fill_2 FILLER_68_367 ();
 sg13g2_fill_1 FILLER_68_369 ();
 sg13g2_decap_4 FILLER_68_374 ();
 sg13g2_fill_2 FILLER_68_378 ();
 sg13g2_fill_2 FILLER_68_384 ();
 sg13g2_fill_1 FILLER_68_429 ();
 sg13g2_fill_1 FILLER_69_0 ();
 sg13g2_decap_8 FILLER_69_6 ();
 sg13g2_fill_2 FILLER_69_17 ();
 sg13g2_fill_2 FILLER_69_28 ();
 sg13g2_fill_1 FILLER_69_35 ();
 sg13g2_fill_1 FILLER_69_50 ();
 sg13g2_fill_1 FILLER_69_65 ();
 sg13g2_fill_2 FILLER_69_71 ();
 sg13g2_fill_2 FILLER_69_77 ();
 sg13g2_decap_4 FILLER_69_84 ();
 sg13g2_fill_2 FILLER_69_97 ();
 sg13g2_fill_1 FILLER_69_99 ();
 sg13g2_decap_4 FILLER_69_108 ();
 sg13g2_fill_2 FILLER_69_117 ();
 sg13g2_fill_1 FILLER_69_119 ();
 sg13g2_decap_8 FILLER_69_124 ();
 sg13g2_decap_4 FILLER_69_131 ();
 sg13g2_fill_2 FILLER_69_135 ();
 sg13g2_decap_4 FILLER_69_146 ();
 sg13g2_fill_2 FILLER_69_165 ();
 sg13g2_fill_2 FILLER_69_190 ();
 sg13g2_fill_1 FILLER_69_192 ();
 sg13g2_fill_1 FILLER_69_198 ();
 sg13g2_fill_2 FILLER_69_203 ();
 sg13g2_fill_1 FILLER_69_209 ();
 sg13g2_decap_4 FILLER_69_218 ();
 sg13g2_fill_1 FILLER_69_222 ();
 sg13g2_fill_1 FILLER_69_248 ();
 sg13g2_decap_4 FILLER_69_253 ();
 sg13g2_fill_2 FILLER_69_257 ();
 sg13g2_fill_1 FILLER_69_263 ();
 sg13g2_fill_2 FILLER_69_290 ();
 sg13g2_fill_1 FILLER_69_292 ();
 sg13g2_decap_8 FILLER_69_297 ();
 sg13g2_fill_2 FILLER_69_304 ();
 sg13g2_fill_1 FILLER_69_306 ();
 sg13g2_fill_2 FILLER_69_336 ();
 sg13g2_fill_1 FILLER_69_338 ();
 sg13g2_fill_1 FILLER_69_349 ();
 sg13g2_fill_2 FILLER_69_354 ();
 sg13g2_fill_1 FILLER_69_356 ();
 sg13g2_fill_2 FILLER_69_391 ();
 sg13g2_decap_8 FILLER_69_397 ();
 sg13g2_fill_2 FILLER_69_404 ();
 sg13g2_decap_8 FILLER_69_410 ();
 sg13g2_fill_2 FILLER_69_417 ();
 sg13g2_fill_1 FILLER_70_0 ();
 sg13g2_fill_1 FILLER_70_56 ();
 sg13g2_fill_1 FILLER_70_61 ();
 sg13g2_fill_1 FILLER_70_67 ();
 sg13g2_fill_1 FILLER_70_75 ();
 sg13g2_fill_2 FILLER_70_81 ();
 sg13g2_fill_2 FILLER_70_87 ();
 sg13g2_fill_1 FILLER_70_93 ();
 sg13g2_fill_2 FILLER_70_100 ();
 sg13g2_fill_2 FILLER_70_114 ();
 sg13g2_decap_4 FILLER_70_167 ();
 sg13g2_fill_2 FILLER_70_171 ();
 sg13g2_fill_2 FILLER_70_178 ();
 sg13g2_fill_1 FILLER_70_180 ();
 sg13g2_fill_1 FILLER_70_186 ();
 sg13g2_fill_1 FILLER_70_192 ();
 sg13g2_fill_2 FILLER_70_228 ();
 sg13g2_decap_8 FILLER_70_234 ();
 sg13g2_decap_4 FILLER_70_241 ();
 sg13g2_fill_2 FILLER_70_245 ();
 sg13g2_decap_4 FILLER_70_256 ();
 sg13g2_fill_2 FILLER_70_260 ();
 sg13g2_decap_4 FILLER_70_292 ();
 sg13g2_decap_8 FILLER_70_300 ();
 sg13g2_fill_1 FILLER_70_307 ();
 sg13g2_fill_2 FILLER_70_317 ();
 sg13g2_fill_1 FILLER_70_328 ();
 sg13g2_fill_1 FILLER_70_355 ();
 sg13g2_fill_1 FILLER_70_373 ();
 sg13g2_decap_8 FILLER_70_378 ();
 sg13g2_fill_1 FILLER_70_385 ();
 sg13g2_fill_1 FILLER_70_417 ();
 sg13g2_fill_2 FILLER_70_427 ();
 sg13g2_fill_1 FILLER_70_429 ();
 sg13g2_fill_2 FILLER_71_25 ();
 sg13g2_fill_2 FILLER_71_55 ();
 sg13g2_fill_2 FILLER_71_69 ();
 sg13g2_fill_1 FILLER_71_80 ();
 sg13g2_fill_1 FILLER_71_90 ();
 sg13g2_decap_4 FILLER_71_106 ();
 sg13g2_fill_2 FILLER_71_110 ();
 sg13g2_decap_4 FILLER_71_116 ();
 sg13g2_decap_4 FILLER_71_125 ();
 sg13g2_fill_2 FILLER_71_129 ();
 sg13g2_decap_8 FILLER_71_139 ();
 sg13g2_decap_8 FILLER_71_146 ();
 sg13g2_decap_4 FILLER_71_157 ();
 sg13g2_fill_2 FILLER_71_166 ();
 sg13g2_fill_1 FILLER_71_171 ();
 sg13g2_fill_1 FILLER_71_188 ();
 sg13g2_fill_2 FILLER_71_202 ();
 sg13g2_fill_1 FILLER_71_225 ();
 sg13g2_decap_4 FILLER_71_230 ();
 sg13g2_fill_1 FILLER_71_234 ();
 sg13g2_fill_2 FILLER_71_270 ();
 sg13g2_fill_1 FILLER_71_272 ();
 sg13g2_fill_1 FILLER_71_278 ();
 sg13g2_fill_1 FILLER_71_284 ();
 sg13g2_decap_4 FILLER_71_326 ();
 sg13g2_fill_2 FILLER_71_330 ();
 sg13g2_fill_1 FILLER_71_336 ();
 sg13g2_fill_2 FILLER_71_347 ();
 sg13g2_fill_2 FILLER_71_354 ();
 sg13g2_fill_2 FILLER_71_396 ();
 sg13g2_fill_2 FILLER_71_402 ();
 sg13g2_decap_8 FILLER_72_0 ();
 sg13g2_decap_8 FILLER_72_7 ();
 sg13g2_fill_2 FILLER_72_14 ();
 sg13g2_fill_1 FILLER_72_16 ();
 sg13g2_fill_2 FILLER_72_29 ();
 sg13g2_fill_2 FILLER_72_36 ();
 sg13g2_fill_2 FILLER_72_43 ();
 sg13g2_fill_1 FILLER_72_45 ();
 sg13g2_decap_4 FILLER_72_54 ();
 sg13g2_fill_2 FILLER_72_70 ();
 sg13g2_fill_2 FILLER_72_76 ();
 sg13g2_fill_1 FILLER_72_78 ();
 sg13g2_fill_1 FILLER_72_84 ();
 sg13g2_fill_2 FILLER_72_95 ();
 sg13g2_decap_4 FILLER_72_101 ();
 sg13g2_fill_1 FILLER_72_127 ();
 sg13g2_fill_1 FILLER_72_137 ();
 sg13g2_fill_2 FILLER_72_143 ();
 sg13g2_fill_1 FILLER_72_145 ();
 sg13g2_fill_1 FILLER_72_189 ();
 sg13g2_fill_2 FILLER_72_193 ();
 sg13g2_decap_8 FILLER_72_199 ();
 sg13g2_decap_4 FILLER_72_206 ();
 sg13g2_fill_1 FILLER_72_241 ();
 sg13g2_fill_1 FILLER_72_268 ();
 sg13g2_fill_1 FILLER_72_279 ();
 sg13g2_fill_1 FILLER_72_283 ();
 sg13g2_fill_2 FILLER_72_310 ();
 sg13g2_decap_4 FILLER_72_331 ();
 sg13g2_fill_1 FILLER_72_335 ();
 sg13g2_fill_1 FILLER_72_349 ();
 sg13g2_fill_1 FILLER_72_395 ();
 sg13g2_fill_2 FILLER_72_399 ();
 sg13g2_decap_4 FILLER_72_405 ();
 sg13g2_fill_2 FILLER_72_412 ();
 sg13g2_fill_1 FILLER_72_418 ();
 sg13g2_fill_2 FILLER_73_0 ();
 sg13g2_fill_2 FILLER_73_15 ();
 sg13g2_fill_1 FILLER_73_17 ();
 sg13g2_fill_1 FILLER_73_27 ();
 sg13g2_fill_1 FILLER_73_33 ();
 sg13g2_fill_1 FILLER_73_39 ();
 sg13g2_decap_4 FILLER_73_50 ();
 sg13g2_fill_1 FILLER_73_54 ();
 sg13g2_decap_4 FILLER_73_60 ();
 sg13g2_fill_1 FILLER_73_64 ();
 sg13g2_fill_1 FILLER_73_85 ();
 sg13g2_decap_8 FILLER_73_94 ();
 sg13g2_fill_1 FILLER_73_101 ();
 sg13g2_fill_1 FILLER_73_107 ();
 sg13g2_fill_2 FILLER_73_112 ();
 sg13g2_fill_1 FILLER_73_122 ();
 sg13g2_fill_1 FILLER_73_127 ();
 sg13g2_decap_4 FILLER_73_132 ();
 sg13g2_decap_8 FILLER_73_140 ();
 sg13g2_decap_4 FILLER_73_147 ();
 sg13g2_fill_2 FILLER_73_156 ();
 sg13g2_fill_1 FILLER_73_158 ();
 sg13g2_fill_2 FILLER_73_164 ();
 sg13g2_fill_1 FILLER_73_166 ();
 sg13g2_decap_8 FILLER_73_189 ();
 sg13g2_decap_4 FILLER_73_196 ();
 sg13g2_fill_1 FILLER_73_214 ();
 sg13g2_fill_2 FILLER_73_220 ();
 sg13g2_decap_8 FILLER_73_227 ();
 sg13g2_decap_4 FILLER_73_234 ();
 sg13g2_fill_1 FILLER_73_238 ();
 sg13g2_fill_1 FILLER_73_243 ();
 sg13g2_fill_1 FILLER_73_248 ();
 sg13g2_decap_8 FILLER_73_257 ();
 sg13g2_fill_2 FILLER_73_264 ();
 sg13g2_fill_1 FILLER_73_266 ();
 sg13g2_fill_1 FILLER_73_272 ();
 sg13g2_fill_1 FILLER_73_277 ();
 sg13g2_fill_1 FILLER_73_283 ();
 sg13g2_fill_2 FILLER_73_288 ();
 sg13g2_fill_2 FILLER_73_294 ();
 sg13g2_fill_1 FILLER_73_296 ();
 sg13g2_fill_2 FILLER_73_302 ();
 sg13g2_fill_1 FILLER_73_304 ();
 sg13g2_fill_2 FILLER_73_310 ();
 sg13g2_fill_1 FILLER_73_312 ();
 sg13g2_fill_1 FILLER_73_317 ();
 sg13g2_fill_1 FILLER_73_344 ();
 sg13g2_fill_1 FILLER_73_348 ();
 sg13g2_fill_1 FILLER_73_356 ();
 sg13g2_fill_2 FILLER_73_362 ();
 sg13g2_decap_4 FILLER_73_368 ();
 sg13g2_decap_4 FILLER_73_376 ();
 sg13g2_fill_2 FILLER_73_384 ();
 sg13g2_decap_8 FILLER_74_0 ();
 sg13g2_fill_2 FILLER_74_7 ();
 sg13g2_fill_1 FILLER_74_9 ();
 sg13g2_fill_1 FILLER_74_19 ();
 sg13g2_fill_2 FILLER_74_29 ();
 sg13g2_fill_1 FILLER_74_31 ();
 sg13g2_fill_2 FILLER_74_35 ();
 sg13g2_fill_1 FILLER_74_37 ();
 sg13g2_fill_2 FILLER_74_43 ();
 sg13g2_fill_1 FILLER_74_64 ();
 sg13g2_fill_1 FILLER_74_70 ();
 sg13g2_fill_1 FILLER_74_75 ();
 sg13g2_fill_2 FILLER_74_90 ();
 sg13g2_decap_4 FILLER_74_101 ();
 sg13g2_fill_1 FILLER_74_114 ();
 sg13g2_fill_2 FILLER_74_121 ();
 sg13g2_fill_1 FILLER_74_123 ();
 sg13g2_decap_4 FILLER_74_128 ();
 sg13g2_fill_1 FILLER_74_132 ();
 sg13g2_fill_1 FILLER_74_167 ();
 sg13g2_decap_4 FILLER_74_185 ();
 sg13g2_fill_1 FILLER_74_189 ();
 sg13g2_fill_2 FILLER_74_194 ();
 sg13g2_decap_4 FILLER_74_205 ();
 sg13g2_fill_2 FILLER_74_214 ();
 sg13g2_fill_1 FILLER_74_242 ();
 sg13g2_fill_2 FILLER_74_269 ();
 sg13g2_fill_2 FILLER_74_274 ();
 sg13g2_fill_2 FILLER_74_281 ();
 sg13g2_decap_4 FILLER_74_291 ();
 sg13g2_fill_1 FILLER_74_295 ();
 sg13g2_fill_1 FILLER_74_306 ();
 sg13g2_fill_1 FILLER_74_312 ();
 sg13g2_fill_2 FILLER_74_322 ();
 sg13g2_decap_8 FILLER_74_333 ();
 sg13g2_fill_2 FILLER_74_340 ();
 sg13g2_fill_2 FILLER_74_412 ();
 sg13g2_fill_1 FILLER_74_414 ();
 sg13g2_fill_2 FILLER_74_428 ();
 sg13g2_decap_8 FILLER_75_0 ();
 sg13g2_decap_8 FILLER_75_7 ();
 sg13g2_fill_2 FILLER_75_23 ();
 sg13g2_fill_1 FILLER_75_25 ();
 sg13g2_fill_1 FILLER_75_34 ();
 sg13g2_fill_2 FILLER_75_57 ();
 sg13g2_fill_2 FILLER_75_67 ();
 sg13g2_fill_2 FILLER_75_73 ();
 sg13g2_fill_2 FILLER_75_82 ();
 sg13g2_fill_1 FILLER_75_88 ();
 sg13g2_fill_2 FILLER_75_94 ();
 sg13g2_fill_1 FILLER_75_109 ();
 sg13g2_decap_8 FILLER_75_131 ();
 sg13g2_decap_4 FILLER_75_138 ();
 sg13g2_fill_2 FILLER_75_142 ();
 sg13g2_decap_8 FILLER_75_153 ();
 sg13g2_fill_1 FILLER_75_160 ();
 sg13g2_decap_4 FILLER_75_164 ();
 sg13g2_fill_1 FILLER_75_171 ();
 sg13g2_fill_2 FILLER_75_224 ();
 sg13g2_decap_4 FILLER_75_230 ();
 sg13g2_fill_1 FILLER_75_234 ();
 sg13g2_decap_8 FILLER_75_239 ();
 sg13g2_decap_8 FILLER_75_246 ();
 sg13g2_decap_8 FILLER_75_258 ();
 sg13g2_fill_1 FILLER_75_265 ();
 sg13g2_fill_1 FILLER_75_312 ();
 sg13g2_fill_1 FILLER_75_325 ();
 sg13g2_fill_1 FILLER_75_331 ();
 sg13g2_fill_2 FILLER_75_338 ();
 sg13g2_fill_2 FILLER_75_344 ();
 sg13g2_fill_1 FILLER_75_346 ();
 sg13g2_decap_4 FILLER_75_373 ();
 sg13g2_fill_2 FILLER_75_377 ();
 sg13g2_decap_8 FILLER_75_389 ();
 sg13g2_fill_2 FILLER_75_396 ();
 sg13g2_fill_1 FILLER_75_398 ();
 sg13g2_decap_4 FILLER_76_0 ();
 sg13g2_fill_2 FILLER_76_4 ();
 sg13g2_fill_1 FILLER_76_19 ();
 sg13g2_fill_1 FILLER_76_24 ();
 sg13g2_fill_2 FILLER_76_80 ();
 sg13g2_fill_2 FILLER_76_86 ();
 sg13g2_fill_1 FILLER_76_93 ();
 sg13g2_fill_1 FILLER_76_107 ();
 sg13g2_fill_1 FILLER_76_111 ();
 sg13g2_decap_8 FILLER_76_116 ();
 sg13g2_decap_8 FILLER_76_128 ();
 sg13g2_fill_2 FILLER_76_161 ();
 sg13g2_fill_1 FILLER_76_172 ();
 sg13g2_fill_1 FILLER_76_177 ();
 sg13g2_fill_1 FILLER_76_187 ();
 sg13g2_fill_2 FILLER_76_192 ();
 sg13g2_fill_1 FILLER_76_199 ();
 sg13g2_fill_1 FILLER_76_209 ();
 sg13g2_decap_8 FILLER_76_220 ();
 sg13g2_fill_1 FILLER_76_227 ();
 sg13g2_fill_2 FILLER_76_293 ();
 sg13g2_fill_1 FILLER_76_295 ();
 sg13g2_fill_2 FILLER_76_306 ();
 sg13g2_fill_2 FILLER_76_357 ();
 sg13g2_decap_4 FILLER_76_385 ();
 sg13g2_decap_8 FILLER_77_0 ();
 sg13g2_decap_8 FILLER_77_7 ();
 sg13g2_decap_8 FILLER_77_14 ();
 sg13g2_fill_2 FILLER_77_21 ();
 sg13g2_fill_2 FILLER_77_44 ();
 sg13g2_fill_1 FILLER_77_50 ();
 sg13g2_fill_1 FILLER_77_55 ();
 sg13g2_fill_1 FILLER_77_60 ();
 sg13g2_fill_1 FILLER_77_83 ();
 sg13g2_fill_1 FILLER_77_88 ();
 sg13g2_fill_1 FILLER_77_105 ();
 sg13g2_fill_2 FILLER_77_111 ();
 sg13g2_decap_8 FILLER_77_117 ();
 sg13g2_decap_8 FILLER_77_124 ();
 sg13g2_fill_1 FILLER_77_131 ();
 sg13g2_fill_1 FILLER_77_167 ();
 sg13g2_fill_1 FILLER_77_254 ();
 sg13g2_decap_4 FILLER_77_264 ();
 sg13g2_fill_2 FILLER_77_271 ();
 sg13g2_fill_1 FILLER_77_313 ();
 sg13g2_decap_4 FILLER_77_345 ();
 sg13g2_fill_2 FILLER_77_357 ();
 sg13g2_fill_1 FILLER_77_359 ();
 sg13g2_decap_4 FILLER_77_375 ();
 sg13g2_fill_1 FILLER_77_387 ();
 sg13g2_decap_4 FILLER_77_406 ();
 sg13g2_fill_1 FILLER_77_410 ();
 sg13g2_decap_8 FILLER_77_419 ();
 sg13g2_decap_4 FILLER_77_426 ();
 sg13g2_decap_8 FILLER_78_0 ();
 sg13g2_decap_8 FILLER_78_7 ();
 sg13g2_fill_2 FILLER_78_14 ();
 sg13g2_fill_2 FILLER_78_39 ();
 sg13g2_decap_4 FILLER_78_46 ();
 sg13g2_fill_2 FILLER_78_54 ();
 sg13g2_fill_1 FILLER_78_87 ();
 sg13g2_fill_1 FILLER_78_93 ();
 sg13g2_fill_1 FILLER_78_109 ();
 sg13g2_fill_1 FILLER_78_115 ();
 sg13g2_fill_2 FILLER_78_172 ();
 sg13g2_decap_8 FILLER_78_182 ();
 sg13g2_fill_2 FILLER_78_189 ();
 sg13g2_fill_1 FILLER_78_191 ();
 sg13g2_decap_8 FILLER_78_222 ();
 sg13g2_fill_2 FILLER_78_229 ();
 sg13g2_fill_1 FILLER_78_264 ();
 sg13g2_fill_1 FILLER_78_284 ();
 sg13g2_fill_1 FILLER_78_290 ();
 sg13g2_fill_1 FILLER_78_296 ();
 sg13g2_fill_2 FILLER_78_302 ();
 sg13g2_decap_8 FILLER_78_309 ();
 sg13g2_fill_1 FILLER_78_316 ();
 sg13g2_decap_4 FILLER_78_325 ();
 sg13g2_fill_1 FILLER_78_329 ();
 sg13g2_fill_1 FILLER_78_349 ();
 sg13g2_fill_1 FILLER_78_353 ();
 sg13g2_fill_1 FILLER_78_384 ();
 sg13g2_fill_1 FILLER_78_388 ();
 sg13g2_fill_1 FILLER_78_394 ();
 sg13g2_fill_1 FILLER_78_403 ();
 sg13g2_decap_8 FILLER_79_0 ();
 sg13g2_decap_8 FILLER_79_7 ();
 sg13g2_decap_8 FILLER_79_14 ();
 sg13g2_decap_4 FILLER_79_21 ();
 sg13g2_fill_1 FILLER_79_25 ();
 sg13g2_fill_2 FILLER_79_44 ();
 sg13g2_fill_1 FILLER_79_77 ();
 sg13g2_fill_1 FILLER_79_83 ();
 sg13g2_fill_2 FILLER_79_89 ();
 sg13g2_fill_1 FILLER_79_91 ();
 sg13g2_fill_2 FILLER_79_101 ();
 sg13g2_fill_1 FILLER_79_108 ();
 sg13g2_fill_1 FILLER_79_113 ();
 sg13g2_fill_2 FILLER_79_122 ();
 sg13g2_decap_4 FILLER_79_128 ();
 sg13g2_fill_1 FILLER_79_132 ();
 sg13g2_fill_2 FILLER_79_137 ();
 sg13g2_fill_1 FILLER_79_143 ();
 sg13g2_fill_1 FILLER_79_148 ();
 sg13g2_fill_1 FILLER_79_153 ();
 sg13g2_fill_2 FILLER_79_180 ();
 sg13g2_fill_1 FILLER_79_182 ();
 sg13g2_decap_4 FILLER_79_209 ();
 sg13g2_fill_2 FILLER_79_213 ();
 sg13g2_fill_1 FILLER_79_266 ();
 sg13g2_decap_4 FILLER_79_272 ();
 sg13g2_fill_2 FILLER_79_276 ();
 sg13g2_decap_8 FILLER_79_282 ();
 sg13g2_fill_2 FILLER_79_298 ();
 sg13g2_fill_1 FILLER_79_300 ();
 sg13g2_fill_1 FILLER_79_305 ();
 sg13g2_fill_2 FILLER_79_337 ();
 sg13g2_fill_1 FILLER_79_339 ();
 sg13g2_decap_8 FILLER_79_344 ();
 sg13g2_fill_1 FILLER_79_351 ();
 sg13g2_fill_2 FILLER_79_356 ();
 sg13g2_fill_1 FILLER_79_372 ();
 sg13g2_fill_2 FILLER_79_390 ();
 sg13g2_fill_2 FILLER_79_409 ();
 sg13g2_decap_8 FILLER_79_419 ();
 sg13g2_decap_4 FILLER_79_426 ();
 sg13g2_decap_8 FILLER_80_0 ();
 sg13g2_decap_8 FILLER_80_7 ();
 sg13g2_decap_8 FILLER_80_14 ();
 sg13g2_decap_8 FILLER_80_21 ();
 sg13g2_decap_8 FILLER_80_28 ();
 sg13g2_decap_8 FILLER_80_35 ();
 sg13g2_fill_2 FILLER_80_42 ();
 sg13g2_fill_1 FILLER_80_57 ();
 sg13g2_fill_2 FILLER_80_62 ();
 sg13g2_fill_1 FILLER_80_64 ();
 sg13g2_decap_4 FILLER_80_133 ();
 sg13g2_decap_4 FILLER_80_209 ();
 sg13g2_fill_1 FILLER_80_243 ();
 sg13g2_decap_8 FILLER_80_322 ();
 sg13g2_decap_4 FILLER_80_329 ();
endmodule
