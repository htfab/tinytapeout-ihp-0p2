module tt_um_urish_giant_ringosc (clk,
    ena,
    rst_n,
    ui_in,
    uio_in,
    uio_oe,
    uio_out,
    uo_out);
 input clk;
 input ena;
 input rst_n;
 input [7:0] ui_in;
 input [7:0] uio_in;
 output [7:0] uio_oe;
 output [7:0] uio_out;
 output [7:0] uo_out;

 wire net18;
 wire \inv_in[1000] ;
 wire \inv_in[1001] ;
 wire \inv_in[1002] ;
 wire \inv_in[1003] ;
 wire \inv_in[1004] ;
 wire \inv_in[1005] ;
 wire \inv_in[1006] ;
 wire \inv_in[1007] ;
 wire \inv_in[1008] ;
 wire \inv_in[1009] ;
 wire \inv_in[100] ;
 wire \inv_in[1010] ;
 wire \inv_in[1011] ;
 wire \inv_in[1012] ;
 wire \inv_in[1013] ;
 wire \inv_in[1014] ;
 wire \inv_in[1015] ;
 wire \inv_in[1016] ;
 wire \inv_in[1017] ;
 wire \inv_in[1018] ;
 wire \inv_in[1019] ;
 wire \inv_in[101] ;
 wire \inv_in[1020] ;
 wire \inv_in[1021] ;
 wire \inv_in[1022] ;
 wire \inv_in[1023] ;
 wire \inv_in[1024] ;
 wire \inv_in[1025] ;
 wire \inv_in[1026] ;
 wire \inv_in[1027] ;
 wire \inv_in[1028] ;
 wire \inv_in[1029] ;
 wire \inv_in[102] ;
 wire \inv_in[1030] ;
 wire \inv_in[1031] ;
 wire \inv_in[1032] ;
 wire \inv_in[1033] ;
 wire \inv_in[1034] ;
 wire \inv_in[1035] ;
 wire \inv_in[1036] ;
 wire \inv_in[1037] ;
 wire \inv_in[1038] ;
 wire \inv_in[1039] ;
 wire \inv_in[103] ;
 wire \inv_in[1040] ;
 wire \inv_in[1041] ;
 wire \inv_in[1042] ;
 wire \inv_in[1043] ;
 wire \inv_in[1044] ;
 wire \inv_in[1045] ;
 wire \inv_in[1046] ;
 wire \inv_in[1047] ;
 wire \inv_in[1048] ;
 wire \inv_in[1049] ;
 wire \inv_in[104] ;
 wire \inv_in[1050] ;
 wire \inv_in[1051] ;
 wire \inv_in[1052] ;
 wire \inv_in[1053] ;
 wire \inv_in[1054] ;
 wire \inv_in[1055] ;
 wire \inv_in[1056] ;
 wire \inv_in[1057] ;
 wire \inv_in[1058] ;
 wire \inv_in[1059] ;
 wire \inv_in[105] ;
 wire \inv_in[1060] ;
 wire \inv_in[1061] ;
 wire \inv_in[1062] ;
 wire \inv_in[1063] ;
 wire \inv_in[1064] ;
 wire \inv_in[1065] ;
 wire \inv_in[1066] ;
 wire \inv_in[1067] ;
 wire \inv_in[1068] ;
 wire \inv_in[1069] ;
 wire \inv_in[106] ;
 wire \inv_in[1070] ;
 wire \inv_in[1071] ;
 wire \inv_in[1072] ;
 wire \inv_in[1073] ;
 wire \inv_in[1074] ;
 wire \inv_in[1075] ;
 wire \inv_in[1076] ;
 wire \inv_in[1077] ;
 wire \inv_in[1078] ;
 wire \inv_in[1079] ;
 wire \inv_in[107] ;
 wire \inv_in[1080] ;
 wire \inv_in[1081] ;
 wire \inv_in[1082] ;
 wire \inv_in[1083] ;
 wire \inv_in[1084] ;
 wire \inv_in[1085] ;
 wire \inv_in[1086] ;
 wire \inv_in[1087] ;
 wire \inv_in[1088] ;
 wire \inv_in[1089] ;
 wire \inv_in[108] ;
 wire \inv_in[1090] ;
 wire \inv_in[1091] ;
 wire \inv_in[1092] ;
 wire \inv_in[1093] ;
 wire \inv_in[1094] ;
 wire \inv_in[1095] ;
 wire \inv_in[1096] ;
 wire \inv_in[1097] ;
 wire \inv_in[1098] ;
 wire \inv_in[1099] ;
 wire \inv_in[109] ;
 wire \inv_in[10] ;
 wire \inv_in[1100] ;
 wire \inv_in[1101] ;
 wire \inv_in[1102] ;
 wire \inv_in[1103] ;
 wire \inv_in[1104] ;
 wire \inv_in[1105] ;
 wire \inv_in[1106] ;
 wire \inv_in[1107] ;
 wire \inv_in[1108] ;
 wire \inv_in[1109] ;
 wire \inv_in[110] ;
 wire \inv_in[1110] ;
 wire \inv_in[1111] ;
 wire \inv_in[1112] ;
 wire \inv_in[1113] ;
 wire \inv_in[1114] ;
 wire \inv_in[1115] ;
 wire \inv_in[1116] ;
 wire \inv_in[1117] ;
 wire \inv_in[1118] ;
 wire \inv_in[1119] ;
 wire \inv_in[111] ;
 wire \inv_in[1120] ;
 wire \inv_in[1121] ;
 wire \inv_in[1122] ;
 wire \inv_in[1123] ;
 wire \inv_in[1124] ;
 wire \inv_in[1125] ;
 wire \inv_in[1126] ;
 wire \inv_in[1127] ;
 wire \inv_in[1128] ;
 wire \inv_in[1129] ;
 wire \inv_in[112] ;
 wire \inv_in[1130] ;
 wire \inv_in[1131] ;
 wire \inv_in[1132] ;
 wire \inv_in[1133] ;
 wire \inv_in[1134] ;
 wire \inv_in[1135] ;
 wire \inv_in[1136] ;
 wire \inv_in[1137] ;
 wire \inv_in[1138] ;
 wire \inv_in[1139] ;
 wire \inv_in[113] ;
 wire \inv_in[1140] ;
 wire \inv_in[1141] ;
 wire \inv_in[1142] ;
 wire \inv_in[1143] ;
 wire \inv_in[1144] ;
 wire \inv_in[1145] ;
 wire \inv_in[1146] ;
 wire \inv_in[1147] ;
 wire \inv_in[1148] ;
 wire \inv_in[1149] ;
 wire \inv_in[114] ;
 wire \inv_in[1150] ;
 wire \inv_in[1151] ;
 wire \inv_in[1152] ;
 wire \inv_in[1153] ;
 wire \inv_in[1154] ;
 wire \inv_in[1155] ;
 wire \inv_in[1156] ;
 wire \inv_in[1157] ;
 wire \inv_in[1158] ;
 wire \inv_in[1159] ;
 wire \inv_in[115] ;
 wire \inv_in[1160] ;
 wire \inv_in[1161] ;
 wire \inv_in[1162] ;
 wire \inv_in[1163] ;
 wire \inv_in[1164] ;
 wire \inv_in[1165] ;
 wire \inv_in[1166] ;
 wire \inv_in[1167] ;
 wire \inv_in[1168] ;
 wire \inv_in[1169] ;
 wire \inv_in[116] ;
 wire \inv_in[1170] ;
 wire \inv_in[1171] ;
 wire \inv_in[1172] ;
 wire \inv_in[1173] ;
 wire \inv_in[1174] ;
 wire \inv_in[1175] ;
 wire \inv_in[1176] ;
 wire \inv_in[1177] ;
 wire \inv_in[1178] ;
 wire \inv_in[1179] ;
 wire \inv_in[117] ;
 wire \inv_in[1180] ;
 wire \inv_in[1181] ;
 wire \inv_in[1182] ;
 wire \inv_in[1183] ;
 wire \inv_in[1184] ;
 wire \inv_in[1185] ;
 wire \inv_in[1186] ;
 wire \inv_in[1187] ;
 wire \inv_in[1188] ;
 wire \inv_in[1189] ;
 wire \inv_in[118] ;
 wire \inv_in[1190] ;
 wire \inv_in[1191] ;
 wire \inv_in[1192] ;
 wire \inv_in[1193] ;
 wire \inv_in[1194] ;
 wire \inv_in[1195] ;
 wire \inv_in[1196] ;
 wire \inv_in[1197] ;
 wire \inv_in[1198] ;
 wire \inv_in[1199] ;
 wire \inv_in[119] ;
 wire \inv_in[11] ;
 wire \inv_in[1200] ;
 wire \inv_in[1201] ;
 wire \inv_in[1202] ;
 wire \inv_in[1203] ;
 wire \inv_in[1204] ;
 wire \inv_in[1205] ;
 wire \inv_in[1206] ;
 wire \inv_in[1207] ;
 wire \inv_in[1208] ;
 wire \inv_in[1209] ;
 wire \inv_in[120] ;
 wire \inv_in[1210] ;
 wire \inv_in[1211] ;
 wire \inv_in[1212] ;
 wire \inv_in[1213] ;
 wire \inv_in[1214] ;
 wire \inv_in[1215] ;
 wire \inv_in[1216] ;
 wire \inv_in[1217] ;
 wire \inv_in[1218] ;
 wire \inv_in[1219] ;
 wire \inv_in[121] ;
 wire \inv_in[1220] ;
 wire \inv_in[1221] ;
 wire \inv_in[1222] ;
 wire \inv_in[1223] ;
 wire \inv_in[1224] ;
 wire \inv_in[1225] ;
 wire \inv_in[1226] ;
 wire \inv_in[1227] ;
 wire \inv_in[1228] ;
 wire \inv_in[1229] ;
 wire \inv_in[122] ;
 wire \inv_in[1230] ;
 wire \inv_in[1231] ;
 wire \inv_in[1232] ;
 wire \inv_in[1233] ;
 wire \inv_in[1234] ;
 wire \inv_in[1235] ;
 wire \inv_in[1236] ;
 wire \inv_in[1237] ;
 wire \inv_in[1238] ;
 wire \inv_in[1239] ;
 wire \inv_in[123] ;
 wire \inv_in[1240] ;
 wire \inv_in[1241] ;
 wire \inv_in[1242] ;
 wire \inv_in[1243] ;
 wire \inv_in[1244] ;
 wire \inv_in[1245] ;
 wire \inv_in[1246] ;
 wire \inv_in[1247] ;
 wire \inv_in[1248] ;
 wire \inv_in[1249] ;
 wire \inv_in[124] ;
 wire \inv_in[1250] ;
 wire \inv_in[1251] ;
 wire \inv_in[1252] ;
 wire \inv_in[1253] ;
 wire \inv_in[1254] ;
 wire \inv_in[1255] ;
 wire \inv_in[1256] ;
 wire \inv_in[1257] ;
 wire \inv_in[1258] ;
 wire \inv_in[1259] ;
 wire \inv_in[125] ;
 wire \inv_in[1260] ;
 wire \inv_in[1261] ;
 wire \inv_in[1262] ;
 wire \inv_in[1263] ;
 wire \inv_in[1264] ;
 wire \inv_in[1265] ;
 wire \inv_in[1266] ;
 wire \inv_in[1267] ;
 wire \inv_in[1268] ;
 wire \inv_in[1269] ;
 wire \inv_in[126] ;
 wire \inv_in[1270] ;
 wire \inv_in[1271] ;
 wire \inv_in[1272] ;
 wire \inv_in[1273] ;
 wire \inv_in[1274] ;
 wire \inv_in[1275] ;
 wire \inv_in[1276] ;
 wire \inv_in[1277] ;
 wire \inv_in[1278] ;
 wire \inv_in[1279] ;
 wire \inv_in[127] ;
 wire \inv_in[1280] ;
 wire \inv_in[1281] ;
 wire \inv_in[1282] ;
 wire \inv_in[1283] ;
 wire \inv_in[1284] ;
 wire \inv_in[1285] ;
 wire \inv_in[1286] ;
 wire \inv_in[1287] ;
 wire \inv_in[1288] ;
 wire \inv_in[1289] ;
 wire \inv_in[128] ;
 wire \inv_in[1290] ;
 wire \inv_in[1291] ;
 wire \inv_in[1292] ;
 wire \inv_in[1293] ;
 wire \inv_in[1294] ;
 wire \inv_in[1295] ;
 wire \inv_in[1296] ;
 wire \inv_in[1297] ;
 wire \inv_in[1298] ;
 wire \inv_in[1299] ;
 wire \inv_in[129] ;
 wire \inv_in[12] ;
 wire \inv_in[1300] ;
 wire \inv_in[1301] ;
 wire \inv_in[1302] ;
 wire \inv_in[1303] ;
 wire \inv_in[1304] ;
 wire \inv_in[1305] ;
 wire \inv_in[1306] ;
 wire \inv_in[1307] ;
 wire \inv_in[1308] ;
 wire \inv_in[1309] ;
 wire \inv_in[130] ;
 wire \inv_in[1310] ;
 wire \inv_in[1311] ;
 wire \inv_in[1312] ;
 wire \inv_in[1313] ;
 wire \inv_in[1314] ;
 wire \inv_in[1315] ;
 wire \inv_in[1316] ;
 wire \inv_in[1317] ;
 wire \inv_in[1318] ;
 wire \inv_in[1319] ;
 wire \inv_in[131] ;
 wire \inv_in[1320] ;
 wire \inv_in[1321] ;
 wire \inv_in[1322] ;
 wire \inv_in[1323] ;
 wire \inv_in[1324] ;
 wire \inv_in[1325] ;
 wire \inv_in[1326] ;
 wire \inv_in[1327] ;
 wire \inv_in[1328] ;
 wire \inv_in[1329] ;
 wire \inv_in[132] ;
 wire \inv_in[1330] ;
 wire \inv_in[1331] ;
 wire \inv_in[1332] ;
 wire \inv_in[1333] ;
 wire \inv_in[1334] ;
 wire \inv_in[1335] ;
 wire \inv_in[1336] ;
 wire \inv_in[1337] ;
 wire \inv_in[1338] ;
 wire \inv_in[1339] ;
 wire \inv_in[133] ;
 wire \inv_in[1340] ;
 wire \inv_in[1341] ;
 wire \inv_in[1342] ;
 wire \inv_in[1343] ;
 wire \inv_in[1344] ;
 wire \inv_in[1345] ;
 wire \inv_in[1346] ;
 wire \inv_in[1347] ;
 wire \inv_in[1348] ;
 wire \inv_in[1349] ;
 wire \inv_in[134] ;
 wire \inv_in[1350] ;
 wire \inv_in[1351] ;
 wire \inv_in[1352] ;
 wire \inv_in[1353] ;
 wire \inv_in[1354] ;
 wire \inv_in[1355] ;
 wire \inv_in[1356] ;
 wire \inv_in[1357] ;
 wire \inv_in[1358] ;
 wire \inv_in[1359] ;
 wire \inv_in[135] ;
 wire \inv_in[1360] ;
 wire \inv_in[1361] ;
 wire \inv_in[1362] ;
 wire \inv_in[1363] ;
 wire \inv_in[1364] ;
 wire \inv_in[1365] ;
 wire \inv_in[1366] ;
 wire \inv_in[1367] ;
 wire \inv_in[1368] ;
 wire \inv_in[1369] ;
 wire \inv_in[136] ;
 wire \inv_in[1370] ;
 wire \inv_in[1371] ;
 wire \inv_in[1372] ;
 wire \inv_in[1373] ;
 wire \inv_in[1374] ;
 wire \inv_in[1375] ;
 wire \inv_in[1376] ;
 wire \inv_in[1377] ;
 wire \inv_in[1378] ;
 wire \inv_in[1379] ;
 wire \inv_in[137] ;
 wire \inv_in[1380] ;
 wire \inv_in[1381] ;
 wire \inv_in[1382] ;
 wire \inv_in[1383] ;
 wire \inv_in[1384] ;
 wire \inv_in[1385] ;
 wire \inv_in[1386] ;
 wire \inv_in[1387] ;
 wire \inv_in[1388] ;
 wire \inv_in[1389] ;
 wire \inv_in[138] ;
 wire \inv_in[1390] ;
 wire \inv_in[1391] ;
 wire \inv_in[1392] ;
 wire \inv_in[1393] ;
 wire \inv_in[1394] ;
 wire \inv_in[1395] ;
 wire \inv_in[1396] ;
 wire \inv_in[1397] ;
 wire \inv_in[1398] ;
 wire \inv_in[1399] ;
 wire \inv_in[139] ;
 wire \inv_in[13] ;
 wire \inv_in[1400] ;
 wire \inv_in[1401] ;
 wire \inv_in[1402] ;
 wire \inv_in[1403] ;
 wire \inv_in[1404] ;
 wire \inv_in[1405] ;
 wire \inv_in[1406] ;
 wire \inv_in[1407] ;
 wire \inv_in[1408] ;
 wire \inv_in[1409] ;
 wire \inv_in[140] ;
 wire \inv_in[1410] ;
 wire \inv_in[1411] ;
 wire \inv_in[1412] ;
 wire \inv_in[1413] ;
 wire \inv_in[1414] ;
 wire \inv_in[1415] ;
 wire \inv_in[1416] ;
 wire \inv_in[1417] ;
 wire \inv_in[1418] ;
 wire \inv_in[1419] ;
 wire \inv_in[141] ;
 wire \inv_in[1420] ;
 wire \inv_in[1421] ;
 wire \inv_in[1422] ;
 wire \inv_in[1423] ;
 wire \inv_in[1424] ;
 wire \inv_in[1425] ;
 wire \inv_in[1426] ;
 wire \inv_in[1427] ;
 wire \inv_in[1428] ;
 wire \inv_in[1429] ;
 wire \inv_in[142] ;
 wire \inv_in[1430] ;
 wire \inv_in[1431] ;
 wire \inv_in[1432] ;
 wire \inv_in[1433] ;
 wire \inv_in[1434] ;
 wire \inv_in[1435] ;
 wire \inv_in[1436] ;
 wire \inv_in[1437] ;
 wire \inv_in[1438] ;
 wire \inv_in[1439] ;
 wire \inv_in[143] ;
 wire \inv_in[1440] ;
 wire \inv_in[1441] ;
 wire \inv_in[1442] ;
 wire \inv_in[1443] ;
 wire \inv_in[1444] ;
 wire \inv_in[1445] ;
 wire \inv_in[1446] ;
 wire \inv_in[1447] ;
 wire \inv_in[1448] ;
 wire \inv_in[1449] ;
 wire \inv_in[144] ;
 wire \inv_in[1450] ;
 wire \inv_in[1451] ;
 wire \inv_in[1452] ;
 wire \inv_in[1453] ;
 wire \inv_in[1454] ;
 wire \inv_in[1455] ;
 wire \inv_in[1456] ;
 wire \inv_in[1457] ;
 wire \inv_in[1458] ;
 wire \inv_in[1459] ;
 wire \inv_in[145] ;
 wire \inv_in[1460] ;
 wire \inv_in[1461] ;
 wire \inv_in[1462] ;
 wire \inv_in[1463] ;
 wire \inv_in[1464] ;
 wire \inv_in[1465] ;
 wire \inv_in[1466] ;
 wire \inv_in[1467] ;
 wire \inv_in[1468] ;
 wire \inv_in[1469] ;
 wire \inv_in[146] ;
 wire \inv_in[1470] ;
 wire \inv_in[1471] ;
 wire \inv_in[1472] ;
 wire \inv_in[1473] ;
 wire \inv_in[1474] ;
 wire \inv_in[1475] ;
 wire \inv_in[1476] ;
 wire \inv_in[1477] ;
 wire \inv_in[1478] ;
 wire \inv_in[1479] ;
 wire \inv_in[147] ;
 wire \inv_in[1480] ;
 wire \inv_in[1481] ;
 wire \inv_in[1482] ;
 wire \inv_in[1483] ;
 wire \inv_in[1484] ;
 wire \inv_in[1485] ;
 wire \inv_in[1486] ;
 wire \inv_in[1487] ;
 wire \inv_in[1488] ;
 wire \inv_in[1489] ;
 wire \inv_in[148] ;
 wire \inv_in[1490] ;
 wire \inv_in[1491] ;
 wire \inv_in[1492] ;
 wire \inv_in[1493] ;
 wire \inv_in[1494] ;
 wire \inv_in[1495] ;
 wire \inv_in[1496] ;
 wire \inv_in[1497] ;
 wire \inv_in[1498] ;
 wire \inv_in[1499] ;
 wire \inv_in[149] ;
 wire \inv_in[14] ;
 wire \inv_in[1500] ;
 wire \inv_in[1501] ;
 wire \inv_in[1502] ;
 wire \inv_in[1503] ;
 wire \inv_in[1504] ;
 wire \inv_in[1505] ;
 wire \inv_in[1506] ;
 wire \inv_in[1507] ;
 wire \inv_in[1508] ;
 wire \inv_in[1509] ;
 wire \inv_in[150] ;
 wire \inv_in[1510] ;
 wire \inv_in[1511] ;
 wire \inv_in[1512] ;
 wire \inv_in[1513] ;
 wire \inv_in[1514] ;
 wire \inv_in[1515] ;
 wire \inv_in[1516] ;
 wire \inv_in[1517] ;
 wire \inv_in[1518] ;
 wire \inv_in[1519] ;
 wire \inv_in[151] ;
 wire \inv_in[1520] ;
 wire \inv_in[1521] ;
 wire \inv_in[1522] ;
 wire \inv_in[1523] ;
 wire \inv_in[1524] ;
 wire \inv_in[1525] ;
 wire \inv_in[1526] ;
 wire \inv_in[1527] ;
 wire \inv_in[1528] ;
 wire \inv_in[1529] ;
 wire \inv_in[152] ;
 wire \inv_in[1530] ;
 wire \inv_in[1531] ;
 wire \inv_in[1532] ;
 wire \inv_in[1533] ;
 wire \inv_in[1534] ;
 wire \inv_in[1535] ;
 wire \inv_in[1536] ;
 wire \inv_in[1537] ;
 wire \inv_in[1538] ;
 wire \inv_in[1539] ;
 wire \inv_in[153] ;
 wire \inv_in[1540] ;
 wire \inv_in[1541] ;
 wire \inv_in[1542] ;
 wire \inv_in[1543] ;
 wire \inv_in[1544] ;
 wire \inv_in[1545] ;
 wire \inv_in[1546] ;
 wire \inv_in[1547] ;
 wire \inv_in[1548] ;
 wire \inv_in[1549] ;
 wire \inv_in[154] ;
 wire \inv_in[1550] ;
 wire \inv_in[1551] ;
 wire \inv_in[1552] ;
 wire \inv_in[1553] ;
 wire \inv_in[1554] ;
 wire \inv_in[1555] ;
 wire \inv_in[1556] ;
 wire \inv_in[1557] ;
 wire \inv_in[1558] ;
 wire \inv_in[1559] ;
 wire \inv_in[155] ;
 wire \inv_in[1560] ;
 wire \inv_in[1561] ;
 wire \inv_in[1562] ;
 wire \inv_in[1563] ;
 wire \inv_in[1564] ;
 wire \inv_in[1565] ;
 wire \inv_in[1566] ;
 wire \inv_in[1567] ;
 wire \inv_in[1568] ;
 wire \inv_in[1569] ;
 wire \inv_in[156] ;
 wire \inv_in[1570] ;
 wire \inv_in[1571] ;
 wire \inv_in[1572] ;
 wire \inv_in[1573] ;
 wire \inv_in[1574] ;
 wire \inv_in[1575] ;
 wire \inv_in[1576] ;
 wire \inv_in[1577] ;
 wire \inv_in[1578] ;
 wire \inv_in[1579] ;
 wire \inv_in[157] ;
 wire \inv_in[1580] ;
 wire \inv_in[1581] ;
 wire \inv_in[1582] ;
 wire \inv_in[1583] ;
 wire \inv_in[1584] ;
 wire \inv_in[1585] ;
 wire \inv_in[1586] ;
 wire \inv_in[1587] ;
 wire \inv_in[1588] ;
 wire \inv_in[1589] ;
 wire \inv_in[158] ;
 wire \inv_in[1590] ;
 wire \inv_in[1591] ;
 wire \inv_in[1592] ;
 wire \inv_in[1593] ;
 wire \inv_in[1594] ;
 wire \inv_in[1595] ;
 wire \inv_in[1596] ;
 wire \inv_in[1597] ;
 wire \inv_in[1598] ;
 wire \inv_in[1599] ;
 wire \inv_in[159] ;
 wire \inv_in[15] ;
 wire \inv_in[1600] ;
 wire \inv_in[1601] ;
 wire \inv_in[1602] ;
 wire \inv_in[1603] ;
 wire \inv_in[1604] ;
 wire \inv_in[1605] ;
 wire \inv_in[1606] ;
 wire \inv_in[1607] ;
 wire \inv_in[1608] ;
 wire \inv_in[1609] ;
 wire \inv_in[160] ;
 wire \inv_in[1610] ;
 wire \inv_in[1611] ;
 wire \inv_in[1612] ;
 wire \inv_in[1613] ;
 wire \inv_in[1614] ;
 wire \inv_in[1615] ;
 wire \inv_in[1616] ;
 wire \inv_in[1617] ;
 wire \inv_in[1618] ;
 wire \inv_in[1619] ;
 wire \inv_in[161] ;
 wire \inv_in[1620] ;
 wire \inv_in[1621] ;
 wire \inv_in[1622] ;
 wire \inv_in[1623] ;
 wire \inv_in[1624] ;
 wire \inv_in[1625] ;
 wire \inv_in[1626] ;
 wire \inv_in[1627] ;
 wire \inv_in[1628] ;
 wire \inv_in[1629] ;
 wire \inv_in[162] ;
 wire \inv_in[1630] ;
 wire \inv_in[1631] ;
 wire \inv_in[1632] ;
 wire \inv_in[1633] ;
 wire \inv_in[1634] ;
 wire \inv_in[1635] ;
 wire \inv_in[1636] ;
 wire \inv_in[1637] ;
 wire \inv_in[1638] ;
 wire \inv_in[1639] ;
 wire \inv_in[163] ;
 wire \inv_in[1640] ;
 wire \inv_in[1641] ;
 wire \inv_in[1642] ;
 wire \inv_in[1643] ;
 wire \inv_in[1644] ;
 wire \inv_in[1645] ;
 wire \inv_in[1646] ;
 wire \inv_in[1647] ;
 wire \inv_in[1648] ;
 wire \inv_in[1649] ;
 wire \inv_in[164] ;
 wire \inv_in[1650] ;
 wire \inv_in[1651] ;
 wire \inv_in[1652] ;
 wire \inv_in[1653] ;
 wire \inv_in[1654] ;
 wire \inv_in[1655] ;
 wire \inv_in[1656] ;
 wire \inv_in[1657] ;
 wire \inv_in[1658] ;
 wire \inv_in[1659] ;
 wire \inv_in[165] ;
 wire \inv_in[1660] ;
 wire \inv_in[1661] ;
 wire \inv_in[1662] ;
 wire \inv_in[1663] ;
 wire \inv_in[1664] ;
 wire \inv_in[1665] ;
 wire \inv_in[1666] ;
 wire \inv_in[1667] ;
 wire \inv_in[1668] ;
 wire \inv_in[1669] ;
 wire \inv_in[166] ;
 wire \inv_in[1670] ;
 wire \inv_in[1671] ;
 wire \inv_in[1672] ;
 wire \inv_in[1673] ;
 wire \inv_in[1674] ;
 wire \inv_in[1675] ;
 wire \inv_in[1676] ;
 wire \inv_in[1677] ;
 wire \inv_in[1678] ;
 wire \inv_in[1679] ;
 wire \inv_in[167] ;
 wire \inv_in[1680] ;
 wire \inv_in[1681] ;
 wire \inv_in[1682] ;
 wire \inv_in[1683] ;
 wire \inv_in[1684] ;
 wire \inv_in[1685] ;
 wire \inv_in[1686] ;
 wire \inv_in[1687] ;
 wire \inv_in[1688] ;
 wire \inv_in[1689] ;
 wire \inv_in[168] ;
 wire \inv_in[1690] ;
 wire \inv_in[1691] ;
 wire \inv_in[1692] ;
 wire \inv_in[1693] ;
 wire \inv_in[1694] ;
 wire \inv_in[1695] ;
 wire \inv_in[1696] ;
 wire \inv_in[1697] ;
 wire \inv_in[1698] ;
 wire \inv_in[1699] ;
 wire \inv_in[169] ;
 wire \inv_in[16] ;
 wire \inv_in[1700] ;
 wire \inv_in[1701] ;
 wire \inv_in[1702] ;
 wire \inv_in[1703] ;
 wire \inv_in[1704] ;
 wire \inv_in[1705] ;
 wire \inv_in[1706] ;
 wire \inv_in[1707] ;
 wire \inv_in[1708] ;
 wire \inv_in[1709] ;
 wire \inv_in[170] ;
 wire \inv_in[1710] ;
 wire \inv_in[1711] ;
 wire \inv_in[1712] ;
 wire \inv_in[1713] ;
 wire \inv_in[1714] ;
 wire \inv_in[1715] ;
 wire \inv_in[1716] ;
 wire \inv_in[1717] ;
 wire \inv_in[1718] ;
 wire \inv_in[1719] ;
 wire \inv_in[171] ;
 wire \inv_in[1720] ;
 wire \inv_in[1721] ;
 wire \inv_in[1722] ;
 wire \inv_in[1723] ;
 wire \inv_in[1724] ;
 wire \inv_in[1725] ;
 wire \inv_in[1726] ;
 wire \inv_in[1727] ;
 wire \inv_in[1728] ;
 wire \inv_in[1729] ;
 wire \inv_in[172] ;
 wire \inv_in[1730] ;
 wire \inv_in[1731] ;
 wire \inv_in[1732] ;
 wire \inv_in[1733] ;
 wire \inv_in[1734] ;
 wire \inv_in[1735] ;
 wire \inv_in[1736] ;
 wire \inv_in[1737] ;
 wire \inv_in[1738] ;
 wire \inv_in[1739] ;
 wire \inv_in[173] ;
 wire \inv_in[1740] ;
 wire \inv_in[1741] ;
 wire \inv_in[1742] ;
 wire \inv_in[1743] ;
 wire \inv_in[1744] ;
 wire \inv_in[1745] ;
 wire \inv_in[1746] ;
 wire \inv_in[1747] ;
 wire \inv_in[1748] ;
 wire \inv_in[1749] ;
 wire \inv_in[174] ;
 wire \inv_in[1750] ;
 wire \inv_in[1751] ;
 wire \inv_in[1752] ;
 wire \inv_in[1753] ;
 wire \inv_in[1754] ;
 wire \inv_in[1755] ;
 wire \inv_in[1756] ;
 wire \inv_in[1757] ;
 wire \inv_in[1758] ;
 wire \inv_in[1759] ;
 wire \inv_in[175] ;
 wire \inv_in[1760] ;
 wire \inv_in[1761] ;
 wire \inv_in[1762] ;
 wire \inv_in[1763] ;
 wire \inv_in[1764] ;
 wire \inv_in[1765] ;
 wire \inv_in[1766] ;
 wire \inv_in[1767] ;
 wire \inv_in[1768] ;
 wire \inv_in[1769] ;
 wire \inv_in[176] ;
 wire \inv_in[1770] ;
 wire \inv_in[1771] ;
 wire \inv_in[1772] ;
 wire \inv_in[1773] ;
 wire \inv_in[1774] ;
 wire \inv_in[1775] ;
 wire \inv_in[1776] ;
 wire \inv_in[1777] ;
 wire \inv_in[1778] ;
 wire \inv_in[1779] ;
 wire \inv_in[177] ;
 wire \inv_in[1780] ;
 wire \inv_in[1781] ;
 wire \inv_in[1782] ;
 wire \inv_in[1783] ;
 wire \inv_in[1784] ;
 wire \inv_in[1785] ;
 wire \inv_in[1786] ;
 wire \inv_in[1787] ;
 wire \inv_in[1788] ;
 wire \inv_in[1789] ;
 wire \inv_in[178] ;
 wire \inv_in[1790] ;
 wire \inv_in[1791] ;
 wire \inv_in[1792] ;
 wire \inv_in[1793] ;
 wire \inv_in[1794] ;
 wire \inv_in[1795] ;
 wire \inv_in[1796] ;
 wire \inv_in[1797] ;
 wire \inv_in[1798] ;
 wire \inv_in[1799] ;
 wire \inv_in[179] ;
 wire \inv_in[17] ;
 wire \inv_in[1800] ;
 wire \inv_in[1801] ;
 wire \inv_in[1802] ;
 wire \inv_in[1803] ;
 wire \inv_in[1804] ;
 wire \inv_in[1805] ;
 wire \inv_in[1806] ;
 wire \inv_in[1807] ;
 wire \inv_in[1808] ;
 wire \inv_in[1809] ;
 wire \inv_in[180] ;
 wire \inv_in[1810] ;
 wire \inv_in[1811] ;
 wire \inv_in[1812] ;
 wire \inv_in[1813] ;
 wire \inv_in[1814] ;
 wire \inv_in[1815] ;
 wire \inv_in[1816] ;
 wire \inv_in[1817] ;
 wire \inv_in[1818] ;
 wire \inv_in[1819] ;
 wire \inv_in[181] ;
 wire \inv_in[1820] ;
 wire \inv_in[1821] ;
 wire \inv_in[1822] ;
 wire \inv_in[1823] ;
 wire \inv_in[1824] ;
 wire \inv_in[1825] ;
 wire \inv_in[1826] ;
 wire \inv_in[1827] ;
 wire \inv_in[1828] ;
 wire \inv_in[1829] ;
 wire \inv_in[182] ;
 wire \inv_in[1830] ;
 wire \inv_in[1831] ;
 wire \inv_in[1832] ;
 wire \inv_in[1833] ;
 wire \inv_in[1834] ;
 wire \inv_in[1835] ;
 wire \inv_in[1836] ;
 wire \inv_in[1837] ;
 wire \inv_in[1838] ;
 wire \inv_in[1839] ;
 wire \inv_in[183] ;
 wire \inv_in[1840] ;
 wire \inv_in[1841] ;
 wire \inv_in[1842] ;
 wire \inv_in[1843] ;
 wire \inv_in[1844] ;
 wire \inv_in[1845] ;
 wire \inv_in[1846] ;
 wire \inv_in[1847] ;
 wire \inv_in[1848] ;
 wire \inv_in[1849] ;
 wire \inv_in[184] ;
 wire \inv_in[1850] ;
 wire \inv_in[1851] ;
 wire \inv_in[1852] ;
 wire \inv_in[1853] ;
 wire \inv_in[1854] ;
 wire \inv_in[1855] ;
 wire \inv_in[1856] ;
 wire \inv_in[1857] ;
 wire \inv_in[1858] ;
 wire \inv_in[1859] ;
 wire \inv_in[185] ;
 wire \inv_in[1860] ;
 wire \inv_in[1861] ;
 wire \inv_in[1862] ;
 wire \inv_in[1863] ;
 wire \inv_in[1864] ;
 wire \inv_in[1865] ;
 wire \inv_in[1866] ;
 wire \inv_in[1867] ;
 wire \inv_in[1868] ;
 wire \inv_in[1869] ;
 wire \inv_in[186] ;
 wire \inv_in[1870] ;
 wire \inv_in[1871] ;
 wire \inv_in[1872] ;
 wire \inv_in[1873] ;
 wire \inv_in[1874] ;
 wire \inv_in[1875] ;
 wire \inv_in[1876] ;
 wire \inv_in[1877] ;
 wire \inv_in[1878] ;
 wire \inv_in[1879] ;
 wire \inv_in[187] ;
 wire \inv_in[1880] ;
 wire \inv_in[1881] ;
 wire \inv_in[1882] ;
 wire \inv_in[1883] ;
 wire \inv_in[1884] ;
 wire \inv_in[1885] ;
 wire \inv_in[1886] ;
 wire \inv_in[1887] ;
 wire \inv_in[1888] ;
 wire \inv_in[1889] ;
 wire \inv_in[188] ;
 wire \inv_in[1890] ;
 wire \inv_in[1891] ;
 wire \inv_in[1892] ;
 wire \inv_in[1893] ;
 wire \inv_in[1894] ;
 wire \inv_in[1895] ;
 wire \inv_in[1896] ;
 wire \inv_in[1897] ;
 wire \inv_in[1898] ;
 wire \inv_in[1899] ;
 wire \inv_in[189] ;
 wire \inv_in[18] ;
 wire \inv_in[1900] ;
 wire \inv_in[1901] ;
 wire \inv_in[1902] ;
 wire \inv_in[1903] ;
 wire \inv_in[1904] ;
 wire \inv_in[1905] ;
 wire \inv_in[1906] ;
 wire \inv_in[1907] ;
 wire \inv_in[1908] ;
 wire \inv_in[1909] ;
 wire \inv_in[190] ;
 wire \inv_in[1910] ;
 wire \inv_in[1911] ;
 wire \inv_in[1912] ;
 wire \inv_in[1913] ;
 wire \inv_in[1914] ;
 wire \inv_in[1915] ;
 wire \inv_in[1916] ;
 wire \inv_in[1917] ;
 wire \inv_in[1918] ;
 wire \inv_in[1919] ;
 wire \inv_in[191] ;
 wire \inv_in[1920] ;
 wire \inv_in[1921] ;
 wire \inv_in[1922] ;
 wire \inv_in[1923] ;
 wire \inv_in[1924] ;
 wire \inv_in[1925] ;
 wire \inv_in[1926] ;
 wire \inv_in[1927] ;
 wire \inv_in[1928] ;
 wire \inv_in[1929] ;
 wire \inv_in[192] ;
 wire \inv_in[1930] ;
 wire \inv_in[1931] ;
 wire \inv_in[1932] ;
 wire \inv_in[1933] ;
 wire \inv_in[1934] ;
 wire \inv_in[1935] ;
 wire \inv_in[1936] ;
 wire \inv_in[1937] ;
 wire \inv_in[1938] ;
 wire \inv_in[1939] ;
 wire \inv_in[193] ;
 wire \inv_in[1940] ;
 wire \inv_in[1941] ;
 wire \inv_in[1942] ;
 wire \inv_in[1943] ;
 wire \inv_in[1944] ;
 wire \inv_in[1945] ;
 wire \inv_in[1946] ;
 wire \inv_in[1947] ;
 wire \inv_in[1948] ;
 wire \inv_in[1949] ;
 wire \inv_in[194] ;
 wire \inv_in[1950] ;
 wire \inv_in[1951] ;
 wire \inv_in[1952] ;
 wire \inv_in[1953] ;
 wire \inv_in[1954] ;
 wire \inv_in[1955] ;
 wire \inv_in[1956] ;
 wire \inv_in[1957] ;
 wire \inv_in[1958] ;
 wire \inv_in[1959] ;
 wire \inv_in[195] ;
 wire \inv_in[1960] ;
 wire \inv_in[1961] ;
 wire \inv_in[1962] ;
 wire \inv_in[1963] ;
 wire \inv_in[1964] ;
 wire \inv_in[1965] ;
 wire \inv_in[1966] ;
 wire \inv_in[1967] ;
 wire \inv_in[1968] ;
 wire \inv_in[1969] ;
 wire \inv_in[196] ;
 wire \inv_in[1970] ;
 wire \inv_in[1971] ;
 wire \inv_in[1972] ;
 wire \inv_in[1973] ;
 wire \inv_in[1974] ;
 wire \inv_in[1975] ;
 wire \inv_in[1976] ;
 wire \inv_in[1977] ;
 wire \inv_in[1978] ;
 wire \inv_in[1979] ;
 wire \inv_in[197] ;
 wire \inv_in[1980] ;
 wire \inv_in[1981] ;
 wire \inv_in[1982] ;
 wire \inv_in[1983] ;
 wire \inv_in[1984] ;
 wire \inv_in[1985] ;
 wire \inv_in[1986] ;
 wire \inv_in[1987] ;
 wire \inv_in[1988] ;
 wire \inv_in[1989] ;
 wire \inv_in[198] ;
 wire \inv_in[1990] ;
 wire \inv_in[1991] ;
 wire \inv_in[1992] ;
 wire \inv_in[1993] ;
 wire \inv_in[1994] ;
 wire \inv_in[1995] ;
 wire \inv_in[1996] ;
 wire \inv_in[1997] ;
 wire \inv_in[1998] ;
 wire \inv_in[1999] ;
 wire \inv_in[199] ;
 wire \inv_in[19] ;
 wire \inv_in[1] ;
 wire \inv_in[2000] ;
 wire \inv_in[2001] ;
 wire \inv_in[2002] ;
 wire \inv_in[2003] ;
 wire \inv_in[2004] ;
 wire \inv_in[2005] ;
 wire \inv_in[2006] ;
 wire \inv_in[2007] ;
 wire \inv_in[2008] ;
 wire \inv_in[2009] ;
 wire \inv_in[200] ;
 wire \inv_in[2010] ;
 wire \inv_in[2011] ;
 wire \inv_in[2012] ;
 wire \inv_in[2013] ;
 wire \inv_in[2014] ;
 wire \inv_in[2015] ;
 wire \inv_in[2016] ;
 wire \inv_in[2017] ;
 wire \inv_in[2018] ;
 wire \inv_in[2019] ;
 wire \inv_in[201] ;
 wire \inv_in[2020] ;
 wire \inv_in[2021] ;
 wire \inv_in[2022] ;
 wire \inv_in[2023] ;
 wire \inv_in[2024] ;
 wire \inv_in[2025] ;
 wire \inv_in[2026] ;
 wire \inv_in[2027] ;
 wire \inv_in[2028] ;
 wire \inv_in[2029] ;
 wire \inv_in[202] ;
 wire \inv_in[2030] ;
 wire \inv_in[2031] ;
 wire \inv_in[2032] ;
 wire \inv_in[2033] ;
 wire \inv_in[2034] ;
 wire \inv_in[2035] ;
 wire \inv_in[2036] ;
 wire \inv_in[2037] ;
 wire \inv_in[2038] ;
 wire \inv_in[2039] ;
 wire \inv_in[203] ;
 wire \inv_in[2040] ;
 wire \inv_in[2041] ;
 wire \inv_in[2042] ;
 wire \inv_in[2043] ;
 wire \inv_in[2044] ;
 wire \inv_in[2045] ;
 wire \inv_in[2046] ;
 wire \inv_in[2047] ;
 wire \inv_in[2048] ;
 wire \inv_in[2049] ;
 wire \inv_in[204] ;
 wire \inv_in[2050] ;
 wire \inv_in[2051] ;
 wire \inv_in[2052] ;
 wire \inv_in[2053] ;
 wire \inv_in[2054] ;
 wire \inv_in[2055] ;
 wire \inv_in[2056] ;
 wire \inv_in[2057] ;
 wire \inv_in[2058] ;
 wire \inv_in[2059] ;
 wire \inv_in[205] ;
 wire \inv_in[2060] ;
 wire \inv_in[2061] ;
 wire \inv_in[2062] ;
 wire \inv_in[2063] ;
 wire \inv_in[2064] ;
 wire \inv_in[2065] ;
 wire \inv_in[2066] ;
 wire \inv_in[2067] ;
 wire \inv_in[2068] ;
 wire \inv_in[2069] ;
 wire \inv_in[206] ;
 wire \inv_in[2070] ;
 wire \inv_in[2071] ;
 wire \inv_in[2072] ;
 wire \inv_in[2073] ;
 wire \inv_in[2074] ;
 wire \inv_in[2075] ;
 wire \inv_in[2076] ;
 wire \inv_in[2077] ;
 wire \inv_in[2078] ;
 wire \inv_in[2079] ;
 wire \inv_in[207] ;
 wire \inv_in[2080] ;
 wire \inv_in[2081] ;
 wire \inv_in[2082] ;
 wire \inv_in[2083] ;
 wire \inv_in[2084] ;
 wire \inv_in[2085] ;
 wire \inv_in[2086] ;
 wire \inv_in[2087] ;
 wire \inv_in[2088] ;
 wire \inv_in[2089] ;
 wire \inv_in[208] ;
 wire \inv_in[2090] ;
 wire \inv_in[2091] ;
 wire \inv_in[2092] ;
 wire \inv_in[2093] ;
 wire \inv_in[2094] ;
 wire \inv_in[2095] ;
 wire \inv_in[2096] ;
 wire \inv_in[2097] ;
 wire \inv_in[2098] ;
 wire \inv_in[2099] ;
 wire \inv_in[209] ;
 wire \inv_in[20] ;
 wire \inv_in[2100] ;
 wire \inv_in[2101] ;
 wire \inv_in[2102] ;
 wire \inv_in[2103] ;
 wire \inv_in[2104] ;
 wire \inv_in[2105] ;
 wire \inv_in[2106] ;
 wire \inv_in[2107] ;
 wire \inv_in[2108] ;
 wire \inv_in[2109] ;
 wire \inv_in[210] ;
 wire \inv_in[2110] ;
 wire \inv_in[2111] ;
 wire \inv_in[2112] ;
 wire \inv_in[2113] ;
 wire \inv_in[2114] ;
 wire \inv_in[2115] ;
 wire \inv_in[2116] ;
 wire \inv_in[2117] ;
 wire \inv_in[2118] ;
 wire \inv_in[2119] ;
 wire \inv_in[211] ;
 wire \inv_in[2120] ;
 wire \inv_in[2121] ;
 wire \inv_in[2122] ;
 wire \inv_in[2123] ;
 wire \inv_in[2124] ;
 wire \inv_in[2125] ;
 wire \inv_in[2126] ;
 wire \inv_in[2127] ;
 wire \inv_in[2128] ;
 wire \inv_in[2129] ;
 wire \inv_in[212] ;
 wire \inv_in[2130] ;
 wire \inv_in[2131] ;
 wire \inv_in[2132] ;
 wire \inv_in[2133] ;
 wire \inv_in[2134] ;
 wire \inv_in[2135] ;
 wire \inv_in[2136] ;
 wire \inv_in[2137] ;
 wire \inv_in[2138] ;
 wire \inv_in[2139] ;
 wire \inv_in[213] ;
 wire \inv_in[2140] ;
 wire \inv_in[2141] ;
 wire \inv_in[2142] ;
 wire \inv_in[2143] ;
 wire \inv_in[2144] ;
 wire \inv_in[2145] ;
 wire \inv_in[2146] ;
 wire \inv_in[2147] ;
 wire \inv_in[2148] ;
 wire \inv_in[2149] ;
 wire \inv_in[214] ;
 wire \inv_in[2150] ;
 wire \inv_in[2151] ;
 wire \inv_in[2152] ;
 wire \inv_in[2153] ;
 wire \inv_in[2154] ;
 wire \inv_in[2155] ;
 wire \inv_in[2156] ;
 wire \inv_in[2157] ;
 wire \inv_in[2158] ;
 wire \inv_in[2159] ;
 wire \inv_in[215] ;
 wire \inv_in[2160] ;
 wire \inv_in[2161] ;
 wire \inv_in[2162] ;
 wire \inv_in[2163] ;
 wire \inv_in[2164] ;
 wire \inv_in[2165] ;
 wire \inv_in[2166] ;
 wire \inv_in[2167] ;
 wire \inv_in[2168] ;
 wire \inv_in[2169] ;
 wire \inv_in[216] ;
 wire \inv_in[2170] ;
 wire \inv_in[2171] ;
 wire \inv_in[2172] ;
 wire \inv_in[2173] ;
 wire \inv_in[2174] ;
 wire \inv_in[2175] ;
 wire \inv_in[2176] ;
 wire \inv_in[2177] ;
 wire \inv_in[2178] ;
 wire \inv_in[2179] ;
 wire \inv_in[217] ;
 wire \inv_in[2180] ;
 wire \inv_in[2181] ;
 wire \inv_in[2182] ;
 wire \inv_in[2183] ;
 wire \inv_in[2184] ;
 wire \inv_in[2185] ;
 wire \inv_in[2186] ;
 wire \inv_in[2187] ;
 wire \inv_in[2188] ;
 wire \inv_in[2189] ;
 wire \inv_in[218] ;
 wire \inv_in[2190] ;
 wire \inv_in[2191] ;
 wire \inv_in[2192] ;
 wire \inv_in[2193] ;
 wire \inv_in[2194] ;
 wire \inv_in[2195] ;
 wire \inv_in[2196] ;
 wire \inv_in[2197] ;
 wire \inv_in[2198] ;
 wire \inv_in[2199] ;
 wire \inv_in[219] ;
 wire \inv_in[21] ;
 wire \inv_in[2200] ;
 wire \inv_in[2201] ;
 wire \inv_in[2202] ;
 wire \inv_in[2203] ;
 wire \inv_in[2204] ;
 wire \inv_in[2205] ;
 wire \inv_in[2206] ;
 wire \inv_in[2207] ;
 wire \inv_in[2208] ;
 wire \inv_in[2209] ;
 wire \inv_in[220] ;
 wire \inv_in[2210] ;
 wire \inv_in[2211] ;
 wire \inv_in[2212] ;
 wire \inv_in[2213] ;
 wire \inv_in[2214] ;
 wire \inv_in[2215] ;
 wire \inv_in[2216] ;
 wire \inv_in[2217] ;
 wire \inv_in[2218] ;
 wire \inv_in[2219] ;
 wire \inv_in[221] ;
 wire \inv_in[2220] ;
 wire \inv_in[2221] ;
 wire \inv_in[2222] ;
 wire \inv_in[2223] ;
 wire \inv_in[2224] ;
 wire \inv_in[2225] ;
 wire \inv_in[2226] ;
 wire \inv_in[2227] ;
 wire \inv_in[2228] ;
 wire \inv_in[2229] ;
 wire \inv_in[222] ;
 wire \inv_in[2230] ;
 wire \inv_in[2231] ;
 wire \inv_in[2232] ;
 wire \inv_in[2233] ;
 wire \inv_in[2234] ;
 wire \inv_in[2235] ;
 wire \inv_in[2236] ;
 wire \inv_in[2237] ;
 wire \inv_in[2238] ;
 wire \inv_in[2239] ;
 wire \inv_in[223] ;
 wire \inv_in[2240] ;
 wire \inv_in[2241] ;
 wire \inv_in[2242] ;
 wire \inv_in[2243] ;
 wire \inv_in[2244] ;
 wire \inv_in[2245] ;
 wire \inv_in[2246] ;
 wire \inv_in[2247] ;
 wire \inv_in[2248] ;
 wire \inv_in[2249] ;
 wire \inv_in[224] ;
 wire \inv_in[2250] ;
 wire \inv_in[2251] ;
 wire \inv_in[2252] ;
 wire \inv_in[2253] ;
 wire \inv_in[2254] ;
 wire \inv_in[2255] ;
 wire \inv_in[2256] ;
 wire \inv_in[2257] ;
 wire \inv_in[2258] ;
 wire \inv_in[2259] ;
 wire \inv_in[225] ;
 wire \inv_in[2260] ;
 wire \inv_in[2261] ;
 wire \inv_in[2262] ;
 wire \inv_in[2263] ;
 wire \inv_in[2264] ;
 wire \inv_in[2265] ;
 wire \inv_in[2266] ;
 wire \inv_in[2267] ;
 wire \inv_in[2268] ;
 wire \inv_in[2269] ;
 wire \inv_in[226] ;
 wire \inv_in[2270] ;
 wire \inv_in[2271] ;
 wire \inv_in[2272] ;
 wire \inv_in[2273] ;
 wire \inv_in[2274] ;
 wire \inv_in[2275] ;
 wire \inv_in[2276] ;
 wire \inv_in[2277] ;
 wire \inv_in[2278] ;
 wire \inv_in[2279] ;
 wire \inv_in[227] ;
 wire \inv_in[2280] ;
 wire \inv_in[2281] ;
 wire \inv_in[2282] ;
 wire \inv_in[2283] ;
 wire \inv_in[2284] ;
 wire \inv_in[2285] ;
 wire \inv_in[2286] ;
 wire \inv_in[2287] ;
 wire \inv_in[2288] ;
 wire \inv_in[2289] ;
 wire \inv_in[228] ;
 wire \inv_in[2290] ;
 wire \inv_in[2291] ;
 wire \inv_in[2292] ;
 wire \inv_in[2293] ;
 wire \inv_in[2294] ;
 wire \inv_in[2295] ;
 wire \inv_in[2296] ;
 wire \inv_in[2297] ;
 wire \inv_in[2298] ;
 wire \inv_in[2299] ;
 wire \inv_in[229] ;
 wire \inv_in[22] ;
 wire \inv_in[2300] ;
 wire \inv_in[2301] ;
 wire \inv_in[2302] ;
 wire \inv_in[2303] ;
 wire \inv_in[2304] ;
 wire \inv_in[2305] ;
 wire \inv_in[2306] ;
 wire \inv_in[2307] ;
 wire \inv_in[2308] ;
 wire \inv_in[2309] ;
 wire \inv_in[230] ;
 wire \inv_in[2310] ;
 wire \inv_in[2311] ;
 wire \inv_in[2312] ;
 wire \inv_in[2313] ;
 wire \inv_in[2314] ;
 wire \inv_in[2315] ;
 wire \inv_in[2316] ;
 wire \inv_in[2317] ;
 wire \inv_in[2318] ;
 wire \inv_in[2319] ;
 wire \inv_in[231] ;
 wire \inv_in[2320] ;
 wire \inv_in[2321] ;
 wire \inv_in[2322] ;
 wire \inv_in[2323] ;
 wire \inv_in[2324] ;
 wire \inv_in[2325] ;
 wire \inv_in[2326] ;
 wire \inv_in[2327] ;
 wire \inv_in[2328] ;
 wire \inv_in[2329] ;
 wire \inv_in[232] ;
 wire \inv_in[2330] ;
 wire \inv_in[2331] ;
 wire \inv_in[2332] ;
 wire \inv_in[2333] ;
 wire \inv_in[2334] ;
 wire \inv_in[2335] ;
 wire \inv_in[2336] ;
 wire \inv_in[2337] ;
 wire \inv_in[2338] ;
 wire \inv_in[2339] ;
 wire \inv_in[233] ;
 wire \inv_in[2340] ;
 wire \inv_in[2341] ;
 wire \inv_in[2342] ;
 wire \inv_in[2343] ;
 wire \inv_in[2344] ;
 wire \inv_in[2345] ;
 wire \inv_in[2346] ;
 wire \inv_in[2347] ;
 wire \inv_in[2348] ;
 wire \inv_in[2349] ;
 wire \inv_in[234] ;
 wire \inv_in[2350] ;
 wire \inv_in[2351] ;
 wire \inv_in[2352] ;
 wire \inv_in[2353] ;
 wire \inv_in[2354] ;
 wire \inv_in[2355] ;
 wire \inv_in[2356] ;
 wire \inv_in[2357] ;
 wire \inv_in[2358] ;
 wire \inv_in[2359] ;
 wire \inv_in[235] ;
 wire \inv_in[2360] ;
 wire \inv_in[2361] ;
 wire \inv_in[2362] ;
 wire \inv_in[2363] ;
 wire \inv_in[2364] ;
 wire \inv_in[2365] ;
 wire \inv_in[2366] ;
 wire \inv_in[2367] ;
 wire \inv_in[2368] ;
 wire \inv_in[2369] ;
 wire \inv_in[236] ;
 wire \inv_in[2370] ;
 wire \inv_in[2371] ;
 wire \inv_in[2372] ;
 wire \inv_in[2373] ;
 wire \inv_in[2374] ;
 wire \inv_in[2375] ;
 wire \inv_in[2376] ;
 wire \inv_in[2377] ;
 wire \inv_in[2378] ;
 wire \inv_in[2379] ;
 wire \inv_in[237] ;
 wire \inv_in[2380] ;
 wire \inv_in[2381] ;
 wire \inv_in[2382] ;
 wire \inv_in[2383] ;
 wire \inv_in[2384] ;
 wire \inv_in[2385] ;
 wire \inv_in[2386] ;
 wire \inv_in[2387] ;
 wire \inv_in[2388] ;
 wire \inv_in[2389] ;
 wire \inv_in[238] ;
 wire \inv_in[2390] ;
 wire \inv_in[2391] ;
 wire \inv_in[2392] ;
 wire \inv_in[2393] ;
 wire \inv_in[2394] ;
 wire \inv_in[2395] ;
 wire \inv_in[2396] ;
 wire \inv_in[2397] ;
 wire \inv_in[2398] ;
 wire \inv_in[2399] ;
 wire \inv_in[239] ;
 wire \inv_in[23] ;
 wire \inv_in[2400] ;
 wire \inv_in[2401] ;
 wire \inv_in[2402] ;
 wire \inv_in[2403] ;
 wire \inv_in[2404] ;
 wire \inv_in[2405] ;
 wire \inv_in[2406] ;
 wire \inv_in[2407] ;
 wire \inv_in[2408] ;
 wire \inv_in[2409] ;
 wire \inv_in[240] ;
 wire \inv_in[2410] ;
 wire \inv_in[2411] ;
 wire \inv_in[2412] ;
 wire \inv_in[2413] ;
 wire \inv_in[2414] ;
 wire \inv_in[2415] ;
 wire \inv_in[2416] ;
 wire \inv_in[2417] ;
 wire \inv_in[2418] ;
 wire \inv_in[2419] ;
 wire \inv_in[241] ;
 wire \inv_in[2420] ;
 wire \inv_in[2421] ;
 wire \inv_in[2422] ;
 wire \inv_in[2423] ;
 wire \inv_in[2424] ;
 wire \inv_in[2425] ;
 wire \inv_in[2426] ;
 wire \inv_in[2427] ;
 wire \inv_in[2428] ;
 wire \inv_in[2429] ;
 wire \inv_in[242] ;
 wire \inv_in[2430] ;
 wire \inv_in[2431] ;
 wire \inv_in[2432] ;
 wire \inv_in[2433] ;
 wire \inv_in[2434] ;
 wire \inv_in[2435] ;
 wire \inv_in[2436] ;
 wire \inv_in[2437] ;
 wire \inv_in[2438] ;
 wire \inv_in[2439] ;
 wire \inv_in[243] ;
 wire \inv_in[2440] ;
 wire \inv_in[2441] ;
 wire \inv_in[2442] ;
 wire \inv_in[2443] ;
 wire \inv_in[2444] ;
 wire \inv_in[2445] ;
 wire \inv_in[2446] ;
 wire \inv_in[2447] ;
 wire \inv_in[2448] ;
 wire \inv_in[2449] ;
 wire \inv_in[244] ;
 wire \inv_in[2450] ;
 wire \inv_in[2451] ;
 wire \inv_in[2452] ;
 wire \inv_in[2453] ;
 wire \inv_in[2454] ;
 wire \inv_in[2455] ;
 wire \inv_in[2456] ;
 wire \inv_in[2457] ;
 wire \inv_in[2458] ;
 wire \inv_in[2459] ;
 wire \inv_in[245] ;
 wire \inv_in[2460] ;
 wire \inv_in[2461] ;
 wire \inv_in[2462] ;
 wire \inv_in[2463] ;
 wire \inv_in[2464] ;
 wire \inv_in[2465] ;
 wire \inv_in[2466] ;
 wire \inv_in[2467] ;
 wire \inv_in[2468] ;
 wire \inv_in[2469] ;
 wire \inv_in[246] ;
 wire \inv_in[2470] ;
 wire \inv_in[2471] ;
 wire \inv_in[2472] ;
 wire \inv_in[2473] ;
 wire \inv_in[2474] ;
 wire \inv_in[2475] ;
 wire \inv_in[2476] ;
 wire \inv_in[2477] ;
 wire \inv_in[2478] ;
 wire \inv_in[2479] ;
 wire \inv_in[247] ;
 wire \inv_in[2480] ;
 wire \inv_in[2481] ;
 wire \inv_in[2482] ;
 wire \inv_in[2483] ;
 wire \inv_in[2484] ;
 wire \inv_in[2485] ;
 wire \inv_in[2486] ;
 wire \inv_in[2487] ;
 wire \inv_in[2488] ;
 wire \inv_in[2489] ;
 wire \inv_in[248] ;
 wire \inv_in[2490] ;
 wire \inv_in[2491] ;
 wire \inv_in[2492] ;
 wire \inv_in[2493] ;
 wire \inv_in[2494] ;
 wire \inv_in[2495] ;
 wire \inv_in[2496] ;
 wire \inv_in[2497] ;
 wire \inv_in[2498] ;
 wire \inv_in[2499] ;
 wire \inv_in[249] ;
 wire \inv_in[24] ;
 wire \inv_in[2500] ;
 wire \inv_in[2501] ;
 wire \inv_in[2502] ;
 wire \inv_in[2503] ;
 wire \inv_in[2504] ;
 wire \inv_in[2505] ;
 wire \inv_in[2506] ;
 wire \inv_in[2507] ;
 wire \inv_in[2508] ;
 wire \inv_in[2509] ;
 wire \inv_in[250] ;
 wire \inv_in[2510] ;
 wire \inv_in[2511] ;
 wire \inv_in[2512] ;
 wire \inv_in[2513] ;
 wire \inv_in[2514] ;
 wire \inv_in[2515] ;
 wire \inv_in[2516] ;
 wire \inv_in[2517] ;
 wire \inv_in[2518] ;
 wire \inv_in[2519] ;
 wire \inv_in[251] ;
 wire \inv_in[2520] ;
 wire \inv_in[2521] ;
 wire \inv_in[2522] ;
 wire \inv_in[2523] ;
 wire \inv_in[2524] ;
 wire \inv_in[2525] ;
 wire \inv_in[2526] ;
 wire \inv_in[2527] ;
 wire \inv_in[2528] ;
 wire \inv_in[2529] ;
 wire \inv_in[252] ;
 wire \inv_in[2530] ;
 wire \inv_in[2531] ;
 wire \inv_in[2532] ;
 wire \inv_in[2533] ;
 wire \inv_in[2534] ;
 wire \inv_in[2535] ;
 wire \inv_in[2536] ;
 wire \inv_in[2537] ;
 wire \inv_in[2538] ;
 wire \inv_in[2539] ;
 wire \inv_in[253] ;
 wire \inv_in[2540] ;
 wire \inv_in[2541] ;
 wire \inv_in[2542] ;
 wire \inv_in[2543] ;
 wire \inv_in[2544] ;
 wire \inv_in[2545] ;
 wire \inv_in[2546] ;
 wire \inv_in[2547] ;
 wire \inv_in[2548] ;
 wire \inv_in[2549] ;
 wire \inv_in[254] ;
 wire \inv_in[2550] ;
 wire \inv_in[2551] ;
 wire \inv_in[2552] ;
 wire \inv_in[2553] ;
 wire \inv_in[2554] ;
 wire \inv_in[2555] ;
 wire \inv_in[2556] ;
 wire \inv_in[2557] ;
 wire \inv_in[2558] ;
 wire \inv_in[2559] ;
 wire \inv_in[255] ;
 wire \inv_in[2560] ;
 wire \inv_in[2561] ;
 wire \inv_in[2562] ;
 wire \inv_in[2563] ;
 wire \inv_in[2564] ;
 wire \inv_in[2565] ;
 wire \inv_in[2566] ;
 wire \inv_in[2567] ;
 wire \inv_in[2568] ;
 wire \inv_in[2569] ;
 wire \inv_in[256] ;
 wire \inv_in[2570] ;
 wire \inv_in[2571] ;
 wire \inv_in[2572] ;
 wire \inv_in[2573] ;
 wire \inv_in[2574] ;
 wire \inv_in[2575] ;
 wire \inv_in[2576] ;
 wire \inv_in[2577] ;
 wire \inv_in[2578] ;
 wire \inv_in[2579] ;
 wire \inv_in[257] ;
 wire \inv_in[2580] ;
 wire \inv_in[2581] ;
 wire \inv_in[2582] ;
 wire \inv_in[2583] ;
 wire \inv_in[2584] ;
 wire \inv_in[2585] ;
 wire \inv_in[2586] ;
 wire \inv_in[2587] ;
 wire \inv_in[2588] ;
 wire \inv_in[2589] ;
 wire \inv_in[258] ;
 wire \inv_in[2590] ;
 wire \inv_in[2591] ;
 wire \inv_in[2592] ;
 wire \inv_in[2593] ;
 wire \inv_in[2594] ;
 wire \inv_in[2595] ;
 wire \inv_in[2596] ;
 wire \inv_in[2597] ;
 wire \inv_in[2598] ;
 wire \inv_in[2599] ;
 wire \inv_in[259] ;
 wire \inv_in[25] ;
 wire \inv_in[2600] ;
 wire \inv_in[2601] ;
 wire \inv_in[2602] ;
 wire \inv_in[2603] ;
 wire \inv_in[2604] ;
 wire \inv_in[2605] ;
 wire \inv_in[2606] ;
 wire \inv_in[2607] ;
 wire \inv_in[2608] ;
 wire \inv_in[2609] ;
 wire \inv_in[260] ;
 wire \inv_in[2610] ;
 wire \inv_in[2611] ;
 wire \inv_in[2612] ;
 wire \inv_in[2613] ;
 wire \inv_in[2614] ;
 wire \inv_in[2615] ;
 wire \inv_in[2616] ;
 wire \inv_in[2617] ;
 wire \inv_in[2618] ;
 wire \inv_in[2619] ;
 wire \inv_in[261] ;
 wire \inv_in[2620] ;
 wire \inv_in[2621] ;
 wire \inv_in[2622] ;
 wire \inv_in[2623] ;
 wire \inv_in[2624] ;
 wire \inv_in[2625] ;
 wire \inv_in[2626] ;
 wire \inv_in[2627] ;
 wire \inv_in[2628] ;
 wire \inv_in[2629] ;
 wire \inv_in[262] ;
 wire \inv_in[2630] ;
 wire \inv_in[2631] ;
 wire \inv_in[2632] ;
 wire \inv_in[2633] ;
 wire \inv_in[2634] ;
 wire \inv_in[2635] ;
 wire \inv_in[2636] ;
 wire \inv_in[2637] ;
 wire \inv_in[2638] ;
 wire \inv_in[2639] ;
 wire \inv_in[263] ;
 wire \inv_in[2640] ;
 wire \inv_in[2641] ;
 wire \inv_in[2642] ;
 wire \inv_in[2643] ;
 wire \inv_in[2644] ;
 wire \inv_in[2645] ;
 wire \inv_in[2646] ;
 wire \inv_in[2647] ;
 wire \inv_in[2648] ;
 wire \inv_in[2649] ;
 wire \inv_in[264] ;
 wire \inv_in[2650] ;
 wire \inv_in[2651] ;
 wire \inv_in[2652] ;
 wire \inv_in[2653] ;
 wire \inv_in[2654] ;
 wire \inv_in[2655] ;
 wire \inv_in[2656] ;
 wire \inv_in[2657] ;
 wire \inv_in[2658] ;
 wire \inv_in[2659] ;
 wire \inv_in[265] ;
 wire \inv_in[2660] ;
 wire \inv_in[2661] ;
 wire \inv_in[2662] ;
 wire \inv_in[2663] ;
 wire \inv_in[2664] ;
 wire \inv_in[2665] ;
 wire \inv_in[2666] ;
 wire \inv_in[2667] ;
 wire \inv_in[2668] ;
 wire \inv_in[2669] ;
 wire \inv_in[266] ;
 wire \inv_in[2670] ;
 wire \inv_in[2671] ;
 wire \inv_in[2672] ;
 wire \inv_in[2673] ;
 wire \inv_in[2674] ;
 wire \inv_in[2675] ;
 wire \inv_in[2676] ;
 wire \inv_in[2677] ;
 wire \inv_in[2678] ;
 wire \inv_in[2679] ;
 wire \inv_in[267] ;
 wire \inv_in[2680] ;
 wire \inv_in[2681] ;
 wire \inv_in[2682] ;
 wire \inv_in[2683] ;
 wire \inv_in[2684] ;
 wire \inv_in[2685] ;
 wire \inv_in[2686] ;
 wire \inv_in[2687] ;
 wire \inv_in[2688] ;
 wire \inv_in[2689] ;
 wire \inv_in[268] ;
 wire \inv_in[2690] ;
 wire \inv_in[2691] ;
 wire \inv_in[2692] ;
 wire \inv_in[2693] ;
 wire \inv_in[2694] ;
 wire \inv_in[2695] ;
 wire \inv_in[2696] ;
 wire \inv_in[2697] ;
 wire \inv_in[2698] ;
 wire \inv_in[2699] ;
 wire \inv_in[269] ;
 wire \inv_in[26] ;
 wire \inv_in[2700] ;
 wire \inv_in[2701] ;
 wire \inv_in[2702] ;
 wire \inv_in[2703] ;
 wire \inv_in[2704] ;
 wire \inv_in[2705] ;
 wire \inv_in[2706] ;
 wire \inv_in[2707] ;
 wire \inv_in[2708] ;
 wire \inv_in[2709] ;
 wire \inv_in[270] ;
 wire \inv_in[2710] ;
 wire \inv_in[2711] ;
 wire \inv_in[2712] ;
 wire \inv_in[2713] ;
 wire \inv_in[2714] ;
 wire \inv_in[2715] ;
 wire \inv_in[2716] ;
 wire \inv_in[2717] ;
 wire \inv_in[2718] ;
 wire \inv_in[2719] ;
 wire \inv_in[271] ;
 wire \inv_in[2720] ;
 wire \inv_in[2721] ;
 wire \inv_in[2722] ;
 wire \inv_in[2723] ;
 wire \inv_in[2724] ;
 wire \inv_in[2725] ;
 wire \inv_in[2726] ;
 wire \inv_in[2727] ;
 wire \inv_in[2728] ;
 wire \inv_in[2729] ;
 wire \inv_in[272] ;
 wire \inv_in[2730] ;
 wire \inv_in[2731] ;
 wire \inv_in[2732] ;
 wire \inv_in[2733] ;
 wire \inv_in[2734] ;
 wire \inv_in[2735] ;
 wire \inv_in[2736] ;
 wire \inv_in[2737] ;
 wire \inv_in[2738] ;
 wire \inv_in[2739] ;
 wire \inv_in[273] ;
 wire \inv_in[2740] ;
 wire \inv_in[2741] ;
 wire \inv_in[2742] ;
 wire \inv_in[2743] ;
 wire \inv_in[2744] ;
 wire \inv_in[2745] ;
 wire \inv_in[2746] ;
 wire \inv_in[2747] ;
 wire \inv_in[2748] ;
 wire \inv_in[2749] ;
 wire \inv_in[274] ;
 wire \inv_in[2750] ;
 wire \inv_in[2751] ;
 wire \inv_in[2752] ;
 wire \inv_in[2753] ;
 wire \inv_in[2754] ;
 wire \inv_in[2755] ;
 wire \inv_in[2756] ;
 wire \inv_in[2757] ;
 wire \inv_in[2758] ;
 wire \inv_in[2759] ;
 wire \inv_in[275] ;
 wire \inv_in[2760] ;
 wire \inv_in[2761] ;
 wire \inv_in[2762] ;
 wire \inv_in[2763] ;
 wire \inv_in[2764] ;
 wire \inv_in[2765] ;
 wire \inv_in[2766] ;
 wire \inv_in[2767] ;
 wire \inv_in[2768] ;
 wire \inv_in[2769] ;
 wire \inv_in[276] ;
 wire \inv_in[2770] ;
 wire \inv_in[2771] ;
 wire \inv_in[2772] ;
 wire \inv_in[2773] ;
 wire \inv_in[2774] ;
 wire \inv_in[2775] ;
 wire \inv_in[2776] ;
 wire \inv_in[2777] ;
 wire \inv_in[2778] ;
 wire \inv_in[2779] ;
 wire \inv_in[277] ;
 wire \inv_in[2780] ;
 wire \inv_in[2781] ;
 wire \inv_in[2782] ;
 wire \inv_in[2783] ;
 wire \inv_in[2784] ;
 wire \inv_in[2785] ;
 wire \inv_in[2786] ;
 wire \inv_in[2787] ;
 wire \inv_in[2788] ;
 wire \inv_in[2789] ;
 wire \inv_in[278] ;
 wire \inv_in[2790] ;
 wire \inv_in[2791] ;
 wire \inv_in[2792] ;
 wire \inv_in[2793] ;
 wire \inv_in[2794] ;
 wire \inv_in[2795] ;
 wire \inv_in[2796] ;
 wire \inv_in[2797] ;
 wire \inv_in[2798] ;
 wire \inv_in[2799] ;
 wire \inv_in[279] ;
 wire \inv_in[27] ;
 wire \inv_in[2800] ;
 wire \inv_in[2801] ;
 wire \inv_in[2802] ;
 wire \inv_in[2803] ;
 wire \inv_in[2804] ;
 wire \inv_in[2805] ;
 wire \inv_in[2806] ;
 wire \inv_in[2807] ;
 wire \inv_in[2808] ;
 wire \inv_in[2809] ;
 wire \inv_in[280] ;
 wire \inv_in[2810] ;
 wire \inv_in[2811] ;
 wire \inv_in[2812] ;
 wire \inv_in[2813] ;
 wire \inv_in[2814] ;
 wire \inv_in[2815] ;
 wire \inv_in[2816] ;
 wire \inv_in[2817] ;
 wire \inv_in[2818] ;
 wire \inv_in[2819] ;
 wire \inv_in[281] ;
 wire \inv_in[2820] ;
 wire \inv_in[2821] ;
 wire \inv_in[2822] ;
 wire \inv_in[2823] ;
 wire \inv_in[2824] ;
 wire \inv_in[2825] ;
 wire \inv_in[2826] ;
 wire \inv_in[2827] ;
 wire \inv_in[2828] ;
 wire \inv_in[2829] ;
 wire \inv_in[282] ;
 wire \inv_in[2830] ;
 wire \inv_in[2831] ;
 wire \inv_in[2832] ;
 wire \inv_in[2833] ;
 wire \inv_in[2834] ;
 wire \inv_in[2835] ;
 wire \inv_in[2836] ;
 wire \inv_in[2837] ;
 wire \inv_in[2838] ;
 wire \inv_in[2839] ;
 wire \inv_in[283] ;
 wire \inv_in[2840] ;
 wire \inv_in[2841] ;
 wire \inv_in[2842] ;
 wire \inv_in[2843] ;
 wire \inv_in[2844] ;
 wire \inv_in[2845] ;
 wire \inv_in[2846] ;
 wire \inv_in[2847] ;
 wire \inv_in[2848] ;
 wire \inv_in[2849] ;
 wire \inv_in[284] ;
 wire \inv_in[2850] ;
 wire \inv_in[2851] ;
 wire \inv_in[2852] ;
 wire \inv_in[2853] ;
 wire \inv_in[2854] ;
 wire \inv_in[2855] ;
 wire \inv_in[2856] ;
 wire \inv_in[2857] ;
 wire \inv_in[2858] ;
 wire \inv_in[2859] ;
 wire \inv_in[285] ;
 wire \inv_in[2860] ;
 wire \inv_in[2861] ;
 wire \inv_in[2862] ;
 wire \inv_in[2863] ;
 wire \inv_in[2864] ;
 wire \inv_in[2865] ;
 wire \inv_in[2866] ;
 wire \inv_in[2867] ;
 wire \inv_in[2868] ;
 wire \inv_in[2869] ;
 wire \inv_in[286] ;
 wire \inv_in[2870] ;
 wire \inv_in[2871] ;
 wire \inv_in[2872] ;
 wire \inv_in[2873] ;
 wire \inv_in[2874] ;
 wire \inv_in[2875] ;
 wire \inv_in[2876] ;
 wire \inv_in[2877] ;
 wire \inv_in[2878] ;
 wire \inv_in[2879] ;
 wire \inv_in[287] ;
 wire \inv_in[2880] ;
 wire \inv_in[2881] ;
 wire \inv_in[2882] ;
 wire \inv_in[2883] ;
 wire \inv_in[2884] ;
 wire \inv_in[2885] ;
 wire \inv_in[2886] ;
 wire \inv_in[2887] ;
 wire \inv_in[2888] ;
 wire \inv_in[2889] ;
 wire \inv_in[288] ;
 wire \inv_in[2890] ;
 wire \inv_in[2891] ;
 wire \inv_in[2892] ;
 wire \inv_in[2893] ;
 wire \inv_in[2894] ;
 wire \inv_in[2895] ;
 wire \inv_in[2896] ;
 wire \inv_in[2897] ;
 wire \inv_in[2898] ;
 wire \inv_in[2899] ;
 wire \inv_in[289] ;
 wire \inv_in[28] ;
 wire \inv_in[2900] ;
 wire \inv_in[2901] ;
 wire \inv_in[2902] ;
 wire \inv_in[2903] ;
 wire \inv_in[2904] ;
 wire \inv_in[2905] ;
 wire \inv_in[2906] ;
 wire \inv_in[2907] ;
 wire \inv_in[2908] ;
 wire \inv_in[2909] ;
 wire \inv_in[290] ;
 wire \inv_in[2910] ;
 wire \inv_in[2911] ;
 wire \inv_in[2912] ;
 wire \inv_in[2913] ;
 wire \inv_in[2914] ;
 wire \inv_in[2915] ;
 wire \inv_in[2916] ;
 wire \inv_in[2917] ;
 wire \inv_in[2918] ;
 wire \inv_in[2919] ;
 wire \inv_in[291] ;
 wire \inv_in[2920] ;
 wire \inv_in[2921] ;
 wire \inv_in[2922] ;
 wire \inv_in[2923] ;
 wire \inv_in[2924] ;
 wire \inv_in[2925] ;
 wire \inv_in[2926] ;
 wire \inv_in[2927] ;
 wire \inv_in[2928] ;
 wire \inv_in[2929] ;
 wire \inv_in[292] ;
 wire \inv_in[2930] ;
 wire \inv_in[2931] ;
 wire \inv_in[2932] ;
 wire \inv_in[2933] ;
 wire \inv_in[2934] ;
 wire \inv_in[2935] ;
 wire \inv_in[2936] ;
 wire \inv_in[2937] ;
 wire \inv_in[2938] ;
 wire \inv_in[2939] ;
 wire \inv_in[293] ;
 wire \inv_in[2940] ;
 wire \inv_in[2941] ;
 wire \inv_in[2942] ;
 wire \inv_in[2943] ;
 wire \inv_in[2944] ;
 wire \inv_in[2945] ;
 wire \inv_in[2946] ;
 wire \inv_in[2947] ;
 wire \inv_in[2948] ;
 wire \inv_in[2949] ;
 wire \inv_in[294] ;
 wire \inv_in[2950] ;
 wire \inv_in[2951] ;
 wire \inv_in[2952] ;
 wire \inv_in[2953] ;
 wire \inv_in[2954] ;
 wire \inv_in[2955] ;
 wire \inv_in[2956] ;
 wire \inv_in[2957] ;
 wire \inv_in[2958] ;
 wire \inv_in[2959] ;
 wire \inv_in[295] ;
 wire \inv_in[2960] ;
 wire \inv_in[2961] ;
 wire \inv_in[2962] ;
 wire \inv_in[2963] ;
 wire \inv_in[2964] ;
 wire \inv_in[2965] ;
 wire \inv_in[2966] ;
 wire \inv_in[2967] ;
 wire \inv_in[2968] ;
 wire \inv_in[2969] ;
 wire \inv_in[296] ;
 wire \inv_in[2970] ;
 wire \inv_in[2971] ;
 wire \inv_in[2972] ;
 wire \inv_in[2973] ;
 wire \inv_in[2974] ;
 wire \inv_in[2975] ;
 wire \inv_in[2976] ;
 wire \inv_in[2977] ;
 wire \inv_in[2978] ;
 wire \inv_in[2979] ;
 wire \inv_in[297] ;
 wire \inv_in[2980] ;
 wire \inv_in[2981] ;
 wire \inv_in[2982] ;
 wire \inv_in[2983] ;
 wire \inv_in[2984] ;
 wire \inv_in[2985] ;
 wire \inv_in[2986] ;
 wire \inv_in[2987] ;
 wire \inv_in[2988] ;
 wire \inv_in[2989] ;
 wire \inv_in[298] ;
 wire \inv_in[2990] ;
 wire \inv_in[2991] ;
 wire \inv_in[2992] ;
 wire \inv_in[2993] ;
 wire \inv_in[2994] ;
 wire \inv_in[2995] ;
 wire \inv_in[2996] ;
 wire \inv_in[2997] ;
 wire \inv_in[2998] ;
 wire \inv_in[2999] ;
 wire \inv_in[299] ;
 wire \inv_in[29] ;
 wire \inv_in[2] ;
 wire \inv_in[3000] ;
 wire \inv_in[3001] ;
 wire \inv_in[3002] ;
 wire \inv_in[3003] ;
 wire \inv_in[3004] ;
 wire \inv_in[3005] ;
 wire \inv_in[3006] ;
 wire \inv_in[3007] ;
 wire \inv_in[3008] ;
 wire \inv_in[3009] ;
 wire \inv_in[300] ;
 wire \inv_in[3010] ;
 wire \inv_in[3011] ;
 wire \inv_in[3012] ;
 wire \inv_in[3013] ;
 wire \inv_in[3014] ;
 wire \inv_in[3015] ;
 wire \inv_in[3016] ;
 wire \inv_in[3017] ;
 wire \inv_in[3018] ;
 wire \inv_in[3019] ;
 wire \inv_in[301] ;
 wire \inv_in[3020] ;
 wire \inv_in[3021] ;
 wire \inv_in[3022] ;
 wire \inv_in[3023] ;
 wire \inv_in[3024] ;
 wire \inv_in[3025] ;
 wire \inv_in[3026] ;
 wire \inv_in[3027] ;
 wire \inv_in[3028] ;
 wire \inv_in[3029] ;
 wire \inv_in[302] ;
 wire \inv_in[3030] ;
 wire \inv_in[3031] ;
 wire \inv_in[3032] ;
 wire \inv_in[3033] ;
 wire \inv_in[3034] ;
 wire \inv_in[3035] ;
 wire \inv_in[3036] ;
 wire \inv_in[3037] ;
 wire \inv_in[3038] ;
 wire \inv_in[3039] ;
 wire \inv_in[303] ;
 wire \inv_in[3040] ;
 wire \inv_in[3041] ;
 wire \inv_in[3042] ;
 wire \inv_in[3043] ;
 wire \inv_in[3044] ;
 wire \inv_in[3045] ;
 wire \inv_in[3046] ;
 wire \inv_in[3047] ;
 wire \inv_in[3048] ;
 wire \inv_in[3049] ;
 wire \inv_in[304] ;
 wire \inv_in[3050] ;
 wire \inv_in[3051] ;
 wire \inv_in[3052] ;
 wire \inv_in[3053] ;
 wire \inv_in[3054] ;
 wire \inv_in[3055] ;
 wire \inv_in[3056] ;
 wire \inv_in[3057] ;
 wire \inv_in[3058] ;
 wire \inv_in[3059] ;
 wire \inv_in[305] ;
 wire \inv_in[3060] ;
 wire \inv_in[3061] ;
 wire \inv_in[3062] ;
 wire \inv_in[3063] ;
 wire \inv_in[3064] ;
 wire \inv_in[3065] ;
 wire \inv_in[3066] ;
 wire \inv_in[3067] ;
 wire \inv_in[3068] ;
 wire \inv_in[3069] ;
 wire \inv_in[306] ;
 wire \inv_in[3070] ;
 wire \inv_in[3071] ;
 wire \inv_in[3072] ;
 wire \inv_in[3073] ;
 wire \inv_in[3074] ;
 wire \inv_in[3075] ;
 wire \inv_in[3076] ;
 wire \inv_in[3077] ;
 wire \inv_in[3078] ;
 wire \inv_in[3079] ;
 wire \inv_in[307] ;
 wire \inv_in[3080] ;
 wire \inv_in[3081] ;
 wire \inv_in[3082] ;
 wire \inv_in[3083] ;
 wire \inv_in[3084] ;
 wire \inv_in[3085] ;
 wire \inv_in[3086] ;
 wire \inv_in[3087] ;
 wire \inv_in[3088] ;
 wire \inv_in[3089] ;
 wire \inv_in[308] ;
 wire \inv_in[3090] ;
 wire \inv_in[3091] ;
 wire \inv_in[3092] ;
 wire \inv_in[3093] ;
 wire \inv_in[3094] ;
 wire \inv_in[3095] ;
 wire \inv_in[3096] ;
 wire \inv_in[3097] ;
 wire \inv_in[3098] ;
 wire \inv_in[3099] ;
 wire \inv_in[309] ;
 wire \inv_in[30] ;
 wire \inv_in[3100] ;
 wire \inv_in[3101] ;
 wire \inv_in[3102] ;
 wire \inv_in[3103] ;
 wire \inv_in[3104] ;
 wire \inv_in[3105] ;
 wire \inv_in[3106] ;
 wire \inv_in[3107] ;
 wire \inv_in[3108] ;
 wire \inv_in[3109] ;
 wire \inv_in[310] ;
 wire \inv_in[3110] ;
 wire \inv_in[3111] ;
 wire \inv_in[3112] ;
 wire \inv_in[3113] ;
 wire \inv_in[3114] ;
 wire \inv_in[3115] ;
 wire \inv_in[3116] ;
 wire \inv_in[3117] ;
 wire \inv_in[3118] ;
 wire \inv_in[3119] ;
 wire \inv_in[311] ;
 wire \inv_in[3120] ;
 wire \inv_in[3121] ;
 wire \inv_in[3122] ;
 wire \inv_in[3123] ;
 wire \inv_in[3124] ;
 wire \inv_in[3125] ;
 wire \inv_in[3126] ;
 wire \inv_in[3127] ;
 wire \inv_in[3128] ;
 wire \inv_in[3129] ;
 wire \inv_in[312] ;
 wire \inv_in[3130] ;
 wire \inv_in[3131] ;
 wire \inv_in[3132] ;
 wire \inv_in[3133] ;
 wire \inv_in[3134] ;
 wire \inv_in[3135] ;
 wire \inv_in[3136] ;
 wire \inv_in[3137] ;
 wire \inv_in[3138] ;
 wire \inv_in[3139] ;
 wire \inv_in[313] ;
 wire \inv_in[3140] ;
 wire \inv_in[3141] ;
 wire \inv_in[3142] ;
 wire \inv_in[3143] ;
 wire \inv_in[3144] ;
 wire \inv_in[3145] ;
 wire \inv_in[3146] ;
 wire \inv_in[3147] ;
 wire \inv_in[3148] ;
 wire \inv_in[3149] ;
 wire \inv_in[314] ;
 wire \inv_in[3150] ;
 wire \inv_in[3151] ;
 wire \inv_in[3152] ;
 wire \inv_in[3153] ;
 wire \inv_in[3154] ;
 wire \inv_in[3155] ;
 wire \inv_in[3156] ;
 wire \inv_in[3157] ;
 wire \inv_in[3158] ;
 wire \inv_in[3159] ;
 wire \inv_in[315] ;
 wire \inv_in[3160] ;
 wire \inv_in[3161] ;
 wire \inv_in[3162] ;
 wire \inv_in[3163] ;
 wire \inv_in[3164] ;
 wire \inv_in[3165] ;
 wire \inv_in[3166] ;
 wire \inv_in[3167] ;
 wire \inv_in[3168] ;
 wire \inv_in[3169] ;
 wire \inv_in[316] ;
 wire \inv_in[3170] ;
 wire \inv_in[3171] ;
 wire \inv_in[3172] ;
 wire \inv_in[3173] ;
 wire \inv_in[3174] ;
 wire \inv_in[3175] ;
 wire \inv_in[3176] ;
 wire \inv_in[3177] ;
 wire \inv_in[3178] ;
 wire \inv_in[3179] ;
 wire \inv_in[317] ;
 wire \inv_in[3180] ;
 wire \inv_in[3181] ;
 wire \inv_in[3182] ;
 wire \inv_in[3183] ;
 wire \inv_in[3184] ;
 wire \inv_in[3185] ;
 wire \inv_in[3186] ;
 wire \inv_in[3187] ;
 wire \inv_in[3188] ;
 wire \inv_in[3189] ;
 wire \inv_in[318] ;
 wire \inv_in[3190] ;
 wire \inv_in[3191] ;
 wire \inv_in[3192] ;
 wire \inv_in[3193] ;
 wire \inv_in[3194] ;
 wire \inv_in[3195] ;
 wire \inv_in[3196] ;
 wire \inv_in[3197] ;
 wire \inv_in[3198] ;
 wire \inv_in[3199] ;
 wire \inv_in[319] ;
 wire \inv_in[31] ;
 wire \inv_in[3200] ;
 wire \inv_in[3201] ;
 wire \inv_in[3202] ;
 wire \inv_in[3203] ;
 wire \inv_in[3204] ;
 wire \inv_in[3205] ;
 wire \inv_in[3206] ;
 wire \inv_in[3207] ;
 wire \inv_in[3208] ;
 wire \inv_in[3209] ;
 wire \inv_in[320] ;
 wire \inv_in[3210] ;
 wire \inv_in[3211] ;
 wire \inv_in[3212] ;
 wire \inv_in[3213] ;
 wire \inv_in[3214] ;
 wire \inv_in[3215] ;
 wire \inv_in[3216] ;
 wire \inv_in[3217] ;
 wire \inv_in[3218] ;
 wire \inv_in[3219] ;
 wire \inv_in[321] ;
 wire \inv_in[3220] ;
 wire \inv_in[3221] ;
 wire \inv_in[3222] ;
 wire \inv_in[3223] ;
 wire \inv_in[3224] ;
 wire \inv_in[3225] ;
 wire \inv_in[3226] ;
 wire \inv_in[3227] ;
 wire \inv_in[3228] ;
 wire \inv_in[3229] ;
 wire \inv_in[322] ;
 wire \inv_in[3230] ;
 wire \inv_in[3231] ;
 wire \inv_in[3232] ;
 wire \inv_in[3233] ;
 wire \inv_in[3234] ;
 wire \inv_in[3235] ;
 wire \inv_in[3236] ;
 wire \inv_in[3237] ;
 wire \inv_in[3238] ;
 wire \inv_in[3239] ;
 wire \inv_in[323] ;
 wire \inv_in[3240] ;
 wire \inv_in[3241] ;
 wire \inv_in[3242] ;
 wire \inv_in[3243] ;
 wire \inv_in[3244] ;
 wire \inv_in[3245] ;
 wire \inv_in[3246] ;
 wire \inv_in[3247] ;
 wire \inv_in[3248] ;
 wire \inv_in[3249] ;
 wire \inv_in[324] ;
 wire \inv_in[3250] ;
 wire \inv_in[3251] ;
 wire \inv_in[3252] ;
 wire \inv_in[3253] ;
 wire \inv_in[3254] ;
 wire \inv_in[3255] ;
 wire \inv_in[3256] ;
 wire \inv_in[3257] ;
 wire \inv_in[3258] ;
 wire \inv_in[3259] ;
 wire \inv_in[325] ;
 wire \inv_in[3260] ;
 wire \inv_in[3261] ;
 wire \inv_in[3262] ;
 wire \inv_in[3263] ;
 wire \inv_in[3264] ;
 wire \inv_in[3265] ;
 wire \inv_in[3266] ;
 wire \inv_in[3267] ;
 wire \inv_in[3268] ;
 wire \inv_in[3269] ;
 wire \inv_in[326] ;
 wire \inv_in[3270] ;
 wire \inv_in[3271] ;
 wire \inv_in[3272] ;
 wire \inv_in[3273] ;
 wire \inv_in[3274] ;
 wire \inv_in[3275] ;
 wire \inv_in[3276] ;
 wire \inv_in[3277] ;
 wire \inv_in[3278] ;
 wire \inv_in[3279] ;
 wire \inv_in[327] ;
 wire \inv_in[3280] ;
 wire \inv_in[3281] ;
 wire \inv_in[3282] ;
 wire \inv_in[3283] ;
 wire \inv_in[3284] ;
 wire \inv_in[3285] ;
 wire \inv_in[3286] ;
 wire \inv_in[3287] ;
 wire \inv_in[3288] ;
 wire \inv_in[3289] ;
 wire \inv_in[328] ;
 wire \inv_in[3290] ;
 wire \inv_in[3291] ;
 wire \inv_in[3292] ;
 wire \inv_in[3293] ;
 wire \inv_in[3294] ;
 wire \inv_in[3295] ;
 wire \inv_in[3296] ;
 wire \inv_in[3297] ;
 wire \inv_in[3298] ;
 wire \inv_in[3299] ;
 wire \inv_in[329] ;
 wire \inv_in[32] ;
 wire \inv_in[3300] ;
 wire \inv_in[3301] ;
 wire \inv_in[3302] ;
 wire \inv_in[3303] ;
 wire \inv_in[3304] ;
 wire \inv_in[3305] ;
 wire \inv_in[3306] ;
 wire \inv_in[3307] ;
 wire \inv_in[3308] ;
 wire \inv_in[3309] ;
 wire \inv_in[330] ;
 wire \inv_in[3310] ;
 wire \inv_in[3311] ;
 wire \inv_in[3312] ;
 wire \inv_in[3313] ;
 wire \inv_in[3314] ;
 wire \inv_in[3315] ;
 wire \inv_in[3316] ;
 wire \inv_in[3317] ;
 wire \inv_in[3318] ;
 wire \inv_in[3319] ;
 wire \inv_in[331] ;
 wire \inv_in[3320] ;
 wire \inv_in[3321] ;
 wire \inv_in[3322] ;
 wire \inv_in[3323] ;
 wire \inv_in[3324] ;
 wire \inv_in[3325] ;
 wire \inv_in[3326] ;
 wire \inv_in[3327] ;
 wire \inv_in[3328] ;
 wire \inv_in[3329] ;
 wire \inv_in[332] ;
 wire \inv_in[3330] ;
 wire \inv_in[3331] ;
 wire \inv_in[3332] ;
 wire \inv_in[3333] ;
 wire \inv_in[3334] ;
 wire \inv_in[3335] ;
 wire \inv_in[3336] ;
 wire \inv_in[3337] ;
 wire \inv_in[3338] ;
 wire \inv_in[3339] ;
 wire \inv_in[333] ;
 wire \inv_in[3340] ;
 wire \inv_in[3341] ;
 wire \inv_in[3342] ;
 wire \inv_in[3343] ;
 wire \inv_in[3344] ;
 wire \inv_in[3345] ;
 wire \inv_in[3346] ;
 wire \inv_in[3347] ;
 wire \inv_in[3348] ;
 wire \inv_in[3349] ;
 wire \inv_in[334] ;
 wire \inv_in[3350] ;
 wire \inv_in[3351] ;
 wire \inv_in[3352] ;
 wire \inv_in[3353] ;
 wire \inv_in[3354] ;
 wire \inv_in[3355] ;
 wire \inv_in[3356] ;
 wire \inv_in[3357] ;
 wire \inv_in[3358] ;
 wire \inv_in[3359] ;
 wire \inv_in[335] ;
 wire \inv_in[3360] ;
 wire \inv_in[3361] ;
 wire \inv_in[3362] ;
 wire \inv_in[3363] ;
 wire \inv_in[3364] ;
 wire \inv_in[3365] ;
 wire \inv_in[3366] ;
 wire \inv_in[3367] ;
 wire \inv_in[3368] ;
 wire \inv_in[3369] ;
 wire \inv_in[336] ;
 wire \inv_in[3370] ;
 wire \inv_in[3371] ;
 wire \inv_in[3372] ;
 wire \inv_in[3373] ;
 wire \inv_in[3374] ;
 wire \inv_in[3375] ;
 wire \inv_in[3376] ;
 wire \inv_in[3377] ;
 wire \inv_in[3378] ;
 wire \inv_in[3379] ;
 wire \inv_in[337] ;
 wire \inv_in[3380] ;
 wire \inv_in[3381] ;
 wire \inv_in[3382] ;
 wire \inv_in[3383] ;
 wire \inv_in[3384] ;
 wire \inv_in[3385] ;
 wire \inv_in[3386] ;
 wire \inv_in[3387] ;
 wire \inv_in[3388] ;
 wire \inv_in[3389] ;
 wire \inv_in[338] ;
 wire \inv_in[3390] ;
 wire \inv_in[3391] ;
 wire \inv_in[3392] ;
 wire \inv_in[3393] ;
 wire \inv_in[3394] ;
 wire \inv_in[3395] ;
 wire \inv_in[3396] ;
 wire \inv_in[3397] ;
 wire \inv_in[3398] ;
 wire \inv_in[3399] ;
 wire \inv_in[339] ;
 wire \inv_in[33] ;
 wire \inv_in[3400] ;
 wire \inv_in[3401] ;
 wire \inv_in[3402] ;
 wire \inv_in[3403] ;
 wire \inv_in[3404] ;
 wire \inv_in[3405] ;
 wire \inv_in[3406] ;
 wire \inv_in[3407] ;
 wire \inv_in[3408] ;
 wire \inv_in[3409] ;
 wire \inv_in[340] ;
 wire \inv_in[3410] ;
 wire \inv_in[3411] ;
 wire \inv_in[3412] ;
 wire \inv_in[3413] ;
 wire \inv_in[3414] ;
 wire \inv_in[3415] ;
 wire \inv_in[3416] ;
 wire \inv_in[3417] ;
 wire \inv_in[3418] ;
 wire \inv_in[3419] ;
 wire \inv_in[341] ;
 wire \inv_in[3420] ;
 wire \inv_in[3421] ;
 wire \inv_in[3422] ;
 wire \inv_in[3423] ;
 wire \inv_in[3424] ;
 wire \inv_in[3425] ;
 wire \inv_in[3426] ;
 wire \inv_in[3427] ;
 wire \inv_in[3428] ;
 wire \inv_in[3429] ;
 wire \inv_in[342] ;
 wire \inv_in[3430] ;
 wire \inv_in[3431] ;
 wire \inv_in[3432] ;
 wire \inv_in[3433] ;
 wire \inv_in[3434] ;
 wire \inv_in[3435] ;
 wire \inv_in[3436] ;
 wire \inv_in[3437] ;
 wire \inv_in[3438] ;
 wire \inv_in[3439] ;
 wire \inv_in[343] ;
 wire \inv_in[3440] ;
 wire \inv_in[3441] ;
 wire \inv_in[3442] ;
 wire \inv_in[3443] ;
 wire \inv_in[3444] ;
 wire \inv_in[3445] ;
 wire \inv_in[3446] ;
 wire \inv_in[3447] ;
 wire \inv_in[3448] ;
 wire \inv_in[3449] ;
 wire \inv_in[344] ;
 wire \inv_in[3450] ;
 wire \inv_in[3451] ;
 wire \inv_in[3452] ;
 wire \inv_in[3453] ;
 wire \inv_in[3454] ;
 wire \inv_in[3455] ;
 wire \inv_in[3456] ;
 wire \inv_in[3457] ;
 wire \inv_in[3458] ;
 wire \inv_in[3459] ;
 wire \inv_in[345] ;
 wire \inv_in[3460] ;
 wire \inv_in[3461] ;
 wire \inv_in[3462] ;
 wire \inv_in[3463] ;
 wire \inv_in[3464] ;
 wire \inv_in[3465] ;
 wire \inv_in[3466] ;
 wire \inv_in[3467] ;
 wire \inv_in[3468] ;
 wire \inv_in[3469] ;
 wire \inv_in[346] ;
 wire \inv_in[3470] ;
 wire \inv_in[3471] ;
 wire \inv_in[3472] ;
 wire \inv_in[3473] ;
 wire \inv_in[3474] ;
 wire \inv_in[3475] ;
 wire \inv_in[3476] ;
 wire \inv_in[3477] ;
 wire \inv_in[3478] ;
 wire \inv_in[3479] ;
 wire \inv_in[347] ;
 wire \inv_in[3480] ;
 wire \inv_in[3481] ;
 wire \inv_in[3482] ;
 wire \inv_in[3483] ;
 wire \inv_in[3484] ;
 wire \inv_in[3485] ;
 wire \inv_in[3486] ;
 wire \inv_in[3487] ;
 wire \inv_in[3488] ;
 wire \inv_in[3489] ;
 wire \inv_in[348] ;
 wire \inv_in[3490] ;
 wire \inv_in[3491] ;
 wire \inv_in[3492] ;
 wire \inv_in[3493] ;
 wire \inv_in[3494] ;
 wire \inv_in[3495] ;
 wire \inv_in[3496] ;
 wire \inv_in[3497] ;
 wire \inv_in[3498] ;
 wire \inv_in[3499] ;
 wire \inv_in[349] ;
 wire \inv_in[34] ;
 wire \inv_in[3500] ;
 wire \inv_in[3501] ;
 wire \inv_in[3502] ;
 wire \inv_in[3503] ;
 wire \inv_in[3504] ;
 wire \inv_in[3505] ;
 wire \inv_in[3506] ;
 wire \inv_in[3507] ;
 wire \inv_in[3508] ;
 wire \inv_in[3509] ;
 wire \inv_in[350] ;
 wire \inv_in[3510] ;
 wire \inv_in[3511] ;
 wire \inv_in[3512] ;
 wire \inv_in[3513] ;
 wire \inv_in[3514] ;
 wire \inv_in[3515] ;
 wire \inv_in[3516] ;
 wire \inv_in[3517] ;
 wire \inv_in[3518] ;
 wire \inv_in[3519] ;
 wire \inv_in[351] ;
 wire \inv_in[3520] ;
 wire \inv_in[3521] ;
 wire \inv_in[3522] ;
 wire \inv_in[3523] ;
 wire \inv_in[3524] ;
 wire \inv_in[3525] ;
 wire \inv_in[3526] ;
 wire \inv_in[3527] ;
 wire \inv_in[3528] ;
 wire \inv_in[3529] ;
 wire \inv_in[352] ;
 wire \inv_in[3530] ;
 wire \inv_in[3531] ;
 wire \inv_in[3532] ;
 wire \inv_in[3533] ;
 wire \inv_in[3534] ;
 wire \inv_in[3535] ;
 wire \inv_in[3536] ;
 wire \inv_in[3537] ;
 wire \inv_in[3538] ;
 wire \inv_in[3539] ;
 wire \inv_in[353] ;
 wire \inv_in[3540] ;
 wire \inv_in[3541] ;
 wire \inv_in[3542] ;
 wire \inv_in[3543] ;
 wire \inv_in[3544] ;
 wire \inv_in[3545] ;
 wire \inv_in[3546] ;
 wire \inv_in[3547] ;
 wire \inv_in[3548] ;
 wire \inv_in[3549] ;
 wire \inv_in[354] ;
 wire \inv_in[3550] ;
 wire \inv_in[3551] ;
 wire \inv_in[3552] ;
 wire \inv_in[3553] ;
 wire \inv_in[3554] ;
 wire \inv_in[3555] ;
 wire \inv_in[3556] ;
 wire \inv_in[3557] ;
 wire \inv_in[3558] ;
 wire \inv_in[3559] ;
 wire \inv_in[355] ;
 wire \inv_in[3560] ;
 wire \inv_in[3561] ;
 wire \inv_in[3562] ;
 wire \inv_in[3563] ;
 wire \inv_in[3564] ;
 wire \inv_in[3565] ;
 wire \inv_in[3566] ;
 wire \inv_in[3567] ;
 wire \inv_in[3568] ;
 wire \inv_in[3569] ;
 wire \inv_in[356] ;
 wire \inv_in[3570] ;
 wire \inv_in[3571] ;
 wire \inv_in[3572] ;
 wire \inv_in[3573] ;
 wire \inv_in[3574] ;
 wire \inv_in[3575] ;
 wire \inv_in[3576] ;
 wire \inv_in[3577] ;
 wire \inv_in[3578] ;
 wire \inv_in[3579] ;
 wire \inv_in[357] ;
 wire \inv_in[3580] ;
 wire \inv_in[3581] ;
 wire \inv_in[3582] ;
 wire \inv_in[3583] ;
 wire \inv_in[3584] ;
 wire \inv_in[3585] ;
 wire \inv_in[3586] ;
 wire \inv_in[3587] ;
 wire \inv_in[3588] ;
 wire \inv_in[3589] ;
 wire \inv_in[358] ;
 wire \inv_in[3590] ;
 wire \inv_in[3591] ;
 wire \inv_in[3592] ;
 wire \inv_in[3593] ;
 wire \inv_in[3594] ;
 wire \inv_in[3595] ;
 wire \inv_in[3596] ;
 wire \inv_in[3597] ;
 wire \inv_in[3598] ;
 wire \inv_in[3599] ;
 wire \inv_in[359] ;
 wire \inv_in[35] ;
 wire \inv_in[3600] ;
 wire \inv_in[3601] ;
 wire \inv_in[3602] ;
 wire \inv_in[3603] ;
 wire \inv_in[3604] ;
 wire \inv_in[3605] ;
 wire \inv_in[3606] ;
 wire \inv_in[3607] ;
 wire \inv_in[3608] ;
 wire \inv_in[3609] ;
 wire \inv_in[360] ;
 wire \inv_in[3610] ;
 wire \inv_in[3611] ;
 wire \inv_in[3612] ;
 wire \inv_in[3613] ;
 wire \inv_in[3614] ;
 wire \inv_in[3615] ;
 wire \inv_in[3616] ;
 wire \inv_in[3617] ;
 wire \inv_in[3618] ;
 wire \inv_in[3619] ;
 wire \inv_in[361] ;
 wire \inv_in[3620] ;
 wire \inv_in[3621] ;
 wire \inv_in[3622] ;
 wire \inv_in[3623] ;
 wire \inv_in[3624] ;
 wire \inv_in[3625] ;
 wire \inv_in[3626] ;
 wire \inv_in[3627] ;
 wire \inv_in[3628] ;
 wire \inv_in[3629] ;
 wire \inv_in[362] ;
 wire \inv_in[3630] ;
 wire \inv_in[3631] ;
 wire \inv_in[3632] ;
 wire \inv_in[3633] ;
 wire \inv_in[3634] ;
 wire \inv_in[3635] ;
 wire \inv_in[3636] ;
 wire \inv_in[3637] ;
 wire \inv_in[3638] ;
 wire \inv_in[3639] ;
 wire \inv_in[363] ;
 wire \inv_in[3640] ;
 wire \inv_in[3641] ;
 wire \inv_in[3642] ;
 wire \inv_in[3643] ;
 wire \inv_in[3644] ;
 wire \inv_in[3645] ;
 wire \inv_in[3646] ;
 wire \inv_in[3647] ;
 wire \inv_in[3648] ;
 wire \inv_in[3649] ;
 wire \inv_in[364] ;
 wire \inv_in[3650] ;
 wire \inv_in[3651] ;
 wire \inv_in[3652] ;
 wire \inv_in[3653] ;
 wire \inv_in[3654] ;
 wire \inv_in[3655] ;
 wire \inv_in[3656] ;
 wire \inv_in[3657] ;
 wire \inv_in[3658] ;
 wire \inv_in[3659] ;
 wire \inv_in[365] ;
 wire \inv_in[3660] ;
 wire \inv_in[3661] ;
 wire \inv_in[3662] ;
 wire \inv_in[3663] ;
 wire \inv_in[3664] ;
 wire \inv_in[3665] ;
 wire \inv_in[3666] ;
 wire \inv_in[3667] ;
 wire \inv_in[3668] ;
 wire \inv_in[3669] ;
 wire \inv_in[366] ;
 wire \inv_in[3670] ;
 wire \inv_in[3671] ;
 wire \inv_in[3672] ;
 wire \inv_in[3673] ;
 wire \inv_in[3674] ;
 wire \inv_in[3675] ;
 wire \inv_in[3676] ;
 wire \inv_in[3677] ;
 wire \inv_in[3678] ;
 wire \inv_in[3679] ;
 wire \inv_in[367] ;
 wire \inv_in[3680] ;
 wire \inv_in[3681] ;
 wire \inv_in[3682] ;
 wire \inv_in[3683] ;
 wire \inv_in[3684] ;
 wire \inv_in[3685] ;
 wire \inv_in[3686] ;
 wire \inv_in[3687] ;
 wire \inv_in[3688] ;
 wire \inv_in[3689] ;
 wire \inv_in[368] ;
 wire \inv_in[3690] ;
 wire \inv_in[3691] ;
 wire \inv_in[3692] ;
 wire \inv_in[3693] ;
 wire \inv_in[3694] ;
 wire \inv_in[3695] ;
 wire \inv_in[3696] ;
 wire \inv_in[3697] ;
 wire \inv_in[3698] ;
 wire \inv_in[3699] ;
 wire \inv_in[369] ;
 wire \inv_in[36] ;
 wire \inv_in[3700] ;
 wire \inv_in[3701] ;
 wire \inv_in[3702] ;
 wire \inv_in[3703] ;
 wire \inv_in[3704] ;
 wire \inv_in[3705] ;
 wire \inv_in[3706] ;
 wire \inv_in[3707] ;
 wire \inv_in[3708] ;
 wire \inv_in[3709] ;
 wire \inv_in[370] ;
 wire \inv_in[3710] ;
 wire \inv_in[3711] ;
 wire \inv_in[3712] ;
 wire \inv_in[3713] ;
 wire \inv_in[3714] ;
 wire \inv_in[3715] ;
 wire \inv_in[3716] ;
 wire \inv_in[3717] ;
 wire \inv_in[3718] ;
 wire \inv_in[3719] ;
 wire \inv_in[371] ;
 wire \inv_in[3720] ;
 wire \inv_in[3721] ;
 wire \inv_in[3722] ;
 wire \inv_in[3723] ;
 wire \inv_in[3724] ;
 wire \inv_in[3725] ;
 wire \inv_in[3726] ;
 wire \inv_in[3727] ;
 wire \inv_in[3728] ;
 wire \inv_in[3729] ;
 wire \inv_in[372] ;
 wire \inv_in[3730] ;
 wire \inv_in[3731] ;
 wire \inv_in[3732] ;
 wire \inv_in[3733] ;
 wire \inv_in[3734] ;
 wire \inv_in[3735] ;
 wire \inv_in[3736] ;
 wire \inv_in[3737] ;
 wire \inv_in[3738] ;
 wire \inv_in[3739] ;
 wire \inv_in[373] ;
 wire \inv_in[3740] ;
 wire \inv_in[3741] ;
 wire \inv_in[3742] ;
 wire \inv_in[3743] ;
 wire \inv_in[3744] ;
 wire \inv_in[3745] ;
 wire \inv_in[3746] ;
 wire \inv_in[3747] ;
 wire \inv_in[3748] ;
 wire \inv_in[3749] ;
 wire \inv_in[374] ;
 wire \inv_in[3750] ;
 wire \inv_in[3751] ;
 wire \inv_in[3752] ;
 wire \inv_in[3753] ;
 wire \inv_in[3754] ;
 wire \inv_in[3755] ;
 wire \inv_in[3756] ;
 wire \inv_in[3757] ;
 wire \inv_in[3758] ;
 wire \inv_in[3759] ;
 wire \inv_in[375] ;
 wire \inv_in[3760] ;
 wire \inv_in[3761] ;
 wire \inv_in[3762] ;
 wire \inv_in[3763] ;
 wire \inv_in[3764] ;
 wire \inv_in[3765] ;
 wire \inv_in[3766] ;
 wire \inv_in[3767] ;
 wire \inv_in[3768] ;
 wire \inv_in[3769] ;
 wire \inv_in[376] ;
 wire \inv_in[3770] ;
 wire \inv_in[3771] ;
 wire \inv_in[3772] ;
 wire \inv_in[3773] ;
 wire \inv_in[3774] ;
 wire \inv_in[3775] ;
 wire \inv_in[3776] ;
 wire \inv_in[3777] ;
 wire \inv_in[3778] ;
 wire \inv_in[3779] ;
 wire \inv_in[377] ;
 wire \inv_in[3780] ;
 wire \inv_in[3781] ;
 wire \inv_in[3782] ;
 wire \inv_in[3783] ;
 wire \inv_in[3784] ;
 wire \inv_in[3785] ;
 wire \inv_in[3786] ;
 wire \inv_in[3787] ;
 wire \inv_in[3788] ;
 wire \inv_in[3789] ;
 wire \inv_in[378] ;
 wire \inv_in[3790] ;
 wire \inv_in[3791] ;
 wire \inv_in[3792] ;
 wire \inv_in[3793] ;
 wire \inv_in[3794] ;
 wire \inv_in[3795] ;
 wire \inv_in[3796] ;
 wire \inv_in[3797] ;
 wire \inv_in[3798] ;
 wire \inv_in[3799] ;
 wire \inv_in[379] ;
 wire \inv_in[37] ;
 wire \inv_in[3800] ;
 wire \inv_in[3801] ;
 wire \inv_in[3802] ;
 wire \inv_in[3803] ;
 wire \inv_in[3804] ;
 wire \inv_in[3805] ;
 wire \inv_in[3806] ;
 wire \inv_in[3807] ;
 wire \inv_in[3808] ;
 wire \inv_in[3809] ;
 wire \inv_in[380] ;
 wire \inv_in[3810] ;
 wire \inv_in[3811] ;
 wire \inv_in[3812] ;
 wire \inv_in[3813] ;
 wire \inv_in[3814] ;
 wire \inv_in[3815] ;
 wire \inv_in[3816] ;
 wire \inv_in[3817] ;
 wire \inv_in[3818] ;
 wire \inv_in[3819] ;
 wire \inv_in[381] ;
 wire \inv_in[3820] ;
 wire \inv_in[3821] ;
 wire \inv_in[3822] ;
 wire \inv_in[3823] ;
 wire \inv_in[3824] ;
 wire \inv_in[3825] ;
 wire \inv_in[3826] ;
 wire \inv_in[3827] ;
 wire \inv_in[3828] ;
 wire \inv_in[3829] ;
 wire \inv_in[382] ;
 wire \inv_in[3830] ;
 wire \inv_in[3831] ;
 wire \inv_in[3832] ;
 wire \inv_in[3833] ;
 wire \inv_in[3834] ;
 wire \inv_in[3835] ;
 wire \inv_in[3836] ;
 wire \inv_in[3837] ;
 wire \inv_in[3838] ;
 wire \inv_in[3839] ;
 wire \inv_in[383] ;
 wire \inv_in[3840] ;
 wire \inv_in[3841] ;
 wire \inv_in[3842] ;
 wire \inv_in[3843] ;
 wire \inv_in[3844] ;
 wire \inv_in[3845] ;
 wire \inv_in[3846] ;
 wire \inv_in[3847] ;
 wire \inv_in[3848] ;
 wire \inv_in[3849] ;
 wire \inv_in[384] ;
 wire \inv_in[3850] ;
 wire \inv_in[3851] ;
 wire \inv_in[3852] ;
 wire \inv_in[385] ;
 wire \inv_in[386] ;
 wire \inv_in[387] ;
 wire \inv_in[388] ;
 wire \inv_in[389] ;
 wire \inv_in[38] ;
 wire \inv_in[390] ;
 wire \inv_in[391] ;
 wire \inv_in[392] ;
 wire \inv_in[393] ;
 wire \inv_in[394] ;
 wire \inv_in[395] ;
 wire \inv_in[396] ;
 wire \inv_in[397] ;
 wire \inv_in[398] ;
 wire \inv_in[399] ;
 wire \inv_in[39] ;
 wire \inv_in[3] ;
 wire \inv_in[400] ;
 wire \inv_in[401] ;
 wire \inv_in[402] ;
 wire \inv_in[403] ;
 wire \inv_in[404] ;
 wire \inv_in[405] ;
 wire \inv_in[406] ;
 wire \inv_in[407] ;
 wire \inv_in[408] ;
 wire \inv_in[409] ;
 wire \inv_in[40] ;
 wire \inv_in[410] ;
 wire \inv_in[411] ;
 wire \inv_in[412] ;
 wire \inv_in[413] ;
 wire \inv_in[414] ;
 wire \inv_in[415] ;
 wire \inv_in[416] ;
 wire \inv_in[417] ;
 wire \inv_in[418] ;
 wire \inv_in[419] ;
 wire \inv_in[41] ;
 wire \inv_in[420] ;
 wire \inv_in[421] ;
 wire \inv_in[422] ;
 wire \inv_in[423] ;
 wire \inv_in[424] ;
 wire \inv_in[425] ;
 wire \inv_in[426] ;
 wire \inv_in[427] ;
 wire \inv_in[428] ;
 wire \inv_in[429] ;
 wire \inv_in[42] ;
 wire \inv_in[430] ;
 wire \inv_in[431] ;
 wire \inv_in[432] ;
 wire \inv_in[433] ;
 wire \inv_in[434] ;
 wire \inv_in[435] ;
 wire \inv_in[436] ;
 wire \inv_in[437] ;
 wire \inv_in[438] ;
 wire \inv_in[439] ;
 wire \inv_in[43] ;
 wire \inv_in[440] ;
 wire \inv_in[441] ;
 wire \inv_in[442] ;
 wire \inv_in[443] ;
 wire \inv_in[444] ;
 wire \inv_in[445] ;
 wire \inv_in[446] ;
 wire \inv_in[447] ;
 wire \inv_in[448] ;
 wire \inv_in[449] ;
 wire \inv_in[44] ;
 wire \inv_in[450] ;
 wire \inv_in[451] ;
 wire \inv_in[452] ;
 wire \inv_in[453] ;
 wire \inv_in[454] ;
 wire \inv_in[455] ;
 wire \inv_in[456] ;
 wire \inv_in[457] ;
 wire \inv_in[458] ;
 wire \inv_in[459] ;
 wire \inv_in[45] ;
 wire \inv_in[460] ;
 wire \inv_in[461] ;
 wire \inv_in[462] ;
 wire \inv_in[463] ;
 wire \inv_in[464] ;
 wire \inv_in[465] ;
 wire \inv_in[466] ;
 wire \inv_in[467] ;
 wire \inv_in[468] ;
 wire \inv_in[469] ;
 wire \inv_in[46] ;
 wire \inv_in[470] ;
 wire \inv_in[471] ;
 wire \inv_in[472] ;
 wire \inv_in[473] ;
 wire \inv_in[474] ;
 wire \inv_in[475] ;
 wire \inv_in[476] ;
 wire \inv_in[477] ;
 wire \inv_in[478] ;
 wire \inv_in[479] ;
 wire \inv_in[47] ;
 wire \inv_in[480] ;
 wire \inv_in[481] ;
 wire \inv_in[482] ;
 wire \inv_in[483] ;
 wire \inv_in[484] ;
 wire \inv_in[485] ;
 wire \inv_in[486] ;
 wire \inv_in[487] ;
 wire \inv_in[488] ;
 wire \inv_in[489] ;
 wire \inv_in[48] ;
 wire \inv_in[490] ;
 wire \inv_in[491] ;
 wire \inv_in[492] ;
 wire \inv_in[493] ;
 wire \inv_in[494] ;
 wire \inv_in[495] ;
 wire \inv_in[496] ;
 wire \inv_in[497] ;
 wire \inv_in[498] ;
 wire \inv_in[499] ;
 wire \inv_in[49] ;
 wire \inv_in[4] ;
 wire \inv_in[500] ;
 wire \inv_in[501] ;
 wire \inv_in[502] ;
 wire \inv_in[503] ;
 wire \inv_in[504] ;
 wire \inv_in[505] ;
 wire \inv_in[506] ;
 wire \inv_in[507] ;
 wire \inv_in[508] ;
 wire \inv_in[509] ;
 wire \inv_in[50] ;
 wire \inv_in[510] ;
 wire \inv_in[511] ;
 wire \inv_in[512] ;
 wire \inv_in[513] ;
 wire \inv_in[514] ;
 wire \inv_in[515] ;
 wire \inv_in[516] ;
 wire \inv_in[517] ;
 wire \inv_in[518] ;
 wire \inv_in[519] ;
 wire \inv_in[51] ;
 wire \inv_in[520] ;
 wire \inv_in[521] ;
 wire \inv_in[522] ;
 wire \inv_in[523] ;
 wire \inv_in[524] ;
 wire \inv_in[525] ;
 wire \inv_in[526] ;
 wire \inv_in[527] ;
 wire \inv_in[528] ;
 wire \inv_in[529] ;
 wire \inv_in[52] ;
 wire \inv_in[530] ;
 wire \inv_in[531] ;
 wire \inv_in[532] ;
 wire \inv_in[533] ;
 wire \inv_in[534] ;
 wire \inv_in[535] ;
 wire \inv_in[536] ;
 wire \inv_in[537] ;
 wire \inv_in[538] ;
 wire \inv_in[539] ;
 wire \inv_in[53] ;
 wire \inv_in[540] ;
 wire \inv_in[541] ;
 wire \inv_in[542] ;
 wire \inv_in[543] ;
 wire \inv_in[544] ;
 wire \inv_in[545] ;
 wire \inv_in[546] ;
 wire \inv_in[547] ;
 wire \inv_in[548] ;
 wire \inv_in[549] ;
 wire \inv_in[54] ;
 wire \inv_in[550] ;
 wire \inv_in[551] ;
 wire \inv_in[552] ;
 wire \inv_in[553] ;
 wire \inv_in[554] ;
 wire \inv_in[555] ;
 wire \inv_in[556] ;
 wire \inv_in[557] ;
 wire \inv_in[558] ;
 wire \inv_in[559] ;
 wire \inv_in[55] ;
 wire \inv_in[560] ;
 wire \inv_in[561] ;
 wire \inv_in[562] ;
 wire \inv_in[563] ;
 wire \inv_in[564] ;
 wire \inv_in[565] ;
 wire \inv_in[566] ;
 wire \inv_in[567] ;
 wire \inv_in[568] ;
 wire \inv_in[569] ;
 wire \inv_in[56] ;
 wire \inv_in[570] ;
 wire \inv_in[571] ;
 wire \inv_in[572] ;
 wire \inv_in[573] ;
 wire \inv_in[574] ;
 wire \inv_in[575] ;
 wire \inv_in[576] ;
 wire \inv_in[577] ;
 wire \inv_in[578] ;
 wire \inv_in[579] ;
 wire \inv_in[57] ;
 wire \inv_in[580] ;
 wire \inv_in[581] ;
 wire \inv_in[582] ;
 wire \inv_in[583] ;
 wire \inv_in[584] ;
 wire \inv_in[585] ;
 wire \inv_in[586] ;
 wire \inv_in[587] ;
 wire \inv_in[588] ;
 wire \inv_in[589] ;
 wire \inv_in[58] ;
 wire \inv_in[590] ;
 wire \inv_in[591] ;
 wire \inv_in[592] ;
 wire \inv_in[593] ;
 wire \inv_in[594] ;
 wire \inv_in[595] ;
 wire \inv_in[596] ;
 wire \inv_in[597] ;
 wire \inv_in[598] ;
 wire \inv_in[599] ;
 wire \inv_in[59] ;
 wire \inv_in[5] ;
 wire \inv_in[600] ;
 wire \inv_in[601] ;
 wire \inv_in[602] ;
 wire \inv_in[603] ;
 wire \inv_in[604] ;
 wire \inv_in[605] ;
 wire \inv_in[606] ;
 wire \inv_in[607] ;
 wire \inv_in[608] ;
 wire \inv_in[609] ;
 wire \inv_in[60] ;
 wire \inv_in[610] ;
 wire \inv_in[611] ;
 wire \inv_in[612] ;
 wire \inv_in[613] ;
 wire \inv_in[614] ;
 wire \inv_in[615] ;
 wire \inv_in[616] ;
 wire \inv_in[617] ;
 wire \inv_in[618] ;
 wire \inv_in[619] ;
 wire \inv_in[61] ;
 wire \inv_in[620] ;
 wire \inv_in[621] ;
 wire \inv_in[622] ;
 wire \inv_in[623] ;
 wire \inv_in[624] ;
 wire \inv_in[625] ;
 wire \inv_in[626] ;
 wire \inv_in[627] ;
 wire \inv_in[628] ;
 wire \inv_in[629] ;
 wire \inv_in[62] ;
 wire \inv_in[630] ;
 wire \inv_in[631] ;
 wire \inv_in[632] ;
 wire \inv_in[633] ;
 wire \inv_in[634] ;
 wire \inv_in[635] ;
 wire \inv_in[636] ;
 wire \inv_in[637] ;
 wire \inv_in[638] ;
 wire \inv_in[639] ;
 wire \inv_in[63] ;
 wire \inv_in[640] ;
 wire \inv_in[641] ;
 wire \inv_in[642] ;
 wire \inv_in[643] ;
 wire \inv_in[644] ;
 wire \inv_in[645] ;
 wire \inv_in[646] ;
 wire \inv_in[647] ;
 wire \inv_in[648] ;
 wire \inv_in[649] ;
 wire \inv_in[64] ;
 wire \inv_in[650] ;
 wire \inv_in[651] ;
 wire \inv_in[652] ;
 wire \inv_in[653] ;
 wire \inv_in[654] ;
 wire \inv_in[655] ;
 wire \inv_in[656] ;
 wire \inv_in[657] ;
 wire \inv_in[658] ;
 wire \inv_in[659] ;
 wire \inv_in[65] ;
 wire \inv_in[660] ;
 wire \inv_in[661] ;
 wire \inv_in[662] ;
 wire \inv_in[663] ;
 wire \inv_in[664] ;
 wire \inv_in[665] ;
 wire \inv_in[666] ;
 wire \inv_in[667] ;
 wire \inv_in[668] ;
 wire \inv_in[669] ;
 wire \inv_in[66] ;
 wire \inv_in[670] ;
 wire \inv_in[671] ;
 wire \inv_in[672] ;
 wire \inv_in[673] ;
 wire \inv_in[674] ;
 wire \inv_in[675] ;
 wire \inv_in[676] ;
 wire \inv_in[677] ;
 wire \inv_in[678] ;
 wire \inv_in[679] ;
 wire \inv_in[67] ;
 wire \inv_in[680] ;
 wire \inv_in[681] ;
 wire \inv_in[682] ;
 wire \inv_in[683] ;
 wire \inv_in[684] ;
 wire \inv_in[685] ;
 wire \inv_in[686] ;
 wire \inv_in[687] ;
 wire \inv_in[688] ;
 wire \inv_in[689] ;
 wire \inv_in[68] ;
 wire \inv_in[690] ;
 wire \inv_in[691] ;
 wire \inv_in[692] ;
 wire \inv_in[693] ;
 wire \inv_in[694] ;
 wire \inv_in[695] ;
 wire \inv_in[696] ;
 wire \inv_in[697] ;
 wire \inv_in[698] ;
 wire \inv_in[699] ;
 wire \inv_in[69] ;
 wire \inv_in[6] ;
 wire \inv_in[700] ;
 wire \inv_in[701] ;
 wire \inv_in[702] ;
 wire \inv_in[703] ;
 wire \inv_in[704] ;
 wire \inv_in[705] ;
 wire \inv_in[706] ;
 wire \inv_in[707] ;
 wire \inv_in[708] ;
 wire \inv_in[709] ;
 wire \inv_in[70] ;
 wire \inv_in[710] ;
 wire \inv_in[711] ;
 wire \inv_in[712] ;
 wire \inv_in[713] ;
 wire \inv_in[714] ;
 wire \inv_in[715] ;
 wire \inv_in[716] ;
 wire \inv_in[717] ;
 wire \inv_in[718] ;
 wire \inv_in[719] ;
 wire \inv_in[71] ;
 wire \inv_in[720] ;
 wire \inv_in[721] ;
 wire \inv_in[722] ;
 wire \inv_in[723] ;
 wire \inv_in[724] ;
 wire \inv_in[725] ;
 wire \inv_in[726] ;
 wire \inv_in[727] ;
 wire \inv_in[728] ;
 wire \inv_in[729] ;
 wire \inv_in[72] ;
 wire \inv_in[730] ;
 wire \inv_in[731] ;
 wire \inv_in[732] ;
 wire \inv_in[733] ;
 wire \inv_in[734] ;
 wire \inv_in[735] ;
 wire \inv_in[736] ;
 wire \inv_in[737] ;
 wire \inv_in[738] ;
 wire \inv_in[739] ;
 wire \inv_in[73] ;
 wire \inv_in[740] ;
 wire \inv_in[741] ;
 wire \inv_in[742] ;
 wire \inv_in[743] ;
 wire \inv_in[744] ;
 wire \inv_in[745] ;
 wire \inv_in[746] ;
 wire \inv_in[747] ;
 wire \inv_in[748] ;
 wire \inv_in[749] ;
 wire \inv_in[74] ;
 wire \inv_in[750] ;
 wire \inv_in[751] ;
 wire \inv_in[752] ;
 wire \inv_in[753] ;
 wire \inv_in[754] ;
 wire \inv_in[755] ;
 wire \inv_in[756] ;
 wire \inv_in[757] ;
 wire \inv_in[758] ;
 wire \inv_in[759] ;
 wire \inv_in[75] ;
 wire \inv_in[760] ;
 wire \inv_in[761] ;
 wire \inv_in[762] ;
 wire \inv_in[763] ;
 wire \inv_in[764] ;
 wire \inv_in[765] ;
 wire \inv_in[766] ;
 wire \inv_in[767] ;
 wire \inv_in[768] ;
 wire \inv_in[769] ;
 wire \inv_in[76] ;
 wire \inv_in[770] ;
 wire \inv_in[771] ;
 wire \inv_in[772] ;
 wire \inv_in[773] ;
 wire \inv_in[774] ;
 wire \inv_in[775] ;
 wire \inv_in[776] ;
 wire \inv_in[777] ;
 wire \inv_in[778] ;
 wire \inv_in[779] ;
 wire \inv_in[77] ;
 wire \inv_in[780] ;
 wire \inv_in[781] ;
 wire \inv_in[782] ;
 wire \inv_in[783] ;
 wire \inv_in[784] ;
 wire \inv_in[785] ;
 wire \inv_in[786] ;
 wire \inv_in[787] ;
 wire \inv_in[788] ;
 wire \inv_in[789] ;
 wire \inv_in[78] ;
 wire \inv_in[790] ;
 wire \inv_in[791] ;
 wire \inv_in[792] ;
 wire \inv_in[793] ;
 wire \inv_in[794] ;
 wire \inv_in[795] ;
 wire \inv_in[796] ;
 wire \inv_in[797] ;
 wire \inv_in[798] ;
 wire \inv_in[799] ;
 wire \inv_in[79] ;
 wire \inv_in[7] ;
 wire \inv_in[800] ;
 wire \inv_in[801] ;
 wire \inv_in[802] ;
 wire \inv_in[803] ;
 wire \inv_in[804] ;
 wire \inv_in[805] ;
 wire \inv_in[806] ;
 wire \inv_in[807] ;
 wire \inv_in[808] ;
 wire \inv_in[809] ;
 wire \inv_in[80] ;
 wire \inv_in[810] ;
 wire \inv_in[811] ;
 wire \inv_in[812] ;
 wire \inv_in[813] ;
 wire \inv_in[814] ;
 wire \inv_in[815] ;
 wire \inv_in[816] ;
 wire \inv_in[817] ;
 wire \inv_in[818] ;
 wire \inv_in[819] ;
 wire \inv_in[81] ;
 wire \inv_in[820] ;
 wire \inv_in[821] ;
 wire \inv_in[822] ;
 wire \inv_in[823] ;
 wire \inv_in[824] ;
 wire \inv_in[825] ;
 wire \inv_in[826] ;
 wire \inv_in[827] ;
 wire \inv_in[828] ;
 wire \inv_in[829] ;
 wire \inv_in[82] ;
 wire \inv_in[830] ;
 wire \inv_in[831] ;
 wire \inv_in[832] ;
 wire \inv_in[833] ;
 wire \inv_in[834] ;
 wire \inv_in[835] ;
 wire \inv_in[836] ;
 wire \inv_in[837] ;
 wire \inv_in[838] ;
 wire \inv_in[839] ;
 wire \inv_in[83] ;
 wire \inv_in[840] ;
 wire \inv_in[841] ;
 wire \inv_in[842] ;
 wire \inv_in[843] ;
 wire \inv_in[844] ;
 wire \inv_in[845] ;
 wire \inv_in[846] ;
 wire \inv_in[847] ;
 wire \inv_in[848] ;
 wire \inv_in[849] ;
 wire \inv_in[84] ;
 wire \inv_in[850] ;
 wire \inv_in[851] ;
 wire \inv_in[852] ;
 wire \inv_in[853] ;
 wire \inv_in[854] ;
 wire \inv_in[855] ;
 wire \inv_in[856] ;
 wire \inv_in[857] ;
 wire \inv_in[858] ;
 wire \inv_in[859] ;
 wire \inv_in[85] ;
 wire \inv_in[860] ;
 wire \inv_in[861] ;
 wire \inv_in[862] ;
 wire \inv_in[863] ;
 wire \inv_in[864] ;
 wire \inv_in[865] ;
 wire \inv_in[866] ;
 wire \inv_in[867] ;
 wire \inv_in[868] ;
 wire \inv_in[869] ;
 wire \inv_in[86] ;
 wire \inv_in[870] ;
 wire \inv_in[871] ;
 wire \inv_in[872] ;
 wire \inv_in[873] ;
 wire \inv_in[874] ;
 wire \inv_in[875] ;
 wire \inv_in[876] ;
 wire \inv_in[877] ;
 wire \inv_in[878] ;
 wire \inv_in[879] ;
 wire \inv_in[87] ;
 wire \inv_in[880] ;
 wire \inv_in[881] ;
 wire \inv_in[882] ;
 wire \inv_in[883] ;
 wire \inv_in[884] ;
 wire \inv_in[885] ;
 wire \inv_in[886] ;
 wire \inv_in[887] ;
 wire \inv_in[888] ;
 wire \inv_in[889] ;
 wire \inv_in[88] ;
 wire \inv_in[890] ;
 wire \inv_in[891] ;
 wire \inv_in[892] ;
 wire \inv_in[893] ;
 wire \inv_in[894] ;
 wire \inv_in[895] ;
 wire \inv_in[896] ;
 wire \inv_in[897] ;
 wire \inv_in[898] ;
 wire \inv_in[899] ;
 wire \inv_in[89] ;
 wire \inv_in[8] ;
 wire \inv_in[900] ;
 wire \inv_in[901] ;
 wire \inv_in[902] ;
 wire \inv_in[903] ;
 wire \inv_in[904] ;
 wire \inv_in[905] ;
 wire \inv_in[906] ;
 wire \inv_in[907] ;
 wire \inv_in[908] ;
 wire \inv_in[909] ;
 wire \inv_in[90] ;
 wire \inv_in[910] ;
 wire \inv_in[911] ;
 wire \inv_in[912] ;
 wire \inv_in[913] ;
 wire \inv_in[914] ;
 wire \inv_in[915] ;
 wire \inv_in[916] ;
 wire \inv_in[917] ;
 wire \inv_in[918] ;
 wire \inv_in[919] ;
 wire \inv_in[91] ;
 wire \inv_in[920] ;
 wire \inv_in[921] ;
 wire \inv_in[922] ;
 wire \inv_in[923] ;
 wire \inv_in[924] ;
 wire \inv_in[925] ;
 wire \inv_in[926] ;
 wire \inv_in[927] ;
 wire \inv_in[928] ;
 wire \inv_in[929] ;
 wire \inv_in[92] ;
 wire \inv_in[930] ;
 wire \inv_in[931] ;
 wire \inv_in[932] ;
 wire \inv_in[933] ;
 wire \inv_in[934] ;
 wire \inv_in[935] ;
 wire \inv_in[936] ;
 wire \inv_in[937] ;
 wire \inv_in[938] ;
 wire \inv_in[939] ;
 wire \inv_in[93] ;
 wire \inv_in[940] ;
 wire \inv_in[941] ;
 wire \inv_in[942] ;
 wire \inv_in[943] ;
 wire \inv_in[944] ;
 wire \inv_in[945] ;
 wire \inv_in[946] ;
 wire \inv_in[947] ;
 wire \inv_in[948] ;
 wire \inv_in[949] ;
 wire \inv_in[94] ;
 wire \inv_in[950] ;
 wire \inv_in[951] ;
 wire \inv_in[952] ;
 wire \inv_in[953] ;
 wire \inv_in[954] ;
 wire \inv_in[955] ;
 wire \inv_in[956] ;
 wire \inv_in[957] ;
 wire \inv_in[958] ;
 wire \inv_in[959] ;
 wire \inv_in[95] ;
 wire \inv_in[960] ;
 wire \inv_in[961] ;
 wire \inv_in[962] ;
 wire \inv_in[963] ;
 wire \inv_in[964] ;
 wire \inv_in[965] ;
 wire \inv_in[966] ;
 wire \inv_in[967] ;
 wire \inv_in[968] ;
 wire \inv_in[969] ;
 wire \inv_in[96] ;
 wire \inv_in[970] ;
 wire \inv_in[971] ;
 wire \inv_in[972] ;
 wire \inv_in[973] ;
 wire \inv_in[974] ;
 wire \inv_in[975] ;
 wire \inv_in[976] ;
 wire \inv_in[977] ;
 wire \inv_in[978] ;
 wire \inv_in[979] ;
 wire \inv_in[97] ;
 wire \inv_in[980] ;
 wire \inv_in[981] ;
 wire \inv_in[982] ;
 wire \inv_in[983] ;
 wire \inv_in[984] ;
 wire \inv_in[985] ;
 wire \inv_in[986] ;
 wire \inv_in[987] ;
 wire \inv_in[988] ;
 wire \inv_in[989] ;
 wire \inv_in[98] ;
 wire \inv_in[990] ;
 wire \inv_in[991] ;
 wire \inv_in[992] ;
 wire \inv_in[993] ;
 wire \inv_in[994] ;
 wire \inv_in[995] ;
 wire \inv_in[996] ;
 wire \inv_in[997] ;
 wire \inv_in[998] ;
 wire \inv_in[999] ;
 wire \inv_in[99] ;
 wire \inv_in[9] ;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;

 sg13g2_fill_2 FILLER_0_0 ();
 sg13g2_tiehi _04__18 (.L_HI(net18));
 sg13g2_buf_1 _04_ (.A(net18),
    .X(uio_oe[1]));
 sg13g2_buf_1 _05_ (.A(net19),
    .X(uio_oe[2]));
 sg13g2_buf_1 _06_ (.A(net20),
    .X(uio_oe[3]));
 sg13g2_buf_1 _07_ (.A(net21),
    .X(uio_oe[4]));
 sg13g2_buf_1 _08_ (.A(net22),
    .X(uio_oe[5]));
 sg13g2_buf_1 _09_ (.A(net23),
    .X(uio_oe[6]));
 sg13g2_buf_1 _10_ (.A(net24),
    .X(uio_oe[7]));
 sg13g2_buf_1 _11_ (.A(\inv_in[201] ),
    .X(net2));
 sg13g2_buf_1 _12_ (.A(\inv_in[501] ),
    .X(net3));
 sg13g2_buf_1 _13_ (.A(\inv_in[1001] ),
    .X(net4));
 sg13g2_buf_1 _14_ (.A(\inv_in[2001] ),
    .X(net5));
 sg13g2_buf_1 _15_ (.A(\inv_in[3001] ),
    .X(net6));
 sg13g2_buf_1 _16_ (.A(net16),
    .X(uio_out[6]));
 sg13g2_buf_1 _17_ (.A(net17),
    .X(uio_out[7]));
 sg13g2_buf_1 _18_ (.A(\inv_in[1] ),
    .X(net8));
 sg13g2_buf_1 _19_ (.A(\inv_in[3] ),
    .X(net9));
 sg13g2_buf_1 _20_ (.A(\inv_in[5] ),
    .X(net10));
 sg13g2_buf_1 _21_ (.A(\inv_in[7] ),
    .X(net11));
 sg13g2_buf_1 _22_ (.A(\inv_in[11] ),
    .X(net12));
 sg13g2_buf_1 _23_ (.A(\inv_in[21] ),
    .X(net13));
 sg13g2_buf_1 _24_ (.A(\inv_in[51] ),
    .X(net14));
 sg13g2_buf_1 _25_ (.A(\inv_in[101] ),
    .X(net15));
 sg13g2_buf_1 _26_ (.A(net25),
    .X(uio_oe[0]));
 sg13g2_inv_16 \inv[0]/_0_  (.A(net1),
    .Y(\inv_in[1] ));
 sg13g2_inv_2 \inv[1000]/_0_  (.Y(\inv_in[1001] ),
    .A(\inv_in[1000] ));
 sg13g2_inv_2 \inv[1001]/_0_  (.Y(\inv_in[1002] ),
    .A(\inv_in[1001] ));
 sg13g2_inv_2 \inv[1002]/_0_  (.Y(\inv_in[1003] ),
    .A(\inv_in[1002] ));
 sg13g2_inv_2 \inv[1003]/_0_  (.Y(\inv_in[1004] ),
    .A(\inv_in[1003] ));
 sg13g2_inv_2 \inv[1004]/_0_  (.Y(\inv_in[1005] ),
    .A(\inv_in[1004] ));
 sg13g2_inv_2 \inv[1005]/_0_  (.Y(\inv_in[1006] ),
    .A(\inv_in[1005] ));
 sg13g2_inv_2 \inv[1006]/_0_  (.Y(\inv_in[1007] ),
    .A(\inv_in[1006] ));
 sg13g2_inv_2 \inv[1007]/_0_  (.Y(\inv_in[1008] ),
    .A(\inv_in[1007] ));
 sg13g2_inv_2 \inv[1008]/_0_  (.Y(\inv_in[1009] ),
    .A(\inv_in[1008] ));
 sg13g2_inv_2 \inv[1009]/_0_  (.Y(\inv_in[1010] ),
    .A(\inv_in[1009] ));
 sg13g2_inv_2 \inv[100]/_0_  (.Y(\inv_in[101] ),
    .A(\inv_in[100] ));
 sg13g2_inv_2 \inv[1010]/_0_  (.Y(\inv_in[1011] ),
    .A(\inv_in[1010] ));
 sg13g2_inv_2 \inv[1011]/_0_  (.Y(\inv_in[1012] ),
    .A(\inv_in[1011] ));
 sg13g2_inv_2 \inv[1012]/_0_  (.Y(\inv_in[1013] ),
    .A(\inv_in[1012] ));
 sg13g2_inv_2 \inv[1013]/_0_  (.Y(\inv_in[1014] ),
    .A(\inv_in[1013] ));
 sg13g2_inv_2 \inv[1014]/_0_  (.Y(\inv_in[1015] ),
    .A(\inv_in[1014] ));
 sg13g2_inv_2 \inv[1015]/_0_  (.Y(\inv_in[1016] ),
    .A(\inv_in[1015] ));
 sg13g2_inv_2 \inv[1016]/_0_  (.Y(\inv_in[1017] ),
    .A(\inv_in[1016] ));
 sg13g2_inv_2 \inv[1017]/_0_  (.Y(\inv_in[1018] ),
    .A(\inv_in[1017] ));
 sg13g2_inv_2 \inv[1018]/_0_  (.Y(\inv_in[1019] ),
    .A(\inv_in[1018] ));
 sg13g2_inv_2 \inv[1019]/_0_  (.Y(\inv_in[1020] ),
    .A(\inv_in[1019] ));
 sg13g2_inv_2 \inv[101]/_0_  (.Y(\inv_in[102] ),
    .A(\inv_in[101] ));
 sg13g2_inv_2 \inv[1020]/_0_  (.Y(\inv_in[1021] ),
    .A(\inv_in[1020] ));
 sg13g2_inv_2 \inv[1021]/_0_  (.Y(\inv_in[1022] ),
    .A(\inv_in[1021] ));
 sg13g2_inv_2 \inv[1022]/_0_  (.Y(\inv_in[1023] ),
    .A(\inv_in[1022] ));
 sg13g2_inv_2 \inv[1023]/_0_  (.Y(\inv_in[1024] ),
    .A(\inv_in[1023] ));
 sg13g2_inv_2 \inv[1024]/_0_  (.Y(\inv_in[1025] ),
    .A(\inv_in[1024] ));
 sg13g2_inv_2 \inv[1025]/_0_  (.Y(\inv_in[1026] ),
    .A(\inv_in[1025] ));
 sg13g2_inv_2 \inv[1026]/_0_  (.Y(\inv_in[1027] ),
    .A(\inv_in[1026] ));
 sg13g2_inv_2 \inv[1027]/_0_  (.Y(\inv_in[1028] ),
    .A(\inv_in[1027] ));
 sg13g2_inv_2 \inv[1028]/_0_  (.Y(\inv_in[1029] ),
    .A(\inv_in[1028] ));
 sg13g2_inv_2 \inv[1029]/_0_  (.Y(\inv_in[1030] ),
    .A(\inv_in[1029] ));
 sg13g2_inv_2 \inv[102]/_0_  (.Y(\inv_in[103] ),
    .A(\inv_in[102] ));
 sg13g2_inv_2 \inv[1030]/_0_  (.Y(\inv_in[1031] ),
    .A(\inv_in[1030] ));
 sg13g2_inv_2 \inv[1031]/_0_  (.Y(\inv_in[1032] ),
    .A(\inv_in[1031] ));
 sg13g2_inv_2 \inv[1032]/_0_  (.Y(\inv_in[1033] ),
    .A(\inv_in[1032] ));
 sg13g2_inv_2 \inv[1033]/_0_  (.Y(\inv_in[1034] ),
    .A(\inv_in[1033] ));
 sg13g2_inv_2 \inv[1034]/_0_  (.Y(\inv_in[1035] ),
    .A(\inv_in[1034] ));
 sg13g2_inv_2 \inv[1035]/_0_  (.Y(\inv_in[1036] ),
    .A(\inv_in[1035] ));
 sg13g2_inv_2 \inv[1036]/_0_  (.Y(\inv_in[1037] ),
    .A(\inv_in[1036] ));
 sg13g2_inv_2 \inv[1037]/_0_  (.Y(\inv_in[1038] ),
    .A(\inv_in[1037] ));
 sg13g2_inv_2 \inv[1038]/_0_  (.Y(\inv_in[1039] ),
    .A(\inv_in[1038] ));
 sg13g2_inv_2 \inv[1039]/_0_  (.Y(\inv_in[1040] ),
    .A(\inv_in[1039] ));
 sg13g2_inv_2 \inv[103]/_0_  (.Y(\inv_in[104] ),
    .A(\inv_in[103] ));
 sg13g2_inv_2 \inv[1040]/_0_  (.Y(\inv_in[1041] ),
    .A(\inv_in[1040] ));
 sg13g2_inv_2 \inv[1041]/_0_  (.Y(\inv_in[1042] ),
    .A(\inv_in[1041] ));
 sg13g2_inv_2 \inv[1042]/_0_  (.Y(\inv_in[1043] ),
    .A(\inv_in[1042] ));
 sg13g2_inv_2 \inv[1043]/_0_  (.Y(\inv_in[1044] ),
    .A(\inv_in[1043] ));
 sg13g2_inv_2 \inv[1044]/_0_  (.Y(\inv_in[1045] ),
    .A(\inv_in[1044] ));
 sg13g2_inv_2 \inv[1045]/_0_  (.Y(\inv_in[1046] ),
    .A(\inv_in[1045] ));
 sg13g2_inv_2 \inv[1046]/_0_  (.Y(\inv_in[1047] ),
    .A(\inv_in[1046] ));
 sg13g2_inv_2 \inv[1047]/_0_  (.Y(\inv_in[1048] ),
    .A(\inv_in[1047] ));
 sg13g2_inv_2 \inv[1048]/_0_  (.Y(\inv_in[1049] ),
    .A(\inv_in[1048] ));
 sg13g2_inv_2 \inv[1049]/_0_  (.Y(\inv_in[1050] ),
    .A(\inv_in[1049] ));
 sg13g2_inv_2 \inv[104]/_0_  (.Y(\inv_in[105] ),
    .A(\inv_in[104] ));
 sg13g2_inv_2 \inv[1050]/_0_  (.Y(\inv_in[1051] ),
    .A(\inv_in[1050] ));
 sg13g2_inv_2 \inv[1051]/_0_  (.Y(\inv_in[1052] ),
    .A(\inv_in[1051] ));
 sg13g2_inv_2 \inv[1052]/_0_  (.Y(\inv_in[1053] ),
    .A(\inv_in[1052] ));
 sg13g2_inv_2 \inv[1053]/_0_  (.Y(\inv_in[1054] ),
    .A(\inv_in[1053] ));
 sg13g2_inv_2 \inv[1054]/_0_  (.Y(\inv_in[1055] ),
    .A(\inv_in[1054] ));
 sg13g2_inv_2 \inv[1055]/_0_  (.Y(\inv_in[1056] ),
    .A(\inv_in[1055] ));
 sg13g2_inv_2 \inv[1056]/_0_  (.Y(\inv_in[1057] ),
    .A(\inv_in[1056] ));
 sg13g2_inv_2 \inv[1057]/_0_  (.Y(\inv_in[1058] ),
    .A(\inv_in[1057] ));
 sg13g2_inv_2 \inv[1058]/_0_  (.Y(\inv_in[1059] ),
    .A(\inv_in[1058] ));
 sg13g2_inv_2 \inv[1059]/_0_  (.Y(\inv_in[1060] ),
    .A(\inv_in[1059] ));
 sg13g2_inv_2 \inv[105]/_0_  (.Y(\inv_in[106] ),
    .A(\inv_in[105] ));
 sg13g2_inv_2 \inv[1060]/_0_  (.Y(\inv_in[1061] ),
    .A(\inv_in[1060] ));
 sg13g2_inv_2 \inv[1061]/_0_  (.Y(\inv_in[1062] ),
    .A(\inv_in[1061] ));
 sg13g2_inv_2 \inv[1062]/_0_  (.Y(\inv_in[1063] ),
    .A(\inv_in[1062] ));
 sg13g2_inv_2 \inv[1063]/_0_  (.Y(\inv_in[1064] ),
    .A(\inv_in[1063] ));
 sg13g2_inv_2 \inv[1064]/_0_  (.Y(\inv_in[1065] ),
    .A(\inv_in[1064] ));
 sg13g2_inv_2 \inv[1065]/_0_  (.Y(\inv_in[1066] ),
    .A(\inv_in[1065] ));
 sg13g2_inv_2 \inv[1066]/_0_  (.Y(\inv_in[1067] ),
    .A(\inv_in[1066] ));
 sg13g2_inv_2 \inv[1067]/_0_  (.Y(\inv_in[1068] ),
    .A(\inv_in[1067] ));
 sg13g2_inv_2 \inv[1068]/_0_  (.Y(\inv_in[1069] ),
    .A(\inv_in[1068] ));
 sg13g2_inv_2 \inv[1069]/_0_  (.Y(\inv_in[1070] ),
    .A(\inv_in[1069] ));
 sg13g2_inv_2 \inv[106]/_0_  (.Y(\inv_in[107] ),
    .A(\inv_in[106] ));
 sg13g2_inv_2 \inv[1070]/_0_  (.Y(\inv_in[1071] ),
    .A(\inv_in[1070] ));
 sg13g2_inv_2 \inv[1071]/_0_  (.Y(\inv_in[1072] ),
    .A(\inv_in[1071] ));
 sg13g2_inv_2 \inv[1072]/_0_  (.Y(\inv_in[1073] ),
    .A(\inv_in[1072] ));
 sg13g2_inv_2 \inv[1073]/_0_  (.Y(\inv_in[1074] ),
    .A(\inv_in[1073] ));
 sg13g2_inv_2 \inv[1074]/_0_  (.Y(\inv_in[1075] ),
    .A(\inv_in[1074] ));
 sg13g2_inv_2 \inv[1075]/_0_  (.Y(\inv_in[1076] ),
    .A(\inv_in[1075] ));
 sg13g2_inv_2 \inv[1076]/_0_  (.Y(\inv_in[1077] ),
    .A(\inv_in[1076] ));
 sg13g2_inv_2 \inv[1077]/_0_  (.Y(\inv_in[1078] ),
    .A(\inv_in[1077] ));
 sg13g2_inv_2 \inv[1078]/_0_  (.Y(\inv_in[1079] ),
    .A(\inv_in[1078] ));
 sg13g2_inv_2 \inv[1079]/_0_  (.Y(\inv_in[1080] ),
    .A(\inv_in[1079] ));
 sg13g2_inv_2 \inv[107]/_0_  (.Y(\inv_in[108] ),
    .A(\inv_in[107] ));
 sg13g2_inv_2 \inv[1080]/_0_  (.Y(\inv_in[1081] ),
    .A(\inv_in[1080] ));
 sg13g2_inv_2 \inv[1081]/_0_  (.Y(\inv_in[1082] ),
    .A(\inv_in[1081] ));
 sg13g2_inv_2 \inv[1082]/_0_  (.Y(\inv_in[1083] ),
    .A(\inv_in[1082] ));
 sg13g2_inv_2 \inv[1083]/_0_  (.Y(\inv_in[1084] ),
    .A(\inv_in[1083] ));
 sg13g2_inv_2 \inv[1084]/_0_  (.Y(\inv_in[1085] ),
    .A(\inv_in[1084] ));
 sg13g2_inv_2 \inv[1085]/_0_  (.Y(\inv_in[1086] ),
    .A(\inv_in[1085] ));
 sg13g2_inv_2 \inv[1086]/_0_  (.Y(\inv_in[1087] ),
    .A(\inv_in[1086] ));
 sg13g2_inv_2 \inv[1087]/_0_  (.Y(\inv_in[1088] ),
    .A(\inv_in[1087] ));
 sg13g2_inv_2 \inv[1088]/_0_  (.Y(\inv_in[1089] ),
    .A(\inv_in[1088] ));
 sg13g2_inv_2 \inv[1089]/_0_  (.Y(\inv_in[1090] ),
    .A(\inv_in[1089] ));
 sg13g2_inv_2 \inv[108]/_0_  (.Y(\inv_in[109] ),
    .A(\inv_in[108] ));
 sg13g2_inv_2 \inv[1090]/_0_  (.Y(\inv_in[1091] ),
    .A(\inv_in[1090] ));
 sg13g2_inv_2 \inv[1091]/_0_  (.Y(\inv_in[1092] ),
    .A(\inv_in[1091] ));
 sg13g2_inv_2 \inv[1092]/_0_  (.Y(\inv_in[1093] ),
    .A(\inv_in[1092] ));
 sg13g2_inv_2 \inv[1093]/_0_  (.Y(\inv_in[1094] ),
    .A(\inv_in[1093] ));
 sg13g2_inv_2 \inv[1094]/_0_  (.Y(\inv_in[1095] ),
    .A(\inv_in[1094] ));
 sg13g2_inv_2 \inv[1095]/_0_  (.Y(\inv_in[1096] ),
    .A(\inv_in[1095] ));
 sg13g2_inv_2 \inv[1096]/_0_  (.Y(\inv_in[1097] ),
    .A(\inv_in[1096] ));
 sg13g2_inv_2 \inv[1097]/_0_  (.Y(\inv_in[1098] ),
    .A(\inv_in[1097] ));
 sg13g2_inv_2 \inv[1098]/_0_  (.Y(\inv_in[1099] ),
    .A(\inv_in[1098] ));
 sg13g2_inv_2 \inv[1099]/_0_  (.Y(\inv_in[1100] ),
    .A(\inv_in[1099] ));
 sg13g2_inv_2 \inv[109]/_0_  (.Y(\inv_in[110] ),
    .A(\inv_in[109] ));
 sg13g2_inv_2 \inv[10]/_0_  (.Y(\inv_in[11] ),
    .A(\inv_in[10] ));
 sg13g2_inv_2 \inv[1100]/_0_  (.Y(\inv_in[1101] ),
    .A(\inv_in[1100] ));
 sg13g2_inv_2 \inv[1101]/_0_  (.Y(\inv_in[1102] ),
    .A(\inv_in[1101] ));
 sg13g2_inv_2 \inv[1102]/_0_  (.Y(\inv_in[1103] ),
    .A(\inv_in[1102] ));
 sg13g2_inv_2 \inv[1103]/_0_  (.Y(\inv_in[1104] ),
    .A(\inv_in[1103] ));
 sg13g2_inv_2 \inv[1104]/_0_  (.Y(\inv_in[1105] ),
    .A(\inv_in[1104] ));
 sg13g2_inv_2 \inv[1105]/_0_  (.Y(\inv_in[1106] ),
    .A(\inv_in[1105] ));
 sg13g2_inv_2 \inv[1106]/_0_  (.Y(\inv_in[1107] ),
    .A(\inv_in[1106] ));
 sg13g2_inv_2 \inv[1107]/_0_  (.Y(\inv_in[1108] ),
    .A(\inv_in[1107] ));
 sg13g2_inv_2 \inv[1108]/_0_  (.Y(\inv_in[1109] ),
    .A(\inv_in[1108] ));
 sg13g2_inv_2 \inv[1109]/_0_  (.Y(\inv_in[1110] ),
    .A(\inv_in[1109] ));
 sg13g2_inv_2 \inv[110]/_0_  (.Y(\inv_in[111] ),
    .A(\inv_in[110] ));
 sg13g2_inv_2 \inv[1110]/_0_  (.Y(\inv_in[1111] ),
    .A(\inv_in[1110] ));
 sg13g2_inv_2 \inv[1111]/_0_  (.Y(\inv_in[1112] ),
    .A(\inv_in[1111] ));
 sg13g2_inv_2 \inv[1112]/_0_  (.Y(\inv_in[1113] ),
    .A(\inv_in[1112] ));
 sg13g2_inv_2 \inv[1113]/_0_  (.Y(\inv_in[1114] ),
    .A(\inv_in[1113] ));
 sg13g2_inv_2 \inv[1114]/_0_  (.Y(\inv_in[1115] ),
    .A(\inv_in[1114] ));
 sg13g2_inv_2 \inv[1115]/_0_  (.Y(\inv_in[1116] ),
    .A(\inv_in[1115] ));
 sg13g2_inv_2 \inv[1116]/_0_  (.Y(\inv_in[1117] ),
    .A(\inv_in[1116] ));
 sg13g2_inv_2 \inv[1117]/_0_  (.Y(\inv_in[1118] ),
    .A(\inv_in[1117] ));
 sg13g2_inv_2 \inv[1118]/_0_  (.Y(\inv_in[1119] ),
    .A(\inv_in[1118] ));
 sg13g2_inv_2 \inv[1119]/_0_  (.Y(\inv_in[1120] ),
    .A(\inv_in[1119] ));
 sg13g2_inv_2 \inv[111]/_0_  (.Y(\inv_in[112] ),
    .A(\inv_in[111] ));
 sg13g2_inv_2 \inv[1120]/_0_  (.Y(\inv_in[1121] ),
    .A(\inv_in[1120] ));
 sg13g2_inv_2 \inv[1121]/_0_  (.Y(\inv_in[1122] ),
    .A(\inv_in[1121] ));
 sg13g2_inv_2 \inv[1122]/_0_  (.Y(\inv_in[1123] ),
    .A(\inv_in[1122] ));
 sg13g2_inv_2 \inv[1123]/_0_  (.Y(\inv_in[1124] ),
    .A(\inv_in[1123] ));
 sg13g2_inv_2 \inv[1124]/_0_  (.Y(\inv_in[1125] ),
    .A(\inv_in[1124] ));
 sg13g2_inv_2 \inv[1125]/_0_  (.Y(\inv_in[1126] ),
    .A(\inv_in[1125] ));
 sg13g2_inv_2 \inv[1126]/_0_  (.Y(\inv_in[1127] ),
    .A(\inv_in[1126] ));
 sg13g2_inv_2 \inv[1127]/_0_  (.Y(\inv_in[1128] ),
    .A(\inv_in[1127] ));
 sg13g2_inv_2 \inv[1128]/_0_  (.Y(\inv_in[1129] ),
    .A(\inv_in[1128] ));
 sg13g2_inv_2 \inv[1129]/_0_  (.Y(\inv_in[1130] ),
    .A(\inv_in[1129] ));
 sg13g2_inv_2 \inv[112]/_0_  (.Y(\inv_in[113] ),
    .A(\inv_in[112] ));
 sg13g2_inv_2 \inv[1130]/_0_  (.Y(\inv_in[1131] ),
    .A(\inv_in[1130] ));
 sg13g2_inv_2 \inv[1131]/_0_  (.Y(\inv_in[1132] ),
    .A(\inv_in[1131] ));
 sg13g2_inv_2 \inv[1132]/_0_  (.Y(\inv_in[1133] ),
    .A(\inv_in[1132] ));
 sg13g2_inv_2 \inv[1133]/_0_  (.Y(\inv_in[1134] ),
    .A(\inv_in[1133] ));
 sg13g2_inv_2 \inv[1134]/_0_  (.Y(\inv_in[1135] ),
    .A(\inv_in[1134] ));
 sg13g2_inv_2 \inv[1135]/_0_  (.Y(\inv_in[1136] ),
    .A(\inv_in[1135] ));
 sg13g2_inv_2 \inv[1136]/_0_  (.Y(\inv_in[1137] ),
    .A(\inv_in[1136] ));
 sg13g2_inv_2 \inv[1137]/_0_  (.Y(\inv_in[1138] ),
    .A(\inv_in[1137] ));
 sg13g2_inv_2 \inv[1138]/_0_  (.Y(\inv_in[1139] ),
    .A(\inv_in[1138] ));
 sg13g2_inv_2 \inv[1139]/_0_  (.Y(\inv_in[1140] ),
    .A(\inv_in[1139] ));
 sg13g2_inv_2 \inv[113]/_0_  (.Y(\inv_in[114] ),
    .A(\inv_in[113] ));
 sg13g2_inv_2 \inv[1140]/_0_  (.Y(\inv_in[1141] ),
    .A(\inv_in[1140] ));
 sg13g2_inv_2 \inv[1141]/_0_  (.Y(\inv_in[1142] ),
    .A(\inv_in[1141] ));
 sg13g2_inv_2 \inv[1142]/_0_  (.Y(\inv_in[1143] ),
    .A(\inv_in[1142] ));
 sg13g2_inv_2 \inv[1143]/_0_  (.Y(\inv_in[1144] ),
    .A(\inv_in[1143] ));
 sg13g2_inv_2 \inv[1144]/_0_  (.Y(\inv_in[1145] ),
    .A(\inv_in[1144] ));
 sg13g2_inv_2 \inv[1145]/_0_  (.Y(\inv_in[1146] ),
    .A(\inv_in[1145] ));
 sg13g2_inv_2 \inv[1146]/_0_  (.Y(\inv_in[1147] ),
    .A(\inv_in[1146] ));
 sg13g2_inv_2 \inv[1147]/_0_  (.Y(\inv_in[1148] ),
    .A(\inv_in[1147] ));
 sg13g2_inv_2 \inv[1148]/_0_  (.Y(\inv_in[1149] ),
    .A(\inv_in[1148] ));
 sg13g2_inv_2 \inv[1149]/_0_  (.Y(\inv_in[1150] ),
    .A(\inv_in[1149] ));
 sg13g2_inv_2 \inv[114]/_0_  (.Y(\inv_in[115] ),
    .A(\inv_in[114] ));
 sg13g2_inv_2 \inv[1150]/_0_  (.Y(\inv_in[1151] ),
    .A(\inv_in[1150] ));
 sg13g2_inv_2 \inv[1151]/_0_  (.Y(\inv_in[1152] ),
    .A(\inv_in[1151] ));
 sg13g2_inv_2 \inv[1152]/_0_  (.Y(\inv_in[1153] ),
    .A(\inv_in[1152] ));
 sg13g2_inv_2 \inv[1153]/_0_  (.Y(\inv_in[1154] ),
    .A(\inv_in[1153] ));
 sg13g2_inv_2 \inv[1154]/_0_  (.Y(\inv_in[1155] ),
    .A(\inv_in[1154] ));
 sg13g2_inv_2 \inv[1155]/_0_  (.Y(\inv_in[1156] ),
    .A(\inv_in[1155] ));
 sg13g2_inv_2 \inv[1156]/_0_  (.Y(\inv_in[1157] ),
    .A(\inv_in[1156] ));
 sg13g2_inv_2 \inv[1157]/_0_  (.Y(\inv_in[1158] ),
    .A(\inv_in[1157] ));
 sg13g2_inv_2 \inv[1158]/_0_  (.Y(\inv_in[1159] ),
    .A(\inv_in[1158] ));
 sg13g2_inv_2 \inv[1159]/_0_  (.Y(\inv_in[1160] ),
    .A(\inv_in[1159] ));
 sg13g2_inv_2 \inv[115]/_0_  (.Y(\inv_in[116] ),
    .A(\inv_in[115] ));
 sg13g2_inv_2 \inv[1160]/_0_  (.Y(\inv_in[1161] ),
    .A(\inv_in[1160] ));
 sg13g2_inv_2 \inv[1161]/_0_  (.Y(\inv_in[1162] ),
    .A(\inv_in[1161] ));
 sg13g2_inv_2 \inv[1162]/_0_  (.Y(\inv_in[1163] ),
    .A(\inv_in[1162] ));
 sg13g2_inv_2 \inv[1163]/_0_  (.Y(\inv_in[1164] ),
    .A(\inv_in[1163] ));
 sg13g2_inv_2 \inv[1164]/_0_  (.Y(\inv_in[1165] ),
    .A(\inv_in[1164] ));
 sg13g2_inv_2 \inv[1165]/_0_  (.Y(\inv_in[1166] ),
    .A(\inv_in[1165] ));
 sg13g2_inv_2 \inv[1166]/_0_  (.Y(\inv_in[1167] ),
    .A(\inv_in[1166] ));
 sg13g2_inv_2 \inv[1167]/_0_  (.Y(\inv_in[1168] ),
    .A(\inv_in[1167] ));
 sg13g2_inv_2 \inv[1168]/_0_  (.Y(\inv_in[1169] ),
    .A(\inv_in[1168] ));
 sg13g2_inv_2 \inv[1169]/_0_  (.Y(\inv_in[1170] ),
    .A(\inv_in[1169] ));
 sg13g2_inv_2 \inv[116]/_0_  (.Y(\inv_in[117] ),
    .A(\inv_in[116] ));
 sg13g2_inv_2 \inv[1170]/_0_  (.Y(\inv_in[1171] ),
    .A(\inv_in[1170] ));
 sg13g2_inv_2 \inv[1171]/_0_  (.Y(\inv_in[1172] ),
    .A(\inv_in[1171] ));
 sg13g2_inv_2 \inv[1172]/_0_  (.Y(\inv_in[1173] ),
    .A(\inv_in[1172] ));
 sg13g2_inv_2 \inv[1173]/_0_  (.Y(\inv_in[1174] ),
    .A(\inv_in[1173] ));
 sg13g2_inv_2 \inv[1174]/_0_  (.Y(\inv_in[1175] ),
    .A(\inv_in[1174] ));
 sg13g2_inv_2 \inv[1175]/_0_  (.Y(\inv_in[1176] ),
    .A(\inv_in[1175] ));
 sg13g2_inv_2 \inv[1176]/_0_  (.Y(\inv_in[1177] ),
    .A(\inv_in[1176] ));
 sg13g2_inv_2 \inv[1177]/_0_  (.Y(\inv_in[1178] ),
    .A(\inv_in[1177] ));
 sg13g2_inv_2 \inv[1178]/_0_  (.Y(\inv_in[1179] ),
    .A(\inv_in[1178] ));
 sg13g2_inv_2 \inv[1179]/_0_  (.Y(\inv_in[1180] ),
    .A(\inv_in[1179] ));
 sg13g2_inv_2 \inv[117]/_0_  (.Y(\inv_in[118] ),
    .A(\inv_in[117] ));
 sg13g2_inv_2 \inv[1180]/_0_  (.Y(\inv_in[1181] ),
    .A(\inv_in[1180] ));
 sg13g2_inv_2 \inv[1181]/_0_  (.Y(\inv_in[1182] ),
    .A(\inv_in[1181] ));
 sg13g2_inv_2 \inv[1182]/_0_  (.Y(\inv_in[1183] ),
    .A(\inv_in[1182] ));
 sg13g2_inv_2 \inv[1183]/_0_  (.Y(\inv_in[1184] ),
    .A(\inv_in[1183] ));
 sg13g2_inv_2 \inv[1184]/_0_  (.Y(\inv_in[1185] ),
    .A(\inv_in[1184] ));
 sg13g2_inv_2 \inv[1185]/_0_  (.Y(\inv_in[1186] ),
    .A(\inv_in[1185] ));
 sg13g2_inv_2 \inv[1186]/_0_  (.Y(\inv_in[1187] ),
    .A(\inv_in[1186] ));
 sg13g2_inv_2 \inv[1187]/_0_  (.Y(\inv_in[1188] ),
    .A(\inv_in[1187] ));
 sg13g2_inv_2 \inv[1188]/_0_  (.Y(\inv_in[1189] ),
    .A(\inv_in[1188] ));
 sg13g2_inv_2 \inv[1189]/_0_  (.Y(\inv_in[1190] ),
    .A(\inv_in[1189] ));
 sg13g2_inv_2 \inv[118]/_0_  (.Y(\inv_in[119] ),
    .A(\inv_in[118] ));
 sg13g2_inv_2 \inv[1190]/_0_  (.Y(\inv_in[1191] ),
    .A(\inv_in[1190] ));
 sg13g2_inv_2 \inv[1191]/_0_  (.Y(\inv_in[1192] ),
    .A(\inv_in[1191] ));
 sg13g2_inv_2 \inv[1192]/_0_  (.Y(\inv_in[1193] ),
    .A(\inv_in[1192] ));
 sg13g2_inv_2 \inv[1193]/_0_  (.Y(\inv_in[1194] ),
    .A(\inv_in[1193] ));
 sg13g2_inv_2 \inv[1194]/_0_  (.Y(\inv_in[1195] ),
    .A(\inv_in[1194] ));
 sg13g2_inv_2 \inv[1195]/_0_  (.Y(\inv_in[1196] ),
    .A(\inv_in[1195] ));
 sg13g2_inv_2 \inv[1196]/_0_  (.Y(\inv_in[1197] ),
    .A(\inv_in[1196] ));
 sg13g2_inv_2 \inv[1197]/_0_  (.Y(\inv_in[1198] ),
    .A(\inv_in[1197] ));
 sg13g2_inv_2 \inv[1198]/_0_  (.Y(\inv_in[1199] ),
    .A(\inv_in[1198] ));
 sg13g2_inv_2 \inv[1199]/_0_  (.Y(\inv_in[1200] ),
    .A(\inv_in[1199] ));
 sg13g2_inv_2 \inv[119]/_0_  (.Y(\inv_in[120] ),
    .A(\inv_in[119] ));
 sg13g2_inv_2 \inv[11]/_0_  (.Y(\inv_in[12] ),
    .A(\inv_in[11] ));
 sg13g2_inv_2 \inv[1200]/_0_  (.Y(\inv_in[1201] ),
    .A(\inv_in[1200] ));
 sg13g2_inv_2 \inv[1201]/_0_  (.Y(\inv_in[1202] ),
    .A(\inv_in[1201] ));
 sg13g2_inv_2 \inv[1202]/_0_  (.Y(\inv_in[1203] ),
    .A(\inv_in[1202] ));
 sg13g2_inv_2 \inv[1203]/_0_  (.Y(\inv_in[1204] ),
    .A(\inv_in[1203] ));
 sg13g2_inv_2 \inv[1204]/_0_  (.Y(\inv_in[1205] ),
    .A(\inv_in[1204] ));
 sg13g2_inv_2 \inv[1205]/_0_  (.Y(\inv_in[1206] ),
    .A(\inv_in[1205] ));
 sg13g2_inv_2 \inv[1206]/_0_  (.Y(\inv_in[1207] ),
    .A(\inv_in[1206] ));
 sg13g2_inv_2 \inv[1207]/_0_  (.Y(\inv_in[1208] ),
    .A(\inv_in[1207] ));
 sg13g2_inv_2 \inv[1208]/_0_  (.Y(\inv_in[1209] ),
    .A(\inv_in[1208] ));
 sg13g2_inv_2 \inv[1209]/_0_  (.Y(\inv_in[1210] ),
    .A(\inv_in[1209] ));
 sg13g2_inv_2 \inv[120]/_0_  (.Y(\inv_in[121] ),
    .A(\inv_in[120] ));
 sg13g2_inv_2 \inv[1210]/_0_  (.Y(\inv_in[1211] ),
    .A(\inv_in[1210] ));
 sg13g2_inv_2 \inv[1211]/_0_  (.Y(\inv_in[1212] ),
    .A(\inv_in[1211] ));
 sg13g2_inv_2 \inv[1212]/_0_  (.Y(\inv_in[1213] ),
    .A(\inv_in[1212] ));
 sg13g2_inv_2 \inv[1213]/_0_  (.Y(\inv_in[1214] ),
    .A(\inv_in[1213] ));
 sg13g2_inv_2 \inv[1214]/_0_  (.Y(\inv_in[1215] ),
    .A(\inv_in[1214] ));
 sg13g2_inv_2 \inv[1215]/_0_  (.Y(\inv_in[1216] ),
    .A(\inv_in[1215] ));
 sg13g2_inv_2 \inv[1216]/_0_  (.Y(\inv_in[1217] ),
    .A(\inv_in[1216] ));
 sg13g2_inv_2 \inv[1217]/_0_  (.Y(\inv_in[1218] ),
    .A(\inv_in[1217] ));
 sg13g2_inv_2 \inv[1218]/_0_  (.Y(\inv_in[1219] ),
    .A(\inv_in[1218] ));
 sg13g2_inv_2 \inv[1219]/_0_  (.Y(\inv_in[1220] ),
    .A(\inv_in[1219] ));
 sg13g2_inv_2 \inv[121]/_0_  (.Y(\inv_in[122] ),
    .A(\inv_in[121] ));
 sg13g2_inv_2 \inv[1220]/_0_  (.Y(\inv_in[1221] ),
    .A(\inv_in[1220] ));
 sg13g2_inv_2 \inv[1221]/_0_  (.Y(\inv_in[1222] ),
    .A(\inv_in[1221] ));
 sg13g2_inv_2 \inv[1222]/_0_  (.Y(\inv_in[1223] ),
    .A(\inv_in[1222] ));
 sg13g2_inv_2 \inv[1223]/_0_  (.Y(\inv_in[1224] ),
    .A(\inv_in[1223] ));
 sg13g2_inv_2 \inv[1224]/_0_  (.Y(\inv_in[1225] ),
    .A(\inv_in[1224] ));
 sg13g2_inv_2 \inv[1225]/_0_  (.Y(\inv_in[1226] ),
    .A(\inv_in[1225] ));
 sg13g2_inv_2 \inv[1226]/_0_  (.Y(\inv_in[1227] ),
    .A(\inv_in[1226] ));
 sg13g2_inv_2 \inv[1227]/_0_  (.Y(\inv_in[1228] ),
    .A(\inv_in[1227] ));
 sg13g2_inv_2 \inv[1228]/_0_  (.Y(\inv_in[1229] ),
    .A(\inv_in[1228] ));
 sg13g2_inv_2 \inv[1229]/_0_  (.Y(\inv_in[1230] ),
    .A(\inv_in[1229] ));
 sg13g2_inv_2 \inv[122]/_0_  (.Y(\inv_in[123] ),
    .A(\inv_in[122] ));
 sg13g2_inv_2 \inv[1230]/_0_  (.Y(\inv_in[1231] ),
    .A(\inv_in[1230] ));
 sg13g2_inv_2 \inv[1231]/_0_  (.Y(\inv_in[1232] ),
    .A(\inv_in[1231] ));
 sg13g2_inv_2 \inv[1232]/_0_  (.Y(\inv_in[1233] ),
    .A(\inv_in[1232] ));
 sg13g2_inv_2 \inv[1233]/_0_  (.Y(\inv_in[1234] ),
    .A(\inv_in[1233] ));
 sg13g2_inv_2 \inv[1234]/_0_  (.Y(\inv_in[1235] ),
    .A(\inv_in[1234] ));
 sg13g2_inv_2 \inv[1235]/_0_  (.Y(\inv_in[1236] ),
    .A(\inv_in[1235] ));
 sg13g2_inv_2 \inv[1236]/_0_  (.Y(\inv_in[1237] ),
    .A(\inv_in[1236] ));
 sg13g2_inv_2 \inv[1237]/_0_  (.Y(\inv_in[1238] ),
    .A(\inv_in[1237] ));
 sg13g2_inv_2 \inv[1238]/_0_  (.Y(\inv_in[1239] ),
    .A(\inv_in[1238] ));
 sg13g2_inv_2 \inv[1239]/_0_  (.Y(\inv_in[1240] ),
    .A(\inv_in[1239] ));
 sg13g2_inv_2 \inv[123]/_0_  (.Y(\inv_in[124] ),
    .A(\inv_in[123] ));
 sg13g2_inv_2 \inv[1240]/_0_  (.Y(\inv_in[1241] ),
    .A(\inv_in[1240] ));
 sg13g2_inv_2 \inv[1241]/_0_  (.Y(\inv_in[1242] ),
    .A(\inv_in[1241] ));
 sg13g2_inv_2 \inv[1242]/_0_  (.Y(\inv_in[1243] ),
    .A(\inv_in[1242] ));
 sg13g2_inv_2 \inv[1243]/_0_  (.Y(\inv_in[1244] ),
    .A(\inv_in[1243] ));
 sg13g2_inv_2 \inv[1244]/_0_  (.Y(\inv_in[1245] ),
    .A(\inv_in[1244] ));
 sg13g2_inv_2 \inv[1245]/_0_  (.Y(\inv_in[1246] ),
    .A(\inv_in[1245] ));
 sg13g2_inv_2 \inv[1246]/_0_  (.Y(\inv_in[1247] ),
    .A(\inv_in[1246] ));
 sg13g2_inv_2 \inv[1247]/_0_  (.Y(\inv_in[1248] ),
    .A(\inv_in[1247] ));
 sg13g2_inv_2 \inv[1248]/_0_  (.Y(\inv_in[1249] ),
    .A(\inv_in[1248] ));
 sg13g2_inv_2 \inv[1249]/_0_  (.Y(\inv_in[1250] ),
    .A(\inv_in[1249] ));
 sg13g2_inv_2 \inv[124]/_0_  (.Y(\inv_in[125] ),
    .A(\inv_in[124] ));
 sg13g2_inv_2 \inv[1250]/_0_  (.Y(\inv_in[1251] ),
    .A(\inv_in[1250] ));
 sg13g2_inv_2 \inv[1251]/_0_  (.Y(\inv_in[1252] ),
    .A(\inv_in[1251] ));
 sg13g2_inv_2 \inv[1252]/_0_  (.Y(\inv_in[1253] ),
    .A(\inv_in[1252] ));
 sg13g2_inv_2 \inv[1253]/_0_  (.Y(\inv_in[1254] ),
    .A(\inv_in[1253] ));
 sg13g2_inv_2 \inv[1254]/_0_  (.Y(\inv_in[1255] ),
    .A(\inv_in[1254] ));
 sg13g2_inv_2 \inv[1255]/_0_  (.Y(\inv_in[1256] ),
    .A(\inv_in[1255] ));
 sg13g2_inv_2 \inv[1256]/_0_  (.Y(\inv_in[1257] ),
    .A(\inv_in[1256] ));
 sg13g2_inv_2 \inv[1257]/_0_  (.Y(\inv_in[1258] ),
    .A(\inv_in[1257] ));
 sg13g2_inv_2 \inv[1258]/_0_  (.Y(\inv_in[1259] ),
    .A(\inv_in[1258] ));
 sg13g2_inv_2 \inv[1259]/_0_  (.Y(\inv_in[1260] ),
    .A(\inv_in[1259] ));
 sg13g2_inv_2 \inv[125]/_0_  (.Y(\inv_in[126] ),
    .A(\inv_in[125] ));
 sg13g2_inv_2 \inv[1260]/_0_  (.Y(\inv_in[1261] ),
    .A(\inv_in[1260] ));
 sg13g2_inv_2 \inv[1261]/_0_  (.Y(\inv_in[1262] ),
    .A(\inv_in[1261] ));
 sg13g2_inv_2 \inv[1262]/_0_  (.Y(\inv_in[1263] ),
    .A(\inv_in[1262] ));
 sg13g2_inv_2 \inv[1263]/_0_  (.Y(\inv_in[1264] ),
    .A(\inv_in[1263] ));
 sg13g2_inv_2 \inv[1264]/_0_  (.Y(\inv_in[1265] ),
    .A(\inv_in[1264] ));
 sg13g2_inv_2 \inv[1265]/_0_  (.Y(\inv_in[1266] ),
    .A(\inv_in[1265] ));
 sg13g2_inv_2 \inv[1266]/_0_  (.Y(\inv_in[1267] ),
    .A(\inv_in[1266] ));
 sg13g2_inv_2 \inv[1267]/_0_  (.Y(\inv_in[1268] ),
    .A(\inv_in[1267] ));
 sg13g2_inv_2 \inv[1268]/_0_  (.Y(\inv_in[1269] ),
    .A(\inv_in[1268] ));
 sg13g2_inv_2 \inv[1269]/_0_  (.Y(\inv_in[1270] ),
    .A(\inv_in[1269] ));
 sg13g2_inv_2 \inv[126]/_0_  (.Y(\inv_in[127] ),
    .A(\inv_in[126] ));
 sg13g2_inv_2 \inv[1270]/_0_  (.Y(\inv_in[1271] ),
    .A(\inv_in[1270] ));
 sg13g2_inv_2 \inv[1271]/_0_  (.Y(\inv_in[1272] ),
    .A(\inv_in[1271] ));
 sg13g2_inv_2 \inv[1272]/_0_  (.Y(\inv_in[1273] ),
    .A(\inv_in[1272] ));
 sg13g2_inv_2 \inv[1273]/_0_  (.Y(\inv_in[1274] ),
    .A(\inv_in[1273] ));
 sg13g2_inv_2 \inv[1274]/_0_  (.Y(\inv_in[1275] ),
    .A(\inv_in[1274] ));
 sg13g2_inv_2 \inv[1275]/_0_  (.Y(\inv_in[1276] ),
    .A(\inv_in[1275] ));
 sg13g2_inv_2 \inv[1276]/_0_  (.Y(\inv_in[1277] ),
    .A(\inv_in[1276] ));
 sg13g2_inv_2 \inv[1277]/_0_  (.Y(\inv_in[1278] ),
    .A(\inv_in[1277] ));
 sg13g2_inv_2 \inv[1278]/_0_  (.Y(\inv_in[1279] ),
    .A(\inv_in[1278] ));
 sg13g2_inv_2 \inv[1279]/_0_  (.Y(\inv_in[1280] ),
    .A(\inv_in[1279] ));
 sg13g2_inv_2 \inv[127]/_0_  (.Y(\inv_in[128] ),
    .A(\inv_in[127] ));
 sg13g2_inv_2 \inv[1280]/_0_  (.Y(\inv_in[1281] ),
    .A(\inv_in[1280] ));
 sg13g2_inv_2 \inv[1281]/_0_  (.Y(\inv_in[1282] ),
    .A(\inv_in[1281] ));
 sg13g2_inv_2 \inv[1282]/_0_  (.Y(\inv_in[1283] ),
    .A(\inv_in[1282] ));
 sg13g2_inv_2 \inv[1283]/_0_  (.Y(\inv_in[1284] ),
    .A(\inv_in[1283] ));
 sg13g2_inv_2 \inv[1284]/_0_  (.Y(\inv_in[1285] ),
    .A(\inv_in[1284] ));
 sg13g2_inv_2 \inv[1285]/_0_  (.Y(\inv_in[1286] ),
    .A(\inv_in[1285] ));
 sg13g2_inv_2 \inv[1286]/_0_  (.Y(\inv_in[1287] ),
    .A(\inv_in[1286] ));
 sg13g2_inv_2 \inv[1287]/_0_  (.Y(\inv_in[1288] ),
    .A(\inv_in[1287] ));
 sg13g2_inv_2 \inv[1288]/_0_  (.Y(\inv_in[1289] ),
    .A(\inv_in[1288] ));
 sg13g2_inv_2 \inv[1289]/_0_  (.Y(\inv_in[1290] ),
    .A(\inv_in[1289] ));
 sg13g2_inv_2 \inv[128]/_0_  (.Y(\inv_in[129] ),
    .A(\inv_in[128] ));
 sg13g2_inv_2 \inv[1290]/_0_  (.Y(\inv_in[1291] ),
    .A(\inv_in[1290] ));
 sg13g2_inv_2 \inv[1291]/_0_  (.Y(\inv_in[1292] ),
    .A(\inv_in[1291] ));
 sg13g2_inv_2 \inv[1292]/_0_  (.Y(\inv_in[1293] ),
    .A(\inv_in[1292] ));
 sg13g2_inv_2 \inv[1293]/_0_  (.Y(\inv_in[1294] ),
    .A(\inv_in[1293] ));
 sg13g2_inv_2 \inv[1294]/_0_  (.Y(\inv_in[1295] ),
    .A(\inv_in[1294] ));
 sg13g2_inv_2 \inv[1295]/_0_  (.Y(\inv_in[1296] ),
    .A(\inv_in[1295] ));
 sg13g2_inv_2 \inv[1296]/_0_  (.Y(\inv_in[1297] ),
    .A(\inv_in[1296] ));
 sg13g2_inv_2 \inv[1297]/_0_  (.Y(\inv_in[1298] ),
    .A(\inv_in[1297] ));
 sg13g2_inv_2 \inv[1298]/_0_  (.Y(\inv_in[1299] ),
    .A(\inv_in[1298] ));
 sg13g2_inv_2 \inv[1299]/_0_  (.Y(\inv_in[1300] ),
    .A(\inv_in[1299] ));
 sg13g2_inv_2 \inv[129]/_0_  (.Y(\inv_in[130] ),
    .A(\inv_in[129] ));
 sg13g2_inv_2 \inv[12]/_0_  (.Y(\inv_in[13] ),
    .A(\inv_in[12] ));
 sg13g2_inv_2 \inv[1300]/_0_  (.Y(\inv_in[1301] ),
    .A(\inv_in[1300] ));
 sg13g2_inv_2 \inv[1301]/_0_  (.Y(\inv_in[1302] ),
    .A(\inv_in[1301] ));
 sg13g2_inv_2 \inv[1302]/_0_  (.Y(\inv_in[1303] ),
    .A(\inv_in[1302] ));
 sg13g2_inv_2 \inv[1303]/_0_  (.Y(\inv_in[1304] ),
    .A(\inv_in[1303] ));
 sg13g2_inv_2 \inv[1304]/_0_  (.Y(\inv_in[1305] ),
    .A(\inv_in[1304] ));
 sg13g2_inv_2 \inv[1305]/_0_  (.Y(\inv_in[1306] ),
    .A(\inv_in[1305] ));
 sg13g2_inv_2 \inv[1306]/_0_  (.Y(\inv_in[1307] ),
    .A(\inv_in[1306] ));
 sg13g2_inv_2 \inv[1307]/_0_  (.Y(\inv_in[1308] ),
    .A(\inv_in[1307] ));
 sg13g2_inv_2 \inv[1308]/_0_  (.Y(\inv_in[1309] ),
    .A(\inv_in[1308] ));
 sg13g2_inv_2 \inv[1309]/_0_  (.Y(\inv_in[1310] ),
    .A(\inv_in[1309] ));
 sg13g2_inv_2 \inv[130]/_0_  (.Y(\inv_in[131] ),
    .A(\inv_in[130] ));
 sg13g2_inv_2 \inv[1310]/_0_  (.Y(\inv_in[1311] ),
    .A(\inv_in[1310] ));
 sg13g2_inv_2 \inv[1311]/_0_  (.Y(\inv_in[1312] ),
    .A(\inv_in[1311] ));
 sg13g2_inv_2 \inv[1312]/_0_  (.Y(\inv_in[1313] ),
    .A(\inv_in[1312] ));
 sg13g2_inv_2 \inv[1313]/_0_  (.Y(\inv_in[1314] ),
    .A(\inv_in[1313] ));
 sg13g2_inv_2 \inv[1314]/_0_  (.Y(\inv_in[1315] ),
    .A(\inv_in[1314] ));
 sg13g2_inv_2 \inv[1315]/_0_  (.Y(\inv_in[1316] ),
    .A(\inv_in[1315] ));
 sg13g2_inv_2 \inv[1316]/_0_  (.Y(\inv_in[1317] ),
    .A(\inv_in[1316] ));
 sg13g2_inv_4 \inv[1317]/_0_  (.A(\inv_in[1317] ),
    .Y(\inv_in[1318] ));
 sg13g2_inv_4 \inv[1318]/_0_  (.A(\inv_in[1318] ),
    .Y(\inv_in[1319] ));
 sg13g2_inv_4 \inv[1319]/_0_  (.A(\inv_in[1319] ),
    .Y(\inv_in[1320] ));
 sg13g2_inv_2 \inv[131]/_0_  (.Y(\inv_in[132] ),
    .A(\inv_in[131] ));
 sg13g2_inv_4 \inv[1320]/_0_  (.A(\inv_in[1320] ),
    .Y(\inv_in[1321] ));
 sg13g2_inv_4 \inv[1321]/_0_  (.A(\inv_in[1321] ),
    .Y(\inv_in[1322] ));
 sg13g2_inv_4 \inv[1322]/_0_  (.A(\inv_in[1322] ),
    .Y(\inv_in[1323] ));
 sg13g2_inv_4 \inv[1323]/_0_  (.A(\inv_in[1323] ),
    .Y(\inv_in[1324] ));
 sg13g2_inv_4 \inv[1324]/_0_  (.A(\inv_in[1324] ),
    .Y(\inv_in[1325] ));
 sg13g2_inv_4 \inv[1325]/_0_  (.A(\inv_in[1325] ),
    .Y(\inv_in[1326] ));
 sg13g2_inv_4 \inv[1326]/_0_  (.A(\inv_in[1326] ),
    .Y(\inv_in[1327] ));
 sg13g2_inv_4 \inv[1327]/_0_  (.A(\inv_in[1327] ),
    .Y(\inv_in[1328] ));
 sg13g2_inv_4 \inv[1328]/_0_  (.A(\inv_in[1328] ),
    .Y(\inv_in[1329] ));
 sg13g2_inv_2 \inv[1329]/_0_  (.Y(\inv_in[1330] ),
    .A(\inv_in[1329] ));
 sg13g2_inv_2 \inv[132]/_0_  (.Y(\inv_in[133] ),
    .A(\inv_in[132] ));
 sg13g2_inv_2 \inv[1330]/_0_  (.Y(\inv_in[1331] ),
    .A(\inv_in[1330] ));
 sg13g2_inv_4 \inv[1331]/_0_  (.A(\inv_in[1331] ),
    .Y(\inv_in[1332] ));
 sg13g2_inv_4 \inv[1332]/_0_  (.A(\inv_in[1332] ),
    .Y(\inv_in[1333] ));
 sg13g2_inv_4 \inv[1333]/_0_  (.A(\inv_in[1333] ),
    .Y(\inv_in[1334] ));
 sg13g2_inv_4 \inv[1334]/_0_  (.A(\inv_in[1334] ),
    .Y(\inv_in[1335] ));
 sg13g2_inv_4 \inv[1335]/_0_  (.A(\inv_in[1335] ),
    .Y(\inv_in[1336] ));
 sg13g2_inv_4 \inv[1336]/_0_  (.A(\inv_in[1336] ),
    .Y(\inv_in[1337] ));
 sg13g2_inv_2 \inv[1337]/_0_  (.Y(\inv_in[1338] ),
    .A(\inv_in[1337] ));
 sg13g2_inv_2 \inv[1338]/_0_  (.Y(\inv_in[1339] ),
    .A(\inv_in[1338] ));
 sg13g2_inv_2 \inv[1339]/_0_  (.Y(\inv_in[1340] ),
    .A(\inv_in[1339] ));
 sg13g2_inv_2 \inv[133]/_0_  (.Y(\inv_in[134] ),
    .A(\inv_in[133] ));
 sg13g2_inv_2 \inv[1340]/_0_  (.Y(\inv_in[1341] ),
    .A(\inv_in[1340] ));
 sg13g2_inv_2 \inv[1341]/_0_  (.Y(\inv_in[1342] ),
    .A(\inv_in[1341] ));
 sg13g2_inv_2 \inv[1342]/_0_  (.Y(\inv_in[1343] ),
    .A(\inv_in[1342] ));
 sg13g2_inv_2 \inv[1343]/_0_  (.Y(\inv_in[1344] ),
    .A(\inv_in[1343] ));
 sg13g2_inv_2 \inv[1344]/_0_  (.Y(\inv_in[1345] ),
    .A(\inv_in[1344] ));
 sg13g2_inv_2 \inv[1345]/_0_  (.Y(\inv_in[1346] ),
    .A(\inv_in[1345] ));
 sg13g2_inv_2 \inv[1346]/_0_  (.Y(\inv_in[1347] ),
    .A(\inv_in[1346] ));
 sg13g2_inv_2 \inv[1347]/_0_  (.Y(\inv_in[1348] ),
    .A(\inv_in[1347] ));
 sg13g2_inv_2 \inv[1348]/_0_  (.Y(\inv_in[1349] ),
    .A(\inv_in[1348] ));
 sg13g2_inv_2 \inv[1349]/_0_  (.Y(\inv_in[1350] ),
    .A(\inv_in[1349] ));
 sg13g2_inv_2 \inv[134]/_0_  (.Y(\inv_in[135] ),
    .A(\inv_in[134] ));
 sg13g2_inv_2 \inv[1350]/_0_  (.Y(\inv_in[1351] ),
    .A(\inv_in[1350] ));
 sg13g2_inv_2 \inv[1351]/_0_  (.Y(\inv_in[1352] ),
    .A(\inv_in[1351] ));
 sg13g2_inv_2 \inv[1352]/_0_  (.Y(\inv_in[1353] ),
    .A(\inv_in[1352] ));
 sg13g2_inv_2 \inv[1353]/_0_  (.Y(\inv_in[1354] ),
    .A(\inv_in[1353] ));
 sg13g2_inv_2 \inv[1354]/_0_  (.Y(\inv_in[1355] ),
    .A(\inv_in[1354] ));
 sg13g2_inv_2 \inv[1355]/_0_  (.Y(\inv_in[1356] ),
    .A(\inv_in[1355] ));
 sg13g2_inv_2 \inv[1356]/_0_  (.Y(\inv_in[1357] ),
    .A(\inv_in[1356] ));
 sg13g2_inv_2 \inv[1357]/_0_  (.Y(\inv_in[1358] ),
    .A(\inv_in[1357] ));
 sg13g2_inv_2 \inv[1358]/_0_  (.Y(\inv_in[1359] ),
    .A(\inv_in[1358] ));
 sg13g2_inv_2 \inv[1359]/_0_  (.Y(\inv_in[1360] ),
    .A(\inv_in[1359] ));
 sg13g2_inv_2 \inv[135]/_0_  (.Y(\inv_in[136] ),
    .A(\inv_in[135] ));
 sg13g2_inv_2 \inv[1360]/_0_  (.Y(\inv_in[1361] ),
    .A(\inv_in[1360] ));
 sg13g2_inv_2 \inv[1361]/_0_  (.Y(\inv_in[1362] ),
    .A(\inv_in[1361] ));
 sg13g2_inv_2 \inv[1362]/_0_  (.Y(\inv_in[1363] ),
    .A(\inv_in[1362] ));
 sg13g2_inv_2 \inv[1363]/_0_  (.Y(\inv_in[1364] ),
    .A(\inv_in[1363] ));
 sg13g2_inv_2 \inv[1364]/_0_  (.Y(\inv_in[1365] ),
    .A(\inv_in[1364] ));
 sg13g2_inv_2 \inv[1365]/_0_  (.Y(\inv_in[1366] ),
    .A(\inv_in[1365] ));
 sg13g2_inv_2 \inv[1366]/_0_  (.Y(\inv_in[1367] ),
    .A(\inv_in[1366] ));
 sg13g2_inv_2 \inv[1367]/_0_  (.Y(\inv_in[1368] ),
    .A(\inv_in[1367] ));
 sg13g2_inv_2 \inv[1368]/_0_  (.Y(\inv_in[1369] ),
    .A(\inv_in[1368] ));
 sg13g2_inv_2 \inv[1369]/_0_  (.Y(\inv_in[1370] ),
    .A(\inv_in[1369] ));
 sg13g2_inv_2 \inv[136]/_0_  (.Y(\inv_in[137] ),
    .A(\inv_in[136] ));
 sg13g2_inv_2 \inv[1370]/_0_  (.Y(\inv_in[1371] ),
    .A(\inv_in[1370] ));
 sg13g2_inv_2 \inv[1371]/_0_  (.Y(\inv_in[1372] ),
    .A(\inv_in[1371] ));
 sg13g2_inv_2 \inv[1372]/_0_  (.Y(\inv_in[1373] ),
    .A(\inv_in[1372] ));
 sg13g2_inv_2 \inv[1373]/_0_  (.Y(\inv_in[1374] ),
    .A(\inv_in[1373] ));
 sg13g2_inv_2 \inv[1374]/_0_  (.Y(\inv_in[1375] ),
    .A(\inv_in[1374] ));
 sg13g2_inv_2 \inv[1375]/_0_  (.Y(\inv_in[1376] ),
    .A(\inv_in[1375] ));
 sg13g2_inv_4 \inv[1376]/_0_  (.A(\inv_in[1376] ),
    .Y(\inv_in[1377] ));
 sg13g2_inv_4 \inv[1377]/_0_  (.A(\inv_in[1377] ),
    .Y(\inv_in[1378] ));
 sg13g2_inv_4 \inv[1378]/_0_  (.A(\inv_in[1378] ),
    .Y(\inv_in[1379] ));
 sg13g2_inv_4 \inv[1379]/_0_  (.A(\inv_in[1379] ),
    .Y(\inv_in[1380] ));
 sg13g2_inv_2 \inv[137]/_0_  (.Y(\inv_in[138] ),
    .A(\inv_in[137] ));
 sg13g2_inv_4 \inv[1380]/_0_  (.A(\inv_in[1380] ),
    .Y(\inv_in[1381] ));
 sg13g2_inv_4 \inv[1381]/_0_  (.A(\inv_in[1381] ),
    .Y(\inv_in[1382] ));
 sg13g2_inv_4 \inv[1382]/_0_  (.A(\inv_in[1382] ),
    .Y(\inv_in[1383] ));
 sg13g2_inv_4 \inv[1383]/_0_  (.A(\inv_in[1383] ),
    .Y(\inv_in[1384] ));
 sg13g2_inv_4 \inv[1384]/_0_  (.A(\inv_in[1384] ),
    .Y(\inv_in[1385] ));
 sg13g2_inv_4 \inv[1385]/_0_  (.A(\inv_in[1385] ),
    .Y(\inv_in[1386] ));
 sg13g2_inv_4 \inv[1386]/_0_  (.A(\inv_in[1386] ),
    .Y(\inv_in[1387] ));
 sg13g2_inv_4 \inv[1387]/_0_  (.A(\inv_in[1387] ),
    .Y(\inv_in[1388] ));
 sg13g2_inv_2 \inv[1388]/_0_  (.Y(\inv_in[1389] ),
    .A(\inv_in[1388] ));
 sg13g2_inv_2 \inv[1389]/_0_  (.Y(\inv_in[1390] ),
    .A(\inv_in[1389] ));
 sg13g2_inv_2 \inv[138]/_0_  (.Y(\inv_in[139] ),
    .A(\inv_in[138] ));
 sg13g2_inv_2 \inv[1390]/_0_  (.Y(\inv_in[1391] ),
    .A(\inv_in[1390] ));
 sg13g2_inv_2 \inv[1391]/_0_  (.Y(\inv_in[1392] ),
    .A(\inv_in[1391] ));
 sg13g2_inv_2 \inv[1392]/_0_  (.Y(\inv_in[1393] ),
    .A(\inv_in[1392] ));
 sg13g2_inv_2 \inv[1393]/_0_  (.Y(\inv_in[1394] ),
    .A(\inv_in[1393] ));
 sg13g2_inv_2 \inv[1394]/_0_  (.Y(\inv_in[1395] ),
    .A(\inv_in[1394] ));
 sg13g2_inv_2 \inv[1395]/_0_  (.Y(\inv_in[1396] ),
    .A(\inv_in[1395] ));
 sg13g2_inv_2 \inv[1396]/_0_  (.Y(\inv_in[1397] ),
    .A(\inv_in[1396] ));
 sg13g2_inv_2 \inv[1397]/_0_  (.Y(\inv_in[1398] ),
    .A(\inv_in[1397] ));
 sg13g2_inv_2 \inv[1398]/_0_  (.Y(\inv_in[1399] ),
    .A(\inv_in[1398] ));
 sg13g2_inv_2 \inv[1399]/_0_  (.Y(\inv_in[1400] ),
    .A(\inv_in[1399] ));
 sg13g2_inv_2 \inv[139]/_0_  (.Y(\inv_in[140] ),
    .A(\inv_in[139] ));
 sg13g2_inv_2 \inv[13]/_0_  (.Y(\inv_in[14] ),
    .A(\inv_in[13] ));
 sg13g2_inv_2 \inv[1400]/_0_  (.Y(\inv_in[1401] ),
    .A(\inv_in[1400] ));
 sg13g2_inv_2 \inv[1401]/_0_  (.Y(\inv_in[1402] ),
    .A(\inv_in[1401] ));
 sg13g2_inv_2 \inv[1402]/_0_  (.Y(\inv_in[1403] ),
    .A(\inv_in[1402] ));
 sg13g2_inv_2 \inv[1403]/_0_  (.Y(\inv_in[1404] ),
    .A(\inv_in[1403] ));
 sg13g2_inv_2 \inv[1404]/_0_  (.Y(\inv_in[1405] ),
    .A(\inv_in[1404] ));
 sg13g2_inv_2 \inv[1405]/_0_  (.Y(\inv_in[1406] ),
    .A(\inv_in[1405] ));
 sg13g2_inv_2 \inv[1406]/_0_  (.Y(\inv_in[1407] ),
    .A(\inv_in[1406] ));
 sg13g2_inv_2 \inv[1407]/_0_  (.Y(\inv_in[1408] ),
    .A(\inv_in[1407] ));
 sg13g2_inv_2 \inv[1408]/_0_  (.Y(\inv_in[1409] ),
    .A(\inv_in[1408] ));
 sg13g2_inv_2 \inv[1409]/_0_  (.Y(\inv_in[1410] ),
    .A(\inv_in[1409] ));
 sg13g2_inv_2 \inv[140]/_0_  (.Y(\inv_in[141] ),
    .A(\inv_in[140] ));
 sg13g2_inv_2 \inv[1410]/_0_  (.Y(\inv_in[1411] ),
    .A(\inv_in[1410] ));
 sg13g2_inv_2 \inv[1411]/_0_  (.Y(\inv_in[1412] ),
    .A(\inv_in[1411] ));
 sg13g2_inv_2 \inv[1412]/_0_  (.Y(\inv_in[1413] ),
    .A(\inv_in[1412] ));
 sg13g2_inv_2 \inv[1413]/_0_  (.Y(\inv_in[1414] ),
    .A(\inv_in[1413] ));
 sg13g2_inv_2 \inv[1414]/_0_  (.Y(\inv_in[1415] ),
    .A(\inv_in[1414] ));
 sg13g2_inv_2 \inv[1415]/_0_  (.Y(\inv_in[1416] ),
    .A(\inv_in[1415] ));
 sg13g2_inv_2 \inv[1416]/_0_  (.Y(\inv_in[1417] ),
    .A(\inv_in[1416] ));
 sg13g2_inv_2 \inv[1417]/_0_  (.Y(\inv_in[1418] ),
    .A(\inv_in[1417] ));
 sg13g2_inv_2 \inv[1418]/_0_  (.Y(\inv_in[1419] ),
    .A(\inv_in[1418] ));
 sg13g2_inv_2 \inv[1419]/_0_  (.Y(\inv_in[1420] ),
    .A(\inv_in[1419] ));
 sg13g2_inv_2 \inv[141]/_0_  (.Y(\inv_in[142] ),
    .A(\inv_in[141] ));
 sg13g2_inv_2 \inv[1420]/_0_  (.Y(\inv_in[1421] ),
    .A(\inv_in[1420] ));
 sg13g2_inv_2 \inv[1421]/_0_  (.Y(\inv_in[1422] ),
    .A(\inv_in[1421] ));
 sg13g2_inv_2 \inv[1422]/_0_  (.Y(\inv_in[1423] ),
    .A(\inv_in[1422] ));
 sg13g2_inv_2 \inv[1423]/_0_  (.Y(\inv_in[1424] ),
    .A(\inv_in[1423] ));
 sg13g2_inv_2 \inv[1424]/_0_  (.Y(\inv_in[1425] ),
    .A(\inv_in[1424] ));
 sg13g2_inv_2 \inv[1425]/_0_  (.Y(\inv_in[1426] ),
    .A(\inv_in[1425] ));
 sg13g2_inv_2 \inv[1426]/_0_  (.Y(\inv_in[1427] ),
    .A(\inv_in[1426] ));
 sg13g2_inv_2 \inv[1427]/_0_  (.Y(\inv_in[1428] ),
    .A(\inv_in[1427] ));
 sg13g2_inv_2 \inv[1428]/_0_  (.Y(\inv_in[1429] ),
    .A(\inv_in[1428] ));
 sg13g2_inv_2 \inv[1429]/_0_  (.Y(\inv_in[1430] ),
    .A(\inv_in[1429] ));
 sg13g2_inv_2 \inv[142]/_0_  (.Y(\inv_in[143] ),
    .A(\inv_in[142] ));
 sg13g2_inv_2 \inv[1430]/_0_  (.Y(\inv_in[1431] ),
    .A(\inv_in[1430] ));
 sg13g2_inv_2 \inv[1431]/_0_  (.Y(\inv_in[1432] ),
    .A(\inv_in[1431] ));
 sg13g2_inv_2 \inv[1432]/_0_  (.Y(\inv_in[1433] ),
    .A(\inv_in[1432] ));
 sg13g2_inv_2 \inv[1433]/_0_  (.Y(\inv_in[1434] ),
    .A(\inv_in[1433] ));
 sg13g2_inv_2 \inv[1434]/_0_  (.Y(\inv_in[1435] ),
    .A(\inv_in[1434] ));
 sg13g2_inv_2 \inv[1435]/_0_  (.Y(\inv_in[1436] ),
    .A(\inv_in[1435] ));
 sg13g2_inv_2 \inv[1436]/_0_  (.Y(\inv_in[1437] ),
    .A(\inv_in[1436] ));
 sg13g2_inv_2 \inv[1437]/_0_  (.Y(\inv_in[1438] ),
    .A(\inv_in[1437] ));
 sg13g2_inv_2 \inv[1438]/_0_  (.Y(\inv_in[1439] ),
    .A(\inv_in[1438] ));
 sg13g2_inv_2 \inv[1439]/_0_  (.Y(\inv_in[1440] ),
    .A(\inv_in[1439] ));
 sg13g2_inv_2 \inv[143]/_0_  (.Y(\inv_in[144] ),
    .A(\inv_in[143] ));
 sg13g2_inv_2 \inv[1440]/_0_  (.Y(\inv_in[1441] ),
    .A(\inv_in[1440] ));
 sg13g2_inv_2 \inv[1441]/_0_  (.Y(\inv_in[1442] ),
    .A(\inv_in[1441] ));
 sg13g2_inv_2 \inv[1442]/_0_  (.Y(\inv_in[1443] ),
    .A(\inv_in[1442] ));
 sg13g2_inv_2 \inv[1443]/_0_  (.Y(\inv_in[1444] ),
    .A(\inv_in[1443] ));
 sg13g2_inv_2 \inv[1444]/_0_  (.Y(\inv_in[1445] ),
    .A(\inv_in[1444] ));
 sg13g2_inv_2 \inv[1445]/_0_  (.Y(\inv_in[1446] ),
    .A(\inv_in[1445] ));
 sg13g2_inv_2 \inv[1446]/_0_  (.Y(\inv_in[1447] ),
    .A(\inv_in[1446] ));
 sg13g2_inv_2 \inv[1447]/_0_  (.Y(\inv_in[1448] ),
    .A(\inv_in[1447] ));
 sg13g2_inv_2 \inv[1448]/_0_  (.Y(\inv_in[1449] ),
    .A(\inv_in[1448] ));
 sg13g2_inv_2 \inv[1449]/_0_  (.Y(\inv_in[1450] ),
    .A(\inv_in[1449] ));
 sg13g2_inv_2 \inv[144]/_0_  (.Y(\inv_in[145] ),
    .A(\inv_in[144] ));
 sg13g2_inv_2 \inv[1450]/_0_  (.Y(\inv_in[1451] ),
    .A(\inv_in[1450] ));
 sg13g2_inv_2 \inv[1451]/_0_  (.Y(\inv_in[1452] ),
    .A(\inv_in[1451] ));
 sg13g2_inv_2 \inv[1452]/_0_  (.Y(\inv_in[1453] ),
    .A(\inv_in[1452] ));
 sg13g2_inv_2 \inv[1453]/_0_  (.Y(\inv_in[1454] ),
    .A(\inv_in[1453] ));
 sg13g2_inv_2 \inv[1454]/_0_  (.Y(\inv_in[1455] ),
    .A(\inv_in[1454] ));
 sg13g2_inv_2 \inv[1455]/_0_  (.Y(\inv_in[1456] ),
    .A(\inv_in[1455] ));
 sg13g2_inv_2 \inv[1456]/_0_  (.Y(\inv_in[1457] ),
    .A(\inv_in[1456] ));
 sg13g2_inv_2 \inv[1457]/_0_  (.Y(\inv_in[1458] ),
    .A(\inv_in[1457] ));
 sg13g2_inv_2 \inv[1458]/_0_  (.Y(\inv_in[1459] ),
    .A(\inv_in[1458] ));
 sg13g2_inv_2 \inv[1459]/_0_  (.Y(\inv_in[1460] ),
    .A(\inv_in[1459] ));
 sg13g2_inv_2 \inv[145]/_0_  (.Y(\inv_in[146] ),
    .A(\inv_in[145] ));
 sg13g2_inv_2 \inv[1460]/_0_  (.Y(\inv_in[1461] ),
    .A(\inv_in[1460] ));
 sg13g2_inv_2 \inv[1461]/_0_  (.Y(\inv_in[1462] ),
    .A(\inv_in[1461] ));
 sg13g2_inv_2 \inv[1462]/_0_  (.Y(\inv_in[1463] ),
    .A(\inv_in[1462] ));
 sg13g2_inv_2 \inv[1463]/_0_  (.Y(\inv_in[1464] ),
    .A(\inv_in[1463] ));
 sg13g2_inv_2 \inv[1464]/_0_  (.Y(\inv_in[1465] ),
    .A(\inv_in[1464] ));
 sg13g2_inv_2 \inv[1465]/_0_  (.Y(\inv_in[1466] ),
    .A(\inv_in[1465] ));
 sg13g2_inv_2 \inv[1466]/_0_  (.Y(\inv_in[1467] ),
    .A(\inv_in[1466] ));
 sg13g2_inv_2 \inv[1467]/_0_  (.Y(\inv_in[1468] ),
    .A(\inv_in[1467] ));
 sg13g2_inv_2 \inv[1468]/_0_  (.Y(\inv_in[1469] ),
    .A(\inv_in[1468] ));
 sg13g2_inv_2 \inv[1469]/_0_  (.Y(\inv_in[1470] ),
    .A(\inv_in[1469] ));
 sg13g2_inv_2 \inv[146]/_0_  (.Y(\inv_in[147] ),
    .A(\inv_in[146] ));
 sg13g2_inv_2 \inv[1470]/_0_  (.Y(\inv_in[1471] ),
    .A(\inv_in[1470] ));
 sg13g2_inv_2 \inv[1471]/_0_  (.Y(\inv_in[1472] ),
    .A(\inv_in[1471] ));
 sg13g2_inv_2 \inv[1472]/_0_  (.Y(\inv_in[1473] ),
    .A(\inv_in[1472] ));
 sg13g2_inv_2 \inv[1473]/_0_  (.Y(\inv_in[1474] ),
    .A(\inv_in[1473] ));
 sg13g2_inv_2 \inv[1474]/_0_  (.Y(\inv_in[1475] ),
    .A(\inv_in[1474] ));
 sg13g2_inv_2 \inv[1475]/_0_  (.Y(\inv_in[1476] ),
    .A(\inv_in[1475] ));
 sg13g2_inv_2 \inv[1476]/_0_  (.Y(\inv_in[1477] ),
    .A(\inv_in[1476] ));
 sg13g2_inv_2 \inv[1477]/_0_  (.Y(\inv_in[1478] ),
    .A(\inv_in[1477] ));
 sg13g2_inv_2 \inv[1478]/_0_  (.Y(\inv_in[1479] ),
    .A(\inv_in[1478] ));
 sg13g2_inv_2 \inv[1479]/_0_  (.Y(\inv_in[1480] ),
    .A(\inv_in[1479] ));
 sg13g2_inv_2 \inv[147]/_0_  (.Y(\inv_in[148] ),
    .A(\inv_in[147] ));
 sg13g2_inv_2 \inv[1480]/_0_  (.Y(\inv_in[1481] ),
    .A(\inv_in[1480] ));
 sg13g2_inv_2 \inv[1481]/_0_  (.Y(\inv_in[1482] ),
    .A(\inv_in[1481] ));
 sg13g2_inv_2 \inv[1482]/_0_  (.Y(\inv_in[1483] ),
    .A(\inv_in[1482] ));
 sg13g2_inv_2 \inv[1483]/_0_  (.Y(\inv_in[1484] ),
    .A(\inv_in[1483] ));
 sg13g2_inv_2 \inv[1484]/_0_  (.Y(\inv_in[1485] ),
    .A(\inv_in[1484] ));
 sg13g2_inv_2 \inv[1485]/_0_  (.Y(\inv_in[1486] ),
    .A(\inv_in[1485] ));
 sg13g2_inv_2 \inv[1486]/_0_  (.Y(\inv_in[1487] ),
    .A(\inv_in[1486] ));
 sg13g2_inv_2 \inv[1487]/_0_  (.Y(\inv_in[1488] ),
    .A(\inv_in[1487] ));
 sg13g2_inv_2 \inv[1488]/_0_  (.Y(\inv_in[1489] ),
    .A(\inv_in[1488] ));
 sg13g2_inv_2 \inv[1489]/_0_  (.Y(\inv_in[1490] ),
    .A(\inv_in[1489] ));
 sg13g2_inv_2 \inv[148]/_0_  (.Y(\inv_in[149] ),
    .A(\inv_in[148] ));
 sg13g2_inv_2 \inv[1490]/_0_  (.Y(\inv_in[1491] ),
    .A(\inv_in[1490] ));
 sg13g2_inv_2 \inv[1491]/_0_  (.Y(\inv_in[1492] ),
    .A(\inv_in[1491] ));
 sg13g2_inv_2 \inv[1492]/_0_  (.Y(\inv_in[1493] ),
    .A(\inv_in[1492] ));
 sg13g2_inv_2 \inv[1493]/_0_  (.Y(\inv_in[1494] ),
    .A(\inv_in[1493] ));
 sg13g2_inv_2 \inv[1494]/_0_  (.Y(\inv_in[1495] ),
    .A(\inv_in[1494] ));
 sg13g2_inv_2 \inv[1495]/_0_  (.Y(\inv_in[1496] ),
    .A(\inv_in[1495] ));
 sg13g2_inv_2 \inv[1496]/_0_  (.Y(\inv_in[1497] ),
    .A(\inv_in[1496] ));
 sg13g2_inv_2 \inv[1497]/_0_  (.Y(\inv_in[1498] ),
    .A(\inv_in[1497] ));
 sg13g2_inv_2 \inv[1498]/_0_  (.Y(\inv_in[1499] ),
    .A(\inv_in[1498] ));
 sg13g2_inv_2 \inv[1499]/_0_  (.Y(\inv_in[1500] ),
    .A(\inv_in[1499] ));
 sg13g2_inv_2 \inv[149]/_0_  (.Y(\inv_in[150] ),
    .A(\inv_in[149] ));
 sg13g2_inv_2 \inv[14]/_0_  (.Y(\inv_in[15] ),
    .A(\inv_in[14] ));
 sg13g2_inv_2 \inv[1500]/_0_  (.Y(\inv_in[1501] ),
    .A(\inv_in[1500] ));
 sg13g2_inv_2 \inv[1501]/_0_  (.Y(\inv_in[1502] ),
    .A(\inv_in[1501] ));
 sg13g2_inv_2 \inv[1502]/_0_  (.Y(\inv_in[1503] ),
    .A(\inv_in[1502] ));
 sg13g2_inv_2 \inv[1503]/_0_  (.Y(\inv_in[1504] ),
    .A(\inv_in[1503] ));
 sg13g2_inv_2 \inv[1504]/_0_  (.Y(\inv_in[1505] ),
    .A(\inv_in[1504] ));
 sg13g2_inv_2 \inv[1505]/_0_  (.Y(\inv_in[1506] ),
    .A(\inv_in[1505] ));
 sg13g2_inv_2 \inv[1506]/_0_  (.Y(\inv_in[1507] ),
    .A(\inv_in[1506] ));
 sg13g2_inv_2 \inv[1507]/_0_  (.Y(\inv_in[1508] ),
    .A(\inv_in[1507] ));
 sg13g2_inv_2 \inv[1508]/_0_  (.Y(\inv_in[1509] ),
    .A(\inv_in[1508] ));
 sg13g2_inv_2 \inv[1509]/_0_  (.Y(\inv_in[1510] ),
    .A(\inv_in[1509] ));
 sg13g2_inv_2 \inv[150]/_0_  (.Y(\inv_in[151] ),
    .A(\inv_in[150] ));
 sg13g2_inv_2 \inv[1510]/_0_  (.Y(\inv_in[1511] ),
    .A(\inv_in[1510] ));
 sg13g2_inv_2 \inv[1511]/_0_  (.Y(\inv_in[1512] ),
    .A(\inv_in[1511] ));
 sg13g2_inv_2 \inv[1512]/_0_  (.Y(\inv_in[1513] ),
    .A(\inv_in[1512] ));
 sg13g2_inv_2 \inv[1513]/_0_  (.Y(\inv_in[1514] ),
    .A(\inv_in[1513] ));
 sg13g2_inv_2 \inv[1514]/_0_  (.Y(\inv_in[1515] ),
    .A(\inv_in[1514] ));
 sg13g2_inv_2 \inv[1515]/_0_  (.Y(\inv_in[1516] ),
    .A(\inv_in[1515] ));
 sg13g2_inv_2 \inv[1516]/_0_  (.Y(\inv_in[1517] ),
    .A(\inv_in[1516] ));
 sg13g2_inv_2 \inv[1517]/_0_  (.Y(\inv_in[1518] ),
    .A(\inv_in[1517] ));
 sg13g2_inv_2 \inv[1518]/_0_  (.Y(\inv_in[1519] ),
    .A(\inv_in[1518] ));
 sg13g2_inv_2 \inv[1519]/_0_  (.Y(\inv_in[1520] ),
    .A(\inv_in[1519] ));
 sg13g2_inv_2 \inv[151]/_0_  (.Y(\inv_in[152] ),
    .A(\inv_in[151] ));
 sg13g2_inv_2 \inv[1520]/_0_  (.Y(\inv_in[1521] ),
    .A(\inv_in[1520] ));
 sg13g2_inv_2 \inv[1521]/_0_  (.Y(\inv_in[1522] ),
    .A(\inv_in[1521] ));
 sg13g2_inv_2 \inv[1522]/_0_  (.Y(\inv_in[1523] ),
    .A(\inv_in[1522] ));
 sg13g2_inv_2 \inv[1523]/_0_  (.Y(\inv_in[1524] ),
    .A(\inv_in[1523] ));
 sg13g2_inv_2 \inv[1524]/_0_  (.Y(\inv_in[1525] ),
    .A(\inv_in[1524] ));
 sg13g2_inv_2 \inv[1525]/_0_  (.Y(\inv_in[1526] ),
    .A(\inv_in[1525] ));
 sg13g2_inv_2 \inv[1526]/_0_  (.Y(\inv_in[1527] ),
    .A(\inv_in[1526] ));
 sg13g2_inv_2 \inv[1527]/_0_  (.Y(\inv_in[1528] ),
    .A(\inv_in[1527] ));
 sg13g2_inv_2 \inv[1528]/_0_  (.Y(\inv_in[1529] ),
    .A(\inv_in[1528] ));
 sg13g2_inv_2 \inv[1529]/_0_  (.Y(\inv_in[1530] ),
    .A(\inv_in[1529] ));
 sg13g2_inv_2 \inv[152]/_0_  (.Y(\inv_in[153] ),
    .A(\inv_in[152] ));
 sg13g2_inv_2 \inv[1530]/_0_  (.Y(\inv_in[1531] ),
    .A(\inv_in[1530] ));
 sg13g2_inv_2 \inv[1531]/_0_  (.Y(\inv_in[1532] ),
    .A(\inv_in[1531] ));
 sg13g2_inv_2 \inv[1532]/_0_  (.Y(\inv_in[1533] ),
    .A(\inv_in[1532] ));
 sg13g2_inv_2 \inv[1533]/_0_  (.Y(\inv_in[1534] ),
    .A(\inv_in[1533] ));
 sg13g2_inv_2 \inv[1534]/_0_  (.Y(\inv_in[1535] ),
    .A(\inv_in[1534] ));
 sg13g2_inv_2 \inv[1535]/_0_  (.Y(\inv_in[1536] ),
    .A(\inv_in[1535] ));
 sg13g2_inv_2 \inv[1536]/_0_  (.Y(\inv_in[1537] ),
    .A(\inv_in[1536] ));
 sg13g2_inv_2 \inv[1537]/_0_  (.Y(\inv_in[1538] ),
    .A(\inv_in[1537] ));
 sg13g2_inv_2 \inv[1538]/_0_  (.Y(\inv_in[1539] ),
    .A(\inv_in[1538] ));
 sg13g2_inv_2 \inv[1539]/_0_  (.Y(\inv_in[1540] ),
    .A(\inv_in[1539] ));
 sg13g2_inv_2 \inv[153]/_0_  (.Y(\inv_in[154] ),
    .A(\inv_in[153] ));
 sg13g2_inv_2 \inv[1540]/_0_  (.Y(\inv_in[1541] ),
    .A(\inv_in[1540] ));
 sg13g2_inv_2 \inv[1541]/_0_  (.Y(\inv_in[1542] ),
    .A(\inv_in[1541] ));
 sg13g2_inv_2 \inv[1542]/_0_  (.Y(\inv_in[1543] ),
    .A(\inv_in[1542] ));
 sg13g2_inv_2 \inv[1543]/_0_  (.Y(\inv_in[1544] ),
    .A(\inv_in[1543] ));
 sg13g2_inv_2 \inv[1544]/_0_  (.Y(\inv_in[1545] ),
    .A(\inv_in[1544] ));
 sg13g2_inv_2 \inv[1545]/_0_  (.Y(\inv_in[1546] ),
    .A(\inv_in[1545] ));
 sg13g2_inv_2 \inv[1546]/_0_  (.Y(\inv_in[1547] ),
    .A(\inv_in[1546] ));
 sg13g2_inv_2 \inv[1547]/_0_  (.Y(\inv_in[1548] ),
    .A(\inv_in[1547] ));
 sg13g2_inv_2 \inv[1548]/_0_  (.Y(\inv_in[1549] ),
    .A(\inv_in[1548] ));
 sg13g2_inv_2 \inv[1549]/_0_  (.Y(\inv_in[1550] ),
    .A(\inv_in[1549] ));
 sg13g2_inv_2 \inv[154]/_0_  (.Y(\inv_in[155] ),
    .A(\inv_in[154] ));
 sg13g2_inv_2 \inv[1550]/_0_  (.Y(\inv_in[1551] ),
    .A(\inv_in[1550] ));
 sg13g2_inv_2 \inv[1551]/_0_  (.Y(\inv_in[1552] ),
    .A(\inv_in[1551] ));
 sg13g2_inv_2 \inv[1552]/_0_  (.Y(\inv_in[1553] ),
    .A(\inv_in[1552] ));
 sg13g2_inv_2 \inv[1553]/_0_  (.Y(\inv_in[1554] ),
    .A(\inv_in[1553] ));
 sg13g2_inv_2 \inv[1554]/_0_  (.Y(\inv_in[1555] ),
    .A(\inv_in[1554] ));
 sg13g2_inv_2 \inv[1555]/_0_  (.Y(\inv_in[1556] ),
    .A(\inv_in[1555] ));
 sg13g2_inv_2 \inv[1556]/_0_  (.Y(\inv_in[1557] ),
    .A(\inv_in[1556] ));
 sg13g2_inv_2 \inv[1557]/_0_  (.Y(\inv_in[1558] ),
    .A(\inv_in[1557] ));
 sg13g2_inv_2 \inv[1558]/_0_  (.Y(\inv_in[1559] ),
    .A(\inv_in[1558] ));
 sg13g2_inv_2 \inv[1559]/_0_  (.Y(\inv_in[1560] ),
    .A(\inv_in[1559] ));
 sg13g2_inv_2 \inv[155]/_0_  (.Y(\inv_in[156] ),
    .A(\inv_in[155] ));
 sg13g2_inv_2 \inv[1560]/_0_  (.Y(\inv_in[1561] ),
    .A(\inv_in[1560] ));
 sg13g2_inv_2 \inv[1561]/_0_  (.Y(\inv_in[1562] ),
    .A(\inv_in[1561] ));
 sg13g2_inv_2 \inv[1562]/_0_  (.Y(\inv_in[1563] ),
    .A(\inv_in[1562] ));
 sg13g2_inv_2 \inv[1563]/_0_  (.Y(\inv_in[1564] ),
    .A(\inv_in[1563] ));
 sg13g2_inv_2 \inv[1564]/_0_  (.Y(\inv_in[1565] ),
    .A(\inv_in[1564] ));
 sg13g2_inv_2 \inv[1565]/_0_  (.Y(\inv_in[1566] ),
    .A(\inv_in[1565] ));
 sg13g2_inv_2 \inv[1566]/_0_  (.Y(\inv_in[1567] ),
    .A(\inv_in[1566] ));
 sg13g2_inv_2 \inv[1567]/_0_  (.Y(\inv_in[1568] ),
    .A(\inv_in[1567] ));
 sg13g2_inv_2 \inv[1568]/_0_  (.Y(\inv_in[1569] ),
    .A(\inv_in[1568] ));
 sg13g2_inv_2 \inv[1569]/_0_  (.Y(\inv_in[1570] ),
    .A(\inv_in[1569] ));
 sg13g2_inv_2 \inv[156]/_0_  (.Y(\inv_in[157] ),
    .A(\inv_in[156] ));
 sg13g2_inv_2 \inv[1570]/_0_  (.Y(\inv_in[1571] ),
    .A(\inv_in[1570] ));
 sg13g2_inv_2 \inv[1571]/_0_  (.Y(\inv_in[1572] ),
    .A(\inv_in[1571] ));
 sg13g2_inv_2 \inv[1572]/_0_  (.Y(\inv_in[1573] ),
    .A(\inv_in[1572] ));
 sg13g2_inv_2 \inv[1573]/_0_  (.Y(\inv_in[1574] ),
    .A(\inv_in[1573] ));
 sg13g2_inv_2 \inv[1574]/_0_  (.Y(\inv_in[1575] ),
    .A(\inv_in[1574] ));
 sg13g2_inv_2 \inv[1575]/_0_  (.Y(\inv_in[1576] ),
    .A(\inv_in[1575] ));
 sg13g2_inv_2 \inv[1576]/_0_  (.Y(\inv_in[1577] ),
    .A(\inv_in[1576] ));
 sg13g2_inv_2 \inv[1577]/_0_  (.Y(\inv_in[1578] ),
    .A(\inv_in[1577] ));
 sg13g2_inv_2 \inv[1578]/_0_  (.Y(\inv_in[1579] ),
    .A(\inv_in[1578] ));
 sg13g2_inv_2 \inv[1579]/_0_  (.Y(\inv_in[1580] ),
    .A(\inv_in[1579] ));
 sg13g2_inv_2 \inv[157]/_0_  (.Y(\inv_in[158] ),
    .A(\inv_in[157] ));
 sg13g2_inv_2 \inv[1580]/_0_  (.Y(\inv_in[1581] ),
    .A(\inv_in[1580] ));
 sg13g2_inv_2 \inv[1581]/_0_  (.Y(\inv_in[1582] ),
    .A(\inv_in[1581] ));
 sg13g2_inv_2 \inv[1582]/_0_  (.Y(\inv_in[1583] ),
    .A(\inv_in[1582] ));
 sg13g2_inv_2 \inv[1583]/_0_  (.Y(\inv_in[1584] ),
    .A(\inv_in[1583] ));
 sg13g2_inv_2 \inv[1584]/_0_  (.Y(\inv_in[1585] ),
    .A(\inv_in[1584] ));
 sg13g2_inv_2 \inv[1585]/_0_  (.Y(\inv_in[1586] ),
    .A(\inv_in[1585] ));
 sg13g2_inv_2 \inv[1586]/_0_  (.Y(\inv_in[1587] ),
    .A(\inv_in[1586] ));
 sg13g2_inv_2 \inv[1587]/_0_  (.Y(\inv_in[1588] ),
    .A(\inv_in[1587] ));
 sg13g2_inv_2 \inv[1588]/_0_  (.Y(\inv_in[1589] ),
    .A(\inv_in[1588] ));
 sg13g2_inv_2 \inv[1589]/_0_  (.Y(\inv_in[1590] ),
    .A(\inv_in[1589] ));
 sg13g2_inv_2 \inv[158]/_0_  (.Y(\inv_in[159] ),
    .A(\inv_in[158] ));
 sg13g2_inv_2 \inv[1590]/_0_  (.Y(\inv_in[1591] ),
    .A(\inv_in[1590] ));
 sg13g2_inv_2 \inv[1591]/_0_  (.Y(\inv_in[1592] ),
    .A(\inv_in[1591] ));
 sg13g2_inv_2 \inv[1592]/_0_  (.Y(\inv_in[1593] ),
    .A(\inv_in[1592] ));
 sg13g2_inv_2 \inv[1593]/_0_  (.Y(\inv_in[1594] ),
    .A(\inv_in[1593] ));
 sg13g2_inv_2 \inv[1594]/_0_  (.Y(\inv_in[1595] ),
    .A(\inv_in[1594] ));
 sg13g2_inv_2 \inv[1595]/_0_  (.Y(\inv_in[1596] ),
    .A(\inv_in[1595] ));
 sg13g2_inv_2 \inv[1596]/_0_  (.Y(\inv_in[1597] ),
    .A(\inv_in[1596] ));
 sg13g2_inv_2 \inv[1597]/_0_  (.Y(\inv_in[1598] ),
    .A(\inv_in[1597] ));
 sg13g2_inv_2 \inv[1598]/_0_  (.Y(\inv_in[1599] ),
    .A(\inv_in[1598] ));
 sg13g2_inv_2 \inv[1599]/_0_  (.Y(\inv_in[1600] ),
    .A(\inv_in[1599] ));
 sg13g2_inv_2 \inv[159]/_0_  (.Y(\inv_in[160] ),
    .A(\inv_in[159] ));
 sg13g2_inv_2 \inv[15]/_0_  (.Y(\inv_in[16] ),
    .A(\inv_in[15] ));
 sg13g2_inv_2 \inv[1600]/_0_  (.Y(\inv_in[1601] ),
    .A(\inv_in[1600] ));
 sg13g2_inv_2 \inv[1601]/_0_  (.Y(\inv_in[1602] ),
    .A(\inv_in[1601] ));
 sg13g2_inv_2 \inv[1602]/_0_  (.Y(\inv_in[1603] ),
    .A(\inv_in[1602] ));
 sg13g2_inv_2 \inv[1603]/_0_  (.Y(\inv_in[1604] ),
    .A(\inv_in[1603] ));
 sg13g2_inv_2 \inv[1604]/_0_  (.Y(\inv_in[1605] ),
    .A(\inv_in[1604] ));
 sg13g2_inv_2 \inv[1605]/_0_  (.Y(\inv_in[1606] ),
    .A(\inv_in[1605] ));
 sg13g2_inv_2 \inv[1606]/_0_  (.Y(\inv_in[1607] ),
    .A(\inv_in[1606] ));
 sg13g2_inv_2 \inv[1607]/_0_  (.Y(\inv_in[1608] ),
    .A(\inv_in[1607] ));
 sg13g2_inv_2 \inv[1608]/_0_  (.Y(\inv_in[1609] ),
    .A(\inv_in[1608] ));
 sg13g2_inv_2 \inv[1609]/_0_  (.Y(\inv_in[1610] ),
    .A(\inv_in[1609] ));
 sg13g2_inv_2 \inv[160]/_0_  (.Y(\inv_in[161] ),
    .A(\inv_in[160] ));
 sg13g2_inv_2 \inv[1610]/_0_  (.Y(\inv_in[1611] ),
    .A(\inv_in[1610] ));
 sg13g2_inv_2 \inv[1611]/_0_  (.Y(\inv_in[1612] ),
    .A(\inv_in[1611] ));
 sg13g2_inv_2 \inv[1612]/_0_  (.Y(\inv_in[1613] ),
    .A(\inv_in[1612] ));
 sg13g2_inv_2 \inv[1613]/_0_  (.Y(\inv_in[1614] ),
    .A(\inv_in[1613] ));
 sg13g2_inv_2 \inv[1614]/_0_  (.Y(\inv_in[1615] ),
    .A(\inv_in[1614] ));
 sg13g2_inv_2 \inv[1615]/_0_  (.Y(\inv_in[1616] ),
    .A(\inv_in[1615] ));
 sg13g2_inv_2 \inv[1616]/_0_  (.Y(\inv_in[1617] ),
    .A(\inv_in[1616] ));
 sg13g2_inv_2 \inv[1617]/_0_  (.Y(\inv_in[1618] ),
    .A(\inv_in[1617] ));
 sg13g2_inv_2 \inv[1618]/_0_  (.Y(\inv_in[1619] ),
    .A(\inv_in[1618] ));
 sg13g2_inv_2 \inv[1619]/_0_  (.Y(\inv_in[1620] ),
    .A(\inv_in[1619] ));
 sg13g2_inv_2 \inv[161]/_0_  (.Y(\inv_in[162] ),
    .A(\inv_in[161] ));
 sg13g2_inv_2 \inv[1620]/_0_  (.Y(\inv_in[1621] ),
    .A(\inv_in[1620] ));
 sg13g2_inv_2 \inv[1621]/_0_  (.Y(\inv_in[1622] ),
    .A(\inv_in[1621] ));
 sg13g2_inv_2 \inv[1622]/_0_  (.Y(\inv_in[1623] ),
    .A(\inv_in[1622] ));
 sg13g2_inv_2 \inv[1623]/_0_  (.Y(\inv_in[1624] ),
    .A(\inv_in[1623] ));
 sg13g2_inv_2 \inv[1624]/_0_  (.Y(\inv_in[1625] ),
    .A(\inv_in[1624] ));
 sg13g2_inv_2 \inv[1625]/_0_  (.Y(\inv_in[1626] ),
    .A(\inv_in[1625] ));
 sg13g2_inv_2 \inv[1626]/_0_  (.Y(\inv_in[1627] ),
    .A(\inv_in[1626] ));
 sg13g2_inv_2 \inv[1627]/_0_  (.Y(\inv_in[1628] ),
    .A(\inv_in[1627] ));
 sg13g2_inv_2 \inv[1628]/_0_  (.Y(\inv_in[1629] ),
    .A(\inv_in[1628] ));
 sg13g2_inv_2 \inv[1629]/_0_  (.Y(\inv_in[1630] ),
    .A(\inv_in[1629] ));
 sg13g2_inv_2 \inv[162]/_0_  (.Y(\inv_in[163] ),
    .A(\inv_in[162] ));
 sg13g2_inv_2 \inv[1630]/_0_  (.Y(\inv_in[1631] ),
    .A(\inv_in[1630] ));
 sg13g2_inv_2 \inv[1631]/_0_  (.Y(\inv_in[1632] ),
    .A(\inv_in[1631] ));
 sg13g2_inv_2 \inv[1632]/_0_  (.Y(\inv_in[1633] ),
    .A(\inv_in[1632] ));
 sg13g2_inv_2 \inv[1633]/_0_  (.Y(\inv_in[1634] ),
    .A(\inv_in[1633] ));
 sg13g2_inv_2 \inv[1634]/_0_  (.Y(\inv_in[1635] ),
    .A(\inv_in[1634] ));
 sg13g2_inv_2 \inv[1635]/_0_  (.Y(\inv_in[1636] ),
    .A(\inv_in[1635] ));
 sg13g2_inv_2 \inv[1636]/_0_  (.Y(\inv_in[1637] ),
    .A(\inv_in[1636] ));
 sg13g2_inv_2 \inv[1637]/_0_  (.Y(\inv_in[1638] ),
    .A(\inv_in[1637] ));
 sg13g2_inv_2 \inv[1638]/_0_  (.Y(\inv_in[1639] ),
    .A(\inv_in[1638] ));
 sg13g2_inv_2 \inv[1639]/_0_  (.Y(\inv_in[1640] ),
    .A(\inv_in[1639] ));
 sg13g2_inv_2 \inv[163]/_0_  (.Y(\inv_in[164] ),
    .A(\inv_in[163] ));
 sg13g2_inv_2 \inv[1640]/_0_  (.Y(\inv_in[1641] ),
    .A(\inv_in[1640] ));
 sg13g2_inv_2 \inv[1641]/_0_  (.Y(\inv_in[1642] ),
    .A(\inv_in[1641] ));
 sg13g2_inv_2 \inv[1642]/_0_  (.Y(\inv_in[1643] ),
    .A(\inv_in[1642] ));
 sg13g2_inv_2 \inv[1643]/_0_  (.Y(\inv_in[1644] ),
    .A(\inv_in[1643] ));
 sg13g2_inv_2 \inv[1644]/_0_  (.Y(\inv_in[1645] ),
    .A(\inv_in[1644] ));
 sg13g2_inv_2 \inv[1645]/_0_  (.Y(\inv_in[1646] ),
    .A(\inv_in[1645] ));
 sg13g2_inv_2 \inv[1646]/_0_  (.Y(\inv_in[1647] ),
    .A(\inv_in[1646] ));
 sg13g2_inv_2 \inv[1647]/_0_  (.Y(\inv_in[1648] ),
    .A(\inv_in[1647] ));
 sg13g2_inv_2 \inv[1648]/_0_  (.Y(\inv_in[1649] ),
    .A(\inv_in[1648] ));
 sg13g2_inv_2 \inv[1649]/_0_  (.Y(\inv_in[1650] ),
    .A(\inv_in[1649] ));
 sg13g2_inv_2 \inv[164]/_0_  (.Y(\inv_in[165] ),
    .A(\inv_in[164] ));
 sg13g2_inv_2 \inv[1650]/_0_  (.Y(\inv_in[1651] ),
    .A(\inv_in[1650] ));
 sg13g2_inv_2 \inv[1651]/_0_  (.Y(\inv_in[1652] ),
    .A(\inv_in[1651] ));
 sg13g2_inv_2 \inv[1652]/_0_  (.Y(\inv_in[1653] ),
    .A(\inv_in[1652] ));
 sg13g2_inv_2 \inv[1653]/_0_  (.Y(\inv_in[1654] ),
    .A(\inv_in[1653] ));
 sg13g2_inv_2 \inv[1654]/_0_  (.Y(\inv_in[1655] ),
    .A(\inv_in[1654] ));
 sg13g2_inv_2 \inv[1655]/_0_  (.Y(\inv_in[1656] ),
    .A(\inv_in[1655] ));
 sg13g2_inv_2 \inv[1656]/_0_  (.Y(\inv_in[1657] ),
    .A(\inv_in[1656] ));
 sg13g2_inv_2 \inv[1657]/_0_  (.Y(\inv_in[1658] ),
    .A(\inv_in[1657] ));
 sg13g2_inv_2 \inv[1658]/_0_  (.Y(\inv_in[1659] ),
    .A(\inv_in[1658] ));
 sg13g2_inv_2 \inv[1659]/_0_  (.Y(\inv_in[1660] ),
    .A(\inv_in[1659] ));
 sg13g2_inv_2 \inv[165]/_0_  (.Y(\inv_in[166] ),
    .A(\inv_in[165] ));
 sg13g2_inv_2 \inv[1660]/_0_  (.Y(\inv_in[1661] ),
    .A(\inv_in[1660] ));
 sg13g2_inv_2 \inv[1661]/_0_  (.Y(\inv_in[1662] ),
    .A(\inv_in[1661] ));
 sg13g2_inv_2 \inv[1662]/_0_  (.Y(\inv_in[1663] ),
    .A(\inv_in[1662] ));
 sg13g2_inv_2 \inv[1663]/_0_  (.Y(\inv_in[1664] ),
    .A(\inv_in[1663] ));
 sg13g2_inv_2 \inv[1664]/_0_  (.Y(\inv_in[1665] ),
    .A(\inv_in[1664] ));
 sg13g2_inv_2 \inv[1665]/_0_  (.Y(\inv_in[1666] ),
    .A(\inv_in[1665] ));
 sg13g2_inv_2 \inv[1666]/_0_  (.Y(\inv_in[1667] ),
    .A(\inv_in[1666] ));
 sg13g2_inv_2 \inv[1667]/_0_  (.Y(\inv_in[1668] ),
    .A(\inv_in[1667] ));
 sg13g2_inv_2 \inv[1668]/_0_  (.Y(\inv_in[1669] ),
    .A(\inv_in[1668] ));
 sg13g2_inv_2 \inv[1669]/_0_  (.Y(\inv_in[1670] ),
    .A(\inv_in[1669] ));
 sg13g2_inv_2 \inv[166]/_0_  (.Y(\inv_in[167] ),
    .A(\inv_in[166] ));
 sg13g2_inv_2 \inv[1670]/_0_  (.Y(\inv_in[1671] ),
    .A(\inv_in[1670] ));
 sg13g2_inv_2 \inv[1671]/_0_  (.Y(\inv_in[1672] ),
    .A(\inv_in[1671] ));
 sg13g2_inv_2 \inv[1672]/_0_  (.Y(\inv_in[1673] ),
    .A(\inv_in[1672] ));
 sg13g2_inv_2 \inv[1673]/_0_  (.Y(\inv_in[1674] ),
    .A(\inv_in[1673] ));
 sg13g2_inv_2 \inv[1674]/_0_  (.Y(\inv_in[1675] ),
    .A(\inv_in[1674] ));
 sg13g2_inv_2 \inv[1675]/_0_  (.Y(\inv_in[1676] ),
    .A(\inv_in[1675] ));
 sg13g2_inv_2 \inv[1676]/_0_  (.Y(\inv_in[1677] ),
    .A(\inv_in[1676] ));
 sg13g2_inv_2 \inv[1677]/_0_  (.Y(\inv_in[1678] ),
    .A(\inv_in[1677] ));
 sg13g2_inv_2 \inv[1678]/_0_  (.Y(\inv_in[1679] ),
    .A(\inv_in[1678] ));
 sg13g2_inv_2 \inv[1679]/_0_  (.Y(\inv_in[1680] ),
    .A(\inv_in[1679] ));
 sg13g2_inv_2 \inv[167]/_0_  (.Y(\inv_in[168] ),
    .A(\inv_in[167] ));
 sg13g2_inv_2 \inv[1680]/_0_  (.Y(\inv_in[1681] ),
    .A(\inv_in[1680] ));
 sg13g2_inv_2 \inv[1681]/_0_  (.Y(\inv_in[1682] ),
    .A(\inv_in[1681] ));
 sg13g2_inv_2 \inv[1682]/_0_  (.Y(\inv_in[1683] ),
    .A(\inv_in[1682] ));
 sg13g2_inv_2 \inv[1683]/_0_  (.Y(\inv_in[1684] ),
    .A(\inv_in[1683] ));
 sg13g2_inv_2 \inv[1684]/_0_  (.Y(\inv_in[1685] ),
    .A(\inv_in[1684] ));
 sg13g2_inv_2 \inv[1685]/_0_  (.Y(\inv_in[1686] ),
    .A(\inv_in[1685] ));
 sg13g2_inv_2 \inv[1686]/_0_  (.Y(\inv_in[1687] ),
    .A(\inv_in[1686] ));
 sg13g2_inv_2 \inv[1687]/_0_  (.Y(\inv_in[1688] ),
    .A(\inv_in[1687] ));
 sg13g2_inv_2 \inv[1688]/_0_  (.Y(\inv_in[1689] ),
    .A(\inv_in[1688] ));
 sg13g2_inv_2 \inv[1689]/_0_  (.Y(\inv_in[1690] ),
    .A(\inv_in[1689] ));
 sg13g2_inv_2 \inv[168]/_0_  (.Y(\inv_in[169] ),
    .A(\inv_in[168] ));
 sg13g2_inv_2 \inv[1690]/_0_  (.Y(\inv_in[1691] ),
    .A(\inv_in[1690] ));
 sg13g2_inv_2 \inv[1691]/_0_  (.Y(\inv_in[1692] ),
    .A(\inv_in[1691] ));
 sg13g2_inv_2 \inv[1692]/_0_  (.Y(\inv_in[1693] ),
    .A(\inv_in[1692] ));
 sg13g2_inv_2 \inv[1693]/_0_  (.Y(\inv_in[1694] ),
    .A(\inv_in[1693] ));
 sg13g2_inv_2 \inv[1694]/_0_  (.Y(\inv_in[1695] ),
    .A(\inv_in[1694] ));
 sg13g2_inv_2 \inv[1695]/_0_  (.Y(\inv_in[1696] ),
    .A(\inv_in[1695] ));
 sg13g2_inv_2 \inv[1696]/_0_  (.Y(\inv_in[1697] ),
    .A(\inv_in[1696] ));
 sg13g2_inv_2 \inv[1697]/_0_  (.Y(\inv_in[1698] ),
    .A(\inv_in[1697] ));
 sg13g2_inv_2 \inv[1698]/_0_  (.Y(\inv_in[1699] ),
    .A(\inv_in[1698] ));
 sg13g2_inv_2 \inv[1699]/_0_  (.Y(\inv_in[1700] ),
    .A(\inv_in[1699] ));
 sg13g2_inv_2 \inv[169]/_0_  (.Y(\inv_in[170] ),
    .A(\inv_in[169] ));
 sg13g2_inv_2 \inv[16]/_0_  (.Y(\inv_in[17] ),
    .A(\inv_in[16] ));
 sg13g2_inv_2 \inv[1700]/_0_  (.Y(\inv_in[1701] ),
    .A(\inv_in[1700] ));
 sg13g2_inv_2 \inv[1701]/_0_  (.Y(\inv_in[1702] ),
    .A(\inv_in[1701] ));
 sg13g2_inv_2 \inv[1702]/_0_  (.Y(\inv_in[1703] ),
    .A(\inv_in[1702] ));
 sg13g2_inv_2 \inv[1703]/_0_  (.Y(\inv_in[1704] ),
    .A(\inv_in[1703] ));
 sg13g2_inv_2 \inv[1704]/_0_  (.Y(\inv_in[1705] ),
    .A(\inv_in[1704] ));
 sg13g2_inv_2 \inv[1705]/_0_  (.Y(\inv_in[1706] ),
    .A(\inv_in[1705] ));
 sg13g2_inv_2 \inv[1706]/_0_  (.Y(\inv_in[1707] ),
    .A(\inv_in[1706] ));
 sg13g2_inv_2 \inv[1707]/_0_  (.Y(\inv_in[1708] ),
    .A(\inv_in[1707] ));
 sg13g2_inv_2 \inv[1708]/_0_  (.Y(\inv_in[1709] ),
    .A(\inv_in[1708] ));
 sg13g2_inv_2 \inv[1709]/_0_  (.Y(\inv_in[1710] ),
    .A(\inv_in[1709] ));
 sg13g2_inv_2 \inv[170]/_0_  (.Y(\inv_in[171] ),
    .A(\inv_in[170] ));
 sg13g2_inv_2 \inv[1710]/_0_  (.Y(\inv_in[1711] ),
    .A(\inv_in[1710] ));
 sg13g2_inv_2 \inv[1711]/_0_  (.Y(\inv_in[1712] ),
    .A(\inv_in[1711] ));
 sg13g2_inv_2 \inv[1712]/_0_  (.Y(\inv_in[1713] ),
    .A(\inv_in[1712] ));
 sg13g2_inv_2 \inv[1713]/_0_  (.Y(\inv_in[1714] ),
    .A(\inv_in[1713] ));
 sg13g2_inv_2 \inv[1714]/_0_  (.Y(\inv_in[1715] ),
    .A(\inv_in[1714] ));
 sg13g2_inv_2 \inv[1715]/_0_  (.Y(\inv_in[1716] ),
    .A(\inv_in[1715] ));
 sg13g2_inv_2 \inv[1716]/_0_  (.Y(\inv_in[1717] ),
    .A(\inv_in[1716] ));
 sg13g2_inv_2 \inv[1717]/_0_  (.Y(\inv_in[1718] ),
    .A(\inv_in[1717] ));
 sg13g2_inv_2 \inv[1718]/_0_  (.Y(\inv_in[1719] ),
    .A(\inv_in[1718] ));
 sg13g2_inv_2 \inv[1719]/_0_  (.Y(\inv_in[1720] ),
    .A(\inv_in[1719] ));
 sg13g2_inv_2 \inv[171]/_0_  (.Y(\inv_in[172] ),
    .A(\inv_in[171] ));
 sg13g2_inv_2 \inv[1720]/_0_  (.Y(\inv_in[1721] ),
    .A(\inv_in[1720] ));
 sg13g2_inv_2 \inv[1721]/_0_  (.Y(\inv_in[1722] ),
    .A(\inv_in[1721] ));
 sg13g2_inv_2 \inv[1722]/_0_  (.Y(\inv_in[1723] ),
    .A(\inv_in[1722] ));
 sg13g2_inv_2 \inv[1723]/_0_  (.Y(\inv_in[1724] ),
    .A(\inv_in[1723] ));
 sg13g2_inv_2 \inv[1724]/_0_  (.Y(\inv_in[1725] ),
    .A(\inv_in[1724] ));
 sg13g2_inv_2 \inv[1725]/_0_  (.Y(\inv_in[1726] ),
    .A(\inv_in[1725] ));
 sg13g2_inv_2 \inv[1726]/_0_  (.Y(\inv_in[1727] ),
    .A(\inv_in[1726] ));
 sg13g2_inv_2 \inv[1727]/_0_  (.Y(\inv_in[1728] ),
    .A(\inv_in[1727] ));
 sg13g2_inv_2 \inv[1728]/_0_  (.Y(\inv_in[1729] ),
    .A(\inv_in[1728] ));
 sg13g2_inv_2 \inv[1729]/_0_  (.Y(\inv_in[1730] ),
    .A(\inv_in[1729] ));
 sg13g2_inv_2 \inv[172]/_0_  (.Y(\inv_in[173] ),
    .A(\inv_in[172] ));
 sg13g2_inv_2 \inv[1730]/_0_  (.Y(\inv_in[1731] ),
    .A(\inv_in[1730] ));
 sg13g2_inv_2 \inv[1731]/_0_  (.Y(\inv_in[1732] ),
    .A(\inv_in[1731] ));
 sg13g2_inv_2 \inv[1732]/_0_  (.Y(\inv_in[1733] ),
    .A(\inv_in[1732] ));
 sg13g2_inv_2 \inv[1733]/_0_  (.Y(\inv_in[1734] ),
    .A(\inv_in[1733] ));
 sg13g2_inv_2 \inv[1734]/_0_  (.Y(\inv_in[1735] ),
    .A(\inv_in[1734] ));
 sg13g2_inv_2 \inv[1735]/_0_  (.Y(\inv_in[1736] ),
    .A(\inv_in[1735] ));
 sg13g2_inv_2 \inv[1736]/_0_  (.Y(\inv_in[1737] ),
    .A(\inv_in[1736] ));
 sg13g2_inv_2 \inv[1737]/_0_  (.Y(\inv_in[1738] ),
    .A(\inv_in[1737] ));
 sg13g2_inv_2 \inv[1738]/_0_  (.Y(\inv_in[1739] ),
    .A(\inv_in[1738] ));
 sg13g2_inv_2 \inv[1739]/_0_  (.Y(\inv_in[1740] ),
    .A(\inv_in[1739] ));
 sg13g2_inv_2 \inv[173]/_0_  (.Y(\inv_in[174] ),
    .A(\inv_in[173] ));
 sg13g2_inv_2 \inv[1740]/_0_  (.Y(\inv_in[1741] ),
    .A(\inv_in[1740] ));
 sg13g2_inv_2 \inv[1741]/_0_  (.Y(\inv_in[1742] ),
    .A(\inv_in[1741] ));
 sg13g2_inv_2 \inv[1742]/_0_  (.Y(\inv_in[1743] ),
    .A(\inv_in[1742] ));
 sg13g2_inv_2 \inv[1743]/_0_  (.Y(\inv_in[1744] ),
    .A(\inv_in[1743] ));
 sg13g2_inv_2 \inv[1744]/_0_  (.Y(\inv_in[1745] ),
    .A(\inv_in[1744] ));
 sg13g2_inv_2 \inv[1745]/_0_  (.Y(\inv_in[1746] ),
    .A(\inv_in[1745] ));
 sg13g2_inv_2 \inv[1746]/_0_  (.Y(\inv_in[1747] ),
    .A(\inv_in[1746] ));
 sg13g2_inv_2 \inv[1747]/_0_  (.Y(\inv_in[1748] ),
    .A(\inv_in[1747] ));
 sg13g2_inv_2 \inv[1748]/_0_  (.Y(\inv_in[1749] ),
    .A(\inv_in[1748] ));
 sg13g2_inv_2 \inv[1749]/_0_  (.Y(\inv_in[1750] ),
    .A(\inv_in[1749] ));
 sg13g2_inv_2 \inv[174]/_0_  (.Y(\inv_in[175] ),
    .A(\inv_in[174] ));
 sg13g2_inv_2 \inv[1750]/_0_  (.Y(\inv_in[1751] ),
    .A(\inv_in[1750] ));
 sg13g2_inv_2 \inv[1751]/_0_  (.Y(\inv_in[1752] ),
    .A(\inv_in[1751] ));
 sg13g2_inv_2 \inv[1752]/_0_  (.Y(\inv_in[1753] ),
    .A(\inv_in[1752] ));
 sg13g2_inv_2 \inv[1753]/_0_  (.Y(\inv_in[1754] ),
    .A(\inv_in[1753] ));
 sg13g2_inv_2 \inv[1754]/_0_  (.Y(\inv_in[1755] ),
    .A(\inv_in[1754] ));
 sg13g2_inv_2 \inv[1755]/_0_  (.Y(\inv_in[1756] ),
    .A(\inv_in[1755] ));
 sg13g2_inv_2 \inv[1756]/_0_  (.Y(\inv_in[1757] ),
    .A(\inv_in[1756] ));
 sg13g2_inv_2 \inv[1757]/_0_  (.Y(\inv_in[1758] ),
    .A(\inv_in[1757] ));
 sg13g2_inv_2 \inv[1758]/_0_  (.Y(\inv_in[1759] ),
    .A(\inv_in[1758] ));
 sg13g2_inv_2 \inv[1759]/_0_  (.Y(\inv_in[1760] ),
    .A(\inv_in[1759] ));
 sg13g2_inv_2 \inv[175]/_0_  (.Y(\inv_in[176] ),
    .A(\inv_in[175] ));
 sg13g2_inv_2 \inv[1760]/_0_  (.Y(\inv_in[1761] ),
    .A(\inv_in[1760] ));
 sg13g2_inv_2 \inv[1761]/_0_  (.Y(\inv_in[1762] ),
    .A(\inv_in[1761] ));
 sg13g2_inv_2 \inv[1762]/_0_  (.Y(\inv_in[1763] ),
    .A(\inv_in[1762] ));
 sg13g2_inv_2 \inv[1763]/_0_  (.Y(\inv_in[1764] ),
    .A(\inv_in[1763] ));
 sg13g2_inv_2 \inv[1764]/_0_  (.Y(\inv_in[1765] ),
    .A(\inv_in[1764] ));
 sg13g2_inv_2 \inv[1765]/_0_  (.Y(\inv_in[1766] ),
    .A(\inv_in[1765] ));
 sg13g2_inv_2 \inv[1766]/_0_  (.Y(\inv_in[1767] ),
    .A(\inv_in[1766] ));
 sg13g2_inv_2 \inv[1767]/_0_  (.Y(\inv_in[1768] ),
    .A(\inv_in[1767] ));
 sg13g2_inv_2 \inv[1768]/_0_  (.Y(\inv_in[1769] ),
    .A(\inv_in[1768] ));
 sg13g2_inv_2 \inv[1769]/_0_  (.Y(\inv_in[1770] ),
    .A(\inv_in[1769] ));
 sg13g2_inv_2 \inv[176]/_0_  (.Y(\inv_in[177] ),
    .A(\inv_in[176] ));
 sg13g2_inv_2 \inv[1770]/_0_  (.Y(\inv_in[1771] ),
    .A(\inv_in[1770] ));
 sg13g2_inv_2 \inv[1771]/_0_  (.Y(\inv_in[1772] ),
    .A(\inv_in[1771] ));
 sg13g2_inv_2 \inv[1772]/_0_  (.Y(\inv_in[1773] ),
    .A(\inv_in[1772] ));
 sg13g2_inv_2 \inv[1773]/_0_  (.Y(\inv_in[1774] ),
    .A(\inv_in[1773] ));
 sg13g2_inv_2 \inv[1774]/_0_  (.Y(\inv_in[1775] ),
    .A(\inv_in[1774] ));
 sg13g2_inv_2 \inv[1775]/_0_  (.Y(\inv_in[1776] ),
    .A(\inv_in[1775] ));
 sg13g2_inv_2 \inv[1776]/_0_  (.Y(\inv_in[1777] ),
    .A(\inv_in[1776] ));
 sg13g2_inv_2 \inv[1777]/_0_  (.Y(\inv_in[1778] ),
    .A(\inv_in[1777] ));
 sg13g2_inv_2 \inv[1778]/_0_  (.Y(\inv_in[1779] ),
    .A(\inv_in[1778] ));
 sg13g2_inv_2 \inv[1779]/_0_  (.Y(\inv_in[1780] ),
    .A(\inv_in[1779] ));
 sg13g2_inv_2 \inv[177]/_0_  (.Y(\inv_in[178] ),
    .A(\inv_in[177] ));
 sg13g2_inv_2 \inv[1780]/_0_  (.Y(\inv_in[1781] ),
    .A(\inv_in[1780] ));
 sg13g2_inv_2 \inv[1781]/_0_  (.Y(\inv_in[1782] ),
    .A(\inv_in[1781] ));
 sg13g2_inv_2 \inv[1782]/_0_  (.Y(\inv_in[1783] ),
    .A(\inv_in[1782] ));
 sg13g2_inv_2 \inv[1783]/_0_  (.Y(\inv_in[1784] ),
    .A(\inv_in[1783] ));
 sg13g2_inv_2 \inv[1784]/_0_  (.Y(\inv_in[1785] ),
    .A(\inv_in[1784] ));
 sg13g2_inv_2 \inv[1785]/_0_  (.Y(\inv_in[1786] ),
    .A(\inv_in[1785] ));
 sg13g2_inv_2 \inv[1786]/_0_  (.Y(\inv_in[1787] ),
    .A(\inv_in[1786] ));
 sg13g2_inv_2 \inv[1787]/_0_  (.Y(\inv_in[1788] ),
    .A(\inv_in[1787] ));
 sg13g2_inv_2 \inv[1788]/_0_  (.Y(\inv_in[1789] ),
    .A(\inv_in[1788] ));
 sg13g2_inv_2 \inv[1789]/_0_  (.Y(\inv_in[1790] ),
    .A(\inv_in[1789] ));
 sg13g2_inv_2 \inv[178]/_0_  (.Y(\inv_in[179] ),
    .A(\inv_in[178] ));
 sg13g2_inv_2 \inv[1790]/_0_  (.Y(\inv_in[1791] ),
    .A(\inv_in[1790] ));
 sg13g2_inv_2 \inv[1791]/_0_  (.Y(\inv_in[1792] ),
    .A(\inv_in[1791] ));
 sg13g2_inv_2 \inv[1792]/_0_  (.Y(\inv_in[1793] ),
    .A(\inv_in[1792] ));
 sg13g2_inv_2 \inv[1793]/_0_  (.Y(\inv_in[1794] ),
    .A(\inv_in[1793] ));
 sg13g2_inv_2 \inv[1794]/_0_  (.Y(\inv_in[1795] ),
    .A(\inv_in[1794] ));
 sg13g2_inv_2 \inv[1795]/_0_  (.Y(\inv_in[1796] ),
    .A(\inv_in[1795] ));
 sg13g2_inv_2 \inv[1796]/_0_  (.Y(\inv_in[1797] ),
    .A(\inv_in[1796] ));
 sg13g2_inv_2 \inv[1797]/_0_  (.Y(\inv_in[1798] ),
    .A(\inv_in[1797] ));
 sg13g2_inv_2 \inv[1798]/_0_  (.Y(\inv_in[1799] ),
    .A(\inv_in[1798] ));
 sg13g2_inv_2 \inv[1799]/_0_  (.Y(\inv_in[1800] ),
    .A(\inv_in[1799] ));
 sg13g2_inv_2 \inv[179]/_0_  (.Y(\inv_in[180] ),
    .A(\inv_in[179] ));
 sg13g2_inv_2 \inv[17]/_0_  (.Y(\inv_in[18] ),
    .A(\inv_in[17] ));
 sg13g2_inv_2 \inv[1800]/_0_  (.Y(\inv_in[1801] ),
    .A(\inv_in[1800] ));
 sg13g2_inv_2 \inv[1801]/_0_  (.Y(\inv_in[1802] ),
    .A(\inv_in[1801] ));
 sg13g2_inv_2 \inv[1802]/_0_  (.Y(\inv_in[1803] ),
    .A(\inv_in[1802] ));
 sg13g2_inv_2 \inv[1803]/_0_  (.Y(\inv_in[1804] ),
    .A(\inv_in[1803] ));
 sg13g2_inv_2 \inv[1804]/_0_  (.Y(\inv_in[1805] ),
    .A(\inv_in[1804] ));
 sg13g2_inv_2 \inv[1805]/_0_  (.Y(\inv_in[1806] ),
    .A(\inv_in[1805] ));
 sg13g2_inv_2 \inv[1806]/_0_  (.Y(\inv_in[1807] ),
    .A(\inv_in[1806] ));
 sg13g2_inv_2 \inv[1807]/_0_  (.Y(\inv_in[1808] ),
    .A(\inv_in[1807] ));
 sg13g2_inv_2 \inv[1808]/_0_  (.Y(\inv_in[1809] ),
    .A(\inv_in[1808] ));
 sg13g2_inv_2 \inv[1809]/_0_  (.Y(\inv_in[1810] ),
    .A(\inv_in[1809] ));
 sg13g2_inv_2 \inv[180]/_0_  (.Y(\inv_in[181] ),
    .A(\inv_in[180] ));
 sg13g2_inv_2 \inv[1810]/_0_  (.Y(\inv_in[1811] ),
    .A(\inv_in[1810] ));
 sg13g2_inv_2 \inv[1811]/_0_  (.Y(\inv_in[1812] ),
    .A(\inv_in[1811] ));
 sg13g2_inv_2 \inv[1812]/_0_  (.Y(\inv_in[1813] ),
    .A(\inv_in[1812] ));
 sg13g2_inv_2 \inv[1813]/_0_  (.Y(\inv_in[1814] ),
    .A(\inv_in[1813] ));
 sg13g2_inv_2 \inv[1814]/_0_  (.Y(\inv_in[1815] ),
    .A(\inv_in[1814] ));
 sg13g2_inv_2 \inv[1815]/_0_  (.Y(\inv_in[1816] ),
    .A(\inv_in[1815] ));
 sg13g2_inv_2 \inv[1816]/_0_  (.Y(\inv_in[1817] ),
    .A(\inv_in[1816] ));
 sg13g2_inv_2 \inv[1817]/_0_  (.Y(\inv_in[1818] ),
    .A(\inv_in[1817] ));
 sg13g2_inv_2 \inv[1818]/_0_  (.Y(\inv_in[1819] ),
    .A(\inv_in[1818] ));
 sg13g2_inv_2 \inv[1819]/_0_  (.Y(\inv_in[1820] ),
    .A(\inv_in[1819] ));
 sg13g2_inv_2 \inv[181]/_0_  (.Y(\inv_in[182] ),
    .A(\inv_in[181] ));
 sg13g2_inv_2 \inv[1820]/_0_  (.Y(\inv_in[1821] ),
    .A(\inv_in[1820] ));
 sg13g2_inv_2 \inv[1821]/_0_  (.Y(\inv_in[1822] ),
    .A(\inv_in[1821] ));
 sg13g2_inv_2 \inv[1822]/_0_  (.Y(\inv_in[1823] ),
    .A(\inv_in[1822] ));
 sg13g2_inv_2 \inv[1823]/_0_  (.Y(\inv_in[1824] ),
    .A(\inv_in[1823] ));
 sg13g2_inv_2 \inv[1824]/_0_  (.Y(\inv_in[1825] ),
    .A(\inv_in[1824] ));
 sg13g2_inv_2 \inv[1825]/_0_  (.Y(\inv_in[1826] ),
    .A(\inv_in[1825] ));
 sg13g2_inv_2 \inv[1826]/_0_  (.Y(\inv_in[1827] ),
    .A(\inv_in[1826] ));
 sg13g2_inv_2 \inv[1827]/_0_  (.Y(\inv_in[1828] ),
    .A(\inv_in[1827] ));
 sg13g2_inv_2 \inv[1828]/_0_  (.Y(\inv_in[1829] ),
    .A(\inv_in[1828] ));
 sg13g2_inv_2 \inv[1829]/_0_  (.Y(\inv_in[1830] ),
    .A(\inv_in[1829] ));
 sg13g2_inv_2 \inv[182]/_0_  (.Y(\inv_in[183] ),
    .A(\inv_in[182] ));
 sg13g2_inv_2 \inv[1830]/_0_  (.Y(\inv_in[1831] ),
    .A(\inv_in[1830] ));
 sg13g2_inv_2 \inv[1831]/_0_  (.Y(\inv_in[1832] ),
    .A(\inv_in[1831] ));
 sg13g2_inv_2 \inv[1832]/_0_  (.Y(\inv_in[1833] ),
    .A(\inv_in[1832] ));
 sg13g2_inv_2 \inv[1833]/_0_  (.Y(\inv_in[1834] ),
    .A(\inv_in[1833] ));
 sg13g2_inv_2 \inv[1834]/_0_  (.Y(\inv_in[1835] ),
    .A(\inv_in[1834] ));
 sg13g2_inv_2 \inv[1835]/_0_  (.Y(\inv_in[1836] ),
    .A(\inv_in[1835] ));
 sg13g2_inv_2 \inv[1836]/_0_  (.Y(\inv_in[1837] ),
    .A(\inv_in[1836] ));
 sg13g2_inv_2 \inv[1837]/_0_  (.Y(\inv_in[1838] ),
    .A(\inv_in[1837] ));
 sg13g2_inv_2 \inv[1838]/_0_  (.Y(\inv_in[1839] ),
    .A(\inv_in[1838] ));
 sg13g2_inv_2 \inv[1839]/_0_  (.Y(\inv_in[1840] ),
    .A(\inv_in[1839] ));
 sg13g2_inv_2 \inv[183]/_0_  (.Y(\inv_in[184] ),
    .A(\inv_in[183] ));
 sg13g2_inv_2 \inv[1840]/_0_  (.Y(\inv_in[1841] ),
    .A(\inv_in[1840] ));
 sg13g2_inv_2 \inv[1841]/_0_  (.Y(\inv_in[1842] ),
    .A(\inv_in[1841] ));
 sg13g2_inv_2 \inv[1842]/_0_  (.Y(\inv_in[1843] ),
    .A(\inv_in[1842] ));
 sg13g2_inv_2 \inv[1843]/_0_  (.Y(\inv_in[1844] ),
    .A(\inv_in[1843] ));
 sg13g2_inv_2 \inv[1844]/_0_  (.Y(\inv_in[1845] ),
    .A(\inv_in[1844] ));
 sg13g2_inv_2 \inv[1845]/_0_  (.Y(\inv_in[1846] ),
    .A(\inv_in[1845] ));
 sg13g2_inv_2 \inv[1846]/_0_  (.Y(\inv_in[1847] ),
    .A(\inv_in[1846] ));
 sg13g2_inv_2 \inv[1847]/_0_  (.Y(\inv_in[1848] ),
    .A(\inv_in[1847] ));
 sg13g2_inv_2 \inv[1848]/_0_  (.Y(\inv_in[1849] ),
    .A(\inv_in[1848] ));
 sg13g2_inv_2 \inv[1849]/_0_  (.Y(\inv_in[1850] ),
    .A(\inv_in[1849] ));
 sg13g2_inv_2 \inv[184]/_0_  (.Y(\inv_in[185] ),
    .A(\inv_in[184] ));
 sg13g2_inv_2 \inv[1850]/_0_  (.Y(\inv_in[1851] ),
    .A(\inv_in[1850] ));
 sg13g2_inv_2 \inv[1851]/_0_  (.Y(\inv_in[1852] ),
    .A(\inv_in[1851] ));
 sg13g2_inv_2 \inv[1852]/_0_  (.Y(\inv_in[1853] ),
    .A(\inv_in[1852] ));
 sg13g2_inv_2 \inv[1853]/_0_  (.Y(\inv_in[1854] ),
    .A(\inv_in[1853] ));
 sg13g2_inv_2 \inv[1854]/_0_  (.Y(\inv_in[1855] ),
    .A(\inv_in[1854] ));
 sg13g2_inv_2 \inv[1855]/_0_  (.Y(\inv_in[1856] ),
    .A(\inv_in[1855] ));
 sg13g2_inv_2 \inv[1856]/_0_  (.Y(\inv_in[1857] ),
    .A(\inv_in[1856] ));
 sg13g2_inv_2 \inv[1857]/_0_  (.Y(\inv_in[1858] ),
    .A(\inv_in[1857] ));
 sg13g2_inv_2 \inv[1858]/_0_  (.Y(\inv_in[1859] ),
    .A(\inv_in[1858] ));
 sg13g2_inv_2 \inv[1859]/_0_  (.Y(\inv_in[1860] ),
    .A(\inv_in[1859] ));
 sg13g2_inv_2 \inv[185]/_0_  (.Y(\inv_in[186] ),
    .A(\inv_in[185] ));
 sg13g2_inv_2 \inv[1860]/_0_  (.Y(\inv_in[1861] ),
    .A(\inv_in[1860] ));
 sg13g2_inv_2 \inv[1861]/_0_  (.Y(\inv_in[1862] ),
    .A(\inv_in[1861] ));
 sg13g2_inv_2 \inv[1862]/_0_  (.Y(\inv_in[1863] ),
    .A(\inv_in[1862] ));
 sg13g2_inv_2 \inv[1863]/_0_  (.Y(\inv_in[1864] ),
    .A(\inv_in[1863] ));
 sg13g2_inv_2 \inv[1864]/_0_  (.Y(\inv_in[1865] ),
    .A(\inv_in[1864] ));
 sg13g2_inv_2 \inv[1865]/_0_  (.Y(\inv_in[1866] ),
    .A(\inv_in[1865] ));
 sg13g2_inv_2 \inv[1866]/_0_  (.Y(\inv_in[1867] ),
    .A(\inv_in[1866] ));
 sg13g2_inv_2 \inv[1867]/_0_  (.Y(\inv_in[1868] ),
    .A(\inv_in[1867] ));
 sg13g2_inv_2 \inv[1868]/_0_  (.Y(\inv_in[1869] ),
    .A(\inv_in[1868] ));
 sg13g2_inv_2 \inv[1869]/_0_  (.Y(\inv_in[1870] ),
    .A(\inv_in[1869] ));
 sg13g2_inv_2 \inv[186]/_0_  (.Y(\inv_in[187] ),
    .A(\inv_in[186] ));
 sg13g2_inv_2 \inv[1870]/_0_  (.Y(\inv_in[1871] ),
    .A(\inv_in[1870] ));
 sg13g2_inv_2 \inv[1871]/_0_  (.Y(\inv_in[1872] ),
    .A(\inv_in[1871] ));
 sg13g2_inv_2 \inv[1872]/_0_  (.Y(\inv_in[1873] ),
    .A(\inv_in[1872] ));
 sg13g2_inv_2 \inv[1873]/_0_  (.Y(\inv_in[1874] ),
    .A(\inv_in[1873] ));
 sg13g2_inv_2 \inv[1874]/_0_  (.Y(\inv_in[1875] ),
    .A(\inv_in[1874] ));
 sg13g2_inv_2 \inv[1875]/_0_  (.Y(\inv_in[1876] ),
    .A(\inv_in[1875] ));
 sg13g2_inv_2 \inv[1876]/_0_  (.Y(\inv_in[1877] ),
    .A(\inv_in[1876] ));
 sg13g2_inv_2 \inv[1877]/_0_  (.Y(\inv_in[1878] ),
    .A(\inv_in[1877] ));
 sg13g2_inv_2 \inv[1878]/_0_  (.Y(\inv_in[1879] ),
    .A(\inv_in[1878] ));
 sg13g2_inv_2 \inv[1879]/_0_  (.Y(\inv_in[1880] ),
    .A(\inv_in[1879] ));
 sg13g2_inv_2 \inv[187]/_0_  (.Y(\inv_in[188] ),
    .A(\inv_in[187] ));
 sg13g2_inv_2 \inv[1880]/_0_  (.Y(\inv_in[1881] ),
    .A(\inv_in[1880] ));
 sg13g2_inv_2 \inv[1881]/_0_  (.Y(\inv_in[1882] ),
    .A(\inv_in[1881] ));
 sg13g2_inv_2 \inv[1882]/_0_  (.Y(\inv_in[1883] ),
    .A(\inv_in[1882] ));
 sg13g2_inv_2 \inv[1883]/_0_  (.Y(\inv_in[1884] ),
    .A(\inv_in[1883] ));
 sg13g2_inv_2 \inv[1884]/_0_  (.Y(\inv_in[1885] ),
    .A(\inv_in[1884] ));
 sg13g2_inv_2 \inv[1885]/_0_  (.Y(\inv_in[1886] ),
    .A(\inv_in[1885] ));
 sg13g2_inv_2 \inv[1886]/_0_  (.Y(\inv_in[1887] ),
    .A(\inv_in[1886] ));
 sg13g2_inv_2 \inv[1887]/_0_  (.Y(\inv_in[1888] ),
    .A(\inv_in[1887] ));
 sg13g2_inv_2 \inv[1888]/_0_  (.Y(\inv_in[1889] ),
    .A(\inv_in[1888] ));
 sg13g2_inv_2 \inv[1889]/_0_  (.Y(\inv_in[1890] ),
    .A(\inv_in[1889] ));
 sg13g2_inv_2 \inv[188]/_0_  (.Y(\inv_in[189] ),
    .A(\inv_in[188] ));
 sg13g2_inv_2 \inv[1890]/_0_  (.Y(\inv_in[1891] ),
    .A(\inv_in[1890] ));
 sg13g2_inv_2 \inv[1891]/_0_  (.Y(\inv_in[1892] ),
    .A(\inv_in[1891] ));
 sg13g2_inv_2 \inv[1892]/_0_  (.Y(\inv_in[1893] ),
    .A(\inv_in[1892] ));
 sg13g2_inv_2 \inv[1893]/_0_  (.Y(\inv_in[1894] ),
    .A(\inv_in[1893] ));
 sg13g2_inv_2 \inv[1894]/_0_  (.Y(\inv_in[1895] ),
    .A(\inv_in[1894] ));
 sg13g2_inv_2 \inv[1895]/_0_  (.Y(\inv_in[1896] ),
    .A(\inv_in[1895] ));
 sg13g2_inv_2 \inv[1896]/_0_  (.Y(\inv_in[1897] ),
    .A(\inv_in[1896] ));
 sg13g2_inv_2 \inv[1897]/_0_  (.Y(\inv_in[1898] ),
    .A(\inv_in[1897] ));
 sg13g2_inv_2 \inv[1898]/_0_  (.Y(\inv_in[1899] ),
    .A(\inv_in[1898] ));
 sg13g2_inv_2 \inv[1899]/_0_  (.Y(\inv_in[1900] ),
    .A(\inv_in[1899] ));
 sg13g2_inv_2 \inv[189]/_0_  (.Y(\inv_in[190] ),
    .A(\inv_in[189] ));
 sg13g2_inv_2 \inv[18]/_0_  (.Y(\inv_in[19] ),
    .A(\inv_in[18] ));
 sg13g2_inv_2 \inv[1900]/_0_  (.Y(\inv_in[1901] ),
    .A(\inv_in[1900] ));
 sg13g2_inv_2 \inv[1901]/_0_  (.Y(\inv_in[1902] ),
    .A(\inv_in[1901] ));
 sg13g2_inv_2 \inv[1902]/_0_  (.Y(\inv_in[1903] ),
    .A(\inv_in[1902] ));
 sg13g2_inv_2 \inv[1903]/_0_  (.Y(\inv_in[1904] ),
    .A(\inv_in[1903] ));
 sg13g2_inv_2 \inv[1904]/_0_  (.Y(\inv_in[1905] ),
    .A(\inv_in[1904] ));
 sg13g2_inv_2 \inv[1905]/_0_  (.Y(\inv_in[1906] ),
    .A(\inv_in[1905] ));
 sg13g2_inv_2 \inv[1906]/_0_  (.Y(\inv_in[1907] ),
    .A(\inv_in[1906] ));
 sg13g2_inv_2 \inv[1907]/_0_  (.Y(\inv_in[1908] ),
    .A(\inv_in[1907] ));
 sg13g2_inv_2 \inv[1908]/_0_  (.Y(\inv_in[1909] ),
    .A(\inv_in[1908] ));
 sg13g2_inv_2 \inv[1909]/_0_  (.Y(\inv_in[1910] ),
    .A(\inv_in[1909] ));
 sg13g2_inv_2 \inv[190]/_0_  (.Y(\inv_in[191] ),
    .A(\inv_in[190] ));
 sg13g2_inv_2 \inv[1910]/_0_  (.Y(\inv_in[1911] ),
    .A(\inv_in[1910] ));
 sg13g2_inv_2 \inv[1911]/_0_  (.Y(\inv_in[1912] ),
    .A(\inv_in[1911] ));
 sg13g2_inv_2 \inv[1912]/_0_  (.Y(\inv_in[1913] ),
    .A(\inv_in[1912] ));
 sg13g2_inv_2 \inv[1913]/_0_  (.Y(\inv_in[1914] ),
    .A(\inv_in[1913] ));
 sg13g2_inv_2 \inv[1914]/_0_  (.Y(\inv_in[1915] ),
    .A(\inv_in[1914] ));
 sg13g2_inv_2 \inv[1915]/_0_  (.Y(\inv_in[1916] ),
    .A(\inv_in[1915] ));
 sg13g2_inv_2 \inv[1916]/_0_  (.Y(\inv_in[1917] ),
    .A(\inv_in[1916] ));
 sg13g2_inv_2 \inv[1917]/_0_  (.Y(\inv_in[1918] ),
    .A(\inv_in[1917] ));
 sg13g2_inv_2 \inv[1918]/_0_  (.Y(\inv_in[1919] ),
    .A(\inv_in[1918] ));
 sg13g2_inv_2 \inv[1919]/_0_  (.Y(\inv_in[1920] ),
    .A(\inv_in[1919] ));
 sg13g2_inv_2 \inv[191]/_0_  (.Y(\inv_in[192] ),
    .A(\inv_in[191] ));
 sg13g2_inv_2 \inv[1920]/_0_  (.Y(\inv_in[1921] ),
    .A(\inv_in[1920] ));
 sg13g2_inv_2 \inv[1921]/_0_  (.Y(\inv_in[1922] ),
    .A(\inv_in[1921] ));
 sg13g2_inv_2 \inv[1922]/_0_  (.Y(\inv_in[1923] ),
    .A(\inv_in[1922] ));
 sg13g2_inv_2 \inv[1923]/_0_  (.Y(\inv_in[1924] ),
    .A(\inv_in[1923] ));
 sg13g2_inv_2 \inv[1924]/_0_  (.Y(\inv_in[1925] ),
    .A(\inv_in[1924] ));
 sg13g2_inv_2 \inv[1925]/_0_  (.Y(\inv_in[1926] ),
    .A(\inv_in[1925] ));
 sg13g2_inv_2 \inv[1926]/_0_  (.Y(\inv_in[1927] ),
    .A(\inv_in[1926] ));
 sg13g2_inv_2 \inv[1927]/_0_  (.Y(\inv_in[1928] ),
    .A(\inv_in[1927] ));
 sg13g2_inv_2 \inv[1928]/_0_  (.Y(\inv_in[1929] ),
    .A(\inv_in[1928] ));
 sg13g2_inv_2 \inv[1929]/_0_  (.Y(\inv_in[1930] ),
    .A(\inv_in[1929] ));
 sg13g2_inv_2 \inv[192]/_0_  (.Y(\inv_in[193] ),
    .A(\inv_in[192] ));
 sg13g2_inv_2 \inv[1930]/_0_  (.Y(\inv_in[1931] ),
    .A(\inv_in[1930] ));
 sg13g2_inv_2 \inv[1931]/_0_  (.Y(\inv_in[1932] ),
    .A(\inv_in[1931] ));
 sg13g2_inv_2 \inv[1932]/_0_  (.Y(\inv_in[1933] ),
    .A(\inv_in[1932] ));
 sg13g2_inv_2 \inv[1933]/_0_  (.Y(\inv_in[1934] ),
    .A(\inv_in[1933] ));
 sg13g2_inv_2 \inv[1934]/_0_  (.Y(\inv_in[1935] ),
    .A(\inv_in[1934] ));
 sg13g2_inv_2 \inv[1935]/_0_  (.Y(\inv_in[1936] ),
    .A(\inv_in[1935] ));
 sg13g2_inv_2 \inv[1936]/_0_  (.Y(\inv_in[1937] ),
    .A(\inv_in[1936] ));
 sg13g2_inv_2 \inv[1937]/_0_  (.Y(\inv_in[1938] ),
    .A(\inv_in[1937] ));
 sg13g2_inv_2 \inv[1938]/_0_  (.Y(\inv_in[1939] ),
    .A(\inv_in[1938] ));
 sg13g2_inv_2 \inv[1939]/_0_  (.Y(\inv_in[1940] ),
    .A(\inv_in[1939] ));
 sg13g2_inv_2 \inv[193]/_0_  (.Y(\inv_in[194] ),
    .A(\inv_in[193] ));
 sg13g2_inv_2 \inv[1940]/_0_  (.Y(\inv_in[1941] ),
    .A(\inv_in[1940] ));
 sg13g2_inv_2 \inv[1941]/_0_  (.Y(\inv_in[1942] ),
    .A(\inv_in[1941] ));
 sg13g2_inv_2 \inv[1942]/_0_  (.Y(\inv_in[1943] ),
    .A(\inv_in[1942] ));
 sg13g2_inv_2 \inv[1943]/_0_  (.Y(\inv_in[1944] ),
    .A(\inv_in[1943] ));
 sg13g2_inv_2 \inv[1944]/_0_  (.Y(\inv_in[1945] ),
    .A(\inv_in[1944] ));
 sg13g2_inv_2 \inv[1945]/_0_  (.Y(\inv_in[1946] ),
    .A(\inv_in[1945] ));
 sg13g2_inv_2 \inv[1946]/_0_  (.Y(\inv_in[1947] ),
    .A(\inv_in[1946] ));
 sg13g2_inv_2 \inv[1947]/_0_  (.Y(\inv_in[1948] ),
    .A(\inv_in[1947] ));
 sg13g2_inv_2 \inv[1948]/_0_  (.Y(\inv_in[1949] ),
    .A(\inv_in[1948] ));
 sg13g2_inv_2 \inv[1949]/_0_  (.Y(\inv_in[1950] ),
    .A(\inv_in[1949] ));
 sg13g2_inv_2 \inv[194]/_0_  (.Y(\inv_in[195] ),
    .A(\inv_in[194] ));
 sg13g2_inv_2 \inv[1950]/_0_  (.Y(\inv_in[1951] ),
    .A(\inv_in[1950] ));
 sg13g2_inv_2 \inv[1951]/_0_  (.Y(\inv_in[1952] ),
    .A(\inv_in[1951] ));
 sg13g2_inv_2 \inv[1952]/_0_  (.Y(\inv_in[1953] ),
    .A(\inv_in[1952] ));
 sg13g2_inv_2 \inv[1953]/_0_  (.Y(\inv_in[1954] ),
    .A(\inv_in[1953] ));
 sg13g2_inv_2 \inv[1954]/_0_  (.Y(\inv_in[1955] ),
    .A(\inv_in[1954] ));
 sg13g2_inv_2 \inv[1955]/_0_  (.Y(\inv_in[1956] ),
    .A(\inv_in[1955] ));
 sg13g2_inv_2 \inv[1956]/_0_  (.Y(\inv_in[1957] ),
    .A(\inv_in[1956] ));
 sg13g2_inv_2 \inv[1957]/_0_  (.Y(\inv_in[1958] ),
    .A(\inv_in[1957] ));
 sg13g2_inv_2 \inv[1958]/_0_  (.Y(\inv_in[1959] ),
    .A(\inv_in[1958] ));
 sg13g2_inv_2 \inv[1959]/_0_  (.Y(\inv_in[1960] ),
    .A(\inv_in[1959] ));
 sg13g2_inv_2 \inv[195]/_0_  (.Y(\inv_in[196] ),
    .A(\inv_in[195] ));
 sg13g2_inv_2 \inv[1960]/_0_  (.Y(\inv_in[1961] ),
    .A(\inv_in[1960] ));
 sg13g2_inv_2 \inv[1961]/_0_  (.Y(\inv_in[1962] ),
    .A(\inv_in[1961] ));
 sg13g2_inv_2 \inv[1962]/_0_  (.Y(\inv_in[1963] ),
    .A(\inv_in[1962] ));
 sg13g2_inv_2 \inv[1963]/_0_  (.Y(\inv_in[1964] ),
    .A(\inv_in[1963] ));
 sg13g2_inv_2 \inv[1964]/_0_  (.Y(\inv_in[1965] ),
    .A(\inv_in[1964] ));
 sg13g2_inv_2 \inv[1965]/_0_  (.Y(\inv_in[1966] ),
    .A(\inv_in[1965] ));
 sg13g2_inv_2 \inv[1966]/_0_  (.Y(\inv_in[1967] ),
    .A(\inv_in[1966] ));
 sg13g2_inv_2 \inv[1967]/_0_  (.Y(\inv_in[1968] ),
    .A(\inv_in[1967] ));
 sg13g2_inv_2 \inv[1968]/_0_  (.Y(\inv_in[1969] ),
    .A(\inv_in[1968] ));
 sg13g2_inv_2 \inv[1969]/_0_  (.Y(\inv_in[1970] ),
    .A(\inv_in[1969] ));
 sg13g2_inv_2 \inv[196]/_0_  (.Y(\inv_in[197] ),
    .A(\inv_in[196] ));
 sg13g2_inv_2 \inv[1970]/_0_  (.Y(\inv_in[1971] ),
    .A(\inv_in[1970] ));
 sg13g2_inv_2 \inv[1971]/_0_  (.Y(\inv_in[1972] ),
    .A(\inv_in[1971] ));
 sg13g2_inv_2 \inv[1972]/_0_  (.Y(\inv_in[1973] ),
    .A(\inv_in[1972] ));
 sg13g2_inv_2 \inv[1973]/_0_  (.Y(\inv_in[1974] ),
    .A(\inv_in[1973] ));
 sg13g2_inv_2 \inv[1974]/_0_  (.Y(\inv_in[1975] ),
    .A(\inv_in[1974] ));
 sg13g2_inv_2 \inv[1975]/_0_  (.Y(\inv_in[1976] ),
    .A(\inv_in[1975] ));
 sg13g2_inv_2 \inv[1976]/_0_  (.Y(\inv_in[1977] ),
    .A(\inv_in[1976] ));
 sg13g2_inv_2 \inv[1977]/_0_  (.Y(\inv_in[1978] ),
    .A(\inv_in[1977] ));
 sg13g2_inv_2 \inv[1978]/_0_  (.Y(\inv_in[1979] ),
    .A(\inv_in[1978] ));
 sg13g2_inv_2 \inv[1979]/_0_  (.Y(\inv_in[1980] ),
    .A(\inv_in[1979] ));
 sg13g2_inv_2 \inv[197]/_0_  (.Y(\inv_in[198] ),
    .A(\inv_in[197] ));
 sg13g2_inv_2 \inv[1980]/_0_  (.Y(\inv_in[1981] ),
    .A(\inv_in[1980] ));
 sg13g2_inv_2 \inv[1981]/_0_  (.Y(\inv_in[1982] ),
    .A(\inv_in[1981] ));
 sg13g2_inv_2 \inv[1982]/_0_  (.Y(\inv_in[1983] ),
    .A(\inv_in[1982] ));
 sg13g2_inv_2 \inv[1983]/_0_  (.Y(\inv_in[1984] ),
    .A(\inv_in[1983] ));
 sg13g2_inv_2 \inv[1984]/_0_  (.Y(\inv_in[1985] ),
    .A(\inv_in[1984] ));
 sg13g2_inv_2 \inv[1985]/_0_  (.Y(\inv_in[1986] ),
    .A(\inv_in[1985] ));
 sg13g2_inv_2 \inv[1986]/_0_  (.Y(\inv_in[1987] ),
    .A(\inv_in[1986] ));
 sg13g2_inv_2 \inv[1987]/_0_  (.Y(\inv_in[1988] ),
    .A(\inv_in[1987] ));
 sg13g2_inv_2 \inv[1988]/_0_  (.Y(\inv_in[1989] ),
    .A(\inv_in[1988] ));
 sg13g2_inv_2 \inv[1989]/_0_  (.Y(\inv_in[1990] ),
    .A(\inv_in[1989] ));
 sg13g2_inv_2 \inv[198]/_0_  (.Y(\inv_in[199] ),
    .A(\inv_in[198] ));
 sg13g2_inv_2 \inv[1990]/_0_  (.Y(\inv_in[1991] ),
    .A(\inv_in[1990] ));
 sg13g2_inv_2 \inv[1991]/_0_  (.Y(\inv_in[1992] ),
    .A(\inv_in[1991] ));
 sg13g2_inv_2 \inv[1992]/_0_  (.Y(\inv_in[1993] ),
    .A(\inv_in[1992] ));
 sg13g2_inv_2 \inv[1993]/_0_  (.Y(\inv_in[1994] ),
    .A(\inv_in[1993] ));
 sg13g2_inv_2 \inv[1994]/_0_  (.Y(\inv_in[1995] ),
    .A(\inv_in[1994] ));
 sg13g2_inv_2 \inv[1995]/_0_  (.Y(\inv_in[1996] ),
    .A(\inv_in[1995] ));
 sg13g2_inv_2 \inv[1996]/_0_  (.Y(\inv_in[1997] ),
    .A(\inv_in[1996] ));
 sg13g2_inv_2 \inv[1997]/_0_  (.Y(\inv_in[1998] ),
    .A(\inv_in[1997] ));
 sg13g2_inv_2 \inv[1998]/_0_  (.Y(\inv_in[1999] ),
    .A(\inv_in[1998] ));
 sg13g2_inv_2 \inv[1999]/_0_  (.Y(\inv_in[2000] ),
    .A(\inv_in[1999] ));
 sg13g2_inv_2 \inv[199]/_0_  (.Y(\inv_in[200] ),
    .A(\inv_in[199] ));
 sg13g2_inv_2 \inv[19]/_0_  (.Y(\inv_in[20] ),
    .A(\inv_in[19] ));
 sg13g2_inv_8 \inv[1]/_0_  (.Y(\inv_in[2] ),
    .A(\inv_in[1] ));
 sg13g2_inv_2 \inv[2000]/_0_  (.Y(\inv_in[2001] ),
    .A(\inv_in[2000] ));
 sg13g2_inv_2 \inv[2001]/_0_  (.Y(\inv_in[2002] ),
    .A(\inv_in[2001] ));
 sg13g2_inv_2 \inv[2002]/_0_  (.Y(\inv_in[2003] ),
    .A(\inv_in[2002] ));
 sg13g2_inv_2 \inv[2003]/_0_  (.Y(\inv_in[2004] ),
    .A(\inv_in[2003] ));
 sg13g2_inv_2 \inv[2004]/_0_  (.Y(\inv_in[2005] ),
    .A(\inv_in[2004] ));
 sg13g2_inv_2 \inv[2005]/_0_  (.Y(\inv_in[2006] ),
    .A(\inv_in[2005] ));
 sg13g2_inv_2 \inv[2006]/_0_  (.Y(\inv_in[2007] ),
    .A(\inv_in[2006] ));
 sg13g2_inv_2 \inv[2007]/_0_  (.Y(\inv_in[2008] ),
    .A(\inv_in[2007] ));
 sg13g2_inv_2 \inv[2008]/_0_  (.Y(\inv_in[2009] ),
    .A(\inv_in[2008] ));
 sg13g2_inv_2 \inv[2009]/_0_  (.Y(\inv_in[2010] ),
    .A(\inv_in[2009] ));
 sg13g2_inv_2 \inv[200]/_0_  (.Y(\inv_in[201] ),
    .A(\inv_in[200] ));
 sg13g2_inv_2 \inv[2010]/_0_  (.Y(\inv_in[2011] ),
    .A(\inv_in[2010] ));
 sg13g2_inv_2 \inv[2011]/_0_  (.Y(\inv_in[2012] ),
    .A(\inv_in[2011] ));
 sg13g2_inv_2 \inv[2012]/_0_  (.Y(\inv_in[2013] ),
    .A(\inv_in[2012] ));
 sg13g2_inv_2 \inv[2013]/_0_  (.Y(\inv_in[2014] ),
    .A(\inv_in[2013] ));
 sg13g2_inv_2 \inv[2014]/_0_  (.Y(\inv_in[2015] ),
    .A(\inv_in[2014] ));
 sg13g2_inv_2 \inv[2015]/_0_  (.Y(\inv_in[2016] ),
    .A(\inv_in[2015] ));
 sg13g2_inv_2 \inv[2016]/_0_  (.Y(\inv_in[2017] ),
    .A(\inv_in[2016] ));
 sg13g2_inv_2 \inv[2017]/_0_  (.Y(\inv_in[2018] ),
    .A(\inv_in[2017] ));
 sg13g2_inv_2 \inv[2018]/_0_  (.Y(\inv_in[2019] ),
    .A(\inv_in[2018] ));
 sg13g2_inv_2 \inv[2019]/_0_  (.Y(\inv_in[2020] ),
    .A(\inv_in[2019] ));
 sg13g2_inv_2 \inv[201]/_0_  (.Y(\inv_in[202] ),
    .A(\inv_in[201] ));
 sg13g2_inv_2 \inv[2020]/_0_  (.Y(\inv_in[2021] ),
    .A(\inv_in[2020] ));
 sg13g2_inv_2 \inv[2021]/_0_  (.Y(\inv_in[2022] ),
    .A(\inv_in[2021] ));
 sg13g2_inv_2 \inv[2022]/_0_  (.Y(\inv_in[2023] ),
    .A(\inv_in[2022] ));
 sg13g2_inv_2 \inv[2023]/_0_  (.Y(\inv_in[2024] ),
    .A(\inv_in[2023] ));
 sg13g2_inv_2 \inv[2024]/_0_  (.Y(\inv_in[2025] ),
    .A(\inv_in[2024] ));
 sg13g2_inv_2 \inv[2025]/_0_  (.Y(\inv_in[2026] ),
    .A(\inv_in[2025] ));
 sg13g2_inv_2 \inv[2026]/_0_  (.Y(\inv_in[2027] ),
    .A(\inv_in[2026] ));
 sg13g2_inv_2 \inv[2027]/_0_  (.Y(\inv_in[2028] ),
    .A(\inv_in[2027] ));
 sg13g2_inv_2 \inv[2028]/_0_  (.Y(\inv_in[2029] ),
    .A(\inv_in[2028] ));
 sg13g2_inv_2 \inv[2029]/_0_  (.Y(\inv_in[2030] ),
    .A(\inv_in[2029] ));
 sg13g2_inv_2 \inv[202]/_0_  (.Y(\inv_in[203] ),
    .A(\inv_in[202] ));
 sg13g2_inv_2 \inv[2030]/_0_  (.Y(\inv_in[2031] ),
    .A(\inv_in[2030] ));
 sg13g2_inv_2 \inv[2031]/_0_  (.Y(\inv_in[2032] ),
    .A(\inv_in[2031] ));
 sg13g2_inv_2 \inv[2032]/_0_  (.Y(\inv_in[2033] ),
    .A(\inv_in[2032] ));
 sg13g2_inv_2 \inv[2033]/_0_  (.Y(\inv_in[2034] ),
    .A(\inv_in[2033] ));
 sg13g2_inv_2 \inv[2034]/_0_  (.Y(\inv_in[2035] ),
    .A(\inv_in[2034] ));
 sg13g2_inv_2 \inv[2035]/_0_  (.Y(\inv_in[2036] ),
    .A(\inv_in[2035] ));
 sg13g2_inv_2 \inv[2036]/_0_  (.Y(\inv_in[2037] ),
    .A(\inv_in[2036] ));
 sg13g2_inv_2 \inv[2037]/_0_  (.Y(\inv_in[2038] ),
    .A(\inv_in[2037] ));
 sg13g2_inv_2 \inv[2038]/_0_  (.Y(\inv_in[2039] ),
    .A(\inv_in[2038] ));
 sg13g2_inv_2 \inv[2039]/_0_  (.Y(\inv_in[2040] ),
    .A(\inv_in[2039] ));
 sg13g2_inv_2 \inv[203]/_0_  (.Y(\inv_in[204] ),
    .A(\inv_in[203] ));
 sg13g2_inv_2 \inv[2040]/_0_  (.Y(\inv_in[2041] ),
    .A(\inv_in[2040] ));
 sg13g2_inv_2 \inv[2041]/_0_  (.Y(\inv_in[2042] ),
    .A(\inv_in[2041] ));
 sg13g2_inv_2 \inv[2042]/_0_  (.Y(\inv_in[2043] ),
    .A(\inv_in[2042] ));
 sg13g2_inv_2 \inv[2043]/_0_  (.Y(\inv_in[2044] ),
    .A(\inv_in[2043] ));
 sg13g2_inv_2 \inv[2044]/_0_  (.Y(\inv_in[2045] ),
    .A(\inv_in[2044] ));
 sg13g2_inv_2 \inv[2045]/_0_  (.Y(\inv_in[2046] ),
    .A(\inv_in[2045] ));
 sg13g2_inv_2 \inv[2046]/_0_  (.Y(\inv_in[2047] ),
    .A(\inv_in[2046] ));
 sg13g2_inv_2 \inv[2047]/_0_  (.Y(\inv_in[2048] ),
    .A(\inv_in[2047] ));
 sg13g2_inv_2 \inv[2048]/_0_  (.Y(\inv_in[2049] ),
    .A(\inv_in[2048] ));
 sg13g2_inv_2 \inv[2049]/_0_  (.Y(\inv_in[2050] ),
    .A(\inv_in[2049] ));
 sg13g2_inv_2 \inv[204]/_0_  (.Y(\inv_in[205] ),
    .A(\inv_in[204] ));
 sg13g2_inv_2 \inv[2050]/_0_  (.Y(\inv_in[2051] ),
    .A(\inv_in[2050] ));
 sg13g2_inv_2 \inv[2051]/_0_  (.Y(\inv_in[2052] ),
    .A(\inv_in[2051] ));
 sg13g2_inv_2 \inv[2052]/_0_  (.Y(\inv_in[2053] ),
    .A(\inv_in[2052] ));
 sg13g2_inv_2 \inv[2053]/_0_  (.Y(\inv_in[2054] ),
    .A(\inv_in[2053] ));
 sg13g2_inv_2 \inv[2054]/_0_  (.Y(\inv_in[2055] ),
    .A(\inv_in[2054] ));
 sg13g2_inv_2 \inv[2055]/_0_  (.Y(\inv_in[2056] ),
    .A(\inv_in[2055] ));
 sg13g2_inv_2 \inv[2056]/_0_  (.Y(\inv_in[2057] ),
    .A(\inv_in[2056] ));
 sg13g2_inv_2 \inv[2057]/_0_  (.Y(\inv_in[2058] ),
    .A(\inv_in[2057] ));
 sg13g2_inv_2 \inv[2058]/_0_  (.Y(\inv_in[2059] ),
    .A(\inv_in[2058] ));
 sg13g2_inv_2 \inv[2059]/_0_  (.Y(\inv_in[2060] ),
    .A(\inv_in[2059] ));
 sg13g2_inv_2 \inv[205]/_0_  (.Y(\inv_in[206] ),
    .A(\inv_in[205] ));
 sg13g2_inv_2 \inv[2060]/_0_  (.Y(\inv_in[2061] ),
    .A(\inv_in[2060] ));
 sg13g2_inv_2 \inv[2061]/_0_  (.Y(\inv_in[2062] ),
    .A(\inv_in[2061] ));
 sg13g2_inv_2 \inv[2062]/_0_  (.Y(\inv_in[2063] ),
    .A(\inv_in[2062] ));
 sg13g2_inv_2 \inv[2063]/_0_  (.Y(\inv_in[2064] ),
    .A(\inv_in[2063] ));
 sg13g2_inv_2 \inv[2064]/_0_  (.Y(\inv_in[2065] ),
    .A(\inv_in[2064] ));
 sg13g2_inv_2 \inv[2065]/_0_  (.Y(\inv_in[2066] ),
    .A(\inv_in[2065] ));
 sg13g2_inv_2 \inv[2066]/_0_  (.Y(\inv_in[2067] ),
    .A(\inv_in[2066] ));
 sg13g2_inv_2 \inv[2067]/_0_  (.Y(\inv_in[2068] ),
    .A(\inv_in[2067] ));
 sg13g2_inv_2 \inv[2068]/_0_  (.Y(\inv_in[2069] ),
    .A(\inv_in[2068] ));
 sg13g2_inv_2 \inv[2069]/_0_  (.Y(\inv_in[2070] ),
    .A(\inv_in[2069] ));
 sg13g2_inv_2 \inv[206]/_0_  (.Y(\inv_in[207] ),
    .A(\inv_in[206] ));
 sg13g2_inv_2 \inv[2070]/_0_  (.Y(\inv_in[2071] ),
    .A(\inv_in[2070] ));
 sg13g2_inv_2 \inv[2071]/_0_  (.Y(\inv_in[2072] ),
    .A(\inv_in[2071] ));
 sg13g2_inv_2 \inv[2072]/_0_  (.Y(\inv_in[2073] ),
    .A(\inv_in[2072] ));
 sg13g2_inv_2 \inv[2073]/_0_  (.Y(\inv_in[2074] ),
    .A(\inv_in[2073] ));
 sg13g2_inv_2 \inv[2074]/_0_  (.Y(\inv_in[2075] ),
    .A(\inv_in[2074] ));
 sg13g2_inv_2 \inv[2075]/_0_  (.Y(\inv_in[2076] ),
    .A(\inv_in[2075] ));
 sg13g2_inv_2 \inv[2076]/_0_  (.Y(\inv_in[2077] ),
    .A(\inv_in[2076] ));
 sg13g2_inv_2 \inv[2077]/_0_  (.Y(\inv_in[2078] ),
    .A(\inv_in[2077] ));
 sg13g2_inv_2 \inv[2078]/_0_  (.Y(\inv_in[2079] ),
    .A(\inv_in[2078] ));
 sg13g2_inv_2 \inv[2079]/_0_  (.Y(\inv_in[2080] ),
    .A(\inv_in[2079] ));
 sg13g2_inv_2 \inv[207]/_0_  (.Y(\inv_in[208] ),
    .A(\inv_in[207] ));
 sg13g2_inv_2 \inv[2080]/_0_  (.Y(\inv_in[2081] ),
    .A(\inv_in[2080] ));
 sg13g2_inv_2 \inv[2081]/_0_  (.Y(\inv_in[2082] ),
    .A(\inv_in[2081] ));
 sg13g2_inv_2 \inv[2082]/_0_  (.Y(\inv_in[2083] ),
    .A(\inv_in[2082] ));
 sg13g2_inv_2 \inv[2083]/_0_  (.Y(\inv_in[2084] ),
    .A(\inv_in[2083] ));
 sg13g2_inv_2 \inv[2084]/_0_  (.Y(\inv_in[2085] ),
    .A(\inv_in[2084] ));
 sg13g2_inv_2 \inv[2085]/_0_  (.Y(\inv_in[2086] ),
    .A(\inv_in[2085] ));
 sg13g2_inv_2 \inv[2086]/_0_  (.Y(\inv_in[2087] ),
    .A(\inv_in[2086] ));
 sg13g2_inv_2 \inv[2087]/_0_  (.Y(\inv_in[2088] ),
    .A(\inv_in[2087] ));
 sg13g2_inv_2 \inv[2088]/_0_  (.Y(\inv_in[2089] ),
    .A(\inv_in[2088] ));
 sg13g2_inv_2 \inv[2089]/_0_  (.Y(\inv_in[2090] ),
    .A(\inv_in[2089] ));
 sg13g2_inv_2 \inv[208]/_0_  (.Y(\inv_in[209] ),
    .A(\inv_in[208] ));
 sg13g2_inv_2 \inv[2090]/_0_  (.Y(\inv_in[2091] ),
    .A(\inv_in[2090] ));
 sg13g2_inv_2 \inv[2091]/_0_  (.Y(\inv_in[2092] ),
    .A(\inv_in[2091] ));
 sg13g2_inv_2 \inv[2092]/_0_  (.Y(\inv_in[2093] ),
    .A(\inv_in[2092] ));
 sg13g2_inv_2 \inv[2093]/_0_  (.Y(\inv_in[2094] ),
    .A(\inv_in[2093] ));
 sg13g2_inv_2 \inv[2094]/_0_  (.Y(\inv_in[2095] ),
    .A(\inv_in[2094] ));
 sg13g2_inv_2 \inv[2095]/_0_  (.Y(\inv_in[2096] ),
    .A(\inv_in[2095] ));
 sg13g2_inv_2 \inv[2096]/_0_  (.Y(\inv_in[2097] ),
    .A(\inv_in[2096] ));
 sg13g2_inv_2 \inv[2097]/_0_  (.Y(\inv_in[2098] ),
    .A(\inv_in[2097] ));
 sg13g2_inv_2 \inv[2098]/_0_  (.Y(\inv_in[2099] ),
    .A(\inv_in[2098] ));
 sg13g2_inv_2 \inv[2099]/_0_  (.Y(\inv_in[2100] ),
    .A(\inv_in[2099] ));
 sg13g2_inv_2 \inv[209]/_0_  (.Y(\inv_in[210] ),
    .A(\inv_in[209] ));
 sg13g2_inv_2 \inv[20]/_0_  (.Y(\inv_in[21] ),
    .A(\inv_in[20] ));
 sg13g2_inv_2 \inv[2100]/_0_  (.Y(\inv_in[2101] ),
    .A(\inv_in[2100] ));
 sg13g2_inv_2 \inv[2101]/_0_  (.Y(\inv_in[2102] ),
    .A(\inv_in[2101] ));
 sg13g2_inv_2 \inv[2102]/_0_  (.Y(\inv_in[2103] ),
    .A(\inv_in[2102] ));
 sg13g2_inv_2 \inv[2103]/_0_  (.Y(\inv_in[2104] ),
    .A(\inv_in[2103] ));
 sg13g2_inv_2 \inv[2104]/_0_  (.Y(\inv_in[2105] ),
    .A(\inv_in[2104] ));
 sg13g2_inv_2 \inv[2105]/_0_  (.Y(\inv_in[2106] ),
    .A(\inv_in[2105] ));
 sg13g2_inv_2 \inv[2106]/_0_  (.Y(\inv_in[2107] ),
    .A(\inv_in[2106] ));
 sg13g2_inv_2 \inv[2107]/_0_  (.Y(\inv_in[2108] ),
    .A(\inv_in[2107] ));
 sg13g2_inv_2 \inv[2108]/_0_  (.Y(\inv_in[2109] ),
    .A(\inv_in[2108] ));
 sg13g2_inv_2 \inv[2109]/_0_  (.Y(\inv_in[2110] ),
    .A(\inv_in[2109] ));
 sg13g2_inv_2 \inv[210]/_0_  (.Y(\inv_in[211] ),
    .A(\inv_in[210] ));
 sg13g2_inv_2 \inv[2110]/_0_  (.Y(\inv_in[2111] ),
    .A(\inv_in[2110] ));
 sg13g2_inv_2 \inv[2111]/_0_  (.Y(\inv_in[2112] ),
    .A(\inv_in[2111] ));
 sg13g2_inv_2 \inv[2112]/_0_  (.Y(\inv_in[2113] ),
    .A(\inv_in[2112] ));
 sg13g2_inv_2 \inv[2113]/_0_  (.Y(\inv_in[2114] ),
    .A(\inv_in[2113] ));
 sg13g2_inv_2 \inv[2114]/_0_  (.Y(\inv_in[2115] ),
    .A(\inv_in[2114] ));
 sg13g2_inv_2 \inv[2115]/_0_  (.Y(\inv_in[2116] ),
    .A(\inv_in[2115] ));
 sg13g2_inv_2 \inv[2116]/_0_  (.Y(\inv_in[2117] ),
    .A(\inv_in[2116] ));
 sg13g2_inv_2 \inv[2117]/_0_  (.Y(\inv_in[2118] ),
    .A(\inv_in[2117] ));
 sg13g2_inv_2 \inv[2118]/_0_  (.Y(\inv_in[2119] ),
    .A(\inv_in[2118] ));
 sg13g2_inv_2 \inv[2119]/_0_  (.Y(\inv_in[2120] ),
    .A(\inv_in[2119] ));
 sg13g2_inv_2 \inv[211]/_0_  (.Y(\inv_in[212] ),
    .A(\inv_in[211] ));
 sg13g2_inv_2 \inv[2120]/_0_  (.Y(\inv_in[2121] ),
    .A(\inv_in[2120] ));
 sg13g2_inv_2 \inv[2121]/_0_  (.Y(\inv_in[2122] ),
    .A(\inv_in[2121] ));
 sg13g2_inv_2 \inv[2122]/_0_  (.Y(\inv_in[2123] ),
    .A(\inv_in[2122] ));
 sg13g2_inv_2 \inv[2123]/_0_  (.Y(\inv_in[2124] ),
    .A(\inv_in[2123] ));
 sg13g2_inv_2 \inv[2124]/_0_  (.Y(\inv_in[2125] ),
    .A(\inv_in[2124] ));
 sg13g2_inv_2 \inv[2125]/_0_  (.Y(\inv_in[2126] ),
    .A(\inv_in[2125] ));
 sg13g2_inv_2 \inv[2126]/_0_  (.Y(\inv_in[2127] ),
    .A(\inv_in[2126] ));
 sg13g2_inv_2 \inv[2127]/_0_  (.Y(\inv_in[2128] ),
    .A(\inv_in[2127] ));
 sg13g2_inv_2 \inv[2128]/_0_  (.Y(\inv_in[2129] ),
    .A(\inv_in[2128] ));
 sg13g2_inv_2 \inv[2129]/_0_  (.Y(\inv_in[2130] ),
    .A(\inv_in[2129] ));
 sg13g2_inv_2 \inv[212]/_0_  (.Y(\inv_in[213] ),
    .A(\inv_in[212] ));
 sg13g2_inv_2 \inv[2130]/_0_  (.Y(\inv_in[2131] ),
    .A(\inv_in[2130] ));
 sg13g2_inv_2 \inv[2131]/_0_  (.Y(\inv_in[2132] ),
    .A(\inv_in[2131] ));
 sg13g2_inv_2 \inv[2132]/_0_  (.Y(\inv_in[2133] ),
    .A(\inv_in[2132] ));
 sg13g2_inv_2 \inv[2133]/_0_  (.Y(\inv_in[2134] ),
    .A(\inv_in[2133] ));
 sg13g2_inv_2 \inv[2134]/_0_  (.Y(\inv_in[2135] ),
    .A(\inv_in[2134] ));
 sg13g2_inv_2 \inv[2135]/_0_  (.Y(\inv_in[2136] ),
    .A(\inv_in[2135] ));
 sg13g2_inv_2 \inv[2136]/_0_  (.Y(\inv_in[2137] ),
    .A(\inv_in[2136] ));
 sg13g2_inv_2 \inv[2137]/_0_  (.Y(\inv_in[2138] ),
    .A(\inv_in[2137] ));
 sg13g2_inv_2 \inv[2138]/_0_  (.Y(\inv_in[2139] ),
    .A(\inv_in[2138] ));
 sg13g2_inv_2 \inv[2139]/_0_  (.Y(\inv_in[2140] ),
    .A(\inv_in[2139] ));
 sg13g2_inv_2 \inv[213]/_0_  (.Y(\inv_in[214] ),
    .A(\inv_in[213] ));
 sg13g2_inv_2 \inv[2140]/_0_  (.Y(\inv_in[2141] ),
    .A(\inv_in[2140] ));
 sg13g2_inv_2 \inv[2141]/_0_  (.Y(\inv_in[2142] ),
    .A(\inv_in[2141] ));
 sg13g2_inv_2 \inv[2142]/_0_  (.Y(\inv_in[2143] ),
    .A(\inv_in[2142] ));
 sg13g2_inv_2 \inv[2143]/_0_  (.Y(\inv_in[2144] ),
    .A(\inv_in[2143] ));
 sg13g2_inv_2 \inv[2144]/_0_  (.Y(\inv_in[2145] ),
    .A(\inv_in[2144] ));
 sg13g2_inv_2 \inv[2145]/_0_  (.Y(\inv_in[2146] ),
    .A(\inv_in[2145] ));
 sg13g2_inv_2 \inv[2146]/_0_  (.Y(\inv_in[2147] ),
    .A(\inv_in[2146] ));
 sg13g2_inv_2 \inv[2147]/_0_  (.Y(\inv_in[2148] ),
    .A(\inv_in[2147] ));
 sg13g2_inv_2 \inv[2148]/_0_  (.Y(\inv_in[2149] ),
    .A(\inv_in[2148] ));
 sg13g2_inv_2 \inv[2149]/_0_  (.Y(\inv_in[2150] ),
    .A(\inv_in[2149] ));
 sg13g2_inv_2 \inv[214]/_0_  (.Y(\inv_in[215] ),
    .A(\inv_in[214] ));
 sg13g2_inv_2 \inv[2150]/_0_  (.Y(\inv_in[2151] ),
    .A(\inv_in[2150] ));
 sg13g2_inv_2 \inv[2151]/_0_  (.Y(\inv_in[2152] ),
    .A(\inv_in[2151] ));
 sg13g2_inv_2 \inv[2152]/_0_  (.Y(\inv_in[2153] ),
    .A(\inv_in[2152] ));
 sg13g2_inv_2 \inv[2153]/_0_  (.Y(\inv_in[2154] ),
    .A(\inv_in[2153] ));
 sg13g2_inv_2 \inv[2154]/_0_  (.Y(\inv_in[2155] ),
    .A(\inv_in[2154] ));
 sg13g2_inv_2 \inv[2155]/_0_  (.Y(\inv_in[2156] ),
    .A(\inv_in[2155] ));
 sg13g2_inv_2 \inv[2156]/_0_  (.Y(\inv_in[2157] ),
    .A(\inv_in[2156] ));
 sg13g2_inv_2 \inv[2157]/_0_  (.Y(\inv_in[2158] ),
    .A(\inv_in[2157] ));
 sg13g2_inv_2 \inv[2158]/_0_  (.Y(\inv_in[2159] ),
    .A(\inv_in[2158] ));
 sg13g2_inv_2 \inv[2159]/_0_  (.Y(\inv_in[2160] ),
    .A(\inv_in[2159] ));
 sg13g2_inv_2 \inv[215]/_0_  (.Y(\inv_in[216] ),
    .A(\inv_in[215] ));
 sg13g2_inv_2 \inv[2160]/_0_  (.Y(\inv_in[2161] ),
    .A(\inv_in[2160] ));
 sg13g2_inv_2 \inv[2161]/_0_  (.Y(\inv_in[2162] ),
    .A(\inv_in[2161] ));
 sg13g2_inv_2 \inv[2162]/_0_  (.Y(\inv_in[2163] ),
    .A(\inv_in[2162] ));
 sg13g2_inv_2 \inv[2163]/_0_  (.Y(\inv_in[2164] ),
    .A(\inv_in[2163] ));
 sg13g2_inv_2 \inv[2164]/_0_  (.Y(\inv_in[2165] ),
    .A(\inv_in[2164] ));
 sg13g2_inv_2 \inv[2165]/_0_  (.Y(\inv_in[2166] ),
    .A(\inv_in[2165] ));
 sg13g2_inv_2 \inv[2166]/_0_  (.Y(\inv_in[2167] ),
    .A(\inv_in[2166] ));
 sg13g2_inv_2 \inv[2167]/_0_  (.Y(\inv_in[2168] ),
    .A(\inv_in[2167] ));
 sg13g2_inv_2 \inv[2168]/_0_  (.Y(\inv_in[2169] ),
    .A(\inv_in[2168] ));
 sg13g2_inv_2 \inv[2169]/_0_  (.Y(\inv_in[2170] ),
    .A(\inv_in[2169] ));
 sg13g2_inv_2 \inv[216]/_0_  (.Y(\inv_in[217] ),
    .A(\inv_in[216] ));
 sg13g2_inv_2 \inv[2170]/_0_  (.Y(\inv_in[2171] ),
    .A(\inv_in[2170] ));
 sg13g2_inv_2 \inv[2171]/_0_  (.Y(\inv_in[2172] ),
    .A(\inv_in[2171] ));
 sg13g2_inv_2 \inv[2172]/_0_  (.Y(\inv_in[2173] ),
    .A(\inv_in[2172] ));
 sg13g2_inv_2 \inv[2173]/_0_  (.Y(\inv_in[2174] ),
    .A(\inv_in[2173] ));
 sg13g2_inv_2 \inv[2174]/_0_  (.Y(\inv_in[2175] ),
    .A(\inv_in[2174] ));
 sg13g2_inv_2 \inv[2175]/_0_  (.Y(\inv_in[2176] ),
    .A(\inv_in[2175] ));
 sg13g2_inv_2 \inv[2176]/_0_  (.Y(\inv_in[2177] ),
    .A(\inv_in[2176] ));
 sg13g2_inv_2 \inv[2177]/_0_  (.Y(\inv_in[2178] ),
    .A(\inv_in[2177] ));
 sg13g2_inv_2 \inv[2178]/_0_  (.Y(\inv_in[2179] ),
    .A(\inv_in[2178] ));
 sg13g2_inv_2 \inv[2179]/_0_  (.Y(\inv_in[2180] ),
    .A(\inv_in[2179] ));
 sg13g2_inv_2 \inv[217]/_0_  (.Y(\inv_in[218] ),
    .A(\inv_in[217] ));
 sg13g2_inv_2 \inv[2180]/_0_  (.Y(\inv_in[2181] ),
    .A(\inv_in[2180] ));
 sg13g2_inv_2 \inv[2181]/_0_  (.Y(\inv_in[2182] ),
    .A(\inv_in[2181] ));
 sg13g2_inv_2 \inv[2182]/_0_  (.Y(\inv_in[2183] ),
    .A(\inv_in[2182] ));
 sg13g2_inv_2 \inv[2183]/_0_  (.Y(\inv_in[2184] ),
    .A(\inv_in[2183] ));
 sg13g2_inv_2 \inv[2184]/_0_  (.Y(\inv_in[2185] ),
    .A(\inv_in[2184] ));
 sg13g2_inv_2 \inv[2185]/_0_  (.Y(\inv_in[2186] ),
    .A(\inv_in[2185] ));
 sg13g2_inv_2 \inv[2186]/_0_  (.Y(\inv_in[2187] ),
    .A(\inv_in[2186] ));
 sg13g2_inv_2 \inv[2187]/_0_  (.Y(\inv_in[2188] ),
    .A(\inv_in[2187] ));
 sg13g2_inv_2 \inv[2188]/_0_  (.Y(\inv_in[2189] ),
    .A(\inv_in[2188] ));
 sg13g2_inv_2 \inv[2189]/_0_  (.Y(\inv_in[2190] ),
    .A(\inv_in[2189] ));
 sg13g2_inv_2 \inv[218]/_0_  (.Y(\inv_in[219] ),
    .A(\inv_in[218] ));
 sg13g2_inv_2 \inv[2190]/_0_  (.Y(\inv_in[2191] ),
    .A(\inv_in[2190] ));
 sg13g2_inv_2 \inv[2191]/_0_  (.Y(\inv_in[2192] ),
    .A(\inv_in[2191] ));
 sg13g2_inv_2 \inv[2192]/_0_  (.Y(\inv_in[2193] ),
    .A(\inv_in[2192] ));
 sg13g2_inv_2 \inv[2193]/_0_  (.Y(\inv_in[2194] ),
    .A(\inv_in[2193] ));
 sg13g2_inv_2 \inv[2194]/_0_  (.Y(\inv_in[2195] ),
    .A(\inv_in[2194] ));
 sg13g2_inv_2 \inv[2195]/_0_  (.Y(\inv_in[2196] ),
    .A(\inv_in[2195] ));
 sg13g2_inv_2 \inv[2196]/_0_  (.Y(\inv_in[2197] ),
    .A(\inv_in[2196] ));
 sg13g2_inv_2 \inv[2197]/_0_  (.Y(\inv_in[2198] ),
    .A(\inv_in[2197] ));
 sg13g2_inv_2 \inv[2198]/_0_  (.Y(\inv_in[2199] ),
    .A(\inv_in[2198] ));
 sg13g2_inv_2 \inv[2199]/_0_  (.Y(\inv_in[2200] ),
    .A(\inv_in[2199] ));
 sg13g2_inv_2 \inv[219]/_0_  (.Y(\inv_in[220] ),
    .A(\inv_in[219] ));
 sg13g2_inv_2 \inv[21]/_0_  (.Y(\inv_in[22] ),
    .A(\inv_in[21] ));
 sg13g2_inv_2 \inv[2200]/_0_  (.Y(\inv_in[2201] ),
    .A(\inv_in[2200] ));
 sg13g2_inv_2 \inv[2201]/_0_  (.Y(\inv_in[2202] ),
    .A(\inv_in[2201] ));
 sg13g2_inv_2 \inv[2202]/_0_  (.Y(\inv_in[2203] ),
    .A(\inv_in[2202] ));
 sg13g2_inv_2 \inv[2203]/_0_  (.Y(\inv_in[2204] ),
    .A(\inv_in[2203] ));
 sg13g2_inv_2 \inv[2204]/_0_  (.Y(\inv_in[2205] ),
    .A(\inv_in[2204] ));
 sg13g2_inv_2 \inv[2205]/_0_  (.Y(\inv_in[2206] ),
    .A(\inv_in[2205] ));
 sg13g2_inv_2 \inv[2206]/_0_  (.Y(\inv_in[2207] ),
    .A(\inv_in[2206] ));
 sg13g2_inv_2 \inv[2207]/_0_  (.Y(\inv_in[2208] ),
    .A(\inv_in[2207] ));
 sg13g2_inv_2 \inv[2208]/_0_  (.Y(\inv_in[2209] ),
    .A(\inv_in[2208] ));
 sg13g2_inv_2 \inv[2209]/_0_  (.Y(\inv_in[2210] ),
    .A(\inv_in[2209] ));
 sg13g2_inv_2 \inv[220]/_0_  (.Y(\inv_in[221] ),
    .A(\inv_in[220] ));
 sg13g2_inv_2 \inv[2210]/_0_  (.Y(\inv_in[2211] ),
    .A(\inv_in[2210] ));
 sg13g2_inv_2 \inv[2211]/_0_  (.Y(\inv_in[2212] ),
    .A(\inv_in[2211] ));
 sg13g2_inv_2 \inv[2212]/_0_  (.Y(\inv_in[2213] ),
    .A(\inv_in[2212] ));
 sg13g2_inv_2 \inv[2213]/_0_  (.Y(\inv_in[2214] ),
    .A(\inv_in[2213] ));
 sg13g2_inv_2 \inv[2214]/_0_  (.Y(\inv_in[2215] ),
    .A(\inv_in[2214] ));
 sg13g2_inv_2 \inv[2215]/_0_  (.Y(\inv_in[2216] ),
    .A(\inv_in[2215] ));
 sg13g2_inv_2 \inv[2216]/_0_  (.Y(\inv_in[2217] ),
    .A(\inv_in[2216] ));
 sg13g2_inv_2 \inv[2217]/_0_  (.Y(\inv_in[2218] ),
    .A(\inv_in[2217] ));
 sg13g2_inv_2 \inv[2218]/_0_  (.Y(\inv_in[2219] ),
    .A(\inv_in[2218] ));
 sg13g2_inv_2 \inv[2219]/_0_  (.Y(\inv_in[2220] ),
    .A(\inv_in[2219] ));
 sg13g2_inv_2 \inv[221]/_0_  (.Y(\inv_in[222] ),
    .A(\inv_in[221] ));
 sg13g2_inv_2 \inv[2220]/_0_  (.Y(\inv_in[2221] ),
    .A(\inv_in[2220] ));
 sg13g2_inv_2 \inv[2221]/_0_  (.Y(\inv_in[2222] ),
    .A(\inv_in[2221] ));
 sg13g2_inv_2 \inv[2222]/_0_  (.Y(\inv_in[2223] ),
    .A(\inv_in[2222] ));
 sg13g2_inv_2 \inv[2223]/_0_  (.Y(\inv_in[2224] ),
    .A(\inv_in[2223] ));
 sg13g2_inv_2 \inv[2224]/_0_  (.Y(\inv_in[2225] ),
    .A(\inv_in[2224] ));
 sg13g2_inv_2 \inv[2225]/_0_  (.Y(\inv_in[2226] ),
    .A(\inv_in[2225] ));
 sg13g2_inv_2 \inv[2226]/_0_  (.Y(\inv_in[2227] ),
    .A(\inv_in[2226] ));
 sg13g2_inv_2 \inv[2227]/_0_  (.Y(\inv_in[2228] ),
    .A(\inv_in[2227] ));
 sg13g2_inv_2 \inv[2228]/_0_  (.Y(\inv_in[2229] ),
    .A(\inv_in[2228] ));
 sg13g2_inv_2 \inv[2229]/_0_  (.Y(\inv_in[2230] ),
    .A(\inv_in[2229] ));
 sg13g2_inv_2 \inv[222]/_0_  (.Y(\inv_in[223] ),
    .A(\inv_in[222] ));
 sg13g2_inv_2 \inv[2230]/_0_  (.Y(\inv_in[2231] ),
    .A(\inv_in[2230] ));
 sg13g2_inv_2 \inv[2231]/_0_  (.Y(\inv_in[2232] ),
    .A(\inv_in[2231] ));
 sg13g2_inv_2 \inv[2232]/_0_  (.Y(\inv_in[2233] ),
    .A(\inv_in[2232] ));
 sg13g2_inv_2 \inv[2233]/_0_  (.Y(\inv_in[2234] ),
    .A(\inv_in[2233] ));
 sg13g2_inv_2 \inv[2234]/_0_  (.Y(\inv_in[2235] ),
    .A(\inv_in[2234] ));
 sg13g2_inv_2 \inv[2235]/_0_  (.Y(\inv_in[2236] ),
    .A(\inv_in[2235] ));
 sg13g2_inv_2 \inv[2236]/_0_  (.Y(\inv_in[2237] ),
    .A(\inv_in[2236] ));
 sg13g2_inv_2 \inv[2237]/_0_  (.Y(\inv_in[2238] ),
    .A(\inv_in[2237] ));
 sg13g2_inv_2 \inv[2238]/_0_  (.Y(\inv_in[2239] ),
    .A(\inv_in[2238] ));
 sg13g2_inv_2 \inv[2239]/_0_  (.Y(\inv_in[2240] ),
    .A(\inv_in[2239] ));
 sg13g2_inv_2 \inv[223]/_0_  (.Y(\inv_in[224] ),
    .A(\inv_in[223] ));
 sg13g2_inv_2 \inv[2240]/_0_  (.Y(\inv_in[2241] ),
    .A(\inv_in[2240] ));
 sg13g2_inv_2 \inv[2241]/_0_  (.Y(\inv_in[2242] ),
    .A(\inv_in[2241] ));
 sg13g2_inv_2 \inv[2242]/_0_  (.Y(\inv_in[2243] ),
    .A(\inv_in[2242] ));
 sg13g2_inv_2 \inv[2243]/_0_  (.Y(\inv_in[2244] ),
    .A(\inv_in[2243] ));
 sg13g2_inv_2 \inv[2244]/_0_  (.Y(\inv_in[2245] ),
    .A(\inv_in[2244] ));
 sg13g2_inv_2 \inv[2245]/_0_  (.Y(\inv_in[2246] ),
    .A(\inv_in[2245] ));
 sg13g2_inv_2 \inv[2246]/_0_  (.Y(\inv_in[2247] ),
    .A(\inv_in[2246] ));
 sg13g2_inv_2 \inv[2247]/_0_  (.Y(\inv_in[2248] ),
    .A(\inv_in[2247] ));
 sg13g2_inv_2 \inv[2248]/_0_  (.Y(\inv_in[2249] ),
    .A(\inv_in[2248] ));
 sg13g2_inv_2 \inv[2249]/_0_  (.Y(\inv_in[2250] ),
    .A(\inv_in[2249] ));
 sg13g2_inv_2 \inv[224]/_0_  (.Y(\inv_in[225] ),
    .A(\inv_in[224] ));
 sg13g2_inv_2 \inv[2250]/_0_  (.Y(\inv_in[2251] ),
    .A(\inv_in[2250] ));
 sg13g2_inv_2 \inv[2251]/_0_  (.Y(\inv_in[2252] ),
    .A(\inv_in[2251] ));
 sg13g2_inv_2 \inv[2252]/_0_  (.Y(\inv_in[2253] ),
    .A(\inv_in[2252] ));
 sg13g2_inv_2 \inv[2253]/_0_  (.Y(\inv_in[2254] ),
    .A(\inv_in[2253] ));
 sg13g2_inv_2 \inv[2254]/_0_  (.Y(\inv_in[2255] ),
    .A(\inv_in[2254] ));
 sg13g2_inv_2 \inv[2255]/_0_  (.Y(\inv_in[2256] ),
    .A(\inv_in[2255] ));
 sg13g2_inv_2 \inv[2256]/_0_  (.Y(\inv_in[2257] ),
    .A(\inv_in[2256] ));
 sg13g2_inv_2 \inv[2257]/_0_  (.Y(\inv_in[2258] ),
    .A(\inv_in[2257] ));
 sg13g2_inv_2 \inv[2258]/_0_  (.Y(\inv_in[2259] ),
    .A(\inv_in[2258] ));
 sg13g2_inv_2 \inv[2259]/_0_  (.Y(\inv_in[2260] ),
    .A(\inv_in[2259] ));
 sg13g2_inv_2 \inv[225]/_0_  (.Y(\inv_in[226] ),
    .A(\inv_in[225] ));
 sg13g2_inv_2 \inv[2260]/_0_  (.Y(\inv_in[2261] ),
    .A(\inv_in[2260] ));
 sg13g2_inv_2 \inv[2261]/_0_  (.Y(\inv_in[2262] ),
    .A(\inv_in[2261] ));
 sg13g2_inv_2 \inv[2262]/_0_  (.Y(\inv_in[2263] ),
    .A(\inv_in[2262] ));
 sg13g2_inv_2 \inv[2263]/_0_  (.Y(\inv_in[2264] ),
    .A(\inv_in[2263] ));
 sg13g2_inv_2 \inv[2264]/_0_  (.Y(\inv_in[2265] ),
    .A(\inv_in[2264] ));
 sg13g2_inv_2 \inv[2265]/_0_  (.Y(\inv_in[2266] ),
    .A(\inv_in[2265] ));
 sg13g2_inv_2 \inv[2266]/_0_  (.Y(\inv_in[2267] ),
    .A(\inv_in[2266] ));
 sg13g2_inv_2 \inv[2267]/_0_  (.Y(\inv_in[2268] ),
    .A(\inv_in[2267] ));
 sg13g2_inv_2 \inv[2268]/_0_  (.Y(\inv_in[2269] ),
    .A(\inv_in[2268] ));
 sg13g2_inv_2 \inv[2269]/_0_  (.Y(\inv_in[2270] ),
    .A(\inv_in[2269] ));
 sg13g2_inv_2 \inv[226]/_0_  (.Y(\inv_in[227] ),
    .A(\inv_in[226] ));
 sg13g2_inv_2 \inv[2270]/_0_  (.Y(\inv_in[2271] ),
    .A(\inv_in[2270] ));
 sg13g2_inv_2 \inv[2271]/_0_  (.Y(\inv_in[2272] ),
    .A(\inv_in[2271] ));
 sg13g2_inv_2 \inv[2272]/_0_  (.Y(\inv_in[2273] ),
    .A(\inv_in[2272] ));
 sg13g2_inv_2 \inv[2273]/_0_  (.Y(\inv_in[2274] ),
    .A(\inv_in[2273] ));
 sg13g2_inv_2 \inv[2274]/_0_  (.Y(\inv_in[2275] ),
    .A(\inv_in[2274] ));
 sg13g2_inv_2 \inv[2275]/_0_  (.Y(\inv_in[2276] ),
    .A(\inv_in[2275] ));
 sg13g2_inv_2 \inv[2276]/_0_  (.Y(\inv_in[2277] ),
    .A(\inv_in[2276] ));
 sg13g2_inv_2 \inv[2277]/_0_  (.Y(\inv_in[2278] ),
    .A(\inv_in[2277] ));
 sg13g2_inv_2 \inv[2278]/_0_  (.Y(\inv_in[2279] ),
    .A(\inv_in[2278] ));
 sg13g2_inv_2 \inv[2279]/_0_  (.Y(\inv_in[2280] ),
    .A(\inv_in[2279] ));
 sg13g2_inv_2 \inv[227]/_0_  (.Y(\inv_in[228] ),
    .A(\inv_in[227] ));
 sg13g2_inv_2 \inv[2280]/_0_  (.Y(\inv_in[2281] ),
    .A(\inv_in[2280] ));
 sg13g2_inv_2 \inv[2281]/_0_  (.Y(\inv_in[2282] ),
    .A(\inv_in[2281] ));
 sg13g2_inv_2 \inv[2282]/_0_  (.Y(\inv_in[2283] ),
    .A(\inv_in[2282] ));
 sg13g2_inv_2 \inv[2283]/_0_  (.Y(\inv_in[2284] ),
    .A(\inv_in[2283] ));
 sg13g2_inv_2 \inv[2284]/_0_  (.Y(\inv_in[2285] ),
    .A(\inv_in[2284] ));
 sg13g2_inv_2 \inv[2285]/_0_  (.Y(\inv_in[2286] ),
    .A(\inv_in[2285] ));
 sg13g2_inv_2 \inv[2286]/_0_  (.Y(\inv_in[2287] ),
    .A(\inv_in[2286] ));
 sg13g2_inv_2 \inv[2287]/_0_  (.Y(\inv_in[2288] ),
    .A(\inv_in[2287] ));
 sg13g2_inv_2 \inv[2288]/_0_  (.Y(\inv_in[2289] ),
    .A(\inv_in[2288] ));
 sg13g2_inv_2 \inv[2289]/_0_  (.Y(\inv_in[2290] ),
    .A(\inv_in[2289] ));
 sg13g2_inv_2 \inv[228]/_0_  (.Y(\inv_in[229] ),
    .A(\inv_in[228] ));
 sg13g2_inv_2 \inv[2290]/_0_  (.Y(\inv_in[2291] ),
    .A(\inv_in[2290] ));
 sg13g2_inv_2 \inv[2291]/_0_  (.Y(\inv_in[2292] ),
    .A(\inv_in[2291] ));
 sg13g2_inv_2 \inv[2292]/_0_  (.Y(\inv_in[2293] ),
    .A(\inv_in[2292] ));
 sg13g2_inv_2 \inv[2293]/_0_  (.Y(\inv_in[2294] ),
    .A(\inv_in[2293] ));
 sg13g2_inv_2 \inv[2294]/_0_  (.Y(\inv_in[2295] ),
    .A(\inv_in[2294] ));
 sg13g2_inv_2 \inv[2295]/_0_  (.Y(\inv_in[2296] ),
    .A(\inv_in[2295] ));
 sg13g2_inv_2 \inv[2296]/_0_  (.Y(\inv_in[2297] ),
    .A(\inv_in[2296] ));
 sg13g2_inv_2 \inv[2297]/_0_  (.Y(\inv_in[2298] ),
    .A(\inv_in[2297] ));
 sg13g2_inv_2 \inv[2298]/_0_  (.Y(\inv_in[2299] ),
    .A(\inv_in[2298] ));
 sg13g2_inv_2 \inv[2299]/_0_  (.Y(\inv_in[2300] ),
    .A(\inv_in[2299] ));
 sg13g2_inv_2 \inv[229]/_0_  (.Y(\inv_in[230] ),
    .A(\inv_in[229] ));
 sg13g2_inv_2 \inv[22]/_0_  (.Y(\inv_in[23] ),
    .A(\inv_in[22] ));
 sg13g2_inv_2 \inv[2300]/_0_  (.Y(\inv_in[2301] ),
    .A(\inv_in[2300] ));
 sg13g2_inv_2 \inv[2301]/_0_  (.Y(\inv_in[2302] ),
    .A(\inv_in[2301] ));
 sg13g2_inv_2 \inv[2302]/_0_  (.Y(\inv_in[2303] ),
    .A(\inv_in[2302] ));
 sg13g2_inv_2 \inv[2303]/_0_  (.Y(\inv_in[2304] ),
    .A(\inv_in[2303] ));
 sg13g2_inv_2 \inv[2304]/_0_  (.Y(\inv_in[2305] ),
    .A(\inv_in[2304] ));
 sg13g2_inv_2 \inv[2305]/_0_  (.Y(\inv_in[2306] ),
    .A(\inv_in[2305] ));
 sg13g2_inv_2 \inv[2306]/_0_  (.Y(\inv_in[2307] ),
    .A(\inv_in[2306] ));
 sg13g2_inv_2 \inv[2307]/_0_  (.Y(\inv_in[2308] ),
    .A(\inv_in[2307] ));
 sg13g2_inv_2 \inv[2308]/_0_  (.Y(\inv_in[2309] ),
    .A(\inv_in[2308] ));
 sg13g2_inv_2 \inv[2309]/_0_  (.Y(\inv_in[2310] ),
    .A(\inv_in[2309] ));
 sg13g2_inv_2 \inv[230]/_0_  (.Y(\inv_in[231] ),
    .A(\inv_in[230] ));
 sg13g2_inv_2 \inv[2310]/_0_  (.Y(\inv_in[2311] ),
    .A(\inv_in[2310] ));
 sg13g2_inv_2 \inv[2311]/_0_  (.Y(\inv_in[2312] ),
    .A(\inv_in[2311] ));
 sg13g2_inv_2 \inv[2312]/_0_  (.Y(\inv_in[2313] ),
    .A(\inv_in[2312] ));
 sg13g2_inv_2 \inv[2313]/_0_  (.Y(\inv_in[2314] ),
    .A(\inv_in[2313] ));
 sg13g2_inv_2 \inv[2314]/_0_  (.Y(\inv_in[2315] ),
    .A(\inv_in[2314] ));
 sg13g2_inv_2 \inv[2315]/_0_  (.Y(\inv_in[2316] ),
    .A(\inv_in[2315] ));
 sg13g2_inv_2 \inv[2316]/_0_  (.Y(\inv_in[2317] ),
    .A(\inv_in[2316] ));
 sg13g2_inv_2 \inv[2317]/_0_  (.Y(\inv_in[2318] ),
    .A(\inv_in[2317] ));
 sg13g2_inv_2 \inv[2318]/_0_  (.Y(\inv_in[2319] ),
    .A(\inv_in[2318] ));
 sg13g2_inv_2 \inv[2319]/_0_  (.Y(\inv_in[2320] ),
    .A(\inv_in[2319] ));
 sg13g2_inv_2 \inv[231]/_0_  (.Y(\inv_in[232] ),
    .A(\inv_in[231] ));
 sg13g2_inv_2 \inv[2320]/_0_  (.Y(\inv_in[2321] ),
    .A(\inv_in[2320] ));
 sg13g2_inv_2 \inv[2321]/_0_  (.Y(\inv_in[2322] ),
    .A(\inv_in[2321] ));
 sg13g2_inv_2 \inv[2322]/_0_  (.Y(\inv_in[2323] ),
    .A(\inv_in[2322] ));
 sg13g2_inv_2 \inv[2323]/_0_  (.Y(\inv_in[2324] ),
    .A(\inv_in[2323] ));
 sg13g2_inv_2 \inv[2324]/_0_  (.Y(\inv_in[2325] ),
    .A(\inv_in[2324] ));
 sg13g2_inv_2 \inv[2325]/_0_  (.Y(\inv_in[2326] ),
    .A(\inv_in[2325] ));
 sg13g2_inv_2 \inv[2326]/_0_  (.Y(\inv_in[2327] ),
    .A(\inv_in[2326] ));
 sg13g2_inv_2 \inv[2327]/_0_  (.Y(\inv_in[2328] ),
    .A(\inv_in[2327] ));
 sg13g2_inv_2 \inv[2328]/_0_  (.Y(\inv_in[2329] ),
    .A(\inv_in[2328] ));
 sg13g2_inv_2 \inv[2329]/_0_  (.Y(\inv_in[2330] ),
    .A(\inv_in[2329] ));
 sg13g2_inv_2 \inv[232]/_0_  (.Y(\inv_in[233] ),
    .A(\inv_in[232] ));
 sg13g2_inv_2 \inv[2330]/_0_  (.Y(\inv_in[2331] ),
    .A(\inv_in[2330] ));
 sg13g2_inv_2 \inv[2331]/_0_  (.Y(\inv_in[2332] ),
    .A(\inv_in[2331] ));
 sg13g2_inv_2 \inv[2332]/_0_  (.Y(\inv_in[2333] ),
    .A(\inv_in[2332] ));
 sg13g2_inv_2 \inv[2333]/_0_  (.Y(\inv_in[2334] ),
    .A(\inv_in[2333] ));
 sg13g2_inv_2 \inv[2334]/_0_  (.Y(\inv_in[2335] ),
    .A(\inv_in[2334] ));
 sg13g2_inv_2 \inv[2335]/_0_  (.Y(\inv_in[2336] ),
    .A(\inv_in[2335] ));
 sg13g2_inv_2 \inv[2336]/_0_  (.Y(\inv_in[2337] ),
    .A(\inv_in[2336] ));
 sg13g2_inv_2 \inv[2337]/_0_  (.Y(\inv_in[2338] ),
    .A(\inv_in[2337] ));
 sg13g2_inv_2 \inv[2338]/_0_  (.Y(\inv_in[2339] ),
    .A(\inv_in[2338] ));
 sg13g2_inv_2 \inv[2339]/_0_  (.Y(\inv_in[2340] ),
    .A(\inv_in[2339] ));
 sg13g2_inv_2 \inv[233]/_0_  (.Y(\inv_in[234] ),
    .A(\inv_in[233] ));
 sg13g2_inv_2 \inv[2340]/_0_  (.Y(\inv_in[2341] ),
    .A(\inv_in[2340] ));
 sg13g2_inv_2 \inv[2341]/_0_  (.Y(\inv_in[2342] ),
    .A(\inv_in[2341] ));
 sg13g2_inv_2 \inv[2342]/_0_  (.Y(\inv_in[2343] ),
    .A(\inv_in[2342] ));
 sg13g2_inv_2 \inv[2343]/_0_  (.Y(\inv_in[2344] ),
    .A(\inv_in[2343] ));
 sg13g2_inv_2 \inv[2344]/_0_  (.Y(\inv_in[2345] ),
    .A(\inv_in[2344] ));
 sg13g2_inv_2 \inv[2345]/_0_  (.Y(\inv_in[2346] ),
    .A(\inv_in[2345] ));
 sg13g2_inv_2 \inv[2346]/_0_  (.Y(\inv_in[2347] ),
    .A(\inv_in[2346] ));
 sg13g2_inv_2 \inv[2347]/_0_  (.Y(\inv_in[2348] ),
    .A(\inv_in[2347] ));
 sg13g2_inv_2 \inv[2348]/_0_  (.Y(\inv_in[2349] ),
    .A(\inv_in[2348] ));
 sg13g2_inv_2 \inv[2349]/_0_  (.Y(\inv_in[2350] ),
    .A(\inv_in[2349] ));
 sg13g2_inv_2 \inv[234]/_0_  (.Y(\inv_in[235] ),
    .A(\inv_in[234] ));
 sg13g2_inv_2 \inv[2350]/_0_  (.Y(\inv_in[2351] ),
    .A(\inv_in[2350] ));
 sg13g2_inv_2 \inv[2351]/_0_  (.Y(\inv_in[2352] ),
    .A(\inv_in[2351] ));
 sg13g2_inv_2 \inv[2352]/_0_  (.Y(\inv_in[2353] ),
    .A(\inv_in[2352] ));
 sg13g2_inv_2 \inv[2353]/_0_  (.Y(\inv_in[2354] ),
    .A(\inv_in[2353] ));
 sg13g2_inv_2 \inv[2354]/_0_  (.Y(\inv_in[2355] ),
    .A(\inv_in[2354] ));
 sg13g2_inv_2 \inv[2355]/_0_  (.Y(\inv_in[2356] ),
    .A(\inv_in[2355] ));
 sg13g2_inv_2 \inv[2356]/_0_  (.Y(\inv_in[2357] ),
    .A(\inv_in[2356] ));
 sg13g2_inv_2 \inv[2357]/_0_  (.Y(\inv_in[2358] ),
    .A(\inv_in[2357] ));
 sg13g2_inv_2 \inv[2358]/_0_  (.Y(\inv_in[2359] ),
    .A(\inv_in[2358] ));
 sg13g2_inv_2 \inv[2359]/_0_  (.Y(\inv_in[2360] ),
    .A(\inv_in[2359] ));
 sg13g2_inv_2 \inv[235]/_0_  (.Y(\inv_in[236] ),
    .A(\inv_in[235] ));
 sg13g2_inv_2 \inv[2360]/_0_  (.Y(\inv_in[2361] ),
    .A(\inv_in[2360] ));
 sg13g2_inv_2 \inv[2361]/_0_  (.Y(\inv_in[2362] ),
    .A(\inv_in[2361] ));
 sg13g2_inv_2 \inv[2362]/_0_  (.Y(\inv_in[2363] ),
    .A(\inv_in[2362] ));
 sg13g2_inv_2 \inv[2363]/_0_  (.Y(\inv_in[2364] ),
    .A(\inv_in[2363] ));
 sg13g2_inv_2 \inv[2364]/_0_  (.Y(\inv_in[2365] ),
    .A(\inv_in[2364] ));
 sg13g2_inv_2 \inv[2365]/_0_  (.Y(\inv_in[2366] ),
    .A(\inv_in[2365] ));
 sg13g2_inv_2 \inv[2366]/_0_  (.Y(\inv_in[2367] ),
    .A(\inv_in[2366] ));
 sg13g2_inv_2 \inv[2367]/_0_  (.Y(\inv_in[2368] ),
    .A(\inv_in[2367] ));
 sg13g2_inv_2 \inv[2368]/_0_  (.Y(\inv_in[2369] ),
    .A(\inv_in[2368] ));
 sg13g2_inv_2 \inv[2369]/_0_  (.Y(\inv_in[2370] ),
    .A(\inv_in[2369] ));
 sg13g2_inv_2 \inv[236]/_0_  (.Y(\inv_in[237] ),
    .A(\inv_in[236] ));
 sg13g2_inv_2 \inv[2370]/_0_  (.Y(\inv_in[2371] ),
    .A(\inv_in[2370] ));
 sg13g2_inv_2 \inv[2371]/_0_  (.Y(\inv_in[2372] ),
    .A(\inv_in[2371] ));
 sg13g2_inv_2 \inv[2372]/_0_  (.Y(\inv_in[2373] ),
    .A(\inv_in[2372] ));
 sg13g2_inv_2 \inv[2373]/_0_  (.Y(\inv_in[2374] ),
    .A(\inv_in[2373] ));
 sg13g2_inv_2 \inv[2374]/_0_  (.Y(\inv_in[2375] ),
    .A(\inv_in[2374] ));
 sg13g2_inv_2 \inv[2375]/_0_  (.Y(\inv_in[2376] ),
    .A(\inv_in[2375] ));
 sg13g2_inv_2 \inv[2376]/_0_  (.Y(\inv_in[2377] ),
    .A(\inv_in[2376] ));
 sg13g2_inv_2 \inv[2377]/_0_  (.Y(\inv_in[2378] ),
    .A(\inv_in[2377] ));
 sg13g2_inv_2 \inv[2378]/_0_  (.Y(\inv_in[2379] ),
    .A(\inv_in[2378] ));
 sg13g2_inv_2 \inv[2379]/_0_  (.Y(\inv_in[2380] ),
    .A(\inv_in[2379] ));
 sg13g2_inv_2 \inv[237]/_0_  (.Y(\inv_in[238] ),
    .A(\inv_in[237] ));
 sg13g2_inv_2 \inv[2380]/_0_  (.Y(\inv_in[2381] ),
    .A(\inv_in[2380] ));
 sg13g2_inv_2 \inv[2381]/_0_  (.Y(\inv_in[2382] ),
    .A(\inv_in[2381] ));
 sg13g2_inv_2 \inv[2382]/_0_  (.Y(\inv_in[2383] ),
    .A(\inv_in[2382] ));
 sg13g2_inv_2 \inv[2383]/_0_  (.Y(\inv_in[2384] ),
    .A(\inv_in[2383] ));
 sg13g2_inv_2 \inv[2384]/_0_  (.Y(\inv_in[2385] ),
    .A(\inv_in[2384] ));
 sg13g2_inv_2 \inv[2385]/_0_  (.Y(\inv_in[2386] ),
    .A(\inv_in[2385] ));
 sg13g2_inv_2 \inv[2386]/_0_  (.Y(\inv_in[2387] ),
    .A(\inv_in[2386] ));
 sg13g2_inv_2 \inv[2387]/_0_  (.Y(\inv_in[2388] ),
    .A(\inv_in[2387] ));
 sg13g2_inv_2 \inv[2388]/_0_  (.Y(\inv_in[2389] ),
    .A(\inv_in[2388] ));
 sg13g2_inv_2 \inv[2389]/_0_  (.Y(\inv_in[2390] ),
    .A(\inv_in[2389] ));
 sg13g2_inv_2 \inv[238]/_0_  (.Y(\inv_in[239] ),
    .A(\inv_in[238] ));
 sg13g2_inv_2 \inv[2390]/_0_  (.Y(\inv_in[2391] ),
    .A(\inv_in[2390] ));
 sg13g2_inv_2 \inv[2391]/_0_  (.Y(\inv_in[2392] ),
    .A(\inv_in[2391] ));
 sg13g2_inv_2 \inv[2392]/_0_  (.Y(\inv_in[2393] ),
    .A(\inv_in[2392] ));
 sg13g2_inv_2 \inv[2393]/_0_  (.Y(\inv_in[2394] ),
    .A(\inv_in[2393] ));
 sg13g2_inv_2 \inv[2394]/_0_  (.Y(\inv_in[2395] ),
    .A(\inv_in[2394] ));
 sg13g2_inv_2 \inv[2395]/_0_  (.Y(\inv_in[2396] ),
    .A(\inv_in[2395] ));
 sg13g2_inv_2 \inv[2396]/_0_  (.Y(\inv_in[2397] ),
    .A(\inv_in[2396] ));
 sg13g2_inv_2 \inv[2397]/_0_  (.Y(\inv_in[2398] ),
    .A(\inv_in[2397] ));
 sg13g2_inv_2 \inv[2398]/_0_  (.Y(\inv_in[2399] ),
    .A(\inv_in[2398] ));
 sg13g2_inv_2 \inv[2399]/_0_  (.Y(\inv_in[2400] ),
    .A(\inv_in[2399] ));
 sg13g2_inv_2 \inv[239]/_0_  (.Y(\inv_in[240] ),
    .A(\inv_in[239] ));
 sg13g2_inv_2 \inv[23]/_0_  (.Y(\inv_in[24] ),
    .A(\inv_in[23] ));
 sg13g2_inv_2 \inv[2400]/_0_  (.Y(\inv_in[2401] ),
    .A(\inv_in[2400] ));
 sg13g2_inv_2 \inv[2401]/_0_  (.Y(\inv_in[2402] ),
    .A(\inv_in[2401] ));
 sg13g2_inv_2 \inv[2402]/_0_  (.Y(\inv_in[2403] ),
    .A(\inv_in[2402] ));
 sg13g2_inv_2 \inv[2403]/_0_  (.Y(\inv_in[2404] ),
    .A(\inv_in[2403] ));
 sg13g2_inv_2 \inv[2404]/_0_  (.Y(\inv_in[2405] ),
    .A(\inv_in[2404] ));
 sg13g2_inv_2 \inv[2405]/_0_  (.Y(\inv_in[2406] ),
    .A(\inv_in[2405] ));
 sg13g2_inv_2 \inv[2406]/_0_  (.Y(\inv_in[2407] ),
    .A(\inv_in[2406] ));
 sg13g2_inv_2 \inv[2407]/_0_  (.Y(\inv_in[2408] ),
    .A(\inv_in[2407] ));
 sg13g2_inv_2 \inv[2408]/_0_  (.Y(\inv_in[2409] ),
    .A(\inv_in[2408] ));
 sg13g2_inv_2 \inv[2409]/_0_  (.Y(\inv_in[2410] ),
    .A(\inv_in[2409] ));
 sg13g2_inv_2 \inv[240]/_0_  (.Y(\inv_in[241] ),
    .A(\inv_in[240] ));
 sg13g2_inv_2 \inv[2410]/_0_  (.Y(\inv_in[2411] ),
    .A(\inv_in[2410] ));
 sg13g2_inv_2 \inv[2411]/_0_  (.Y(\inv_in[2412] ),
    .A(\inv_in[2411] ));
 sg13g2_inv_2 \inv[2412]/_0_  (.Y(\inv_in[2413] ),
    .A(\inv_in[2412] ));
 sg13g2_inv_2 \inv[2413]/_0_  (.Y(\inv_in[2414] ),
    .A(\inv_in[2413] ));
 sg13g2_inv_2 \inv[2414]/_0_  (.Y(\inv_in[2415] ),
    .A(\inv_in[2414] ));
 sg13g2_inv_2 \inv[2415]/_0_  (.Y(\inv_in[2416] ),
    .A(\inv_in[2415] ));
 sg13g2_inv_2 \inv[2416]/_0_  (.Y(\inv_in[2417] ),
    .A(\inv_in[2416] ));
 sg13g2_inv_2 \inv[2417]/_0_  (.Y(\inv_in[2418] ),
    .A(\inv_in[2417] ));
 sg13g2_inv_2 \inv[2418]/_0_  (.Y(\inv_in[2419] ),
    .A(\inv_in[2418] ));
 sg13g2_inv_2 \inv[2419]/_0_  (.Y(\inv_in[2420] ),
    .A(\inv_in[2419] ));
 sg13g2_inv_2 \inv[241]/_0_  (.Y(\inv_in[242] ),
    .A(\inv_in[241] ));
 sg13g2_inv_2 \inv[2420]/_0_  (.Y(\inv_in[2421] ),
    .A(\inv_in[2420] ));
 sg13g2_inv_2 \inv[2421]/_0_  (.Y(\inv_in[2422] ),
    .A(\inv_in[2421] ));
 sg13g2_inv_2 \inv[2422]/_0_  (.Y(\inv_in[2423] ),
    .A(\inv_in[2422] ));
 sg13g2_inv_2 \inv[2423]/_0_  (.Y(\inv_in[2424] ),
    .A(\inv_in[2423] ));
 sg13g2_inv_2 \inv[2424]/_0_  (.Y(\inv_in[2425] ),
    .A(\inv_in[2424] ));
 sg13g2_inv_2 \inv[2425]/_0_  (.Y(\inv_in[2426] ),
    .A(\inv_in[2425] ));
 sg13g2_inv_2 \inv[2426]/_0_  (.Y(\inv_in[2427] ),
    .A(\inv_in[2426] ));
 sg13g2_inv_2 \inv[2427]/_0_  (.Y(\inv_in[2428] ),
    .A(\inv_in[2427] ));
 sg13g2_inv_2 \inv[2428]/_0_  (.Y(\inv_in[2429] ),
    .A(\inv_in[2428] ));
 sg13g2_inv_2 \inv[2429]/_0_  (.Y(\inv_in[2430] ),
    .A(\inv_in[2429] ));
 sg13g2_inv_2 \inv[242]/_0_  (.Y(\inv_in[243] ),
    .A(\inv_in[242] ));
 sg13g2_inv_2 \inv[2430]/_0_  (.Y(\inv_in[2431] ),
    .A(\inv_in[2430] ));
 sg13g2_inv_2 \inv[2431]/_0_  (.Y(\inv_in[2432] ),
    .A(\inv_in[2431] ));
 sg13g2_inv_2 \inv[2432]/_0_  (.Y(\inv_in[2433] ),
    .A(\inv_in[2432] ));
 sg13g2_inv_2 \inv[2433]/_0_  (.Y(\inv_in[2434] ),
    .A(\inv_in[2433] ));
 sg13g2_inv_2 \inv[2434]/_0_  (.Y(\inv_in[2435] ),
    .A(\inv_in[2434] ));
 sg13g2_inv_2 \inv[2435]/_0_  (.Y(\inv_in[2436] ),
    .A(\inv_in[2435] ));
 sg13g2_inv_2 \inv[2436]/_0_  (.Y(\inv_in[2437] ),
    .A(\inv_in[2436] ));
 sg13g2_inv_2 \inv[2437]/_0_  (.Y(\inv_in[2438] ),
    .A(\inv_in[2437] ));
 sg13g2_inv_2 \inv[2438]/_0_  (.Y(\inv_in[2439] ),
    .A(\inv_in[2438] ));
 sg13g2_inv_2 \inv[2439]/_0_  (.Y(\inv_in[2440] ),
    .A(\inv_in[2439] ));
 sg13g2_inv_2 \inv[243]/_0_  (.Y(\inv_in[244] ),
    .A(\inv_in[243] ));
 sg13g2_inv_2 \inv[2440]/_0_  (.Y(\inv_in[2441] ),
    .A(\inv_in[2440] ));
 sg13g2_inv_2 \inv[2441]/_0_  (.Y(\inv_in[2442] ),
    .A(\inv_in[2441] ));
 sg13g2_inv_2 \inv[2442]/_0_  (.Y(\inv_in[2443] ),
    .A(\inv_in[2442] ));
 sg13g2_inv_2 \inv[2443]/_0_  (.Y(\inv_in[2444] ),
    .A(\inv_in[2443] ));
 sg13g2_inv_2 \inv[2444]/_0_  (.Y(\inv_in[2445] ),
    .A(\inv_in[2444] ));
 sg13g2_inv_2 \inv[2445]/_0_  (.Y(\inv_in[2446] ),
    .A(\inv_in[2445] ));
 sg13g2_inv_2 \inv[2446]/_0_  (.Y(\inv_in[2447] ),
    .A(\inv_in[2446] ));
 sg13g2_inv_2 \inv[2447]/_0_  (.Y(\inv_in[2448] ),
    .A(\inv_in[2447] ));
 sg13g2_inv_2 \inv[2448]/_0_  (.Y(\inv_in[2449] ),
    .A(\inv_in[2448] ));
 sg13g2_inv_2 \inv[2449]/_0_  (.Y(\inv_in[2450] ),
    .A(\inv_in[2449] ));
 sg13g2_inv_2 \inv[244]/_0_  (.Y(\inv_in[245] ),
    .A(\inv_in[244] ));
 sg13g2_inv_2 \inv[2450]/_0_  (.Y(\inv_in[2451] ),
    .A(\inv_in[2450] ));
 sg13g2_inv_2 \inv[2451]/_0_  (.Y(\inv_in[2452] ),
    .A(\inv_in[2451] ));
 sg13g2_inv_2 \inv[2452]/_0_  (.Y(\inv_in[2453] ),
    .A(\inv_in[2452] ));
 sg13g2_inv_2 \inv[2453]/_0_  (.Y(\inv_in[2454] ),
    .A(\inv_in[2453] ));
 sg13g2_inv_2 \inv[2454]/_0_  (.Y(\inv_in[2455] ),
    .A(\inv_in[2454] ));
 sg13g2_inv_2 \inv[2455]/_0_  (.Y(\inv_in[2456] ),
    .A(\inv_in[2455] ));
 sg13g2_inv_2 \inv[2456]/_0_  (.Y(\inv_in[2457] ),
    .A(\inv_in[2456] ));
 sg13g2_inv_2 \inv[2457]/_0_  (.Y(\inv_in[2458] ),
    .A(\inv_in[2457] ));
 sg13g2_inv_2 \inv[2458]/_0_  (.Y(\inv_in[2459] ),
    .A(\inv_in[2458] ));
 sg13g2_inv_2 \inv[2459]/_0_  (.Y(\inv_in[2460] ),
    .A(\inv_in[2459] ));
 sg13g2_inv_2 \inv[245]/_0_  (.Y(\inv_in[246] ),
    .A(\inv_in[245] ));
 sg13g2_inv_2 \inv[2460]/_0_  (.Y(\inv_in[2461] ),
    .A(\inv_in[2460] ));
 sg13g2_inv_2 \inv[2461]/_0_  (.Y(\inv_in[2462] ),
    .A(\inv_in[2461] ));
 sg13g2_inv_2 \inv[2462]/_0_  (.Y(\inv_in[2463] ),
    .A(\inv_in[2462] ));
 sg13g2_inv_2 \inv[2463]/_0_  (.Y(\inv_in[2464] ),
    .A(\inv_in[2463] ));
 sg13g2_inv_2 \inv[2464]/_0_  (.Y(\inv_in[2465] ),
    .A(\inv_in[2464] ));
 sg13g2_inv_2 \inv[2465]/_0_  (.Y(\inv_in[2466] ),
    .A(\inv_in[2465] ));
 sg13g2_inv_2 \inv[2466]/_0_  (.Y(\inv_in[2467] ),
    .A(\inv_in[2466] ));
 sg13g2_inv_2 \inv[2467]/_0_  (.Y(\inv_in[2468] ),
    .A(\inv_in[2467] ));
 sg13g2_inv_2 \inv[2468]/_0_  (.Y(\inv_in[2469] ),
    .A(\inv_in[2468] ));
 sg13g2_inv_2 \inv[2469]/_0_  (.Y(\inv_in[2470] ),
    .A(\inv_in[2469] ));
 sg13g2_inv_2 \inv[246]/_0_  (.Y(\inv_in[247] ),
    .A(\inv_in[246] ));
 sg13g2_inv_2 \inv[2470]/_0_  (.Y(\inv_in[2471] ),
    .A(\inv_in[2470] ));
 sg13g2_inv_2 \inv[2471]/_0_  (.Y(\inv_in[2472] ),
    .A(\inv_in[2471] ));
 sg13g2_inv_2 \inv[2472]/_0_  (.Y(\inv_in[2473] ),
    .A(\inv_in[2472] ));
 sg13g2_inv_2 \inv[2473]/_0_  (.Y(\inv_in[2474] ),
    .A(\inv_in[2473] ));
 sg13g2_inv_2 \inv[2474]/_0_  (.Y(\inv_in[2475] ),
    .A(\inv_in[2474] ));
 sg13g2_inv_2 \inv[2475]/_0_  (.Y(\inv_in[2476] ),
    .A(\inv_in[2475] ));
 sg13g2_inv_2 \inv[2476]/_0_  (.Y(\inv_in[2477] ),
    .A(\inv_in[2476] ));
 sg13g2_inv_2 \inv[2477]/_0_  (.Y(\inv_in[2478] ),
    .A(\inv_in[2477] ));
 sg13g2_inv_2 \inv[2478]/_0_  (.Y(\inv_in[2479] ),
    .A(\inv_in[2478] ));
 sg13g2_inv_2 \inv[2479]/_0_  (.Y(\inv_in[2480] ),
    .A(\inv_in[2479] ));
 sg13g2_inv_2 \inv[247]/_0_  (.Y(\inv_in[248] ),
    .A(\inv_in[247] ));
 sg13g2_inv_2 \inv[2480]/_0_  (.Y(\inv_in[2481] ),
    .A(\inv_in[2480] ));
 sg13g2_inv_2 \inv[2481]/_0_  (.Y(\inv_in[2482] ),
    .A(\inv_in[2481] ));
 sg13g2_inv_2 \inv[2482]/_0_  (.Y(\inv_in[2483] ),
    .A(\inv_in[2482] ));
 sg13g2_inv_2 \inv[2483]/_0_  (.Y(\inv_in[2484] ),
    .A(\inv_in[2483] ));
 sg13g2_inv_2 \inv[2484]/_0_  (.Y(\inv_in[2485] ),
    .A(\inv_in[2484] ));
 sg13g2_inv_2 \inv[2485]/_0_  (.Y(\inv_in[2486] ),
    .A(\inv_in[2485] ));
 sg13g2_inv_2 \inv[2486]/_0_  (.Y(\inv_in[2487] ),
    .A(\inv_in[2486] ));
 sg13g2_inv_2 \inv[2487]/_0_  (.Y(\inv_in[2488] ),
    .A(\inv_in[2487] ));
 sg13g2_inv_2 \inv[2488]/_0_  (.Y(\inv_in[2489] ),
    .A(\inv_in[2488] ));
 sg13g2_inv_2 \inv[2489]/_0_  (.Y(\inv_in[2490] ),
    .A(\inv_in[2489] ));
 sg13g2_inv_2 \inv[248]/_0_  (.Y(\inv_in[249] ),
    .A(\inv_in[248] ));
 sg13g2_inv_2 \inv[2490]/_0_  (.Y(\inv_in[2491] ),
    .A(\inv_in[2490] ));
 sg13g2_inv_2 \inv[2491]/_0_  (.Y(\inv_in[2492] ),
    .A(\inv_in[2491] ));
 sg13g2_inv_2 \inv[2492]/_0_  (.Y(\inv_in[2493] ),
    .A(\inv_in[2492] ));
 sg13g2_inv_2 \inv[2493]/_0_  (.Y(\inv_in[2494] ),
    .A(\inv_in[2493] ));
 sg13g2_inv_2 \inv[2494]/_0_  (.Y(\inv_in[2495] ),
    .A(\inv_in[2494] ));
 sg13g2_inv_2 \inv[2495]/_0_  (.Y(\inv_in[2496] ),
    .A(\inv_in[2495] ));
 sg13g2_inv_2 \inv[2496]/_0_  (.Y(\inv_in[2497] ),
    .A(\inv_in[2496] ));
 sg13g2_inv_2 \inv[2497]/_0_  (.Y(\inv_in[2498] ),
    .A(\inv_in[2497] ));
 sg13g2_inv_2 \inv[2498]/_0_  (.Y(\inv_in[2499] ),
    .A(\inv_in[2498] ));
 sg13g2_inv_2 \inv[2499]/_0_  (.Y(\inv_in[2500] ),
    .A(\inv_in[2499] ));
 sg13g2_inv_2 \inv[249]/_0_  (.Y(\inv_in[250] ),
    .A(\inv_in[249] ));
 sg13g2_inv_2 \inv[24]/_0_  (.Y(\inv_in[25] ),
    .A(\inv_in[24] ));
 sg13g2_inv_2 \inv[2500]/_0_  (.Y(\inv_in[2501] ),
    .A(\inv_in[2500] ));
 sg13g2_inv_2 \inv[2501]/_0_  (.Y(\inv_in[2502] ),
    .A(\inv_in[2501] ));
 sg13g2_inv_2 \inv[2502]/_0_  (.Y(\inv_in[2503] ),
    .A(\inv_in[2502] ));
 sg13g2_inv_2 \inv[2503]/_0_  (.Y(\inv_in[2504] ),
    .A(\inv_in[2503] ));
 sg13g2_inv_2 \inv[2504]/_0_  (.Y(\inv_in[2505] ),
    .A(\inv_in[2504] ));
 sg13g2_inv_2 \inv[2505]/_0_  (.Y(\inv_in[2506] ),
    .A(\inv_in[2505] ));
 sg13g2_inv_2 \inv[2506]/_0_  (.Y(\inv_in[2507] ),
    .A(\inv_in[2506] ));
 sg13g2_inv_2 \inv[2507]/_0_  (.Y(\inv_in[2508] ),
    .A(\inv_in[2507] ));
 sg13g2_inv_2 \inv[2508]/_0_  (.Y(\inv_in[2509] ),
    .A(\inv_in[2508] ));
 sg13g2_inv_2 \inv[2509]/_0_  (.Y(\inv_in[2510] ),
    .A(\inv_in[2509] ));
 sg13g2_inv_2 \inv[250]/_0_  (.Y(\inv_in[251] ),
    .A(\inv_in[250] ));
 sg13g2_inv_2 \inv[2510]/_0_  (.Y(\inv_in[2511] ),
    .A(\inv_in[2510] ));
 sg13g2_inv_2 \inv[2511]/_0_  (.Y(\inv_in[2512] ),
    .A(\inv_in[2511] ));
 sg13g2_inv_2 \inv[2512]/_0_  (.Y(\inv_in[2513] ),
    .A(\inv_in[2512] ));
 sg13g2_inv_2 \inv[2513]/_0_  (.Y(\inv_in[2514] ),
    .A(\inv_in[2513] ));
 sg13g2_inv_2 \inv[2514]/_0_  (.Y(\inv_in[2515] ),
    .A(\inv_in[2514] ));
 sg13g2_inv_2 \inv[2515]/_0_  (.Y(\inv_in[2516] ),
    .A(\inv_in[2515] ));
 sg13g2_inv_2 \inv[2516]/_0_  (.Y(\inv_in[2517] ),
    .A(\inv_in[2516] ));
 sg13g2_inv_2 \inv[2517]/_0_  (.Y(\inv_in[2518] ),
    .A(\inv_in[2517] ));
 sg13g2_inv_2 \inv[2518]/_0_  (.Y(\inv_in[2519] ),
    .A(\inv_in[2518] ));
 sg13g2_inv_2 \inv[2519]/_0_  (.Y(\inv_in[2520] ),
    .A(\inv_in[2519] ));
 sg13g2_inv_2 \inv[251]/_0_  (.Y(\inv_in[252] ),
    .A(\inv_in[251] ));
 sg13g2_inv_2 \inv[2520]/_0_  (.Y(\inv_in[2521] ),
    .A(\inv_in[2520] ));
 sg13g2_inv_2 \inv[2521]/_0_  (.Y(\inv_in[2522] ),
    .A(\inv_in[2521] ));
 sg13g2_inv_2 \inv[2522]/_0_  (.Y(\inv_in[2523] ),
    .A(\inv_in[2522] ));
 sg13g2_inv_2 \inv[2523]/_0_  (.Y(\inv_in[2524] ),
    .A(\inv_in[2523] ));
 sg13g2_inv_2 \inv[2524]/_0_  (.Y(\inv_in[2525] ),
    .A(\inv_in[2524] ));
 sg13g2_inv_2 \inv[2525]/_0_  (.Y(\inv_in[2526] ),
    .A(\inv_in[2525] ));
 sg13g2_inv_2 \inv[2526]/_0_  (.Y(\inv_in[2527] ),
    .A(\inv_in[2526] ));
 sg13g2_inv_2 \inv[2527]/_0_  (.Y(\inv_in[2528] ),
    .A(\inv_in[2527] ));
 sg13g2_inv_2 \inv[2528]/_0_  (.Y(\inv_in[2529] ),
    .A(\inv_in[2528] ));
 sg13g2_inv_2 \inv[2529]/_0_  (.Y(\inv_in[2530] ),
    .A(\inv_in[2529] ));
 sg13g2_inv_2 \inv[252]/_0_  (.Y(\inv_in[253] ),
    .A(\inv_in[252] ));
 sg13g2_inv_2 \inv[2530]/_0_  (.Y(\inv_in[2531] ),
    .A(\inv_in[2530] ));
 sg13g2_inv_2 \inv[2531]/_0_  (.Y(\inv_in[2532] ),
    .A(\inv_in[2531] ));
 sg13g2_inv_2 \inv[2532]/_0_  (.Y(\inv_in[2533] ),
    .A(\inv_in[2532] ));
 sg13g2_inv_2 \inv[2533]/_0_  (.Y(\inv_in[2534] ),
    .A(\inv_in[2533] ));
 sg13g2_inv_2 \inv[2534]/_0_  (.Y(\inv_in[2535] ),
    .A(\inv_in[2534] ));
 sg13g2_inv_2 \inv[2535]/_0_  (.Y(\inv_in[2536] ),
    .A(\inv_in[2535] ));
 sg13g2_inv_2 \inv[2536]/_0_  (.Y(\inv_in[2537] ),
    .A(\inv_in[2536] ));
 sg13g2_inv_2 \inv[2537]/_0_  (.Y(\inv_in[2538] ),
    .A(\inv_in[2537] ));
 sg13g2_inv_2 \inv[2538]/_0_  (.Y(\inv_in[2539] ),
    .A(\inv_in[2538] ));
 sg13g2_inv_2 \inv[2539]/_0_  (.Y(\inv_in[2540] ),
    .A(\inv_in[2539] ));
 sg13g2_inv_2 \inv[253]/_0_  (.Y(\inv_in[254] ),
    .A(\inv_in[253] ));
 sg13g2_inv_2 \inv[2540]/_0_  (.Y(\inv_in[2541] ),
    .A(\inv_in[2540] ));
 sg13g2_inv_2 \inv[2541]/_0_  (.Y(\inv_in[2542] ),
    .A(\inv_in[2541] ));
 sg13g2_inv_2 \inv[2542]/_0_  (.Y(\inv_in[2543] ),
    .A(\inv_in[2542] ));
 sg13g2_inv_2 \inv[2543]/_0_  (.Y(\inv_in[2544] ),
    .A(\inv_in[2543] ));
 sg13g2_inv_2 \inv[2544]/_0_  (.Y(\inv_in[2545] ),
    .A(\inv_in[2544] ));
 sg13g2_inv_2 \inv[2545]/_0_  (.Y(\inv_in[2546] ),
    .A(\inv_in[2545] ));
 sg13g2_inv_2 \inv[2546]/_0_  (.Y(\inv_in[2547] ),
    .A(\inv_in[2546] ));
 sg13g2_inv_2 \inv[2547]/_0_  (.Y(\inv_in[2548] ),
    .A(\inv_in[2547] ));
 sg13g2_inv_2 \inv[2548]/_0_  (.Y(\inv_in[2549] ),
    .A(\inv_in[2548] ));
 sg13g2_inv_2 \inv[2549]/_0_  (.Y(\inv_in[2550] ),
    .A(\inv_in[2549] ));
 sg13g2_inv_2 \inv[254]/_0_  (.Y(\inv_in[255] ),
    .A(\inv_in[254] ));
 sg13g2_inv_2 \inv[2550]/_0_  (.Y(\inv_in[2551] ),
    .A(\inv_in[2550] ));
 sg13g2_inv_2 \inv[2551]/_0_  (.Y(\inv_in[2552] ),
    .A(\inv_in[2551] ));
 sg13g2_inv_2 \inv[2552]/_0_  (.Y(\inv_in[2553] ),
    .A(\inv_in[2552] ));
 sg13g2_inv_2 \inv[2553]/_0_  (.Y(\inv_in[2554] ),
    .A(\inv_in[2553] ));
 sg13g2_inv_2 \inv[2554]/_0_  (.Y(\inv_in[2555] ),
    .A(\inv_in[2554] ));
 sg13g2_inv_2 \inv[2555]/_0_  (.Y(\inv_in[2556] ),
    .A(\inv_in[2555] ));
 sg13g2_inv_2 \inv[2556]/_0_  (.Y(\inv_in[2557] ),
    .A(\inv_in[2556] ));
 sg13g2_inv_2 \inv[2557]/_0_  (.Y(\inv_in[2558] ),
    .A(\inv_in[2557] ));
 sg13g2_inv_2 \inv[2558]/_0_  (.Y(\inv_in[2559] ),
    .A(\inv_in[2558] ));
 sg13g2_inv_2 \inv[2559]/_0_  (.Y(\inv_in[2560] ),
    .A(\inv_in[2559] ));
 sg13g2_inv_2 \inv[255]/_0_  (.Y(\inv_in[256] ),
    .A(\inv_in[255] ));
 sg13g2_inv_2 \inv[2560]/_0_  (.Y(\inv_in[2561] ),
    .A(\inv_in[2560] ));
 sg13g2_inv_2 \inv[2561]/_0_  (.Y(\inv_in[2562] ),
    .A(\inv_in[2561] ));
 sg13g2_inv_2 \inv[2562]/_0_  (.Y(\inv_in[2563] ),
    .A(\inv_in[2562] ));
 sg13g2_inv_2 \inv[2563]/_0_  (.Y(\inv_in[2564] ),
    .A(\inv_in[2563] ));
 sg13g2_inv_2 \inv[2564]/_0_  (.Y(\inv_in[2565] ),
    .A(\inv_in[2564] ));
 sg13g2_inv_2 \inv[2565]/_0_  (.Y(\inv_in[2566] ),
    .A(\inv_in[2565] ));
 sg13g2_inv_2 \inv[2566]/_0_  (.Y(\inv_in[2567] ),
    .A(\inv_in[2566] ));
 sg13g2_inv_2 \inv[2567]/_0_  (.Y(\inv_in[2568] ),
    .A(\inv_in[2567] ));
 sg13g2_inv_2 \inv[2568]/_0_  (.Y(\inv_in[2569] ),
    .A(\inv_in[2568] ));
 sg13g2_inv_2 \inv[2569]/_0_  (.Y(\inv_in[2570] ),
    .A(\inv_in[2569] ));
 sg13g2_inv_2 \inv[256]/_0_  (.Y(\inv_in[257] ),
    .A(\inv_in[256] ));
 sg13g2_inv_2 \inv[2570]/_0_  (.Y(\inv_in[2571] ),
    .A(\inv_in[2570] ));
 sg13g2_inv_2 \inv[2571]/_0_  (.Y(\inv_in[2572] ),
    .A(\inv_in[2571] ));
 sg13g2_inv_2 \inv[2572]/_0_  (.Y(\inv_in[2573] ),
    .A(\inv_in[2572] ));
 sg13g2_inv_2 \inv[2573]/_0_  (.Y(\inv_in[2574] ),
    .A(\inv_in[2573] ));
 sg13g2_inv_2 \inv[2574]/_0_  (.Y(\inv_in[2575] ),
    .A(\inv_in[2574] ));
 sg13g2_inv_2 \inv[2575]/_0_  (.Y(\inv_in[2576] ),
    .A(\inv_in[2575] ));
 sg13g2_inv_2 \inv[2576]/_0_  (.Y(\inv_in[2577] ),
    .A(\inv_in[2576] ));
 sg13g2_inv_2 \inv[2577]/_0_  (.Y(\inv_in[2578] ),
    .A(\inv_in[2577] ));
 sg13g2_inv_2 \inv[2578]/_0_  (.Y(\inv_in[2579] ),
    .A(\inv_in[2578] ));
 sg13g2_inv_2 \inv[2579]/_0_  (.Y(\inv_in[2580] ),
    .A(\inv_in[2579] ));
 sg13g2_inv_2 \inv[257]/_0_  (.Y(\inv_in[258] ),
    .A(\inv_in[257] ));
 sg13g2_inv_2 \inv[2580]/_0_  (.Y(\inv_in[2581] ),
    .A(\inv_in[2580] ));
 sg13g2_inv_2 \inv[2581]/_0_  (.Y(\inv_in[2582] ),
    .A(\inv_in[2581] ));
 sg13g2_inv_2 \inv[2582]/_0_  (.Y(\inv_in[2583] ),
    .A(\inv_in[2582] ));
 sg13g2_inv_2 \inv[2583]/_0_  (.Y(\inv_in[2584] ),
    .A(\inv_in[2583] ));
 sg13g2_inv_2 \inv[2584]/_0_  (.Y(\inv_in[2585] ),
    .A(\inv_in[2584] ));
 sg13g2_inv_2 \inv[2585]/_0_  (.Y(\inv_in[2586] ),
    .A(\inv_in[2585] ));
 sg13g2_inv_2 \inv[2586]/_0_  (.Y(\inv_in[2587] ),
    .A(\inv_in[2586] ));
 sg13g2_inv_2 \inv[2587]/_0_  (.Y(\inv_in[2588] ),
    .A(\inv_in[2587] ));
 sg13g2_inv_2 \inv[2588]/_0_  (.Y(\inv_in[2589] ),
    .A(\inv_in[2588] ));
 sg13g2_inv_2 \inv[2589]/_0_  (.Y(\inv_in[2590] ),
    .A(\inv_in[2589] ));
 sg13g2_inv_2 \inv[258]/_0_  (.Y(\inv_in[259] ),
    .A(\inv_in[258] ));
 sg13g2_inv_2 \inv[2590]/_0_  (.Y(\inv_in[2591] ),
    .A(\inv_in[2590] ));
 sg13g2_inv_2 \inv[2591]/_0_  (.Y(\inv_in[2592] ),
    .A(\inv_in[2591] ));
 sg13g2_inv_2 \inv[2592]/_0_  (.Y(\inv_in[2593] ),
    .A(\inv_in[2592] ));
 sg13g2_inv_2 \inv[2593]/_0_  (.Y(\inv_in[2594] ),
    .A(\inv_in[2593] ));
 sg13g2_inv_2 \inv[2594]/_0_  (.Y(\inv_in[2595] ),
    .A(\inv_in[2594] ));
 sg13g2_inv_2 \inv[2595]/_0_  (.Y(\inv_in[2596] ),
    .A(\inv_in[2595] ));
 sg13g2_inv_2 \inv[2596]/_0_  (.Y(\inv_in[2597] ),
    .A(\inv_in[2596] ));
 sg13g2_inv_2 \inv[2597]/_0_  (.Y(\inv_in[2598] ),
    .A(\inv_in[2597] ));
 sg13g2_inv_2 \inv[2598]/_0_  (.Y(\inv_in[2599] ),
    .A(\inv_in[2598] ));
 sg13g2_inv_2 \inv[2599]/_0_  (.Y(\inv_in[2600] ),
    .A(\inv_in[2599] ));
 sg13g2_inv_2 \inv[259]/_0_  (.Y(\inv_in[260] ),
    .A(\inv_in[259] ));
 sg13g2_inv_2 \inv[25]/_0_  (.Y(\inv_in[26] ),
    .A(\inv_in[25] ));
 sg13g2_inv_2 \inv[2600]/_0_  (.Y(\inv_in[2601] ),
    .A(\inv_in[2600] ));
 sg13g2_inv_2 \inv[2601]/_0_  (.Y(\inv_in[2602] ),
    .A(\inv_in[2601] ));
 sg13g2_inv_2 \inv[2602]/_0_  (.Y(\inv_in[2603] ),
    .A(\inv_in[2602] ));
 sg13g2_inv_2 \inv[2603]/_0_  (.Y(\inv_in[2604] ),
    .A(\inv_in[2603] ));
 sg13g2_inv_2 \inv[2604]/_0_  (.Y(\inv_in[2605] ),
    .A(\inv_in[2604] ));
 sg13g2_inv_2 \inv[2605]/_0_  (.Y(\inv_in[2606] ),
    .A(\inv_in[2605] ));
 sg13g2_inv_2 \inv[2606]/_0_  (.Y(\inv_in[2607] ),
    .A(\inv_in[2606] ));
 sg13g2_inv_2 \inv[2607]/_0_  (.Y(\inv_in[2608] ),
    .A(\inv_in[2607] ));
 sg13g2_inv_2 \inv[2608]/_0_  (.Y(\inv_in[2609] ),
    .A(\inv_in[2608] ));
 sg13g2_inv_2 \inv[2609]/_0_  (.Y(\inv_in[2610] ),
    .A(\inv_in[2609] ));
 sg13g2_inv_4 \inv[260]/_0_  (.A(\inv_in[260] ),
    .Y(\inv_in[261] ));
 sg13g2_inv_2 \inv[2610]/_0_  (.Y(\inv_in[2611] ),
    .A(\inv_in[2610] ));
 sg13g2_inv_2 \inv[2611]/_0_  (.Y(\inv_in[2612] ),
    .A(\inv_in[2611] ));
 sg13g2_inv_2 \inv[2612]/_0_  (.Y(\inv_in[2613] ),
    .A(\inv_in[2612] ));
 sg13g2_inv_2 \inv[2613]/_0_  (.Y(\inv_in[2614] ),
    .A(\inv_in[2613] ));
 sg13g2_inv_2 \inv[2614]/_0_  (.Y(\inv_in[2615] ),
    .A(\inv_in[2614] ));
 sg13g2_inv_2 \inv[2615]/_0_  (.Y(\inv_in[2616] ),
    .A(\inv_in[2615] ));
 sg13g2_inv_2 \inv[2616]/_0_  (.Y(\inv_in[2617] ),
    .A(\inv_in[2616] ));
 sg13g2_inv_2 \inv[2617]/_0_  (.Y(\inv_in[2618] ),
    .A(\inv_in[2617] ));
 sg13g2_inv_2 \inv[2618]/_0_  (.Y(\inv_in[2619] ),
    .A(\inv_in[2618] ));
 sg13g2_inv_2 \inv[2619]/_0_  (.Y(\inv_in[2620] ),
    .A(\inv_in[2619] ));
 sg13g2_inv_4 \inv[261]/_0_  (.A(\inv_in[261] ),
    .Y(\inv_in[262] ));
 sg13g2_inv_2 \inv[2620]/_0_  (.Y(\inv_in[2621] ),
    .A(\inv_in[2620] ));
 sg13g2_inv_2 \inv[2621]/_0_  (.Y(\inv_in[2622] ),
    .A(\inv_in[2621] ));
 sg13g2_inv_2 \inv[2622]/_0_  (.Y(\inv_in[2623] ),
    .A(\inv_in[2622] ));
 sg13g2_inv_2 \inv[2623]/_0_  (.Y(\inv_in[2624] ),
    .A(\inv_in[2623] ));
 sg13g2_inv_2 \inv[2624]/_0_  (.Y(\inv_in[2625] ),
    .A(\inv_in[2624] ));
 sg13g2_inv_2 \inv[2625]/_0_  (.Y(\inv_in[2626] ),
    .A(\inv_in[2625] ));
 sg13g2_inv_2 \inv[2626]/_0_  (.Y(\inv_in[2627] ),
    .A(\inv_in[2626] ));
 sg13g2_inv_2 \inv[2627]/_0_  (.Y(\inv_in[2628] ),
    .A(\inv_in[2627] ));
 sg13g2_inv_2 \inv[2628]/_0_  (.Y(\inv_in[2629] ),
    .A(\inv_in[2628] ));
 sg13g2_inv_2 \inv[2629]/_0_  (.Y(\inv_in[2630] ),
    .A(\inv_in[2629] ));
 sg13g2_inv_4 \inv[262]/_0_  (.A(\inv_in[262] ),
    .Y(\inv_in[263] ));
 sg13g2_inv_2 \inv[2630]/_0_  (.Y(\inv_in[2631] ),
    .A(\inv_in[2630] ));
 sg13g2_inv_2 \inv[2631]/_0_  (.Y(\inv_in[2632] ),
    .A(\inv_in[2631] ));
 sg13g2_inv_2 \inv[2632]/_0_  (.Y(\inv_in[2633] ),
    .A(\inv_in[2632] ));
 sg13g2_inv_2 \inv[2633]/_0_  (.Y(\inv_in[2634] ),
    .A(\inv_in[2633] ));
 sg13g2_inv_2 \inv[2634]/_0_  (.Y(\inv_in[2635] ),
    .A(\inv_in[2634] ));
 sg13g2_inv_2 \inv[2635]/_0_  (.Y(\inv_in[2636] ),
    .A(\inv_in[2635] ));
 sg13g2_inv_2 \inv[2636]/_0_  (.Y(\inv_in[2637] ),
    .A(\inv_in[2636] ));
 sg13g2_inv_2 \inv[2637]/_0_  (.Y(\inv_in[2638] ),
    .A(\inv_in[2637] ));
 sg13g2_inv_2 \inv[2638]/_0_  (.Y(\inv_in[2639] ),
    .A(\inv_in[2638] ));
 sg13g2_inv_2 \inv[2639]/_0_  (.Y(\inv_in[2640] ),
    .A(\inv_in[2639] ));
 sg13g2_inv_4 \inv[263]/_0_  (.A(\inv_in[263] ),
    .Y(\inv_in[264] ));
 sg13g2_inv_2 \inv[2640]/_0_  (.Y(\inv_in[2641] ),
    .A(\inv_in[2640] ));
 sg13g2_inv_2 \inv[2641]/_0_  (.Y(\inv_in[2642] ),
    .A(\inv_in[2641] ));
 sg13g2_inv_2 \inv[2642]/_0_  (.Y(\inv_in[2643] ),
    .A(\inv_in[2642] ));
 sg13g2_inv_2 \inv[2643]/_0_  (.Y(\inv_in[2644] ),
    .A(\inv_in[2643] ));
 sg13g2_inv_2 \inv[2644]/_0_  (.Y(\inv_in[2645] ),
    .A(\inv_in[2644] ));
 sg13g2_inv_2 \inv[2645]/_0_  (.Y(\inv_in[2646] ),
    .A(\inv_in[2645] ));
 sg13g2_inv_2 \inv[2646]/_0_  (.Y(\inv_in[2647] ),
    .A(\inv_in[2646] ));
 sg13g2_inv_2 \inv[2647]/_0_  (.Y(\inv_in[2648] ),
    .A(\inv_in[2647] ));
 sg13g2_inv_2 \inv[2648]/_0_  (.Y(\inv_in[2649] ),
    .A(\inv_in[2648] ));
 sg13g2_inv_2 \inv[2649]/_0_  (.Y(\inv_in[2650] ),
    .A(\inv_in[2649] ));
 sg13g2_inv_4 \inv[264]/_0_  (.A(\inv_in[264] ),
    .Y(\inv_in[265] ));
 sg13g2_inv_2 \inv[2650]/_0_  (.Y(\inv_in[2651] ),
    .A(\inv_in[2650] ));
 sg13g2_inv_2 \inv[2651]/_0_  (.Y(\inv_in[2652] ),
    .A(\inv_in[2651] ));
 sg13g2_inv_2 \inv[2652]/_0_  (.Y(\inv_in[2653] ),
    .A(\inv_in[2652] ));
 sg13g2_inv_2 \inv[2653]/_0_  (.Y(\inv_in[2654] ),
    .A(\inv_in[2653] ));
 sg13g2_inv_2 \inv[2654]/_0_  (.Y(\inv_in[2655] ),
    .A(\inv_in[2654] ));
 sg13g2_inv_2 \inv[2655]/_0_  (.Y(\inv_in[2656] ),
    .A(\inv_in[2655] ));
 sg13g2_inv_2 \inv[2656]/_0_  (.Y(\inv_in[2657] ),
    .A(\inv_in[2656] ));
 sg13g2_inv_2 \inv[2657]/_0_  (.Y(\inv_in[2658] ),
    .A(\inv_in[2657] ));
 sg13g2_inv_2 \inv[2658]/_0_  (.Y(\inv_in[2659] ),
    .A(\inv_in[2658] ));
 sg13g2_inv_2 \inv[2659]/_0_  (.Y(\inv_in[2660] ),
    .A(\inv_in[2659] ));
 sg13g2_inv_4 \inv[265]/_0_  (.A(\inv_in[265] ),
    .Y(\inv_in[266] ));
 sg13g2_inv_2 \inv[2660]/_0_  (.Y(\inv_in[2661] ),
    .A(\inv_in[2660] ));
 sg13g2_inv_2 \inv[2661]/_0_  (.Y(\inv_in[2662] ),
    .A(\inv_in[2661] ));
 sg13g2_inv_2 \inv[2662]/_0_  (.Y(\inv_in[2663] ),
    .A(\inv_in[2662] ));
 sg13g2_inv_2 \inv[2663]/_0_  (.Y(\inv_in[2664] ),
    .A(\inv_in[2663] ));
 sg13g2_inv_2 \inv[2664]/_0_  (.Y(\inv_in[2665] ),
    .A(\inv_in[2664] ));
 sg13g2_inv_2 \inv[2665]/_0_  (.Y(\inv_in[2666] ),
    .A(\inv_in[2665] ));
 sg13g2_inv_2 \inv[2666]/_0_  (.Y(\inv_in[2667] ),
    .A(\inv_in[2666] ));
 sg13g2_inv_2 \inv[2667]/_0_  (.Y(\inv_in[2668] ),
    .A(\inv_in[2667] ));
 sg13g2_inv_2 \inv[2668]/_0_  (.Y(\inv_in[2669] ),
    .A(\inv_in[2668] ));
 sg13g2_inv_2 \inv[2669]/_0_  (.Y(\inv_in[2670] ),
    .A(\inv_in[2669] ));
 sg13g2_inv_4 \inv[266]/_0_  (.A(\inv_in[266] ),
    .Y(\inv_in[267] ));
 sg13g2_inv_2 \inv[2670]/_0_  (.Y(\inv_in[2671] ),
    .A(\inv_in[2670] ));
 sg13g2_inv_2 \inv[2671]/_0_  (.Y(\inv_in[2672] ),
    .A(\inv_in[2671] ));
 sg13g2_inv_2 \inv[2672]/_0_  (.Y(\inv_in[2673] ),
    .A(\inv_in[2672] ));
 sg13g2_inv_2 \inv[2673]/_0_  (.Y(\inv_in[2674] ),
    .A(\inv_in[2673] ));
 sg13g2_inv_2 \inv[2674]/_0_  (.Y(\inv_in[2675] ),
    .A(\inv_in[2674] ));
 sg13g2_inv_2 \inv[2675]/_0_  (.Y(\inv_in[2676] ),
    .A(\inv_in[2675] ));
 sg13g2_inv_2 \inv[2676]/_0_  (.Y(\inv_in[2677] ),
    .A(\inv_in[2676] ));
 sg13g2_inv_2 \inv[2677]/_0_  (.Y(\inv_in[2678] ),
    .A(\inv_in[2677] ));
 sg13g2_inv_2 \inv[2678]/_0_  (.Y(\inv_in[2679] ),
    .A(\inv_in[2678] ));
 sg13g2_inv_2 \inv[2679]/_0_  (.Y(\inv_in[2680] ),
    .A(\inv_in[2679] ));
 sg13g2_inv_4 \inv[267]/_0_  (.A(\inv_in[267] ),
    .Y(\inv_in[268] ));
 sg13g2_inv_2 \inv[2680]/_0_  (.Y(\inv_in[2681] ),
    .A(\inv_in[2680] ));
 sg13g2_inv_2 \inv[2681]/_0_  (.Y(\inv_in[2682] ),
    .A(\inv_in[2681] ));
 sg13g2_inv_2 \inv[2682]/_0_  (.Y(\inv_in[2683] ),
    .A(\inv_in[2682] ));
 sg13g2_inv_2 \inv[2683]/_0_  (.Y(\inv_in[2684] ),
    .A(\inv_in[2683] ));
 sg13g2_inv_2 \inv[2684]/_0_  (.Y(\inv_in[2685] ),
    .A(\inv_in[2684] ));
 sg13g2_inv_2 \inv[2685]/_0_  (.Y(\inv_in[2686] ),
    .A(\inv_in[2685] ));
 sg13g2_inv_2 \inv[2686]/_0_  (.Y(\inv_in[2687] ),
    .A(\inv_in[2686] ));
 sg13g2_inv_2 \inv[2687]/_0_  (.Y(\inv_in[2688] ),
    .A(\inv_in[2687] ));
 sg13g2_inv_2 \inv[2688]/_0_  (.Y(\inv_in[2689] ),
    .A(\inv_in[2688] ));
 sg13g2_inv_2 \inv[2689]/_0_  (.Y(\inv_in[2690] ),
    .A(\inv_in[2689] ));
 sg13g2_inv_4 \inv[268]/_0_  (.A(\inv_in[268] ),
    .Y(\inv_in[269] ));
 sg13g2_inv_2 \inv[2690]/_0_  (.Y(\inv_in[2691] ),
    .A(\inv_in[2690] ));
 sg13g2_inv_2 \inv[2691]/_0_  (.Y(\inv_in[2692] ),
    .A(\inv_in[2691] ));
 sg13g2_inv_2 \inv[2692]/_0_  (.Y(\inv_in[2693] ),
    .A(\inv_in[2692] ));
 sg13g2_inv_2 \inv[2693]/_0_  (.Y(\inv_in[2694] ),
    .A(\inv_in[2693] ));
 sg13g2_inv_2 \inv[2694]/_0_  (.Y(\inv_in[2695] ),
    .A(\inv_in[2694] ));
 sg13g2_inv_2 \inv[2695]/_0_  (.Y(\inv_in[2696] ),
    .A(\inv_in[2695] ));
 sg13g2_inv_2 \inv[2696]/_0_  (.Y(\inv_in[2697] ),
    .A(\inv_in[2696] ));
 sg13g2_inv_2 \inv[2697]/_0_  (.Y(\inv_in[2698] ),
    .A(\inv_in[2697] ));
 sg13g2_inv_2 \inv[2698]/_0_  (.Y(\inv_in[2699] ),
    .A(\inv_in[2698] ));
 sg13g2_inv_2 \inv[2699]/_0_  (.Y(\inv_in[2700] ),
    .A(\inv_in[2699] ));
 sg13g2_inv_4 \inv[269]/_0_  (.A(\inv_in[269] ),
    .Y(\inv_in[270] ));
 sg13g2_inv_2 \inv[26]/_0_  (.Y(\inv_in[27] ),
    .A(\inv_in[26] ));
 sg13g2_inv_2 \inv[2700]/_0_  (.Y(\inv_in[2701] ),
    .A(\inv_in[2700] ));
 sg13g2_inv_2 \inv[2701]/_0_  (.Y(\inv_in[2702] ),
    .A(\inv_in[2701] ));
 sg13g2_inv_2 \inv[2702]/_0_  (.Y(\inv_in[2703] ),
    .A(\inv_in[2702] ));
 sg13g2_inv_2 \inv[2703]/_0_  (.Y(\inv_in[2704] ),
    .A(\inv_in[2703] ));
 sg13g2_inv_2 \inv[2704]/_0_  (.Y(\inv_in[2705] ),
    .A(\inv_in[2704] ));
 sg13g2_inv_2 \inv[2705]/_0_  (.Y(\inv_in[2706] ),
    .A(\inv_in[2705] ));
 sg13g2_inv_2 \inv[2706]/_0_  (.Y(\inv_in[2707] ),
    .A(\inv_in[2706] ));
 sg13g2_inv_2 \inv[2707]/_0_  (.Y(\inv_in[2708] ),
    .A(\inv_in[2707] ));
 sg13g2_inv_2 \inv[2708]/_0_  (.Y(\inv_in[2709] ),
    .A(\inv_in[2708] ));
 sg13g2_inv_2 \inv[2709]/_0_  (.Y(\inv_in[2710] ),
    .A(\inv_in[2709] ));
 sg13g2_inv_2 \inv[270]/_0_  (.Y(\inv_in[271] ),
    .A(\inv_in[270] ));
 sg13g2_inv_2 \inv[2710]/_0_  (.Y(\inv_in[2711] ),
    .A(\inv_in[2710] ));
 sg13g2_inv_2 \inv[2711]/_0_  (.Y(\inv_in[2712] ),
    .A(\inv_in[2711] ));
 sg13g2_inv_2 \inv[2712]/_0_  (.Y(\inv_in[2713] ),
    .A(\inv_in[2712] ));
 sg13g2_inv_2 \inv[2713]/_0_  (.Y(\inv_in[2714] ),
    .A(\inv_in[2713] ));
 sg13g2_inv_2 \inv[2714]/_0_  (.Y(\inv_in[2715] ),
    .A(\inv_in[2714] ));
 sg13g2_inv_4 \inv[2715]/_0_  (.A(\inv_in[2715] ),
    .Y(\inv_in[2716] ));
 sg13g2_inv_4 \inv[2716]/_0_  (.A(\inv_in[2716] ),
    .Y(\inv_in[2717] ));
 sg13g2_inv_4 \inv[2717]/_0_  (.A(\inv_in[2717] ),
    .Y(\inv_in[2718] ));
 sg13g2_inv_2 \inv[2718]/_0_  (.Y(\inv_in[2719] ),
    .A(\inv_in[2718] ));
 sg13g2_inv_2 \inv[2719]/_0_  (.Y(\inv_in[2720] ),
    .A(\inv_in[2719] ));
 sg13g2_inv_2 \inv[271]/_0_  (.Y(\inv_in[272] ),
    .A(\inv_in[271] ));
 sg13g2_inv_2 \inv[2720]/_0_  (.Y(\inv_in[2721] ),
    .A(\inv_in[2720] ));
 sg13g2_inv_2 \inv[2721]/_0_  (.Y(\inv_in[2722] ),
    .A(\inv_in[2721] ));
 sg13g2_inv_2 \inv[2722]/_0_  (.Y(\inv_in[2723] ),
    .A(\inv_in[2722] ));
 sg13g2_inv_2 \inv[2723]/_0_  (.Y(\inv_in[2724] ),
    .A(\inv_in[2723] ));
 sg13g2_inv_2 \inv[2724]/_0_  (.Y(\inv_in[2725] ),
    .A(\inv_in[2724] ));
 sg13g2_inv_2 \inv[2725]/_0_  (.Y(\inv_in[2726] ),
    .A(\inv_in[2725] ));
 sg13g2_inv_2 \inv[2726]/_0_  (.Y(\inv_in[2727] ),
    .A(\inv_in[2726] ));
 sg13g2_inv_2 \inv[2727]/_0_  (.Y(\inv_in[2728] ),
    .A(\inv_in[2727] ));
 sg13g2_inv_2 \inv[2728]/_0_  (.Y(\inv_in[2729] ),
    .A(\inv_in[2728] ));
 sg13g2_inv_2 \inv[2729]/_0_  (.Y(\inv_in[2730] ),
    .A(\inv_in[2729] ));
 sg13g2_inv_4 \inv[272]/_0_  (.A(\inv_in[272] ),
    .Y(\inv_in[273] ));
 sg13g2_inv_2 \inv[2730]/_0_  (.Y(\inv_in[2731] ),
    .A(\inv_in[2730] ));
 sg13g2_inv_2 \inv[2731]/_0_  (.Y(\inv_in[2732] ),
    .A(\inv_in[2731] ));
 sg13g2_inv_2 \inv[2732]/_0_  (.Y(\inv_in[2733] ),
    .A(\inv_in[2732] ));
 sg13g2_inv_2 \inv[2733]/_0_  (.Y(\inv_in[2734] ),
    .A(\inv_in[2733] ));
 sg13g2_inv_2 \inv[2734]/_0_  (.Y(\inv_in[2735] ),
    .A(\inv_in[2734] ));
 sg13g2_inv_2 \inv[2735]/_0_  (.Y(\inv_in[2736] ),
    .A(\inv_in[2735] ));
 sg13g2_inv_2 \inv[2736]/_0_  (.Y(\inv_in[2737] ),
    .A(\inv_in[2736] ));
 sg13g2_inv_2 \inv[2737]/_0_  (.Y(\inv_in[2738] ),
    .A(\inv_in[2737] ));
 sg13g2_inv_2 \inv[2738]/_0_  (.Y(\inv_in[2739] ),
    .A(\inv_in[2738] ));
 sg13g2_inv_2 \inv[2739]/_0_  (.Y(\inv_in[2740] ),
    .A(\inv_in[2739] ));
 sg13g2_inv_4 \inv[273]/_0_  (.A(\inv_in[273] ),
    .Y(\inv_in[274] ));
 sg13g2_inv_2 \inv[2740]/_0_  (.Y(\inv_in[2741] ),
    .A(\inv_in[2740] ));
 sg13g2_inv_2 \inv[2741]/_0_  (.Y(\inv_in[2742] ),
    .A(\inv_in[2741] ));
 sg13g2_inv_2 \inv[2742]/_0_  (.Y(\inv_in[2743] ),
    .A(\inv_in[2742] ));
 sg13g2_inv_2 \inv[2743]/_0_  (.Y(\inv_in[2744] ),
    .A(\inv_in[2743] ));
 sg13g2_inv_2 \inv[2744]/_0_  (.Y(\inv_in[2745] ),
    .A(\inv_in[2744] ));
 sg13g2_inv_2 \inv[2745]/_0_  (.Y(\inv_in[2746] ),
    .A(\inv_in[2745] ));
 sg13g2_inv_2 \inv[2746]/_0_  (.Y(\inv_in[2747] ),
    .A(\inv_in[2746] ));
 sg13g2_inv_2 \inv[2747]/_0_  (.Y(\inv_in[2748] ),
    .A(\inv_in[2747] ));
 sg13g2_inv_2 \inv[2748]/_0_  (.Y(\inv_in[2749] ),
    .A(\inv_in[2748] ));
 sg13g2_inv_2 \inv[2749]/_0_  (.Y(\inv_in[2750] ),
    .A(\inv_in[2749] ));
 sg13g2_inv_4 \inv[274]/_0_  (.A(\inv_in[274] ),
    .Y(\inv_in[275] ));
 sg13g2_inv_2 \inv[2750]/_0_  (.Y(\inv_in[2751] ),
    .A(\inv_in[2750] ));
 sg13g2_inv_2 \inv[2751]/_0_  (.Y(\inv_in[2752] ),
    .A(\inv_in[2751] ));
 sg13g2_inv_2 \inv[2752]/_0_  (.Y(\inv_in[2753] ),
    .A(\inv_in[2752] ));
 sg13g2_inv_2 \inv[2753]/_0_  (.Y(\inv_in[2754] ),
    .A(\inv_in[2753] ));
 sg13g2_inv_2 \inv[2754]/_0_  (.Y(\inv_in[2755] ),
    .A(\inv_in[2754] ));
 sg13g2_inv_2 \inv[2755]/_0_  (.Y(\inv_in[2756] ),
    .A(\inv_in[2755] ));
 sg13g2_inv_2 \inv[2756]/_0_  (.Y(\inv_in[2757] ),
    .A(\inv_in[2756] ));
 sg13g2_inv_2 \inv[2757]/_0_  (.Y(\inv_in[2758] ),
    .A(\inv_in[2757] ));
 sg13g2_inv_2 \inv[2758]/_0_  (.Y(\inv_in[2759] ),
    .A(\inv_in[2758] ));
 sg13g2_inv_2 \inv[2759]/_0_  (.Y(\inv_in[2760] ),
    .A(\inv_in[2759] ));
 sg13g2_inv_4 \inv[275]/_0_  (.A(\inv_in[275] ),
    .Y(\inv_in[276] ));
 sg13g2_inv_2 \inv[2760]/_0_  (.Y(\inv_in[2761] ),
    .A(\inv_in[2760] ));
 sg13g2_inv_2 \inv[2761]/_0_  (.Y(\inv_in[2762] ),
    .A(\inv_in[2761] ));
 sg13g2_inv_2 \inv[2762]/_0_  (.Y(\inv_in[2763] ),
    .A(\inv_in[2762] ));
 sg13g2_inv_2 \inv[2763]/_0_  (.Y(\inv_in[2764] ),
    .A(\inv_in[2763] ));
 sg13g2_inv_2 \inv[2764]/_0_  (.Y(\inv_in[2765] ),
    .A(\inv_in[2764] ));
 sg13g2_inv_2 \inv[2765]/_0_  (.Y(\inv_in[2766] ),
    .A(\inv_in[2765] ));
 sg13g2_inv_2 \inv[2766]/_0_  (.Y(\inv_in[2767] ),
    .A(\inv_in[2766] ));
 sg13g2_inv_2 \inv[2767]/_0_  (.Y(\inv_in[2768] ),
    .A(\inv_in[2767] ));
 sg13g2_inv_2 \inv[2768]/_0_  (.Y(\inv_in[2769] ),
    .A(\inv_in[2768] ));
 sg13g2_inv_2 \inv[2769]/_0_  (.Y(\inv_in[2770] ),
    .A(\inv_in[2769] ));
 sg13g2_inv_4 \inv[276]/_0_  (.A(\inv_in[276] ),
    .Y(\inv_in[277] ));
 sg13g2_inv_2 \inv[2770]/_0_  (.Y(\inv_in[2771] ),
    .A(\inv_in[2770] ));
 sg13g2_inv_2 \inv[2771]/_0_  (.Y(\inv_in[2772] ),
    .A(\inv_in[2771] ));
 sg13g2_inv_2 \inv[2772]/_0_  (.Y(\inv_in[2773] ),
    .A(\inv_in[2772] ));
 sg13g2_inv_2 \inv[2773]/_0_  (.Y(\inv_in[2774] ),
    .A(\inv_in[2773] ));
 sg13g2_inv_2 \inv[2774]/_0_  (.Y(\inv_in[2775] ),
    .A(\inv_in[2774] ));
 sg13g2_inv_2 \inv[2775]/_0_  (.Y(\inv_in[2776] ),
    .A(\inv_in[2775] ));
 sg13g2_inv_2 \inv[2776]/_0_  (.Y(\inv_in[2777] ),
    .A(\inv_in[2776] ));
 sg13g2_inv_2 \inv[2777]/_0_  (.Y(\inv_in[2778] ),
    .A(\inv_in[2777] ));
 sg13g2_inv_2 \inv[2778]/_0_  (.Y(\inv_in[2779] ),
    .A(\inv_in[2778] ));
 sg13g2_inv_2 \inv[2779]/_0_  (.Y(\inv_in[2780] ),
    .A(\inv_in[2779] ));
 sg13g2_inv_2 \inv[277]/_0_  (.Y(\inv_in[278] ),
    .A(\inv_in[277] ));
 sg13g2_inv_2 \inv[2780]/_0_  (.Y(\inv_in[2781] ),
    .A(\inv_in[2780] ));
 sg13g2_inv_2 \inv[2781]/_0_  (.Y(\inv_in[2782] ),
    .A(\inv_in[2781] ));
 sg13g2_inv_2 \inv[2782]/_0_  (.Y(\inv_in[2783] ),
    .A(\inv_in[2782] ));
 sg13g2_inv_2 \inv[2783]/_0_  (.Y(\inv_in[2784] ),
    .A(\inv_in[2783] ));
 sg13g2_inv_2 \inv[2784]/_0_  (.Y(\inv_in[2785] ),
    .A(\inv_in[2784] ));
 sg13g2_inv_2 \inv[2785]/_0_  (.Y(\inv_in[2786] ),
    .A(\inv_in[2785] ));
 sg13g2_inv_2 \inv[2786]/_0_  (.Y(\inv_in[2787] ),
    .A(\inv_in[2786] ));
 sg13g2_inv_2 \inv[2787]/_0_  (.Y(\inv_in[2788] ),
    .A(\inv_in[2787] ));
 sg13g2_inv_2 \inv[2788]/_0_  (.Y(\inv_in[2789] ),
    .A(\inv_in[2788] ));
 sg13g2_inv_2 \inv[2789]/_0_  (.Y(\inv_in[2790] ),
    .A(\inv_in[2789] ));
 sg13g2_inv_2 \inv[278]/_0_  (.Y(\inv_in[279] ),
    .A(\inv_in[278] ));
 sg13g2_inv_2 \inv[2790]/_0_  (.Y(\inv_in[2791] ),
    .A(\inv_in[2790] ));
 sg13g2_inv_2 \inv[2791]/_0_  (.Y(\inv_in[2792] ),
    .A(\inv_in[2791] ));
 sg13g2_inv_2 \inv[2792]/_0_  (.Y(\inv_in[2793] ),
    .A(\inv_in[2792] ));
 sg13g2_inv_2 \inv[2793]/_0_  (.Y(\inv_in[2794] ),
    .A(\inv_in[2793] ));
 sg13g2_inv_2 \inv[2794]/_0_  (.Y(\inv_in[2795] ),
    .A(\inv_in[2794] ));
 sg13g2_inv_2 \inv[2795]/_0_  (.Y(\inv_in[2796] ),
    .A(\inv_in[2795] ));
 sg13g2_inv_2 \inv[2796]/_0_  (.Y(\inv_in[2797] ),
    .A(\inv_in[2796] ));
 sg13g2_inv_2 \inv[2797]/_0_  (.Y(\inv_in[2798] ),
    .A(\inv_in[2797] ));
 sg13g2_inv_2 \inv[2798]/_0_  (.Y(\inv_in[2799] ),
    .A(\inv_in[2798] ));
 sg13g2_inv_2 \inv[2799]/_0_  (.Y(\inv_in[2800] ),
    .A(\inv_in[2799] ));
 sg13g2_inv_2 \inv[279]/_0_  (.Y(\inv_in[280] ),
    .A(\inv_in[279] ));
 sg13g2_inv_2 \inv[27]/_0_  (.Y(\inv_in[28] ),
    .A(\inv_in[27] ));
 sg13g2_inv_2 \inv[2800]/_0_  (.Y(\inv_in[2801] ),
    .A(\inv_in[2800] ));
 sg13g2_inv_2 \inv[2801]/_0_  (.Y(\inv_in[2802] ),
    .A(\inv_in[2801] ));
 sg13g2_inv_2 \inv[2802]/_0_  (.Y(\inv_in[2803] ),
    .A(\inv_in[2802] ));
 sg13g2_inv_2 \inv[2803]/_0_  (.Y(\inv_in[2804] ),
    .A(\inv_in[2803] ));
 sg13g2_inv_2 \inv[2804]/_0_  (.Y(\inv_in[2805] ),
    .A(\inv_in[2804] ));
 sg13g2_inv_2 \inv[2805]/_0_  (.Y(\inv_in[2806] ),
    .A(\inv_in[2805] ));
 sg13g2_inv_2 \inv[2806]/_0_  (.Y(\inv_in[2807] ),
    .A(\inv_in[2806] ));
 sg13g2_inv_2 \inv[2807]/_0_  (.Y(\inv_in[2808] ),
    .A(\inv_in[2807] ));
 sg13g2_inv_2 \inv[2808]/_0_  (.Y(\inv_in[2809] ),
    .A(\inv_in[2808] ));
 sg13g2_inv_2 \inv[2809]/_0_  (.Y(\inv_in[2810] ),
    .A(\inv_in[2809] ));
 sg13g2_inv_2 \inv[280]/_0_  (.Y(\inv_in[281] ),
    .A(\inv_in[280] ));
 sg13g2_inv_2 \inv[2810]/_0_  (.Y(\inv_in[2811] ),
    .A(\inv_in[2810] ));
 sg13g2_inv_2 \inv[2811]/_0_  (.Y(\inv_in[2812] ),
    .A(\inv_in[2811] ));
 sg13g2_inv_2 \inv[2812]/_0_  (.Y(\inv_in[2813] ),
    .A(\inv_in[2812] ));
 sg13g2_inv_2 \inv[2813]/_0_  (.Y(\inv_in[2814] ),
    .A(\inv_in[2813] ));
 sg13g2_inv_2 \inv[2814]/_0_  (.Y(\inv_in[2815] ),
    .A(\inv_in[2814] ));
 sg13g2_inv_2 \inv[2815]/_0_  (.Y(\inv_in[2816] ),
    .A(\inv_in[2815] ));
 sg13g2_inv_2 \inv[2816]/_0_  (.Y(\inv_in[2817] ),
    .A(\inv_in[2816] ));
 sg13g2_inv_2 \inv[2817]/_0_  (.Y(\inv_in[2818] ),
    .A(\inv_in[2817] ));
 sg13g2_inv_2 \inv[2818]/_0_  (.Y(\inv_in[2819] ),
    .A(\inv_in[2818] ));
 sg13g2_inv_2 \inv[2819]/_0_  (.Y(\inv_in[2820] ),
    .A(\inv_in[2819] ));
 sg13g2_inv_2 \inv[281]/_0_  (.Y(\inv_in[282] ),
    .A(\inv_in[281] ));
 sg13g2_inv_2 \inv[2820]/_0_  (.Y(\inv_in[2821] ),
    .A(\inv_in[2820] ));
 sg13g2_inv_2 \inv[2821]/_0_  (.Y(\inv_in[2822] ),
    .A(\inv_in[2821] ));
 sg13g2_inv_2 \inv[2822]/_0_  (.Y(\inv_in[2823] ),
    .A(\inv_in[2822] ));
 sg13g2_inv_2 \inv[2823]/_0_  (.Y(\inv_in[2824] ),
    .A(\inv_in[2823] ));
 sg13g2_inv_2 \inv[2824]/_0_  (.Y(\inv_in[2825] ),
    .A(\inv_in[2824] ));
 sg13g2_inv_2 \inv[2825]/_0_  (.Y(\inv_in[2826] ),
    .A(\inv_in[2825] ));
 sg13g2_inv_2 \inv[2826]/_0_  (.Y(\inv_in[2827] ),
    .A(\inv_in[2826] ));
 sg13g2_inv_2 \inv[2827]/_0_  (.Y(\inv_in[2828] ),
    .A(\inv_in[2827] ));
 sg13g2_inv_2 \inv[2828]/_0_  (.Y(\inv_in[2829] ),
    .A(\inv_in[2828] ));
 sg13g2_inv_2 \inv[2829]/_0_  (.Y(\inv_in[2830] ),
    .A(\inv_in[2829] ));
 sg13g2_inv_2 \inv[282]/_0_  (.Y(\inv_in[283] ),
    .A(\inv_in[282] ));
 sg13g2_inv_2 \inv[2830]/_0_  (.Y(\inv_in[2831] ),
    .A(\inv_in[2830] ));
 sg13g2_inv_2 \inv[2831]/_0_  (.Y(\inv_in[2832] ),
    .A(\inv_in[2831] ));
 sg13g2_inv_2 \inv[2832]/_0_  (.Y(\inv_in[2833] ),
    .A(\inv_in[2832] ));
 sg13g2_inv_2 \inv[2833]/_0_  (.Y(\inv_in[2834] ),
    .A(\inv_in[2833] ));
 sg13g2_inv_2 \inv[2834]/_0_  (.Y(\inv_in[2835] ),
    .A(\inv_in[2834] ));
 sg13g2_inv_2 \inv[2835]/_0_  (.Y(\inv_in[2836] ),
    .A(\inv_in[2835] ));
 sg13g2_inv_2 \inv[2836]/_0_  (.Y(\inv_in[2837] ),
    .A(\inv_in[2836] ));
 sg13g2_inv_2 \inv[2837]/_0_  (.Y(\inv_in[2838] ),
    .A(\inv_in[2837] ));
 sg13g2_inv_2 \inv[2838]/_0_  (.Y(\inv_in[2839] ),
    .A(\inv_in[2838] ));
 sg13g2_inv_2 \inv[2839]/_0_  (.Y(\inv_in[2840] ),
    .A(\inv_in[2839] ));
 sg13g2_inv_2 \inv[283]/_0_  (.Y(\inv_in[284] ),
    .A(\inv_in[283] ));
 sg13g2_inv_2 \inv[2840]/_0_  (.Y(\inv_in[2841] ),
    .A(\inv_in[2840] ));
 sg13g2_inv_2 \inv[2841]/_0_  (.Y(\inv_in[2842] ),
    .A(\inv_in[2841] ));
 sg13g2_inv_2 \inv[2842]/_0_  (.Y(\inv_in[2843] ),
    .A(\inv_in[2842] ));
 sg13g2_inv_2 \inv[2843]/_0_  (.Y(\inv_in[2844] ),
    .A(\inv_in[2843] ));
 sg13g2_inv_2 \inv[2844]/_0_  (.Y(\inv_in[2845] ),
    .A(\inv_in[2844] ));
 sg13g2_inv_2 \inv[2845]/_0_  (.Y(\inv_in[2846] ),
    .A(\inv_in[2845] ));
 sg13g2_inv_2 \inv[2846]/_0_  (.Y(\inv_in[2847] ),
    .A(\inv_in[2846] ));
 sg13g2_inv_2 \inv[2847]/_0_  (.Y(\inv_in[2848] ),
    .A(\inv_in[2847] ));
 sg13g2_inv_2 \inv[2848]/_0_  (.Y(\inv_in[2849] ),
    .A(\inv_in[2848] ));
 sg13g2_inv_2 \inv[2849]/_0_  (.Y(\inv_in[2850] ),
    .A(\inv_in[2849] ));
 sg13g2_inv_2 \inv[284]/_0_  (.Y(\inv_in[285] ),
    .A(\inv_in[284] ));
 sg13g2_inv_2 \inv[2850]/_0_  (.Y(\inv_in[2851] ),
    .A(\inv_in[2850] ));
 sg13g2_inv_2 \inv[2851]/_0_  (.Y(\inv_in[2852] ),
    .A(\inv_in[2851] ));
 sg13g2_inv_2 \inv[2852]/_0_  (.Y(\inv_in[2853] ),
    .A(\inv_in[2852] ));
 sg13g2_inv_2 \inv[2853]/_0_  (.Y(\inv_in[2854] ),
    .A(\inv_in[2853] ));
 sg13g2_inv_2 \inv[2854]/_0_  (.Y(\inv_in[2855] ),
    .A(\inv_in[2854] ));
 sg13g2_inv_2 \inv[2855]/_0_  (.Y(\inv_in[2856] ),
    .A(\inv_in[2855] ));
 sg13g2_inv_2 \inv[2856]/_0_  (.Y(\inv_in[2857] ),
    .A(\inv_in[2856] ));
 sg13g2_inv_2 \inv[2857]/_0_  (.Y(\inv_in[2858] ),
    .A(\inv_in[2857] ));
 sg13g2_inv_2 \inv[2858]/_0_  (.Y(\inv_in[2859] ),
    .A(\inv_in[2858] ));
 sg13g2_inv_2 \inv[2859]/_0_  (.Y(\inv_in[2860] ),
    .A(\inv_in[2859] ));
 sg13g2_inv_2 \inv[285]/_0_  (.Y(\inv_in[286] ),
    .A(\inv_in[285] ));
 sg13g2_inv_2 \inv[2860]/_0_  (.Y(\inv_in[2861] ),
    .A(\inv_in[2860] ));
 sg13g2_inv_2 \inv[2861]/_0_  (.Y(\inv_in[2862] ),
    .A(\inv_in[2861] ));
 sg13g2_inv_2 \inv[2862]/_0_  (.Y(\inv_in[2863] ),
    .A(\inv_in[2862] ));
 sg13g2_inv_2 \inv[2863]/_0_  (.Y(\inv_in[2864] ),
    .A(\inv_in[2863] ));
 sg13g2_inv_2 \inv[2864]/_0_  (.Y(\inv_in[2865] ),
    .A(\inv_in[2864] ));
 sg13g2_inv_2 \inv[2865]/_0_  (.Y(\inv_in[2866] ),
    .A(\inv_in[2865] ));
 sg13g2_inv_2 \inv[2866]/_0_  (.Y(\inv_in[2867] ),
    .A(\inv_in[2866] ));
 sg13g2_inv_2 \inv[2867]/_0_  (.Y(\inv_in[2868] ),
    .A(\inv_in[2867] ));
 sg13g2_inv_2 \inv[2868]/_0_  (.Y(\inv_in[2869] ),
    .A(\inv_in[2868] ));
 sg13g2_inv_2 \inv[2869]/_0_  (.Y(\inv_in[2870] ),
    .A(\inv_in[2869] ));
 sg13g2_inv_2 \inv[286]/_0_  (.Y(\inv_in[287] ),
    .A(\inv_in[286] ));
 sg13g2_inv_2 \inv[2870]/_0_  (.Y(\inv_in[2871] ),
    .A(\inv_in[2870] ));
 sg13g2_inv_2 \inv[2871]/_0_  (.Y(\inv_in[2872] ),
    .A(\inv_in[2871] ));
 sg13g2_inv_2 \inv[2872]/_0_  (.Y(\inv_in[2873] ),
    .A(\inv_in[2872] ));
 sg13g2_inv_2 \inv[2873]/_0_  (.Y(\inv_in[2874] ),
    .A(\inv_in[2873] ));
 sg13g2_inv_2 \inv[2874]/_0_  (.Y(\inv_in[2875] ),
    .A(\inv_in[2874] ));
 sg13g2_inv_2 \inv[2875]/_0_  (.Y(\inv_in[2876] ),
    .A(\inv_in[2875] ));
 sg13g2_inv_2 \inv[2876]/_0_  (.Y(\inv_in[2877] ),
    .A(\inv_in[2876] ));
 sg13g2_inv_2 \inv[2877]/_0_  (.Y(\inv_in[2878] ),
    .A(\inv_in[2877] ));
 sg13g2_inv_2 \inv[2878]/_0_  (.Y(\inv_in[2879] ),
    .A(\inv_in[2878] ));
 sg13g2_inv_2 \inv[2879]/_0_  (.Y(\inv_in[2880] ),
    .A(\inv_in[2879] ));
 sg13g2_inv_2 \inv[287]/_0_  (.Y(\inv_in[288] ),
    .A(\inv_in[287] ));
 sg13g2_inv_2 \inv[2880]/_0_  (.Y(\inv_in[2881] ),
    .A(\inv_in[2880] ));
 sg13g2_inv_2 \inv[2881]/_0_  (.Y(\inv_in[2882] ),
    .A(\inv_in[2881] ));
 sg13g2_inv_2 \inv[2882]/_0_  (.Y(\inv_in[2883] ),
    .A(\inv_in[2882] ));
 sg13g2_inv_2 \inv[2883]/_0_  (.Y(\inv_in[2884] ),
    .A(\inv_in[2883] ));
 sg13g2_inv_2 \inv[2884]/_0_  (.Y(\inv_in[2885] ),
    .A(\inv_in[2884] ));
 sg13g2_inv_2 \inv[2885]/_0_  (.Y(\inv_in[2886] ),
    .A(\inv_in[2885] ));
 sg13g2_inv_2 \inv[2886]/_0_  (.Y(\inv_in[2887] ),
    .A(\inv_in[2886] ));
 sg13g2_inv_2 \inv[2887]/_0_  (.Y(\inv_in[2888] ),
    .A(\inv_in[2887] ));
 sg13g2_inv_2 \inv[2888]/_0_  (.Y(\inv_in[2889] ),
    .A(\inv_in[2888] ));
 sg13g2_inv_2 \inv[2889]/_0_  (.Y(\inv_in[2890] ),
    .A(\inv_in[2889] ));
 sg13g2_inv_2 \inv[288]/_0_  (.Y(\inv_in[289] ),
    .A(\inv_in[288] ));
 sg13g2_inv_2 \inv[2890]/_0_  (.Y(\inv_in[2891] ),
    .A(\inv_in[2890] ));
 sg13g2_inv_2 \inv[2891]/_0_  (.Y(\inv_in[2892] ),
    .A(\inv_in[2891] ));
 sg13g2_inv_2 \inv[2892]/_0_  (.Y(\inv_in[2893] ),
    .A(\inv_in[2892] ));
 sg13g2_inv_2 \inv[2893]/_0_  (.Y(\inv_in[2894] ),
    .A(\inv_in[2893] ));
 sg13g2_inv_2 \inv[2894]/_0_  (.Y(\inv_in[2895] ),
    .A(\inv_in[2894] ));
 sg13g2_inv_2 \inv[2895]/_0_  (.Y(\inv_in[2896] ),
    .A(\inv_in[2895] ));
 sg13g2_inv_2 \inv[2896]/_0_  (.Y(\inv_in[2897] ),
    .A(\inv_in[2896] ));
 sg13g2_inv_2 \inv[2897]/_0_  (.Y(\inv_in[2898] ),
    .A(\inv_in[2897] ));
 sg13g2_inv_2 \inv[2898]/_0_  (.Y(\inv_in[2899] ),
    .A(\inv_in[2898] ));
 sg13g2_inv_2 \inv[2899]/_0_  (.Y(\inv_in[2900] ),
    .A(\inv_in[2899] ));
 sg13g2_inv_2 \inv[289]/_0_  (.Y(\inv_in[290] ),
    .A(\inv_in[289] ));
 sg13g2_inv_2 \inv[28]/_0_  (.Y(\inv_in[29] ),
    .A(\inv_in[28] ));
 sg13g2_inv_2 \inv[2900]/_0_  (.Y(\inv_in[2901] ),
    .A(\inv_in[2900] ));
 sg13g2_inv_2 \inv[2901]/_0_  (.Y(\inv_in[2902] ),
    .A(\inv_in[2901] ));
 sg13g2_inv_2 \inv[2902]/_0_  (.Y(\inv_in[2903] ),
    .A(\inv_in[2902] ));
 sg13g2_inv_2 \inv[2903]/_0_  (.Y(\inv_in[2904] ),
    .A(\inv_in[2903] ));
 sg13g2_inv_2 \inv[2904]/_0_  (.Y(\inv_in[2905] ),
    .A(\inv_in[2904] ));
 sg13g2_inv_2 \inv[2905]/_0_  (.Y(\inv_in[2906] ),
    .A(\inv_in[2905] ));
 sg13g2_inv_2 \inv[2906]/_0_  (.Y(\inv_in[2907] ),
    .A(\inv_in[2906] ));
 sg13g2_inv_2 \inv[2907]/_0_  (.Y(\inv_in[2908] ),
    .A(\inv_in[2907] ));
 sg13g2_inv_2 \inv[2908]/_0_  (.Y(\inv_in[2909] ),
    .A(\inv_in[2908] ));
 sg13g2_inv_2 \inv[2909]/_0_  (.Y(\inv_in[2910] ),
    .A(\inv_in[2909] ));
 sg13g2_inv_2 \inv[290]/_0_  (.Y(\inv_in[291] ),
    .A(\inv_in[290] ));
 sg13g2_inv_2 \inv[2910]/_0_  (.Y(\inv_in[2911] ),
    .A(\inv_in[2910] ));
 sg13g2_inv_2 \inv[2911]/_0_  (.Y(\inv_in[2912] ),
    .A(\inv_in[2911] ));
 sg13g2_inv_2 \inv[2912]/_0_  (.Y(\inv_in[2913] ),
    .A(\inv_in[2912] ));
 sg13g2_inv_2 \inv[2913]/_0_  (.Y(\inv_in[2914] ),
    .A(\inv_in[2913] ));
 sg13g2_inv_2 \inv[2914]/_0_  (.Y(\inv_in[2915] ),
    .A(\inv_in[2914] ));
 sg13g2_inv_2 \inv[2915]/_0_  (.Y(\inv_in[2916] ),
    .A(\inv_in[2915] ));
 sg13g2_inv_2 \inv[2916]/_0_  (.Y(\inv_in[2917] ),
    .A(\inv_in[2916] ));
 sg13g2_inv_2 \inv[2917]/_0_  (.Y(\inv_in[2918] ),
    .A(\inv_in[2917] ));
 sg13g2_inv_2 \inv[2918]/_0_  (.Y(\inv_in[2919] ),
    .A(\inv_in[2918] ));
 sg13g2_inv_2 \inv[2919]/_0_  (.Y(\inv_in[2920] ),
    .A(\inv_in[2919] ));
 sg13g2_inv_2 \inv[291]/_0_  (.Y(\inv_in[292] ),
    .A(\inv_in[291] ));
 sg13g2_inv_2 \inv[2920]/_0_  (.Y(\inv_in[2921] ),
    .A(\inv_in[2920] ));
 sg13g2_inv_2 \inv[2921]/_0_  (.Y(\inv_in[2922] ),
    .A(\inv_in[2921] ));
 sg13g2_inv_2 \inv[2922]/_0_  (.Y(\inv_in[2923] ),
    .A(\inv_in[2922] ));
 sg13g2_inv_2 \inv[2923]/_0_  (.Y(\inv_in[2924] ),
    .A(\inv_in[2923] ));
 sg13g2_inv_2 \inv[2924]/_0_  (.Y(\inv_in[2925] ),
    .A(\inv_in[2924] ));
 sg13g2_inv_2 \inv[2925]/_0_  (.Y(\inv_in[2926] ),
    .A(\inv_in[2925] ));
 sg13g2_inv_2 \inv[2926]/_0_  (.Y(\inv_in[2927] ),
    .A(\inv_in[2926] ));
 sg13g2_inv_2 \inv[2927]/_0_  (.Y(\inv_in[2928] ),
    .A(\inv_in[2927] ));
 sg13g2_inv_2 \inv[2928]/_0_  (.Y(\inv_in[2929] ),
    .A(\inv_in[2928] ));
 sg13g2_inv_2 \inv[2929]/_0_  (.Y(\inv_in[2930] ),
    .A(\inv_in[2929] ));
 sg13g2_inv_2 \inv[292]/_0_  (.Y(\inv_in[293] ),
    .A(\inv_in[292] ));
 sg13g2_inv_2 \inv[2930]/_0_  (.Y(\inv_in[2931] ),
    .A(\inv_in[2930] ));
 sg13g2_inv_2 \inv[2931]/_0_  (.Y(\inv_in[2932] ),
    .A(\inv_in[2931] ));
 sg13g2_inv_2 \inv[2932]/_0_  (.Y(\inv_in[2933] ),
    .A(\inv_in[2932] ));
 sg13g2_inv_2 \inv[2933]/_0_  (.Y(\inv_in[2934] ),
    .A(\inv_in[2933] ));
 sg13g2_inv_2 \inv[2934]/_0_  (.Y(\inv_in[2935] ),
    .A(\inv_in[2934] ));
 sg13g2_inv_2 \inv[2935]/_0_  (.Y(\inv_in[2936] ),
    .A(\inv_in[2935] ));
 sg13g2_inv_2 \inv[2936]/_0_  (.Y(\inv_in[2937] ),
    .A(\inv_in[2936] ));
 sg13g2_inv_2 \inv[2937]/_0_  (.Y(\inv_in[2938] ),
    .A(\inv_in[2937] ));
 sg13g2_inv_2 \inv[2938]/_0_  (.Y(\inv_in[2939] ),
    .A(\inv_in[2938] ));
 sg13g2_inv_2 \inv[2939]/_0_  (.Y(\inv_in[2940] ),
    .A(\inv_in[2939] ));
 sg13g2_inv_2 \inv[293]/_0_  (.Y(\inv_in[294] ),
    .A(\inv_in[293] ));
 sg13g2_inv_2 \inv[2940]/_0_  (.Y(\inv_in[2941] ),
    .A(\inv_in[2940] ));
 sg13g2_inv_2 \inv[2941]/_0_  (.Y(\inv_in[2942] ),
    .A(\inv_in[2941] ));
 sg13g2_inv_2 \inv[2942]/_0_  (.Y(\inv_in[2943] ),
    .A(\inv_in[2942] ));
 sg13g2_inv_2 \inv[2943]/_0_  (.Y(\inv_in[2944] ),
    .A(\inv_in[2943] ));
 sg13g2_inv_2 \inv[2944]/_0_  (.Y(\inv_in[2945] ),
    .A(\inv_in[2944] ));
 sg13g2_inv_2 \inv[2945]/_0_  (.Y(\inv_in[2946] ),
    .A(\inv_in[2945] ));
 sg13g2_inv_2 \inv[2946]/_0_  (.Y(\inv_in[2947] ),
    .A(\inv_in[2946] ));
 sg13g2_inv_2 \inv[2947]/_0_  (.Y(\inv_in[2948] ),
    .A(\inv_in[2947] ));
 sg13g2_inv_2 \inv[2948]/_0_  (.Y(\inv_in[2949] ),
    .A(\inv_in[2948] ));
 sg13g2_inv_2 \inv[2949]/_0_  (.Y(\inv_in[2950] ),
    .A(\inv_in[2949] ));
 sg13g2_inv_2 \inv[294]/_0_  (.Y(\inv_in[295] ),
    .A(\inv_in[294] ));
 sg13g2_inv_2 \inv[2950]/_0_  (.Y(\inv_in[2951] ),
    .A(\inv_in[2950] ));
 sg13g2_inv_2 \inv[2951]/_0_  (.Y(\inv_in[2952] ),
    .A(\inv_in[2951] ));
 sg13g2_inv_2 \inv[2952]/_0_  (.Y(\inv_in[2953] ),
    .A(\inv_in[2952] ));
 sg13g2_inv_2 \inv[2953]/_0_  (.Y(\inv_in[2954] ),
    .A(\inv_in[2953] ));
 sg13g2_inv_2 \inv[2954]/_0_  (.Y(\inv_in[2955] ),
    .A(\inv_in[2954] ));
 sg13g2_inv_2 \inv[2955]/_0_  (.Y(\inv_in[2956] ),
    .A(\inv_in[2955] ));
 sg13g2_inv_2 \inv[2956]/_0_  (.Y(\inv_in[2957] ),
    .A(\inv_in[2956] ));
 sg13g2_inv_2 \inv[2957]/_0_  (.Y(\inv_in[2958] ),
    .A(\inv_in[2957] ));
 sg13g2_inv_2 \inv[2958]/_0_  (.Y(\inv_in[2959] ),
    .A(\inv_in[2958] ));
 sg13g2_inv_2 \inv[2959]/_0_  (.Y(\inv_in[2960] ),
    .A(\inv_in[2959] ));
 sg13g2_inv_2 \inv[295]/_0_  (.Y(\inv_in[296] ),
    .A(\inv_in[295] ));
 sg13g2_inv_2 \inv[2960]/_0_  (.Y(\inv_in[2961] ),
    .A(\inv_in[2960] ));
 sg13g2_inv_2 \inv[2961]/_0_  (.Y(\inv_in[2962] ),
    .A(\inv_in[2961] ));
 sg13g2_inv_2 \inv[2962]/_0_  (.Y(\inv_in[2963] ),
    .A(\inv_in[2962] ));
 sg13g2_inv_2 \inv[2963]/_0_  (.Y(\inv_in[2964] ),
    .A(\inv_in[2963] ));
 sg13g2_inv_2 \inv[2964]/_0_  (.Y(\inv_in[2965] ),
    .A(\inv_in[2964] ));
 sg13g2_inv_2 \inv[2965]/_0_  (.Y(\inv_in[2966] ),
    .A(\inv_in[2965] ));
 sg13g2_inv_2 \inv[2966]/_0_  (.Y(\inv_in[2967] ),
    .A(\inv_in[2966] ));
 sg13g2_inv_2 \inv[2967]/_0_  (.Y(\inv_in[2968] ),
    .A(\inv_in[2967] ));
 sg13g2_inv_2 \inv[2968]/_0_  (.Y(\inv_in[2969] ),
    .A(\inv_in[2968] ));
 sg13g2_inv_2 \inv[2969]/_0_  (.Y(\inv_in[2970] ),
    .A(\inv_in[2969] ));
 sg13g2_inv_2 \inv[296]/_0_  (.Y(\inv_in[297] ),
    .A(\inv_in[296] ));
 sg13g2_inv_2 \inv[2970]/_0_  (.Y(\inv_in[2971] ),
    .A(\inv_in[2970] ));
 sg13g2_inv_2 \inv[2971]/_0_  (.Y(\inv_in[2972] ),
    .A(\inv_in[2971] ));
 sg13g2_inv_2 \inv[2972]/_0_  (.Y(\inv_in[2973] ),
    .A(\inv_in[2972] ));
 sg13g2_inv_2 \inv[2973]/_0_  (.Y(\inv_in[2974] ),
    .A(\inv_in[2973] ));
 sg13g2_inv_2 \inv[2974]/_0_  (.Y(\inv_in[2975] ),
    .A(\inv_in[2974] ));
 sg13g2_inv_2 \inv[2975]/_0_  (.Y(\inv_in[2976] ),
    .A(\inv_in[2975] ));
 sg13g2_inv_2 \inv[2976]/_0_  (.Y(\inv_in[2977] ),
    .A(\inv_in[2976] ));
 sg13g2_inv_2 \inv[2977]/_0_  (.Y(\inv_in[2978] ),
    .A(\inv_in[2977] ));
 sg13g2_inv_2 \inv[2978]/_0_  (.Y(\inv_in[2979] ),
    .A(\inv_in[2978] ));
 sg13g2_inv_2 \inv[2979]/_0_  (.Y(\inv_in[2980] ),
    .A(\inv_in[2979] ));
 sg13g2_inv_2 \inv[297]/_0_  (.Y(\inv_in[298] ),
    .A(\inv_in[297] ));
 sg13g2_inv_2 \inv[2980]/_0_  (.Y(\inv_in[2981] ),
    .A(\inv_in[2980] ));
 sg13g2_inv_2 \inv[2981]/_0_  (.Y(\inv_in[2982] ),
    .A(\inv_in[2981] ));
 sg13g2_inv_2 \inv[2982]/_0_  (.Y(\inv_in[2983] ),
    .A(\inv_in[2982] ));
 sg13g2_inv_2 \inv[2983]/_0_  (.Y(\inv_in[2984] ),
    .A(\inv_in[2983] ));
 sg13g2_inv_2 \inv[2984]/_0_  (.Y(\inv_in[2985] ),
    .A(\inv_in[2984] ));
 sg13g2_inv_2 \inv[2985]/_0_  (.Y(\inv_in[2986] ),
    .A(\inv_in[2985] ));
 sg13g2_inv_2 \inv[2986]/_0_  (.Y(\inv_in[2987] ),
    .A(\inv_in[2986] ));
 sg13g2_inv_2 \inv[2987]/_0_  (.Y(\inv_in[2988] ),
    .A(\inv_in[2987] ));
 sg13g2_inv_2 \inv[2988]/_0_  (.Y(\inv_in[2989] ),
    .A(\inv_in[2988] ));
 sg13g2_inv_2 \inv[2989]/_0_  (.Y(\inv_in[2990] ),
    .A(\inv_in[2989] ));
 sg13g2_inv_2 \inv[298]/_0_  (.Y(\inv_in[299] ),
    .A(\inv_in[298] ));
 sg13g2_inv_2 \inv[2990]/_0_  (.Y(\inv_in[2991] ),
    .A(\inv_in[2990] ));
 sg13g2_inv_2 \inv[2991]/_0_  (.Y(\inv_in[2992] ),
    .A(\inv_in[2991] ));
 sg13g2_inv_2 \inv[2992]/_0_  (.Y(\inv_in[2993] ),
    .A(\inv_in[2992] ));
 sg13g2_inv_2 \inv[2993]/_0_  (.Y(\inv_in[2994] ),
    .A(\inv_in[2993] ));
 sg13g2_inv_2 \inv[2994]/_0_  (.Y(\inv_in[2995] ),
    .A(\inv_in[2994] ));
 sg13g2_inv_2 \inv[2995]/_0_  (.Y(\inv_in[2996] ),
    .A(\inv_in[2995] ));
 sg13g2_inv_2 \inv[2996]/_0_  (.Y(\inv_in[2997] ),
    .A(\inv_in[2996] ));
 sg13g2_inv_2 \inv[2997]/_0_  (.Y(\inv_in[2998] ),
    .A(\inv_in[2997] ));
 sg13g2_inv_2 \inv[2998]/_0_  (.Y(\inv_in[2999] ),
    .A(\inv_in[2998] ));
 sg13g2_inv_2 \inv[2999]/_0_  (.Y(\inv_in[3000] ),
    .A(\inv_in[2999] ));
 sg13g2_inv_2 \inv[299]/_0_  (.Y(\inv_in[300] ),
    .A(\inv_in[299] ));
 sg13g2_inv_2 \inv[29]/_0_  (.Y(\inv_in[30] ),
    .A(\inv_in[29] ));
 sg13g2_inv_4 \inv[2]/_0_  (.A(\inv_in[2] ),
    .Y(\inv_in[3] ));
 sg13g2_inv_2 \inv[3000]/_0_  (.Y(\inv_in[3001] ),
    .A(\inv_in[3000] ));
 sg13g2_inv_2 \inv[3001]/_0_  (.Y(\inv_in[3002] ),
    .A(\inv_in[3001] ));
 sg13g2_inv_2 \inv[3002]/_0_  (.Y(\inv_in[3003] ),
    .A(\inv_in[3002] ));
 sg13g2_inv_2 \inv[3003]/_0_  (.Y(\inv_in[3004] ),
    .A(\inv_in[3003] ));
 sg13g2_inv_2 \inv[3004]/_0_  (.Y(\inv_in[3005] ),
    .A(\inv_in[3004] ));
 sg13g2_inv_2 \inv[3005]/_0_  (.Y(\inv_in[3006] ),
    .A(\inv_in[3005] ));
 sg13g2_inv_2 \inv[3006]/_0_  (.Y(\inv_in[3007] ),
    .A(\inv_in[3006] ));
 sg13g2_inv_2 \inv[3007]/_0_  (.Y(\inv_in[3008] ),
    .A(\inv_in[3007] ));
 sg13g2_inv_2 \inv[3008]/_0_  (.Y(\inv_in[3009] ),
    .A(\inv_in[3008] ));
 sg13g2_inv_2 \inv[3009]/_0_  (.Y(\inv_in[3010] ),
    .A(\inv_in[3009] ));
 sg13g2_inv_2 \inv[300]/_0_  (.Y(\inv_in[301] ),
    .A(\inv_in[300] ));
 sg13g2_inv_2 \inv[3010]/_0_  (.Y(\inv_in[3011] ),
    .A(\inv_in[3010] ));
 sg13g2_inv_2 \inv[3011]/_0_  (.Y(\inv_in[3012] ),
    .A(\inv_in[3011] ));
 sg13g2_inv_2 \inv[3012]/_0_  (.Y(\inv_in[3013] ),
    .A(\inv_in[3012] ));
 sg13g2_inv_2 \inv[3013]/_0_  (.Y(\inv_in[3014] ),
    .A(\inv_in[3013] ));
 sg13g2_inv_2 \inv[3014]/_0_  (.Y(\inv_in[3015] ),
    .A(\inv_in[3014] ));
 sg13g2_inv_2 \inv[3015]/_0_  (.Y(\inv_in[3016] ),
    .A(\inv_in[3015] ));
 sg13g2_inv_2 \inv[3016]/_0_  (.Y(\inv_in[3017] ),
    .A(\inv_in[3016] ));
 sg13g2_inv_2 \inv[3017]/_0_  (.Y(\inv_in[3018] ),
    .A(\inv_in[3017] ));
 sg13g2_inv_2 \inv[3018]/_0_  (.Y(\inv_in[3019] ),
    .A(\inv_in[3018] ));
 sg13g2_inv_2 \inv[3019]/_0_  (.Y(\inv_in[3020] ),
    .A(\inv_in[3019] ));
 sg13g2_inv_2 \inv[301]/_0_  (.Y(\inv_in[302] ),
    .A(\inv_in[301] ));
 sg13g2_inv_2 \inv[3020]/_0_  (.Y(\inv_in[3021] ),
    .A(\inv_in[3020] ));
 sg13g2_inv_2 \inv[3021]/_0_  (.Y(\inv_in[3022] ),
    .A(\inv_in[3021] ));
 sg13g2_inv_2 \inv[3022]/_0_  (.Y(\inv_in[3023] ),
    .A(\inv_in[3022] ));
 sg13g2_inv_2 \inv[3023]/_0_  (.Y(\inv_in[3024] ),
    .A(\inv_in[3023] ));
 sg13g2_inv_2 \inv[3024]/_0_  (.Y(\inv_in[3025] ),
    .A(\inv_in[3024] ));
 sg13g2_inv_2 \inv[3025]/_0_  (.Y(\inv_in[3026] ),
    .A(\inv_in[3025] ));
 sg13g2_inv_2 \inv[3026]/_0_  (.Y(\inv_in[3027] ),
    .A(\inv_in[3026] ));
 sg13g2_inv_2 \inv[3027]/_0_  (.Y(\inv_in[3028] ),
    .A(\inv_in[3027] ));
 sg13g2_inv_2 \inv[3028]/_0_  (.Y(\inv_in[3029] ),
    .A(\inv_in[3028] ));
 sg13g2_inv_2 \inv[3029]/_0_  (.Y(\inv_in[3030] ),
    .A(\inv_in[3029] ));
 sg13g2_inv_2 \inv[302]/_0_  (.Y(\inv_in[303] ),
    .A(\inv_in[302] ));
 sg13g2_inv_2 \inv[3030]/_0_  (.Y(\inv_in[3031] ),
    .A(\inv_in[3030] ));
 sg13g2_inv_2 \inv[3031]/_0_  (.Y(\inv_in[3032] ),
    .A(\inv_in[3031] ));
 sg13g2_inv_2 \inv[3032]/_0_  (.Y(\inv_in[3033] ),
    .A(\inv_in[3032] ));
 sg13g2_inv_2 \inv[3033]/_0_  (.Y(\inv_in[3034] ),
    .A(\inv_in[3033] ));
 sg13g2_inv_2 \inv[3034]/_0_  (.Y(\inv_in[3035] ),
    .A(\inv_in[3034] ));
 sg13g2_inv_2 \inv[3035]/_0_  (.Y(\inv_in[3036] ),
    .A(\inv_in[3035] ));
 sg13g2_inv_2 \inv[3036]/_0_  (.Y(\inv_in[3037] ),
    .A(\inv_in[3036] ));
 sg13g2_inv_2 \inv[3037]/_0_  (.Y(\inv_in[3038] ),
    .A(\inv_in[3037] ));
 sg13g2_inv_2 \inv[3038]/_0_  (.Y(\inv_in[3039] ),
    .A(\inv_in[3038] ));
 sg13g2_inv_2 \inv[3039]/_0_  (.Y(\inv_in[3040] ),
    .A(\inv_in[3039] ));
 sg13g2_inv_2 \inv[303]/_0_  (.Y(\inv_in[304] ),
    .A(\inv_in[303] ));
 sg13g2_inv_2 \inv[3040]/_0_  (.Y(\inv_in[3041] ),
    .A(\inv_in[3040] ));
 sg13g2_inv_2 \inv[3041]/_0_  (.Y(\inv_in[3042] ),
    .A(\inv_in[3041] ));
 sg13g2_inv_2 \inv[3042]/_0_  (.Y(\inv_in[3043] ),
    .A(\inv_in[3042] ));
 sg13g2_inv_2 \inv[3043]/_0_  (.Y(\inv_in[3044] ),
    .A(\inv_in[3043] ));
 sg13g2_inv_2 \inv[3044]/_0_  (.Y(\inv_in[3045] ),
    .A(\inv_in[3044] ));
 sg13g2_inv_2 \inv[3045]/_0_  (.Y(\inv_in[3046] ),
    .A(\inv_in[3045] ));
 sg13g2_inv_2 \inv[3046]/_0_  (.Y(\inv_in[3047] ),
    .A(\inv_in[3046] ));
 sg13g2_inv_2 \inv[3047]/_0_  (.Y(\inv_in[3048] ),
    .A(\inv_in[3047] ));
 sg13g2_inv_2 \inv[3048]/_0_  (.Y(\inv_in[3049] ),
    .A(\inv_in[3048] ));
 sg13g2_inv_2 \inv[3049]/_0_  (.Y(\inv_in[3050] ),
    .A(\inv_in[3049] ));
 sg13g2_inv_2 \inv[304]/_0_  (.Y(\inv_in[305] ),
    .A(\inv_in[304] ));
 sg13g2_inv_2 \inv[3050]/_0_  (.Y(\inv_in[3051] ),
    .A(\inv_in[3050] ));
 sg13g2_inv_2 \inv[3051]/_0_  (.Y(\inv_in[3052] ),
    .A(\inv_in[3051] ));
 sg13g2_inv_2 \inv[3052]/_0_  (.Y(\inv_in[3053] ),
    .A(\inv_in[3052] ));
 sg13g2_inv_2 \inv[3053]/_0_  (.Y(\inv_in[3054] ),
    .A(\inv_in[3053] ));
 sg13g2_inv_2 \inv[3054]/_0_  (.Y(\inv_in[3055] ),
    .A(\inv_in[3054] ));
 sg13g2_inv_2 \inv[3055]/_0_  (.Y(\inv_in[3056] ),
    .A(\inv_in[3055] ));
 sg13g2_inv_2 \inv[3056]/_0_  (.Y(\inv_in[3057] ),
    .A(\inv_in[3056] ));
 sg13g2_inv_2 \inv[3057]/_0_  (.Y(\inv_in[3058] ),
    .A(\inv_in[3057] ));
 sg13g2_inv_2 \inv[3058]/_0_  (.Y(\inv_in[3059] ),
    .A(\inv_in[3058] ));
 sg13g2_inv_2 \inv[3059]/_0_  (.Y(\inv_in[3060] ),
    .A(\inv_in[3059] ));
 sg13g2_inv_2 \inv[305]/_0_  (.Y(\inv_in[306] ),
    .A(\inv_in[305] ));
 sg13g2_inv_2 \inv[3060]/_0_  (.Y(\inv_in[3061] ),
    .A(\inv_in[3060] ));
 sg13g2_inv_2 \inv[3061]/_0_  (.Y(\inv_in[3062] ),
    .A(\inv_in[3061] ));
 sg13g2_inv_2 \inv[3062]/_0_  (.Y(\inv_in[3063] ),
    .A(\inv_in[3062] ));
 sg13g2_inv_2 \inv[3063]/_0_  (.Y(\inv_in[3064] ),
    .A(\inv_in[3063] ));
 sg13g2_inv_2 \inv[3064]/_0_  (.Y(\inv_in[3065] ),
    .A(\inv_in[3064] ));
 sg13g2_inv_2 \inv[3065]/_0_  (.Y(\inv_in[3066] ),
    .A(\inv_in[3065] ));
 sg13g2_inv_2 \inv[3066]/_0_  (.Y(\inv_in[3067] ),
    .A(\inv_in[3066] ));
 sg13g2_inv_2 \inv[3067]/_0_  (.Y(\inv_in[3068] ),
    .A(\inv_in[3067] ));
 sg13g2_inv_2 \inv[3068]/_0_  (.Y(\inv_in[3069] ),
    .A(\inv_in[3068] ));
 sg13g2_inv_2 \inv[3069]/_0_  (.Y(\inv_in[3070] ),
    .A(\inv_in[3069] ));
 sg13g2_inv_2 \inv[306]/_0_  (.Y(\inv_in[307] ),
    .A(\inv_in[306] ));
 sg13g2_inv_2 \inv[3070]/_0_  (.Y(\inv_in[3071] ),
    .A(\inv_in[3070] ));
 sg13g2_inv_2 \inv[3071]/_0_  (.Y(\inv_in[3072] ),
    .A(\inv_in[3071] ));
 sg13g2_inv_2 \inv[3072]/_0_  (.Y(\inv_in[3073] ),
    .A(\inv_in[3072] ));
 sg13g2_inv_2 \inv[3073]/_0_  (.Y(\inv_in[3074] ),
    .A(\inv_in[3073] ));
 sg13g2_inv_2 \inv[3074]/_0_  (.Y(\inv_in[3075] ),
    .A(\inv_in[3074] ));
 sg13g2_inv_2 \inv[3075]/_0_  (.Y(\inv_in[3076] ),
    .A(\inv_in[3075] ));
 sg13g2_inv_2 \inv[3076]/_0_  (.Y(\inv_in[3077] ),
    .A(\inv_in[3076] ));
 sg13g2_inv_2 \inv[3077]/_0_  (.Y(\inv_in[3078] ),
    .A(\inv_in[3077] ));
 sg13g2_inv_2 \inv[3078]/_0_  (.Y(\inv_in[3079] ),
    .A(\inv_in[3078] ));
 sg13g2_inv_2 \inv[3079]/_0_  (.Y(\inv_in[3080] ),
    .A(\inv_in[3079] ));
 sg13g2_inv_2 \inv[307]/_0_  (.Y(\inv_in[308] ),
    .A(\inv_in[307] ));
 sg13g2_inv_2 \inv[3080]/_0_  (.Y(\inv_in[3081] ),
    .A(\inv_in[3080] ));
 sg13g2_inv_2 \inv[3081]/_0_  (.Y(\inv_in[3082] ),
    .A(\inv_in[3081] ));
 sg13g2_inv_2 \inv[3082]/_0_  (.Y(\inv_in[3083] ),
    .A(\inv_in[3082] ));
 sg13g2_inv_2 \inv[3083]/_0_  (.Y(\inv_in[3084] ),
    .A(\inv_in[3083] ));
 sg13g2_inv_2 \inv[3084]/_0_  (.Y(\inv_in[3085] ),
    .A(\inv_in[3084] ));
 sg13g2_inv_2 \inv[3085]/_0_  (.Y(\inv_in[3086] ),
    .A(\inv_in[3085] ));
 sg13g2_inv_2 \inv[3086]/_0_  (.Y(\inv_in[3087] ),
    .A(\inv_in[3086] ));
 sg13g2_inv_2 \inv[3087]/_0_  (.Y(\inv_in[3088] ),
    .A(\inv_in[3087] ));
 sg13g2_inv_2 \inv[3088]/_0_  (.Y(\inv_in[3089] ),
    .A(\inv_in[3088] ));
 sg13g2_inv_2 \inv[3089]/_0_  (.Y(\inv_in[3090] ),
    .A(\inv_in[3089] ));
 sg13g2_inv_2 \inv[308]/_0_  (.Y(\inv_in[309] ),
    .A(\inv_in[308] ));
 sg13g2_inv_2 \inv[3090]/_0_  (.Y(\inv_in[3091] ),
    .A(\inv_in[3090] ));
 sg13g2_inv_2 \inv[3091]/_0_  (.Y(\inv_in[3092] ),
    .A(\inv_in[3091] ));
 sg13g2_inv_2 \inv[3092]/_0_  (.Y(\inv_in[3093] ),
    .A(\inv_in[3092] ));
 sg13g2_inv_2 \inv[3093]/_0_  (.Y(\inv_in[3094] ),
    .A(\inv_in[3093] ));
 sg13g2_inv_2 \inv[3094]/_0_  (.Y(\inv_in[3095] ),
    .A(\inv_in[3094] ));
 sg13g2_inv_2 \inv[3095]/_0_  (.Y(\inv_in[3096] ),
    .A(\inv_in[3095] ));
 sg13g2_inv_2 \inv[3096]/_0_  (.Y(\inv_in[3097] ),
    .A(\inv_in[3096] ));
 sg13g2_inv_2 \inv[3097]/_0_  (.Y(\inv_in[3098] ),
    .A(\inv_in[3097] ));
 sg13g2_inv_2 \inv[3098]/_0_  (.Y(\inv_in[3099] ),
    .A(\inv_in[3098] ));
 sg13g2_inv_2 \inv[3099]/_0_  (.Y(\inv_in[3100] ),
    .A(\inv_in[3099] ));
 sg13g2_inv_2 \inv[309]/_0_  (.Y(\inv_in[310] ),
    .A(\inv_in[309] ));
 sg13g2_inv_2 \inv[30]/_0_  (.Y(\inv_in[31] ),
    .A(\inv_in[30] ));
 sg13g2_inv_2 \inv[3100]/_0_  (.Y(\inv_in[3101] ),
    .A(\inv_in[3100] ));
 sg13g2_inv_2 \inv[3101]/_0_  (.Y(\inv_in[3102] ),
    .A(\inv_in[3101] ));
 sg13g2_inv_2 \inv[3102]/_0_  (.Y(\inv_in[3103] ),
    .A(\inv_in[3102] ));
 sg13g2_inv_2 \inv[3103]/_0_  (.Y(\inv_in[3104] ),
    .A(\inv_in[3103] ));
 sg13g2_inv_2 \inv[3104]/_0_  (.Y(\inv_in[3105] ),
    .A(\inv_in[3104] ));
 sg13g2_inv_2 \inv[3105]/_0_  (.Y(\inv_in[3106] ),
    .A(\inv_in[3105] ));
 sg13g2_inv_2 \inv[3106]/_0_  (.Y(\inv_in[3107] ),
    .A(\inv_in[3106] ));
 sg13g2_inv_2 \inv[3107]/_0_  (.Y(\inv_in[3108] ),
    .A(\inv_in[3107] ));
 sg13g2_inv_2 \inv[3108]/_0_  (.Y(\inv_in[3109] ),
    .A(\inv_in[3108] ));
 sg13g2_inv_2 \inv[3109]/_0_  (.Y(\inv_in[3110] ),
    .A(\inv_in[3109] ));
 sg13g2_inv_2 \inv[310]/_0_  (.Y(\inv_in[311] ),
    .A(\inv_in[310] ));
 sg13g2_inv_2 \inv[3110]/_0_  (.Y(\inv_in[3111] ),
    .A(\inv_in[3110] ));
 sg13g2_inv_2 \inv[3111]/_0_  (.Y(\inv_in[3112] ),
    .A(\inv_in[3111] ));
 sg13g2_inv_2 \inv[3112]/_0_  (.Y(\inv_in[3113] ),
    .A(\inv_in[3112] ));
 sg13g2_inv_2 \inv[3113]/_0_  (.Y(\inv_in[3114] ),
    .A(\inv_in[3113] ));
 sg13g2_inv_2 \inv[3114]/_0_  (.Y(\inv_in[3115] ),
    .A(\inv_in[3114] ));
 sg13g2_inv_2 \inv[3115]/_0_  (.Y(\inv_in[3116] ),
    .A(\inv_in[3115] ));
 sg13g2_inv_2 \inv[3116]/_0_  (.Y(\inv_in[3117] ),
    .A(\inv_in[3116] ));
 sg13g2_inv_2 \inv[3117]/_0_  (.Y(\inv_in[3118] ),
    .A(\inv_in[3117] ));
 sg13g2_inv_2 \inv[3118]/_0_  (.Y(\inv_in[3119] ),
    .A(\inv_in[3118] ));
 sg13g2_inv_2 \inv[3119]/_0_  (.Y(\inv_in[3120] ),
    .A(\inv_in[3119] ));
 sg13g2_inv_2 \inv[311]/_0_  (.Y(\inv_in[312] ),
    .A(\inv_in[311] ));
 sg13g2_inv_2 \inv[3120]/_0_  (.Y(\inv_in[3121] ),
    .A(\inv_in[3120] ));
 sg13g2_inv_2 \inv[3121]/_0_  (.Y(\inv_in[3122] ),
    .A(\inv_in[3121] ));
 sg13g2_inv_2 \inv[3122]/_0_  (.Y(\inv_in[3123] ),
    .A(\inv_in[3122] ));
 sg13g2_inv_2 \inv[3123]/_0_  (.Y(\inv_in[3124] ),
    .A(\inv_in[3123] ));
 sg13g2_inv_2 \inv[3124]/_0_  (.Y(\inv_in[3125] ),
    .A(\inv_in[3124] ));
 sg13g2_inv_2 \inv[3125]/_0_  (.Y(\inv_in[3126] ),
    .A(\inv_in[3125] ));
 sg13g2_inv_2 \inv[3126]/_0_  (.Y(\inv_in[3127] ),
    .A(\inv_in[3126] ));
 sg13g2_inv_2 \inv[3127]/_0_  (.Y(\inv_in[3128] ),
    .A(\inv_in[3127] ));
 sg13g2_inv_2 \inv[3128]/_0_  (.Y(\inv_in[3129] ),
    .A(\inv_in[3128] ));
 sg13g2_inv_2 \inv[3129]/_0_  (.Y(\inv_in[3130] ),
    .A(\inv_in[3129] ));
 sg13g2_inv_2 \inv[312]/_0_  (.Y(\inv_in[313] ),
    .A(\inv_in[312] ));
 sg13g2_inv_2 \inv[3130]/_0_  (.Y(\inv_in[3131] ),
    .A(\inv_in[3130] ));
 sg13g2_inv_2 \inv[3131]/_0_  (.Y(\inv_in[3132] ),
    .A(\inv_in[3131] ));
 sg13g2_inv_2 \inv[3132]/_0_  (.Y(\inv_in[3133] ),
    .A(\inv_in[3132] ));
 sg13g2_inv_2 \inv[3133]/_0_  (.Y(\inv_in[3134] ),
    .A(\inv_in[3133] ));
 sg13g2_inv_2 \inv[3134]/_0_  (.Y(\inv_in[3135] ),
    .A(\inv_in[3134] ));
 sg13g2_inv_2 \inv[3135]/_0_  (.Y(\inv_in[3136] ),
    .A(\inv_in[3135] ));
 sg13g2_inv_2 \inv[3136]/_0_  (.Y(\inv_in[3137] ),
    .A(\inv_in[3136] ));
 sg13g2_inv_2 \inv[3137]/_0_  (.Y(\inv_in[3138] ),
    .A(\inv_in[3137] ));
 sg13g2_inv_2 \inv[3138]/_0_  (.Y(\inv_in[3139] ),
    .A(\inv_in[3138] ));
 sg13g2_inv_2 \inv[3139]/_0_  (.Y(\inv_in[3140] ),
    .A(\inv_in[3139] ));
 sg13g2_inv_2 \inv[313]/_0_  (.Y(\inv_in[314] ),
    .A(\inv_in[313] ));
 sg13g2_inv_2 \inv[3140]/_0_  (.Y(\inv_in[3141] ),
    .A(\inv_in[3140] ));
 sg13g2_inv_2 \inv[3141]/_0_  (.Y(\inv_in[3142] ),
    .A(\inv_in[3141] ));
 sg13g2_inv_2 \inv[3142]/_0_  (.Y(\inv_in[3143] ),
    .A(\inv_in[3142] ));
 sg13g2_inv_2 \inv[3143]/_0_  (.Y(\inv_in[3144] ),
    .A(\inv_in[3143] ));
 sg13g2_inv_2 \inv[3144]/_0_  (.Y(\inv_in[3145] ),
    .A(\inv_in[3144] ));
 sg13g2_inv_2 \inv[3145]/_0_  (.Y(\inv_in[3146] ),
    .A(\inv_in[3145] ));
 sg13g2_inv_2 \inv[3146]/_0_  (.Y(\inv_in[3147] ),
    .A(\inv_in[3146] ));
 sg13g2_inv_2 \inv[3147]/_0_  (.Y(\inv_in[3148] ),
    .A(\inv_in[3147] ));
 sg13g2_inv_2 \inv[3148]/_0_  (.Y(\inv_in[3149] ),
    .A(\inv_in[3148] ));
 sg13g2_inv_2 \inv[3149]/_0_  (.Y(\inv_in[3150] ),
    .A(\inv_in[3149] ));
 sg13g2_inv_2 \inv[314]/_0_  (.Y(\inv_in[315] ),
    .A(\inv_in[314] ));
 sg13g2_inv_2 \inv[3150]/_0_  (.Y(\inv_in[3151] ),
    .A(\inv_in[3150] ));
 sg13g2_inv_2 \inv[3151]/_0_  (.Y(\inv_in[3152] ),
    .A(\inv_in[3151] ));
 sg13g2_inv_2 \inv[3152]/_0_  (.Y(\inv_in[3153] ),
    .A(\inv_in[3152] ));
 sg13g2_inv_2 \inv[3153]/_0_  (.Y(\inv_in[3154] ),
    .A(\inv_in[3153] ));
 sg13g2_inv_2 \inv[3154]/_0_  (.Y(\inv_in[3155] ),
    .A(\inv_in[3154] ));
 sg13g2_inv_2 \inv[3155]/_0_  (.Y(\inv_in[3156] ),
    .A(\inv_in[3155] ));
 sg13g2_inv_2 \inv[3156]/_0_  (.Y(\inv_in[3157] ),
    .A(\inv_in[3156] ));
 sg13g2_inv_2 \inv[3157]/_0_  (.Y(\inv_in[3158] ),
    .A(\inv_in[3157] ));
 sg13g2_inv_2 \inv[3158]/_0_  (.Y(\inv_in[3159] ),
    .A(\inv_in[3158] ));
 sg13g2_inv_2 \inv[3159]/_0_  (.Y(\inv_in[3160] ),
    .A(\inv_in[3159] ));
 sg13g2_inv_2 \inv[315]/_0_  (.Y(\inv_in[316] ),
    .A(\inv_in[315] ));
 sg13g2_inv_2 \inv[3160]/_0_  (.Y(\inv_in[3161] ),
    .A(\inv_in[3160] ));
 sg13g2_inv_2 \inv[3161]/_0_  (.Y(\inv_in[3162] ),
    .A(\inv_in[3161] ));
 sg13g2_inv_2 \inv[3162]/_0_  (.Y(\inv_in[3163] ),
    .A(\inv_in[3162] ));
 sg13g2_inv_2 \inv[3163]/_0_  (.Y(\inv_in[3164] ),
    .A(\inv_in[3163] ));
 sg13g2_inv_2 \inv[3164]/_0_  (.Y(\inv_in[3165] ),
    .A(\inv_in[3164] ));
 sg13g2_inv_2 \inv[3165]/_0_  (.Y(\inv_in[3166] ),
    .A(\inv_in[3165] ));
 sg13g2_inv_2 \inv[3166]/_0_  (.Y(\inv_in[3167] ),
    .A(\inv_in[3166] ));
 sg13g2_inv_2 \inv[3167]/_0_  (.Y(\inv_in[3168] ),
    .A(\inv_in[3167] ));
 sg13g2_inv_2 \inv[3168]/_0_  (.Y(\inv_in[3169] ),
    .A(\inv_in[3168] ));
 sg13g2_inv_2 \inv[3169]/_0_  (.Y(\inv_in[3170] ),
    .A(\inv_in[3169] ));
 sg13g2_inv_2 \inv[316]/_0_  (.Y(\inv_in[317] ),
    .A(\inv_in[316] ));
 sg13g2_inv_2 \inv[3170]/_0_  (.Y(\inv_in[3171] ),
    .A(\inv_in[3170] ));
 sg13g2_inv_2 \inv[3171]/_0_  (.Y(\inv_in[3172] ),
    .A(\inv_in[3171] ));
 sg13g2_inv_2 \inv[3172]/_0_  (.Y(\inv_in[3173] ),
    .A(\inv_in[3172] ));
 sg13g2_inv_2 \inv[3173]/_0_  (.Y(\inv_in[3174] ),
    .A(\inv_in[3173] ));
 sg13g2_inv_2 \inv[3174]/_0_  (.Y(\inv_in[3175] ),
    .A(\inv_in[3174] ));
 sg13g2_inv_2 \inv[3175]/_0_  (.Y(\inv_in[3176] ),
    .A(\inv_in[3175] ));
 sg13g2_inv_2 \inv[3176]/_0_  (.Y(\inv_in[3177] ),
    .A(\inv_in[3176] ));
 sg13g2_inv_2 \inv[3177]/_0_  (.Y(\inv_in[3178] ),
    .A(\inv_in[3177] ));
 sg13g2_inv_2 \inv[3178]/_0_  (.Y(\inv_in[3179] ),
    .A(\inv_in[3178] ));
 sg13g2_inv_2 \inv[3179]/_0_  (.Y(\inv_in[3180] ),
    .A(\inv_in[3179] ));
 sg13g2_inv_2 \inv[317]/_0_  (.Y(\inv_in[318] ),
    .A(\inv_in[317] ));
 sg13g2_inv_2 \inv[3180]/_0_  (.Y(\inv_in[3181] ),
    .A(\inv_in[3180] ));
 sg13g2_inv_2 \inv[3181]/_0_  (.Y(\inv_in[3182] ),
    .A(\inv_in[3181] ));
 sg13g2_inv_2 \inv[3182]/_0_  (.Y(\inv_in[3183] ),
    .A(\inv_in[3182] ));
 sg13g2_inv_2 \inv[3183]/_0_  (.Y(\inv_in[3184] ),
    .A(\inv_in[3183] ));
 sg13g2_inv_2 \inv[3184]/_0_  (.Y(\inv_in[3185] ),
    .A(\inv_in[3184] ));
 sg13g2_inv_2 \inv[3185]/_0_  (.Y(\inv_in[3186] ),
    .A(\inv_in[3185] ));
 sg13g2_inv_2 \inv[3186]/_0_  (.Y(\inv_in[3187] ),
    .A(\inv_in[3186] ));
 sg13g2_inv_2 \inv[3187]/_0_  (.Y(\inv_in[3188] ),
    .A(\inv_in[3187] ));
 sg13g2_inv_2 \inv[3188]/_0_  (.Y(\inv_in[3189] ),
    .A(\inv_in[3188] ));
 sg13g2_inv_2 \inv[3189]/_0_  (.Y(\inv_in[3190] ),
    .A(\inv_in[3189] ));
 sg13g2_inv_2 \inv[318]/_0_  (.Y(\inv_in[319] ),
    .A(\inv_in[318] ));
 sg13g2_inv_2 \inv[3190]/_0_  (.Y(\inv_in[3191] ),
    .A(\inv_in[3190] ));
 sg13g2_inv_2 \inv[3191]/_0_  (.Y(\inv_in[3192] ),
    .A(\inv_in[3191] ));
 sg13g2_inv_2 \inv[3192]/_0_  (.Y(\inv_in[3193] ),
    .A(\inv_in[3192] ));
 sg13g2_inv_2 \inv[3193]/_0_  (.Y(\inv_in[3194] ),
    .A(\inv_in[3193] ));
 sg13g2_inv_2 \inv[3194]/_0_  (.Y(\inv_in[3195] ),
    .A(\inv_in[3194] ));
 sg13g2_inv_2 \inv[3195]/_0_  (.Y(\inv_in[3196] ),
    .A(\inv_in[3195] ));
 sg13g2_inv_2 \inv[3196]/_0_  (.Y(\inv_in[3197] ),
    .A(\inv_in[3196] ));
 sg13g2_inv_2 \inv[3197]/_0_  (.Y(\inv_in[3198] ),
    .A(\inv_in[3197] ));
 sg13g2_inv_2 \inv[3198]/_0_  (.Y(\inv_in[3199] ),
    .A(\inv_in[3198] ));
 sg13g2_inv_2 \inv[3199]/_0_  (.Y(\inv_in[3200] ),
    .A(\inv_in[3199] ));
 sg13g2_inv_2 \inv[319]/_0_  (.Y(\inv_in[320] ),
    .A(\inv_in[319] ));
 sg13g2_inv_2 \inv[31]/_0_  (.Y(\inv_in[32] ),
    .A(\inv_in[31] ));
 sg13g2_inv_2 \inv[3200]/_0_  (.Y(\inv_in[3201] ),
    .A(\inv_in[3200] ));
 sg13g2_inv_2 \inv[3201]/_0_  (.Y(\inv_in[3202] ),
    .A(\inv_in[3201] ));
 sg13g2_inv_2 \inv[3202]/_0_  (.Y(\inv_in[3203] ),
    .A(\inv_in[3202] ));
 sg13g2_inv_2 \inv[3203]/_0_  (.Y(\inv_in[3204] ),
    .A(\inv_in[3203] ));
 sg13g2_inv_2 \inv[3204]/_0_  (.Y(\inv_in[3205] ),
    .A(\inv_in[3204] ));
 sg13g2_inv_2 \inv[3205]/_0_  (.Y(\inv_in[3206] ),
    .A(\inv_in[3205] ));
 sg13g2_inv_2 \inv[3206]/_0_  (.Y(\inv_in[3207] ),
    .A(\inv_in[3206] ));
 sg13g2_inv_2 \inv[3207]/_0_  (.Y(\inv_in[3208] ),
    .A(\inv_in[3207] ));
 sg13g2_inv_2 \inv[3208]/_0_  (.Y(\inv_in[3209] ),
    .A(\inv_in[3208] ));
 sg13g2_inv_2 \inv[3209]/_0_  (.Y(\inv_in[3210] ),
    .A(\inv_in[3209] ));
 sg13g2_inv_2 \inv[320]/_0_  (.Y(\inv_in[321] ),
    .A(\inv_in[320] ));
 sg13g2_inv_2 \inv[3210]/_0_  (.Y(\inv_in[3211] ),
    .A(\inv_in[3210] ));
 sg13g2_inv_2 \inv[3211]/_0_  (.Y(\inv_in[3212] ),
    .A(\inv_in[3211] ));
 sg13g2_inv_2 \inv[3212]/_0_  (.Y(\inv_in[3213] ),
    .A(\inv_in[3212] ));
 sg13g2_inv_2 \inv[3213]/_0_  (.Y(\inv_in[3214] ),
    .A(\inv_in[3213] ));
 sg13g2_inv_2 \inv[3214]/_0_  (.Y(\inv_in[3215] ),
    .A(\inv_in[3214] ));
 sg13g2_inv_2 \inv[3215]/_0_  (.Y(\inv_in[3216] ),
    .A(\inv_in[3215] ));
 sg13g2_inv_2 \inv[3216]/_0_  (.Y(\inv_in[3217] ),
    .A(\inv_in[3216] ));
 sg13g2_inv_2 \inv[3217]/_0_  (.Y(\inv_in[3218] ),
    .A(\inv_in[3217] ));
 sg13g2_inv_2 \inv[3218]/_0_  (.Y(\inv_in[3219] ),
    .A(\inv_in[3218] ));
 sg13g2_inv_2 \inv[3219]/_0_  (.Y(\inv_in[3220] ),
    .A(\inv_in[3219] ));
 sg13g2_inv_2 \inv[321]/_0_  (.Y(\inv_in[322] ),
    .A(\inv_in[321] ));
 sg13g2_inv_2 \inv[3220]/_0_  (.Y(\inv_in[3221] ),
    .A(\inv_in[3220] ));
 sg13g2_inv_2 \inv[3221]/_0_  (.Y(\inv_in[3222] ),
    .A(\inv_in[3221] ));
 sg13g2_inv_2 \inv[3222]/_0_  (.Y(\inv_in[3223] ),
    .A(\inv_in[3222] ));
 sg13g2_inv_2 \inv[3223]/_0_  (.Y(\inv_in[3224] ),
    .A(\inv_in[3223] ));
 sg13g2_inv_2 \inv[3224]/_0_  (.Y(\inv_in[3225] ),
    .A(\inv_in[3224] ));
 sg13g2_inv_2 \inv[3225]/_0_  (.Y(\inv_in[3226] ),
    .A(\inv_in[3225] ));
 sg13g2_inv_2 \inv[3226]/_0_  (.Y(\inv_in[3227] ),
    .A(\inv_in[3226] ));
 sg13g2_inv_2 \inv[3227]/_0_  (.Y(\inv_in[3228] ),
    .A(\inv_in[3227] ));
 sg13g2_inv_2 \inv[3228]/_0_  (.Y(\inv_in[3229] ),
    .A(\inv_in[3228] ));
 sg13g2_inv_2 \inv[3229]/_0_  (.Y(\inv_in[3230] ),
    .A(\inv_in[3229] ));
 sg13g2_inv_2 \inv[322]/_0_  (.Y(\inv_in[323] ),
    .A(\inv_in[322] ));
 sg13g2_inv_2 \inv[3230]/_0_  (.Y(\inv_in[3231] ),
    .A(\inv_in[3230] ));
 sg13g2_inv_2 \inv[3231]/_0_  (.Y(\inv_in[3232] ),
    .A(\inv_in[3231] ));
 sg13g2_inv_2 \inv[3232]/_0_  (.Y(\inv_in[3233] ),
    .A(\inv_in[3232] ));
 sg13g2_inv_2 \inv[3233]/_0_  (.Y(\inv_in[3234] ),
    .A(\inv_in[3233] ));
 sg13g2_inv_2 \inv[3234]/_0_  (.Y(\inv_in[3235] ),
    .A(\inv_in[3234] ));
 sg13g2_inv_2 \inv[3235]/_0_  (.Y(\inv_in[3236] ),
    .A(\inv_in[3235] ));
 sg13g2_inv_2 \inv[3236]/_0_  (.Y(\inv_in[3237] ),
    .A(\inv_in[3236] ));
 sg13g2_inv_2 \inv[3237]/_0_  (.Y(\inv_in[3238] ),
    .A(\inv_in[3237] ));
 sg13g2_inv_2 \inv[3238]/_0_  (.Y(\inv_in[3239] ),
    .A(\inv_in[3238] ));
 sg13g2_inv_2 \inv[3239]/_0_  (.Y(\inv_in[3240] ),
    .A(\inv_in[3239] ));
 sg13g2_inv_2 \inv[323]/_0_  (.Y(\inv_in[324] ),
    .A(\inv_in[323] ));
 sg13g2_inv_2 \inv[3240]/_0_  (.Y(\inv_in[3241] ),
    .A(\inv_in[3240] ));
 sg13g2_inv_2 \inv[3241]/_0_  (.Y(\inv_in[3242] ),
    .A(\inv_in[3241] ));
 sg13g2_inv_2 \inv[3242]/_0_  (.Y(\inv_in[3243] ),
    .A(\inv_in[3242] ));
 sg13g2_inv_2 \inv[3243]/_0_  (.Y(\inv_in[3244] ),
    .A(\inv_in[3243] ));
 sg13g2_inv_2 \inv[3244]/_0_  (.Y(\inv_in[3245] ),
    .A(\inv_in[3244] ));
 sg13g2_inv_2 \inv[3245]/_0_  (.Y(\inv_in[3246] ),
    .A(\inv_in[3245] ));
 sg13g2_inv_2 \inv[3246]/_0_  (.Y(\inv_in[3247] ),
    .A(\inv_in[3246] ));
 sg13g2_inv_2 \inv[3247]/_0_  (.Y(\inv_in[3248] ),
    .A(\inv_in[3247] ));
 sg13g2_inv_2 \inv[3248]/_0_  (.Y(\inv_in[3249] ),
    .A(\inv_in[3248] ));
 sg13g2_inv_2 \inv[3249]/_0_  (.Y(\inv_in[3250] ),
    .A(\inv_in[3249] ));
 sg13g2_inv_2 \inv[324]/_0_  (.Y(\inv_in[325] ),
    .A(\inv_in[324] ));
 sg13g2_inv_2 \inv[3250]/_0_  (.Y(\inv_in[3251] ),
    .A(\inv_in[3250] ));
 sg13g2_inv_2 \inv[3251]/_0_  (.Y(\inv_in[3252] ),
    .A(\inv_in[3251] ));
 sg13g2_inv_2 \inv[3252]/_0_  (.Y(\inv_in[3253] ),
    .A(\inv_in[3252] ));
 sg13g2_inv_2 \inv[3253]/_0_  (.Y(\inv_in[3254] ),
    .A(\inv_in[3253] ));
 sg13g2_inv_2 \inv[3254]/_0_  (.Y(\inv_in[3255] ),
    .A(\inv_in[3254] ));
 sg13g2_inv_2 \inv[3255]/_0_  (.Y(\inv_in[3256] ),
    .A(\inv_in[3255] ));
 sg13g2_inv_2 \inv[3256]/_0_  (.Y(\inv_in[3257] ),
    .A(\inv_in[3256] ));
 sg13g2_inv_2 \inv[3257]/_0_  (.Y(\inv_in[3258] ),
    .A(\inv_in[3257] ));
 sg13g2_inv_2 \inv[3258]/_0_  (.Y(\inv_in[3259] ),
    .A(\inv_in[3258] ));
 sg13g2_inv_2 \inv[3259]/_0_  (.Y(\inv_in[3260] ),
    .A(\inv_in[3259] ));
 sg13g2_inv_2 \inv[325]/_0_  (.Y(\inv_in[326] ),
    .A(\inv_in[325] ));
 sg13g2_inv_2 \inv[3260]/_0_  (.Y(\inv_in[3261] ),
    .A(\inv_in[3260] ));
 sg13g2_inv_2 \inv[3261]/_0_  (.Y(\inv_in[3262] ),
    .A(\inv_in[3261] ));
 sg13g2_inv_2 \inv[3262]/_0_  (.Y(\inv_in[3263] ),
    .A(\inv_in[3262] ));
 sg13g2_inv_2 \inv[3263]/_0_  (.Y(\inv_in[3264] ),
    .A(\inv_in[3263] ));
 sg13g2_inv_2 \inv[3264]/_0_  (.Y(\inv_in[3265] ),
    .A(\inv_in[3264] ));
 sg13g2_inv_2 \inv[3265]/_0_  (.Y(\inv_in[3266] ),
    .A(\inv_in[3265] ));
 sg13g2_inv_2 \inv[3266]/_0_  (.Y(\inv_in[3267] ),
    .A(\inv_in[3266] ));
 sg13g2_inv_2 \inv[3267]/_0_  (.Y(\inv_in[3268] ),
    .A(\inv_in[3267] ));
 sg13g2_inv_2 \inv[3268]/_0_  (.Y(\inv_in[3269] ),
    .A(\inv_in[3268] ));
 sg13g2_inv_2 \inv[3269]/_0_  (.Y(\inv_in[3270] ),
    .A(\inv_in[3269] ));
 sg13g2_inv_2 \inv[326]/_0_  (.Y(\inv_in[327] ),
    .A(\inv_in[326] ));
 sg13g2_inv_2 \inv[3270]/_0_  (.Y(\inv_in[3271] ),
    .A(\inv_in[3270] ));
 sg13g2_inv_2 \inv[3271]/_0_  (.Y(\inv_in[3272] ),
    .A(\inv_in[3271] ));
 sg13g2_inv_2 \inv[3272]/_0_  (.Y(\inv_in[3273] ),
    .A(\inv_in[3272] ));
 sg13g2_inv_2 \inv[3273]/_0_  (.Y(\inv_in[3274] ),
    .A(\inv_in[3273] ));
 sg13g2_inv_2 \inv[3274]/_0_  (.Y(\inv_in[3275] ),
    .A(\inv_in[3274] ));
 sg13g2_inv_2 \inv[3275]/_0_  (.Y(\inv_in[3276] ),
    .A(\inv_in[3275] ));
 sg13g2_inv_2 \inv[3276]/_0_  (.Y(\inv_in[3277] ),
    .A(\inv_in[3276] ));
 sg13g2_inv_2 \inv[3277]/_0_  (.Y(\inv_in[3278] ),
    .A(\inv_in[3277] ));
 sg13g2_inv_2 \inv[3278]/_0_  (.Y(\inv_in[3279] ),
    .A(\inv_in[3278] ));
 sg13g2_inv_2 \inv[3279]/_0_  (.Y(\inv_in[3280] ),
    .A(\inv_in[3279] ));
 sg13g2_inv_2 \inv[327]/_0_  (.Y(\inv_in[328] ),
    .A(\inv_in[327] ));
 sg13g2_inv_2 \inv[3280]/_0_  (.Y(\inv_in[3281] ),
    .A(\inv_in[3280] ));
 sg13g2_inv_2 \inv[3281]/_0_  (.Y(\inv_in[3282] ),
    .A(\inv_in[3281] ));
 sg13g2_inv_2 \inv[3282]/_0_  (.Y(\inv_in[3283] ),
    .A(\inv_in[3282] ));
 sg13g2_inv_2 \inv[3283]/_0_  (.Y(\inv_in[3284] ),
    .A(\inv_in[3283] ));
 sg13g2_inv_2 \inv[3284]/_0_  (.Y(\inv_in[3285] ),
    .A(\inv_in[3284] ));
 sg13g2_inv_2 \inv[3285]/_0_  (.Y(\inv_in[3286] ),
    .A(\inv_in[3285] ));
 sg13g2_inv_2 \inv[3286]/_0_  (.Y(\inv_in[3287] ),
    .A(\inv_in[3286] ));
 sg13g2_inv_2 \inv[3287]/_0_  (.Y(\inv_in[3288] ),
    .A(\inv_in[3287] ));
 sg13g2_inv_2 \inv[3288]/_0_  (.Y(\inv_in[3289] ),
    .A(\inv_in[3288] ));
 sg13g2_inv_2 \inv[3289]/_0_  (.Y(\inv_in[3290] ),
    .A(\inv_in[3289] ));
 sg13g2_inv_2 \inv[328]/_0_  (.Y(\inv_in[329] ),
    .A(\inv_in[328] ));
 sg13g2_inv_2 \inv[3290]/_0_  (.Y(\inv_in[3291] ),
    .A(\inv_in[3290] ));
 sg13g2_inv_2 \inv[3291]/_0_  (.Y(\inv_in[3292] ),
    .A(\inv_in[3291] ));
 sg13g2_inv_2 \inv[3292]/_0_  (.Y(\inv_in[3293] ),
    .A(\inv_in[3292] ));
 sg13g2_inv_2 \inv[3293]/_0_  (.Y(\inv_in[3294] ),
    .A(\inv_in[3293] ));
 sg13g2_inv_2 \inv[3294]/_0_  (.Y(\inv_in[3295] ),
    .A(\inv_in[3294] ));
 sg13g2_inv_2 \inv[3295]/_0_  (.Y(\inv_in[3296] ),
    .A(\inv_in[3295] ));
 sg13g2_inv_2 \inv[3296]/_0_  (.Y(\inv_in[3297] ),
    .A(\inv_in[3296] ));
 sg13g2_inv_2 \inv[3297]/_0_  (.Y(\inv_in[3298] ),
    .A(\inv_in[3297] ));
 sg13g2_inv_2 \inv[3298]/_0_  (.Y(\inv_in[3299] ),
    .A(\inv_in[3298] ));
 sg13g2_inv_2 \inv[3299]/_0_  (.Y(\inv_in[3300] ),
    .A(\inv_in[3299] ));
 sg13g2_inv_2 \inv[329]/_0_  (.Y(\inv_in[330] ),
    .A(\inv_in[329] ));
 sg13g2_inv_2 \inv[32]/_0_  (.Y(\inv_in[33] ),
    .A(\inv_in[32] ));
 sg13g2_inv_2 \inv[3300]/_0_  (.Y(\inv_in[3301] ),
    .A(\inv_in[3300] ));
 sg13g2_inv_2 \inv[3301]/_0_  (.Y(\inv_in[3302] ),
    .A(\inv_in[3301] ));
 sg13g2_inv_2 \inv[3302]/_0_  (.Y(\inv_in[3303] ),
    .A(\inv_in[3302] ));
 sg13g2_inv_2 \inv[3303]/_0_  (.Y(\inv_in[3304] ),
    .A(\inv_in[3303] ));
 sg13g2_inv_2 \inv[3304]/_0_  (.Y(\inv_in[3305] ),
    .A(\inv_in[3304] ));
 sg13g2_inv_2 \inv[3305]/_0_  (.Y(\inv_in[3306] ),
    .A(\inv_in[3305] ));
 sg13g2_inv_2 \inv[3306]/_0_  (.Y(\inv_in[3307] ),
    .A(\inv_in[3306] ));
 sg13g2_inv_2 \inv[3307]/_0_  (.Y(\inv_in[3308] ),
    .A(\inv_in[3307] ));
 sg13g2_inv_2 \inv[3308]/_0_  (.Y(\inv_in[3309] ),
    .A(\inv_in[3308] ));
 sg13g2_inv_2 \inv[3309]/_0_  (.Y(\inv_in[3310] ),
    .A(\inv_in[3309] ));
 sg13g2_inv_2 \inv[330]/_0_  (.Y(\inv_in[331] ),
    .A(\inv_in[330] ));
 sg13g2_inv_2 \inv[3310]/_0_  (.Y(\inv_in[3311] ),
    .A(\inv_in[3310] ));
 sg13g2_inv_2 \inv[3311]/_0_  (.Y(\inv_in[3312] ),
    .A(\inv_in[3311] ));
 sg13g2_inv_2 \inv[3312]/_0_  (.Y(\inv_in[3313] ),
    .A(\inv_in[3312] ));
 sg13g2_inv_2 \inv[3313]/_0_  (.Y(\inv_in[3314] ),
    .A(\inv_in[3313] ));
 sg13g2_inv_2 \inv[3314]/_0_  (.Y(\inv_in[3315] ),
    .A(\inv_in[3314] ));
 sg13g2_inv_2 \inv[3315]/_0_  (.Y(\inv_in[3316] ),
    .A(\inv_in[3315] ));
 sg13g2_inv_2 \inv[3316]/_0_  (.Y(\inv_in[3317] ),
    .A(\inv_in[3316] ));
 sg13g2_inv_2 \inv[3317]/_0_  (.Y(\inv_in[3318] ),
    .A(\inv_in[3317] ));
 sg13g2_inv_2 \inv[3318]/_0_  (.Y(\inv_in[3319] ),
    .A(\inv_in[3318] ));
 sg13g2_inv_2 \inv[3319]/_0_  (.Y(\inv_in[3320] ),
    .A(\inv_in[3319] ));
 sg13g2_inv_2 \inv[331]/_0_  (.Y(\inv_in[332] ),
    .A(\inv_in[331] ));
 sg13g2_inv_2 \inv[3320]/_0_  (.Y(\inv_in[3321] ),
    .A(\inv_in[3320] ));
 sg13g2_inv_2 \inv[3321]/_0_  (.Y(\inv_in[3322] ),
    .A(\inv_in[3321] ));
 sg13g2_inv_2 \inv[3322]/_0_  (.Y(\inv_in[3323] ),
    .A(\inv_in[3322] ));
 sg13g2_inv_2 \inv[3323]/_0_  (.Y(\inv_in[3324] ),
    .A(\inv_in[3323] ));
 sg13g2_inv_2 \inv[3324]/_0_  (.Y(\inv_in[3325] ),
    .A(\inv_in[3324] ));
 sg13g2_inv_2 \inv[3325]/_0_  (.Y(\inv_in[3326] ),
    .A(\inv_in[3325] ));
 sg13g2_inv_2 \inv[3326]/_0_  (.Y(\inv_in[3327] ),
    .A(\inv_in[3326] ));
 sg13g2_inv_2 \inv[3327]/_0_  (.Y(\inv_in[3328] ),
    .A(\inv_in[3327] ));
 sg13g2_inv_2 \inv[3328]/_0_  (.Y(\inv_in[3329] ),
    .A(\inv_in[3328] ));
 sg13g2_inv_2 \inv[3329]/_0_  (.Y(\inv_in[3330] ),
    .A(\inv_in[3329] ));
 sg13g2_inv_2 \inv[332]/_0_  (.Y(\inv_in[333] ),
    .A(\inv_in[332] ));
 sg13g2_inv_2 \inv[3330]/_0_  (.Y(\inv_in[3331] ),
    .A(\inv_in[3330] ));
 sg13g2_inv_2 \inv[3331]/_0_  (.Y(\inv_in[3332] ),
    .A(\inv_in[3331] ));
 sg13g2_inv_2 \inv[3332]/_0_  (.Y(\inv_in[3333] ),
    .A(\inv_in[3332] ));
 sg13g2_inv_2 \inv[3333]/_0_  (.Y(\inv_in[3334] ),
    .A(\inv_in[3333] ));
 sg13g2_inv_2 \inv[3334]/_0_  (.Y(\inv_in[3335] ),
    .A(\inv_in[3334] ));
 sg13g2_inv_2 \inv[3335]/_0_  (.Y(\inv_in[3336] ),
    .A(\inv_in[3335] ));
 sg13g2_inv_2 \inv[3336]/_0_  (.Y(\inv_in[3337] ),
    .A(\inv_in[3336] ));
 sg13g2_inv_2 \inv[3337]/_0_  (.Y(\inv_in[3338] ),
    .A(\inv_in[3337] ));
 sg13g2_inv_2 \inv[3338]/_0_  (.Y(\inv_in[3339] ),
    .A(\inv_in[3338] ));
 sg13g2_inv_2 \inv[3339]/_0_  (.Y(\inv_in[3340] ),
    .A(\inv_in[3339] ));
 sg13g2_inv_2 \inv[333]/_0_  (.Y(\inv_in[334] ),
    .A(\inv_in[333] ));
 sg13g2_inv_2 \inv[3340]/_0_  (.Y(\inv_in[3341] ),
    .A(\inv_in[3340] ));
 sg13g2_inv_2 \inv[3341]/_0_  (.Y(\inv_in[3342] ),
    .A(\inv_in[3341] ));
 sg13g2_inv_2 \inv[3342]/_0_  (.Y(\inv_in[3343] ),
    .A(\inv_in[3342] ));
 sg13g2_inv_2 \inv[3343]/_0_  (.Y(\inv_in[3344] ),
    .A(\inv_in[3343] ));
 sg13g2_inv_2 \inv[3344]/_0_  (.Y(\inv_in[3345] ),
    .A(\inv_in[3344] ));
 sg13g2_inv_2 \inv[3345]/_0_  (.Y(\inv_in[3346] ),
    .A(\inv_in[3345] ));
 sg13g2_inv_2 \inv[3346]/_0_  (.Y(\inv_in[3347] ),
    .A(\inv_in[3346] ));
 sg13g2_inv_2 \inv[3347]/_0_  (.Y(\inv_in[3348] ),
    .A(\inv_in[3347] ));
 sg13g2_inv_2 \inv[3348]/_0_  (.Y(\inv_in[3349] ),
    .A(\inv_in[3348] ));
 sg13g2_inv_2 \inv[3349]/_0_  (.Y(\inv_in[3350] ),
    .A(\inv_in[3349] ));
 sg13g2_inv_2 \inv[334]/_0_  (.Y(\inv_in[335] ),
    .A(\inv_in[334] ));
 sg13g2_inv_2 \inv[3350]/_0_  (.Y(\inv_in[3351] ),
    .A(\inv_in[3350] ));
 sg13g2_inv_2 \inv[3351]/_0_  (.Y(\inv_in[3352] ),
    .A(\inv_in[3351] ));
 sg13g2_inv_2 \inv[3352]/_0_  (.Y(\inv_in[3353] ),
    .A(\inv_in[3352] ));
 sg13g2_inv_2 \inv[3353]/_0_  (.Y(\inv_in[3354] ),
    .A(\inv_in[3353] ));
 sg13g2_inv_2 \inv[3354]/_0_  (.Y(\inv_in[3355] ),
    .A(\inv_in[3354] ));
 sg13g2_inv_2 \inv[3355]/_0_  (.Y(\inv_in[3356] ),
    .A(\inv_in[3355] ));
 sg13g2_inv_2 \inv[3356]/_0_  (.Y(\inv_in[3357] ),
    .A(\inv_in[3356] ));
 sg13g2_inv_2 \inv[3357]/_0_  (.Y(\inv_in[3358] ),
    .A(\inv_in[3357] ));
 sg13g2_inv_2 \inv[3358]/_0_  (.Y(\inv_in[3359] ),
    .A(\inv_in[3358] ));
 sg13g2_inv_2 \inv[3359]/_0_  (.Y(\inv_in[3360] ),
    .A(\inv_in[3359] ));
 sg13g2_inv_2 \inv[335]/_0_  (.Y(\inv_in[336] ),
    .A(\inv_in[335] ));
 sg13g2_inv_2 \inv[3360]/_0_  (.Y(\inv_in[3361] ),
    .A(\inv_in[3360] ));
 sg13g2_inv_2 \inv[3361]/_0_  (.Y(\inv_in[3362] ),
    .A(\inv_in[3361] ));
 sg13g2_inv_2 \inv[3362]/_0_  (.Y(\inv_in[3363] ),
    .A(\inv_in[3362] ));
 sg13g2_inv_2 \inv[3363]/_0_  (.Y(\inv_in[3364] ),
    .A(\inv_in[3363] ));
 sg13g2_inv_2 \inv[3364]/_0_  (.Y(\inv_in[3365] ),
    .A(\inv_in[3364] ));
 sg13g2_inv_2 \inv[3365]/_0_  (.Y(\inv_in[3366] ),
    .A(\inv_in[3365] ));
 sg13g2_inv_2 \inv[3366]/_0_  (.Y(\inv_in[3367] ),
    .A(\inv_in[3366] ));
 sg13g2_inv_2 \inv[3367]/_0_  (.Y(\inv_in[3368] ),
    .A(\inv_in[3367] ));
 sg13g2_inv_2 \inv[3368]/_0_  (.Y(\inv_in[3369] ),
    .A(\inv_in[3368] ));
 sg13g2_inv_2 \inv[3369]/_0_  (.Y(\inv_in[3370] ),
    .A(\inv_in[3369] ));
 sg13g2_inv_2 \inv[336]/_0_  (.Y(\inv_in[337] ),
    .A(\inv_in[336] ));
 sg13g2_inv_2 \inv[3370]/_0_  (.Y(\inv_in[3371] ),
    .A(\inv_in[3370] ));
 sg13g2_inv_2 \inv[3371]/_0_  (.Y(\inv_in[3372] ),
    .A(\inv_in[3371] ));
 sg13g2_inv_2 \inv[3372]/_0_  (.Y(\inv_in[3373] ),
    .A(\inv_in[3372] ));
 sg13g2_inv_2 \inv[3373]/_0_  (.Y(\inv_in[3374] ),
    .A(\inv_in[3373] ));
 sg13g2_inv_2 \inv[3374]/_0_  (.Y(\inv_in[3375] ),
    .A(\inv_in[3374] ));
 sg13g2_inv_2 \inv[3375]/_0_  (.Y(\inv_in[3376] ),
    .A(\inv_in[3375] ));
 sg13g2_inv_2 \inv[3376]/_0_  (.Y(\inv_in[3377] ),
    .A(\inv_in[3376] ));
 sg13g2_inv_2 \inv[3377]/_0_  (.Y(\inv_in[3378] ),
    .A(\inv_in[3377] ));
 sg13g2_inv_2 \inv[3378]/_0_  (.Y(\inv_in[3379] ),
    .A(\inv_in[3378] ));
 sg13g2_inv_2 \inv[3379]/_0_  (.Y(\inv_in[3380] ),
    .A(\inv_in[3379] ));
 sg13g2_inv_2 \inv[337]/_0_  (.Y(\inv_in[338] ),
    .A(\inv_in[337] ));
 sg13g2_inv_2 \inv[3380]/_0_  (.Y(\inv_in[3381] ),
    .A(\inv_in[3380] ));
 sg13g2_inv_2 \inv[3381]/_0_  (.Y(\inv_in[3382] ),
    .A(\inv_in[3381] ));
 sg13g2_inv_2 \inv[3382]/_0_  (.Y(\inv_in[3383] ),
    .A(\inv_in[3382] ));
 sg13g2_inv_2 \inv[3383]/_0_  (.Y(\inv_in[3384] ),
    .A(\inv_in[3383] ));
 sg13g2_inv_2 \inv[3384]/_0_  (.Y(\inv_in[3385] ),
    .A(\inv_in[3384] ));
 sg13g2_inv_2 \inv[3385]/_0_  (.Y(\inv_in[3386] ),
    .A(\inv_in[3385] ));
 sg13g2_inv_2 \inv[3386]/_0_  (.Y(\inv_in[3387] ),
    .A(\inv_in[3386] ));
 sg13g2_inv_2 \inv[3387]/_0_  (.Y(\inv_in[3388] ),
    .A(\inv_in[3387] ));
 sg13g2_inv_2 \inv[3388]/_0_  (.Y(\inv_in[3389] ),
    .A(\inv_in[3388] ));
 sg13g2_inv_2 \inv[3389]/_0_  (.Y(\inv_in[3390] ),
    .A(\inv_in[3389] ));
 sg13g2_inv_2 \inv[338]/_0_  (.Y(\inv_in[339] ),
    .A(\inv_in[338] ));
 sg13g2_inv_2 \inv[3390]/_0_  (.Y(\inv_in[3391] ),
    .A(\inv_in[3390] ));
 sg13g2_inv_2 \inv[3391]/_0_  (.Y(\inv_in[3392] ),
    .A(\inv_in[3391] ));
 sg13g2_inv_2 \inv[3392]/_0_  (.Y(\inv_in[3393] ),
    .A(\inv_in[3392] ));
 sg13g2_inv_2 \inv[3393]/_0_  (.Y(\inv_in[3394] ),
    .A(\inv_in[3393] ));
 sg13g2_inv_2 \inv[3394]/_0_  (.Y(\inv_in[3395] ),
    .A(\inv_in[3394] ));
 sg13g2_inv_2 \inv[3395]/_0_  (.Y(\inv_in[3396] ),
    .A(\inv_in[3395] ));
 sg13g2_inv_2 \inv[3396]/_0_  (.Y(\inv_in[3397] ),
    .A(\inv_in[3396] ));
 sg13g2_inv_2 \inv[3397]/_0_  (.Y(\inv_in[3398] ),
    .A(\inv_in[3397] ));
 sg13g2_inv_2 \inv[3398]/_0_  (.Y(\inv_in[3399] ),
    .A(\inv_in[3398] ));
 sg13g2_inv_2 \inv[3399]/_0_  (.Y(\inv_in[3400] ),
    .A(\inv_in[3399] ));
 sg13g2_inv_2 \inv[339]/_0_  (.Y(\inv_in[340] ),
    .A(\inv_in[339] ));
 sg13g2_inv_2 \inv[33]/_0_  (.Y(\inv_in[34] ),
    .A(\inv_in[33] ));
 sg13g2_inv_2 \inv[3400]/_0_  (.Y(\inv_in[3401] ),
    .A(\inv_in[3400] ));
 sg13g2_inv_2 \inv[3401]/_0_  (.Y(\inv_in[3402] ),
    .A(\inv_in[3401] ));
 sg13g2_inv_2 \inv[3402]/_0_  (.Y(\inv_in[3403] ),
    .A(\inv_in[3402] ));
 sg13g2_inv_2 \inv[3403]/_0_  (.Y(\inv_in[3404] ),
    .A(\inv_in[3403] ));
 sg13g2_inv_2 \inv[3404]/_0_  (.Y(\inv_in[3405] ),
    .A(\inv_in[3404] ));
 sg13g2_inv_2 \inv[3405]/_0_  (.Y(\inv_in[3406] ),
    .A(\inv_in[3405] ));
 sg13g2_inv_2 \inv[3406]/_0_  (.Y(\inv_in[3407] ),
    .A(\inv_in[3406] ));
 sg13g2_inv_2 \inv[3407]/_0_  (.Y(\inv_in[3408] ),
    .A(\inv_in[3407] ));
 sg13g2_inv_2 \inv[3408]/_0_  (.Y(\inv_in[3409] ),
    .A(\inv_in[3408] ));
 sg13g2_inv_2 \inv[3409]/_0_  (.Y(\inv_in[3410] ),
    .A(\inv_in[3409] ));
 sg13g2_inv_2 \inv[340]/_0_  (.Y(\inv_in[341] ),
    .A(\inv_in[340] ));
 sg13g2_inv_2 \inv[3410]/_0_  (.Y(\inv_in[3411] ),
    .A(\inv_in[3410] ));
 sg13g2_inv_2 \inv[3411]/_0_  (.Y(\inv_in[3412] ),
    .A(\inv_in[3411] ));
 sg13g2_inv_2 \inv[3412]/_0_  (.Y(\inv_in[3413] ),
    .A(\inv_in[3412] ));
 sg13g2_inv_2 \inv[3413]/_0_  (.Y(\inv_in[3414] ),
    .A(\inv_in[3413] ));
 sg13g2_inv_2 \inv[3414]/_0_  (.Y(\inv_in[3415] ),
    .A(\inv_in[3414] ));
 sg13g2_inv_2 \inv[3415]/_0_  (.Y(\inv_in[3416] ),
    .A(\inv_in[3415] ));
 sg13g2_inv_2 \inv[3416]/_0_  (.Y(\inv_in[3417] ),
    .A(\inv_in[3416] ));
 sg13g2_inv_2 \inv[3417]/_0_  (.Y(\inv_in[3418] ),
    .A(\inv_in[3417] ));
 sg13g2_inv_2 \inv[3418]/_0_  (.Y(\inv_in[3419] ),
    .A(\inv_in[3418] ));
 sg13g2_inv_2 \inv[3419]/_0_  (.Y(\inv_in[3420] ),
    .A(\inv_in[3419] ));
 sg13g2_inv_2 \inv[341]/_0_  (.Y(\inv_in[342] ),
    .A(\inv_in[341] ));
 sg13g2_inv_2 \inv[3420]/_0_  (.Y(\inv_in[3421] ),
    .A(\inv_in[3420] ));
 sg13g2_inv_2 \inv[3421]/_0_  (.Y(\inv_in[3422] ),
    .A(\inv_in[3421] ));
 sg13g2_inv_2 \inv[3422]/_0_  (.Y(\inv_in[3423] ),
    .A(\inv_in[3422] ));
 sg13g2_inv_2 \inv[3423]/_0_  (.Y(\inv_in[3424] ),
    .A(\inv_in[3423] ));
 sg13g2_inv_2 \inv[3424]/_0_  (.Y(\inv_in[3425] ),
    .A(\inv_in[3424] ));
 sg13g2_inv_2 \inv[3425]/_0_  (.Y(\inv_in[3426] ),
    .A(\inv_in[3425] ));
 sg13g2_inv_2 \inv[3426]/_0_  (.Y(\inv_in[3427] ),
    .A(\inv_in[3426] ));
 sg13g2_inv_2 \inv[3427]/_0_  (.Y(\inv_in[3428] ),
    .A(\inv_in[3427] ));
 sg13g2_inv_2 \inv[3428]/_0_  (.Y(\inv_in[3429] ),
    .A(\inv_in[3428] ));
 sg13g2_inv_2 \inv[3429]/_0_  (.Y(\inv_in[3430] ),
    .A(\inv_in[3429] ));
 sg13g2_inv_2 \inv[342]/_0_  (.Y(\inv_in[343] ),
    .A(\inv_in[342] ));
 sg13g2_inv_2 \inv[3430]/_0_  (.Y(\inv_in[3431] ),
    .A(\inv_in[3430] ));
 sg13g2_inv_2 \inv[3431]/_0_  (.Y(\inv_in[3432] ),
    .A(\inv_in[3431] ));
 sg13g2_inv_2 \inv[3432]/_0_  (.Y(\inv_in[3433] ),
    .A(\inv_in[3432] ));
 sg13g2_inv_2 \inv[3433]/_0_  (.Y(\inv_in[3434] ),
    .A(\inv_in[3433] ));
 sg13g2_inv_2 \inv[3434]/_0_  (.Y(\inv_in[3435] ),
    .A(\inv_in[3434] ));
 sg13g2_inv_2 \inv[3435]/_0_  (.Y(\inv_in[3436] ),
    .A(\inv_in[3435] ));
 sg13g2_inv_2 \inv[3436]/_0_  (.Y(\inv_in[3437] ),
    .A(\inv_in[3436] ));
 sg13g2_inv_2 \inv[3437]/_0_  (.Y(\inv_in[3438] ),
    .A(\inv_in[3437] ));
 sg13g2_inv_2 \inv[3438]/_0_  (.Y(\inv_in[3439] ),
    .A(\inv_in[3438] ));
 sg13g2_inv_2 \inv[3439]/_0_  (.Y(\inv_in[3440] ),
    .A(\inv_in[3439] ));
 sg13g2_inv_2 \inv[343]/_0_  (.Y(\inv_in[344] ),
    .A(\inv_in[343] ));
 sg13g2_inv_2 \inv[3440]/_0_  (.Y(\inv_in[3441] ),
    .A(\inv_in[3440] ));
 sg13g2_inv_2 \inv[3441]/_0_  (.Y(\inv_in[3442] ),
    .A(\inv_in[3441] ));
 sg13g2_inv_2 \inv[3442]/_0_  (.Y(\inv_in[3443] ),
    .A(\inv_in[3442] ));
 sg13g2_inv_2 \inv[3443]/_0_  (.Y(\inv_in[3444] ),
    .A(\inv_in[3443] ));
 sg13g2_inv_2 \inv[3444]/_0_  (.Y(\inv_in[3445] ),
    .A(\inv_in[3444] ));
 sg13g2_inv_2 \inv[3445]/_0_  (.Y(\inv_in[3446] ),
    .A(\inv_in[3445] ));
 sg13g2_inv_2 \inv[3446]/_0_  (.Y(\inv_in[3447] ),
    .A(\inv_in[3446] ));
 sg13g2_inv_2 \inv[3447]/_0_  (.Y(\inv_in[3448] ),
    .A(\inv_in[3447] ));
 sg13g2_inv_2 \inv[3448]/_0_  (.Y(\inv_in[3449] ),
    .A(\inv_in[3448] ));
 sg13g2_inv_2 \inv[3449]/_0_  (.Y(\inv_in[3450] ),
    .A(\inv_in[3449] ));
 sg13g2_inv_2 \inv[344]/_0_  (.Y(\inv_in[345] ),
    .A(\inv_in[344] ));
 sg13g2_inv_2 \inv[3450]/_0_  (.Y(\inv_in[3451] ),
    .A(\inv_in[3450] ));
 sg13g2_inv_2 \inv[3451]/_0_  (.Y(\inv_in[3452] ),
    .A(\inv_in[3451] ));
 sg13g2_inv_2 \inv[3452]/_0_  (.Y(\inv_in[3453] ),
    .A(\inv_in[3452] ));
 sg13g2_inv_2 \inv[3453]/_0_  (.Y(\inv_in[3454] ),
    .A(\inv_in[3453] ));
 sg13g2_inv_2 \inv[3454]/_0_  (.Y(\inv_in[3455] ),
    .A(\inv_in[3454] ));
 sg13g2_inv_2 \inv[3455]/_0_  (.Y(\inv_in[3456] ),
    .A(\inv_in[3455] ));
 sg13g2_inv_2 \inv[3456]/_0_  (.Y(\inv_in[3457] ),
    .A(\inv_in[3456] ));
 sg13g2_inv_2 \inv[3457]/_0_  (.Y(\inv_in[3458] ),
    .A(\inv_in[3457] ));
 sg13g2_inv_2 \inv[3458]/_0_  (.Y(\inv_in[3459] ),
    .A(\inv_in[3458] ));
 sg13g2_inv_2 \inv[3459]/_0_  (.Y(\inv_in[3460] ),
    .A(\inv_in[3459] ));
 sg13g2_inv_2 \inv[345]/_0_  (.Y(\inv_in[346] ),
    .A(\inv_in[345] ));
 sg13g2_inv_2 \inv[3460]/_0_  (.Y(\inv_in[3461] ),
    .A(\inv_in[3460] ));
 sg13g2_inv_2 \inv[3461]/_0_  (.Y(\inv_in[3462] ),
    .A(\inv_in[3461] ));
 sg13g2_inv_2 \inv[3462]/_0_  (.Y(\inv_in[3463] ),
    .A(\inv_in[3462] ));
 sg13g2_inv_2 \inv[3463]/_0_  (.Y(\inv_in[3464] ),
    .A(\inv_in[3463] ));
 sg13g2_inv_2 \inv[3464]/_0_  (.Y(\inv_in[3465] ),
    .A(\inv_in[3464] ));
 sg13g2_inv_2 \inv[3465]/_0_  (.Y(\inv_in[3466] ),
    .A(\inv_in[3465] ));
 sg13g2_inv_2 \inv[3466]/_0_  (.Y(\inv_in[3467] ),
    .A(\inv_in[3466] ));
 sg13g2_inv_2 \inv[3467]/_0_  (.Y(\inv_in[3468] ),
    .A(\inv_in[3467] ));
 sg13g2_inv_2 \inv[3468]/_0_  (.Y(\inv_in[3469] ),
    .A(\inv_in[3468] ));
 sg13g2_inv_2 \inv[3469]/_0_  (.Y(\inv_in[3470] ),
    .A(\inv_in[3469] ));
 sg13g2_inv_2 \inv[346]/_0_  (.Y(\inv_in[347] ),
    .A(\inv_in[346] ));
 sg13g2_inv_2 \inv[3470]/_0_  (.Y(\inv_in[3471] ),
    .A(\inv_in[3470] ));
 sg13g2_inv_2 \inv[3471]/_0_  (.Y(\inv_in[3472] ),
    .A(\inv_in[3471] ));
 sg13g2_inv_2 \inv[3472]/_0_  (.Y(\inv_in[3473] ),
    .A(\inv_in[3472] ));
 sg13g2_inv_2 \inv[3473]/_0_  (.Y(\inv_in[3474] ),
    .A(\inv_in[3473] ));
 sg13g2_inv_2 \inv[3474]/_0_  (.Y(\inv_in[3475] ),
    .A(\inv_in[3474] ));
 sg13g2_inv_2 \inv[3475]/_0_  (.Y(\inv_in[3476] ),
    .A(\inv_in[3475] ));
 sg13g2_inv_2 \inv[3476]/_0_  (.Y(\inv_in[3477] ),
    .A(\inv_in[3476] ));
 sg13g2_inv_2 \inv[3477]/_0_  (.Y(\inv_in[3478] ),
    .A(\inv_in[3477] ));
 sg13g2_inv_2 \inv[3478]/_0_  (.Y(\inv_in[3479] ),
    .A(\inv_in[3478] ));
 sg13g2_inv_2 \inv[3479]/_0_  (.Y(\inv_in[3480] ),
    .A(\inv_in[3479] ));
 sg13g2_inv_2 \inv[347]/_0_  (.Y(\inv_in[348] ),
    .A(\inv_in[347] ));
 sg13g2_inv_2 \inv[3480]/_0_  (.Y(\inv_in[3481] ),
    .A(\inv_in[3480] ));
 sg13g2_inv_2 \inv[3481]/_0_  (.Y(\inv_in[3482] ),
    .A(\inv_in[3481] ));
 sg13g2_inv_2 \inv[3482]/_0_  (.Y(\inv_in[3483] ),
    .A(\inv_in[3482] ));
 sg13g2_inv_2 \inv[3483]/_0_  (.Y(\inv_in[3484] ),
    .A(\inv_in[3483] ));
 sg13g2_inv_2 \inv[3484]/_0_  (.Y(\inv_in[3485] ),
    .A(\inv_in[3484] ));
 sg13g2_inv_2 \inv[3485]/_0_  (.Y(\inv_in[3486] ),
    .A(\inv_in[3485] ));
 sg13g2_inv_2 \inv[3486]/_0_  (.Y(\inv_in[3487] ),
    .A(\inv_in[3486] ));
 sg13g2_inv_2 \inv[3487]/_0_  (.Y(\inv_in[3488] ),
    .A(\inv_in[3487] ));
 sg13g2_inv_2 \inv[3488]/_0_  (.Y(\inv_in[3489] ),
    .A(\inv_in[3488] ));
 sg13g2_inv_2 \inv[3489]/_0_  (.Y(\inv_in[3490] ),
    .A(\inv_in[3489] ));
 sg13g2_inv_2 \inv[348]/_0_  (.Y(\inv_in[349] ),
    .A(\inv_in[348] ));
 sg13g2_inv_2 \inv[3490]/_0_  (.Y(\inv_in[3491] ),
    .A(\inv_in[3490] ));
 sg13g2_inv_2 \inv[3491]/_0_  (.Y(\inv_in[3492] ),
    .A(\inv_in[3491] ));
 sg13g2_inv_2 \inv[3492]/_0_  (.Y(\inv_in[3493] ),
    .A(\inv_in[3492] ));
 sg13g2_inv_2 \inv[3493]/_0_  (.Y(\inv_in[3494] ),
    .A(\inv_in[3493] ));
 sg13g2_inv_2 \inv[3494]/_0_  (.Y(\inv_in[3495] ),
    .A(\inv_in[3494] ));
 sg13g2_inv_2 \inv[3495]/_0_  (.Y(\inv_in[3496] ),
    .A(\inv_in[3495] ));
 sg13g2_inv_2 \inv[3496]/_0_  (.Y(\inv_in[3497] ),
    .A(\inv_in[3496] ));
 sg13g2_inv_2 \inv[3497]/_0_  (.Y(\inv_in[3498] ),
    .A(\inv_in[3497] ));
 sg13g2_inv_2 \inv[3498]/_0_  (.Y(\inv_in[3499] ),
    .A(\inv_in[3498] ));
 sg13g2_inv_2 \inv[3499]/_0_  (.Y(\inv_in[3500] ),
    .A(\inv_in[3499] ));
 sg13g2_inv_2 \inv[349]/_0_  (.Y(\inv_in[350] ),
    .A(\inv_in[349] ));
 sg13g2_inv_2 \inv[34]/_0_  (.Y(\inv_in[35] ),
    .A(\inv_in[34] ));
 sg13g2_inv_2 \inv[3500]/_0_  (.Y(\inv_in[3501] ),
    .A(\inv_in[3500] ));
 sg13g2_inv_2 \inv[3501]/_0_  (.Y(\inv_in[3502] ),
    .A(\inv_in[3501] ));
 sg13g2_inv_2 \inv[3502]/_0_  (.Y(\inv_in[3503] ),
    .A(\inv_in[3502] ));
 sg13g2_inv_2 \inv[3503]/_0_  (.Y(\inv_in[3504] ),
    .A(\inv_in[3503] ));
 sg13g2_inv_2 \inv[3504]/_0_  (.Y(\inv_in[3505] ),
    .A(\inv_in[3504] ));
 sg13g2_inv_2 \inv[3505]/_0_  (.Y(\inv_in[3506] ),
    .A(\inv_in[3505] ));
 sg13g2_inv_2 \inv[3506]/_0_  (.Y(\inv_in[3507] ),
    .A(\inv_in[3506] ));
 sg13g2_inv_2 \inv[3507]/_0_  (.Y(\inv_in[3508] ),
    .A(\inv_in[3507] ));
 sg13g2_inv_2 \inv[3508]/_0_  (.Y(\inv_in[3509] ),
    .A(\inv_in[3508] ));
 sg13g2_inv_2 \inv[3509]/_0_  (.Y(\inv_in[3510] ),
    .A(\inv_in[3509] ));
 sg13g2_inv_2 \inv[350]/_0_  (.Y(\inv_in[351] ),
    .A(\inv_in[350] ));
 sg13g2_inv_2 \inv[3510]/_0_  (.Y(\inv_in[3511] ),
    .A(\inv_in[3510] ));
 sg13g2_inv_2 \inv[3511]/_0_  (.Y(\inv_in[3512] ),
    .A(\inv_in[3511] ));
 sg13g2_inv_2 \inv[3512]/_0_  (.Y(\inv_in[3513] ),
    .A(\inv_in[3512] ));
 sg13g2_inv_2 \inv[3513]/_0_  (.Y(\inv_in[3514] ),
    .A(\inv_in[3513] ));
 sg13g2_inv_2 \inv[3514]/_0_  (.Y(\inv_in[3515] ),
    .A(\inv_in[3514] ));
 sg13g2_inv_2 \inv[3515]/_0_  (.Y(\inv_in[3516] ),
    .A(\inv_in[3515] ));
 sg13g2_inv_2 \inv[3516]/_0_  (.Y(\inv_in[3517] ),
    .A(\inv_in[3516] ));
 sg13g2_inv_2 \inv[3517]/_0_  (.Y(\inv_in[3518] ),
    .A(\inv_in[3517] ));
 sg13g2_inv_2 \inv[3518]/_0_  (.Y(\inv_in[3519] ),
    .A(\inv_in[3518] ));
 sg13g2_inv_2 \inv[3519]/_0_  (.Y(\inv_in[3520] ),
    .A(\inv_in[3519] ));
 sg13g2_inv_2 \inv[351]/_0_  (.Y(\inv_in[352] ),
    .A(\inv_in[351] ));
 sg13g2_inv_2 \inv[3520]/_0_  (.Y(\inv_in[3521] ),
    .A(\inv_in[3520] ));
 sg13g2_inv_2 \inv[3521]/_0_  (.Y(\inv_in[3522] ),
    .A(\inv_in[3521] ));
 sg13g2_inv_2 \inv[3522]/_0_  (.Y(\inv_in[3523] ),
    .A(\inv_in[3522] ));
 sg13g2_inv_2 \inv[3523]/_0_  (.Y(\inv_in[3524] ),
    .A(\inv_in[3523] ));
 sg13g2_inv_2 \inv[3524]/_0_  (.Y(\inv_in[3525] ),
    .A(\inv_in[3524] ));
 sg13g2_inv_2 \inv[3525]/_0_  (.Y(\inv_in[3526] ),
    .A(\inv_in[3525] ));
 sg13g2_inv_2 \inv[3526]/_0_  (.Y(\inv_in[3527] ),
    .A(\inv_in[3526] ));
 sg13g2_inv_2 \inv[3527]/_0_  (.Y(\inv_in[3528] ),
    .A(\inv_in[3527] ));
 sg13g2_inv_2 \inv[3528]/_0_  (.Y(\inv_in[3529] ),
    .A(\inv_in[3528] ));
 sg13g2_inv_2 \inv[3529]/_0_  (.Y(\inv_in[3530] ),
    .A(\inv_in[3529] ));
 sg13g2_inv_2 \inv[352]/_0_  (.Y(\inv_in[353] ),
    .A(\inv_in[352] ));
 sg13g2_inv_2 \inv[3530]/_0_  (.Y(\inv_in[3531] ),
    .A(\inv_in[3530] ));
 sg13g2_inv_2 \inv[3531]/_0_  (.Y(\inv_in[3532] ),
    .A(\inv_in[3531] ));
 sg13g2_inv_2 \inv[3532]/_0_  (.Y(\inv_in[3533] ),
    .A(\inv_in[3532] ));
 sg13g2_inv_2 \inv[3533]/_0_  (.Y(\inv_in[3534] ),
    .A(\inv_in[3533] ));
 sg13g2_inv_2 \inv[3534]/_0_  (.Y(\inv_in[3535] ),
    .A(\inv_in[3534] ));
 sg13g2_inv_2 \inv[3535]/_0_  (.Y(\inv_in[3536] ),
    .A(\inv_in[3535] ));
 sg13g2_inv_2 \inv[3536]/_0_  (.Y(\inv_in[3537] ),
    .A(\inv_in[3536] ));
 sg13g2_inv_2 \inv[3537]/_0_  (.Y(\inv_in[3538] ),
    .A(\inv_in[3537] ));
 sg13g2_inv_2 \inv[3538]/_0_  (.Y(\inv_in[3539] ),
    .A(\inv_in[3538] ));
 sg13g2_inv_2 \inv[3539]/_0_  (.Y(\inv_in[3540] ),
    .A(\inv_in[3539] ));
 sg13g2_inv_2 \inv[353]/_0_  (.Y(\inv_in[354] ),
    .A(\inv_in[353] ));
 sg13g2_inv_2 \inv[3540]/_0_  (.Y(\inv_in[3541] ),
    .A(\inv_in[3540] ));
 sg13g2_inv_2 \inv[3541]/_0_  (.Y(\inv_in[3542] ),
    .A(\inv_in[3541] ));
 sg13g2_inv_2 \inv[3542]/_0_  (.Y(\inv_in[3543] ),
    .A(\inv_in[3542] ));
 sg13g2_inv_2 \inv[3543]/_0_  (.Y(\inv_in[3544] ),
    .A(\inv_in[3543] ));
 sg13g2_inv_2 \inv[3544]/_0_  (.Y(\inv_in[3545] ),
    .A(\inv_in[3544] ));
 sg13g2_inv_2 \inv[3545]/_0_  (.Y(\inv_in[3546] ),
    .A(\inv_in[3545] ));
 sg13g2_inv_2 \inv[3546]/_0_  (.Y(\inv_in[3547] ),
    .A(\inv_in[3546] ));
 sg13g2_inv_2 \inv[3547]/_0_  (.Y(\inv_in[3548] ),
    .A(\inv_in[3547] ));
 sg13g2_inv_2 \inv[3548]/_0_  (.Y(\inv_in[3549] ),
    .A(\inv_in[3548] ));
 sg13g2_inv_2 \inv[3549]/_0_  (.Y(\inv_in[3550] ),
    .A(\inv_in[3549] ));
 sg13g2_inv_2 \inv[354]/_0_  (.Y(\inv_in[355] ),
    .A(\inv_in[354] ));
 sg13g2_inv_2 \inv[3550]/_0_  (.Y(\inv_in[3551] ),
    .A(\inv_in[3550] ));
 sg13g2_inv_2 \inv[3551]/_0_  (.Y(\inv_in[3552] ),
    .A(\inv_in[3551] ));
 sg13g2_inv_2 \inv[3552]/_0_  (.Y(\inv_in[3553] ),
    .A(\inv_in[3552] ));
 sg13g2_inv_2 \inv[3553]/_0_  (.Y(\inv_in[3554] ),
    .A(\inv_in[3553] ));
 sg13g2_inv_2 \inv[3554]/_0_  (.Y(\inv_in[3555] ),
    .A(\inv_in[3554] ));
 sg13g2_inv_2 \inv[3555]/_0_  (.Y(\inv_in[3556] ),
    .A(\inv_in[3555] ));
 sg13g2_inv_2 \inv[3556]/_0_  (.Y(\inv_in[3557] ),
    .A(\inv_in[3556] ));
 sg13g2_inv_2 \inv[3557]/_0_  (.Y(\inv_in[3558] ),
    .A(\inv_in[3557] ));
 sg13g2_inv_2 \inv[3558]/_0_  (.Y(\inv_in[3559] ),
    .A(\inv_in[3558] ));
 sg13g2_inv_2 \inv[3559]/_0_  (.Y(\inv_in[3560] ),
    .A(\inv_in[3559] ));
 sg13g2_inv_2 \inv[355]/_0_  (.Y(\inv_in[356] ),
    .A(\inv_in[355] ));
 sg13g2_inv_2 \inv[3560]/_0_  (.Y(\inv_in[3561] ),
    .A(\inv_in[3560] ));
 sg13g2_inv_2 \inv[3561]/_0_  (.Y(\inv_in[3562] ),
    .A(\inv_in[3561] ));
 sg13g2_inv_2 \inv[3562]/_0_  (.Y(\inv_in[3563] ),
    .A(\inv_in[3562] ));
 sg13g2_inv_2 \inv[3563]/_0_  (.Y(\inv_in[3564] ),
    .A(\inv_in[3563] ));
 sg13g2_inv_2 \inv[3564]/_0_  (.Y(\inv_in[3565] ),
    .A(\inv_in[3564] ));
 sg13g2_inv_2 \inv[3565]/_0_  (.Y(\inv_in[3566] ),
    .A(\inv_in[3565] ));
 sg13g2_inv_2 \inv[3566]/_0_  (.Y(\inv_in[3567] ),
    .A(\inv_in[3566] ));
 sg13g2_inv_2 \inv[3567]/_0_  (.Y(\inv_in[3568] ),
    .A(\inv_in[3567] ));
 sg13g2_inv_2 \inv[3568]/_0_  (.Y(\inv_in[3569] ),
    .A(\inv_in[3568] ));
 sg13g2_inv_2 \inv[3569]/_0_  (.Y(\inv_in[3570] ),
    .A(\inv_in[3569] ));
 sg13g2_inv_2 \inv[356]/_0_  (.Y(\inv_in[357] ),
    .A(\inv_in[356] ));
 sg13g2_inv_2 \inv[3570]/_0_  (.Y(\inv_in[3571] ),
    .A(\inv_in[3570] ));
 sg13g2_inv_2 \inv[3571]/_0_  (.Y(\inv_in[3572] ),
    .A(\inv_in[3571] ));
 sg13g2_inv_2 \inv[3572]/_0_  (.Y(\inv_in[3573] ),
    .A(\inv_in[3572] ));
 sg13g2_inv_2 \inv[3573]/_0_  (.Y(\inv_in[3574] ),
    .A(\inv_in[3573] ));
 sg13g2_inv_2 \inv[3574]/_0_  (.Y(\inv_in[3575] ),
    .A(\inv_in[3574] ));
 sg13g2_inv_2 \inv[3575]/_0_  (.Y(\inv_in[3576] ),
    .A(\inv_in[3575] ));
 sg13g2_inv_2 \inv[3576]/_0_  (.Y(\inv_in[3577] ),
    .A(\inv_in[3576] ));
 sg13g2_inv_2 \inv[3577]/_0_  (.Y(\inv_in[3578] ),
    .A(\inv_in[3577] ));
 sg13g2_inv_2 \inv[3578]/_0_  (.Y(\inv_in[3579] ),
    .A(\inv_in[3578] ));
 sg13g2_inv_2 \inv[3579]/_0_  (.Y(\inv_in[3580] ),
    .A(\inv_in[3579] ));
 sg13g2_inv_2 \inv[357]/_0_  (.Y(\inv_in[358] ),
    .A(\inv_in[357] ));
 sg13g2_inv_2 \inv[3580]/_0_  (.Y(\inv_in[3581] ),
    .A(\inv_in[3580] ));
 sg13g2_inv_2 \inv[3581]/_0_  (.Y(\inv_in[3582] ),
    .A(\inv_in[3581] ));
 sg13g2_inv_2 \inv[3582]/_0_  (.Y(\inv_in[3583] ),
    .A(\inv_in[3582] ));
 sg13g2_inv_2 \inv[3583]/_0_  (.Y(\inv_in[3584] ),
    .A(\inv_in[3583] ));
 sg13g2_inv_2 \inv[3584]/_0_  (.Y(\inv_in[3585] ),
    .A(\inv_in[3584] ));
 sg13g2_inv_2 \inv[3585]/_0_  (.Y(\inv_in[3586] ),
    .A(\inv_in[3585] ));
 sg13g2_inv_2 \inv[3586]/_0_  (.Y(\inv_in[3587] ),
    .A(\inv_in[3586] ));
 sg13g2_inv_2 \inv[3587]/_0_  (.Y(\inv_in[3588] ),
    .A(\inv_in[3587] ));
 sg13g2_inv_2 \inv[3588]/_0_  (.Y(\inv_in[3589] ),
    .A(\inv_in[3588] ));
 sg13g2_inv_2 \inv[3589]/_0_  (.Y(\inv_in[3590] ),
    .A(\inv_in[3589] ));
 sg13g2_inv_2 \inv[358]/_0_  (.Y(\inv_in[359] ),
    .A(\inv_in[358] ));
 sg13g2_inv_2 \inv[3590]/_0_  (.Y(\inv_in[3591] ),
    .A(\inv_in[3590] ));
 sg13g2_inv_2 \inv[3591]/_0_  (.Y(\inv_in[3592] ),
    .A(\inv_in[3591] ));
 sg13g2_inv_2 \inv[3592]/_0_  (.Y(\inv_in[3593] ),
    .A(\inv_in[3592] ));
 sg13g2_inv_2 \inv[3593]/_0_  (.Y(\inv_in[3594] ),
    .A(\inv_in[3593] ));
 sg13g2_inv_2 \inv[3594]/_0_  (.Y(\inv_in[3595] ),
    .A(\inv_in[3594] ));
 sg13g2_inv_2 \inv[3595]/_0_  (.Y(\inv_in[3596] ),
    .A(\inv_in[3595] ));
 sg13g2_inv_2 \inv[3596]/_0_  (.Y(\inv_in[3597] ),
    .A(\inv_in[3596] ));
 sg13g2_inv_2 \inv[3597]/_0_  (.Y(\inv_in[3598] ),
    .A(\inv_in[3597] ));
 sg13g2_inv_2 \inv[3598]/_0_  (.Y(\inv_in[3599] ),
    .A(\inv_in[3598] ));
 sg13g2_inv_2 \inv[3599]/_0_  (.Y(\inv_in[3600] ),
    .A(\inv_in[3599] ));
 sg13g2_inv_2 \inv[359]/_0_  (.Y(\inv_in[360] ),
    .A(\inv_in[359] ));
 sg13g2_inv_2 \inv[35]/_0_  (.Y(\inv_in[36] ),
    .A(\inv_in[35] ));
 sg13g2_inv_2 \inv[3600]/_0_  (.Y(\inv_in[3601] ),
    .A(\inv_in[3600] ));
 sg13g2_inv_2 \inv[3601]/_0_  (.Y(\inv_in[3602] ),
    .A(\inv_in[3601] ));
 sg13g2_inv_2 \inv[3602]/_0_  (.Y(\inv_in[3603] ),
    .A(\inv_in[3602] ));
 sg13g2_inv_2 \inv[3603]/_0_  (.Y(\inv_in[3604] ),
    .A(\inv_in[3603] ));
 sg13g2_inv_2 \inv[3604]/_0_  (.Y(\inv_in[3605] ),
    .A(\inv_in[3604] ));
 sg13g2_inv_2 \inv[3605]/_0_  (.Y(\inv_in[3606] ),
    .A(\inv_in[3605] ));
 sg13g2_inv_2 \inv[3606]/_0_  (.Y(\inv_in[3607] ),
    .A(\inv_in[3606] ));
 sg13g2_inv_2 \inv[3607]/_0_  (.Y(\inv_in[3608] ),
    .A(\inv_in[3607] ));
 sg13g2_inv_2 \inv[3608]/_0_  (.Y(\inv_in[3609] ),
    .A(\inv_in[3608] ));
 sg13g2_inv_2 \inv[3609]/_0_  (.Y(\inv_in[3610] ),
    .A(\inv_in[3609] ));
 sg13g2_inv_2 \inv[360]/_0_  (.Y(\inv_in[361] ),
    .A(\inv_in[360] ));
 sg13g2_inv_2 \inv[3610]/_0_  (.Y(\inv_in[3611] ),
    .A(\inv_in[3610] ));
 sg13g2_inv_2 \inv[3611]/_0_  (.Y(\inv_in[3612] ),
    .A(\inv_in[3611] ));
 sg13g2_inv_2 \inv[3612]/_0_  (.Y(\inv_in[3613] ),
    .A(\inv_in[3612] ));
 sg13g2_inv_2 \inv[3613]/_0_  (.Y(\inv_in[3614] ),
    .A(\inv_in[3613] ));
 sg13g2_inv_2 \inv[3614]/_0_  (.Y(\inv_in[3615] ),
    .A(\inv_in[3614] ));
 sg13g2_inv_2 \inv[3615]/_0_  (.Y(\inv_in[3616] ),
    .A(\inv_in[3615] ));
 sg13g2_inv_2 \inv[3616]/_0_  (.Y(\inv_in[3617] ),
    .A(\inv_in[3616] ));
 sg13g2_inv_2 \inv[3617]/_0_  (.Y(\inv_in[3618] ),
    .A(\inv_in[3617] ));
 sg13g2_inv_2 \inv[3618]/_0_  (.Y(\inv_in[3619] ),
    .A(\inv_in[3618] ));
 sg13g2_inv_2 \inv[3619]/_0_  (.Y(\inv_in[3620] ),
    .A(\inv_in[3619] ));
 sg13g2_inv_2 \inv[361]/_0_  (.Y(\inv_in[362] ),
    .A(\inv_in[361] ));
 sg13g2_inv_2 \inv[3620]/_0_  (.Y(\inv_in[3621] ),
    .A(\inv_in[3620] ));
 sg13g2_inv_2 \inv[3621]/_0_  (.Y(\inv_in[3622] ),
    .A(\inv_in[3621] ));
 sg13g2_inv_2 \inv[3622]/_0_  (.Y(\inv_in[3623] ),
    .A(\inv_in[3622] ));
 sg13g2_inv_2 \inv[3623]/_0_  (.Y(\inv_in[3624] ),
    .A(\inv_in[3623] ));
 sg13g2_inv_2 \inv[3624]/_0_  (.Y(\inv_in[3625] ),
    .A(\inv_in[3624] ));
 sg13g2_inv_2 \inv[3625]/_0_  (.Y(\inv_in[3626] ),
    .A(\inv_in[3625] ));
 sg13g2_inv_2 \inv[3626]/_0_  (.Y(\inv_in[3627] ),
    .A(\inv_in[3626] ));
 sg13g2_inv_2 \inv[3627]/_0_  (.Y(\inv_in[3628] ),
    .A(\inv_in[3627] ));
 sg13g2_inv_2 \inv[3628]/_0_  (.Y(\inv_in[3629] ),
    .A(\inv_in[3628] ));
 sg13g2_inv_2 \inv[3629]/_0_  (.Y(\inv_in[3630] ),
    .A(\inv_in[3629] ));
 sg13g2_inv_2 \inv[362]/_0_  (.Y(\inv_in[363] ),
    .A(\inv_in[362] ));
 sg13g2_inv_2 \inv[3630]/_0_  (.Y(\inv_in[3631] ),
    .A(\inv_in[3630] ));
 sg13g2_inv_2 \inv[3631]/_0_  (.Y(\inv_in[3632] ),
    .A(\inv_in[3631] ));
 sg13g2_inv_2 \inv[3632]/_0_  (.Y(\inv_in[3633] ),
    .A(\inv_in[3632] ));
 sg13g2_inv_2 \inv[3633]/_0_  (.Y(\inv_in[3634] ),
    .A(\inv_in[3633] ));
 sg13g2_inv_2 \inv[3634]/_0_  (.Y(\inv_in[3635] ),
    .A(\inv_in[3634] ));
 sg13g2_inv_2 \inv[3635]/_0_  (.Y(\inv_in[3636] ),
    .A(\inv_in[3635] ));
 sg13g2_inv_2 \inv[3636]/_0_  (.Y(\inv_in[3637] ),
    .A(\inv_in[3636] ));
 sg13g2_inv_2 \inv[3637]/_0_  (.Y(\inv_in[3638] ),
    .A(\inv_in[3637] ));
 sg13g2_inv_2 \inv[3638]/_0_  (.Y(\inv_in[3639] ),
    .A(\inv_in[3638] ));
 sg13g2_inv_2 \inv[3639]/_0_  (.Y(\inv_in[3640] ),
    .A(\inv_in[3639] ));
 sg13g2_inv_2 \inv[363]/_0_  (.Y(\inv_in[364] ),
    .A(\inv_in[363] ));
 sg13g2_inv_2 \inv[3640]/_0_  (.Y(\inv_in[3641] ),
    .A(\inv_in[3640] ));
 sg13g2_inv_2 \inv[3641]/_0_  (.Y(\inv_in[3642] ),
    .A(\inv_in[3641] ));
 sg13g2_inv_2 \inv[3642]/_0_  (.Y(\inv_in[3643] ),
    .A(\inv_in[3642] ));
 sg13g2_inv_2 \inv[3643]/_0_  (.Y(\inv_in[3644] ),
    .A(\inv_in[3643] ));
 sg13g2_inv_2 \inv[3644]/_0_  (.Y(\inv_in[3645] ),
    .A(\inv_in[3644] ));
 sg13g2_inv_2 \inv[3645]/_0_  (.Y(\inv_in[3646] ),
    .A(\inv_in[3645] ));
 sg13g2_inv_2 \inv[3646]/_0_  (.Y(\inv_in[3647] ),
    .A(\inv_in[3646] ));
 sg13g2_inv_2 \inv[3647]/_0_  (.Y(\inv_in[3648] ),
    .A(\inv_in[3647] ));
 sg13g2_inv_2 \inv[3648]/_0_  (.Y(\inv_in[3649] ),
    .A(\inv_in[3648] ));
 sg13g2_inv_2 \inv[3649]/_0_  (.Y(\inv_in[3650] ),
    .A(\inv_in[3649] ));
 sg13g2_inv_2 \inv[364]/_0_  (.Y(\inv_in[365] ),
    .A(\inv_in[364] ));
 sg13g2_inv_2 \inv[3650]/_0_  (.Y(\inv_in[3651] ),
    .A(\inv_in[3650] ));
 sg13g2_inv_2 \inv[3651]/_0_  (.Y(\inv_in[3652] ),
    .A(\inv_in[3651] ));
 sg13g2_inv_2 \inv[3652]/_0_  (.Y(\inv_in[3653] ),
    .A(\inv_in[3652] ));
 sg13g2_inv_2 \inv[3653]/_0_  (.Y(\inv_in[3654] ),
    .A(\inv_in[3653] ));
 sg13g2_inv_2 \inv[3654]/_0_  (.Y(\inv_in[3655] ),
    .A(\inv_in[3654] ));
 sg13g2_inv_2 \inv[3655]/_0_  (.Y(\inv_in[3656] ),
    .A(\inv_in[3655] ));
 sg13g2_inv_2 \inv[3656]/_0_  (.Y(\inv_in[3657] ),
    .A(\inv_in[3656] ));
 sg13g2_inv_2 \inv[3657]/_0_  (.Y(\inv_in[3658] ),
    .A(\inv_in[3657] ));
 sg13g2_inv_2 \inv[3658]/_0_  (.Y(\inv_in[3659] ),
    .A(\inv_in[3658] ));
 sg13g2_inv_2 \inv[3659]/_0_  (.Y(\inv_in[3660] ),
    .A(\inv_in[3659] ));
 sg13g2_inv_2 \inv[365]/_0_  (.Y(\inv_in[366] ),
    .A(\inv_in[365] ));
 sg13g2_inv_2 \inv[3660]/_0_  (.Y(\inv_in[3661] ),
    .A(\inv_in[3660] ));
 sg13g2_inv_2 \inv[3661]/_0_  (.Y(\inv_in[3662] ),
    .A(\inv_in[3661] ));
 sg13g2_inv_2 \inv[3662]/_0_  (.Y(\inv_in[3663] ),
    .A(\inv_in[3662] ));
 sg13g2_inv_2 \inv[3663]/_0_  (.Y(\inv_in[3664] ),
    .A(\inv_in[3663] ));
 sg13g2_inv_2 \inv[3664]/_0_  (.Y(\inv_in[3665] ),
    .A(\inv_in[3664] ));
 sg13g2_inv_2 \inv[3665]/_0_  (.Y(\inv_in[3666] ),
    .A(\inv_in[3665] ));
 sg13g2_inv_2 \inv[3666]/_0_  (.Y(\inv_in[3667] ),
    .A(\inv_in[3666] ));
 sg13g2_inv_2 \inv[3667]/_0_  (.Y(\inv_in[3668] ),
    .A(\inv_in[3667] ));
 sg13g2_inv_2 \inv[3668]/_0_  (.Y(\inv_in[3669] ),
    .A(\inv_in[3668] ));
 sg13g2_inv_2 \inv[3669]/_0_  (.Y(\inv_in[3670] ),
    .A(\inv_in[3669] ));
 sg13g2_inv_2 \inv[366]/_0_  (.Y(\inv_in[367] ),
    .A(\inv_in[366] ));
 sg13g2_inv_2 \inv[3670]/_0_  (.Y(\inv_in[3671] ),
    .A(\inv_in[3670] ));
 sg13g2_inv_2 \inv[3671]/_0_  (.Y(\inv_in[3672] ),
    .A(\inv_in[3671] ));
 sg13g2_inv_2 \inv[3672]/_0_  (.Y(\inv_in[3673] ),
    .A(\inv_in[3672] ));
 sg13g2_inv_2 \inv[3673]/_0_  (.Y(\inv_in[3674] ),
    .A(\inv_in[3673] ));
 sg13g2_inv_2 \inv[3674]/_0_  (.Y(\inv_in[3675] ),
    .A(\inv_in[3674] ));
 sg13g2_inv_2 \inv[3675]/_0_  (.Y(\inv_in[3676] ),
    .A(\inv_in[3675] ));
 sg13g2_inv_2 \inv[3676]/_0_  (.Y(\inv_in[3677] ),
    .A(\inv_in[3676] ));
 sg13g2_inv_2 \inv[3677]/_0_  (.Y(\inv_in[3678] ),
    .A(\inv_in[3677] ));
 sg13g2_inv_2 \inv[3678]/_0_  (.Y(\inv_in[3679] ),
    .A(\inv_in[3678] ));
 sg13g2_inv_2 \inv[3679]/_0_  (.Y(\inv_in[3680] ),
    .A(\inv_in[3679] ));
 sg13g2_inv_2 \inv[367]/_0_  (.Y(\inv_in[368] ),
    .A(\inv_in[367] ));
 sg13g2_inv_2 \inv[3680]/_0_  (.Y(\inv_in[3681] ),
    .A(\inv_in[3680] ));
 sg13g2_inv_2 \inv[3681]/_0_  (.Y(\inv_in[3682] ),
    .A(\inv_in[3681] ));
 sg13g2_inv_2 \inv[3682]/_0_  (.Y(\inv_in[3683] ),
    .A(\inv_in[3682] ));
 sg13g2_inv_2 \inv[3683]/_0_  (.Y(\inv_in[3684] ),
    .A(\inv_in[3683] ));
 sg13g2_inv_2 \inv[3684]/_0_  (.Y(\inv_in[3685] ),
    .A(\inv_in[3684] ));
 sg13g2_inv_2 \inv[3685]/_0_  (.Y(\inv_in[3686] ),
    .A(\inv_in[3685] ));
 sg13g2_inv_2 \inv[3686]/_0_  (.Y(\inv_in[3687] ),
    .A(\inv_in[3686] ));
 sg13g2_inv_2 \inv[3687]/_0_  (.Y(\inv_in[3688] ),
    .A(\inv_in[3687] ));
 sg13g2_inv_2 \inv[3688]/_0_  (.Y(\inv_in[3689] ),
    .A(\inv_in[3688] ));
 sg13g2_inv_2 \inv[3689]/_0_  (.Y(\inv_in[3690] ),
    .A(\inv_in[3689] ));
 sg13g2_inv_2 \inv[368]/_0_  (.Y(\inv_in[369] ),
    .A(\inv_in[368] ));
 sg13g2_inv_2 \inv[3690]/_0_  (.Y(\inv_in[3691] ),
    .A(\inv_in[3690] ));
 sg13g2_inv_2 \inv[3691]/_0_  (.Y(\inv_in[3692] ),
    .A(\inv_in[3691] ));
 sg13g2_inv_2 \inv[3692]/_0_  (.Y(\inv_in[3693] ),
    .A(\inv_in[3692] ));
 sg13g2_inv_2 \inv[3693]/_0_  (.Y(\inv_in[3694] ),
    .A(\inv_in[3693] ));
 sg13g2_inv_2 \inv[3694]/_0_  (.Y(\inv_in[3695] ),
    .A(\inv_in[3694] ));
 sg13g2_inv_2 \inv[3695]/_0_  (.Y(\inv_in[3696] ),
    .A(\inv_in[3695] ));
 sg13g2_inv_2 \inv[3696]/_0_  (.Y(\inv_in[3697] ),
    .A(\inv_in[3696] ));
 sg13g2_inv_2 \inv[3697]/_0_  (.Y(\inv_in[3698] ),
    .A(\inv_in[3697] ));
 sg13g2_inv_2 \inv[3698]/_0_  (.Y(\inv_in[3699] ),
    .A(\inv_in[3698] ));
 sg13g2_inv_2 \inv[3699]/_0_  (.Y(\inv_in[3700] ),
    .A(\inv_in[3699] ));
 sg13g2_inv_2 \inv[369]/_0_  (.Y(\inv_in[370] ),
    .A(\inv_in[369] ));
 sg13g2_inv_2 \inv[36]/_0_  (.Y(\inv_in[37] ),
    .A(\inv_in[36] ));
 sg13g2_inv_2 \inv[3700]/_0_  (.Y(\inv_in[3701] ),
    .A(\inv_in[3700] ));
 sg13g2_inv_2 \inv[3701]/_0_  (.Y(\inv_in[3702] ),
    .A(\inv_in[3701] ));
 sg13g2_inv_2 \inv[3702]/_0_  (.Y(\inv_in[3703] ),
    .A(\inv_in[3702] ));
 sg13g2_inv_2 \inv[3703]/_0_  (.Y(\inv_in[3704] ),
    .A(\inv_in[3703] ));
 sg13g2_inv_2 \inv[3704]/_0_  (.Y(\inv_in[3705] ),
    .A(\inv_in[3704] ));
 sg13g2_inv_2 \inv[3705]/_0_  (.Y(\inv_in[3706] ),
    .A(\inv_in[3705] ));
 sg13g2_inv_2 \inv[3706]/_0_  (.Y(\inv_in[3707] ),
    .A(\inv_in[3706] ));
 sg13g2_inv_2 \inv[3707]/_0_  (.Y(\inv_in[3708] ),
    .A(\inv_in[3707] ));
 sg13g2_inv_2 \inv[3708]/_0_  (.Y(\inv_in[3709] ),
    .A(\inv_in[3708] ));
 sg13g2_inv_2 \inv[3709]/_0_  (.Y(\inv_in[3710] ),
    .A(\inv_in[3709] ));
 sg13g2_inv_2 \inv[370]/_0_  (.Y(\inv_in[371] ),
    .A(\inv_in[370] ));
 sg13g2_inv_2 \inv[3710]/_0_  (.Y(\inv_in[3711] ),
    .A(\inv_in[3710] ));
 sg13g2_inv_2 \inv[3711]/_0_  (.Y(\inv_in[3712] ),
    .A(\inv_in[3711] ));
 sg13g2_inv_2 \inv[3712]/_0_  (.Y(\inv_in[3713] ),
    .A(\inv_in[3712] ));
 sg13g2_inv_2 \inv[3713]/_0_  (.Y(\inv_in[3714] ),
    .A(\inv_in[3713] ));
 sg13g2_inv_2 \inv[3714]/_0_  (.Y(\inv_in[3715] ),
    .A(\inv_in[3714] ));
 sg13g2_inv_2 \inv[3715]/_0_  (.Y(\inv_in[3716] ),
    .A(\inv_in[3715] ));
 sg13g2_inv_2 \inv[3716]/_0_  (.Y(\inv_in[3717] ),
    .A(\inv_in[3716] ));
 sg13g2_inv_2 \inv[3717]/_0_  (.Y(\inv_in[3718] ),
    .A(\inv_in[3717] ));
 sg13g2_inv_2 \inv[3718]/_0_  (.Y(\inv_in[3719] ),
    .A(\inv_in[3718] ));
 sg13g2_inv_2 \inv[3719]/_0_  (.Y(\inv_in[3720] ),
    .A(\inv_in[3719] ));
 sg13g2_inv_2 \inv[371]/_0_  (.Y(\inv_in[372] ),
    .A(\inv_in[371] ));
 sg13g2_inv_2 \inv[3720]/_0_  (.Y(\inv_in[3721] ),
    .A(\inv_in[3720] ));
 sg13g2_inv_2 \inv[3721]/_0_  (.Y(\inv_in[3722] ),
    .A(\inv_in[3721] ));
 sg13g2_inv_2 \inv[3722]/_0_  (.Y(\inv_in[3723] ),
    .A(\inv_in[3722] ));
 sg13g2_inv_2 \inv[3723]/_0_  (.Y(\inv_in[3724] ),
    .A(\inv_in[3723] ));
 sg13g2_inv_2 \inv[3724]/_0_  (.Y(\inv_in[3725] ),
    .A(\inv_in[3724] ));
 sg13g2_inv_2 \inv[3725]/_0_  (.Y(\inv_in[3726] ),
    .A(\inv_in[3725] ));
 sg13g2_inv_2 \inv[3726]/_0_  (.Y(\inv_in[3727] ),
    .A(\inv_in[3726] ));
 sg13g2_inv_2 \inv[3727]/_0_  (.Y(\inv_in[3728] ),
    .A(\inv_in[3727] ));
 sg13g2_inv_2 \inv[3728]/_0_  (.Y(\inv_in[3729] ),
    .A(\inv_in[3728] ));
 sg13g2_inv_2 \inv[3729]/_0_  (.Y(\inv_in[3730] ),
    .A(\inv_in[3729] ));
 sg13g2_inv_2 \inv[372]/_0_  (.Y(\inv_in[373] ),
    .A(\inv_in[372] ));
 sg13g2_inv_2 \inv[3730]/_0_  (.Y(\inv_in[3731] ),
    .A(\inv_in[3730] ));
 sg13g2_inv_2 \inv[3731]/_0_  (.Y(\inv_in[3732] ),
    .A(\inv_in[3731] ));
 sg13g2_inv_2 \inv[3732]/_0_  (.Y(\inv_in[3733] ),
    .A(\inv_in[3732] ));
 sg13g2_inv_2 \inv[3733]/_0_  (.Y(\inv_in[3734] ),
    .A(\inv_in[3733] ));
 sg13g2_inv_2 \inv[3734]/_0_  (.Y(\inv_in[3735] ),
    .A(\inv_in[3734] ));
 sg13g2_inv_2 \inv[3735]/_0_  (.Y(\inv_in[3736] ),
    .A(\inv_in[3735] ));
 sg13g2_inv_2 \inv[3736]/_0_  (.Y(\inv_in[3737] ),
    .A(\inv_in[3736] ));
 sg13g2_inv_2 \inv[3737]/_0_  (.Y(\inv_in[3738] ),
    .A(\inv_in[3737] ));
 sg13g2_inv_2 \inv[3738]/_0_  (.Y(\inv_in[3739] ),
    .A(\inv_in[3738] ));
 sg13g2_inv_2 \inv[3739]/_0_  (.Y(\inv_in[3740] ),
    .A(\inv_in[3739] ));
 sg13g2_inv_2 \inv[373]/_0_  (.Y(\inv_in[374] ),
    .A(\inv_in[373] ));
 sg13g2_inv_2 \inv[3740]/_0_  (.Y(\inv_in[3741] ),
    .A(\inv_in[3740] ));
 sg13g2_inv_2 \inv[3741]/_0_  (.Y(\inv_in[3742] ),
    .A(\inv_in[3741] ));
 sg13g2_inv_2 \inv[3742]/_0_  (.Y(\inv_in[3743] ),
    .A(\inv_in[3742] ));
 sg13g2_inv_2 \inv[3743]/_0_  (.Y(\inv_in[3744] ),
    .A(\inv_in[3743] ));
 sg13g2_inv_2 \inv[3744]/_0_  (.Y(\inv_in[3745] ),
    .A(\inv_in[3744] ));
 sg13g2_inv_2 \inv[3745]/_0_  (.Y(\inv_in[3746] ),
    .A(\inv_in[3745] ));
 sg13g2_inv_2 \inv[3746]/_0_  (.Y(\inv_in[3747] ),
    .A(\inv_in[3746] ));
 sg13g2_inv_2 \inv[3747]/_0_  (.Y(\inv_in[3748] ),
    .A(\inv_in[3747] ));
 sg13g2_inv_2 \inv[3748]/_0_  (.Y(\inv_in[3749] ),
    .A(\inv_in[3748] ));
 sg13g2_inv_2 \inv[3749]/_0_  (.Y(\inv_in[3750] ),
    .A(\inv_in[3749] ));
 sg13g2_inv_2 \inv[374]/_0_  (.Y(\inv_in[375] ),
    .A(\inv_in[374] ));
 sg13g2_inv_2 \inv[3750]/_0_  (.Y(\inv_in[3751] ),
    .A(\inv_in[3750] ));
 sg13g2_inv_2 \inv[3751]/_0_  (.Y(\inv_in[3752] ),
    .A(\inv_in[3751] ));
 sg13g2_inv_2 \inv[3752]/_0_  (.Y(\inv_in[3753] ),
    .A(\inv_in[3752] ));
 sg13g2_inv_2 \inv[3753]/_0_  (.Y(\inv_in[3754] ),
    .A(\inv_in[3753] ));
 sg13g2_inv_2 \inv[3754]/_0_  (.Y(\inv_in[3755] ),
    .A(\inv_in[3754] ));
 sg13g2_inv_2 \inv[3755]/_0_  (.Y(\inv_in[3756] ),
    .A(\inv_in[3755] ));
 sg13g2_inv_2 \inv[3756]/_0_  (.Y(\inv_in[3757] ),
    .A(\inv_in[3756] ));
 sg13g2_inv_2 \inv[3757]/_0_  (.Y(\inv_in[3758] ),
    .A(\inv_in[3757] ));
 sg13g2_inv_2 \inv[3758]/_0_  (.Y(\inv_in[3759] ),
    .A(\inv_in[3758] ));
 sg13g2_inv_2 \inv[3759]/_0_  (.Y(\inv_in[3760] ),
    .A(\inv_in[3759] ));
 sg13g2_inv_2 \inv[375]/_0_  (.Y(\inv_in[376] ),
    .A(\inv_in[375] ));
 sg13g2_inv_2 \inv[3760]/_0_  (.Y(\inv_in[3761] ),
    .A(\inv_in[3760] ));
 sg13g2_inv_2 \inv[3761]/_0_  (.Y(\inv_in[3762] ),
    .A(\inv_in[3761] ));
 sg13g2_inv_4 \inv[3762]/_0_  (.A(\inv_in[3762] ),
    .Y(\inv_in[3763] ));
 sg13g2_inv_4 \inv[3763]/_0_  (.A(\inv_in[3763] ),
    .Y(\inv_in[3764] ));
 sg13g2_inv_4 \inv[3764]/_0_  (.A(\inv_in[3764] ),
    .Y(\inv_in[3765] ));
 sg13g2_inv_4 \inv[3765]/_0_  (.A(\inv_in[3765] ),
    .Y(\inv_in[3766] ));
 sg13g2_inv_4 \inv[3766]/_0_  (.A(\inv_in[3766] ),
    .Y(\inv_in[3767] ));
 sg13g2_inv_4 \inv[3767]/_0_  (.A(\inv_in[3767] ),
    .Y(\inv_in[3768] ));
 sg13g2_inv_2 \inv[3768]/_0_  (.Y(\inv_in[3769] ),
    .A(\inv_in[3768] ));
 sg13g2_inv_2 \inv[3769]/_0_  (.Y(\inv_in[3770] ),
    .A(\inv_in[3769] ));
 sg13g2_inv_2 \inv[376]/_0_  (.Y(\inv_in[377] ),
    .A(\inv_in[376] ));
 sg13g2_inv_4 \inv[3770]/_0_  (.A(\inv_in[3770] ),
    .Y(\inv_in[3771] ));
 sg13g2_inv_4 \inv[3771]/_0_  (.A(\inv_in[3771] ),
    .Y(\inv_in[3772] ));
 sg13g2_inv_4 \inv[3772]/_0_  (.A(\inv_in[3772] ),
    .Y(\inv_in[3773] ));
 sg13g2_inv_2 \inv[3773]/_0_  (.Y(\inv_in[3774] ),
    .A(\inv_in[3773] ));
 sg13g2_inv_2 \inv[3774]/_0_  (.Y(\inv_in[3775] ),
    .A(\inv_in[3774] ));
 sg13g2_inv_2 \inv[3775]/_0_  (.Y(\inv_in[3776] ),
    .A(\inv_in[3775] ));
 sg13g2_inv_2 \inv[3776]/_0_  (.Y(\inv_in[3777] ),
    .A(\inv_in[3776] ));
 sg13g2_inv_2 \inv[3777]/_0_  (.Y(\inv_in[3778] ),
    .A(\inv_in[3777] ));
 sg13g2_inv_2 \inv[3778]/_0_  (.Y(\inv_in[3779] ),
    .A(\inv_in[3778] ));
 sg13g2_inv_2 \inv[3779]/_0_  (.Y(\inv_in[3780] ),
    .A(\inv_in[3779] ));
 sg13g2_inv_2 \inv[377]/_0_  (.Y(\inv_in[378] ),
    .A(\inv_in[377] ));
 sg13g2_inv_4 \inv[3780]/_0_  (.A(\inv_in[3780] ),
    .Y(\inv_in[3781] ));
 sg13g2_inv_4 \inv[3781]/_0_  (.A(\inv_in[3781] ),
    .Y(\inv_in[3782] ));
 sg13g2_inv_2 \inv[3782]/_0_  (.Y(\inv_in[3783] ),
    .A(\inv_in[3782] ));
 sg13g2_inv_2 \inv[3783]/_0_  (.Y(\inv_in[3784] ),
    .A(\inv_in[3783] ));
 sg13g2_inv_2 \inv[3784]/_0_  (.Y(\inv_in[3785] ),
    .A(\inv_in[3784] ));
 sg13g2_inv_2 \inv[3785]/_0_  (.Y(\inv_in[3786] ),
    .A(\inv_in[3785] ));
 sg13g2_inv_2 \inv[3786]/_0_  (.Y(\inv_in[3787] ),
    .A(\inv_in[3786] ));
 sg13g2_inv_4 \inv[3787]/_0_  (.A(\inv_in[3787] ),
    .Y(\inv_in[3788] ));
 sg13g2_inv_4 \inv[3788]/_0_  (.A(\inv_in[3788] ),
    .Y(\inv_in[3789] ));
 sg13g2_inv_2 \inv[3789]/_0_  (.Y(\inv_in[3790] ),
    .A(\inv_in[3789] ));
 sg13g2_inv_2 \inv[378]/_0_  (.Y(\inv_in[379] ),
    .A(\inv_in[378] ));
 sg13g2_inv_2 \inv[3790]/_0_  (.Y(\inv_in[3791] ),
    .A(\inv_in[3790] ));
 sg13g2_inv_2 \inv[3791]/_0_  (.Y(\inv_in[3792] ),
    .A(\inv_in[3791] ));
 sg13g2_inv_2 \inv[3792]/_0_  (.Y(\inv_in[3793] ),
    .A(\inv_in[3792] ));
 sg13g2_inv_2 \inv[3793]/_0_  (.Y(\inv_in[3794] ),
    .A(\inv_in[3793] ));
 sg13g2_inv_2 \inv[3794]/_0_  (.Y(\inv_in[3795] ),
    .A(\inv_in[3794] ));
 sg13g2_inv_2 \inv[3795]/_0_  (.Y(\inv_in[3796] ),
    .A(\inv_in[3795] ));
 sg13g2_inv_2 \inv[3796]/_0_  (.Y(\inv_in[3797] ),
    .A(\inv_in[3796] ));
 sg13g2_inv_2 \inv[3797]/_0_  (.Y(\inv_in[3798] ),
    .A(\inv_in[3797] ));
 sg13g2_inv_2 \inv[3798]/_0_  (.Y(\inv_in[3799] ),
    .A(\inv_in[3798] ));
 sg13g2_inv_2 \inv[3799]/_0_  (.Y(\inv_in[3800] ),
    .A(\inv_in[3799] ));
 sg13g2_inv_2 \inv[379]/_0_  (.Y(\inv_in[380] ),
    .A(\inv_in[379] ));
 sg13g2_inv_2 \inv[37]/_0_  (.Y(\inv_in[38] ),
    .A(\inv_in[37] ));
 sg13g2_inv_2 \inv[3800]/_0_  (.Y(\inv_in[3801] ),
    .A(\inv_in[3800] ));
 sg13g2_inv_2 \inv[3801]/_0_  (.Y(\inv_in[3802] ),
    .A(\inv_in[3801] ));
 sg13g2_inv_2 \inv[3802]/_0_  (.Y(\inv_in[3803] ),
    .A(\inv_in[3802] ));
 sg13g2_inv_2 \inv[3803]/_0_  (.Y(\inv_in[3804] ),
    .A(\inv_in[3803] ));
 sg13g2_inv_2 \inv[3804]/_0_  (.Y(\inv_in[3805] ),
    .A(\inv_in[3804] ));
 sg13g2_inv_2 \inv[3805]/_0_  (.Y(\inv_in[3806] ),
    .A(\inv_in[3805] ));
 sg13g2_inv_2 \inv[3806]/_0_  (.Y(\inv_in[3807] ),
    .A(\inv_in[3806] ));
 sg13g2_inv_2 \inv[3807]/_0_  (.Y(\inv_in[3808] ),
    .A(\inv_in[3807] ));
 sg13g2_inv_2 \inv[3808]/_0_  (.Y(\inv_in[3809] ),
    .A(\inv_in[3808] ));
 sg13g2_inv_2 \inv[3809]/_0_  (.Y(\inv_in[3810] ),
    .A(\inv_in[3809] ));
 sg13g2_inv_2 \inv[380]/_0_  (.Y(\inv_in[381] ),
    .A(\inv_in[380] ));
 sg13g2_inv_2 \inv[3810]/_0_  (.Y(\inv_in[3811] ),
    .A(\inv_in[3810] ));
 sg13g2_inv_2 \inv[3811]/_0_  (.Y(\inv_in[3812] ),
    .A(\inv_in[3811] ));
 sg13g2_inv_2 \inv[3812]/_0_  (.Y(\inv_in[3813] ),
    .A(\inv_in[3812] ));
 sg13g2_inv_2 \inv[3813]/_0_  (.Y(\inv_in[3814] ),
    .A(\inv_in[3813] ));
 sg13g2_inv_2 \inv[3814]/_0_  (.Y(\inv_in[3815] ),
    .A(\inv_in[3814] ));
 sg13g2_inv_2 \inv[3815]/_0_  (.Y(\inv_in[3816] ),
    .A(\inv_in[3815] ));
 sg13g2_inv_2 \inv[3816]/_0_  (.Y(\inv_in[3817] ),
    .A(\inv_in[3816] ));
 sg13g2_inv_2 \inv[3817]/_0_  (.Y(\inv_in[3818] ),
    .A(\inv_in[3817] ));
 sg13g2_inv_2 \inv[3818]/_0_  (.Y(\inv_in[3819] ),
    .A(\inv_in[3818] ));
 sg13g2_inv_2 \inv[3819]/_0_  (.Y(\inv_in[3820] ),
    .A(\inv_in[3819] ));
 sg13g2_inv_2 \inv[381]/_0_  (.Y(\inv_in[382] ),
    .A(\inv_in[381] ));
 sg13g2_inv_2 \inv[3820]/_0_  (.Y(\inv_in[3821] ),
    .A(\inv_in[3820] ));
 sg13g2_inv_2 \inv[3821]/_0_  (.Y(\inv_in[3822] ),
    .A(\inv_in[3821] ));
 sg13g2_inv_2 \inv[3822]/_0_  (.Y(\inv_in[3823] ),
    .A(\inv_in[3822] ));
 sg13g2_inv_2 \inv[3823]/_0_  (.Y(\inv_in[3824] ),
    .A(\inv_in[3823] ));
 sg13g2_inv_2 \inv[3824]/_0_  (.Y(\inv_in[3825] ),
    .A(\inv_in[3824] ));
 sg13g2_inv_2 \inv[3825]/_0_  (.Y(\inv_in[3826] ),
    .A(\inv_in[3825] ));
 sg13g2_inv_2 \inv[3826]/_0_  (.Y(\inv_in[3827] ),
    .A(\inv_in[3826] ));
 sg13g2_inv_2 \inv[3827]/_0_  (.Y(\inv_in[3828] ),
    .A(\inv_in[3827] ));
 sg13g2_inv_2 \inv[3828]/_0_  (.Y(\inv_in[3829] ),
    .A(\inv_in[3828] ));
 sg13g2_inv_2 \inv[3829]/_0_  (.Y(\inv_in[3830] ),
    .A(\inv_in[3829] ));
 sg13g2_inv_2 \inv[382]/_0_  (.Y(\inv_in[383] ),
    .A(\inv_in[382] ));
 sg13g2_inv_2 \inv[3830]/_0_  (.Y(\inv_in[3831] ),
    .A(\inv_in[3830] ));
 sg13g2_inv_2 \inv[3831]/_0_  (.Y(\inv_in[3832] ),
    .A(\inv_in[3831] ));
 sg13g2_inv_2 \inv[3832]/_0_  (.Y(\inv_in[3833] ),
    .A(\inv_in[3832] ));
 sg13g2_inv_2 \inv[3833]/_0_  (.Y(\inv_in[3834] ),
    .A(\inv_in[3833] ));
 sg13g2_inv_2 \inv[3834]/_0_  (.Y(\inv_in[3835] ),
    .A(\inv_in[3834] ));
 sg13g2_inv_2 \inv[3835]/_0_  (.Y(\inv_in[3836] ),
    .A(\inv_in[3835] ));
 sg13g2_inv_2 \inv[3836]/_0_  (.Y(\inv_in[3837] ),
    .A(\inv_in[3836] ));
 sg13g2_inv_2 \inv[3837]/_0_  (.Y(\inv_in[3838] ),
    .A(\inv_in[3837] ));
 sg13g2_inv_2 \inv[3838]/_0_  (.Y(\inv_in[3839] ),
    .A(\inv_in[3838] ));
 sg13g2_inv_2 \inv[3839]/_0_  (.Y(\inv_in[3840] ),
    .A(\inv_in[3839] ));
 sg13g2_inv_2 \inv[383]/_0_  (.Y(\inv_in[384] ),
    .A(\inv_in[383] ));
 sg13g2_inv_2 \inv[3840]/_0_  (.Y(\inv_in[3841] ),
    .A(\inv_in[3840] ));
 sg13g2_inv_2 \inv[3841]/_0_  (.Y(\inv_in[3842] ),
    .A(\inv_in[3841] ));
 sg13g2_inv_2 \inv[3842]/_0_  (.Y(\inv_in[3843] ),
    .A(\inv_in[3842] ));
 sg13g2_inv_2 \inv[3843]/_0_  (.Y(\inv_in[3844] ),
    .A(\inv_in[3843] ));
 sg13g2_inv_2 \inv[3844]/_0_  (.Y(\inv_in[3845] ),
    .A(\inv_in[3844] ));
 sg13g2_inv_2 \inv[3845]/_0_  (.Y(\inv_in[3846] ),
    .A(\inv_in[3845] ));
 sg13g2_inv_2 \inv[3846]/_0_  (.Y(\inv_in[3847] ),
    .A(\inv_in[3846] ));
 sg13g2_inv_2 \inv[3847]/_0_  (.Y(\inv_in[3848] ),
    .A(\inv_in[3847] ));
 sg13g2_inv_2 \inv[3848]/_0_  (.Y(\inv_in[3849] ),
    .A(\inv_in[3848] ));
 sg13g2_inv_2 \inv[3849]/_0_  (.Y(\inv_in[3850] ),
    .A(\inv_in[3849] ));
 sg13g2_inv_2 \inv[384]/_0_  (.Y(\inv_in[385] ),
    .A(\inv_in[384] ));
 sg13g2_inv_2 \inv[3850]/_0_  (.Y(\inv_in[3851] ),
    .A(\inv_in[3850] ));
 sg13g2_inv_2 \inv[3851]/_0_  (.Y(\inv_in[3852] ),
    .A(\inv_in[3851] ));
 sg13g2_inv_2 \inv[3852]/_0_  (.Y(net7),
    .A(\inv_in[3852] ));
 sg13g2_inv_2 \inv[385]/_0_  (.Y(\inv_in[386] ),
    .A(\inv_in[385] ));
 sg13g2_inv_2 \inv[386]/_0_  (.Y(\inv_in[387] ),
    .A(\inv_in[386] ));
 sg13g2_inv_2 \inv[387]/_0_  (.Y(\inv_in[388] ),
    .A(\inv_in[387] ));
 sg13g2_inv_2 \inv[388]/_0_  (.Y(\inv_in[389] ),
    .A(\inv_in[388] ));
 sg13g2_inv_2 \inv[389]/_0_  (.Y(\inv_in[390] ),
    .A(\inv_in[389] ));
 sg13g2_inv_2 \inv[38]/_0_  (.Y(\inv_in[39] ),
    .A(\inv_in[38] ));
 sg13g2_inv_2 \inv[390]/_0_  (.Y(\inv_in[391] ),
    .A(\inv_in[390] ));
 sg13g2_inv_2 \inv[391]/_0_  (.Y(\inv_in[392] ),
    .A(\inv_in[391] ));
 sg13g2_inv_2 \inv[392]/_0_  (.Y(\inv_in[393] ),
    .A(\inv_in[392] ));
 sg13g2_inv_2 \inv[393]/_0_  (.Y(\inv_in[394] ),
    .A(\inv_in[393] ));
 sg13g2_inv_2 \inv[394]/_0_  (.Y(\inv_in[395] ),
    .A(\inv_in[394] ));
 sg13g2_inv_2 \inv[395]/_0_  (.Y(\inv_in[396] ),
    .A(\inv_in[395] ));
 sg13g2_inv_2 \inv[396]/_0_  (.Y(\inv_in[397] ),
    .A(\inv_in[396] ));
 sg13g2_inv_2 \inv[397]/_0_  (.Y(\inv_in[398] ),
    .A(\inv_in[397] ));
 sg13g2_inv_2 \inv[398]/_0_  (.Y(\inv_in[399] ),
    .A(\inv_in[398] ));
 sg13g2_inv_2 \inv[399]/_0_  (.Y(\inv_in[400] ),
    .A(\inv_in[399] ));
 sg13g2_inv_2 \inv[39]/_0_  (.Y(\inv_in[40] ),
    .A(\inv_in[39] ));
 sg13g2_inv_2 \inv[3]/_0_  (.Y(\inv_in[4] ),
    .A(\inv_in[3] ));
 sg13g2_inv_2 \inv[400]/_0_  (.Y(\inv_in[401] ),
    .A(\inv_in[400] ));
 sg13g2_inv_2 \inv[401]/_0_  (.Y(\inv_in[402] ),
    .A(\inv_in[401] ));
 sg13g2_inv_2 \inv[402]/_0_  (.Y(\inv_in[403] ),
    .A(\inv_in[402] ));
 sg13g2_inv_2 \inv[403]/_0_  (.Y(\inv_in[404] ),
    .A(\inv_in[403] ));
 sg13g2_inv_2 \inv[404]/_0_  (.Y(\inv_in[405] ),
    .A(\inv_in[404] ));
 sg13g2_inv_2 \inv[405]/_0_  (.Y(\inv_in[406] ),
    .A(\inv_in[405] ));
 sg13g2_inv_2 \inv[406]/_0_  (.Y(\inv_in[407] ),
    .A(\inv_in[406] ));
 sg13g2_inv_2 \inv[407]/_0_  (.Y(\inv_in[408] ),
    .A(\inv_in[407] ));
 sg13g2_inv_2 \inv[408]/_0_  (.Y(\inv_in[409] ),
    .A(\inv_in[408] ));
 sg13g2_inv_2 \inv[409]/_0_  (.Y(\inv_in[410] ),
    .A(\inv_in[409] ));
 sg13g2_inv_2 \inv[40]/_0_  (.Y(\inv_in[41] ),
    .A(\inv_in[40] ));
 sg13g2_inv_2 \inv[410]/_0_  (.Y(\inv_in[411] ),
    .A(\inv_in[410] ));
 sg13g2_inv_2 \inv[411]/_0_  (.Y(\inv_in[412] ),
    .A(\inv_in[411] ));
 sg13g2_inv_2 \inv[412]/_0_  (.Y(\inv_in[413] ),
    .A(\inv_in[412] ));
 sg13g2_inv_2 \inv[413]/_0_  (.Y(\inv_in[414] ),
    .A(\inv_in[413] ));
 sg13g2_inv_2 \inv[414]/_0_  (.Y(\inv_in[415] ),
    .A(\inv_in[414] ));
 sg13g2_inv_2 \inv[415]/_0_  (.Y(\inv_in[416] ),
    .A(\inv_in[415] ));
 sg13g2_inv_2 \inv[416]/_0_  (.Y(\inv_in[417] ),
    .A(\inv_in[416] ));
 sg13g2_inv_2 \inv[417]/_0_  (.Y(\inv_in[418] ),
    .A(\inv_in[417] ));
 sg13g2_inv_2 \inv[418]/_0_  (.Y(\inv_in[419] ),
    .A(\inv_in[418] ));
 sg13g2_inv_2 \inv[419]/_0_  (.Y(\inv_in[420] ),
    .A(\inv_in[419] ));
 sg13g2_inv_2 \inv[41]/_0_  (.Y(\inv_in[42] ),
    .A(\inv_in[41] ));
 sg13g2_inv_2 \inv[420]/_0_  (.Y(\inv_in[421] ),
    .A(\inv_in[420] ));
 sg13g2_inv_2 \inv[421]/_0_  (.Y(\inv_in[422] ),
    .A(\inv_in[421] ));
 sg13g2_inv_2 \inv[422]/_0_  (.Y(\inv_in[423] ),
    .A(\inv_in[422] ));
 sg13g2_inv_2 \inv[423]/_0_  (.Y(\inv_in[424] ),
    .A(\inv_in[423] ));
 sg13g2_inv_2 \inv[424]/_0_  (.Y(\inv_in[425] ),
    .A(\inv_in[424] ));
 sg13g2_inv_2 \inv[425]/_0_  (.Y(\inv_in[426] ),
    .A(\inv_in[425] ));
 sg13g2_inv_2 \inv[426]/_0_  (.Y(\inv_in[427] ),
    .A(\inv_in[426] ));
 sg13g2_inv_2 \inv[427]/_0_  (.Y(\inv_in[428] ),
    .A(\inv_in[427] ));
 sg13g2_inv_2 \inv[428]/_0_  (.Y(\inv_in[429] ),
    .A(\inv_in[428] ));
 sg13g2_inv_2 \inv[429]/_0_  (.Y(\inv_in[430] ),
    .A(\inv_in[429] ));
 sg13g2_inv_2 \inv[42]/_0_  (.Y(\inv_in[43] ),
    .A(\inv_in[42] ));
 sg13g2_inv_2 \inv[430]/_0_  (.Y(\inv_in[431] ),
    .A(\inv_in[430] ));
 sg13g2_inv_2 \inv[431]/_0_  (.Y(\inv_in[432] ),
    .A(\inv_in[431] ));
 sg13g2_inv_2 \inv[432]/_0_  (.Y(\inv_in[433] ),
    .A(\inv_in[432] ));
 sg13g2_inv_2 \inv[433]/_0_  (.Y(\inv_in[434] ),
    .A(\inv_in[433] ));
 sg13g2_inv_2 \inv[434]/_0_  (.Y(\inv_in[435] ),
    .A(\inv_in[434] ));
 sg13g2_inv_2 \inv[435]/_0_  (.Y(\inv_in[436] ),
    .A(\inv_in[435] ));
 sg13g2_inv_2 \inv[436]/_0_  (.Y(\inv_in[437] ),
    .A(\inv_in[436] ));
 sg13g2_inv_2 \inv[437]/_0_  (.Y(\inv_in[438] ),
    .A(\inv_in[437] ));
 sg13g2_inv_2 \inv[438]/_0_  (.Y(\inv_in[439] ),
    .A(\inv_in[438] ));
 sg13g2_inv_2 \inv[439]/_0_  (.Y(\inv_in[440] ),
    .A(\inv_in[439] ));
 sg13g2_inv_2 \inv[43]/_0_  (.Y(\inv_in[44] ),
    .A(\inv_in[43] ));
 sg13g2_inv_2 \inv[440]/_0_  (.Y(\inv_in[441] ),
    .A(\inv_in[440] ));
 sg13g2_inv_2 \inv[441]/_0_  (.Y(\inv_in[442] ),
    .A(\inv_in[441] ));
 sg13g2_inv_2 \inv[442]/_0_  (.Y(\inv_in[443] ),
    .A(\inv_in[442] ));
 sg13g2_inv_2 \inv[443]/_0_  (.Y(\inv_in[444] ),
    .A(\inv_in[443] ));
 sg13g2_inv_2 \inv[444]/_0_  (.Y(\inv_in[445] ),
    .A(\inv_in[444] ));
 sg13g2_inv_2 \inv[445]/_0_  (.Y(\inv_in[446] ),
    .A(\inv_in[445] ));
 sg13g2_inv_2 \inv[446]/_0_  (.Y(\inv_in[447] ),
    .A(\inv_in[446] ));
 sg13g2_inv_2 \inv[447]/_0_  (.Y(\inv_in[448] ),
    .A(\inv_in[447] ));
 sg13g2_inv_2 \inv[448]/_0_  (.Y(\inv_in[449] ),
    .A(\inv_in[448] ));
 sg13g2_inv_2 \inv[449]/_0_  (.Y(\inv_in[450] ),
    .A(\inv_in[449] ));
 sg13g2_inv_2 \inv[44]/_0_  (.Y(\inv_in[45] ),
    .A(\inv_in[44] ));
 sg13g2_inv_2 \inv[450]/_0_  (.Y(\inv_in[451] ),
    .A(\inv_in[450] ));
 sg13g2_inv_2 \inv[451]/_0_  (.Y(\inv_in[452] ),
    .A(\inv_in[451] ));
 sg13g2_inv_2 \inv[452]/_0_  (.Y(\inv_in[453] ),
    .A(\inv_in[452] ));
 sg13g2_inv_2 \inv[453]/_0_  (.Y(\inv_in[454] ),
    .A(\inv_in[453] ));
 sg13g2_inv_2 \inv[454]/_0_  (.Y(\inv_in[455] ),
    .A(\inv_in[454] ));
 sg13g2_inv_2 \inv[455]/_0_  (.Y(\inv_in[456] ),
    .A(\inv_in[455] ));
 sg13g2_inv_2 \inv[456]/_0_  (.Y(\inv_in[457] ),
    .A(\inv_in[456] ));
 sg13g2_inv_2 \inv[457]/_0_  (.Y(\inv_in[458] ),
    .A(\inv_in[457] ));
 sg13g2_inv_2 \inv[458]/_0_  (.Y(\inv_in[459] ),
    .A(\inv_in[458] ));
 sg13g2_inv_2 \inv[459]/_0_  (.Y(\inv_in[460] ),
    .A(\inv_in[459] ));
 sg13g2_inv_2 \inv[45]/_0_  (.Y(\inv_in[46] ),
    .A(\inv_in[45] ));
 sg13g2_inv_2 \inv[460]/_0_  (.Y(\inv_in[461] ),
    .A(\inv_in[460] ));
 sg13g2_inv_2 \inv[461]/_0_  (.Y(\inv_in[462] ),
    .A(\inv_in[461] ));
 sg13g2_inv_2 \inv[462]/_0_  (.Y(\inv_in[463] ),
    .A(\inv_in[462] ));
 sg13g2_inv_2 \inv[463]/_0_  (.Y(\inv_in[464] ),
    .A(\inv_in[463] ));
 sg13g2_inv_2 \inv[464]/_0_  (.Y(\inv_in[465] ),
    .A(\inv_in[464] ));
 sg13g2_inv_2 \inv[465]/_0_  (.Y(\inv_in[466] ),
    .A(\inv_in[465] ));
 sg13g2_inv_2 \inv[466]/_0_  (.Y(\inv_in[467] ),
    .A(\inv_in[466] ));
 sg13g2_inv_2 \inv[467]/_0_  (.Y(\inv_in[468] ),
    .A(\inv_in[467] ));
 sg13g2_inv_2 \inv[468]/_0_  (.Y(\inv_in[469] ),
    .A(\inv_in[468] ));
 sg13g2_inv_2 \inv[469]/_0_  (.Y(\inv_in[470] ),
    .A(\inv_in[469] ));
 sg13g2_inv_2 \inv[46]/_0_  (.Y(\inv_in[47] ),
    .A(\inv_in[46] ));
 sg13g2_inv_2 \inv[470]/_0_  (.Y(\inv_in[471] ),
    .A(\inv_in[470] ));
 sg13g2_inv_2 \inv[471]/_0_  (.Y(\inv_in[472] ),
    .A(\inv_in[471] ));
 sg13g2_inv_2 \inv[472]/_0_  (.Y(\inv_in[473] ),
    .A(\inv_in[472] ));
 sg13g2_inv_2 \inv[473]/_0_  (.Y(\inv_in[474] ),
    .A(\inv_in[473] ));
 sg13g2_inv_2 \inv[474]/_0_  (.Y(\inv_in[475] ),
    .A(\inv_in[474] ));
 sg13g2_inv_2 \inv[475]/_0_  (.Y(\inv_in[476] ),
    .A(\inv_in[475] ));
 sg13g2_inv_2 \inv[476]/_0_  (.Y(\inv_in[477] ),
    .A(\inv_in[476] ));
 sg13g2_inv_2 \inv[477]/_0_  (.Y(\inv_in[478] ),
    .A(\inv_in[477] ));
 sg13g2_inv_2 \inv[478]/_0_  (.Y(\inv_in[479] ),
    .A(\inv_in[478] ));
 sg13g2_inv_2 \inv[479]/_0_  (.Y(\inv_in[480] ),
    .A(\inv_in[479] ));
 sg13g2_inv_2 \inv[47]/_0_  (.Y(\inv_in[48] ),
    .A(\inv_in[47] ));
 sg13g2_inv_2 \inv[480]/_0_  (.Y(\inv_in[481] ),
    .A(\inv_in[480] ));
 sg13g2_inv_2 \inv[481]/_0_  (.Y(\inv_in[482] ),
    .A(\inv_in[481] ));
 sg13g2_inv_2 \inv[482]/_0_  (.Y(\inv_in[483] ),
    .A(\inv_in[482] ));
 sg13g2_inv_2 \inv[483]/_0_  (.Y(\inv_in[484] ),
    .A(\inv_in[483] ));
 sg13g2_inv_2 \inv[484]/_0_  (.Y(\inv_in[485] ),
    .A(\inv_in[484] ));
 sg13g2_inv_2 \inv[485]/_0_  (.Y(\inv_in[486] ),
    .A(\inv_in[485] ));
 sg13g2_inv_2 \inv[486]/_0_  (.Y(\inv_in[487] ),
    .A(\inv_in[486] ));
 sg13g2_inv_2 \inv[487]/_0_  (.Y(\inv_in[488] ),
    .A(\inv_in[487] ));
 sg13g2_inv_2 \inv[488]/_0_  (.Y(\inv_in[489] ),
    .A(\inv_in[488] ));
 sg13g2_inv_2 \inv[489]/_0_  (.Y(\inv_in[490] ),
    .A(\inv_in[489] ));
 sg13g2_inv_2 \inv[48]/_0_  (.Y(\inv_in[49] ),
    .A(\inv_in[48] ));
 sg13g2_inv_2 \inv[490]/_0_  (.Y(\inv_in[491] ),
    .A(\inv_in[490] ));
 sg13g2_inv_2 \inv[491]/_0_  (.Y(\inv_in[492] ),
    .A(\inv_in[491] ));
 sg13g2_inv_2 \inv[492]/_0_  (.Y(\inv_in[493] ),
    .A(\inv_in[492] ));
 sg13g2_inv_2 \inv[493]/_0_  (.Y(\inv_in[494] ),
    .A(\inv_in[493] ));
 sg13g2_inv_2 \inv[494]/_0_  (.Y(\inv_in[495] ),
    .A(\inv_in[494] ));
 sg13g2_inv_2 \inv[495]/_0_  (.Y(\inv_in[496] ),
    .A(\inv_in[495] ));
 sg13g2_inv_2 \inv[496]/_0_  (.Y(\inv_in[497] ),
    .A(\inv_in[496] ));
 sg13g2_inv_2 \inv[497]/_0_  (.Y(\inv_in[498] ),
    .A(\inv_in[497] ));
 sg13g2_inv_2 \inv[498]/_0_  (.Y(\inv_in[499] ),
    .A(\inv_in[498] ));
 sg13g2_inv_2 \inv[499]/_0_  (.Y(\inv_in[500] ),
    .A(\inv_in[499] ));
 sg13g2_inv_2 \inv[49]/_0_  (.Y(\inv_in[50] ),
    .A(\inv_in[49] ));
 sg13g2_inv_2 \inv[4]/_0_  (.Y(\inv_in[5] ),
    .A(\inv_in[4] ));
 sg13g2_inv_2 \inv[500]/_0_  (.Y(\inv_in[501] ),
    .A(\inv_in[500] ));
 sg13g2_inv_2 \inv[501]/_0_  (.Y(\inv_in[502] ),
    .A(\inv_in[501] ));
 sg13g2_inv_2 \inv[502]/_0_  (.Y(\inv_in[503] ),
    .A(\inv_in[502] ));
 sg13g2_inv_2 \inv[503]/_0_  (.Y(\inv_in[504] ),
    .A(\inv_in[503] ));
 sg13g2_inv_2 \inv[504]/_0_  (.Y(\inv_in[505] ),
    .A(\inv_in[504] ));
 sg13g2_inv_2 \inv[505]/_0_  (.Y(\inv_in[506] ),
    .A(\inv_in[505] ));
 sg13g2_inv_2 \inv[506]/_0_  (.Y(\inv_in[507] ),
    .A(\inv_in[506] ));
 sg13g2_inv_2 \inv[507]/_0_  (.Y(\inv_in[508] ),
    .A(\inv_in[507] ));
 sg13g2_inv_2 \inv[508]/_0_  (.Y(\inv_in[509] ),
    .A(\inv_in[508] ));
 sg13g2_inv_2 \inv[509]/_0_  (.Y(\inv_in[510] ),
    .A(\inv_in[509] ));
 sg13g2_inv_2 \inv[50]/_0_  (.Y(\inv_in[51] ),
    .A(\inv_in[50] ));
 sg13g2_inv_2 \inv[510]/_0_  (.Y(\inv_in[511] ),
    .A(\inv_in[510] ));
 sg13g2_inv_2 \inv[511]/_0_  (.Y(\inv_in[512] ),
    .A(\inv_in[511] ));
 sg13g2_inv_2 \inv[512]/_0_  (.Y(\inv_in[513] ),
    .A(\inv_in[512] ));
 sg13g2_inv_2 \inv[513]/_0_  (.Y(\inv_in[514] ),
    .A(\inv_in[513] ));
 sg13g2_inv_2 \inv[514]/_0_  (.Y(\inv_in[515] ),
    .A(\inv_in[514] ));
 sg13g2_inv_2 \inv[515]/_0_  (.Y(\inv_in[516] ),
    .A(\inv_in[515] ));
 sg13g2_inv_2 \inv[516]/_0_  (.Y(\inv_in[517] ),
    .A(\inv_in[516] ));
 sg13g2_inv_2 \inv[517]/_0_  (.Y(\inv_in[518] ),
    .A(\inv_in[517] ));
 sg13g2_inv_2 \inv[518]/_0_  (.Y(\inv_in[519] ),
    .A(\inv_in[518] ));
 sg13g2_inv_2 \inv[519]/_0_  (.Y(\inv_in[520] ),
    .A(\inv_in[519] ));
 sg13g2_inv_2 \inv[51]/_0_  (.Y(\inv_in[52] ),
    .A(\inv_in[51] ));
 sg13g2_inv_2 \inv[520]/_0_  (.Y(\inv_in[521] ),
    .A(\inv_in[520] ));
 sg13g2_inv_2 \inv[521]/_0_  (.Y(\inv_in[522] ),
    .A(\inv_in[521] ));
 sg13g2_inv_2 \inv[522]/_0_  (.Y(\inv_in[523] ),
    .A(\inv_in[522] ));
 sg13g2_inv_2 \inv[523]/_0_  (.Y(\inv_in[524] ),
    .A(\inv_in[523] ));
 sg13g2_inv_2 \inv[524]/_0_  (.Y(\inv_in[525] ),
    .A(\inv_in[524] ));
 sg13g2_inv_2 \inv[525]/_0_  (.Y(\inv_in[526] ),
    .A(\inv_in[525] ));
 sg13g2_inv_2 \inv[526]/_0_  (.Y(\inv_in[527] ),
    .A(\inv_in[526] ));
 sg13g2_inv_2 \inv[527]/_0_  (.Y(\inv_in[528] ),
    .A(\inv_in[527] ));
 sg13g2_inv_2 \inv[528]/_0_  (.Y(\inv_in[529] ),
    .A(\inv_in[528] ));
 sg13g2_inv_2 \inv[529]/_0_  (.Y(\inv_in[530] ),
    .A(\inv_in[529] ));
 sg13g2_inv_2 \inv[52]/_0_  (.Y(\inv_in[53] ),
    .A(\inv_in[52] ));
 sg13g2_inv_2 \inv[530]/_0_  (.Y(\inv_in[531] ),
    .A(\inv_in[530] ));
 sg13g2_inv_2 \inv[531]/_0_  (.Y(\inv_in[532] ),
    .A(\inv_in[531] ));
 sg13g2_inv_2 \inv[532]/_0_  (.Y(\inv_in[533] ),
    .A(\inv_in[532] ));
 sg13g2_inv_2 \inv[533]/_0_  (.Y(\inv_in[534] ),
    .A(\inv_in[533] ));
 sg13g2_inv_2 \inv[534]/_0_  (.Y(\inv_in[535] ),
    .A(\inv_in[534] ));
 sg13g2_inv_2 \inv[535]/_0_  (.Y(\inv_in[536] ),
    .A(\inv_in[535] ));
 sg13g2_inv_2 \inv[536]/_0_  (.Y(\inv_in[537] ),
    .A(\inv_in[536] ));
 sg13g2_inv_2 \inv[537]/_0_  (.Y(\inv_in[538] ),
    .A(\inv_in[537] ));
 sg13g2_inv_2 \inv[538]/_0_  (.Y(\inv_in[539] ),
    .A(\inv_in[538] ));
 sg13g2_inv_2 \inv[539]/_0_  (.Y(\inv_in[540] ),
    .A(\inv_in[539] ));
 sg13g2_inv_2 \inv[53]/_0_  (.Y(\inv_in[54] ),
    .A(\inv_in[53] ));
 sg13g2_inv_2 \inv[540]/_0_  (.Y(\inv_in[541] ),
    .A(\inv_in[540] ));
 sg13g2_inv_2 \inv[541]/_0_  (.Y(\inv_in[542] ),
    .A(\inv_in[541] ));
 sg13g2_inv_2 \inv[542]/_0_  (.Y(\inv_in[543] ),
    .A(\inv_in[542] ));
 sg13g2_inv_2 \inv[543]/_0_  (.Y(\inv_in[544] ),
    .A(\inv_in[543] ));
 sg13g2_inv_2 \inv[544]/_0_  (.Y(\inv_in[545] ),
    .A(\inv_in[544] ));
 sg13g2_inv_2 \inv[545]/_0_  (.Y(\inv_in[546] ),
    .A(\inv_in[545] ));
 sg13g2_inv_2 \inv[546]/_0_  (.Y(\inv_in[547] ),
    .A(\inv_in[546] ));
 sg13g2_inv_2 \inv[547]/_0_  (.Y(\inv_in[548] ),
    .A(\inv_in[547] ));
 sg13g2_inv_2 \inv[548]/_0_  (.Y(\inv_in[549] ),
    .A(\inv_in[548] ));
 sg13g2_inv_2 \inv[549]/_0_  (.Y(\inv_in[550] ),
    .A(\inv_in[549] ));
 sg13g2_inv_2 \inv[54]/_0_  (.Y(\inv_in[55] ),
    .A(\inv_in[54] ));
 sg13g2_inv_2 \inv[550]/_0_  (.Y(\inv_in[551] ),
    .A(\inv_in[550] ));
 sg13g2_inv_2 \inv[551]/_0_  (.Y(\inv_in[552] ),
    .A(\inv_in[551] ));
 sg13g2_inv_2 \inv[552]/_0_  (.Y(\inv_in[553] ),
    .A(\inv_in[552] ));
 sg13g2_inv_2 \inv[553]/_0_  (.Y(\inv_in[554] ),
    .A(\inv_in[553] ));
 sg13g2_inv_2 \inv[554]/_0_  (.Y(\inv_in[555] ),
    .A(\inv_in[554] ));
 sg13g2_inv_2 \inv[555]/_0_  (.Y(\inv_in[556] ),
    .A(\inv_in[555] ));
 sg13g2_inv_2 \inv[556]/_0_  (.Y(\inv_in[557] ),
    .A(\inv_in[556] ));
 sg13g2_inv_2 \inv[557]/_0_  (.Y(\inv_in[558] ),
    .A(\inv_in[557] ));
 sg13g2_inv_2 \inv[558]/_0_  (.Y(\inv_in[559] ),
    .A(\inv_in[558] ));
 sg13g2_inv_2 \inv[559]/_0_  (.Y(\inv_in[560] ),
    .A(\inv_in[559] ));
 sg13g2_inv_2 \inv[55]/_0_  (.Y(\inv_in[56] ),
    .A(\inv_in[55] ));
 sg13g2_inv_2 \inv[560]/_0_  (.Y(\inv_in[561] ),
    .A(\inv_in[560] ));
 sg13g2_inv_2 \inv[561]/_0_  (.Y(\inv_in[562] ),
    .A(\inv_in[561] ));
 sg13g2_inv_2 \inv[562]/_0_  (.Y(\inv_in[563] ),
    .A(\inv_in[562] ));
 sg13g2_inv_2 \inv[563]/_0_  (.Y(\inv_in[564] ),
    .A(\inv_in[563] ));
 sg13g2_inv_2 \inv[564]/_0_  (.Y(\inv_in[565] ),
    .A(\inv_in[564] ));
 sg13g2_inv_2 \inv[565]/_0_  (.Y(\inv_in[566] ),
    .A(\inv_in[565] ));
 sg13g2_inv_2 \inv[566]/_0_  (.Y(\inv_in[567] ),
    .A(\inv_in[566] ));
 sg13g2_inv_2 \inv[567]/_0_  (.Y(\inv_in[568] ),
    .A(\inv_in[567] ));
 sg13g2_inv_2 \inv[568]/_0_  (.Y(\inv_in[569] ),
    .A(\inv_in[568] ));
 sg13g2_inv_2 \inv[569]/_0_  (.Y(\inv_in[570] ),
    .A(\inv_in[569] ));
 sg13g2_inv_2 \inv[56]/_0_  (.Y(\inv_in[57] ),
    .A(\inv_in[56] ));
 sg13g2_inv_2 \inv[570]/_0_  (.Y(\inv_in[571] ),
    .A(\inv_in[570] ));
 sg13g2_inv_2 \inv[571]/_0_  (.Y(\inv_in[572] ),
    .A(\inv_in[571] ));
 sg13g2_inv_2 \inv[572]/_0_  (.Y(\inv_in[573] ),
    .A(\inv_in[572] ));
 sg13g2_inv_2 \inv[573]/_0_  (.Y(\inv_in[574] ),
    .A(\inv_in[573] ));
 sg13g2_inv_2 \inv[574]/_0_  (.Y(\inv_in[575] ),
    .A(\inv_in[574] ));
 sg13g2_inv_2 \inv[575]/_0_  (.Y(\inv_in[576] ),
    .A(\inv_in[575] ));
 sg13g2_inv_2 \inv[576]/_0_  (.Y(\inv_in[577] ),
    .A(\inv_in[576] ));
 sg13g2_inv_2 \inv[577]/_0_  (.Y(\inv_in[578] ),
    .A(\inv_in[577] ));
 sg13g2_inv_2 \inv[578]/_0_  (.Y(\inv_in[579] ),
    .A(\inv_in[578] ));
 sg13g2_inv_2 \inv[579]/_0_  (.Y(\inv_in[580] ),
    .A(\inv_in[579] ));
 sg13g2_inv_2 \inv[57]/_0_  (.Y(\inv_in[58] ),
    .A(\inv_in[57] ));
 sg13g2_inv_2 \inv[580]/_0_  (.Y(\inv_in[581] ),
    .A(\inv_in[580] ));
 sg13g2_inv_2 \inv[581]/_0_  (.Y(\inv_in[582] ),
    .A(\inv_in[581] ));
 sg13g2_inv_2 \inv[582]/_0_  (.Y(\inv_in[583] ),
    .A(\inv_in[582] ));
 sg13g2_inv_2 \inv[583]/_0_  (.Y(\inv_in[584] ),
    .A(\inv_in[583] ));
 sg13g2_inv_2 \inv[584]/_0_  (.Y(\inv_in[585] ),
    .A(\inv_in[584] ));
 sg13g2_inv_2 \inv[585]/_0_  (.Y(\inv_in[586] ),
    .A(\inv_in[585] ));
 sg13g2_inv_2 \inv[586]/_0_  (.Y(\inv_in[587] ),
    .A(\inv_in[586] ));
 sg13g2_inv_2 \inv[587]/_0_  (.Y(\inv_in[588] ),
    .A(\inv_in[587] ));
 sg13g2_inv_2 \inv[588]/_0_  (.Y(\inv_in[589] ),
    .A(\inv_in[588] ));
 sg13g2_inv_2 \inv[589]/_0_  (.Y(\inv_in[590] ),
    .A(\inv_in[589] ));
 sg13g2_inv_2 \inv[58]/_0_  (.Y(\inv_in[59] ),
    .A(\inv_in[58] ));
 sg13g2_inv_2 \inv[590]/_0_  (.Y(\inv_in[591] ),
    .A(\inv_in[590] ));
 sg13g2_inv_2 \inv[591]/_0_  (.Y(\inv_in[592] ),
    .A(\inv_in[591] ));
 sg13g2_inv_2 \inv[592]/_0_  (.Y(\inv_in[593] ),
    .A(\inv_in[592] ));
 sg13g2_inv_2 \inv[593]/_0_  (.Y(\inv_in[594] ),
    .A(\inv_in[593] ));
 sg13g2_inv_2 \inv[594]/_0_  (.Y(\inv_in[595] ),
    .A(\inv_in[594] ));
 sg13g2_inv_2 \inv[595]/_0_  (.Y(\inv_in[596] ),
    .A(\inv_in[595] ));
 sg13g2_inv_2 \inv[596]/_0_  (.Y(\inv_in[597] ),
    .A(\inv_in[596] ));
 sg13g2_inv_2 \inv[597]/_0_  (.Y(\inv_in[598] ),
    .A(\inv_in[597] ));
 sg13g2_inv_2 \inv[598]/_0_  (.Y(\inv_in[599] ),
    .A(\inv_in[598] ));
 sg13g2_inv_2 \inv[599]/_0_  (.Y(\inv_in[600] ),
    .A(\inv_in[599] ));
 sg13g2_inv_2 \inv[59]/_0_  (.Y(\inv_in[60] ),
    .A(\inv_in[59] ));
 sg13g2_inv_2 \inv[5]/_0_  (.Y(\inv_in[6] ),
    .A(\inv_in[5] ));
 sg13g2_inv_2 \inv[600]/_0_  (.Y(\inv_in[601] ),
    .A(\inv_in[600] ));
 sg13g2_inv_2 \inv[601]/_0_  (.Y(\inv_in[602] ),
    .A(\inv_in[601] ));
 sg13g2_inv_2 \inv[602]/_0_  (.Y(\inv_in[603] ),
    .A(\inv_in[602] ));
 sg13g2_inv_2 \inv[603]/_0_  (.Y(\inv_in[604] ),
    .A(\inv_in[603] ));
 sg13g2_inv_2 \inv[604]/_0_  (.Y(\inv_in[605] ),
    .A(\inv_in[604] ));
 sg13g2_inv_2 \inv[605]/_0_  (.Y(\inv_in[606] ),
    .A(\inv_in[605] ));
 sg13g2_inv_2 \inv[606]/_0_  (.Y(\inv_in[607] ),
    .A(\inv_in[606] ));
 sg13g2_inv_2 \inv[607]/_0_  (.Y(\inv_in[608] ),
    .A(\inv_in[607] ));
 sg13g2_inv_2 \inv[608]/_0_  (.Y(\inv_in[609] ),
    .A(\inv_in[608] ));
 sg13g2_inv_2 \inv[609]/_0_  (.Y(\inv_in[610] ),
    .A(\inv_in[609] ));
 sg13g2_inv_2 \inv[60]/_0_  (.Y(\inv_in[61] ),
    .A(\inv_in[60] ));
 sg13g2_inv_2 \inv[610]/_0_  (.Y(\inv_in[611] ),
    .A(\inv_in[610] ));
 sg13g2_inv_2 \inv[611]/_0_  (.Y(\inv_in[612] ),
    .A(\inv_in[611] ));
 sg13g2_inv_2 \inv[612]/_0_  (.Y(\inv_in[613] ),
    .A(\inv_in[612] ));
 sg13g2_inv_2 \inv[613]/_0_  (.Y(\inv_in[614] ),
    .A(\inv_in[613] ));
 sg13g2_inv_2 \inv[614]/_0_  (.Y(\inv_in[615] ),
    .A(\inv_in[614] ));
 sg13g2_inv_2 \inv[615]/_0_  (.Y(\inv_in[616] ),
    .A(\inv_in[615] ));
 sg13g2_inv_2 \inv[616]/_0_  (.Y(\inv_in[617] ),
    .A(\inv_in[616] ));
 sg13g2_inv_2 \inv[617]/_0_  (.Y(\inv_in[618] ),
    .A(\inv_in[617] ));
 sg13g2_inv_2 \inv[618]/_0_  (.Y(\inv_in[619] ),
    .A(\inv_in[618] ));
 sg13g2_inv_2 \inv[619]/_0_  (.Y(\inv_in[620] ),
    .A(\inv_in[619] ));
 sg13g2_inv_2 \inv[61]/_0_  (.Y(\inv_in[62] ),
    .A(\inv_in[61] ));
 sg13g2_inv_2 \inv[620]/_0_  (.Y(\inv_in[621] ),
    .A(\inv_in[620] ));
 sg13g2_inv_2 \inv[621]/_0_  (.Y(\inv_in[622] ),
    .A(\inv_in[621] ));
 sg13g2_inv_2 \inv[622]/_0_  (.Y(\inv_in[623] ),
    .A(\inv_in[622] ));
 sg13g2_inv_2 \inv[623]/_0_  (.Y(\inv_in[624] ),
    .A(\inv_in[623] ));
 sg13g2_inv_2 \inv[624]/_0_  (.Y(\inv_in[625] ),
    .A(\inv_in[624] ));
 sg13g2_inv_2 \inv[625]/_0_  (.Y(\inv_in[626] ),
    .A(\inv_in[625] ));
 sg13g2_inv_2 \inv[626]/_0_  (.Y(\inv_in[627] ),
    .A(\inv_in[626] ));
 sg13g2_inv_2 \inv[627]/_0_  (.Y(\inv_in[628] ),
    .A(\inv_in[627] ));
 sg13g2_inv_2 \inv[628]/_0_  (.Y(\inv_in[629] ),
    .A(\inv_in[628] ));
 sg13g2_inv_2 \inv[629]/_0_  (.Y(\inv_in[630] ),
    .A(\inv_in[629] ));
 sg13g2_inv_2 \inv[62]/_0_  (.Y(\inv_in[63] ),
    .A(\inv_in[62] ));
 sg13g2_inv_2 \inv[630]/_0_  (.Y(\inv_in[631] ),
    .A(\inv_in[630] ));
 sg13g2_inv_2 \inv[631]/_0_  (.Y(\inv_in[632] ),
    .A(\inv_in[631] ));
 sg13g2_inv_2 \inv[632]/_0_  (.Y(\inv_in[633] ),
    .A(\inv_in[632] ));
 sg13g2_inv_2 \inv[633]/_0_  (.Y(\inv_in[634] ),
    .A(\inv_in[633] ));
 sg13g2_inv_2 \inv[634]/_0_  (.Y(\inv_in[635] ),
    .A(\inv_in[634] ));
 sg13g2_inv_2 \inv[635]/_0_  (.Y(\inv_in[636] ),
    .A(\inv_in[635] ));
 sg13g2_inv_2 \inv[636]/_0_  (.Y(\inv_in[637] ),
    .A(\inv_in[636] ));
 sg13g2_inv_2 \inv[637]/_0_  (.Y(\inv_in[638] ),
    .A(\inv_in[637] ));
 sg13g2_inv_2 \inv[638]/_0_  (.Y(\inv_in[639] ),
    .A(\inv_in[638] ));
 sg13g2_inv_2 \inv[639]/_0_  (.Y(\inv_in[640] ),
    .A(\inv_in[639] ));
 sg13g2_inv_2 \inv[63]/_0_  (.Y(\inv_in[64] ),
    .A(\inv_in[63] ));
 sg13g2_inv_2 \inv[640]/_0_  (.Y(\inv_in[641] ),
    .A(\inv_in[640] ));
 sg13g2_inv_2 \inv[641]/_0_  (.Y(\inv_in[642] ),
    .A(\inv_in[641] ));
 sg13g2_inv_2 \inv[642]/_0_  (.Y(\inv_in[643] ),
    .A(\inv_in[642] ));
 sg13g2_inv_2 \inv[643]/_0_  (.Y(\inv_in[644] ),
    .A(\inv_in[643] ));
 sg13g2_inv_2 \inv[644]/_0_  (.Y(\inv_in[645] ),
    .A(\inv_in[644] ));
 sg13g2_inv_2 \inv[645]/_0_  (.Y(\inv_in[646] ),
    .A(\inv_in[645] ));
 sg13g2_inv_2 \inv[646]/_0_  (.Y(\inv_in[647] ),
    .A(\inv_in[646] ));
 sg13g2_inv_2 \inv[647]/_0_  (.Y(\inv_in[648] ),
    .A(\inv_in[647] ));
 sg13g2_inv_2 \inv[648]/_0_  (.Y(\inv_in[649] ),
    .A(\inv_in[648] ));
 sg13g2_inv_2 \inv[649]/_0_  (.Y(\inv_in[650] ),
    .A(\inv_in[649] ));
 sg13g2_inv_2 \inv[64]/_0_  (.Y(\inv_in[65] ),
    .A(\inv_in[64] ));
 sg13g2_inv_2 \inv[650]/_0_  (.Y(\inv_in[651] ),
    .A(\inv_in[650] ));
 sg13g2_inv_2 \inv[651]/_0_  (.Y(\inv_in[652] ),
    .A(\inv_in[651] ));
 sg13g2_inv_2 \inv[652]/_0_  (.Y(\inv_in[653] ),
    .A(\inv_in[652] ));
 sg13g2_inv_2 \inv[653]/_0_  (.Y(\inv_in[654] ),
    .A(\inv_in[653] ));
 sg13g2_inv_2 \inv[654]/_0_  (.Y(\inv_in[655] ),
    .A(\inv_in[654] ));
 sg13g2_inv_2 \inv[655]/_0_  (.Y(\inv_in[656] ),
    .A(\inv_in[655] ));
 sg13g2_inv_2 \inv[656]/_0_  (.Y(\inv_in[657] ),
    .A(\inv_in[656] ));
 sg13g2_inv_2 \inv[657]/_0_  (.Y(\inv_in[658] ),
    .A(\inv_in[657] ));
 sg13g2_inv_2 \inv[658]/_0_  (.Y(\inv_in[659] ),
    .A(\inv_in[658] ));
 sg13g2_inv_2 \inv[659]/_0_  (.Y(\inv_in[660] ),
    .A(\inv_in[659] ));
 sg13g2_inv_2 \inv[65]/_0_  (.Y(\inv_in[66] ),
    .A(\inv_in[65] ));
 sg13g2_inv_2 \inv[660]/_0_  (.Y(\inv_in[661] ),
    .A(\inv_in[660] ));
 sg13g2_inv_2 \inv[661]/_0_  (.Y(\inv_in[662] ),
    .A(\inv_in[661] ));
 sg13g2_inv_2 \inv[662]/_0_  (.Y(\inv_in[663] ),
    .A(\inv_in[662] ));
 sg13g2_inv_2 \inv[663]/_0_  (.Y(\inv_in[664] ),
    .A(\inv_in[663] ));
 sg13g2_inv_2 \inv[664]/_0_  (.Y(\inv_in[665] ),
    .A(\inv_in[664] ));
 sg13g2_inv_2 \inv[665]/_0_  (.Y(\inv_in[666] ),
    .A(\inv_in[665] ));
 sg13g2_inv_2 \inv[666]/_0_  (.Y(\inv_in[667] ),
    .A(\inv_in[666] ));
 sg13g2_inv_2 \inv[667]/_0_  (.Y(\inv_in[668] ),
    .A(\inv_in[667] ));
 sg13g2_inv_2 \inv[668]/_0_  (.Y(\inv_in[669] ),
    .A(\inv_in[668] ));
 sg13g2_inv_2 \inv[669]/_0_  (.Y(\inv_in[670] ),
    .A(\inv_in[669] ));
 sg13g2_inv_2 \inv[66]/_0_  (.Y(\inv_in[67] ),
    .A(\inv_in[66] ));
 sg13g2_inv_2 \inv[670]/_0_  (.Y(\inv_in[671] ),
    .A(\inv_in[670] ));
 sg13g2_inv_2 \inv[671]/_0_  (.Y(\inv_in[672] ),
    .A(\inv_in[671] ));
 sg13g2_inv_2 \inv[672]/_0_  (.Y(\inv_in[673] ),
    .A(\inv_in[672] ));
 sg13g2_inv_2 \inv[673]/_0_  (.Y(\inv_in[674] ),
    .A(\inv_in[673] ));
 sg13g2_inv_2 \inv[674]/_0_  (.Y(\inv_in[675] ),
    .A(\inv_in[674] ));
 sg13g2_inv_2 \inv[675]/_0_  (.Y(\inv_in[676] ),
    .A(\inv_in[675] ));
 sg13g2_inv_2 \inv[676]/_0_  (.Y(\inv_in[677] ),
    .A(\inv_in[676] ));
 sg13g2_inv_2 \inv[677]/_0_  (.Y(\inv_in[678] ),
    .A(\inv_in[677] ));
 sg13g2_inv_2 \inv[678]/_0_  (.Y(\inv_in[679] ),
    .A(\inv_in[678] ));
 sg13g2_inv_2 \inv[679]/_0_  (.Y(\inv_in[680] ),
    .A(\inv_in[679] ));
 sg13g2_inv_2 \inv[67]/_0_  (.Y(\inv_in[68] ),
    .A(\inv_in[67] ));
 sg13g2_inv_2 \inv[680]/_0_  (.Y(\inv_in[681] ),
    .A(\inv_in[680] ));
 sg13g2_inv_2 \inv[681]/_0_  (.Y(\inv_in[682] ),
    .A(\inv_in[681] ));
 sg13g2_inv_2 \inv[682]/_0_  (.Y(\inv_in[683] ),
    .A(\inv_in[682] ));
 sg13g2_inv_2 \inv[683]/_0_  (.Y(\inv_in[684] ),
    .A(\inv_in[683] ));
 sg13g2_inv_2 \inv[684]/_0_  (.Y(\inv_in[685] ),
    .A(\inv_in[684] ));
 sg13g2_inv_2 \inv[685]/_0_  (.Y(\inv_in[686] ),
    .A(\inv_in[685] ));
 sg13g2_inv_2 \inv[686]/_0_  (.Y(\inv_in[687] ),
    .A(\inv_in[686] ));
 sg13g2_inv_2 \inv[687]/_0_  (.Y(\inv_in[688] ),
    .A(\inv_in[687] ));
 sg13g2_inv_2 \inv[688]/_0_  (.Y(\inv_in[689] ),
    .A(\inv_in[688] ));
 sg13g2_inv_2 \inv[689]/_0_  (.Y(\inv_in[690] ),
    .A(\inv_in[689] ));
 sg13g2_inv_2 \inv[68]/_0_  (.Y(\inv_in[69] ),
    .A(\inv_in[68] ));
 sg13g2_inv_2 \inv[690]/_0_  (.Y(\inv_in[691] ),
    .A(\inv_in[690] ));
 sg13g2_inv_2 \inv[691]/_0_  (.Y(\inv_in[692] ),
    .A(\inv_in[691] ));
 sg13g2_inv_2 \inv[692]/_0_  (.Y(\inv_in[693] ),
    .A(\inv_in[692] ));
 sg13g2_inv_2 \inv[693]/_0_  (.Y(\inv_in[694] ),
    .A(\inv_in[693] ));
 sg13g2_inv_2 \inv[694]/_0_  (.Y(\inv_in[695] ),
    .A(\inv_in[694] ));
 sg13g2_inv_2 \inv[695]/_0_  (.Y(\inv_in[696] ),
    .A(\inv_in[695] ));
 sg13g2_inv_2 \inv[696]/_0_  (.Y(\inv_in[697] ),
    .A(\inv_in[696] ));
 sg13g2_inv_2 \inv[697]/_0_  (.Y(\inv_in[698] ),
    .A(\inv_in[697] ));
 sg13g2_inv_2 \inv[698]/_0_  (.Y(\inv_in[699] ),
    .A(\inv_in[698] ));
 sg13g2_inv_2 \inv[699]/_0_  (.Y(\inv_in[700] ),
    .A(\inv_in[699] ));
 sg13g2_inv_2 \inv[69]/_0_  (.Y(\inv_in[70] ),
    .A(\inv_in[69] ));
 sg13g2_inv_2 \inv[6]/_0_  (.Y(\inv_in[7] ),
    .A(\inv_in[6] ));
 sg13g2_inv_2 \inv[700]/_0_  (.Y(\inv_in[701] ),
    .A(\inv_in[700] ));
 sg13g2_inv_2 \inv[701]/_0_  (.Y(\inv_in[702] ),
    .A(\inv_in[701] ));
 sg13g2_inv_2 \inv[702]/_0_  (.Y(\inv_in[703] ),
    .A(\inv_in[702] ));
 sg13g2_inv_2 \inv[703]/_0_  (.Y(\inv_in[704] ),
    .A(\inv_in[703] ));
 sg13g2_inv_2 \inv[704]/_0_  (.Y(\inv_in[705] ),
    .A(\inv_in[704] ));
 sg13g2_inv_2 \inv[705]/_0_  (.Y(\inv_in[706] ),
    .A(\inv_in[705] ));
 sg13g2_inv_2 \inv[706]/_0_  (.Y(\inv_in[707] ),
    .A(\inv_in[706] ));
 sg13g2_inv_2 \inv[707]/_0_  (.Y(\inv_in[708] ),
    .A(\inv_in[707] ));
 sg13g2_inv_2 \inv[708]/_0_  (.Y(\inv_in[709] ),
    .A(\inv_in[708] ));
 sg13g2_inv_2 \inv[709]/_0_  (.Y(\inv_in[710] ),
    .A(\inv_in[709] ));
 sg13g2_inv_2 \inv[70]/_0_  (.Y(\inv_in[71] ),
    .A(\inv_in[70] ));
 sg13g2_inv_2 \inv[710]/_0_  (.Y(\inv_in[711] ),
    .A(\inv_in[710] ));
 sg13g2_inv_2 \inv[711]/_0_  (.Y(\inv_in[712] ),
    .A(\inv_in[711] ));
 sg13g2_inv_2 \inv[712]/_0_  (.Y(\inv_in[713] ),
    .A(\inv_in[712] ));
 sg13g2_inv_2 \inv[713]/_0_  (.Y(\inv_in[714] ),
    .A(\inv_in[713] ));
 sg13g2_inv_2 \inv[714]/_0_  (.Y(\inv_in[715] ),
    .A(\inv_in[714] ));
 sg13g2_inv_2 \inv[715]/_0_  (.Y(\inv_in[716] ),
    .A(\inv_in[715] ));
 sg13g2_inv_2 \inv[716]/_0_  (.Y(\inv_in[717] ),
    .A(\inv_in[716] ));
 sg13g2_inv_2 \inv[717]/_0_  (.Y(\inv_in[718] ),
    .A(\inv_in[717] ));
 sg13g2_inv_2 \inv[718]/_0_  (.Y(\inv_in[719] ),
    .A(\inv_in[718] ));
 sg13g2_inv_2 \inv[719]/_0_  (.Y(\inv_in[720] ),
    .A(\inv_in[719] ));
 sg13g2_inv_2 \inv[71]/_0_  (.Y(\inv_in[72] ),
    .A(\inv_in[71] ));
 sg13g2_inv_2 \inv[720]/_0_  (.Y(\inv_in[721] ),
    .A(\inv_in[720] ));
 sg13g2_inv_2 \inv[721]/_0_  (.Y(\inv_in[722] ),
    .A(\inv_in[721] ));
 sg13g2_inv_2 \inv[722]/_0_  (.Y(\inv_in[723] ),
    .A(\inv_in[722] ));
 sg13g2_inv_2 \inv[723]/_0_  (.Y(\inv_in[724] ),
    .A(\inv_in[723] ));
 sg13g2_inv_2 \inv[724]/_0_  (.Y(\inv_in[725] ),
    .A(\inv_in[724] ));
 sg13g2_inv_2 \inv[725]/_0_  (.Y(\inv_in[726] ),
    .A(\inv_in[725] ));
 sg13g2_inv_2 \inv[726]/_0_  (.Y(\inv_in[727] ),
    .A(\inv_in[726] ));
 sg13g2_inv_2 \inv[727]/_0_  (.Y(\inv_in[728] ),
    .A(\inv_in[727] ));
 sg13g2_inv_2 \inv[728]/_0_  (.Y(\inv_in[729] ),
    .A(\inv_in[728] ));
 sg13g2_inv_2 \inv[729]/_0_  (.Y(\inv_in[730] ),
    .A(\inv_in[729] ));
 sg13g2_inv_2 \inv[72]/_0_  (.Y(\inv_in[73] ),
    .A(\inv_in[72] ));
 sg13g2_inv_2 \inv[730]/_0_  (.Y(\inv_in[731] ),
    .A(\inv_in[730] ));
 sg13g2_inv_2 \inv[731]/_0_  (.Y(\inv_in[732] ),
    .A(\inv_in[731] ));
 sg13g2_inv_2 \inv[732]/_0_  (.Y(\inv_in[733] ),
    .A(\inv_in[732] ));
 sg13g2_inv_2 \inv[733]/_0_  (.Y(\inv_in[734] ),
    .A(\inv_in[733] ));
 sg13g2_inv_2 \inv[734]/_0_  (.Y(\inv_in[735] ),
    .A(\inv_in[734] ));
 sg13g2_inv_2 \inv[735]/_0_  (.Y(\inv_in[736] ),
    .A(\inv_in[735] ));
 sg13g2_inv_2 \inv[736]/_0_  (.Y(\inv_in[737] ),
    .A(\inv_in[736] ));
 sg13g2_inv_2 \inv[737]/_0_  (.Y(\inv_in[738] ),
    .A(\inv_in[737] ));
 sg13g2_inv_2 \inv[738]/_0_  (.Y(\inv_in[739] ),
    .A(\inv_in[738] ));
 sg13g2_inv_2 \inv[739]/_0_  (.Y(\inv_in[740] ),
    .A(\inv_in[739] ));
 sg13g2_inv_2 \inv[73]/_0_  (.Y(\inv_in[74] ),
    .A(\inv_in[73] ));
 sg13g2_inv_2 \inv[740]/_0_  (.Y(\inv_in[741] ),
    .A(\inv_in[740] ));
 sg13g2_inv_2 \inv[741]/_0_  (.Y(\inv_in[742] ),
    .A(\inv_in[741] ));
 sg13g2_inv_2 \inv[742]/_0_  (.Y(\inv_in[743] ),
    .A(\inv_in[742] ));
 sg13g2_inv_2 \inv[743]/_0_  (.Y(\inv_in[744] ),
    .A(\inv_in[743] ));
 sg13g2_inv_2 \inv[744]/_0_  (.Y(\inv_in[745] ),
    .A(\inv_in[744] ));
 sg13g2_inv_2 \inv[745]/_0_  (.Y(\inv_in[746] ),
    .A(\inv_in[745] ));
 sg13g2_inv_2 \inv[746]/_0_  (.Y(\inv_in[747] ),
    .A(\inv_in[746] ));
 sg13g2_inv_2 \inv[747]/_0_  (.Y(\inv_in[748] ),
    .A(\inv_in[747] ));
 sg13g2_inv_2 \inv[748]/_0_  (.Y(\inv_in[749] ),
    .A(\inv_in[748] ));
 sg13g2_inv_2 \inv[749]/_0_  (.Y(\inv_in[750] ),
    .A(\inv_in[749] ));
 sg13g2_inv_2 \inv[74]/_0_  (.Y(\inv_in[75] ),
    .A(\inv_in[74] ));
 sg13g2_inv_2 \inv[750]/_0_  (.Y(\inv_in[751] ),
    .A(\inv_in[750] ));
 sg13g2_inv_2 \inv[751]/_0_  (.Y(\inv_in[752] ),
    .A(\inv_in[751] ));
 sg13g2_inv_2 \inv[752]/_0_  (.Y(\inv_in[753] ),
    .A(\inv_in[752] ));
 sg13g2_inv_2 \inv[753]/_0_  (.Y(\inv_in[754] ),
    .A(\inv_in[753] ));
 sg13g2_inv_2 \inv[754]/_0_  (.Y(\inv_in[755] ),
    .A(\inv_in[754] ));
 sg13g2_inv_2 \inv[755]/_0_  (.Y(\inv_in[756] ),
    .A(\inv_in[755] ));
 sg13g2_inv_2 \inv[756]/_0_  (.Y(\inv_in[757] ),
    .A(\inv_in[756] ));
 sg13g2_inv_2 \inv[757]/_0_  (.Y(\inv_in[758] ),
    .A(\inv_in[757] ));
 sg13g2_inv_2 \inv[758]/_0_  (.Y(\inv_in[759] ),
    .A(\inv_in[758] ));
 sg13g2_inv_2 \inv[759]/_0_  (.Y(\inv_in[760] ),
    .A(\inv_in[759] ));
 sg13g2_inv_2 \inv[75]/_0_  (.Y(\inv_in[76] ),
    .A(\inv_in[75] ));
 sg13g2_inv_2 \inv[760]/_0_  (.Y(\inv_in[761] ),
    .A(\inv_in[760] ));
 sg13g2_inv_2 \inv[761]/_0_  (.Y(\inv_in[762] ),
    .A(\inv_in[761] ));
 sg13g2_inv_2 \inv[762]/_0_  (.Y(\inv_in[763] ),
    .A(\inv_in[762] ));
 sg13g2_inv_2 \inv[763]/_0_  (.Y(\inv_in[764] ),
    .A(\inv_in[763] ));
 sg13g2_inv_2 \inv[764]/_0_  (.Y(\inv_in[765] ),
    .A(\inv_in[764] ));
 sg13g2_inv_2 \inv[765]/_0_  (.Y(\inv_in[766] ),
    .A(\inv_in[765] ));
 sg13g2_inv_2 \inv[766]/_0_  (.Y(\inv_in[767] ),
    .A(\inv_in[766] ));
 sg13g2_inv_2 \inv[767]/_0_  (.Y(\inv_in[768] ),
    .A(\inv_in[767] ));
 sg13g2_inv_2 \inv[768]/_0_  (.Y(\inv_in[769] ),
    .A(\inv_in[768] ));
 sg13g2_inv_2 \inv[769]/_0_  (.Y(\inv_in[770] ),
    .A(\inv_in[769] ));
 sg13g2_inv_2 \inv[76]/_0_  (.Y(\inv_in[77] ),
    .A(\inv_in[76] ));
 sg13g2_inv_2 \inv[770]/_0_  (.Y(\inv_in[771] ),
    .A(\inv_in[770] ));
 sg13g2_inv_2 \inv[771]/_0_  (.Y(\inv_in[772] ),
    .A(\inv_in[771] ));
 sg13g2_inv_2 \inv[772]/_0_  (.Y(\inv_in[773] ),
    .A(\inv_in[772] ));
 sg13g2_inv_2 \inv[773]/_0_  (.Y(\inv_in[774] ),
    .A(\inv_in[773] ));
 sg13g2_inv_2 \inv[774]/_0_  (.Y(\inv_in[775] ),
    .A(\inv_in[774] ));
 sg13g2_inv_2 \inv[775]/_0_  (.Y(\inv_in[776] ),
    .A(\inv_in[775] ));
 sg13g2_inv_2 \inv[776]/_0_  (.Y(\inv_in[777] ),
    .A(\inv_in[776] ));
 sg13g2_inv_2 \inv[777]/_0_  (.Y(\inv_in[778] ),
    .A(\inv_in[777] ));
 sg13g2_inv_2 \inv[778]/_0_  (.Y(\inv_in[779] ),
    .A(\inv_in[778] ));
 sg13g2_inv_2 \inv[779]/_0_  (.Y(\inv_in[780] ),
    .A(\inv_in[779] ));
 sg13g2_inv_2 \inv[77]/_0_  (.Y(\inv_in[78] ),
    .A(\inv_in[77] ));
 sg13g2_inv_2 \inv[780]/_0_  (.Y(\inv_in[781] ),
    .A(\inv_in[780] ));
 sg13g2_inv_2 \inv[781]/_0_  (.Y(\inv_in[782] ),
    .A(\inv_in[781] ));
 sg13g2_inv_2 \inv[782]/_0_  (.Y(\inv_in[783] ),
    .A(\inv_in[782] ));
 sg13g2_inv_2 \inv[783]/_0_  (.Y(\inv_in[784] ),
    .A(\inv_in[783] ));
 sg13g2_inv_2 \inv[784]/_0_  (.Y(\inv_in[785] ),
    .A(\inv_in[784] ));
 sg13g2_inv_2 \inv[785]/_0_  (.Y(\inv_in[786] ),
    .A(\inv_in[785] ));
 sg13g2_inv_2 \inv[786]/_0_  (.Y(\inv_in[787] ),
    .A(\inv_in[786] ));
 sg13g2_inv_2 \inv[787]/_0_  (.Y(\inv_in[788] ),
    .A(\inv_in[787] ));
 sg13g2_inv_2 \inv[788]/_0_  (.Y(\inv_in[789] ),
    .A(\inv_in[788] ));
 sg13g2_inv_2 \inv[789]/_0_  (.Y(\inv_in[790] ),
    .A(\inv_in[789] ));
 sg13g2_inv_2 \inv[78]/_0_  (.Y(\inv_in[79] ),
    .A(\inv_in[78] ));
 sg13g2_inv_2 \inv[790]/_0_  (.Y(\inv_in[791] ),
    .A(\inv_in[790] ));
 sg13g2_inv_2 \inv[791]/_0_  (.Y(\inv_in[792] ),
    .A(\inv_in[791] ));
 sg13g2_inv_2 \inv[792]/_0_  (.Y(\inv_in[793] ),
    .A(\inv_in[792] ));
 sg13g2_inv_2 \inv[793]/_0_  (.Y(\inv_in[794] ),
    .A(\inv_in[793] ));
 sg13g2_inv_2 \inv[794]/_0_  (.Y(\inv_in[795] ),
    .A(\inv_in[794] ));
 sg13g2_inv_2 \inv[795]/_0_  (.Y(\inv_in[796] ),
    .A(\inv_in[795] ));
 sg13g2_inv_2 \inv[796]/_0_  (.Y(\inv_in[797] ),
    .A(\inv_in[796] ));
 sg13g2_inv_2 \inv[797]/_0_  (.Y(\inv_in[798] ),
    .A(\inv_in[797] ));
 sg13g2_inv_2 \inv[798]/_0_  (.Y(\inv_in[799] ),
    .A(\inv_in[798] ));
 sg13g2_inv_2 \inv[799]/_0_  (.Y(\inv_in[800] ),
    .A(\inv_in[799] ));
 sg13g2_inv_2 \inv[79]/_0_  (.Y(\inv_in[80] ),
    .A(\inv_in[79] ));
 sg13g2_inv_2 \inv[7]/_0_  (.Y(\inv_in[8] ),
    .A(\inv_in[7] ));
 sg13g2_inv_2 \inv[800]/_0_  (.Y(\inv_in[801] ),
    .A(\inv_in[800] ));
 sg13g2_inv_2 \inv[801]/_0_  (.Y(\inv_in[802] ),
    .A(\inv_in[801] ));
 sg13g2_inv_2 \inv[802]/_0_  (.Y(\inv_in[803] ),
    .A(\inv_in[802] ));
 sg13g2_inv_2 \inv[803]/_0_  (.Y(\inv_in[804] ),
    .A(\inv_in[803] ));
 sg13g2_inv_2 \inv[804]/_0_  (.Y(\inv_in[805] ),
    .A(\inv_in[804] ));
 sg13g2_inv_2 \inv[805]/_0_  (.Y(\inv_in[806] ),
    .A(\inv_in[805] ));
 sg13g2_inv_2 \inv[806]/_0_  (.Y(\inv_in[807] ),
    .A(\inv_in[806] ));
 sg13g2_inv_2 \inv[807]/_0_  (.Y(\inv_in[808] ),
    .A(\inv_in[807] ));
 sg13g2_inv_2 \inv[808]/_0_  (.Y(\inv_in[809] ),
    .A(\inv_in[808] ));
 sg13g2_inv_2 \inv[809]/_0_  (.Y(\inv_in[810] ),
    .A(\inv_in[809] ));
 sg13g2_inv_2 \inv[80]/_0_  (.Y(\inv_in[81] ),
    .A(\inv_in[80] ));
 sg13g2_inv_2 \inv[810]/_0_  (.Y(\inv_in[811] ),
    .A(\inv_in[810] ));
 sg13g2_inv_2 \inv[811]/_0_  (.Y(\inv_in[812] ),
    .A(\inv_in[811] ));
 sg13g2_inv_2 \inv[812]/_0_  (.Y(\inv_in[813] ),
    .A(\inv_in[812] ));
 sg13g2_inv_2 \inv[813]/_0_  (.Y(\inv_in[814] ),
    .A(\inv_in[813] ));
 sg13g2_inv_2 \inv[814]/_0_  (.Y(\inv_in[815] ),
    .A(\inv_in[814] ));
 sg13g2_inv_2 \inv[815]/_0_  (.Y(\inv_in[816] ),
    .A(\inv_in[815] ));
 sg13g2_inv_2 \inv[816]/_0_  (.Y(\inv_in[817] ),
    .A(\inv_in[816] ));
 sg13g2_inv_2 \inv[817]/_0_  (.Y(\inv_in[818] ),
    .A(\inv_in[817] ));
 sg13g2_inv_2 \inv[818]/_0_  (.Y(\inv_in[819] ),
    .A(\inv_in[818] ));
 sg13g2_inv_2 \inv[819]/_0_  (.Y(\inv_in[820] ),
    .A(\inv_in[819] ));
 sg13g2_inv_2 \inv[81]/_0_  (.Y(\inv_in[82] ),
    .A(\inv_in[81] ));
 sg13g2_inv_2 \inv[820]/_0_  (.Y(\inv_in[821] ),
    .A(\inv_in[820] ));
 sg13g2_inv_2 \inv[821]/_0_  (.Y(\inv_in[822] ),
    .A(\inv_in[821] ));
 sg13g2_inv_2 \inv[822]/_0_  (.Y(\inv_in[823] ),
    .A(\inv_in[822] ));
 sg13g2_inv_2 \inv[823]/_0_  (.Y(\inv_in[824] ),
    .A(\inv_in[823] ));
 sg13g2_inv_2 \inv[824]/_0_  (.Y(\inv_in[825] ),
    .A(\inv_in[824] ));
 sg13g2_inv_2 \inv[825]/_0_  (.Y(\inv_in[826] ),
    .A(\inv_in[825] ));
 sg13g2_inv_2 \inv[826]/_0_  (.Y(\inv_in[827] ),
    .A(\inv_in[826] ));
 sg13g2_inv_2 \inv[827]/_0_  (.Y(\inv_in[828] ),
    .A(\inv_in[827] ));
 sg13g2_inv_2 \inv[828]/_0_  (.Y(\inv_in[829] ),
    .A(\inv_in[828] ));
 sg13g2_inv_2 \inv[829]/_0_  (.Y(\inv_in[830] ),
    .A(\inv_in[829] ));
 sg13g2_inv_2 \inv[82]/_0_  (.Y(\inv_in[83] ),
    .A(\inv_in[82] ));
 sg13g2_inv_2 \inv[830]/_0_  (.Y(\inv_in[831] ),
    .A(\inv_in[830] ));
 sg13g2_inv_2 \inv[831]/_0_  (.Y(\inv_in[832] ),
    .A(\inv_in[831] ));
 sg13g2_inv_2 \inv[832]/_0_  (.Y(\inv_in[833] ),
    .A(\inv_in[832] ));
 sg13g2_inv_2 \inv[833]/_0_  (.Y(\inv_in[834] ),
    .A(\inv_in[833] ));
 sg13g2_inv_2 \inv[834]/_0_  (.Y(\inv_in[835] ),
    .A(\inv_in[834] ));
 sg13g2_inv_2 \inv[835]/_0_  (.Y(\inv_in[836] ),
    .A(\inv_in[835] ));
 sg13g2_inv_2 \inv[836]/_0_  (.Y(\inv_in[837] ),
    .A(\inv_in[836] ));
 sg13g2_inv_2 \inv[837]/_0_  (.Y(\inv_in[838] ),
    .A(\inv_in[837] ));
 sg13g2_inv_2 \inv[838]/_0_  (.Y(\inv_in[839] ),
    .A(\inv_in[838] ));
 sg13g2_inv_2 \inv[839]/_0_  (.Y(\inv_in[840] ),
    .A(\inv_in[839] ));
 sg13g2_inv_2 \inv[83]/_0_  (.Y(\inv_in[84] ),
    .A(\inv_in[83] ));
 sg13g2_inv_2 \inv[840]/_0_  (.Y(\inv_in[841] ),
    .A(\inv_in[840] ));
 sg13g2_inv_2 \inv[841]/_0_  (.Y(\inv_in[842] ),
    .A(\inv_in[841] ));
 sg13g2_inv_2 \inv[842]/_0_  (.Y(\inv_in[843] ),
    .A(\inv_in[842] ));
 sg13g2_inv_2 \inv[843]/_0_  (.Y(\inv_in[844] ),
    .A(\inv_in[843] ));
 sg13g2_inv_2 \inv[844]/_0_  (.Y(\inv_in[845] ),
    .A(\inv_in[844] ));
 sg13g2_inv_2 \inv[845]/_0_  (.Y(\inv_in[846] ),
    .A(\inv_in[845] ));
 sg13g2_inv_2 \inv[846]/_0_  (.Y(\inv_in[847] ),
    .A(\inv_in[846] ));
 sg13g2_inv_2 \inv[847]/_0_  (.Y(\inv_in[848] ),
    .A(\inv_in[847] ));
 sg13g2_inv_2 \inv[848]/_0_  (.Y(\inv_in[849] ),
    .A(\inv_in[848] ));
 sg13g2_inv_2 \inv[849]/_0_  (.Y(\inv_in[850] ),
    .A(\inv_in[849] ));
 sg13g2_inv_2 \inv[84]/_0_  (.Y(\inv_in[85] ),
    .A(\inv_in[84] ));
 sg13g2_inv_2 \inv[850]/_0_  (.Y(\inv_in[851] ),
    .A(\inv_in[850] ));
 sg13g2_inv_2 \inv[851]/_0_  (.Y(\inv_in[852] ),
    .A(\inv_in[851] ));
 sg13g2_inv_2 \inv[852]/_0_  (.Y(\inv_in[853] ),
    .A(\inv_in[852] ));
 sg13g2_inv_2 \inv[853]/_0_  (.Y(\inv_in[854] ),
    .A(\inv_in[853] ));
 sg13g2_inv_2 \inv[854]/_0_  (.Y(\inv_in[855] ),
    .A(\inv_in[854] ));
 sg13g2_inv_2 \inv[855]/_0_  (.Y(\inv_in[856] ),
    .A(\inv_in[855] ));
 sg13g2_inv_2 \inv[856]/_0_  (.Y(\inv_in[857] ),
    .A(\inv_in[856] ));
 sg13g2_inv_2 \inv[857]/_0_  (.Y(\inv_in[858] ),
    .A(\inv_in[857] ));
 sg13g2_inv_2 \inv[858]/_0_  (.Y(\inv_in[859] ),
    .A(\inv_in[858] ));
 sg13g2_inv_2 \inv[859]/_0_  (.Y(\inv_in[860] ),
    .A(\inv_in[859] ));
 sg13g2_inv_2 \inv[85]/_0_  (.Y(\inv_in[86] ),
    .A(\inv_in[85] ));
 sg13g2_inv_2 \inv[860]/_0_  (.Y(\inv_in[861] ),
    .A(\inv_in[860] ));
 sg13g2_inv_2 \inv[861]/_0_  (.Y(\inv_in[862] ),
    .A(\inv_in[861] ));
 sg13g2_inv_2 \inv[862]/_0_  (.Y(\inv_in[863] ),
    .A(\inv_in[862] ));
 sg13g2_inv_2 \inv[863]/_0_  (.Y(\inv_in[864] ),
    .A(\inv_in[863] ));
 sg13g2_inv_2 \inv[864]/_0_  (.Y(\inv_in[865] ),
    .A(\inv_in[864] ));
 sg13g2_inv_2 \inv[865]/_0_  (.Y(\inv_in[866] ),
    .A(\inv_in[865] ));
 sg13g2_inv_2 \inv[866]/_0_  (.Y(\inv_in[867] ),
    .A(\inv_in[866] ));
 sg13g2_inv_2 \inv[867]/_0_  (.Y(\inv_in[868] ),
    .A(\inv_in[867] ));
 sg13g2_inv_2 \inv[868]/_0_  (.Y(\inv_in[869] ),
    .A(\inv_in[868] ));
 sg13g2_inv_2 \inv[869]/_0_  (.Y(\inv_in[870] ),
    .A(\inv_in[869] ));
 sg13g2_inv_2 \inv[86]/_0_  (.Y(\inv_in[87] ),
    .A(\inv_in[86] ));
 sg13g2_inv_2 \inv[870]/_0_  (.Y(\inv_in[871] ),
    .A(\inv_in[870] ));
 sg13g2_inv_2 \inv[871]/_0_  (.Y(\inv_in[872] ),
    .A(\inv_in[871] ));
 sg13g2_inv_2 \inv[872]/_0_  (.Y(\inv_in[873] ),
    .A(\inv_in[872] ));
 sg13g2_inv_2 \inv[873]/_0_  (.Y(\inv_in[874] ),
    .A(\inv_in[873] ));
 sg13g2_inv_2 \inv[874]/_0_  (.Y(\inv_in[875] ),
    .A(\inv_in[874] ));
 sg13g2_inv_2 \inv[875]/_0_  (.Y(\inv_in[876] ),
    .A(\inv_in[875] ));
 sg13g2_inv_2 \inv[876]/_0_  (.Y(\inv_in[877] ),
    .A(\inv_in[876] ));
 sg13g2_inv_2 \inv[877]/_0_  (.Y(\inv_in[878] ),
    .A(\inv_in[877] ));
 sg13g2_inv_2 \inv[878]/_0_  (.Y(\inv_in[879] ),
    .A(\inv_in[878] ));
 sg13g2_inv_2 \inv[879]/_0_  (.Y(\inv_in[880] ),
    .A(\inv_in[879] ));
 sg13g2_inv_2 \inv[87]/_0_  (.Y(\inv_in[88] ),
    .A(\inv_in[87] ));
 sg13g2_inv_2 \inv[880]/_0_  (.Y(\inv_in[881] ),
    .A(\inv_in[880] ));
 sg13g2_inv_2 \inv[881]/_0_  (.Y(\inv_in[882] ),
    .A(\inv_in[881] ));
 sg13g2_inv_2 \inv[882]/_0_  (.Y(\inv_in[883] ),
    .A(\inv_in[882] ));
 sg13g2_inv_2 \inv[883]/_0_  (.Y(\inv_in[884] ),
    .A(\inv_in[883] ));
 sg13g2_inv_2 \inv[884]/_0_  (.Y(\inv_in[885] ),
    .A(\inv_in[884] ));
 sg13g2_inv_2 \inv[885]/_0_  (.Y(\inv_in[886] ),
    .A(\inv_in[885] ));
 sg13g2_inv_2 \inv[886]/_0_  (.Y(\inv_in[887] ),
    .A(\inv_in[886] ));
 sg13g2_inv_2 \inv[887]/_0_  (.Y(\inv_in[888] ),
    .A(\inv_in[887] ));
 sg13g2_inv_2 \inv[888]/_0_  (.Y(\inv_in[889] ),
    .A(\inv_in[888] ));
 sg13g2_inv_2 \inv[889]/_0_  (.Y(\inv_in[890] ),
    .A(\inv_in[889] ));
 sg13g2_inv_2 \inv[88]/_0_  (.Y(\inv_in[89] ),
    .A(\inv_in[88] ));
 sg13g2_inv_2 \inv[890]/_0_  (.Y(\inv_in[891] ),
    .A(\inv_in[890] ));
 sg13g2_inv_2 \inv[891]/_0_  (.Y(\inv_in[892] ),
    .A(\inv_in[891] ));
 sg13g2_inv_2 \inv[892]/_0_  (.Y(\inv_in[893] ),
    .A(\inv_in[892] ));
 sg13g2_inv_2 \inv[893]/_0_  (.Y(\inv_in[894] ),
    .A(\inv_in[893] ));
 sg13g2_inv_2 \inv[894]/_0_  (.Y(\inv_in[895] ),
    .A(\inv_in[894] ));
 sg13g2_inv_2 \inv[895]/_0_  (.Y(\inv_in[896] ),
    .A(\inv_in[895] ));
 sg13g2_inv_2 \inv[896]/_0_  (.Y(\inv_in[897] ),
    .A(\inv_in[896] ));
 sg13g2_inv_2 \inv[897]/_0_  (.Y(\inv_in[898] ),
    .A(\inv_in[897] ));
 sg13g2_inv_2 \inv[898]/_0_  (.Y(\inv_in[899] ),
    .A(\inv_in[898] ));
 sg13g2_inv_2 \inv[899]/_0_  (.Y(\inv_in[900] ),
    .A(\inv_in[899] ));
 sg13g2_inv_2 \inv[89]/_0_  (.Y(\inv_in[90] ),
    .A(\inv_in[89] ));
 sg13g2_inv_2 \inv[8]/_0_  (.Y(\inv_in[9] ),
    .A(\inv_in[8] ));
 sg13g2_inv_2 \inv[900]/_0_  (.Y(\inv_in[901] ),
    .A(\inv_in[900] ));
 sg13g2_inv_2 \inv[901]/_0_  (.Y(\inv_in[902] ),
    .A(\inv_in[901] ));
 sg13g2_inv_2 \inv[902]/_0_  (.Y(\inv_in[903] ),
    .A(\inv_in[902] ));
 sg13g2_inv_2 \inv[903]/_0_  (.Y(\inv_in[904] ),
    .A(\inv_in[903] ));
 sg13g2_inv_2 \inv[904]/_0_  (.Y(\inv_in[905] ),
    .A(\inv_in[904] ));
 sg13g2_inv_2 \inv[905]/_0_  (.Y(\inv_in[906] ),
    .A(\inv_in[905] ));
 sg13g2_inv_2 \inv[906]/_0_  (.Y(\inv_in[907] ),
    .A(\inv_in[906] ));
 sg13g2_inv_2 \inv[907]/_0_  (.Y(\inv_in[908] ),
    .A(\inv_in[907] ));
 sg13g2_inv_2 \inv[908]/_0_  (.Y(\inv_in[909] ),
    .A(\inv_in[908] ));
 sg13g2_inv_2 \inv[909]/_0_  (.Y(\inv_in[910] ),
    .A(\inv_in[909] ));
 sg13g2_inv_2 \inv[90]/_0_  (.Y(\inv_in[91] ),
    .A(\inv_in[90] ));
 sg13g2_inv_2 \inv[910]/_0_  (.Y(\inv_in[911] ),
    .A(\inv_in[910] ));
 sg13g2_inv_2 \inv[911]/_0_  (.Y(\inv_in[912] ),
    .A(\inv_in[911] ));
 sg13g2_inv_2 \inv[912]/_0_  (.Y(\inv_in[913] ),
    .A(\inv_in[912] ));
 sg13g2_inv_2 \inv[913]/_0_  (.Y(\inv_in[914] ),
    .A(\inv_in[913] ));
 sg13g2_inv_2 \inv[914]/_0_  (.Y(\inv_in[915] ),
    .A(\inv_in[914] ));
 sg13g2_inv_2 \inv[915]/_0_  (.Y(\inv_in[916] ),
    .A(\inv_in[915] ));
 sg13g2_inv_2 \inv[916]/_0_  (.Y(\inv_in[917] ),
    .A(\inv_in[916] ));
 sg13g2_inv_2 \inv[917]/_0_  (.Y(\inv_in[918] ),
    .A(\inv_in[917] ));
 sg13g2_inv_2 \inv[918]/_0_  (.Y(\inv_in[919] ),
    .A(\inv_in[918] ));
 sg13g2_inv_2 \inv[919]/_0_  (.Y(\inv_in[920] ),
    .A(\inv_in[919] ));
 sg13g2_inv_2 \inv[91]/_0_  (.Y(\inv_in[92] ),
    .A(\inv_in[91] ));
 sg13g2_inv_2 \inv[920]/_0_  (.Y(\inv_in[921] ),
    .A(\inv_in[920] ));
 sg13g2_inv_2 \inv[921]/_0_  (.Y(\inv_in[922] ),
    .A(\inv_in[921] ));
 sg13g2_inv_2 \inv[922]/_0_  (.Y(\inv_in[923] ),
    .A(\inv_in[922] ));
 sg13g2_inv_2 \inv[923]/_0_  (.Y(\inv_in[924] ),
    .A(\inv_in[923] ));
 sg13g2_inv_2 \inv[924]/_0_  (.Y(\inv_in[925] ),
    .A(\inv_in[924] ));
 sg13g2_inv_2 \inv[925]/_0_  (.Y(\inv_in[926] ),
    .A(\inv_in[925] ));
 sg13g2_inv_2 \inv[926]/_0_  (.Y(\inv_in[927] ),
    .A(\inv_in[926] ));
 sg13g2_inv_2 \inv[927]/_0_  (.Y(\inv_in[928] ),
    .A(\inv_in[927] ));
 sg13g2_inv_2 \inv[928]/_0_  (.Y(\inv_in[929] ),
    .A(\inv_in[928] ));
 sg13g2_inv_2 \inv[929]/_0_  (.Y(\inv_in[930] ),
    .A(\inv_in[929] ));
 sg13g2_inv_2 \inv[92]/_0_  (.Y(\inv_in[93] ),
    .A(\inv_in[92] ));
 sg13g2_inv_2 \inv[930]/_0_  (.Y(\inv_in[931] ),
    .A(\inv_in[930] ));
 sg13g2_inv_2 \inv[931]/_0_  (.Y(\inv_in[932] ),
    .A(\inv_in[931] ));
 sg13g2_inv_2 \inv[932]/_0_  (.Y(\inv_in[933] ),
    .A(\inv_in[932] ));
 sg13g2_inv_2 \inv[933]/_0_  (.Y(\inv_in[934] ),
    .A(\inv_in[933] ));
 sg13g2_inv_2 \inv[934]/_0_  (.Y(\inv_in[935] ),
    .A(\inv_in[934] ));
 sg13g2_inv_2 \inv[935]/_0_  (.Y(\inv_in[936] ),
    .A(\inv_in[935] ));
 sg13g2_inv_2 \inv[936]/_0_  (.Y(\inv_in[937] ),
    .A(\inv_in[936] ));
 sg13g2_inv_2 \inv[937]/_0_  (.Y(\inv_in[938] ),
    .A(\inv_in[937] ));
 sg13g2_inv_2 \inv[938]/_0_  (.Y(\inv_in[939] ),
    .A(\inv_in[938] ));
 sg13g2_inv_2 \inv[939]/_0_  (.Y(\inv_in[940] ),
    .A(\inv_in[939] ));
 sg13g2_inv_2 \inv[93]/_0_  (.Y(\inv_in[94] ),
    .A(\inv_in[93] ));
 sg13g2_inv_2 \inv[940]/_0_  (.Y(\inv_in[941] ),
    .A(\inv_in[940] ));
 sg13g2_inv_2 \inv[941]/_0_  (.Y(\inv_in[942] ),
    .A(\inv_in[941] ));
 sg13g2_inv_2 \inv[942]/_0_  (.Y(\inv_in[943] ),
    .A(\inv_in[942] ));
 sg13g2_inv_2 \inv[943]/_0_  (.Y(\inv_in[944] ),
    .A(\inv_in[943] ));
 sg13g2_inv_2 \inv[944]/_0_  (.Y(\inv_in[945] ),
    .A(\inv_in[944] ));
 sg13g2_inv_2 \inv[945]/_0_  (.Y(\inv_in[946] ),
    .A(\inv_in[945] ));
 sg13g2_inv_2 \inv[946]/_0_  (.Y(\inv_in[947] ),
    .A(\inv_in[946] ));
 sg13g2_inv_2 \inv[947]/_0_  (.Y(\inv_in[948] ),
    .A(\inv_in[947] ));
 sg13g2_inv_2 \inv[948]/_0_  (.Y(\inv_in[949] ),
    .A(\inv_in[948] ));
 sg13g2_inv_2 \inv[949]/_0_  (.Y(\inv_in[950] ),
    .A(\inv_in[949] ));
 sg13g2_inv_2 \inv[94]/_0_  (.Y(\inv_in[95] ),
    .A(\inv_in[94] ));
 sg13g2_inv_2 \inv[950]/_0_  (.Y(\inv_in[951] ),
    .A(\inv_in[950] ));
 sg13g2_inv_2 \inv[951]/_0_  (.Y(\inv_in[952] ),
    .A(\inv_in[951] ));
 sg13g2_inv_2 \inv[952]/_0_  (.Y(\inv_in[953] ),
    .A(\inv_in[952] ));
 sg13g2_inv_2 \inv[953]/_0_  (.Y(\inv_in[954] ),
    .A(\inv_in[953] ));
 sg13g2_inv_2 \inv[954]/_0_  (.Y(\inv_in[955] ),
    .A(\inv_in[954] ));
 sg13g2_inv_2 \inv[955]/_0_  (.Y(\inv_in[956] ),
    .A(\inv_in[955] ));
 sg13g2_inv_2 \inv[956]/_0_  (.Y(\inv_in[957] ),
    .A(\inv_in[956] ));
 sg13g2_inv_2 \inv[957]/_0_  (.Y(\inv_in[958] ),
    .A(\inv_in[957] ));
 sg13g2_inv_2 \inv[958]/_0_  (.Y(\inv_in[959] ),
    .A(\inv_in[958] ));
 sg13g2_inv_2 \inv[959]/_0_  (.Y(\inv_in[960] ),
    .A(\inv_in[959] ));
 sg13g2_inv_2 \inv[95]/_0_  (.Y(\inv_in[96] ),
    .A(\inv_in[95] ));
 sg13g2_inv_2 \inv[960]/_0_  (.Y(\inv_in[961] ),
    .A(\inv_in[960] ));
 sg13g2_inv_2 \inv[961]/_0_  (.Y(\inv_in[962] ),
    .A(\inv_in[961] ));
 sg13g2_inv_2 \inv[962]/_0_  (.Y(\inv_in[963] ),
    .A(\inv_in[962] ));
 sg13g2_inv_2 \inv[963]/_0_  (.Y(\inv_in[964] ),
    .A(\inv_in[963] ));
 sg13g2_inv_2 \inv[964]/_0_  (.Y(\inv_in[965] ),
    .A(\inv_in[964] ));
 sg13g2_inv_2 \inv[965]/_0_  (.Y(\inv_in[966] ),
    .A(\inv_in[965] ));
 sg13g2_inv_2 \inv[966]/_0_  (.Y(\inv_in[967] ),
    .A(\inv_in[966] ));
 sg13g2_inv_2 \inv[967]/_0_  (.Y(\inv_in[968] ),
    .A(\inv_in[967] ));
 sg13g2_inv_2 \inv[968]/_0_  (.Y(\inv_in[969] ),
    .A(\inv_in[968] ));
 sg13g2_inv_2 \inv[969]/_0_  (.Y(\inv_in[970] ),
    .A(\inv_in[969] ));
 sg13g2_inv_2 \inv[96]/_0_  (.Y(\inv_in[97] ),
    .A(\inv_in[96] ));
 sg13g2_inv_2 \inv[970]/_0_  (.Y(\inv_in[971] ),
    .A(\inv_in[970] ));
 sg13g2_inv_2 \inv[971]/_0_  (.Y(\inv_in[972] ),
    .A(\inv_in[971] ));
 sg13g2_inv_2 \inv[972]/_0_  (.Y(\inv_in[973] ),
    .A(\inv_in[972] ));
 sg13g2_inv_2 \inv[973]/_0_  (.Y(\inv_in[974] ),
    .A(\inv_in[973] ));
 sg13g2_inv_2 \inv[974]/_0_  (.Y(\inv_in[975] ),
    .A(\inv_in[974] ));
 sg13g2_inv_2 \inv[975]/_0_  (.Y(\inv_in[976] ),
    .A(\inv_in[975] ));
 sg13g2_inv_2 \inv[976]/_0_  (.Y(\inv_in[977] ),
    .A(\inv_in[976] ));
 sg13g2_inv_2 \inv[977]/_0_  (.Y(\inv_in[978] ),
    .A(\inv_in[977] ));
 sg13g2_inv_2 \inv[978]/_0_  (.Y(\inv_in[979] ),
    .A(\inv_in[978] ));
 sg13g2_inv_2 \inv[979]/_0_  (.Y(\inv_in[980] ),
    .A(\inv_in[979] ));
 sg13g2_inv_2 \inv[97]/_0_  (.Y(\inv_in[98] ),
    .A(\inv_in[97] ));
 sg13g2_inv_2 \inv[980]/_0_  (.Y(\inv_in[981] ),
    .A(\inv_in[980] ));
 sg13g2_inv_2 \inv[981]/_0_  (.Y(\inv_in[982] ),
    .A(\inv_in[981] ));
 sg13g2_inv_2 \inv[982]/_0_  (.Y(\inv_in[983] ),
    .A(\inv_in[982] ));
 sg13g2_inv_2 \inv[983]/_0_  (.Y(\inv_in[984] ),
    .A(\inv_in[983] ));
 sg13g2_inv_2 \inv[984]/_0_  (.Y(\inv_in[985] ),
    .A(\inv_in[984] ));
 sg13g2_inv_2 \inv[985]/_0_  (.Y(\inv_in[986] ),
    .A(\inv_in[985] ));
 sg13g2_inv_2 \inv[986]/_0_  (.Y(\inv_in[987] ),
    .A(\inv_in[986] ));
 sg13g2_inv_2 \inv[987]/_0_  (.Y(\inv_in[988] ),
    .A(\inv_in[987] ));
 sg13g2_inv_2 \inv[988]/_0_  (.Y(\inv_in[989] ),
    .A(\inv_in[988] ));
 sg13g2_inv_2 \inv[989]/_0_  (.Y(\inv_in[990] ),
    .A(\inv_in[989] ));
 sg13g2_inv_2 \inv[98]/_0_  (.Y(\inv_in[99] ),
    .A(\inv_in[98] ));
 sg13g2_inv_2 \inv[990]/_0_  (.Y(\inv_in[991] ),
    .A(\inv_in[990] ));
 sg13g2_inv_2 \inv[991]/_0_  (.Y(\inv_in[992] ),
    .A(\inv_in[991] ));
 sg13g2_inv_2 \inv[992]/_0_  (.Y(\inv_in[993] ),
    .A(\inv_in[992] ));
 sg13g2_inv_2 \inv[993]/_0_  (.Y(\inv_in[994] ),
    .A(\inv_in[993] ));
 sg13g2_inv_2 \inv[994]/_0_  (.Y(\inv_in[995] ),
    .A(\inv_in[994] ));
 sg13g2_inv_2 \inv[995]/_0_  (.Y(\inv_in[996] ),
    .A(\inv_in[995] ));
 sg13g2_inv_2 \inv[996]/_0_  (.Y(\inv_in[997] ),
    .A(\inv_in[996] ));
 sg13g2_inv_2 \inv[997]/_0_  (.Y(\inv_in[998] ),
    .A(\inv_in[997] ));
 sg13g2_inv_2 \inv[998]/_0_  (.Y(\inv_in[999] ),
    .A(\inv_in[998] ));
 sg13g2_inv_2 \inv[999]/_0_  (.Y(\inv_in[1000] ),
    .A(\inv_in[999] ));
 sg13g2_inv_2 \inv[99]/_0_  (.Y(\inv_in[100] ),
    .A(\inv_in[99] ));
 sg13g2_inv_2 \inv[9]/_0_  (.Y(\inv_in[10] ),
    .A(\inv_in[9] ));
 sg13g2_buf_16 input1 (.X(net1),
    .A(ui_in[0]));
 sg13g2_buf_1 output2 (.A(net2),
    .X(uio_out[0]));
 sg13g2_buf_1 output3 (.A(net3),
    .X(uio_out[1]));
 sg13g2_buf_1 output4 (.A(net4),
    .X(uio_out[2]));
 sg13g2_buf_1 output5 (.A(net5),
    .X(uio_out[3]));
 sg13g2_buf_1 output6 (.A(net6),
    .X(uio_out[4]));
 sg13g2_buf_1 output7 (.A(net7),
    .X(uio_out[5]));
 sg13g2_buf_1 output8 (.A(net8),
    .X(uo_out[0]));
 sg13g2_buf_1 output9 (.A(net9),
    .X(uo_out[1]));
 sg13g2_buf_1 output10 (.A(net10),
    .X(uo_out[2]));
 sg13g2_buf_1 output11 (.A(net11),
    .X(uo_out[3]));
 sg13g2_buf_1 output12 (.A(net12),
    .X(uo_out[4]));
 sg13g2_buf_1 output13 (.A(net13),
    .X(uo_out[5]));
 sg13g2_buf_1 output14 (.A(net14),
    .X(uo_out[6]));
 sg13g2_buf_1 output15 (.A(net15),
    .X(uo_out[7]));
 sg13g2_tielo _16__16 (.L_LO(net16));
 sg13g2_tielo _17__17 (.L_LO(net17));
 sg13g2_tiehi _05__19 (.L_HI(net19));
 sg13g2_tiehi _06__20 (.L_HI(net20));
 sg13g2_tiehi _07__21 (.L_HI(net21));
 sg13g2_tiehi _08__22 (.L_HI(net22));
 sg13g2_tiehi _09__23 (.L_HI(net23));
 sg13g2_tiehi _10__24 (.L_HI(net24));
 sg13g2_tiehi _26__25 (.L_HI(net25));
 sg13g2_fill_1 FILLER_0_14 ();
 sg13g2_fill_1 FILLER_0_19 ();
 sg13g2_fill_1 FILLER_0_164 ();
 sg13g2_fill_2 FILLER_0_397 ();
 sg13g2_fill_1 FILLER_0_403 ();
 sg13g2_fill_2 FILLER_0_412 ();
 sg13g2_fill_2 FILLER_1_12 ();
 sg13g2_fill_1 FILLER_1_18 ();
 sg13g2_fill_1 FILLER_1_23 ();
 sg13g2_fill_1 FILLER_1_92 ();
 sg13g2_fill_1 FILLER_1_97 ();
 sg13g2_fill_1 FILLER_1_106 ();
 sg13g2_fill_1 FILLER_1_115 ();
 sg13g2_fill_1 FILLER_1_120 ();
 sg13g2_fill_2 FILLER_1_141 ();
 sg13g2_fill_1 FILLER_1_143 ();
 sg13g2_fill_1 FILLER_1_208 ();
 sg13g2_fill_1 FILLER_1_213 ();
 sg13g2_fill_2 FILLER_1_396 ();
 sg13g2_fill_1 FILLER_1_398 ();
 sg13g2_fill_1 FILLER_1_425 ();
 sg13g2_fill_2 FILLER_2_8 ();
 sg13g2_fill_1 FILLER_2_10 ();
 sg13g2_fill_1 FILLER_2_59 ();
 sg13g2_fill_2 FILLER_2_96 ();
 sg13g2_fill_1 FILLER_2_126 ();
 sg13g2_fill_2 FILLER_2_187 ();
 sg13g2_fill_2 FILLER_2_193 ();
 sg13g2_fill_1 FILLER_2_235 ();
 sg13g2_fill_1 FILLER_2_266 ();
 sg13g2_fill_1 FILLER_2_279 ();
 sg13g2_fill_1 FILLER_2_284 ();
 sg13g2_fill_1 FILLER_2_293 ();
 sg13g2_fill_1 FILLER_2_298 ();
 sg13g2_fill_1 FILLER_2_303 ();
 sg13g2_fill_1 FILLER_2_320 ();
 sg13g2_fill_2 FILLER_2_345 ();
 sg13g2_fill_1 FILLER_2_351 ();
 sg13g2_fill_1 FILLER_2_356 ();
 sg13g2_fill_2 FILLER_2_393 ();
 sg13g2_fill_2 FILLER_2_399 ();
 sg13g2_fill_2 FILLER_2_405 ();
 sg13g2_fill_1 FILLER_2_407 ();
 sg13g2_fill_2 FILLER_2_416 ();
 sg13g2_fill_1 FILLER_3_0 ();
 sg13g2_fill_2 FILLER_3_5 ();
 sg13g2_fill_1 FILLER_3_7 ();
 sg13g2_fill_2 FILLER_3_20 ();
 sg13g2_fill_1 FILLER_3_22 ();
 sg13g2_fill_1 FILLER_3_27 ();
 sg13g2_fill_1 FILLER_3_32 ();
 sg13g2_fill_1 FILLER_3_69 ();
 sg13g2_fill_2 FILLER_3_86 ();
 sg13g2_fill_2 FILLER_3_92 ();
 sg13g2_fill_1 FILLER_3_94 ();
 sg13g2_fill_2 FILLER_3_119 ();
 sg13g2_fill_2 FILLER_3_145 ();
 sg13g2_fill_2 FILLER_3_391 ();
 sg13g2_fill_2 FILLER_3_401 ();
 sg13g2_fill_1 FILLER_3_403 ();
 sg13g2_fill_2 FILLER_3_408 ();
 sg13g2_fill_2 FILLER_3_418 ();
 sg13g2_fill_2 FILLER_3_428 ();
 sg13g2_fill_1 FILLER_4_4 ();
 sg13g2_fill_2 FILLER_4_17 ();
 sg13g2_fill_1 FILLER_4_19 ();
 sg13g2_fill_1 FILLER_4_24 ();
 sg13g2_fill_2 FILLER_4_93 ();
 sg13g2_fill_1 FILLER_4_95 ();
 sg13g2_fill_2 FILLER_4_164 ();
 sg13g2_fill_2 FILLER_4_182 ();
 sg13g2_fill_1 FILLER_4_184 ();
 sg13g2_fill_1 FILLER_4_209 ();
 sg13g2_fill_1 FILLER_4_214 ();
 sg13g2_fill_2 FILLER_4_305 ();
 sg13g2_fill_1 FILLER_4_307 ();
 sg13g2_fill_2 FILLER_4_340 ();
 sg13g2_fill_1 FILLER_4_342 ();
 sg13g2_fill_1 FILLER_4_409 ();
 sg13g2_fill_2 FILLER_4_418 ();
 sg13g2_fill_1 FILLER_4_420 ();
 sg13g2_fill_1 FILLER_4_425 ();
 sg13g2_fill_2 FILLER_5_4 ();
 sg13g2_fill_1 FILLER_5_6 ();
 sg13g2_fill_2 FILLER_5_15 ();
 sg13g2_fill_1 FILLER_5_33 ();
 sg13g2_fill_1 FILLER_5_58 ();
 sg13g2_fill_1 FILLER_5_63 ();
 sg13g2_fill_1 FILLER_5_88 ();
 sg13g2_fill_1 FILLER_5_97 ();
 sg13g2_fill_2 FILLER_5_122 ();
 sg13g2_fill_1 FILLER_5_124 ();
 sg13g2_fill_1 FILLER_5_169 ();
 sg13g2_fill_2 FILLER_5_174 ();
 sg13g2_fill_1 FILLER_5_200 ();
 sg13g2_fill_1 FILLER_5_229 ();
 sg13g2_fill_1 FILLER_5_238 ();
 sg13g2_fill_1 FILLER_5_247 ();
 sg13g2_fill_1 FILLER_5_252 ();
 sg13g2_fill_1 FILLER_5_261 ();
 sg13g2_fill_1 FILLER_5_276 ();
 sg13g2_fill_1 FILLER_5_397 ();
 sg13g2_fill_2 FILLER_5_410 ();
 sg13g2_fill_1 FILLER_5_412 ();
 sg13g2_fill_2 FILLER_5_421 ();
 sg13g2_fill_1 FILLER_5_423 ();
 sg13g2_fill_2 FILLER_5_428 ();
 sg13g2_fill_1 FILLER_6_16 ();
 sg13g2_fill_2 FILLER_6_21 ();
 sg13g2_fill_1 FILLER_6_23 ();
 sg13g2_fill_1 FILLER_6_96 ();
 sg13g2_fill_1 FILLER_6_101 ();
 sg13g2_fill_1 FILLER_6_122 ();
 sg13g2_fill_2 FILLER_6_155 ();
 sg13g2_fill_2 FILLER_6_163 ();
 sg13g2_fill_2 FILLER_6_399 ();
 sg13g2_fill_1 FILLER_6_401 ();
 sg13g2_fill_1 FILLER_6_410 ();
 sg13g2_fill_1 FILLER_6_419 ();
 sg13g2_fill_1 FILLER_6_424 ();
 sg13g2_fill_1 FILLER_6_429 ();
 sg13g2_fill_1 FILLER_7_0 ();
 sg13g2_fill_1 FILLER_7_9 ();
 sg13g2_fill_2 FILLER_7_18 ();
 sg13g2_fill_1 FILLER_7_20 ();
 sg13g2_fill_2 FILLER_7_53 ();
 sg13g2_fill_2 FILLER_7_107 ();
 sg13g2_fill_2 FILLER_7_141 ();
 sg13g2_fill_2 FILLER_7_159 ();
 sg13g2_fill_1 FILLER_7_169 ();
 sg13g2_fill_1 FILLER_7_174 ();
 sg13g2_fill_2 FILLER_7_261 ();
 sg13g2_fill_2 FILLER_7_285 ();
 sg13g2_fill_1 FILLER_7_297 ();
 sg13g2_fill_1 FILLER_7_402 ();
 sg13g2_fill_2 FILLER_7_415 ();
 sg13g2_fill_1 FILLER_7_429 ();
 sg13g2_fill_2 FILLER_8_16 ();
 sg13g2_fill_1 FILLER_8_22 ();
 sg13g2_fill_2 FILLER_8_27 ();
 sg13g2_fill_2 FILLER_8_85 ();
 sg13g2_fill_1 FILLER_8_87 ();
 sg13g2_fill_2 FILLER_8_116 ();
 sg13g2_fill_1 FILLER_8_118 ();
 sg13g2_fill_2 FILLER_8_139 ();
 sg13g2_fill_2 FILLER_8_193 ();
 sg13g2_fill_1 FILLER_8_301 ();
 sg13g2_fill_2 FILLER_8_348 ();
 sg13g2_fill_2 FILLER_8_418 ();
 sg13g2_fill_2 FILLER_8_428 ();
 sg13g2_fill_1 FILLER_9_0 ();
 sg13g2_fill_2 FILLER_9_13 ();
 sg13g2_fill_1 FILLER_9_15 ();
 sg13g2_fill_1 FILLER_9_36 ();
 sg13g2_fill_2 FILLER_9_45 ();
 sg13g2_fill_1 FILLER_9_47 ();
 sg13g2_fill_1 FILLER_9_52 ();
 sg13g2_fill_2 FILLER_9_85 ();
 sg13g2_fill_1 FILLER_9_87 ();
 sg13g2_fill_1 FILLER_9_112 ();
 sg13g2_fill_1 FILLER_9_121 ();
 sg13g2_fill_1 FILLER_9_126 ();
 sg13g2_fill_1 FILLER_9_135 ();
 sg13g2_fill_2 FILLER_9_168 ();
 sg13g2_fill_1 FILLER_9_186 ();
 sg13g2_fill_1 FILLER_9_195 ();
 sg13g2_fill_1 FILLER_9_204 ();
 sg13g2_fill_2 FILLER_9_241 ();
 sg13g2_fill_1 FILLER_9_259 ();
 sg13g2_fill_2 FILLER_9_272 ();
 sg13g2_fill_1 FILLER_9_352 ();
 sg13g2_fill_2 FILLER_9_409 ();
 sg13g2_fill_1 FILLER_9_411 ();
 sg13g2_fill_1 FILLER_9_420 ();
 sg13g2_fill_1 FILLER_9_429 ();
 sg13g2_fill_1 FILLER_10_4 ();
 sg13g2_fill_2 FILLER_10_37 ();
 sg13g2_fill_1 FILLER_10_59 ();
 sg13g2_fill_1 FILLER_10_72 ();
 sg13g2_fill_2 FILLER_10_77 ();
 sg13g2_fill_2 FILLER_10_87 ();
 sg13g2_fill_1 FILLER_10_89 ();
 sg13g2_fill_2 FILLER_10_148 ();
 sg13g2_fill_1 FILLER_10_202 ();
 sg13g2_fill_1 FILLER_10_211 ();
 sg13g2_fill_1 FILLER_10_216 ();
 sg13g2_fill_2 FILLER_10_221 ();
 sg13g2_fill_1 FILLER_10_227 ();
 sg13g2_fill_2 FILLER_10_232 ();
 sg13g2_fill_2 FILLER_10_254 ();
 sg13g2_fill_1 FILLER_10_360 ();
 sg13g2_fill_2 FILLER_10_421 ();
 sg13g2_fill_1 FILLER_10_423 ();
 sg13g2_fill_2 FILLER_10_428 ();
 sg13g2_fill_2 FILLER_11_0 ();
 sg13g2_fill_1 FILLER_11_2 ();
 sg13g2_fill_2 FILLER_11_11 ();
 sg13g2_fill_2 FILLER_11_33 ();
 sg13g2_fill_1 FILLER_11_35 ();
 sg13g2_fill_1 FILLER_11_84 ();
 sg13g2_fill_1 FILLER_11_89 ();
 sg13g2_fill_1 FILLER_11_114 ();
 sg13g2_fill_1 FILLER_11_119 ();
 sg13g2_fill_2 FILLER_11_192 ();
 sg13g2_fill_2 FILLER_11_198 ();
 sg13g2_fill_1 FILLER_11_200 ();
 sg13g2_fill_2 FILLER_11_269 ();
 sg13g2_fill_1 FILLER_11_271 ();
 sg13g2_fill_2 FILLER_11_342 ();
 sg13g2_fill_2 FILLER_11_370 ();
 sg13g2_fill_1 FILLER_11_372 ();
 sg13g2_fill_1 FILLER_11_419 ();
 sg13g2_fill_2 FILLER_11_428 ();
 sg13g2_fill_2 FILLER_12_0 ();
 sg13g2_fill_1 FILLER_12_10 ();
 sg13g2_fill_1 FILLER_12_23 ();
 sg13g2_fill_1 FILLER_12_36 ();
 sg13g2_fill_2 FILLER_12_41 ();
 sg13g2_fill_1 FILLER_12_43 ();
 sg13g2_fill_1 FILLER_12_104 ();
 sg13g2_fill_2 FILLER_12_141 ();
 sg13g2_fill_1 FILLER_12_167 ();
 sg13g2_fill_1 FILLER_12_176 ();
 sg13g2_fill_1 FILLER_12_181 ();
 sg13g2_fill_1 FILLER_12_294 ();
 sg13g2_fill_2 FILLER_12_371 ();
 sg13g2_fill_1 FILLER_12_373 ();
 sg13g2_fill_2 FILLER_12_394 ();
 sg13g2_fill_2 FILLER_12_428 ();
 sg13g2_fill_2 FILLER_13_0 ();
 sg13g2_fill_2 FILLER_13_14 ();
 sg13g2_fill_1 FILLER_13_120 ();
 sg13g2_fill_1 FILLER_13_153 ();
 sg13g2_fill_1 FILLER_13_158 ();
 sg13g2_fill_1 FILLER_13_163 ();
 sg13g2_fill_2 FILLER_13_176 ();
 sg13g2_fill_2 FILLER_13_210 ();
 sg13g2_fill_1 FILLER_13_280 ();
 sg13g2_fill_1 FILLER_13_313 ();
 sg13g2_fill_1 FILLER_13_326 ();
 sg13g2_fill_1 FILLER_13_335 ();
 sg13g2_fill_1 FILLER_13_348 ();
 sg13g2_fill_2 FILLER_13_373 ();
 sg13g2_fill_1 FILLER_13_417 ();
 sg13g2_fill_2 FILLER_14_8 ();
 sg13g2_fill_2 FILLER_14_22 ();
 sg13g2_fill_2 FILLER_14_40 ();
 sg13g2_fill_1 FILLER_14_46 ();
 sg13g2_fill_1 FILLER_14_51 ();
 sg13g2_fill_2 FILLER_14_140 ();
 sg13g2_fill_1 FILLER_14_142 ();
 sg13g2_fill_2 FILLER_14_179 ();
 sg13g2_fill_2 FILLER_14_233 ();
 sg13g2_fill_1 FILLER_14_235 ();
 sg13g2_fill_1 FILLER_14_292 ();
 sg13g2_fill_1 FILLER_14_355 ();
 sg13g2_fill_1 FILLER_14_376 ();
 sg13g2_fill_1 FILLER_14_409 ();
 sg13g2_fill_2 FILLER_14_418 ();
 sg13g2_fill_1 FILLER_14_420 ();
 sg13g2_fill_1 FILLER_14_429 ();
 sg13g2_fill_2 FILLER_15_0 ();
 sg13g2_fill_2 FILLER_15_6 ();
 sg13g2_fill_1 FILLER_15_12 ();
 sg13g2_fill_1 FILLER_15_41 ();
 sg13g2_fill_2 FILLER_15_110 ();
 sg13g2_fill_1 FILLER_15_120 ();
 sg13g2_fill_2 FILLER_15_165 ();
 sg13g2_fill_2 FILLER_15_203 ();
 sg13g2_fill_1 FILLER_15_213 ();
 sg13g2_fill_1 FILLER_15_218 ();
 sg13g2_fill_1 FILLER_15_223 ();
 sg13g2_fill_2 FILLER_15_240 ();
 sg13g2_fill_2 FILLER_15_274 ();
 sg13g2_fill_2 FILLER_15_308 ();
 sg13g2_fill_2 FILLER_15_366 ();
 sg13g2_fill_2 FILLER_15_380 ();
 sg13g2_fill_2 FILLER_15_394 ();
 sg13g2_fill_1 FILLER_15_408 ();
 sg13g2_fill_1 FILLER_15_425 ();
 sg13g2_fill_2 FILLER_16_0 ();
 sg13g2_fill_1 FILLER_16_26 ();
 sg13g2_fill_1 FILLER_16_31 ();
 sg13g2_fill_1 FILLER_16_40 ();
 sg13g2_fill_1 FILLER_16_57 ();
 sg13g2_fill_2 FILLER_16_86 ();
 sg13g2_fill_1 FILLER_16_88 ();
 sg13g2_fill_2 FILLER_16_163 ();
 sg13g2_fill_1 FILLER_16_169 ();
 sg13g2_fill_1 FILLER_16_190 ();
 sg13g2_fill_1 FILLER_16_195 ();
 sg13g2_fill_2 FILLER_16_288 ();
 sg13g2_fill_2 FILLER_16_314 ();
 sg13g2_fill_1 FILLER_16_316 ();
 sg13g2_fill_2 FILLER_16_341 ();
 sg13g2_fill_1 FILLER_16_343 ();
 sg13g2_fill_1 FILLER_16_420 ();
 sg13g2_fill_1 FILLER_16_425 ();
 sg13g2_fill_2 FILLER_17_0 ();
 sg13g2_fill_1 FILLER_17_42 ();
 sg13g2_fill_1 FILLER_17_51 ();
 sg13g2_fill_1 FILLER_17_92 ();
 sg13g2_fill_1 FILLER_17_209 ();
 sg13g2_fill_1 FILLER_17_234 ();
 sg13g2_fill_2 FILLER_17_255 ();
 sg13g2_fill_2 FILLER_17_277 ();
 sg13g2_fill_1 FILLER_17_279 ();
 sg13g2_fill_2 FILLER_17_296 ();
 sg13g2_fill_1 FILLER_17_298 ();
 sg13g2_fill_1 FILLER_17_319 ();
 sg13g2_fill_2 FILLER_17_324 ();
 sg13g2_fill_1 FILLER_17_408 ();
 sg13g2_fill_2 FILLER_17_421 ();
 sg13g2_fill_2 FILLER_17_427 ();
 sg13g2_fill_1 FILLER_17_429 ();
 sg13g2_fill_1 FILLER_18_0 ();
 sg13g2_fill_1 FILLER_18_25 ();
 sg13g2_fill_2 FILLER_18_40 ();
 sg13g2_fill_2 FILLER_18_46 ();
 sg13g2_fill_2 FILLER_18_68 ();
 sg13g2_fill_1 FILLER_18_90 ();
 sg13g2_fill_2 FILLER_18_103 ();
 sg13g2_fill_1 FILLER_18_121 ();
 sg13g2_fill_1 FILLER_18_158 ();
 sg13g2_fill_2 FILLER_18_163 ();
 sg13g2_fill_2 FILLER_18_233 ();
 sg13g2_fill_1 FILLER_18_239 ();
 sg13g2_fill_1 FILLER_18_244 ();
 sg13g2_fill_1 FILLER_18_249 ();
 sg13g2_fill_1 FILLER_18_290 ();
 sg13g2_fill_2 FILLER_18_329 ();
 sg13g2_fill_2 FILLER_18_427 ();
 sg13g2_fill_1 FILLER_18_429 ();
 sg13g2_fill_2 FILLER_19_20 ();
 sg13g2_fill_1 FILLER_19_30 ();
 sg13g2_fill_2 FILLER_19_35 ();
 sg13g2_fill_2 FILLER_19_77 ();
 sg13g2_fill_1 FILLER_19_95 ();
 sg13g2_fill_1 FILLER_19_122 ();
 sg13g2_fill_1 FILLER_19_147 ();
 sg13g2_fill_1 FILLER_19_200 ();
 sg13g2_fill_2 FILLER_19_225 ();
 sg13g2_fill_1 FILLER_19_227 ();
 sg13g2_fill_2 FILLER_19_256 ();
 sg13g2_fill_1 FILLER_19_262 ();
 sg13g2_fill_2 FILLER_19_267 ();
 sg13g2_fill_2 FILLER_19_289 ();
 sg13g2_fill_2 FILLER_19_333 ();
 sg13g2_fill_1 FILLER_19_353 ();
 sg13g2_fill_1 FILLER_19_378 ();
 sg13g2_fill_2 FILLER_19_391 ();
 sg13g2_fill_1 FILLER_19_397 ();
 sg13g2_fill_2 FILLER_19_410 ();
 sg13g2_fill_1 FILLER_19_412 ();
 sg13g2_fill_1 FILLER_19_429 ();
 sg13g2_fill_1 FILLER_20_0 ();
 sg13g2_fill_1 FILLER_20_5 ();
 sg13g2_fill_1 FILLER_20_10 ();
 sg13g2_fill_1 FILLER_20_15 ();
 sg13g2_fill_1 FILLER_20_24 ();
 sg13g2_fill_2 FILLER_20_29 ();
 sg13g2_fill_2 FILLER_20_55 ();
 sg13g2_fill_1 FILLER_20_97 ();
 sg13g2_fill_2 FILLER_20_102 ();
 sg13g2_fill_2 FILLER_20_124 ();
 sg13g2_fill_1 FILLER_20_138 ();
 sg13g2_fill_1 FILLER_20_155 ();
 sg13g2_fill_1 FILLER_20_160 ();
 sg13g2_fill_2 FILLER_20_165 ();
 sg13g2_fill_1 FILLER_20_183 ();
 sg13g2_fill_1 FILLER_20_192 ();
 sg13g2_fill_2 FILLER_20_269 ();
 sg13g2_fill_2 FILLER_20_279 ();
 sg13g2_fill_1 FILLER_20_285 ();
 sg13g2_fill_1 FILLER_20_290 ();
 sg13g2_fill_1 FILLER_20_307 ();
 sg13g2_fill_2 FILLER_20_318 ();
 sg13g2_fill_1 FILLER_20_350 ();
 sg13g2_fill_2 FILLER_20_367 ();
 sg13g2_fill_2 FILLER_20_409 ();
 sg13g2_fill_2 FILLER_20_415 ();
 sg13g2_fill_1 FILLER_20_417 ();
 sg13g2_fill_1 FILLER_21_8 ();
 sg13g2_fill_1 FILLER_21_13 ();
 sg13g2_fill_1 FILLER_21_18 ();
 sg13g2_fill_1 FILLER_21_23 ();
 sg13g2_fill_1 FILLER_21_28 ();
 sg13g2_fill_1 FILLER_21_33 ();
 sg13g2_fill_1 FILLER_21_38 ();
 sg13g2_fill_1 FILLER_21_43 ();
 sg13g2_fill_2 FILLER_21_48 ();
 sg13g2_fill_2 FILLER_21_74 ();
 sg13g2_fill_2 FILLER_21_112 ();
 sg13g2_fill_1 FILLER_21_140 ();
 sg13g2_fill_1 FILLER_21_145 ();
 sg13g2_fill_2 FILLER_21_150 ();
 sg13g2_fill_1 FILLER_21_192 ();
 sg13g2_fill_1 FILLER_21_233 ();
 sg13g2_fill_1 FILLER_21_338 ();
 sg13g2_fill_2 FILLER_21_351 ();
 sg13g2_fill_2 FILLER_21_411 ();
 sg13g2_fill_1 FILLER_21_413 ();
 sg13g2_fill_2 FILLER_22_38 ();
 sg13g2_fill_1 FILLER_22_64 ();
 sg13g2_fill_2 FILLER_22_89 ();
 sg13g2_fill_1 FILLER_22_91 ();
 sg13g2_fill_1 FILLER_22_148 ();
 sg13g2_fill_1 FILLER_22_193 ();
 sg13g2_fill_2 FILLER_22_206 ();
 sg13g2_fill_2 FILLER_22_248 ();
 sg13g2_fill_2 FILLER_22_258 ();
 sg13g2_fill_1 FILLER_22_260 ();
 sg13g2_fill_2 FILLER_22_273 ();
 sg13g2_fill_1 FILLER_22_275 ();
 sg13g2_fill_2 FILLER_22_292 ();
 sg13g2_fill_1 FILLER_22_310 ();
 sg13g2_fill_1 FILLER_22_335 ();
 sg13g2_fill_1 FILLER_22_402 ();
 sg13g2_fill_2 FILLER_22_415 ();
 sg13g2_fill_1 FILLER_22_417 ();
 sg13g2_fill_2 FILLER_23_40 ();
 sg13g2_fill_1 FILLER_23_42 ();
 sg13g2_fill_1 FILLER_23_47 ();
 sg13g2_fill_2 FILLER_23_52 ();
 sg13g2_fill_1 FILLER_23_58 ();
 sg13g2_fill_1 FILLER_23_67 ();
 sg13g2_fill_1 FILLER_23_72 ();
 sg13g2_fill_2 FILLER_23_77 ();
 sg13g2_fill_2 FILLER_23_99 ();
 sg13g2_fill_1 FILLER_23_101 ();
 sg13g2_fill_2 FILLER_23_106 ();
 sg13g2_fill_1 FILLER_23_160 ();
 sg13g2_fill_2 FILLER_23_165 ();
 sg13g2_fill_1 FILLER_23_179 ();
 sg13g2_fill_1 FILLER_23_184 ();
 sg13g2_fill_2 FILLER_23_305 ();
 sg13g2_fill_1 FILLER_23_319 ();
 sg13g2_fill_2 FILLER_23_348 ();
 sg13g2_fill_1 FILLER_23_418 ();
 sg13g2_fill_2 FILLER_23_427 ();
 sg13g2_fill_1 FILLER_23_429 ();
 sg13g2_fill_1 FILLER_24_0 ();
 sg13g2_fill_2 FILLER_24_5 ();
 sg13g2_fill_1 FILLER_24_7 ();
 sg13g2_fill_2 FILLER_24_26 ();
 sg13g2_fill_1 FILLER_24_28 ();
 sg13g2_fill_2 FILLER_24_47 ();
 sg13g2_fill_1 FILLER_24_69 ();
 sg13g2_fill_1 FILLER_24_114 ();
 sg13g2_fill_1 FILLER_24_123 ();
 sg13g2_fill_1 FILLER_24_128 ();
 sg13g2_fill_1 FILLER_24_133 ();
 sg13g2_fill_1 FILLER_24_138 ();
 sg13g2_fill_1 FILLER_24_143 ();
 sg13g2_fill_1 FILLER_24_148 ();
 sg13g2_fill_2 FILLER_24_153 ();
 sg13g2_fill_2 FILLER_24_207 ();
 sg13g2_fill_1 FILLER_24_237 ();
 sg13g2_fill_2 FILLER_24_242 ();
 sg13g2_fill_1 FILLER_24_244 ();
 sg13g2_fill_1 FILLER_24_265 ();
 sg13g2_fill_2 FILLER_24_270 ();
 sg13g2_fill_1 FILLER_24_284 ();
 sg13g2_fill_2 FILLER_24_309 ();
 sg13g2_fill_2 FILLER_24_421 ();
 sg13g2_fill_2 FILLER_24_427 ();
 sg13g2_fill_1 FILLER_24_429 ();
 sg13g2_fill_1 FILLER_25_28 ();
 sg13g2_fill_1 FILLER_25_45 ();
 sg13g2_fill_2 FILLER_25_52 ();
 sg13g2_fill_1 FILLER_25_54 ();
 sg13g2_fill_1 FILLER_25_71 ();
 sg13g2_fill_2 FILLER_25_80 ();
 sg13g2_fill_1 FILLER_25_86 ();
 sg13g2_fill_2 FILLER_25_103 ();
 sg13g2_fill_2 FILLER_25_125 ();
 sg13g2_fill_1 FILLER_25_127 ();
 sg13g2_fill_2 FILLER_25_134 ();
 sg13g2_fill_1 FILLER_25_164 ();
 sg13g2_fill_2 FILLER_25_169 ();
 sg13g2_fill_1 FILLER_25_175 ();
 sg13g2_fill_2 FILLER_25_180 ();
 sg13g2_fill_2 FILLER_25_198 ();
 sg13g2_fill_1 FILLER_25_204 ();
 sg13g2_fill_1 FILLER_25_233 ();
 sg13g2_fill_1 FILLER_25_250 ();
 sg13g2_fill_2 FILLER_25_327 ();
 sg13g2_fill_1 FILLER_25_381 ();
 sg13g2_fill_2 FILLER_25_406 ();
 sg13g2_fill_2 FILLER_25_416 ();
 sg13g2_fill_1 FILLER_25_418 ();
 sg13g2_fill_2 FILLER_25_427 ();
 sg13g2_fill_1 FILLER_25_429 ();
 sg13g2_fill_2 FILLER_26_4 ();
 sg13g2_fill_1 FILLER_26_12 ();
 sg13g2_fill_2 FILLER_26_33 ();
 sg13g2_fill_1 FILLER_26_35 ();
 sg13g2_fill_2 FILLER_26_136 ();
 sg13g2_fill_1 FILLER_26_138 ();
 sg13g2_fill_2 FILLER_26_147 ();
 sg13g2_fill_1 FILLER_26_197 ();
 sg13g2_fill_1 FILLER_26_242 ();
 sg13g2_fill_2 FILLER_26_247 ();
 sg13g2_fill_1 FILLER_26_249 ();
 sg13g2_fill_2 FILLER_26_262 ();
 sg13g2_fill_1 FILLER_26_290 ();
 sg13g2_fill_1 FILLER_26_299 ();
 sg13g2_fill_1 FILLER_26_316 ();
 sg13g2_fill_2 FILLER_26_333 ();
 sg13g2_fill_1 FILLER_26_379 ();
 sg13g2_fill_2 FILLER_26_408 ();
 sg13g2_fill_2 FILLER_27_8 ();
 sg13g2_fill_1 FILLER_27_18 ();
 sg13g2_fill_2 FILLER_27_51 ();
 sg13g2_fill_1 FILLER_27_57 ();
 sg13g2_fill_1 FILLER_27_90 ();
 sg13g2_fill_1 FILLER_27_99 ();
 sg13g2_fill_1 FILLER_27_104 ();
 sg13g2_fill_2 FILLER_27_137 ();
 sg13g2_fill_2 FILLER_27_155 ();
 sg13g2_fill_1 FILLER_27_161 ();
 sg13g2_fill_1 FILLER_27_190 ();
 sg13g2_fill_2 FILLER_27_203 ();
 sg13g2_fill_1 FILLER_27_205 ();
 sg13g2_fill_2 FILLER_27_214 ();
 sg13g2_fill_1 FILLER_27_216 ();
 sg13g2_fill_2 FILLER_27_237 ();
 sg13g2_fill_1 FILLER_27_251 ();
 sg13g2_fill_2 FILLER_27_268 ();
 sg13g2_fill_1 FILLER_27_316 ();
 sg13g2_fill_2 FILLER_27_357 ();
 sg13g2_fill_2 FILLER_27_403 ();
 sg13g2_fill_1 FILLER_27_429 ();
 sg13g2_fill_2 FILLER_28_0 ();
 sg13g2_fill_1 FILLER_28_22 ();
 sg13g2_fill_2 FILLER_28_51 ();
 sg13g2_fill_1 FILLER_28_57 ();
 sg13g2_fill_2 FILLER_28_74 ();
 sg13g2_fill_1 FILLER_28_96 ();
 sg13g2_fill_1 FILLER_28_129 ();
 sg13g2_fill_2 FILLER_28_166 ();
 sg13g2_fill_2 FILLER_28_188 ();
 sg13g2_fill_1 FILLER_28_226 ();
 sg13g2_fill_2 FILLER_28_247 ();
 sg13g2_fill_1 FILLER_28_249 ();
 sg13g2_fill_2 FILLER_28_282 ();
 sg13g2_fill_2 FILLER_28_288 ();
 sg13g2_fill_1 FILLER_28_290 ();
 sg13g2_fill_2 FILLER_28_311 ();
 sg13g2_fill_2 FILLER_28_345 ();
 sg13g2_fill_2 FILLER_28_363 ();
 sg13g2_fill_1 FILLER_28_373 ();
 sg13g2_fill_1 FILLER_28_378 ();
 sg13g2_fill_1 FILLER_28_403 ();
 sg13g2_fill_2 FILLER_28_428 ();
 sg13g2_fill_2 FILLER_29_0 ();
 sg13g2_fill_1 FILLER_29_6 ();
 sg13g2_fill_1 FILLER_29_23 ();
 sg13g2_fill_1 FILLER_29_44 ();
 sg13g2_fill_2 FILLER_29_57 ();
 sg13g2_fill_2 FILLER_29_95 ();
 sg13g2_fill_1 FILLER_29_125 ();
 sg13g2_fill_1 FILLER_29_130 ();
 sg13g2_fill_2 FILLER_29_143 ();
 sg13g2_fill_1 FILLER_29_145 ();
 sg13g2_fill_2 FILLER_29_158 ();
 sg13g2_fill_2 FILLER_29_180 ();
 sg13g2_fill_2 FILLER_29_222 ();
 sg13g2_fill_2 FILLER_29_256 ();
 sg13g2_fill_1 FILLER_29_258 ();
 sg13g2_fill_1 FILLER_29_329 ();
 sg13g2_fill_1 FILLER_29_382 ();
 sg13g2_fill_1 FILLER_29_403 ();
 sg13g2_fill_1 FILLER_29_408 ();
 sg13g2_fill_1 FILLER_29_429 ();
 sg13g2_fill_2 FILLER_30_0 ();
 sg13g2_fill_1 FILLER_30_2 ();
 sg13g2_fill_1 FILLER_30_19 ();
 sg13g2_fill_2 FILLER_30_24 ();
 sg13g2_fill_1 FILLER_30_54 ();
 sg13g2_fill_2 FILLER_30_71 ();
 sg13g2_fill_1 FILLER_30_101 ();
 sg13g2_fill_2 FILLER_30_118 ();
 sg13g2_fill_2 FILLER_30_140 ();
 sg13g2_fill_1 FILLER_30_142 ();
 sg13g2_fill_1 FILLER_30_207 ();
 sg13g2_fill_1 FILLER_30_212 ();
 sg13g2_fill_1 FILLER_30_221 ();
 sg13g2_fill_1 FILLER_30_226 ();
 sg13g2_fill_2 FILLER_30_231 ();
 sg13g2_fill_1 FILLER_30_233 ();
 sg13g2_fill_1 FILLER_30_330 ();
 sg13g2_fill_1 FILLER_30_343 ();
 sg13g2_fill_2 FILLER_30_396 ();
 sg13g2_fill_1 FILLER_30_414 ();
 sg13g2_fill_2 FILLER_30_427 ();
 sg13g2_fill_1 FILLER_30_429 ();
 sg13g2_fill_2 FILLER_31_0 ();
 sg13g2_fill_1 FILLER_31_2 ();
 sg13g2_fill_1 FILLER_31_47 ();
 sg13g2_fill_2 FILLER_31_52 ();
 sg13g2_fill_2 FILLER_31_96 ();
 sg13g2_fill_2 FILLER_31_110 ();
 sg13g2_fill_1 FILLER_31_132 ();
 sg13g2_fill_1 FILLER_31_193 ();
 sg13g2_fill_1 FILLER_31_218 ();
 sg13g2_fill_1 FILLER_31_235 ();
 sg13g2_fill_2 FILLER_31_248 ();
 sg13g2_fill_1 FILLER_31_254 ();
 sg13g2_fill_1 FILLER_31_271 ();
 sg13g2_fill_2 FILLER_31_276 ();
 sg13g2_fill_1 FILLER_31_378 ();
 sg13g2_fill_1 FILLER_31_409 ();
 sg13g2_fill_2 FILLER_32_0 ();
 sg13g2_fill_1 FILLER_32_2 ();
 sg13g2_fill_2 FILLER_32_23 ();
 sg13g2_fill_1 FILLER_32_25 ();
 sg13g2_fill_1 FILLER_32_98 ();
 sg13g2_fill_1 FILLER_32_103 ();
 sg13g2_fill_1 FILLER_32_120 ();
 sg13g2_fill_1 FILLER_32_125 ();
 sg13g2_fill_1 FILLER_32_158 ();
 sg13g2_fill_2 FILLER_32_177 ();
 sg13g2_fill_1 FILLER_32_191 ();
 sg13g2_fill_2 FILLER_32_220 ();
 sg13g2_fill_1 FILLER_32_222 ();
 sg13g2_fill_2 FILLER_32_227 ();
 sg13g2_fill_2 FILLER_32_269 ();
 sg13g2_fill_1 FILLER_32_271 ();
 sg13g2_fill_2 FILLER_32_288 ();
 sg13g2_fill_1 FILLER_32_290 ();
 sg13g2_fill_1 FILLER_32_359 ();
 sg13g2_fill_1 FILLER_32_372 ();
 sg13g2_fill_1 FILLER_32_429 ();
 sg13g2_fill_2 FILLER_33_28 ();
 sg13g2_fill_1 FILLER_33_30 ();
 sg13g2_fill_2 FILLER_33_179 ();
 sg13g2_fill_1 FILLER_33_181 ();
 sg13g2_fill_1 FILLER_33_186 ();
 sg13g2_fill_2 FILLER_33_211 ();
 sg13g2_fill_2 FILLER_33_241 ();
 sg13g2_fill_2 FILLER_33_327 ();
 sg13g2_fill_2 FILLER_33_397 ();
 sg13g2_fill_2 FILLER_33_427 ();
 sg13g2_fill_1 FILLER_33_429 ();
 sg13g2_fill_2 FILLER_34_8 ();
 sg13g2_fill_1 FILLER_34_10 ();
 sg13g2_fill_1 FILLER_34_31 ();
 sg13g2_fill_2 FILLER_34_40 ();
 sg13g2_fill_2 FILLER_34_110 ();
 sg13g2_fill_2 FILLER_34_116 ();
 sg13g2_fill_2 FILLER_34_158 ();
 sg13g2_fill_1 FILLER_34_160 ();
 sg13g2_fill_2 FILLER_34_173 ();
 sg13g2_fill_1 FILLER_34_175 ();
 sg13g2_fill_2 FILLER_34_208 ();
 sg13g2_fill_1 FILLER_34_230 ();
 sg13g2_fill_1 FILLER_34_239 ();
 sg13g2_fill_1 FILLER_34_244 ();
 sg13g2_fill_1 FILLER_34_249 ();
 sg13g2_fill_1 FILLER_34_258 ();
 sg13g2_fill_2 FILLER_34_267 ();
 sg13g2_fill_1 FILLER_34_269 ();
 sg13g2_fill_2 FILLER_35_32 ();
 sg13g2_fill_2 FILLER_35_102 ();
 sg13g2_fill_2 FILLER_35_184 ();
 sg13g2_fill_2 FILLER_35_202 ();
 sg13g2_fill_1 FILLER_35_208 ();
 sg13g2_fill_2 FILLER_35_377 ();
 sg13g2_fill_1 FILLER_35_379 ();
 sg13g2_fill_1 FILLER_35_404 ();
 sg13g2_fill_1 FILLER_35_429 ();
 sg13g2_fill_1 FILLER_36_4 ();
 sg13g2_fill_2 FILLER_36_9 ();
 sg13g2_fill_1 FILLER_36_23 ();
 sg13g2_fill_1 FILLER_36_156 ();
 sg13g2_fill_1 FILLER_36_213 ();
 sg13g2_fill_2 FILLER_36_282 ();
 sg13g2_fill_2 FILLER_36_352 ();
 sg13g2_fill_1 FILLER_36_378 ();
 sg13g2_fill_1 FILLER_36_383 ();
 sg13g2_fill_1 FILLER_36_404 ();
 sg13g2_fill_2 FILLER_36_409 ();
 sg13g2_fill_1 FILLER_36_423 ();
 sg13g2_fill_2 FILLER_36_428 ();
 sg13g2_fill_2 FILLER_37_0 ();
 sg13g2_fill_1 FILLER_37_2 ();
 sg13g2_fill_1 FILLER_37_11 ();
 sg13g2_fill_2 FILLER_37_24 ();
 sg13g2_fill_2 FILLER_37_44 ();
 sg13g2_fill_2 FILLER_37_214 ();
 sg13g2_fill_1 FILLER_37_216 ();
 sg13g2_fill_2 FILLER_37_427 ();
 sg13g2_fill_1 FILLER_37_429 ();
 sg13g2_fill_2 FILLER_38_0 ();
 sg13g2_fill_2 FILLER_38_12 ();
 sg13g2_fill_1 FILLER_38_210 ();
 sg13g2_fill_1 FILLER_38_215 ();
 sg13g2_fill_1 FILLER_38_224 ();
 sg13g2_fill_2 FILLER_38_253 ();
 sg13g2_fill_2 FILLER_38_307 ();
 sg13g2_fill_2 FILLER_38_421 ();
 sg13g2_fill_1 FILLER_38_423 ();
endmodule
