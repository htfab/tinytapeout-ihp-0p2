module tt_um_brandonramos_VGA_Pong_with_NES_Controllers (clk,
    ena,
    rst_n,
    ui_in,
    uio_in,
    uio_oe,
    uio_out,
    uo_out);
 input clk;
 input ena;
 input rst_n;
 input [7:0] ui_in;
 input [7:0] uio_in;
 output [7:0] uio_oe;
 output [7:0] uio_out;
 output [7:0] uo_out;

 wire \Pong.b ;
 wire \Pong.control_unit.NES_Controller_Left.state_NESController[0] ;
 wire \Pong.control_unit.NES_Controller_Left.state_NESController[10] ;
 wire \Pong.control_unit.NES_Controller_Left.state_NESController[11] ;
 wire \Pong.control_unit.NES_Controller_Left.state_NESController[12] ;
 wire \Pong.control_unit.NES_Controller_Left.state_NESController[13] ;
 wire \Pong.control_unit.NES_Controller_Left.state_NESController[14] ;
 wire \Pong.control_unit.NES_Controller_Left.state_NESController[15] ;
 wire \Pong.control_unit.NES_Controller_Left.state_NESController[16] ;
 wire \Pong.control_unit.NES_Controller_Left.state_NESController[17] ;
 wire \Pong.control_unit.NES_Controller_Left.state_NESController[18] ;
 wire \Pong.control_unit.NES_Controller_Left.state_NESController[1] ;
 wire \Pong.control_unit.NES_Controller_Left.state_NESController[2] ;
 wire \Pong.control_unit.NES_Controller_Left.state_NESController[3] ;
 wire \Pong.control_unit.NES_Controller_Left.state_NESController[4] ;
 wire \Pong.control_unit.NES_Controller_Left.state_NESController[5] ;
 wire \Pong.control_unit.NES_Controller_Left.state_NESController[6] ;
 wire \Pong.control_unit.NES_Controller_Left.state_NESController[7] ;
 wire \Pong.control_unit.NES_Controller_Left.state_NESController[8] ;
 wire \Pong.control_unit.NES_Controller_Left.state_NESController[9] ;
 wire \Pong.control_unit.NES_Controller_Right.state_NESController[0] ;
 wire \Pong.control_unit.NES_Controller_Right.state_NESController[10] ;
 wire \Pong.control_unit.NES_Controller_Right.state_NESController[11] ;
 wire \Pong.control_unit.NES_Controller_Right.state_NESController[12] ;
 wire \Pong.control_unit.NES_Controller_Right.state_NESController[13] ;
 wire \Pong.control_unit.NES_Controller_Right.state_NESController[14] ;
 wire \Pong.control_unit.NES_Controller_Right.state_NESController[15] ;
 wire \Pong.control_unit.NES_Controller_Right.state_NESController[16] ;
 wire \Pong.control_unit.NES_Controller_Right.state_NESController[17] ;
 wire \Pong.control_unit.NES_Controller_Right.state_NESController[18] ;
 wire \Pong.control_unit.NES_Controller_Right.state_NESController[1] ;
 wire \Pong.control_unit.NES_Controller_Right.state_NESController[2] ;
 wire \Pong.control_unit.NES_Controller_Right.state_NESController[3] ;
 wire \Pong.control_unit.NES_Controller_Right.state_NESController[4] ;
 wire \Pong.control_unit.NES_Controller_Right.state_NESController[5] ;
 wire \Pong.control_unit.NES_Controller_Right.state_NESController[6] ;
 wire \Pong.control_unit.NES_Controller_Right.state_NESController[7] ;
 wire \Pong.control_unit.NES_Controller_Right.state_NESController[8] ;
 wire \Pong.control_unit.NES_Controller_Right.state_NESController[9] ;
 wire \Pong.control_unit.state_ballMovement[0] ;
 wire \Pong.control_unit.state_ballMovement[1] ;
 wire \Pong.control_unit.state_ballMovement[2] ;
 wire \Pong.control_unit.state_ballMovement[3] ;
 wire \Pong.control_unit.state_ballMovement[4] ;
 wire \Pong.datapath.Ball_Clock.Q[0] ;
 wire \Pong.datapath.Ball_Clock.Q[10] ;
 wire \Pong.datapath.Ball_Clock.Q[11] ;
 wire \Pong.datapath.Ball_Clock.Q[12] ;
 wire \Pong.datapath.Ball_Clock.Q[13] ;
 wire \Pong.datapath.Ball_Clock.Q[14] ;
 wire \Pong.datapath.Ball_Clock.Q[15] ;
 wire \Pong.datapath.Ball_Clock.Q[16] ;
 wire \Pong.datapath.Ball_Clock.Q[1] ;
 wire \Pong.datapath.Ball_Clock.Q[2] ;
 wire \Pong.datapath.Ball_Clock.Q[3] ;
 wire \Pong.datapath.Ball_Clock.Q[4] ;
 wire \Pong.datapath.Ball_Clock.Q[5] ;
 wire \Pong.datapath.Ball_Clock.Q[6] ;
 wire \Pong.datapath.Ball_Clock.Q[7] ;
 wire \Pong.datapath.Ball_Clock.Q[8] ;
 wire \Pong.datapath.Ball_Clock.Q[9] ;
 wire \Pong.datapath.Ball_Clock.roll ;
 wire \Pong.datapath.NES_activity_Left[2] ;
 wire \Pong.datapath.NES_activity_Left[3] ;
 wire \Pong.datapath.NES_activity_Left[4] ;
 wire \Pong.datapath.NES_activity_Left[5] ;
 wire \Pong.datapath.NES_activity_Right[2] ;
 wire \Pong.datapath.NES_activity_Right[3] ;
 wire \Pong.datapath.NES_activity_Right[4] ;
 wire \Pong.datapath.NES_activity_Right[5] ;
 wire \Pong.datapath.NES_counter_left.Q[0] ;
 wire \Pong.datapath.NES_counter_left.Q[1] ;
 wire \Pong.datapath.NES_counter_left.Q[2] ;
 wire \Pong.datapath.NES_counter_left.Q[3] ;
 wire \Pong.datapath.NES_counter_left.Q[4] ;
 wire \Pong.datapath.NES_counter_left.Q[5] ;
 wire \Pong.datapath.NES_counter_left.Q[6] ;
 wire \Pong.datapath.NES_counter_left.Q[7] ;
 wire \Pong.datapath.NES_counter_right.Q[0] ;
 wire \Pong.datapath.NES_counter_right.Q[1] ;
 wire \Pong.datapath.NES_counter_right.Q[2] ;
 wire \Pong.datapath.NES_counter_right.Q[3] ;
 wire \Pong.datapath.NES_counter_right.Q[4] ;
 wire \Pong.datapath.NES_counter_right.Q[5] ;
 wire \Pong.datapath.NES_counter_right.Q[6] ;
 wire \Pong.datapath.NES_counter_right.Q[7] ;
 wire \Pong.datapath.NES_delay_counter_left.Q[0] ;
 wire \Pong.datapath.NES_delay_counter_left.Q[10] ;
 wire \Pong.datapath.NES_delay_counter_left.Q[11] ;
 wire \Pong.datapath.NES_delay_counter_left.Q[12] ;
 wire \Pong.datapath.NES_delay_counter_left.Q[13] ;
 wire \Pong.datapath.NES_delay_counter_left.Q[14] ;
 wire \Pong.datapath.NES_delay_counter_left.Q[15] ;
 wire \Pong.datapath.NES_delay_counter_left.Q[16] ;
 wire \Pong.datapath.NES_delay_counter_left.Q[17] ;
 wire \Pong.datapath.NES_delay_counter_left.Q[18] ;
 wire \Pong.datapath.NES_delay_counter_left.Q[1] ;
 wire \Pong.datapath.NES_delay_counter_left.Q[2] ;
 wire \Pong.datapath.NES_delay_counter_left.Q[3] ;
 wire \Pong.datapath.NES_delay_counter_left.Q[4] ;
 wire \Pong.datapath.NES_delay_counter_left.Q[5] ;
 wire \Pong.datapath.NES_delay_counter_left.Q[6] ;
 wire \Pong.datapath.NES_delay_counter_left.Q[7] ;
 wire \Pong.datapath.NES_delay_counter_left.Q[8] ;
 wire \Pong.datapath.NES_delay_counter_left.Q[9] ;
 wire \Pong.datapath.NES_delay_counter_right.Q[0] ;
 wire \Pong.datapath.NES_delay_counter_right.Q[10] ;
 wire \Pong.datapath.NES_delay_counter_right.Q[11] ;
 wire \Pong.datapath.NES_delay_counter_right.Q[12] ;
 wire \Pong.datapath.NES_delay_counter_right.Q[13] ;
 wire \Pong.datapath.NES_delay_counter_right.Q[14] ;
 wire \Pong.datapath.NES_delay_counter_right.Q[15] ;
 wire \Pong.datapath.NES_delay_counter_right.Q[16] ;
 wire \Pong.datapath.NES_delay_counter_right.Q[17] ;
 wire \Pong.datapath.NES_delay_counter_right.Q[18] ;
 wire \Pong.datapath.NES_delay_counter_right.Q[1] ;
 wire \Pong.datapath.NES_delay_counter_right.Q[2] ;
 wire \Pong.datapath.NES_delay_counter_right.Q[3] ;
 wire \Pong.datapath.NES_delay_counter_right.Q[4] ;
 wire \Pong.datapath.NES_delay_counter_right.Q[5] ;
 wire \Pong.datapath.NES_delay_counter_right.Q[6] ;
 wire \Pong.datapath.NES_delay_counter_right.Q[7] ;
 wire \Pong.datapath.NES_delay_counter_right.Q[8] ;
 wire \Pong.datapath.NES_delay_counter_right.Q[9] ;
 wire \Pong.datapath.NES_wire_Left[2] ;
 wire \Pong.datapath.NES_wire_Left[3] ;
 wire \Pong.datapath.NES_wire_Left[4] ;
 wire \Pong.datapath.NES_wire_Left[5] ;
 wire \Pong.datapath.NES_wire_Right[2] ;
 wire \Pong.datapath.NES_wire_Right[3] ;
 wire \Pong.datapath.NES_wire_Right[4] ;
 wire \Pong.datapath.NES_wire_Right[5] ;
 wire \Pong.datapath.ballFunction.ball_center_x[0] ;
 wire \Pong.datapath.ballFunction.ball_center_x[1] ;
 wire \Pong.datapath.ballFunction.ball_center_x[2] ;
 wire \Pong.datapath.ballFunction.ball_center_x[3] ;
 wire \Pong.datapath.ballFunction.ball_center_x[4] ;
 wire \Pong.datapath.ballFunction.ball_center_x[5] ;
 wire \Pong.datapath.ballFunction.ball_center_x[6] ;
 wire \Pong.datapath.ballFunction.ball_center_x[7] ;
 wire \Pong.datapath.ballFunction.ball_center_x[8] ;
 wire \Pong.datapath.ballFunction.ball_center_x[9] ;
 wire \Pong.datapath.ballFunction.ball_center_y[0] ;
 wire \Pong.datapath.ballFunction.ball_center_y[1] ;
 wire \Pong.datapath.ballFunction.ball_center_y[2] ;
 wire \Pong.datapath.ballFunction.ball_center_y[3] ;
 wire \Pong.datapath.ballFunction.ball_center_y[4] ;
 wire \Pong.datapath.ballFunction.ball_center_y[5] ;
 wire \Pong.datapath.ballFunction.ball_center_y[6] ;
 wire \Pong.datapath.ballFunction.ball_center_y[7] ;
 wire \Pong.datapath.ballFunction.ball_center_y[8] ;
 wire \Pong.datapath.ballFunction.ball_center_y[9] ;
 wire \Pong.datapath.ballFunction.reset_n ;
 wire \Pong.datapath.h_sync ;
 wire \Pong.datapath.leftPaddle[0] ;
 wire \Pong.datapath.leftPaddle[1] ;
 wire \Pong.datapath.leftPaddle[2] ;
 wire \Pong.datapath.leftPaddle[3] ;
 wire \Pong.datapath.leftPaddle[4] ;
 wire \Pong.datapath.leftPaddle[5] ;
 wire \Pong.datapath.leftPaddle[6] ;
 wire \Pong.datapath.leftPaddle[7] ;
 wire \Pong.datapath.leftPaddle[8] ;
 wire \Pong.datapath.leftPaddle[9] ;
 wire \Pong.datapath.old_NES_Left[2] ;
 wire \Pong.datapath.old_NES_Left[3] ;
 wire \Pong.datapath.old_NES_Left[4] ;
 wire \Pong.datapath.old_NES_Left[5] ;
 wire \Pong.datapath.old_NES_Right[2] ;
 wire \Pong.datapath.old_NES_Right[3] ;
 wire \Pong.datapath.old_NES_Right[4] ;
 wire \Pong.datapath.old_NES_Right[5] ;
 wire \Pong.datapath.rightPaddle[0] ;
 wire \Pong.datapath.rightPaddle[1] ;
 wire \Pong.datapath.rightPaddle[2] ;
 wire \Pong.datapath.rightPaddle[3] ;
 wire \Pong.datapath.rightPaddle[4] ;
 wire \Pong.datapath.rightPaddle[5] ;
 wire \Pong.datapath.rightPaddle[6] ;
 wire \Pong.datapath.rightPaddle[7] ;
 wire \Pong.datapath.rightPaddle[8] ;
 wire \Pong.datapath.rightPaddle[9] ;
 wire \Pong.datapath.scoreLeft[0] ;
 wire \Pong.datapath.scoreLeft[1] ;
 wire \Pong.datapath.scoreLeft[2] ;
 wire \Pong.datapath.scoreLeft[3] ;
 wire \Pong.datapath.scoreRight[0] ;
 wire \Pong.datapath.scoreRight[1] ;
 wire \Pong.datapath.scoreRight[2] ;
 wire \Pong.datapath.scoreRight[3] ;
 wire \Pong.datapath.score_flag ;
 wire \Pong.datapath.sw_ballMovement_reg[0] ;
 wire \Pong.datapath.sw_ballMovement_reg[2] ;
 wire \Pong.datapath.sw_ballMovement_reg[3] ;
 wire \Pong.datapath.sw_ballMovement_reg[4] ;
 wire \Pong.datapath.sw_ballMovement_reg[5] ;
 wire \Pong.datapath.v_sync ;
 wire \Pong.datapath.vga.Column_Counter.Q[0] ;
 wire \Pong.datapath.vga.Column_Counter.Q[1] ;
 wire \Pong.datapath.vga.Column_Counter.Q[2] ;
 wire \Pong.datapath.vga.Column_Counter.Q[3] ;
 wire \Pong.datapath.vga.Column_Counter.Q[4] ;
 wire \Pong.datapath.vga.Column_Counter.Q[5] ;
 wire \Pong.datapath.vga.Column_Counter.Q[6] ;
 wire \Pong.datapath.vga.Column_Counter.Q[7] ;
 wire \Pong.datapath.vga.Column_Counter.Q[8] ;
 wire \Pong.datapath.vga.Column_Counter.Q[9] ;
 wire \Pong.datapath.vga.Row_Counter.Q[0] ;
 wire \Pong.datapath.vga.Row_Counter.Q[1] ;
 wire \Pong.datapath.vga.Row_Counter.Q[2] ;
 wire \Pong.datapath.vga.Row_Counter.Q[3] ;
 wire \Pong.datapath.vga.Row_Counter.Q[4] ;
 wire \Pong.datapath.vga.Row_Counter.Q[5] ;
 wire \Pong.datapath.vga.Row_Counter.Q[6] ;
 wire \Pong.datapath.vga.Row_Counter.Q[7] ;
 wire \Pong.datapath.vga.Row_Counter.Q[8] ;
 wire \Pong.datapath.vga.Row_Counter.Q[9] ;
 wire _0000_;
 wire _0001_;
 wire _0002_;
 wire _0003_;
 wire _0004_;
 wire _0005_;
 wire _0006_;
 wire _0007_;
 wire _0008_;
 wire _0009_;
 wire _0010_;
 wire _0011_;
 wire _0012_;
 wire _0013_;
 wire _0014_;
 wire _0015_;
 wire _0016_;
 wire _0017_;
 wire _0018_;
 wire _0019_;
 wire _0020_;
 wire _0021_;
 wire _0022_;
 wire _0023_;
 wire _0024_;
 wire _0025_;
 wire _0026_;
 wire _0027_;
 wire _0028_;
 wire _0029_;
 wire _0030_;
 wire _0031_;
 wire _0032_;
 wire _0033_;
 wire _0034_;
 wire _0035_;
 wire _0036_;
 wire _0037_;
 wire _0038_;
 wire _0039_;
 wire _0040_;
 wire _0041_;
 wire _0042_;
 wire _0043_;
 wire _0044_;
 wire _0045_;
 wire _0046_;
 wire _0047_;
 wire _0048_;
 wire _0049_;
 wire _0050_;
 wire _0051_;
 wire _0052_;
 wire _0053_;
 wire _0054_;
 wire _0055_;
 wire _0056_;
 wire _0057_;
 wire _0058_;
 wire _0059_;
 wire _0060_;
 wire _0061_;
 wire _0062_;
 wire _0063_;
 wire _0064_;
 wire _0065_;
 wire _0066_;
 wire _0067_;
 wire _0068_;
 wire _0069_;
 wire _0070_;
 wire _0071_;
 wire _0072_;
 wire _0073_;
 wire _0074_;
 wire _0075_;
 wire _0076_;
 wire _0077_;
 wire _0078_;
 wire _0079_;
 wire _0080_;
 wire _0081_;
 wire _0082_;
 wire _0083_;
 wire _0084_;
 wire _0085_;
 wire _0086_;
 wire _0087_;
 wire _0088_;
 wire _0089_;
 wire _0090_;
 wire _0091_;
 wire _0092_;
 wire _0093_;
 wire _0094_;
 wire _0095_;
 wire _0096_;
 wire _0097_;
 wire _0098_;
 wire _0099_;
 wire _0100_;
 wire _0101_;
 wire _0102_;
 wire _0103_;
 wire _0104_;
 wire _0105_;
 wire _0106_;
 wire _0107_;
 wire _0108_;
 wire _0109_;
 wire _0110_;
 wire _0111_;
 wire _0112_;
 wire _0113_;
 wire _0114_;
 wire _0115_;
 wire _0116_;
 wire _0117_;
 wire _0118_;
 wire _0119_;
 wire _0120_;
 wire _0121_;
 wire _0122_;
 wire _0123_;
 wire _0124_;
 wire _0125_;
 wire _0126_;
 wire _0127_;
 wire _0128_;
 wire _0129_;
 wire _0130_;
 wire _0131_;
 wire _0132_;
 wire _0133_;
 wire _0134_;
 wire _0135_;
 wire _0136_;
 wire _0137_;
 wire _0138_;
 wire _0139_;
 wire _0140_;
 wire _0141_;
 wire _0142_;
 wire _0143_;
 wire _0144_;
 wire _0145_;
 wire _0146_;
 wire _0147_;
 wire _0148_;
 wire _0149_;
 wire _0150_;
 wire _0151_;
 wire _0152_;
 wire _0153_;
 wire _0154_;
 wire _0155_;
 wire _0156_;
 wire _0157_;
 wire _0158_;
 wire _0159_;
 wire _0160_;
 wire _0161_;
 wire _0162_;
 wire _0163_;
 wire _0164_;
 wire _0165_;
 wire _0166_;
 wire _0167_;
 wire _0168_;
 wire _0169_;
 wire _0170_;
 wire _0171_;
 wire _0172_;
 wire _0173_;
 wire _0174_;
 wire _0175_;
 wire _0176_;
 wire _0177_;
 wire _0178_;
 wire _0179_;
 wire _0180_;
 wire _0181_;
 wire _0182_;
 wire _0183_;
 wire _0184_;
 wire _0185_;
 wire _0186_;
 wire _0187_;
 wire _0188_;
 wire _0189_;
 wire _0190_;
 wire _0191_;
 wire _0192_;
 wire _0193_;
 wire _0194_;
 wire _0195_;
 wire _0196_;
 wire _0197_;
 wire _0198_;
 wire _0199_;
 wire _0200_;
 wire _0201_;
 wire _0202_;
 wire _0203_;
 wire _0204_;
 wire _0205_;
 wire _0206_;
 wire _0207_;
 wire _0208_;
 wire _0209_;
 wire _0210_;
 wire _0211_;
 wire _0212_;
 wire _0213_;
 wire _0214_;
 wire _0215_;
 wire _0216_;
 wire _0217_;
 wire _0218_;
 wire _0219_;
 wire _0220_;
 wire _0221_;
 wire _0222_;
 wire _0223_;
 wire _0224_;
 wire _0225_;
 wire _0226_;
 wire _0227_;
 wire _0228_;
 wire _0229_;
 wire _0230_;
 wire _0231_;
 wire _0232_;
 wire _0233_;
 wire _0234_;
 wire _0235_;
 wire _0236_;
 wire _0237_;
 wire _0238_;
 wire _0239_;
 wire _0240_;
 wire _0241_;
 wire _0242_;
 wire _0243_;
 wire _0244_;
 wire _0245_;
 wire _0246_;
 wire _0247_;
 wire _0248_;
 wire _0249_;
 wire _0250_;
 wire _0251_;
 wire _0252_;
 wire _0253_;
 wire _0254_;
 wire _0255_;
 wire _0256_;
 wire _0257_;
 wire _0258_;
 wire _0259_;
 wire _0260_;
 wire _0261_;
 wire _0262_;
 wire _0263_;
 wire _0264_;
 wire _0265_;
 wire _0266_;
 wire _0267_;
 wire _0268_;
 wire _0269_;
 wire _0270_;
 wire _0271_;
 wire _0272_;
 wire _0273_;
 wire _0274_;
 wire _0275_;
 wire _0276_;
 wire _0277_;
 wire _0278_;
 wire _0279_;
 wire _0280_;
 wire _0281_;
 wire _0282_;
 wire _0283_;
 wire _0284_;
 wire _0285_;
 wire _0286_;
 wire _0287_;
 wire _0288_;
 wire _0289_;
 wire _0290_;
 wire _0291_;
 wire _0292_;
 wire _0293_;
 wire _0294_;
 wire _0295_;
 wire _0296_;
 wire _0297_;
 wire _0298_;
 wire _0299_;
 wire _0300_;
 wire _0301_;
 wire _0302_;
 wire _0303_;
 wire _0304_;
 wire _0305_;
 wire _0306_;
 wire _0307_;
 wire _0308_;
 wire _0309_;
 wire _0310_;
 wire _0311_;
 wire _0312_;
 wire _0313_;
 wire _0314_;
 wire _0315_;
 wire _0316_;
 wire _0317_;
 wire _0318_;
 wire _0319_;
 wire _0320_;
 wire _0321_;
 wire _0322_;
 wire _0323_;
 wire _0324_;
 wire _0325_;
 wire _0326_;
 wire _0327_;
 wire _0328_;
 wire _0329_;
 wire _0330_;
 wire _0331_;
 wire _0332_;
 wire _0333_;
 wire _0334_;
 wire _0335_;
 wire _0336_;
 wire _0337_;
 wire _0338_;
 wire _0339_;
 wire _0340_;
 wire _0341_;
 wire _0342_;
 wire _0343_;
 wire _0344_;
 wire _0345_;
 wire _0346_;
 wire _0347_;
 wire _0348_;
 wire _0349_;
 wire _0350_;
 wire _0351_;
 wire _0352_;
 wire _0353_;
 wire _0354_;
 wire _0355_;
 wire _0356_;
 wire _0357_;
 wire _0358_;
 wire _0359_;
 wire _0360_;
 wire _0361_;
 wire _0362_;
 wire _0363_;
 wire _0364_;
 wire _0365_;
 wire _0366_;
 wire _0367_;
 wire _0368_;
 wire _0369_;
 wire _0370_;
 wire _0371_;
 wire _0372_;
 wire _0373_;
 wire _0374_;
 wire _0375_;
 wire _0376_;
 wire _0377_;
 wire _0378_;
 wire _0379_;
 wire _0380_;
 wire _0381_;
 wire _0382_;
 wire _0383_;
 wire _0384_;
 wire _0385_;
 wire _0386_;
 wire _0387_;
 wire _0388_;
 wire _0389_;
 wire _0390_;
 wire _0391_;
 wire _0392_;
 wire _0393_;
 wire _0394_;
 wire _0395_;
 wire _0396_;
 wire _0397_;
 wire _0398_;
 wire _0399_;
 wire _0400_;
 wire _0401_;
 wire _0402_;
 wire _0403_;
 wire _0404_;
 wire _0405_;
 wire _0406_;
 wire _0407_;
 wire _0408_;
 wire _0409_;
 wire _0410_;
 wire _0411_;
 wire _0412_;
 wire _0413_;
 wire _0414_;
 wire _0415_;
 wire _0416_;
 wire _0417_;
 wire _0418_;
 wire _0419_;
 wire _0420_;
 wire _0421_;
 wire _0422_;
 wire _0423_;
 wire _0424_;
 wire _0425_;
 wire _0426_;
 wire _0427_;
 wire _0428_;
 wire _0429_;
 wire _0430_;
 wire _0431_;
 wire _0432_;
 wire _0433_;
 wire _0434_;
 wire _0435_;
 wire _0436_;
 wire _0437_;
 wire _0438_;
 wire _0439_;
 wire _0440_;
 wire _0441_;
 wire _0442_;
 wire _0443_;
 wire _0444_;
 wire _0445_;
 wire _0446_;
 wire _0447_;
 wire _0448_;
 wire _0449_;
 wire _0450_;
 wire _0451_;
 wire _0452_;
 wire _0453_;
 wire _0454_;
 wire _0455_;
 wire _0456_;
 wire _0457_;
 wire _0458_;
 wire _0459_;
 wire _0460_;
 wire _0461_;
 wire _0462_;
 wire _0463_;
 wire _0464_;
 wire _0465_;
 wire _0466_;
 wire _0467_;
 wire _0468_;
 wire _0469_;
 wire _0470_;
 wire _0471_;
 wire _0472_;
 wire _0473_;
 wire _0474_;
 wire _0475_;
 wire _0476_;
 wire _0477_;
 wire _0478_;
 wire _0479_;
 wire _0480_;
 wire _0481_;
 wire _0482_;
 wire _0483_;
 wire _0484_;
 wire _0485_;
 wire _0486_;
 wire _0487_;
 wire _0488_;
 wire _0489_;
 wire _0490_;
 wire _0491_;
 wire _0492_;
 wire _0493_;
 wire _0494_;
 wire _0495_;
 wire _0496_;
 wire _0497_;
 wire _0498_;
 wire _0499_;
 wire _0500_;
 wire _0501_;
 wire _0502_;
 wire _0503_;
 wire _0504_;
 wire _0505_;
 wire _0506_;
 wire _0507_;
 wire _0508_;
 wire _0509_;
 wire _0510_;
 wire _0511_;
 wire _0512_;
 wire _0513_;
 wire _0514_;
 wire _0515_;
 wire _0516_;
 wire _0517_;
 wire _0518_;
 wire _0519_;
 wire _0520_;
 wire _0521_;
 wire _0522_;
 wire _0523_;
 wire _0524_;
 wire _0525_;
 wire _0526_;
 wire _0527_;
 wire _0528_;
 wire _0529_;
 wire _0530_;
 wire _0531_;
 wire _0532_;
 wire _0533_;
 wire _0534_;
 wire _0535_;
 wire _0536_;
 wire _0537_;
 wire _0538_;
 wire _0539_;
 wire _0540_;
 wire _0541_;
 wire _0542_;
 wire _0543_;
 wire _0544_;
 wire _0545_;
 wire _0546_;
 wire _0547_;
 wire _0548_;
 wire _0549_;
 wire _0550_;
 wire _0551_;
 wire _0552_;
 wire _0553_;
 wire _0554_;
 wire _0555_;
 wire _0556_;
 wire _0557_;
 wire _0558_;
 wire _0559_;
 wire _0560_;
 wire _0561_;
 wire _0562_;
 wire _0563_;
 wire _0564_;
 wire _0565_;
 wire _0566_;
 wire _0567_;
 wire _0568_;
 wire _0569_;
 wire _0570_;
 wire _0571_;
 wire _0572_;
 wire _0573_;
 wire _0574_;
 wire _0575_;
 wire _0576_;
 wire _0577_;
 wire _0578_;
 wire _0579_;
 wire _0580_;
 wire _0581_;
 wire _0582_;
 wire _0583_;
 wire _0584_;
 wire _0585_;
 wire _0586_;
 wire _0587_;
 wire _0588_;
 wire _0589_;
 wire _0590_;
 wire _0591_;
 wire _0592_;
 wire _0593_;
 wire _0594_;
 wire _0595_;
 wire _0596_;
 wire _0597_;
 wire _0598_;
 wire _0599_;
 wire _0600_;
 wire _0601_;
 wire _0602_;
 wire _0603_;
 wire _0604_;
 wire _0605_;
 wire _0606_;
 wire _0607_;
 wire _0608_;
 wire _0609_;
 wire _0610_;
 wire _0611_;
 wire _0612_;
 wire _0613_;
 wire _0614_;
 wire _0615_;
 wire _0616_;
 wire _0617_;
 wire _0618_;
 wire _0619_;
 wire _0620_;
 wire _0621_;
 wire _0622_;
 wire _0623_;
 wire _0624_;
 wire _0625_;
 wire _0626_;
 wire _0627_;
 wire _0628_;
 wire _0629_;
 wire _0630_;
 wire _0631_;
 wire _0632_;
 wire _0633_;
 wire _0634_;
 wire _0635_;
 wire _0636_;
 wire _0637_;
 wire _0638_;
 wire _0639_;
 wire _0640_;
 wire _0641_;
 wire _0642_;
 wire _0643_;
 wire _0644_;
 wire _0645_;
 wire _0646_;
 wire _0647_;
 wire _0648_;
 wire _0649_;
 wire _0650_;
 wire _0651_;
 wire _0652_;
 wire _0653_;
 wire _0654_;
 wire _0655_;
 wire _0656_;
 wire _0657_;
 wire _0658_;
 wire _0659_;
 wire _0660_;
 wire _0661_;
 wire _0662_;
 wire _0663_;
 wire _0664_;
 wire _0665_;
 wire _0666_;
 wire _0667_;
 wire _0668_;
 wire _0669_;
 wire _0670_;
 wire _0671_;
 wire _0672_;
 wire _0673_;
 wire _0674_;
 wire _0675_;
 wire _0676_;
 wire _0677_;
 wire _0678_;
 wire _0679_;
 wire _0680_;
 wire _0681_;
 wire _0682_;
 wire _0683_;
 wire _0684_;
 wire _0685_;
 wire _0686_;
 wire _0687_;
 wire _0688_;
 wire _0689_;
 wire _0690_;
 wire _0691_;
 wire _0692_;
 wire _0693_;
 wire _0694_;
 wire _0695_;
 wire _0696_;
 wire _0697_;
 wire _0698_;
 wire _0699_;
 wire _0700_;
 wire _0701_;
 wire _0702_;
 wire _0703_;
 wire _0704_;
 wire _0705_;
 wire _0706_;
 wire _0707_;
 wire _0708_;
 wire _0709_;
 wire _0710_;
 wire _0711_;
 wire _0712_;
 wire _0713_;
 wire _0714_;
 wire _0715_;
 wire _0716_;
 wire _0717_;
 wire _0718_;
 wire _0719_;
 wire _0720_;
 wire _0721_;
 wire _0722_;
 wire _0723_;
 wire _0724_;
 wire _0725_;
 wire _0726_;
 wire _0727_;
 wire _0728_;
 wire _0729_;
 wire _0730_;
 wire _0731_;
 wire _0732_;
 wire _0733_;
 wire _0734_;
 wire _0735_;
 wire _0736_;
 wire _0737_;
 wire _0738_;
 wire _0739_;
 wire _0740_;
 wire _0741_;
 wire _0742_;
 wire _0743_;
 wire _0744_;
 wire _0745_;
 wire _0746_;
 wire _0747_;
 wire _0748_;
 wire _0749_;
 wire _0750_;
 wire _0751_;
 wire _0752_;
 wire _0753_;
 wire _0754_;
 wire _0755_;
 wire _0756_;
 wire _0757_;
 wire _0758_;
 wire _0759_;
 wire _0760_;
 wire _0761_;
 wire _0762_;
 wire _0763_;
 wire _0764_;
 wire _0765_;
 wire _0766_;
 wire _0767_;
 wire _0768_;
 wire _0769_;
 wire _0770_;
 wire _0771_;
 wire _0772_;
 wire _0773_;
 wire _0774_;
 wire _0775_;
 wire _0776_;
 wire _0777_;
 wire _0778_;
 wire _0779_;
 wire _0780_;
 wire _0781_;
 wire _0782_;
 wire _0783_;
 wire _0784_;
 wire _0785_;
 wire _0786_;
 wire _0787_;
 wire _0788_;
 wire _0789_;
 wire _0790_;
 wire _0791_;
 wire _0792_;
 wire _0793_;
 wire _0794_;
 wire _0795_;
 wire _0796_;
 wire _0797_;
 wire _0798_;
 wire _0799_;
 wire _0800_;
 wire _0801_;
 wire _0802_;
 wire _0803_;
 wire _0804_;
 wire _0805_;
 wire _0806_;
 wire _0807_;
 wire _0808_;
 wire _0809_;
 wire _0810_;
 wire _0811_;
 wire _0812_;
 wire _0813_;
 wire _0814_;
 wire _0815_;
 wire _0816_;
 wire _0817_;
 wire _0818_;
 wire _0819_;
 wire _0820_;
 wire _0821_;
 wire _0822_;
 wire _0823_;
 wire _0824_;
 wire _0825_;
 wire _0826_;
 wire _0827_;
 wire _0828_;
 wire _0829_;
 wire _0830_;
 wire _0831_;
 wire _0832_;
 wire _0833_;
 wire _0834_;
 wire _0835_;
 wire _0836_;
 wire _0837_;
 wire _0838_;
 wire _0839_;
 wire _0840_;
 wire _0841_;
 wire _0842_;
 wire _0843_;
 wire _0844_;
 wire _0845_;
 wire _0846_;
 wire _0847_;
 wire _0848_;
 wire _0849_;
 wire _0850_;
 wire _0851_;
 wire _0852_;
 wire _0853_;
 wire _0854_;
 wire _0855_;
 wire _0856_;
 wire _0857_;
 wire _0858_;
 wire _0859_;
 wire _0860_;
 wire _0861_;
 wire _0862_;
 wire _0863_;
 wire _0864_;
 wire _0865_;
 wire _0866_;
 wire _0867_;
 wire _0868_;
 wire _0869_;
 wire _0870_;
 wire _0871_;
 wire _0872_;
 wire _0873_;
 wire _0874_;
 wire _0875_;
 wire _0876_;
 wire _0877_;
 wire _0878_;
 wire _0879_;
 wire _0880_;
 wire _0881_;
 wire _0882_;
 wire _0883_;
 wire _0884_;
 wire _0885_;
 wire _0886_;
 wire _0887_;
 wire _0888_;
 wire _0889_;
 wire _0890_;
 wire _0891_;
 wire _0892_;
 wire _0893_;
 wire _0894_;
 wire _0895_;
 wire _0896_;
 wire _0897_;
 wire _0898_;
 wire _0899_;
 wire _0900_;
 wire _0901_;
 wire _0902_;
 wire _0903_;
 wire _0904_;
 wire _0905_;
 wire _0906_;
 wire _0907_;
 wire _0908_;
 wire _0909_;
 wire _0910_;
 wire _0911_;
 wire _0912_;
 wire _0913_;
 wire _0914_;
 wire _0915_;
 wire _0916_;
 wire _0917_;
 wire _0918_;
 wire _0919_;
 wire _0920_;
 wire _0921_;
 wire _0922_;
 wire _0923_;
 wire _0924_;
 wire _0925_;
 wire _0926_;
 wire _0927_;
 wire _0928_;
 wire _0929_;
 wire _0930_;
 wire _0931_;
 wire _0932_;
 wire _0933_;
 wire _0934_;
 wire _0935_;
 wire _0936_;
 wire _0937_;
 wire _0938_;
 wire _0939_;
 wire _0940_;
 wire _0941_;
 wire _0942_;
 wire _0943_;
 wire _0944_;
 wire _0945_;
 wire _0946_;
 wire _0947_;
 wire _0948_;
 wire _0949_;
 wire _0950_;
 wire _0951_;
 wire _0952_;
 wire _0953_;
 wire _0954_;
 wire _0955_;
 wire _0956_;
 wire _0957_;
 wire _0958_;
 wire _0959_;
 wire _0960_;
 wire _0961_;
 wire _0962_;
 wire _0963_;
 wire _0964_;
 wire _0965_;
 wire _0966_;
 wire _0967_;
 wire _0968_;
 wire _0969_;
 wire _0970_;
 wire _0971_;
 wire _0972_;
 wire _0973_;
 wire _0974_;
 wire _0975_;
 wire _0976_;
 wire _0977_;
 wire _0978_;
 wire _0979_;
 wire _0980_;
 wire _0981_;
 wire _0982_;
 wire _0983_;
 wire _0984_;
 wire _0985_;
 wire _0986_;
 wire _0987_;
 wire _0988_;
 wire _0989_;
 wire _0990_;
 wire _0991_;
 wire _0992_;
 wire _0993_;
 wire _0994_;
 wire _0995_;
 wire _0996_;
 wire _0997_;
 wire _0998_;
 wire _0999_;
 wire _1000_;
 wire _1001_;
 wire _1002_;
 wire _1003_;
 wire _1004_;
 wire _1005_;
 wire _1006_;
 wire _1007_;
 wire _1008_;
 wire _1009_;
 wire _1010_;
 wire _1011_;
 wire _1012_;
 wire _1013_;
 wire _1014_;
 wire _1015_;
 wire _1016_;
 wire _1017_;
 wire _1018_;
 wire _1019_;
 wire _1020_;
 wire _1021_;
 wire _1022_;
 wire _1023_;
 wire _1024_;
 wire _1025_;
 wire _1026_;
 wire _1027_;
 wire _1028_;
 wire _1029_;
 wire _1030_;
 wire _1031_;
 wire _1032_;
 wire _1033_;
 wire _1034_;
 wire _1035_;
 wire _1036_;
 wire _1037_;
 wire _1038_;
 wire _1039_;
 wire _1040_;
 wire _1041_;
 wire _1042_;
 wire _1043_;
 wire _1044_;
 wire _1045_;
 wire _1046_;
 wire _1047_;
 wire _1048_;
 wire _1049_;
 wire _1050_;
 wire _1051_;
 wire _1052_;
 wire _1053_;
 wire _1054_;
 wire _1055_;
 wire _1056_;
 wire _1057_;
 wire _1058_;
 wire _1059_;
 wire _1060_;
 wire _1061_;
 wire _1062_;
 wire _1063_;
 wire _1064_;
 wire _1065_;
 wire _1066_;
 wire _1067_;
 wire _1068_;
 wire _1069_;
 wire _1070_;
 wire _1071_;
 wire _1072_;
 wire _1073_;
 wire _1074_;
 wire _1075_;
 wire _1076_;
 wire _1077_;
 wire _1078_;
 wire _1079_;
 wire _1080_;
 wire _1081_;
 wire _1082_;
 wire _1083_;
 wire _1084_;
 wire _1085_;
 wire _1086_;
 wire _1087_;
 wire _1088_;
 wire _1089_;
 wire _1090_;
 wire _1091_;
 wire _1092_;
 wire _1093_;
 wire _1094_;
 wire _1095_;
 wire _1096_;
 wire _1097_;
 wire _1098_;
 wire _1099_;
 wire _1100_;
 wire _1101_;
 wire _1102_;
 wire _1103_;
 wire _1104_;
 wire _1105_;
 wire _1106_;
 wire _1107_;
 wire _1108_;
 wire _1109_;
 wire _1110_;
 wire _1111_;
 wire _1112_;
 wire _1113_;
 wire _1114_;
 wire _1115_;
 wire _1116_;
 wire _1117_;
 wire _1118_;
 wire _1119_;
 wire _1120_;
 wire _1121_;
 wire _1122_;
 wire _1123_;
 wire _1124_;
 wire _1125_;
 wire _1126_;
 wire _1127_;
 wire _1128_;
 wire _1129_;
 wire _1130_;
 wire _1131_;
 wire _1132_;
 wire _1133_;
 wire _1134_;
 wire _1135_;
 wire _1136_;
 wire _1137_;
 wire _1138_;
 wire _1139_;
 wire _1140_;
 wire _1141_;
 wire _1142_;
 wire _1143_;
 wire _1144_;
 wire _1145_;
 wire _1146_;
 wire _1147_;
 wire _1148_;
 wire _1149_;
 wire _1150_;
 wire _1151_;
 wire _1152_;
 wire _1153_;
 wire _1154_;
 wire _1155_;
 wire _1156_;
 wire _1157_;
 wire _1158_;
 wire _1159_;
 wire _1160_;
 wire _1161_;
 wire _1162_;
 wire _1163_;
 wire _1164_;
 wire _1165_;
 wire _1166_;
 wire _1167_;
 wire _1168_;
 wire _1169_;
 wire _1170_;
 wire _1171_;
 wire _1172_;
 wire _1173_;
 wire _1174_;
 wire _1175_;
 wire _1176_;
 wire _1177_;
 wire _1178_;
 wire _1179_;
 wire _1180_;
 wire _1181_;
 wire _1182_;
 wire _1183_;
 wire _1184_;
 wire _1185_;
 wire _1186_;
 wire _1187_;
 wire _1188_;
 wire _1189_;
 wire _1190_;
 wire _1191_;
 wire _1192_;
 wire _1193_;
 wire _1194_;
 wire _1195_;
 wire _1196_;
 wire _1197_;
 wire _1198_;
 wire _1199_;
 wire _1200_;
 wire _1201_;
 wire _1202_;
 wire _1203_;
 wire _1204_;
 wire _1205_;
 wire _1206_;
 wire _1207_;
 wire _1208_;
 wire _1209_;
 wire _1210_;
 wire _1211_;
 wire _1212_;
 wire _1213_;
 wire _1214_;
 wire _1215_;
 wire _1216_;
 wire _1217_;
 wire _1218_;
 wire _1219_;
 wire _1220_;
 wire _1221_;
 wire _1222_;
 wire _1223_;
 wire _1224_;
 wire _1225_;
 wire _1226_;
 wire _1227_;
 wire _1228_;
 wire _1229_;
 wire _1230_;
 wire _1231_;
 wire _1232_;
 wire _1233_;
 wire _1234_;
 wire _1235_;
 wire _1236_;
 wire _1237_;
 wire _1238_;
 wire _1239_;
 wire _1240_;
 wire _1241_;
 wire _1242_;
 wire _1243_;
 wire _1244_;
 wire _1245_;
 wire _1246_;
 wire _1247_;
 wire _1248_;
 wire _1249_;
 wire _1250_;
 wire _1251_;
 wire _1252_;
 wire _1253_;
 wire _1254_;
 wire _1255_;
 wire _1256_;
 wire _1257_;
 wire _1258_;
 wire _1259_;
 wire _1260_;
 wire _1261_;
 wire _1262_;
 wire _1263_;
 wire _1264_;
 wire _1265_;
 wire _1266_;
 wire _1267_;
 wire _1268_;
 wire _1269_;
 wire _1270_;
 wire _1271_;
 wire _1272_;
 wire _1273_;
 wire _1274_;
 wire _1275_;
 wire _1276_;
 wire _1277_;
 wire _1278_;
 wire _1279_;
 wire _1280_;
 wire _1281_;
 wire _1282_;
 wire _1283_;
 wire _1284_;
 wire _1285_;
 wire _1286_;
 wire _1287_;
 wire _1288_;
 wire _1289_;
 wire _1290_;
 wire _1291_;
 wire _1292_;
 wire _1293_;
 wire _1294_;
 wire _1295_;
 wire _1296_;
 wire _1297_;
 wire _1298_;
 wire _1299_;
 wire _1300_;
 wire _1301_;
 wire _1302_;
 wire _1303_;
 wire _1304_;
 wire _1305_;
 wire _1306_;
 wire _1307_;
 wire _1308_;
 wire _1309_;
 wire _1310_;
 wire _1311_;
 wire _1312_;
 wire _1313_;
 wire _1314_;
 wire _1315_;
 wire _1316_;
 wire _1317_;
 wire _1318_;
 wire _1319_;
 wire _1320_;
 wire _1321_;
 wire _1322_;
 wire _1323_;
 wire _1324_;
 wire _1325_;
 wire _1326_;
 wire _1327_;
 wire _1328_;
 wire _1329_;
 wire _1330_;
 wire _1331_;
 wire _1332_;
 wire _1333_;
 wire _1334_;
 wire _1335_;
 wire _1336_;
 wire _1337_;
 wire _1338_;
 wire _1339_;
 wire _1340_;
 wire _1341_;
 wire _1342_;
 wire _1343_;
 wire _1344_;
 wire _1345_;
 wire _1346_;
 wire _1347_;
 wire _1348_;
 wire _1349_;
 wire _1350_;
 wire _1351_;
 wire _1352_;
 wire _1353_;
 wire _1354_;
 wire _1355_;
 wire _1356_;
 wire _1357_;
 wire _1358_;
 wire _1359_;
 wire _1360_;
 wire _1361_;
 wire _1362_;
 wire _1363_;
 wire _1364_;
 wire _1365_;
 wire _1366_;
 wire _1367_;
 wire _1368_;
 wire _1369_;
 wire _1370_;
 wire _1371_;
 wire _1372_;
 wire _1373_;
 wire _1374_;
 wire _1375_;
 wire _1376_;
 wire _1377_;
 wire _1378_;
 wire _1379_;
 wire _1380_;
 wire _1381_;
 wire _1382_;
 wire _1383_;
 wire _1384_;
 wire _1385_;
 wire _1386_;
 wire _1387_;
 wire _1388_;
 wire _1389_;
 wire _1390_;
 wire _1391_;
 wire _1392_;
 wire _1393_;
 wire _1394_;
 wire _1395_;
 wire _1396_;
 wire _1397_;
 wire _1398_;
 wire _1399_;
 wire _1400_;
 wire _1401_;
 wire _1402_;
 wire _1403_;
 wire _1404_;
 wire _1405_;
 wire _1406_;
 wire _1407_;
 wire _1408_;
 wire _1409_;
 wire _1410_;
 wire _1411_;
 wire _1412_;
 wire _1413_;
 wire _1414_;
 wire _1415_;
 wire _1416_;
 wire _1417_;
 wire _1418_;
 wire _1419_;
 wire _1420_;
 wire _1421_;
 wire _1422_;
 wire _1423_;
 wire _1424_;
 wire _1425_;
 wire _1426_;
 wire _1427_;
 wire _1428_;
 wire _1429_;
 wire _1430_;
 wire _1431_;
 wire _1432_;
 wire _1433_;
 wire _1434_;
 wire _1435_;
 wire _1436_;
 wire _1437_;
 wire _1438_;
 wire _1439_;
 wire _1440_;
 wire _1441_;
 wire _1442_;
 wire _1443_;
 wire _1444_;
 wire _1445_;
 wire _1446_;
 wire _1447_;
 wire _1448_;
 wire _1449_;
 wire _1450_;
 wire _1451_;
 wire _1452_;
 wire _1453_;
 wire _1454_;
 wire _1455_;
 wire _1456_;
 wire _1457_;
 wire _1458_;
 wire _1459_;
 wire _1460_;
 wire _1461_;
 wire _1462_;
 wire _1463_;
 wire _1464_;
 wire _1465_;
 wire _1466_;
 wire _1467_;
 wire _1468_;
 wire _1469_;
 wire _1470_;
 wire _1471_;
 wire _1472_;
 wire _1473_;
 wire _1474_;
 wire _1475_;
 wire _1476_;
 wire _1477_;
 wire _1478_;
 wire _1479_;
 wire _1480_;
 wire _1481_;
 wire _1482_;
 wire _1483_;
 wire _1484_;
 wire _1485_;
 wire _1486_;
 wire _1487_;
 wire _1488_;
 wire _1489_;
 wire _1490_;
 wire _1491_;
 wire _1492_;
 wire _1493_;
 wire _1494_;
 wire _1495_;
 wire _1496_;
 wire _1497_;
 wire _1498_;
 wire _1499_;
 wire _1500_;
 wire _1501_;
 wire _1502_;
 wire _1503_;
 wire _1504_;
 wire _1505_;
 wire _1506_;
 wire _1507_;
 wire _1508_;
 wire _1509_;
 wire _1510_;
 wire _1511_;
 wire _1512_;
 wire _1513_;
 wire _1514_;
 wire _1515_;
 wire _1516_;
 wire _1517_;
 wire _1518_;
 wire _1519_;
 wire _1520_;
 wire _1521_;
 wire _1522_;
 wire _1523_;
 wire _1524_;
 wire _1525_;
 wire _1526_;
 wire _1527_;
 wire _1528_;
 wire _1529_;
 wire _1530_;
 wire _1531_;
 wire _1532_;
 wire _1533_;
 wire _1534_;
 wire _1535_;
 wire _1536_;
 wire _1537_;
 wire _1538_;
 wire _1539_;
 wire _1540_;
 wire _1541_;
 wire _1542_;
 wire _1543_;
 wire _1544_;
 wire _1545_;
 wire _1546_;
 wire _1547_;
 wire _1548_;
 wire _1549_;
 wire _1550_;
 wire _1551_;
 wire _1552_;
 wire _1553_;
 wire _1554_;
 wire _1555_;
 wire _1556_;
 wire _1557_;
 wire _1558_;
 wire _1559_;
 wire _1560_;
 wire _1561_;
 wire _1562_;
 wire _1563_;
 wire _1564_;
 wire _1565_;
 wire _1566_;
 wire _1567_;
 wire _1568_;
 wire _1569_;
 wire _1570_;
 wire _1571_;
 wire _1572_;
 wire _1573_;
 wire _1574_;
 wire _1575_;
 wire _1576_;
 wire _1577_;
 wire _1578_;
 wire _1579_;
 wire _1580_;
 wire _1581_;
 wire _1582_;
 wire _1583_;
 wire _1584_;
 wire _1585_;
 wire _1586_;
 wire _1587_;
 wire _1588_;
 wire _1589_;
 wire _1590_;
 wire _1591_;
 wire _1592_;
 wire _1593_;
 wire _1594_;
 wire _1595_;
 wire _1596_;
 wire _1597_;
 wire _1598_;
 wire _1599_;
 wire _1600_;
 wire _1601_;
 wire _1602_;
 wire _1603_;
 wire _1604_;
 wire _1605_;
 wire _1606_;
 wire _1607_;
 wire _1608_;
 wire _1609_;
 wire _1610_;
 wire _1611_;
 wire _1612_;
 wire _1613_;
 wire _1614_;
 wire _1615_;
 wire _1616_;
 wire _1617_;
 wire _1618_;
 wire _1619_;
 wire _1620_;
 wire _1621_;
 wire _1622_;
 wire _1623_;
 wire _1624_;
 wire _1625_;
 wire _1626_;
 wire _1627_;
 wire _1628_;
 wire _1629_;
 wire _1630_;
 wire _1631_;
 wire _1632_;
 wire _1633_;
 wire _1634_;
 wire _1635_;
 wire _1636_;
 wire _1637_;
 wire _1638_;
 wire _1639_;
 wire _1640_;
 wire _1641_;
 wire _1642_;
 wire _1643_;
 wire _1644_;
 wire _1645_;
 wire _1646_;
 wire _1647_;
 wire _1648_;
 wire _1649_;
 wire _1650_;
 wire _1651_;
 wire _1652_;
 wire _1653_;
 wire _1654_;
 wire _1655_;
 wire _1656_;
 wire _1657_;
 wire _1658_;
 wire _1659_;
 wire _1660_;
 wire _1661_;
 wire _1662_;
 wire _1663_;
 wire _1664_;
 wire _1665_;
 wire _1666_;
 wire _1667_;
 wire _1668_;
 wire _1669_;
 wire _1670_;
 wire _1671_;
 wire _1672_;
 wire _1673_;
 wire _1674_;
 wire _1675_;
 wire _1676_;
 wire _1677_;
 wire _1678_;
 wire _1679_;
 wire _1680_;
 wire _1681_;
 wire _1682_;
 wire _1683_;
 wire _1684_;
 wire _1685_;
 wire _1686_;
 wire _1687_;
 wire _1688_;
 wire _1689_;
 wire _1690_;
 wire _1691_;
 wire _1692_;
 wire _1693_;
 wire _1694_;
 wire _1695_;
 wire _1696_;
 wire _1697_;
 wire _1698_;
 wire _1699_;
 wire _1700_;
 wire _1701_;
 wire _1702_;
 wire _1703_;
 wire _1704_;
 wire _1705_;
 wire _1706_;
 wire _1707_;
 wire _1708_;
 wire _1709_;
 wire _1710_;
 wire _1711_;
 wire _1712_;
 wire _1713_;
 wire _1714_;
 wire _1715_;
 wire _1716_;
 wire _1717_;
 wire _1718_;
 wire _1719_;
 wire _1720_;
 wire _1721_;
 wire _1722_;
 wire _1723_;
 wire _1724_;
 wire _1725_;
 wire _1726_;
 wire _1727_;
 wire _1728_;
 wire _1729_;
 wire _1730_;
 wire _1731_;
 wire _1732_;
 wire _1733_;
 wire _1734_;
 wire _1735_;
 wire _1736_;
 wire _1737_;
 wire _1738_;
 wire _1739_;
 wire _1740_;
 wire _1741_;
 wire _1742_;
 wire _1743_;
 wire _1744_;
 wire _1745_;
 wire _1746_;
 wire _1747_;
 wire _1748_;
 wire _1749_;
 wire _1750_;
 wire _1751_;
 wire _1752_;
 wire _1753_;
 wire _1754_;
 wire _1755_;
 wire _1756_;
 wire _1757_;
 wire _1758_;
 wire _1759_;
 wire _1760_;
 wire _1761_;
 wire _1762_;
 wire _1763_;
 wire _1764_;
 wire _1765_;
 wire _1766_;
 wire _1767_;
 wire _1768_;
 wire _1769_;
 wire _1770_;
 wire _1771_;
 wire _1772_;
 wire _1773_;
 wire _1774_;
 wire _1775_;
 wire _1776_;
 wire _1777_;
 wire _1778_;
 wire _1779_;
 wire _1780_;
 wire _1781_;
 wire _1782_;
 wire _1783_;
 wire _1784_;
 wire _1785_;
 wire _1786_;
 wire _1787_;
 wire _1788_;
 wire _1789_;
 wire _1790_;
 wire _1791_;
 wire _1792_;
 wire _1793_;
 wire _1794_;
 wire _1795_;
 wire _1796_;
 wire _1797_;
 wire _1798_;
 wire _1799_;
 wire _1800_;
 wire _1801_;
 wire _1802_;
 wire _1803_;
 wire _1804_;
 wire _1805_;
 wire _1806_;
 wire _1807_;
 wire _1808_;
 wire _1809_;
 wire _1810_;
 wire _1811_;
 wire _1812_;
 wire _1813_;
 wire _1814_;
 wire _1815_;
 wire _1816_;
 wire _1817_;
 wire _1818_;
 wire _1819_;
 wire _1820_;
 wire _1821_;
 wire _1822_;
 wire _1823_;
 wire _1824_;
 wire _1825_;
 wire _1826_;
 wire _1827_;
 wire _1828_;
 wire _1829_;
 wire _1830_;
 wire _1831_;
 wire _1832_;
 wire _1833_;
 wire _1834_;
 wire _1835_;
 wire _1836_;
 wire _1837_;
 wire _1838_;
 wire _1839_;
 wire _1840_;
 wire _1841_;
 wire _1842_;
 wire _1843_;
 wire _1844_;
 wire _1845_;
 wire _1846_;
 wire _1847_;
 wire _1848_;
 wire _1849_;
 wire _1850_;
 wire _1851_;
 wire _1852_;
 wire _1853_;
 wire _1854_;
 wire _1855_;
 wire _1856_;
 wire _1857_;
 wire _1858_;
 wire _1859_;
 wire _1860_;
 wire _1861_;
 wire _1862_;
 wire _1863_;
 wire _1864_;
 wire _1865_;
 wire _1866_;
 wire _1867_;
 wire _1868_;
 wire _1869_;
 wire _1870_;
 wire _1871_;
 wire _1872_;
 wire _1873_;
 wire _1874_;
 wire _1875_;
 wire _1876_;
 wire _1877_;
 wire _1878_;
 wire _1879_;
 wire _1880_;
 wire _1881_;
 wire _1882_;
 wire _1883_;
 wire _1884_;
 wire _1885_;
 wire _1886_;
 wire _1887_;
 wire _1888_;
 wire _1889_;
 wire _1890_;
 wire _1891_;
 wire _1892_;
 wire _1893_;
 wire _1894_;
 wire _1895_;
 wire _1896_;
 wire _1897_;
 wire _1898_;
 wire _1899_;
 wire _1900_;
 wire _1901_;
 wire _1902_;
 wire _1903_;
 wire _1904_;
 wire _1905_;
 wire _1906_;
 wire _1907_;
 wire _1908_;
 wire _1909_;
 wire _1910_;
 wire _1911_;
 wire _1912_;
 wire _1913_;
 wire _1914_;
 wire _1915_;
 wire _1916_;
 wire _1917_;
 wire _1918_;
 wire _1919_;
 wire _1920_;
 wire _1921_;
 wire _1922_;
 wire _1923_;
 wire _1924_;
 wire _1925_;
 wire _1926_;
 wire _1927_;
 wire _1928_;
 wire _1929_;
 wire _1930_;
 wire _1931_;
 wire _1932_;
 wire _1933_;
 wire _1934_;
 wire _1935_;
 wire _1936_;
 wire _1937_;
 wire _1938_;
 wire _1939_;
 wire _1940_;
 wire _1941_;
 wire _1942_;
 wire _1943_;
 wire _1944_;
 wire _1945_;
 wire _1946_;
 wire _1947_;
 wire _1948_;
 wire _1949_;
 wire _1950_;
 wire _1951_;
 wire _1952_;
 wire _1953_;
 wire _1954_;
 wire _1955_;
 wire _1956_;
 wire _1957_;
 wire _1958_;
 wire _1959_;
 wire _1960_;
 wire _1961_;
 wire _1962_;
 wire _1963_;
 wire _1964_;
 wire _1965_;
 wire _1966_;
 wire _1967_;
 wire _1968_;
 wire _1969_;
 wire _1970_;
 wire _1971_;
 wire _1972_;
 wire _1973_;
 wire _1974_;
 wire _1975_;
 wire _1976_;
 wire _1977_;
 wire _1978_;
 wire _1979_;
 wire _1980_;
 wire _1981_;
 wire _1982_;
 wire _1983_;
 wire _1984_;
 wire _1985_;
 wire _1986_;
 wire _1987_;
 wire _1988_;
 wire _1989_;
 wire _1990_;
 wire _1991_;
 wire _1992_;
 wire _1993_;
 wire _1994_;
 wire _1995_;
 wire _1996_;
 wire _1997_;
 wire _1998_;
 wire _1999_;
 wire _2000_;
 wire _2001_;
 wire _2002_;
 wire _2003_;
 wire _2004_;
 wire _2005_;
 wire _2006_;
 wire _2007_;
 wire _2008_;
 wire _2009_;
 wire _2010_;
 wire _2011_;
 wire _2012_;
 wire _2013_;
 wire _2014_;
 wire _2015_;
 wire _2016_;
 wire _2017_;
 wire _2018_;
 wire _2019_;
 wire _2020_;
 wire _2021_;
 wire _2022_;
 wire _2023_;
 wire _2024_;
 wire _2025_;
 wire _2026_;
 wire _2027_;
 wire _2028_;
 wire _2029_;
 wire _2030_;
 wire _2031_;
 wire _2032_;
 wire _2033_;
 wire _2034_;
 wire _2035_;
 wire _2036_;
 wire _2037_;
 wire _2038_;
 wire _2039_;
 wire _2040_;
 wire _2041_;
 wire _2042_;
 wire _2043_;
 wire _2044_;
 wire _2045_;
 wire _2046_;
 wire _2047_;
 wire _2048_;
 wire _2049_;
 wire _2050_;
 wire _2051_;
 wire _2052_;
 wire _2053_;
 wire _2054_;
 wire _2055_;
 wire _2056_;
 wire _2057_;
 wire _2058_;
 wire _2059_;
 wire _2060_;
 wire _2061_;
 wire _2062_;
 wire _2063_;
 wire _2064_;
 wire _2065_;
 wire _2066_;
 wire _2067_;
 wire _2068_;
 wire _2069_;
 wire _2070_;
 wire _2071_;
 wire _2072_;
 wire _2073_;
 wire _2074_;
 wire _2075_;
 wire _2076_;
 wire _2077_;
 wire _2078_;
 wire _2079_;
 wire _2080_;
 wire _2081_;
 wire _2082_;
 wire _2083_;
 wire _2084_;
 wire _2085_;
 wire _2086_;
 wire _2087_;
 wire _2088_;
 wire _2089_;
 wire _2090_;
 wire _2091_;
 wire _2092_;
 wire _2093_;
 wire _2094_;
 wire _2095_;
 wire _2096_;
 wire _2097_;
 wire _2098_;
 wire _2099_;
 wire _2100_;
 wire _2101_;
 wire _2102_;
 wire _2103_;
 wire _2104_;
 wire _2105_;
 wire _2106_;
 wire _2107_;
 wire _2108_;
 wire _2109_;
 wire _2110_;
 wire _2111_;
 wire _2112_;
 wire _2113_;
 wire _2114_;
 wire _2115_;
 wire _2116_;
 wire _2117_;
 wire _2118_;
 wire _2119_;
 wire _2120_;
 wire _2121_;
 wire _2122_;
 wire _2123_;
 wire _2124_;
 wire _2125_;
 wire _2126_;
 wire _2127_;
 wire _2128_;
 wire _2129_;
 wire _2130_;
 wire _2131_;
 wire _2132_;
 wire _2133_;
 wire _2134_;
 wire _2135_;
 wire _2136_;
 wire _2137_;
 wire _2138_;
 wire _2139_;
 wire _2140_;
 wire _2141_;
 wire _2142_;
 wire _2143_;
 wire _2144_;
 wire _2145_;
 wire _2146_;
 wire _2147_;
 wire _2148_;
 wire _2149_;
 wire _2150_;
 wire _2151_;
 wire _2152_;
 wire _2153_;
 wire _2154_;
 wire _2155_;
 wire _2156_;
 wire _2157_;
 wire _2158_;
 wire _2159_;
 wire _2160_;
 wire _2161_;
 wire _2162_;
 wire _2163_;
 wire _2164_;
 wire _2165_;
 wire _2166_;
 wire _2167_;
 wire _2168_;
 wire _2169_;
 wire _2170_;
 wire _2171_;
 wire _2172_;
 wire _2173_;
 wire _2174_;
 wire _2175_;
 wire _2176_;
 wire _2177_;
 wire _2178_;
 wire _2179_;
 wire _2180_;
 wire _2181_;
 wire _2182_;
 wire _2183_;
 wire _2184_;
 wire _2185_;
 wire _2186_;
 wire _2187_;
 wire _2188_;
 wire _2189_;
 wire _2190_;
 wire _2191_;
 wire _2192_;
 wire _2193_;
 wire _2194_;
 wire _2195_;
 wire _2196_;
 wire _2197_;
 wire _2198_;
 wire _2199_;
 wire _2200_;
 wire _2201_;
 wire _2202_;
 wire _2203_;
 wire _2204_;
 wire _2205_;
 wire _2206_;
 wire _2207_;
 wire _2208_;
 wire _2209_;
 wire _2210_;
 wire _2211_;
 wire _2212_;
 wire _2213_;
 wire _2214_;
 wire _2215_;
 wire _2216_;
 wire _2217_;
 wire _2218_;
 wire _2219_;
 wire _2220_;
 wire _2221_;
 wire _2222_;
 wire _2223_;
 wire _2224_;
 wire _2225_;
 wire _2226_;
 wire _2227_;
 wire _2228_;
 wire _2229_;
 wire _2230_;
 wire _2231_;
 wire _2232_;
 wire _2233_;
 wire _2234_;
 wire _2235_;
 wire _2236_;
 wire _2237_;
 wire _2238_;
 wire _2239_;
 wire _2240_;
 wire _2241_;
 wire _2242_;
 wire _2243_;
 wire _2244_;
 wire _2245_;
 wire _2246_;
 wire _2247_;
 wire _2248_;
 wire _2249_;
 wire _2250_;
 wire _2251_;
 wire _2252_;
 wire _2253_;
 wire _2254_;
 wire _2255_;
 wire _2256_;
 wire _2257_;
 wire _2258_;
 wire _2259_;
 wire _2260_;
 wire _2261_;
 wire _2262_;
 wire _2263_;
 wire _2264_;
 wire _2265_;
 wire _2266_;
 wire _2267_;
 wire _2268_;
 wire _2269_;
 wire _2270_;
 wire _2271_;
 wire _2272_;
 wire _2273_;
 wire _2274_;
 wire _2275_;
 wire _2276_;
 wire _2277_;
 wire _2278_;
 wire _2279_;
 wire _2280_;
 wire _2281_;
 wire _2282_;
 wire _2283_;
 wire _2284_;
 wire _2285_;
 wire _2286_;
 wire _2287_;
 wire _2288_;
 wire _2289_;
 wire _2290_;
 wire _2291_;
 wire _2292_;
 wire _2293_;
 wire _2294_;
 wire _2295_;
 wire _2296_;
 wire _2297_;
 wire _2298_;
 wire _2299_;
 wire _2300_;
 wire _2301_;
 wire _2302_;
 wire _2303_;
 wire _2304_;
 wire _2305_;
 wire _2306_;
 wire _2307_;
 wire _2308_;
 wire _2309_;
 wire _2310_;
 wire _2311_;
 wire _2312_;
 wire _2313_;
 wire _2314_;
 wire _2315_;
 wire _2316_;
 wire _2317_;
 wire _2318_;
 wire _2319_;
 wire _2320_;
 wire _2321_;
 wire _2322_;
 wire _2323_;
 wire _2324_;
 wire _2325_;
 wire _2326_;
 wire _2327_;
 wire _2328_;
 wire _2329_;
 wire _2330_;
 wire _2331_;
 wire _2332_;
 wire _2333_;
 wire _2334_;
 wire _2335_;
 wire _2336_;
 wire _2337_;
 wire _2338_;
 wire _2339_;
 wire _2340_;
 wire _2341_;
 wire _2342_;
 wire _2343_;
 wire _2344_;
 wire _2345_;
 wire _2346_;
 wire _2347_;
 wire _2348_;
 wire _2349_;
 wire _2350_;
 wire _2351_;
 wire _2352_;
 wire _2353_;
 wire _2354_;
 wire _2355_;
 wire _2356_;
 wire _2357_;
 wire _2358_;
 wire _2359_;
 wire _2360_;
 wire _2361_;
 wire _2362_;
 wire _2363_;
 wire _2364_;
 wire _2365_;
 wire _2366_;
 wire _2367_;
 wire _2368_;
 wire _2369_;
 wire _2370_;
 wire _2371_;
 wire _2372_;
 wire _2373_;
 wire _2374_;
 wire _2375_;
 wire _2376_;
 wire _2377_;
 wire _2378_;
 wire _2379_;
 wire _2380_;
 wire _2381_;
 wire _2382_;
 wire _2383_;
 wire _2384_;
 wire _2385_;
 wire _2386_;
 wire _2387_;
 wire _2388_;
 wire _2389_;
 wire _2390_;
 wire _2391_;
 wire _2392_;
 wire _2393_;
 wire _2394_;
 wire _2395_;
 wire _2396_;
 wire _2397_;
 wire _2398_;
 wire _2399_;
 wire _2400_;
 wire _2401_;
 wire _2402_;
 wire _2403_;
 wire _2404_;
 wire _2405_;
 wire _2406_;
 wire _2407_;
 wire _2408_;
 wire _2409_;
 wire _2410_;
 wire _2411_;
 wire _2412_;
 wire _2413_;
 wire _2414_;
 wire _2415_;
 wire _2416_;
 wire _2417_;
 wire _2418_;
 wire _2419_;
 wire _2420_;
 wire _2421_;
 wire _2422_;
 wire _2423_;
 wire _2424_;
 wire _2425_;
 wire _2426_;
 wire _2427_;
 wire _2428_;
 wire _2429_;
 wire _2430_;
 wire _2431_;
 wire _2432_;
 wire _2433_;
 wire _2434_;
 wire _2435_;
 wire _2436_;
 wire _2437_;
 wire _2438_;
 wire _2439_;
 wire _2440_;
 wire _2441_;
 wire _2442_;
 wire _2443_;
 wire _2444_;
 wire _2445_;
 wire _2446_;
 wire _2447_;
 wire _2448_;
 wire _2449_;
 wire _2450_;
 wire _2451_;
 wire _2452_;
 wire _2453_;
 wire _2454_;
 wire _2455_;
 wire _2456_;
 wire _2457_;
 wire _2458_;
 wire _2459_;
 wire _2460_;
 wire _2461_;
 wire _2462_;
 wire _2463_;
 wire _2464_;
 wire _2465_;
 wire _2466_;
 wire _2467_;
 wire _2468_;
 wire _2469_;
 wire _2470_;
 wire _2471_;
 wire _2472_;
 wire _2473_;
 wire _2474_;
 wire _2475_;
 wire _2476_;
 wire _2477_;
 wire _2478_;
 wire _2479_;
 wire _2480_;
 wire _2481_;
 wire _2482_;
 wire _2483_;
 wire _2484_;
 wire _2485_;
 wire _2486_;
 wire _2487_;
 wire _2488_;
 wire _2489_;
 wire _2490_;
 wire _2491_;
 wire _2492_;
 wire _2493_;
 wire _2494_;
 wire _2495_;
 wire _2496_;
 wire _2497_;
 wire _2498_;
 wire _2499_;
 wire _2500_;
 wire _2501_;
 wire _2502_;
 wire _2503_;
 wire _2504_;
 wire _2505_;
 wire _2506_;
 wire _2507_;
 wire _2508_;
 wire _2509_;
 wire _2510_;
 wire _2511_;
 wire _2512_;
 wire _2513_;
 wire _2514_;
 wire _2515_;
 wire _2516_;
 wire _2517_;
 wire _2518_;
 wire _2519_;
 wire _2520_;
 wire _2521_;
 wire _2522_;
 wire _2523_;
 wire _2524_;
 wire _2525_;
 wire _2526_;
 wire _2527_;
 wire _2528_;
 wire _2529_;
 wire _2530_;
 wire _2531_;
 wire _2532_;
 wire _2533_;
 wire _2534_;
 wire _2535_;
 wire _2536_;
 wire _2537_;
 wire _2538_;
 wire _2539_;
 wire _2540_;
 wire _2541_;
 wire _2542_;
 wire _2543_;
 wire _2544_;
 wire _2545_;
 wire _2546_;
 wire _2547_;
 wire _2548_;
 wire _2549_;
 wire _2550_;
 wire _2551_;
 wire _2552_;
 wire _2553_;
 wire _2554_;
 wire _2555_;
 wire _2556_;
 wire _2557_;
 wire _2558_;
 wire _2559_;
 wire _2560_;
 wire _2561_;
 wire _2562_;
 wire _2563_;
 wire _2564_;
 wire _2565_;
 wire _2566_;
 wire _2567_;
 wire _2568_;
 wire _2569_;
 wire _2570_;
 wire _2571_;
 wire _2572_;
 wire _2573_;
 wire _2574_;
 wire _2575_;
 wire _2576_;
 wire _2577_;
 wire _2578_;
 wire _2579_;
 wire _2580_;
 wire _2581_;
 wire _2582_;
 wire _2583_;
 wire _2584_;
 wire _2585_;
 wire _2586_;
 wire _2587_;
 wire _2588_;
 wire _2589_;
 wire _2590_;
 wire _2591_;
 wire _2592_;
 wire _2593_;
 wire _2594_;
 wire _2595_;
 wire _2596_;
 wire _2597_;
 wire _2598_;
 wire _2599_;
 wire _2600_;
 wire _2601_;
 wire _2602_;
 wire _2603_;
 wire _2604_;
 wire _2605_;
 wire _2606_;
 wire _2607_;
 wire _2608_;
 wire _2609_;
 wire _2610_;
 wire _2611_;
 wire _2612_;
 wire _2613_;
 wire _2614_;
 wire _2615_;
 wire _2616_;
 wire _2617_;
 wire _2618_;
 wire _2619_;
 wire _2620_;
 wire _2621_;
 wire _2622_;
 wire _2623_;
 wire _2624_;
 wire _2625_;
 wire _2626_;
 wire _2627_;
 wire _2628_;
 wire _2629_;
 wire _2630_;
 wire _2631_;
 wire _2632_;
 wire _2633_;
 wire _2634_;
 wire _2635_;
 wire _2636_;
 wire _2637_;
 wire _2638_;
 wire _2639_;
 wire _2640_;
 wire _2641_;
 wire _2642_;
 wire _2643_;
 wire _2644_;
 wire _2645_;
 wire _2646_;
 wire _2647_;
 wire _2648_;
 wire _2649_;
 wire _2650_;
 wire _2651_;
 wire _2652_;
 wire _2653_;
 wire _2654_;
 wire _2655_;
 wire _2656_;
 wire _2657_;
 wire _2658_;
 wire _2659_;
 wire _2660_;
 wire _2661_;
 wire _2662_;
 wire _2663_;
 wire _2664_;
 wire _2665_;
 wire _2666_;
 wire _2667_;
 wire _2668_;
 wire _2669_;
 wire _2670_;
 wire _2671_;
 wire _2672_;
 wire _2673_;
 wire _2674_;
 wire _2675_;
 wire _2676_;
 wire _2677_;
 wire _2678_;
 wire _2679_;
 wire _2680_;
 wire _2681_;
 wire _2682_;
 wire _2683_;
 wire _2684_;
 wire _2685_;
 wire _2686_;
 wire _2687_;
 wire _2688_;
 wire _2689_;
 wire _2690_;
 wire _2691_;
 wire _2692_;
 wire _2693_;
 wire _2694_;
 wire _2695_;
 wire _2696_;
 wire _2697_;
 wire _2698_;
 wire _2699_;
 wire _2700_;
 wire _2701_;
 wire _2702_;
 wire _2703_;
 wire _2704_;
 wire _2705_;
 wire _2706_;
 wire _2707_;
 wire _2708_;
 wire _2709_;
 wire _2710_;
 wire _2711_;
 wire _2712_;
 wire _2713_;
 wire _2714_;
 wire _2715_;
 wire _2716_;
 wire _2717_;
 wire _2718_;
 wire _2719_;
 wire _2720_;
 wire _2721_;
 wire _2722_;
 wire _2723_;
 wire _2724_;
 wire _2725_;
 wire _2726_;
 wire _2727_;
 wire _2728_;
 wire _2729_;
 wire _2730_;
 wire _2731_;
 wire _2732_;
 wire _2733_;
 wire _2734_;
 wire _2735_;
 wire _2736_;
 wire _2737_;
 wire _2738_;
 wire _2739_;
 wire _2740_;
 wire _2741_;
 wire _2742_;
 wire _2743_;
 wire _2744_;
 wire _2745_;
 wire _2746_;
 wire _2747_;
 wire _2748_;
 wire _2749_;
 wire _2750_;
 wire _2751_;
 wire _2752_;
 wire _2753_;
 wire _2754_;
 wire _2755_;
 wire _2756_;
 wire _2757_;
 wire _2758_;
 wire _2759_;
 wire _2760_;
 wire _2761_;
 wire _2762_;
 wire _2763_;
 wire _2764_;
 wire _2765_;
 wire _2766_;
 wire _2767_;
 wire _2768_;
 wire _2769_;
 wire _2770_;
 wire _2771_;
 wire _2772_;
 wire _2773_;
 wire _2774_;
 wire _2775_;
 wire _2776_;
 wire _2777_;
 wire _2778_;
 wire _2779_;
 wire _2780_;
 wire _2781_;
 wire _2782_;
 wire _2783_;
 wire _2784_;
 wire _2785_;
 wire _2786_;
 wire _2787_;
 wire _2788_;
 wire _2789_;
 wire _2790_;
 wire _2791_;
 wire _2792_;
 wire _2793_;
 wire _2794_;
 wire _2795_;
 wire _2796_;
 wire _2797_;
 wire _2798_;
 wire _2799_;
 wire _2800_;
 wire _2801_;
 wire _2802_;
 wire _2803_;
 wire _2804_;
 wire _2805_;
 wire _2806_;
 wire _2807_;
 wire _2808_;
 wire _2809_;
 wire _2810_;
 wire _2811_;
 wire _2812_;
 wire _2813_;
 wire _2814_;
 wire _2815_;
 wire _2816_;
 wire _2817_;
 wire _2818_;
 wire _2819_;
 wire _2820_;
 wire _2821_;
 wire _2822_;
 wire _2823_;
 wire _2824_;
 wire _2825_;
 wire _2826_;
 wire _2827_;
 wire _2828_;
 wire _2829_;
 wire _2830_;
 wire _2831_;
 wire _2832_;
 wire _2833_;
 wire _2834_;
 wire _2835_;
 wire _2836_;
 wire _2837_;
 wire _2838_;
 wire _2839_;
 wire _2840_;
 wire _2841_;
 wire _2842_;
 wire _2843_;
 wire _2844_;
 wire _2845_;
 wire _2846_;
 wire _2847_;
 wire _2848_;
 wire _2849_;
 wire _2850_;
 wire _2851_;
 wire _2852_;
 wire _2853_;
 wire _2854_;
 wire _2855_;
 wire _2856_;
 wire _2857_;
 wire _2858_;
 wire _2859_;
 wire _2860_;
 wire _2861_;
 wire _2862_;
 wire _2863_;
 wire _2864_;
 wire _2865_;
 wire _2866_;
 wire _2867_;
 wire _2868_;
 wire _2869_;
 wire _2870_;
 wire _2871_;
 wire _2872_;
 wire _2873_;
 wire _2874_;
 wire _2875_;
 wire _2876_;
 wire _2877_;
 wire _2878_;
 wire _2879_;
 wire _2880_;
 wire _2881_;
 wire _2882_;
 wire _2883_;
 wire _2884_;
 wire _2885_;
 wire _2886_;
 wire _2887_;
 wire _2888_;
 wire _2889_;
 wire _2890_;
 wire _2891_;
 wire _2892_;
 wire _2893_;
 wire _2894_;
 wire _2895_;
 wire _2896_;
 wire _2897_;
 wire _2898_;
 wire _2899_;
 wire _2900_;
 wire _2901_;
 wire _2902_;
 wire _2903_;
 wire _2904_;
 wire _2905_;
 wire _2906_;
 wire _2907_;
 wire _2908_;
 wire _2909_;
 wire _2910_;
 wire _2911_;
 wire _2912_;
 wire _2913_;
 wire _2914_;
 wire _2915_;
 wire _2916_;
 wire _2917_;
 wire _2918_;
 wire _2919_;
 wire _2920_;
 wire _2921_;
 wire _2922_;
 wire _2923_;
 wire _2924_;
 wire _2925_;
 wire _2926_;
 wire _2927_;
 wire _2928_;
 wire _2929_;
 wire _2930_;
 wire _2931_;
 wire _2932_;
 wire _2933_;
 wire _2934_;
 wire _2935_;
 wire _2936_;
 wire _2937_;
 wire _2938_;
 wire _2939_;
 wire _2940_;
 wire _2941_;
 wire _2942_;
 wire _2943_;
 wire _2944_;
 wire _2945_;
 wire _2946_;
 wire _2947_;
 wire _2948_;
 wire _2949_;
 wire _2950_;
 wire _2951_;
 wire _2952_;
 wire _2953_;
 wire _2954_;
 wire _2955_;
 wire _2956_;
 wire _2957_;
 wire _2958_;
 wire _2959_;
 wire _2960_;
 wire _2961_;
 wire _2962_;
 wire _2963_;
 wire _2964_;
 wire _2965_;
 wire _2966_;
 wire _2967_;
 wire _2968_;
 wire _2969_;
 wire _2970_;
 wire _2971_;
 wire _2972_;
 wire _2973_;
 wire _2974_;
 wire _2975_;
 wire _2976_;
 wire _2977_;
 wire _2978_;
 wire _2979_;
 wire _2980_;
 wire _2981_;
 wire _2982_;
 wire _2983_;
 wire _2984_;
 wire _2985_;
 wire _2986_;
 wire _2987_;
 wire _2988_;
 wire _2989_;
 wire _2990_;
 wire _2991_;
 wire _2992_;
 wire _2993_;
 wire _2994_;
 wire _2995_;
 wire _2996_;
 wire _2997_;
 wire _2998_;
 wire _2999_;
 wire _3000_;
 wire _3001_;
 wire _3002_;
 wire _3003_;
 wire _3004_;
 wire _3005_;
 wire _3006_;
 wire _3007_;
 wire _3008_;
 wire _3009_;
 wire _3010_;
 wire _3011_;
 wire _3012_;
 wire _3013_;
 wire _3014_;
 wire _3015_;
 wire _3016_;
 wire _3017_;
 wire _3018_;
 wire _3019_;
 wire _3020_;
 wire _3021_;
 wire _3022_;
 wire _3023_;
 wire _3024_;
 wire _3025_;
 wire _3026_;
 wire _3027_;
 wire _3028_;
 wire _3029_;
 wire _3030_;
 wire _3031_;
 wire _3032_;
 wire _3033_;
 wire _3034_;
 wire _3035_;
 wire _3036_;
 wire _3037_;
 wire _3038_;
 wire _3039_;
 wire _3040_;
 wire _3041_;
 wire _3042_;
 wire _3043_;
 wire _3044_;
 wire _3045_;
 wire _3046_;
 wire _3047_;
 wire _3048_;
 wire _3049_;
 wire _3050_;
 wire _3051_;
 wire _3052_;
 wire _3053_;
 wire _3054_;
 wire _3055_;
 wire _3056_;
 wire _3057_;
 wire _3058_;
 wire _3059_;
 wire _3060_;
 wire _3061_;
 wire _3062_;
 wire _3063_;
 wire _3064_;
 wire _3065_;
 wire _3066_;
 wire _3067_;
 wire _3068_;
 wire _3069_;
 wire _3070_;
 wire _3071_;
 wire _3072_;
 wire _3073_;
 wire _3074_;
 wire _3075_;
 wire _3076_;
 wire _3077_;
 wire _3078_;
 wire _3079_;
 wire _3080_;
 wire _3081_;
 wire _3082_;
 wire _3083_;
 wire _3084_;
 wire _3085_;
 wire _3086_;
 wire _3087_;
 wire _3088_;
 wire _3089_;
 wire _3090_;
 wire _3091_;
 wire _3092_;
 wire _3093_;
 wire _3094_;
 wire _3095_;
 wire _3096_;
 wire _3097_;
 wire _3098_;
 wire _3099_;
 wire _3100_;
 wire _3101_;
 wire _3102_;
 wire _3103_;
 wire _3104_;
 wire _3105_;
 wire _3106_;
 wire _3107_;
 wire _3108_;
 wire _3109_;
 wire _3110_;
 wire _3111_;
 wire _3112_;
 wire _3113_;
 wire _3114_;
 wire _3115_;
 wire _3116_;
 wire _3117_;
 wire _3118_;
 wire _3119_;
 wire _3120_;
 wire _3121_;
 wire _3122_;
 wire _3123_;
 wire _3124_;
 wire _3125_;
 wire _3126_;
 wire _3127_;
 wire _3128_;
 wire _3129_;
 wire _3130_;
 wire _3131_;
 wire _3132_;
 wire _3133_;
 wire _3134_;
 wire _3135_;
 wire _3136_;
 wire _3137_;
 wire _3138_;
 wire _3139_;
 wire _3140_;
 wire _3141_;
 wire _3142_;
 wire _3143_;
 wire _3144_;
 wire _3145_;
 wire _3146_;
 wire _3147_;
 wire _3148_;
 wire _3149_;
 wire _3150_;
 wire _3151_;
 wire _3152_;
 wire _3153_;
 wire _3154_;
 wire _3155_;
 wire _3156_;
 wire _3157_;
 wire _3158_;
 wire _3159_;
 wire _3160_;
 wire _3161_;
 wire _3162_;
 wire _3163_;
 wire _3164_;
 wire _3165_;
 wire _3166_;
 wire _3167_;
 wire _3168_;
 wire _3169_;
 wire _3170_;
 wire _3171_;
 wire _3172_;
 wire _3173_;
 wire _3174_;
 wire _3175_;
 wire _3176_;
 wire _3177_;
 wire _3178_;
 wire _3179_;
 wire _3180_;
 wire _3181_;
 wire _3182_;
 wire _3183_;
 wire _3184_;
 wire _3185_;
 wire _3186_;
 wire _3187_;
 wire _3188_;
 wire _3189_;
 wire _3190_;
 wire _3191_;
 wire _3192_;
 wire _3193_;
 wire _3194_;
 wire clknet_0_clk;
 wire net197;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net180;
 wire net181;
 wire net182;
 wire net183;
 wire net184;
 wire net185;
 wire net186;
 wire net187;
 wire net188;
 wire net189;
 wire net190;
 wire net191;
 wire net192;
 wire net193;
 wire net194;
 wire net195;
 wire net196;
 wire net198;
 wire net199;
 wire net200;
 wire net201;
 wire net202;
 wire net203;
 wire net204;
 wire net205;
 wire net206;
 wire net207;
 wire net208;
 wire net209;
 wire net210;
 wire net211;
 wire net212;
 wire net213;
 wire net214;
 wire net215;
 wire net216;
 wire net217;
 wire net218;
 wire net219;
 wire net220;
 wire net221;
 wire net222;
 wire net223;
 wire net224;
 wire net225;
 wire net226;
 wire net227;
 wire net228;
 wire net229;
 wire net230;
 wire net231;
 wire net232;
 wire net233;
 wire net234;
 wire net235;
 wire net236;
 wire net237;
 wire net238;
 wire net239;
 wire net240;
 wire net241;
 wire net242;
 wire net243;
 wire net244;
 wire net245;
 wire net246;
 wire net247;
 wire net248;
 wire net249;
 wire net250;
 wire net251;
 wire net252;
 wire net253;
 wire net254;
 wire net255;
 wire net256;
 wire net257;
 wire net258;
 wire net259;
 wire net260;
 wire net261;
 wire net262;
 wire net263;
 wire net264;
 wire net265;
 wire net266;
 wire net267;
 wire net268;
 wire net269;
 wire net270;
 wire net271;
 wire net272;
 wire net273;
 wire net274;
 wire net275;
 wire net276;
 wire net277;
 wire net278;
 wire net279;
 wire net280;
 wire net281;
 wire net282;
 wire net283;
 wire net284;
 wire net285;
 wire net286;
 wire net287;
 wire net288;
 wire net289;
 wire net290;
 wire net291;
 wire net292;
 wire net293;
 wire net294;
 wire net295;
 wire net296;
 wire net297;
 wire net298;
 wire net299;
 wire net300;
 wire net301;
 wire net302;
 wire net303;
 wire net304;
 wire net305;
 wire net306;
 wire net307;
 wire net308;
 wire net309;
 wire net310;
 wire net311;
 wire net312;
 wire net313;
 wire net314;
 wire net315;
 wire net316;
 wire net317;
 wire net318;
 wire net319;
 wire net320;
 wire net321;
 wire net322;
 wire net323;
 wire net324;
 wire net325;
 wire net326;
 wire net327;
 wire net328;
 wire net329;
 wire net330;
 wire net331;
 wire net332;
 wire net333;
 wire net334;
 wire net335;
 wire net336;
 wire net337;
 wire net338;
 wire net339;
 wire net340;
 wire net341;
 wire net342;
 wire net343;
 wire net344;
 wire net345;
 wire net346;
 wire net347;
 wire net348;
 wire net349;
 wire net350;
 wire net351;
 wire net352;
 wire net353;
 wire net354;
 wire net355;
 wire net356;
 wire net357;
 wire net358;
 wire net359;
 wire net360;
 wire net361;
 wire net362;
 wire net363;
 wire net364;
 wire net365;
 wire net366;
 wire net367;
 wire net368;
 wire net369;
 wire net370;
 wire net371;
 wire net372;
 wire net373;
 wire net374;
 wire net375;
 wire net376;
 wire net377;
 wire net378;
 wire net379;
 wire net380;
 wire net381;
 wire net382;
 wire net383;
 wire net384;
 wire net385;
 wire net386;
 wire net387;
 wire net388;
 wire net389;
 wire net390;
 wire net391;
 wire net392;
 wire net393;
 wire net394;
 wire net395;
 wire net396;
 wire net397;
 wire net398;
 wire net399;
 wire net400;
 wire net401;
 wire net402;
 wire net403;
 wire net404;
 wire net405;
 wire net406;
 wire net407;
 wire net408;
 wire net409;
 wire net410;
 wire net411;
 wire net412;
 wire net413;
 wire clknet_4_0_0_clk;
 wire clknet_4_1_0_clk;
 wire clknet_4_2_0_clk;
 wire clknet_4_3_0_clk;
 wire clknet_4_4_0_clk;
 wire clknet_4_5_0_clk;
 wire clknet_4_6_0_clk;
 wire clknet_4_7_0_clk;
 wire clknet_4_8_0_clk;
 wire clknet_4_9_0_clk;
 wire clknet_4_10_0_clk;
 wire clknet_4_11_0_clk;
 wire clknet_4_12_0_clk;
 wire clknet_4_13_0_clk;
 wire clknet_4_14_0_clk;
 wire clknet_4_15_0_clk;
 wire clknet_5_0__leaf_clk;
 wire clknet_5_1__leaf_clk;
 wire clknet_5_2__leaf_clk;
 wire clknet_5_3__leaf_clk;
 wire clknet_5_4__leaf_clk;
 wire clknet_5_5__leaf_clk;
 wire clknet_5_6__leaf_clk;
 wire clknet_5_7__leaf_clk;
 wire clknet_5_8__leaf_clk;
 wire clknet_5_9__leaf_clk;
 wire clknet_5_10__leaf_clk;
 wire clknet_5_11__leaf_clk;
 wire clknet_5_12__leaf_clk;
 wire clknet_5_13__leaf_clk;
 wire clknet_5_14__leaf_clk;
 wire clknet_5_15__leaf_clk;
 wire clknet_5_16__leaf_clk;
 wire clknet_5_17__leaf_clk;
 wire clknet_5_18__leaf_clk;
 wire clknet_5_19__leaf_clk;
 wire clknet_5_20__leaf_clk;
 wire clknet_5_21__leaf_clk;
 wire clknet_5_22__leaf_clk;
 wire clknet_5_23__leaf_clk;
 wire clknet_5_24__leaf_clk;
 wire clknet_5_25__leaf_clk;
 wire clknet_5_26__leaf_clk;
 wire clknet_5_27__leaf_clk;
 wire clknet_5_28__leaf_clk;
 wire clknet_5_29__leaf_clk;
 wire clknet_5_30__leaf_clk;
 wire clknet_5_31__leaf_clk;

 sg13g2_dfrbp_1 \Pong.control_unit.NES_Controller_Left.state_NESController[0]$_DFF_P_  (.CLK(clknet_5_0__leaf_clk),
    .RESET_B(net197),
    .D(_0000_),
    .Q_N(_0119_),
    .Q(\Pong.control_unit.NES_Controller_Left.state_NESController[0] ));
 sg13g2_dfrbp_1 \Pong.control_unit.NES_Controller_Left.state_NESController[10]$_DFF_P_  (.CLK(clknet_5_5__leaf_clk),
    .RESET_B(net198),
    .D(_0001_),
    .Q_N(_3166_),
    .Q(\Pong.control_unit.NES_Controller_Left.state_NESController[10] ));
 sg13g2_dfrbp_1 \Pong.control_unit.NES_Controller_Left.state_NESController[11]$_DFF_P_  (.CLK(clknet_5_4__leaf_clk),
    .RESET_B(net199),
    .D(_0002_),
    .Q_N(_3167_),
    .Q(\Pong.control_unit.NES_Controller_Left.state_NESController[11] ));
 sg13g2_dfrbp_1 \Pong.control_unit.NES_Controller_Left.state_NESController[12]$_DFF_P_  (.CLK(clknet_5_7__leaf_clk),
    .RESET_B(net200),
    .D(_0003_),
    .Q_N(_0125_),
    .Q(\Pong.control_unit.NES_Controller_Left.state_NESController[12] ));
 sg13g2_dfrbp_1 \Pong.control_unit.NES_Controller_Left.state_NESController[13]$_DFF_P_  (.CLK(clknet_5_18__leaf_clk),
    .RESET_B(net201),
    .D(_0004_),
    .Q_N(_3168_),
    .Q(\Pong.control_unit.NES_Controller_Left.state_NESController[13] ));
 sg13g2_dfrbp_1 \Pong.control_unit.NES_Controller_Left.state_NESController[14]$_DFF_P_  (.CLK(clknet_5_6__leaf_clk),
    .RESET_B(net202),
    .D(_0005_),
    .Q_N(_0124_),
    .Q(\Pong.control_unit.NES_Controller_Left.state_NESController[14] ));
 sg13g2_dfrbp_1 \Pong.control_unit.NES_Controller_Left.state_NESController[15]$_DFF_P_  (.CLK(clknet_5_18__leaf_clk),
    .RESET_B(net203),
    .D(_0006_),
    .Q_N(_3169_),
    .Q(\Pong.control_unit.NES_Controller_Left.state_NESController[15] ));
 sg13g2_dfrbp_1 \Pong.control_unit.NES_Controller_Left.state_NESController[16]$_DFF_P_  (.CLK(clknet_5_5__leaf_clk),
    .RESET_B(net204),
    .D(_0007_),
    .Q_N(_0122_),
    .Q(\Pong.control_unit.NES_Controller_Left.state_NESController[16] ));
 sg13g2_dfrbp_1 \Pong.control_unit.NES_Controller_Left.state_NESController[17]$_DFF_P_  (.CLK(clknet_5_18__leaf_clk),
    .RESET_B(net205),
    .D(_0008_),
    .Q_N(_0120_),
    .Q(\Pong.control_unit.NES_Controller_Left.state_NESController[17] ));
 sg13g2_dfrbp_1 \Pong.control_unit.NES_Controller_Left.state_NESController[18]$_DFF_P_  (.CLK(clknet_5_0__leaf_clk),
    .RESET_B(net206),
    .D(_0009_),
    .Q_N(_3170_),
    .Q(\Pong.control_unit.NES_Controller_Left.state_NESController[18] ));
 sg13g2_dfrbp_1 \Pong.control_unit.NES_Controller_Left.state_NESController[1]$_DFF_P_  (.CLK(clknet_5_4__leaf_clk),
    .RESET_B(net207),
    .D(_0010_),
    .Q_N(_3171_),
    .Q(\Pong.control_unit.NES_Controller_Left.state_NESController[1] ));
 sg13g2_dfrbp_1 \Pong.control_unit.NES_Controller_Left.state_NESController[2]$_DFF_P_  (.CLK(clknet_5_7__leaf_clk),
    .RESET_B(net208),
    .D(_0011_),
    .Q_N(_0121_),
    .Q(\Pong.control_unit.NES_Controller_Left.state_NESController[2] ));
 sg13g2_dfrbp_1 \Pong.control_unit.NES_Controller_Left.state_NESController[3]$_DFF_P_  (.CLK(clknet_5_18__leaf_clk),
    .RESET_B(net209),
    .D(_0012_),
    .Q_N(_3172_),
    .Q(\Pong.control_unit.NES_Controller_Left.state_NESController[3] ));
 sg13g2_dfrbp_1 \Pong.control_unit.NES_Controller_Left.state_NESController[4]$_DFF_P_  (.CLK(clknet_5_6__leaf_clk),
    .RESET_B(net210),
    .D(_0013_),
    .Q_N(_0123_),
    .Q(\Pong.control_unit.NES_Controller_Left.state_NESController[4] ));
 sg13g2_dfrbp_1 \Pong.control_unit.NES_Controller_Left.state_NESController[5]$_DFF_P_  (.CLK(clknet_5_5__leaf_clk),
    .RESET_B(net211),
    .D(_0014_),
    .Q_N(_3173_),
    .Q(\Pong.control_unit.NES_Controller_Left.state_NESController[5] ));
 sg13g2_dfrbp_1 \Pong.control_unit.NES_Controller_Left.state_NESController[6]$_DFF_P_  (.CLK(clknet_5_0__leaf_clk),
    .RESET_B(net212),
    .D(_0015_),
    .Q_N(_3174_),
    .Q(\Pong.control_unit.NES_Controller_Left.state_NESController[6] ));
 sg13g2_dfrbp_1 \Pong.control_unit.NES_Controller_Left.state_NESController[7]$_DFF_P_  (.CLK(clknet_5_7__leaf_clk),
    .RESET_B(net213),
    .D(_0016_),
    .Q_N(_0126_),
    .Q(\Pong.control_unit.NES_Controller_Left.state_NESController[7] ));
 sg13g2_dfrbp_1 \Pong.control_unit.NES_Controller_Left.state_NESController[8]$_DFF_P_  (.CLK(clknet_5_7__leaf_clk),
    .RESET_B(net214),
    .D(_0017_),
    .Q_N(_3175_),
    .Q(\Pong.control_unit.NES_Controller_Left.state_NESController[8] ));
 sg13g2_dfrbp_1 \Pong.control_unit.NES_Controller_Left.state_NESController[9]$_DFF_P_  (.CLK(clknet_5_0__leaf_clk),
    .RESET_B(net215),
    .D(_0018_),
    .Q_N(_3176_),
    .Q(\Pong.control_unit.NES_Controller_Left.state_NESController[9] ));
 sg13g2_dfrbp_1 \Pong.control_unit.NES_Controller_Right.state_NESController[0]$_DFF_P_  (.CLK(clknet_5_20__leaf_clk),
    .RESET_B(net216),
    .D(_0019_),
    .Q_N(_0127_),
    .Q(\Pong.control_unit.NES_Controller_Right.state_NESController[0] ));
 sg13g2_dfrbp_1 \Pong.control_unit.NES_Controller_Right.state_NESController[10]$_DFF_P_  (.CLK(clknet_5_22__leaf_clk),
    .RESET_B(net217),
    .D(_0020_),
    .Q_N(_3177_),
    .Q(\Pong.control_unit.NES_Controller_Right.state_NESController[10] ));
 sg13g2_dfrbp_1 \Pong.control_unit.NES_Controller_Right.state_NESController[11]$_DFF_P_  (.CLK(clknet_5_19__leaf_clk),
    .RESET_B(net218),
    .D(_0021_),
    .Q_N(_3178_),
    .Q(\Pong.control_unit.NES_Controller_Right.state_NESController[11] ));
 sg13g2_dfrbp_1 \Pong.control_unit.NES_Controller_Right.state_NESController[12]$_DFF_P_  (.CLK(clknet_5_22__leaf_clk),
    .RESET_B(net219),
    .D(_0022_),
    .Q_N(_0133_),
    .Q(\Pong.control_unit.NES_Controller_Right.state_NESController[12] ));
 sg13g2_dfrbp_1 \Pong.control_unit.NES_Controller_Right.state_NESController[13]$_DFF_P_  (.CLK(clknet_5_23__leaf_clk),
    .RESET_B(net220),
    .D(_0023_),
    .Q_N(_3179_),
    .Q(\Pong.control_unit.NES_Controller_Right.state_NESController[13] ));
 sg13g2_dfrbp_1 \Pong.control_unit.NES_Controller_Right.state_NESController[14]$_DFF_P_  (.CLK(clknet_5_19__leaf_clk),
    .RESET_B(net221),
    .D(_0024_),
    .Q_N(_0132_),
    .Q(\Pong.control_unit.NES_Controller_Right.state_NESController[14] ));
 sg13g2_dfrbp_1 \Pong.control_unit.NES_Controller_Right.state_NESController[15]$_DFF_P_  (.CLK(clknet_5_23__leaf_clk),
    .RESET_B(net222),
    .D(_0025_),
    .Q_N(_3180_),
    .Q(\Pong.control_unit.NES_Controller_Right.state_NESController[15] ));
 sg13g2_dfrbp_1 \Pong.control_unit.NES_Controller_Right.state_NESController[16]$_DFF_P_  (.CLK(clknet_5_25__leaf_clk),
    .RESET_B(net223),
    .D(_0026_),
    .Q_N(_0130_),
    .Q(\Pong.control_unit.NES_Controller_Right.state_NESController[16] ));
 sg13g2_dfrbp_1 \Pong.control_unit.NES_Controller_Right.state_NESController[17]$_DFF_P_  (.CLK(clknet_5_23__leaf_clk),
    .RESET_B(net224),
    .D(_0027_),
    .Q_N(_0128_),
    .Q(\Pong.control_unit.NES_Controller_Right.state_NESController[17] ));
 sg13g2_dfrbp_1 \Pong.control_unit.NES_Controller_Right.state_NESController[18]$_DFF_P_  (.CLK(clknet_5_19__leaf_clk),
    .RESET_B(net225),
    .D(_0028_),
    .Q_N(_3181_),
    .Q(\Pong.control_unit.NES_Controller_Right.state_NESController[18] ));
 sg13g2_dfrbp_1 \Pong.control_unit.NES_Controller_Right.state_NESController[1]$_DFF_P_  (.CLK(clknet_5_18__leaf_clk),
    .RESET_B(net226),
    .D(_0029_),
    .Q_N(_3182_),
    .Q(\Pong.control_unit.NES_Controller_Right.state_NESController[1] ));
 sg13g2_dfrbp_1 \Pong.control_unit.NES_Controller_Right.state_NESController[2]$_DFF_P_  (.CLK(clknet_5_22__leaf_clk),
    .RESET_B(net227),
    .D(_0030_),
    .Q_N(_0129_),
    .Q(\Pong.control_unit.NES_Controller_Right.state_NESController[2] ));
 sg13g2_dfrbp_1 \Pong.control_unit.NES_Controller_Right.state_NESController[3]$_DFF_P_  (.CLK(clknet_5_23__leaf_clk),
    .RESET_B(net228),
    .D(_0031_),
    .Q_N(_3183_),
    .Q(\Pong.control_unit.NES_Controller_Right.state_NESController[3] ));
 sg13g2_dfrbp_1 \Pong.control_unit.NES_Controller_Right.state_NESController[4]$_DFF_P_  (.CLK(clknet_5_19__leaf_clk),
    .RESET_B(net229),
    .D(_0032_),
    .Q_N(_0131_),
    .Q(\Pong.control_unit.NES_Controller_Right.state_NESController[4] ));
 sg13g2_dfrbp_1 \Pong.control_unit.NES_Controller_Right.state_NESController[5]$_DFF_P_  (.CLK(clknet_5_22__leaf_clk),
    .RESET_B(net230),
    .D(_0033_),
    .Q_N(_3184_),
    .Q(\Pong.control_unit.NES_Controller_Right.state_NESController[5] ));
 sg13g2_dfrbp_1 \Pong.control_unit.NES_Controller_Right.state_NESController[6]$_DFF_P_  (.CLK(clknet_5_19__leaf_clk),
    .RESET_B(net231),
    .D(_0034_),
    .Q_N(_3185_),
    .Q(\Pong.control_unit.NES_Controller_Right.state_NESController[6] ));
 sg13g2_dfrbp_1 \Pong.control_unit.NES_Controller_Right.state_NESController[7]$_DFF_P_  (.CLK(clknet_5_22__leaf_clk),
    .RESET_B(net232),
    .D(_0035_),
    .Q_N(_0134_),
    .Q(\Pong.control_unit.NES_Controller_Right.state_NESController[7] ));
 sg13g2_dfrbp_1 \Pong.control_unit.NES_Controller_Right.state_NESController[8]$_DFF_P_  (.CLK(clknet_5_22__leaf_clk),
    .RESET_B(net233),
    .D(_0036_),
    .Q_N(_3186_),
    .Q(\Pong.control_unit.NES_Controller_Right.state_NESController[8] ));
 sg13g2_dfrbp_1 \Pong.control_unit.NES_Controller_Right.state_NESController[9]$_DFF_P_  (.CLK(clknet_5_19__leaf_clk),
    .RESET_B(net234),
    .D(_0037_),
    .Q_N(_3187_),
    .Q(\Pong.control_unit.NES_Controller_Right.state_NESController[9] ));
 sg13g2_dfrbp_1 \Pong.control_unit.state_ballMovement[0]$_DFF_P_  (.CLK(clknet_5_10__leaf_clk),
    .RESET_B(net235),
    .D(_0038_),
    .Q_N(_3188_),
    .Q(\Pong.control_unit.state_ballMovement[0] ));
 sg13g2_dfrbp_1 \Pong.control_unit.state_ballMovement[1]$_DFF_P_  (.CLK(clknet_5_10__leaf_clk),
    .RESET_B(net236),
    .D(_0039_),
    .Q_N(_3189_),
    .Q(\Pong.control_unit.state_ballMovement[1] ));
 sg13g2_dfrbp_1 \Pong.control_unit.state_ballMovement[2]$_DFF_P_  (.CLK(clknet_5_10__leaf_clk),
    .RESET_B(net237),
    .D(_0040_),
    .Q_N(_3190_),
    .Q(\Pong.control_unit.state_ballMovement[2] ));
 sg13g2_dfrbp_1 \Pong.control_unit.state_ballMovement[3]$_DFF_P_  (.CLK(clknet_5_11__leaf_clk),
    .RESET_B(net238),
    .D(_0041_),
    .Q_N(_0115_),
    .Q(\Pong.control_unit.state_ballMovement[3] ));
 sg13g2_dfrbp_1 \Pong.control_unit.state_ballMovement[4]$_DFF_P_  (.CLK(clknet_5_11__leaf_clk),
    .RESET_B(net239),
    .D(_0042_),
    .Q_N(_3165_),
    .Q(\Pong.control_unit.state_ballMovement[4] ));
 sg13g2_dfrbp_1 \Pong.datapath.Ball_Clock.processQ[0]$_SDFFE_PN0P_  (.CLK(clknet_5_3__leaf_clk),
    .RESET_B(net240),
    .D(_0135_),
    .Q_N(_3164_),
    .Q(\Pong.datapath.Ball_Clock.Q[0] ));
 sg13g2_dfrbp_1 \Pong.datapath.Ball_Clock.processQ[10]$_SDFFE_PN0P_  (.CLK(clknet_5_8__leaf_clk),
    .RESET_B(net241),
    .D(_0136_),
    .Q_N(_3163_),
    .Q(\Pong.datapath.Ball_Clock.Q[10] ));
 sg13g2_dfrbp_1 \Pong.datapath.Ball_Clock.processQ[11]$_SDFFE_PN0P_  (.CLK(clknet_5_8__leaf_clk),
    .RESET_B(net242),
    .D(_0137_),
    .Q_N(_3162_),
    .Q(\Pong.datapath.Ball_Clock.Q[11] ));
 sg13g2_dfrbp_1 \Pong.datapath.Ball_Clock.processQ[12]$_SDFFE_PN0P_  (.CLK(clknet_5_8__leaf_clk),
    .RESET_B(net243),
    .D(_0138_),
    .Q_N(_3161_),
    .Q(\Pong.datapath.Ball_Clock.Q[12] ));
 sg13g2_dfrbp_1 \Pong.datapath.Ball_Clock.processQ[13]$_SDFFE_PN0P_  (.CLK(clknet_5_8__leaf_clk),
    .RESET_B(net244),
    .D(_0139_),
    .Q_N(_3160_),
    .Q(\Pong.datapath.Ball_Clock.Q[13] ));
 sg13g2_dfrbp_1 \Pong.datapath.Ball_Clock.processQ[14]$_SDFFE_PN0P_  (.CLK(clknet_5_10__leaf_clk),
    .RESET_B(net245),
    .D(_0140_),
    .Q_N(_3159_),
    .Q(\Pong.datapath.Ball_Clock.Q[14] ));
 sg13g2_dfrbp_1 \Pong.datapath.Ball_Clock.processQ[15]$_SDFFE_PN0P_  (.CLK(clknet_5_9__leaf_clk),
    .RESET_B(net246),
    .D(_0141_),
    .Q_N(_3158_),
    .Q(\Pong.datapath.Ball_Clock.Q[15] ));
 sg13g2_dfrbp_1 \Pong.datapath.Ball_Clock.processQ[16]$_SDFFE_PN0P_  (.CLK(clknet_5_9__leaf_clk),
    .RESET_B(net247),
    .D(_0142_),
    .Q_N(_3157_),
    .Q(\Pong.datapath.Ball_Clock.Q[16] ));
 sg13g2_dfrbp_1 \Pong.datapath.Ball_Clock.processQ[1]$_SDFFE_PN0P_  (.CLK(clknet_5_3__leaf_clk),
    .RESET_B(net248),
    .D(_0143_),
    .Q_N(_3156_),
    .Q(\Pong.datapath.Ball_Clock.Q[1] ));
 sg13g2_dfrbp_1 \Pong.datapath.Ball_Clock.processQ[2]$_SDFFE_PN0P_  (.CLK(clknet_5_2__leaf_clk),
    .RESET_B(net249),
    .D(_0144_),
    .Q_N(_3155_),
    .Q(\Pong.datapath.Ball_Clock.Q[2] ));
 sg13g2_dfrbp_1 \Pong.datapath.Ball_Clock.processQ[3]$_SDFFE_PN0P_  (.CLK(clknet_5_2__leaf_clk),
    .RESET_B(net250),
    .D(_0145_),
    .Q_N(_3154_),
    .Q(\Pong.datapath.Ball_Clock.Q[3] ));
 sg13g2_dfrbp_1 \Pong.datapath.Ball_Clock.processQ[4]$_SDFFE_PN0P_  (.CLK(clknet_5_2__leaf_clk),
    .RESET_B(net251),
    .D(_0146_),
    .Q_N(_3153_),
    .Q(\Pong.datapath.Ball_Clock.Q[4] ));
 sg13g2_dfrbp_1 \Pong.datapath.Ball_Clock.processQ[5]$_SDFFE_PN0P_  (.CLK(clknet_5_2__leaf_clk),
    .RESET_B(net252),
    .D(_0147_),
    .Q_N(_3152_),
    .Q(\Pong.datapath.Ball_Clock.Q[5] ));
 sg13g2_dfrbp_1 \Pong.datapath.Ball_Clock.processQ[6]$_SDFFE_PN0P_  (.CLK(clknet_5_2__leaf_clk),
    .RESET_B(net253),
    .D(_0148_),
    .Q_N(_3151_),
    .Q(\Pong.datapath.Ball_Clock.Q[6] ));
 sg13g2_dfrbp_1 \Pong.datapath.Ball_Clock.processQ[7]$_SDFFE_PN0P_  (.CLK(clknet_5_2__leaf_clk),
    .RESET_B(net254),
    .D(_0149_),
    .Q_N(_3150_),
    .Q(\Pong.datapath.Ball_Clock.Q[7] ));
 sg13g2_dfrbp_1 \Pong.datapath.Ball_Clock.processQ[8]$_SDFFE_PN0P_  (.CLK(clknet_5_9__leaf_clk),
    .RESET_B(net255),
    .D(_0150_),
    .Q_N(_0056_),
    .Q(\Pong.datapath.Ball_Clock.Q[8] ));
 sg13g2_dfrbp_1 \Pong.datapath.Ball_Clock.processQ[9]$_SDFFE_PN0P_  (.CLK(clknet_5_8__leaf_clk),
    .RESET_B(net256),
    .D(_0151_),
    .Q_N(_3149_),
    .Q(\Pong.datapath.Ball_Clock.Q[9] ));
 sg13g2_dfrbp_1 \Pong.datapath.NES_activity_Left[2]$_SDFF_PP0_  (.CLK(clknet_5_30__leaf_clk),
    .RESET_B(net257),
    .D(_0152_),
    .Q_N(_3148_),
    .Q(\Pong.datapath.NES_activity_Left[2] ));
 sg13g2_dfrbp_1 \Pong.datapath.NES_activity_Left[3]$_SDFF_PP0_  (.CLK(clknet_5_29__leaf_clk),
    .RESET_B(net258),
    .D(_0153_),
    .Q_N(_3147_),
    .Q(\Pong.datapath.NES_activity_Left[3] ));
 sg13g2_dfrbp_1 \Pong.datapath.NES_activity_Left[4]$_SDFF_PP0_  (.CLK(clknet_5_25__leaf_clk),
    .RESET_B(net259),
    .D(_0154_),
    .Q_N(_3146_),
    .Q(\Pong.datapath.NES_activity_Left[4] ));
 sg13g2_dfrbp_1 \Pong.datapath.NES_activity_Left[5]$_SDFF_PP0_  (.CLK(clknet_5_26__leaf_clk),
    .RESET_B(net260),
    .D(_0155_),
    .Q_N(_3145_),
    .Q(\Pong.datapath.NES_activity_Left[5] ));
 sg13g2_dfrbp_1 \Pong.datapath.NES_activity_Right[2]$_SDFF_PP0_  (.CLK(clknet_5_27__leaf_clk),
    .RESET_B(net261),
    .D(_0156_),
    .Q_N(_3144_),
    .Q(\Pong.datapath.NES_activity_Right[2] ));
 sg13g2_dfrbp_1 \Pong.datapath.NES_activity_Right[3]$_SDFF_PP0_  (.CLK(clknet_5_29__leaf_clk),
    .RESET_B(net262),
    .D(_0157_),
    .Q_N(_3143_),
    .Q(\Pong.datapath.NES_activity_Right[3] ));
 sg13g2_dfrbp_1 \Pong.datapath.NES_activity_Right[4]$_SDFF_PP0_  (.CLK(clknet_5_27__leaf_clk),
    .RESET_B(net263),
    .D(_0158_),
    .Q_N(_3142_),
    .Q(\Pong.datapath.NES_activity_Right[4] ));
 sg13g2_dfrbp_1 \Pong.datapath.NES_activity_Right[5]$_SDFF_PP0_  (.CLK(clknet_5_26__leaf_clk),
    .RESET_B(net264),
    .D(_0159_),
    .Q_N(_0081_),
    .Q(\Pong.datapath.NES_activity_Right[5] ));
 sg13g2_dfrbp_1 \Pong.datapath.NES_counter_left.processQ[0]$_SDFFE_PP0P_  (.CLK(clknet_5_13__leaf_clk),
    .RESET_B(net265),
    .D(_0160_),
    .Q_N(_3141_),
    .Q(\Pong.datapath.NES_counter_left.Q[0] ));
 sg13g2_dfrbp_1 \Pong.datapath.NES_counter_left.processQ[1]$_SDFFE_PP0P_  (.CLK(clknet_5_9__leaf_clk),
    .RESET_B(net266),
    .D(_0161_),
    .Q_N(_3140_),
    .Q(\Pong.datapath.NES_counter_left.Q[1] ));
 sg13g2_dfrbp_1 \Pong.datapath.NES_counter_left.processQ[2]$_SDFFE_PP0P_  (.CLK(clknet_5_12__leaf_clk),
    .RESET_B(net267),
    .D(_0162_),
    .Q_N(_3139_),
    .Q(\Pong.datapath.NES_counter_left.Q[2] ));
 sg13g2_dfrbp_1 \Pong.datapath.NES_counter_left.processQ[3]$_SDFFE_PP0P_  (.CLK(clknet_5_13__leaf_clk),
    .RESET_B(net268),
    .D(_0163_),
    .Q_N(_3138_),
    .Q(\Pong.datapath.NES_counter_left.Q[3] ));
 sg13g2_dfrbp_1 \Pong.datapath.NES_counter_left.processQ[4]$_SDFFE_PP0P_  (.CLK(clknet_5_12__leaf_clk),
    .RESET_B(net269),
    .D(_0164_),
    .Q_N(_3137_),
    .Q(\Pong.datapath.NES_counter_left.Q[4] ));
 sg13g2_dfrbp_1 \Pong.datapath.NES_counter_left.processQ[5]$_SDFFE_PP0P_  (.CLK(clknet_5_13__leaf_clk),
    .RESET_B(net270),
    .D(_0165_),
    .Q_N(_3136_),
    .Q(\Pong.datapath.NES_counter_left.Q[5] ));
 sg13g2_dfrbp_1 \Pong.datapath.NES_counter_left.processQ[6]$_SDFFE_PP0P_  (.CLK(clknet_5_0__leaf_clk),
    .RESET_B(net271),
    .D(_0166_),
    .Q_N(_3135_),
    .Q(\Pong.datapath.NES_counter_left.Q[6] ));
 sg13g2_dfrbp_1 \Pong.datapath.NES_counter_left.processQ[7]$_SDFFE_PP0P_  (.CLK(clknet_5_0__leaf_clk),
    .RESET_B(net272),
    .D(_0167_),
    .Q_N(_3134_),
    .Q(\Pong.datapath.NES_counter_left.Q[7] ));
 sg13g2_dfrbp_1 \Pong.datapath.NES_counter_right.processQ[0]$_SDFFE_PP0P_  (.CLK(clknet_5_21__leaf_clk),
    .RESET_B(net273),
    .D(_0168_),
    .Q_N(_3133_),
    .Q(\Pong.datapath.NES_counter_right.Q[0] ));
 sg13g2_dfrbp_1 \Pong.datapath.NES_counter_right.processQ[1]$_SDFFE_PP0P_  (.CLK(clknet_5_21__leaf_clk),
    .RESET_B(net274),
    .D(_0169_),
    .Q_N(_3132_),
    .Q(\Pong.datapath.NES_counter_right.Q[1] ));
 sg13g2_dfrbp_1 \Pong.datapath.NES_counter_right.processQ[2]$_SDFFE_PP0P_  (.CLK(clknet_5_21__leaf_clk),
    .RESET_B(net275),
    .D(_0170_),
    .Q_N(_3131_),
    .Q(\Pong.datapath.NES_counter_right.Q[2] ));
 sg13g2_dfrbp_1 \Pong.datapath.NES_counter_right.processQ[3]$_SDFFE_PP0P_  (.CLK(clknet_5_20__leaf_clk),
    .RESET_B(net276),
    .D(_0171_),
    .Q_N(_3130_),
    .Q(\Pong.datapath.NES_counter_right.Q[3] ));
 sg13g2_dfrbp_1 \Pong.datapath.NES_counter_right.processQ[4]$_SDFFE_PP0P_  (.CLK(clknet_5_21__leaf_clk),
    .RESET_B(net277),
    .D(_0172_),
    .Q_N(_3129_),
    .Q(\Pong.datapath.NES_counter_right.Q[4] ));
 sg13g2_dfrbp_1 \Pong.datapath.NES_counter_right.processQ[5]$_SDFFE_PP0P_  (.CLK(clknet_5_21__leaf_clk),
    .RESET_B(net278),
    .D(_0173_),
    .Q_N(_3128_),
    .Q(\Pong.datapath.NES_counter_right.Q[5] ));
 sg13g2_dfrbp_1 \Pong.datapath.NES_counter_right.processQ[6]$_SDFFE_PP0P_  (.CLK(clknet_5_21__leaf_clk),
    .RESET_B(net279),
    .D(_0174_),
    .Q_N(_3127_),
    .Q(\Pong.datapath.NES_counter_right.Q[6] ));
 sg13g2_dfrbp_1 \Pong.datapath.NES_counter_right.processQ[7]$_SDFFE_PP0P_  (.CLK(clknet_5_23__leaf_clk),
    .RESET_B(net280),
    .D(_0175_),
    .Q_N(_3126_),
    .Q(\Pong.datapath.NES_counter_right.Q[7] ));
 sg13g2_dfrbp_1 \Pong.datapath.NES_delay_counter_left.processQ[0]$_SDFFE_PN0P_  (.CLK(clknet_5_4__leaf_clk),
    .RESET_B(net281),
    .D(_0176_),
    .Q_N(_3125_),
    .Q(\Pong.datapath.NES_delay_counter_left.Q[0] ));
 sg13g2_dfrbp_1 \Pong.datapath.NES_delay_counter_left.processQ[10]$_SDFFE_PN0P_  (.CLK(clknet_5_1__leaf_clk),
    .RESET_B(net282),
    .D(_0177_),
    .Q_N(_3124_),
    .Q(\Pong.datapath.NES_delay_counter_left.Q[10] ));
 sg13g2_dfrbp_1 \Pong.datapath.NES_delay_counter_left.processQ[11]$_SDFFE_PN0P_  (.CLK(clknet_5_3__leaf_clk),
    .RESET_B(net283),
    .D(_0178_),
    .Q_N(_3123_),
    .Q(\Pong.datapath.NES_delay_counter_left.Q[11] ));
 sg13g2_dfrbp_1 \Pong.datapath.NES_delay_counter_left.processQ[12]$_SDFFE_PN0P_  (.CLK(clknet_5_3__leaf_clk),
    .RESET_B(net284),
    .D(_0179_),
    .Q_N(_3122_),
    .Q(\Pong.datapath.NES_delay_counter_left.Q[12] ));
 sg13g2_dfrbp_1 \Pong.datapath.NES_delay_counter_left.processQ[13]$_SDFFE_PN0P_  (.CLK(clknet_5_3__leaf_clk),
    .RESET_B(net285),
    .D(_0180_),
    .Q_N(_3121_),
    .Q(\Pong.datapath.NES_delay_counter_left.Q[13] ));
 sg13g2_dfrbp_1 \Pong.datapath.NES_delay_counter_left.processQ[14]$_SDFFE_PN0P_  (.CLK(clknet_5_9__leaf_clk),
    .RESET_B(net286),
    .D(_0181_),
    .Q_N(_3120_),
    .Q(\Pong.datapath.NES_delay_counter_left.Q[14] ));
 sg13g2_dfrbp_1 \Pong.datapath.NES_delay_counter_left.processQ[15]$_SDFFE_PN0P_  (.CLK(clknet_5_9__leaf_clk),
    .RESET_B(net287),
    .D(_0182_),
    .Q_N(_3119_),
    .Q(\Pong.datapath.NES_delay_counter_left.Q[15] ));
 sg13g2_dfrbp_1 \Pong.datapath.NES_delay_counter_left.processQ[16]$_SDFFE_PN0P_  (.CLK(clknet_5_13__leaf_clk),
    .RESET_B(net288),
    .D(_0183_),
    .Q_N(_3118_),
    .Q(\Pong.datapath.NES_delay_counter_left.Q[16] ));
 sg13g2_dfrbp_1 \Pong.datapath.NES_delay_counter_left.processQ[17]$_SDFFE_PN0P_  (.CLK(clknet_5_3__leaf_clk),
    .RESET_B(net289),
    .D(_0184_),
    .Q_N(_3117_),
    .Q(\Pong.datapath.NES_delay_counter_left.Q[17] ));
 sg13g2_dfrbp_1 \Pong.datapath.NES_delay_counter_left.processQ[18]$_SDFFE_PN0P_  (.CLK(clknet_5_0__leaf_clk),
    .RESET_B(net290),
    .D(_0185_),
    .Q_N(_0117_),
    .Q(\Pong.datapath.NES_delay_counter_left.Q[18] ));
 sg13g2_dfrbp_1 \Pong.datapath.NES_delay_counter_left.processQ[1]$_SDFFE_PN0P_  (.CLK(clknet_5_4__leaf_clk),
    .RESET_B(net291),
    .D(_0186_),
    .Q_N(_3116_),
    .Q(\Pong.datapath.NES_delay_counter_left.Q[1] ));
 sg13g2_dfrbp_1 \Pong.datapath.NES_delay_counter_left.processQ[2]$_SDFFE_PN0P_  (.CLK(clknet_5_1__leaf_clk),
    .RESET_B(net292),
    .D(_0187_),
    .Q_N(_3115_),
    .Q(\Pong.datapath.NES_delay_counter_left.Q[2] ));
 sg13g2_dfrbp_1 \Pong.datapath.NES_delay_counter_left.processQ[3]$_SDFFE_PN0P_  (.CLK(clknet_5_5__leaf_clk),
    .RESET_B(net293),
    .D(_0188_),
    .Q_N(_3114_),
    .Q(\Pong.datapath.NES_delay_counter_left.Q[3] ));
 sg13g2_dfrbp_1 \Pong.datapath.NES_delay_counter_left.processQ[4]$_SDFFE_PN0P_  (.CLK(clknet_5_4__leaf_clk),
    .RESET_B(net294),
    .D(_0189_),
    .Q_N(_3113_),
    .Q(\Pong.datapath.NES_delay_counter_left.Q[4] ));
 sg13g2_dfrbp_1 \Pong.datapath.NES_delay_counter_left.processQ[5]$_SDFFE_PN0P_  (.CLK(clknet_5_4__leaf_clk),
    .RESET_B(net295),
    .D(_0190_),
    .Q_N(_3112_),
    .Q(\Pong.datapath.NES_delay_counter_left.Q[5] ));
 sg13g2_dfrbp_1 \Pong.datapath.NES_delay_counter_left.processQ[6]$_SDFFE_PN0P_  (.CLK(clknet_5_1__leaf_clk),
    .RESET_B(net296),
    .D(_0191_),
    .Q_N(_3111_),
    .Q(\Pong.datapath.NES_delay_counter_left.Q[6] ));
 sg13g2_dfrbp_1 \Pong.datapath.NES_delay_counter_left.processQ[7]$_SDFFE_PN0P_  (.CLK(clknet_5_1__leaf_clk),
    .RESET_B(net297),
    .D(_0192_),
    .Q_N(_3110_),
    .Q(\Pong.datapath.NES_delay_counter_left.Q[7] ));
 sg13g2_dfrbp_1 \Pong.datapath.NES_delay_counter_left.processQ[8]$_SDFFE_PN0P_  (.CLK(clknet_5_1__leaf_clk),
    .RESET_B(net298),
    .D(_0193_),
    .Q_N(_0118_),
    .Q(\Pong.datapath.NES_delay_counter_left.Q[8] ));
 sg13g2_dfrbp_1 \Pong.datapath.NES_delay_counter_left.processQ[9]$_SDFFE_PN0P_  (.CLK(clknet_5_1__leaf_clk),
    .RESET_B(net299),
    .D(_0194_),
    .Q_N(_3109_),
    .Q(\Pong.datapath.NES_delay_counter_left.Q[9] ));
 sg13g2_dfrbp_1 \Pong.datapath.NES_delay_counter_right.processQ[0]$_SDFFE_PN0P_  (.CLK(clknet_5_16__leaf_clk),
    .RESET_B(net300),
    .D(_0195_),
    .Q_N(_3108_),
    .Q(\Pong.datapath.NES_delay_counter_right.Q[0] ));
 sg13g2_dfrbp_1 \Pong.datapath.NES_delay_counter_right.processQ[10]$_SDFFE_PN0P_  (.CLK(clknet_5_20__leaf_clk),
    .RESET_B(net301),
    .D(_0196_),
    .Q_N(_3107_),
    .Q(\Pong.datapath.NES_delay_counter_right.Q[10] ));
 sg13g2_dfrbp_1 \Pong.datapath.NES_delay_counter_right.processQ[11]$_SDFFE_PN0P_  (.CLK(clknet_5_20__leaf_clk),
    .RESET_B(net302),
    .D(_0197_),
    .Q_N(_3106_),
    .Q(\Pong.datapath.NES_delay_counter_right.Q[11] ));
 sg13g2_dfrbp_1 \Pong.datapath.NES_delay_counter_right.processQ[12]$_SDFFE_PN0P_  (.CLK(clknet_5_20__leaf_clk),
    .RESET_B(net303),
    .D(_0198_),
    .Q_N(_3105_),
    .Q(\Pong.datapath.NES_delay_counter_right.Q[12] ));
 sg13g2_dfrbp_1 \Pong.datapath.NES_delay_counter_right.processQ[13]$_SDFFE_PN0P_  (.CLK(clknet_5_20__leaf_clk),
    .RESET_B(net304),
    .D(_0199_),
    .Q_N(_3104_),
    .Q(\Pong.datapath.NES_delay_counter_right.Q[13] ));
 sg13g2_dfrbp_1 \Pong.datapath.NES_delay_counter_right.processQ[14]$_SDFFE_PN0P_  (.CLK(clknet_5_17__leaf_clk),
    .RESET_B(net305),
    .D(_0200_),
    .Q_N(_3103_),
    .Q(\Pong.datapath.NES_delay_counter_right.Q[14] ));
 sg13g2_dfrbp_1 \Pong.datapath.NES_delay_counter_right.processQ[15]$_SDFFE_PN0P_  (.CLK(clknet_5_17__leaf_clk),
    .RESET_B(net306),
    .D(_0201_),
    .Q_N(_3102_),
    .Q(\Pong.datapath.NES_delay_counter_right.Q[15] ));
 sg13g2_dfrbp_1 \Pong.datapath.NES_delay_counter_right.processQ[16]$_SDFFE_PN0P_  (.CLK(clknet_5_17__leaf_clk),
    .RESET_B(net307),
    .D(_0202_),
    .Q_N(_3101_),
    .Q(\Pong.datapath.NES_delay_counter_right.Q[16] ));
 sg13g2_dfrbp_1 \Pong.datapath.NES_delay_counter_right.processQ[17]$_SDFFE_PN0P_  (.CLK(clknet_5_18__leaf_clk),
    .RESET_B(net308),
    .D(_0203_),
    .Q_N(_3100_),
    .Q(\Pong.datapath.NES_delay_counter_right.Q[17] ));
 sg13g2_dfrbp_1 \Pong.datapath.NES_delay_counter_right.processQ[18]$_SDFFE_PN0P_  (.CLK(clknet_5_17__leaf_clk),
    .RESET_B(net309),
    .D(_0204_),
    .Q_N(_0110_),
    .Q(\Pong.datapath.NES_delay_counter_right.Q[18] ));
 sg13g2_dfrbp_1 \Pong.datapath.NES_delay_counter_right.processQ[1]$_SDFFE_PN0P_  (.CLK(clknet_5_16__leaf_clk),
    .RESET_B(net310),
    .D(_0205_),
    .Q_N(_3099_),
    .Q(\Pong.datapath.NES_delay_counter_right.Q[1] ));
 sg13g2_dfrbp_1 \Pong.datapath.NES_delay_counter_right.processQ[2]$_SDFFE_PN0P_  (.CLK(clknet_5_16__leaf_clk),
    .RESET_B(net311),
    .D(_0206_),
    .Q_N(_3098_),
    .Q(\Pong.datapath.NES_delay_counter_right.Q[2] ));
 sg13g2_dfrbp_1 \Pong.datapath.NES_delay_counter_right.processQ[3]$_SDFFE_PN0P_  (.CLK(clknet_5_5__leaf_clk),
    .RESET_B(net312),
    .D(_0207_),
    .Q_N(_3097_),
    .Q(\Pong.datapath.NES_delay_counter_right.Q[3] ));
 sg13g2_dfrbp_1 \Pong.datapath.NES_delay_counter_right.processQ[4]$_SDFFE_PN0P_  (.CLK(clknet_5_5__leaf_clk),
    .RESET_B(net313),
    .D(_0208_),
    .Q_N(_3096_),
    .Q(\Pong.datapath.NES_delay_counter_right.Q[4] ));
 sg13g2_dfrbp_1 \Pong.datapath.NES_delay_counter_right.processQ[5]$_SDFFE_PN0P_  (.CLK(clknet_5_16__leaf_clk),
    .RESET_B(net314),
    .D(_0209_),
    .Q_N(_3095_),
    .Q(\Pong.datapath.NES_delay_counter_right.Q[5] ));
 sg13g2_dfrbp_1 \Pong.datapath.NES_delay_counter_right.processQ[6]$_SDFFE_PN0P_  (.CLK(clknet_5_16__leaf_clk),
    .RESET_B(net315),
    .D(_0210_),
    .Q_N(_3094_),
    .Q(\Pong.datapath.NES_delay_counter_right.Q[6] ));
 sg13g2_dfrbp_1 \Pong.datapath.NES_delay_counter_right.processQ[7]$_SDFFE_PN0P_  (.CLK(clknet_5_16__leaf_clk),
    .RESET_B(net316),
    .D(_0211_),
    .Q_N(_3093_),
    .Q(\Pong.datapath.NES_delay_counter_right.Q[7] ));
 sg13g2_dfrbp_1 \Pong.datapath.NES_delay_counter_right.processQ[8]$_SDFFE_PN0P_  (.CLK(clknet_5_17__leaf_clk),
    .RESET_B(net317),
    .D(_0212_),
    .Q_N(_0116_),
    .Q(\Pong.datapath.NES_delay_counter_right.Q[8] ));
 sg13g2_dfrbp_1 \Pong.datapath.NES_delay_counter_right.processQ[9]$_SDFFE_PN0P_  (.CLK(clknet_5_17__leaf_clk),
    .RESET_B(net318),
    .D(_0213_),
    .Q_N(_3092_),
    .Q(\Pong.datapath.NES_delay_counter_right.Q[9] ));
 sg13g2_dfrbp_1 \Pong.datapath.NES_wire_Left[2]$_SDFFE_PN0N_  (.CLK(clknet_5_24__leaf_clk),
    .RESET_B(net319),
    .D(_0214_),
    .Q_N(_0048_),
    .Q(\Pong.datapath.NES_wire_Left[2] ));
 sg13g2_dfrbp_1 \Pong.datapath.NES_wire_Left[3]$_SDFFE_PN0N_  (.CLK(clknet_5_24__leaf_clk),
    .RESET_B(net320),
    .D(_0215_),
    .Q_N(_0049_),
    .Q(\Pong.datapath.NES_wire_Left[3] ));
 sg13g2_dfrbp_1 \Pong.datapath.NES_wire_Left[4]$_SDFFE_PN0N_  (.CLK(clknet_5_24__leaf_clk),
    .RESET_B(net321),
    .D(_0216_),
    .Q_N(_0050_),
    .Q(\Pong.datapath.NES_wire_Left[4] ));
 sg13g2_dfrbp_1 \Pong.datapath.NES_wire_Left[5]$_SDFFE_PN0N_  (.CLK(clknet_5_25__leaf_clk),
    .RESET_B(net322),
    .D(_0217_),
    .Q_N(_0051_),
    .Q(\Pong.datapath.NES_wire_Left[5] ));
 sg13g2_dfrbp_1 \Pong.datapath.NES_wire_Right[2]$_SDFFE_PN0N_  (.CLK(clknet_5_26__leaf_clk),
    .RESET_B(net323),
    .D(_0218_),
    .Q_N(_0052_),
    .Q(\Pong.datapath.NES_wire_Right[2] ));
 sg13g2_dfrbp_1 \Pong.datapath.NES_wire_Right[3]$_SDFFE_PN0N_  (.CLK(clknet_5_27__leaf_clk),
    .RESET_B(net324),
    .D(_0219_),
    .Q_N(_0053_),
    .Q(\Pong.datapath.NES_wire_Right[3] ));
 sg13g2_dfrbp_1 \Pong.datapath.NES_wire_Right[4]$_SDFFE_PN0N_  (.CLK(clknet_5_23__leaf_clk),
    .RESET_B(net325),
    .D(_0220_),
    .Q_N(_0054_),
    .Q(\Pong.datapath.NES_wire_Right[4] ));
 sg13g2_dfrbp_1 \Pong.datapath.NES_wire_Right[5]$_SDFFE_PN0N_  (.CLK(clknet_5_26__leaf_clk),
    .RESET_B(net326),
    .D(_0221_),
    .Q_N(_0055_),
    .Q(\Pong.datapath.NES_wire_Right[5] ));
 sg13g2_dfrbp_1 \Pong.datapath.ballFunction.ball_center_x_proc[0]$_SDFFE_PN0P_  (.CLK(net82),
    .RESET_B(net327),
    .D(_0222_),
    .Q_N(_0085_),
    .Q(\Pong.datapath.ballFunction.ball_center_x[0] ));
 sg13g2_dfrbp_1 \Pong.datapath.ballFunction.ball_center_x_proc[1]$_SDFFE_PN0P_  (.CLK(net82),
    .RESET_B(net328),
    .D(_0223_),
    .Q_N(_3091_),
    .Q(\Pong.datapath.ballFunction.ball_center_x[1] ));
 sg13g2_dfrbp_1 \Pong.datapath.ballFunction.ball_center_x_proc[2]$_SDFFE_PN0P_  (.CLK(net82),
    .RESET_B(net329),
    .D(_0224_),
    .Q_N(_0086_),
    .Q(\Pong.datapath.ballFunction.ball_center_x[2] ));
 sg13g2_dfrbp_1 \Pong.datapath.ballFunction.ball_center_x_proc[3]$_SDFFE_PN0P_  (.CLK(net82),
    .RESET_B(net330),
    .D(_0225_),
    .Q_N(_0080_),
    .Q(\Pong.datapath.ballFunction.ball_center_x[3] ));
 sg13g2_dfrbp_1 \Pong.datapath.ballFunction.ball_center_x_proc[4]$_SDFFE_PN0P_  (.CLK(net82),
    .RESET_B(net331),
    .D(_0226_),
    .Q_N(_0087_),
    .Q(\Pong.datapath.ballFunction.ball_center_x[4] ));
 sg13g2_dfrbp_1 \Pong.datapath.ballFunction.ball_center_x_proc[5]$_SDFFE_PN0P_  (.CLK(net82),
    .RESET_B(net332),
    .D(_0227_),
    .Q_N(_0088_),
    .Q(\Pong.datapath.ballFunction.ball_center_x[5] ));
 sg13g2_dfrbp_1 \Pong.datapath.ballFunction.ball_center_x_proc[6]$_SDFFE_PN1P_  (.CLK(net80),
    .RESET_B(net333),
    .D(_0228_),
    .Q_N(_0089_),
    .Q(\Pong.datapath.ballFunction.ball_center_x[6] ));
 sg13g2_dfrbp_1 \Pong.datapath.ballFunction.ball_center_x_proc[7]$_SDFFE_PN0P_  (.CLK(net80),
    .RESET_B(net334),
    .D(_0229_),
    .Q_N(_0079_),
    .Q(\Pong.datapath.ballFunction.ball_center_x[7] ));
 sg13g2_dfrbp_1 \Pong.datapath.ballFunction.ball_center_x_proc[8]$_SDFFE_PN1P_  (.CLK(net80),
    .RESET_B(net335),
    .D(_0230_),
    .Q_N(_0090_),
    .Q(\Pong.datapath.ballFunction.ball_center_x[8] ));
 sg13g2_dfrbp_1 \Pong.datapath.ballFunction.ball_center_x_proc[9]$_SDFFE_PN0P_  (.CLK(net80),
    .RESET_B(net336),
    .D(_0231_),
    .Q_N(_0091_),
    .Q(\Pong.datapath.ballFunction.ball_center_x[9] ));
 sg13g2_dfrbp_1 \Pong.datapath.ballFunction.ball_center_y_proc[0]$_SDFFE_PN0P_  (.CLK(net81),
    .RESET_B(net337),
    .D(_0232_),
    .Q_N(_0092_),
    .Q(\Pong.datapath.ballFunction.ball_center_y[0] ));
 sg13g2_dfrbp_1 \Pong.datapath.ballFunction.ball_center_y_proc[1]$_SDFFE_PN0P_  (.CLK(net81),
    .RESET_B(net338),
    .D(_0233_),
    .Q_N(_0113_),
    .Q(\Pong.datapath.ballFunction.ball_center_y[1] ));
 sg13g2_dfrbp_1 \Pong.datapath.ballFunction.ball_center_y_proc[2]$_SDFFE_PN1P_  (.CLK(net81),
    .RESET_B(net339),
    .D(_0234_),
    .Q_N(_0069_),
    .Q(\Pong.datapath.ballFunction.ball_center_y[2] ));
 sg13g2_dfrbp_1 \Pong.datapath.ballFunction.ball_center_y_proc[3]$_SDFFE_PN1P_  (.CLK(net81),
    .RESET_B(net340),
    .D(_0235_),
    .Q_N(_0112_),
    .Q(\Pong.datapath.ballFunction.ball_center_y[3] ));
 sg13g2_dfrbp_1 \Pong.datapath.ballFunction.ball_center_y_proc[4]$_SDFFE_PN1P_  (.CLK(net81),
    .RESET_B(net341),
    .D(_0236_),
    .Q_N(_0066_),
    .Q(\Pong.datapath.ballFunction.ball_center_y[4] ));
 sg13g2_dfrbp_1 \Pong.datapath.ballFunction.ball_center_y_proc[5]$_SDFFE_PN0P_  (.CLK(net80),
    .RESET_B(net342),
    .D(_0237_),
    .Q_N(_0065_),
    .Q(\Pong.datapath.ballFunction.ball_center_y[5] ));
 sg13g2_dfrbp_1 \Pong.datapath.ballFunction.ball_center_y_proc[6]$_SDFFE_PN1P_  (.CLK(net81),
    .RESET_B(net343),
    .D(_0238_),
    .Q_N(_0064_),
    .Q(\Pong.datapath.ballFunction.ball_center_y[6] ));
 sg13g2_dfrbp_1 \Pong.datapath.ballFunction.ball_center_y_proc[7]$_SDFFE_PN1P_  (.CLK(net80),
    .RESET_B(net344),
    .D(_0239_),
    .Q_N(_0070_),
    .Q(\Pong.datapath.ballFunction.ball_center_y[7] ));
 sg13g2_dfrbp_1 \Pong.datapath.ballFunction.ball_center_y_proc[8]$_SDFFE_PN0P_  (.CLK(net80),
    .RESET_B(net345),
    .D(_0240_),
    .Q_N(_0060_),
    .Q(\Pong.datapath.ballFunction.ball_center_y[8] ));
 sg13g2_dfrbp_1 \Pong.datapath.ballFunction.ball_center_y_proc[9]$_SDFFE_PN0P_  (.CLK(net80),
    .RESET_B(net346),
    .D(_0241_),
    .Q_N(_0059_),
    .Q(\Pong.datapath.ballFunction.ball_center_y[9] ));
 sg13g2_dfrbp_1 \Pong.datapath.ballReset$_SDFF_PN0_  (.CLK(clknet_5_31__leaf_clk),
    .RESET_B(net347),
    .D(_0242_),
    .Q_N(_3090_),
    .Q(\Pong.datapath.ballFunction.reset_n ));
 sg13g2_dfrbp_1 \Pong.datapath.leftPaddle[0]$_SDFF_PN0_  (.CLK(clknet_5_30__leaf_clk),
    .RESET_B(net348),
    .D(_0243_),
    .Q_N(_0083_),
    .Q(\Pong.datapath.leftPaddle[0] ));
 sg13g2_dfrbp_1 \Pong.datapath.leftPaddle[1]$_SDFF_PN0_  (.CLK(clknet_5_31__leaf_clk),
    .RESET_B(net349),
    .D(_0244_),
    .Q_N(_0076_),
    .Q(\Pong.datapath.leftPaddle[1] ));
 sg13g2_dfrbp_1 \Pong.datapath.leftPaddle[2]$_SDFF_PN1_  (.CLK(clknet_5_30__leaf_clk),
    .RESET_B(net350),
    .D(_0245_),
    .Q_N(_0084_),
    .Q(\Pong.datapath.leftPaddle[2] ));
 sg13g2_dfrbp_1 \Pong.datapath.leftPaddle[3]$_SDFF_PN1_  (.CLK(clknet_5_30__leaf_clk),
    .RESET_B(net351),
    .D(_0246_),
    .Q_N(_0078_),
    .Q(\Pong.datapath.leftPaddle[3] ));
 sg13g2_dfrbp_1 \Pong.datapath.leftPaddle[4]$_SDFF_PN1_  (.CLK(clknet_5_31__leaf_clk),
    .RESET_B(net352),
    .D(_0247_),
    .Q_N(_0077_),
    .Q(\Pong.datapath.leftPaddle[4] ));
 sg13g2_dfrbp_1 \Pong.datapath.leftPaddle[5]$_SDFF_PN0_  (.CLK(clknet_5_31__leaf_clk),
    .RESET_B(net353),
    .D(_0248_),
    .Q_N(_0071_),
    .Q(\Pong.datapath.leftPaddle[5] ));
 sg13g2_dfrbp_1 \Pong.datapath.leftPaddle[6]$_SDFF_PN1_  (.CLK(clknet_5_30__leaf_clk),
    .RESET_B(net354),
    .D(_0249_),
    .Q_N(_0075_),
    .Q(\Pong.datapath.leftPaddle[6] ));
 sg13g2_dfrbp_1 \Pong.datapath.leftPaddle[7]$_SDFF_PN1_  (.CLK(clknet_5_28__leaf_clk),
    .RESET_B(net355),
    .D(_0250_),
    .Q_N(_0074_),
    .Q(\Pong.datapath.leftPaddle[7] ));
 sg13g2_dfrbp_1 \Pong.datapath.leftPaddle[8]$_SDFF_PN0_  (.CLK(clknet_5_31__leaf_clk),
    .RESET_B(net356),
    .D(_0251_),
    .Q_N(_0073_),
    .Q(\Pong.datapath.leftPaddle[8] ));
 sg13g2_dfrbp_1 \Pong.datapath.leftPaddle[9]$_SDFF_PN0_  (.CLK(clknet_5_30__leaf_clk),
    .RESET_B(net357),
    .D(_0252_),
    .Q_N(_0072_),
    .Q(\Pong.datapath.leftPaddle[9] ));
 sg13g2_dfrbp_1 \Pong.datapath.old_NES_Left[2]$_SDFF_PN0_  (.CLK(clknet_5_25__leaf_clk),
    .RESET_B(net358),
    .D(_0253_),
    .Q_N(_3089_),
    .Q(\Pong.datapath.old_NES_Left[2] ));
 sg13g2_dfrbp_1 \Pong.datapath.old_NES_Left[3]$_SDFF_PN0_  (.CLK(clknet_5_24__leaf_clk),
    .RESET_B(net359),
    .D(_0254_),
    .Q_N(_3088_),
    .Q(\Pong.datapath.old_NES_Left[3] ));
 sg13g2_dfrbp_1 \Pong.datapath.old_NES_Left[4]$_SDFF_PN0_  (.CLK(clknet_5_24__leaf_clk),
    .RESET_B(net360),
    .D(_0255_),
    .Q_N(_3087_),
    .Q(\Pong.datapath.old_NES_Left[4] ));
 sg13g2_dfrbp_1 \Pong.datapath.old_NES_Left[5]$_SDFF_PN0_  (.CLK(clknet_5_26__leaf_clk),
    .RESET_B(net361),
    .D(_0256_),
    .Q_N(_3086_),
    .Q(\Pong.datapath.old_NES_Left[5] ));
 sg13g2_dfrbp_1 \Pong.datapath.old_NES_Right[2]$_SDFF_PN0_  (.CLK(clknet_5_27__leaf_clk),
    .RESET_B(net362),
    .D(_0257_),
    .Q_N(_3085_),
    .Q(\Pong.datapath.old_NES_Right[2] ));
 sg13g2_dfrbp_1 \Pong.datapath.old_NES_Right[3]$_SDFF_PN0_  (.CLK(clknet_5_27__leaf_clk),
    .RESET_B(net363),
    .D(_0258_),
    .Q_N(_3084_),
    .Q(\Pong.datapath.old_NES_Right[3] ));
 sg13g2_dfrbp_1 \Pong.datapath.old_NES_Right[4]$_SDFF_PN0_  (.CLK(clknet_5_27__leaf_clk),
    .RESET_B(net364),
    .D(_0259_),
    .Q_N(_3083_),
    .Q(\Pong.datapath.old_NES_Right[4] ));
 sg13g2_dfrbp_1 \Pong.datapath.old_NES_Right[5]$_SDFF_PN0_  (.CLK(clknet_5_26__leaf_clk),
    .RESET_B(net365),
    .D(_0260_),
    .Q_N(_3082_),
    .Q(\Pong.datapath.old_NES_Right[5] ));
 sg13g2_dfrbp_1 \Pong.datapath.rightPaddle[0]$_SDFF_PN0_  (.CLK(clknet_5_31__leaf_clk),
    .RESET_B(net366),
    .D(_0261_),
    .Q_N(_3081_),
    .Q(\Pong.datapath.rightPaddle[0] ));
 sg13g2_dfrbp_1 \Pong.datapath.rightPaddle[1]$_SDFF_PN0_  (.CLK(clknet_5_29__leaf_clk),
    .RESET_B(net367),
    .D(_0262_),
    .Q_N(_3080_),
    .Q(\Pong.datapath.rightPaddle[1] ));
 sg13g2_dfrbp_1 \Pong.datapath.rightPaddle[2]$_SDFF_PN1_  (.CLK(clknet_5_28__leaf_clk),
    .RESET_B(net368),
    .D(_0263_),
    .Q_N(_0082_),
    .Q(\Pong.datapath.rightPaddle[2] ));
 sg13g2_dfrbp_1 \Pong.datapath.rightPaddle[3]$_SDFF_PN1_  (.CLK(clknet_5_29__leaf_clk),
    .RESET_B(net369),
    .D(_0264_),
    .Q_N(_0068_),
    .Q(\Pong.datapath.rightPaddle[3] ));
 sg13g2_dfrbp_1 \Pong.datapath.rightPaddle[4]$_SDFF_PN1_  (.CLK(clknet_5_29__leaf_clk),
    .RESET_B(net370),
    .D(_0265_),
    .Q_N(_0067_),
    .Q(\Pong.datapath.rightPaddle[4] ));
 sg13g2_dfrbp_1 \Pong.datapath.rightPaddle[5]$_SDFF_PN0_  (.CLK(clknet_5_28__leaf_clk),
    .RESET_B(net371),
    .D(_0266_),
    .Q_N(_0057_),
    .Q(\Pong.datapath.rightPaddle[5] ));
 sg13g2_dfrbp_1 \Pong.datapath.rightPaddle[6]$_SDFF_PN1_  (.CLK(clknet_5_29__leaf_clk),
    .RESET_B(net372),
    .D(_0267_),
    .Q_N(_0063_),
    .Q(\Pong.datapath.rightPaddle[6] ));
 sg13g2_dfrbp_1 \Pong.datapath.rightPaddle[7]$_SDFF_PN1_  (.CLK(clknet_5_28__leaf_clk),
    .RESET_B(net373),
    .D(_0268_),
    .Q_N(_0062_),
    .Q(\Pong.datapath.rightPaddle[7] ));
 sg13g2_dfrbp_1 \Pong.datapath.rightPaddle[8]$_SDFF_PN0_  (.CLK(clknet_5_28__leaf_clk),
    .RESET_B(net374),
    .D(_0269_),
    .Q_N(_0061_),
    .Q(\Pong.datapath.rightPaddle[8] ));
 sg13g2_dfrbp_1 \Pong.datapath.rightPaddle[9]$_SDFF_PN0_  (.CLK(clknet_5_28__leaf_clk),
    .RESET_B(net375),
    .D(_0270_),
    .Q_N(_0058_),
    .Q(\Pong.datapath.rightPaddle[9] ));
 sg13g2_dfrbp_1 \Pong.datapath.scoreLeftProc[0]$_SDFF_PN0_  (.CLK(clknet_5_15__leaf_clk),
    .RESET_B(net376),
    .D(_0271_),
    .Q_N(_3079_),
    .Q(\Pong.datapath.scoreLeft[0] ));
 sg13g2_dfrbp_1 \Pong.datapath.scoreLeftProc[1]$_SDFF_PN0_  (.CLK(clknet_5_7__leaf_clk),
    .RESET_B(net377),
    .D(_0272_),
    .Q_N(_3078_),
    .Q(\Pong.datapath.scoreLeft[1] ));
 sg13g2_dfrbp_1 \Pong.datapath.scoreLeftProc[2]$_SDFF_PN0_  (.CLK(clknet_5_25__leaf_clk),
    .RESET_B(net378),
    .D(_0273_),
    .Q_N(_3077_),
    .Q(\Pong.datapath.scoreLeft[2] ));
 sg13g2_dfrbp_1 \Pong.datapath.scoreLeftProc[3]$_SDFF_PN0_  (.CLK(clknet_5_24__leaf_clk),
    .RESET_B(net379),
    .D(_0274_),
    .Q_N(_3076_),
    .Q(\Pong.datapath.scoreLeft[3] ));
 sg13g2_dfrbp_1 \Pong.datapath.scoreRightProc[0]$_SDFF_PN0_  (.CLK(clknet_5_6__leaf_clk),
    .RESET_B(net380),
    .D(_0275_),
    .Q_N(_3075_),
    .Q(\Pong.datapath.scoreRight[0] ));
 sg13g2_dfrbp_1 \Pong.datapath.scoreRightProc[1]$_SDFF_PN0_  (.CLK(clknet_5_6__leaf_clk),
    .RESET_B(net381),
    .D(_0276_),
    .Q_N(_3074_),
    .Q(\Pong.datapath.scoreRight[1] ));
 sg13g2_dfrbp_1 \Pong.datapath.scoreRightProc[2]$_SDFF_PN0_  (.CLK(clknet_5_6__leaf_clk),
    .RESET_B(net382),
    .D(_0277_),
    .Q_N(_3073_),
    .Q(\Pong.datapath.scoreRight[2] ));
 sg13g2_dfrbp_1 \Pong.datapath.scoreRightProc[3]$_SDFF_PN0_  (.CLK(clknet_5_7__leaf_clk),
    .RESET_B(net383),
    .D(_0278_),
    .Q_N(_3072_),
    .Q(\Pong.datapath.scoreRight[3] ));
 sg13g2_dfrbp_1 \Pong.datapath.score_flag$_SDFF_PN1_  (.CLK(clknet_5_25__leaf_clk),
    .RESET_B(net384),
    .D(_0279_),
    .Q_N(_3191_),
    .Q(\Pong.datapath.score_flag ));
 sg13g2_dfrbp_1 \Pong.datapath.sw_ballMovement_reg[0]$_DFF_P_  (.CLK(clknet_5_10__leaf_clk),
    .RESET_B(net385),
    .D(_0043_),
    .Q_N(_0111_),
    .Q(\Pong.datapath.sw_ballMovement_reg[0] ));
 sg13g2_dfrbp_1 \Pong.datapath.sw_ballMovement_reg[2]$_DFF_P_  (.CLK(clknet_5_11__leaf_clk),
    .RESET_B(net386),
    .D(_0044_),
    .Q_N(_3192_),
    .Q(\Pong.datapath.sw_ballMovement_reg[2] ));
 sg13g2_dfrbp_1 \Pong.datapath.sw_ballMovement_reg[3]$_DFF_P_  (.CLK(clknet_5_11__leaf_clk),
    .RESET_B(net387),
    .D(_0045_),
    .Q_N(_3193_),
    .Q(\Pong.datapath.sw_ballMovement_reg[3] ));
 sg13g2_dfrbp_1 \Pong.datapath.sw_ballMovement_reg[4]$_DFF_P_  (.CLK(clknet_5_11__leaf_clk),
    .RESET_B(net388),
    .D(_0046_),
    .Q_N(_3194_),
    .Q(\Pong.datapath.sw_ballMovement_reg[4] ));
 sg13g2_dfrbp_1 \Pong.datapath.sw_ballMovement_reg[5]$_DFF_P_  (.CLK(clknet_5_11__leaf_clk),
    .RESET_B(net389),
    .D(_0047_),
    .Q_N(_3071_),
    .Q(\Pong.datapath.sw_ballMovement_reg[5] ));
 sg13g2_dfrbp_1 \Pong.datapath.vga.Column_Counter.processQ[0]$_SDFFE_PN0P_  (.CLK(clknet_5_10__leaf_clk),
    .RESET_B(net390),
    .D(_0280_),
    .Q_N(_3070_),
    .Q(\Pong.datapath.vga.Column_Counter.Q[0] ));
 sg13g2_dfrbp_1 \Pong.datapath.vga.Column_Counter.processQ[1]$_SDFFE_PN0P_  (.CLK(clknet_5_8__leaf_clk),
    .RESET_B(net391),
    .D(_0281_),
    .Q_N(_0109_),
    .Q(\Pong.datapath.vga.Column_Counter.Q[1] ));
 sg13g2_dfrbp_1 \Pong.datapath.vga.Column_Counter.processQ[2]$_SDFFE_PN0P_  (.CLK(clknet_5_12__leaf_clk),
    .RESET_B(net392),
    .D(_0282_),
    .Q_N(_0101_),
    .Q(\Pong.datapath.vga.Column_Counter.Q[2] ));
 sg13g2_dfrbp_1 \Pong.datapath.vga.Column_Counter.processQ[3]$_SDFFE_PN0P_  (.CLK(clknet_5_14__leaf_clk),
    .RESET_B(net393),
    .D(_0283_),
    .Q_N(_0102_),
    .Q(\Pong.datapath.vga.Column_Counter.Q[3] ));
 sg13g2_dfrbp_1 \Pong.datapath.vga.Column_Counter.processQ[4]$_SDFFE_PN0P_  (.CLK(clknet_5_6__leaf_clk),
    .RESET_B(net394),
    .D(_0284_),
    .Q_N(_0103_),
    .Q(\Pong.datapath.vga.Column_Counter.Q[4] ));
 sg13g2_dfrbp_1 \Pong.datapath.vga.Column_Counter.processQ[5]$_SDFFE_PN0P_  (.CLK(clknet_5_13__leaf_clk),
    .RESET_B(net395),
    .D(_0285_),
    .Q_N(_0114_),
    .Q(\Pong.datapath.vga.Column_Counter.Q[5] ));
 sg13g2_dfrbp_1 \Pong.datapath.vga.Column_Counter.processQ[6]$_SDFFE_PN0P_  (.CLK(clknet_5_13__leaf_clk),
    .RESET_B(net396),
    .D(_0286_),
    .Q_N(_0104_),
    .Q(\Pong.datapath.vga.Column_Counter.Q[6] ));
 sg13g2_dfrbp_1 \Pong.datapath.vga.Column_Counter.processQ[7]$_SDFFE_PN0P_  (.CLK(clknet_5_12__leaf_clk),
    .RESET_B(net397),
    .D(_0287_),
    .Q_N(_0105_),
    .Q(\Pong.datapath.vga.Column_Counter.Q[7] ));
 sg13g2_dfrbp_1 \Pong.datapath.vga.Column_Counter.processQ[8]$_SDFFE_PN0P_  (.CLK(clknet_5_12__leaf_clk),
    .RESET_B(net398),
    .D(_0288_),
    .Q_N(_0106_),
    .Q(\Pong.datapath.vga.Column_Counter.Q[8] ));
 sg13g2_dfrbp_1 \Pong.datapath.vga.Column_Counter.processQ[9]$_SDFFE_PN0P_  (.CLK(clknet_5_12__leaf_clk),
    .RESET_B(net399),
    .D(_0289_),
    .Q_N(_0107_),
    .Q(\Pong.datapath.vga.Column_Counter.Q[9] ));
 sg13g2_dfrbp_1 \Pong.datapath.vga.Row_Counter.processQ[0]$_SDFFE_PN0P_  (.CLK(clknet_5_15__leaf_clk),
    .RESET_B(net400),
    .D(_0290_),
    .Q_N(_3069_),
    .Q(\Pong.datapath.vga.Row_Counter.Q[0] ));
 sg13g2_dfrbp_1 \Pong.datapath.vga.Row_Counter.processQ[1]$_SDFFE_PN0P_  (.CLK(clknet_5_15__leaf_clk),
    .RESET_B(net401),
    .D(_0291_),
    .Q_N(_0108_),
    .Q(\Pong.datapath.vga.Row_Counter.Q[1] ));
 sg13g2_dfrbp_1 \Pong.datapath.vga.Row_Counter.processQ[2]$_SDFFE_PN0P_  (.CLK(clknet_5_15__leaf_clk),
    .RESET_B(net402),
    .D(_0292_),
    .Q_N(_0093_),
    .Q(\Pong.datapath.vga.Row_Counter.Q[2] ));
 sg13g2_dfrbp_1 \Pong.datapath.vga.Row_Counter.processQ[3]$_SDFFE_PN0P_  (.CLK(clknet_5_15__leaf_clk),
    .RESET_B(net403),
    .D(_0293_),
    .Q_N(_0094_),
    .Q(\Pong.datapath.vga.Row_Counter.Q[3] ));
 sg13g2_dfrbp_1 \Pong.datapath.vga.Row_Counter.processQ[4]$_SDFFE_PN0P_  (.CLK(clknet_5_15__leaf_clk),
    .RESET_B(net404),
    .D(_0294_),
    .Q_N(_0095_),
    .Q(\Pong.datapath.vga.Row_Counter.Q[4] ));
 sg13g2_dfrbp_1 \Pong.datapath.vga.Row_Counter.processQ[5]$_SDFFE_PN0P_  (.CLK(clknet_5_14__leaf_clk),
    .RESET_B(net405),
    .D(_0295_),
    .Q_N(_0096_),
    .Q(\Pong.datapath.vga.Row_Counter.Q[5] ));
 sg13g2_dfrbp_1 \Pong.datapath.vga.Row_Counter.processQ[6]$_SDFFE_PN0P_  (.CLK(clknet_5_14__leaf_clk),
    .RESET_B(net406),
    .D(_0296_),
    .Q_N(_0097_),
    .Q(\Pong.datapath.vga.Row_Counter.Q[6] ));
 sg13g2_dfrbp_1 \Pong.datapath.vga.Row_Counter.processQ[7]$_SDFFE_PN0P_  (.CLK(clknet_5_14__leaf_clk),
    .RESET_B(net407),
    .D(_0297_),
    .Q_N(_0098_),
    .Q(\Pong.datapath.vga.Row_Counter.Q[7] ));
 sg13g2_dfrbp_1 \Pong.datapath.vga.Row_Counter.processQ[8]$_SDFFE_PN0P_  (.CLK(clknet_5_14__leaf_clk),
    .RESET_B(net408),
    .D(_0298_),
    .Q_N(_0099_),
    .Q(\Pong.datapath.vga.Row_Counter.Q[8] ));
 sg13g2_dfrbp_1 \Pong.datapath.vga.Row_Counter.processQ[9]$_SDFFE_PN0P_  (.CLK(clknet_5_14__leaf_clk),
    .RESET_B(net409),
    .D(_0299_),
    .Q_N(_0100_),
    .Q(\Pong.datapath.vga.Row_Counter.Q[9] ));
 sg13g2_buf_1 _3197_ (.A(\Pong.datapath.NES_counter_right.Q[3] ),
    .X(_2640_));
 sg13g2_buf_2 _3198_ (.A(\Pong.datapath.NES_counter_right.Q[4] ),
    .X(_2641_));
 sg13g2_buf_1 _3199_ (.A(\Pong.datapath.NES_counter_right.Q[5] ),
    .X(_2642_));
 sg13g2_nor2_1 _3200_ (.A(\Pong.datapath.NES_counter_right.Q[6] ),
    .B(_2642_),
    .Y(_2643_));
 sg13g2_buf_1 _3201_ (.A(\Pong.datapath.NES_counter_right.Q[1] ),
    .X(_2644_));
 sg13g2_buf_1 _3202_ (.A(\Pong.datapath.NES_counter_right.Q[0] ),
    .X(_2645_));
 sg13g2_inv_1 _3203_ (.Y(_2646_),
    .A(\Pong.datapath.NES_counter_right.Q[7] ));
 sg13g2_nor4_1 _3204_ (.A(_2644_),
    .B(_2645_),
    .C(\Pong.datapath.NES_counter_right.Q[2] ),
    .D(_2646_),
    .Y(_2647_));
 sg13g2_nand4_1 _3205_ (.B(_2641_),
    .C(_2643_),
    .A(_2640_),
    .Y(_2648_),
    .D(_2647_));
 sg13g2_buf_1 _3206_ (.A(_2648_),
    .X(_2649_));
 sg13g2_inv_1 _3207_ (.Y(_2650_),
    .A(_2649_));
 sg13g2_buf_1 _3208_ (.A(net93),
    .X(_2651_));
 sg13g2_nand2_1 _3209_ (.Y(_2652_),
    .A(\Pong.control_unit.NES_Controller_Right.state_NESController[10] ),
    .B(net85));
 sg13g2_buf_1 _3210_ (.A(_2649_),
    .X(_2653_));
 sg13g2_buf_1 _3211_ (.A(net92),
    .X(_2654_));
 sg13g2_nand2_1 _3212_ (.Y(_2655_),
    .A(\Pong.control_unit.NES_Controller_Right.state_NESController[5] ),
    .B(net84));
 sg13g2_buf_2 _3213_ (.A(rst_n),
    .X(_2656_));
 sg13g2_inv_1 _3214_ (.Y(_2657_),
    .A(_2656_));
 sg13g2_buf_1 _3215_ (.A(_2657_),
    .X(_2658_));
 sg13g2_a21oi_1 _3216_ (.A1(_2652_),
    .A2(_2655_),
    .Y(_0033_),
    .B1(net158));
 sg13g2_nand2_1 _3217_ (.Y(_2659_),
    .A(\Pong.control_unit.NES_Controller_Right.state_NESController[11] ),
    .B(net85));
 sg13g2_nand2_1 _3218_ (.Y(_2660_),
    .A(\Pong.control_unit.NES_Controller_Right.state_NESController[6] ),
    .B(net84));
 sg13g2_a21oi_1 _3219_ (.A1(_2659_),
    .A2(_2660_),
    .Y(_0034_),
    .B1(net158));
 sg13g2_nand2_1 _3220_ (.Y(_2661_),
    .A(\Pong.control_unit.NES_Controller_Right.state_NESController[12] ),
    .B(net85));
 sg13g2_nand2_1 _3221_ (.Y(_2662_),
    .A(\Pong.control_unit.NES_Controller_Right.state_NESController[7] ),
    .B(net84));
 sg13g2_a21oi_1 _3222_ (.A1(_2661_),
    .A2(_2662_),
    .Y(_0035_),
    .B1(net158));
 sg13g2_buf_1 _3223_ (.A(_2657_),
    .X(_2663_));
 sg13g2_buf_1 _3224_ (.A(net157),
    .X(_2664_));
 sg13g2_buf_1 _3225_ (.A(\Pong.control_unit.NES_Controller_Right.state_NESController[8] ),
    .X(_2665_));
 sg13g2_buf_1 _3226_ (.A(\Pong.control_unit.NES_Controller_Right.state_NESController[13] ),
    .X(_2666_));
 sg13g2_inv_1 _3227_ (.Y(_2667_),
    .A(_2666_));
 sg13g2_nor2_1 _3228_ (.A(_2667_),
    .B(net92),
    .Y(_2668_));
 sg13g2_a21oi_1 _3229_ (.A1(_2665_),
    .A2(net84),
    .Y(_2669_),
    .B1(_2668_));
 sg13g2_nor2_1 _3230_ (.A(_2664_),
    .B(_2669_),
    .Y(_0036_));
 sg13g2_nand2_1 _3231_ (.Y(_2670_),
    .A(\Pong.control_unit.NES_Controller_Right.state_NESController[14] ),
    .B(net85));
 sg13g2_buf_1 _3232_ (.A(\Pong.control_unit.NES_Controller_Right.state_NESController[9] ),
    .X(_2671_));
 sg13g2_nand2_1 _3233_ (.Y(_2672_),
    .A(_2671_),
    .B(net84));
 sg13g2_a21oi_1 _3234_ (.A1(_2670_),
    .A2(_2672_),
    .Y(_0037_),
    .B1(_2658_));
 sg13g2_nand2_1 _3235_ (.Y(_2673_),
    .A(\Pong.control_unit.NES_Controller_Right.state_NESController[10] ),
    .B(_2654_));
 sg13g2_buf_2 _3236_ (.A(\Pong.datapath.NES_delay_counter_right.Q[6] ),
    .X(_2674_));
 sg13g2_buf_8 _3237_ (.A(\Pong.datapath.NES_delay_counter_right.Q[0] ),
    .X(_2675_));
 sg13g2_and3_1 _3238_ (.X(_2676_),
    .A(\Pong.datapath.NES_delay_counter_right.Q[2] ),
    .B(\Pong.datapath.NES_delay_counter_right.Q[1] ),
    .C(_2675_));
 sg13g2_buf_8 _3239_ (.A(_2676_),
    .X(_2677_));
 sg13g2_buf_8 _3240_ (.A(\Pong.datapath.NES_delay_counter_right.Q[3] ),
    .X(_2678_));
 sg13g2_and3_1 _3241_ (.X(_2679_),
    .A(\Pong.datapath.NES_delay_counter_right.Q[4] ),
    .B(\Pong.datapath.NES_delay_counter_right.Q[5] ),
    .C(_2678_));
 sg13g2_buf_1 _3242_ (.A(_2679_),
    .X(_2680_));
 sg13g2_nand4_1 _3243_ (.B(_2674_),
    .C(_2677_),
    .A(\Pong.datapath.NES_delay_counter_right.Q[7] ),
    .Y(_2681_),
    .D(_2680_));
 sg13g2_buf_2 _3244_ (.A(_2681_),
    .X(_2682_));
 sg13g2_inv_1 _3245_ (.Y(_2683_),
    .A(\Pong.datapath.NES_delay_counter_right.Q[8] ));
 sg13g2_nand2b_1 _3246_ (.Y(_2684_),
    .B(_2683_),
    .A_N(_2682_));
 sg13g2_buf_8 _3247_ (.A(\Pong.datapath.NES_delay_counter_right.Q[17] ),
    .X(_2685_));
 sg13g2_nand2b_1 _3248_ (.Y(_2686_),
    .B(_2685_),
    .A_N(_0110_));
 sg13g2_buf_1 _3249_ (.A(\Pong.datapath.NES_delay_counter_right.Q[12] ),
    .X(_2687_));
 sg13g2_buf_1 _3250_ (.A(\Pong.datapath.NES_delay_counter_right.Q[11] ),
    .X(_2688_));
 sg13g2_or2_1 _3251_ (.X(_2689_),
    .B(_2688_),
    .A(_2687_));
 sg13g2_buf_2 _3252_ (.A(\Pong.datapath.NES_delay_counter_right.Q[14] ),
    .X(_2690_));
 sg13g2_buf_2 _3253_ (.A(\Pong.datapath.NES_delay_counter_right.Q[13] ),
    .X(_2691_));
 sg13g2_nor2_1 _3254_ (.A(\Pong.datapath.NES_delay_counter_right.Q[15] ),
    .B(\Pong.datapath.NES_delay_counter_right.Q[16] ),
    .Y(_2692_));
 sg13g2_buf_1 _3255_ (.A(\Pong.datapath.NES_delay_counter_right.Q[9] ),
    .X(_2693_));
 sg13g2_and2_1 _3256_ (.A(\Pong.datapath.NES_delay_counter_right.Q[10] ),
    .B(_2693_),
    .X(_2694_));
 sg13g2_nand4_1 _3257_ (.B(_2691_),
    .C(_2692_),
    .A(_2690_),
    .Y(_2695_),
    .D(_2694_));
 sg13g2_nor4_1 _3258_ (.A(_2684_),
    .B(_2686_),
    .C(_2689_),
    .D(_2695_),
    .Y(_2696_));
 sg13g2_nand2_1 _3259_ (.Y(_2697_),
    .A(\Pong.control_unit.NES_Controller_Right.state_NESController[0] ),
    .B(_2696_));
 sg13g2_buf_1 _3260_ (.A(_2697_),
    .X(_2698_));
 sg13g2_a21oi_1 _3261_ (.A1(_2673_),
    .A2(_2698_),
    .Y(_0020_),
    .B1(_2658_));
 sg13g2_nand2_1 _3262_ (.Y(_2699_),
    .A(\Pong.control_unit.NES_Controller_Right.state_NESController[1] ),
    .B(net85));
 sg13g2_nand2_1 _3263_ (.Y(_2700_),
    .A(\Pong.control_unit.NES_Controller_Right.state_NESController[11] ),
    .B(net84));
 sg13g2_buf_1 _3264_ (.A(net157),
    .X(_2701_));
 sg13g2_a21oi_1 _3265_ (.A1(_2699_),
    .A2(_2700_),
    .Y(_0021_),
    .B1(net108));
 sg13g2_nand2_1 _3266_ (.Y(_2702_),
    .A(\Pong.control_unit.NES_Controller_Right.state_NESController[2] ),
    .B(net85));
 sg13g2_nand2_1 _3267_ (.Y(_2703_),
    .A(\Pong.control_unit.NES_Controller_Right.state_NESController[12] ),
    .B(net84));
 sg13g2_a21oi_1 _3268_ (.A1(_2702_),
    .A2(_2703_),
    .Y(_0022_),
    .B1(net108));
 sg13g2_buf_1 _3269_ (.A(\Pong.control_unit.NES_Controller_Right.state_NESController[3] ),
    .X(_2704_));
 sg13g2_nand2_1 _3270_ (.Y(_2705_),
    .A(_2704_),
    .B(net85));
 sg13g2_nand2_1 _3271_ (.Y(_2706_),
    .A(_2666_),
    .B(_2654_));
 sg13g2_a21oi_1 _3272_ (.A1(_2705_),
    .A2(_2706_),
    .Y(_0023_),
    .B1(net108));
 sg13g2_buf_1 _3273_ (.A(\Pong.control_unit.NES_Controller_Right.state_NESController[4] ),
    .X(_2707_));
 sg13g2_nand2_1 _3274_ (.Y(_2708_),
    .A(_2707_),
    .B(net85));
 sg13g2_nand2_1 _3275_ (.Y(_2709_),
    .A(\Pong.control_unit.NES_Controller_Right.state_NESController[14] ),
    .B(net84));
 sg13g2_a21oi_1 _3276_ (.A1(_2708_),
    .A2(_2709_),
    .Y(_0024_),
    .B1(net108));
 sg13g2_nand2_1 _3277_ (.Y(_2710_),
    .A(\Pong.control_unit.NES_Controller_Right.state_NESController[5] ),
    .B(_2651_));
 sg13g2_nand2_1 _3278_ (.Y(_2711_),
    .A(\Pong.control_unit.NES_Controller_Right.state_NESController[15] ),
    .B(net92));
 sg13g2_a21oi_1 _3279_ (.A1(_2710_),
    .A2(_2711_),
    .Y(_0025_),
    .B1(net108));
 sg13g2_nand2_1 _3280_ (.Y(_2712_),
    .A(\Pong.control_unit.NES_Controller_Right.state_NESController[7] ),
    .B(net93));
 sg13g2_buf_1 _3281_ (.A(\Pong.control_unit.NES_Controller_Right.state_NESController[16] ),
    .X(_2713_));
 sg13g2_nand2_1 _3282_ (.Y(_2714_),
    .A(_2713_),
    .B(net92));
 sg13g2_a21oi_1 _3283_ (.A1(_2712_),
    .A2(_2714_),
    .Y(_0026_),
    .B1(net108));
 sg13g2_nand2_1 _3284_ (.Y(_2715_),
    .A(_2665_),
    .B(net93));
 sg13g2_nand2_1 _3285_ (.Y(_2716_),
    .A(\Pong.control_unit.NES_Controller_Right.state_NESController[17] ),
    .B(_2653_));
 sg13g2_a21oi_1 _3286_ (.A1(_2715_),
    .A2(_2716_),
    .Y(_0027_),
    .B1(_2701_));
 sg13g2_buf_1 _3287_ (.A(_2656_),
    .X(_2717_));
 sg13g2_buf_1 _3288_ (.A(\Pong.datapath.sw_ballMovement_reg[4] ),
    .X(_2718_));
 sg13g2_inv_1 _3289_ (.Y(_2719_),
    .A(\Pong.datapath.sw_ballMovement_reg[2] ));
 sg13g2_buf_1 _3290_ (.A(\Pong.control_unit.state_ballMovement[3] ),
    .X(_2720_));
 sg13g2_inv_1 _3291_ (.Y(_2721_),
    .A(\Pong.datapath.sw_ballMovement_reg[0] ));
 sg13g2_a22oi_1 _3292_ (.Y(_2722_),
    .B1(net187),
    .B2(_2721_),
    .A2(\Pong.control_unit.state_ballMovement[4] ),
    .A1(_2719_));
 sg13g2_buf_1 _3293_ (.A(\Pong.datapath.sw_ballMovement_reg[3] ),
    .X(_2723_));
 sg13g2_buf_2 _3294_ (.A(\Pong.control_unit.state_ballMovement[2] ),
    .X(_2724_));
 sg13g2_buf_2 _3295_ (.A(\Pong.control_unit.state_ballMovement[0] ),
    .X(_2725_));
 sg13g2_a22oi_1 _3296_ (.Y(_2726_),
    .B1(_2721_),
    .B2(_2725_),
    .A2(_2724_),
    .A1(_2719_));
 sg13g2_or2_1 _3297_ (.X(_2727_),
    .B(_2726_),
    .A(_2723_));
 sg13g2_o21ai_1 _3298_ (.B1(_2727_),
    .Y(_2728_),
    .A1(_2718_),
    .A2(_2722_));
 sg13g2_and3_1 _3299_ (.X(_0039_),
    .A(net188),
    .B(\Pong.datapath.sw_ballMovement_reg[5] ),
    .C(_2728_));
 sg13g2_inv_1 _3300_ (.Y(_2729_),
    .A(_0111_));
 sg13g2_nor2_1 _3301_ (.A(\Pong.datapath.sw_ballMovement_reg[2] ),
    .B(\Pong.datapath.sw_ballMovement_reg[5] ),
    .Y(_2730_));
 sg13g2_a22oi_1 _3302_ (.Y(_2731_),
    .B1(_2730_),
    .B2(_2724_),
    .A2(_2729_),
    .A1(_2725_));
 sg13g2_nor2_1 _3303_ (.A(_2723_),
    .B(_2731_),
    .Y(_2732_));
 sg13g2_a21oi_1 _3304_ (.A1(_2718_),
    .A2(\Pong.control_unit.state_ballMovement[4] ),
    .Y(_2733_),
    .B1(_2732_));
 sg13g2_nor2_1 _3305_ (.A(net109),
    .B(_2733_),
    .Y(_0040_));
 sg13g2_nand2_1 _3306_ (.Y(_2734_),
    .A(_2721_),
    .B(_2725_));
 sg13g2_nor2_1 _3307_ (.A(\Pong.datapath.sw_ballMovement_reg[5] ),
    .B(_2734_),
    .Y(_2735_));
 sg13g2_a21oi_1 _3308_ (.A1(\Pong.datapath.sw_ballMovement_reg[2] ),
    .A2(_2724_),
    .Y(_2736_),
    .B1(_2735_));
 sg13g2_buf_1 _3309_ (.A(_2656_),
    .X(_2737_));
 sg13g2_inv_1 _3310_ (.Y(_2738_),
    .A(\Pong.control_unit.state_ballMovement[1] ));
 sg13g2_nand2_1 _3311_ (.Y(_2739_),
    .A(net186),
    .B(_2738_));
 sg13g2_a21oi_1 _3312_ (.A1(_2718_),
    .A2(net187),
    .Y(_2740_),
    .B1(_2739_));
 sg13g2_o21ai_1 _3313_ (.B1(_2740_),
    .Y(_0038_),
    .A1(_2723_),
    .A2(_2736_));
 sg13g2_inv_1 _3314_ (.Y(_2741_),
    .A(net187));
 sg13g2_nor3_1 _3315_ (.A(\Pong.datapath.sw_ballMovement_reg[5] ),
    .B(\Pong.datapath.sw_ballMovement_reg[0] ),
    .C(_2741_),
    .Y(_2742_));
 sg13g2_a21oi_1 _3316_ (.A1(\Pong.datapath.sw_ballMovement_reg[2] ),
    .A2(\Pong.control_unit.state_ballMovement[4] ),
    .Y(_2743_),
    .B1(_2742_));
 sg13g2_nor2_1 _3317_ (.A(_2718_),
    .B(_2743_),
    .Y(_2744_));
 sg13g2_a21oi_1 _3318_ (.A1(_2723_),
    .A2(_2725_),
    .Y(_2745_),
    .B1(_2744_));
 sg13g2_nor2_1 _3319_ (.A(net109),
    .B(_2745_),
    .Y(_0041_));
 sg13g2_a22oi_1 _3320_ (.Y(_2746_),
    .B1(_2730_),
    .B2(\Pong.control_unit.state_ballMovement[4] ),
    .A2(_2729_),
    .A1(net187));
 sg13g2_nor2_1 _3321_ (.A(_2718_),
    .B(_2746_),
    .Y(_2747_));
 sg13g2_a21oi_1 _3322_ (.A1(_2723_),
    .A2(_2724_),
    .Y(_2748_),
    .B1(_2747_));
 sg13g2_nor2_1 _3323_ (.A(net109),
    .B(_2748_),
    .Y(_0042_));
 sg13g2_buf_2 _3324_ (.A(\Pong.datapath.ballFunction.ball_center_y[5] ),
    .X(_2749_));
 sg13g2_buf_1 _3325_ (.A(_2749_),
    .X(_2750_));
 sg13g2_inv_1 _3326_ (.Y(_2751_),
    .A(net61));
 sg13g2_buf_1 _3327_ (.A(\Pong.datapath.ballFunction.ball_center_y[4] ),
    .X(_2752_));
 sg13g2_buf_1 _3328_ (.A(_2752_),
    .X(_2753_));
 sg13g2_buf_1 _3329_ (.A(net60),
    .X(_2754_));
 sg13g2_buf_2 _3330_ (.A(_0112_),
    .X(_2755_));
 sg13g2_inv_1 _3331_ (.Y(_2756_),
    .A(_2755_));
 sg13g2_buf_2 _3332_ (.A(_0113_),
    .X(_2757_));
 sg13g2_buf_1 _3333_ (.A(\Pong.datapath.ballFunction.ball_center_y[1] ),
    .X(_2758_));
 sg13g2_buf_1 _3334_ (.A(net74),
    .X(_2759_));
 sg13g2_buf_1 _3335_ (.A(\Pong.datapath.ballFunction.ball_center_y[0] ),
    .X(_2760_));
 sg13g2_buf_1 _3336_ (.A(_2760_),
    .X(_2761_));
 sg13g2_nor2b_1 _3337_ (.A(net59),
    .B_N(net58),
    .Y(_2762_));
 sg13g2_buf_1 _3338_ (.A(\Pong.datapath.ballFunction.ball_center_y[2] ),
    .X(_2763_));
 sg13g2_buf_1 _3339_ (.A(_2763_),
    .X(_2764_));
 sg13g2_buf_2 _3340_ (.A(\Pong.datapath.ballFunction.ball_center_y[3] ),
    .X(_2765_));
 sg13g2_buf_1 _3341_ (.A(_2765_),
    .X(_2766_));
 sg13g2_inv_2 _3342_ (.Y(_2767_),
    .A(net56));
 sg13g2_nor2_1 _3343_ (.A(net57),
    .B(_2767_),
    .Y(_2768_));
 sg13g2_o21ai_1 _3344_ (.B1(_2768_),
    .Y(_2769_),
    .A1(_2757_),
    .A2(_2762_));
 sg13g2_nand3_1 _3345_ (.B(_2756_),
    .C(_2769_),
    .A(net38),
    .Y(_2770_));
 sg13g2_buf_1 _3346_ (.A(\Pong.datapath.ballFunction.ball_center_y[7] ),
    .X(_2771_));
 sg13g2_buf_1 _3347_ (.A(\Pong.datapath.ballFunction.ball_center_y[6] ),
    .X(_2772_));
 sg13g2_buf_1 _3348_ (.A(\Pong.datapath.ballFunction.ball_center_y[8] ),
    .X(_2773_));
 sg13g2_buf_1 _3349_ (.A(\Pong.datapath.ballFunction.ball_center_y[9] ),
    .X(_2774_));
 sg13g2_nor4_2 _3350_ (.A(_2771_),
    .B(_2772_),
    .C(_2773_),
    .Y(_2775_),
    .D(net72));
 sg13g2_and3_1 _3351_ (.X(_0043_),
    .A(_2751_),
    .B(_2770_),
    .C(_2775_));
 sg13g2_nand2_1 _3352_ (.Y(_2776_),
    .A(_2671_),
    .B(net93));
 sg13g2_nand2_1 _3353_ (.Y(_2777_),
    .A(\Pong.control_unit.NES_Controller_Right.state_NESController[18] ),
    .B(net92));
 sg13g2_a21oi_1 _3354_ (.A1(_2776_),
    .A2(_2777_),
    .Y(_0028_),
    .B1(_2701_));
 sg13g2_and2_1 _3355_ (.A(\Pong.datapath.NES_counter_left.Q[3] ),
    .B(\Pong.datapath.NES_counter_left.Q[4] ),
    .X(_2778_));
 sg13g2_buf_1 _3356_ (.A(_2778_),
    .X(_2779_));
 sg13g2_nor2_1 _3357_ (.A(\Pong.datapath.NES_counter_left.Q[6] ),
    .B(\Pong.datapath.NES_counter_left.Q[5] ),
    .Y(_2780_));
 sg13g2_buf_1 _3358_ (.A(\Pong.datapath.NES_counter_left.Q[0] ),
    .X(_2781_));
 sg13g2_inv_1 _3359_ (.Y(_2782_),
    .A(\Pong.datapath.NES_counter_left.Q[7] ));
 sg13g2_nor4_1 _3360_ (.A(\Pong.datapath.NES_counter_left.Q[1] ),
    .B(_2781_),
    .C(\Pong.datapath.NES_counter_left.Q[2] ),
    .D(_2782_),
    .Y(_2783_));
 sg13g2_nand3_1 _3361_ (.B(_2780_),
    .C(_2783_),
    .A(_2779_),
    .Y(_2784_));
 sg13g2_buf_1 _3362_ (.A(_2784_),
    .X(_2785_));
 sg13g2_inv_1 _3363_ (.Y(_2786_),
    .A(_2785_));
 sg13g2_buf_1 _3364_ (.A(net91),
    .X(_2787_));
 sg13g2_nand2_1 _3365_ (.Y(_2788_),
    .A(\Pong.control_unit.NES_Controller_Left.state_NESController[16] ),
    .B(net83));
 sg13g2_buf_1 _3366_ (.A(_2785_),
    .X(_2789_));
 sg13g2_nand2_1 _3367_ (.Y(_2790_),
    .A(\Pong.control_unit.NES_Controller_Left.state_NESController[4] ),
    .B(net90));
 sg13g2_a21oi_1 _3368_ (.A1(_2788_),
    .A2(_2790_),
    .Y(_0013_),
    .B1(net108));
 sg13g2_nand2_1 _3369_ (.Y(_2791_),
    .A(\Pong.control_unit.NES_Controller_Left.state_NESController[1] ),
    .B(net83));
 sg13g2_buf_1 _3370_ (.A(\Pong.control_unit.NES_Controller_Left.state_NESController[11] ),
    .X(_2792_));
 sg13g2_nand2_1 _3371_ (.Y(_2793_),
    .A(_2792_),
    .B(net90));
 sg13g2_a21oi_1 _3372_ (.A1(_2791_),
    .A2(_2793_),
    .Y(_0002_),
    .B1(net108));
 sg13g2_nand2_1 _3373_ (.Y(_2794_),
    .A(\Pong.control_unit.NES_Controller_Left.state_NESController[10] ),
    .B(net83));
 sg13g2_nand2_1 _3374_ (.Y(_2795_),
    .A(\Pong.control_unit.NES_Controller_Left.state_NESController[5] ),
    .B(net90));
 sg13g2_buf_1 _3375_ (.A(net157),
    .X(_2796_));
 sg13g2_a21oi_1 _3376_ (.A1(_2794_),
    .A2(_2795_),
    .Y(_0014_),
    .B1(net107));
 sg13g2_buf_1 _3377_ (.A(\Pong.control_unit.NES_Controller_Left.state_NESController[8] ),
    .X(_2797_));
 sg13g2_buf_1 _3378_ (.A(\Pong.control_unit.NES_Controller_Left.state_NESController[13] ),
    .X(_2798_));
 sg13g2_inv_1 _3379_ (.Y(_2799_),
    .A(_2798_));
 sg13g2_buf_1 _3380_ (.A(_2785_),
    .X(_2800_));
 sg13g2_nor2_1 _3381_ (.A(_2799_),
    .B(net89),
    .Y(_2801_));
 sg13g2_a21oi_1 _3382_ (.A1(_2797_),
    .A2(_2789_),
    .Y(_2802_),
    .B1(_2801_));
 sg13g2_nor2_1 _3383_ (.A(_2664_),
    .B(_2802_),
    .Y(_0017_));
 sg13g2_nand2_1 _3384_ (.Y(_2803_),
    .A(\Pong.control_unit.NES_Controller_Left.state_NESController[12] ),
    .B(net83));
 sg13g2_nand2_1 _3385_ (.Y(_2804_),
    .A(\Pong.control_unit.NES_Controller_Left.state_NESController[7] ),
    .B(_2789_));
 sg13g2_a21oi_1 _3386_ (.A1(_2803_),
    .A2(_2804_),
    .Y(_0016_),
    .B1(net107));
 sg13g2_nand2_1 _3387_ (.Y(_2805_),
    .A(\Pong.control_unit.NES_Controller_Left.state_NESController[15] ),
    .B(_2787_));
 sg13g2_buf_1 _3388_ (.A(\Pong.control_unit.NES_Controller_Left.state_NESController[3] ),
    .X(_2806_));
 sg13g2_nand2_1 _3389_ (.Y(_2807_),
    .A(_2806_),
    .B(net90));
 sg13g2_a21oi_1 _3390_ (.A1(_2805_),
    .A2(_2807_),
    .Y(_0012_),
    .B1(net107));
 sg13g2_nand2_1 _3391_ (.Y(_2808_),
    .A(_2792_),
    .B(net83));
 sg13g2_nand2_1 _3392_ (.Y(_2809_),
    .A(\Pong.control_unit.NES_Controller_Left.state_NESController[6] ),
    .B(net90));
 sg13g2_a21oi_1 _3393_ (.A1(_2808_),
    .A2(_2809_),
    .Y(_0015_),
    .B1(net107));
 sg13g2_nand2_1 _3394_ (.Y(_2810_),
    .A(\Pong.control_unit.NES_Controller_Left.state_NESController[10] ),
    .B(net90));
 sg13g2_buf_2 _3395_ (.A(\Pong.control_unit.NES_Controller_Left.state_NESController[0] ),
    .X(_2811_));
 sg13g2_inv_1 _3396_ (.Y(_2812_),
    .A(\Pong.datapath.NES_delay_counter_left.Q[8] ));
 sg13g2_buf_1 _3397_ (.A(\Pong.datapath.NES_delay_counter_left.Q[0] ),
    .X(_2813_));
 sg13g2_and3_1 _3398_ (.X(_2814_),
    .A(\Pong.datapath.NES_delay_counter_left.Q[2] ),
    .B(\Pong.datapath.NES_delay_counter_left.Q[1] ),
    .C(_2813_));
 sg13g2_buf_2 _3399_ (.A(_2814_),
    .X(_2815_));
 sg13g2_buf_1 _3400_ (.A(\Pong.datapath.NES_delay_counter_left.Q[3] ),
    .X(_2816_));
 sg13g2_and3_1 _3401_ (.X(_2817_),
    .A(\Pong.datapath.NES_delay_counter_left.Q[5] ),
    .B(\Pong.datapath.NES_delay_counter_left.Q[4] ),
    .C(_2816_));
 sg13g2_buf_1 _3402_ (.A(_2817_),
    .X(_2818_));
 sg13g2_buf_1 _3403_ (.A(\Pong.datapath.NES_delay_counter_left.Q[6] ),
    .X(_2819_));
 sg13g2_and2_1 _3404_ (.A(\Pong.datapath.NES_delay_counter_left.Q[7] ),
    .B(_2819_),
    .X(_2820_));
 sg13g2_buf_1 _3405_ (.A(_2820_),
    .X(_2821_));
 sg13g2_nand4_1 _3406_ (.B(_2815_),
    .C(_2818_),
    .A(_2812_),
    .Y(_2822_),
    .D(_2821_));
 sg13g2_or2_1 _3407_ (.X(_2823_),
    .B(\Pong.datapath.NES_delay_counter_left.Q[11] ),
    .A(\Pong.datapath.NES_delay_counter_left.Q[12] ));
 sg13g2_buf_1 _3408_ (.A(_2823_),
    .X(_2824_));
 sg13g2_buf_1 _3409_ (.A(\Pong.datapath.NES_delay_counter_left.Q[10] ),
    .X(_2825_));
 sg13g2_buf_1 _3410_ (.A(\Pong.datapath.NES_delay_counter_left.Q[9] ),
    .X(_2826_));
 sg13g2_inv_1 _3411_ (.Y(_2827_),
    .A(\Pong.datapath.NES_delay_counter_left.Q[17] ));
 sg13g2_nor2_1 _3412_ (.A(_2827_),
    .B(_0117_),
    .Y(_2828_));
 sg13g2_nor2_1 _3413_ (.A(\Pong.datapath.NES_delay_counter_left.Q[15] ),
    .B(\Pong.datapath.NES_delay_counter_left.Q[16] ),
    .Y(_2829_));
 sg13g2_and2_1 _3414_ (.A(\Pong.datapath.NES_delay_counter_left.Q[14] ),
    .B(\Pong.datapath.NES_delay_counter_left.Q[13] ),
    .X(_2830_));
 sg13g2_and2_1 _3415_ (.A(_2829_),
    .B(_2830_),
    .X(_2831_));
 sg13g2_nand4_1 _3416_ (.B(_2826_),
    .C(_2828_),
    .A(_2825_),
    .Y(_2832_),
    .D(_2831_));
 sg13g2_nor3_1 _3417_ (.A(_2822_),
    .B(_2824_),
    .C(_2832_),
    .Y(_2833_));
 sg13g2_nand2_1 _3418_ (.Y(_2834_),
    .A(_2811_),
    .B(_2833_));
 sg13g2_buf_2 _3419_ (.A(_2834_),
    .X(_2835_));
 sg13g2_a21oi_1 _3420_ (.A1(_2810_),
    .A2(_2835_),
    .Y(_0001_),
    .B1(net107));
 sg13g2_inv_1 _3421_ (.Y(_2836_),
    .A(_2811_));
 sg13g2_a21oi_1 _3422_ (.A1(\Pong.control_unit.NES_Controller_Left.state_NESController[6] ),
    .A2(net91),
    .Y(_2837_),
    .B1(net157));
 sg13g2_o21ai_1 _3423_ (.B1(_2837_),
    .Y(_0000_),
    .A1(_2836_),
    .A2(_2833_));
 sg13g2_inv_1 _3424_ (.Y(_2838_),
    .A(\Pong.control_unit.NES_Controller_Left.state_NESController[14] ));
 sg13g2_nor2_1 _3425_ (.A(_2838_),
    .B(net89),
    .Y(_2839_));
 sg13g2_a21oi_1 _3426_ (.A1(\Pong.control_unit.NES_Controller_Left.state_NESController[9] ),
    .A2(net90),
    .Y(_2840_),
    .B1(_2839_));
 sg13g2_nor2_1 _3427_ (.A(net109),
    .B(_2840_),
    .Y(_0018_));
 sg13g2_buf_1 _3428_ (.A(\Pong.control_unit.NES_Controller_Left.state_NESController[18] ),
    .X(_2841_));
 sg13g2_nand2_1 _3429_ (.Y(_2842_),
    .A(_2841_),
    .B(net83));
 sg13g2_nand2_1 _3430_ (.Y(_2843_),
    .A(\Pong.control_unit.NES_Controller_Left.state_NESController[1] ),
    .B(net90));
 sg13g2_a21oi_1 _3431_ (.A1(_2842_),
    .A2(_2843_),
    .Y(_0010_),
    .B1(net107));
 sg13g2_buf_1 _3432_ (.A(\Pong.control_unit.NES_Controller_Left.state_NESController[17] ),
    .X(_2844_));
 sg13g2_nand2_1 _3433_ (.Y(_2845_),
    .A(_2844_),
    .B(_2787_));
 sg13g2_nand2_1 _3434_ (.Y(_2846_),
    .A(\Pong.control_unit.NES_Controller_Left.state_NESController[2] ),
    .B(net89));
 sg13g2_a21oi_1 _3435_ (.A1(_2845_),
    .A2(_2846_),
    .Y(_0011_),
    .B1(net107));
 sg13g2_nand2_1 _3436_ (.Y(_2847_),
    .A(_2713_),
    .B(net93));
 sg13g2_nand2_1 _3437_ (.Y(_2848_),
    .A(_2707_),
    .B(net92));
 sg13g2_a21oi_1 _3438_ (.A1(_2847_),
    .A2(_2848_),
    .Y(_0032_),
    .B1(net107));
 sg13g2_nand2_1 _3439_ (.Y(_2849_),
    .A(\Pong.control_unit.NES_Controller_Right.state_NESController[15] ),
    .B(_2650_));
 sg13g2_nand2_1 _3440_ (.Y(_2850_),
    .A(_2704_),
    .B(_2653_));
 sg13g2_a21oi_1 _3441_ (.A1(_2849_),
    .A2(_2850_),
    .Y(_0031_),
    .B1(_2796_));
 sg13g2_nand2_1 _3442_ (.Y(_2851_),
    .A(\Pong.control_unit.NES_Controller_Right.state_NESController[17] ),
    .B(_2650_));
 sg13g2_nand2_1 _3443_ (.Y(_2852_),
    .A(\Pong.control_unit.NES_Controller_Right.state_NESController[2] ),
    .B(net92));
 sg13g2_a21oi_1 _3444_ (.A1(_2851_),
    .A2(_2852_),
    .Y(_0030_),
    .B1(_2796_));
 sg13g2_nand2_1 _3445_ (.Y(_2853_),
    .A(\Pong.control_unit.NES_Controller_Right.state_NESController[18] ),
    .B(net93));
 sg13g2_nand2_1 _3446_ (.Y(_2854_),
    .A(\Pong.control_unit.NES_Controller_Right.state_NESController[1] ),
    .B(net92));
 sg13g2_buf_1 _3447_ (.A(net157),
    .X(_2855_));
 sg13g2_a21oi_1 _3448_ (.A1(_2853_),
    .A2(_2854_),
    .Y(_0029_),
    .B1(net106));
 sg13g2_inv_1 _3449_ (.Y(_2856_),
    .A(\Pong.control_unit.NES_Controller_Right.state_NESController[0] ));
 sg13g2_a21oi_1 _3450_ (.A1(\Pong.control_unit.NES_Controller_Right.state_NESController[6] ),
    .A2(net93),
    .Y(_2857_),
    .B1(net157));
 sg13g2_o21ai_1 _3451_ (.B1(_2857_),
    .Y(_0019_),
    .A1(_2856_),
    .A2(_2696_));
 sg13g2_nand2_1 _3452_ (.Y(_2858_),
    .A(\Pong.control_unit.NES_Controller_Left.state_NESController[9] ),
    .B(net91));
 sg13g2_nand2_1 _3453_ (.Y(_2859_),
    .A(_2841_),
    .B(net89));
 sg13g2_a21oi_1 _3454_ (.A1(_2858_),
    .A2(_2859_),
    .Y(_0009_),
    .B1(net106));
 sg13g2_nand2_1 _3455_ (.Y(_2860_),
    .A(_2797_),
    .B(net91));
 sg13g2_nand2_1 _3456_ (.Y(_2861_),
    .A(_2844_),
    .B(net89));
 sg13g2_a21oi_1 _3457_ (.A1(_2860_),
    .A2(_2861_),
    .Y(_0008_),
    .B1(net106));
 sg13g2_nor4_1 _3458_ (.A(\Pong.datapath.Ball_Clock.Q[14] ),
    .B(\Pong.datapath.Ball_Clock.Q[13] ),
    .C(\Pong.datapath.Ball_Clock.Q[12] ),
    .D(\Pong.datapath.Ball_Clock.Q[11] ),
    .Y(_2862_));
 sg13g2_buf_2 _3459_ (.A(\Pong.datapath.Ball_Clock.Q[0] ),
    .X(_2863_));
 sg13g2_nor4_1 _3460_ (.A(\Pong.datapath.Ball_Clock.Q[1] ),
    .B(_2863_),
    .C(\Pong.datapath.Ball_Clock.Q[3] ),
    .D(\Pong.datapath.Ball_Clock.Q[2] ),
    .Y(_2864_));
 sg13g2_buf_1 _3461_ (.A(\Pong.datapath.Ball_Clock.Q[5] ),
    .X(_2865_));
 sg13g2_inv_1 _3462_ (.Y(_2866_),
    .A(_2865_));
 sg13g2_buf_1 _3463_ (.A(\Pong.datapath.Ball_Clock.Q[6] ),
    .X(_2867_));
 sg13g2_nor3_1 _3464_ (.A(\Pong.datapath.Ball_Clock.Q[4] ),
    .B(_2866_),
    .C(_2867_),
    .Y(_2868_));
 sg13g2_nand2_1 _3465_ (.Y(_2869_),
    .A(\Pong.datapath.Ball_Clock.Q[10] ),
    .B(\Pong.datapath.Ball_Clock.Q[9] ));
 sg13g2_nand2b_1 _3466_ (.Y(_2870_),
    .B(\Pong.datapath.Ball_Clock.Q[7] ),
    .A_N(\Pong.datapath.Ball_Clock.Q[8] ));
 sg13g2_nand2_1 _3467_ (.Y(_2871_),
    .A(\Pong.datapath.Ball_Clock.Q[15] ),
    .B(\Pong.datapath.Ball_Clock.Q[16] ));
 sg13g2_nor3_1 _3468_ (.A(_2869_),
    .B(_2870_),
    .C(_2871_),
    .Y(_2872_));
 sg13g2_nand4_1 _3469_ (.B(_2864_),
    .C(_2868_),
    .A(_2862_),
    .Y(_2873_),
    .D(_2872_));
 sg13g2_buf_1 _3470_ (.A(_2873_),
    .X(_2874_));
 sg13g2_inv_1 _3471_ (.Y(\Pong.datapath.Ball_Clock.roll ),
    .A(_2874_));
 sg13g2_nand2_1 _3472_ (.Y(_2875_),
    .A(\Pong.control_unit.NES_Controller_Left.state_NESController[7] ),
    .B(net91));
 sg13g2_nand2_1 _3473_ (.Y(_2876_),
    .A(\Pong.control_unit.NES_Controller_Left.state_NESController[16] ),
    .B(net89));
 sg13g2_a21oi_1 _3474_ (.A1(_2875_),
    .A2(_2876_),
    .Y(_0007_),
    .B1(net106));
 sg13g2_nand2_1 _3475_ (.Y(_2877_),
    .A(\Pong.control_unit.NES_Controller_Left.state_NESController[5] ),
    .B(net91));
 sg13g2_nand2_1 _3476_ (.Y(_2878_),
    .A(\Pong.control_unit.NES_Controller_Left.state_NESController[15] ),
    .B(net89));
 sg13g2_a21oi_1 _3477_ (.A1(_2877_),
    .A2(_2878_),
    .Y(_0006_),
    .B1(net106));
 sg13g2_nand2_1 _3478_ (.Y(_2879_),
    .A(\Pong.control_unit.NES_Controller_Left.state_NESController[4] ),
    .B(net91));
 sg13g2_nand2_1 _3479_ (.Y(_2880_),
    .A(\Pong.control_unit.NES_Controller_Left.state_NESController[14] ),
    .B(net89));
 sg13g2_a21oi_1 _3480_ (.A1(_2879_),
    .A2(_2880_),
    .Y(_0005_),
    .B1(net106));
 sg13g2_nand2_1 _3481_ (.Y(_2881_),
    .A(_2806_),
    .B(net91));
 sg13g2_nand2_1 _3482_ (.Y(_2882_),
    .A(_2798_),
    .B(_2800_));
 sg13g2_a21oi_1 _3483_ (.A1(_2881_),
    .A2(_2882_),
    .Y(_0004_),
    .B1(_2855_));
 sg13g2_nand2_1 _3484_ (.Y(_2883_),
    .A(\Pong.control_unit.NES_Controller_Left.state_NESController[2] ),
    .B(_2786_));
 sg13g2_nand2_1 _3485_ (.Y(_2884_),
    .A(\Pong.control_unit.NES_Controller_Left.state_NESController[12] ),
    .B(_2800_));
 sg13g2_a21oi_1 _3486_ (.A1(_2883_),
    .A2(_2884_),
    .Y(_0003_),
    .B1(_2855_));
 sg13g2_buf_1 _3487_ (.A(_2771_),
    .X(_2885_));
 sg13g2_buf_1 _3488_ (.A(_2773_),
    .X(_2886_));
 sg13g2_buf_1 _3489_ (.A(net57),
    .X(_2887_));
 sg13g2_or2_1 _3490_ (.X(_2888_),
    .B(_2758_),
    .A(_2760_));
 sg13g2_buf_1 _3491_ (.A(_2888_),
    .X(_2889_));
 sg13g2_nor2_1 _3492_ (.A(net37),
    .B(_2889_),
    .Y(_2890_));
 sg13g2_nand4_1 _3493_ (.B(net61),
    .C(net54),
    .A(net55),
    .Y(_2891_),
    .D(_2890_));
 sg13g2_buf_1 _3494_ (.A(net56),
    .X(_2892_));
 sg13g2_buf_1 _3495_ (.A(_2772_),
    .X(_2893_));
 sg13g2_nor4_1 _3496_ (.A(net36),
    .B(net53),
    .C(net38),
    .D(net72),
    .Y(_2894_));
 sg13g2_nor2b_1 _3497_ (.A(_2891_),
    .B_N(_2894_),
    .Y(_0044_));
 sg13g2_buf_1 _3498_ (.A(\Pong.datapath.leftPaddle[8] ),
    .X(_2895_));
 sg13g2_buf_1 _3499_ (.A(_0060_),
    .X(_2896_));
 sg13g2_buf_1 _3500_ (.A(_2896_),
    .X(_2897_));
 sg13g2_nor2b_1 _3501_ (.A(net54),
    .B_N(net52),
    .Y(_2898_));
 sg13g2_buf_1 _3502_ (.A(_0070_),
    .X(_2899_));
 sg13g2_o21ai_1 _3503_ (.B1(net71),
    .Y(_2900_),
    .A1(net185),
    .A2(_2898_));
 sg13g2_buf_1 _3504_ (.A(\Pong.datapath.leftPaddle[2] ),
    .X(_2901_));
 sg13g2_buf_1 _3505_ (.A(net184),
    .X(_2902_));
 sg13g2_buf_2 _3506_ (.A(\Pong.datapath.leftPaddle[1] ),
    .X(_2903_));
 sg13g2_buf_8 _3507_ (.A(_2903_),
    .X(_2904_));
 sg13g2_buf_1 _3508_ (.A(net155),
    .X(_2905_));
 sg13g2_nor2_2 _3509_ (.A(net156),
    .B(net105),
    .Y(_2906_));
 sg13g2_buf_2 _3510_ (.A(\Pong.datapath.leftPaddle[4] ),
    .X(_2907_));
 sg13g2_buf_1 _3511_ (.A(\Pong.datapath.leftPaddle[3] ),
    .X(_2908_));
 sg13g2_nor2_1 _3512_ (.A(_2907_),
    .B(net183),
    .Y(_2909_));
 sg13g2_buf_1 _3513_ (.A(_2909_),
    .X(_2910_));
 sg13g2_buf_1 _3514_ (.A(\Pong.datapath.leftPaddle[6] ),
    .X(_2911_));
 sg13g2_buf_1 _3515_ (.A(\Pong.datapath.leftPaddle[5] ),
    .X(_2912_));
 sg13g2_nand2_1 _3516_ (.Y(_2913_),
    .A(_2911_),
    .B(net182));
 sg13g2_a21oi_2 _3517_ (.B1(_2913_),
    .Y(_2914_),
    .A2(net104),
    .A1(_2906_));
 sg13g2_nand2_1 _3518_ (.Y(_2915_),
    .A(net185),
    .B(_2914_));
 sg13g2_nand2b_1 _3519_ (.Y(_2916_),
    .B(_2914_),
    .A_N(_2900_));
 sg13g2_buf_1 _3520_ (.A(\Pong.datapath.leftPaddle[7] ),
    .X(_2917_));
 sg13g2_buf_1 _3521_ (.A(_2917_),
    .X(_2918_));
 sg13g2_inv_1 _3522_ (.Y(_2919_),
    .A(net154));
 sg13g2_buf_2 _3523_ (.A(_0059_),
    .X(_2920_));
 sg13g2_buf_2 _3524_ (.A(_0072_),
    .X(_2921_));
 sg13g2_xor2_1 _3525_ (.B(_2921_),
    .A(_2920_),
    .X(_2922_));
 sg13g2_a221oi_1 _3526_ (.B2(_2919_),
    .C1(_2922_),
    .B1(_2916_),
    .A1(_2900_),
    .Y(_2923_),
    .A2(_2915_));
 sg13g2_buf_1 _3527_ (.A(\Pong.datapath.leftPaddle[9] ),
    .X(_2924_));
 sg13g2_and2_1 _3528_ (.A(net154),
    .B(_2914_),
    .X(_2925_));
 sg13g2_buf_2 _3529_ (.A(_2925_),
    .X(_2926_));
 sg13g2_nand2_1 _3530_ (.Y(_2927_),
    .A(net185),
    .B(_2926_));
 sg13g2_o21ai_1 _3531_ (.B1(_2922_),
    .Y(_2928_),
    .A1(net181),
    .A2(_2927_));
 sg13g2_nor2b_1 _3532_ (.A(_2923_),
    .B_N(_2928_),
    .Y(_2929_));
 sg13g2_buf_1 _3533_ (.A(_2911_),
    .X(_2930_));
 sg13g2_nand2_2 _3534_ (.Y(_2931_),
    .A(_2906_),
    .B(net104));
 sg13g2_buf_1 _3535_ (.A(_0065_),
    .X(_2932_));
 sg13g2_buf_1 _3536_ (.A(net182),
    .X(_2933_));
 sg13g2_xnor2_1 _3537_ (.Y(_2934_),
    .A(net70),
    .B(net152));
 sg13g2_nand2_1 _3538_ (.Y(_2935_),
    .A(_2931_),
    .B(_2934_));
 sg13g2_or2_1 _3539_ (.X(_2936_),
    .B(_2934_),
    .A(_2931_));
 sg13g2_buf_1 _3540_ (.A(net183),
    .X(_2937_));
 sg13g2_or2_1 _3541_ (.X(_2938_),
    .B(net155),
    .A(net156));
 sg13g2_nor2_1 _3542_ (.A(net151),
    .B(_2938_),
    .Y(_2939_));
 sg13g2_xnor2_1 _3543_ (.Y(_2940_),
    .A(_0077_),
    .B(_2939_));
 sg13g2_nand2b_1 _3544_ (.Y(_2941_),
    .B(net38),
    .A_N(_2940_));
 sg13g2_buf_2 _3545_ (.A(_0066_),
    .X(_2942_));
 sg13g2_inv_2 _3546_ (.Y(_2943_),
    .A(_2942_));
 sg13g2_xnor2_1 _3547_ (.Y(_2944_),
    .A(_2943_),
    .B(_2940_));
 sg13g2_buf_1 _3548_ (.A(\Pong.datapath.leftPaddle[0] ),
    .X(_2945_));
 sg13g2_buf_1 _3549_ (.A(net180),
    .X(_2946_));
 sg13g2_nor2b_1 _3550_ (.A(net58),
    .B_N(net150),
    .Y(_2947_));
 sg13g2_xor2_1 _3551_ (.B(net156),
    .A(_0069_),
    .X(_2948_));
 sg13g2_nor3_1 _3552_ (.A(net105),
    .B(_2947_),
    .C(_2948_),
    .Y(_2949_));
 sg13g2_inv_1 _3553_ (.Y(_2950_),
    .A(_2905_));
 sg13g2_buf_1 _3554_ (.A(_0069_),
    .X(_2951_));
 sg13g2_xnor2_1 _3555_ (.Y(_2952_),
    .A(net69),
    .B(net156));
 sg13g2_nor2_1 _3556_ (.A(_2950_),
    .B(_2952_),
    .Y(_2953_));
 sg13g2_buf_1 _3557_ (.A(net59),
    .X(_2954_));
 sg13g2_o21ai_1 _3558_ (.B1(net35),
    .Y(_2955_),
    .A1(_2949_),
    .A2(_2953_));
 sg13g2_nor2_1 _3559_ (.A(_2950_),
    .B(_2947_),
    .Y(_2956_));
 sg13g2_xor2_1 _3560_ (.B(net105),
    .A(net156),
    .X(_2957_));
 sg13g2_a22oi_1 _3561_ (.Y(_2958_),
    .B1(_2957_),
    .B2(net37),
    .A2(_2956_),
    .A1(_2948_));
 sg13g2_buf_2 _3562_ (.A(_0078_),
    .X(_2959_));
 sg13g2_xnor2_1 _3563_ (.Y(_2960_),
    .A(_2959_),
    .B(_2906_));
 sg13g2_nand3_1 _3564_ (.B(_2958_),
    .C(_2960_),
    .A(_2955_),
    .Y(_2961_));
 sg13g2_nand3_1 _3565_ (.B(_2955_),
    .C(_2958_),
    .A(_2755_),
    .Y(_2962_));
 sg13g2_nand2_1 _3566_ (.Y(_2963_),
    .A(_2755_),
    .B(_2960_));
 sg13g2_nand4_1 _3567_ (.B(_2961_),
    .C(_2962_),
    .A(_2944_),
    .Y(_2964_),
    .D(_2963_));
 sg13g2_a22oi_1 _3568_ (.Y(_2965_),
    .B1(_2941_),
    .B2(_2964_),
    .A2(_2936_),
    .A1(_2935_));
 sg13g2_nor3_1 _3569_ (.A(_2751_),
    .B(net152),
    .C(_2931_),
    .Y(_2966_));
 sg13g2_buf_1 _3570_ (.A(net53),
    .X(_2967_));
 sg13g2_o21ai_1 _3571_ (.B1(net34),
    .Y(_2968_),
    .A1(_2965_),
    .A2(_2966_));
 sg13g2_nand2_1 _3572_ (.Y(_2969_),
    .A(net152),
    .B(_2931_));
 sg13g2_nand3_1 _3573_ (.B(_2968_),
    .C(_2969_),
    .A(net153),
    .Y(_2970_));
 sg13g2_o21ai_1 _3574_ (.B1(net34),
    .Y(_2971_),
    .A1(net153),
    .A2(_2969_));
 sg13g2_nand2_1 _3575_ (.Y(_2972_),
    .A(_2751_),
    .B(_2971_));
 sg13g2_nor2_1 _3576_ (.A(net34),
    .B(net153),
    .Y(_2973_));
 sg13g2_o21ai_1 _3577_ (.B1(_2973_),
    .Y(_2974_),
    .A1(net152),
    .A2(_2931_));
 sg13g2_a21oi_1 _3578_ (.A1(_2972_),
    .A2(_2974_),
    .Y(_2975_),
    .B1(_2965_));
 sg13g2_nor2b_1 _3579_ (.A(_2969_),
    .B_N(_2973_),
    .Y(_2976_));
 sg13g2_xnor2_1 _3580_ (.Y(_2977_),
    .A(net52),
    .B(net185));
 sg13g2_xor2_1 _3581_ (.B(_2977_),
    .A(_2926_),
    .X(_2978_));
 sg13g2_nor3_1 _3582_ (.A(_2975_),
    .B(_2976_),
    .C(_2978_),
    .Y(_2979_));
 sg13g2_nor3_1 _3583_ (.A(net154),
    .B(_2914_),
    .C(_2977_),
    .Y(_2980_));
 sg13g2_a21oi_1 _3584_ (.A1(_2926_),
    .A2(_2977_),
    .Y(_2981_),
    .B1(_2980_));
 sg13g2_nor2_1 _3585_ (.A(net71),
    .B(_2981_),
    .Y(_2982_));
 sg13g2_a21o_1 _3586_ (.A2(_2979_),
    .A1(_2970_),
    .B1(_2982_),
    .X(_2983_));
 sg13g2_buf_1 _3587_ (.A(_0073_),
    .X(_2984_));
 sg13g2_nand2_1 _3588_ (.Y(_2985_),
    .A(net184),
    .B(net155));
 sg13g2_nand2_2 _3589_ (.Y(_2986_),
    .A(_2907_),
    .B(net183));
 sg13g2_or2_1 _3590_ (.X(_2987_),
    .B(_2986_),
    .A(_2985_));
 sg13g2_buf_2 _3591_ (.A(_2987_),
    .X(_2988_));
 sg13g2_nor2_1 _3592_ (.A(net182),
    .B(_2988_),
    .Y(_2989_));
 sg13g2_buf_1 _3593_ (.A(_0071_),
    .X(_2990_));
 sg13g2_buf_1 _3594_ (.A(_2990_),
    .X(_2991_));
 sg13g2_nor2_1 _3595_ (.A(net154),
    .B(net153),
    .Y(_2992_));
 sg13g2_nand2_1 _3596_ (.Y(_2993_),
    .A(net149),
    .B(_2992_));
 sg13g2_nor2_1 _3597_ (.A(_2989_),
    .B(_2993_),
    .Y(_2994_));
 sg13g2_xnor2_1 _3598_ (.Y(_2995_),
    .A(net179),
    .B(_2994_));
 sg13g2_or2_1 _3599_ (.X(_2996_),
    .B(net182),
    .A(_2911_));
 sg13g2_buf_1 _3600_ (.A(_2996_),
    .X(_2997_));
 sg13g2_nor2b_1 _3601_ (.A(_2997_),
    .B_N(_2988_),
    .Y(_2998_));
 sg13g2_xnor2_1 _3602_ (.Y(_2999_),
    .A(_0074_),
    .B(_2998_));
 sg13g2_inv_1 _3603_ (.Y(_3000_),
    .A(net55));
 sg13g2_nor3_1 _3604_ (.A(_2895_),
    .B(net154),
    .C(_2997_),
    .Y(_3001_));
 sg13g2_nand2_1 _3605_ (.Y(_3002_),
    .A(_2988_),
    .B(_3001_));
 sg13g2_xnor2_1 _3606_ (.Y(_3003_),
    .A(_2921_),
    .B(_3002_));
 sg13g2_xor2_1 _3607_ (.B(_3003_),
    .A(_2920_),
    .X(_3004_));
 sg13g2_a221oi_1 _3608_ (.B2(_3000_),
    .C1(_3004_),
    .B1(_2999_),
    .A1(_2897_),
    .Y(_3005_),
    .A2(_2995_));
 sg13g2_inv_1 _3609_ (.Y(_3006_),
    .A(_0075_));
 sg13g2_inv_1 _3610_ (.Y(_3007_),
    .A(net184));
 sg13g2_nor4_1 _3611_ (.A(net152),
    .B(_3007_),
    .C(_0076_),
    .D(_2986_),
    .Y(_3008_));
 sg13g2_nor2b_1 _3612_ (.A(_3008_),
    .B_N(net149),
    .Y(_3009_));
 sg13g2_xnor2_1 _3613_ (.Y(_3010_),
    .A(_3006_),
    .B(_3009_));
 sg13g2_nand3_1 _3614_ (.B(_3005_),
    .C(_3010_),
    .A(net34),
    .Y(_3011_));
 sg13g2_inv_1 _3615_ (.Y(_3012_),
    .A(_3004_));
 sg13g2_nand2b_1 _3616_ (.Y(_3013_),
    .B(net55),
    .A_N(_2999_));
 sg13g2_a21o_1 _3617_ (.A2(_3013_),
    .A1(_2995_),
    .B1(net52),
    .X(_3014_));
 sg13g2_o21ai_1 _3618_ (.B1(_3014_),
    .Y(_3015_),
    .A1(_2995_),
    .A2(_3013_));
 sg13g2_xnor2_1 _3619_ (.Y(_3016_),
    .A(net152),
    .B(_2988_));
 sg13g2_inv_2 _3620_ (.Y(_3017_),
    .A(_0077_));
 sg13g2_nand3_1 _3621_ (.B(net156),
    .C(net105),
    .A(net151),
    .Y(_3018_));
 sg13g2_xnor2_1 _3622_ (.Y(_3019_),
    .A(_3017_),
    .B(_3018_));
 sg13g2_xor2_1 _3623_ (.B(_2988_),
    .A(_2934_),
    .X(_3020_));
 sg13g2_a21oi_1 _3624_ (.A1(_2942_),
    .A2(_3019_),
    .Y(_3021_),
    .B1(_3020_));
 sg13g2_nor2_1 _3625_ (.A(_2942_),
    .B(_3019_),
    .Y(_3022_));
 sg13g2_a22oi_1 _3626_ (.Y(_3023_),
    .B1(_3021_),
    .B2(_3022_),
    .A2(_3016_),
    .A1(net61));
 sg13g2_or3_1 _3627_ (.A(net105),
    .B(_2947_),
    .C(_2952_),
    .X(_3024_));
 sg13g2_o21ai_1 _3628_ (.B1(_3024_),
    .Y(_3025_),
    .A1(_2950_),
    .A2(_2948_));
 sg13g2_inv_2 _3629_ (.Y(_3026_),
    .A(net57));
 sg13g2_nor2_1 _3630_ (.A(_3026_),
    .B(_2957_),
    .Y(_3027_));
 sg13g2_a221oi_1 _3631_ (.B2(net35),
    .C1(_3027_),
    .B1(_3025_),
    .A1(_2952_),
    .Y(_3028_),
    .A2(_2956_));
 sg13g2_xor2_1 _3632_ (.B(_2985_),
    .A(_2959_),
    .X(_3029_));
 sg13g2_nand2_1 _3633_ (.Y(_3030_),
    .A(_3028_),
    .B(_3029_));
 sg13g2_o21ai_1 _3634_ (.B1(_2767_),
    .Y(_3031_),
    .A1(_3028_),
    .A2(_3029_));
 sg13g2_nand3_1 _3635_ (.B(_3030_),
    .C(_3031_),
    .A(_3021_),
    .Y(_3032_));
 sg13g2_buf_2 _3636_ (.A(_0064_),
    .X(_3033_));
 sg13g2_xnor2_1 _3637_ (.Y(_3034_),
    .A(_3033_),
    .B(_3010_));
 sg13g2_nand2_1 _3638_ (.Y(_3035_),
    .A(_3005_),
    .B(_3034_));
 sg13g2_a21oi_1 _3639_ (.A1(_3023_),
    .A2(_3032_),
    .Y(_3036_),
    .B1(_3035_));
 sg13g2_a221oi_1 _3640_ (.B2(_3015_),
    .C1(_3036_),
    .B1(_3012_),
    .A1(net72),
    .Y(_3037_),
    .A2(_3003_));
 sg13g2_or2_1 _3641_ (.X(_3038_),
    .B(_0044_),
    .A(_0043_));
 sg13g2_buf_1 _3642_ (.A(_3038_),
    .X(_3039_));
 sg13g2_nor4_1 _3643_ (.A(net181),
    .B(net185),
    .C(_2989_),
    .D(_2993_),
    .Y(_3040_));
 sg13g2_buf_2 _3644_ (.A(\Pong.datapath.ballFunction.ball_center_x[6] ),
    .X(_3041_));
 sg13g2_buf_1 _3645_ (.A(\Pong.datapath.ballFunction.ball_center_x[7] ),
    .X(_3042_));
 sg13g2_buf_1 _3646_ (.A(\Pong.datapath.ballFunction.ball_center_x[8] ),
    .X(_3043_));
 sg13g2_buf_1 _3647_ (.A(\Pong.datapath.ballFunction.ball_center_x[9] ),
    .X(_3044_));
 sg13g2_nor4_2 _3648_ (.A(_3041_),
    .B(net68),
    .C(_3043_),
    .Y(_3045_),
    .D(_3044_));
 sg13g2_buf_2 _3649_ (.A(\Pong.datapath.ballFunction.ball_center_x[3] ),
    .X(_3046_));
 sg13g2_buf_8 _3650_ (.A(_3046_),
    .X(_3047_));
 sg13g2_buf_1 _3651_ (.A(\Pong.datapath.ballFunction.ball_center_x[2] ),
    .X(_3048_));
 sg13g2_buf_1 _3652_ (.A(net67),
    .X(_3049_));
 sg13g2_buf_2 _3653_ (.A(\Pong.datapath.ballFunction.ball_center_x[0] ),
    .X(_3050_));
 sg13g2_buf_1 _3654_ (.A(\Pong.datapath.ballFunction.ball_center_x[1] ),
    .X(_3051_));
 sg13g2_and2_1 _3655_ (.A(_3050_),
    .B(_3051_),
    .X(_3052_));
 sg13g2_buf_2 _3656_ (.A(_3052_),
    .X(_3053_));
 sg13g2_nand3_1 _3657_ (.B(net50),
    .C(_3053_),
    .A(net51),
    .Y(_3054_));
 sg13g2_inv_1 _3658_ (.Y(_3055_),
    .A(_3054_));
 sg13g2_buf_2 _3659_ (.A(\Pong.datapath.ballFunction.ball_center_x[5] ),
    .X(_3056_));
 sg13g2_inv_2 _3660_ (.Y(_3057_),
    .A(_3056_));
 sg13g2_buf_1 _3661_ (.A(\Pong.datapath.ballFunction.ball_center_x[4] ),
    .X(_3058_));
 sg13g2_nor2_1 _3662_ (.A(_3057_),
    .B(_3058_),
    .Y(_3059_));
 sg13g2_nand3_1 _3663_ (.B(_3055_),
    .C(_3059_),
    .A(_3045_),
    .Y(_3060_));
 sg13g2_nor3_1 _3664_ (.A(_3039_),
    .B(_3040_),
    .C(_3060_),
    .Y(_3061_));
 sg13g2_nor3_1 _3665_ (.A(net181),
    .B(_2921_),
    .C(_2927_),
    .Y(_3062_));
 sg13g2_inv_1 _3666_ (.Y(_3063_),
    .A(_2921_));
 sg13g2_a21oi_1 _3667_ (.A1(net185),
    .A2(_2926_),
    .Y(_3064_),
    .B1(_3063_));
 sg13g2_o21ai_1 _3668_ (.B1(net72),
    .Y(_3065_),
    .A1(_3062_),
    .A2(_3064_));
 sg13g2_xnor2_1 _3669_ (.Y(_3066_),
    .A(net185),
    .B(_2926_));
 sg13g2_nand3_1 _3670_ (.B(_2929_),
    .C(_3066_),
    .A(net54),
    .Y(_3067_));
 sg13g2_nand3_1 _3671_ (.B(_2950_),
    .C(_2948_),
    .A(net35),
    .Y(_3068_));
 sg13g2_inv_1 _3672_ (.Y(_0300_),
    .A(net35));
 sg13g2_nand3_1 _3673_ (.B(net105),
    .C(_2952_),
    .A(_0300_),
    .Y(_0301_));
 sg13g2_xnor2_1 _3674_ (.Y(_0302_),
    .A(_2767_),
    .B(_3029_));
 sg13g2_a21oi_1 _3675_ (.A1(_3068_),
    .A2(_0301_),
    .Y(_0303_),
    .B1(_0302_));
 sg13g2_inv_1 _3676_ (.Y(_0304_),
    .A(net58));
 sg13g2_nor2_1 _3677_ (.A(_0304_),
    .B(net150),
    .Y(_0305_));
 sg13g2_nor3_1 _3678_ (.A(_2947_),
    .B(_3022_),
    .C(_0305_),
    .Y(_0306_));
 sg13g2_nand4_1 _3679_ (.B(_3013_),
    .C(_0303_),
    .A(_3021_),
    .Y(_0307_),
    .D(_0306_));
 sg13g2_nor2_1 _3680_ (.A(net52),
    .B(_2995_),
    .Y(_0308_));
 sg13g2_or3_1 _3681_ (.A(_3035_),
    .B(_0307_),
    .C(_0308_),
    .X(_0309_));
 sg13g2_nand4_1 _3682_ (.B(_3065_),
    .C(_3067_),
    .A(_3061_),
    .Y(_0310_),
    .D(_0309_));
 sg13g2_a221oi_1 _3683_ (.B2(_3037_),
    .C1(_0310_),
    .B1(_3011_),
    .A1(_2929_),
    .Y(_0045_),
    .A2(_2983_));
 sg13g2_buf_2 _3684_ (.A(\Pong.datapath.rightPaddle[5] ),
    .X(_0311_));
 sg13g2_buf_1 _3685_ (.A(_0311_),
    .X(_0312_));
 sg13g2_inv_2 _3686_ (.Y(_0313_),
    .A(net148));
 sg13g2_buf_1 _3687_ (.A(\Pong.datapath.rightPaddle[4] ),
    .X(_0314_));
 sg13g2_buf_2 _3688_ (.A(\Pong.datapath.rightPaddle[2] ),
    .X(_0315_));
 sg13g2_buf_8 _3689_ (.A(_0315_),
    .X(_0316_));
 sg13g2_buf_1 _3690_ (.A(\Pong.datapath.rightPaddle[3] ),
    .X(_0317_));
 sg13g2_buf_1 _3691_ (.A(\Pong.datapath.rightPaddle[1] ),
    .X(_0318_));
 sg13g2_nand4_1 _3692_ (.B(net147),
    .C(_0317_),
    .A(net178),
    .Y(_0319_),
    .D(net177));
 sg13g2_buf_1 _3693_ (.A(_0319_),
    .X(_0320_));
 sg13g2_xnor2_1 _3694_ (.Y(_0321_),
    .A(_0313_),
    .B(_0320_));
 sg13g2_buf_2 _3695_ (.A(_0067_),
    .X(_0322_));
 sg13g2_inv_1 _3696_ (.Y(_0323_),
    .A(_0322_));
 sg13g2_buf_1 _3697_ (.A(net147),
    .X(_0324_));
 sg13g2_buf_1 _3698_ (.A(_0317_),
    .X(_0325_));
 sg13g2_buf_2 _3699_ (.A(net177),
    .X(_0326_));
 sg13g2_buf_1 _3700_ (.A(net145),
    .X(_0327_));
 sg13g2_nand3_1 _3701_ (.B(net146),
    .C(_0327_),
    .A(_0324_),
    .Y(_0328_));
 sg13g2_xnor2_1 _3702_ (.Y(_0329_),
    .A(_0323_),
    .B(_0328_));
 sg13g2_inv_1 _3703_ (.Y(_0330_),
    .A(_0329_));
 sg13g2_nor2_1 _3704_ (.A(_2943_),
    .B(_0330_),
    .Y(_0331_));
 sg13g2_buf_1 _3705_ (.A(_0068_),
    .X(_0332_));
 sg13g2_buf_1 _3706_ (.A(_0332_),
    .X(_0333_));
 sg13g2_nand2_1 _3707_ (.Y(_0334_),
    .A(net56),
    .B(net144));
 sg13g2_nor2b_1 _3708_ (.A(net102),
    .B_N(net57),
    .Y(_0335_));
 sg13g2_o21ai_1 _3709_ (.B1(_0335_),
    .Y(_0336_),
    .A1(net36),
    .A2(net144));
 sg13g2_a21oi_1 _3710_ (.A1(_0334_),
    .A2(_0336_),
    .Y(_0337_),
    .B1(net103));
 sg13g2_nand2_1 _3711_ (.Y(_0338_),
    .A(net147),
    .B(net145));
 sg13g2_nand2b_1 _3712_ (.Y(_0339_),
    .B(net144),
    .A_N(net56));
 sg13g2_nor2b_1 _3713_ (.A(net144),
    .B_N(_2766_),
    .Y(_0340_));
 sg13g2_a21oi_1 _3714_ (.A1(net57),
    .A2(_0339_),
    .Y(_0341_),
    .B1(_0340_));
 sg13g2_inv_1 _3715_ (.Y(_0342_),
    .A(net145));
 sg13g2_nand2b_1 _3716_ (.Y(_0343_),
    .B(_0342_),
    .A_N(_0334_));
 sg13g2_o21ai_1 _3717_ (.B1(_0343_),
    .Y(_0344_),
    .A1(_0338_),
    .A2(_0341_));
 sg13g2_inv_1 _3718_ (.Y(_0345_),
    .A(_0332_));
 sg13g2_xnor2_1 _3719_ (.Y(_0346_),
    .A(_0345_),
    .B(_0338_));
 sg13g2_buf_1 _3720_ (.A(\Pong.datapath.rightPaddle[0] ),
    .X(_0347_));
 sg13g2_buf_1 _3721_ (.A(net176),
    .X(_0348_));
 sg13g2_nand2b_1 _3722_ (.Y(_0349_),
    .B(net143),
    .A_N(net58));
 sg13g2_nand2_1 _3723_ (.Y(_0350_),
    .A(net102),
    .B(_0349_));
 sg13g2_o21ai_1 _3724_ (.B1(net59),
    .Y(_0351_),
    .A1(net102),
    .A2(_0349_));
 sg13g2_xor2_1 _3725_ (.B(net145),
    .A(net147),
    .X(_0352_));
 sg13g2_xnor2_1 _3726_ (.Y(_0353_),
    .A(net69),
    .B(_0352_));
 sg13g2_a221oi_1 _3727_ (.B2(_0351_),
    .C1(_0353_),
    .B1(_0350_),
    .A1(_2767_),
    .Y(_0354_),
    .A2(_0346_));
 sg13g2_nor4_1 _3728_ (.A(_0330_),
    .B(_0337_),
    .C(_0344_),
    .D(_0354_),
    .Y(_0355_));
 sg13g2_nor4_1 _3729_ (.A(_2943_),
    .B(_0337_),
    .C(_0344_),
    .D(_0354_),
    .Y(_0356_));
 sg13g2_nor3_1 _3730_ (.A(_0331_),
    .B(_0355_),
    .C(_0356_),
    .Y(_0357_));
 sg13g2_nand2b_1 _3731_ (.Y(_0358_),
    .B(_0357_),
    .A_N(net70));
 sg13g2_nor2_1 _3732_ (.A(net61),
    .B(_0321_),
    .Y(_0359_));
 sg13g2_nand2_1 _3733_ (.Y(_0360_),
    .A(net70),
    .B(_0357_));
 sg13g2_buf_2 _3734_ (.A(_0061_),
    .X(_0361_));
 sg13g2_nor2_1 _3735_ (.A(net148),
    .B(_0320_),
    .Y(_0362_));
 sg13g2_buf_1 _3736_ (.A(\Pong.datapath.rightPaddle[7] ),
    .X(_0363_));
 sg13g2_buf_2 _3737_ (.A(\Pong.datapath.rightPaddle[6] ),
    .X(_0364_));
 sg13g2_buf_1 _3738_ (.A(_0364_),
    .X(_0365_));
 sg13g2_nor2_1 _3739_ (.A(_0363_),
    .B(net142),
    .Y(_0366_));
 sg13g2_nand2_2 _3740_ (.Y(_0367_),
    .A(_0057_),
    .B(_0366_));
 sg13g2_nor2_1 _3741_ (.A(_0362_),
    .B(_0367_),
    .Y(_0368_));
 sg13g2_xnor2_1 _3742_ (.Y(_0369_),
    .A(_0361_),
    .B(_0368_));
 sg13g2_buf_1 _3743_ (.A(\Pong.datapath.rightPaddle[8] ),
    .X(_0370_));
 sg13g2_nor4_2 _3744_ (.A(_0370_),
    .B(_0363_),
    .C(_0364_),
    .Y(_0371_),
    .D(_0311_));
 sg13g2_nand2_1 _3745_ (.Y(_0372_),
    .A(_0320_),
    .B(_0371_));
 sg13g2_buf_2 _3746_ (.A(_0058_),
    .X(_0373_));
 sg13g2_xnor2_1 _3747_ (.Y(_0374_),
    .A(_0373_),
    .B(_2920_));
 sg13g2_xor2_1 _3748_ (.B(_0374_),
    .A(_0372_),
    .X(_0375_));
 sg13g2_a21o_1 _3749_ (.A2(_0369_),
    .A1(net52),
    .B1(_0375_),
    .X(_0376_));
 sg13g2_nor2_1 _3750_ (.A(net142),
    .B(net148),
    .Y(_0377_));
 sg13g2_nand2_1 _3751_ (.Y(_0378_),
    .A(_0320_),
    .B(_0377_));
 sg13g2_xnor2_1 _3752_ (.Y(_0379_),
    .A(_0062_),
    .B(_0378_));
 sg13g2_nor2_1 _3753_ (.A(net55),
    .B(_0379_),
    .Y(_0380_));
 sg13g2_buf_2 _3754_ (.A(_0063_),
    .X(_0381_));
 sg13g2_buf_1 _3755_ (.A(net148),
    .X(_0382_));
 sg13g2_buf_1 _3756_ (.A(_0057_),
    .X(_0383_));
 sg13g2_o21ai_1 _3757_ (.B1(net175),
    .Y(_0384_),
    .A1(net101),
    .A2(_0320_));
 sg13g2_xor2_1 _3758_ (.B(_0384_),
    .A(_0381_),
    .X(_0385_));
 sg13g2_xnor2_1 _3759_ (.Y(_0386_),
    .A(_3033_),
    .B(_0385_));
 sg13g2_or3_1 _3760_ (.A(_0376_),
    .B(_0380_),
    .C(_0386_),
    .X(_0387_));
 sg13g2_a221oi_1 _3761_ (.B2(_0360_),
    .C1(_0387_),
    .B1(_0359_),
    .A1(_0321_),
    .Y(_0388_),
    .A2(_0358_));
 sg13g2_nor2_1 _3762_ (.A(_2897_),
    .B(_0369_),
    .Y(_0389_));
 sg13g2_a21o_1 _3763_ (.A2(_0389_),
    .A1(_2920_),
    .B1(_2774_),
    .X(_0390_));
 sg13g2_xnor2_1 _3764_ (.Y(_0391_),
    .A(_0373_),
    .B(_0372_));
 sg13g2_nor2_1 _3765_ (.A(_2920_),
    .B(_0391_),
    .Y(_0392_));
 sg13g2_a22oi_1 _3766_ (.Y(_0393_),
    .B1(_0392_),
    .B2(_0389_),
    .A2(_0391_),
    .A1(_0390_));
 sg13g2_nand2_1 _3767_ (.Y(_0394_),
    .A(net55),
    .B(_0379_));
 sg13g2_nor2b_1 _3768_ (.A(_0385_),
    .B_N(net34),
    .Y(_0395_));
 sg13g2_o21ai_1 _3769_ (.B1(_0395_),
    .Y(_0396_),
    .A1(net55),
    .A2(_0379_));
 sg13g2_a21o_1 _3770_ (.A2(_0396_),
    .A1(_0394_),
    .B1(_0376_),
    .X(_0397_));
 sg13g2_nand3b_1 _3771_ (.B(_0393_),
    .C(_0397_),
    .Y(_0398_),
    .A_N(_0388_));
 sg13g2_buf_1 _3772_ (.A(_0370_),
    .X(_0399_));
 sg13g2_buf_1 _3773_ (.A(_0363_),
    .X(_0400_));
 sg13g2_nor2_2 _3774_ (.A(net147),
    .B(net145),
    .Y(_0401_));
 sg13g2_nor2_1 _3775_ (.A(net178),
    .B(_0317_),
    .Y(_0402_));
 sg13g2_buf_1 _3776_ (.A(_0402_),
    .X(_0403_));
 sg13g2_nand2_1 _3777_ (.Y(_0404_),
    .A(_0364_),
    .B(_0311_));
 sg13g2_a21oi_2 _3778_ (.B1(_0404_),
    .Y(_0405_),
    .A2(net100),
    .A1(_0401_));
 sg13g2_and2_1 _3779_ (.A(net140),
    .B(_0405_),
    .X(_0406_));
 sg13g2_buf_1 _3780_ (.A(_0406_),
    .X(_0407_));
 sg13g2_nand2_1 _3781_ (.Y(_0408_),
    .A(net141),
    .B(_0407_));
 sg13g2_buf_1 _3782_ (.A(\Pong.datapath.rightPaddle[9] ),
    .X(_0409_));
 sg13g2_nor3_1 _3783_ (.A(net174),
    .B(_0374_),
    .C(_0408_),
    .Y(_0410_));
 sg13g2_a21oi_1 _3784_ (.A1(_0374_),
    .A2(_0408_),
    .Y(_0411_),
    .B1(_0410_));
 sg13g2_or2_1 _3785_ (.X(_0412_),
    .B(net145),
    .A(net147));
 sg13g2_buf_1 _3786_ (.A(_0412_),
    .X(_0413_));
 sg13g2_or2_1 _3787_ (.X(_0414_),
    .B(net146),
    .A(net178));
 sg13g2_o21ai_1 _3788_ (.B1(net148),
    .Y(_0415_),
    .A1(_0413_),
    .A2(_0414_));
 sg13g2_xor2_1 _3789_ (.B(_0415_),
    .A(net142),
    .X(_0416_));
 sg13g2_nor2_1 _3790_ (.A(_2967_),
    .B(_0416_),
    .Y(_0417_));
 sg13g2_nor2_1 _3791_ (.A(_2750_),
    .B(net70),
    .Y(_0418_));
 sg13g2_nand3_1 _3792_ (.B(_0401_),
    .C(net100),
    .A(_0313_),
    .Y(_0419_));
 sg13g2_nand2_1 _3793_ (.Y(_0420_),
    .A(_0415_),
    .B(_0419_));
 sg13g2_mux2_1 _3794_ (.A0(net70),
    .A1(_0418_),
    .S(_0420_),
    .X(_0421_));
 sg13g2_nor3_1 _3795_ (.A(_0411_),
    .B(_0417_),
    .C(_0421_),
    .Y(_0422_));
 sg13g2_xnor2_1 _3796_ (.Y(_0423_),
    .A(net141),
    .B(net52));
 sg13g2_a21oi_1 _3797_ (.A1(net71),
    .A2(_0405_),
    .Y(_0424_),
    .B1(net140));
 sg13g2_nor2_1 _3798_ (.A(net71),
    .B(_0405_),
    .Y(_0425_));
 sg13g2_nor2_1 _3799_ (.A(_0424_),
    .B(_0425_),
    .Y(_0426_));
 sg13g2_nand2_1 _3800_ (.Y(_0427_),
    .A(_0407_),
    .B(_0423_));
 sg13g2_o21ai_1 _3801_ (.B1(_0427_),
    .Y(_0428_),
    .A1(_0423_),
    .A2(_0426_));
 sg13g2_nor2b_1 _3802_ (.A(net58),
    .B_N(net143),
    .Y(_0429_));
 sg13g2_xor2_1 _3803_ (.B(net69),
    .A(net103),
    .X(_0430_));
 sg13g2_nor3_1 _3804_ (.A(net102),
    .B(_0429_),
    .C(_0430_),
    .Y(_0431_));
 sg13g2_and2_1 _3805_ (.A(net102),
    .B(_0430_),
    .X(_0432_));
 sg13g2_o21ai_1 _3806_ (.B1(_2954_),
    .Y(_0433_),
    .A1(_0431_),
    .A2(_0432_));
 sg13g2_nor2_1 _3807_ (.A(_0342_),
    .B(_0429_),
    .Y(_0434_));
 sg13g2_a22oi_1 _3808_ (.Y(_0435_),
    .B1(_0434_),
    .B2(_0430_),
    .A2(_0352_),
    .A1(net37));
 sg13g2_xnor2_1 _3809_ (.Y(_0436_),
    .A(net144),
    .B(_0401_));
 sg13g2_nand3_1 _3810_ (.B(_0435_),
    .C(_0436_),
    .A(_0433_),
    .Y(_0437_));
 sg13g2_nand2_1 _3811_ (.Y(_0438_),
    .A(_2756_),
    .B(_0437_));
 sg13g2_a21o_1 _3812_ (.A2(_0435_),
    .A1(_0433_),
    .B1(_0436_),
    .X(_0439_));
 sg13g2_buf_1 _3813_ (.A(net146),
    .X(_0440_));
 sg13g2_nor2_1 _3814_ (.A(net99),
    .B(_0413_),
    .Y(_0441_));
 sg13g2_xnor2_1 _3815_ (.Y(_0442_),
    .A(_0322_),
    .B(_0441_));
 sg13g2_xnor2_1 _3816_ (.Y(_0443_),
    .A(_2942_),
    .B(_0442_));
 sg13g2_a21oi_1 _3817_ (.A1(_0438_),
    .A2(_0439_),
    .Y(_0444_),
    .B1(_0443_));
 sg13g2_nor2b_1 _3818_ (.A(_0442_),
    .B_N(net38),
    .Y(_0445_));
 sg13g2_a21oi_1 _3819_ (.A1(_2750_),
    .A2(_0420_),
    .Y(_0446_),
    .B1(_0445_));
 sg13g2_nand2b_1 _3820_ (.Y(_0447_),
    .B(_0446_),
    .A_N(_0444_));
 sg13g2_nand3_1 _3821_ (.B(_0428_),
    .C(_0447_),
    .A(_0422_),
    .Y(_0448_));
 sg13g2_xnor2_1 _3822_ (.Y(_0449_),
    .A(net141),
    .B(_0407_));
 sg13g2_or2_1 _3823_ (.X(_0450_),
    .B(_0423_),
    .A(net140));
 sg13g2_o21ai_1 _3824_ (.B1(_0427_),
    .Y(_0451_),
    .A1(_0405_),
    .A2(_0450_));
 sg13g2_nand2_1 _3825_ (.Y(_0452_),
    .A(_2967_),
    .B(_0416_));
 sg13g2_nand2_1 _3826_ (.Y(_0453_),
    .A(net71),
    .B(_0452_));
 sg13g2_nor4_1 _3827_ (.A(_2899_),
    .B(_0407_),
    .C(_0423_),
    .D(_0452_),
    .Y(_0454_));
 sg13g2_a221oi_1 _3828_ (.B2(_0453_),
    .C1(_0454_),
    .B1(_0451_),
    .A1(_2886_),
    .Y(_0455_),
    .A2(_0449_));
 sg13g2_nor2_1 _3829_ (.A(_0411_),
    .B(_0455_),
    .Y(_0456_));
 sg13g2_nor3_1 _3830_ (.A(net174),
    .B(_0373_),
    .C(_0408_),
    .Y(_0457_));
 sg13g2_a21oi_1 _3831_ (.A1(_0373_),
    .A2(_0408_),
    .Y(_0458_),
    .B1(_0457_));
 sg13g2_nor2b_1 _3832_ (.A(_0458_),
    .B_N(_2774_),
    .Y(_0459_));
 sg13g2_buf_1 _3833_ (.A(_3050_),
    .X(_0460_));
 sg13g2_nor2_2 _3834_ (.A(net68),
    .B(_3043_),
    .Y(_0461_));
 sg13g2_or2_1 _3835_ (.X(_0462_),
    .B(net67),
    .A(_3051_));
 sg13g2_buf_1 _3836_ (.A(_0462_),
    .X(_0463_));
 sg13g2_nor2_1 _3837_ (.A(_3047_),
    .B(_0463_),
    .Y(_0464_));
 sg13g2_buf_1 _3838_ (.A(_3041_),
    .X(_0465_));
 sg13g2_buf_1 _3839_ (.A(_3044_),
    .X(_0466_));
 sg13g2_buf_1 _3840_ (.A(_3058_),
    .X(_0467_));
 sg13g2_nor2b_1 _3841_ (.A(_3056_),
    .B_N(_0467_),
    .Y(_0468_));
 sg13g2_and3_1 _3842_ (.X(_0469_),
    .A(net48),
    .B(net47),
    .C(_0468_));
 sg13g2_nand4_1 _3843_ (.B(_0461_),
    .C(_0464_),
    .A(net49),
    .Y(_0470_),
    .D(_0469_));
 sg13g2_nor4_1 _3844_ (.A(net174),
    .B(net141),
    .C(_0362_),
    .D(_0367_),
    .Y(_0471_));
 sg13g2_nor4_1 _3845_ (.A(_0456_),
    .B(_0459_),
    .C(_0470_),
    .D(_0471_),
    .Y(_0472_));
 sg13g2_xor2_1 _3846_ (.B(_0321_),
    .A(_2932_),
    .X(_0473_));
 sg13g2_xnor2_1 _3847_ (.Y(_0474_),
    .A(_2943_),
    .B(_0329_));
 sg13g2_a21o_1 _3848_ (.A2(_0346_),
    .A1(_2767_),
    .B1(_0353_),
    .X(_0475_));
 sg13g2_xnor2_1 _3849_ (.Y(_0476_),
    .A(net58),
    .B(net143));
 sg13g2_o21ai_1 _3850_ (.B1(_0476_),
    .Y(_0477_),
    .A1(net103),
    .A2(_0334_));
 sg13g2_nand2_1 _3851_ (.Y(_0478_),
    .A(net103),
    .B(_0340_));
 sg13g2_nor2_1 _3852_ (.A(_2954_),
    .B(_0342_),
    .Y(_0479_));
 sg13g2_nor2_1 _3853_ (.A(_0300_),
    .B(net102),
    .Y(_0480_));
 sg13g2_a22oi_1 _3854_ (.Y(_0481_),
    .B1(_0480_),
    .B2(_0334_),
    .A2(_0479_),
    .A1(_0478_));
 sg13g2_nor4_1 _3855_ (.A(_0389_),
    .B(_0475_),
    .C(_0477_),
    .D(_0481_),
    .Y(_0482_));
 sg13g2_nand4_1 _3856_ (.B(_0473_),
    .C(_0474_),
    .A(_0394_),
    .Y(_0483_),
    .D(_0482_));
 sg13g2_or2_1 _3857_ (.X(_0484_),
    .B(_0483_),
    .A(_0387_));
 sg13g2_nand4_1 _3858_ (.B(_0448_),
    .C(_0472_),
    .A(_0398_),
    .Y(_0485_),
    .D(_0484_));
 sg13g2_nor2_1 _3859_ (.A(_3039_),
    .B(_0485_),
    .Y(_0046_));
 sg13g2_buf_1 _3860_ (.A(net51),
    .X(_0486_));
 sg13g2_buf_1 _3861_ (.A(net46),
    .X(_0487_));
 sg13g2_and2_1 _3862_ (.A(_3056_),
    .B(_3041_),
    .X(_0488_));
 sg13g2_buf_1 _3863_ (.A(_0488_),
    .X(_0489_));
 sg13g2_o21ai_1 _3864_ (.B1(_0489_),
    .Y(_0490_),
    .A1(net33),
    .A2(net32));
 sg13g2_buf_1 _3865_ (.A(_3043_),
    .X(_0491_));
 sg13g2_buf_1 _3866_ (.A(_0079_),
    .X(_0492_));
 sg13g2_nor2b_1 _3867_ (.A(_0491_),
    .B_N(_0492_),
    .Y(_0493_));
 sg13g2_o21ai_1 _3868_ (.B1(_0493_),
    .Y(_0494_),
    .A1(net68),
    .A2(_0490_));
 sg13g2_and2_1 _3869_ (.A(_3057_),
    .B(_3045_),
    .X(_0495_));
 sg13g2_buf_2 _3870_ (.A(_0080_),
    .X(_0496_));
 sg13g2_nand2b_1 _3871_ (.Y(_0497_),
    .B(net32),
    .A_N(_0496_));
 sg13g2_nor2_1 _3872_ (.A(_3041_),
    .B(_3044_),
    .Y(_0498_));
 sg13g2_nand2_1 _3873_ (.Y(_0499_),
    .A(_0498_),
    .B(_0468_));
 sg13g2_nand3_1 _3874_ (.B(_3044_),
    .C(_3059_),
    .A(_3041_),
    .Y(_0500_));
 sg13g2_nor3_1 _3875_ (.A(_3050_),
    .B(_3051_),
    .C(net67),
    .Y(_0501_));
 sg13g2_nand3_1 _3876_ (.B(_0461_),
    .C(_0501_),
    .A(_3047_),
    .Y(_0502_));
 sg13g2_a21oi_1 _3877_ (.A1(_0499_),
    .A2(_0500_),
    .Y(_0503_),
    .B1(_0502_));
 sg13g2_a221oi_1 _3878_ (.B2(_0497_),
    .C1(_0503_),
    .B1(_0495_),
    .A1(_0466_),
    .Y(_0504_),
    .A2(_0494_));
 sg13g2_nor2_1 _3879_ (.A(_3039_),
    .B(_0504_),
    .Y(_0505_));
 sg13g2_and2_1 _3880_ (.A(_0485_),
    .B(_0505_),
    .X(_0047_));
 sg13g2_buf_2 _3881_ (.A(\Pong.datapath.NES_activity_Left[5] ),
    .X(_0506_));
 sg13g2_inv_2 _3882_ (.Y(_0507_),
    .A(_0506_));
 sg13g2_nand2_1 _3883_ (.Y(_0508_),
    .A(net186),
    .B(_0507_));
 sg13g2_nor3_1 _3884_ (.A(\Pong.datapath.old_NES_Left[2] ),
    .B(\Pong.datapath.NES_wire_Left[2] ),
    .C(_0508_),
    .Y(_0152_));
 sg13g2_nor3_1 _3885_ (.A(\Pong.datapath.old_NES_Left[3] ),
    .B(\Pong.datapath.NES_wire_Left[3] ),
    .C(_0508_),
    .Y(_0153_));
 sg13g2_nor3_1 _3886_ (.A(\Pong.datapath.old_NES_Left[4] ),
    .B(\Pong.datapath.NES_wire_Left[4] ),
    .C(_0508_),
    .Y(_0154_));
 sg13g2_nor3_1 _3887_ (.A(\Pong.datapath.old_NES_Left[5] ),
    .B(\Pong.datapath.NES_wire_Left[5] ),
    .C(_0508_),
    .Y(_0155_));
 sg13g2_inv_1 _3888_ (.Y(_0509_),
    .A(\Pong.datapath.NES_activity_Right[5] ));
 sg13g2_nand2_1 _3889_ (.Y(_0510_),
    .A(_2737_),
    .B(_0509_));
 sg13g2_nor3_1 _3890_ (.A(\Pong.datapath.old_NES_Right[2] ),
    .B(\Pong.datapath.NES_wire_Right[2] ),
    .C(_0510_),
    .Y(_0156_));
 sg13g2_nor3_1 _3891_ (.A(\Pong.datapath.old_NES_Right[3] ),
    .B(\Pong.datapath.NES_wire_Right[3] ),
    .C(_0510_),
    .Y(_0157_));
 sg13g2_nor3_1 _3892_ (.A(\Pong.datapath.old_NES_Right[4] ),
    .B(\Pong.datapath.NES_wire_Right[4] ),
    .C(_0510_),
    .Y(_0158_));
 sg13g2_nor3_1 _3893_ (.A(\Pong.datapath.old_NES_Right[5] ),
    .B(\Pong.datapath.NES_wire_Right[5] ),
    .C(_0510_),
    .Y(_0159_));
 sg13g2_nand2b_1 _3894_ (.Y(_0511_),
    .B(_2656_),
    .A_N(_2811_));
 sg13g2_buf_2 _3895_ (.A(_0511_),
    .X(_0512_));
 sg13g2_nand2b_1 _3896_ (.Y(_0513_),
    .B(_2780_),
    .A_N(_2779_));
 sg13g2_inv_1 _3897_ (.Y(_0514_),
    .A(_0119_));
 sg13g2_a21oi_1 _3898_ (.A1(\Pong.datapath.NES_counter_left.Q[7] ),
    .A2(_0513_),
    .Y(_0515_),
    .B1(_0514_));
 sg13g2_xnor2_1 _3899_ (.Y(_0516_),
    .A(_2781_),
    .B(_0515_));
 sg13g2_nor2_1 _3900_ (.A(_0512_),
    .B(_0516_),
    .Y(_0160_));
 sg13g2_nand2_1 _3901_ (.Y(_0517_),
    .A(_2781_),
    .B(_0515_));
 sg13g2_xor2_1 _3902_ (.B(_0517_),
    .A(\Pong.datapath.NES_counter_left.Q[1] ),
    .X(_0518_));
 sg13g2_nor2_1 _3903_ (.A(_0512_),
    .B(_0518_),
    .Y(_0161_));
 sg13g2_inv_1 _3904_ (.Y(_0519_),
    .A(\Pong.datapath.NES_counter_left.Q[2] ));
 sg13g2_nand3_1 _3905_ (.B(_2781_),
    .C(_0515_),
    .A(\Pong.datapath.NES_counter_left.Q[1] ),
    .Y(_0520_));
 sg13g2_xnor2_1 _3906_ (.Y(_0521_),
    .A(_0519_),
    .B(_0520_));
 sg13g2_nor2_1 _3907_ (.A(_0512_),
    .B(_0521_),
    .Y(_0162_));
 sg13g2_or2_1 _3908_ (.X(_0522_),
    .B(_0520_),
    .A(_0519_));
 sg13g2_nand2_1 _3909_ (.Y(_0523_),
    .A(_2785_),
    .B(_0522_));
 sg13g2_mux2_1 _3910_ (.A0(_0522_),
    .A1(_0523_),
    .S(\Pong.datapath.NES_counter_left.Q[3] ),
    .X(_0524_));
 sg13g2_nor2_1 _3911_ (.A(_0512_),
    .B(_0524_),
    .Y(_0163_));
 sg13g2_nor2_1 _3912_ (.A(_0519_),
    .B(_0520_),
    .Y(_0525_));
 sg13g2_nand2_1 _3913_ (.Y(_0526_),
    .A(\Pong.datapath.NES_counter_left.Q[3] ),
    .B(_0525_));
 sg13g2_inv_1 _3914_ (.Y(_0527_),
    .A(\Pong.datapath.NES_counter_left.Q[4] ));
 sg13g2_a221oi_1 _3915_ (.B2(_0527_),
    .C1(_0512_),
    .B1(_0526_),
    .A1(_2779_),
    .Y(_0164_),
    .A2(_0523_));
 sg13g2_o21ai_1 _3916_ (.B1(_0526_),
    .Y(_0528_),
    .A1(_2811_),
    .A2(_2785_));
 sg13g2_and3_1 _3917_ (.X(_0529_),
    .A(\Pong.datapath.NES_counter_left.Q[5] ),
    .B(\Pong.datapath.NES_counter_left.Q[4] ),
    .C(_0528_));
 sg13g2_buf_1 _3918_ (.A(_0529_),
    .X(_0530_));
 sg13g2_a21oi_1 _3919_ (.A1(_2779_),
    .A2(_0525_),
    .Y(_0531_),
    .B1(\Pong.datapath.NES_counter_left.Q[5] ));
 sg13g2_nor3_1 _3920_ (.A(_0512_),
    .B(_0530_),
    .C(_0531_),
    .Y(_0165_));
 sg13g2_xnor2_1 _3921_ (.Y(_0532_),
    .A(\Pong.datapath.NES_counter_left.Q[6] ),
    .B(_0530_));
 sg13g2_nor3_1 _3922_ (.A(net83),
    .B(_0512_),
    .C(_0532_),
    .Y(_0166_));
 sg13g2_a21oi_1 _3923_ (.A1(\Pong.datapath.NES_counter_left.Q[6] ),
    .A2(_0530_),
    .Y(_0533_),
    .B1(\Pong.datapath.NES_counter_left.Q[7] ));
 sg13g2_nor3_1 _3924_ (.A(net83),
    .B(_0512_),
    .C(_0533_),
    .Y(_0167_));
 sg13g2_nand2_1 _3925_ (.Y(_0534_),
    .A(_2656_),
    .B(_2856_));
 sg13g2_buf_2 _3926_ (.A(_0534_),
    .X(_0535_));
 sg13g2_nand2_1 _3927_ (.Y(_0536_),
    .A(_2640_),
    .B(_2641_));
 sg13g2_a21oi_1 _3928_ (.A1(_2643_),
    .A2(_0536_),
    .Y(_0537_),
    .B1(_2646_));
 sg13g2_buf_1 _3929_ (.A(_0127_),
    .X(_0538_));
 sg13g2_nor2b_1 _3930_ (.A(_0537_),
    .B_N(_0538_),
    .Y(_0539_));
 sg13g2_buf_2 _3931_ (.A(_0539_),
    .X(_0540_));
 sg13g2_xnor2_1 _3932_ (.Y(_0541_),
    .A(_2645_),
    .B(_0540_));
 sg13g2_nor2_1 _3933_ (.A(_0535_),
    .B(_0541_),
    .Y(_0168_));
 sg13g2_nand2_1 _3934_ (.Y(_0542_),
    .A(_2645_),
    .B(_0540_));
 sg13g2_xor2_1 _3935_ (.B(_0542_),
    .A(_2644_),
    .X(_0543_));
 sg13g2_nor2_1 _3936_ (.A(_0535_),
    .B(_0543_),
    .Y(_0169_));
 sg13g2_nand3_1 _3937_ (.B(_2645_),
    .C(_0540_),
    .A(_2644_),
    .Y(_0544_));
 sg13g2_xor2_1 _3938_ (.B(_0544_),
    .A(\Pong.datapath.NES_counter_right.Q[2] ),
    .X(_0545_));
 sg13g2_nor2_1 _3939_ (.A(_0535_),
    .B(_0545_),
    .Y(_0170_));
 sg13g2_nand3_1 _3940_ (.B(_2645_),
    .C(\Pong.datapath.NES_counter_right.Q[2] ),
    .A(_2644_),
    .Y(_0546_));
 sg13g2_mux2_1 _3941_ (.A0(_2649_),
    .A1(_0546_),
    .S(_0540_),
    .X(_0547_));
 sg13g2_nor2_1 _3942_ (.A(_2640_),
    .B(_0546_),
    .Y(_0548_));
 sg13g2_a22oi_1 _3943_ (.Y(_0549_),
    .B1(_0548_),
    .B2(_0540_),
    .A2(_0547_),
    .A1(_2640_));
 sg13g2_nor2_1 _3944_ (.A(_0535_),
    .B(_0549_),
    .Y(_0171_));
 sg13g2_inv_1 _3945_ (.Y(_0550_),
    .A(_2640_));
 sg13g2_nor2_1 _3946_ (.A(_0550_),
    .B(_0546_),
    .Y(_0551_));
 sg13g2_mux2_1 _3947_ (.A0(net93),
    .A1(_0551_),
    .S(_0540_),
    .X(_0552_));
 sg13g2_and2_1 _3948_ (.A(_0540_),
    .B(_0551_),
    .X(_0553_));
 sg13g2_inv_1 _3949_ (.Y(_0554_),
    .A(_0535_));
 sg13g2_o21ai_1 _3950_ (.B1(_0554_),
    .Y(_0555_),
    .A1(_2641_),
    .A2(_0553_));
 sg13g2_a21oi_1 _3951_ (.A1(_2641_),
    .A2(_0552_),
    .Y(_0172_),
    .B1(_0555_));
 sg13g2_nand2_1 _3952_ (.Y(_0556_),
    .A(_2641_),
    .B(_0553_));
 sg13g2_xor2_1 _3953_ (.B(_0556_),
    .A(_2642_),
    .X(_0557_));
 sg13g2_nor2_1 _3954_ (.A(_0535_),
    .B(_0557_),
    .Y(_0173_));
 sg13g2_nand4_1 _3955_ (.B(_2641_),
    .C(_0540_),
    .A(_2642_),
    .Y(_0558_),
    .D(_0551_));
 sg13g2_xor2_1 _3956_ (.B(_0558_),
    .A(\Pong.datapath.NES_counter_right.Q[6] ),
    .X(_0559_));
 sg13g2_nor2_1 _3957_ (.A(_0535_),
    .B(_0559_),
    .Y(_0174_));
 sg13g2_and2_1 _3958_ (.A(\Pong.datapath.NES_counter_right.Q[6] ),
    .B(_0538_),
    .X(_0560_));
 sg13g2_nand4_1 _3959_ (.B(_2641_),
    .C(_0551_),
    .A(_2642_),
    .Y(_0561_),
    .D(_0560_));
 sg13g2_and2_1 _3960_ (.A(_2646_),
    .B(_0561_),
    .X(_0562_));
 sg13g2_nor3_1 _3961_ (.A(_2651_),
    .B(_0535_),
    .C(_0562_),
    .Y(_0175_));
 sg13g2_nor2_1 _3962_ (.A(_2865_),
    .B(_2867_),
    .Y(_0563_));
 sg13g2_o21ai_1 _3963_ (.B1(_0056_),
    .Y(_0564_),
    .A1(_2870_),
    .A2(_0563_));
 sg13g2_nand2b_1 _3964_ (.Y(_0565_),
    .B(_0564_),
    .A_N(_2869_));
 sg13g2_a21oi_1 _3965_ (.A1(_2862_),
    .A2(_0565_),
    .Y(_0566_),
    .B1(_2871_));
 sg13g2_buf_1 _3966_ (.A(_0566_),
    .X(_0567_));
 sg13g2_nand2b_1 _3967_ (.Y(_0568_),
    .B(_0567_),
    .A_N(_2863_));
 sg13g2_inv_2 _3968_ (.Y(_0569_),
    .A(_0566_));
 sg13g2_nand2_1 _3969_ (.Y(_0570_),
    .A(_2863_),
    .B(_0569_));
 sg13g2_and3_1 _3970_ (.X(_0135_),
    .A(net188),
    .B(_0568_),
    .C(_0570_));
 sg13g2_nand2_1 _3971_ (.Y(_0571_),
    .A(net186),
    .B(_2874_));
 sg13g2_inv_1 _3972_ (.Y(_0572_),
    .A(\Pong.datapath.Ball_Clock.Q[9] ));
 sg13g2_and3_1 _3973_ (.X(_0573_),
    .A(\Pong.datapath.Ball_Clock.Q[1] ),
    .B(_2863_),
    .C(\Pong.datapath.Ball_Clock.Q[2] ));
 sg13g2_and2_1 _3974_ (.A(\Pong.datapath.Ball_Clock.Q[3] ),
    .B(_0573_),
    .X(_0574_));
 sg13g2_and2_1 _3975_ (.A(\Pong.datapath.Ball_Clock.Q[4] ),
    .B(_0574_),
    .X(_0575_));
 sg13g2_buf_1 _3976_ (.A(_0575_),
    .X(_0576_));
 sg13g2_nand3_1 _3977_ (.B(_2867_),
    .C(_0576_),
    .A(_2865_),
    .Y(_0577_));
 sg13g2_inv_1 _3978_ (.Y(_0578_),
    .A(_0577_));
 sg13g2_and2_1 _3979_ (.A(\Pong.datapath.Ball_Clock.Q[7] ),
    .B(_0578_),
    .X(_0579_));
 sg13g2_buf_1 _3980_ (.A(_0579_),
    .X(_0580_));
 sg13g2_nand3_1 _3981_ (.B(_0569_),
    .C(_0580_),
    .A(\Pong.datapath.Ball_Clock.Q[8] ),
    .Y(_0581_));
 sg13g2_buf_2 _3982_ (.A(_0581_),
    .X(_0582_));
 sg13g2_nor2_1 _3983_ (.A(_0572_),
    .B(_0582_),
    .Y(_0583_));
 sg13g2_xnor2_1 _3984_ (.Y(_0584_),
    .A(\Pong.datapath.Ball_Clock.Q[10] ),
    .B(_0583_));
 sg13g2_nor2_1 _3985_ (.A(_0571_),
    .B(_0584_),
    .Y(_0136_));
 sg13g2_nor2_1 _3986_ (.A(_2869_),
    .B(_0582_),
    .Y(_0585_));
 sg13g2_xnor2_1 _3987_ (.Y(_0586_),
    .A(\Pong.datapath.Ball_Clock.Q[11] ),
    .B(_0585_));
 sg13g2_nor2_1 _3988_ (.A(net109),
    .B(_0586_),
    .Y(_0137_));
 sg13g2_inv_1 _3989_ (.Y(_0587_),
    .A(\Pong.datapath.Ball_Clock.Q[11] ));
 sg13g2_nor3_1 _3990_ (.A(_0587_),
    .B(_2869_),
    .C(_0582_),
    .Y(_0588_));
 sg13g2_xnor2_1 _3991_ (.Y(_0589_),
    .A(\Pong.datapath.Ball_Clock.Q[12] ),
    .B(_0588_));
 sg13g2_nor2_1 _3992_ (.A(net109),
    .B(_0589_),
    .Y(_0138_));
 sg13g2_nand4_1 _3993_ (.B(\Pong.datapath.Ball_Clock.Q[11] ),
    .C(\Pong.datapath.Ball_Clock.Q[10] ),
    .A(\Pong.datapath.Ball_Clock.Q[12] ),
    .Y(_0590_),
    .D(\Pong.datapath.Ball_Clock.Q[9] ));
 sg13g2_nor2_1 _3994_ (.A(_0582_),
    .B(_0590_),
    .Y(_0591_));
 sg13g2_xnor2_1 _3995_ (.Y(_0592_),
    .A(\Pong.datapath.Ball_Clock.Q[13] ),
    .B(_0591_));
 sg13g2_nor2_1 _3996_ (.A(net109),
    .B(_0592_),
    .Y(_0139_));
 sg13g2_inv_1 _3997_ (.Y(_0593_),
    .A(\Pong.datapath.Ball_Clock.Q[13] ));
 sg13g2_or2_1 _3998_ (.X(_0594_),
    .B(_0590_),
    .A(_0593_));
 sg13g2_nor2_1 _3999_ (.A(_0582_),
    .B(_0594_),
    .Y(_0595_));
 sg13g2_xnor2_1 _4000_ (.Y(_0596_),
    .A(\Pong.datapath.Ball_Clock.Q[14] ),
    .B(_0595_));
 sg13g2_nor2_1 _4001_ (.A(net109),
    .B(_0596_),
    .Y(_0140_));
 sg13g2_inv_1 _4002_ (.Y(_0597_),
    .A(\Pong.datapath.Ball_Clock.Q[14] ));
 sg13g2_nand2_1 _4003_ (.Y(_0598_),
    .A(\Pong.datapath.Ball_Clock.Q[8] ),
    .B(_0580_));
 sg13g2_nor3_1 _4004_ (.A(_0597_),
    .B(_0598_),
    .C(_0594_),
    .Y(_0599_));
 sg13g2_xnor2_1 _4005_ (.Y(_0600_),
    .A(\Pong.datapath.Ball_Clock.Q[15] ),
    .B(_0599_));
 sg13g2_a21oi_1 _4006_ (.A1(_0569_),
    .A2(_0600_),
    .Y(_0141_),
    .B1(_0571_));
 sg13g2_a21oi_1 _4007_ (.A1(\Pong.datapath.Ball_Clock.Q[15] ),
    .A2(_0599_),
    .Y(_0601_),
    .B1(\Pong.datapath.Ball_Clock.Q[16] ));
 sg13g2_nor2_1 _4008_ (.A(_0571_),
    .B(_0601_),
    .Y(_0142_));
 sg13g2_buf_1 _4009_ (.A(net157),
    .X(_0602_));
 sg13g2_xor2_1 _4010_ (.B(_0570_),
    .A(\Pong.datapath.Ball_Clock.Q[1] ),
    .X(_0603_));
 sg13g2_nor2_1 _4011_ (.A(net98),
    .B(_0603_),
    .Y(_0143_));
 sg13g2_nand3_1 _4012_ (.B(_2863_),
    .C(_0569_),
    .A(\Pong.datapath.Ball_Clock.Q[1] ),
    .Y(_0604_));
 sg13g2_xor2_1 _4013_ (.B(_0604_),
    .A(\Pong.datapath.Ball_Clock.Q[2] ),
    .X(_0605_));
 sg13g2_nor2_1 _4014_ (.A(net98),
    .B(_0605_),
    .Y(_0144_));
 sg13g2_nand2_2 _4015_ (.Y(_0606_),
    .A(_2874_),
    .B(net79));
 sg13g2_o21ai_1 _4016_ (.B1(_0606_),
    .Y(_0607_),
    .A1(net79),
    .A2(_0573_));
 sg13g2_nor2b_1 _4017_ (.A(\Pong.datapath.Ball_Clock.Q[3] ),
    .B_N(_0573_),
    .Y(_0608_));
 sg13g2_a22oi_1 _4018_ (.Y(_0609_),
    .B1(_0608_),
    .B2(_0569_),
    .A2(_0607_),
    .A1(\Pong.datapath.Ball_Clock.Q[3] ));
 sg13g2_nor2_1 _4019_ (.A(net98),
    .B(_0609_),
    .Y(_0145_));
 sg13g2_o21ai_1 _4020_ (.B1(_0606_),
    .Y(_0610_),
    .A1(net79),
    .A2(_0574_));
 sg13g2_nor2b_1 _4021_ (.A(\Pong.datapath.Ball_Clock.Q[4] ),
    .B_N(_0574_),
    .Y(_0611_));
 sg13g2_a22oi_1 _4022_ (.Y(_0612_),
    .B1(_0611_),
    .B2(_0569_),
    .A2(_0610_),
    .A1(\Pong.datapath.Ball_Clock.Q[4] ));
 sg13g2_nor2_1 _4023_ (.A(net98),
    .B(_0612_),
    .Y(_0146_));
 sg13g2_o21ai_1 _4024_ (.B1(_0606_),
    .Y(_0613_),
    .A1(net79),
    .A2(_0576_));
 sg13g2_inv_1 _4025_ (.Y(_0614_),
    .A(_0576_));
 sg13g2_nor3_1 _4026_ (.A(_2865_),
    .B(net79),
    .C(_0614_),
    .Y(_0615_));
 sg13g2_a21oi_1 _4027_ (.A1(_2865_),
    .A2(_0613_),
    .Y(_0616_),
    .B1(_0615_));
 sg13g2_nor2_1 _4028_ (.A(net98),
    .B(_0616_),
    .Y(_0147_));
 sg13g2_nor2_1 _4029_ (.A(_2866_),
    .B(_0614_),
    .Y(_0617_));
 sg13g2_o21ai_1 _4030_ (.B1(_0606_),
    .Y(_0618_),
    .A1(net79),
    .A2(_0617_));
 sg13g2_nor4_1 _4031_ (.A(_2866_),
    .B(_2867_),
    .C(net79),
    .D(_0614_),
    .Y(_0619_));
 sg13g2_a21oi_1 _4032_ (.A1(_2867_),
    .A2(_0618_),
    .Y(_0620_),
    .B1(_0619_));
 sg13g2_nor2_1 _4033_ (.A(net98),
    .B(_0620_),
    .Y(_0148_));
 sg13g2_o21ai_1 _4034_ (.B1(_0606_),
    .Y(_0621_),
    .A1(_0567_),
    .A2(_0578_));
 sg13g2_nor2_1 _4035_ (.A(\Pong.datapath.Ball_Clock.Q[7] ),
    .B(_0577_),
    .Y(_0622_));
 sg13g2_a22oi_1 _4036_ (.Y(_0623_),
    .B1(_0622_),
    .B2(_0569_),
    .A2(_0621_),
    .A1(\Pong.datapath.Ball_Clock.Q[7] ));
 sg13g2_nor2_1 _4037_ (.A(net98),
    .B(_0623_),
    .Y(_0149_));
 sg13g2_nand2_1 _4038_ (.Y(_0624_),
    .A(\Pong.datapath.Ball_Clock.Q[8] ),
    .B(net79));
 sg13g2_xnor2_1 _4039_ (.Y(_0625_),
    .A(_0056_),
    .B(_0580_));
 sg13g2_nand2_1 _4040_ (.Y(_0626_),
    .A(_0569_),
    .B(_0625_));
 sg13g2_a21oi_1 _4041_ (.A1(_0624_),
    .A2(_0626_),
    .Y(_0150_),
    .B1(net106));
 sg13g2_xnor2_1 _4042_ (.Y(_0627_),
    .A(_0572_),
    .B(_0582_));
 sg13g2_nor2_1 _4043_ (.A(_0571_),
    .B(_0627_),
    .Y(_0151_));
 sg13g2_buf_1 _4044_ (.A(net186),
    .X(_0628_));
 sg13g2_nand2_1 _4045_ (.Y(_0629_),
    .A(_2825_),
    .B(_2826_));
 sg13g2_a21oi_1 _4046_ (.A1(_0118_),
    .A2(_2822_),
    .Y(_0630_),
    .B1(_0629_));
 sg13g2_o21ai_1 _4047_ (.B1(_2830_),
    .Y(_0631_),
    .A1(_2824_),
    .A2(_0630_));
 sg13g2_nand2_1 _4048_ (.Y(_0632_),
    .A(\Pong.datapath.NES_delay_counter_left.Q[17] ),
    .B(\Pong.datapath.NES_delay_counter_left.Q[18] ));
 sg13g2_a21o_1 _4049_ (.A2(_0631_),
    .A1(_2829_),
    .B1(_0632_),
    .X(_0633_));
 sg13g2_nand2_1 _4050_ (.Y(_0634_),
    .A(_2811_),
    .B(_0633_));
 sg13g2_buf_1 _4051_ (.A(_0634_),
    .X(_0635_));
 sg13g2_nand3_1 _4052_ (.B(_2835_),
    .C(net44),
    .A(_2813_),
    .Y(_0636_));
 sg13g2_o21ai_1 _4053_ (.B1(_0636_),
    .Y(_0637_),
    .A1(_2813_),
    .A2(net44));
 sg13g2_and2_1 _4054_ (.A(net139),
    .B(_0637_),
    .X(_0176_));
 sg13g2_and2_1 _4055_ (.A(_2815_),
    .B(_2818_),
    .X(_0638_));
 sg13g2_buf_1 _4056_ (.A(_0638_),
    .X(_0639_));
 sg13g2_nand2_1 _4057_ (.Y(_0640_),
    .A(_0639_),
    .B(_2821_));
 sg13g2_nor2_1 _4058_ (.A(_2812_),
    .B(_0640_),
    .Y(_0641_));
 sg13g2_and2_1 _4059_ (.A(_2826_),
    .B(_0641_),
    .X(_0642_));
 sg13g2_and2_1 _4060_ (.A(_2811_),
    .B(_0633_),
    .X(_0643_));
 sg13g2_buf_1 _4061_ (.A(_0643_),
    .X(_0644_));
 sg13g2_nand2_1 _4062_ (.Y(_0645_),
    .A(_2656_),
    .B(_0644_));
 sg13g2_buf_1 _4063_ (.A(_0645_),
    .X(_0646_));
 sg13g2_nor3_1 _4064_ (.A(_2827_),
    .B(_0117_),
    .C(_2824_),
    .Y(_0647_));
 sg13g2_nand4_1 _4065_ (.B(_2826_),
    .C(_0647_),
    .A(_2825_),
    .Y(_0648_),
    .D(_2831_));
 sg13g2_nor2_1 _4066_ (.A(_2822_),
    .B(_0648_),
    .Y(_0649_));
 sg13g2_o21ai_1 _4067_ (.B1(_2811_),
    .Y(_0650_),
    .A1(_0649_),
    .A2(_0633_));
 sg13g2_nand2_1 _4068_ (.Y(_0651_),
    .A(_2656_),
    .B(_0650_));
 sg13g2_buf_1 _4069_ (.A(_0651_),
    .X(_0652_));
 sg13g2_o21ai_1 _4070_ (.B1(net31),
    .Y(_0653_),
    .A1(_0642_),
    .A2(net20));
 sg13g2_inv_1 _4071_ (.Y(_0654_),
    .A(_0642_));
 sg13g2_nor3_1 _4072_ (.A(_2825_),
    .B(_0654_),
    .C(net20),
    .Y(_0655_));
 sg13g2_a21o_1 _4073_ (.A2(_0653_),
    .A1(_2825_),
    .B1(_0655_),
    .X(_0177_));
 sg13g2_buf_1 _4074_ (.A(_0644_),
    .X(_0656_));
 sg13g2_nand4_1 _4075_ (.B(_2815_),
    .C(_2818_),
    .A(\Pong.datapath.NES_delay_counter_left.Q[8] ),
    .Y(_0657_),
    .D(_2821_));
 sg13g2_nor2_1 _4076_ (.A(_0629_),
    .B(_0657_),
    .Y(_0658_));
 sg13g2_nand2_1 _4077_ (.Y(_0659_),
    .A(net30),
    .B(_0658_));
 sg13g2_xor2_1 _4078_ (.B(_0659_),
    .A(\Pong.datapath.NES_delay_counter_left.Q[11] ),
    .X(_0660_));
 sg13g2_nor2_1 _4079_ (.A(_0602_),
    .B(_0660_),
    .Y(_0178_));
 sg13g2_and3_1 _4080_ (.X(_0661_),
    .A(\Pong.datapath.NES_delay_counter_left.Q[11] ),
    .B(_2825_),
    .C(_0642_));
 sg13g2_nand3_1 _4081_ (.B(net30),
    .C(_0661_),
    .A(net186),
    .Y(_0662_));
 sg13g2_o21ai_1 _4082_ (.B1(net31),
    .Y(_0663_),
    .A1(net20),
    .A2(_0661_));
 sg13g2_nand2_1 _4083_ (.Y(_0664_),
    .A(\Pong.datapath.NES_delay_counter_left.Q[12] ),
    .B(_0663_));
 sg13g2_o21ai_1 _4084_ (.B1(_0664_),
    .Y(_0179_),
    .A1(\Pong.datapath.NES_delay_counter_left.Q[12] ),
    .A2(_0662_));
 sg13g2_and3_1 _4085_ (.X(_0665_),
    .A(\Pong.datapath.NES_delay_counter_left.Q[12] ),
    .B(\Pong.datapath.NES_delay_counter_left.Q[11] ),
    .C(_0658_));
 sg13g2_buf_1 _4086_ (.A(_0665_),
    .X(_0666_));
 sg13g2_nand3_1 _4087_ (.B(net30),
    .C(_0666_),
    .A(net186),
    .Y(_0667_));
 sg13g2_o21ai_1 _4088_ (.B1(net31),
    .Y(_0668_),
    .A1(_0645_),
    .A2(_0666_));
 sg13g2_nand2_1 _4089_ (.Y(_0669_),
    .A(\Pong.datapath.NES_delay_counter_left.Q[13] ),
    .B(_0668_));
 sg13g2_o21ai_1 _4090_ (.B1(_0669_),
    .Y(_0180_),
    .A1(\Pong.datapath.NES_delay_counter_left.Q[13] ),
    .A2(_0667_));
 sg13g2_and2_1 _4091_ (.A(\Pong.datapath.NES_delay_counter_left.Q[13] ),
    .B(_0666_),
    .X(_0670_));
 sg13g2_nand3_1 _4092_ (.B(net30),
    .C(_0670_),
    .A(net186),
    .Y(_0671_));
 sg13g2_o21ai_1 _4093_ (.B1(net31),
    .Y(_0672_),
    .A1(_0645_),
    .A2(_0670_));
 sg13g2_nand2_1 _4094_ (.Y(_0673_),
    .A(\Pong.datapath.NES_delay_counter_left.Q[14] ),
    .B(_0672_));
 sg13g2_o21ai_1 _4095_ (.B1(_0673_),
    .Y(_0181_),
    .A1(\Pong.datapath.NES_delay_counter_left.Q[14] ),
    .A2(_0671_));
 sg13g2_nand3_1 _4096_ (.B(_0644_),
    .C(_0666_),
    .A(_2830_),
    .Y(_0674_));
 sg13g2_xor2_1 _4097_ (.B(_0674_),
    .A(\Pong.datapath.NES_delay_counter_left.Q[15] ),
    .X(_0675_));
 sg13g2_nor2_1 _4098_ (.A(_0602_),
    .B(_0675_),
    .Y(_0182_));
 sg13g2_and3_1 _4099_ (.X(_0676_),
    .A(\Pong.datapath.NES_delay_counter_left.Q[15] ),
    .B(\Pong.datapath.NES_delay_counter_left.Q[14] ),
    .C(_0670_));
 sg13g2_buf_1 _4100_ (.A(_0676_),
    .X(_0677_));
 sg13g2_nand2b_1 _4101_ (.Y(_0678_),
    .B(_0677_),
    .A_N(\Pong.datapath.NES_delay_counter_left.Q[16] ));
 sg13g2_o21ai_1 _4102_ (.B1(net31),
    .Y(_0679_),
    .A1(_0645_),
    .A2(_0677_));
 sg13g2_nand2_1 _4103_ (.Y(_0680_),
    .A(\Pong.datapath.NES_delay_counter_left.Q[16] ),
    .B(_0679_));
 sg13g2_o21ai_1 _4104_ (.B1(_0680_),
    .Y(_0183_),
    .A1(net20),
    .A2(_0678_));
 sg13g2_and2_1 _4105_ (.A(\Pong.datapath.NES_delay_counter_left.Q[16] ),
    .B(_0677_),
    .X(_0681_));
 sg13g2_nor3_1 _4106_ (.A(_2827_),
    .B(_0634_),
    .C(_0681_),
    .Y(_0682_));
 sg13g2_and3_1 _4107_ (.X(_0683_),
    .A(_2827_),
    .B(_2811_),
    .C(_0681_));
 sg13g2_o21ai_1 _4108_ (.B1(net188),
    .Y(_0684_),
    .A1(_0682_),
    .A2(_0683_));
 sg13g2_o21ai_1 _4109_ (.B1(_0684_),
    .Y(_0184_),
    .A1(_2827_),
    .A2(_0652_));
 sg13g2_nand2_1 _4110_ (.Y(_0685_),
    .A(\Pong.datapath.NES_delay_counter_left.Q[17] ),
    .B(_0681_));
 sg13g2_xnor2_1 _4111_ (.Y(_0686_),
    .A(_0117_),
    .B(_0685_));
 sg13g2_nand4_1 _4112_ (.B(\Pong.datapath.NES_delay_counter_left.Q[18] ),
    .C(_2835_),
    .A(net188),
    .Y(_0687_),
    .D(net44));
 sg13g2_o21ai_1 _4113_ (.B1(_0687_),
    .Y(_0185_),
    .A1(net20),
    .A2(_0686_));
 sg13g2_nand3_1 _4114_ (.B(_2835_),
    .C(_0635_),
    .A(\Pong.datapath.NES_delay_counter_left.Q[1] ),
    .Y(_0688_));
 sg13g2_xor2_1 _4115_ (.B(_2813_),
    .A(\Pong.datapath.NES_delay_counter_left.Q[1] ),
    .X(_0689_));
 sg13g2_nand2_1 _4116_ (.Y(_0690_),
    .A(_0656_),
    .B(_0689_));
 sg13g2_a21oi_1 _4117_ (.A1(_0688_),
    .A2(_0690_),
    .Y(_0186_),
    .B1(net106));
 sg13g2_nand3_1 _4118_ (.B(_2835_),
    .C(_0635_),
    .A(\Pong.datapath.NES_delay_counter_left.Q[2] ),
    .Y(_0691_));
 sg13g2_nand2_1 _4119_ (.Y(_0692_),
    .A(\Pong.datapath.NES_delay_counter_left.Q[1] ),
    .B(_2813_));
 sg13g2_xnor2_1 _4120_ (.Y(_0693_),
    .A(\Pong.datapath.NES_delay_counter_left.Q[2] ),
    .B(_0692_));
 sg13g2_nand2_1 _4121_ (.Y(_0694_),
    .A(_0656_),
    .B(_0693_));
 sg13g2_buf_1 _4122_ (.A(net157),
    .X(_0695_));
 sg13g2_a21oi_1 _4123_ (.A1(_0691_),
    .A2(_0694_),
    .Y(_0187_),
    .B1(net97));
 sg13g2_nand3_1 _4124_ (.B(_2835_),
    .C(net44),
    .A(_2816_),
    .Y(_0696_));
 sg13g2_xor2_1 _4125_ (.B(_2815_),
    .A(_2816_),
    .X(_0697_));
 sg13g2_nand2_1 _4126_ (.Y(_0698_),
    .A(net30),
    .B(_0697_));
 sg13g2_a21oi_1 _4127_ (.A1(_0696_),
    .A2(_0698_),
    .Y(_0188_),
    .B1(net97));
 sg13g2_nand3_1 _4128_ (.B(_2835_),
    .C(net44),
    .A(\Pong.datapath.NES_delay_counter_left.Q[4] ),
    .Y(_0699_));
 sg13g2_nand2_1 _4129_ (.Y(_0700_),
    .A(_2816_),
    .B(_2815_));
 sg13g2_xnor2_1 _4130_ (.Y(_0701_),
    .A(\Pong.datapath.NES_delay_counter_left.Q[4] ),
    .B(_0700_));
 sg13g2_nand2_1 _4131_ (.Y(_0702_),
    .A(net30),
    .B(_0701_));
 sg13g2_a21oi_1 _4132_ (.A1(_0699_),
    .A2(_0702_),
    .Y(_0189_),
    .B1(net97));
 sg13g2_nand3_1 _4133_ (.B(_2816_),
    .C(_2815_),
    .A(\Pong.datapath.NES_delay_counter_left.Q[4] ),
    .Y(_0703_));
 sg13g2_xnor2_1 _4134_ (.Y(_0704_),
    .A(\Pong.datapath.NES_delay_counter_left.Q[5] ),
    .B(_0703_));
 sg13g2_nand2_1 _4135_ (.Y(_0705_),
    .A(net30),
    .B(_0704_));
 sg13g2_nand3_1 _4136_ (.B(_2835_),
    .C(net44),
    .A(\Pong.datapath.NES_delay_counter_left.Q[5] ),
    .Y(_0706_));
 sg13g2_a21oi_1 _4137_ (.A1(_0705_),
    .A2(_0706_),
    .Y(_0190_),
    .B1(net97));
 sg13g2_nand3_1 _4138_ (.B(_0639_),
    .C(net30),
    .A(net186),
    .Y(_0707_));
 sg13g2_o21ai_1 _4139_ (.B1(net31),
    .Y(_0708_),
    .A1(_0639_),
    .A2(net20));
 sg13g2_nand2_1 _4140_ (.Y(_0709_),
    .A(_2819_),
    .B(_0708_));
 sg13g2_o21ai_1 _4141_ (.B1(_0709_),
    .Y(_0191_),
    .A1(_2819_),
    .A2(_0707_));
 sg13g2_and2_1 _4142_ (.A(_2819_),
    .B(_0639_),
    .X(_0710_));
 sg13g2_o21ai_1 _4143_ (.B1(net31),
    .Y(_0711_),
    .A1(_0710_),
    .A2(net20));
 sg13g2_nand2_1 _4144_ (.Y(_0712_),
    .A(_2819_),
    .B(_0639_));
 sg13g2_nor3_1 _4145_ (.A(\Pong.datapath.NES_delay_counter_left.Q[7] ),
    .B(_0712_),
    .C(net20),
    .Y(_0713_));
 sg13g2_a21o_1 _4146_ (.A2(_0711_),
    .A1(\Pong.datapath.NES_delay_counter_left.Q[7] ),
    .B1(_0713_),
    .X(_0192_));
 sg13g2_xnor2_1 _4147_ (.Y(_0714_),
    .A(_0118_),
    .B(_0640_));
 sg13g2_nor2_1 _4148_ (.A(net44),
    .B(_0714_),
    .Y(_0715_));
 sg13g2_a21oi_1 _4149_ (.A1(\Pong.datapath.NES_delay_counter_left.Q[8] ),
    .A2(net44),
    .Y(_0716_),
    .B1(_0715_));
 sg13g2_nor2_1 _4150_ (.A(net98),
    .B(_0716_),
    .Y(_0193_));
 sg13g2_o21ai_1 _4151_ (.B1(net31),
    .Y(_0717_),
    .A1(_0641_),
    .A2(_0646_));
 sg13g2_nor3_1 _4152_ (.A(_2826_),
    .B(_0657_),
    .C(_0646_),
    .Y(_0718_));
 sg13g2_a21o_1 _4153_ (.A2(_0717_),
    .A1(_2826_),
    .B1(_0718_),
    .X(_0194_));
 sg13g2_nand2_1 _4154_ (.Y(_0719_),
    .A(_2690_),
    .B(_2691_));
 sg13g2_o21ai_1 _4155_ (.B1(_0116_),
    .Y(_0720_),
    .A1(\Pong.datapath.NES_delay_counter_right.Q[8] ),
    .A2(_2682_));
 sg13g2_a21oi_1 _4156_ (.A1(_2694_),
    .A2(_0720_),
    .Y(_0721_),
    .B1(_2689_));
 sg13g2_o21ai_1 _4157_ (.B1(_2692_),
    .Y(_0722_),
    .A1(_0719_),
    .A2(_0721_));
 sg13g2_and2_1 _4158_ (.A(_2685_),
    .B(\Pong.datapath.NES_delay_counter_right.Q[18] ),
    .X(_0723_));
 sg13g2_a21o_1 _4159_ (.A2(_0723_),
    .A1(_0722_),
    .B1(_2856_),
    .X(_0724_));
 sg13g2_buf_1 _4160_ (.A(_0724_),
    .X(_0725_));
 sg13g2_buf_1 _4161_ (.A(net29),
    .X(_0726_));
 sg13g2_nand3_1 _4162_ (.B(net62),
    .C(net19),
    .A(_2675_),
    .Y(_0727_));
 sg13g2_buf_1 _4163_ (.A(net29),
    .X(_0728_));
 sg13g2_or2_1 _4164_ (.X(_0729_),
    .B(net18),
    .A(_2675_));
 sg13g2_a21oi_1 _4165_ (.A1(_0727_),
    .A2(_0729_),
    .Y(_0195_),
    .B1(net97));
 sg13g2_buf_1 _4166_ (.A(_2663_),
    .X(_0730_));
 sg13g2_nor2_1 _4167_ (.A(_2683_),
    .B(_2682_),
    .Y(_0731_));
 sg13g2_nand2_1 _4168_ (.Y(_0732_),
    .A(_2693_),
    .B(_0731_));
 sg13g2_mux2_1 _4169_ (.A0(_0732_),
    .A1(_2697_),
    .S(net29),
    .X(_0733_));
 sg13g2_buf_1 _4170_ (.A(net29),
    .X(_0734_));
 sg13g2_nor3_1 _4171_ (.A(\Pong.datapath.NES_delay_counter_right.Q[10] ),
    .B(net17),
    .C(_0732_),
    .Y(_0735_));
 sg13g2_a21oi_1 _4172_ (.A1(\Pong.datapath.NES_delay_counter_right.Q[10] ),
    .A2(_0733_),
    .Y(_0736_),
    .B1(_0735_));
 sg13g2_nor2_1 _4173_ (.A(net96),
    .B(_0736_),
    .Y(_0196_));
 sg13g2_nand2_1 _4174_ (.Y(_0737_),
    .A(\Pong.datapath.NES_delay_counter_right.Q[10] ),
    .B(_2693_));
 sg13g2_nor3_2 _4175_ (.A(_2683_),
    .B(_2682_),
    .C(_0737_),
    .Y(_0738_));
 sg13g2_nand2_1 _4176_ (.Y(_0739_),
    .A(_2697_),
    .B(net29));
 sg13g2_buf_2 _4177_ (.A(_0739_),
    .X(_0740_));
 sg13g2_o21ai_1 _4178_ (.B1(_0740_),
    .Y(_0741_),
    .A1(_0734_),
    .A2(_0738_));
 sg13g2_inv_1 _4179_ (.Y(_0742_),
    .A(_0738_));
 sg13g2_nor3_1 _4180_ (.A(_2688_),
    .B(net17),
    .C(_0742_),
    .Y(_0743_));
 sg13g2_a21oi_1 _4181_ (.A1(_2688_),
    .A2(_0741_),
    .Y(_0744_),
    .B1(_0743_));
 sg13g2_nor2_1 _4182_ (.A(net96),
    .B(_0744_),
    .Y(_0197_));
 sg13g2_and2_1 _4183_ (.A(_2688_),
    .B(_0738_),
    .X(_0745_));
 sg13g2_buf_1 _4184_ (.A(_0745_),
    .X(_0746_));
 sg13g2_o21ai_1 _4185_ (.B1(_0740_),
    .Y(_0747_),
    .A1(net17),
    .A2(_0746_));
 sg13g2_inv_1 _4186_ (.Y(_0748_),
    .A(_0746_));
 sg13g2_nor3_1 _4187_ (.A(_2687_),
    .B(net17),
    .C(_0748_),
    .Y(_0749_));
 sg13g2_a21oi_1 _4188_ (.A1(_2687_),
    .A2(_0747_),
    .Y(_0750_),
    .B1(_0749_));
 sg13g2_nor2_1 _4189_ (.A(_0730_),
    .B(_0750_),
    .Y(_0198_));
 sg13g2_and3_1 _4190_ (.X(_0751_),
    .A(_2687_),
    .B(_2688_),
    .C(_0738_));
 sg13g2_buf_1 _4191_ (.A(_0751_),
    .X(_0752_));
 sg13g2_o21ai_1 _4192_ (.B1(_0740_),
    .Y(_0753_),
    .A1(_0725_),
    .A2(_0752_));
 sg13g2_nand2_1 _4193_ (.Y(_0754_),
    .A(_2687_),
    .B(_0746_));
 sg13g2_nor3_1 _4194_ (.A(_2691_),
    .B(_0734_),
    .C(_0754_),
    .Y(_0755_));
 sg13g2_a21oi_1 _4195_ (.A1(_2691_),
    .A2(_0753_),
    .Y(_0756_),
    .B1(_0755_));
 sg13g2_nor2_1 _4196_ (.A(net96),
    .B(_0756_),
    .Y(_0199_));
 sg13g2_nand2_1 _4197_ (.Y(_0757_),
    .A(_2691_),
    .B(_0752_));
 sg13g2_inv_1 _4198_ (.Y(_0758_),
    .A(_0757_));
 sg13g2_o21ai_1 _4199_ (.B1(_0740_),
    .Y(_0759_),
    .A1(_0725_),
    .A2(_0758_));
 sg13g2_nor3_1 _4200_ (.A(_2690_),
    .B(net17),
    .C(_0757_),
    .Y(_0760_));
 sg13g2_a21oi_1 _4201_ (.A1(_2690_),
    .A2(_0759_),
    .Y(_0761_),
    .B1(_0760_));
 sg13g2_nor2_1 _4202_ (.A(net96),
    .B(_0761_),
    .Y(_0200_));
 sg13g2_nor3_1 _4203_ (.A(_0719_),
    .B(net29),
    .C(_0754_),
    .Y(_0762_));
 sg13g2_xnor2_1 _4204_ (.Y(_0763_),
    .A(\Pong.datapath.NES_delay_counter_right.Q[15] ),
    .B(_0762_));
 sg13g2_nor2_1 _4205_ (.A(net96),
    .B(_0763_),
    .Y(_0201_));
 sg13g2_and4_1 _4206_ (.A(\Pong.datapath.NES_delay_counter_right.Q[15] ),
    .B(_2690_),
    .C(_2691_),
    .D(_0752_),
    .X(_0764_));
 sg13g2_buf_8 _4207_ (.A(_0764_),
    .X(_0765_));
 sg13g2_o21ai_1 _4208_ (.B1(_0740_),
    .Y(_0766_),
    .A1(net29),
    .A2(_0765_));
 sg13g2_nand2b_1 _4209_ (.Y(_0767_),
    .B(_0765_),
    .A_N(\Pong.datapath.NES_delay_counter_right.Q[16] ));
 sg13g2_nor2_1 _4210_ (.A(net18),
    .B(_0767_),
    .Y(_0768_));
 sg13g2_a21oi_1 _4211_ (.A1(\Pong.datapath.NES_delay_counter_right.Q[16] ),
    .A2(_0766_),
    .Y(_0769_),
    .B1(_0768_));
 sg13g2_nor2_1 _4212_ (.A(net96),
    .B(_0769_),
    .Y(_0202_));
 sg13g2_and2_1 _4213_ (.A(\Pong.datapath.NES_delay_counter_right.Q[16] ),
    .B(_0765_),
    .X(_0770_));
 sg13g2_buf_8 _4214_ (.A(_0770_),
    .X(_0771_));
 sg13g2_o21ai_1 _4215_ (.B1(_0740_),
    .Y(_0772_),
    .A1(net29),
    .A2(_0771_));
 sg13g2_nor2_1 _4216_ (.A(_2685_),
    .B(_2856_),
    .Y(_0773_));
 sg13g2_a22oi_1 _4217_ (.Y(_0774_),
    .B1(_0773_),
    .B2(_0771_),
    .A2(_0772_),
    .A1(_2685_));
 sg13g2_nor2_1 _4218_ (.A(net96),
    .B(_0774_),
    .Y(_0203_));
 sg13g2_nand2_1 _4219_ (.Y(_0775_),
    .A(_2685_),
    .B(_0771_));
 sg13g2_xnor2_1 _4220_ (.Y(_0776_),
    .A(_0110_),
    .B(_0775_));
 sg13g2_nand3_1 _4221_ (.B(_2698_),
    .C(net17),
    .A(\Pong.datapath.NES_delay_counter_right.Q[18] ),
    .Y(_0777_));
 sg13g2_o21ai_1 _4222_ (.B1(_0777_),
    .Y(_0778_),
    .A1(net18),
    .A2(_0776_));
 sg13g2_and2_1 _4223_ (.A(net139),
    .B(_0778_),
    .X(_0204_));
 sg13g2_nand3_1 _4224_ (.B(net62),
    .C(net19),
    .A(\Pong.datapath.NES_delay_counter_right.Q[1] ),
    .Y(_0779_));
 sg13g2_xor2_1 _4225_ (.B(_2675_),
    .A(\Pong.datapath.NES_delay_counter_right.Q[1] ),
    .X(_0780_));
 sg13g2_nand2b_1 _4226_ (.Y(_0781_),
    .B(_0780_),
    .A_N(net19));
 sg13g2_a21oi_1 _4227_ (.A1(_0779_),
    .A2(_0781_),
    .Y(_0205_),
    .B1(net97));
 sg13g2_nand3_1 _4228_ (.B(net62),
    .C(net19),
    .A(\Pong.datapath.NES_delay_counter_right.Q[2] ),
    .Y(_0782_));
 sg13g2_nand2_1 _4229_ (.Y(_0783_),
    .A(\Pong.datapath.NES_delay_counter_right.Q[1] ),
    .B(_2675_));
 sg13g2_xnor2_1 _4230_ (.Y(_0784_),
    .A(\Pong.datapath.NES_delay_counter_right.Q[2] ),
    .B(_0783_));
 sg13g2_nand2b_1 _4231_ (.Y(_0785_),
    .B(_0784_),
    .A_N(net18));
 sg13g2_a21oi_1 _4232_ (.A1(_0782_),
    .A2(_0785_),
    .Y(_0206_),
    .B1(net97));
 sg13g2_nand3_1 _4233_ (.B(net62),
    .C(net19),
    .A(_2678_),
    .Y(_0786_));
 sg13g2_xor2_1 _4234_ (.B(_2677_),
    .A(_2678_),
    .X(_0787_));
 sg13g2_nand2b_1 _4235_ (.Y(_0788_),
    .B(_0787_),
    .A_N(net18));
 sg13g2_a21oi_1 _4236_ (.A1(_0786_),
    .A2(_0788_),
    .Y(_0207_),
    .B1(net97));
 sg13g2_nand3_1 _4237_ (.B(net62),
    .C(net19),
    .A(\Pong.datapath.NES_delay_counter_right.Q[4] ),
    .Y(_0789_));
 sg13g2_nand2_1 _4238_ (.Y(_0790_),
    .A(_2678_),
    .B(_2677_));
 sg13g2_xnor2_1 _4239_ (.Y(_0791_),
    .A(\Pong.datapath.NES_delay_counter_right.Q[4] ),
    .B(_0790_));
 sg13g2_nand2b_1 _4240_ (.Y(_0792_),
    .B(_0791_),
    .A_N(net18));
 sg13g2_a21oi_1 _4241_ (.A1(_0789_),
    .A2(_0792_),
    .Y(_0208_),
    .B1(_0695_));
 sg13g2_nand3_1 _4242_ (.B(net62),
    .C(net19),
    .A(\Pong.datapath.NES_delay_counter_right.Q[5] ),
    .Y(_0793_));
 sg13g2_nand3_1 _4243_ (.B(_2678_),
    .C(_2677_),
    .A(\Pong.datapath.NES_delay_counter_right.Q[4] ),
    .Y(_0794_));
 sg13g2_xnor2_1 _4244_ (.Y(_0795_),
    .A(\Pong.datapath.NES_delay_counter_right.Q[5] ),
    .B(_0794_));
 sg13g2_nand2b_1 _4245_ (.Y(_0796_),
    .B(_0795_),
    .A_N(net18));
 sg13g2_a21oi_1 _4246_ (.A1(_0793_),
    .A2(_0796_),
    .Y(_0209_),
    .B1(_0695_));
 sg13g2_nand3_1 _4247_ (.B(net62),
    .C(_0726_),
    .A(_2674_),
    .Y(_0797_));
 sg13g2_nand2_1 _4248_ (.Y(_0798_),
    .A(_2677_),
    .B(_2680_));
 sg13g2_xnor2_1 _4249_ (.Y(_0799_),
    .A(_2674_),
    .B(_0798_));
 sg13g2_nand2b_1 _4250_ (.Y(_0800_),
    .B(_0799_),
    .A_N(_0728_));
 sg13g2_buf_1 _4251_ (.A(_2657_),
    .X(_0801_));
 sg13g2_a21oi_1 _4252_ (.A1(_0797_),
    .A2(_0800_),
    .Y(_0210_),
    .B1(_0801_));
 sg13g2_nand3_1 _4253_ (.B(net62),
    .C(_0726_),
    .A(\Pong.datapath.NES_delay_counter_right.Q[7] ),
    .Y(_0802_));
 sg13g2_nand3_1 _4254_ (.B(_2677_),
    .C(_2680_),
    .A(_2674_),
    .Y(_0803_));
 sg13g2_xnor2_1 _4255_ (.Y(_0804_),
    .A(\Pong.datapath.NES_delay_counter_right.Q[7] ),
    .B(_0803_));
 sg13g2_nand2b_1 _4256_ (.Y(_0805_),
    .B(_0804_),
    .A_N(net18));
 sg13g2_a21oi_1 _4257_ (.A1(_0802_),
    .A2(_0805_),
    .Y(_0211_),
    .B1(_0801_));
 sg13g2_xnor2_1 _4258_ (.Y(_0806_),
    .A(_0116_),
    .B(_2682_));
 sg13g2_nor2_1 _4259_ (.A(_0728_),
    .B(_0806_),
    .Y(_0807_));
 sg13g2_a21oi_1 _4260_ (.A1(\Pong.datapath.NES_delay_counter_right.Q[8] ),
    .A2(net19),
    .Y(_0808_),
    .B1(_0807_));
 sg13g2_nor2_1 _4261_ (.A(net96),
    .B(_0808_),
    .Y(_0212_));
 sg13g2_o21ai_1 _4262_ (.B1(_0740_),
    .Y(_0809_),
    .A1(net17),
    .A2(_0731_));
 sg13g2_inv_1 _4263_ (.Y(_0810_),
    .A(_0809_));
 sg13g2_nor2b_1 _4264_ (.A(net17),
    .B_N(_0731_),
    .Y(_0811_));
 sg13g2_o21ai_1 _4265_ (.B1(net188),
    .Y(_0812_),
    .A1(_2693_),
    .A2(_0811_));
 sg13g2_a21oi_1 _4266_ (.A1(_2693_),
    .A2(_0810_),
    .Y(_0213_),
    .B1(_0812_));
 sg13g2_inv_1 _4267_ (.Y(_0813_),
    .A(\Pong.datapath.NES_wire_Left[2] ));
 sg13g2_inv_1 _4268_ (.Y(_0814_),
    .A(\Pong.control_unit.NES_Controller_Left.state_NESController[15] ));
 sg13g2_nand2b_1 _4269_ (.Y(_0815_),
    .B(_2841_),
    .A_N(\Pong.control_unit.NES_Controller_Left.state_NESController[9] ));
 sg13g2_nand2_1 _4270_ (.Y(_0816_),
    .A(_0124_),
    .B(_0123_));
 sg13g2_o21ai_1 _4271_ (.B1(_0122_),
    .Y(_0817_),
    .A1(_0815_),
    .A2(_0816_));
 sg13g2_nor2_1 _4272_ (.A(\Pong.control_unit.NES_Controller_Left.state_NESController[12] ),
    .B(\Pong.control_unit.NES_Controller_Left.state_NESController[7] ),
    .Y(_0818_));
 sg13g2_nand3_1 _4273_ (.B(_0817_),
    .C(_0818_),
    .A(_0121_),
    .Y(_0819_));
 sg13g2_or3_1 _4274_ (.A(_2798_),
    .B(_2797_),
    .C(_2806_),
    .X(_0820_));
 sg13g2_a21o_1 _4275_ (.A2(_0819_),
    .A1(_0120_),
    .B1(_0820_),
    .X(_0821_));
 sg13g2_nor2_1 _4276_ (.A(\Pong.control_unit.NES_Controller_Left.state_NESController[5] ),
    .B(\Pong.control_unit.NES_Controller_Left.state_NESController[10] ),
    .Y(_0822_));
 sg13g2_nand2_1 _4277_ (.Y(_0823_),
    .A(_0119_),
    .B(_0822_));
 sg13g2_a21oi_1 _4278_ (.A1(_0814_),
    .A2(_0821_),
    .Y(_0824_),
    .B1(_0823_));
 sg13g2_buf_2 _4279_ (.A(_0824_),
    .X(_0825_));
 sg13g2_nor4_2 _4280_ (.A(\Pong.control_unit.NES_Controller_Left.state_NESController[16] ),
    .B(\Pong.control_unit.NES_Controller_Left.state_NESController[4] ),
    .C(\Pong.control_unit.NES_Controller_Left.state_NESController[12] ),
    .Y(_0826_),
    .D(\Pong.control_unit.NES_Controller_Left.state_NESController[7] ));
 sg13g2_nor2_1 _4281_ (.A(\Pong.control_unit.NES_Controller_Left.state_NESController[1] ),
    .B(\Pong.control_unit.NES_Controller_Left.state_NESController[9] ),
    .Y(_0827_));
 sg13g2_nor2_1 _4282_ (.A(\Pong.control_unit.NES_Controller_Left.state_NESController[14] ),
    .B(_2841_),
    .Y(_0828_));
 sg13g2_nand4_1 _4283_ (.B(_0826_),
    .C(_0827_),
    .A(_2792_),
    .Y(_0829_),
    .D(_0828_));
 sg13g2_nand3_1 _4284_ (.B(_0119_),
    .C(_0822_),
    .A(_0814_),
    .Y(_0830_));
 sg13g2_nor2_1 _4285_ (.A(_2806_),
    .B(_0830_),
    .Y(_0831_));
 sg13g2_nor4_1 _4286_ (.A(_2798_),
    .B(_2797_),
    .C(\Pong.control_unit.NES_Controller_Left.state_NESController[2] ),
    .D(_2844_),
    .Y(_0832_));
 sg13g2_and2_1 _4287_ (.A(_0831_),
    .B(_0832_),
    .X(_0833_));
 sg13g2_nor2b_1 _4288_ (.A(_0829_),
    .B_N(_0833_),
    .Y(_0834_));
 sg13g2_inv_1 _4289_ (.Y(_0835_),
    .A(_0834_));
 sg13g2_nand2_1 _4290_ (.Y(_0836_),
    .A(_0825_),
    .B(_0835_));
 sg13g2_nor4_2 _4291_ (.A(\Pong.control_unit.NES_Controller_Left.state_NESController[2] ),
    .B(_2844_),
    .C(_0820_),
    .Y(_0837_),
    .D(_0830_));
 sg13g2_nand2_1 _4292_ (.Y(_0838_),
    .A(_0124_),
    .B(_0815_));
 sg13g2_nand3_1 _4293_ (.B(_0826_),
    .C(_0838_),
    .A(_0121_),
    .Y(_0839_));
 sg13g2_a21oi_1 _4294_ (.A1(_0120_),
    .A2(_0839_),
    .Y(_0840_),
    .B1(_2797_));
 sg13g2_o21ai_1 _4295_ (.B1(_0831_),
    .Y(_0841_),
    .A1(_2798_),
    .A2(_0840_));
 sg13g2_buf_1 _4296_ (.A(_0841_),
    .X(_0842_));
 sg13g2_nand4_1 _4297_ (.B(_2838_),
    .C(_0826_),
    .A(_2792_),
    .Y(_0843_),
    .D(_0827_));
 sg13g2_nor2_1 _4298_ (.A(_2841_),
    .B(_0843_),
    .Y(_0844_));
 sg13g2_a21oi_1 _4299_ (.A1(_0124_),
    .A2(_0815_),
    .Y(_0845_),
    .B1(\Pong.control_unit.NES_Controller_Left.state_NESController[4] ));
 sg13g2_o21ai_1 _4300_ (.B1(_0126_),
    .Y(_0846_),
    .A1(\Pong.control_unit.NES_Controller_Left.state_NESController[16] ),
    .A2(_0845_));
 sg13g2_and2_1 _4301_ (.A(_0125_),
    .B(_0846_),
    .X(_0847_));
 sg13g2_nand2_1 _4302_ (.Y(_0848_),
    .A(_0844_),
    .B(_0847_));
 sg13g2_nand2_1 _4303_ (.Y(_0849_),
    .A(_0125_),
    .B(_0846_));
 sg13g2_nand2_1 _4304_ (.Y(_0850_),
    .A(_0829_),
    .B(_0849_));
 sg13g2_o21ai_1 _4305_ (.B1(_0850_),
    .Y(_0851_),
    .A1(_0825_),
    .A2(_0848_));
 sg13g2_nand3_1 _4306_ (.B(_0842_),
    .C(_0851_),
    .A(_0837_),
    .Y(_0852_));
 sg13g2_inv_1 _4307_ (.Y(_0853_),
    .A(_0842_));
 sg13g2_o21ai_1 _4308_ (.B1(_0837_),
    .Y(_0854_),
    .A1(_0844_),
    .A2(_0849_));
 sg13g2_nand2_1 _4309_ (.Y(_0855_),
    .A(_0853_),
    .B(_0854_));
 sg13g2_nand3_1 _4310_ (.B(_0852_),
    .C(_0855_),
    .A(_0836_),
    .Y(_0856_));
 sg13g2_or2_1 _4311_ (.X(_0857_),
    .B(_0842_),
    .A(_0825_));
 sg13g2_inv_1 _4312_ (.Y(_0858_),
    .A(net1));
 sg13g2_nand4_1 _4313_ (.B(_0829_),
    .C(_0833_),
    .A(_0858_),
    .Y(_0859_),
    .D(_0849_));
 sg13g2_o21ai_1 _4314_ (.B1(net188),
    .Y(_0860_),
    .A1(_0857_),
    .A2(_0859_));
 sg13g2_a21oi_1 _4315_ (.A1(_0813_),
    .A2(_0856_),
    .Y(_0214_),
    .B1(_0860_));
 sg13g2_o21ai_1 _4316_ (.B1(_0850_),
    .Y(_0861_),
    .A1(_0853_),
    .A2(_0848_));
 sg13g2_nand3b_1 _4317_ (.B(_0837_),
    .C(_0861_),
    .Y(_0862_),
    .A_N(_0825_));
 sg13g2_a22oi_1 _4318_ (.Y(_0863_),
    .B1(_0854_),
    .B2(_0825_),
    .A2(_0853_),
    .A1(_0835_));
 sg13g2_a21oi_1 _4319_ (.A1(_0862_),
    .A2(_0863_),
    .Y(_0864_),
    .B1(\Pong.datapath.NES_wire_Left[3] ));
 sg13g2_nand2_1 _4320_ (.Y(_0865_),
    .A(_0825_),
    .B(_0842_));
 sg13g2_o21ai_1 _4321_ (.B1(net188),
    .Y(_0866_),
    .A1(_0859_),
    .A2(_0865_));
 sg13g2_nor2_1 _4322_ (.A(_0864_),
    .B(_0866_),
    .Y(_0215_));
 sg13g2_nand2b_1 _4323_ (.Y(_0867_),
    .B(_0842_),
    .A_N(_0825_));
 sg13g2_nand2_1 _4324_ (.Y(_0868_),
    .A(_0834_),
    .B(_0847_));
 sg13g2_o21ai_1 _4325_ (.B1(_0859_),
    .Y(_0869_),
    .A1(\Pong.datapath.NES_wire_Left[4] ),
    .A2(_0868_));
 sg13g2_o21ai_1 _4326_ (.B1(_0867_),
    .Y(_0870_),
    .A1(\Pong.datapath.NES_wire_Left[4] ),
    .A2(_0834_));
 sg13g2_o21ai_1 _4327_ (.B1(_0870_),
    .Y(_0871_),
    .A1(_0867_),
    .A2(_0869_));
 sg13g2_and2_1 _4328_ (.A(net139),
    .B(_0871_),
    .X(_0216_));
 sg13g2_nand2_1 _4329_ (.Y(_0872_),
    .A(_0857_),
    .B(_0865_));
 sg13g2_o21ai_1 _4330_ (.B1(_0850_),
    .Y(_0873_),
    .A1(_0867_),
    .A2(_0848_));
 sg13g2_a22oi_1 _4331_ (.Y(_0874_),
    .B1(_0873_),
    .B2(_0833_),
    .A2(_0872_),
    .A1(_0835_));
 sg13g2_nor2_1 _4332_ (.A(\Pong.datapath.NES_wire_Left[5] ),
    .B(_0874_),
    .Y(_0875_));
 sg13g2_nand2_1 _4333_ (.Y(_0876_),
    .A(_0858_),
    .B(_0825_));
 sg13g2_o21ai_1 _4334_ (.B1(net188),
    .Y(_0877_),
    .A1(_0855_),
    .A2(_0876_));
 sg13g2_nor2_1 _4335_ (.A(_0875_),
    .B(_0877_),
    .Y(_0217_));
 sg13g2_nor2_1 _4336_ (.A(\Pong.control_unit.NES_Controller_Right.state_NESController[5] ),
    .B(\Pong.control_unit.NES_Controller_Right.state_NESController[10] ),
    .Y(_0878_));
 sg13g2_nand2_1 _4337_ (.Y(_0879_),
    .A(_0538_),
    .B(_0878_));
 sg13g2_nor2_1 _4338_ (.A(\Pong.control_unit.NES_Controller_Right.state_NESController[7] ),
    .B(\Pong.control_unit.NES_Controller_Right.state_NESController[12] ),
    .Y(_0880_));
 sg13g2_nand2b_1 _4339_ (.Y(_0881_),
    .B(\Pong.control_unit.NES_Controller_Right.state_NESController[18] ),
    .A_N(_2671_));
 sg13g2_nand2_1 _4340_ (.Y(_0882_),
    .A(_0132_),
    .B(_0131_));
 sg13g2_o21ai_1 _4341_ (.B1(_0130_),
    .Y(_0883_),
    .A1(_0881_),
    .A2(_0882_));
 sg13g2_nand3_1 _4342_ (.B(_0880_),
    .C(_0883_),
    .A(_0129_),
    .Y(_0884_));
 sg13g2_nand2_1 _4343_ (.Y(_0885_),
    .A(_0128_),
    .B(_0884_));
 sg13g2_nor3_1 _4344_ (.A(_2665_),
    .B(_2666_),
    .C(_2704_),
    .Y(_0886_));
 sg13g2_a21oi_1 _4345_ (.A1(_0885_),
    .A2(_0886_),
    .Y(_0887_),
    .B1(\Pong.control_unit.NES_Controller_Right.state_NESController[15] ));
 sg13g2_nor2_1 _4346_ (.A(_0879_),
    .B(_0887_),
    .Y(_0888_));
 sg13g2_buf_2 _4347_ (.A(_0888_),
    .X(_0889_));
 sg13g2_nor2_1 _4348_ (.A(_2707_),
    .B(_2713_),
    .Y(_0890_));
 sg13g2_nand2_1 _4349_ (.Y(_0891_),
    .A(_0132_),
    .B(_0881_));
 sg13g2_nand4_1 _4350_ (.B(_0880_),
    .C(_0890_),
    .A(_0129_),
    .Y(_0892_),
    .D(_0891_));
 sg13g2_a21oi_1 _4351_ (.A1(_0128_),
    .A2(_0892_),
    .Y(_0893_),
    .B1(_2665_));
 sg13g2_nand3b_1 _4352_ (.B(_0538_),
    .C(_0878_),
    .Y(_0894_),
    .A_N(\Pong.control_unit.NES_Controller_Right.state_NESController[15] ));
 sg13g2_nor2_1 _4353_ (.A(_2704_),
    .B(_0894_),
    .Y(_0895_));
 sg13g2_o21ai_1 _4354_ (.B1(_0895_),
    .Y(_0896_),
    .A1(_2666_),
    .A2(_0893_));
 sg13g2_buf_2 _4355_ (.A(_0896_),
    .X(_0897_));
 sg13g2_a21oi_1 _4356_ (.A1(_0132_),
    .A2(_0881_),
    .Y(_0898_),
    .B1(_2707_));
 sg13g2_o21ai_1 _4357_ (.B1(_0134_),
    .Y(_0899_),
    .A1(_2713_),
    .A2(_0898_));
 sg13g2_nor4_1 _4358_ (.A(_2665_),
    .B(_2666_),
    .C(\Pong.control_unit.NES_Controller_Right.state_NESController[2] ),
    .D(\Pong.control_unit.NES_Controller_Right.state_NESController[17] ),
    .Y(_0900_));
 sg13g2_nand2_1 _4359_ (.Y(_0901_),
    .A(_0895_),
    .B(_0900_));
 sg13g2_a21oi_1 _4360_ (.A1(_0133_),
    .A2(_0899_),
    .Y(_0902_),
    .B1(_0901_));
 sg13g2_buf_1 _4361_ (.A(_0902_),
    .X(_0903_));
 sg13g2_nor2_1 _4362_ (.A(_0897_),
    .B(_0903_),
    .Y(_0904_));
 sg13g2_nor2_1 _4363_ (.A(\Pong.control_unit.NES_Controller_Right.state_NESController[14] ),
    .B(\Pong.control_unit.NES_Controller_Right.state_NESController[18] ),
    .Y(_0905_));
 sg13g2_nor4_1 _4364_ (.A(_2671_),
    .B(\Pong.control_unit.NES_Controller_Right.state_NESController[1] ),
    .C(_2707_),
    .D(_2713_),
    .Y(_0906_));
 sg13g2_nand4_1 _4365_ (.B(_0880_),
    .C(_0905_),
    .A(\Pong.control_unit.NES_Controller_Right.state_NESController[11] ),
    .Y(_0907_),
    .D(_0906_));
 sg13g2_nor2_1 _4366_ (.A(_0901_),
    .B(_0907_),
    .Y(_0908_));
 sg13g2_buf_1 _4367_ (.A(_0908_),
    .X(_0909_));
 sg13g2_inv_1 _4368_ (.Y(_0910_),
    .A(_0909_));
 sg13g2_o21ai_1 _4369_ (.B1(_0910_),
    .Y(_0911_),
    .A1(_0889_),
    .A2(_0904_));
 sg13g2_nand2b_1 _4370_ (.Y(_0912_),
    .B(_0903_),
    .A_N(_0909_));
 sg13g2_inv_1 _4371_ (.Y(_0913_),
    .A(_0912_));
 sg13g2_nand2b_1 _4372_ (.Y(_0914_),
    .B(_0909_),
    .A_N(_0903_));
 sg13g2_nor2_1 _4373_ (.A(_0889_),
    .B(_0914_),
    .Y(_0915_));
 sg13g2_o21ai_1 _4374_ (.B1(_0897_),
    .Y(_0916_),
    .A1(_0913_),
    .A2(_0915_));
 sg13g2_a21oi_1 _4375_ (.A1(_0911_),
    .A2(_0916_),
    .Y(_0917_),
    .B1(\Pong.datapath.NES_wire_Right[2] ));
 sg13g2_nor2_1 _4376_ (.A(_0889_),
    .B(_0897_),
    .Y(_0918_));
 sg13g2_nor2_1 _4377_ (.A(net2),
    .B(_0909_),
    .Y(_0919_));
 sg13g2_and3_1 _4378_ (.X(_0920_),
    .A(_0903_),
    .B(_0918_),
    .C(_0919_));
 sg13g2_nor3_1 _4379_ (.A(net138),
    .B(_0917_),
    .C(_0920_),
    .Y(_0218_));
 sg13g2_nand2b_1 _4380_ (.Y(_0921_),
    .B(_0889_),
    .A_N(_0903_));
 sg13g2_a21oi_1 _4381_ (.A1(_0897_),
    .A2(_0921_),
    .Y(_0922_),
    .B1(_0909_));
 sg13g2_nand2b_1 _4382_ (.Y(_0923_),
    .B(_0897_),
    .A_N(_0914_));
 sg13g2_a21oi_1 _4383_ (.A1(_0912_),
    .A2(_0923_),
    .Y(_0924_),
    .B1(_0889_));
 sg13g2_inv_1 _4384_ (.Y(_0925_),
    .A(\Pong.datapath.NES_wire_Right[3] ));
 sg13g2_o21ai_1 _4385_ (.B1(_0925_),
    .Y(_0926_),
    .A1(_0922_),
    .A2(_0924_));
 sg13g2_nand4_1 _4386_ (.B(_0897_),
    .C(_0903_),
    .A(_0889_),
    .Y(_0927_),
    .D(_0919_));
 sg13g2_and3_1 _4387_ (.X(_0219_),
    .A(_2717_),
    .B(_0926_),
    .C(_0927_));
 sg13g2_nor2_1 _4388_ (.A(\Pong.datapath.NES_wire_Right[4] ),
    .B(_0909_),
    .Y(_0928_));
 sg13g2_or2_1 _4389_ (.X(_0929_),
    .B(_0912_),
    .A(net2));
 sg13g2_o21ai_1 _4390_ (.B1(_0929_),
    .Y(_0930_),
    .A1(\Pong.datapath.NES_wire_Right[4] ),
    .A2(_0914_));
 sg13g2_nor2b_1 _4391_ (.A(_0889_),
    .B_N(_0897_),
    .Y(_0931_));
 sg13g2_mux2_1 _4392_ (.A0(_0928_),
    .A1(_0930_),
    .S(_0931_),
    .X(_0932_));
 sg13g2_nor2_1 _4393_ (.A(_0730_),
    .B(_0932_),
    .Y(_0220_));
 sg13g2_nor3_1 _4394_ (.A(_0879_),
    .B(_0887_),
    .C(_0909_),
    .Y(_0933_));
 sg13g2_o21ai_1 _4395_ (.B1(_0897_),
    .Y(_0934_),
    .A1(_0915_),
    .A2(_0933_));
 sg13g2_o21ai_1 _4396_ (.B1(_0910_),
    .Y(_0935_),
    .A1(_0903_),
    .A2(_0918_));
 sg13g2_a21oi_1 _4397_ (.A1(_0934_),
    .A2(_0935_),
    .Y(_0936_),
    .B1(\Pong.datapath.NES_wire_Right[5] ));
 sg13g2_and3_1 _4398_ (.X(_0937_),
    .A(_0889_),
    .B(_0904_),
    .C(_0919_));
 sg13g2_nor3_1 _4399_ (.A(_2663_),
    .B(_0936_),
    .C(_0937_),
    .Y(_0221_));
 sg13g2_buf_1 _4400_ (.A(\Pong.datapath.ballFunction.reset_n ),
    .X(_0938_));
 sg13g2_buf_1 _4401_ (.A(_0938_),
    .X(_0939_));
 sg13g2_inv_2 _4402_ (.Y(_0940_),
    .A(net49));
 sg13g2_buf_2 _4403_ (.A(_0115_),
    .X(_0941_));
 sg13g2_nor2_1 _4404_ (.A(_2724_),
    .B(_2725_),
    .Y(_0942_));
 sg13g2_nand2_1 _4405_ (.Y(_0943_),
    .A(\Pong.control_unit.state_ballMovement[1] ),
    .B(_0942_));
 sg13g2_and3_1 _4406_ (.X(_0944_),
    .A(net187),
    .B(_0941_),
    .C(_0943_));
 sg13g2_buf_1 _4407_ (.A(_0944_),
    .X(_0945_));
 sg13g2_buf_1 _4408_ (.A(net88),
    .X(_0946_));
 sg13g2_or2_1 _4409_ (.X(_0947_),
    .B(_2720_),
    .A(_2725_));
 sg13g2_buf_1 _4410_ (.A(_0947_),
    .X(_0948_));
 sg13g2_a21o_1 _4411_ (.A2(_0941_),
    .A1(_2724_),
    .B1(_0948_),
    .X(_0949_));
 sg13g2_nand2b_1 _4412_ (.Y(_0950_),
    .B(_0941_),
    .A_N(\Pong.control_unit.state_ballMovement[1] ));
 sg13g2_nor2_1 _4413_ (.A(_0949_),
    .B(_0950_),
    .Y(_0951_));
 sg13g2_a221oi_1 _4414_ (.B2(_0940_),
    .C1(net88),
    .B1(_0951_),
    .A1(_0085_),
    .Y(_0952_),
    .A2(_0949_));
 sg13g2_a21oi_1 _4415_ (.A1(_0940_),
    .A2(net78),
    .Y(_0953_),
    .B1(_0952_));
 sg13g2_and2_1 _4416_ (.A(net137),
    .B(_0953_),
    .X(_0222_));
 sg13g2_nand2_1 _4417_ (.Y(_0954_),
    .A(\Pong.control_unit.state_ballMovement[3] ),
    .B(\Pong.control_unit.state_ballMovement[1] ));
 sg13g2_o21ai_1 _4418_ (.B1(_0954_),
    .Y(_0955_),
    .A1(\Pong.control_unit.state_ballMovement[3] ),
    .A2(_0950_));
 sg13g2_nand2_1 _4419_ (.Y(_0956_),
    .A(_0942_),
    .B(_0955_));
 sg13g2_o21ai_1 _4420_ (.B1(_0956_),
    .Y(_0957_),
    .A1(_2741_),
    .A2(_0941_));
 sg13g2_buf_2 _4421_ (.A(_0957_),
    .X(_0958_));
 sg13g2_buf_1 _4422_ (.A(_0958_),
    .X(_0959_));
 sg13g2_a21oi_1 _4423_ (.A1(_2724_),
    .A2(_0941_),
    .Y(_0960_),
    .B1(_2725_));
 sg13g2_nor2_1 _4424_ (.A(net187),
    .B(_0960_),
    .Y(_0961_));
 sg13g2_buf_1 _4425_ (.A(_0961_),
    .X(_0962_));
 sg13g2_nand3_1 _4426_ (.B(_0941_),
    .C(_0943_),
    .A(net187),
    .Y(_0963_));
 sg13g2_buf_1 _4427_ (.A(_0963_),
    .X(_0964_));
 sg13g2_or2_1 _4428_ (.X(_0965_),
    .B(_0960_),
    .A(net187));
 sg13g2_buf_2 _4429_ (.A(_0965_),
    .X(_0966_));
 sg13g2_nand2_1 _4430_ (.Y(_0967_),
    .A(net87),
    .B(_0966_));
 sg13g2_nand2b_1 _4431_ (.Y(_0968_),
    .B(net87),
    .A_N(_0958_));
 sg13g2_buf_1 _4432_ (.A(_3051_),
    .X(_0969_));
 sg13g2_buf_1 _4433_ (.A(net43),
    .X(_0970_));
 sg13g2_mux4_1 _4434_ (.S0(_0940_),
    .A0(net77),
    .A1(net94),
    .A2(_0967_),
    .A3(_0968_),
    .S1(net28),
    .X(_0971_));
 sg13g2_and2_1 _4435_ (.A(net137),
    .B(_0971_),
    .X(_0223_));
 sg13g2_buf_1 _4436_ (.A(net50),
    .X(_0972_));
 sg13g2_nor2_1 _4437_ (.A(net28),
    .B(net77),
    .Y(_0973_));
 sg13g2_a21oi_1 _4438_ (.A1(net28),
    .A2(_0966_),
    .Y(_0974_),
    .B1(_0973_));
 sg13g2_buf_1 _4439_ (.A(_0086_),
    .X(_0975_));
 sg13g2_inv_1 _4440_ (.Y(_0976_),
    .A(net66));
 sg13g2_o21ai_1 _4441_ (.B1(net66),
    .Y(_0977_),
    .A1(net28),
    .A2(_0966_));
 sg13g2_o21ai_1 _4442_ (.B1(_0977_),
    .Y(_0978_),
    .A1(net66),
    .A2(net77));
 sg13g2_and2_1 _4443_ (.A(net28),
    .B(_0975_),
    .X(_0979_));
 sg13g2_a221oi_1 _4444_ (.B2(_0958_),
    .C1(_0940_),
    .B1(_0979_),
    .A1(_0976_),
    .Y(_0980_),
    .A2(net94));
 sg13g2_a21oi_1 _4445_ (.A1(_0940_),
    .A2(_0978_),
    .Y(_0981_),
    .B1(_0980_));
 sg13g2_a221oi_1 _4446_ (.B2(_0976_),
    .C1(_0981_),
    .B1(_0974_),
    .A1(_0972_),
    .Y(_0982_),
    .A2(net78));
 sg13g2_buf_1 _4447_ (.A(_0938_),
    .X(_0983_));
 sg13g2_nor2b_1 _4448_ (.A(_0982_),
    .B_N(net136),
    .Y(_0224_));
 sg13g2_nand4_1 _4449_ (.B(_0972_),
    .C(_0496_),
    .A(net28),
    .Y(_0984_),
    .D(_0958_));
 sg13g2_o21ai_1 _4450_ (.B1(_0984_),
    .Y(_0985_),
    .A1(_0496_),
    .A2(_0966_));
 sg13g2_o21ai_1 _4451_ (.B1(_0496_),
    .Y(_0986_),
    .A1(_0463_),
    .A2(_0966_));
 sg13g2_o21ai_1 _4452_ (.B1(_0986_),
    .Y(_0987_),
    .A1(_0496_),
    .A2(_0958_));
 sg13g2_nand2_1 _4453_ (.Y(_0988_),
    .A(net28),
    .B(net50));
 sg13g2_a22oi_1 _4454_ (.Y(_0989_),
    .B1(_0988_),
    .B2(_0958_),
    .A2(net94),
    .A1(_0463_));
 sg13g2_or2_1 _4455_ (.X(_0990_),
    .B(_0989_),
    .A(_0496_));
 sg13g2_o21ai_1 _4456_ (.B1(_0990_),
    .Y(_0991_),
    .A1(net49),
    .A2(_0987_));
 sg13g2_a21oi_1 _4457_ (.A1(net49),
    .A2(_0985_),
    .Y(_0992_),
    .B1(_0991_));
 sg13g2_nor2_1 _4458_ (.A(net33),
    .B(net87),
    .Y(_0993_));
 sg13g2_a21oi_1 _4459_ (.A1(net87),
    .A2(_0992_),
    .Y(_0994_),
    .B1(_0993_));
 sg13g2_and2_1 _4460_ (.A(net137),
    .B(_0994_),
    .X(_0225_));
 sg13g2_buf_1 _4461_ (.A(_0087_),
    .X(_0995_));
 sg13g2_nor2_1 _4462_ (.A(_3050_),
    .B(net43),
    .Y(_0996_));
 sg13g2_buf_1 _4463_ (.A(_0996_),
    .X(_0997_));
 sg13g2_nor2_2 _4464_ (.A(_3046_),
    .B(net67),
    .Y(_0998_));
 sg13g2_and2_1 _4465_ (.A(net16),
    .B(_0998_),
    .X(_0999_));
 sg13g2_buf_1 _4466_ (.A(_0999_),
    .X(_1000_));
 sg13g2_a22oi_1 _4467_ (.Y(_1001_),
    .B1(net94),
    .B2(_1000_),
    .A2(net77),
    .A1(_3055_));
 sg13g2_nand2_1 _4468_ (.Y(_1002_),
    .A(net16),
    .B(_0998_));
 sg13g2_a221oi_1 _4469_ (.B2(_1002_),
    .C1(_0995_),
    .B1(net94),
    .A1(_3054_),
    .Y(_1003_),
    .A2(_0958_));
 sg13g2_a21oi_1 _4470_ (.A1(_0995_),
    .A2(_1001_),
    .Y(_1004_),
    .B1(_1003_));
 sg13g2_a21oi_1 _4471_ (.A1(net32),
    .A2(net78),
    .Y(_1005_),
    .B1(_1004_));
 sg13g2_nor2b_1 _4472_ (.A(_1005_),
    .B_N(net136),
    .Y(_0226_));
 sg13g2_buf_1 _4473_ (.A(_3056_),
    .X(_1006_));
 sg13g2_buf_1 _4474_ (.A(_0088_),
    .X(_1007_));
 sg13g2_or2_1 _4475_ (.X(_1008_),
    .B(net43),
    .A(_3050_));
 sg13g2_buf_1 _4476_ (.A(_1008_),
    .X(_1009_));
 sg13g2_or3_1 _4477_ (.A(_3046_),
    .B(_3048_),
    .C(net46),
    .X(_1010_));
 sg13g2_nor2_1 _4478_ (.A(_1009_),
    .B(_1010_),
    .Y(_1011_));
 sg13g2_nand2_1 _4479_ (.Y(_1012_),
    .A(_3050_),
    .B(net43));
 sg13g2_buf_2 _4480_ (.A(_1012_),
    .X(_1013_));
 sg13g2_nand3_1 _4481_ (.B(net67),
    .C(net46),
    .A(_3046_),
    .Y(_1014_));
 sg13g2_buf_2 _4482_ (.A(_1014_),
    .X(_1015_));
 sg13g2_nor2_1 _4483_ (.A(_1013_),
    .B(_1015_),
    .Y(_1016_));
 sg13g2_a22oi_1 _4484_ (.Y(_1017_),
    .B1(_1016_),
    .B2(net77),
    .A2(_1011_),
    .A1(net94));
 sg13g2_nand2_1 _4485_ (.Y(_1018_),
    .A(_1007_),
    .B(_1017_));
 sg13g2_o21ai_1 _4486_ (.B1(_0958_),
    .Y(_1019_),
    .A1(_1013_),
    .A2(_1015_));
 sg13g2_o21ai_1 _4487_ (.B1(_1019_),
    .Y(_1020_),
    .A1(_0966_),
    .A2(_1011_));
 sg13g2_or2_1 _4488_ (.X(_1021_),
    .B(_1020_),
    .A(_1007_));
 sg13g2_a22oi_1 _4489_ (.Y(_1022_),
    .B1(_1018_),
    .B2(_1021_),
    .A2(net78),
    .A1(net42));
 sg13g2_nor2b_1 _4490_ (.A(_1022_),
    .B_N(net136),
    .Y(_0227_));
 sg13g2_buf_2 _4491_ (.A(_0089_),
    .X(_1023_));
 sg13g2_nand4_1 _4492_ (.B(net67),
    .C(_3056_),
    .A(net51),
    .Y(_1024_),
    .D(net46));
 sg13g2_nor2_1 _4493_ (.A(_1013_),
    .B(_1024_),
    .Y(_1025_));
 sg13g2_xor2_1 _4494_ (.B(_1025_),
    .A(_1023_),
    .X(_1026_));
 sg13g2_nor4_1 _4495_ (.A(_3046_),
    .B(net67),
    .C(_3056_),
    .D(net46),
    .Y(_1027_));
 sg13g2_buf_2 _4496_ (.A(_1027_),
    .X(_1028_));
 sg13g2_nand2_1 _4497_ (.Y(_1029_),
    .A(_0997_),
    .B(_1028_));
 sg13g2_xnor2_1 _4498_ (.Y(_1030_),
    .A(_1023_),
    .B(_1029_));
 sg13g2_a22oi_1 _4499_ (.Y(_1031_),
    .B1(_1030_),
    .B2(net94),
    .A2(_1026_),
    .A1(net77));
 sg13g2_o21ai_1 _4500_ (.B1(_1031_),
    .Y(_1032_),
    .A1(net48),
    .A2(_0964_));
 sg13g2_nand2_1 _4501_ (.Y(_0228_),
    .A(_0939_),
    .B(_1032_));
 sg13g2_nor3_2 _4502_ (.A(net42),
    .B(net46),
    .C(net48),
    .Y(_1033_));
 sg13g2_nand2_1 _4503_ (.Y(_1034_),
    .A(_1000_),
    .B(_1033_));
 sg13g2_nand2_1 _4504_ (.Y(_1035_),
    .A(_0489_),
    .B(_1016_));
 sg13g2_nand2b_1 _4505_ (.Y(_1036_),
    .B(_0959_),
    .A_N(_1035_));
 sg13g2_o21ai_1 _4506_ (.B1(_1036_),
    .Y(_1037_),
    .A1(_0966_),
    .A2(_1034_));
 sg13g2_a22oi_1 _4507_ (.Y(_1038_),
    .B1(_1034_),
    .B2(_0962_),
    .A2(_1035_),
    .A1(_0959_));
 sg13g2_nor2_1 _4508_ (.A(_0492_),
    .B(_1038_),
    .Y(_1039_));
 sg13g2_a221oi_1 _4509_ (.B2(_0492_),
    .C1(_1039_),
    .B1(_1037_),
    .A1(net68),
    .Y(_1040_),
    .A2(net88));
 sg13g2_nor2b_1 _4510_ (.A(_1040_),
    .B_N(_0983_),
    .Y(_0229_));
 sg13g2_nor2_1 _4511_ (.A(_3041_),
    .B(net68),
    .Y(_1041_));
 sg13g2_nand2_1 _4512_ (.Y(_1042_),
    .A(_1041_),
    .B(_1028_));
 sg13g2_nor2_1 _4513_ (.A(_1009_),
    .B(_1042_),
    .Y(_1043_));
 sg13g2_xor2_1 _4514_ (.B(_1043_),
    .A(_0090_),
    .X(_1044_));
 sg13g2_and4_1 _4515_ (.A(_0969_),
    .B(net51),
    .C(net67),
    .D(net46),
    .X(_1045_));
 sg13g2_buf_2 _4516_ (.A(_1045_),
    .X(_1046_));
 sg13g2_and3_1 _4517_ (.X(_1047_),
    .A(_3056_),
    .B(_3041_),
    .C(\Pong.datapath.ballFunction.ball_center_x[7] ));
 sg13g2_buf_1 _4518_ (.A(_1047_),
    .X(_1048_));
 sg13g2_nand3_1 _4519_ (.B(_1046_),
    .C(_1048_),
    .A(_0460_),
    .Y(_1049_));
 sg13g2_xnor2_1 _4520_ (.Y(_1050_),
    .A(_0090_),
    .B(_1049_));
 sg13g2_a22oi_1 _4521_ (.Y(_1051_),
    .B1(_1050_),
    .B2(net77),
    .A2(_1044_),
    .A1(net94));
 sg13g2_o21ai_1 _4522_ (.B1(_1051_),
    .Y(_1052_),
    .A1(net45),
    .A2(_0964_));
 sg13g2_nand2_1 _4523_ (.Y(_0230_),
    .A(_0939_),
    .B(_1052_));
 sg13g2_buf_2 _4524_ (.A(_0091_),
    .X(_1053_));
 sg13g2_and3_1 _4525_ (.X(_1054_),
    .A(_3046_),
    .B(_3048_),
    .C(_3058_));
 sg13g2_buf_1 _4526_ (.A(_1054_),
    .X(_1055_));
 sg13g2_nand4_1 _4527_ (.B(_3053_),
    .C(_1055_),
    .A(net45),
    .Y(_1056_),
    .D(_1048_));
 sg13g2_xor2_1 _4528_ (.B(_1056_),
    .A(_1053_),
    .X(_1057_));
 sg13g2_nand3_1 _4529_ (.B(_1000_),
    .C(_1033_),
    .A(_0461_),
    .Y(_1058_));
 sg13g2_xnor2_1 _4530_ (.Y(_1059_),
    .A(_1053_),
    .B(_1058_));
 sg13g2_nor2_1 _4531_ (.A(_0966_),
    .B(_1059_),
    .Y(_1060_));
 sg13g2_a221oi_1 _4532_ (.B2(_1057_),
    .C1(_1060_),
    .B1(net77),
    .A1(_0466_),
    .Y(_1061_),
    .A2(net88));
 sg13g2_nor2b_1 _4533_ (.A(_1061_),
    .B_N(_0983_),
    .Y(_0231_));
 sg13g2_a221oi_1 _4534_ (.B2(_0304_),
    .C1(_0945_),
    .B1(_0951_),
    .A1(_0092_),
    .Y(_1062_),
    .A2(_0949_));
 sg13g2_a21oi_1 _4535_ (.A1(_0304_),
    .A2(net78),
    .Y(_1063_),
    .B1(_1062_));
 sg13g2_and2_1 _4536_ (.A(net136),
    .B(_1063_),
    .X(_0232_));
 sg13g2_nor2_2 _4537_ (.A(_2725_),
    .B(_2720_),
    .Y(_1064_));
 sg13g2_o21ai_1 _4538_ (.B1(_0941_),
    .Y(_1065_),
    .A1(_2724_),
    .A2(_2738_));
 sg13g2_a21oi_1 _4539_ (.A1(_1064_),
    .A2(_1065_),
    .Y(_1066_),
    .B1(_0945_));
 sg13g2_buf_1 _4540_ (.A(_1066_),
    .X(_1067_));
 sg13g2_xnor2_1 _4541_ (.Y(_1068_),
    .A(_0304_),
    .B(_1064_));
 sg13g2_a21o_1 _4542_ (.A2(_1068_),
    .A1(net76),
    .B1(net88),
    .X(_1069_));
 sg13g2_nor3_1 _4543_ (.A(net35),
    .B(net88),
    .C(_1068_),
    .Y(_1070_));
 sg13g2_a22oi_1 _4544_ (.Y(_1071_),
    .B1(_1070_),
    .B2(net76),
    .A2(_1069_),
    .A1(net35));
 sg13g2_nor2b_1 _4545_ (.A(_1071_),
    .B_N(net136),
    .Y(_0233_));
 sg13g2_nor2_1 _4546_ (.A(net58),
    .B(net74),
    .Y(_1072_));
 sg13g2_buf_2 _4547_ (.A(_1072_),
    .X(_1073_));
 sg13g2_nor2_1 _4548_ (.A(net88),
    .B(_1064_),
    .Y(_1074_));
 sg13g2_buf_1 _4549_ (.A(_1074_),
    .X(_1075_));
 sg13g2_nand2_1 _4550_ (.Y(_1076_),
    .A(net58),
    .B(net74));
 sg13g2_buf_1 _4551_ (.A(_1076_),
    .X(_1077_));
 sg13g2_nor2_1 _4552_ (.A(net75),
    .B(net15),
    .Y(_1078_));
 sg13g2_a21oi_1 _4553_ (.A1(_1073_),
    .A2(net75),
    .Y(_1079_),
    .B1(_1078_));
 sg13g2_xnor2_1 _4554_ (.Y(_1080_),
    .A(net69),
    .B(_1079_));
 sg13g2_a22oi_1 _4555_ (.Y(_1081_),
    .B1(_1067_),
    .B2(_1080_),
    .A2(net78),
    .A1(_3026_));
 sg13g2_nand2b_1 _4556_ (.Y(_0234_),
    .B(net137),
    .A_N(_1081_));
 sg13g2_nand2_1 _4557_ (.Y(_1082_),
    .A(net74),
    .B(net73));
 sg13g2_nor2_1 _4558_ (.A(_0092_),
    .B(_1082_),
    .Y(_1083_));
 sg13g2_a221oi_1 _4559_ (.B2(_1064_),
    .C1(_2756_),
    .B1(_1083_),
    .A1(_2890_),
    .Y(_1084_),
    .A2(_1075_));
 sg13g2_nand2_1 _4560_ (.Y(_1085_),
    .A(_3026_),
    .B(_1073_));
 sg13g2_or2_1 _4561_ (.X(_1086_),
    .B(_1082_),
    .A(_0092_));
 sg13g2_buf_1 _4562_ (.A(_1086_),
    .X(_1087_));
 sg13g2_a221oi_1 _4563_ (.B2(_1064_),
    .C1(_2755_),
    .B1(_1087_),
    .A1(_1085_),
    .Y(_1088_),
    .A2(net75));
 sg13g2_o21ai_1 _4564_ (.B1(_1067_),
    .Y(_1089_),
    .A1(_1084_),
    .A2(_1088_));
 sg13g2_o21ai_1 _4565_ (.B1(_1089_),
    .Y(_1090_),
    .A1(net36),
    .A2(net87));
 sg13g2_nand2_1 _4566_ (.Y(_0235_),
    .A(net137),
    .B(_1090_));
 sg13g2_nor2_2 _4567_ (.A(_2763_),
    .B(net56),
    .Y(_1091_));
 sg13g2_and2_1 _4568_ (.A(_1073_),
    .B(_1091_),
    .X(_1092_));
 sg13g2_buf_1 _4569_ (.A(_1092_),
    .X(_1093_));
 sg13g2_xnor2_1 _4570_ (.Y(_1094_),
    .A(_2942_),
    .B(_1093_));
 sg13g2_nand2_1 _4571_ (.Y(_1095_),
    .A(net73),
    .B(_2765_));
 sg13g2_buf_2 _4572_ (.A(_1095_),
    .X(_1096_));
 sg13g2_nor2_1 _4573_ (.A(net15),
    .B(_1096_),
    .Y(_1097_));
 sg13g2_xnor2_1 _4574_ (.Y(_1098_),
    .A(_2943_),
    .B(_1097_));
 sg13g2_o21ai_1 _4575_ (.B1(net76),
    .Y(_1099_),
    .A1(net75),
    .A2(_1098_));
 sg13g2_a21oi_1 _4576_ (.A1(_0948_),
    .A2(_1094_),
    .Y(_1100_),
    .B1(_1099_));
 sg13g2_nor2_1 _4577_ (.A(net38),
    .B(net87),
    .Y(_1101_));
 sg13g2_o21ai_1 _4578_ (.B1(net137),
    .Y(_0236_),
    .A1(_1100_),
    .A2(_1101_));
 sg13g2_nand2_1 _4579_ (.Y(_1102_),
    .A(net36),
    .B(net60));
 sg13g2_or2_1 _4580_ (.X(_1103_),
    .B(_1102_),
    .A(_1087_));
 sg13g2_buf_1 _4581_ (.A(_1103_),
    .X(_1104_));
 sg13g2_nor3_2 _4582_ (.A(net73),
    .B(net56),
    .C(net60),
    .Y(_1105_));
 sg13g2_nand3_1 _4583_ (.B(net75),
    .C(_1105_),
    .A(_1073_),
    .Y(_1106_));
 sg13g2_o21ai_1 _4584_ (.B1(_1106_),
    .Y(_1107_),
    .A1(net75),
    .A2(_1104_));
 sg13g2_xnor2_1 _4585_ (.Y(_1108_),
    .A(net70),
    .B(_1107_));
 sg13g2_a22oi_1 _4586_ (.Y(_1109_),
    .B1(net76),
    .B2(_1108_),
    .A2(net78),
    .A1(net61));
 sg13g2_nor2b_1 _4587_ (.A(_1109_),
    .B_N(net136),
    .Y(_0237_));
 sg13g2_nand4_1 _4588_ (.B(_2765_),
    .C(_2749_),
    .A(net73),
    .Y(_1110_),
    .D(net60));
 sg13g2_buf_1 _4589_ (.A(_1110_),
    .X(_1111_));
 sg13g2_or3_1 _4590_ (.A(_0948_),
    .B(net15),
    .C(_1111_),
    .X(_1112_));
 sg13g2_or4_1 _4591_ (.A(\Pong.datapath.ballFunction.ball_center_y[2] ),
    .B(_2765_),
    .C(_2749_),
    .D(_2752_),
    .X(_1113_));
 sg13g2_buf_1 _4592_ (.A(_1113_),
    .X(_1114_));
 sg13g2_nor2_2 _4593_ (.A(_2889_),
    .B(_1114_),
    .Y(_1115_));
 sg13g2_nand3_1 _4594_ (.B(_0948_),
    .C(_1115_),
    .A(net87),
    .Y(_1116_));
 sg13g2_and3_1 _4595_ (.X(_1117_),
    .A(_3033_),
    .B(_1112_),
    .C(_1116_));
 sg13g2_o21ai_1 _4596_ (.B1(_0948_),
    .Y(_1118_),
    .A1(net88),
    .A2(_1115_));
 sg13g2_a21oi_1 _4597_ (.A1(_1112_),
    .A2(_1118_),
    .Y(_1119_),
    .B1(_3033_));
 sg13g2_o21ai_1 _4598_ (.B1(net76),
    .Y(_1120_),
    .A1(_1117_),
    .A2(_1119_));
 sg13g2_o21ai_1 _4599_ (.B1(_1120_),
    .Y(_1121_),
    .A1(net34),
    .A2(net87));
 sg13g2_nand2_1 _4600_ (.Y(_0238_),
    .A(net137),
    .B(_1121_));
 sg13g2_nor4_2 _4601_ (.A(net73),
    .B(_2765_),
    .C(_2749_),
    .Y(_1122_),
    .D(net60));
 sg13g2_nand2_1 _4602_ (.Y(_1123_),
    .A(_1073_),
    .B(_1122_));
 sg13g2_nor2_1 _4603_ (.A(net34),
    .B(_1123_),
    .Y(_1124_));
 sg13g2_nand4_1 _4604_ (.B(net53),
    .C(_2749_),
    .A(net56),
    .Y(_1125_),
    .D(net60));
 sg13g2_buf_1 _4605_ (.A(_1125_),
    .X(_1126_));
 sg13g2_nor3_1 _4606_ (.A(_1074_),
    .B(_1087_),
    .C(_1126_),
    .Y(_1127_));
 sg13g2_a21oi_1 _4607_ (.A1(net75),
    .A2(_1124_),
    .Y(_1128_),
    .B1(_1127_));
 sg13g2_xnor2_1 _4608_ (.Y(_1129_),
    .A(net71),
    .B(_1128_));
 sg13g2_a22oi_1 _4609_ (.Y(_1130_),
    .B1(net76),
    .B2(_1129_),
    .A2(net78),
    .A1(_3000_));
 sg13g2_nand2b_1 _4610_ (.Y(_0239_),
    .B(net137),
    .A_N(_1130_));
 sg13g2_nand4_1 _4611_ (.B(_2772_),
    .C(_2749_),
    .A(_2771_),
    .Y(_1131_),
    .D(_2752_));
 sg13g2_buf_1 _4612_ (.A(_1131_),
    .X(_1132_));
 sg13g2_or2_1 _4613_ (.X(_1133_),
    .B(_1132_),
    .A(_1096_));
 sg13g2_nor2_1 _4614_ (.A(net15),
    .B(_1133_),
    .Y(_1134_));
 sg13g2_xor2_1 _4615_ (.B(_1134_),
    .A(net52),
    .X(_1135_));
 sg13g2_nor2_2 _4616_ (.A(_2771_),
    .B(net53),
    .Y(_1136_));
 sg13g2_nand2_1 _4617_ (.Y(_1137_),
    .A(_1136_),
    .B(_1115_));
 sg13g2_xnor2_1 _4618_ (.Y(_1138_),
    .A(net52),
    .B(_1137_));
 sg13g2_a22oi_1 _4619_ (.Y(_1139_),
    .B1(_1138_),
    .B2(_1075_),
    .A2(_1135_),
    .A1(_1064_));
 sg13g2_a22oi_1 _4620_ (.Y(_1140_),
    .B1(net76),
    .B2(_1139_),
    .A2(_0946_),
    .A1(net54));
 sg13g2_nor2b_1 _4621_ (.A(_1140_),
    .B_N(net136),
    .Y(_0240_));
 sg13g2_nor3_1 _4622_ (.A(_2885_),
    .B(net53),
    .C(net54),
    .Y(_1141_));
 sg13g2_and2_1 _4623_ (.A(_1141_),
    .B(_1115_),
    .X(_1142_));
 sg13g2_nand4_1 _4624_ (.B(net53),
    .C(_2749_),
    .A(_2771_),
    .Y(_1143_),
    .D(_2773_));
 sg13g2_buf_1 _4625_ (.A(_1143_),
    .X(_1144_));
 sg13g2_nor3_1 _4626_ (.A(_1074_),
    .B(_1104_),
    .C(_1144_),
    .Y(_1145_));
 sg13g2_a21oi_1 _4627_ (.A1(net75),
    .A2(_1142_),
    .Y(_1146_),
    .B1(_1145_));
 sg13g2_xor2_1 _4628_ (.B(_1146_),
    .A(_2920_),
    .X(_1147_));
 sg13g2_a22oi_1 _4629_ (.Y(_1148_),
    .B1(net76),
    .B2(_1147_),
    .A2(_0946_),
    .A1(net72));
 sg13g2_nor2b_1 _4630_ (.A(_1148_),
    .B_N(net136),
    .Y(_0241_));
 sg13g2_buf_1 _4631_ (.A(\Pong.datapath.NES_activity_Right[4] ),
    .X(_1149_));
 sg13g2_inv_2 _4632_ (.Y(_1150_),
    .A(_1149_));
 sg13g2_buf_2 _4633_ (.A(\Pong.datapath.NES_activity_Left[4] ),
    .X(_1151_));
 sg13g2_buf_1 _4634_ (.A(_1151_),
    .X(_1152_));
 sg13g2_o21ai_1 _4635_ (.B1(_0507_),
    .Y(_1153_),
    .A1(net135),
    .A2(_0938_));
 sg13g2_buf_1 _4636_ (.A(\Pong.datapath.score_flag ),
    .X(_1154_));
 sg13g2_buf_1 _4637_ (.A(\Pong.datapath.scoreLeft[3] ),
    .X(_1155_));
 sg13g2_buf_1 _4638_ (.A(\Pong.datapath.scoreLeft[2] ),
    .X(_1156_));
 sg13g2_buf_1 _4639_ (.A(\Pong.datapath.scoreLeft[1] ),
    .X(_1157_));
 sg13g2_nor2_1 _4640_ (.A(_1156_),
    .B(net171),
    .Y(_1158_));
 sg13g2_nand3_1 _4641_ (.B(\Pong.datapath.scoreLeft[0] ),
    .C(_1158_),
    .A(_1155_),
    .Y(_1159_));
 sg13g2_buf_1 _4642_ (.A(\Pong.datapath.scoreRight[3] ),
    .X(_1160_));
 sg13g2_buf_2 _4643_ (.A(\Pong.datapath.scoreRight[0] ),
    .X(_1161_));
 sg13g2_buf_1 _4644_ (.A(\Pong.datapath.scoreRight[1] ),
    .X(_1162_));
 sg13g2_nor2_1 _4645_ (.A(\Pong.datapath.scoreRight[2] ),
    .B(net170),
    .Y(_1163_));
 sg13g2_nand3_1 _4646_ (.B(_1161_),
    .C(_1163_),
    .A(_1160_),
    .Y(_1164_));
 sg13g2_a221oi_1 _4647_ (.B2(_1164_),
    .C1(_0502_),
    .B1(_1159_),
    .A1(_0499_),
    .Y(_1165_),
    .A2(_0500_));
 sg13g2_buf_2 _4648_ (.A(_1165_),
    .X(_1166_));
 sg13g2_a21o_1 _4649_ (.A2(_1166_),
    .A1(net173),
    .B1(_2657_),
    .X(_1167_));
 sg13g2_buf_2 _4650_ (.A(_1167_),
    .X(_1168_));
 sg13g2_nand2_1 _4651_ (.Y(_1169_),
    .A(_3057_),
    .B(_3045_));
 sg13g2_or2_1 _4652_ (.X(_1170_),
    .B(\Pong.datapath.scoreRight[1] ),
    .A(\Pong.datapath.scoreRight[2] ));
 sg13g2_buf_1 _4653_ (.A(_1170_),
    .X(_1171_));
 sg13g2_o21ai_1 _4654_ (.B1(_1160_),
    .Y(_1172_),
    .A1(_1161_),
    .A2(_1171_));
 sg13g2_nand4_1 _4655_ (.B(net32),
    .C(_0501_),
    .A(_0486_),
    .Y(_1173_),
    .D(_1172_));
 sg13g2_nor2_2 _4656_ (.A(_1169_),
    .B(_1173_),
    .Y(_1174_));
 sg13g2_buf_1 _4657_ (.A(\Pong.datapath.scoreLeft[0] ),
    .X(_1175_));
 sg13g2_inv_1 _4658_ (.Y(_1176_),
    .A(_1175_));
 sg13g2_inv_1 _4659_ (.Y(_1177_),
    .A(net172));
 sg13g2_a21oi_1 _4660_ (.A1(_1176_),
    .A2(_1158_),
    .Y(_1178_),
    .B1(_1177_));
 sg13g2_nor3_2 _4661_ (.A(_0502_),
    .B(_0500_),
    .C(_1178_),
    .Y(_1179_));
 sg13g2_o21ai_1 _4662_ (.B1(net173),
    .Y(_1180_),
    .A1(_1174_),
    .A2(_1179_));
 sg13g2_nor2b_1 _4663_ (.A(_1168_),
    .B_N(_1180_),
    .Y(_1181_));
 sg13g2_nand2_1 _4664_ (.Y(_1182_),
    .A(_0081_),
    .B(_1181_));
 sg13g2_buf_2 _4665_ (.A(_1182_),
    .X(_1183_));
 sg13g2_a21oi_1 _4666_ (.A1(_1150_),
    .A2(_1153_),
    .Y(_0242_),
    .B1(_1183_));
 sg13g2_inv_1 _4667_ (.Y(_1184_),
    .A(_1151_));
 sg13g2_inv_1 _4668_ (.Y(_1185_),
    .A(net150));
 sg13g2_buf_1 _4669_ (.A(\Pong.datapath.NES_activity_Left[3] ),
    .X(_1186_));
 sg13g2_buf_1 _4670_ (.A(_1186_),
    .X(_1187_));
 sg13g2_o21ai_1 _4671_ (.B1(net183),
    .Y(_1188_),
    .A1(net155),
    .A2(net180));
 sg13g2_o21ai_1 _4672_ (.B1(_2938_),
    .Y(_1189_),
    .A1(_3007_),
    .A2(_1188_));
 sg13g2_buf_1 _4673_ (.A(_2907_),
    .X(_1190_));
 sg13g2_nand2b_1 _4674_ (.Y(_1191_),
    .B(net133),
    .A_N(_2990_));
 sg13g2_a21oi_1 _4675_ (.A1(_2959_),
    .A2(_1189_),
    .Y(_1192_),
    .B1(_1191_));
 sg13g2_inv_1 _4676_ (.Y(_1193_),
    .A(net182));
 sg13g2_o21ai_1 _4677_ (.B1(net184),
    .Y(_1194_),
    .A1(_2903_),
    .A2(net180));
 sg13g2_buf_2 _4678_ (.A(_1194_),
    .X(_1195_));
 sg13g2_and3_1 _4679_ (.X(_1196_),
    .A(_1193_),
    .B(_2909_),
    .C(_1195_));
 sg13g2_buf_1 _4680_ (.A(_1196_),
    .X(_1197_));
 sg13g2_xor2_1 _4681_ (.B(_1197_),
    .A(net153),
    .X(_1198_));
 sg13g2_nand2b_1 _4682_ (.Y(_1199_),
    .B(_2921_),
    .A_N(net154));
 sg13g2_inv_1 _4683_ (.Y(_1200_),
    .A(net183));
 sg13g2_nand3_1 _4684_ (.B(_1200_),
    .C(_1195_),
    .A(_2990_),
    .Y(_1201_));
 sg13g2_nand2b_1 _4685_ (.Y(_1202_),
    .B(net151),
    .A_N(_2990_));
 sg13g2_nand2b_1 _4686_ (.Y(_1203_),
    .B(_2959_),
    .A_N(net133));
 sg13g2_a21oi_1 _4687_ (.A1(_1201_),
    .A2(_1202_),
    .Y(_1204_),
    .B1(_1203_));
 sg13g2_or4_1 _4688_ (.A(_1192_),
    .B(_1198_),
    .C(_1199_),
    .D(_1204_),
    .X(_1205_));
 sg13g2_buf_1 _4689_ (.A(_1205_),
    .X(_1206_));
 sg13g2_o21ai_1 _4690_ (.B1(_2959_),
    .Y(_1207_),
    .A1(_2908_),
    .A2(_1195_));
 sg13g2_or4_1 _4691_ (.A(net154),
    .B(net133),
    .C(_2997_),
    .D(_1207_),
    .X(_1208_));
 sg13g2_buf_1 _4692_ (.A(_1208_),
    .X(_1209_));
 sg13g2_xor2_1 _4693_ (.B(_1209_),
    .A(net179),
    .X(_1210_));
 sg13g2_nor2_2 _4694_ (.A(_1206_),
    .B(_1210_),
    .Y(_1211_));
 sg13g2_inv_1 _4695_ (.Y(_1212_),
    .A(\Pong.datapath.NES_activity_Left[2] ));
 sg13g2_and2_1 _4696_ (.A(_2903_),
    .B(net180),
    .X(_1213_));
 sg13g2_buf_1 _4697_ (.A(_0084_),
    .X(_1214_));
 sg13g2_nand3_1 _4698_ (.B(net180),
    .C(net168),
    .A(net155),
    .Y(_1215_));
 sg13g2_mux2_1 _4699_ (.A0(_1213_),
    .A1(_1215_),
    .S(net184),
    .X(_1216_));
 sg13g2_a21o_1 _4700_ (.A2(net180),
    .A1(_2903_),
    .B1(net184),
    .X(_1217_));
 sg13g2_nor3_1 _4701_ (.A(_3017_),
    .B(net168),
    .C(_1217_),
    .Y(_1218_));
 sg13g2_a21o_1 _4702_ (.A2(_1216_),
    .A1(_3017_),
    .B1(_1218_),
    .X(_1219_));
 sg13g2_nand3_1 _4703_ (.B(_2903_),
    .C(net180),
    .A(net184),
    .Y(_1220_));
 sg13g2_buf_1 _4704_ (.A(_1220_),
    .X(_1221_));
 sg13g2_a21oi_1 _4705_ (.A1(_1217_),
    .A2(_1221_),
    .Y(_1222_),
    .B1(net168));
 sg13g2_nor3_1 _4706_ (.A(_2937_),
    .B(_3017_),
    .C(_1222_),
    .Y(_1223_));
 sg13g2_a21oi_1 _4707_ (.A1(_2937_),
    .A2(_1219_),
    .Y(_1224_),
    .B1(_1223_));
 sg13g2_nand4_1 _4708_ (.B(net133),
    .C(net183),
    .A(net182),
    .Y(_1225_),
    .D(_1217_));
 sg13g2_nor2_1 _4709_ (.A(_0075_),
    .B(_1225_),
    .Y(_1226_));
 sg13g2_a21oi_2 _4710_ (.B1(_2901_),
    .Y(_1227_),
    .A2(_2945_),
    .A1(_2903_));
 sg13g2_nor2_2 _4711_ (.A(_2986_),
    .B(_1227_),
    .Y(_1228_));
 sg13g2_nor3_1 _4712_ (.A(net182),
    .B(_3006_),
    .C(_1228_),
    .Y(_1229_));
 sg13g2_nor2_1 _4713_ (.A(_1226_),
    .B(_1229_),
    .Y(_1230_));
 sg13g2_nand4_1 _4714_ (.B(net182),
    .C(_2907_),
    .A(_2911_),
    .Y(_1231_),
    .D(net183));
 sg13g2_buf_1 _4715_ (.A(_1231_),
    .X(_1232_));
 sg13g2_a21o_1 _4716_ (.A2(_1227_),
    .A1(net168),
    .B1(_1232_),
    .X(_1233_));
 sg13g2_nand2_1 _4717_ (.Y(_1234_),
    .A(_2904_),
    .B(net180));
 sg13g2_o21ai_1 _4718_ (.B1(net168),
    .Y(_1235_),
    .A1(net156),
    .A2(_1234_));
 sg13g2_nor2_1 _4719_ (.A(_2917_),
    .B(_1232_),
    .Y(_1236_));
 sg13g2_a22oi_1 _4720_ (.Y(_1237_),
    .B1(_1235_),
    .B2(_1236_),
    .A2(_1233_),
    .A1(_2918_));
 sg13g2_nand4_1 _4721_ (.B(_2902_),
    .C(net179),
    .A(_2917_),
    .Y(_1238_),
    .D(_1214_));
 sg13g2_or2_1 _4722_ (.X(_1239_),
    .B(_1238_),
    .A(_1232_));
 sg13g2_o21ai_1 _4723_ (.B1(_1239_),
    .Y(_1240_),
    .A1(net179),
    .A2(_1237_));
 sg13g2_o21ai_1 _4724_ (.B1(_1240_),
    .Y(_1241_),
    .A1(_1224_),
    .A2(_1230_));
 sg13g2_and3_1 _4725_ (.X(_1242_),
    .A(_2917_),
    .B(_2911_),
    .C(_2912_));
 sg13g2_buf_1 _4726_ (.A(_1242_),
    .X(_1243_));
 sg13g2_and2_1 _4727_ (.A(\Pong.datapath.leftPaddle[8] ),
    .B(_1243_),
    .X(_1244_));
 sg13g2_a21oi_1 _4728_ (.A1(_1228_),
    .A2(_1244_),
    .Y(_1245_),
    .B1(net181));
 sg13g2_and2_1 _4729_ (.A(_1241_),
    .B(_1245_),
    .X(_1246_));
 sg13g2_nor3_1 _4730_ (.A(_1212_),
    .B(_1186_),
    .C(_1246_),
    .Y(_1247_));
 sg13g2_a21oi_1 _4731_ (.A1(net134),
    .A2(_1211_),
    .Y(_1248_),
    .B1(_1247_));
 sg13g2_nand3_1 _4732_ (.B(_1241_),
    .C(_1245_),
    .A(\Pong.datapath.NES_activity_Left[2] ),
    .Y(_1249_));
 sg13g2_buf_1 _4733_ (.A(_1249_),
    .X(_1250_));
 sg13g2_inv_1 _4734_ (.Y(_1251_),
    .A(_1186_));
 sg13g2_nand2b_1 _4735_ (.Y(_1252_),
    .B(_1251_),
    .A_N(net41));
 sg13g2_buf_2 _4736_ (.A(_1252_),
    .X(_1253_));
 sg13g2_o21ai_1 _4737_ (.B1(_1186_),
    .Y(_1254_),
    .A1(_1206_),
    .A2(_1210_));
 sg13g2_buf_2 _4738_ (.A(_1254_),
    .X(_1255_));
 sg13g2_and2_1 _4739_ (.A(net150),
    .B(_1255_),
    .X(_1256_));
 sg13g2_a22oi_1 _4740_ (.Y(_1257_),
    .B1(_1253_),
    .B2(_1256_),
    .A2(_1248_),
    .A1(_1185_));
 sg13g2_o21ai_1 _4741_ (.B1(_1184_),
    .Y(_1258_),
    .A1(\Pong.datapath.NES_activity_Left[2] ),
    .A2(net134));
 sg13g2_nand3_1 _4742_ (.B(_0081_),
    .C(_1181_),
    .A(_0507_),
    .Y(_1259_));
 sg13g2_a221oi_1 _4743_ (.B2(_0083_),
    .C1(_1259_),
    .B1(_1258_),
    .A1(_1184_),
    .Y(_0243_),
    .A2(_1257_));
 sg13g2_buf_1 _4744_ (.A(_0506_),
    .X(_1260_));
 sg13g2_nor2_1 _4745_ (.A(_1260_),
    .B(_1183_),
    .Y(_1261_));
 sg13g2_nand2b_1 _4746_ (.Y(_1262_),
    .B(net150),
    .A_N(net155));
 sg13g2_nand2b_1 _4747_ (.Y(_1263_),
    .B(net155),
    .A_N(_2946_));
 sg13g2_and2_1 _4748_ (.A(_1262_),
    .B(_1263_),
    .X(_1264_));
 sg13g2_mux2_1 _4749_ (.A0(_1255_),
    .A1(_1253_),
    .S(_1264_),
    .X(_1265_));
 sg13g2_or2_1 _4750_ (.X(_1266_),
    .B(_1265_),
    .A(net135));
 sg13g2_mux2_1 _4751_ (.A0(_1253_),
    .A1(_1255_),
    .S(_1264_),
    .X(_1267_));
 sg13g2_o21ai_1 _4752_ (.B1(_0076_),
    .Y(_1268_),
    .A1(net135),
    .A2(_1267_));
 sg13g2_and3_1 _4753_ (.X(_0244_),
    .A(_1261_),
    .B(_1266_),
    .C(_1268_));
 sg13g2_inv_1 _4754_ (.Y(_1269_),
    .A(_1168_));
 sg13g2_nand2_1 _4755_ (.Y(_1270_),
    .A(_1269_),
    .B(_1180_));
 sg13g2_nor3_2 _4756_ (.A(\Pong.datapath.NES_activity_Right[5] ),
    .B(net132),
    .C(_1270_),
    .Y(_1271_));
 sg13g2_nor2_2 _4757_ (.A(_2904_),
    .B(_2946_),
    .Y(_1272_));
 sg13g2_or2_1 _4758_ (.X(_1273_),
    .B(_1255_),
    .A(_1272_));
 sg13g2_a221oi_1 _4759_ (.B2(_1253_),
    .C1(_1151_),
    .B1(_1273_),
    .A1(_1213_),
    .Y(_1274_),
    .A2(_1255_));
 sg13g2_xnor2_1 _4760_ (.Y(_1275_),
    .A(_2902_),
    .B(_1274_));
 sg13g2_nand2_1 _4761_ (.Y(_0245_),
    .A(_1271_),
    .B(_1275_));
 sg13g2_xor2_1 _4762_ (.B(_1195_),
    .A(_2959_),
    .X(_1276_));
 sg13g2_nor2_1 _4763_ (.A(_1211_),
    .B(_1276_),
    .Y(_1277_));
 sg13g2_a21oi_1 _4764_ (.A1(net151),
    .A2(_1211_),
    .Y(_1278_),
    .B1(_1277_));
 sg13g2_inv_1 _4765_ (.Y(_1279_),
    .A(_1235_));
 sg13g2_nor4_1 _4766_ (.A(_1200_),
    .B(net134),
    .C(_1279_),
    .D(net41),
    .Y(_1280_));
 sg13g2_a21oi_1 _4767_ (.A1(net134),
    .A2(_1278_),
    .Y(_1281_),
    .B1(_1280_));
 sg13g2_nor2_1 _4768_ (.A(_1152_),
    .B(_1281_),
    .Y(_1282_));
 sg13g2_o21ai_1 _4769_ (.B1(_1251_),
    .Y(_1283_),
    .A1(_1279_),
    .A2(_1250_));
 sg13g2_a21oi_1 _4770_ (.A1(_1184_),
    .A2(_1283_),
    .Y(_1284_),
    .B1(net151));
 sg13g2_o21ai_1 _4771_ (.B1(_1271_),
    .Y(_0246_),
    .A1(_1282_),
    .A2(_1284_));
 sg13g2_nor2_1 _4772_ (.A(_1200_),
    .B(_1227_),
    .Y(_1285_));
 sg13g2_xnor2_1 _4773_ (.Y(_1286_),
    .A(_3017_),
    .B(_1285_));
 sg13g2_nand2_1 _4774_ (.Y(_1287_),
    .A(net133),
    .B(net41));
 sg13g2_o21ai_1 _4775_ (.B1(_1287_),
    .Y(_1288_),
    .A1(net41),
    .A2(_1286_));
 sg13g2_nor2_1 _4776_ (.A(_1207_),
    .B(_1255_),
    .Y(_1289_));
 sg13g2_o21ai_1 _4777_ (.B1(_1186_),
    .Y(_1290_),
    .A1(_1207_),
    .A2(_1211_));
 sg13g2_a21oi_1 _4778_ (.A1(_1184_),
    .A2(_1290_),
    .Y(_1291_),
    .B1(net133));
 sg13g2_a21oi_1 _4779_ (.A1(_1190_),
    .A2(_1289_),
    .Y(_1292_),
    .B1(_1291_));
 sg13g2_o21ai_1 _4780_ (.B1(_1292_),
    .Y(_1293_),
    .A1(net134),
    .A2(_1288_));
 sg13g2_nand2_1 _4781_ (.Y(_1294_),
    .A(_1190_),
    .B(net135));
 sg13g2_nand3_1 _4782_ (.B(_1293_),
    .C(_1294_),
    .A(_1271_),
    .Y(_0247_));
 sg13g2_nand2_1 _4783_ (.Y(_1295_),
    .A(net149),
    .B(net41));
 sg13g2_xnor2_1 _4784_ (.Y(_1296_),
    .A(net152),
    .B(_1228_));
 sg13g2_nand2b_1 _4785_ (.Y(_1297_),
    .B(_1296_),
    .A_N(net41));
 sg13g2_nand3_1 _4786_ (.B(_1295_),
    .C(_1297_),
    .A(_1251_),
    .Y(_1298_));
 sg13g2_nand2_1 _4787_ (.Y(_1299_),
    .A(net104),
    .B(_1195_));
 sg13g2_nor2_1 _4788_ (.A(_1299_),
    .B(_1255_),
    .Y(_1300_));
 sg13g2_o21ai_1 _4789_ (.B1(net134),
    .Y(_1301_),
    .A1(_1299_),
    .A2(_1211_));
 sg13g2_a21oi_1 _4790_ (.A1(_1184_),
    .A2(_1301_),
    .Y(_1302_),
    .B1(net149));
 sg13g2_a21oi_1 _4791_ (.A1(_2991_),
    .A2(_1300_),
    .Y(_1303_),
    .B1(_1302_));
 sg13g2_a221oi_1 _4792_ (.B2(_1303_),
    .C1(_1259_),
    .B1(_1298_),
    .A1(_2991_),
    .Y(_0248_),
    .A2(_1152_));
 sg13g2_xnor2_1 _4793_ (.Y(_1304_),
    .A(_3006_),
    .B(_1225_));
 sg13g2_nand2_1 _4794_ (.Y(_1305_),
    .A(net153),
    .B(_1197_));
 sg13g2_or2_1 _4795_ (.X(_1306_),
    .B(_1255_),
    .A(_1305_));
 sg13g2_o21ai_1 _4796_ (.B1(_1306_),
    .Y(_1307_),
    .A1(_1253_),
    .A2(_1304_));
 sg13g2_and2_1 _4797_ (.A(_1184_),
    .B(_1307_),
    .X(_1308_));
 sg13g2_nand2_1 _4798_ (.Y(_1309_),
    .A(net134),
    .B(_1197_));
 sg13g2_a21oi_1 _4799_ (.A1(_1253_),
    .A2(_1309_),
    .Y(_1310_),
    .B1(net135));
 sg13g2_nor2_1 _4800_ (.A(net153),
    .B(_1310_),
    .Y(_1311_));
 sg13g2_o21ai_1 _4801_ (.B1(_1271_),
    .Y(_0249_),
    .A1(_1308_),
    .A2(_1311_));
 sg13g2_nand3b_1 _4802_ (.B(net134),
    .C(_1197_),
    .Y(_1312_),
    .A_N(_2930_));
 sg13g2_or4_1 _4803_ (.A(_1186_),
    .B(_1232_),
    .C(_1279_),
    .D(net41),
    .X(_1313_));
 sg13g2_a21oi_1 _4804_ (.A1(_1312_),
    .A2(_1313_),
    .Y(_1314_),
    .B1(net135));
 sg13g2_xnor2_1 _4805_ (.Y(_1315_),
    .A(_2918_),
    .B(_1314_));
 sg13g2_nand2_1 _4806_ (.Y(_0250_),
    .A(_1271_),
    .B(_1315_));
 sg13g2_nor2_1 _4807_ (.A(net179),
    .B(net135),
    .Y(_1316_));
 sg13g2_nand4_1 _4808_ (.B(_1228_),
    .C(_1243_),
    .A(\Pong.datapath.NES_activity_Left[2] ),
    .Y(_1317_),
    .D(_1246_));
 sg13g2_mux2_1 _4809_ (.A0(_1316_),
    .A1(net179),
    .S(_1317_),
    .X(_1318_));
 sg13g2_nor4_1 _4810_ (.A(net179),
    .B(_1151_),
    .C(_1251_),
    .D(_1209_),
    .Y(_1319_));
 sg13g2_a21o_1 _4811_ (.A2(_1209_),
    .A1(_1187_),
    .B1(_1151_),
    .X(_1320_));
 sg13g2_a22oi_1 _4812_ (.Y(_1321_),
    .B1(_1320_),
    .B2(_2984_),
    .A2(_1319_),
    .A1(_1206_));
 sg13g2_nand2_1 _4813_ (.Y(_1322_),
    .A(_1261_),
    .B(_1321_));
 sg13g2_a21oi_1 _4814_ (.A1(_1251_),
    .A2(_1318_),
    .Y(_0251_),
    .B1(_1322_));
 sg13g2_a21oi_1 _4815_ (.A1(_1251_),
    .A2(net41),
    .Y(_1323_),
    .B1(net135));
 sg13g2_nand3_1 _4816_ (.B(_3001_),
    .C(_1195_),
    .A(net104),
    .Y(_1324_));
 sg13g2_nor3_1 _4817_ (.A(_3063_),
    .B(_1151_),
    .C(_1324_),
    .Y(_1325_));
 sg13g2_a21oi_1 _4818_ (.A1(_3063_),
    .A2(_1324_),
    .Y(_1326_),
    .B1(_1325_));
 sg13g2_nand2b_1 _4819_ (.Y(_1327_),
    .B(_1187_),
    .A_N(_1326_));
 sg13g2_o21ai_1 _4820_ (.B1(_1327_),
    .Y(_1328_),
    .A1(_2921_),
    .A2(_1323_));
 sg13g2_and2_1 _4821_ (.A(_1261_),
    .B(_1328_),
    .X(_0252_));
 sg13g2_and2_1 _4822_ (.A(net139),
    .B(_0048_),
    .X(_0253_));
 sg13g2_and2_1 _4823_ (.A(net139),
    .B(_0049_),
    .X(_0254_));
 sg13g2_and2_1 _4824_ (.A(net139),
    .B(_0050_),
    .X(_0255_));
 sg13g2_and2_1 _4825_ (.A(net139),
    .B(_0051_),
    .X(_0256_));
 sg13g2_and2_1 _4826_ (.A(net139),
    .B(_0052_),
    .X(_0257_));
 sg13g2_and2_1 _4827_ (.A(_0628_),
    .B(_0053_),
    .X(_0258_));
 sg13g2_and2_1 _4828_ (.A(_0628_),
    .B(_0054_),
    .X(_0259_));
 sg13g2_and2_1 _4829_ (.A(_2717_),
    .B(_0055_),
    .X(_0260_));
 sg13g2_nand2_1 _4830_ (.Y(_1329_),
    .A(_0507_),
    .B(net143));
 sg13g2_or2_1 _4831_ (.X(_1330_),
    .B(net148),
    .A(net142));
 sg13g2_buf_1 _4832_ (.A(_1330_),
    .X(_1331_));
 sg13g2_o21ai_1 _4833_ (.B1(net147),
    .Y(_1332_),
    .A1(net177),
    .A2(net176));
 sg13g2_buf_2 _4834_ (.A(_1332_),
    .X(_1333_));
 sg13g2_nor2_1 _4835_ (.A(net146),
    .B(_1333_),
    .Y(_1334_));
 sg13g2_inv_1 _4836_ (.Y(_1335_),
    .A(_0314_));
 sg13g2_nand2_1 _4837_ (.Y(_1336_),
    .A(_1335_),
    .B(net144));
 sg13g2_nor4_1 _4838_ (.A(net140),
    .B(_1331_),
    .C(_1334_),
    .D(_1336_),
    .Y(_1337_));
 sg13g2_xnor2_1 _4839_ (.Y(_1338_),
    .A(_0361_),
    .B(_1337_));
 sg13g2_or2_1 _4840_ (.X(_1339_),
    .B(net176),
    .A(net177));
 sg13g2_buf_1 _4841_ (.A(_1339_),
    .X(_1340_));
 sg13g2_nand3_1 _4842_ (.B(net146),
    .C(_1340_),
    .A(net103),
    .Y(_1341_));
 sg13g2_a21oi_1 _4843_ (.A1(_0413_),
    .A2(_1341_),
    .Y(_1342_),
    .B1(_0345_));
 sg13g2_nand2b_1 _4844_ (.Y(_1343_),
    .B(net178),
    .A_N(_0057_));
 sg13g2_nor2b_1 _4845_ (.A(net140),
    .B_N(_0373_),
    .Y(_1344_));
 sg13g2_o21ai_1 _4846_ (.B1(_1344_),
    .Y(_1345_),
    .A1(_1342_),
    .A2(_1343_));
 sg13g2_nand2_2 _4847_ (.Y(_1346_),
    .A(net100),
    .B(_1333_));
 sg13g2_o21ai_1 _4848_ (.B1(_0365_),
    .Y(_1347_),
    .A1(_0382_),
    .A2(_1346_));
 sg13g2_o21ai_1 _4849_ (.B1(_1347_),
    .Y(_1348_),
    .A1(_1331_),
    .A2(_1346_));
 sg13g2_inv_2 _4850_ (.Y(_1349_),
    .A(net146));
 sg13g2_nand3_1 _4851_ (.B(_1349_),
    .C(_1333_),
    .A(net175),
    .Y(_1350_));
 sg13g2_nand2b_1 _4852_ (.Y(_1351_),
    .B(net99),
    .A_N(_0383_));
 sg13g2_a21oi_1 _4853_ (.A1(_1350_),
    .A2(_1351_),
    .Y(_1352_),
    .B1(_1336_));
 sg13g2_nor4_2 _4854_ (.A(_1338_),
    .B(_1345_),
    .C(_1348_),
    .Y(_1353_),
    .D(_1352_));
 sg13g2_buf_1 _4855_ (.A(\Pong.datapath.NES_activity_Right[3] ),
    .X(_1354_));
 sg13g2_nand2b_1 _4856_ (.Y(_1355_),
    .B(_1354_),
    .A_N(_1353_));
 sg13g2_nand2_1 _4857_ (.Y(_1356_),
    .A(\Pong.datapath.rightPaddle[4] ),
    .B(_0317_));
 sg13g2_buf_1 _4858_ (.A(_1356_),
    .X(_1357_));
 sg13g2_a21oi_2 _4859_ (.B1(_0315_),
    .Y(_1358_),
    .A2(net176),
    .A1(net177));
 sg13g2_nand3_1 _4860_ (.B(_0364_),
    .C(_0311_),
    .A(_0363_),
    .Y(_1359_));
 sg13g2_nor3_1 _4861_ (.A(net95),
    .B(_1358_),
    .C(_1359_),
    .Y(_1360_));
 sg13g2_xnor2_1 _4862_ (.Y(_1361_),
    .A(_0361_),
    .B(_1360_));
 sg13g2_buf_2 _4863_ (.A(_0082_),
    .X(_1362_));
 sg13g2_nand3b_1 _4864_ (.B(net177),
    .C(net176),
    .Y(_1363_),
    .A_N(_0315_));
 sg13g2_and2_1 _4865_ (.A(_1362_),
    .B(_1363_),
    .X(_1364_));
 sg13g2_nor3_1 _4866_ (.A(net95),
    .B(_0404_),
    .C(_1364_),
    .Y(_1365_));
 sg13g2_xnor2_1 _4867_ (.Y(_1366_),
    .A(_0062_),
    .B(_1365_));
 sg13g2_and2_1 _4868_ (.A(_1361_),
    .B(_1366_),
    .X(_1367_));
 sg13g2_inv_1 _4869_ (.Y(_1368_),
    .A(_1362_));
 sg13g2_nand2_2 _4870_ (.Y(_1369_),
    .A(_0318_),
    .B(_0347_));
 sg13g2_o21ai_1 _4871_ (.B1(_0316_),
    .Y(_1370_),
    .A1(_1368_),
    .A2(_1369_));
 sg13g2_nand3_1 _4872_ (.B(_1363_),
    .C(_1370_),
    .A(_0323_),
    .Y(_1371_));
 sg13g2_nand2b_1 _4873_ (.Y(_1372_),
    .B(_1369_),
    .A_N(net147));
 sg13g2_o21ai_1 _4874_ (.B1(_0322_),
    .Y(_1373_),
    .A1(_1362_),
    .A2(_1372_));
 sg13g2_and3_1 _4875_ (.X(_1374_),
    .A(_0325_),
    .B(_1371_),
    .C(_1373_));
 sg13g2_nand3_1 _4876_ (.B(net177),
    .C(\Pong.datapath.rightPaddle[0] ),
    .A(_0315_),
    .Y(_1375_));
 sg13g2_buf_2 _4877_ (.A(_1375_),
    .X(_1376_));
 sg13g2_a21oi_1 _4878_ (.A1(_1372_),
    .A2(_1376_),
    .Y(_1377_),
    .B1(_1362_));
 sg13g2_nor3_1 _4879_ (.A(_0325_),
    .B(_0323_),
    .C(_1377_),
    .Y(_1378_));
 sg13g2_nor2_1 _4880_ (.A(net95),
    .B(_1358_),
    .Y(_1379_));
 sg13g2_nand2_1 _4881_ (.Y(_1380_),
    .A(_0312_),
    .B(_1379_));
 sg13g2_nor2b_1 _4882_ (.A(_0312_),
    .B_N(_0381_),
    .Y(_1381_));
 sg13g2_o21ai_1 _4883_ (.B1(_1381_),
    .Y(_1382_),
    .A1(net95),
    .A2(_1358_));
 sg13g2_o21ai_1 _4884_ (.B1(_1382_),
    .Y(_1383_),
    .A1(_0381_),
    .A2(_1380_));
 sg13g2_o21ai_1 _4885_ (.B1(_1383_),
    .Y(_1384_),
    .A1(_1374_),
    .A2(_1378_));
 sg13g2_and4_1 _4886_ (.A(_0370_),
    .B(_0363_),
    .C(_0364_),
    .D(_0311_),
    .X(_1385_));
 sg13g2_buf_1 _4887_ (.A(_1385_),
    .X(_1386_));
 sg13g2_nand2b_1 _4888_ (.Y(_1387_),
    .B(\Pong.datapath.NES_activity_Right[2] ),
    .A_N(_0409_));
 sg13g2_a221oi_1 _4889_ (.B2(_1379_),
    .C1(_1387_),
    .B1(_1386_),
    .A1(_1367_),
    .Y(_1388_),
    .A2(_1384_));
 sg13g2_buf_2 _4890_ (.A(_1388_),
    .X(_1389_));
 sg13g2_nand2b_1 _4891_ (.Y(_1390_),
    .B(_1389_),
    .A_N(_1354_));
 sg13g2_buf_2 _4892_ (.A(_1390_),
    .X(_1391_));
 sg13g2_a21oi_1 _4893_ (.A1(_1355_),
    .A2(_1391_),
    .Y(_1392_),
    .B1(_1149_));
 sg13g2_mux2_1 _4894_ (.A0(_1329_),
    .A1(net143),
    .S(_1392_),
    .X(_1393_));
 sg13g2_nor2_1 _4895_ (.A(_1183_),
    .B(_1393_),
    .Y(_0261_));
 sg13g2_buf_1 _4896_ (.A(_1149_),
    .X(_1394_));
 sg13g2_mux2_1 _4897_ (.A0(_1355_),
    .A1(_1391_),
    .S(_0348_),
    .X(_1395_));
 sg13g2_nor2_1 _4898_ (.A(_1260_),
    .B(_0342_),
    .Y(_1396_));
 sg13g2_o21ai_1 _4899_ (.B1(_1396_),
    .Y(_1397_),
    .A1(_1394_),
    .A2(_1395_));
 sg13g2_xor2_1 _4900_ (.B(_0348_),
    .A(_0327_),
    .X(_1398_));
 sg13g2_mux2_1 _4901_ (.A0(_1355_),
    .A1(_1391_),
    .S(_1398_),
    .X(_1399_));
 sg13g2_or2_1 _4902_ (.X(_1400_),
    .B(_1399_),
    .A(net131));
 sg13g2_a21oi_1 _4903_ (.A1(_1397_),
    .A2(_1400_),
    .Y(_0262_),
    .B1(_1183_));
 sg13g2_nor3_1 _4904_ (.A(net132),
    .B(net103),
    .C(_1150_),
    .Y(_1401_));
 sg13g2_and2_1 _4905_ (.A(_0326_),
    .B(net176),
    .X(_1402_));
 sg13g2_mux2_1 _4906_ (.A0(_0507_),
    .A1(_1402_),
    .S(_1389_),
    .X(_1403_));
 sg13g2_nand2b_1 _4907_ (.Y(_1404_),
    .B(_1403_),
    .A_N(net103));
 sg13g2_and2_1 _4908_ (.A(_0324_),
    .B(_1369_),
    .X(_1405_));
 sg13g2_buf_8 _4909_ (.A(_1389_),
    .X(_1406_));
 sg13g2_buf_1 _4910_ (.A(_1354_),
    .X(_1407_));
 sg13g2_a21oi_1 _4911_ (.A1(_1405_),
    .A2(_1406_),
    .Y(_1408_),
    .B1(net130));
 sg13g2_mux2_1 _4912_ (.A0(_1340_),
    .A1(_0506_),
    .S(_1353_),
    .X(_1409_));
 sg13g2_nor2_1 _4913_ (.A(net103),
    .B(_1409_),
    .Y(_1410_));
 sg13g2_buf_1 _4914_ (.A(_1353_),
    .X(_1411_));
 sg13g2_nor2_1 _4915_ (.A(_1333_),
    .B(net40),
    .Y(_1412_));
 sg13g2_nor2_1 _4916_ (.A(_1410_),
    .B(_1412_),
    .Y(_1413_));
 sg13g2_a221oi_1 _4917_ (.B2(net130),
    .C1(net131),
    .B1(_1413_),
    .A1(_1404_),
    .Y(_1414_),
    .A2(_1408_));
 sg13g2_nor2_2 _4918_ (.A(\Pong.datapath.NES_activity_Right[5] ),
    .B(_1270_),
    .Y(_1415_));
 sg13g2_o21ai_1 _4919_ (.B1(_1415_),
    .Y(_0263_),
    .A1(_1401_),
    .A2(_1414_));
 sg13g2_nor2_1 _4920_ (.A(_0506_),
    .B(net99),
    .Y(_1416_));
 sg13g2_and2_1 _4921_ (.A(net131),
    .B(_1416_),
    .X(_1417_));
 sg13g2_mux2_1 _4922_ (.A0(_0507_),
    .A1(_1364_),
    .S(_1406_),
    .X(_1418_));
 sg13g2_nand2_1 _4923_ (.Y(_1419_),
    .A(_1349_),
    .B(_1418_));
 sg13g2_nor2_1 _4924_ (.A(_1349_),
    .B(_1364_),
    .Y(_1420_));
 sg13g2_a21oi_1 _4925_ (.A1(net26),
    .A2(_1420_),
    .Y(_1421_),
    .B1(_1407_));
 sg13g2_xnor2_1 _4926_ (.Y(_1422_),
    .A(net144),
    .B(_1333_));
 sg13g2_nor2_1 _4927_ (.A(net40),
    .B(_1422_),
    .Y(_1423_));
 sg13g2_a21oi_1 _4928_ (.A1(net40),
    .A2(_1416_),
    .Y(_1424_),
    .B1(_1423_));
 sg13g2_a221oi_1 _4929_ (.B2(net130),
    .C1(_1394_),
    .B1(_1424_),
    .A1(_1419_),
    .Y(_1425_),
    .A2(_1421_));
 sg13g2_o21ai_1 _4930_ (.B1(_1415_),
    .Y(_0264_),
    .A1(_1417_),
    .A2(_1425_));
 sg13g2_o21ai_1 _4931_ (.B1(net144),
    .Y(_1426_),
    .A1(_0440_),
    .A2(_1333_));
 sg13g2_nor2_1 _4932_ (.A(_1353_),
    .B(_1426_),
    .Y(_1427_));
 sg13g2_a21oi_1 _4933_ (.A1(net132),
    .A2(_1411_),
    .Y(_1428_),
    .B1(_1427_));
 sg13g2_o21ai_1 _4934_ (.B1(net178),
    .Y(_1429_),
    .A1(_1411_),
    .A2(_1426_));
 sg13g2_o21ai_1 _4935_ (.B1(_1429_),
    .Y(_1430_),
    .A1(_0314_),
    .A2(_1428_));
 sg13g2_nor2_1 _4936_ (.A(_1349_),
    .B(_1358_),
    .Y(_1431_));
 sg13g2_xnor2_1 _4937_ (.Y(_1432_),
    .A(_0322_),
    .B(_1431_));
 sg13g2_inv_1 _4938_ (.Y(_1433_),
    .A(_1391_));
 sg13g2_a22oi_1 _4939_ (.Y(_1434_),
    .B1(_1432_),
    .B2(_1433_),
    .A2(_1430_),
    .A1(_1407_));
 sg13g2_o21ai_1 _4940_ (.B1(_1150_),
    .Y(_1435_),
    .A1(_1354_),
    .A2(net26));
 sg13g2_o21ai_1 _4941_ (.B1(_1435_),
    .Y(_1436_),
    .A1(net132),
    .A2(net178));
 sg13g2_and2_1 _4942_ (.A(_1415_),
    .B(_1436_),
    .X(_1437_));
 sg13g2_o21ai_1 _4943_ (.B1(_1437_),
    .Y(_0265_),
    .A1(net131),
    .A2(_1434_));
 sg13g2_nor2_1 _4944_ (.A(_0506_),
    .B(_0313_),
    .Y(_1438_));
 sg13g2_nand2_1 _4945_ (.Y(_1439_),
    .A(net131),
    .B(_1438_));
 sg13g2_mux2_1 _4946_ (.A0(_0506_),
    .A1(_1379_),
    .S(net26),
    .X(_1440_));
 sg13g2_nor3_1 _4947_ (.A(_0382_),
    .B(_1357_),
    .C(_1358_),
    .Y(_1441_));
 sg13g2_a21oi_1 _4948_ (.A1(net26),
    .A2(_1441_),
    .Y(_1442_),
    .B1(_1354_));
 sg13g2_o21ai_1 _4949_ (.B1(_1442_),
    .Y(_1443_),
    .A1(_0313_),
    .A2(_1440_));
 sg13g2_xnor2_1 _4950_ (.Y(_1444_),
    .A(_0383_),
    .B(_1346_));
 sg13g2_nor2_1 _4951_ (.A(net40),
    .B(_1444_),
    .Y(_1445_));
 sg13g2_a21oi_1 _4952_ (.A1(net40),
    .A2(_1438_),
    .Y(_1446_),
    .B1(_1445_));
 sg13g2_nand2_1 _4953_ (.Y(_1447_),
    .A(net130),
    .B(_1446_));
 sg13g2_nand3_1 _4954_ (.B(_1443_),
    .C(_1447_),
    .A(_1150_),
    .Y(_1448_));
 sg13g2_a21oi_1 _4955_ (.A1(_1439_),
    .A2(_1448_),
    .Y(_0266_),
    .B1(_1183_));
 sg13g2_nor2_1 _4956_ (.A(net132),
    .B(_0365_),
    .Y(_1449_));
 sg13g2_xor2_1 _4957_ (.B(_1380_),
    .A(_0381_),
    .X(_1450_));
 sg13g2_nand2_1 _4958_ (.Y(_1451_),
    .A(net26),
    .B(_1450_));
 sg13g2_o21ai_1 _4959_ (.B1(_1451_),
    .Y(_1452_),
    .A1(net26),
    .A2(_1449_));
 sg13g2_inv_1 _4960_ (.Y(_1453_),
    .A(_1348_));
 sg13g2_a21oi_1 _4961_ (.A1(net130),
    .A2(_1453_),
    .Y(_1454_),
    .B1(net131));
 sg13g2_o21ai_1 _4962_ (.B1(_1454_),
    .Y(_1455_),
    .A1(net130),
    .A2(_1452_));
 sg13g2_o21ai_1 _4963_ (.B1(net40),
    .Y(_1456_),
    .A1(_1391_),
    .A2(_1450_));
 sg13g2_a21o_1 _4964_ (.A2(_1456_),
    .A1(_1150_),
    .B1(_1449_),
    .X(_1457_));
 sg13g2_nand3_1 _4965_ (.B(_1455_),
    .C(_1457_),
    .A(_1415_),
    .Y(_0267_));
 sg13g2_nor2_1 _4966_ (.A(_1331_),
    .B(_1346_),
    .Y(_1458_));
 sg13g2_or2_1 _4967_ (.X(_1459_),
    .B(_1458_),
    .A(net140));
 sg13g2_a21oi_1 _4968_ (.A1(net132),
    .A2(net40),
    .Y(_1460_),
    .B1(_1459_));
 sg13g2_a21oi_1 _4969_ (.A1(net140),
    .A2(_1458_),
    .Y(_1461_),
    .B1(_1460_));
 sg13g2_a22oi_1 _4970_ (.Y(_1462_),
    .B1(_1461_),
    .B2(net130),
    .A2(_1433_),
    .A1(_1366_));
 sg13g2_o21ai_1 _4971_ (.B1(_1435_),
    .Y(_1463_),
    .A1(net132),
    .A2(_0400_));
 sg13g2_and2_1 _4972_ (.A(_1415_),
    .B(_1463_),
    .X(_1464_));
 sg13g2_o21ai_1 _4973_ (.B1(_1464_),
    .Y(_0268_),
    .A1(net131),
    .A2(_1462_));
 sg13g2_nor2b_1 _4974_ (.A(_0506_),
    .B_N(net141),
    .Y(_1465_));
 sg13g2_nor3_1 _4975_ (.A(_1345_),
    .B(_1348_),
    .C(_1352_),
    .Y(_1466_));
 sg13g2_nand2b_1 _4976_ (.Y(_1467_),
    .B(_1354_),
    .A_N(_1338_));
 sg13g2_a22oi_1 _4977_ (.Y(_1468_),
    .B1(_1467_),
    .B2(_1150_),
    .A2(_1465_),
    .A1(_1466_));
 sg13g2_o21ai_1 _4978_ (.B1(_1150_),
    .Y(_1469_),
    .A1(net26),
    .A2(_1468_));
 sg13g2_a21oi_1 _4979_ (.A1(_1361_),
    .A2(net26),
    .Y(_1470_),
    .B1(net130));
 sg13g2_nor2_1 _4980_ (.A(_1468_),
    .B(_1470_),
    .Y(_1471_));
 sg13g2_a21oi_1 _4981_ (.A1(_1465_),
    .A2(_1469_),
    .Y(_1472_),
    .B1(_1471_));
 sg13g2_nor2_1 _4982_ (.A(_1183_),
    .B(_1472_),
    .Y(_0269_));
 sg13g2_nand2_1 _4983_ (.Y(_1473_),
    .A(_1150_),
    .B(_1354_));
 sg13g2_nand3_1 _4984_ (.B(net100),
    .C(_1333_),
    .A(_0371_),
    .Y(_1474_));
 sg13g2_xnor2_1 _4985_ (.Y(_1475_),
    .A(_0373_),
    .B(_1474_));
 sg13g2_nor2b_1 _4986_ (.A(net132),
    .B_N(_0409_),
    .Y(_1476_));
 sg13g2_o21ai_1 _4987_ (.B1(_1476_),
    .Y(_1477_),
    .A1(net40),
    .A2(_1473_));
 sg13g2_o21ai_1 _4988_ (.B1(_1477_),
    .Y(_1478_),
    .A1(_1473_),
    .A2(_1475_));
 sg13g2_nor2b_1 _4989_ (.A(_1183_),
    .B_N(_1478_),
    .Y(_0270_));
 sg13g2_o21ai_1 _4990_ (.B1(net173),
    .Y(_1479_),
    .A1(_1166_),
    .A2(_1179_));
 sg13g2_nor2b_1 _4991_ (.A(_0506_),
    .B_N(_0081_),
    .Y(_1480_));
 sg13g2_buf_1 _4992_ (.A(_1480_),
    .X(_1481_));
 sg13g2_nand3_1 _4993_ (.B(_1479_),
    .C(_1481_),
    .A(net169),
    .Y(_1482_));
 sg13g2_nand2_1 _4994_ (.Y(_1483_),
    .A(net173),
    .B(_1179_));
 sg13g2_or3_1 _4995_ (.A(net169),
    .B(_1166_),
    .C(_1483_),
    .X(_1484_));
 sg13g2_a21oi_1 _4996_ (.A1(_1482_),
    .A2(_1484_),
    .Y(_0271_),
    .B1(net138));
 sg13g2_nand2_1 _4997_ (.Y(_1485_),
    .A(_1481_),
    .B(_1483_));
 sg13g2_o21ai_1 _4998_ (.B1(_1485_),
    .Y(_1486_),
    .A1(_1175_),
    .A2(_1483_));
 sg13g2_nor2_1 _4999_ (.A(net171),
    .B(_1176_),
    .Y(_1487_));
 sg13g2_and2_1 _5000_ (.A(net173),
    .B(_1179_),
    .X(_1488_));
 sg13g2_buf_1 _5001_ (.A(_1488_),
    .X(_1489_));
 sg13g2_a22oi_1 _5002_ (.Y(_1490_),
    .B1(_1487_),
    .B2(_1489_),
    .A2(_1486_),
    .A1(net171));
 sg13g2_nor2_1 _5003_ (.A(_1168_),
    .B(_1490_),
    .Y(_0272_));
 sg13g2_buf_1 _5004_ (.A(_1156_),
    .X(_1491_));
 sg13g2_nand2_1 _5005_ (.Y(_1492_),
    .A(net171),
    .B(net169));
 sg13g2_nor2_1 _5006_ (.A(_1483_),
    .B(_1492_),
    .Y(_1493_));
 sg13g2_o21ai_1 _5007_ (.B1(_1269_),
    .Y(_1494_),
    .A1(net129),
    .A2(_1493_));
 sg13g2_nand2_1 _5008_ (.Y(_1495_),
    .A(_1489_),
    .B(_1492_));
 sg13g2_nand3_1 _5009_ (.B(_1485_),
    .C(_1495_),
    .A(_1491_),
    .Y(_1496_));
 sg13g2_nor2b_1 _5010_ (.A(_1494_),
    .B_N(_1496_),
    .Y(_0273_));
 sg13g2_o21ai_1 _5011_ (.B1(net172),
    .Y(_1497_),
    .A1(_1481_),
    .A2(_1489_));
 sg13g2_nand2_1 _5012_ (.Y(_1498_),
    .A(_1491_),
    .B(_1493_));
 sg13g2_a21oi_1 _5013_ (.A1(_1497_),
    .A2(_1498_),
    .Y(_0274_),
    .B1(_1168_));
 sg13g2_inv_1 _5014_ (.Y(_1499_),
    .A(_1161_));
 sg13g2_nand2_2 _5015_ (.Y(_1500_),
    .A(net173),
    .B(_1174_));
 sg13g2_inv_1 _5016_ (.Y(_1501_),
    .A(_1500_));
 sg13g2_nand2_1 _5017_ (.Y(_1502_),
    .A(_1499_),
    .B(_1501_));
 sg13g2_nand3_1 _5018_ (.B(_1481_),
    .C(_1500_),
    .A(_1161_),
    .Y(_1503_));
 sg13g2_a21oi_1 _5019_ (.A1(_1502_),
    .A2(_1503_),
    .Y(_0275_),
    .B1(_1168_));
 sg13g2_nor2_1 _5020_ (.A(_1499_),
    .B(net170),
    .Y(_1504_));
 sg13g2_nand2_1 _5021_ (.Y(_1505_),
    .A(_1481_),
    .B(_1500_));
 sg13g2_nand2_1 _5022_ (.Y(_1506_),
    .A(_1502_),
    .B(_1505_));
 sg13g2_a22oi_1 _5023_ (.Y(_1507_),
    .B1(_1506_),
    .B2(net170),
    .A2(_1504_),
    .A1(_1501_));
 sg13g2_nor2_1 _5024_ (.A(_1168_),
    .B(_1507_),
    .Y(_0276_));
 sg13g2_buf_1 _5025_ (.A(\Pong.datapath.scoreRight[2] ),
    .X(_1508_));
 sg13g2_and2_1 _5026_ (.A(_1161_),
    .B(net170),
    .X(_1509_));
 sg13g2_buf_1 _5027_ (.A(_1509_),
    .X(_1510_));
 sg13g2_o21ai_1 _5028_ (.B1(_1505_),
    .Y(_1511_),
    .A1(_1500_),
    .A2(_1510_));
 sg13g2_nand2_1 _5029_ (.Y(_1512_),
    .A(_1161_),
    .B(net170));
 sg13g2_nor2_1 _5030_ (.A(net167),
    .B(_1512_),
    .Y(_1513_));
 sg13g2_a22oi_1 _5031_ (.Y(_1514_),
    .B1(_1513_),
    .B2(_1501_),
    .A2(_1511_),
    .A1(net167));
 sg13g2_nor2_1 _5032_ (.A(_1168_),
    .B(_1514_),
    .Y(_0277_));
 sg13g2_buf_1 _5033_ (.A(_1160_),
    .X(_1515_));
 sg13g2_a21oi_1 _5034_ (.A1(net167),
    .A2(_1510_),
    .Y(_1516_),
    .B1(_1515_));
 sg13g2_or3_1 _5035_ (.A(_1166_),
    .B(_1500_),
    .C(_1516_),
    .X(_1517_));
 sg13g2_nand2_1 _5036_ (.Y(_1518_),
    .A(net173),
    .B(_1166_));
 sg13g2_nand3_1 _5037_ (.B(_1518_),
    .C(_1481_),
    .A(_1515_),
    .Y(_1519_));
 sg13g2_a21oi_1 _5038_ (.A1(_1517_),
    .A2(_1519_),
    .Y(_0278_),
    .B1(net138));
 sg13g2_nor3_1 _5039_ (.A(_1166_),
    .B(_1174_),
    .C(_1179_),
    .Y(_1520_));
 sg13g2_a22oi_1 _5040_ (.Y(_1521_),
    .B1(net131),
    .B2(_0509_),
    .A2(_1151_),
    .A1(_0507_));
 sg13g2_o21ai_1 _5041_ (.B1(_2737_),
    .Y(_1522_),
    .A1(net173),
    .A2(_1521_));
 sg13g2_a21o_1 _5042_ (.A2(_1520_),
    .A1(_1154_),
    .B1(_1522_),
    .X(_0279_));
 sg13g2_buf_1 _5043_ (.A(\Pong.datapath.vga.Column_Counter.Q[4] ),
    .X(_1523_));
 sg13g2_buf_1 _5044_ (.A(_1523_),
    .X(_1524_));
 sg13g2_inv_1 _5045_ (.Y(_1525_),
    .A(\Pong.datapath.vga.Column_Counter.Q[5] ));
 sg13g2_nand2_2 _5046_ (.Y(_1526_),
    .A(net127),
    .B(_1525_));
 sg13g2_buf_2 _5047_ (.A(\Pong.datapath.vga.Column_Counter.Q[1] ),
    .X(_1527_));
 sg13g2_buf_1 _5048_ (.A(\Pong.datapath.vga.Column_Counter.Q[0] ),
    .X(_1528_));
 sg13g2_buf_1 _5049_ (.A(_1528_),
    .X(_1529_));
 sg13g2_nand2_1 _5050_ (.Y(_1530_),
    .A(_1527_),
    .B(net126));
 sg13g2_buf_2 _5051_ (.A(\Pong.datapath.vga.Column_Counter.Q[3] ),
    .X(_1531_));
 sg13g2_buf_1 _5052_ (.A(\Pong.datapath.vga.Column_Counter.Q[2] ),
    .X(_1532_));
 sg13g2_buf_1 _5053_ (.A(_1532_),
    .X(_1533_));
 sg13g2_nand2_1 _5054_ (.Y(_1534_),
    .A(_1531_),
    .B(_1533_));
 sg13g2_or2_1 _5055_ (.X(_1535_),
    .B(_1534_),
    .A(_1530_));
 sg13g2_buf_1 _5056_ (.A(_1535_),
    .X(_1536_));
 sg13g2_buf_1 _5057_ (.A(\Pong.datapath.vga.Column_Counter.Q[8] ),
    .X(_1537_));
 sg13g2_buf_1 _5058_ (.A(_1537_),
    .X(_1538_));
 sg13g2_buf_1 _5059_ (.A(\Pong.datapath.vga.Column_Counter.Q[9] ),
    .X(_1539_));
 sg13g2_nand2_1 _5060_ (.Y(_1540_),
    .A(net124),
    .B(net166));
 sg13g2_buf_2 _5061_ (.A(\Pong.datapath.vga.Column_Counter.Q[7] ),
    .X(_1541_));
 sg13g2_buf_2 _5062_ (.A(\Pong.datapath.vga.Column_Counter.Q[6] ),
    .X(_1542_));
 sg13g2_or2_1 _5063_ (.X(_1543_),
    .B(_1542_),
    .A(net165));
 sg13g2_buf_2 _5064_ (.A(_1543_),
    .X(_1544_));
 sg13g2_or4_1 _5065_ (.A(_1526_),
    .B(_1536_),
    .C(_1540_),
    .D(_1544_),
    .X(_1545_));
 sg13g2_nand2_1 _5066_ (.Y(_1546_),
    .A(_2656_),
    .B(_1545_));
 sg13g2_buf_1 _5067_ (.A(_1546_),
    .X(_1547_));
 sg13g2_buf_2 _5068_ (.A(_0114_),
    .X(_1548_));
 sg13g2_nor2_1 _5069_ (.A(net165),
    .B(_1542_),
    .Y(_1549_));
 sg13g2_a21oi_2 _5070_ (.B1(_1540_),
    .Y(_1550_),
    .A2(_1549_),
    .A1(_1548_));
 sg13g2_inv_1 _5071_ (.Y(_1551_),
    .A(_1550_));
 sg13g2_nor2_1 _5072_ (.A(net126),
    .B(_1551_),
    .Y(_1552_));
 sg13g2_nor2b_1 _5073_ (.A(_1550_),
    .B_N(net126),
    .Y(_1553_));
 sg13g2_nor3_1 _5074_ (.A(net65),
    .B(_1552_),
    .C(_1553_),
    .Y(_0280_));
 sg13g2_xnor2_1 _5075_ (.Y(_1554_),
    .A(_1527_),
    .B(_1553_));
 sg13g2_nor2_1 _5076_ (.A(net65),
    .B(_1554_),
    .Y(_0281_));
 sg13g2_buf_1 _5077_ (.A(_1550_),
    .X(_1555_));
 sg13g2_buf_1 _5078_ (.A(_0101_),
    .X(_1556_));
 sg13g2_xnor2_1 _5079_ (.Y(_1557_),
    .A(_1556_),
    .B(_1530_));
 sg13g2_nor2_1 _5080_ (.A(net86),
    .B(_1557_),
    .Y(_1558_));
 sg13g2_a21oi_1 _5081_ (.A1(net125),
    .A2(net86),
    .Y(_1559_),
    .B1(_1558_));
 sg13g2_nor2_1 _5082_ (.A(net65),
    .B(_1559_),
    .Y(_0282_));
 sg13g2_buf_1 _5083_ (.A(_1531_),
    .X(_1560_));
 sg13g2_buf_1 _5084_ (.A(_0102_),
    .X(_1561_));
 sg13g2_nand3_1 _5085_ (.B(_1527_),
    .C(net126),
    .A(_1533_),
    .Y(_1562_));
 sg13g2_xnor2_1 _5086_ (.Y(_1563_),
    .A(net163),
    .B(_1562_));
 sg13g2_nor2_1 _5087_ (.A(net86),
    .B(_1563_),
    .Y(_1564_));
 sg13g2_a21oi_1 _5088_ (.A1(net123),
    .A2(_1555_),
    .Y(_1565_),
    .B1(_1564_));
 sg13g2_nor2_1 _5089_ (.A(net65),
    .B(_1565_),
    .Y(_0283_));
 sg13g2_buf_2 _5090_ (.A(_0103_),
    .X(_1566_));
 sg13g2_xnor2_1 _5091_ (.Y(_1567_),
    .A(_1566_),
    .B(_1536_));
 sg13g2_nor2_1 _5092_ (.A(net86),
    .B(_1567_),
    .Y(_1568_));
 sg13g2_a21oi_1 _5093_ (.A1(_1524_),
    .A2(_1555_),
    .Y(_1569_),
    .B1(_1568_));
 sg13g2_nor2_1 _5094_ (.A(_1547_),
    .B(_1569_),
    .Y(_0284_));
 sg13g2_buf_1 _5095_ (.A(\Pong.datapath.vga.Column_Counter.Q[5] ),
    .X(_1570_));
 sg13g2_nor2_1 _5096_ (.A(_1530_),
    .B(_1534_),
    .Y(_1571_));
 sg13g2_nand2_1 _5097_ (.Y(_1572_),
    .A(net127),
    .B(_1571_));
 sg13g2_xnor2_1 _5098_ (.Y(_1573_),
    .A(_1548_),
    .B(_1572_));
 sg13g2_nor2_1 _5099_ (.A(net86),
    .B(_1573_),
    .Y(_1574_));
 sg13g2_a21oi_1 _5100_ (.A1(net162),
    .A2(net86),
    .Y(_1575_),
    .B1(_1574_));
 sg13g2_nor2_1 _5101_ (.A(_1547_),
    .B(_1575_),
    .Y(_0285_));
 sg13g2_buf_2 _5102_ (.A(_0104_),
    .X(_1576_));
 sg13g2_nor2_1 _5103_ (.A(_1525_),
    .B(_1572_),
    .Y(_1577_));
 sg13g2_xor2_1 _5104_ (.B(_1577_),
    .A(_1576_),
    .X(_1578_));
 sg13g2_nor2_1 _5105_ (.A(_1550_),
    .B(_1578_),
    .Y(_1579_));
 sg13g2_a21oi_1 _5106_ (.A1(_1542_),
    .A2(net86),
    .Y(_1580_),
    .B1(_1579_));
 sg13g2_nor2_1 _5107_ (.A(net65),
    .B(_1580_),
    .Y(_0286_));
 sg13g2_buf_1 _5108_ (.A(_0105_),
    .X(_1581_));
 sg13g2_inv_1 _5109_ (.Y(_1582_),
    .A(_1542_));
 sg13g2_nor3_2 _5110_ (.A(_1582_),
    .B(_1525_),
    .C(_1572_),
    .Y(_1583_));
 sg13g2_xor2_1 _5111_ (.B(_1583_),
    .A(_1581_),
    .X(_1584_));
 sg13g2_nor2_1 _5112_ (.A(_1550_),
    .B(_1584_),
    .Y(_1585_));
 sg13g2_a21oi_1 _5113_ (.A1(net165),
    .A2(net86),
    .Y(_1586_),
    .B1(_1585_));
 sg13g2_nor2_1 _5114_ (.A(net65),
    .B(_1586_),
    .Y(_0287_));
 sg13g2_nand2_1 _5115_ (.Y(_1587_),
    .A(net165),
    .B(_1583_));
 sg13g2_xnor2_1 _5116_ (.Y(_1588_),
    .A(_0106_),
    .B(_1587_));
 sg13g2_a21oi_1 _5117_ (.A1(_1551_),
    .A2(_1588_),
    .Y(_0288_),
    .B1(net65));
 sg13g2_buf_2 _5118_ (.A(_0107_),
    .X(_1589_));
 sg13g2_nand3_1 _5119_ (.B(net124),
    .C(_1583_),
    .A(net165),
    .Y(_1590_));
 sg13g2_xnor2_1 _5120_ (.Y(_1591_),
    .A(_1589_),
    .B(_1590_));
 sg13g2_a21oi_1 _5121_ (.A1(_1551_),
    .A2(_1591_),
    .Y(_0289_),
    .B1(net65));
 sg13g2_buf_2 _5122_ (.A(\Pong.datapath.vga.Row_Counter.Q[0] ),
    .X(_1592_));
 sg13g2_buf_1 _5123_ (.A(_1592_),
    .X(_1593_));
 sg13g2_nor4_1 _5124_ (.A(_1526_),
    .B(_1536_),
    .C(_1540_),
    .D(_1544_),
    .Y(_1594_));
 sg13g2_buf_1 _5125_ (.A(\Pong.datapath.vga.Row_Counter.Q[1] ),
    .X(_1595_));
 sg13g2_buf_1 _5126_ (.A(_1595_),
    .X(_1596_));
 sg13g2_nor2_1 _5127_ (.A(net121),
    .B(net122),
    .Y(_1597_));
 sg13g2_buf_1 _5128_ (.A(\Pong.datapath.vga.Row_Counter.Q[3] ),
    .X(_1598_));
 sg13g2_buf_2 _5129_ (.A(\Pong.datapath.vga.Row_Counter.Q[2] ),
    .X(_1599_));
 sg13g2_nand2_1 _5130_ (.Y(_1600_),
    .A(_1598_),
    .B(_1599_));
 sg13g2_buf_1 _5131_ (.A(\Pong.datapath.vga.Row_Counter.Q[5] ),
    .X(_1601_));
 sg13g2_buf_1 _5132_ (.A(\Pong.datapath.vga.Row_Counter.Q[4] ),
    .X(_1602_));
 sg13g2_nor2_1 _5133_ (.A(_1601_),
    .B(_1602_),
    .Y(_1603_));
 sg13g2_o21ai_1 _5134_ (.B1(_1603_),
    .Y(_1604_),
    .A1(_1597_),
    .A2(_1600_));
 sg13g2_buf_2 _5135_ (.A(\Pong.datapath.vga.Row_Counter.Q[8] ),
    .X(_1605_));
 sg13g2_buf_1 _5136_ (.A(\Pong.datapath.vga.Row_Counter.Q[7] ),
    .X(_1606_));
 sg13g2_buf_1 _5137_ (.A(\Pong.datapath.vga.Row_Counter.Q[6] ),
    .X(_1607_));
 sg13g2_nor3_1 _5138_ (.A(_1605_),
    .B(net161),
    .C(net160),
    .Y(_1608_));
 sg13g2_inv_1 _5139_ (.Y(_1609_),
    .A(_1608_));
 sg13g2_buf_1 _5140_ (.A(\Pong.datapath.vga.Row_Counter.Q[9] ),
    .X(_1610_));
 sg13g2_buf_1 _5141_ (.A(_1610_),
    .X(_1611_));
 sg13g2_o21ai_1 _5142_ (.B1(net120),
    .Y(_1612_),
    .A1(_1604_),
    .A2(_1609_));
 sg13g2_nand2_1 _5143_ (.Y(_1613_),
    .A(_1594_),
    .B(_1612_));
 sg13g2_buf_1 _5144_ (.A(_1613_),
    .X(_1614_));
 sg13g2_nand2_1 _5145_ (.Y(_1615_),
    .A(net122),
    .B(net64));
 sg13g2_inv_1 _5146_ (.Y(_1616_),
    .A(_1592_));
 sg13g2_nand3_1 _5147_ (.B(_1600_),
    .C(_1608_),
    .A(_1603_),
    .Y(_1617_));
 sg13g2_a21oi_1 _5148_ (.A1(net120),
    .A2(_1617_),
    .Y(_1618_),
    .B1(_1545_));
 sg13g2_buf_1 _5149_ (.A(_1618_),
    .X(_1619_));
 sg13g2_nand2_1 _5150_ (.Y(_1620_),
    .A(_1616_),
    .B(net63));
 sg13g2_a21oi_1 _5151_ (.A1(_1615_),
    .A2(_1620_),
    .Y(_0290_),
    .B1(net138));
 sg13g2_xor2_1 _5152_ (.B(net122),
    .A(net121),
    .X(_1621_));
 sg13g2_a22oi_1 _5153_ (.Y(_1622_),
    .B1(net63),
    .B2(_1621_),
    .A2(_1614_),
    .A1(net121));
 sg13g2_nor2_1 _5154_ (.A(net158),
    .B(_1622_),
    .Y(_0291_));
 sg13g2_buf_1 _5155_ (.A(_1599_),
    .X(_1623_));
 sg13g2_nand2_1 _5156_ (.Y(_1624_),
    .A(net119),
    .B(net64));
 sg13g2_buf_2 _5157_ (.A(_0093_),
    .X(_1625_));
 sg13g2_buf_1 _5158_ (.A(_1625_),
    .X(_1626_));
 sg13g2_nand2_1 _5159_ (.Y(_1627_),
    .A(net121),
    .B(net122));
 sg13g2_xor2_1 _5160_ (.B(_1627_),
    .A(net118),
    .X(_1628_));
 sg13g2_nand2_1 _5161_ (.Y(_1629_),
    .A(_1619_),
    .B(_1628_));
 sg13g2_a21oi_1 _5162_ (.A1(_1624_),
    .A2(_1629_),
    .Y(_0292_),
    .B1(net138));
 sg13g2_buf_1 _5163_ (.A(_1598_),
    .X(_1630_));
 sg13g2_nand2_1 _5164_ (.Y(_1631_),
    .A(net117),
    .B(net64));
 sg13g2_buf_1 _5165_ (.A(_0094_),
    .X(_1632_));
 sg13g2_inv_2 _5166_ (.Y(_1633_),
    .A(net159));
 sg13g2_nand3_1 _5167_ (.B(_1596_),
    .C(net122),
    .A(net119),
    .Y(_1634_));
 sg13g2_xnor2_1 _5168_ (.Y(_1635_),
    .A(_1633_),
    .B(_1634_));
 sg13g2_nand2_1 _5169_ (.Y(_1636_),
    .A(net63),
    .B(_1635_));
 sg13g2_a21oi_1 _5170_ (.A1(_1631_),
    .A2(_1636_),
    .Y(_0293_),
    .B1(net138));
 sg13g2_buf_1 _5171_ (.A(_1602_),
    .X(_1637_));
 sg13g2_nand2_1 _5172_ (.Y(_1638_),
    .A(net116),
    .B(_1614_));
 sg13g2_buf_1 _5173_ (.A(_0095_),
    .X(_1639_));
 sg13g2_buf_1 _5174_ (.A(_1639_),
    .X(_1640_));
 sg13g2_nor2_1 _5175_ (.A(_1600_),
    .B(_1627_),
    .Y(_1641_));
 sg13g2_xnor2_1 _5176_ (.Y(_1642_),
    .A(net115),
    .B(_1641_));
 sg13g2_nand2_1 _5177_ (.Y(_1643_),
    .A(_1619_),
    .B(_1642_));
 sg13g2_a21oi_1 _5178_ (.A1(_1638_),
    .A2(_1643_),
    .Y(_0294_),
    .B1(net138));
 sg13g2_buf_1 _5179_ (.A(_1601_),
    .X(_1644_));
 sg13g2_buf_2 _5180_ (.A(_0096_),
    .X(_1645_));
 sg13g2_buf_1 _5181_ (.A(_1645_),
    .X(_1646_));
 sg13g2_inv_1 _5182_ (.Y(_1647_),
    .A(net116));
 sg13g2_nor3_1 _5183_ (.A(_1647_),
    .B(_1600_),
    .C(_1627_),
    .Y(_1648_));
 sg13g2_xnor2_1 _5184_ (.Y(_1649_),
    .A(net113),
    .B(_1648_));
 sg13g2_a22oi_1 _5185_ (.Y(_1650_),
    .B1(net63),
    .B2(_1649_),
    .A2(net64),
    .A1(net114));
 sg13g2_nor2_1 _5186_ (.A(net158),
    .B(_1650_),
    .Y(_0295_));
 sg13g2_buf_2 _5187_ (.A(_0097_),
    .X(_1651_));
 sg13g2_nand2_1 _5188_ (.Y(_1652_),
    .A(net114),
    .B(_1648_));
 sg13g2_xor2_1 _5189_ (.B(_1652_),
    .A(_1651_),
    .X(_1653_));
 sg13g2_a22oi_1 _5190_ (.Y(_1654_),
    .B1(net63),
    .B2(_1653_),
    .A2(net64),
    .A1(net160));
 sg13g2_nor2_1 _5191_ (.A(net158),
    .B(_1654_),
    .Y(_0296_));
 sg13g2_buf_1 _5192_ (.A(_0098_),
    .X(_1655_));
 sg13g2_inv_1 _5193_ (.Y(_1656_),
    .A(net160));
 sg13g2_nor2_1 _5194_ (.A(_1656_),
    .B(_1652_),
    .Y(_1657_));
 sg13g2_xnor2_1 _5195_ (.Y(_1658_),
    .A(_1655_),
    .B(_1657_));
 sg13g2_a22oi_1 _5196_ (.Y(_1659_),
    .B1(net63),
    .B2(_1658_),
    .A2(net64),
    .A1(net161));
 sg13g2_nor2_1 _5197_ (.A(net158),
    .B(_1659_),
    .Y(_0297_));
 sg13g2_nand2_1 _5198_ (.Y(_1660_),
    .A(_1605_),
    .B(net64));
 sg13g2_buf_2 _5199_ (.A(_0099_),
    .X(_1661_));
 sg13g2_inv_1 _5200_ (.Y(_1662_),
    .A(_1661_));
 sg13g2_nand2_1 _5201_ (.Y(_1663_),
    .A(net161),
    .B(_1657_));
 sg13g2_xnor2_1 _5202_ (.Y(_1664_),
    .A(_1662_),
    .B(_1663_));
 sg13g2_nand2_1 _5203_ (.Y(_1665_),
    .A(net63),
    .B(_1664_));
 sg13g2_a21oi_1 _5204_ (.A1(_1660_),
    .A2(_1665_),
    .Y(_0298_),
    .B1(net138));
 sg13g2_buf_1 _5205_ (.A(_0100_),
    .X(_1666_));
 sg13g2_buf_1 _5206_ (.A(_1666_),
    .X(_1667_));
 sg13g2_nand2_1 _5207_ (.Y(_1668_),
    .A(_1605_),
    .B(net161));
 sg13g2_nor3_1 _5208_ (.A(_1656_),
    .B(_1652_),
    .C(_1668_),
    .Y(_1669_));
 sg13g2_xnor2_1 _5209_ (.Y(_1670_),
    .A(_1667_),
    .B(_1669_));
 sg13g2_a22oi_1 _5210_ (.Y(_1671_),
    .B1(net63),
    .B2(_1670_),
    .A2(net64),
    .A1(net120));
 sg13g2_nor2_1 _5211_ (.A(net158),
    .B(_1671_),
    .Y(_0299_));
 sg13g2_nand3_1 _5212_ (.B(net161),
    .C(\Pong.datapath.vga.Row_Counter.Q[6] ),
    .A(_1605_),
    .Y(_1672_));
 sg13g2_inv_1 _5213_ (.Y(_1673_),
    .A(_1672_));
 sg13g2_nand2b_1 _5214_ (.Y(_1674_),
    .B(_1581_),
    .A_N(net124));
 sg13g2_nand2b_1 _5215_ (.Y(_1675_),
    .B(net166),
    .A_N(_1537_));
 sg13g2_nand3b_1 _5216_ (.B(_1542_),
    .C(\Pong.datapath.vga.Column_Counter.Q[5] ),
    .Y(_1676_),
    .A_N(net165));
 sg13g2_buf_1 _5217_ (.A(_1676_),
    .X(_1677_));
 sg13g2_a21oi_1 _5218_ (.A1(_1531_),
    .A2(net125),
    .Y(_1678_),
    .B1(_1523_));
 sg13g2_nor3_1 _5219_ (.A(_1675_),
    .B(_1677_),
    .C(_1678_),
    .Y(_1679_));
 sg13g2_a21oi_1 _5220_ (.A1(net166),
    .A2(_1674_),
    .Y(_1680_),
    .B1(_1679_));
 sg13g2_or2_1 _5221_ (.X(_1681_),
    .B(_1677_),
    .A(_1675_));
 sg13g2_or2_1 _5222_ (.X(_1682_),
    .B(_1528_),
    .A(_1527_));
 sg13g2_buf_1 _5223_ (.A(_1682_),
    .X(_1683_));
 sg13g2_nor4_1 _5224_ (.A(net127),
    .B(_1534_),
    .C(_1681_),
    .D(_1683_),
    .Y(_1684_));
 sg13g2_inv_1 _5225_ (.Y(_1685_),
    .A(_1523_));
 sg13g2_nor2_1 _5226_ (.A(_1531_),
    .B(net125),
    .Y(_1686_));
 sg13g2_nor4_1 _5227_ (.A(net162),
    .B(net124),
    .C(net166),
    .D(_1544_),
    .Y(_1687_));
 sg13g2_o21ai_1 _5228_ (.B1(_1687_),
    .Y(_1688_),
    .A1(_1685_),
    .A2(_1686_));
 sg13g2_o21ai_1 _5229_ (.B1(_1688_),
    .Y(_1689_),
    .A1(_1680_),
    .A2(_1684_));
 sg13g2_inv_1 _5230_ (.Y(_1690_),
    .A(net114));
 sg13g2_or2_1 _5231_ (.X(_1691_),
    .B(_1599_),
    .A(_1598_));
 sg13g2_buf_1 _5232_ (.A(_1691_),
    .X(_1692_));
 sg13g2_nand2_1 _5233_ (.Y(_1693_),
    .A(net116),
    .B(_1692_));
 sg13g2_nand3_1 _5234_ (.B(_1608_),
    .C(_1693_),
    .A(_1690_),
    .Y(_1694_));
 sg13g2_nand2_1 _5235_ (.Y(_1695_),
    .A(_1604_),
    .B(_1673_));
 sg13g2_nand2_1 _5236_ (.Y(_1696_),
    .A(_1694_),
    .B(_1695_));
 sg13g2_o21ai_1 _5237_ (.B1(net166),
    .Y(_1697_),
    .A1(net165),
    .A2(net124));
 sg13g2_nand2b_1 _5238_ (.Y(_1698_),
    .B(_1697_),
    .A_N(net120));
 sg13g2_a221oi_1 _5239_ (.B2(_1696_),
    .C1(_1698_),
    .B1(_1689_),
    .A1(net114),
    .Y(_1699_),
    .A2(_1673_));
 sg13g2_xor2_1 _5240_ (.B(_1645_),
    .A(net70),
    .X(_1700_));
 sg13g2_xnor2_1 _5241_ (.Y(_1701_),
    .A(_2920_),
    .B(_1666_));
 sg13g2_buf_2 _5242_ (.A(_1701_),
    .X(_1702_));
 sg13g2_xnor2_1 _5243_ (.Y(_1703_),
    .A(_1144_),
    .B(_1702_));
 sg13g2_nand2_1 _5244_ (.Y(_1704_),
    .A(_1700_),
    .B(_1703_));
 sg13g2_xnor2_1 _5245_ (.Y(_1705_),
    .A(net70),
    .B(_1645_));
 sg13g2_buf_2 _5246_ (.A(_1705_),
    .X(_1706_));
 sg13g2_nand2_1 _5247_ (.Y(_1707_),
    .A(_1702_),
    .B(_1706_));
 sg13g2_inv_1 _5248_ (.Y(_1708_),
    .A(_1707_));
 sg13g2_nand2_1 _5249_ (.Y(_1709_),
    .A(_1104_),
    .B(_1708_));
 sg13g2_o21ai_1 _5250_ (.B1(_1709_),
    .Y(_1710_),
    .A1(_1104_),
    .A2(_1704_));
 sg13g2_and2_1 _5251_ (.A(_2761_),
    .B(net74),
    .X(_1711_));
 sg13g2_buf_1 _5252_ (.A(_1711_),
    .X(_1712_));
 sg13g2_xor2_1 _5253_ (.B(_1651_),
    .A(_3033_),
    .X(_1713_));
 sg13g2_buf_2 _5254_ (.A(_1713_),
    .X(_1714_));
 sg13g2_xor2_1 _5255_ (.B(net118),
    .A(net69),
    .X(_1715_));
 sg13g2_xor2_1 _5256_ (.B(_1639_),
    .A(_2942_),
    .X(_1716_));
 sg13g2_buf_1 _5257_ (.A(_1716_),
    .X(_1717_));
 sg13g2_nor4_1 _5258_ (.A(_1712_),
    .B(_1714_),
    .C(_1715_),
    .D(net25),
    .Y(_1718_));
 sg13g2_xnor2_1 _5259_ (.Y(_1719_),
    .A(net69),
    .B(net118));
 sg13g2_xor2_1 _5260_ (.B(_1661_),
    .A(_2896_),
    .X(_1720_));
 sg13g2_buf_1 _5261_ (.A(_1720_),
    .X(_1721_));
 sg13g2_nand2_1 _5262_ (.Y(_1722_),
    .A(net54),
    .B(net72));
 sg13g2_a21oi_1 _5263_ (.A1(net24),
    .A2(_1722_),
    .Y(_1723_),
    .B1(_1133_));
 sg13g2_nor2_1 _5264_ (.A(_1111_),
    .B(_1714_),
    .Y(_1724_));
 sg13g2_nor4_1 _5265_ (.A(net15),
    .B(_1719_),
    .C(_1723_),
    .D(_1724_),
    .Y(_1725_));
 sg13g2_nor2_1 _5266_ (.A(_1718_),
    .B(_1725_),
    .Y(_1726_));
 sg13g2_xnor2_1 _5267_ (.Y(_1727_),
    .A(_2942_),
    .B(_1639_));
 sg13g2_nand2_1 _5268_ (.Y(_1728_),
    .A(_1097_),
    .B(_1727_));
 sg13g2_a22oi_1 _5269_ (.Y(_1729_),
    .B1(net25),
    .B2(_1096_),
    .A2(_1714_),
    .A1(_1111_));
 sg13g2_xnor2_1 _5270_ (.Y(_1730_),
    .A(_2755_),
    .B(net159));
 sg13g2_buf_2 _5271_ (.A(_1730_),
    .X(_1731_));
 sg13g2_xor2_1 _5272_ (.B(_1655_),
    .A(net71),
    .X(_1732_));
 sg13g2_buf_1 _5273_ (.A(_1732_),
    .X(_1733_));
 sg13g2_xnor2_1 _5274_ (.Y(_1734_),
    .A(_1126_),
    .B(net23));
 sg13g2_o21ai_1 _5275_ (.B1(_1083_),
    .Y(_1735_),
    .A1(_1731_),
    .A2(_1734_));
 sg13g2_xor2_1 _5276_ (.B(_0094_),
    .A(_2755_),
    .X(_1736_));
 sg13g2_buf_2 _5277_ (.A(_1736_),
    .X(_1737_));
 sg13g2_o21ai_1 _5278_ (.B1(_1087_),
    .Y(_1738_),
    .A1(net23),
    .A2(_1737_));
 sg13g2_nand4_1 _5279_ (.B(_1729_),
    .C(_1735_),
    .A(_1728_),
    .Y(_1739_),
    .D(_1738_));
 sg13g2_buf_1 _5280_ (.A(_0108_),
    .X(_1740_));
 sg13g2_buf_1 _5281_ (.A(_1740_),
    .X(_1741_));
 sg13g2_nor2b_2 _5282_ (.A(net122),
    .B_N(net111),
    .Y(_1742_));
 sg13g2_nor2b_1 _5283_ (.A(_1592_),
    .B_N(_2760_),
    .Y(_1743_));
 sg13g2_nor2b_2 _5284_ (.A(_2760_),
    .B_N(_1592_),
    .Y(_1744_));
 sg13g2_xor2_1 _5285_ (.B(_1740_),
    .A(net74),
    .X(_1745_));
 sg13g2_mux2_1 _5286_ (.A0(_1743_),
    .A1(_1744_),
    .S(_1745_),
    .X(_1746_));
 sg13g2_xnor2_1 _5287_ (.Y(_1747_),
    .A(_2896_),
    .B(_1661_));
 sg13g2_a22oi_1 _5288_ (.Y(_1748_),
    .B1(_1746_),
    .B2(_1747_),
    .A2(_1742_),
    .A1(_1134_));
 sg13g2_nor3_1 _5289_ (.A(_1726_),
    .B(_1739_),
    .C(_1748_),
    .Y(_1749_));
 sg13g2_xnor2_1 _5290_ (.Y(_1750_),
    .A(net71),
    .B(_1655_));
 sg13g2_nor2_1 _5291_ (.A(net24),
    .B(_1714_),
    .Y(_1751_));
 sg13g2_and2_1 _5292_ (.A(_1123_),
    .B(_1751_),
    .X(_1752_));
 sg13g2_xnor2_1 _5293_ (.Y(_1753_),
    .A(_3033_),
    .B(_1651_));
 sg13g2_nor2_1 _5294_ (.A(net23),
    .B(net24),
    .Y(_1754_));
 sg13g2_xnor2_1 _5295_ (.Y(_1755_),
    .A(net55),
    .B(_1747_));
 sg13g2_nor2_1 _5296_ (.A(net53),
    .B(_1750_),
    .Y(_1756_));
 sg13g2_a22oi_1 _5297_ (.Y(_1757_),
    .B1(_1755_),
    .B2(_1756_),
    .A2(_1754_),
    .A1(net34));
 sg13g2_nor2_1 _5298_ (.A(_1753_),
    .B(_1757_),
    .Y(_1758_));
 sg13g2_a22oi_1 _5299_ (.Y(_1759_),
    .B1(_1758_),
    .B2(_1115_),
    .A2(_1752_),
    .A1(_1750_));
 sg13g2_nand3_1 _5300_ (.B(_1731_),
    .C(_1719_),
    .A(_2889_),
    .Y(_1760_));
 sg13g2_nand2_1 _5301_ (.Y(_1761_),
    .A(_2775_),
    .B(_1122_));
 sg13g2_xnor2_1 _5302_ (.Y(_1762_),
    .A(net57),
    .B(_1731_));
 sg13g2_nand4_1 _5303_ (.B(_1715_),
    .C(_1761_),
    .A(_1073_),
    .Y(_1763_),
    .D(_1762_));
 sg13g2_nand2_1 _5304_ (.Y(_1764_),
    .A(_1760_),
    .B(_1763_));
 sg13g2_mux2_1 _5305_ (.A0(_1744_),
    .A1(_1743_),
    .S(_1745_),
    .X(_1765_));
 sg13g2_xor2_1 _5306_ (.B(_1702_),
    .A(_1142_),
    .X(_1766_));
 sg13g2_nand2_1 _5307_ (.Y(_1767_),
    .A(_1706_),
    .B(_1727_));
 sg13g2_xnor2_1 _5308_ (.Y(_1768_),
    .A(_2753_),
    .B(_1706_));
 sg13g2_nand3_1 _5309_ (.B(net25),
    .C(_1768_),
    .A(_1093_),
    .Y(_1769_));
 sg13g2_o21ai_1 _5310_ (.B1(_1769_),
    .Y(_1770_),
    .A1(_1093_),
    .A2(_1767_));
 sg13g2_nand4_1 _5311_ (.B(_1765_),
    .C(_1766_),
    .A(_1764_),
    .Y(_1771_),
    .D(_1770_));
 sg13g2_xnor2_1 _5312_ (.Y(_1772_),
    .A(net37),
    .B(_1623_));
 sg13g2_xnor2_1 _5313_ (.Y(_1773_),
    .A(net72),
    .B(net120));
 sg13g2_or2_1 _5314_ (.X(_1774_),
    .B(_1744_),
    .A(_1743_));
 sg13g2_buf_1 _5315_ (.A(_1774_),
    .X(_1775_));
 sg13g2_xor2_1 _5316_ (.B(_1595_),
    .A(net74),
    .X(_1776_));
 sg13g2_xor2_1 _5317_ (.B(net114),
    .A(net61),
    .X(_1777_));
 sg13g2_xor2_1 _5318_ (.B(_1605_),
    .A(net54),
    .X(_1778_));
 sg13g2_nor4_1 _5319_ (.A(_1775_),
    .B(_1776_),
    .C(_1777_),
    .D(_1778_),
    .Y(_1779_));
 sg13g2_xor2_1 _5320_ (.B(_1637_),
    .A(net38),
    .X(_1780_));
 sg13g2_xor2_1 _5321_ (.B(net161),
    .A(net55),
    .X(_1781_));
 sg13g2_xor2_1 _5322_ (.B(net160),
    .A(_2893_),
    .X(_1782_));
 sg13g2_xor2_1 _5323_ (.B(net117),
    .A(net36),
    .X(_1783_));
 sg13g2_nor4_1 _5324_ (.A(_1780_),
    .B(_1781_),
    .C(_1782_),
    .D(_1783_),
    .Y(_1784_));
 sg13g2_nand4_1 _5325_ (.B(_1773_),
    .C(_1779_),
    .A(_1772_),
    .Y(_1785_),
    .D(_1784_));
 sg13g2_o21ai_1 _5326_ (.B1(_1785_),
    .Y(_1786_),
    .A1(_1759_),
    .A2(_1771_));
 sg13g2_a21oi_1 _5327_ (.A1(_1710_),
    .A2(_1749_),
    .Y(_1787_),
    .B1(_1786_));
 sg13g2_inv_1 _5328_ (.Y(_1788_),
    .A(net69));
 sg13g2_xnor2_1 _5329_ (.Y(_1789_),
    .A(_1788_),
    .B(_1731_));
 sg13g2_nand3_1 _5330_ (.B(_1091_),
    .C(net25),
    .A(net15),
    .Y(_1790_));
 sg13g2_o21ai_1 _5331_ (.B1(_1790_),
    .Y(_1791_),
    .A1(_3026_),
    .A2(net25));
 sg13g2_nand3_1 _5332_ (.B(net15),
    .C(_1737_),
    .A(_2951_),
    .Y(_1792_));
 sg13g2_o21ai_1 _5333_ (.B1(_1792_),
    .Y(_1793_),
    .A1(_2951_),
    .A2(_1737_));
 sg13g2_nor3_1 _5334_ (.A(net37),
    .B(net15),
    .C(_1737_),
    .Y(_1794_));
 sg13g2_a21o_1 _5335_ (.A2(_1793_),
    .A1(_2892_),
    .B1(_1794_),
    .X(_1795_));
 sg13g2_a22oi_1 _5336_ (.Y(_1796_),
    .B1(_1795_),
    .B2(_1727_),
    .A2(_1791_),
    .A1(_1789_));
 sg13g2_nand2_1 _5337_ (.Y(_1797_),
    .A(_1077_),
    .B(_1122_));
 sg13g2_xnor2_1 _5338_ (.Y(_1798_),
    .A(_1136_),
    .B(_1721_));
 sg13g2_nor2_1 _5339_ (.A(_2775_),
    .B(_1753_),
    .Y(_1799_));
 sg13g2_nor2b_1 _5340_ (.A(_1797_),
    .B_N(_1799_),
    .Y(_1800_));
 sg13g2_a22oi_1 _5341_ (.Y(_1801_),
    .B1(_1798_),
    .B2(_1800_),
    .A2(_1797_),
    .A1(_1751_));
 sg13g2_or4_1 _5342_ (.A(_2766_),
    .B(_2893_),
    .C(net61),
    .D(net60),
    .X(_1802_));
 sg13g2_nor2_1 _5343_ (.A(_1788_),
    .B(_1802_),
    .Y(_1803_));
 sg13g2_xnor2_1 _5344_ (.Y(_1804_),
    .A(net23),
    .B(_1803_));
 sg13g2_xnor2_1 _5345_ (.Y(_1805_),
    .A(net118),
    .B(_1712_));
 sg13g2_or3_1 _5346_ (.A(net57),
    .B(net118),
    .C(_1712_),
    .X(_1806_));
 sg13g2_o21ai_1 _5347_ (.B1(_1806_),
    .Y(_1807_),
    .A1(_3026_),
    .A2(_1805_));
 sg13g2_nor3_1 _5348_ (.A(net37),
    .B(_1077_),
    .C(net23),
    .Y(_1808_));
 sg13g2_a22oi_1 _5349_ (.Y(_1809_),
    .B1(_1808_),
    .B2(net118),
    .A2(_1807_),
    .A1(_1804_));
 sg13g2_nor2_2 _5350_ (.A(net122),
    .B(net111),
    .Y(_1810_));
 sg13g2_a22oi_1 _5351_ (.Y(_1811_),
    .B1(_1810_),
    .B2(_2762_),
    .A2(_1745_),
    .A1(_1744_));
 sg13g2_xnor2_1 _5352_ (.Y(_1812_),
    .A(_1105_),
    .B(_1706_));
 sg13g2_nand3_1 _5353_ (.B(_1706_),
    .C(_1742_),
    .A(_1712_),
    .Y(_1813_));
 sg13g2_o21ai_1 _5354_ (.B1(_1813_),
    .Y(_1814_),
    .A1(_1811_),
    .A2(_1812_));
 sg13g2_nand3_1 _5355_ (.B(_1076_),
    .C(_1122_),
    .A(_1141_),
    .Y(_1815_));
 sg13g2_xnor2_1 _5356_ (.Y(_1816_),
    .A(_1702_),
    .B(_1815_));
 sg13g2_nand2_1 _5357_ (.Y(_1817_),
    .A(_1814_),
    .B(_1816_));
 sg13g2_or3_1 _5358_ (.A(_1801_),
    .B(_1809_),
    .C(_1817_),
    .X(_1818_));
 sg13g2_nor2_1 _5359_ (.A(_1073_),
    .B(_1096_),
    .Y(_1819_));
 sg13g2_nand2b_1 _5360_ (.Y(_1820_),
    .B(_1747_),
    .A_N(_1132_));
 sg13g2_nand3_1 _5361_ (.B(net25),
    .C(_1820_),
    .A(net159),
    .Y(_1821_));
 sg13g2_nand2_1 _5362_ (.Y(_1822_),
    .A(_1132_),
    .B(net24));
 sg13g2_nor2_1 _5363_ (.A(net24),
    .B(net25),
    .Y(_1823_));
 sg13g2_a21oi_1 _5364_ (.A1(_1819_),
    .A2(_1822_),
    .Y(_1824_),
    .B1(_1823_));
 sg13g2_a21oi_1 _5365_ (.A1(_1819_),
    .A2(_1821_),
    .Y(_1825_),
    .B1(_1824_));
 sg13g2_and2_1 _5366_ (.A(_2759_),
    .B(net111),
    .X(_1826_));
 sg13g2_a22oi_1 _5367_ (.Y(_1827_),
    .B1(_1826_),
    .B2(_1744_),
    .A2(_1745_),
    .A1(_1743_));
 sg13g2_nor2b_1 _5368_ (.A(net36),
    .B_N(net159),
    .Y(_1828_));
 sg13g2_nand2b_1 _5369_ (.Y(_1829_),
    .B(net57),
    .A_N(_1828_));
 sg13g2_o21ai_1 _5370_ (.B1(_2764_),
    .Y(_1830_),
    .A1(_2761_),
    .A2(net59));
 sg13g2_nor2b_1 _5371_ (.A(net159),
    .B_N(net36),
    .Y(_1831_));
 sg13g2_a21oi_1 _5372_ (.A1(_1828_),
    .A2(_1830_),
    .Y(_1832_),
    .B1(_1831_));
 sg13g2_o21ai_1 _5373_ (.B1(_1832_),
    .Y(_1833_),
    .A1(_1827_),
    .A2(_1829_));
 sg13g2_nor2_1 _5374_ (.A(_1126_),
    .B(_1830_),
    .Y(_1834_));
 sg13g2_xnor2_1 _5375_ (.Y(_1835_),
    .A(net23),
    .B(_1834_));
 sg13g2_and3_1 _5376_ (.X(_1836_),
    .A(_1765_),
    .B(_1833_),
    .C(_1835_));
 sg13g2_xor2_1 _5377_ (.B(_1625_),
    .A(net73),
    .X(_1837_));
 sg13g2_or3_1 _5378_ (.A(_1096_),
    .B(_1132_),
    .C(_1722_),
    .X(_1838_));
 sg13g2_buf_1 _5379_ (.A(_1838_),
    .X(_1839_));
 sg13g2_xnor2_1 _5380_ (.Y(_1840_),
    .A(_1111_),
    .B(_1753_));
 sg13g2_nand3_1 _5381_ (.B(_1839_),
    .C(_1840_),
    .A(_2889_),
    .Y(_1841_));
 sg13g2_nand3_1 _5382_ (.B(_1753_),
    .C(_1837_),
    .A(_1073_),
    .Y(_1842_));
 sg13g2_o21ai_1 _5383_ (.B1(_1842_),
    .Y(_1843_),
    .A1(_1837_),
    .A2(_1841_));
 sg13g2_xor2_1 _5384_ (.B(_1666_),
    .A(net72),
    .X(_1844_));
 sg13g2_xor2_1 _5385_ (.B(_1844_),
    .A(_1144_),
    .X(_1845_));
 sg13g2_xor2_1 _5386_ (.B(net113),
    .A(net61),
    .X(_1846_));
 sg13g2_and2_1 _5387_ (.A(net73),
    .B(net56),
    .X(_1847_));
 sg13g2_buf_1 _5388_ (.A(_1847_),
    .X(_1848_));
 sg13g2_nand2b_1 _5389_ (.Y(_1849_),
    .B(_0092_),
    .A_N(net59));
 sg13g2_nand3_1 _5390_ (.B(_1848_),
    .C(_1849_),
    .A(net60),
    .Y(_1850_));
 sg13g2_nor3_1 _5391_ (.A(_1845_),
    .B(_1846_),
    .C(_1850_),
    .Y(_1851_));
 sg13g2_nand3_1 _5392_ (.B(_1846_),
    .C(_1850_),
    .A(_1844_),
    .Y(_1852_));
 sg13g2_nand2b_1 _5393_ (.Y(_1853_),
    .B(_1852_),
    .A_N(_1851_));
 sg13g2_nand4_1 _5394_ (.B(_1836_),
    .C(_1843_),
    .A(_1825_),
    .Y(_1854_),
    .D(_1853_));
 sg13g2_o21ai_1 _5395_ (.B1(_1854_),
    .Y(_1855_),
    .A1(_1796_),
    .A2(_1818_));
 sg13g2_nand2_1 _5396_ (.Y(_1856_),
    .A(net38),
    .B(_1848_));
 sg13g2_a21oi_1 _5397_ (.A1(_1700_),
    .A2(_1703_),
    .Y(_1857_),
    .B1(_1856_));
 sg13g2_and3_1 _5398_ (.X(_1858_),
    .A(_2764_),
    .B(net118),
    .C(_1737_));
 sg13g2_nor3_1 _5399_ (.A(net37),
    .B(net118),
    .C(_1737_),
    .Y(_1859_));
 sg13g2_o21ai_1 _5400_ (.B1(_1839_),
    .Y(_1860_),
    .A1(_1858_),
    .A2(_1859_));
 sg13g2_o21ai_1 _5401_ (.B1(net35),
    .Y(_1861_),
    .A1(_1857_),
    .A2(_1860_));
 sg13g2_o21ai_1 _5402_ (.B1(net25),
    .Y(_1862_),
    .A1(_1132_),
    .A2(_1720_));
 sg13g2_a21oi_1 _5403_ (.A1(_1848_),
    .A2(_1862_),
    .Y(_1863_),
    .B1(_1724_));
 sg13g2_nor2_1 _5404_ (.A(_2757_),
    .B(_1863_),
    .Y(_1864_));
 sg13g2_o21ai_1 _5405_ (.B1(_1707_),
    .Y(_1865_),
    .A1(_1082_),
    .A2(_1102_));
 sg13g2_inv_1 _5406_ (.Y(_1866_),
    .A(_1776_));
 sg13g2_a21oi_1 _5407_ (.A1(_1731_),
    .A2(_1837_),
    .Y(_1867_),
    .B1(net59));
 sg13g2_nor3_1 _5408_ (.A(_1775_),
    .B(_1866_),
    .C(_1867_),
    .Y(_1868_));
 sg13g2_nand2_1 _5409_ (.Y(_1869_),
    .A(_1865_),
    .B(_1868_));
 sg13g2_a21oi_1 _5410_ (.A1(_1111_),
    .A2(_1714_),
    .Y(_1870_),
    .B1(_2757_));
 sg13g2_a21oi_1 _5411_ (.A1(_1753_),
    .A2(_1823_),
    .Y(_1871_),
    .B1(_1870_));
 sg13g2_a21oi_1 _5412_ (.A1(_1132_),
    .A2(net24),
    .Y(_1872_),
    .B1(_1096_));
 sg13g2_nor2_1 _5413_ (.A(_1082_),
    .B(_1126_),
    .Y(_1873_));
 sg13g2_xnor2_1 _5414_ (.Y(_1874_),
    .A(net23),
    .B(_1873_));
 sg13g2_o21ai_1 _5415_ (.B1(_1874_),
    .Y(_1875_),
    .A1(_1823_),
    .A2(_1872_));
 sg13g2_nor4_1 _5416_ (.A(_1864_),
    .B(_1869_),
    .C(_1871_),
    .D(_1875_),
    .Y(_1876_));
 sg13g2_inv_1 _5417_ (.Y(_1877_),
    .A(net121));
 sg13g2_nand2_1 _5418_ (.Y(_1878_),
    .A(_1877_),
    .B(_1837_));
 sg13g2_a21oi_1 _5419_ (.A1(net23),
    .A2(_1802_),
    .Y(_1879_),
    .B1(_1731_));
 sg13g2_nor3_1 _5420_ (.A(net59),
    .B(_1877_),
    .C(_1837_),
    .Y(_1880_));
 sg13g2_o21ai_1 _5421_ (.B1(_1880_),
    .Y(_1881_),
    .A1(net37),
    .A2(_1879_));
 sg13g2_o21ai_1 _5422_ (.B1(_1881_),
    .Y(_1882_),
    .A1(_0300_),
    .A2(_1878_));
 sg13g2_and3_1 _5423_ (.X(_1883_),
    .A(_2757_),
    .B(_1136_),
    .C(_1122_));
 sg13g2_a21oi_1 _5424_ (.A1(_2757_),
    .A2(_1136_),
    .Y(_1884_),
    .B1(_1720_));
 sg13g2_a21oi_1 _5425_ (.A1(net24),
    .A2(_1883_),
    .Y(_1885_),
    .B1(_1884_));
 sg13g2_nor2_1 _5426_ (.A(net53),
    .B(_2749_),
    .Y(_1886_));
 sg13g2_nand3_1 _5427_ (.B(_1750_),
    .C(_1886_),
    .A(_1105_),
    .Y(_1887_));
 sg13g2_a21oi_1 _5428_ (.A1(_1799_),
    .A2(_1887_),
    .Y(_1888_),
    .B1(net35));
 sg13g2_nand2_1 _5429_ (.Y(_1889_),
    .A(_1114_),
    .B(_1747_));
 sg13g2_o21ai_1 _5430_ (.B1(_1889_),
    .Y(_1890_),
    .A1(_1885_),
    .A2(_1888_));
 sg13g2_o21ai_1 _5431_ (.B1(_1714_),
    .Y(_1891_),
    .A1(net59),
    .A2(_1114_));
 sg13g2_or2_1 _5432_ (.X(_1892_),
    .B(net73),
    .A(net74));
 sg13g2_o21ai_1 _5433_ (.B1(_1892_),
    .Y(_1893_),
    .A1(_1733_),
    .A2(_1737_));
 sg13g2_a21o_1 _5434_ (.A2(_1091_),
    .A1(_2757_),
    .B1(_1727_),
    .X(_1894_));
 sg13g2_nand3_1 _5435_ (.B(_1091_),
    .C(_1727_),
    .A(_2757_),
    .Y(_1895_));
 sg13g2_nand4_1 _5436_ (.B(_1893_),
    .C(_1894_),
    .A(_1891_),
    .Y(_1896_),
    .D(_1895_));
 sg13g2_nor3_1 _5437_ (.A(net36),
    .B(_2753_),
    .C(_1892_),
    .Y(_1897_));
 sg13g2_xnor2_1 _5438_ (.Y(_1898_),
    .A(_1706_),
    .B(_1897_));
 sg13g2_nor3_1 _5439_ (.A(_2759_),
    .B(_2885_),
    .C(_2886_),
    .Y(_1899_));
 sg13g2_nand3_1 _5440_ (.B(_1886_),
    .C(_1899_),
    .A(_1105_),
    .Y(_1900_));
 sg13g2_xor2_1 _5441_ (.B(_1900_),
    .A(_1702_),
    .X(_1901_));
 sg13g2_nor4_1 _5442_ (.A(_1775_),
    .B(_1896_),
    .C(_1898_),
    .D(_1901_),
    .Y(_1902_));
 sg13g2_and3_1 _5443_ (.X(_1903_),
    .A(_1882_),
    .B(_1890_),
    .C(_1902_));
 sg13g2_a21o_1 _5444_ (.A2(_1876_),
    .A1(_1861_),
    .B1(_1903_),
    .X(_1904_));
 sg13g2_xnor2_1 _5445_ (.Y(_1905_),
    .A(_0492_),
    .B(_1581_));
 sg13g2_buf_2 _5446_ (.A(_1905_),
    .X(_1906_));
 sg13g2_xor2_1 _5447_ (.B(_1576_),
    .A(_1023_),
    .X(_1907_));
 sg13g2_buf_2 _5448_ (.A(_1907_),
    .X(_1908_));
 sg13g2_o21ai_1 _5449_ (.B1(_1908_),
    .Y(_1909_),
    .A1(net48),
    .A2(_1906_));
 sg13g2_xnor2_1 _5450_ (.Y(_1910_),
    .A(_0090_),
    .B(_0106_));
 sg13g2_inv_1 _5451_ (.Y(_1911_),
    .A(_1910_));
 sg13g2_xor2_1 _5452_ (.B(_1581_),
    .A(_0492_),
    .X(_1912_));
 sg13g2_buf_2 _5453_ (.A(_1912_),
    .X(_1913_));
 sg13g2_nor2_1 _5454_ (.A(_1913_),
    .B(_1908_),
    .Y(_1914_));
 sg13g2_buf_1 _5455_ (.A(_1910_),
    .X(_1915_));
 sg13g2_nand4_1 _5456_ (.B(_1046_),
    .C(_1048_),
    .A(net49),
    .Y(_1916_),
    .D(net39));
 sg13g2_o21ai_1 _5457_ (.B1(_1916_),
    .Y(_1917_),
    .A1(_1025_),
    .A2(_1914_));
 sg13g2_a221oi_1 _5458_ (.B2(_1049_),
    .C1(_1917_),
    .B1(_1911_),
    .A1(_1025_),
    .Y(_1918_),
    .A2(_1909_));
 sg13g2_xor2_1 _5459_ (.B(_1007_),
    .A(_1548_),
    .X(_1919_));
 sg13g2_buf_2 _5460_ (.A(_1919_),
    .X(_1920_));
 sg13g2_nand2_1 _5461_ (.Y(_1921_),
    .A(net42),
    .B(net48));
 sg13g2_o21ai_1 _5462_ (.B1(_1920_),
    .Y(_1922_),
    .A1(_1921_),
    .A2(_1913_));
 sg13g2_mux2_1 _5463_ (.A0(_1920_),
    .A1(_1922_),
    .S(_1016_),
    .X(_1923_));
 sg13g2_nor2b_1 _5464_ (.A(_3050_),
    .B_N(_1528_),
    .Y(_1924_));
 sg13g2_buf_1 _5465_ (.A(_0109_),
    .X(_1925_));
 sg13g2_xor2_1 _5466_ (.B(_1925_),
    .A(net43),
    .X(_1926_));
 sg13g2_nor2b_1 _5467_ (.A(net126),
    .B_N(_3050_),
    .Y(_1927_));
 sg13g2_nor2b_1 _5468_ (.A(_1926_),
    .B_N(_1927_),
    .Y(_1928_));
 sg13g2_a21oi_1 _5469_ (.A1(_1924_),
    .A2(_1926_),
    .Y(_1929_),
    .B1(_1928_));
 sg13g2_xor2_1 _5470_ (.B(_1566_),
    .A(_0995_),
    .X(_1930_));
 sg13g2_buf_1 _5471_ (.A(_1930_),
    .X(_1931_));
 sg13g2_xnor2_1 _5472_ (.Y(_1932_),
    .A(_3054_),
    .B(net22));
 sg13g2_nor3_1 _5473_ (.A(_1923_),
    .B(_1929_),
    .C(_1932_),
    .Y(_1933_));
 sg13g2_xnor2_1 _5474_ (.Y(_1934_),
    .A(_1053_),
    .B(_1589_));
 sg13g2_buf_1 _5475_ (.A(_1934_),
    .X(_1935_));
 sg13g2_or3_1 _5476_ (.A(net47),
    .B(_1056_),
    .C(net21),
    .X(_1936_));
 sg13g2_nand2_1 _5477_ (.Y(_1937_),
    .A(_1056_),
    .B(net21));
 sg13g2_xnor2_1 _5478_ (.Y(_1938_),
    .A(_0496_),
    .B(net163));
 sg13g2_buf_2 _5479_ (.A(_1938_),
    .X(_1939_));
 sg13g2_xnor2_1 _5480_ (.Y(_1940_),
    .A(net66),
    .B(net164));
 sg13g2_nand3_1 _5481_ (.B(_1939_),
    .C(_1940_),
    .A(_1013_),
    .Y(_1941_));
 sg13g2_xor2_1 _5482_ (.B(net164),
    .A(net66),
    .X(_1942_));
 sg13g2_xor2_1 _5483_ (.B(_1939_),
    .A(net27),
    .X(_1943_));
 sg13g2_nand3_1 _5484_ (.B(_1942_),
    .C(_1943_),
    .A(_3053_),
    .Y(_1944_));
 sg13g2_a22oi_1 _5485_ (.Y(_1945_),
    .B1(_1941_),
    .B2(_1944_),
    .A2(_1937_),
    .A1(_1936_));
 sg13g2_nand3_1 _5486_ (.B(_1933_),
    .C(_1945_),
    .A(_1918_),
    .Y(_1946_));
 sg13g2_xnor2_1 _5487_ (.Y(_1947_),
    .A(_1548_),
    .B(_1007_));
 sg13g2_buf_2 _5488_ (.A(_1947_),
    .X(_1948_));
 sg13g2_nor3_2 _5489_ (.A(net51),
    .B(net50),
    .C(net46),
    .Y(_1949_));
 sg13g2_nor2_1 _5490_ (.A(_1949_),
    .B(_1920_),
    .Y(_1950_));
 sg13g2_a221oi_1 _5491_ (.B2(_1009_),
    .C1(_1950_),
    .B1(_1948_),
    .A1(_1169_),
    .Y(_1951_),
    .A2(_1011_));
 sg13g2_nor2_1 _5492_ (.A(net16),
    .B(_1920_),
    .Y(_1952_));
 sg13g2_o21ai_1 _5493_ (.B1(_1939_),
    .Y(_1953_),
    .A1(net27),
    .A2(_1952_));
 sg13g2_a21oi_1 _5494_ (.A1(_3057_),
    .A2(_3045_),
    .Y(_1954_),
    .B1(_1010_));
 sg13g2_nor2b_1 _5495_ (.A(_1939_),
    .B_N(_0501_),
    .Y(_1955_));
 sg13g2_o21ai_1 _5496_ (.B1(_1955_),
    .Y(_1956_),
    .A1(_1950_),
    .A2(_1954_));
 sg13g2_o21ai_1 _5497_ (.B1(_1956_),
    .Y(_1957_),
    .A1(_1951_),
    .A2(_1953_));
 sg13g2_nand2_1 _5498_ (.Y(_1958_),
    .A(net21),
    .B(_1906_));
 sg13g2_o21ai_1 _5499_ (.B1(_1913_),
    .Y(_1959_),
    .A1(_0461_),
    .A2(net21));
 sg13g2_mux2_1 _5500_ (.A0(_1958_),
    .A1(_1959_),
    .S(_1033_),
    .X(_1960_));
 sg13g2_nand2b_1 _5501_ (.Y(_1961_),
    .B(_1948_),
    .A_N(net32));
 sg13g2_nand3_1 _5502_ (.B(net22),
    .C(_1961_),
    .A(_1000_),
    .Y(_1962_));
 sg13g2_xnor2_1 _5503_ (.Y(_1963_),
    .A(_0995_),
    .B(_1566_));
 sg13g2_nand4_1 _5504_ (.B(net21),
    .C(_1906_),
    .A(_1002_),
    .Y(_1964_),
    .D(_1963_));
 sg13g2_o21ai_1 _5505_ (.B1(_1964_),
    .Y(_1965_),
    .A1(_1960_),
    .A2(_1962_));
 sg13g2_xnor2_1 _5506_ (.Y(_1966_),
    .A(_1042_),
    .B(_1911_));
 sg13g2_nor3_1 _5507_ (.A(_0465_),
    .B(net68),
    .C(_3043_),
    .Y(_1967_));
 sg13g2_xnor2_1 _5508_ (.Y(_1968_),
    .A(_1023_),
    .B(_1576_));
 sg13g2_a21oi_1 _5509_ (.A1(_1967_),
    .A2(net21),
    .Y(_1969_),
    .B1(_1968_));
 sg13g2_nand2b_1 _5510_ (.Y(_1970_),
    .B(_1969_),
    .A_N(_1029_));
 sg13g2_nand3_1 _5511_ (.B(_1968_),
    .C(net39),
    .A(_1029_),
    .Y(_1971_));
 sg13g2_o21ai_1 _5512_ (.B1(_1971_),
    .Y(_1972_),
    .A1(_1966_),
    .A2(_1970_));
 sg13g2_nand3_1 _5513_ (.B(_1926_),
    .C(_1940_),
    .A(net49),
    .Y(_1973_));
 sg13g2_and2_1 _5514_ (.A(_0969_),
    .B(_1925_),
    .X(_1974_));
 sg13g2_nor2_1 _5515_ (.A(net43),
    .B(_1925_),
    .Y(_1975_));
 sg13g2_mux2_1 _5516_ (.A0(_1974_),
    .A1(_1975_),
    .S(_1942_),
    .X(_1976_));
 sg13g2_nand2_1 _5517_ (.Y(_1977_),
    .A(_1924_),
    .B(_1976_));
 sg13g2_o21ai_1 _5518_ (.B1(_1977_),
    .Y(_1978_),
    .A1(net126),
    .A2(_1973_));
 sg13g2_nand4_1 _5519_ (.B(_1965_),
    .C(_1972_),
    .A(_1957_),
    .Y(_1979_),
    .D(_1978_));
 sg13g2_nor2_1 _5520_ (.A(_1924_),
    .B(_1927_),
    .Y(_1980_));
 sg13g2_nor4_1 _5521_ (.A(_0486_),
    .B(net42),
    .C(net32),
    .D(_0463_),
    .Y(_1981_));
 sg13g2_xnor2_1 _5522_ (.Y(_1982_),
    .A(_0465_),
    .B(_1906_));
 sg13g2_nand2_1 _5523_ (.Y(_1983_),
    .A(_1969_),
    .B(_1982_));
 sg13g2_nand2_1 _5524_ (.Y(_1984_),
    .A(_0487_),
    .B(_1920_));
 sg13g2_nor2_1 _5525_ (.A(_1006_),
    .B(_0467_),
    .Y(_1985_));
 sg13g2_a21o_1 _5526_ (.A2(_1985_),
    .A1(_1967_),
    .B1(_1935_),
    .X(_1986_));
 sg13g2_nand4_1 _5527_ (.B(_1931_),
    .C(_1984_),
    .A(_0464_),
    .Y(_1987_),
    .D(_1986_));
 sg13g2_xor2_1 _5528_ (.B(_1589_),
    .A(_1053_),
    .X(_1988_));
 sg13g2_or4_1 _5529_ (.A(_0464_),
    .B(_1988_),
    .C(_1920_),
    .D(_1931_),
    .X(_1989_));
 sg13g2_nand2b_1 _5530_ (.Y(_1990_),
    .B(_1527_),
    .A_N(net43));
 sg13g2_xor2_1 _5531_ (.B(net164),
    .A(net50),
    .X(_1991_));
 sg13g2_nor2_1 _5532_ (.A(_1990_),
    .B(_1991_),
    .Y(_1992_));
 sg13g2_a22oi_1 _5533_ (.Y(_1993_),
    .B1(_1948_),
    .B2(_1949_),
    .A2(_1028_),
    .A1(_3045_));
 sg13g2_nand2b_1 _5534_ (.Y(_1994_),
    .B(net43),
    .A_N(_1527_));
 sg13g2_xnor2_1 _5535_ (.Y(_1995_),
    .A(net50),
    .B(net164));
 sg13g2_nor2_1 _5536_ (.A(_1994_),
    .B(_1995_),
    .Y(_1996_));
 sg13g2_a21oi_1 _5537_ (.A1(_1992_),
    .A2(_1993_),
    .Y(_1997_),
    .B1(_1996_));
 sg13g2_a221oi_1 _5538_ (.B2(_1989_),
    .C1(_1997_),
    .B1(_1987_),
    .A1(_1981_),
    .Y(_1998_),
    .A2(_1983_));
 sg13g2_nor2_1 _5539_ (.A(_1914_),
    .B(_1981_),
    .Y(_1999_));
 sg13g2_xnor2_1 _5540_ (.Y(_2000_),
    .A(net51),
    .B(net163));
 sg13g2_xnor2_1 _5541_ (.Y(_2001_),
    .A(_0463_),
    .B(_2000_));
 sg13g2_nor2_1 _5542_ (.A(_1999_),
    .B(_2001_),
    .Y(_2002_));
 sg13g2_nor2_1 _5543_ (.A(_0970_),
    .B(_1042_),
    .Y(_2003_));
 sg13g2_xnor2_1 _5544_ (.Y(_2004_),
    .A(_1911_),
    .B(_2003_));
 sg13g2_nand4_1 _5545_ (.B(_1998_),
    .C(_2002_),
    .A(_1980_),
    .Y(_2005_),
    .D(_2004_));
 sg13g2_and3_1 _5546_ (.X(_2006_),
    .A(net42),
    .B(_1046_),
    .C(_1908_));
 sg13g2_nor3_1 _5547_ (.A(net42),
    .B(_1046_),
    .C(_1908_),
    .Y(_2007_));
 sg13g2_o21ai_1 _5548_ (.B1(_1548_),
    .Y(_2008_),
    .A1(_2006_),
    .A2(_2007_));
 sg13g2_xnor2_1 _5549_ (.Y(_2009_),
    .A(_3057_),
    .B(_1046_));
 sg13g2_nand3b_1 _5550_ (.B(_1968_),
    .C(_2009_),
    .Y(_2010_),
    .A_N(_1548_));
 sg13g2_nand2_1 _5551_ (.Y(_2011_),
    .A(_0489_),
    .B(_1046_));
 sg13g2_nand3_1 _5552_ (.B(_1906_),
    .C(_1915_),
    .A(_2011_),
    .Y(_2012_));
 sg13g2_xor2_1 _5553_ (.B(_1915_),
    .A(_3042_),
    .X(_2013_));
 sg13g2_nand4_1 _5554_ (.B(_1046_),
    .C(_1913_),
    .A(_0489_),
    .Y(_2014_),
    .D(_2013_));
 sg13g2_a22oi_1 _5555_ (.Y(_2015_),
    .B1(_2012_),
    .B2(_2014_),
    .A2(_2010_),
    .A1(_2008_));
 sg13g2_nand3_1 _5556_ (.B(net163),
    .C(_1930_),
    .A(net33),
    .Y(_2016_));
 sg13g2_inv_1 _5557_ (.Y(_2017_),
    .A(net51));
 sg13g2_inv_1 _5558_ (.Y(_2018_),
    .A(net163));
 sg13g2_nand3_1 _5559_ (.B(_2018_),
    .C(_1963_),
    .A(_2017_),
    .Y(_2019_));
 sg13g2_a21o_1 _5560_ (.A2(_2019_),
    .A1(_2016_),
    .B1(_0988_),
    .X(_2020_));
 sg13g2_nor2_1 _5561_ (.A(net22),
    .B(_2000_),
    .Y(_2021_));
 sg13g2_nand2_1 _5562_ (.Y(_2022_),
    .A(_0988_),
    .B(_2021_));
 sg13g2_nand3_1 _5563_ (.B(_1055_),
    .C(_1048_),
    .A(net45),
    .Y(_2023_));
 sg13g2_or2_1 _5564_ (.X(_2024_),
    .B(_1589_),
    .A(net47));
 sg13g2_buf_1 _5565_ (.A(_2024_),
    .X(_2025_));
 sg13g2_nand2_1 _5566_ (.Y(_2026_),
    .A(_0970_),
    .B(_2025_));
 sg13g2_nand3b_1 _5567_ (.B(_1980_),
    .C(_2026_),
    .Y(_2027_),
    .A_N(_2023_));
 sg13g2_nand3_1 _5568_ (.B(_1980_),
    .C(_2025_),
    .A(_2023_),
    .Y(_2028_));
 sg13g2_a21oi_1 _5569_ (.A1(net47),
    .A2(_1589_),
    .Y(_2029_),
    .B1(_1994_));
 sg13g2_xor2_1 _5570_ (.B(_1589_),
    .A(net47),
    .X(_2030_));
 sg13g2_nor2_1 _5571_ (.A(_1990_),
    .B(_1995_),
    .Y(_2031_));
 sg13g2_a22oi_1 _5572_ (.Y(_2032_),
    .B1(_2030_),
    .B2(_2031_),
    .A2(_2029_),
    .A1(_1995_));
 sg13g2_a221oi_1 _5573_ (.B2(_2028_),
    .C1(_2032_),
    .B1(_2027_),
    .A1(_2020_),
    .Y(_2033_),
    .A2(_2022_));
 sg13g2_nand3_1 _5574_ (.B(_1990_),
    .C(_1994_),
    .A(_1980_),
    .Y(_2034_));
 sg13g2_xnor2_1 _5575_ (.Y(_2035_),
    .A(net125),
    .B(_3049_));
 sg13g2_xnor2_1 _5576_ (.Y(_2036_),
    .A(_1537_),
    .B(_0491_));
 sg13g2_xnor2_1 _5577_ (.Y(_2037_),
    .A(net166),
    .B(net47));
 sg13g2_xnor2_1 _5578_ (.Y(_2038_),
    .A(_1531_),
    .B(net51));
 sg13g2_nand4_1 _5579_ (.B(_2036_),
    .C(_2037_),
    .A(_2035_),
    .Y(_2039_),
    .D(_2038_));
 sg13g2_xnor2_1 _5580_ (.Y(_2040_),
    .A(_1541_),
    .B(_3042_));
 sg13g2_xnor2_1 _5581_ (.Y(_2041_),
    .A(net162),
    .B(_1006_));
 sg13g2_xnor2_1 _5582_ (.Y(_2042_),
    .A(_1542_),
    .B(net48));
 sg13g2_xnor2_1 _5583_ (.Y(_2043_),
    .A(net127),
    .B(_0487_));
 sg13g2_nand4_1 _5584_ (.B(_2041_),
    .C(_2042_),
    .A(_2040_),
    .Y(_2044_),
    .D(_2043_));
 sg13g2_nor3_1 _5585_ (.A(_2034_),
    .B(_2039_),
    .C(_2044_),
    .Y(_2045_));
 sg13g2_a21oi_1 _5586_ (.A1(_2015_),
    .A2(_2033_),
    .Y(_2046_),
    .B1(_2045_));
 sg13g2_nand4_1 _5587_ (.B(_1979_),
    .C(_2005_),
    .A(_1946_),
    .Y(_2047_),
    .D(_2046_));
 sg13g2_o21ai_1 _5588_ (.B1(_2047_),
    .Y(_2048_),
    .A1(_1855_),
    .A2(_1904_));
 sg13g2_a21oi_1 _5589_ (.A1(_0489_),
    .A2(_1055_),
    .Y(_2049_),
    .B1(_1913_));
 sg13g2_nor3_1 _5590_ (.A(_1921_),
    .B(_1015_),
    .C(_1906_),
    .Y(_2050_));
 sg13g2_o21ai_1 _5591_ (.B1(_1995_),
    .Y(_2051_),
    .A1(_2049_),
    .A2(_2050_));
 sg13g2_nand3_1 _5592_ (.B(_1906_),
    .C(_1991_),
    .A(net16),
    .Y(_2052_));
 sg13g2_o21ai_1 _5593_ (.B1(_2052_),
    .Y(_2053_),
    .A1(net16),
    .A2(_2051_));
 sg13g2_a21oi_1 _5594_ (.A1(net27),
    .A2(_1009_),
    .Y(_2054_),
    .B1(net163));
 sg13g2_nor2_1 _5595_ (.A(net22),
    .B(_2054_),
    .Y(_2055_));
 sg13g2_xnor2_1 _5596_ (.Y(_2056_),
    .A(_2017_),
    .B(_2055_));
 sg13g2_nor2_1 _5597_ (.A(net16),
    .B(_1024_),
    .Y(_2057_));
 sg13g2_xnor2_1 _5598_ (.Y(_2058_),
    .A(_1908_),
    .B(_2057_));
 sg13g2_nand3b_1 _5599_ (.B(net49),
    .C(_1926_),
    .Y(_2059_),
    .A_N(net126));
 sg13g2_nor2_1 _5600_ (.A(_0460_),
    .B(_1926_),
    .Y(_2060_));
 sg13g2_nand2_1 _5601_ (.Y(_2061_),
    .A(net126),
    .B(_2060_));
 sg13g2_a22oi_1 _5602_ (.Y(_2062_),
    .B1(_2059_),
    .B2(_2061_),
    .A2(_1589_),
    .A1(net47));
 sg13g2_nand4_1 _5603_ (.B(_2056_),
    .C(_2058_),
    .A(_2053_),
    .Y(_2063_),
    .D(_2062_));
 sg13g2_nand2_1 _5604_ (.Y(_2064_),
    .A(_1055_),
    .B(_1048_));
 sg13g2_o21ai_1 _5605_ (.B1(net39),
    .Y(_2065_),
    .A1(net16),
    .A2(_2064_));
 sg13g2_nand3_1 _5606_ (.B(net48),
    .C(net68),
    .A(net42),
    .Y(_2066_));
 sg13g2_nor4_1 _5607_ (.A(_0997_),
    .B(_1015_),
    .C(_2066_),
    .D(_1910_),
    .Y(_2067_));
 sg13g2_nand2b_1 _5608_ (.Y(_2068_),
    .B(_2067_),
    .A_N(net45));
 sg13g2_nand3_1 _5609_ (.B(_2065_),
    .C(_2068_),
    .A(_2025_),
    .Y(_2069_));
 sg13g2_a21o_1 _5610_ (.A2(_2067_),
    .A1(net45),
    .B1(_2025_),
    .X(_2070_));
 sg13g2_xor2_1 _5611_ (.B(net42),
    .A(_1548_),
    .X(_2071_));
 sg13g2_xnor2_1 _5612_ (.Y(_2072_),
    .A(_1015_),
    .B(_2071_));
 sg13g2_and2_1 _5613_ (.A(net50),
    .B(net163),
    .X(_2073_));
 sg13g2_buf_1 _5614_ (.A(_2073_),
    .X(_2074_));
 sg13g2_and2_1 _5615_ (.A(net22),
    .B(_2074_),
    .X(_2075_));
 sg13g2_nor4_1 _5616_ (.A(_1015_),
    .B(net22),
    .C(_2074_),
    .D(_2071_),
    .Y(_2076_));
 sg13g2_a21oi_1 _5617_ (.A1(_2072_),
    .A2(_2075_),
    .Y(_2077_),
    .B1(_2076_));
 sg13g2_o21ai_1 _5618_ (.B1(_1009_),
    .Y(_2078_),
    .A1(_1055_),
    .A2(_2074_));
 sg13g2_nand3_1 _5619_ (.B(_2071_),
    .C(_2078_),
    .A(_1963_),
    .Y(_2079_));
 sg13g2_o21ai_1 _5620_ (.B1(_2079_),
    .Y(_2080_),
    .A1(net16),
    .A2(_2077_));
 sg13g2_nand3_1 _5621_ (.B(_2070_),
    .C(_2080_),
    .A(_2069_),
    .Y(_2081_));
 sg13g2_nand4_1 _5622_ (.B(_1028_),
    .C(_1908_),
    .A(_1041_),
    .Y(_2082_),
    .D(net39));
 sg13g2_a21oi_1 _5623_ (.A1(_3053_),
    .A2(_2082_),
    .Y(_2083_),
    .B1(_1010_));
 sg13g2_nand3_1 _5624_ (.B(_1028_),
    .C(net39),
    .A(_1041_),
    .Y(_2084_));
 sg13g2_a21oi_1 _5625_ (.A1(_3057_),
    .A2(_3045_),
    .Y(_2085_),
    .B1(_1948_));
 sg13g2_nand4_1 _5626_ (.B(_1949_),
    .C(_2084_),
    .A(_1013_),
    .Y(_2086_),
    .D(_2085_));
 sg13g2_o21ai_1 _5627_ (.B1(_2086_),
    .Y(_2087_),
    .A1(_1920_),
    .A2(_2083_));
 sg13g2_nor2b_1 _5628_ (.A(net164),
    .B_N(net27),
    .Y(_2088_));
 sg13g2_a22oi_1 _5629_ (.Y(_2089_),
    .B1(_1927_),
    .B2(_1975_),
    .A2(_1926_),
    .A1(_1924_));
 sg13g2_nand2_1 _5630_ (.Y(_2090_),
    .A(net27),
    .B(net164));
 sg13g2_nand3_1 _5631_ (.B(_1974_),
    .C(_2090_),
    .A(_1927_),
    .Y(_2091_));
 sg13g2_o21ai_1 _5632_ (.B1(_2091_),
    .Y(_2092_),
    .A1(_2088_),
    .A2(_2089_));
 sg13g2_or2_1 _5633_ (.X(_2093_),
    .B(_1939_),
    .A(net66));
 sg13g2_nand2_1 _5634_ (.Y(_2094_),
    .A(_1013_),
    .B(_1028_));
 sg13g2_xnor2_1 _5635_ (.Y(_2095_),
    .A(_1968_),
    .B(_2094_));
 sg13g2_and3_1 _5636_ (.X(_2096_),
    .A(_2092_),
    .B(_2093_),
    .C(_2095_));
 sg13g2_nand2_1 _5637_ (.Y(_2097_),
    .A(net66),
    .B(_1939_));
 sg13g2_nor3_1 _5638_ (.A(net33),
    .B(_3053_),
    .C(_1963_),
    .Y(_2098_));
 sg13g2_a22oi_1 _5639_ (.Y(_2099_),
    .B1(_2097_),
    .B2(_2098_),
    .A2(_1963_),
    .A1(_3053_));
 sg13g2_nand3b_1 _5640_ (.B(_1963_),
    .C(_2097_),
    .Y(_2100_),
    .A_N(_0998_));
 sg13g2_o21ai_1 _5641_ (.B1(_2100_),
    .Y(_2101_),
    .A1(net27),
    .A2(_2099_));
 sg13g2_nand3_1 _5642_ (.B(_1013_),
    .C(_1028_),
    .A(_1041_),
    .Y(_2102_));
 sg13g2_nand3_1 _5643_ (.B(net39),
    .C(_2102_),
    .A(net21),
    .Y(_2103_));
 sg13g2_xnor2_1 _5644_ (.Y(_2104_),
    .A(net45),
    .B(net21));
 sg13g2_nand2b_1 _5645_ (.Y(_2105_),
    .B(_2104_),
    .A_N(_2102_));
 sg13g2_nand3_1 _5646_ (.B(_3053_),
    .C(_1939_),
    .A(net164),
    .Y(_2106_));
 sg13g2_inv_1 _5647_ (.Y(_2107_),
    .A(net164));
 sg13g2_a21oi_1 _5648_ (.A1(_2107_),
    .A2(_1013_),
    .Y(_2108_),
    .B1(net27));
 sg13g2_nand3b_1 _5649_ (.B(net28),
    .C(net49),
    .Y(_2109_),
    .A_N(net50));
 sg13g2_nand4_1 _5650_ (.B(net66),
    .C(_1033_),
    .A(_2017_),
    .Y(_2110_),
    .D(_2109_));
 sg13g2_xnor2_1 _5651_ (.Y(_2111_),
    .A(_1913_),
    .B(_2110_));
 sg13g2_a221oi_1 _5652_ (.B2(_2108_),
    .C1(_2111_),
    .B1(_2106_),
    .A1(_2103_),
    .Y(_2112_),
    .A2(_2105_));
 sg13g2_nand4_1 _5653_ (.B(_2096_),
    .C(_2101_),
    .A(_2087_),
    .Y(_2113_),
    .D(_2112_));
 sg13g2_o21ai_1 _5654_ (.B1(_2113_),
    .Y(_2114_),
    .A1(_2063_),
    .A2(_2081_));
 sg13g2_xnor2_1 _5655_ (.Y(_2115_),
    .A(net48),
    .B(_1576_));
 sg13g2_xnor2_1 _5656_ (.Y(_2116_),
    .A(_1024_),
    .B(_2115_));
 sg13g2_and2_1 _5657_ (.A(net45),
    .B(net47),
    .X(_2117_));
 sg13g2_nor3_1 _5658_ (.A(_2064_),
    .B(net39),
    .C(_2117_),
    .Y(_2118_));
 sg13g2_a21oi_1 _5659_ (.A1(_2064_),
    .A2(net39),
    .Y(_2119_),
    .B1(_2118_));
 sg13g2_or4_1 _5660_ (.A(_2035_),
    .B(_2034_),
    .C(_2116_),
    .D(_2119_),
    .X(_2120_));
 sg13g2_nor2_1 _5661_ (.A(_3049_),
    .B(_1561_),
    .Y(_2121_));
 sg13g2_xnor2_1 _5662_ (.Y(_2122_),
    .A(net32),
    .B(_1566_));
 sg13g2_mux2_1 _5663_ (.A0(_2121_),
    .A1(_2074_),
    .S(_2122_),
    .X(_2123_));
 sg13g2_xnor2_1 _5664_ (.Y(_2124_),
    .A(net27),
    .B(net163));
 sg13g2_nor3_1 _5665_ (.A(net33),
    .B(_2122_),
    .C(_2124_),
    .Y(_2125_));
 sg13g2_a21oi_1 _5666_ (.A1(net33),
    .A2(_2123_),
    .Y(_2126_),
    .B1(_2125_));
 sg13g2_xnor2_1 _5667_ (.Y(_2127_),
    .A(_2023_),
    .B(_1988_));
 sg13g2_nor2_1 _5668_ (.A(_1055_),
    .B(_1913_),
    .Y(_2128_));
 sg13g2_xnor2_1 _5669_ (.Y(_2129_),
    .A(_1921_),
    .B(_1906_));
 sg13g2_nor2_1 _5670_ (.A(_1015_),
    .B(_1948_),
    .Y(_2130_));
 sg13g2_a22oi_1 _5671_ (.Y(_2131_),
    .B1(_2129_),
    .B2(_2130_),
    .A2(_2128_),
    .A1(_1948_));
 sg13g2_nor4_1 _5672_ (.A(_2120_),
    .B(_2126_),
    .C(_2127_),
    .D(_2131_),
    .Y(_2132_));
 sg13g2_and2_1 _5673_ (.A(_0998_),
    .B(net22),
    .X(_2133_));
 sg13g2_o21ai_1 _5674_ (.B1(_2133_),
    .Y(_2134_),
    .A1(net32),
    .A2(_2085_));
 sg13g2_o21ai_1 _5675_ (.B1(_2134_),
    .Y(_2135_),
    .A1(_0998_),
    .A2(net22));
 sg13g2_nor2b_1 _5676_ (.A(_1985_),
    .B_N(_2121_),
    .Y(_2136_));
 sg13g2_nor3_1 _5677_ (.A(net33),
    .B(_2074_),
    .C(_2136_),
    .Y(_2137_));
 sg13g2_a21o_1 _5678_ (.A2(_2124_),
    .A1(net33),
    .B1(_2137_),
    .X(_2138_));
 sg13g2_or2_1 _5679_ (.X(_2139_),
    .B(net45),
    .A(net68));
 sg13g2_xnor2_1 _5680_ (.Y(_2140_),
    .A(_2139_),
    .B(_1935_));
 sg13g2_nand2_1 _5681_ (.Y(_2141_),
    .A(_0998_),
    .B(_1033_));
 sg13g2_a21oi_1 _5682_ (.A1(_1913_),
    .A2(_2140_),
    .Y(_2142_),
    .B1(_2141_));
 sg13g2_a21oi_1 _5683_ (.A1(_1968_),
    .A2(_2138_),
    .Y(_2143_),
    .B1(_2142_));
 sg13g2_nand2_1 _5684_ (.Y(_2144_),
    .A(_2018_),
    .B(_1028_));
 sg13g2_a22oi_1 _5685_ (.Y(_2145_),
    .B1(_2144_),
    .B2(_1908_),
    .A2(_2141_),
    .A1(_1958_));
 sg13g2_nor2_1 _5686_ (.A(_1949_),
    .B(_1948_),
    .Y(_2146_));
 sg13g2_nor4_1 _5687_ (.A(_2035_),
    .B(_2034_),
    .C(_1966_),
    .D(_2146_),
    .Y(_2147_));
 sg13g2_and4_1 _5688_ (.A(_2135_),
    .B(_2143_),
    .C(_2145_),
    .D(_2147_),
    .X(_2148_));
 sg13g2_nor4_1 _5689_ (.A(_2047_),
    .B(_2114_),
    .C(_2132_),
    .D(_2148_),
    .Y(_2149_));
 sg13g2_a21o_1 _5690_ (.A2(_2048_),
    .A1(_1787_),
    .B1(_2149_),
    .X(_2150_));
 sg13g2_or2_1 _5691_ (.X(_2151_),
    .B(_1856_),
    .A(_1704_));
 sg13g2_o21ai_1 _5692_ (.B1(_2151_),
    .Y(_2152_),
    .A1(net38),
    .A2(_1707_));
 sg13g2_a22oi_1 _5693_ (.Y(_2153_),
    .B1(_1820_),
    .B2(_2152_),
    .A2(_1708_),
    .A1(_1096_));
 sg13g2_nor2_1 _5694_ (.A(_1831_),
    .B(_1828_),
    .Y(_2154_));
 sg13g2_nor3_1 _5695_ (.A(_2887_),
    .B(_1717_),
    .C(_2154_),
    .Y(_2155_));
 sg13g2_nor3_1 _5696_ (.A(_2767_),
    .B(_1633_),
    .C(_1727_),
    .Y(_2156_));
 sg13g2_nor3_1 _5697_ (.A(_2892_),
    .B(net159),
    .C(_1717_),
    .Y(_2157_));
 sg13g2_o21ai_1 _5698_ (.B1(_2887_),
    .Y(_2158_),
    .A1(_2156_),
    .A2(_2157_));
 sg13g2_nor2b_1 _5699_ (.A(_2155_),
    .B_N(_2158_),
    .Y(_2159_));
 sg13g2_nor3_1 _5700_ (.A(_1772_),
    .B(_1775_),
    .C(_1776_),
    .Y(_2160_));
 sg13g2_o21ai_1 _5701_ (.B1(_1721_),
    .Y(_2161_),
    .A1(_1096_),
    .A2(_1132_));
 sg13g2_nand4_1 _5702_ (.B(_1840_),
    .C(_2160_),
    .A(_1839_),
    .Y(_2162_),
    .D(_2161_));
 sg13g2_nor2_1 _5703_ (.A(net69),
    .B(_1126_),
    .Y(_2163_));
 sg13g2_xnor2_1 _5704_ (.Y(_2164_),
    .A(_1750_),
    .B(_2163_));
 sg13g2_nor4_1 _5705_ (.A(_2153_),
    .B(_2159_),
    .C(_2162_),
    .D(_2164_),
    .Y(_2165_));
 sg13g2_nand2_1 _5706_ (.Y(_2166_),
    .A(_1747_),
    .B(_1702_));
 sg13g2_xnor2_1 _5707_ (.Y(_2167_),
    .A(net54),
    .B(_1702_));
 sg13g2_nand3_1 _5708_ (.B(net24),
    .C(_2167_),
    .A(_1136_),
    .Y(_2168_));
 sg13g2_o21ai_1 _5709_ (.B1(_2168_),
    .Y(_2169_),
    .A1(_1136_),
    .A2(_2166_));
 sg13g2_nand3_1 _5710_ (.B(_1714_),
    .C(_2169_),
    .A(_1122_),
    .Y(_2170_));
 sg13g2_nand3_1 _5711_ (.B(_1751_),
    .C(_1702_),
    .A(_1114_),
    .Y(_2171_));
 sg13g2_inv_1 _5712_ (.Y(_2172_),
    .A(_1639_));
 sg13g2_nand3_1 _5713_ (.B(_1105_),
    .C(_1700_),
    .A(net110),
    .Y(_2173_));
 sg13g2_xnor2_1 _5714_ (.Y(_2174_),
    .A(net115),
    .B(_1091_));
 sg13g2_nor3_1 _5715_ (.A(_2754_),
    .B(net110),
    .C(_1091_),
    .Y(_2175_));
 sg13g2_a21oi_1 _5716_ (.A1(_2754_),
    .A2(_2174_),
    .Y(_2176_),
    .B1(_2175_));
 sg13g2_nand2b_1 _5717_ (.Y(_2177_),
    .B(_1706_),
    .A_N(_2176_));
 sg13g2_nand2_1 _5718_ (.Y(_2178_),
    .A(_1105_),
    .B(_1886_));
 sg13g2_xnor2_1 _5719_ (.Y(_2179_),
    .A(_1750_),
    .B(_2178_));
 sg13g2_xnor2_1 _5720_ (.Y(_2180_),
    .A(_3026_),
    .B(_2154_));
 sg13g2_nand4_1 _5721_ (.B(_2160_),
    .C(_2179_),
    .A(_1761_),
    .Y(_2181_),
    .D(_2180_));
 sg13g2_a221oi_1 _5722_ (.B2(_2177_),
    .C1(_2181_),
    .B1(_2173_),
    .A1(_2170_),
    .Y(_2182_),
    .A2(_2171_));
 sg13g2_inv_1 _5723_ (.Y(_2183_),
    .A(_2045_));
 sg13g2_nand3_1 _5724_ (.B(_2183_),
    .C(_1979_),
    .A(_1946_),
    .Y(_2184_));
 sg13g2_o21ai_1 _5725_ (.B1(_2184_),
    .Y(_2185_),
    .A1(_2165_),
    .A2(_2182_));
 sg13g2_nand2b_1 _5726_ (.Y(_2186_),
    .B(_1537_),
    .A_N(\Pong.datapath.vga.Column_Counter.Q[9] ));
 sg13g2_or2_1 _5727_ (.X(_2187_),
    .B(_2186_),
    .A(_1677_));
 sg13g2_nor2b_1 _5728_ (.A(_1532_),
    .B_N(_1531_),
    .Y(_2188_));
 sg13g2_nand2_1 _5729_ (.Y(_2189_),
    .A(_1685_),
    .B(_2188_));
 sg13g2_nor2_1 _5730_ (.A(_2187_),
    .B(_2189_),
    .Y(_2190_));
 sg13g2_nand2_1 _5731_ (.Y(_2191_),
    .A(_1499_),
    .B(net170));
 sg13g2_nand2b_1 _5732_ (.Y(_2192_),
    .B(_2191_),
    .A_N(_1504_));
 sg13g2_nand2b_1 _5733_ (.Y(_2193_),
    .B(_1925_),
    .A_N(_1532_));
 sg13g2_nand4_1 _5734_ (.B(_1538_),
    .C(_1544_),
    .A(net123),
    .Y(_2194_),
    .D(_2193_));
 sg13g2_nor2b_1 _5735_ (.A(_1527_),
    .B_N(_1529_),
    .Y(_2195_));
 sg13g2_and2_1 _5736_ (.A(_1531_),
    .B(net166),
    .X(_2196_));
 sg13g2_a22oi_1 _5737_ (.Y(_2197_),
    .B1(_2196_),
    .B2(_2193_),
    .A2(_2188_),
    .A1(_2195_));
 sg13g2_nor2_1 _5738_ (.A(_1527_),
    .B(_1529_),
    .Y(_2198_));
 sg13g2_nor2_1 _5739_ (.A(_1534_),
    .B(_2198_),
    .Y(_2199_));
 sg13g2_a21o_1 _5740_ (.A2(_1544_),
    .A1(_1537_),
    .B1(net166),
    .X(_2200_));
 sg13g2_or3_1 _5741_ (.A(_1685_),
    .B(_1677_),
    .C(_2186_),
    .X(_2201_));
 sg13g2_a221oi_1 _5742_ (.B2(_2200_),
    .C1(_2201_),
    .B1(_2199_),
    .A1(_2194_),
    .Y(_2202_),
    .A2(_2197_));
 sg13g2_inv_1 _5743_ (.Y(_2203_),
    .A(_2202_));
 sg13g2_a21oi_1 _5744_ (.A1(net167),
    .A2(_2192_),
    .Y(_2204_),
    .B1(_2203_));
 sg13g2_nor2_1 _5745_ (.A(net128),
    .B(_1499_),
    .Y(_2205_));
 sg13g2_inv_1 _5746_ (.Y(_2206_),
    .A(_1508_));
 sg13g2_o21ai_1 _5747_ (.B1(_2206_),
    .Y(_2207_),
    .A1(net170),
    .A2(_2205_));
 sg13g2_nand2_1 _5748_ (.Y(_2208_),
    .A(_1512_),
    .B(_2207_));
 sg13g2_a22oi_1 _5749_ (.Y(_2209_),
    .B1(_2203_),
    .B2(_2208_),
    .A2(_1171_),
    .A1(net128));
 sg13g2_o21ai_1 _5750_ (.B1(_2209_),
    .Y(_2210_),
    .A1(_2190_),
    .A2(_2204_));
 sg13g2_nor3_1 _5751_ (.A(net127),
    .B(net162),
    .C(_1686_),
    .Y(_2211_));
 sg13g2_o21ai_1 _5752_ (.B1(_2018_),
    .Y(_2212_),
    .A1(_1560_),
    .A2(_1530_));
 sg13g2_nor2_1 _5753_ (.A(_1544_),
    .B(_2186_),
    .Y(_2213_));
 sg13g2_and3_1 _5754_ (.X(_2214_),
    .A(_2211_),
    .B(_2212_),
    .C(_2213_));
 sg13g2_nor2_1 _5755_ (.A(net172),
    .B(_1176_),
    .Y(_2215_));
 sg13g2_inv_1 _5756_ (.Y(_2216_),
    .A(net129));
 sg13g2_o21ai_1 _5757_ (.B1(_2216_),
    .Y(_2217_),
    .A1(net171),
    .A2(_2215_));
 sg13g2_and3_1 _5758_ (.X(_2218_),
    .A(_1492_),
    .B(_2214_),
    .C(_2217_));
 sg13g2_nand2_1 _5759_ (.Y(_2219_),
    .A(_1531_),
    .B(_1523_));
 sg13g2_nor2_1 _5760_ (.A(_1532_),
    .B(net162),
    .Y(_2220_));
 sg13g2_a22oi_1 _5761_ (.Y(_2221_),
    .B1(_2220_),
    .B2(_2198_),
    .A2(_2219_),
    .A1(_1525_));
 sg13g2_inv_1 _5762_ (.Y(_2222_),
    .A(_1925_));
 sg13g2_a21oi_1 _5763_ (.A1(net125),
    .A2(_2222_),
    .Y(_2223_),
    .B1(net123));
 sg13g2_nor2_1 _5764_ (.A(_1685_),
    .B(_2223_),
    .Y(_2224_));
 sg13g2_o21ai_1 _5765_ (.B1(net124),
    .Y(_2225_),
    .A1(_1570_),
    .A2(_2224_));
 sg13g2_inv_1 _5766_ (.Y(_2226_),
    .A(_1526_));
 sg13g2_inv_1 _5767_ (.Y(_2227_),
    .A(net125));
 sg13g2_nor2_1 _5768_ (.A(net123),
    .B(_2227_),
    .Y(_2228_));
 sg13g2_nand4_1 _5769_ (.B(_2195_),
    .C(_2213_),
    .A(_2226_),
    .Y(_2229_),
    .D(_2228_));
 sg13g2_a221oi_1 _5770_ (.B2(_2229_),
    .C1(_2200_),
    .B1(_2225_),
    .A1(net124),
    .Y(_2230_),
    .A2(_2221_));
 sg13g2_or2_1 _5771_ (.X(_2231_),
    .B(net171),
    .A(net129));
 sg13g2_nor2b_1 _5772_ (.A(net169),
    .B_N(net171),
    .Y(_2232_));
 sg13g2_o21ai_1 _5773_ (.B1(net129),
    .Y(_2233_),
    .A1(_1487_),
    .A2(_2232_));
 sg13g2_nor2_1 _5774_ (.A(_2214_),
    .B(_2233_),
    .Y(_2234_));
 sg13g2_a21oi_1 _5775_ (.A1(net172),
    .A2(_2231_),
    .Y(_2235_),
    .B1(_2234_));
 sg13g2_o21ai_1 _5776_ (.B1(_2235_),
    .Y(_2236_),
    .A1(_2218_),
    .A2(_2230_));
 sg13g2_nor2_1 _5777_ (.A(net160),
    .B(net116),
    .Y(_2237_));
 sg13g2_nand3_1 _5778_ (.B(net119),
    .C(net121),
    .A(net117),
    .Y(_2238_));
 sg13g2_a21oi_1 _5779_ (.A1(_2237_),
    .A2(_2238_),
    .Y(_2239_),
    .B1(_1668_));
 sg13g2_nor3_1 _5780_ (.A(_1610_),
    .B(_1601_),
    .C(_1672_),
    .Y(_2240_));
 sg13g2_nor2_1 _5781_ (.A(_1602_),
    .B(_1692_),
    .Y(_2241_));
 sg13g2_nand2_1 _5782_ (.Y(_2242_),
    .A(_2240_),
    .B(_2241_));
 sg13g2_nor2b_1 _5783_ (.A(_1596_),
    .B_N(_1592_),
    .Y(_2243_));
 sg13g2_nor2_1 _5784_ (.A(net111),
    .B(_2243_),
    .Y(_2244_));
 sg13g2_nor2_1 _5785_ (.A(_1610_),
    .B(net160),
    .Y(_2245_));
 sg13g2_nand2_1 _5786_ (.Y(_2246_),
    .A(net114),
    .B(_2245_));
 sg13g2_o21ai_1 _5787_ (.B1(_2246_),
    .Y(_2247_),
    .A1(_2242_),
    .A2(_2244_));
 sg13g2_nand2_1 _5788_ (.Y(_2248_),
    .A(_2239_),
    .B(_2247_));
 sg13g2_a21oi_1 _5789_ (.A1(_2210_),
    .A2(_2236_),
    .Y(_2249_),
    .B1(_2248_));
 sg13g2_a21oi_1 _5790_ (.A1(net119),
    .A2(_2244_),
    .Y(_2250_),
    .B1(net117));
 sg13g2_and2_1 _5791_ (.A(_1877_),
    .B(_2241_),
    .X(_2251_));
 sg13g2_nor2b_1 _5792_ (.A(_2251_),
    .B_N(_2240_),
    .Y(_2252_));
 sg13g2_o21ai_1 _5793_ (.B1(_2252_),
    .Y(_2253_),
    .A1(_1647_),
    .A2(_2250_));
 sg13g2_nor2_1 _5794_ (.A(net128),
    .B(_2191_),
    .Y(_2254_));
 sg13g2_nor2_1 _5795_ (.A(net129),
    .B(net169),
    .Y(_2255_));
 sg13g2_o21ai_1 _5796_ (.B1(_2231_),
    .Y(_2256_),
    .A1(net172),
    .A2(_2255_));
 sg13g2_a21oi_1 _5797_ (.A1(_1499_),
    .A2(_2190_),
    .Y(_2257_),
    .B1(_2202_));
 sg13g2_a21oi_1 _5798_ (.A1(_2206_),
    .A2(_1499_),
    .Y(_2258_),
    .B1(net128));
 sg13g2_a21oi_1 _5799_ (.A1(_2202_),
    .A2(_2258_),
    .Y(_2259_),
    .B1(_1163_));
 sg13g2_nor2_1 _5800_ (.A(_2257_),
    .B(_2259_),
    .Y(_2260_));
 sg13g2_a221oi_1 _5801_ (.B2(_2230_),
    .C1(_2260_),
    .B1(_2256_),
    .A1(_2190_),
    .Y(_2261_),
    .A2(_2254_));
 sg13g2_nor2_1 _5802_ (.A(_2253_),
    .B(_2261_),
    .Y(_2262_));
 sg13g2_and2_1 _5803_ (.A(_2114_),
    .B(_1904_),
    .X(_2263_));
 sg13g2_nor3_1 _5804_ (.A(net123),
    .B(net125),
    .C(net127),
    .Y(_2264_));
 sg13g2_nor4_2 _5805_ (.A(_1544_),
    .B(_2186_),
    .C(_2221_),
    .Y(_2265_),
    .D(_2264_));
 sg13g2_a21oi_1 _5806_ (.A1(net129),
    .A2(net169),
    .Y(_2266_),
    .B1(_1157_));
 sg13g2_and2_1 _5807_ (.A(net172),
    .B(net171),
    .X(_2267_));
 sg13g2_buf_1 _5808_ (.A(_2267_),
    .X(_2268_));
 sg13g2_or3_1 _5809_ (.A(_1156_),
    .B(_2215_),
    .C(_2268_),
    .X(_2269_));
 sg13g2_o21ai_1 _5810_ (.B1(_2269_),
    .Y(_2270_),
    .A1(net172),
    .A2(_2266_));
 sg13g2_and4_1 _5811_ (.A(_1560_),
    .B(net125),
    .C(_1523_),
    .D(_1683_),
    .X(_2271_));
 sg13g2_nor2_1 _5812_ (.A(net123),
    .B(net127),
    .Y(_2272_));
 sg13g2_nor3_2 _5813_ (.A(_2187_),
    .B(_2271_),
    .C(_2272_),
    .Y(_2273_));
 sg13g2_a21oi_1 _5814_ (.A1(net167),
    .A2(_1161_),
    .Y(_2274_),
    .B1(net170));
 sg13g2_and2_1 _5815_ (.A(_1160_),
    .B(_1162_),
    .X(_2275_));
 sg13g2_or3_1 _5816_ (.A(net167),
    .B(_2205_),
    .C(_2275_),
    .X(_2276_));
 sg13g2_o21ai_1 _5817_ (.B1(_2276_),
    .Y(_2277_),
    .A1(net128),
    .A2(_2274_));
 sg13g2_a22oi_1 _5818_ (.Y(_2278_),
    .B1(_2273_),
    .B2(_2277_),
    .A2(_2270_),
    .A1(_2265_));
 sg13g2_o21ai_1 _5819_ (.B1(net116),
    .Y(_2279_),
    .A1(_1692_),
    .A2(_2244_));
 sg13g2_nand4_1 _5820_ (.B(_2239_),
    .C(_2245_),
    .A(net114),
    .Y(_2280_),
    .D(_2279_));
 sg13g2_or2_1 _5821_ (.X(_2281_),
    .B(_2280_),
    .A(_2278_));
 sg13g2_nor2b_1 _5822_ (.A(_1157_),
    .B_N(_1156_),
    .Y(_2282_));
 sg13g2_nor3_1 _5823_ (.A(net169),
    .B(_2268_),
    .C(_2282_),
    .Y(_2283_));
 sg13g2_and2_1 _5824_ (.A(_2214_),
    .B(_2283_),
    .X(_2284_));
 sg13g2_nand2b_1 _5825_ (.Y(_2285_),
    .B(_2284_),
    .A_N(_2253_));
 sg13g2_o21ai_1 _5826_ (.B1(net119),
    .Y(_2286_),
    .A1(net121),
    .A2(net122));
 sg13g2_nor3_1 _5827_ (.A(net160),
    .B(_1602_),
    .C(net117),
    .Y(_2287_));
 sg13g2_a221oi_1 _5828_ (.B2(_2287_),
    .C1(_1668_),
    .B1(_2286_),
    .A1(_1656_),
    .Y(_2288_),
    .A2(_1690_));
 sg13g2_or4_1 _5829_ (.A(_2227_),
    .B(_1610_),
    .C(_1683_),
    .D(_2288_),
    .X(_2289_));
 sg13g2_nand2_1 _5830_ (.Y(_2290_),
    .A(_1524_),
    .B(_1687_));
 sg13g2_nor3_2 _5831_ (.A(_1541_),
    .B(_1582_),
    .C(_1675_),
    .Y(_2291_));
 sg13g2_nand4_1 _5832_ (.B(_1685_),
    .C(net162),
    .A(net123),
    .Y(_2292_),
    .D(_2291_));
 sg13g2_o21ai_1 _5833_ (.B1(_2292_),
    .Y(_2293_),
    .A1(net123),
    .A2(_2290_));
 sg13g2_nand3b_1 _5834_ (.B(_2293_),
    .C(_1694_),
    .Y(_2294_),
    .A_N(_2289_));
 sg13g2_nand2b_1 _5835_ (.Y(_2295_),
    .B(_1171_),
    .A_N(net128));
 sg13g2_nand2_1 _5836_ (.Y(_2296_),
    .A(net128),
    .B(_1163_));
 sg13g2_a22oi_1 _5837_ (.Y(_2297_),
    .B1(_2295_),
    .B2(_2296_),
    .A2(_1510_),
    .A1(net167));
 sg13g2_nand2_1 _5838_ (.Y(_2298_),
    .A(_1177_),
    .B(_1492_));
 sg13g2_a221oi_1 _5839_ (.B2(net129),
    .C1(_2268_),
    .B1(_2298_),
    .A1(_1177_),
    .Y(_2299_),
    .A2(_1158_));
 sg13g2_a22oi_1 _5840_ (.Y(_2300_),
    .B1(_2299_),
    .B2(_2265_),
    .A2(_2297_),
    .A1(_2273_));
 sg13g2_nor2_1 _5841_ (.A(_2242_),
    .B(_2300_),
    .Y(_2301_));
 sg13g2_inv_2 _5842_ (.Y(_2302_),
    .A(_1598_));
 sg13g2_nand4_1 _5843_ (.B(net119),
    .C(_1597_),
    .A(_2302_),
    .Y(_2303_),
    .D(_2245_));
 sg13g2_nor4_1 _5844_ (.A(_1605_),
    .B(net161),
    .C(net114),
    .D(_1647_),
    .Y(_2304_));
 sg13g2_nor3_1 _5845_ (.A(_1690_),
    .B(net116),
    .C(_1668_),
    .Y(_2305_));
 sg13g2_nor2_1 _5846_ (.A(_2304_),
    .B(_2305_),
    .Y(_2306_));
 sg13g2_nor3_1 _5847_ (.A(_1689_),
    .B(_2303_),
    .C(_2306_),
    .Y(_2307_));
 sg13g2_nand3b_1 _5848_ (.B(_1161_),
    .C(_1508_),
    .Y(_2308_),
    .A_N(_1162_));
 sg13g2_a21oi_1 _5849_ (.A1(_2191_),
    .A2(_2308_),
    .Y(_2309_),
    .B1(net128));
 sg13g2_nor3_1 _5850_ (.A(net167),
    .B(_1504_),
    .C(_2275_),
    .Y(_2310_));
 sg13g2_o21ai_1 _5851_ (.B1(_2273_),
    .Y(_2311_),
    .A1(_2309_),
    .A2(_2310_));
 sg13g2_nor3_1 _5852_ (.A(net129),
    .B(_1487_),
    .C(_2268_),
    .Y(_2312_));
 sg13g2_a21oi_1 _5853_ (.A1(net169),
    .A2(_2282_),
    .Y(_2313_),
    .B1(_2232_));
 sg13g2_nor2_1 _5854_ (.A(net172),
    .B(_2313_),
    .Y(_2314_));
 sg13g2_o21ai_1 _5855_ (.B1(_2265_),
    .Y(_2315_),
    .A1(_2312_),
    .A2(_2314_));
 sg13g2_or2_1 _5856_ (.X(_2316_),
    .B(net121),
    .A(net119));
 sg13g2_nand4_1 _5857_ (.B(_2240_),
    .C(_2316_),
    .A(net116),
    .Y(_2317_),
    .D(_2250_));
 sg13g2_a21oi_1 _5858_ (.A1(_2311_),
    .A2(_2315_),
    .Y(_2318_),
    .B1(_2317_));
 sg13g2_nor3_1 _5859_ (.A(_2301_),
    .B(_2307_),
    .C(_2318_),
    .Y(_2319_));
 sg13g2_nand4_1 _5860_ (.B(_2285_),
    .C(_2294_),
    .A(_2281_),
    .Y(_2320_),
    .D(_2319_));
 sg13g2_nor4_1 _5861_ (.A(_2249_),
    .B(_2262_),
    .C(_2263_),
    .D(_2320_),
    .Y(_2321_));
 sg13g2_nor3_1 _5862_ (.A(_0315_),
    .B(net177),
    .C(_0347_),
    .Y(_2322_));
 sg13g2_buf_2 _5863_ (.A(_2322_),
    .X(_2323_));
 sg13g2_o21ai_1 _5864_ (.B1(_0371_),
    .Y(_2324_),
    .A1(net95),
    .A2(_2323_));
 sg13g2_xor2_1 _5865_ (.B(_2324_),
    .A(_0373_),
    .X(_2325_));
 sg13g2_nor2b_1 _5866_ (.A(_2325_),
    .B_N(net120),
    .Y(_2326_));
 sg13g2_nor3_2 _5867_ (.A(net148),
    .B(net95),
    .C(_2323_),
    .Y(_2327_));
 sg13g2_o21ai_1 _5868_ (.B1(_0361_),
    .Y(_2328_),
    .A1(_0367_),
    .A2(_2327_));
 sg13g2_or3_1 _5869_ (.A(_0361_),
    .B(_0367_),
    .C(_2327_),
    .X(_2329_));
 sg13g2_and2_1 _5870_ (.A(_2328_),
    .B(_2329_),
    .X(_2330_));
 sg13g2_o21ai_1 _5871_ (.B1(_0377_),
    .Y(_2331_),
    .A1(net95),
    .A2(_2323_));
 sg13g2_xor2_1 _5872_ (.B(_2331_),
    .A(_0062_),
    .X(_2332_));
 sg13g2_nand2b_1 _5873_ (.Y(_2333_),
    .B(net161),
    .A_N(_2332_));
 sg13g2_a21o_1 _5874_ (.A2(_2333_),
    .A1(_2330_),
    .B1(_1661_),
    .X(_2334_));
 sg13g2_or2_1 _5875_ (.X(_2335_),
    .B(_2333_),
    .A(_2330_));
 sg13g2_xnor2_1 _5876_ (.Y(_2336_),
    .A(net112),
    .B(_2325_));
 sg13g2_a21oi_1 _5877_ (.A1(_2334_),
    .A2(_2335_),
    .Y(_2337_),
    .B1(_2336_));
 sg13g2_nand3_1 _5878_ (.B(_2328_),
    .C(_2329_),
    .A(_1661_),
    .Y(_2338_));
 sg13g2_inv_1 _5879_ (.Y(_2339_),
    .A(_1606_));
 sg13g2_nand2_1 _5880_ (.Y(_2340_),
    .A(_2339_),
    .B(_2332_));
 sg13g2_nand3b_1 _5881_ (.B(_2338_),
    .C(_2340_),
    .Y(_2341_),
    .A_N(_2336_));
 sg13g2_nor2_1 _5882_ (.A(net95),
    .B(_2323_),
    .Y(_2342_));
 sg13g2_buf_2 _5883_ (.A(_2342_),
    .X(_2343_));
 sg13g2_xor2_1 _5884_ (.B(_1651_),
    .A(_0381_),
    .X(_2344_));
 sg13g2_or2_1 _5885_ (.X(_2345_),
    .B(_2344_),
    .A(net175));
 sg13g2_xnor2_1 _5886_ (.Y(_2346_),
    .A(net101),
    .B(_2344_));
 sg13g2_nand3_1 _5887_ (.B(_2343_),
    .C(_2346_),
    .A(net175),
    .Y(_2347_));
 sg13g2_o21ai_1 _5888_ (.B1(_2347_),
    .Y(_2348_),
    .A1(_2343_),
    .A2(_2345_));
 sg13g2_nand2b_1 _5889_ (.Y(_2349_),
    .B(net175),
    .A_N(_2327_));
 sg13g2_xnor2_1 _5890_ (.Y(_2350_),
    .A(_0381_),
    .B(_2349_));
 sg13g2_a22oi_1 _5891_ (.Y(_2351_),
    .B1(_2350_),
    .B2(net160),
    .A2(_2348_),
    .A1(_1644_));
 sg13g2_nor2_1 _5892_ (.A(_2341_),
    .B(_2351_),
    .Y(_2352_));
 sg13g2_a21oi_1 _5893_ (.A1(_1630_),
    .A2(_1349_),
    .Y(_2353_),
    .B1(net110));
 sg13g2_nand2_1 _5894_ (.Y(_2354_),
    .A(_2302_),
    .B(net99));
 sg13g2_nand2_1 _5895_ (.Y(_2355_),
    .A(_2323_),
    .B(_2354_));
 sg13g2_xnor2_1 _5896_ (.Y(_2356_),
    .A(_1362_),
    .B(_1340_));
 sg13g2_inv_1 _5897_ (.Y(_2357_),
    .A(_1740_));
 sg13g2_nor2_1 _5898_ (.A(_1595_),
    .B(net143),
    .Y(_2358_));
 sg13g2_o21ai_1 _5899_ (.B1(_2358_),
    .Y(_2359_),
    .A1(_1616_),
    .A2(_2357_));
 sg13g2_o21ai_1 _5900_ (.B1(net143),
    .Y(_2360_),
    .A1(_1595_),
    .A2(_1740_));
 sg13g2_xor2_1 _5901_ (.B(_1625_),
    .A(_1362_),
    .X(_2361_));
 sg13g2_a221oi_1 _5902_ (.B2(_0342_),
    .C1(_2361_),
    .B1(_2360_),
    .A1(net111),
    .Y(_2362_),
    .A2(_1402_));
 sg13g2_nand2b_1 _5903_ (.Y(_2363_),
    .B(_1592_),
    .A_N(net176));
 sg13g2_xnor2_1 _5904_ (.Y(_2364_),
    .A(_1362_),
    .B(_1625_));
 sg13g2_or2_1 _5905_ (.X(_2365_),
    .B(_1740_),
    .A(net145));
 sg13g2_nor3_1 _5906_ (.A(_2363_),
    .B(_2364_),
    .C(_2365_),
    .Y(_2366_));
 sg13g2_a221oi_1 _5907_ (.B2(_2362_),
    .C1(_2366_),
    .B1(_2359_),
    .A1(_1599_),
    .Y(_2367_),
    .A2(_2356_));
 sg13g2_a21o_1 _5908_ (.A2(_2355_),
    .A1(_2353_),
    .B1(_2367_),
    .X(_2368_));
 sg13g2_o21ai_1 _5909_ (.B1(_1639_),
    .Y(_2369_),
    .A1(_2302_),
    .A2(net99));
 sg13g2_a22oi_1 _5910_ (.Y(_2370_),
    .B1(_2354_),
    .B2(net110),
    .A2(_2369_),
    .A1(_2323_));
 sg13g2_a21o_1 _5911_ (.A2(_2370_),
    .A1(_2368_),
    .B1(net178),
    .X(_2371_));
 sg13g2_nor2_1 _5912_ (.A(_1630_),
    .B(net110),
    .Y(_2372_));
 sg13g2_nand2_1 _5913_ (.Y(_2373_),
    .A(_2367_),
    .B(_2372_));
 sg13g2_a21oi_1 _5914_ (.A1(_1349_),
    .A2(_2323_),
    .Y(_2374_),
    .B1(net117));
 sg13g2_nor2_1 _5915_ (.A(_1640_),
    .B(_2374_),
    .Y(_2375_));
 sg13g2_xnor2_1 _5916_ (.Y(_2376_),
    .A(net99),
    .B(_2323_));
 sg13g2_o21ai_1 _5917_ (.B1(_2367_),
    .Y(_2377_),
    .A1(_2302_),
    .A2(_2376_));
 sg13g2_a22oi_1 _5918_ (.Y(_2378_),
    .B1(_2375_),
    .B2(_2377_),
    .A2(_2373_),
    .A1(_2343_));
 sg13g2_xnor2_1 _5919_ (.Y(_2379_),
    .A(net113),
    .B(_2343_));
 sg13g2_nand4_1 _5920_ (.B(_0313_),
    .C(net113),
    .A(net175),
    .Y(_2380_),
    .D(_2343_));
 sg13g2_o21ai_1 _5921_ (.B1(_2380_),
    .Y(_2381_),
    .A1(net175),
    .A2(_2379_));
 sg13g2_nand2b_1 _5922_ (.Y(_2382_),
    .B(_2381_),
    .A_N(_2344_));
 sg13g2_nand3_1 _5923_ (.B(net113),
    .C(_2343_),
    .A(net101),
    .Y(_2383_));
 sg13g2_o21ai_1 _5924_ (.B1(_2383_),
    .Y(_2384_),
    .A1(net113),
    .A2(_2343_));
 sg13g2_nand3_1 _5925_ (.B(_2344_),
    .C(_2384_),
    .A(net175),
    .Y(_2385_));
 sg13g2_a221oi_1 _5926_ (.B2(_2385_),
    .C1(_2341_),
    .B1(_2382_),
    .A1(_2371_),
    .Y(_2386_),
    .A2(_2378_));
 sg13g2_or4_1 _5927_ (.A(_2326_),
    .B(_2337_),
    .C(_2352_),
    .D(_2386_),
    .X(_2387_));
 sg13g2_nand4_1 _5928_ (.B(_0400_),
    .C(net142),
    .A(net141),
    .Y(_2388_),
    .D(net148));
 sg13g2_a21oi_1 _5929_ (.A1(net100),
    .A2(_1376_),
    .Y(_2389_),
    .B1(_2388_));
 sg13g2_nand4_1 _5930_ (.B(net99),
    .C(_0333_),
    .A(_1335_),
    .Y(_2390_),
    .D(_1386_));
 sg13g2_mux2_1 _5931_ (.A0(_2389_),
    .A1(_2390_),
    .S(net174),
    .X(_2391_));
 sg13g2_nand2b_1 _5932_ (.Y(_2392_),
    .B(_1610_),
    .A_N(_2391_));
 sg13g2_and3_1 _5933_ (.X(_2393_),
    .A(_0316_),
    .B(_0326_),
    .C(net176));
 sg13g2_buf_1 _5934_ (.A(_2393_),
    .X(_2394_));
 sg13g2_nand2_1 _5935_ (.Y(_2395_),
    .A(_1349_),
    .B(_2394_));
 sg13g2_nor2b_1 _5936_ (.A(net178),
    .B_N(_0332_),
    .Y(_2396_));
 sg13g2_and2_1 _5937_ (.A(net141),
    .B(_2396_),
    .X(_2397_));
 sg13g2_nor2_1 _5938_ (.A(_0399_),
    .B(_1359_),
    .Y(_2398_));
 sg13g2_o21ai_1 _5939_ (.B1(_2396_),
    .Y(_2399_),
    .A1(net146),
    .A2(_1376_));
 sg13g2_buf_2 _5940_ (.A(_2399_),
    .X(_2400_));
 sg13g2_and2_1 _5941_ (.A(_0399_),
    .B(_1359_),
    .X(_2401_));
 sg13g2_a221oi_1 _5942_ (.B2(_2400_),
    .C1(_2401_),
    .B1(_2398_),
    .A1(_2395_),
    .Y(_2402_),
    .A2(_2397_));
 sg13g2_nand2_1 _5943_ (.Y(_2403_),
    .A(_1605_),
    .B(_2402_));
 sg13g2_nand2_1 _5944_ (.Y(_2404_),
    .A(_2392_),
    .B(_2403_));
 sg13g2_xnor2_1 _5945_ (.Y(_2405_),
    .A(net142),
    .B(_1651_));
 sg13g2_nand2_1 _5946_ (.Y(_2406_),
    .A(net100),
    .B(_1376_));
 sg13g2_nand4_1 _5947_ (.B(_2400_),
    .C(_2405_),
    .A(net101),
    .Y(_2407_),
    .D(_2406_));
 sg13g2_nor2_1 _5948_ (.A(net101),
    .B(_2405_),
    .Y(_2408_));
 sg13g2_nand2b_1 _5949_ (.Y(_2409_),
    .B(_2408_),
    .A_N(_2406_));
 sg13g2_a21o_1 _5950_ (.A2(_2409_),
    .A1(_2407_),
    .B1(net113),
    .X(_2410_));
 sg13g2_and3_1 _5951_ (.X(_2411_),
    .A(net142),
    .B(net101),
    .C(_2400_));
 sg13g2_a21oi_1 _5952_ (.A1(net101),
    .A2(_2400_),
    .Y(_2412_),
    .B1(net142));
 sg13g2_o21ai_1 _5953_ (.B1(_1607_),
    .Y(_2413_),
    .A1(_2411_),
    .A2(_2412_));
 sg13g2_inv_1 _5954_ (.Y(_2414_),
    .A(_1655_));
 sg13g2_a21oi_1 _5955_ (.A1(net100),
    .A2(_1376_),
    .Y(_2415_),
    .B1(_0404_));
 sg13g2_xnor2_1 _5956_ (.Y(_2416_),
    .A(net140),
    .B(_2415_));
 sg13g2_nand2_1 _5957_ (.Y(_2417_),
    .A(_2414_),
    .B(_2416_));
 sg13g2_nand3_1 _5958_ (.B(_0440_),
    .C(_2396_),
    .A(net101),
    .Y(_2418_));
 sg13g2_or3_1 _5959_ (.A(net113),
    .B(_2405_),
    .C(_2418_),
    .X(_2419_));
 sg13g2_nand4_1 _5960_ (.B(_2413_),
    .C(_2417_),
    .A(_2410_),
    .Y(_2420_),
    .D(_2419_));
 sg13g2_xnor2_1 _5961_ (.Y(_2421_),
    .A(_1362_),
    .B(_1369_));
 sg13g2_and2_1 _5962_ (.A(net145),
    .B(_1740_),
    .X(_2422_));
 sg13g2_o21ai_1 _5963_ (.B1(_2365_),
    .Y(_2423_),
    .A1(_2363_),
    .A2(_2422_));
 sg13g2_nor2_1 _5964_ (.A(_1369_),
    .B(_2364_),
    .Y(_2424_));
 sg13g2_a221oi_1 _5965_ (.B2(_2364_),
    .C1(_2424_),
    .B1(_2423_),
    .A1(_1599_),
    .Y(_2425_),
    .A2(_2421_));
 sg13g2_xnor2_1 _5966_ (.Y(_2426_),
    .A(net99),
    .B(_2394_));
 sg13g2_a21o_1 _5967_ (.A2(_2425_),
    .A1(net159),
    .B1(_2426_),
    .X(_2427_));
 sg13g2_or2_1 _5968_ (.X(_2428_),
    .B(_2425_),
    .A(net159));
 sg13g2_o21ai_1 _5969_ (.B1(_0333_),
    .Y(_2429_),
    .A1(net146),
    .A2(_1376_));
 sg13g2_xor2_1 _5970_ (.B(_2429_),
    .A(_0322_),
    .X(_2430_));
 sg13g2_nand2b_1 _5971_ (.Y(_2431_),
    .B(net115),
    .A_N(_2430_));
 sg13g2_nand2_1 _5972_ (.Y(_2432_),
    .A(net110),
    .B(_2430_));
 sg13g2_xnor2_1 _5973_ (.Y(_2433_),
    .A(_2400_),
    .B(_2405_));
 sg13g2_o21ai_1 _5974_ (.B1(_1645_),
    .Y(_2434_),
    .A1(_0414_),
    .A2(_2394_));
 sg13g2_nand3b_1 _5975_ (.B(net100),
    .C(_1376_),
    .Y(_2435_),
    .A_N(_1645_));
 sg13g2_a21oi_1 _5976_ (.A1(_2434_),
    .A2(_2435_),
    .Y(_2436_),
    .B1(_0313_));
 sg13g2_and2_1 _5977_ (.A(_2434_),
    .B(_2435_),
    .X(_2437_));
 sg13g2_a22oi_1 _5978_ (.Y(_2438_),
    .B1(_2408_),
    .B2(_2437_),
    .A2(_2436_),
    .A1(_2433_));
 sg13g2_a221oi_1 _5979_ (.B2(_2432_),
    .C1(_2438_),
    .B1(_2431_),
    .A1(_2427_),
    .Y(_2439_),
    .A2(_2428_));
 sg13g2_nor3_1 _5980_ (.A(_1647_),
    .B(_2438_),
    .C(_2430_),
    .Y(_2440_));
 sg13g2_or4_1 _5981_ (.A(_2404_),
    .B(_2420_),
    .C(_2439_),
    .D(_2440_),
    .X(_2441_));
 sg13g2_xnor2_1 _5982_ (.Y(_2442_),
    .A(_1661_),
    .B(_2402_));
 sg13g2_o21ai_1 _5983_ (.B1(_2442_),
    .Y(_2443_),
    .A1(_2414_),
    .A2(_2416_));
 sg13g2_nand2b_1 _5984_ (.Y(_2444_),
    .B(_2443_),
    .A_N(_2404_));
 sg13g2_nand2_1 _5985_ (.Y(_2445_),
    .A(net174),
    .B(net112));
 sg13g2_or2_1 _5986_ (.X(_2446_),
    .B(net112),
    .A(\Pong.datapath.rightPaddle[9] ));
 sg13g2_o21ai_1 _5987_ (.B1(_2446_),
    .Y(_2447_),
    .A1(_2400_),
    .A2(_2445_));
 sg13g2_nand3_1 _5988_ (.B(_2396_),
    .C(_1376_),
    .A(_0403_),
    .Y(_2448_));
 sg13g2_a21oi_1 _5989_ (.A1(_1386_),
    .A2(_2448_),
    .Y(_2449_),
    .B1(net112));
 sg13g2_inv_1 _5990_ (.Y(_2450_),
    .A(net112));
 sg13g2_nor3_1 _5991_ (.A(net174),
    .B(_2450_),
    .C(_2389_),
    .Y(_2451_));
 sg13g2_a221oi_1 _5992_ (.B2(net174),
    .C1(_2451_),
    .B1(_2449_),
    .A1(_2389_),
    .Y(_2452_),
    .A2(_2447_));
 sg13g2_nand2_1 _5993_ (.Y(_2453_),
    .A(_2392_),
    .B(_2452_));
 sg13g2_xnor2_1 _5994_ (.Y(_2454_),
    .A(net110),
    .B(_2430_));
 sg13g2_xnor2_1 _5995_ (.Y(_2455_),
    .A(_1633_),
    .B(_2426_));
 sg13g2_nor2b_1 _5996_ (.A(net102),
    .B_N(net143),
    .Y(_2456_));
 sg13g2_xnor2_1 _5997_ (.Y(_2457_),
    .A(net102),
    .B(net111));
 sg13g2_nor2_1 _5998_ (.A(_2363_),
    .B(_2457_),
    .Y(_2458_));
 sg13g2_a21oi_1 _5999_ (.A1(_2456_),
    .A2(_1810_),
    .Y(_2459_),
    .B1(_2458_));
 sg13g2_nand2_1 _6000_ (.Y(_2460_),
    .A(_1742_),
    .B(_2424_));
 sg13g2_o21ai_1 _6001_ (.B1(_2460_),
    .Y(_2461_),
    .A1(_2361_),
    .A2(_2459_));
 sg13g2_nand4_1 _6002_ (.B(_2417_),
    .C(_2455_),
    .A(_2454_),
    .Y(_2462_),
    .D(_2461_));
 sg13g2_or4_1 _6003_ (.A(_2438_),
    .B(_2452_),
    .C(_2443_),
    .D(_2462_),
    .X(_2463_));
 sg13g2_nand4_1 _6004_ (.B(_2444_),
    .C(_2453_),
    .A(_2441_),
    .Y(_2464_),
    .D(_2463_));
 sg13g2_inv_1 _6005_ (.Y(_2465_),
    .A(_2291_));
 sg13g2_nand2_1 _6006_ (.Y(_2466_),
    .A(_2198_),
    .B(_2188_));
 sg13g2_nand2_1 _6007_ (.Y(_2467_),
    .A(_1683_),
    .B(_2228_));
 sg13g2_o21ai_1 _6008_ (.B1(_1548_),
    .Y(_2468_),
    .A1(_1561_),
    .A2(_1526_));
 sg13g2_a22oi_1 _6009_ (.Y(_2469_),
    .B1(_2291_),
    .B2(_2468_),
    .A2(_1674_),
    .A1(_1539_));
 sg13g2_mux2_1 _6010_ (.A0(_2466_),
    .A1(_2467_),
    .S(_2469_),
    .X(_2470_));
 sg13g2_nor4_1 _6011_ (.A(net174),
    .B(net141),
    .C(_0367_),
    .D(_2327_),
    .Y(_2471_));
 sg13g2_nor4_1 _6012_ (.A(_1526_),
    .B(_2465_),
    .C(_2470_),
    .D(_2471_),
    .Y(_2472_));
 sg13g2_nand3_1 _6013_ (.B(_2464_),
    .C(_2472_),
    .A(_2387_),
    .Y(_2473_));
 sg13g2_nand4_1 _6014_ (.B(_2185_),
    .C(_2321_),
    .A(_2150_),
    .Y(_2474_),
    .D(_2473_));
 sg13g2_xnor2_1 _6015_ (.Y(_2475_),
    .A(net153),
    .B(_1651_));
 sg13g2_inv_1 _6016_ (.Y(_2476_),
    .A(_2475_));
 sg13g2_nand3b_1 _6017_ (.B(_2903_),
    .C(net184),
    .Y(_2477_),
    .A_N(_0083_));
 sg13g2_buf_1 _6018_ (.A(_2477_),
    .X(_2478_));
 sg13g2_nand2_1 _6019_ (.Y(_2479_),
    .A(net104),
    .B(_2478_));
 sg13g2_xor2_1 _6020_ (.B(_2479_),
    .A(_1645_),
    .X(_2480_));
 sg13g2_nor2b_1 _6021_ (.A(_2907_),
    .B_N(_2959_),
    .Y(_2481_));
 sg13g2_o21ai_1 _6022_ (.B1(_2481_),
    .Y(_2482_),
    .A1(net183),
    .A2(_1221_));
 sg13g2_buf_1 _6023_ (.A(_2482_),
    .X(_2483_));
 sg13g2_nor3_1 _6024_ (.A(_1193_),
    .B(_2483_),
    .C(_2480_),
    .Y(_2484_));
 sg13g2_a21o_1 _6025_ (.A2(_2480_),
    .A1(_1193_),
    .B1(_2484_),
    .X(_2485_));
 sg13g2_nand2_1 _6026_ (.Y(_2486_),
    .A(_2933_),
    .B(_2483_));
 sg13g2_nor2_1 _6027_ (.A(_2476_),
    .B(_2486_),
    .Y(_2487_));
 sg13g2_nor2b_1 _6028_ (.A(_2480_),
    .B_N(_2487_),
    .Y(_2488_));
 sg13g2_a21oi_1 _6029_ (.A1(_2476_),
    .A2(_2485_),
    .Y(_2489_),
    .B1(_2488_));
 sg13g2_o21ai_1 _6030_ (.B1(_2959_),
    .Y(_2490_),
    .A1(net151),
    .A2(_1221_));
 sg13g2_xnor2_1 _6031_ (.Y(_2491_),
    .A(_3017_),
    .B(_2490_));
 sg13g2_inv_1 _6032_ (.Y(_2492_),
    .A(_2491_));
 sg13g2_xnor2_1 _6033_ (.Y(_2493_),
    .A(_1200_),
    .B(_2478_));
 sg13g2_and2_1 _6034_ (.A(_1632_),
    .B(_2493_),
    .X(_2494_));
 sg13g2_nor2_1 _6035_ (.A(net115),
    .B(_2494_),
    .Y(_2495_));
 sg13g2_nor3_1 _6036_ (.A(net110),
    .B(_2491_),
    .C(_2494_),
    .Y(_2496_));
 sg13g2_a21o_1 _6037_ (.A2(_2495_),
    .A1(_2491_),
    .B1(_2496_),
    .X(_2497_));
 sg13g2_xnor2_1 _6038_ (.Y(_2498_),
    .A(net168),
    .B(_1625_));
 sg13g2_nor2_1 _6039_ (.A(_1234_),
    .B(_2498_),
    .Y(_2499_));
 sg13g2_xnor2_1 _6040_ (.Y(_2500_),
    .A(net168),
    .B(_1234_));
 sg13g2_nand2_1 _6041_ (.Y(_2501_),
    .A(_1593_),
    .B(_1185_));
 sg13g2_a21oi_1 _6042_ (.A1(net105),
    .A2(net111),
    .Y(_2502_),
    .B1(_2501_));
 sg13g2_a21o_1 _6043_ (.A2(_2357_),
    .A1(_2950_),
    .B1(_2502_),
    .X(_2503_));
 sg13g2_nor2_1 _6044_ (.A(_1632_),
    .B(_2493_),
    .Y(_2504_));
 sg13g2_a221oi_1 _6045_ (.B2(_2503_),
    .C1(_2504_),
    .B1(_2498_),
    .A1(_1623_),
    .Y(_2505_),
    .A2(_2500_));
 sg13g2_nand2b_1 _6046_ (.Y(_2506_),
    .B(_2505_),
    .A_N(_2499_));
 sg13g2_a22oi_1 _6047_ (.Y(_2507_),
    .B1(_2497_),
    .B2(_2506_),
    .A2(_2492_),
    .A1(_1637_));
 sg13g2_a21oi_1 _6048_ (.A1(net104),
    .A2(_2478_),
    .Y(_2508_),
    .B1(_1193_));
 sg13g2_nand2b_1 _6049_ (.Y(_2509_),
    .B(_2508_),
    .A_N(_2483_));
 sg13g2_o21ai_1 _6050_ (.B1(_2509_),
    .Y(_2510_),
    .A1(_2933_),
    .A2(_2479_));
 sg13g2_a22oi_1 _6051_ (.Y(_2511_),
    .B1(_2487_),
    .B2(_2479_),
    .A2(_2510_),
    .A1(_2476_));
 sg13g2_nor2_1 _6052_ (.A(_1646_),
    .B(_2511_),
    .Y(_2512_));
 sg13g2_a21oi_1 _6053_ (.A1(_2910_),
    .A2(_2478_),
    .Y(_2513_),
    .B1(_2913_));
 sg13g2_xnor2_1 _6054_ (.Y(_2514_),
    .A(net154),
    .B(_2513_));
 sg13g2_and2_1 _6055_ (.A(_2414_),
    .B(_2514_),
    .X(_2515_));
 sg13g2_xnor2_1 _6056_ (.Y(_2516_),
    .A(_2930_),
    .B(_2486_));
 sg13g2_nand2_1 _6057_ (.Y(_2517_),
    .A(_1243_),
    .B(_2483_));
 sg13g2_xor2_1 _6058_ (.B(_2517_),
    .A(_2895_),
    .X(_2518_));
 sg13g2_and2_1 _6059_ (.A(_2910_),
    .B(_1221_),
    .X(_2519_));
 sg13g2_nor2b_1 _6060_ (.A(_2519_),
    .B_N(_1244_),
    .Y(_2520_));
 sg13g2_xnor2_1 _6061_ (.Y(_2521_),
    .A(net181),
    .B(_2520_));
 sg13g2_a22oi_1 _6062_ (.Y(_2522_),
    .B1(_2521_),
    .B2(net120),
    .A2(_2518_),
    .A1(_1605_));
 sg13g2_o21ai_1 _6063_ (.B1(_2522_),
    .Y(_2523_),
    .A1(_1656_),
    .A2(_2516_));
 sg13g2_nor3_1 _6064_ (.A(_2512_),
    .B(_2515_),
    .C(_2523_),
    .Y(_2524_));
 sg13g2_o21ai_1 _6065_ (.B1(_2524_),
    .Y(_2525_),
    .A1(_2489_),
    .A2(_2507_));
 sg13g2_nand2b_1 _6066_ (.Y(_2526_),
    .B(net112),
    .A_N(_2519_));
 sg13g2_nor3_1 _6067_ (.A(_1610_),
    .B(net112),
    .C(_2519_),
    .Y(_2527_));
 sg13g2_o21ai_1 _6068_ (.B1(net181),
    .Y(_2528_),
    .A1(_2483_),
    .A2(_2527_));
 sg13g2_o21ai_1 _6069_ (.B1(_2528_),
    .Y(_2529_),
    .A1(net181),
    .A2(_2526_));
 sg13g2_nor2_1 _6070_ (.A(_2414_),
    .B(_2514_),
    .Y(_2530_));
 sg13g2_xnor2_1 _6071_ (.Y(_2531_),
    .A(_1661_),
    .B(_2518_));
 sg13g2_nand2b_1 _6072_ (.Y(_2532_),
    .B(_2531_),
    .A_N(_2530_));
 sg13g2_nor3_1 _6073_ (.A(_1611_),
    .B(_2924_),
    .C(net112),
    .Y(_2533_));
 sg13g2_a21oi_1 _6074_ (.A1(_2924_),
    .A2(_1667_),
    .Y(_2534_),
    .B1(_2533_));
 sg13g2_nor2_1 _6075_ (.A(_2520_),
    .B(_2534_),
    .Y(_2535_));
 sg13g2_a221oi_1 _6076_ (.B2(_2522_),
    .C1(_2535_),
    .B1(_2532_),
    .A1(_1244_),
    .Y(_2536_),
    .A2(_2529_));
 sg13g2_xnor2_1 _6077_ (.Y(_2537_),
    .A(net105),
    .B(net111));
 sg13g2_nand2b_1 _6078_ (.Y(_2538_),
    .B(_1810_),
    .A_N(_1262_));
 sg13g2_o21ai_1 _6079_ (.B1(_2538_),
    .Y(_2539_),
    .A1(_2501_),
    .A2(_2537_));
 sg13g2_a22oi_1 _6080_ (.Y(_2540_),
    .B1(_2539_),
    .B2(_2498_),
    .A2(_2499_),
    .A1(_1742_));
 sg13g2_xnor2_1 _6081_ (.Y(_2541_),
    .A(_2450_),
    .B(_2521_));
 sg13g2_or4_1 _6082_ (.A(_2515_),
    .B(_2530_),
    .C(_2540_),
    .D(_2541_),
    .X(_2542_));
 sg13g2_nand2_1 _6083_ (.Y(_2543_),
    .A(_2497_),
    .B(_2531_));
 sg13g2_or4_1 _6084_ (.A(_2489_),
    .B(_2504_),
    .C(_2542_),
    .D(_2543_),
    .X(_2544_));
 sg13g2_and2_1 _6085_ (.A(_2536_),
    .B(_2544_),
    .X(_2545_));
 sg13g2_nor3_2 _6086_ (.A(net156),
    .B(net155),
    .C(net150),
    .Y(_2546_));
 sg13g2_nor2_2 _6087_ (.A(_2986_),
    .B(_2546_),
    .Y(_2547_));
 sg13g2_xnor2_1 _6088_ (.Y(_2548_),
    .A(_0075_),
    .B(_1651_));
 sg13g2_nand2b_1 _6089_ (.Y(_2549_),
    .B(_2548_),
    .A_N(net149));
 sg13g2_nor3_2 _6090_ (.A(net152),
    .B(_2986_),
    .C(_2546_),
    .Y(_2550_));
 sg13g2_xnor2_1 _6091_ (.Y(_2551_),
    .A(_2550_),
    .B(_2548_));
 sg13g2_nand3_1 _6092_ (.B(_2547_),
    .C(_2551_),
    .A(net149),
    .Y(_2552_));
 sg13g2_o21ai_1 _6093_ (.B1(_2552_),
    .Y(_2553_),
    .A1(_2547_),
    .A2(_2549_));
 sg13g2_nand2b_1 _6094_ (.Y(_2554_),
    .B(_3001_),
    .A_N(_2547_));
 sg13g2_xor2_1 _6095_ (.B(_2554_),
    .A(_2921_),
    .X(_2555_));
 sg13g2_nand2b_1 _6096_ (.Y(_2556_),
    .B(_1611_),
    .A_N(_2555_));
 sg13g2_nor2_1 _6097_ (.A(_2993_),
    .B(_2550_),
    .Y(_2557_));
 sg13g2_xor2_1 _6098_ (.B(_2557_),
    .A(net179),
    .X(_2558_));
 sg13g2_nand2_1 _6099_ (.Y(_2559_),
    .A(_1662_),
    .B(_2558_));
 sg13g2_nor2b_1 _6100_ (.A(_2550_),
    .B_N(net149),
    .Y(_2560_));
 sg13g2_xnor2_1 _6101_ (.Y(_2561_),
    .A(_3006_),
    .B(_2560_));
 sg13g2_nor2_1 _6102_ (.A(_2997_),
    .B(_2547_),
    .Y(_2562_));
 sg13g2_xnor2_1 _6103_ (.Y(_2563_),
    .A(_0074_),
    .B(_2562_));
 sg13g2_nor2_1 _6104_ (.A(_2339_),
    .B(_2563_),
    .Y(_2564_));
 sg13g2_a21oi_1 _6105_ (.A1(_1607_),
    .A2(_2561_),
    .Y(_2565_),
    .B1(_2564_));
 sg13g2_nand3_1 _6106_ (.B(_2559_),
    .C(_2565_),
    .A(_2556_),
    .Y(_2566_));
 sg13g2_a21oi_1 _6107_ (.A1(_1644_),
    .A2(_2553_),
    .Y(_2567_),
    .B1(_2566_));
 sg13g2_xnor2_1 _6108_ (.Y(_2568_),
    .A(_1646_),
    .B(_2547_));
 sg13g2_nor2_1 _6109_ (.A(_2549_),
    .B(_2568_),
    .Y(_2569_));
 sg13g2_nand3_1 _6110_ (.B(_2551_),
    .C(_2568_),
    .A(net149),
    .Y(_2570_));
 sg13g2_nor2b_1 _6111_ (.A(_2569_),
    .B_N(_2570_),
    .Y(_2571_));
 sg13g2_a21oi_1 _6112_ (.A1(_1593_),
    .A2(_1272_),
    .Y(_2572_),
    .B1(_1213_));
 sg13g2_nand3b_1 _6113_ (.B(_2905_),
    .C(_1592_),
    .Y(_2573_),
    .A_N(net150));
 sg13g2_a21o_1 _6114_ (.A2(_2573_),
    .A1(_1262_),
    .B1(_2357_),
    .X(_2574_));
 sg13g2_o21ai_1 _6115_ (.B1(_2574_),
    .Y(_2575_),
    .A1(_1741_),
    .A2(_2572_));
 sg13g2_nand2b_1 _6116_ (.Y(_2576_),
    .B(net150),
    .A_N(_1741_));
 sg13g2_a21oi_1 _6117_ (.A1(_1263_),
    .A2(_2576_),
    .Y(_2577_),
    .B1(_1877_));
 sg13g2_or2_1 _6118_ (.X(_2578_),
    .B(_2577_),
    .A(_1599_));
 sg13g2_xnor2_1 _6119_ (.Y(_2579_),
    .A(net168),
    .B(_1272_));
 sg13g2_nor2_1 _6120_ (.A(_1599_),
    .B(_1626_),
    .Y(_2580_));
 sg13g2_nor2_1 _6121_ (.A(_2579_),
    .B(_2580_),
    .Y(_2581_));
 sg13g2_o21ai_1 _6122_ (.B1(_2581_),
    .Y(_2582_),
    .A1(_2575_),
    .A2(_2578_));
 sg13g2_nor2b_1 _6123_ (.A(_1626_),
    .B_N(_2579_),
    .Y(_2583_));
 sg13g2_o21ai_1 _6124_ (.B1(_2583_),
    .Y(_2584_),
    .A1(_2575_),
    .A2(_2577_));
 sg13g2_nand3_1 _6125_ (.B(_2582_),
    .C(_2584_),
    .A(_2372_),
    .Y(_2585_));
 sg13g2_nand2_1 _6126_ (.Y(_2586_),
    .A(_3007_),
    .B(_1272_));
 sg13g2_nor3_1 _6127_ (.A(net151),
    .B(net115),
    .C(_2586_),
    .Y(_2587_));
 sg13g2_nand2b_1 _6128_ (.Y(_2588_),
    .B(net117),
    .A_N(net133));
 sg13g2_nor2_1 _6129_ (.A(_2586_),
    .B(_2588_),
    .Y(_2589_));
 sg13g2_nand2_1 _6130_ (.Y(_2590_),
    .A(_2582_),
    .B(_2584_));
 sg13g2_o21ai_1 _6131_ (.B1(_2590_),
    .Y(_2591_),
    .A1(_2587_),
    .A2(_2589_));
 sg13g2_nor2_1 _6132_ (.A(net133),
    .B(net115),
    .Y(_2592_));
 sg13g2_nor2_1 _6133_ (.A(_2302_),
    .B(net115),
    .Y(_2593_));
 sg13g2_o21ai_1 _6134_ (.B1(_2590_),
    .Y(_2594_),
    .A1(_2592_),
    .A2(_2593_));
 sg13g2_nand3b_1 _6135_ (.B(_2590_),
    .C(_1200_),
    .Y(_2595_),
    .A_N(_2588_));
 sg13g2_nor3_1 _6136_ (.A(_2302_),
    .B(net151),
    .C(_1640_),
    .Y(_2596_));
 sg13g2_a21oi_1 _6137_ (.A1(_2546_),
    .A2(_2596_),
    .Y(_2597_),
    .B1(_2547_));
 sg13g2_o21ai_1 _6138_ (.B1(_2546_),
    .Y(_2598_),
    .A1(net104),
    .A2(_2592_));
 sg13g2_nor2_1 _6139_ (.A(net115),
    .B(_2588_),
    .Y(_2599_));
 sg13g2_a21oi_1 _6140_ (.A1(_2172_),
    .A2(net104),
    .Y(_2600_),
    .B1(_2599_));
 sg13g2_and3_1 _6141_ (.X(_2601_),
    .A(_2597_),
    .B(_2598_),
    .C(_2600_));
 sg13g2_nand4_1 _6142_ (.B(_2594_),
    .C(_2595_),
    .A(_2591_),
    .Y(_2602_),
    .D(_2601_));
 sg13g2_nand3b_1 _6143_ (.B(_2585_),
    .C(_2602_),
    .Y(_2603_),
    .A_N(_2571_));
 sg13g2_nor2_1 _6144_ (.A(_1662_),
    .B(_2558_),
    .Y(_2604_));
 sg13g2_nand3_1 _6145_ (.B(_2559_),
    .C(_2563_),
    .A(_2339_),
    .Y(_2605_));
 sg13g2_xnor2_1 _6146_ (.Y(_2606_),
    .A(_2450_),
    .B(_2555_));
 sg13g2_nand3b_1 _6147_ (.B(_2605_),
    .C(_2606_),
    .Y(_2607_),
    .A_N(_2604_));
 sg13g2_or4_1 _6148_ (.A(net181),
    .B(net185),
    .C(_2993_),
    .D(_2550_),
    .X(_2608_));
 sg13g2_nor4_1 _6149_ (.A(_1538_),
    .B(_1539_),
    .C(_1544_),
    .D(_2189_),
    .Y(_2609_));
 sg13g2_nand4_1 _6150_ (.B(_1699_),
    .C(_2608_),
    .A(_1570_),
    .Y(_2610_),
    .D(_2609_));
 sg13g2_a21o_1 _6151_ (.A2(_2607_),
    .A1(_2556_),
    .B1(_2610_),
    .X(_2611_));
 sg13g2_a221oi_1 _6152_ (.B2(_2603_),
    .C1(_2611_),
    .B1(_2567_),
    .A1(_2525_),
    .Y(_2612_),
    .A2(_2545_));
 sg13g2_a21o_1 _6153_ (.A2(_2474_),
    .A1(_1699_),
    .B1(_2612_),
    .X(\Pong.b ));
 sg13g2_inv_1 _6154_ (.Y(_2613_),
    .A(net165));
 sg13g2_nor4_1 _6155_ (.A(_1542_),
    .B(net127),
    .C(net162),
    .D(_1571_),
    .Y(_2614_));
 sg13g2_nor3_1 _6156_ (.A(_2613_),
    .B(_1675_),
    .C(_2614_),
    .Y(_2615_));
 sg13g2_o21ai_1 _6157_ (.B1(_1685_),
    .Y(_2616_),
    .A1(net124),
    .A2(_1536_));
 sg13g2_nand3_1 _6158_ (.B(net162),
    .C(_2616_),
    .A(_1542_),
    .Y(_2617_));
 sg13g2_nand2_1 _6159_ (.Y(\Pong.datapath.h_sync ),
    .A(_2615_),
    .B(_2617_));
 sg13g2_a22oi_1 _6160_ (.Y(_2618_),
    .B1(_1810_),
    .B2(_1633_),
    .A2(_2243_),
    .A1(net117));
 sg13g2_nand2_1 _6161_ (.Y(_2619_),
    .A(_2302_),
    .B(_1633_));
 sg13g2_o21ai_1 _6162_ (.B1(_2619_),
    .Y(_2620_),
    .A1(net119),
    .A2(_2618_));
 sg13g2_nor3_1 _6163_ (.A(net120),
    .B(_1690_),
    .C(net116),
    .Y(_2621_));
 sg13g2_nand3_1 _6164_ (.B(_2620_),
    .C(_2621_),
    .A(_1673_),
    .Y(\Pong.datapath.v_sync ));
 sg13g2_inv_1 _6165_ (.Y(_2622_),
    .A(_2806_));
 sg13g2_nand2b_1 _6166_ (.Y(_2623_),
    .B(\Pong.control_unit.NES_Controller_Left.state_NESController[6] ),
    .A_N(_2792_));
 sg13g2_and2_1 _6167_ (.A(_0827_),
    .B(_2623_),
    .X(_2624_));
 sg13g2_o21ai_1 _6168_ (.B1(_0123_),
    .Y(_2625_),
    .A1(_0838_),
    .A2(_2624_));
 sg13g2_nand2_1 _6169_ (.Y(_2626_),
    .A(_0122_),
    .B(_2625_));
 sg13g2_nand2_1 _6170_ (.Y(_2627_),
    .A(_0126_),
    .B(_2626_));
 sg13g2_nand2_1 _6171_ (.Y(_2628_),
    .A(_0125_),
    .B(_2627_));
 sg13g2_a21oi_1 _6172_ (.A1(_0121_),
    .A2(_2628_),
    .Y(_2629_),
    .B1(_2844_));
 sg13g2_o21ai_1 _6173_ (.B1(_2799_),
    .Y(_2630_),
    .A1(_2797_),
    .A2(_2629_));
 sg13g2_a21oi_1 _6174_ (.A1(_2622_),
    .A2(_2630_),
    .Y(net3),
    .B1(_0830_));
 sg13g2_nor2b_1 _6175_ (.A(_0822_),
    .B_N(_0119_),
    .Y(net4));
 sg13g2_inv_1 _6176_ (.Y(_2631_),
    .A(_2704_));
 sg13g2_nor2b_1 _6177_ (.A(\Pong.control_unit.NES_Controller_Right.state_NESController[11] ),
    .B_N(\Pong.control_unit.NES_Controller_Right.state_NESController[6] ),
    .Y(_2632_));
 sg13g2_nor3_1 _6178_ (.A(_2671_),
    .B(\Pong.control_unit.NES_Controller_Right.state_NESController[1] ),
    .C(_2632_),
    .Y(_2633_));
 sg13g2_o21ai_1 _6179_ (.B1(_0131_),
    .Y(_2634_),
    .A1(_0891_),
    .A2(_2633_));
 sg13g2_nand2_1 _6180_ (.Y(_2635_),
    .A(_0130_),
    .B(_2634_));
 sg13g2_nand2_1 _6181_ (.Y(_2636_),
    .A(_0134_),
    .B(_2635_));
 sg13g2_nand2_1 _6182_ (.Y(_2637_),
    .A(_0133_),
    .B(_2636_));
 sg13g2_a21oi_1 _6183_ (.A1(_0129_),
    .A2(_2637_),
    .Y(_2638_),
    .B1(\Pong.control_unit.NES_Controller_Right.state_NESController[17] ));
 sg13g2_o21ai_1 _6184_ (.B1(_2667_),
    .Y(_2639_),
    .A1(_2665_),
    .A2(_2638_));
 sg13g2_a21oi_1 _6185_ (.A1(_2631_),
    .A2(_2639_),
    .Y(net5),
    .B1(_0894_));
 sg13g2_nor2b_1 _6186_ (.A(_0878_),
    .B_N(_0538_),
    .Y(net6));
 sg13g2_buf_1 clkbuf_0_clk (.A(clk),
    .X(clknet_0_clk));
 sg13g2_tiehi \Pong.control_unit.NES_Controller_Left.state_NESController[0]$_DFF_P__197  (.L_HI(net197));
 sg13g2_buf_1 _6189_ (.A(net189),
    .X(uio_oe[0]));
 sg13g2_buf_1 _6190_ (.A(net410),
    .X(uio_oe[1]));
 sg13g2_buf_1 _6191_ (.A(net411),
    .X(uio_oe[2]));
 sg13g2_buf_1 _6192_ (.A(net190),
    .X(uio_oe[3]));
 sg13g2_buf_1 _6193_ (.A(net412),
    .X(uio_oe[4]));
 sg13g2_buf_1 _6194_ (.A(net413),
    .X(uio_oe[5]));
 sg13g2_buf_1 _6195_ (.A(net191),
    .X(uio_oe[6]));
 sg13g2_buf_1 _6196_ (.A(net192),
    .X(uio_oe[7]));
 sg13g2_buf_1 _6197_ (.A(net193),
    .X(uio_out[0]));
 sg13g2_buf_1 _6198_ (.A(net194),
    .X(uio_out[3]));
 sg13g2_buf_1 _6199_ (.A(net195),
    .X(uio_out[6]));
 sg13g2_buf_1 _6200_ (.A(net196),
    .X(uio_out[7]));
 sg13g2_buf_1 _6201_ (.A(\Pong.b ),
    .X(net7));
 sg13g2_buf_1 _6202_ (.A(\Pong.b ),
    .X(net8));
 sg13g2_buf_1 _6203_ (.A(\Pong.b ),
    .X(net9));
 sg13g2_buf_1 _6204_ (.A(\Pong.datapath.v_sync ),
    .X(net10));
 sg13g2_buf_1 _6205_ (.A(\Pong.b ),
    .X(net11));
 sg13g2_buf_1 _6206_ (.A(\Pong.b ),
    .X(net12));
 sg13g2_buf_1 _6207_ (.A(\Pong.b ),
    .X(net13));
 sg13g2_buf_1 _6208_ (.A(\Pong.datapath.h_sync ),
    .X(net14));
 sg13g2_buf_1 input1 (.A(uio_in[0]),
    .X(net1));
 sg13g2_buf_1 input2 (.A(uio_in[3]),
    .X(net2));
 sg13g2_buf_1 output3 (.A(net3),
    .X(uio_out[1]));
 sg13g2_buf_1 output4 (.A(net4),
    .X(uio_out[2]));
 sg13g2_buf_1 output5 (.A(net5),
    .X(uio_out[4]));
 sg13g2_buf_1 output6 (.A(net6),
    .X(uio_out[5]));
 sg13g2_buf_1 output7 (.A(net7),
    .X(uo_out[0]));
 sg13g2_buf_1 output8 (.A(net8),
    .X(uo_out[1]));
 sg13g2_buf_1 output9 (.A(net9),
    .X(uo_out[2]));
 sg13g2_buf_1 output10 (.A(net10),
    .X(uo_out[3]));
 sg13g2_buf_1 output11 (.A(net11),
    .X(uo_out[4]));
 sg13g2_buf_1 output12 (.A(net12),
    .X(uo_out[5]));
 sg13g2_buf_1 output13 (.A(net13),
    .X(uo_out[6]));
 sg13g2_buf_1 output14 (.A(net14),
    .X(uo_out[7]));
 sg13g2_buf_2 fanout15 (.A(_1077_),
    .X(net15));
 sg13g2_buf_2 fanout16 (.A(_0997_),
    .X(net16));
 sg13g2_buf_2 fanout17 (.A(_0734_),
    .X(net17));
 sg13g2_buf_2 fanout18 (.A(_0728_),
    .X(net18));
 sg13g2_buf_2 fanout19 (.A(_0726_),
    .X(net19));
 sg13g2_buf_2 fanout20 (.A(_0646_),
    .X(net20));
 sg13g2_buf_2 fanout21 (.A(_1935_),
    .X(net21));
 sg13g2_buf_2 fanout22 (.A(_1931_),
    .X(net22));
 sg13g2_buf_2 fanout23 (.A(_1733_),
    .X(net23));
 sg13g2_buf_2 fanout24 (.A(_1721_),
    .X(net24));
 sg13g2_buf_2 fanout25 (.A(_1717_),
    .X(net25));
 sg13g2_buf_2 fanout26 (.A(_1406_),
    .X(net26));
 sg13g2_buf_2 fanout27 (.A(_0972_),
    .X(net27));
 sg13g2_buf_2 fanout28 (.A(_0970_),
    .X(net28));
 sg13g2_buf_2 fanout29 (.A(_0725_),
    .X(net29));
 sg13g2_buf_2 fanout30 (.A(_0656_),
    .X(net30));
 sg13g2_buf_2 fanout31 (.A(_0652_),
    .X(net31));
 sg13g2_buf_2 fanout32 (.A(_0487_),
    .X(net32));
 sg13g2_buf_2 fanout33 (.A(_0486_),
    .X(net33));
 sg13g2_buf_2 fanout34 (.A(_2967_),
    .X(net34));
 sg13g2_buf_2 fanout35 (.A(_2954_),
    .X(net35));
 sg13g2_buf_2 fanout36 (.A(_2892_),
    .X(net36));
 sg13g2_buf_2 fanout37 (.A(_2887_),
    .X(net37));
 sg13g2_buf_2 fanout38 (.A(_2754_),
    .X(net38));
 sg13g2_buf_2 fanout39 (.A(_1915_),
    .X(net39));
 sg13g2_buf_2 fanout40 (.A(_1411_),
    .X(net40));
 sg13g2_buf_2 fanout41 (.A(_1250_),
    .X(net41));
 sg13g2_buf_2 fanout42 (.A(_1006_),
    .X(net42));
 sg13g2_buf_2 fanout43 (.A(_0969_),
    .X(net43));
 sg13g2_buf_2 fanout44 (.A(_0635_),
    .X(net44));
 sg13g2_buf_2 fanout45 (.A(_0491_),
    .X(net45));
 sg13g2_buf_2 fanout46 (.A(_0467_),
    .X(net46));
 sg13g2_buf_2 fanout47 (.A(_0466_),
    .X(net47));
 sg13g2_buf_2 fanout48 (.A(_0465_),
    .X(net48));
 sg13g2_buf_2 fanout49 (.A(_0460_),
    .X(net49));
 sg13g2_buf_2 fanout50 (.A(_3049_),
    .X(net50));
 sg13g2_buf_2 fanout51 (.A(_3047_),
    .X(net51));
 sg13g2_buf_2 fanout52 (.A(_2897_),
    .X(net52));
 sg13g2_buf_2 fanout53 (.A(_2893_),
    .X(net53));
 sg13g2_buf_2 fanout54 (.A(_2886_),
    .X(net54));
 sg13g2_buf_2 fanout55 (.A(_2885_),
    .X(net55));
 sg13g2_buf_2 fanout56 (.A(_2766_),
    .X(net56));
 sg13g2_buf_2 fanout57 (.A(_2764_),
    .X(net57));
 sg13g2_buf_2 fanout58 (.A(_2761_),
    .X(net58));
 sg13g2_buf_2 fanout59 (.A(_2759_),
    .X(net59));
 sg13g2_buf_2 fanout60 (.A(_2753_),
    .X(net60));
 sg13g2_buf_2 fanout61 (.A(_2750_),
    .X(net61));
 sg13g2_buf_2 fanout62 (.A(_2698_),
    .X(net62));
 sg13g2_buf_2 fanout63 (.A(_1619_),
    .X(net63));
 sg13g2_buf_2 fanout64 (.A(_1614_),
    .X(net64));
 sg13g2_buf_2 fanout65 (.A(_1547_),
    .X(net65));
 sg13g2_buf_2 fanout66 (.A(_0975_),
    .X(net66));
 sg13g2_buf_2 fanout67 (.A(_3048_),
    .X(net67));
 sg13g2_buf_2 fanout68 (.A(_3042_),
    .X(net68));
 sg13g2_buf_4 fanout69 (.X(net69),
    .A(_2951_));
 sg13g2_buf_2 fanout70 (.A(_2932_),
    .X(net70));
 sg13g2_buf_2 fanout71 (.A(_2899_),
    .X(net71));
 sg13g2_buf_2 fanout72 (.A(_2774_),
    .X(net72));
 sg13g2_buf_2 fanout73 (.A(_2763_),
    .X(net73));
 sg13g2_buf_2 fanout74 (.A(_2758_),
    .X(net74));
 sg13g2_buf_2 fanout75 (.A(_1075_),
    .X(net75));
 sg13g2_buf_2 fanout76 (.A(_1067_),
    .X(net76));
 sg13g2_buf_2 fanout77 (.A(_0959_),
    .X(net77));
 sg13g2_buf_2 fanout78 (.A(_0946_),
    .X(net78));
 sg13g2_buf_2 fanout79 (.A(_0567_),
    .X(net79));
 sg13g2_buf_2 fanout80 (.A(net82),
    .X(net80));
 sg13g2_buf_1 fanout81 (.A(net82),
    .X(net81));
 sg13g2_buf_2 fanout82 (.A(\Pong.datapath.Ball_Clock.roll ),
    .X(net82));
 sg13g2_buf_2 fanout83 (.A(_2787_),
    .X(net83));
 sg13g2_buf_2 fanout84 (.A(_2654_),
    .X(net84));
 sg13g2_buf_2 fanout85 (.A(_2651_),
    .X(net85));
 sg13g2_buf_2 fanout86 (.A(_1555_),
    .X(net86));
 sg13g2_buf_2 fanout87 (.A(_0964_),
    .X(net87));
 sg13g2_buf_2 fanout88 (.A(_0945_),
    .X(net88));
 sg13g2_buf_2 fanout89 (.A(_2800_),
    .X(net89));
 sg13g2_buf_2 fanout90 (.A(_2789_),
    .X(net90));
 sg13g2_buf_2 fanout91 (.A(_2786_),
    .X(net91));
 sg13g2_buf_2 fanout92 (.A(_2653_),
    .X(net92));
 sg13g2_buf_2 fanout93 (.A(_2650_),
    .X(net93));
 sg13g2_buf_2 fanout94 (.A(_0962_),
    .X(net94));
 sg13g2_buf_2 fanout95 (.A(_1357_),
    .X(net95));
 sg13g2_buf_2 fanout96 (.A(_0730_),
    .X(net96));
 sg13g2_buf_2 fanout97 (.A(_0695_),
    .X(net97));
 sg13g2_buf_2 fanout98 (.A(_0602_),
    .X(net98));
 sg13g2_buf_2 fanout99 (.A(_0440_),
    .X(net99));
 sg13g2_buf_2 fanout100 (.A(_0403_),
    .X(net100));
 sg13g2_buf_2 fanout101 (.A(_0382_),
    .X(net101));
 sg13g2_buf_2 fanout102 (.A(_0327_),
    .X(net102));
 sg13g2_buf_2 fanout103 (.A(_0324_),
    .X(net103));
 sg13g2_buf_2 fanout104 (.A(_2910_),
    .X(net104));
 sg13g2_buf_2 fanout105 (.A(_2905_),
    .X(net105));
 sg13g2_buf_2 fanout106 (.A(_2855_),
    .X(net106));
 sg13g2_buf_2 fanout107 (.A(_2796_),
    .X(net107));
 sg13g2_buf_2 fanout108 (.A(_2701_),
    .X(net108));
 sg13g2_buf_2 fanout109 (.A(_2664_),
    .X(net109));
 sg13g2_buf_2 fanout110 (.A(_2172_),
    .X(net110));
 sg13g2_buf_2 fanout111 (.A(_1741_),
    .X(net111));
 sg13g2_buf_2 fanout112 (.A(_1667_),
    .X(net112));
 sg13g2_buf_2 fanout113 (.A(_1646_),
    .X(net113));
 sg13g2_buf_2 fanout114 (.A(_1644_),
    .X(net114));
 sg13g2_buf_2 fanout115 (.A(_1640_),
    .X(net115));
 sg13g2_buf_2 fanout116 (.A(_1637_),
    .X(net116));
 sg13g2_buf_2 fanout117 (.A(_1630_),
    .X(net117));
 sg13g2_buf_2 fanout118 (.A(_1626_),
    .X(net118));
 sg13g2_buf_2 fanout119 (.A(_1623_),
    .X(net119));
 sg13g2_buf_2 fanout120 (.A(_1611_),
    .X(net120));
 sg13g2_buf_2 fanout121 (.A(_1596_),
    .X(net121));
 sg13g2_buf_2 fanout122 (.A(_1593_),
    .X(net122));
 sg13g2_buf_2 fanout123 (.A(_1560_),
    .X(net123));
 sg13g2_buf_2 fanout124 (.A(_1538_),
    .X(net124));
 sg13g2_buf_2 fanout125 (.A(_1533_),
    .X(net125));
 sg13g2_buf_2 fanout126 (.A(_1529_),
    .X(net126));
 sg13g2_buf_2 fanout127 (.A(_1524_),
    .X(net127));
 sg13g2_buf_2 fanout128 (.A(_1515_),
    .X(net128));
 sg13g2_buf_2 fanout129 (.A(_1491_),
    .X(net129));
 sg13g2_buf_2 fanout130 (.A(_1407_),
    .X(net130));
 sg13g2_buf_2 fanout131 (.A(_1394_),
    .X(net131));
 sg13g2_buf_2 fanout132 (.A(_1260_),
    .X(net132));
 sg13g2_buf_2 fanout133 (.A(_1190_),
    .X(net133));
 sg13g2_buf_2 fanout134 (.A(_1187_),
    .X(net134));
 sg13g2_buf_2 fanout135 (.A(_1152_),
    .X(net135));
 sg13g2_buf_1 fanout136 (.A(_0983_),
    .X(net136));
 sg13g2_buf_2 fanout137 (.A(_0939_),
    .X(net137));
 sg13g2_buf_2 fanout138 (.A(_0801_),
    .X(net138));
 sg13g2_buf_2 fanout139 (.A(_0628_),
    .X(net139));
 sg13g2_buf_2 fanout140 (.A(_0400_),
    .X(net140));
 sg13g2_buf_2 fanout141 (.A(_0399_),
    .X(net141));
 sg13g2_buf_2 fanout142 (.A(_0365_),
    .X(net142));
 sg13g2_buf_2 fanout143 (.A(_0348_),
    .X(net143));
 sg13g2_buf_2 fanout144 (.A(_0333_),
    .X(net144));
 sg13g2_buf_2 fanout145 (.A(_0326_),
    .X(net145));
 sg13g2_buf_2 fanout146 (.A(_0325_),
    .X(net146));
 sg13g2_buf_2 fanout147 (.A(_0316_),
    .X(net147));
 sg13g2_buf_2 fanout148 (.A(_0312_),
    .X(net148));
 sg13g2_buf_2 fanout149 (.A(_2991_),
    .X(net149));
 sg13g2_buf_2 fanout150 (.A(_2946_),
    .X(net150));
 sg13g2_buf_2 fanout151 (.A(_2937_),
    .X(net151));
 sg13g2_buf_2 fanout152 (.A(_2933_),
    .X(net152));
 sg13g2_buf_2 fanout153 (.A(_2930_),
    .X(net153));
 sg13g2_buf_2 fanout154 (.A(_2918_),
    .X(net154));
 sg13g2_buf_2 fanout155 (.A(_2904_),
    .X(net155));
 sg13g2_buf_2 fanout156 (.A(_2902_),
    .X(net156));
 sg13g2_buf_2 fanout157 (.A(_2663_),
    .X(net157));
 sg13g2_buf_2 fanout158 (.A(_2658_),
    .X(net158));
 sg13g2_buf_2 fanout159 (.A(_1632_),
    .X(net159));
 sg13g2_buf_2 fanout160 (.A(_1607_),
    .X(net160));
 sg13g2_buf_2 fanout161 (.A(_1606_),
    .X(net161));
 sg13g2_buf_2 fanout162 (.A(_1570_),
    .X(net162));
 sg13g2_buf_2 fanout163 (.A(_1561_),
    .X(net163));
 sg13g2_buf_2 fanout164 (.A(_1556_),
    .X(net164));
 sg13g2_buf_2 fanout165 (.A(_1541_),
    .X(net165));
 sg13g2_buf_2 fanout166 (.A(_1539_),
    .X(net166));
 sg13g2_buf_2 fanout167 (.A(_1508_),
    .X(net167));
 sg13g2_buf_2 fanout168 (.A(_1214_),
    .X(net168));
 sg13g2_buf_2 fanout169 (.A(_1175_),
    .X(net169));
 sg13g2_buf_2 fanout170 (.A(_1162_),
    .X(net170));
 sg13g2_buf_2 fanout171 (.A(_1157_),
    .X(net171));
 sg13g2_buf_2 fanout172 (.A(_1155_),
    .X(net172));
 sg13g2_buf_2 fanout173 (.A(_1154_),
    .X(net173));
 sg13g2_buf_2 fanout174 (.A(_0409_),
    .X(net174));
 sg13g2_buf_2 fanout175 (.A(_0383_),
    .X(net175));
 sg13g2_buf_2 fanout176 (.A(_0347_),
    .X(net176));
 sg13g2_buf_2 fanout177 (.A(_0318_),
    .X(net177));
 sg13g2_buf_2 fanout178 (.A(_0314_),
    .X(net178));
 sg13g2_buf_2 fanout179 (.A(_2984_),
    .X(net179));
 sg13g2_buf_2 fanout180 (.A(_2945_),
    .X(net180));
 sg13g2_buf_2 fanout181 (.A(_2924_),
    .X(net181));
 sg13g2_buf_2 fanout182 (.A(_2912_),
    .X(net182));
 sg13g2_buf_2 fanout183 (.A(_2908_),
    .X(net183));
 sg13g2_buf_2 fanout184 (.A(_2901_),
    .X(net184));
 sg13g2_buf_2 fanout185 (.A(_2895_),
    .X(net185));
 sg13g2_buf_2 fanout186 (.A(_2737_),
    .X(net186));
 sg13g2_buf_2 fanout187 (.A(_2720_),
    .X(net187));
 sg13g2_buf_2 fanout188 (.A(_2717_),
    .X(net188));
 sg13g2_tielo _6189__189 (.L_LO(net189));
 sg13g2_tielo _6192__190 (.L_LO(net190));
 sg13g2_tielo _6195__191 (.L_LO(net191));
 sg13g2_tielo _6196__192 (.L_LO(net192));
 sg13g2_tielo _6197__193 (.L_LO(net193));
 sg13g2_tielo _6198__194 (.L_LO(net194));
 sg13g2_tielo _6199__195 (.L_LO(net195));
 sg13g2_tielo _6200__196 (.L_LO(net196));
 sg13g2_tiehi \Pong.control_unit.NES_Controller_Left.state_NESController[10]$_DFF_P__198  (.L_HI(net198));
 sg13g2_tiehi \Pong.control_unit.NES_Controller_Left.state_NESController[11]$_DFF_P__199  (.L_HI(net199));
 sg13g2_tiehi \Pong.control_unit.NES_Controller_Left.state_NESController[12]$_DFF_P__200  (.L_HI(net200));
 sg13g2_tiehi \Pong.control_unit.NES_Controller_Left.state_NESController[13]$_DFF_P__201  (.L_HI(net201));
 sg13g2_tiehi \Pong.control_unit.NES_Controller_Left.state_NESController[14]$_DFF_P__202  (.L_HI(net202));
 sg13g2_tiehi \Pong.control_unit.NES_Controller_Left.state_NESController[15]$_DFF_P__203  (.L_HI(net203));
 sg13g2_tiehi \Pong.control_unit.NES_Controller_Left.state_NESController[16]$_DFF_P__204  (.L_HI(net204));
 sg13g2_tiehi \Pong.control_unit.NES_Controller_Left.state_NESController[17]$_DFF_P__205  (.L_HI(net205));
 sg13g2_tiehi \Pong.control_unit.NES_Controller_Left.state_NESController[18]$_DFF_P__206  (.L_HI(net206));
 sg13g2_tiehi \Pong.control_unit.NES_Controller_Left.state_NESController[1]$_DFF_P__207  (.L_HI(net207));
 sg13g2_tiehi \Pong.control_unit.NES_Controller_Left.state_NESController[2]$_DFF_P__208  (.L_HI(net208));
 sg13g2_tiehi \Pong.control_unit.NES_Controller_Left.state_NESController[3]$_DFF_P__209  (.L_HI(net209));
 sg13g2_tiehi \Pong.control_unit.NES_Controller_Left.state_NESController[4]$_DFF_P__210  (.L_HI(net210));
 sg13g2_tiehi \Pong.control_unit.NES_Controller_Left.state_NESController[5]$_DFF_P__211  (.L_HI(net211));
 sg13g2_tiehi \Pong.control_unit.NES_Controller_Left.state_NESController[6]$_DFF_P__212  (.L_HI(net212));
 sg13g2_tiehi \Pong.control_unit.NES_Controller_Left.state_NESController[7]$_DFF_P__213  (.L_HI(net213));
 sg13g2_tiehi \Pong.control_unit.NES_Controller_Left.state_NESController[8]$_DFF_P__214  (.L_HI(net214));
 sg13g2_tiehi \Pong.control_unit.NES_Controller_Left.state_NESController[9]$_DFF_P__215  (.L_HI(net215));
 sg13g2_tiehi \Pong.control_unit.NES_Controller_Right.state_NESController[0]$_DFF_P__216  (.L_HI(net216));
 sg13g2_tiehi \Pong.control_unit.NES_Controller_Right.state_NESController[10]$_DFF_P__217  (.L_HI(net217));
 sg13g2_tiehi \Pong.control_unit.NES_Controller_Right.state_NESController[11]$_DFF_P__218  (.L_HI(net218));
 sg13g2_tiehi \Pong.control_unit.NES_Controller_Right.state_NESController[12]$_DFF_P__219  (.L_HI(net219));
 sg13g2_tiehi \Pong.control_unit.NES_Controller_Right.state_NESController[13]$_DFF_P__220  (.L_HI(net220));
 sg13g2_tiehi \Pong.control_unit.NES_Controller_Right.state_NESController[14]$_DFF_P__221  (.L_HI(net221));
 sg13g2_tiehi \Pong.control_unit.NES_Controller_Right.state_NESController[15]$_DFF_P__222  (.L_HI(net222));
 sg13g2_tiehi \Pong.control_unit.NES_Controller_Right.state_NESController[16]$_DFF_P__223  (.L_HI(net223));
 sg13g2_tiehi \Pong.control_unit.NES_Controller_Right.state_NESController[17]$_DFF_P__224  (.L_HI(net224));
 sg13g2_tiehi \Pong.control_unit.NES_Controller_Right.state_NESController[18]$_DFF_P__225  (.L_HI(net225));
 sg13g2_tiehi \Pong.control_unit.NES_Controller_Right.state_NESController[1]$_DFF_P__226  (.L_HI(net226));
 sg13g2_tiehi \Pong.control_unit.NES_Controller_Right.state_NESController[2]$_DFF_P__227  (.L_HI(net227));
 sg13g2_tiehi \Pong.control_unit.NES_Controller_Right.state_NESController[3]$_DFF_P__228  (.L_HI(net228));
 sg13g2_tiehi \Pong.control_unit.NES_Controller_Right.state_NESController[4]$_DFF_P__229  (.L_HI(net229));
 sg13g2_tiehi \Pong.control_unit.NES_Controller_Right.state_NESController[5]$_DFF_P__230  (.L_HI(net230));
 sg13g2_tiehi \Pong.control_unit.NES_Controller_Right.state_NESController[6]$_DFF_P__231  (.L_HI(net231));
 sg13g2_tiehi \Pong.control_unit.NES_Controller_Right.state_NESController[7]$_DFF_P__232  (.L_HI(net232));
 sg13g2_tiehi \Pong.control_unit.NES_Controller_Right.state_NESController[8]$_DFF_P__233  (.L_HI(net233));
 sg13g2_tiehi \Pong.control_unit.NES_Controller_Right.state_NESController[9]$_DFF_P__234  (.L_HI(net234));
 sg13g2_tiehi \Pong.control_unit.state_ballMovement[0]$_DFF_P__235  (.L_HI(net235));
 sg13g2_tiehi \Pong.control_unit.state_ballMovement[1]$_DFF_P__236  (.L_HI(net236));
 sg13g2_tiehi \Pong.control_unit.state_ballMovement[2]$_DFF_P__237  (.L_HI(net237));
 sg13g2_tiehi \Pong.control_unit.state_ballMovement[3]$_DFF_P__238  (.L_HI(net238));
 sg13g2_tiehi \Pong.control_unit.state_ballMovement[4]$_DFF_P__239  (.L_HI(net239));
 sg13g2_tiehi \Pong.datapath.Ball_Clock.processQ[0]$_SDFFE_PN0P__240  (.L_HI(net240));
 sg13g2_tiehi \Pong.datapath.Ball_Clock.processQ[10]$_SDFFE_PN0P__241  (.L_HI(net241));
 sg13g2_tiehi \Pong.datapath.Ball_Clock.processQ[11]$_SDFFE_PN0P__242  (.L_HI(net242));
 sg13g2_tiehi \Pong.datapath.Ball_Clock.processQ[12]$_SDFFE_PN0P__243  (.L_HI(net243));
 sg13g2_tiehi \Pong.datapath.Ball_Clock.processQ[13]$_SDFFE_PN0P__244  (.L_HI(net244));
 sg13g2_tiehi \Pong.datapath.Ball_Clock.processQ[14]$_SDFFE_PN0P__245  (.L_HI(net245));
 sg13g2_tiehi \Pong.datapath.Ball_Clock.processQ[15]$_SDFFE_PN0P__246  (.L_HI(net246));
 sg13g2_tiehi \Pong.datapath.Ball_Clock.processQ[16]$_SDFFE_PN0P__247  (.L_HI(net247));
 sg13g2_tiehi \Pong.datapath.Ball_Clock.processQ[1]$_SDFFE_PN0P__248  (.L_HI(net248));
 sg13g2_tiehi \Pong.datapath.Ball_Clock.processQ[2]$_SDFFE_PN0P__249  (.L_HI(net249));
 sg13g2_tiehi \Pong.datapath.Ball_Clock.processQ[3]$_SDFFE_PN0P__250  (.L_HI(net250));
 sg13g2_tiehi \Pong.datapath.Ball_Clock.processQ[4]$_SDFFE_PN0P__251  (.L_HI(net251));
 sg13g2_tiehi \Pong.datapath.Ball_Clock.processQ[5]$_SDFFE_PN0P__252  (.L_HI(net252));
 sg13g2_tiehi \Pong.datapath.Ball_Clock.processQ[6]$_SDFFE_PN0P__253  (.L_HI(net253));
 sg13g2_tiehi \Pong.datapath.Ball_Clock.processQ[7]$_SDFFE_PN0P__254  (.L_HI(net254));
 sg13g2_tiehi \Pong.datapath.Ball_Clock.processQ[8]$_SDFFE_PN0P__255  (.L_HI(net255));
 sg13g2_tiehi \Pong.datapath.Ball_Clock.processQ[9]$_SDFFE_PN0P__256  (.L_HI(net256));
 sg13g2_tiehi \Pong.datapath.NES_activity_Left[2]$_SDFF_PP0__257  (.L_HI(net257));
 sg13g2_tiehi \Pong.datapath.NES_activity_Left[3]$_SDFF_PP0__258  (.L_HI(net258));
 sg13g2_tiehi \Pong.datapath.NES_activity_Left[4]$_SDFF_PP0__259  (.L_HI(net259));
 sg13g2_tiehi \Pong.datapath.NES_activity_Left[5]$_SDFF_PP0__260  (.L_HI(net260));
 sg13g2_tiehi \Pong.datapath.NES_activity_Right[2]$_SDFF_PP0__261  (.L_HI(net261));
 sg13g2_tiehi \Pong.datapath.NES_activity_Right[3]$_SDFF_PP0__262  (.L_HI(net262));
 sg13g2_tiehi \Pong.datapath.NES_activity_Right[4]$_SDFF_PP0__263  (.L_HI(net263));
 sg13g2_tiehi \Pong.datapath.NES_activity_Right[5]$_SDFF_PP0__264  (.L_HI(net264));
 sg13g2_tiehi \Pong.datapath.NES_counter_left.processQ[0]$_SDFFE_PP0P__265  (.L_HI(net265));
 sg13g2_tiehi \Pong.datapath.NES_counter_left.processQ[1]$_SDFFE_PP0P__266  (.L_HI(net266));
 sg13g2_tiehi \Pong.datapath.NES_counter_left.processQ[2]$_SDFFE_PP0P__267  (.L_HI(net267));
 sg13g2_tiehi \Pong.datapath.NES_counter_left.processQ[3]$_SDFFE_PP0P__268  (.L_HI(net268));
 sg13g2_tiehi \Pong.datapath.NES_counter_left.processQ[4]$_SDFFE_PP0P__269  (.L_HI(net269));
 sg13g2_tiehi \Pong.datapath.NES_counter_left.processQ[5]$_SDFFE_PP0P__270  (.L_HI(net270));
 sg13g2_tiehi \Pong.datapath.NES_counter_left.processQ[6]$_SDFFE_PP0P__271  (.L_HI(net271));
 sg13g2_tiehi \Pong.datapath.NES_counter_left.processQ[7]$_SDFFE_PP0P__272  (.L_HI(net272));
 sg13g2_tiehi \Pong.datapath.NES_counter_right.processQ[0]$_SDFFE_PP0P__273  (.L_HI(net273));
 sg13g2_tiehi \Pong.datapath.NES_counter_right.processQ[1]$_SDFFE_PP0P__274  (.L_HI(net274));
 sg13g2_tiehi \Pong.datapath.NES_counter_right.processQ[2]$_SDFFE_PP0P__275  (.L_HI(net275));
 sg13g2_tiehi \Pong.datapath.NES_counter_right.processQ[3]$_SDFFE_PP0P__276  (.L_HI(net276));
 sg13g2_tiehi \Pong.datapath.NES_counter_right.processQ[4]$_SDFFE_PP0P__277  (.L_HI(net277));
 sg13g2_tiehi \Pong.datapath.NES_counter_right.processQ[5]$_SDFFE_PP0P__278  (.L_HI(net278));
 sg13g2_tiehi \Pong.datapath.NES_counter_right.processQ[6]$_SDFFE_PP0P__279  (.L_HI(net279));
 sg13g2_tiehi \Pong.datapath.NES_counter_right.processQ[7]$_SDFFE_PP0P__280  (.L_HI(net280));
 sg13g2_tiehi \Pong.datapath.NES_delay_counter_left.processQ[0]$_SDFFE_PN0P__281  (.L_HI(net281));
 sg13g2_tiehi \Pong.datapath.NES_delay_counter_left.processQ[10]$_SDFFE_PN0P__282  (.L_HI(net282));
 sg13g2_tiehi \Pong.datapath.NES_delay_counter_left.processQ[11]$_SDFFE_PN0P__283  (.L_HI(net283));
 sg13g2_tiehi \Pong.datapath.NES_delay_counter_left.processQ[12]$_SDFFE_PN0P__284  (.L_HI(net284));
 sg13g2_tiehi \Pong.datapath.NES_delay_counter_left.processQ[13]$_SDFFE_PN0P__285  (.L_HI(net285));
 sg13g2_tiehi \Pong.datapath.NES_delay_counter_left.processQ[14]$_SDFFE_PN0P__286  (.L_HI(net286));
 sg13g2_tiehi \Pong.datapath.NES_delay_counter_left.processQ[15]$_SDFFE_PN0P__287  (.L_HI(net287));
 sg13g2_tiehi \Pong.datapath.NES_delay_counter_left.processQ[16]$_SDFFE_PN0P__288  (.L_HI(net288));
 sg13g2_tiehi \Pong.datapath.NES_delay_counter_left.processQ[17]$_SDFFE_PN0P__289  (.L_HI(net289));
 sg13g2_tiehi \Pong.datapath.NES_delay_counter_left.processQ[18]$_SDFFE_PN0P__290  (.L_HI(net290));
 sg13g2_tiehi \Pong.datapath.NES_delay_counter_left.processQ[1]$_SDFFE_PN0P__291  (.L_HI(net291));
 sg13g2_tiehi \Pong.datapath.NES_delay_counter_left.processQ[2]$_SDFFE_PN0P__292  (.L_HI(net292));
 sg13g2_tiehi \Pong.datapath.NES_delay_counter_left.processQ[3]$_SDFFE_PN0P__293  (.L_HI(net293));
 sg13g2_tiehi \Pong.datapath.NES_delay_counter_left.processQ[4]$_SDFFE_PN0P__294  (.L_HI(net294));
 sg13g2_tiehi \Pong.datapath.NES_delay_counter_left.processQ[5]$_SDFFE_PN0P__295  (.L_HI(net295));
 sg13g2_tiehi \Pong.datapath.NES_delay_counter_left.processQ[6]$_SDFFE_PN0P__296  (.L_HI(net296));
 sg13g2_tiehi \Pong.datapath.NES_delay_counter_left.processQ[7]$_SDFFE_PN0P__297  (.L_HI(net297));
 sg13g2_tiehi \Pong.datapath.NES_delay_counter_left.processQ[8]$_SDFFE_PN0P__298  (.L_HI(net298));
 sg13g2_tiehi \Pong.datapath.NES_delay_counter_left.processQ[9]$_SDFFE_PN0P__299  (.L_HI(net299));
 sg13g2_tiehi \Pong.datapath.NES_delay_counter_right.processQ[0]$_SDFFE_PN0P__300  (.L_HI(net300));
 sg13g2_tiehi \Pong.datapath.NES_delay_counter_right.processQ[10]$_SDFFE_PN0P__301  (.L_HI(net301));
 sg13g2_tiehi \Pong.datapath.NES_delay_counter_right.processQ[11]$_SDFFE_PN0P__302  (.L_HI(net302));
 sg13g2_tiehi \Pong.datapath.NES_delay_counter_right.processQ[12]$_SDFFE_PN0P__303  (.L_HI(net303));
 sg13g2_tiehi \Pong.datapath.NES_delay_counter_right.processQ[13]$_SDFFE_PN0P__304  (.L_HI(net304));
 sg13g2_tiehi \Pong.datapath.NES_delay_counter_right.processQ[14]$_SDFFE_PN0P__305  (.L_HI(net305));
 sg13g2_tiehi \Pong.datapath.NES_delay_counter_right.processQ[15]$_SDFFE_PN0P__306  (.L_HI(net306));
 sg13g2_tiehi \Pong.datapath.NES_delay_counter_right.processQ[16]$_SDFFE_PN0P__307  (.L_HI(net307));
 sg13g2_tiehi \Pong.datapath.NES_delay_counter_right.processQ[17]$_SDFFE_PN0P__308  (.L_HI(net308));
 sg13g2_tiehi \Pong.datapath.NES_delay_counter_right.processQ[18]$_SDFFE_PN0P__309  (.L_HI(net309));
 sg13g2_tiehi \Pong.datapath.NES_delay_counter_right.processQ[1]$_SDFFE_PN0P__310  (.L_HI(net310));
 sg13g2_tiehi \Pong.datapath.NES_delay_counter_right.processQ[2]$_SDFFE_PN0P__311  (.L_HI(net311));
 sg13g2_tiehi \Pong.datapath.NES_delay_counter_right.processQ[3]$_SDFFE_PN0P__312  (.L_HI(net312));
 sg13g2_tiehi \Pong.datapath.NES_delay_counter_right.processQ[4]$_SDFFE_PN0P__313  (.L_HI(net313));
 sg13g2_tiehi \Pong.datapath.NES_delay_counter_right.processQ[5]$_SDFFE_PN0P__314  (.L_HI(net314));
 sg13g2_tiehi \Pong.datapath.NES_delay_counter_right.processQ[6]$_SDFFE_PN0P__315  (.L_HI(net315));
 sg13g2_tiehi \Pong.datapath.NES_delay_counter_right.processQ[7]$_SDFFE_PN0P__316  (.L_HI(net316));
 sg13g2_tiehi \Pong.datapath.NES_delay_counter_right.processQ[8]$_SDFFE_PN0P__317  (.L_HI(net317));
 sg13g2_tiehi \Pong.datapath.NES_delay_counter_right.processQ[9]$_SDFFE_PN0P__318  (.L_HI(net318));
 sg13g2_tiehi \Pong.datapath.NES_wire_Left[2]$_SDFFE_PN0N__319  (.L_HI(net319));
 sg13g2_tiehi \Pong.datapath.NES_wire_Left[3]$_SDFFE_PN0N__320  (.L_HI(net320));
 sg13g2_tiehi \Pong.datapath.NES_wire_Left[4]$_SDFFE_PN0N__321  (.L_HI(net321));
 sg13g2_tiehi \Pong.datapath.NES_wire_Left[5]$_SDFFE_PN0N__322  (.L_HI(net322));
 sg13g2_tiehi \Pong.datapath.NES_wire_Right[2]$_SDFFE_PN0N__323  (.L_HI(net323));
 sg13g2_tiehi \Pong.datapath.NES_wire_Right[3]$_SDFFE_PN0N__324  (.L_HI(net324));
 sg13g2_tiehi \Pong.datapath.NES_wire_Right[4]$_SDFFE_PN0N__325  (.L_HI(net325));
 sg13g2_tiehi \Pong.datapath.NES_wire_Right[5]$_SDFFE_PN0N__326  (.L_HI(net326));
 sg13g2_tiehi \Pong.datapath.ballFunction.ball_center_x_proc[0]$_SDFFE_PN0P__327  (.L_HI(net327));
 sg13g2_tiehi \Pong.datapath.ballFunction.ball_center_x_proc[1]$_SDFFE_PN0P__328  (.L_HI(net328));
 sg13g2_tiehi \Pong.datapath.ballFunction.ball_center_x_proc[2]$_SDFFE_PN0P__329  (.L_HI(net329));
 sg13g2_tiehi \Pong.datapath.ballFunction.ball_center_x_proc[3]$_SDFFE_PN0P__330  (.L_HI(net330));
 sg13g2_tiehi \Pong.datapath.ballFunction.ball_center_x_proc[4]$_SDFFE_PN0P__331  (.L_HI(net331));
 sg13g2_tiehi \Pong.datapath.ballFunction.ball_center_x_proc[5]$_SDFFE_PN0P__332  (.L_HI(net332));
 sg13g2_tiehi \Pong.datapath.ballFunction.ball_center_x_proc[6]$_SDFFE_PN1P__333  (.L_HI(net333));
 sg13g2_tiehi \Pong.datapath.ballFunction.ball_center_x_proc[7]$_SDFFE_PN0P__334  (.L_HI(net334));
 sg13g2_tiehi \Pong.datapath.ballFunction.ball_center_x_proc[8]$_SDFFE_PN1P__335  (.L_HI(net335));
 sg13g2_tiehi \Pong.datapath.ballFunction.ball_center_x_proc[9]$_SDFFE_PN0P__336  (.L_HI(net336));
 sg13g2_tiehi \Pong.datapath.ballFunction.ball_center_y_proc[0]$_SDFFE_PN0P__337  (.L_HI(net337));
 sg13g2_tiehi \Pong.datapath.ballFunction.ball_center_y_proc[1]$_SDFFE_PN0P__338  (.L_HI(net338));
 sg13g2_tiehi \Pong.datapath.ballFunction.ball_center_y_proc[2]$_SDFFE_PN1P__339  (.L_HI(net339));
 sg13g2_tiehi \Pong.datapath.ballFunction.ball_center_y_proc[3]$_SDFFE_PN1P__340  (.L_HI(net340));
 sg13g2_tiehi \Pong.datapath.ballFunction.ball_center_y_proc[4]$_SDFFE_PN1P__341  (.L_HI(net341));
 sg13g2_tiehi \Pong.datapath.ballFunction.ball_center_y_proc[5]$_SDFFE_PN0P__342  (.L_HI(net342));
 sg13g2_tiehi \Pong.datapath.ballFunction.ball_center_y_proc[6]$_SDFFE_PN1P__343  (.L_HI(net343));
 sg13g2_tiehi \Pong.datapath.ballFunction.ball_center_y_proc[7]$_SDFFE_PN1P__344  (.L_HI(net344));
 sg13g2_tiehi \Pong.datapath.ballFunction.ball_center_y_proc[8]$_SDFFE_PN0P__345  (.L_HI(net345));
 sg13g2_tiehi \Pong.datapath.ballFunction.ball_center_y_proc[9]$_SDFFE_PN0P__346  (.L_HI(net346));
 sg13g2_tiehi \Pong.datapath.ballReset$_SDFF_PN0__347  (.L_HI(net347));
 sg13g2_tiehi \Pong.datapath.leftPaddle[0]$_SDFF_PN0__348  (.L_HI(net348));
 sg13g2_tiehi \Pong.datapath.leftPaddle[1]$_SDFF_PN0__349  (.L_HI(net349));
 sg13g2_tiehi \Pong.datapath.leftPaddle[2]$_SDFF_PN1__350  (.L_HI(net350));
 sg13g2_tiehi \Pong.datapath.leftPaddle[3]$_SDFF_PN1__351  (.L_HI(net351));
 sg13g2_tiehi \Pong.datapath.leftPaddle[4]$_SDFF_PN1__352  (.L_HI(net352));
 sg13g2_tiehi \Pong.datapath.leftPaddle[5]$_SDFF_PN0__353  (.L_HI(net353));
 sg13g2_tiehi \Pong.datapath.leftPaddle[6]$_SDFF_PN1__354  (.L_HI(net354));
 sg13g2_tiehi \Pong.datapath.leftPaddle[7]$_SDFF_PN1__355  (.L_HI(net355));
 sg13g2_tiehi \Pong.datapath.leftPaddle[8]$_SDFF_PN0__356  (.L_HI(net356));
 sg13g2_tiehi \Pong.datapath.leftPaddle[9]$_SDFF_PN0__357  (.L_HI(net357));
 sg13g2_tiehi \Pong.datapath.old_NES_Left[2]$_SDFF_PN0__358  (.L_HI(net358));
 sg13g2_tiehi \Pong.datapath.old_NES_Left[3]$_SDFF_PN0__359  (.L_HI(net359));
 sg13g2_tiehi \Pong.datapath.old_NES_Left[4]$_SDFF_PN0__360  (.L_HI(net360));
 sg13g2_tiehi \Pong.datapath.old_NES_Left[5]$_SDFF_PN0__361  (.L_HI(net361));
 sg13g2_tiehi \Pong.datapath.old_NES_Right[2]$_SDFF_PN0__362  (.L_HI(net362));
 sg13g2_tiehi \Pong.datapath.old_NES_Right[3]$_SDFF_PN0__363  (.L_HI(net363));
 sg13g2_tiehi \Pong.datapath.old_NES_Right[4]$_SDFF_PN0__364  (.L_HI(net364));
 sg13g2_tiehi \Pong.datapath.old_NES_Right[5]$_SDFF_PN0__365  (.L_HI(net365));
 sg13g2_tiehi \Pong.datapath.rightPaddle[0]$_SDFF_PN0__366  (.L_HI(net366));
 sg13g2_tiehi \Pong.datapath.rightPaddle[1]$_SDFF_PN0__367  (.L_HI(net367));
 sg13g2_tiehi \Pong.datapath.rightPaddle[2]$_SDFF_PN1__368  (.L_HI(net368));
 sg13g2_tiehi \Pong.datapath.rightPaddle[3]$_SDFF_PN1__369  (.L_HI(net369));
 sg13g2_tiehi \Pong.datapath.rightPaddle[4]$_SDFF_PN1__370  (.L_HI(net370));
 sg13g2_tiehi \Pong.datapath.rightPaddle[5]$_SDFF_PN0__371  (.L_HI(net371));
 sg13g2_tiehi \Pong.datapath.rightPaddle[6]$_SDFF_PN1__372  (.L_HI(net372));
 sg13g2_tiehi \Pong.datapath.rightPaddle[7]$_SDFF_PN1__373  (.L_HI(net373));
 sg13g2_tiehi \Pong.datapath.rightPaddle[8]$_SDFF_PN0__374  (.L_HI(net374));
 sg13g2_tiehi \Pong.datapath.rightPaddle[9]$_SDFF_PN0__375  (.L_HI(net375));
 sg13g2_tiehi \Pong.datapath.scoreLeftProc[0]$_SDFF_PN0__376  (.L_HI(net376));
 sg13g2_tiehi \Pong.datapath.scoreLeftProc[1]$_SDFF_PN0__377  (.L_HI(net377));
 sg13g2_tiehi \Pong.datapath.scoreLeftProc[2]$_SDFF_PN0__378  (.L_HI(net378));
 sg13g2_tiehi \Pong.datapath.scoreLeftProc[3]$_SDFF_PN0__379  (.L_HI(net379));
 sg13g2_tiehi \Pong.datapath.scoreRightProc[0]$_SDFF_PN0__380  (.L_HI(net380));
 sg13g2_tiehi \Pong.datapath.scoreRightProc[1]$_SDFF_PN0__381  (.L_HI(net381));
 sg13g2_tiehi \Pong.datapath.scoreRightProc[2]$_SDFF_PN0__382  (.L_HI(net382));
 sg13g2_tiehi \Pong.datapath.scoreRightProc[3]$_SDFF_PN0__383  (.L_HI(net383));
 sg13g2_tiehi \Pong.datapath.score_flag$_SDFF_PN1__384  (.L_HI(net384));
 sg13g2_tiehi \Pong.datapath.sw_ballMovement_reg[0]$_DFF_P__385  (.L_HI(net385));
 sg13g2_tiehi \Pong.datapath.sw_ballMovement_reg[2]$_DFF_P__386  (.L_HI(net386));
 sg13g2_tiehi \Pong.datapath.sw_ballMovement_reg[3]$_DFF_P__387  (.L_HI(net387));
 sg13g2_tiehi \Pong.datapath.sw_ballMovement_reg[4]$_DFF_P__388  (.L_HI(net388));
 sg13g2_tiehi \Pong.datapath.sw_ballMovement_reg[5]$_DFF_P__389  (.L_HI(net389));
 sg13g2_tiehi \Pong.datapath.vga.Column_Counter.processQ[0]$_SDFFE_PN0P__390  (.L_HI(net390));
 sg13g2_tiehi \Pong.datapath.vga.Column_Counter.processQ[1]$_SDFFE_PN0P__391  (.L_HI(net391));
 sg13g2_tiehi \Pong.datapath.vga.Column_Counter.processQ[2]$_SDFFE_PN0P__392  (.L_HI(net392));
 sg13g2_tiehi \Pong.datapath.vga.Column_Counter.processQ[3]$_SDFFE_PN0P__393  (.L_HI(net393));
 sg13g2_tiehi \Pong.datapath.vga.Column_Counter.processQ[4]$_SDFFE_PN0P__394  (.L_HI(net394));
 sg13g2_tiehi \Pong.datapath.vga.Column_Counter.processQ[5]$_SDFFE_PN0P__395  (.L_HI(net395));
 sg13g2_tiehi \Pong.datapath.vga.Column_Counter.processQ[6]$_SDFFE_PN0P__396  (.L_HI(net396));
 sg13g2_tiehi \Pong.datapath.vga.Column_Counter.processQ[7]$_SDFFE_PN0P__397  (.L_HI(net397));
 sg13g2_tiehi \Pong.datapath.vga.Column_Counter.processQ[8]$_SDFFE_PN0P__398  (.L_HI(net398));
 sg13g2_tiehi \Pong.datapath.vga.Column_Counter.processQ[9]$_SDFFE_PN0P__399  (.L_HI(net399));
 sg13g2_tiehi \Pong.datapath.vga.Row_Counter.processQ[0]$_SDFFE_PN0P__400  (.L_HI(net400));
 sg13g2_tiehi \Pong.datapath.vga.Row_Counter.processQ[1]$_SDFFE_PN0P__401  (.L_HI(net401));
 sg13g2_tiehi \Pong.datapath.vga.Row_Counter.processQ[2]$_SDFFE_PN0P__402  (.L_HI(net402));
 sg13g2_tiehi \Pong.datapath.vga.Row_Counter.processQ[3]$_SDFFE_PN0P__403  (.L_HI(net403));
 sg13g2_tiehi \Pong.datapath.vga.Row_Counter.processQ[4]$_SDFFE_PN0P__404  (.L_HI(net404));
 sg13g2_tiehi \Pong.datapath.vga.Row_Counter.processQ[5]$_SDFFE_PN0P__405  (.L_HI(net405));
 sg13g2_tiehi \Pong.datapath.vga.Row_Counter.processQ[6]$_SDFFE_PN0P__406  (.L_HI(net406));
 sg13g2_tiehi \Pong.datapath.vga.Row_Counter.processQ[7]$_SDFFE_PN0P__407  (.L_HI(net407));
 sg13g2_tiehi \Pong.datapath.vga.Row_Counter.processQ[8]$_SDFFE_PN0P__408  (.L_HI(net408));
 sg13g2_tiehi \Pong.datapath.vga.Row_Counter.processQ[9]$_SDFFE_PN0P__409  (.L_HI(net409));
 sg13g2_tiehi _6190__410 (.L_HI(net410));
 sg13g2_tiehi _6191__411 (.L_HI(net411));
 sg13g2_tiehi _6193__412 (.L_HI(net412));
 sg13g2_tiehi _6194__413 (.L_HI(net413));
 sg13g2_buf_2 clkbuf_4_0_0_clk (.A(clknet_0_clk),
    .X(clknet_4_0_0_clk));
 sg13g2_buf_2 clkbuf_4_1_0_clk (.A(clknet_0_clk),
    .X(clknet_4_1_0_clk));
 sg13g2_buf_2 clkbuf_4_2_0_clk (.A(clknet_0_clk),
    .X(clknet_4_2_0_clk));
 sg13g2_buf_2 clkbuf_4_3_0_clk (.A(clknet_0_clk),
    .X(clknet_4_3_0_clk));
 sg13g2_buf_2 clkbuf_4_4_0_clk (.A(clknet_0_clk),
    .X(clknet_4_4_0_clk));
 sg13g2_buf_2 clkbuf_4_5_0_clk (.A(clknet_0_clk),
    .X(clknet_4_5_0_clk));
 sg13g2_buf_2 clkbuf_4_6_0_clk (.A(clknet_0_clk),
    .X(clknet_4_6_0_clk));
 sg13g2_buf_2 clkbuf_4_7_0_clk (.A(clknet_0_clk),
    .X(clknet_4_7_0_clk));
 sg13g2_buf_2 clkbuf_4_8_0_clk (.A(clknet_0_clk),
    .X(clknet_4_8_0_clk));
 sg13g2_buf_2 clkbuf_4_9_0_clk (.A(clknet_0_clk),
    .X(clknet_4_9_0_clk));
 sg13g2_buf_2 clkbuf_4_10_0_clk (.A(clknet_0_clk),
    .X(clknet_4_10_0_clk));
 sg13g2_buf_2 clkbuf_4_11_0_clk (.A(clknet_0_clk),
    .X(clknet_4_11_0_clk));
 sg13g2_buf_2 clkbuf_4_12_0_clk (.A(clknet_0_clk),
    .X(clknet_4_12_0_clk));
 sg13g2_buf_2 clkbuf_4_13_0_clk (.A(clknet_0_clk),
    .X(clknet_4_13_0_clk));
 sg13g2_buf_2 clkbuf_4_14_0_clk (.A(clknet_0_clk),
    .X(clknet_4_14_0_clk));
 sg13g2_buf_2 clkbuf_4_15_0_clk (.A(clknet_0_clk),
    .X(clknet_4_15_0_clk));
 sg13g2_buf_1 clkbuf_5_0__f_clk (.A(clknet_4_0_0_clk),
    .X(clknet_5_0__leaf_clk));
 sg13g2_buf_1 clkbuf_5_1__f_clk (.A(clknet_4_0_0_clk),
    .X(clknet_5_1__leaf_clk));
 sg13g2_buf_1 clkbuf_5_2__f_clk (.A(clknet_4_1_0_clk),
    .X(clknet_5_2__leaf_clk));
 sg13g2_buf_1 clkbuf_5_3__f_clk (.A(clknet_4_1_0_clk),
    .X(clknet_5_3__leaf_clk));
 sg13g2_buf_1 clkbuf_5_4__f_clk (.A(clknet_4_2_0_clk),
    .X(clknet_5_4__leaf_clk));
 sg13g2_buf_1 clkbuf_5_5__f_clk (.A(clknet_4_2_0_clk),
    .X(clknet_5_5__leaf_clk));
 sg13g2_buf_1 clkbuf_5_6__f_clk (.A(clknet_4_3_0_clk),
    .X(clknet_5_6__leaf_clk));
 sg13g2_buf_1 clkbuf_5_7__f_clk (.A(clknet_4_3_0_clk),
    .X(clknet_5_7__leaf_clk));
 sg13g2_buf_1 clkbuf_5_8__f_clk (.A(clknet_4_4_0_clk),
    .X(clknet_5_8__leaf_clk));
 sg13g2_buf_1 clkbuf_5_9__f_clk (.A(clknet_4_4_0_clk),
    .X(clknet_5_9__leaf_clk));
 sg13g2_buf_1 clkbuf_5_10__f_clk (.A(clknet_4_5_0_clk),
    .X(clknet_5_10__leaf_clk));
 sg13g2_buf_1 clkbuf_5_11__f_clk (.A(clknet_4_5_0_clk),
    .X(clknet_5_11__leaf_clk));
 sg13g2_buf_1 clkbuf_5_12__f_clk (.A(clknet_4_6_0_clk),
    .X(clknet_5_12__leaf_clk));
 sg13g2_buf_1 clkbuf_5_13__f_clk (.A(clknet_4_6_0_clk),
    .X(clknet_5_13__leaf_clk));
 sg13g2_buf_1 clkbuf_5_14__f_clk (.A(clknet_4_7_0_clk),
    .X(clknet_5_14__leaf_clk));
 sg13g2_buf_1 clkbuf_5_15__f_clk (.A(clknet_4_7_0_clk),
    .X(clknet_5_15__leaf_clk));
 sg13g2_buf_1 clkbuf_5_16__f_clk (.A(clknet_4_8_0_clk),
    .X(clknet_5_16__leaf_clk));
 sg13g2_buf_1 clkbuf_5_17__f_clk (.A(clknet_4_8_0_clk),
    .X(clknet_5_17__leaf_clk));
 sg13g2_buf_1 clkbuf_5_18__f_clk (.A(clknet_4_9_0_clk),
    .X(clknet_5_18__leaf_clk));
 sg13g2_buf_1 clkbuf_5_19__f_clk (.A(clknet_4_9_0_clk),
    .X(clknet_5_19__leaf_clk));
 sg13g2_buf_1 clkbuf_5_20__f_clk (.A(clknet_4_10_0_clk),
    .X(clknet_5_20__leaf_clk));
 sg13g2_buf_1 clkbuf_5_21__f_clk (.A(clknet_4_10_0_clk),
    .X(clknet_5_21__leaf_clk));
 sg13g2_buf_1 clkbuf_5_22__f_clk (.A(clknet_4_11_0_clk),
    .X(clknet_5_22__leaf_clk));
 sg13g2_buf_1 clkbuf_5_23__f_clk (.A(clknet_4_11_0_clk),
    .X(clknet_5_23__leaf_clk));
 sg13g2_buf_1 clkbuf_5_24__f_clk (.A(clknet_4_12_0_clk),
    .X(clknet_5_24__leaf_clk));
 sg13g2_buf_1 clkbuf_5_25__f_clk (.A(clknet_4_12_0_clk),
    .X(clknet_5_25__leaf_clk));
 sg13g2_buf_1 clkbuf_5_26__f_clk (.A(clknet_4_13_0_clk),
    .X(clknet_5_26__leaf_clk));
 sg13g2_buf_1 clkbuf_5_27__f_clk (.A(clknet_4_13_0_clk),
    .X(clknet_5_27__leaf_clk));
 sg13g2_buf_1 clkbuf_5_28__f_clk (.A(clknet_4_14_0_clk),
    .X(clknet_5_28__leaf_clk));
 sg13g2_buf_1 clkbuf_5_29__f_clk (.A(clknet_4_14_0_clk),
    .X(clknet_5_29__leaf_clk));
 sg13g2_buf_1 clkbuf_5_30__f_clk (.A(clknet_4_15_0_clk),
    .X(clknet_5_30__leaf_clk));
 sg13g2_buf_1 clkbuf_5_31__f_clk (.A(clknet_4_15_0_clk),
    .X(clknet_5_31__leaf_clk));
 sg13g2_inv_1 clkload0 (.A(clknet_5_1__leaf_clk));
 sg13g2_antennanp ANTENNA_1 (.A(_0045_));
 sg13g2_antennanp ANTENNA_2 (.A(clk));
 sg13g2_antennanp ANTENNA_3 (.A(clk));
 sg13g2_antennanp ANTENNA_4 (.A(_0045_));
 sg13g2_antennanp ANTENNA_5 (.A(clk));
 sg13g2_antennanp ANTENNA_6 (.A(clk));
 sg13g2_antennanp ANTENNA_7 (.A(clk));
 sg13g2_antennanp ANTENNA_8 (.A(clk));
 sg13g2_decap_8 FILLER_0_0 ();
 sg13g2_decap_8 FILLER_0_7 ();
 sg13g2_decap_8 FILLER_0_14 ();
 sg13g2_decap_8 FILLER_0_21 ();
 sg13g2_decap_8 FILLER_0_28 ();
 sg13g2_decap_8 FILLER_0_35 ();
 sg13g2_decap_8 FILLER_0_42 ();
 sg13g2_decap_8 FILLER_0_49 ();
 sg13g2_decap_8 FILLER_0_56 ();
 sg13g2_decap_8 FILLER_0_63 ();
 sg13g2_decap_8 FILLER_0_70 ();
 sg13g2_decap_8 FILLER_0_77 ();
 sg13g2_decap_8 FILLER_0_84 ();
 sg13g2_decap_8 FILLER_0_91 ();
 sg13g2_decap_8 FILLER_0_98 ();
 sg13g2_decap_8 FILLER_0_105 ();
 sg13g2_decap_8 FILLER_0_112 ();
 sg13g2_decap_8 FILLER_0_119 ();
 sg13g2_decap_8 FILLER_0_126 ();
 sg13g2_decap_8 FILLER_0_133 ();
 sg13g2_decap_8 FILLER_0_140 ();
 sg13g2_decap_8 FILLER_0_147 ();
 sg13g2_decap_8 FILLER_0_154 ();
 sg13g2_decap_8 FILLER_0_161 ();
 sg13g2_decap_8 FILLER_0_168 ();
 sg13g2_decap_8 FILLER_0_175 ();
 sg13g2_decap_8 FILLER_0_182 ();
 sg13g2_decap_8 FILLER_0_189 ();
 sg13g2_decap_8 FILLER_0_196 ();
 sg13g2_decap_8 FILLER_0_203 ();
 sg13g2_decap_8 FILLER_0_210 ();
 sg13g2_decap_8 FILLER_0_217 ();
 sg13g2_fill_2 FILLER_0_224 ();
 sg13g2_fill_1 FILLER_0_226 ();
 sg13g2_decap_8 FILLER_0_231 ();
 sg13g2_decap_8 FILLER_0_238 ();
 sg13g2_fill_1 FILLER_0_245 ();
 sg13g2_decap_8 FILLER_0_259 ();
 sg13g2_decap_8 FILLER_0_266 ();
 sg13g2_fill_1 FILLER_0_273 ();
 sg13g2_decap_8 FILLER_0_278 ();
 sg13g2_decap_8 FILLER_0_285 ();
 sg13g2_decap_8 FILLER_0_292 ();
 sg13g2_decap_8 FILLER_0_299 ();
 sg13g2_decap_8 FILLER_0_306 ();
 sg13g2_decap_8 FILLER_0_313 ();
 sg13g2_decap_8 FILLER_0_320 ();
 sg13g2_decap_8 FILLER_0_327 ();
 sg13g2_decap_8 FILLER_0_334 ();
 sg13g2_decap_8 FILLER_0_341 ();
 sg13g2_decap_8 FILLER_0_348 ();
 sg13g2_decap_8 FILLER_0_355 ();
 sg13g2_decap_8 FILLER_0_362 ();
 sg13g2_decap_8 FILLER_0_369 ();
 sg13g2_decap_8 FILLER_0_376 ();
 sg13g2_decap_8 FILLER_0_383 ();
 sg13g2_decap_8 FILLER_0_390 ();
 sg13g2_decap_8 FILLER_0_397 ();
 sg13g2_decap_8 FILLER_0_404 ();
 sg13g2_decap_8 FILLER_0_411 ();
 sg13g2_decap_8 FILLER_0_418 ();
 sg13g2_decap_4 FILLER_0_425 ();
 sg13g2_fill_1 FILLER_0_429 ();
 sg13g2_decap_8 FILLER_1_0 ();
 sg13g2_decap_8 FILLER_1_7 ();
 sg13g2_decap_8 FILLER_1_14 ();
 sg13g2_decap_8 FILLER_1_21 ();
 sg13g2_decap_8 FILLER_1_28 ();
 sg13g2_decap_8 FILLER_1_35 ();
 sg13g2_decap_8 FILLER_1_42 ();
 sg13g2_decap_8 FILLER_1_49 ();
 sg13g2_decap_8 FILLER_1_56 ();
 sg13g2_decap_8 FILLER_1_63 ();
 sg13g2_decap_8 FILLER_1_70 ();
 sg13g2_decap_8 FILLER_1_77 ();
 sg13g2_decap_8 FILLER_1_84 ();
 sg13g2_decap_8 FILLER_1_91 ();
 sg13g2_decap_8 FILLER_1_98 ();
 sg13g2_decap_8 FILLER_1_105 ();
 sg13g2_decap_8 FILLER_1_112 ();
 sg13g2_decap_8 FILLER_1_119 ();
 sg13g2_decap_8 FILLER_1_126 ();
 sg13g2_decap_8 FILLER_1_133 ();
 sg13g2_decap_8 FILLER_1_140 ();
 sg13g2_decap_8 FILLER_1_147 ();
 sg13g2_decap_8 FILLER_1_154 ();
 sg13g2_decap_8 FILLER_1_161 ();
 sg13g2_decap_8 FILLER_1_168 ();
 sg13g2_decap_8 FILLER_1_175 ();
 sg13g2_decap_8 FILLER_1_182 ();
 sg13g2_decap_8 FILLER_1_189 ();
 sg13g2_decap_8 FILLER_1_196 ();
 sg13g2_decap_4 FILLER_1_203 ();
 sg13g2_fill_2 FILLER_1_210 ();
 sg13g2_fill_2 FILLER_1_216 ();
 sg13g2_fill_1 FILLER_1_218 ();
 sg13g2_fill_1 FILLER_1_224 ();
 sg13g2_fill_1 FILLER_1_230 ();
 sg13g2_decap_4 FILLER_1_239 ();
 sg13g2_fill_2 FILLER_1_243 ();
 sg13g2_fill_2 FILLER_1_250 ();
 sg13g2_fill_2 FILLER_1_265 ();
 sg13g2_decap_8 FILLER_1_331 ();
 sg13g2_decap_8 FILLER_1_338 ();
 sg13g2_decap_8 FILLER_1_345 ();
 sg13g2_decap_8 FILLER_1_352 ();
 sg13g2_decap_8 FILLER_1_359 ();
 sg13g2_decap_8 FILLER_1_366 ();
 sg13g2_decap_8 FILLER_1_373 ();
 sg13g2_decap_8 FILLER_1_380 ();
 sg13g2_decap_8 FILLER_1_387 ();
 sg13g2_decap_8 FILLER_1_394 ();
 sg13g2_decap_8 FILLER_1_401 ();
 sg13g2_decap_8 FILLER_1_408 ();
 sg13g2_decap_8 FILLER_1_415 ();
 sg13g2_decap_8 FILLER_1_422 ();
 sg13g2_fill_1 FILLER_1_429 ();
 sg13g2_decap_8 FILLER_2_0 ();
 sg13g2_decap_8 FILLER_2_7 ();
 sg13g2_decap_8 FILLER_2_14 ();
 sg13g2_decap_8 FILLER_2_21 ();
 sg13g2_decap_8 FILLER_2_28 ();
 sg13g2_decap_8 FILLER_2_35 ();
 sg13g2_decap_8 FILLER_2_42 ();
 sg13g2_decap_8 FILLER_2_49 ();
 sg13g2_decap_8 FILLER_2_56 ();
 sg13g2_decap_8 FILLER_2_63 ();
 sg13g2_decap_8 FILLER_2_70 ();
 sg13g2_decap_8 FILLER_2_77 ();
 sg13g2_decap_8 FILLER_2_84 ();
 sg13g2_decap_8 FILLER_2_91 ();
 sg13g2_decap_8 FILLER_2_98 ();
 sg13g2_decap_8 FILLER_2_105 ();
 sg13g2_decap_8 FILLER_2_112 ();
 sg13g2_decap_8 FILLER_2_119 ();
 sg13g2_decap_8 FILLER_2_126 ();
 sg13g2_decap_8 FILLER_2_133 ();
 sg13g2_decap_8 FILLER_2_140 ();
 sg13g2_decap_8 FILLER_2_147 ();
 sg13g2_decap_8 FILLER_2_154 ();
 sg13g2_decap_8 FILLER_2_161 ();
 sg13g2_decap_8 FILLER_2_168 ();
 sg13g2_decap_8 FILLER_2_175 ();
 sg13g2_decap_8 FILLER_2_182 ();
 sg13g2_decap_8 FILLER_2_189 ();
 sg13g2_fill_1 FILLER_2_196 ();
 sg13g2_fill_2 FILLER_2_201 ();
 sg13g2_fill_1 FILLER_2_203 ();
 sg13g2_fill_1 FILLER_2_212 ();
 sg13g2_fill_2 FILLER_2_221 ();
 sg13g2_fill_2 FILLER_2_227 ();
 sg13g2_fill_2 FILLER_2_233 ();
 sg13g2_fill_1 FILLER_2_235 ();
 sg13g2_decap_4 FILLER_2_248 ();
 sg13g2_fill_2 FILLER_2_252 ();
 sg13g2_fill_1 FILLER_2_264 ();
 sg13g2_fill_1 FILLER_2_270 ();
 sg13g2_fill_1 FILLER_2_281 ();
 sg13g2_fill_2 FILLER_2_312 ();
 sg13g2_fill_1 FILLER_2_314 ();
 sg13g2_decap_8 FILLER_2_319 ();
 sg13g2_decap_8 FILLER_2_326 ();
 sg13g2_decap_8 FILLER_2_333 ();
 sg13g2_decap_8 FILLER_2_340 ();
 sg13g2_decap_8 FILLER_2_347 ();
 sg13g2_decap_8 FILLER_2_354 ();
 sg13g2_decap_8 FILLER_2_361 ();
 sg13g2_decap_8 FILLER_2_368 ();
 sg13g2_decap_8 FILLER_2_375 ();
 sg13g2_decap_8 FILLER_2_382 ();
 sg13g2_decap_8 FILLER_2_389 ();
 sg13g2_decap_8 FILLER_2_396 ();
 sg13g2_decap_8 FILLER_2_403 ();
 sg13g2_decap_8 FILLER_2_410 ();
 sg13g2_decap_8 FILLER_2_417 ();
 sg13g2_decap_4 FILLER_2_424 ();
 sg13g2_fill_2 FILLER_2_428 ();
 sg13g2_decap_8 FILLER_3_0 ();
 sg13g2_decap_8 FILLER_3_7 ();
 sg13g2_decap_8 FILLER_3_14 ();
 sg13g2_decap_8 FILLER_3_21 ();
 sg13g2_decap_8 FILLER_3_28 ();
 sg13g2_decap_8 FILLER_3_35 ();
 sg13g2_decap_8 FILLER_3_42 ();
 sg13g2_decap_8 FILLER_3_49 ();
 sg13g2_decap_8 FILLER_3_56 ();
 sg13g2_decap_8 FILLER_3_63 ();
 sg13g2_decap_8 FILLER_3_70 ();
 sg13g2_decap_8 FILLER_3_77 ();
 sg13g2_decap_8 FILLER_3_84 ();
 sg13g2_decap_8 FILLER_3_91 ();
 sg13g2_decap_8 FILLER_3_98 ();
 sg13g2_decap_8 FILLER_3_105 ();
 sg13g2_decap_8 FILLER_3_112 ();
 sg13g2_decap_8 FILLER_3_119 ();
 sg13g2_decap_8 FILLER_3_126 ();
 sg13g2_decap_8 FILLER_3_133 ();
 sg13g2_decap_8 FILLER_3_140 ();
 sg13g2_decap_8 FILLER_3_147 ();
 sg13g2_decap_8 FILLER_3_154 ();
 sg13g2_decap_8 FILLER_3_161 ();
 sg13g2_decap_8 FILLER_3_168 ();
 sg13g2_decap_8 FILLER_3_175 ();
 sg13g2_decap_4 FILLER_3_182 ();
 sg13g2_fill_2 FILLER_3_186 ();
 sg13g2_decap_4 FILLER_3_203 ();
 sg13g2_fill_2 FILLER_3_207 ();
 sg13g2_fill_1 FILLER_3_217 ();
 sg13g2_decap_4 FILLER_3_228 ();
 sg13g2_fill_1 FILLER_3_232 ();
 sg13g2_fill_2 FILLER_3_246 ();
 sg13g2_fill_1 FILLER_3_263 ();
 sg13g2_fill_2 FILLER_3_274 ();
 sg13g2_fill_1 FILLER_3_281 ();
 sg13g2_decap_8 FILLER_3_313 ();
 sg13g2_decap_8 FILLER_3_320 ();
 sg13g2_decap_8 FILLER_3_327 ();
 sg13g2_decap_4 FILLER_3_334 ();
 sg13g2_decap_8 FILLER_3_364 ();
 sg13g2_decap_8 FILLER_3_371 ();
 sg13g2_decap_8 FILLER_3_378 ();
 sg13g2_decap_8 FILLER_3_385 ();
 sg13g2_decap_8 FILLER_3_392 ();
 sg13g2_decap_8 FILLER_3_399 ();
 sg13g2_decap_8 FILLER_3_406 ();
 sg13g2_decap_8 FILLER_3_413 ();
 sg13g2_decap_8 FILLER_3_420 ();
 sg13g2_fill_2 FILLER_3_427 ();
 sg13g2_fill_1 FILLER_3_429 ();
 sg13g2_decap_8 FILLER_4_0 ();
 sg13g2_decap_8 FILLER_4_7 ();
 sg13g2_decap_8 FILLER_4_14 ();
 sg13g2_decap_8 FILLER_4_21 ();
 sg13g2_decap_8 FILLER_4_28 ();
 sg13g2_decap_8 FILLER_4_35 ();
 sg13g2_decap_8 FILLER_4_42 ();
 sg13g2_decap_8 FILLER_4_49 ();
 sg13g2_decap_8 FILLER_4_56 ();
 sg13g2_decap_8 FILLER_4_63 ();
 sg13g2_decap_8 FILLER_4_70 ();
 sg13g2_decap_8 FILLER_4_77 ();
 sg13g2_decap_8 FILLER_4_84 ();
 sg13g2_decap_8 FILLER_4_91 ();
 sg13g2_decap_8 FILLER_4_98 ();
 sg13g2_decap_8 FILLER_4_105 ();
 sg13g2_decap_8 FILLER_4_112 ();
 sg13g2_decap_8 FILLER_4_119 ();
 sg13g2_decap_8 FILLER_4_126 ();
 sg13g2_decap_8 FILLER_4_133 ();
 sg13g2_decap_8 FILLER_4_140 ();
 sg13g2_decap_8 FILLER_4_147 ();
 sg13g2_decap_8 FILLER_4_154 ();
 sg13g2_decap_8 FILLER_4_161 ();
 sg13g2_decap_8 FILLER_4_168 ();
 sg13g2_decap_8 FILLER_4_175 ();
 sg13g2_fill_2 FILLER_4_182 ();
 sg13g2_fill_1 FILLER_4_200 ();
 sg13g2_fill_1 FILLER_4_209 ();
 sg13g2_fill_1 FILLER_4_215 ();
 sg13g2_fill_2 FILLER_4_257 ();
 sg13g2_fill_1 FILLER_4_276 ();
 sg13g2_fill_2 FILLER_4_286 ();
 sg13g2_fill_1 FILLER_4_288 ();
 sg13g2_fill_2 FILLER_4_303 ();
 sg13g2_decap_8 FILLER_4_310 ();
 sg13g2_decap_8 FILLER_4_317 ();
 sg13g2_decap_8 FILLER_4_324 ();
 sg13g2_decap_8 FILLER_4_331 ();
 sg13g2_fill_2 FILLER_4_338 ();
 sg13g2_fill_1 FILLER_4_340 ();
 sg13g2_fill_2 FILLER_4_345 ();
 sg13g2_decap_4 FILLER_4_351 ();
 sg13g2_fill_2 FILLER_4_355 ();
 sg13g2_decap_8 FILLER_4_362 ();
 sg13g2_decap_8 FILLER_4_369 ();
 sg13g2_decap_8 FILLER_4_376 ();
 sg13g2_decap_8 FILLER_4_383 ();
 sg13g2_decap_8 FILLER_4_390 ();
 sg13g2_decap_8 FILLER_4_397 ();
 sg13g2_decap_8 FILLER_4_404 ();
 sg13g2_decap_8 FILLER_4_411 ();
 sg13g2_decap_8 FILLER_4_418 ();
 sg13g2_decap_4 FILLER_4_425 ();
 sg13g2_fill_1 FILLER_4_429 ();
 sg13g2_decap_8 FILLER_5_0 ();
 sg13g2_decap_8 FILLER_5_7 ();
 sg13g2_decap_8 FILLER_5_14 ();
 sg13g2_decap_8 FILLER_5_21 ();
 sg13g2_decap_8 FILLER_5_28 ();
 sg13g2_decap_8 FILLER_5_35 ();
 sg13g2_decap_8 FILLER_5_42 ();
 sg13g2_decap_8 FILLER_5_49 ();
 sg13g2_decap_8 FILLER_5_56 ();
 sg13g2_decap_8 FILLER_5_63 ();
 sg13g2_decap_8 FILLER_5_70 ();
 sg13g2_decap_8 FILLER_5_77 ();
 sg13g2_decap_8 FILLER_5_84 ();
 sg13g2_fill_2 FILLER_5_91 ();
 sg13g2_decap_8 FILLER_5_97 ();
 sg13g2_decap_8 FILLER_5_104 ();
 sg13g2_decap_4 FILLER_5_111 ();
 sg13g2_fill_1 FILLER_5_115 ();
 sg13g2_decap_8 FILLER_5_128 ();
 sg13g2_decap_8 FILLER_5_135 ();
 sg13g2_decap_8 FILLER_5_142 ();
 sg13g2_decap_8 FILLER_5_149 ();
 sg13g2_decap_8 FILLER_5_156 ();
 sg13g2_decap_8 FILLER_5_163 ();
 sg13g2_decap_8 FILLER_5_170 ();
 sg13g2_decap_8 FILLER_5_177 ();
 sg13g2_decap_8 FILLER_5_184 ();
 sg13g2_decap_4 FILLER_5_191 ();
 sg13g2_fill_1 FILLER_5_195 ();
 sg13g2_fill_1 FILLER_5_205 ();
 sg13g2_fill_1 FILLER_5_211 ();
 sg13g2_fill_1 FILLER_5_225 ();
 sg13g2_fill_1 FILLER_5_230 ();
 sg13g2_fill_1 FILLER_5_240 ();
 sg13g2_decap_8 FILLER_5_249 ();
 sg13g2_decap_8 FILLER_5_278 ();
 sg13g2_fill_2 FILLER_5_285 ();
 sg13g2_fill_1 FILLER_5_295 ();
 sg13g2_decap_8 FILLER_5_311 ();
 sg13g2_decap_8 FILLER_5_322 ();
 sg13g2_fill_1 FILLER_5_329 ();
 sg13g2_decap_8 FILLER_5_360 ();
 sg13g2_decap_8 FILLER_5_367 ();
 sg13g2_decap_8 FILLER_5_374 ();
 sg13g2_decap_8 FILLER_5_381 ();
 sg13g2_decap_8 FILLER_5_388 ();
 sg13g2_decap_8 FILLER_5_395 ();
 sg13g2_decap_8 FILLER_5_402 ();
 sg13g2_decap_8 FILLER_5_409 ();
 sg13g2_decap_8 FILLER_5_416 ();
 sg13g2_decap_8 FILLER_5_423 ();
 sg13g2_decap_8 FILLER_6_0 ();
 sg13g2_decap_8 FILLER_6_7 ();
 sg13g2_decap_8 FILLER_6_14 ();
 sg13g2_decap_8 FILLER_6_21 ();
 sg13g2_decap_8 FILLER_6_28 ();
 sg13g2_decap_8 FILLER_6_35 ();
 sg13g2_decap_8 FILLER_6_42 ();
 sg13g2_decap_8 FILLER_6_49 ();
 sg13g2_decap_8 FILLER_6_56 ();
 sg13g2_decap_8 FILLER_6_63 ();
 sg13g2_decap_8 FILLER_6_70 ();
 sg13g2_decap_8 FILLER_6_77 ();
 sg13g2_fill_2 FILLER_6_84 ();
 sg13g2_fill_2 FILLER_6_112 ();
 sg13g2_fill_1 FILLER_6_114 ();
 sg13g2_decap_8 FILLER_6_141 ();
 sg13g2_decap_8 FILLER_6_148 ();
 sg13g2_decap_8 FILLER_6_155 ();
 sg13g2_decap_8 FILLER_6_162 ();
 sg13g2_decap_8 FILLER_6_169 ();
 sg13g2_decap_8 FILLER_6_176 ();
 sg13g2_decap_4 FILLER_6_183 ();
 sg13g2_decap_8 FILLER_6_191 ();
 sg13g2_fill_1 FILLER_6_246 ();
 sg13g2_fill_1 FILLER_6_252 ();
 sg13g2_decap_8 FILLER_6_257 ();
 sg13g2_decap_4 FILLER_6_264 ();
 sg13g2_fill_2 FILLER_6_268 ();
 sg13g2_fill_1 FILLER_6_280 ();
 sg13g2_fill_2 FILLER_6_333 ();
 sg13g2_decap_8 FILLER_6_357 ();
 sg13g2_decap_8 FILLER_6_364 ();
 sg13g2_decap_8 FILLER_6_371 ();
 sg13g2_decap_8 FILLER_6_378 ();
 sg13g2_decap_8 FILLER_6_385 ();
 sg13g2_decap_8 FILLER_6_392 ();
 sg13g2_decap_8 FILLER_6_399 ();
 sg13g2_decap_8 FILLER_6_406 ();
 sg13g2_decap_8 FILLER_6_413 ();
 sg13g2_decap_8 FILLER_6_420 ();
 sg13g2_fill_2 FILLER_6_427 ();
 sg13g2_fill_1 FILLER_6_429 ();
 sg13g2_decap_8 FILLER_7_0 ();
 sg13g2_decap_8 FILLER_7_7 ();
 sg13g2_decap_8 FILLER_7_14 ();
 sg13g2_decap_8 FILLER_7_21 ();
 sg13g2_decap_8 FILLER_7_28 ();
 sg13g2_decap_8 FILLER_7_35 ();
 sg13g2_decap_8 FILLER_7_42 ();
 sg13g2_decap_8 FILLER_7_49 ();
 sg13g2_decap_8 FILLER_7_56 ();
 sg13g2_decap_8 FILLER_7_63 ();
 sg13g2_decap_8 FILLER_7_70 ();
 sg13g2_decap_8 FILLER_7_77 ();
 sg13g2_fill_1 FILLER_7_84 ();
 sg13g2_fill_2 FILLER_7_111 ();
 sg13g2_decap_4 FILLER_7_169 ();
 sg13g2_fill_2 FILLER_7_181 ();
 sg13g2_fill_1 FILLER_7_183 ();
 sg13g2_decap_8 FILLER_7_199 ();
 sg13g2_fill_2 FILLER_7_206 ();
 sg13g2_fill_1 FILLER_7_208 ();
 sg13g2_fill_1 FILLER_7_223 ();
 sg13g2_fill_2 FILLER_7_306 ();
 sg13g2_fill_1 FILLER_7_312 ();
 sg13g2_fill_1 FILLER_7_331 ();
 sg13g2_decap_8 FILLER_7_365 ();
 sg13g2_decap_8 FILLER_7_372 ();
 sg13g2_decap_8 FILLER_7_379 ();
 sg13g2_decap_8 FILLER_7_386 ();
 sg13g2_decap_8 FILLER_7_393 ();
 sg13g2_decap_8 FILLER_7_400 ();
 sg13g2_decap_8 FILLER_7_407 ();
 sg13g2_decap_8 FILLER_7_414 ();
 sg13g2_decap_8 FILLER_7_421 ();
 sg13g2_fill_2 FILLER_7_428 ();
 sg13g2_decap_8 FILLER_8_0 ();
 sg13g2_decap_8 FILLER_8_7 ();
 sg13g2_decap_8 FILLER_8_14 ();
 sg13g2_decap_8 FILLER_8_21 ();
 sg13g2_decap_8 FILLER_8_28 ();
 sg13g2_decap_8 FILLER_8_35 ();
 sg13g2_decap_8 FILLER_8_42 ();
 sg13g2_decap_8 FILLER_8_49 ();
 sg13g2_decap_8 FILLER_8_56 ();
 sg13g2_decap_4 FILLER_8_63 ();
 sg13g2_decap_8 FILLER_8_97 ();
 sg13g2_decap_4 FILLER_8_148 ();
 sg13g2_decap_8 FILLER_8_156 ();
 sg13g2_decap_8 FILLER_8_163 ();
 sg13g2_fill_2 FILLER_8_170 ();
 sg13g2_decap_4 FILLER_8_180 ();
 sg13g2_fill_2 FILLER_8_187 ();
 sg13g2_fill_1 FILLER_8_194 ();
 sg13g2_fill_1 FILLER_8_203 ();
 sg13g2_fill_1 FILLER_8_253 ();
 sg13g2_fill_2 FILLER_8_262 ();
 sg13g2_fill_2 FILLER_8_286 ();
 sg13g2_fill_2 FILLER_8_296 ();
 sg13g2_decap_4 FILLER_8_306 ();
 sg13g2_fill_2 FILLER_8_310 ();
 sg13g2_decap_4 FILLER_8_317 ();
 sg13g2_fill_1 FILLER_8_334 ();
 sg13g2_fill_1 FILLER_8_344 ();
 sg13g2_decap_8 FILLER_8_374 ();
 sg13g2_decap_8 FILLER_8_381 ();
 sg13g2_decap_8 FILLER_8_388 ();
 sg13g2_decap_8 FILLER_8_395 ();
 sg13g2_decap_8 FILLER_8_402 ();
 sg13g2_decap_8 FILLER_8_409 ();
 sg13g2_decap_8 FILLER_8_416 ();
 sg13g2_decap_8 FILLER_8_423 ();
 sg13g2_decap_8 FILLER_9_0 ();
 sg13g2_decap_8 FILLER_9_7 ();
 sg13g2_decap_8 FILLER_9_14 ();
 sg13g2_decap_8 FILLER_9_21 ();
 sg13g2_decap_8 FILLER_9_28 ();
 sg13g2_decap_8 FILLER_9_35 ();
 sg13g2_decap_8 FILLER_9_42 ();
 sg13g2_decap_8 FILLER_9_49 ();
 sg13g2_decap_8 FILLER_9_56 ();
 sg13g2_decap_8 FILLER_9_63 ();
 sg13g2_decap_4 FILLER_9_70 ();
 sg13g2_fill_2 FILLER_9_74 ();
 sg13g2_decap_4 FILLER_9_80 ();
 sg13g2_fill_1 FILLER_9_108 ();
 sg13g2_decap_8 FILLER_9_112 ();
 sg13g2_decap_4 FILLER_9_119 ();
 sg13g2_fill_2 FILLER_9_130 ();
 sg13g2_decap_4 FILLER_9_166 ();
 sg13g2_fill_2 FILLER_9_170 ();
 sg13g2_decap_4 FILLER_9_189 ();
 sg13g2_fill_2 FILLER_9_193 ();
 sg13g2_decap_4 FILLER_9_208 ();
 sg13g2_fill_1 FILLER_9_212 ();
 sg13g2_fill_2 FILLER_9_221 ();
 sg13g2_fill_1 FILLER_9_223 ();
 sg13g2_fill_1 FILLER_9_240 ();
 sg13g2_fill_1 FILLER_9_271 ();
 sg13g2_decap_4 FILLER_9_288 ();
 sg13g2_fill_2 FILLER_9_292 ();
 sg13g2_decap_8 FILLER_9_298 ();
 sg13g2_decap_8 FILLER_9_305 ();
 sg13g2_decap_4 FILLER_9_312 ();
 sg13g2_fill_2 FILLER_9_316 ();
 sg13g2_fill_2 FILLER_9_338 ();
 sg13g2_decap_8 FILLER_9_363 ();
 sg13g2_decap_8 FILLER_9_370 ();
 sg13g2_decap_8 FILLER_9_377 ();
 sg13g2_decap_8 FILLER_9_384 ();
 sg13g2_decap_8 FILLER_9_391 ();
 sg13g2_decap_8 FILLER_9_398 ();
 sg13g2_decap_8 FILLER_9_405 ();
 sg13g2_decap_8 FILLER_9_412 ();
 sg13g2_decap_8 FILLER_9_419 ();
 sg13g2_decap_4 FILLER_9_426 ();
 sg13g2_decap_8 FILLER_10_0 ();
 sg13g2_decap_8 FILLER_10_7 ();
 sg13g2_decap_8 FILLER_10_14 ();
 sg13g2_decap_8 FILLER_10_21 ();
 sg13g2_decap_8 FILLER_10_28 ();
 sg13g2_decap_8 FILLER_10_35 ();
 sg13g2_decap_8 FILLER_10_42 ();
 sg13g2_decap_8 FILLER_10_49 ();
 sg13g2_decap_8 FILLER_10_56 ();
 sg13g2_fill_2 FILLER_10_63 ();
 sg13g2_fill_2 FILLER_10_69 ();
 sg13g2_fill_1 FILLER_10_71 ();
 sg13g2_decap_4 FILLER_10_76 ();
 sg13g2_decap_8 FILLER_10_118 ();
 sg13g2_fill_1 FILLER_10_125 ();
 sg13g2_fill_1 FILLER_10_135 ();
 sg13g2_fill_2 FILLER_10_145 ();
 sg13g2_decap_8 FILLER_10_151 ();
 sg13g2_decap_8 FILLER_10_158 ();
 sg13g2_fill_2 FILLER_10_165 ();
 sg13g2_decap_4 FILLER_10_192 ();
 sg13g2_fill_1 FILLER_10_196 ();
 sg13g2_decap_8 FILLER_10_211 ();
 sg13g2_decap_4 FILLER_10_218 ();
 sg13g2_decap_8 FILLER_10_246 ();
 sg13g2_fill_1 FILLER_10_264 ();
 sg13g2_fill_2 FILLER_10_306 ();
 sg13g2_fill_1 FILLER_10_343 ();
 sg13g2_fill_2 FILLER_10_348 ();
 sg13g2_decap_8 FILLER_10_365 ();
 sg13g2_decap_8 FILLER_10_372 ();
 sg13g2_decap_8 FILLER_10_379 ();
 sg13g2_decap_8 FILLER_10_386 ();
 sg13g2_decap_8 FILLER_10_393 ();
 sg13g2_decap_8 FILLER_10_400 ();
 sg13g2_decap_8 FILLER_10_407 ();
 sg13g2_decap_8 FILLER_10_414 ();
 sg13g2_decap_8 FILLER_10_421 ();
 sg13g2_fill_2 FILLER_10_428 ();
 sg13g2_decap_8 FILLER_11_0 ();
 sg13g2_decap_8 FILLER_11_7 ();
 sg13g2_decap_8 FILLER_11_14 ();
 sg13g2_decap_8 FILLER_11_21 ();
 sg13g2_decap_8 FILLER_11_28 ();
 sg13g2_decap_8 FILLER_11_35 ();
 sg13g2_decap_8 FILLER_11_42 ();
 sg13g2_decap_8 FILLER_11_49 ();
 sg13g2_fill_2 FILLER_11_56 ();
 sg13g2_fill_1 FILLER_11_108 ();
 sg13g2_fill_1 FILLER_11_119 ();
 sg13g2_decap_8 FILLER_11_124 ();
 sg13g2_fill_1 FILLER_11_131 ();
 sg13g2_decap_8 FILLER_11_138 ();
 sg13g2_decap_8 FILLER_11_148 ();
 sg13g2_decap_8 FILLER_11_155 ();
 sg13g2_fill_2 FILLER_11_162 ();
 sg13g2_fill_1 FILLER_11_164 ();
 sg13g2_decap_8 FILLER_11_190 ();
 sg13g2_decap_4 FILLER_11_213 ();
 sg13g2_fill_2 FILLER_11_217 ();
 sg13g2_fill_2 FILLER_11_227 ();
 sg13g2_fill_1 FILLER_11_229 ();
 sg13g2_fill_1 FILLER_11_235 ();
 sg13g2_fill_2 FILLER_11_246 ();
 sg13g2_fill_1 FILLER_11_248 ();
 sg13g2_fill_2 FILLER_11_254 ();
 sg13g2_decap_8 FILLER_11_273 ();
 sg13g2_decap_8 FILLER_11_280 ();
 sg13g2_fill_2 FILLER_11_287 ();
 sg13g2_fill_2 FILLER_11_293 ();
 sg13g2_decap_8 FILLER_11_300 ();
 sg13g2_decap_8 FILLER_11_307 ();
 sg13g2_fill_1 FILLER_11_314 ();
 sg13g2_decap_8 FILLER_11_319 ();
 sg13g2_fill_1 FILLER_11_326 ();
 sg13g2_fill_1 FILLER_11_332 ();
 sg13g2_fill_1 FILLER_11_350 ();
 sg13g2_decap_8 FILLER_11_377 ();
 sg13g2_decap_8 FILLER_11_384 ();
 sg13g2_decap_8 FILLER_11_391 ();
 sg13g2_decap_8 FILLER_11_398 ();
 sg13g2_decap_8 FILLER_11_405 ();
 sg13g2_decap_8 FILLER_11_412 ();
 sg13g2_decap_8 FILLER_11_419 ();
 sg13g2_decap_4 FILLER_11_426 ();
 sg13g2_decap_8 FILLER_12_0 ();
 sg13g2_decap_8 FILLER_12_7 ();
 sg13g2_decap_8 FILLER_12_14 ();
 sg13g2_decap_8 FILLER_12_21 ();
 sg13g2_decap_8 FILLER_12_28 ();
 sg13g2_decap_8 FILLER_12_35 ();
 sg13g2_decap_8 FILLER_12_42 ();
 sg13g2_fill_1 FILLER_12_96 ();
 sg13g2_fill_1 FILLER_12_101 ();
 sg13g2_fill_1 FILLER_12_127 ();
 sg13g2_fill_2 FILLER_12_136 ();
 sg13g2_fill_2 FILLER_12_164 ();
 sg13g2_fill_1 FILLER_12_166 ();
 sg13g2_fill_1 FILLER_12_172 ();
 sg13g2_fill_1 FILLER_12_178 ();
 sg13g2_fill_1 FILLER_12_189 ();
 sg13g2_decap_4 FILLER_12_200 ();
 sg13g2_fill_2 FILLER_12_204 ();
 sg13g2_fill_1 FILLER_12_210 ();
 sg13g2_fill_1 FILLER_12_237 ();
 sg13g2_fill_1 FILLER_12_243 ();
 sg13g2_fill_1 FILLER_12_249 ();
 sg13g2_fill_1 FILLER_12_258 ();
 sg13g2_decap_8 FILLER_12_264 ();
 sg13g2_fill_2 FILLER_12_276 ();
 sg13g2_decap_8 FILLER_12_282 ();
 sg13g2_fill_1 FILLER_12_289 ();
 sg13g2_decap_8 FILLER_12_295 ();
 sg13g2_fill_2 FILLER_12_302 ();
 sg13g2_decap_4 FILLER_12_314 ();
 sg13g2_fill_1 FILLER_12_322 ();
 sg13g2_decap_8 FILLER_12_374 ();
 sg13g2_decap_8 FILLER_12_381 ();
 sg13g2_decap_8 FILLER_12_388 ();
 sg13g2_decap_8 FILLER_12_395 ();
 sg13g2_decap_8 FILLER_12_402 ();
 sg13g2_decap_8 FILLER_12_409 ();
 sg13g2_decap_8 FILLER_12_416 ();
 sg13g2_decap_8 FILLER_12_423 ();
 sg13g2_decap_8 FILLER_13_0 ();
 sg13g2_decap_8 FILLER_13_7 ();
 sg13g2_decap_8 FILLER_13_14 ();
 sg13g2_decap_8 FILLER_13_21 ();
 sg13g2_decap_8 FILLER_13_28 ();
 sg13g2_decap_8 FILLER_13_35 ();
 sg13g2_decap_8 FILLER_13_42 ();
 sg13g2_decap_8 FILLER_13_49 ();
 sg13g2_decap_4 FILLER_13_56 ();
 sg13g2_fill_1 FILLER_13_68 ();
 sg13g2_fill_1 FILLER_13_77 ();
 sg13g2_fill_1 FILLER_13_83 ();
 sg13g2_fill_1 FILLER_13_91 ();
 sg13g2_fill_2 FILLER_13_97 ();
 sg13g2_fill_1 FILLER_13_103 ();
 sg13g2_fill_2 FILLER_13_109 ();
 sg13g2_decap_4 FILLER_13_120 ();
 sg13g2_fill_2 FILLER_13_124 ();
 sg13g2_fill_2 FILLER_13_164 ();
 sg13g2_decap_8 FILLER_13_221 ();
 sg13g2_decap_4 FILLER_13_228 ();
 sg13g2_decap_4 FILLER_13_263 ();
 sg13g2_fill_2 FILLER_13_267 ();
 sg13g2_decap_4 FILLER_13_282 ();
 sg13g2_decap_4 FILLER_13_318 ();
 sg13g2_fill_1 FILLER_13_326 ();
 sg13g2_fill_2 FILLER_13_331 ();
 sg13g2_fill_2 FILLER_13_337 ();
 sg13g2_fill_2 FILLER_13_346 ();
 sg13g2_decap_8 FILLER_13_374 ();
 sg13g2_decap_8 FILLER_13_381 ();
 sg13g2_decap_8 FILLER_13_388 ();
 sg13g2_decap_8 FILLER_13_395 ();
 sg13g2_decap_8 FILLER_13_402 ();
 sg13g2_decap_8 FILLER_13_409 ();
 sg13g2_decap_8 FILLER_13_416 ();
 sg13g2_decap_8 FILLER_13_423 ();
 sg13g2_decap_8 FILLER_14_0 ();
 sg13g2_decap_8 FILLER_14_7 ();
 sg13g2_decap_8 FILLER_14_14 ();
 sg13g2_decap_8 FILLER_14_21 ();
 sg13g2_decap_8 FILLER_14_28 ();
 sg13g2_decap_8 FILLER_14_35 ();
 sg13g2_decap_8 FILLER_14_42 ();
 sg13g2_decap_8 FILLER_14_49 ();
 sg13g2_decap_8 FILLER_14_56 ();
 sg13g2_decap_8 FILLER_14_63 ();
 sg13g2_decap_8 FILLER_14_70 ();
 sg13g2_decap_8 FILLER_14_77 ();
 sg13g2_decap_8 FILLER_14_84 ();
 sg13g2_fill_2 FILLER_14_109 ();
 sg13g2_fill_1 FILLER_14_116 ();
 sg13g2_fill_2 FILLER_14_142 ();
 sg13g2_fill_2 FILLER_14_147 ();
 sg13g2_decap_8 FILLER_14_161 ();
 sg13g2_decap_8 FILLER_14_168 ();
 sg13g2_decap_4 FILLER_14_192 ();
 sg13g2_fill_1 FILLER_14_216 ();
 sg13g2_decap_4 FILLER_14_233 ();
 sg13g2_fill_2 FILLER_14_237 ();
 sg13g2_fill_1 FILLER_14_244 ();
 sg13g2_fill_2 FILLER_14_263 ();
 sg13g2_fill_1 FILLER_14_281 ();
 sg13g2_decap_4 FILLER_14_296 ();
 sg13g2_fill_1 FILLER_14_300 ();
 sg13g2_fill_2 FILLER_14_305 ();
 sg13g2_fill_1 FILLER_14_307 ();
 sg13g2_decap_8 FILLER_14_344 ();
 sg13g2_fill_2 FILLER_14_351 ();
 sg13g2_fill_2 FILLER_14_357 ();
 sg13g2_fill_1 FILLER_14_359 ();
 sg13g2_decap_8 FILLER_14_364 ();
 sg13g2_decap_8 FILLER_14_371 ();
 sg13g2_decap_8 FILLER_14_378 ();
 sg13g2_decap_8 FILLER_14_385 ();
 sg13g2_decap_8 FILLER_14_392 ();
 sg13g2_decap_8 FILLER_14_399 ();
 sg13g2_decap_8 FILLER_14_406 ();
 sg13g2_decap_8 FILLER_14_413 ();
 sg13g2_decap_8 FILLER_14_420 ();
 sg13g2_fill_2 FILLER_14_427 ();
 sg13g2_fill_1 FILLER_14_429 ();
 sg13g2_decap_8 FILLER_15_0 ();
 sg13g2_decap_8 FILLER_15_7 ();
 sg13g2_decap_8 FILLER_15_14 ();
 sg13g2_decap_8 FILLER_15_21 ();
 sg13g2_decap_8 FILLER_15_28 ();
 sg13g2_decap_8 FILLER_15_35 ();
 sg13g2_decap_8 FILLER_15_42 ();
 sg13g2_decap_8 FILLER_15_49 ();
 sg13g2_decap_8 FILLER_15_56 ();
 sg13g2_decap_8 FILLER_15_63 ();
 sg13g2_decap_8 FILLER_15_70 ();
 sg13g2_fill_1 FILLER_15_81 ();
 sg13g2_fill_2 FILLER_15_87 ();
 sg13g2_fill_2 FILLER_15_93 ();
 sg13g2_fill_1 FILLER_15_99 ();
 sg13g2_fill_1 FILLER_15_105 ();
 sg13g2_fill_2 FILLER_15_118 ();
 sg13g2_decap_4 FILLER_15_124 ();
 sg13g2_decap_4 FILLER_15_133 ();
 sg13g2_fill_2 FILLER_15_137 ();
 sg13g2_decap_8 FILLER_15_148 ();
 sg13g2_decap_8 FILLER_15_155 ();
 sg13g2_decap_4 FILLER_15_162 ();
 sg13g2_decap_8 FILLER_15_175 ();
 sg13g2_decap_8 FILLER_15_182 ();
 sg13g2_decap_8 FILLER_15_189 ();
 sg13g2_fill_1 FILLER_15_201 ();
 sg13g2_decap_4 FILLER_15_214 ();
 sg13g2_fill_1 FILLER_15_223 ();
 sg13g2_fill_1 FILLER_15_230 ();
 sg13g2_fill_1 FILLER_15_239 ();
 sg13g2_fill_2 FILLER_15_249 ();
 sg13g2_fill_2 FILLER_15_259 ();
 sg13g2_decap_8 FILLER_15_265 ();
 sg13g2_decap_8 FILLER_15_272 ();
 sg13g2_fill_1 FILLER_15_279 ();
 sg13g2_decap_8 FILLER_15_292 ();
 sg13g2_decap_8 FILLER_15_299 ();
 sg13g2_fill_1 FILLER_15_306 ();
 sg13g2_decap_8 FILLER_15_311 ();
 sg13g2_fill_2 FILLER_15_318 ();
 sg13g2_fill_1 FILLER_15_320 ();
 sg13g2_fill_2 FILLER_15_325 ();
 sg13g2_fill_1 FILLER_15_327 ();
 sg13g2_fill_1 FILLER_15_333 ();
 sg13g2_decap_8 FILLER_15_342 ();
 sg13g2_fill_1 FILLER_15_353 ();
 sg13g2_decap_8 FILLER_15_380 ();
 sg13g2_decap_8 FILLER_15_387 ();
 sg13g2_decap_8 FILLER_15_394 ();
 sg13g2_decap_8 FILLER_15_401 ();
 sg13g2_decap_8 FILLER_15_408 ();
 sg13g2_decap_8 FILLER_15_415 ();
 sg13g2_decap_8 FILLER_15_422 ();
 sg13g2_fill_1 FILLER_15_429 ();
 sg13g2_decap_8 FILLER_16_0 ();
 sg13g2_decap_8 FILLER_16_7 ();
 sg13g2_decap_8 FILLER_16_14 ();
 sg13g2_decap_8 FILLER_16_21 ();
 sg13g2_decap_8 FILLER_16_28 ();
 sg13g2_decap_8 FILLER_16_35 ();
 sg13g2_decap_8 FILLER_16_42 ();
 sg13g2_decap_8 FILLER_16_49 ();
 sg13g2_decap_8 FILLER_16_56 ();
 sg13g2_fill_1 FILLER_16_67 ();
 sg13g2_fill_1 FILLER_16_76 ();
 sg13g2_fill_1 FILLER_16_84 ();
 sg13g2_fill_2 FILLER_16_111 ();
 sg13g2_fill_1 FILLER_16_117 ();
 sg13g2_fill_2 FILLER_16_123 ();
 sg13g2_fill_1 FILLER_16_125 ();
 sg13g2_decap_8 FILLER_16_173 ();
 sg13g2_fill_1 FILLER_16_180 ();
 sg13g2_decap_4 FILLER_16_186 ();
 sg13g2_fill_1 FILLER_16_203 ();
 sg13g2_fill_1 FILLER_16_253 ();
 sg13g2_fill_2 FILLER_16_273 ();
 sg13g2_fill_2 FILLER_16_279 ();
 sg13g2_decap_4 FILLER_16_294 ();
 sg13g2_decap_8 FILLER_16_324 ();
 sg13g2_decap_4 FILLER_16_357 ();
 sg13g2_decap_8 FILLER_16_365 ();
 sg13g2_decap_4 FILLER_16_372 ();
 sg13g2_decap_8 FILLER_16_380 ();
 sg13g2_decap_8 FILLER_16_387 ();
 sg13g2_decap_8 FILLER_16_394 ();
 sg13g2_decap_8 FILLER_16_401 ();
 sg13g2_decap_8 FILLER_16_408 ();
 sg13g2_decap_8 FILLER_16_415 ();
 sg13g2_decap_8 FILLER_16_422 ();
 sg13g2_fill_1 FILLER_16_429 ();
 sg13g2_decap_8 FILLER_17_0 ();
 sg13g2_decap_8 FILLER_17_7 ();
 sg13g2_decap_8 FILLER_17_14 ();
 sg13g2_decap_8 FILLER_17_21 ();
 sg13g2_decap_8 FILLER_17_28 ();
 sg13g2_decap_8 FILLER_17_35 ();
 sg13g2_decap_8 FILLER_17_42 ();
 sg13g2_decap_8 FILLER_17_49 ();
 sg13g2_fill_1 FILLER_17_56 ();
 sg13g2_fill_2 FILLER_17_61 ();
 sg13g2_fill_1 FILLER_17_63 ();
 sg13g2_decap_8 FILLER_17_168 ();
 sg13g2_fill_1 FILLER_17_188 ();
 sg13g2_fill_2 FILLER_17_197 ();
 sg13g2_fill_1 FILLER_17_203 ();
 sg13g2_fill_1 FILLER_17_221 ();
 sg13g2_fill_2 FILLER_17_266 ();
 sg13g2_fill_2 FILLER_17_309 ();
 sg13g2_decap_8 FILLER_17_337 ();
 sg13g2_decap_8 FILLER_17_344 ();
 sg13g2_decap_4 FILLER_17_351 ();
 sg13g2_decap_8 FILLER_17_385 ();
 sg13g2_decap_8 FILLER_17_392 ();
 sg13g2_decap_8 FILLER_17_399 ();
 sg13g2_decap_8 FILLER_17_406 ();
 sg13g2_decap_8 FILLER_17_413 ();
 sg13g2_decap_8 FILLER_17_420 ();
 sg13g2_fill_2 FILLER_17_427 ();
 sg13g2_fill_1 FILLER_17_429 ();
 sg13g2_decap_8 FILLER_18_0 ();
 sg13g2_decap_8 FILLER_18_7 ();
 sg13g2_decap_8 FILLER_18_14 ();
 sg13g2_decap_8 FILLER_18_21 ();
 sg13g2_decap_8 FILLER_18_28 ();
 sg13g2_decap_8 FILLER_18_35 ();
 sg13g2_decap_8 FILLER_18_42 ();
 sg13g2_decap_8 FILLER_18_49 ();
 sg13g2_decap_4 FILLER_18_56 ();
 sg13g2_fill_1 FILLER_18_60 ();
 sg13g2_fill_2 FILLER_18_87 ();
 sg13g2_decap_4 FILLER_18_94 ();
 sg13g2_fill_2 FILLER_18_102 ();
 sg13g2_decap_4 FILLER_18_109 ();
 sg13g2_fill_1 FILLER_18_117 ();
 sg13g2_decap_4 FILLER_18_144 ();
 sg13g2_fill_2 FILLER_18_148 ();
 sg13g2_fill_2 FILLER_18_158 ();
 sg13g2_fill_1 FILLER_18_160 ();
 sg13g2_fill_1 FILLER_18_175 ();
 sg13g2_fill_2 FILLER_18_186 ();
 sg13g2_fill_1 FILLER_18_188 ();
 sg13g2_fill_2 FILLER_18_193 ();
 sg13g2_fill_2 FILLER_18_204 ();
 sg13g2_decap_8 FILLER_18_232 ();
 sg13g2_decap_4 FILLER_18_239 ();
 sg13g2_fill_1 FILLER_18_243 ();
 sg13g2_fill_1 FILLER_18_298 ();
 sg13g2_fill_2 FILLER_18_303 ();
 sg13g2_fill_1 FILLER_18_310 ();
 sg13g2_fill_2 FILLER_18_315 ();
 sg13g2_decap_8 FILLER_18_337 ();
 sg13g2_fill_2 FILLER_18_373 ();
 sg13g2_decap_8 FILLER_18_401 ();
 sg13g2_decap_8 FILLER_18_408 ();
 sg13g2_decap_8 FILLER_18_415 ();
 sg13g2_decap_8 FILLER_18_422 ();
 sg13g2_fill_1 FILLER_18_429 ();
 sg13g2_decap_8 FILLER_19_0 ();
 sg13g2_decap_8 FILLER_19_7 ();
 sg13g2_decap_8 FILLER_19_14 ();
 sg13g2_decap_8 FILLER_19_21 ();
 sg13g2_decap_8 FILLER_19_28 ();
 sg13g2_decap_8 FILLER_19_35 ();
 sg13g2_decap_8 FILLER_19_42 ();
 sg13g2_decap_8 FILLER_19_49 ();
 sg13g2_decap_4 FILLER_19_56 ();
 sg13g2_fill_2 FILLER_19_60 ();
 sg13g2_fill_2 FILLER_19_66 ();
 sg13g2_fill_1 FILLER_19_68 ();
 sg13g2_decap_8 FILLER_19_77 ();
 sg13g2_decap_8 FILLER_19_84 ();
 sg13g2_decap_8 FILLER_19_91 ();
 sg13g2_decap_8 FILLER_19_98 ();
 sg13g2_decap_8 FILLER_19_105 ();
 sg13g2_decap_8 FILLER_19_112 ();
 sg13g2_decap_4 FILLER_19_119 ();
 sg13g2_fill_1 FILLER_19_123 ();
 sg13g2_decap_8 FILLER_19_132 ();
 sg13g2_decap_8 FILLER_19_156 ();
 sg13g2_decap_8 FILLER_19_163 ();
 sg13g2_fill_1 FILLER_19_170 ();
 sg13g2_fill_1 FILLER_19_180 ();
 sg13g2_fill_1 FILLER_19_195 ();
 sg13g2_decap_8 FILLER_19_201 ();
 sg13g2_fill_2 FILLER_19_216 ();
 sg13g2_decap_8 FILLER_19_226 ();
 sg13g2_fill_2 FILLER_19_233 ();
 sg13g2_decap_8 FILLER_19_249 ();
 sg13g2_decap_8 FILLER_19_256 ();
 sg13g2_fill_2 FILLER_19_263 ();
 sg13g2_decap_8 FILLER_19_296 ();
 sg13g2_fill_2 FILLER_19_303 ();
 sg13g2_fill_1 FILLER_19_305 ();
 sg13g2_fill_1 FILLER_19_310 ();
 sg13g2_fill_2 FILLER_19_360 ();
 sg13g2_fill_1 FILLER_19_367 ();
 sg13g2_decap_8 FILLER_19_403 ();
 sg13g2_decap_8 FILLER_19_410 ();
 sg13g2_decap_8 FILLER_19_417 ();
 sg13g2_decap_4 FILLER_19_424 ();
 sg13g2_fill_2 FILLER_19_428 ();
 sg13g2_decap_8 FILLER_20_0 ();
 sg13g2_decap_8 FILLER_20_7 ();
 sg13g2_decap_8 FILLER_20_14 ();
 sg13g2_decap_8 FILLER_20_21 ();
 sg13g2_decap_4 FILLER_20_28 ();
 sg13g2_fill_2 FILLER_20_32 ();
 sg13g2_fill_1 FILLER_20_64 ();
 sg13g2_decap_8 FILLER_20_117 ();
 sg13g2_decap_8 FILLER_20_124 ();
 sg13g2_decap_8 FILLER_20_131 ();
 sg13g2_decap_8 FILLER_20_138 ();
 sg13g2_fill_2 FILLER_20_145 ();
 sg13g2_decap_8 FILLER_20_186 ();
 sg13g2_decap_4 FILLER_20_193 ();
 sg13g2_fill_2 FILLER_20_197 ();
 sg13g2_fill_2 FILLER_20_212 ();
 sg13g2_fill_2 FILLER_20_227 ();
 sg13g2_fill_1 FILLER_20_229 ();
 sg13g2_fill_2 FILLER_20_260 ();
 sg13g2_fill_1 FILLER_20_276 ();
 sg13g2_decap_4 FILLER_20_281 ();
 sg13g2_fill_2 FILLER_20_285 ();
 sg13g2_decap_4 FILLER_20_291 ();
 sg13g2_decap_4 FILLER_20_300 ();
 sg13g2_decap_8 FILLER_20_308 ();
 sg13g2_decap_8 FILLER_20_315 ();
 sg13g2_fill_1 FILLER_20_322 ();
 sg13g2_decap_8 FILLER_20_332 ();
 sg13g2_fill_2 FILLER_20_339 ();
 sg13g2_decap_4 FILLER_20_345 ();
 sg13g2_fill_1 FILLER_20_349 ();
 sg13g2_fill_2 FILLER_20_355 ();
 sg13g2_fill_2 FILLER_20_390 ();
 sg13g2_decap_8 FILLER_20_401 ();
 sg13g2_decap_8 FILLER_20_408 ();
 sg13g2_decap_8 FILLER_20_415 ();
 sg13g2_decap_8 FILLER_20_422 ();
 sg13g2_fill_1 FILLER_20_429 ();
 sg13g2_decap_8 FILLER_21_0 ();
 sg13g2_decap_8 FILLER_21_7 ();
 sg13g2_decap_8 FILLER_21_14 ();
 sg13g2_decap_8 FILLER_21_21 ();
 sg13g2_decap_8 FILLER_21_28 ();
 sg13g2_decap_8 FILLER_21_35 ();
 sg13g2_fill_1 FILLER_21_56 ();
 sg13g2_fill_1 FILLER_21_67 ();
 sg13g2_fill_1 FILLER_21_94 ();
 sg13g2_fill_1 FILLER_21_103 ();
 sg13g2_fill_2 FILLER_21_124 ();
 sg13g2_fill_1 FILLER_21_126 ();
 sg13g2_decap_4 FILLER_21_131 ();
 sg13g2_decap_8 FILLER_21_139 ();
 sg13g2_decap_4 FILLER_21_146 ();
 sg13g2_fill_1 FILLER_21_150 ();
 sg13g2_fill_2 FILLER_21_179 ();
 sg13g2_fill_1 FILLER_21_181 ();
 sg13g2_decap_8 FILLER_21_187 ();
 sg13g2_fill_1 FILLER_21_194 ();
 sg13g2_fill_2 FILLER_21_207 ();
 sg13g2_fill_1 FILLER_21_217 ();
 sg13g2_decap_8 FILLER_21_223 ();
 sg13g2_decap_8 FILLER_21_230 ();
 sg13g2_fill_1 FILLER_21_252 ();
 sg13g2_fill_2 FILLER_21_257 ();
 sg13g2_fill_1 FILLER_21_278 ();
 sg13g2_fill_1 FILLER_21_283 ();
 sg13g2_fill_2 FILLER_21_289 ();
 sg13g2_fill_2 FILLER_21_300 ();
 sg13g2_fill_1 FILLER_21_302 ();
 sg13g2_fill_1 FILLER_21_329 ();
 sg13g2_decap_8 FILLER_21_339 ();
 sg13g2_fill_2 FILLER_21_346 ();
 sg13g2_fill_1 FILLER_21_348 ();
 sg13g2_fill_2 FILLER_21_353 ();
 sg13g2_fill_1 FILLER_21_355 ();
 sg13g2_fill_1 FILLER_21_365 ();
 sg13g2_fill_2 FILLER_21_376 ();
 sg13g2_fill_1 FILLER_21_378 ();
 sg13g2_decap_8 FILLER_21_405 ();
 sg13g2_decap_8 FILLER_21_412 ();
 sg13g2_decap_8 FILLER_21_419 ();
 sg13g2_decap_4 FILLER_21_426 ();
 sg13g2_decap_8 FILLER_22_0 ();
 sg13g2_decap_8 FILLER_22_7 ();
 sg13g2_decap_8 FILLER_22_14 ();
 sg13g2_decap_8 FILLER_22_21 ();
 sg13g2_fill_2 FILLER_22_28 ();
 sg13g2_decap_4 FILLER_22_38 ();
 sg13g2_fill_2 FILLER_22_85 ();
 sg13g2_fill_1 FILLER_22_148 ();
 sg13g2_fill_2 FILLER_22_154 ();
 sg13g2_decap_8 FILLER_22_187 ();
 sg13g2_fill_2 FILLER_22_204 ();
 sg13g2_decap_8 FILLER_22_211 ();
 sg13g2_fill_2 FILLER_22_218 ();
 sg13g2_fill_2 FILLER_22_244 ();
 sg13g2_fill_1 FILLER_22_246 ();
 sg13g2_fill_1 FILLER_22_267 ();
 sg13g2_fill_2 FILLER_22_279 ();
 sg13g2_fill_1 FILLER_22_316 ();
 sg13g2_fill_1 FILLER_22_321 ();
 sg13g2_fill_1 FILLER_22_326 ();
 sg13g2_fill_2 FILLER_22_332 ();
 sg13g2_fill_2 FILLER_22_339 ();
 sg13g2_fill_1 FILLER_22_345 ();
 sg13g2_fill_1 FILLER_22_351 ();
 sg13g2_fill_1 FILLER_22_362 ();
 sg13g2_decap_4 FILLER_22_378 ();
 sg13g2_fill_2 FILLER_22_386 ();
 sg13g2_fill_2 FILLER_22_392 ();
 sg13g2_fill_2 FILLER_22_400 ();
 sg13g2_fill_1 FILLER_22_402 ();
 sg13g2_decap_8 FILLER_22_407 ();
 sg13g2_decap_8 FILLER_22_414 ();
 sg13g2_decap_8 FILLER_22_421 ();
 sg13g2_fill_2 FILLER_22_428 ();
 sg13g2_decap_8 FILLER_23_0 ();
 sg13g2_decap_8 FILLER_23_7 ();
 sg13g2_decap_8 FILLER_23_14 ();
 sg13g2_fill_2 FILLER_23_21 ();
 sg13g2_fill_2 FILLER_23_62 ();
 sg13g2_fill_2 FILLER_23_69 ();
 sg13g2_fill_1 FILLER_23_71 ();
 sg13g2_decap_8 FILLER_23_80 ();
 sg13g2_decap_4 FILLER_23_87 ();
 sg13g2_fill_1 FILLER_23_91 ();
 sg13g2_fill_2 FILLER_23_112 ();
 sg13g2_fill_2 FILLER_23_125 ();
 sg13g2_fill_1 FILLER_23_127 ();
 sg13g2_fill_2 FILLER_23_158 ();
 sg13g2_fill_1 FILLER_23_160 ();
 sg13g2_fill_2 FILLER_23_173 ();
 sg13g2_decap_8 FILLER_23_179 ();
 sg13g2_decap_4 FILLER_23_186 ();
 sg13g2_fill_2 FILLER_23_190 ();
 sg13g2_fill_1 FILLER_23_200 ();
 sg13g2_fill_1 FILLER_23_247 ();
 sg13g2_fill_2 FILLER_23_262 ();
 sg13g2_fill_1 FILLER_23_264 ();
 sg13g2_fill_1 FILLER_23_290 ();
 sg13g2_fill_1 FILLER_23_300 ();
 sg13g2_fill_1 FILLER_23_305 ();
 sg13g2_fill_1 FILLER_23_310 ();
 sg13g2_fill_1 FILLER_23_316 ();
 sg13g2_fill_2 FILLER_23_328 ();
 sg13g2_fill_1 FILLER_23_330 ();
 sg13g2_fill_1 FILLER_23_377 ();
 sg13g2_fill_2 FILLER_23_401 ();
 sg13g2_decap_8 FILLER_23_407 ();
 sg13g2_decap_8 FILLER_23_414 ();
 sg13g2_decap_8 FILLER_23_421 ();
 sg13g2_fill_2 FILLER_23_428 ();
 sg13g2_decap_8 FILLER_24_0 ();
 sg13g2_decap_8 FILLER_24_7 ();
 sg13g2_decap_8 FILLER_24_14 ();
 sg13g2_decap_4 FILLER_24_21 ();
 sg13g2_fill_1 FILLER_24_25 ();
 sg13g2_decap_8 FILLER_24_30 ();
 sg13g2_fill_1 FILLER_24_47 ();
 sg13g2_fill_1 FILLER_24_66 ();
 sg13g2_fill_1 FILLER_24_75 ();
 sg13g2_decap_8 FILLER_24_84 ();
 sg13g2_decap_8 FILLER_24_91 ();
 sg13g2_fill_2 FILLER_24_98 ();
 sg13g2_fill_1 FILLER_24_100 ();
 sg13g2_fill_2 FILLER_24_113 ();
 sg13g2_decap_8 FILLER_24_118 ();
 sg13g2_decap_8 FILLER_24_125 ();
 sg13g2_decap_4 FILLER_24_132 ();
 sg13g2_fill_1 FILLER_24_136 ();
 sg13g2_fill_2 FILLER_24_145 ();
 sg13g2_fill_2 FILLER_24_179 ();
 sg13g2_fill_2 FILLER_24_186 ();
 sg13g2_fill_1 FILLER_24_188 ();
 sg13g2_fill_2 FILLER_24_203 ();
 sg13g2_fill_1 FILLER_24_205 ();
 sg13g2_decap_8 FILLER_24_227 ();
 sg13g2_fill_2 FILLER_24_234 ();
 sg13g2_fill_1 FILLER_24_266 ();
 sg13g2_fill_1 FILLER_24_286 ();
 sg13g2_fill_1 FILLER_24_296 ();
 sg13g2_fill_1 FILLER_24_331 ();
 sg13g2_fill_1 FILLER_24_352 ();
 sg13g2_decap_4 FILLER_24_358 ();
 sg13g2_fill_2 FILLER_24_370 ();
 sg13g2_fill_1 FILLER_24_372 ();
 sg13g2_fill_2 FILLER_24_382 ();
 sg13g2_fill_1 FILLER_24_384 ();
 sg13g2_fill_2 FILLER_24_401 ();
 sg13g2_fill_1 FILLER_24_403 ();
 sg13g2_decap_8 FILLER_24_409 ();
 sg13g2_decap_8 FILLER_24_416 ();
 sg13g2_decap_8 FILLER_24_423 ();
 sg13g2_decap_8 FILLER_25_0 ();
 sg13g2_decap_8 FILLER_25_7 ();
 sg13g2_decap_4 FILLER_25_14 ();
 sg13g2_fill_1 FILLER_25_18 ();
 sg13g2_decap_4 FILLER_25_52 ();
 sg13g2_fill_2 FILLER_25_96 ();
 sg13g2_fill_1 FILLER_25_121 ();
 sg13g2_fill_2 FILLER_25_127 ();
 sg13g2_fill_1 FILLER_25_129 ();
 sg13g2_fill_1 FILLER_25_161 ();
 sg13g2_fill_2 FILLER_25_167 ();
 sg13g2_fill_2 FILLER_25_173 ();
 sg13g2_fill_1 FILLER_25_187 ();
 sg13g2_decap_4 FILLER_25_193 ();
 sg13g2_fill_2 FILLER_25_197 ();
 sg13g2_fill_1 FILLER_25_207 ();
 sg13g2_decap_4 FILLER_25_221 ();
 sg13g2_fill_1 FILLER_25_225 ();
 sg13g2_fill_1 FILLER_25_264 ();
 sg13g2_decap_8 FILLER_25_270 ();
 sg13g2_fill_2 FILLER_25_277 ();
 sg13g2_fill_1 FILLER_25_279 ();
 sg13g2_fill_2 FILLER_25_285 ();
 sg13g2_fill_1 FILLER_25_287 ();
 sg13g2_decap_8 FILLER_25_296 ();
 sg13g2_decap_4 FILLER_25_303 ();
 sg13g2_fill_1 FILLER_25_307 ();
 sg13g2_fill_2 FILLER_25_314 ();
 sg13g2_fill_2 FILLER_25_347 ();
 sg13g2_fill_1 FILLER_25_349 ();
 sg13g2_fill_1 FILLER_25_355 ();
 sg13g2_fill_2 FILLER_25_360 ();
 sg13g2_fill_1 FILLER_25_366 ();
 sg13g2_fill_1 FILLER_25_372 ();
 sg13g2_fill_1 FILLER_25_377 ();
 sg13g2_fill_2 FILLER_25_382 ();
 sg13g2_fill_2 FILLER_25_390 ();
 sg13g2_decap_8 FILLER_25_405 ();
 sg13g2_decap_8 FILLER_25_412 ();
 sg13g2_decap_8 FILLER_25_419 ();
 sg13g2_decap_4 FILLER_25_426 ();
 sg13g2_decap_8 FILLER_26_0 ();
 sg13g2_decap_8 FILLER_26_7 ();
 sg13g2_decap_8 FILLER_26_14 ();
 sg13g2_decap_8 FILLER_26_21 ();
 sg13g2_decap_4 FILLER_26_28 ();
 sg13g2_fill_2 FILLER_26_32 ();
 sg13g2_fill_2 FILLER_26_43 ();
 sg13g2_decap_8 FILLER_26_59 ();
 sg13g2_fill_1 FILLER_26_79 ();
 sg13g2_decap_4 FILLER_26_140 ();
 sg13g2_fill_2 FILLER_26_148 ();
 sg13g2_fill_1 FILLER_26_150 ();
 sg13g2_decap_4 FILLER_26_176 ();
 sg13g2_fill_2 FILLER_26_180 ();
 sg13g2_decap_4 FILLER_26_186 ();
 sg13g2_decap_4 FILLER_26_194 ();
 sg13g2_decap_4 FILLER_26_203 ();
 sg13g2_decap_4 FILLER_26_215 ();
 sg13g2_fill_1 FILLER_26_219 ();
 sg13g2_decap_8 FILLER_26_226 ();
 sg13g2_decap_8 FILLER_26_233 ();
 sg13g2_fill_1 FILLER_26_255 ();
 sg13g2_fill_1 FILLER_26_261 ();
 sg13g2_fill_1 FILLER_26_288 ();
 sg13g2_fill_2 FILLER_26_294 ();
 sg13g2_fill_1 FILLER_26_296 ();
 sg13g2_fill_1 FILLER_26_322 ();
 sg13g2_fill_1 FILLER_26_328 ();
 sg13g2_fill_1 FILLER_26_335 ();
 sg13g2_fill_1 FILLER_26_342 ();
 sg13g2_fill_1 FILLER_26_360 ();
 sg13g2_fill_2 FILLER_26_366 ();
 sg13g2_fill_2 FILLER_26_377 ();
 sg13g2_fill_2 FILLER_26_387 ();
 sg13g2_fill_2 FILLER_26_393 ();
 sg13g2_decap_8 FILLER_26_400 ();
 sg13g2_decap_8 FILLER_26_407 ();
 sg13g2_decap_8 FILLER_26_414 ();
 sg13g2_decap_8 FILLER_26_421 ();
 sg13g2_fill_2 FILLER_26_428 ();
 sg13g2_decap_8 FILLER_27_0 ();
 sg13g2_decap_8 FILLER_27_7 ();
 sg13g2_decap_8 FILLER_27_14 ();
 sg13g2_decap_8 FILLER_27_21 ();
 sg13g2_decap_4 FILLER_27_28 ();
 sg13g2_fill_2 FILLER_27_32 ();
 sg13g2_decap_8 FILLER_27_69 ();
 sg13g2_decap_8 FILLER_27_76 ();
 sg13g2_decap_4 FILLER_27_83 ();
 sg13g2_decap_8 FILLER_27_91 ();
 sg13g2_decap_4 FILLER_27_98 ();
 sg13g2_fill_2 FILLER_27_102 ();
 sg13g2_fill_2 FILLER_27_129 ();
 sg13g2_fill_1 FILLER_27_131 ();
 sg13g2_decap_4 FILLER_27_185 ();
 sg13g2_fill_1 FILLER_27_189 ();
 sg13g2_fill_2 FILLER_27_199 ();
 sg13g2_fill_1 FILLER_27_201 ();
 sg13g2_fill_2 FILLER_27_232 ();
 sg13g2_decap_8 FILLER_27_262 ();
 sg13g2_fill_2 FILLER_27_269 ();
 sg13g2_fill_2 FILLER_27_331 ();
 sg13g2_fill_1 FILLER_27_345 ();
 sg13g2_fill_1 FILLER_27_358 ();
 sg13g2_fill_1 FILLER_27_367 ();
 sg13g2_fill_1 FILLER_27_373 ();
 sg13g2_fill_1 FILLER_27_379 ();
 sg13g2_fill_1 FILLER_27_386 ();
 sg13g2_fill_2 FILLER_27_400 ();
 sg13g2_fill_1 FILLER_27_402 ();
 sg13g2_decap_8 FILLER_27_416 ();
 sg13g2_decap_8 FILLER_27_423 ();
 sg13g2_decap_8 FILLER_28_0 ();
 sg13g2_decap_8 FILLER_28_7 ();
 sg13g2_decap_8 FILLER_28_14 ();
 sg13g2_fill_2 FILLER_28_21 ();
 sg13g2_fill_1 FILLER_28_23 ();
 sg13g2_fill_1 FILLER_28_50 ();
 sg13g2_fill_1 FILLER_28_76 ();
 sg13g2_decap_8 FILLER_28_81 ();
 sg13g2_decap_8 FILLER_28_88 ();
 sg13g2_decap_8 FILLER_28_95 ();
 sg13g2_fill_1 FILLER_28_118 ();
 sg13g2_decap_8 FILLER_28_128 ();
 sg13g2_decap_8 FILLER_28_135 ();
 sg13g2_decap_4 FILLER_28_146 ();
 sg13g2_fill_1 FILLER_28_150 ();
 sg13g2_fill_1 FILLER_28_160 ();
 sg13g2_fill_1 FILLER_28_166 ();
 sg13g2_fill_1 FILLER_28_174 ();
 sg13g2_fill_2 FILLER_28_179 ();
 sg13g2_fill_1 FILLER_28_187 ();
 sg13g2_decap_4 FILLER_28_211 ();
 sg13g2_fill_1 FILLER_28_215 ();
 sg13g2_fill_1 FILLER_28_240 ();
 sg13g2_decap_8 FILLER_28_253 ();
 sg13g2_decap_8 FILLER_28_260 ();
 sg13g2_decap_8 FILLER_28_267 ();
 sg13g2_decap_8 FILLER_28_274 ();
 sg13g2_decap_4 FILLER_28_285 ();
 sg13g2_fill_1 FILLER_28_289 ();
 sg13g2_fill_2 FILLER_28_295 ();
 sg13g2_decap_8 FILLER_28_301 ();
 sg13g2_fill_2 FILLER_28_312 ();
 sg13g2_fill_2 FILLER_28_319 ();
 sg13g2_fill_2 FILLER_28_325 ();
 sg13g2_decap_4 FILLER_28_337 ();
 sg13g2_fill_2 FILLER_28_345 ();
 sg13g2_fill_1 FILLER_28_347 ();
 sg13g2_fill_2 FILLER_28_356 ();
 sg13g2_decap_8 FILLER_28_382 ();
 sg13g2_fill_2 FILLER_28_389 ();
 sg13g2_fill_1 FILLER_28_391 ();
 sg13g2_fill_1 FILLER_28_401 ();
 sg13g2_fill_1 FILLER_28_406 ();
 sg13g2_decap_4 FILLER_28_425 ();
 sg13g2_fill_1 FILLER_28_429 ();
 sg13g2_decap_8 FILLER_29_0 ();
 sg13g2_decap_8 FILLER_29_7 ();
 sg13g2_decap_8 FILLER_29_14 ();
 sg13g2_decap_8 FILLER_29_21 ();
 sg13g2_fill_2 FILLER_29_28 ();
 sg13g2_fill_1 FILLER_29_30 ();
 sg13g2_fill_1 FILLER_29_42 ();
 sg13g2_fill_1 FILLER_29_48 ();
 sg13g2_fill_2 FILLER_29_60 ();
 sg13g2_fill_2 FILLER_29_98 ();
 sg13g2_fill_1 FILLER_29_100 ();
 sg13g2_fill_2 FILLER_29_109 ();
 sg13g2_fill_1 FILLER_29_111 ();
 sg13g2_fill_1 FILLER_29_117 ();
 sg13g2_fill_1 FILLER_29_152 ();
 sg13g2_fill_2 FILLER_29_158 ();
 sg13g2_fill_1 FILLER_29_164 ();
 sg13g2_fill_2 FILLER_29_177 ();
 sg13g2_fill_1 FILLER_29_190 ();
 sg13g2_decap_4 FILLER_29_205 ();
 sg13g2_decap_8 FILLER_29_212 ();
 sg13g2_decap_8 FILLER_29_219 ();
 sg13g2_decap_4 FILLER_29_226 ();
 sg13g2_fill_1 FILLER_29_230 ();
 sg13g2_decap_8 FILLER_29_236 ();
 sg13g2_decap_4 FILLER_29_243 ();
 sg13g2_fill_2 FILLER_29_247 ();
 sg13g2_decap_8 FILLER_29_254 ();
 sg13g2_decap_8 FILLER_29_261 ();
 sg13g2_decap_8 FILLER_29_272 ();
 sg13g2_decap_8 FILLER_29_279 ();
 sg13g2_decap_8 FILLER_29_286 ();
 sg13g2_decap_4 FILLER_29_293 ();
 sg13g2_fill_2 FILLER_29_297 ();
 sg13g2_decap_8 FILLER_29_304 ();
 sg13g2_decap_8 FILLER_29_311 ();
 sg13g2_fill_2 FILLER_29_318 ();
 sg13g2_decap_8 FILLER_29_324 ();
 sg13g2_fill_1 FILLER_29_331 ();
 sg13g2_decap_4 FILLER_29_335 ();
 sg13g2_fill_1 FILLER_29_339 ();
 sg13g2_fill_1 FILLER_29_345 ();
 sg13g2_fill_2 FILLER_29_350 ();
 sg13g2_decap_8 FILLER_29_423 ();
 sg13g2_decap_8 FILLER_30_0 ();
 sg13g2_decap_8 FILLER_30_7 ();
 sg13g2_decap_8 FILLER_30_14 ();
 sg13g2_fill_2 FILLER_30_21 ();
 sg13g2_fill_1 FILLER_30_23 ();
 sg13g2_fill_1 FILLER_30_50 ();
 sg13g2_fill_1 FILLER_30_78 ();
 sg13g2_decap_4 FILLER_30_119 ();
 sg13g2_fill_1 FILLER_30_123 ();
 sg13g2_fill_2 FILLER_30_128 ();
 sg13g2_fill_1 FILLER_30_130 ();
 sg13g2_decap_4 FILLER_30_157 ();
 sg13g2_fill_1 FILLER_30_161 ();
 sg13g2_fill_2 FILLER_30_167 ();
 sg13g2_fill_1 FILLER_30_169 ();
 sg13g2_fill_1 FILLER_30_186 ();
 sg13g2_fill_2 FILLER_30_197 ();
 sg13g2_fill_1 FILLER_30_204 ();
 sg13g2_decap_8 FILLER_30_210 ();
 sg13g2_decap_8 FILLER_30_217 ();
 sg13g2_decap_8 FILLER_30_224 ();
 sg13g2_decap_8 FILLER_30_231 ();
 sg13g2_decap_8 FILLER_30_238 ();
 sg13g2_fill_2 FILLER_30_245 ();
 sg13g2_fill_2 FILLER_30_254 ();
 sg13g2_fill_1 FILLER_30_260 ();
 sg13g2_fill_1 FILLER_30_295 ();
 sg13g2_fill_2 FILLER_30_306 ();
 sg13g2_fill_1 FILLER_30_308 ();
 sg13g2_fill_2 FILLER_30_325 ();
 sg13g2_fill_2 FILLER_30_335 ();
 sg13g2_fill_1 FILLER_30_345 ();
 sg13g2_fill_2 FILLER_30_389 ();
 sg13g2_fill_2 FILLER_30_401 ();
 sg13g2_fill_1 FILLER_30_422 ();
 sg13g2_decap_8 FILLER_31_0 ();
 sg13g2_decap_8 FILLER_31_7 ();
 sg13g2_decap_8 FILLER_31_14 ();
 sg13g2_decap_8 FILLER_31_21 ();
 sg13g2_decap_4 FILLER_31_28 ();
 sg13g2_decap_4 FILLER_31_36 ();
 sg13g2_fill_1 FILLER_31_40 ();
 sg13g2_fill_1 FILLER_31_63 ();
 sg13g2_fill_1 FILLER_31_69 ();
 sg13g2_fill_2 FILLER_31_88 ();
 sg13g2_fill_2 FILLER_31_95 ();
 sg13g2_fill_1 FILLER_31_128 ();
 sg13g2_fill_1 FILLER_31_133 ();
 sg13g2_fill_2 FILLER_31_159 ();
 sg13g2_decap_4 FILLER_31_224 ();
 sg13g2_fill_1 FILLER_31_228 ();
 sg13g2_fill_2 FILLER_31_233 ();
 sg13g2_fill_1 FILLER_31_235 ();
 sg13g2_fill_1 FILLER_31_240 ();
 sg13g2_fill_1 FILLER_31_267 ();
 sg13g2_fill_1 FILLER_31_276 ();
 sg13g2_fill_1 FILLER_31_315 ();
 sg13g2_fill_2 FILLER_31_320 ();
 sg13g2_fill_1 FILLER_31_330 ();
 sg13g2_fill_1 FILLER_31_339 ();
 sg13g2_decap_8 FILLER_31_353 ();
 sg13g2_fill_1 FILLER_31_360 ();
 sg13g2_decap_8 FILLER_31_370 ();
 sg13g2_fill_1 FILLER_31_399 ();
 sg13g2_fill_1 FILLER_31_408 ();
 sg13g2_fill_1 FILLER_31_419 ();
 sg13g2_fill_2 FILLER_31_424 ();
 sg13g2_decap_8 FILLER_32_0 ();
 sg13g2_decap_8 FILLER_32_7 ();
 sg13g2_decap_8 FILLER_32_14 ();
 sg13g2_decap_8 FILLER_32_21 ();
 sg13g2_fill_2 FILLER_32_32 ();
 sg13g2_fill_1 FILLER_32_47 ();
 sg13g2_decap_8 FILLER_32_52 ();
 sg13g2_fill_1 FILLER_32_59 ();
 sg13g2_fill_1 FILLER_32_69 ();
 sg13g2_decap_8 FILLER_32_82 ();
 sg13g2_fill_2 FILLER_32_89 ();
 sg13g2_fill_2 FILLER_32_96 ();
 sg13g2_fill_1 FILLER_32_98 ();
 sg13g2_decap_4 FILLER_32_103 ();
 sg13g2_fill_2 FILLER_32_107 ();
 sg13g2_decap_4 FILLER_32_113 ();
 sg13g2_decap_8 FILLER_32_120 ();
 sg13g2_fill_2 FILLER_32_127 ();
 sg13g2_fill_1 FILLER_32_129 ();
 sg13g2_fill_1 FILLER_32_156 ();
 sg13g2_fill_1 FILLER_32_170 ();
 sg13g2_fill_1 FILLER_32_194 ();
 sg13g2_decap_4 FILLER_32_203 ();
 sg13g2_fill_2 FILLER_32_207 ();
 sg13g2_fill_2 FILLER_32_256 ();
 sg13g2_fill_1 FILLER_32_258 ();
 sg13g2_decap_4 FILLER_32_312 ();
 sg13g2_fill_1 FILLER_32_324 ();
 sg13g2_fill_1 FILLER_32_349 ();
 sg13g2_fill_1 FILLER_32_377 ();
 sg13g2_decap_8 FILLER_32_391 ();
 sg13g2_fill_1 FILLER_32_398 ();
 sg13g2_fill_2 FILLER_32_405 ();
 sg13g2_decap_8 FILLER_32_412 ();
 sg13g2_decap_4 FILLER_32_424 ();
 sg13g2_fill_2 FILLER_32_428 ();
 sg13g2_decap_8 FILLER_33_0 ();
 sg13g2_decap_8 FILLER_33_7 ();
 sg13g2_decap_8 FILLER_33_14 ();
 sg13g2_fill_1 FILLER_33_28 ();
 sg13g2_fill_1 FILLER_33_47 ();
 sg13g2_fill_2 FILLER_33_52 ();
 sg13g2_fill_1 FILLER_33_54 ();
 sg13g2_fill_1 FILLER_33_60 ();
 sg13g2_fill_1 FILLER_33_69 ();
 sg13g2_fill_2 FILLER_33_74 ();
 sg13g2_fill_2 FILLER_33_80 ();
 sg13g2_fill_1 FILLER_33_87 ();
 sg13g2_fill_2 FILLER_33_96 ();
 sg13g2_fill_1 FILLER_33_102 ();
 sg13g2_fill_2 FILLER_33_125 ();
 sg13g2_fill_1 FILLER_33_127 ();
 sg13g2_decap_4 FILLER_33_132 ();
 sg13g2_fill_1 FILLER_33_136 ();
 sg13g2_fill_1 FILLER_33_141 ();
 sg13g2_fill_2 FILLER_33_155 ();
 sg13g2_fill_1 FILLER_33_169 ();
 sg13g2_fill_1 FILLER_33_179 ();
 sg13g2_fill_2 FILLER_33_185 ();
 sg13g2_decap_8 FILLER_33_211 ();
 sg13g2_fill_2 FILLER_33_218 ();
 sg13g2_fill_1 FILLER_33_224 ();
 sg13g2_decap_4 FILLER_33_229 ();
 sg13g2_fill_1 FILLER_33_233 ();
 sg13g2_fill_1 FILLER_33_239 ();
 sg13g2_fill_1 FILLER_33_269 ();
 sg13g2_fill_2 FILLER_33_290 ();
 sg13g2_fill_1 FILLER_33_296 ();
 sg13g2_fill_2 FILLER_33_301 ();
 sg13g2_fill_1 FILLER_33_329 ();
 sg13g2_fill_2 FILLER_33_335 ();
 sg13g2_fill_1 FILLER_33_343 ();
 sg13g2_decap_4 FILLER_33_367 ();
 sg13g2_fill_1 FILLER_33_391 ();
 sg13g2_fill_1 FILLER_33_397 ();
 sg13g2_fill_2 FILLER_33_417 ();
 sg13g2_decap_4 FILLER_33_424 ();
 sg13g2_fill_2 FILLER_33_428 ();
 sg13g2_decap_4 FILLER_34_0 ();
 sg13g2_fill_1 FILLER_34_4 ();
 sg13g2_fill_2 FILLER_34_36 ();
 sg13g2_fill_1 FILLER_34_42 ();
 sg13g2_decap_4 FILLER_34_138 ();
 sg13g2_fill_1 FILLER_34_142 ();
 sg13g2_decap_8 FILLER_34_147 ();
 sg13g2_decap_4 FILLER_34_189 ();
 sg13g2_fill_2 FILLER_34_200 ();
 sg13g2_fill_1 FILLER_34_217 ();
 sg13g2_decap_8 FILLER_34_228 ();
 sg13g2_fill_1 FILLER_34_270 ();
 sg13g2_fill_1 FILLER_34_282 ();
 sg13g2_fill_2 FILLER_34_287 ();
 sg13g2_decap_8 FILLER_34_294 ();
 sg13g2_fill_1 FILLER_34_301 ();
 sg13g2_decap_4 FILLER_34_305 ();
 sg13g2_fill_1 FILLER_34_309 ();
 sg13g2_decap_8 FILLER_34_314 ();
 sg13g2_decap_8 FILLER_34_321 ();
 sg13g2_fill_2 FILLER_34_336 ();
 sg13g2_fill_1 FILLER_34_338 ();
 sg13g2_fill_1 FILLER_34_344 ();
 sg13g2_decap_4 FILLER_34_350 ();
 sg13g2_fill_2 FILLER_34_354 ();
 sg13g2_decap_4 FILLER_34_369 ();
 sg13g2_fill_2 FILLER_34_373 ();
 sg13g2_fill_2 FILLER_34_390 ();
 sg13g2_decap_4 FILLER_34_397 ();
 sg13g2_fill_1 FILLER_34_401 ();
 sg13g2_decap_8 FILLER_34_421 ();
 sg13g2_fill_2 FILLER_34_428 ();
 sg13g2_fill_1 FILLER_35_0 ();
 sg13g2_fill_2 FILLER_35_110 ();
 sg13g2_fill_1 FILLER_35_196 ();
 sg13g2_fill_2 FILLER_35_202 ();
 sg13g2_decap_8 FILLER_35_214 ();
 sg13g2_fill_2 FILLER_35_221 ();
 sg13g2_fill_1 FILLER_35_235 ();
 sg13g2_fill_1 FILLER_35_258 ();
 sg13g2_decap_4 FILLER_35_263 ();
 sg13g2_decap_8 FILLER_35_271 ();
 sg13g2_decap_4 FILLER_35_304 ();
 sg13g2_fill_2 FILLER_35_308 ();
 sg13g2_decap_8 FILLER_35_313 ();
 sg13g2_fill_1 FILLER_35_320 ();
 sg13g2_fill_2 FILLER_35_326 ();
 sg13g2_fill_1 FILLER_35_345 ();
 sg13g2_fill_1 FILLER_35_354 ();
 sg13g2_fill_1 FILLER_35_360 ();
 sg13g2_fill_1 FILLER_35_369 ();
 sg13g2_fill_1 FILLER_35_374 ();
 sg13g2_decap_4 FILLER_35_386 ();
 sg13g2_decap_8 FILLER_35_412 ();
 sg13g2_decap_8 FILLER_35_419 ();
 sg13g2_decap_4 FILLER_35_426 ();
 sg13g2_decap_8 FILLER_36_0 ();
 sg13g2_decap_8 FILLER_36_7 ();
 sg13g2_fill_2 FILLER_36_14 ();
 sg13g2_decap_4 FILLER_36_20 ();
 sg13g2_fill_1 FILLER_36_28 ();
 sg13g2_fill_2 FILLER_36_38 ();
 sg13g2_fill_1 FILLER_36_40 ();
 sg13g2_fill_2 FILLER_36_63 ();
 sg13g2_fill_2 FILLER_36_70 ();
 sg13g2_fill_1 FILLER_36_72 ();
 sg13g2_fill_2 FILLER_36_77 ();
 sg13g2_fill_1 FILLER_36_79 ();
 sg13g2_fill_2 FILLER_36_84 ();
 sg13g2_fill_1 FILLER_36_86 ();
 sg13g2_fill_1 FILLER_36_92 ();
 sg13g2_fill_1 FILLER_36_98 ();
 sg13g2_fill_2 FILLER_36_125 ();
 sg13g2_fill_1 FILLER_36_131 ();
 sg13g2_decap_4 FILLER_36_141 ();
 sg13g2_decap_8 FILLER_36_149 ();
 sg13g2_decap_8 FILLER_36_156 ();
 sg13g2_fill_1 FILLER_36_167 ();
 sg13g2_fill_2 FILLER_36_208 ();
 sg13g2_fill_1 FILLER_36_234 ();
 sg13g2_fill_1 FILLER_36_249 ();
 sg13g2_decap_8 FILLER_36_255 ();
 sg13g2_fill_1 FILLER_36_307 ();
 sg13g2_decap_8 FILLER_36_316 ();
 sg13g2_decap_8 FILLER_36_323 ();
 sg13g2_decap_8 FILLER_36_330 ();
 sg13g2_fill_2 FILLER_36_337 ();
 sg13g2_fill_1 FILLER_36_387 ();
 sg13g2_fill_2 FILLER_36_413 ();
 sg13g2_fill_2 FILLER_36_427 ();
 sg13g2_fill_1 FILLER_36_429 ();
 sg13g2_decap_8 FILLER_37_0 ();
 sg13g2_decap_8 FILLER_37_7 ();
 sg13g2_decap_8 FILLER_37_14 ();
 sg13g2_decap_8 FILLER_37_21 ();
 sg13g2_decap_8 FILLER_37_28 ();
 sg13g2_decap_8 FILLER_37_35 ();
 sg13g2_fill_2 FILLER_37_42 ();
 sg13g2_decap_4 FILLER_37_50 ();
 sg13g2_fill_2 FILLER_37_54 ();
 sg13g2_decap_8 FILLER_37_60 ();
 sg13g2_decap_8 FILLER_37_67 ();
 sg13g2_decap_8 FILLER_37_74 ();
 sg13g2_fill_1 FILLER_37_90 ();
 sg13g2_fill_1 FILLER_37_95 ();
 sg13g2_fill_2 FILLER_37_105 ();
 sg13g2_fill_1 FILLER_37_107 ();
 sg13g2_fill_1 FILLER_37_113 ();
 sg13g2_fill_2 FILLER_37_124 ();
 sg13g2_fill_1 FILLER_37_126 ();
 sg13g2_decap_8 FILLER_37_131 ();
 sg13g2_decap_8 FILLER_37_138 ();
 sg13g2_decap_8 FILLER_37_145 ();
 sg13g2_decap_8 FILLER_37_152 ();
 sg13g2_decap_8 FILLER_37_159 ();
 sg13g2_fill_1 FILLER_37_166 ();
 sg13g2_fill_2 FILLER_37_187 ();
 sg13g2_fill_1 FILLER_37_193 ();
 sg13g2_fill_1 FILLER_37_198 ();
 sg13g2_fill_1 FILLER_37_208 ();
 sg13g2_fill_1 FILLER_37_212 ();
 sg13g2_fill_2 FILLER_37_228 ();
 sg13g2_fill_1 FILLER_37_230 ();
 sg13g2_fill_1 FILLER_37_242 ();
 sg13g2_fill_1 FILLER_37_248 ();
 sg13g2_fill_1 FILLER_37_254 ();
 sg13g2_fill_2 FILLER_37_289 ();
 sg13g2_fill_1 FILLER_37_300 ();
 sg13g2_fill_1 FILLER_37_331 ();
 sg13g2_fill_1 FILLER_37_338 ();
 sg13g2_fill_1 FILLER_37_362 ();
 sg13g2_fill_2 FILLER_37_371 ();
 sg13g2_fill_1 FILLER_37_419 ();
 sg13g2_decap_4 FILLER_37_425 ();
 sg13g2_fill_1 FILLER_37_429 ();
 sg13g2_decap_8 FILLER_38_0 ();
 sg13g2_decap_8 FILLER_38_7 ();
 sg13g2_decap_8 FILLER_38_14 ();
 sg13g2_decap_8 FILLER_38_21 ();
 sg13g2_decap_8 FILLER_38_28 ();
 sg13g2_fill_1 FILLER_38_35 ();
 sg13g2_decap_8 FILLER_38_40 ();
 sg13g2_fill_2 FILLER_38_47 ();
 sg13g2_fill_1 FILLER_38_49 ();
 sg13g2_fill_2 FILLER_38_58 ();
 sg13g2_fill_1 FILLER_38_60 ();
 sg13g2_decap_8 FILLER_38_75 ();
 sg13g2_fill_1 FILLER_38_82 ();
 sg13g2_fill_1 FILLER_38_109 ();
 sg13g2_fill_1 FILLER_38_114 ();
 sg13g2_fill_1 FILLER_38_119 ();
 sg13g2_fill_1 FILLER_38_125 ();
 sg13g2_fill_1 FILLER_38_135 ();
 sg13g2_decap_8 FILLER_38_166 ();
 sg13g2_decap_8 FILLER_38_173 ();
 sg13g2_fill_1 FILLER_38_180 ();
 sg13g2_fill_1 FILLER_38_203 ();
 sg13g2_decap_8 FILLER_38_208 ();
 sg13g2_decap_4 FILLER_38_215 ();
 sg13g2_fill_1 FILLER_38_219 ();
 sg13g2_fill_1 FILLER_38_224 ();
 sg13g2_fill_1 FILLER_38_241 ();
 sg13g2_fill_2 FILLER_38_259 ();
 sg13g2_fill_2 FILLER_38_294 ();
 sg13g2_fill_1 FILLER_38_304 ();
 sg13g2_decap_4 FILLER_38_318 ();
 sg13g2_fill_2 FILLER_38_336 ();
 sg13g2_fill_2 FILLER_38_343 ();
 sg13g2_decap_4 FILLER_38_350 ();
 sg13g2_fill_1 FILLER_38_354 ();
 sg13g2_fill_2 FILLER_38_360 ();
 sg13g2_decap_4 FILLER_38_425 ();
 sg13g2_fill_1 FILLER_38_429 ();
 sg13g2_decap_8 FILLER_39_0 ();
 sg13g2_decap_8 FILLER_39_7 ();
 sg13g2_decap_4 FILLER_39_14 ();
 sg13g2_fill_1 FILLER_39_18 ();
 sg13g2_fill_2 FILLER_39_50 ();
 sg13g2_fill_1 FILLER_39_52 ();
 sg13g2_fill_1 FILLER_39_83 ();
 sg13g2_fill_2 FILLER_39_171 ();
 sg13g2_fill_1 FILLER_39_173 ();
 sg13g2_decap_4 FILLER_39_177 ();
 sg13g2_decap_8 FILLER_39_184 ();
 sg13g2_decap_8 FILLER_39_191 ();
 sg13g2_decap_8 FILLER_39_198 ();
 sg13g2_decap_8 FILLER_39_205 ();
 sg13g2_decap_8 FILLER_39_212 ();
 sg13g2_decap_8 FILLER_39_219 ();
 sg13g2_decap_4 FILLER_39_226 ();
 sg13g2_fill_1 FILLER_39_230 ();
 sg13g2_fill_1 FILLER_39_270 ();
 sg13g2_decap_8 FILLER_39_302 ();
 sg13g2_decap_4 FILLER_39_309 ();
 sg13g2_decap_4 FILLER_39_321 ();
 sg13g2_decap_8 FILLER_39_337 ();
 sg13g2_fill_2 FILLER_39_344 ();
 sg13g2_fill_1 FILLER_39_355 ();
 sg13g2_fill_1 FILLER_39_379 ();
 sg13g2_decap_8 FILLER_39_396 ();
 sg13g2_fill_2 FILLER_39_403 ();
 sg13g2_fill_1 FILLER_39_405 ();
 sg13g2_fill_1 FILLER_39_411 ();
 sg13g2_fill_1 FILLER_39_424 ();
 sg13g2_fill_2 FILLER_39_428 ();
 sg13g2_decap_8 FILLER_40_0 ();
 sg13g2_decap_8 FILLER_40_7 ();
 sg13g2_decap_8 FILLER_40_14 ();
 sg13g2_decap_4 FILLER_40_21 ();
 sg13g2_fill_1 FILLER_40_54 ();
 sg13g2_fill_1 FILLER_40_63 ();
 sg13g2_decap_4 FILLER_40_83 ();
 sg13g2_fill_1 FILLER_40_105 ();
 sg13g2_fill_1 FILLER_40_110 ();
 sg13g2_fill_2 FILLER_40_135 ();
 sg13g2_fill_1 FILLER_40_145 ();
 sg13g2_decap_4 FILLER_40_150 ();
 sg13g2_fill_2 FILLER_40_154 ();
 sg13g2_decap_8 FILLER_40_191 ();
 sg13g2_decap_4 FILLER_40_198 ();
 sg13g2_decap_8 FILLER_40_206 ();
 sg13g2_fill_2 FILLER_40_213 ();
 sg13g2_decap_8 FILLER_40_219 ();
 sg13g2_fill_1 FILLER_40_226 ();
 sg13g2_fill_1 FILLER_40_232 ();
 sg13g2_fill_1 FILLER_40_237 ();
 sg13g2_fill_2 FILLER_40_244 ();
 sg13g2_fill_2 FILLER_40_273 ();
 sg13g2_fill_2 FILLER_40_280 ();
 sg13g2_fill_1 FILLER_40_282 ();
 sg13g2_decap_4 FILLER_40_287 ();
 sg13g2_fill_2 FILLER_40_296 ();
 sg13g2_decap_8 FILLER_40_324 ();
 sg13g2_fill_2 FILLER_40_331 ();
 sg13g2_decap_4 FILLER_40_365 ();
 sg13g2_fill_1 FILLER_40_374 ();
 sg13g2_decap_8 FILLER_40_400 ();
 sg13g2_fill_2 FILLER_40_407 ();
 sg13g2_decap_4 FILLER_40_415 ();
 sg13g2_fill_2 FILLER_40_419 ();
 sg13g2_fill_1 FILLER_40_429 ();
 sg13g2_decap_8 FILLER_41_0 ();
 sg13g2_decap_8 FILLER_41_7 ();
 sg13g2_decap_8 FILLER_41_14 ();
 sg13g2_fill_2 FILLER_41_55 ();
 sg13g2_fill_1 FILLER_41_66 ();
 sg13g2_decap_4 FILLER_41_105 ();
 sg13g2_fill_1 FILLER_41_109 ();
 sg13g2_decap_8 FILLER_41_114 ();
 sg13g2_decap_8 FILLER_41_121 ();
 sg13g2_fill_2 FILLER_41_128 ();
 sg13g2_fill_1 FILLER_41_130 ();
 sg13g2_decap_8 FILLER_41_135 ();
 sg13g2_decap_8 FILLER_41_142 ();
 sg13g2_fill_2 FILLER_41_149 ();
 sg13g2_fill_1 FILLER_41_151 ();
 sg13g2_fill_1 FILLER_41_198 ();
 sg13g2_fill_2 FILLER_41_222 ();
 sg13g2_fill_1 FILLER_41_228 ();
 sg13g2_fill_2 FILLER_41_233 ();
 sg13g2_decap_8 FILLER_41_254 ();
 sg13g2_fill_2 FILLER_41_261 ();
 sg13g2_fill_2 FILLER_41_289 ();
 sg13g2_decap_4 FILLER_41_300 ();
 sg13g2_fill_2 FILLER_41_304 ();
 sg13g2_decap_8 FILLER_41_310 ();
 sg13g2_decap_4 FILLER_41_317 ();
 sg13g2_decap_8 FILLER_41_326 ();
 sg13g2_decap_4 FILLER_41_333 ();
 sg13g2_fill_2 FILLER_41_337 ();
 sg13g2_fill_2 FILLER_41_352 ();
 sg13g2_decap_8 FILLER_41_371 ();
 sg13g2_fill_1 FILLER_41_378 ();
 sg13g2_fill_1 FILLER_41_422 ();
 sg13g2_decap_8 FILLER_42_0 ();
 sg13g2_decap_8 FILLER_42_7 ();
 sg13g2_decap_8 FILLER_42_14 ();
 sg13g2_decap_8 FILLER_42_21 ();
 sg13g2_fill_2 FILLER_42_28 ();
 sg13g2_decap_8 FILLER_42_60 ();
 sg13g2_fill_1 FILLER_42_77 ();
 sg13g2_decap_8 FILLER_42_82 ();
 sg13g2_decap_8 FILLER_42_89 ();
 sg13g2_fill_1 FILLER_42_96 ();
 sg13g2_decap_8 FILLER_42_131 ();
 sg13g2_fill_1 FILLER_42_138 ();
 sg13g2_fill_1 FILLER_42_180 ();
 sg13g2_fill_1 FILLER_42_206 ();
 sg13g2_fill_1 FILLER_42_227 ();
 sg13g2_fill_1 FILLER_42_232 ();
 sg13g2_fill_1 FILLER_42_239 ();
 sg13g2_fill_1 FILLER_42_245 ();
 sg13g2_fill_1 FILLER_42_276 ();
 sg13g2_fill_2 FILLER_42_281 ();
 sg13g2_fill_2 FILLER_42_287 ();
 sg13g2_fill_2 FILLER_42_299 ();
 sg13g2_fill_1 FILLER_42_312 ();
 sg13g2_fill_2 FILLER_42_319 ();
 sg13g2_fill_1 FILLER_42_334 ();
 sg13g2_fill_2 FILLER_42_347 ();
 sg13g2_fill_1 FILLER_42_349 ();
 sg13g2_fill_1 FILLER_42_368 ();
 sg13g2_fill_1 FILLER_42_384 ();
 sg13g2_fill_1 FILLER_42_390 ();
 sg13g2_fill_1 FILLER_42_396 ();
 sg13g2_fill_1 FILLER_42_401 ();
 sg13g2_fill_1 FILLER_42_409 ();
 sg13g2_decap_8 FILLER_42_423 ();
 sg13g2_decap_8 FILLER_43_0 ();
 sg13g2_decap_8 FILLER_43_7 ();
 sg13g2_decap_8 FILLER_43_14 ();
 sg13g2_decap_8 FILLER_43_21 ();
 sg13g2_decap_8 FILLER_43_28 ();
 sg13g2_decap_8 FILLER_43_35 ();
 sg13g2_fill_2 FILLER_43_42 ();
 sg13g2_decap_8 FILLER_43_54 ();
 sg13g2_fill_2 FILLER_43_61 ();
 sg13g2_fill_1 FILLER_43_63 ();
 sg13g2_decap_4 FILLER_43_69 ();
 sg13g2_fill_1 FILLER_43_73 ();
 sg13g2_fill_1 FILLER_43_78 ();
 sg13g2_fill_2 FILLER_43_89 ();
 sg13g2_fill_2 FILLER_43_99 ();
 sg13g2_fill_1 FILLER_43_101 ();
 sg13g2_fill_1 FILLER_43_111 ();
 sg13g2_fill_1 FILLER_43_135 ();
 sg13g2_fill_2 FILLER_43_185 ();
 sg13g2_fill_2 FILLER_43_192 ();
 sg13g2_fill_2 FILLER_43_215 ();
 sg13g2_decap_4 FILLER_43_248 ();
 sg13g2_fill_1 FILLER_43_252 ();
 sg13g2_decap_8 FILLER_43_257 ();
 sg13g2_fill_1 FILLER_43_264 ();
 sg13g2_decap_8 FILLER_43_272 ();
 sg13g2_decap_8 FILLER_43_279 ();
 sg13g2_decap_8 FILLER_43_286 ();
 sg13g2_fill_2 FILLER_43_293 ();
 sg13g2_fill_1 FILLER_43_295 ();
 sg13g2_decap_8 FILLER_43_299 ();
 sg13g2_decap_8 FILLER_43_306 ();
 sg13g2_decap_4 FILLER_43_313 ();
 sg13g2_decap_4 FILLER_43_322 ();
 sg13g2_fill_1 FILLER_43_326 ();
 sg13g2_fill_2 FILLER_43_342 ();
 sg13g2_fill_1 FILLER_43_357 ();
 sg13g2_fill_1 FILLER_43_390 ();
 sg13g2_fill_1 FILLER_43_416 ();
 sg13g2_decap_8 FILLER_43_422 ();
 sg13g2_fill_1 FILLER_43_429 ();
 sg13g2_decap_8 FILLER_44_0 ();
 sg13g2_decap_8 FILLER_44_7 ();
 sg13g2_decap_8 FILLER_44_14 ();
 sg13g2_decap_8 FILLER_44_21 ();
 sg13g2_decap_4 FILLER_44_28 ();
 sg13g2_fill_1 FILLER_44_84 ();
 sg13g2_fill_2 FILLER_44_142 ();
 sg13g2_fill_1 FILLER_44_144 ();
 sg13g2_fill_1 FILLER_44_154 ();
 sg13g2_fill_1 FILLER_44_160 ();
 sg13g2_fill_2 FILLER_44_171 ();
 sg13g2_fill_1 FILLER_44_185 ();
 sg13g2_fill_2 FILLER_44_191 ();
 sg13g2_fill_2 FILLER_44_202 ();
 sg13g2_fill_2 FILLER_44_212 ();
 sg13g2_decap_8 FILLER_44_219 ();
 sg13g2_decap_4 FILLER_44_226 ();
 sg13g2_fill_1 FILLER_44_230 ();
 sg13g2_fill_1 FILLER_44_235 ();
 sg13g2_decap_8 FILLER_44_251 ();
 sg13g2_decap_8 FILLER_44_258 ();
 sg13g2_decap_4 FILLER_44_265 ();
 sg13g2_decap_4 FILLER_44_283 ();
 sg13g2_fill_1 FILLER_44_291 ();
 sg13g2_fill_1 FILLER_44_297 ();
 sg13g2_fill_1 FILLER_44_301 ();
 sg13g2_fill_1 FILLER_44_306 ();
 sg13g2_fill_2 FILLER_44_312 ();
 sg13g2_fill_2 FILLER_44_323 ();
 sg13g2_fill_2 FILLER_44_338 ();
 sg13g2_decap_4 FILLER_44_347 ();
 sg13g2_fill_2 FILLER_44_351 ();
 sg13g2_decap_4 FILLER_44_360 ();
 sg13g2_fill_1 FILLER_44_364 ();
 sg13g2_fill_1 FILLER_44_399 ();
 sg13g2_fill_1 FILLER_44_409 ();
 sg13g2_decap_8 FILLER_44_419 ();
 sg13g2_decap_4 FILLER_44_426 ();
 sg13g2_decap_8 FILLER_45_0 ();
 sg13g2_decap_8 FILLER_45_7 ();
 sg13g2_decap_8 FILLER_45_14 ();
 sg13g2_decap_8 FILLER_45_21 ();
 sg13g2_decap_8 FILLER_45_28 ();
 sg13g2_fill_2 FILLER_45_35 ();
 sg13g2_decap_8 FILLER_45_41 ();
 sg13g2_decap_4 FILLER_45_48 ();
 sg13g2_fill_2 FILLER_45_52 ();
 sg13g2_decap_4 FILLER_45_58 ();
 sg13g2_fill_2 FILLER_45_62 ();
 sg13g2_fill_1 FILLER_45_107 ();
 sg13g2_fill_1 FILLER_45_164 ();
 sg13g2_fill_2 FILLER_45_170 ();
 sg13g2_decap_8 FILLER_45_176 ();
 sg13g2_decap_4 FILLER_45_183 ();
 sg13g2_fill_2 FILLER_45_197 ();
 sg13g2_decap_8 FILLER_45_208 ();
 sg13g2_decap_8 FILLER_45_215 ();
 sg13g2_decap_8 FILLER_45_222 ();
 sg13g2_decap_8 FILLER_45_229 ();
 sg13g2_fill_2 FILLER_45_236 ();
 sg13g2_fill_1 FILLER_45_238 ();
 sg13g2_decap_8 FILLER_45_242 ();
 sg13g2_decap_8 FILLER_45_249 ();
 sg13g2_decap_8 FILLER_45_256 ();
 sg13g2_decap_4 FILLER_45_263 ();
 sg13g2_fill_1 FILLER_45_267 ();
 sg13g2_fill_2 FILLER_45_300 ();
 sg13g2_decap_8 FILLER_45_333 ();
 sg13g2_fill_2 FILLER_45_340 ();
 sg13g2_decap_8 FILLER_45_367 ();
 sg13g2_decap_8 FILLER_45_374 ();
 sg13g2_decap_8 FILLER_45_386 ();
 sg13g2_fill_2 FILLER_45_393 ();
 sg13g2_fill_1 FILLER_45_395 ();
 sg13g2_decap_8 FILLER_45_399 ();
 sg13g2_decap_4 FILLER_45_406 ();
 sg13g2_fill_1 FILLER_45_410 ();
 sg13g2_decap_8 FILLER_45_419 ();
 sg13g2_decap_4 FILLER_45_426 ();
 sg13g2_decap_8 FILLER_46_0 ();
 sg13g2_decap_8 FILLER_46_7 ();
 sg13g2_decap_8 FILLER_46_14 ();
 sg13g2_fill_2 FILLER_46_21 ();
 sg13g2_decap_8 FILLER_46_53 ();
 sg13g2_fill_2 FILLER_46_60 ();
 sg13g2_fill_1 FILLER_46_62 ();
 sg13g2_decap_8 FILLER_46_68 ();
 sg13g2_fill_2 FILLER_46_75 ();
 sg13g2_fill_1 FILLER_46_77 ();
 sg13g2_decap_8 FILLER_46_82 ();
 sg13g2_fill_2 FILLER_46_89 ();
 sg13g2_fill_2 FILLER_46_104 ();
 sg13g2_fill_1 FILLER_46_138 ();
 sg13g2_fill_2 FILLER_46_143 ();
 sg13g2_decap_4 FILLER_46_149 ();
 sg13g2_fill_2 FILLER_46_153 ();
 sg13g2_fill_1 FILLER_46_160 ();
 sg13g2_fill_2 FILLER_46_168 ();
 sg13g2_fill_2 FILLER_46_174 ();
 sg13g2_fill_1 FILLER_46_176 ();
 sg13g2_fill_1 FILLER_46_187 ();
 sg13g2_fill_1 FILLER_46_209 ();
 sg13g2_decap_8 FILLER_46_218 ();
 sg13g2_decap_8 FILLER_46_225 ();
 sg13g2_decap_4 FILLER_46_232 ();
 sg13g2_fill_2 FILLER_46_236 ();
 sg13g2_decap_4 FILLER_46_242 ();
 sg13g2_fill_1 FILLER_46_274 ();
 sg13g2_fill_1 FILLER_46_294 ();
 sg13g2_fill_1 FILLER_46_301 ();
 sg13g2_fill_1 FILLER_46_307 ();
 sg13g2_fill_2 FILLER_46_317 ();
 sg13g2_fill_2 FILLER_46_325 ();
 sg13g2_fill_1 FILLER_46_346 ();
 sg13g2_fill_2 FILLER_46_355 ();
 sg13g2_fill_1 FILLER_46_357 ();
 sg13g2_fill_1 FILLER_46_362 ();
 sg13g2_fill_2 FILLER_46_377 ();
 sg13g2_fill_1 FILLER_46_379 ();
 sg13g2_decap_8 FILLER_46_383 ();
 sg13g2_decap_8 FILLER_46_390 ();
 sg13g2_decap_8 FILLER_46_397 ();
 sg13g2_decap_8 FILLER_46_404 ();
 sg13g2_decap_8 FILLER_46_416 ();
 sg13g2_decap_8 FILLER_46_423 ();
 sg13g2_decap_8 FILLER_47_0 ();
 sg13g2_decap_8 FILLER_47_7 ();
 sg13g2_decap_4 FILLER_47_14 ();
 sg13g2_fill_2 FILLER_47_18 ();
 sg13g2_fill_1 FILLER_47_33 ();
 sg13g2_fill_1 FILLER_47_52 ();
 sg13g2_decap_8 FILLER_47_57 ();
 sg13g2_fill_2 FILLER_47_64 ();
 sg13g2_fill_1 FILLER_47_66 ();
 sg13g2_decap_4 FILLER_47_71 ();
 sg13g2_fill_2 FILLER_47_114 ();
 sg13g2_decap_8 FILLER_47_120 ();
 sg13g2_decap_8 FILLER_47_127 ();
 sg13g2_decap_8 FILLER_47_134 ();
 sg13g2_decap_8 FILLER_47_141 ();
 sg13g2_decap_8 FILLER_47_148 ();
 sg13g2_fill_2 FILLER_47_155 ();
 sg13g2_fill_1 FILLER_47_157 ();
 sg13g2_fill_1 FILLER_47_163 ();
 sg13g2_fill_1 FILLER_47_169 ();
 sg13g2_decap_8 FILLER_47_174 ();
 sg13g2_decap_8 FILLER_47_181 ();
 sg13g2_decap_4 FILLER_47_188 ();
 sg13g2_fill_1 FILLER_47_192 ();
 sg13g2_decap_8 FILLER_47_218 ();
 sg13g2_fill_1 FILLER_47_225 ();
 sg13g2_fill_1 FILLER_47_248 ();
 sg13g2_fill_2 FILLER_47_254 ();
 sg13g2_fill_2 FILLER_47_290 ();
 sg13g2_fill_1 FILLER_47_300 ();
 sg13g2_decap_4 FILLER_47_327 ();
 sg13g2_fill_2 FILLER_47_331 ();
 sg13g2_fill_2 FILLER_47_344 ();
 sg13g2_decap_8 FILLER_47_354 ();
 sg13g2_fill_1 FILLER_47_361 ();
 sg13g2_decap_8 FILLER_47_373 ();
 sg13g2_decap_4 FILLER_47_380 ();
 sg13g2_fill_2 FILLER_47_399 ();
 sg13g2_fill_2 FILLER_47_427 ();
 sg13g2_fill_1 FILLER_47_429 ();
 sg13g2_fill_1 FILLER_48_0 ();
 sg13g2_fill_1 FILLER_48_27 ();
 sg13g2_fill_2 FILLER_48_80 ();
 sg13g2_decap_4 FILLER_48_86 ();
 sg13g2_fill_1 FILLER_48_90 ();
 sg13g2_fill_1 FILLER_48_95 ();
 sg13g2_fill_1 FILLER_48_100 ();
 sg13g2_fill_1 FILLER_48_109 ();
 sg13g2_fill_2 FILLER_48_145 ();
 sg13g2_decap_8 FILLER_48_173 ();
 sg13g2_decap_8 FILLER_48_180 ();
 sg13g2_fill_2 FILLER_48_187 ();
 sg13g2_decap_4 FILLER_48_225 ();
 sg13g2_fill_2 FILLER_48_233 ();
 sg13g2_fill_1 FILLER_48_235 ();
 sg13g2_fill_1 FILLER_48_251 ();
 sg13g2_fill_2 FILLER_48_265 ();
 sg13g2_decap_4 FILLER_48_280 ();
 sg13g2_decap_8 FILLER_48_291 ();
 sg13g2_decap_8 FILLER_48_298 ();
 sg13g2_decap_4 FILLER_48_322 ();
 sg13g2_decap_4 FILLER_48_331 ();
 sg13g2_fill_2 FILLER_48_335 ();
 sg13g2_fill_2 FILLER_48_350 ();
 sg13g2_fill_2 FILLER_48_428 ();
 sg13g2_decap_8 FILLER_49_0 ();
 sg13g2_fill_2 FILLER_49_7 ();
 sg13g2_fill_1 FILLER_49_9 ();
 sg13g2_decap_4 FILLER_49_14 ();
 sg13g2_fill_1 FILLER_49_18 ();
 sg13g2_decap_4 FILLER_49_57 ();
 sg13g2_decap_8 FILLER_49_65 ();
 sg13g2_decap_4 FILLER_49_85 ();
 sg13g2_fill_1 FILLER_49_98 ();
 sg13g2_fill_1 FILLER_49_103 ();
 sg13g2_fill_1 FILLER_49_135 ();
 sg13g2_decap_8 FILLER_49_145 ();
 sg13g2_fill_1 FILLER_49_152 ();
 sg13g2_decap_8 FILLER_49_161 ();
 sg13g2_decap_4 FILLER_49_168 ();
 sg13g2_fill_1 FILLER_49_172 ();
 sg13g2_fill_1 FILLER_49_187 ();
 sg13g2_fill_1 FILLER_49_216 ();
 sg13g2_fill_1 FILLER_49_224 ();
 sg13g2_fill_2 FILLER_49_245 ();
 sg13g2_fill_1 FILLER_49_273 ();
 sg13g2_fill_1 FILLER_49_278 ();
 sg13g2_fill_1 FILLER_49_289 ();
 sg13g2_decap_4 FILLER_49_298 ();
 sg13g2_fill_1 FILLER_49_302 ();
 sg13g2_decap_4 FILLER_49_322 ();
 sg13g2_fill_2 FILLER_49_326 ();
 sg13g2_fill_1 FILLER_49_341 ();
 sg13g2_fill_1 FILLER_49_347 ();
 sg13g2_fill_1 FILLER_49_356 ();
 sg13g2_fill_1 FILLER_49_362 ();
 sg13g2_fill_2 FILLER_49_377 ();
 sg13g2_fill_1 FILLER_49_391 ();
 sg13g2_decap_8 FILLER_49_396 ();
 sg13g2_fill_2 FILLER_49_403 ();
 sg13g2_fill_1 FILLER_49_429 ();
 sg13g2_decap_8 FILLER_50_0 ();
 sg13g2_decap_8 FILLER_50_7 ();
 sg13g2_decap_4 FILLER_50_14 ();
 sg13g2_fill_1 FILLER_50_18 ();
 sg13g2_fill_2 FILLER_50_29 ();
 sg13g2_decap_4 FILLER_50_70 ();
 sg13g2_decap_4 FILLER_50_125 ();
 sg13g2_fill_2 FILLER_50_129 ();
 sg13g2_decap_8 FILLER_50_139 ();
 sg13g2_fill_1 FILLER_50_150 ();
 sg13g2_fill_2 FILLER_50_192 ();
 sg13g2_fill_1 FILLER_50_194 ();
 sg13g2_fill_1 FILLER_50_204 ();
 sg13g2_fill_1 FILLER_50_208 ();
 sg13g2_decap_8 FILLER_50_214 ();
 sg13g2_fill_2 FILLER_50_221 ();
 sg13g2_fill_2 FILLER_50_246 ();
 sg13g2_fill_1 FILLER_50_248 ();
 sg13g2_fill_1 FILLER_50_254 ();
 sg13g2_decap_4 FILLER_50_268 ();
 sg13g2_fill_2 FILLER_50_303 ();
 sg13g2_fill_2 FILLER_50_324 ();
 sg13g2_fill_1 FILLER_50_326 ();
 sg13g2_fill_2 FILLER_50_351 ();
 sg13g2_fill_2 FILLER_50_378 ();
 sg13g2_fill_1 FILLER_50_388 ();
 sg13g2_fill_1 FILLER_50_399 ();
 sg13g2_fill_1 FILLER_50_408 ();
 sg13g2_fill_2 FILLER_50_419 ();
 sg13g2_fill_1 FILLER_50_421 ();
 sg13g2_fill_1 FILLER_51_0 ();
 sg13g2_decap_4 FILLER_51_46 ();
 sg13g2_fill_2 FILLER_51_50 ();
 sg13g2_fill_2 FILLER_51_56 ();
 sg13g2_fill_1 FILLER_51_58 ();
 sg13g2_decap_8 FILLER_51_64 ();
 sg13g2_decap_8 FILLER_51_71 ();
 sg13g2_decap_8 FILLER_51_78 ();
 sg13g2_fill_2 FILLER_51_85 ();
 sg13g2_fill_1 FILLER_51_87 ();
 sg13g2_decap_4 FILLER_51_93 ();
 sg13g2_fill_1 FILLER_51_105 ();
 sg13g2_decap_8 FILLER_51_109 ();
 sg13g2_decap_4 FILLER_51_116 ();
 sg13g2_fill_1 FILLER_51_129 ();
 sg13g2_fill_2 FILLER_51_156 ();
 sg13g2_fill_2 FILLER_51_162 ();
 sg13g2_fill_2 FILLER_51_168 ();
 sg13g2_fill_1 FILLER_51_170 ();
 sg13g2_decap_8 FILLER_51_213 ();
 sg13g2_decap_4 FILLER_51_220 ();
 sg13g2_decap_4 FILLER_51_232 ();
 sg13g2_decap_4 FILLER_51_241 ();
 sg13g2_decap_4 FILLER_51_249 ();
 sg13g2_fill_2 FILLER_51_261 ();
 sg13g2_fill_2 FILLER_51_268 ();
 sg13g2_decap_4 FILLER_51_278 ();
 sg13g2_fill_1 FILLER_51_282 ();
 sg13g2_decap_8 FILLER_51_293 ();
 sg13g2_fill_1 FILLER_51_300 ();
 sg13g2_decap_4 FILLER_51_321 ();
 sg13g2_fill_2 FILLER_51_325 ();
 sg13g2_fill_2 FILLER_51_356 ();
 sg13g2_fill_1 FILLER_51_363 ();
 sg13g2_fill_2 FILLER_51_383 ();
 sg13g2_decap_4 FILLER_51_391 ();
 sg13g2_fill_2 FILLER_51_395 ();
 sg13g2_fill_2 FILLER_51_427 ();
 sg13g2_fill_1 FILLER_51_429 ();
 sg13g2_decap_8 FILLER_52_0 ();
 sg13g2_decap_8 FILLER_52_7 ();
 sg13g2_decap_8 FILLER_52_14 ();
 sg13g2_fill_1 FILLER_52_21 ();
 sg13g2_fill_2 FILLER_52_65 ();
 sg13g2_fill_2 FILLER_52_71 ();
 sg13g2_fill_1 FILLER_52_73 ();
 sg13g2_fill_1 FILLER_52_122 ();
 sg13g2_fill_1 FILLER_52_127 ();
 sg13g2_fill_1 FILLER_52_131 ();
 sg13g2_fill_2 FILLER_52_137 ();
 sg13g2_fill_2 FILLER_52_143 ();
 sg13g2_fill_1 FILLER_52_145 ();
 sg13g2_decap_8 FILLER_52_151 ();
 sg13g2_decap_8 FILLER_52_158 ();
 sg13g2_fill_1 FILLER_52_197 ();
 sg13g2_decap_8 FILLER_52_202 ();
 sg13g2_decap_8 FILLER_52_209 ();
 sg13g2_fill_2 FILLER_52_229 ();
 sg13g2_fill_2 FILLER_52_260 ();
 sg13g2_fill_1 FILLER_52_262 ();
 sg13g2_decap_8 FILLER_52_271 ();
 sg13g2_decap_4 FILLER_52_278 ();
 sg13g2_decap_8 FILLER_52_287 ();
 sg13g2_decap_8 FILLER_52_294 ();
 sg13g2_fill_2 FILLER_52_301 ();
 sg13g2_fill_1 FILLER_52_303 ();
 sg13g2_decap_8 FILLER_52_316 ();
 sg13g2_decap_8 FILLER_52_323 ();
 sg13g2_decap_8 FILLER_52_330 ();
 sg13g2_decap_4 FILLER_52_337 ();
 sg13g2_decap_8 FILLER_52_349 ();
 sg13g2_decap_8 FILLER_52_356 ();
 sg13g2_decap_8 FILLER_52_363 ();
 sg13g2_decap_8 FILLER_52_370 ();
 sg13g2_decap_8 FILLER_52_377 ();
 sg13g2_decap_8 FILLER_52_384 ();
 sg13g2_decap_8 FILLER_52_399 ();
 sg13g2_decap_8 FILLER_52_406 ();
 sg13g2_decap_8 FILLER_52_413 ();
 sg13g2_decap_8 FILLER_52_420 ();
 sg13g2_fill_2 FILLER_52_427 ();
 sg13g2_fill_1 FILLER_52_429 ();
 sg13g2_fill_1 FILLER_53_0 ();
 sg13g2_fill_2 FILLER_53_27 ();
 sg13g2_fill_1 FILLER_53_36 ();
 sg13g2_decap_8 FILLER_53_87 ();
 sg13g2_decap_4 FILLER_53_94 ();
 sg13g2_decap_8 FILLER_53_148 ();
 sg13g2_fill_1 FILLER_53_158 ();
 sg13g2_fill_1 FILLER_53_164 ();
 sg13g2_fill_1 FILLER_53_172 ();
 sg13g2_fill_1 FILLER_53_183 ();
 sg13g2_fill_2 FILLER_53_189 ();
 sg13g2_decap_4 FILLER_53_200 ();
 sg13g2_fill_1 FILLER_53_204 ();
 sg13g2_decap_8 FILLER_53_210 ();
 sg13g2_fill_2 FILLER_53_217 ();
 sg13g2_fill_1 FILLER_53_219 ();
 sg13g2_fill_1 FILLER_53_248 ();
 sg13g2_decap_4 FILLER_53_259 ();
 sg13g2_fill_1 FILLER_53_263 ();
 sg13g2_decap_8 FILLER_53_268 ();
 sg13g2_fill_2 FILLER_53_289 ();
 sg13g2_fill_1 FILLER_53_291 ();
 sg13g2_decap_8 FILLER_53_304 ();
 sg13g2_decap_4 FILLER_53_311 ();
 sg13g2_fill_1 FILLER_53_315 ();
 sg13g2_decap_8 FILLER_53_320 ();
 sg13g2_fill_2 FILLER_53_327 ();
 sg13g2_fill_1 FILLER_53_329 ();
 sg13g2_decap_8 FILLER_53_338 ();
 sg13g2_fill_1 FILLER_53_345 ();
 sg13g2_fill_2 FILLER_53_350 ();
 sg13g2_fill_1 FILLER_53_356 ();
 sg13g2_fill_2 FILLER_53_365 ();
 sg13g2_fill_1 FILLER_53_378 ();
 sg13g2_decap_4 FILLER_53_383 ();
 sg13g2_decap_8 FILLER_53_405 ();
 sg13g2_decap_8 FILLER_53_412 ();
 sg13g2_decap_8 FILLER_53_419 ();
 sg13g2_decap_4 FILLER_53_426 ();
 sg13g2_decap_8 FILLER_54_0 ();
 sg13g2_decap_8 FILLER_54_15 ();
 sg13g2_decap_4 FILLER_54_22 ();
 sg13g2_decap_4 FILLER_54_39 ();
 sg13g2_fill_1 FILLER_54_82 ();
 sg13g2_fill_1 FILLER_54_130 ();
 sg13g2_fill_1 FILLER_54_144 ();
 sg13g2_decap_8 FILLER_54_154 ();
 sg13g2_decap_8 FILLER_54_161 ();
 sg13g2_fill_2 FILLER_54_177 ();
 sg13g2_fill_1 FILLER_54_179 ();
 sg13g2_fill_1 FILLER_54_188 ();
 sg13g2_fill_1 FILLER_54_194 ();
 sg13g2_fill_1 FILLER_54_199 ();
 sg13g2_fill_2 FILLER_54_204 ();
 sg13g2_decap_8 FILLER_54_210 ();
 sg13g2_fill_1 FILLER_54_222 ();
 sg13g2_decap_8 FILLER_54_232 ();
 sg13g2_fill_2 FILLER_54_239 ();
 sg13g2_fill_1 FILLER_54_241 ();
 sg13g2_decap_8 FILLER_54_250 ();
 sg13g2_fill_2 FILLER_54_257 ();
 sg13g2_fill_1 FILLER_54_259 ();
 sg13g2_fill_2 FILLER_54_296 ();
 sg13g2_fill_2 FILLER_54_310 ();
 sg13g2_fill_1 FILLER_54_312 ();
 sg13g2_fill_1 FILLER_54_321 ();
 sg13g2_fill_2 FILLER_54_327 ();
 sg13g2_fill_1 FILLER_54_329 ();
 sg13g2_fill_2 FILLER_54_340 ();
 sg13g2_decap_8 FILLER_54_358 ();
 sg13g2_fill_2 FILLER_54_365 ();
 sg13g2_fill_1 FILLER_54_389 ();
 sg13g2_fill_1 FILLER_54_400 ();
 sg13g2_decap_8 FILLER_54_414 ();
 sg13g2_decap_8 FILLER_54_421 ();
 sg13g2_fill_2 FILLER_54_428 ();
 sg13g2_decap_8 FILLER_55_0 ();
 sg13g2_decap_8 FILLER_55_7 ();
 sg13g2_decap_8 FILLER_55_14 ();
 sg13g2_decap_8 FILLER_55_21 ();
 sg13g2_decap_8 FILLER_55_28 ();
 sg13g2_decap_8 FILLER_55_35 ();
 sg13g2_decap_4 FILLER_55_42 ();
 sg13g2_fill_2 FILLER_55_46 ();
 sg13g2_decap_4 FILLER_55_72 ();
 sg13g2_fill_2 FILLER_55_81 ();
 sg13g2_fill_1 FILLER_55_83 ();
 sg13g2_decap_4 FILLER_55_88 ();
 sg13g2_decap_4 FILLER_55_96 ();
 sg13g2_fill_2 FILLER_55_100 ();
 sg13g2_fill_2 FILLER_55_124 ();
 sg13g2_fill_1 FILLER_55_130 ();
 sg13g2_fill_1 FILLER_55_136 ();
 sg13g2_fill_1 FILLER_55_159 ();
 sg13g2_decap_8 FILLER_55_164 ();
 sg13g2_decap_4 FILLER_55_171 ();
 sg13g2_fill_2 FILLER_55_175 ();
 sg13g2_fill_1 FILLER_55_207 ();
 sg13g2_fill_1 FILLER_55_214 ();
 sg13g2_fill_1 FILLER_55_229 ();
 sg13g2_fill_2 FILLER_55_238 ();
 sg13g2_decap_4 FILLER_55_249 ();
 sg13g2_fill_2 FILLER_55_253 ();
 sg13g2_fill_2 FILLER_55_289 ();
 sg13g2_fill_1 FILLER_55_296 ();
 sg13g2_fill_2 FILLER_55_302 ();
 sg13g2_fill_2 FILLER_55_308 ();
 sg13g2_fill_1 FILLER_55_310 ();
 sg13g2_fill_1 FILLER_55_328 ();
 sg13g2_fill_1 FILLER_55_345 ();
 sg13g2_fill_1 FILLER_55_351 ();
 sg13g2_fill_1 FILLER_55_360 ();
 sg13g2_fill_2 FILLER_55_403 ();
 sg13g2_fill_1 FILLER_55_420 ();
 sg13g2_decap_4 FILLER_55_424 ();
 sg13g2_fill_2 FILLER_55_428 ();
 sg13g2_decap_8 FILLER_56_0 ();
 sg13g2_decap_4 FILLER_56_7 ();
 sg13g2_decap_4 FILLER_56_15 ();
 sg13g2_fill_2 FILLER_56_28 ();
 sg13g2_fill_2 FILLER_56_42 ();
 sg13g2_fill_1 FILLER_56_44 ();
 sg13g2_decap_8 FILLER_56_63 ();
 sg13g2_decap_8 FILLER_56_70 ();
 sg13g2_decap_8 FILLER_56_77 ();
 sg13g2_decap_8 FILLER_56_84 ();
 sg13g2_decap_8 FILLER_56_91 ();
 sg13g2_decap_4 FILLER_56_98 ();
 sg13g2_fill_1 FILLER_56_128 ();
 sg13g2_fill_1 FILLER_56_136 ();
 sg13g2_decap_4 FILLER_56_166 ();
 sg13g2_fill_1 FILLER_56_170 ();
 sg13g2_fill_2 FILLER_56_215 ();
 sg13g2_fill_1 FILLER_56_217 ();
 sg13g2_fill_2 FILLER_56_228 ();
 sg13g2_fill_1 FILLER_56_235 ();
 sg13g2_fill_2 FILLER_56_251 ();
 sg13g2_decap_8 FILLER_56_258 ();
 sg13g2_decap_8 FILLER_56_265 ();
 sg13g2_decap_8 FILLER_56_272 ();
 sg13g2_decap_4 FILLER_56_279 ();
 sg13g2_fill_1 FILLER_56_283 ();
 sg13g2_fill_1 FILLER_56_348 ();
 sg13g2_fill_2 FILLER_56_374 ();
 sg13g2_fill_1 FILLER_56_376 ();
 sg13g2_decap_4 FILLER_56_407 ();
 sg13g2_decap_4 FILLER_57_0 ();
 sg13g2_fill_2 FILLER_57_4 ();
 sg13g2_fill_2 FILLER_57_41 ();
 sg13g2_fill_1 FILLER_57_43 ();
 sg13g2_decap_8 FILLER_57_62 ();
 sg13g2_decap_8 FILLER_57_69 ();
 sg13g2_fill_1 FILLER_57_76 ();
 sg13g2_decap_4 FILLER_57_103 ();
 sg13g2_fill_1 FILLER_57_107 ();
 sg13g2_decap_8 FILLER_57_112 ();
 sg13g2_decap_8 FILLER_57_119 ();
 sg13g2_fill_1 FILLER_57_126 ();
 sg13g2_fill_1 FILLER_57_153 ();
 sg13g2_decap_8 FILLER_57_196 ();
 sg13g2_decap_4 FILLER_57_203 ();
 sg13g2_decap_8 FILLER_57_247 ();
 sg13g2_fill_2 FILLER_57_254 ();
 sg13g2_fill_1 FILLER_57_256 ();
 sg13g2_decap_8 FILLER_57_268 ();
 sg13g2_decap_8 FILLER_57_275 ();
 sg13g2_decap_4 FILLER_57_282 ();
 sg13g2_fill_2 FILLER_57_286 ();
 sg13g2_decap_4 FILLER_57_306 ();
 sg13g2_fill_1 FILLER_57_310 ();
 sg13g2_fill_2 FILLER_57_319 ();
 sg13g2_fill_1 FILLER_57_321 ();
 sg13g2_fill_2 FILLER_57_330 ();
 sg13g2_fill_2 FILLER_57_340 ();
 sg13g2_fill_1 FILLER_57_346 ();
 sg13g2_fill_1 FILLER_57_351 ();
 sg13g2_fill_2 FILLER_57_357 ();
 sg13g2_fill_1 FILLER_57_364 ();
 sg13g2_fill_2 FILLER_57_374 ();
 sg13g2_fill_1 FILLER_57_376 ();
 sg13g2_fill_2 FILLER_57_383 ();
 sg13g2_fill_1 FILLER_57_385 ();
 sg13g2_fill_1 FILLER_57_390 ();
 sg13g2_fill_2 FILLER_57_400 ();
 sg13g2_fill_1 FILLER_57_402 ();
 sg13g2_decap_4 FILLER_57_426 ();
 sg13g2_fill_1 FILLER_58_49 ();
 sg13g2_fill_2 FILLER_58_107 ();
 sg13g2_decap_8 FILLER_58_113 ();
 sg13g2_decap_8 FILLER_58_120 ();
 sg13g2_fill_1 FILLER_58_127 ();
 sg13g2_decap_8 FILLER_58_166 ();
 sg13g2_fill_1 FILLER_58_173 ();
 sg13g2_decap_8 FILLER_58_208 ();
 sg13g2_decap_8 FILLER_58_215 ();
 sg13g2_decap_8 FILLER_58_222 ();
 sg13g2_fill_2 FILLER_58_229 ();
 sg13g2_fill_1 FILLER_58_231 ();
 sg13g2_fill_2 FILLER_58_247 ();
 sg13g2_fill_2 FILLER_58_253 ();
 sg13g2_fill_2 FILLER_58_261 ();
 sg13g2_fill_2 FILLER_58_285 ();
 sg13g2_decap_8 FILLER_58_295 ();
 sg13g2_fill_1 FILLER_58_302 ();
 sg13g2_decap_8 FILLER_58_315 ();
 sg13g2_decap_8 FILLER_58_322 ();
 sg13g2_decap_8 FILLER_58_329 ();
 sg13g2_decap_4 FILLER_58_336 ();
 sg13g2_decap_8 FILLER_58_356 ();
 sg13g2_decap_8 FILLER_58_363 ();
 sg13g2_fill_2 FILLER_58_370 ();
 sg13g2_decap_8 FILLER_58_376 ();
 sg13g2_decap_4 FILLER_58_383 ();
 sg13g2_fill_2 FILLER_58_387 ();
 sg13g2_decap_4 FILLER_58_414 ();
 sg13g2_fill_2 FILLER_58_427 ();
 sg13g2_fill_1 FILLER_58_429 ();
 sg13g2_decap_8 FILLER_59_0 ();
 sg13g2_decap_4 FILLER_59_11 ();
 sg13g2_fill_2 FILLER_59_15 ();
 sg13g2_fill_1 FILLER_59_26 ();
 sg13g2_fill_2 FILLER_59_32 ();
 sg13g2_fill_1 FILLER_59_39 ();
 sg13g2_fill_2 FILLER_59_66 ();
 sg13g2_fill_2 FILLER_59_81 ();
 sg13g2_fill_1 FILLER_59_101 ();
 sg13g2_decap_4 FILLER_59_128 ();
 sg13g2_fill_2 FILLER_59_146 ();
 sg13g2_fill_1 FILLER_59_153 ();
 sg13g2_fill_2 FILLER_59_159 ();
 sg13g2_fill_1 FILLER_59_161 ();
 sg13g2_fill_1 FILLER_59_167 ();
 sg13g2_decap_8 FILLER_59_176 ();
 sg13g2_decap_4 FILLER_59_183 ();
 sg13g2_fill_1 FILLER_59_187 ();
 sg13g2_decap_8 FILLER_59_193 ();
 sg13g2_decap_8 FILLER_59_200 ();
 sg13g2_decap_8 FILLER_59_207 ();
 sg13g2_decap_4 FILLER_59_214 ();
 sg13g2_fill_1 FILLER_59_218 ();
 sg13g2_decap_8 FILLER_59_224 ();
 sg13g2_decap_4 FILLER_59_231 ();
 sg13g2_fill_1 FILLER_59_235 ();
 sg13g2_fill_1 FILLER_59_287 ();
 sg13g2_fill_2 FILLER_59_300 ();
 sg13g2_fill_1 FILLER_59_302 ();
 sg13g2_fill_2 FILLER_59_308 ();
 sg13g2_decap_8 FILLER_59_319 ();
 sg13g2_fill_1 FILLER_59_326 ();
 sg13g2_fill_1 FILLER_59_336 ();
 sg13g2_decap_4 FILLER_59_342 ();
 sg13g2_decap_4 FILLER_59_349 ();
 sg13g2_fill_2 FILLER_59_353 ();
 sg13g2_fill_2 FILLER_59_361 ();
 sg13g2_fill_1 FILLER_59_363 ();
 sg13g2_fill_2 FILLER_59_367 ();
 sg13g2_fill_1 FILLER_59_374 ();
 sg13g2_fill_1 FILLER_59_379 ();
 sg13g2_fill_1 FILLER_59_403 ();
 sg13g2_fill_2 FILLER_59_409 ();
 sg13g2_fill_1 FILLER_59_411 ();
 sg13g2_decap_4 FILLER_59_425 ();
 sg13g2_fill_1 FILLER_59_429 ();
 sg13g2_decap_8 FILLER_60_0 ();
 sg13g2_fill_1 FILLER_60_32 ();
 sg13g2_fill_1 FILLER_60_47 ();
 sg13g2_fill_1 FILLER_60_58 ();
 sg13g2_fill_1 FILLER_60_77 ();
 sg13g2_fill_1 FILLER_60_99 ();
 sg13g2_fill_1 FILLER_60_104 ();
 sg13g2_fill_1 FILLER_60_109 ();
 sg13g2_decap_8 FILLER_60_114 ();
 sg13g2_decap_4 FILLER_60_121 ();
 sg13g2_fill_1 FILLER_60_125 ();
 sg13g2_fill_2 FILLER_60_135 ();
 sg13g2_fill_1 FILLER_60_137 ();
 sg13g2_decap_8 FILLER_60_143 ();
 sg13g2_fill_2 FILLER_60_150 ();
 sg13g2_decap_4 FILLER_60_217 ();
 sg13g2_fill_2 FILLER_60_221 ();
 sg13g2_decap_4 FILLER_60_272 ();
 sg13g2_fill_1 FILLER_60_276 ();
 sg13g2_fill_1 FILLER_60_313 ();
 sg13g2_fill_2 FILLER_60_352 ();
 sg13g2_fill_1 FILLER_60_358 ();
 sg13g2_fill_1 FILLER_60_367 ();
 sg13g2_fill_1 FILLER_60_375 ();
 sg13g2_fill_1 FILLER_60_389 ();
 sg13g2_decap_8 FILLER_60_416 ();
 sg13g2_decap_8 FILLER_60_423 ();
 sg13g2_fill_2 FILLER_61_46 ();
 sg13g2_fill_2 FILLER_61_62 ();
 sg13g2_fill_1 FILLER_61_64 ();
 sg13g2_fill_2 FILLER_61_70 ();
 sg13g2_fill_1 FILLER_61_72 ();
 sg13g2_decap_4 FILLER_61_78 ();
 sg13g2_fill_1 FILLER_61_82 ();
 sg13g2_fill_2 FILLER_61_121 ();
 sg13g2_fill_1 FILLER_61_123 ();
 sg13g2_decap_4 FILLER_61_176 ();
 sg13g2_decap_4 FILLER_61_185 ();
 sg13g2_decap_4 FILLER_61_193 ();
 sg13g2_decap_8 FILLER_61_201 ();
 sg13g2_fill_1 FILLER_61_232 ();
 sg13g2_fill_1 FILLER_61_243 ();
 sg13g2_fill_2 FILLER_61_248 ();
 sg13g2_fill_2 FILLER_61_275 ();
 sg13g2_decap_4 FILLER_61_285 ();
 sg13g2_fill_1 FILLER_61_289 ();
 sg13g2_fill_1 FILLER_61_294 ();
 sg13g2_decap_4 FILLER_61_300 ();
 sg13g2_fill_1 FILLER_61_304 ();
 sg13g2_fill_1 FILLER_61_320 ();
 sg13g2_fill_1 FILLER_61_335 ();
 sg13g2_fill_1 FILLER_61_341 ();
 sg13g2_fill_1 FILLER_61_355 ();
 sg13g2_fill_1 FILLER_61_360 ();
 sg13g2_fill_1 FILLER_61_366 ();
 sg13g2_fill_1 FILLER_61_372 ();
 sg13g2_fill_1 FILLER_61_378 ();
 sg13g2_decap_8 FILLER_61_387 ();
 sg13g2_fill_2 FILLER_61_394 ();
 sg13g2_decap_8 FILLER_61_415 ();
 sg13g2_decap_8 FILLER_61_422 ();
 sg13g2_fill_1 FILLER_61_429 ();
 sg13g2_decap_8 FILLER_62_0 ();
 sg13g2_fill_1 FILLER_62_27 ();
 sg13g2_fill_2 FILLER_62_46 ();
 sg13g2_fill_1 FILLER_62_48 ();
 sg13g2_decap_4 FILLER_62_56 ();
 sg13g2_fill_2 FILLER_62_60 ();
 sg13g2_fill_1 FILLER_62_66 ();
 sg13g2_fill_1 FILLER_62_93 ();
 sg13g2_fill_1 FILLER_62_99 ();
 sg13g2_fill_1 FILLER_62_105 ();
 sg13g2_fill_1 FILLER_62_110 ();
 sg13g2_fill_2 FILLER_62_137 ();
 sg13g2_fill_1 FILLER_62_231 ();
 sg13g2_fill_1 FILLER_62_236 ();
 sg13g2_fill_1 FILLER_62_246 ();
 sg13g2_fill_2 FILLER_62_255 ();
 sg13g2_fill_1 FILLER_62_257 ();
 sg13g2_fill_1 FILLER_62_262 ();
 sg13g2_fill_1 FILLER_62_267 ();
 sg13g2_decap_4 FILLER_62_273 ();
 sg13g2_fill_2 FILLER_62_288 ();
 sg13g2_fill_1 FILLER_62_290 ();
 sg13g2_decap_8 FILLER_62_303 ();
 sg13g2_fill_2 FILLER_62_310 ();
 sg13g2_fill_1 FILLER_62_312 ();
 sg13g2_fill_1 FILLER_62_318 ();
 sg13g2_fill_1 FILLER_62_327 ();
 sg13g2_fill_1 FILLER_62_333 ();
 sg13g2_fill_2 FILLER_62_339 ();
 sg13g2_fill_2 FILLER_62_362 ();
 sg13g2_fill_1 FILLER_62_374 ();
 sg13g2_decap_4 FILLER_62_383 ();
 sg13g2_fill_2 FILLER_62_397 ();
 sg13g2_fill_1 FILLER_62_399 ();
 sg13g2_fill_2 FILLER_62_407 ();
 sg13g2_fill_1 FILLER_62_409 ();
 sg13g2_fill_2 FILLER_62_414 ();
 sg13g2_fill_1 FILLER_62_416 ();
 sg13g2_decap_8 FILLER_62_423 ();
 sg13g2_fill_2 FILLER_63_31 ();
 sg13g2_fill_1 FILLER_63_33 ();
 sg13g2_fill_1 FILLER_63_40 ();
 sg13g2_fill_1 FILLER_63_47 ();
 sg13g2_decap_4 FILLER_63_61 ();
 sg13g2_fill_1 FILLER_63_86 ();
 sg13g2_fill_2 FILLER_63_106 ();
 sg13g2_fill_1 FILLER_63_144 ();
 sg13g2_fill_2 FILLER_63_150 ();
 sg13g2_fill_1 FILLER_63_156 ();
 sg13g2_fill_2 FILLER_63_207 ();
 sg13g2_fill_1 FILLER_63_218 ();
 sg13g2_fill_2 FILLER_63_263 ();
 sg13g2_fill_2 FILLER_63_270 ();
 sg13g2_fill_1 FILLER_63_280 ();
 sg13g2_fill_1 FILLER_63_294 ();
 sg13g2_decap_8 FILLER_63_302 ();
 sg13g2_decap_4 FILLER_63_309 ();
 sg13g2_fill_1 FILLER_63_313 ();
 sg13g2_fill_1 FILLER_63_323 ();
 sg13g2_fill_2 FILLER_63_346 ();
 sg13g2_fill_2 FILLER_63_366 ();
 sg13g2_fill_2 FILLER_63_373 ();
 sg13g2_fill_1 FILLER_63_375 ();
 sg13g2_decap_8 FILLER_63_381 ();
 sg13g2_fill_1 FILLER_63_388 ();
 sg13g2_fill_2 FILLER_63_411 ();
 sg13g2_fill_1 FILLER_63_413 ();
 sg13g2_fill_2 FILLER_63_427 ();
 sg13g2_fill_1 FILLER_63_429 ();
 sg13g2_decap_8 FILLER_64_0 ();
 sg13g2_fill_2 FILLER_64_43 ();
 sg13g2_fill_1 FILLER_64_108 ();
 sg13g2_fill_1 FILLER_64_113 ();
 sg13g2_decap_8 FILLER_64_133 ();
 sg13g2_fill_2 FILLER_64_140 ();
 sg13g2_fill_1 FILLER_64_142 ();
 sg13g2_decap_8 FILLER_64_151 ();
 sg13g2_decap_8 FILLER_64_158 ();
 sg13g2_decap_4 FILLER_64_165 ();
 sg13g2_fill_1 FILLER_64_169 ();
 sg13g2_fill_2 FILLER_64_177 ();
 sg13g2_fill_2 FILLER_64_183 ();
 sg13g2_fill_2 FILLER_64_211 ();
 sg13g2_fill_1 FILLER_64_213 ();
 sg13g2_fill_2 FILLER_64_276 ();
 sg13g2_decap_4 FILLER_64_292 ();
 sg13g2_fill_2 FILLER_64_296 ();
 sg13g2_decap_8 FILLER_64_306 ();
 sg13g2_decap_4 FILLER_64_313 ();
 sg13g2_fill_2 FILLER_64_317 ();
 sg13g2_decap_8 FILLER_64_334 ();
 sg13g2_fill_1 FILLER_64_341 ();
 sg13g2_decap_8 FILLER_64_369 ();
 sg13g2_decap_8 FILLER_64_376 ();
 sg13g2_decap_4 FILLER_64_383 ();
 sg13g2_fill_1 FILLER_64_391 ();
 sg13g2_fill_1 FILLER_64_402 ();
 sg13g2_fill_1 FILLER_64_408 ();
 sg13g2_decap_8 FILLER_64_423 ();
 sg13g2_decap_8 FILLER_65_0 ();
 sg13g2_decap_4 FILLER_65_7 ();
 sg13g2_fill_1 FILLER_65_11 ();
 sg13g2_fill_2 FILLER_65_40 ();
 sg13g2_fill_1 FILLER_65_46 ();
 sg13g2_fill_2 FILLER_65_52 ();
 sg13g2_decap_8 FILLER_65_59 ();
 sg13g2_decap_8 FILLER_65_66 ();
 sg13g2_decap_4 FILLER_65_73 ();
 sg13g2_fill_1 FILLER_65_89 ();
 sg13g2_decap_4 FILLER_65_95 ();
 sg13g2_fill_1 FILLER_65_103 ();
 sg13g2_decap_8 FILLER_65_112 ();
 sg13g2_fill_2 FILLER_65_128 ();
 sg13g2_decap_8 FILLER_65_160 ();
 sg13g2_decap_8 FILLER_65_167 ();
 sg13g2_decap_8 FILLER_65_174 ();
 sg13g2_decap_8 FILLER_65_181 ();
 sg13g2_decap_4 FILLER_65_188 ();
 sg13g2_fill_1 FILLER_65_196 ();
 sg13g2_fill_1 FILLER_65_223 ();
 sg13g2_decap_8 FILLER_65_238 ();
 sg13g2_fill_2 FILLER_65_245 ();
 sg13g2_fill_1 FILLER_65_252 ();
 sg13g2_fill_2 FILLER_65_258 ();
 sg13g2_fill_1 FILLER_65_260 ();
 sg13g2_fill_2 FILLER_65_266 ();
 sg13g2_fill_2 FILLER_65_273 ();
 sg13g2_fill_1 FILLER_65_279 ();
 sg13g2_decap_8 FILLER_65_302 ();
 sg13g2_decap_8 FILLER_65_309 ();
 sg13g2_decap_8 FILLER_65_316 ();
 sg13g2_fill_1 FILLER_65_323 ();
 sg13g2_fill_1 FILLER_65_336 ();
 sg13g2_decap_8 FILLER_65_344 ();
 sg13g2_fill_1 FILLER_65_351 ();
 sg13g2_fill_2 FILLER_65_392 ();
 sg13g2_fill_1 FILLER_65_406 ();
 sg13g2_fill_2 FILLER_65_428 ();
 sg13g2_fill_1 FILLER_66_0 ();
 sg13g2_fill_2 FILLER_66_31 ();
 sg13g2_decap_8 FILLER_66_42 ();
 sg13g2_decap_4 FILLER_66_49 ();
 sg13g2_decap_8 FILLER_66_57 ();
 sg13g2_fill_2 FILLER_66_64 ();
 sg13g2_decap_4 FILLER_66_71 ();
 sg13g2_fill_1 FILLER_66_75 ();
 sg13g2_decap_8 FILLER_66_81 ();
 sg13g2_fill_1 FILLER_66_88 ();
 sg13g2_fill_1 FILLER_66_99 ();
 sg13g2_fill_2 FILLER_66_126 ();
 sg13g2_fill_1 FILLER_66_128 ();
 sg13g2_fill_2 FILLER_66_134 ();
 sg13g2_decap_4 FILLER_66_176 ();
 sg13g2_decap_8 FILLER_66_184 ();
 sg13g2_decap_4 FILLER_66_200 ();
 sg13g2_fill_1 FILLER_66_204 ();
 sg13g2_fill_2 FILLER_66_209 ();
 sg13g2_fill_1 FILLER_66_211 ();
 sg13g2_decap_8 FILLER_66_221 ();
 sg13g2_decap_4 FILLER_66_228 ();
 sg13g2_fill_1 FILLER_66_236 ();
 sg13g2_decap_8 FILLER_66_263 ();
 sg13g2_decap_4 FILLER_66_270 ();
 sg13g2_fill_1 FILLER_66_283 ();
 sg13g2_decap_8 FILLER_66_305 ();
 sg13g2_decap_8 FILLER_66_312 ();
 sg13g2_decap_8 FILLER_66_319 ();
 sg13g2_decap_8 FILLER_66_326 ();
 sg13g2_fill_2 FILLER_66_333 ();
 sg13g2_fill_1 FILLER_66_335 ();
 sg13g2_fill_1 FILLER_66_341 ();
 sg13g2_decap_4 FILLER_66_374 ();
 sg13g2_decap_4 FILLER_66_396 ();
 sg13g2_fill_2 FILLER_66_400 ();
 sg13g2_decap_4 FILLER_66_412 ();
 sg13g2_decap_8 FILLER_66_421 ();
 sg13g2_fill_2 FILLER_66_428 ();
 sg13g2_decap_8 FILLER_67_0 ();
 sg13g2_fill_2 FILLER_67_11 ();
 sg13g2_fill_2 FILLER_67_53 ();
 sg13g2_fill_2 FILLER_67_60 ();
 sg13g2_fill_1 FILLER_67_62 ();
 sg13g2_fill_1 FILLER_67_66 ();
 sg13g2_fill_2 FILLER_67_93 ();
 sg13g2_fill_1 FILLER_67_95 ();
 sg13g2_fill_2 FILLER_67_104 ();
 sg13g2_fill_1 FILLER_67_106 ();
 sg13g2_decap_4 FILLER_67_111 ();
 sg13g2_fill_1 FILLER_67_115 ();
 sg13g2_fill_2 FILLER_67_120 ();
 sg13g2_fill_1 FILLER_67_122 ();
 sg13g2_fill_1 FILLER_67_149 ();
 sg13g2_fill_2 FILLER_67_163 ();
 sg13g2_decap_4 FILLER_67_200 ();
 sg13g2_fill_1 FILLER_67_204 ();
 sg13g2_decap_4 FILLER_67_218 ();
 sg13g2_fill_2 FILLER_67_222 ();
 sg13g2_fill_2 FILLER_67_247 ();
 sg13g2_fill_1 FILLER_67_255 ();
 sg13g2_decap_4 FILLER_67_265 ();
 sg13g2_decap_8 FILLER_67_278 ();
 sg13g2_fill_2 FILLER_67_285 ();
 sg13g2_fill_1 FILLER_67_297 ();
 sg13g2_fill_1 FILLER_67_303 ();
 sg13g2_fill_2 FILLER_67_335 ();
 sg13g2_decap_4 FILLER_67_350 ();
 sg13g2_fill_2 FILLER_67_381 ();
 sg13g2_fill_1 FILLER_67_387 ();
 sg13g2_fill_1 FILLER_67_393 ();
 sg13g2_fill_1 FILLER_67_425 ();
 sg13g2_decap_8 FILLER_68_0 ();
 sg13g2_fill_2 FILLER_68_7 ();
 sg13g2_fill_2 FILLER_68_48 ();
 sg13g2_fill_2 FILLER_68_85 ();
 sg13g2_fill_1 FILLER_68_87 ();
 sg13g2_decap_4 FILLER_68_119 ();
 sg13g2_decap_4 FILLER_68_127 ();
 sg13g2_decap_8 FILLER_68_135 ();
 sg13g2_fill_1 FILLER_68_142 ();
 sg13g2_fill_2 FILLER_68_147 ();
 sg13g2_fill_1 FILLER_68_149 ();
 sg13g2_fill_1 FILLER_68_180 ();
 sg13g2_fill_1 FILLER_68_186 ();
 sg13g2_fill_2 FILLER_68_203 ();
 sg13g2_fill_1 FILLER_68_205 ();
 sg13g2_decap_8 FILLER_68_211 ();
 sg13g2_fill_1 FILLER_68_239 ();
 sg13g2_fill_1 FILLER_68_245 ();
 sg13g2_fill_1 FILLER_68_250 ();
 sg13g2_fill_2 FILLER_68_260 ();
 sg13g2_fill_1 FILLER_68_267 ();
 sg13g2_fill_1 FILLER_68_288 ();
 sg13g2_fill_1 FILLER_68_294 ();
 sg13g2_fill_1 FILLER_68_313 ();
 sg13g2_decap_8 FILLER_68_318 ();
 sg13g2_fill_2 FILLER_68_341 ();
 sg13g2_fill_1 FILLER_68_347 ();
 sg13g2_fill_2 FILLER_68_353 ();
 sg13g2_fill_1 FILLER_68_355 ();
 sg13g2_fill_1 FILLER_68_360 ();
 sg13g2_fill_1 FILLER_68_371 ();
 sg13g2_fill_2 FILLER_69_60 ();
 sg13g2_fill_1 FILLER_69_62 ();
 sg13g2_fill_2 FILLER_69_84 ();
 sg13g2_fill_1 FILLER_69_86 ();
 sg13g2_fill_2 FILLER_69_109 ();
 sg13g2_fill_1 FILLER_69_115 ();
 sg13g2_fill_2 FILLER_69_121 ();
 sg13g2_decap_8 FILLER_69_128 ();
 sg13g2_fill_2 FILLER_69_135 ();
 sg13g2_fill_2 FILLER_69_167 ();
 sg13g2_fill_1 FILLER_69_195 ();
 sg13g2_decap_4 FILLER_69_199 ();
 sg13g2_fill_1 FILLER_69_207 ();
 sg13g2_fill_1 FILLER_69_213 ();
 sg13g2_fill_1 FILLER_69_259 ();
 sg13g2_fill_1 FILLER_69_272 ();
 sg13g2_fill_1 FILLER_69_280 ();
 sg13g2_fill_1 FILLER_69_302 ();
 sg13g2_fill_2 FILLER_69_308 ();
 sg13g2_decap_8 FILLER_69_315 ();
 sg13g2_decap_4 FILLER_69_322 ();
 sg13g2_fill_2 FILLER_69_326 ();
 sg13g2_fill_2 FILLER_69_371 ();
 sg13g2_fill_1 FILLER_69_383 ();
 sg13g2_fill_2 FILLER_69_392 ();
 sg13g2_fill_2 FILLER_69_424 ();
 sg13g2_fill_2 FILLER_70_39 ();
 sg13g2_decap_4 FILLER_70_45 ();
 sg13g2_fill_1 FILLER_70_92 ();
 sg13g2_fill_1 FILLER_70_119 ();
 sg13g2_fill_2 FILLER_70_129 ();
 sg13g2_fill_2 FILLER_70_135 ();
 sg13g2_fill_1 FILLER_70_137 ();
 sg13g2_fill_2 FILLER_70_143 ();
 sg13g2_fill_2 FILLER_70_150 ();
 sg13g2_fill_1 FILLER_70_152 ();
 sg13g2_fill_1 FILLER_70_158 ();
 sg13g2_fill_2 FILLER_70_164 ();
 sg13g2_fill_1 FILLER_70_166 ();
 sg13g2_fill_2 FILLER_70_172 ();
 sg13g2_fill_1 FILLER_70_174 ();
 sg13g2_fill_2 FILLER_70_179 ();
 sg13g2_fill_1 FILLER_70_181 ();
 sg13g2_fill_2 FILLER_70_186 ();
 sg13g2_fill_1 FILLER_70_188 ();
 sg13g2_fill_1 FILLER_70_193 ();
 sg13g2_fill_1 FILLER_70_200 ();
 sg13g2_fill_1 FILLER_70_215 ();
 sg13g2_decap_4 FILLER_70_225 ();
 sg13g2_fill_2 FILLER_70_241 ();
 sg13g2_fill_2 FILLER_70_249 ();
 sg13g2_fill_2 FILLER_70_256 ();
 sg13g2_fill_1 FILLER_70_258 ();
 sg13g2_fill_2 FILLER_70_296 ();
 sg13g2_fill_2 FILLER_70_376 ();
 sg13g2_fill_1 FILLER_70_378 ();
 sg13g2_fill_1 FILLER_70_384 ();
 sg13g2_decap_8 FILLER_70_389 ();
 sg13g2_fill_2 FILLER_70_396 ();
 sg13g2_fill_1 FILLER_70_398 ();
 sg13g2_fill_1 FILLER_70_404 ();
 sg13g2_fill_2 FILLER_70_427 ();
 sg13g2_fill_1 FILLER_70_429 ();
 sg13g2_decap_4 FILLER_71_0 ();
 sg13g2_fill_1 FILLER_71_12 ();
 sg13g2_decap_4 FILLER_71_17 ();
 sg13g2_fill_1 FILLER_71_21 ();
 sg13g2_decap_8 FILLER_71_33 ();
 sg13g2_fill_2 FILLER_71_40 ();
 sg13g2_fill_1 FILLER_71_42 ();
 sg13g2_decap_8 FILLER_71_47 ();
 sg13g2_decap_8 FILLER_71_54 ();
 sg13g2_decap_8 FILLER_71_61 ();
 sg13g2_decap_8 FILLER_71_68 ();
 sg13g2_fill_2 FILLER_71_75 ();
 sg13g2_decap_4 FILLER_71_90 ();
 sg13g2_fill_1 FILLER_71_98 ();
 sg13g2_fill_1 FILLER_71_103 ();
 sg13g2_fill_1 FILLER_71_108 ();
 sg13g2_fill_1 FILLER_71_112 ();
 sg13g2_fill_1 FILLER_71_119 ();
 sg13g2_fill_2 FILLER_71_125 ();
 sg13g2_decap_4 FILLER_71_131 ();
 sg13g2_fill_1 FILLER_71_135 ();
 sg13g2_fill_2 FILLER_71_148 ();
 sg13g2_decap_8 FILLER_71_180 ();
 sg13g2_decap_8 FILLER_71_187 ();
 sg13g2_fill_1 FILLER_71_203 ();
 sg13g2_fill_1 FILLER_71_209 ();
 sg13g2_fill_1 FILLER_71_222 ();
 sg13g2_fill_2 FILLER_71_228 ();
 sg13g2_fill_2 FILLER_71_235 ();
 sg13g2_decap_8 FILLER_71_250 ();
 sg13g2_decap_8 FILLER_71_257 ();
 sg13g2_fill_1 FILLER_71_264 ();
 sg13g2_fill_2 FILLER_71_278 ();
 sg13g2_fill_1 FILLER_71_285 ();
 sg13g2_fill_1 FILLER_71_296 ();
 sg13g2_fill_1 FILLER_71_302 ();
 sg13g2_decap_4 FILLER_71_313 ();
 sg13g2_fill_2 FILLER_71_317 ();
 sg13g2_decap_4 FILLER_71_327 ();
 sg13g2_fill_2 FILLER_71_331 ();
 sg13g2_fill_1 FILLER_71_336 ();
 sg13g2_fill_2 FILLER_71_342 ();
 sg13g2_fill_2 FILLER_71_348 ();
 sg13g2_fill_1 FILLER_71_372 ();
 sg13g2_fill_1 FILLER_71_377 ();
 sg13g2_fill_2 FILLER_71_391 ();
 sg13g2_decap_8 FILLER_71_402 ();
 sg13g2_decap_4 FILLER_71_409 ();
 sg13g2_fill_2 FILLER_71_413 ();
 sg13g2_decap_8 FILLER_71_420 ();
 sg13g2_fill_2 FILLER_71_427 ();
 sg13g2_fill_1 FILLER_71_429 ();
 sg13g2_decap_4 FILLER_72_0 ();
 sg13g2_decap_8 FILLER_72_8 ();
 sg13g2_decap_8 FILLER_72_15 ();
 sg13g2_decap_8 FILLER_72_22 ();
 sg13g2_decap_4 FILLER_72_29 ();
 sg13g2_fill_1 FILLER_72_63 ();
 sg13g2_fill_1 FILLER_72_68 ();
 sg13g2_decap_4 FILLER_72_104 ();
 sg13g2_decap_4 FILLER_72_112 ();
 sg13g2_fill_1 FILLER_72_130 ();
 sg13g2_fill_1 FILLER_72_136 ();
 sg13g2_fill_1 FILLER_72_154 ();
 sg13g2_fill_1 FILLER_72_186 ();
 sg13g2_fill_1 FILLER_72_204 ();
 sg13g2_fill_1 FILLER_72_209 ();
 sg13g2_decap_8 FILLER_72_240 ();
 sg13g2_fill_1 FILLER_72_247 ();
 sg13g2_fill_2 FILLER_72_269 ();
 sg13g2_fill_2 FILLER_72_283 ();
 sg13g2_fill_1 FILLER_72_285 ();
 sg13g2_fill_1 FILLER_72_312 ();
 sg13g2_decap_8 FILLER_72_317 ();
 sg13g2_decap_8 FILLER_72_324 ();
 sg13g2_decap_4 FILLER_72_331 ();
 sg13g2_fill_1 FILLER_72_335 ();
 sg13g2_fill_1 FILLER_72_341 ();
 sg13g2_fill_2 FILLER_72_346 ();
 sg13g2_fill_2 FILLER_72_365 ();
 sg13g2_fill_2 FILLER_72_380 ();
 sg13g2_decap_8 FILLER_72_413 ();
 sg13g2_decap_8 FILLER_72_420 ();
 sg13g2_fill_2 FILLER_72_427 ();
 sg13g2_fill_1 FILLER_72_429 ();
 sg13g2_fill_2 FILLER_73_26 ();
 sg13g2_fill_1 FILLER_73_28 ();
 sg13g2_decap_4 FILLER_73_66 ();
 sg13g2_fill_2 FILLER_73_74 ();
 sg13g2_fill_1 FILLER_73_89 ();
 sg13g2_decap_8 FILLER_73_129 ();
 sg13g2_decap_4 FILLER_73_147 ();
 sg13g2_fill_1 FILLER_73_151 ();
 sg13g2_decap_4 FILLER_73_161 ();
 sg13g2_fill_1 FILLER_73_165 ();
 sg13g2_fill_2 FILLER_73_205 ();
 sg13g2_fill_1 FILLER_73_222 ();
 sg13g2_fill_1 FILLER_73_228 ();
 sg13g2_fill_1 FILLER_73_233 ();
 sg13g2_fill_1 FILLER_73_239 ();
 sg13g2_fill_1 FILLER_73_250 ();
 sg13g2_fill_2 FILLER_73_265 ();
 sg13g2_fill_1 FILLER_73_267 ();
 sg13g2_decap_4 FILLER_73_272 ();
 sg13g2_fill_1 FILLER_73_276 ();
 sg13g2_fill_1 FILLER_73_287 ();
 sg13g2_fill_2 FILLER_73_305 ();
 sg13g2_decap_8 FILLER_73_311 ();
 sg13g2_decap_8 FILLER_73_318 ();
 sg13g2_decap_4 FILLER_73_325 ();
 sg13g2_fill_2 FILLER_73_329 ();
 sg13g2_decap_8 FILLER_73_335 ();
 sg13g2_fill_2 FILLER_73_342 ();
 sg13g2_fill_1 FILLER_73_344 ();
 sg13g2_fill_1 FILLER_73_350 ();
 sg13g2_fill_2 FILLER_73_360 ();
 sg13g2_fill_2 FILLER_73_370 ();
 sg13g2_fill_1 FILLER_73_377 ();
 sg13g2_fill_1 FILLER_73_383 ();
 sg13g2_fill_1 FILLER_73_389 ();
 sg13g2_fill_2 FILLER_73_394 ();
 sg13g2_decap_8 FILLER_73_422 ();
 sg13g2_fill_1 FILLER_73_429 ();
 sg13g2_decap_8 FILLER_74_0 ();
 sg13g2_decap_4 FILLER_74_71 ();
 sg13g2_fill_1 FILLER_74_75 ();
 sg13g2_fill_1 FILLER_74_79 ();
 sg13g2_fill_2 FILLER_74_84 ();
 sg13g2_fill_1 FILLER_74_86 ();
 sg13g2_fill_1 FILLER_74_91 ();
 sg13g2_decap_4 FILLER_74_121 ();
 sg13g2_fill_1 FILLER_74_134 ();
 sg13g2_fill_2 FILLER_74_140 ();
 sg13g2_fill_1 FILLER_74_142 ();
 sg13g2_fill_2 FILLER_74_148 ();
 sg13g2_fill_1 FILLER_74_150 ();
 sg13g2_decap_8 FILLER_74_159 ();
 sg13g2_decap_8 FILLER_74_166 ();
 sg13g2_decap_8 FILLER_74_173 ();
 sg13g2_fill_1 FILLER_74_180 ();
 sg13g2_decap_4 FILLER_74_207 ();
 sg13g2_fill_2 FILLER_74_211 ();
 sg13g2_decap_8 FILLER_74_217 ();
 sg13g2_decap_4 FILLER_74_224 ();
 sg13g2_fill_1 FILLER_74_228 ();
 sg13g2_fill_2 FILLER_74_241 ();
 sg13g2_fill_1 FILLER_74_253 ();
 sg13g2_fill_1 FILLER_74_259 ();
 sg13g2_decap_8 FILLER_74_282 ();
 sg13g2_fill_2 FILLER_74_289 ();
 sg13g2_fill_1 FILLER_74_291 ();
 sg13g2_fill_2 FILLER_74_322 ();
 sg13g2_fill_2 FILLER_74_329 ();
 sg13g2_fill_1 FILLER_74_331 ();
 sg13g2_decap_4 FILLER_74_337 ();
 sg13g2_fill_1 FILLER_74_341 ();
 sg13g2_decap_8 FILLER_74_347 ();
 sg13g2_fill_1 FILLER_74_354 ();
 sg13g2_decap_8 FILLER_74_368 ();
 sg13g2_fill_1 FILLER_74_375 ();
 sg13g2_fill_1 FILLER_74_413 ();
 sg13g2_decap_8 FILLER_74_418 ();
 sg13g2_decap_4 FILLER_74_425 ();
 sg13g2_fill_1 FILLER_74_429 ();
 sg13g2_decap_8 FILLER_75_0 ();
 sg13g2_decap_8 FILLER_75_7 ();
 sg13g2_fill_2 FILLER_75_14 ();
 sg13g2_fill_1 FILLER_75_16 ();
 sg13g2_decap_8 FILLER_75_38 ();
 sg13g2_fill_2 FILLER_75_45 ();
 sg13g2_fill_2 FILLER_75_54 ();
 sg13g2_fill_1 FILLER_75_56 ();
 sg13g2_fill_2 FILLER_75_62 ();
 sg13g2_decap_4 FILLER_75_69 ();
 sg13g2_fill_2 FILLER_75_91 ();
 sg13g2_fill_1 FILLER_75_93 ();
 sg13g2_fill_2 FILLER_75_99 ();
 sg13g2_fill_2 FILLER_75_106 ();
 sg13g2_fill_2 FILLER_75_112 ();
 sg13g2_decap_4 FILLER_75_130 ();
 sg13g2_decap_8 FILLER_75_155 ();
 sg13g2_decap_4 FILLER_75_162 ();
 sg13g2_decap_8 FILLER_75_170 ();
 sg13g2_decap_8 FILLER_75_177 ();
 sg13g2_decap_4 FILLER_75_184 ();
 sg13g2_fill_2 FILLER_75_188 ();
 sg13g2_decap_8 FILLER_75_194 ();
 sg13g2_decap_8 FILLER_75_201 ();
 sg13g2_fill_1 FILLER_75_208 ();
 sg13g2_fill_2 FILLER_75_214 ();
 sg13g2_fill_1 FILLER_75_216 ();
 sg13g2_fill_2 FILLER_75_220 ();
 sg13g2_fill_1 FILLER_75_222 ();
 sg13g2_decap_4 FILLER_75_235 ();
 sg13g2_fill_2 FILLER_75_244 ();
 sg13g2_decap_4 FILLER_75_251 ();
 sg13g2_fill_2 FILLER_75_255 ();
 sg13g2_fill_1 FILLER_75_275 ();
 sg13g2_fill_2 FILLER_75_280 ();
 sg13g2_fill_1 FILLER_75_282 ();
 sg13g2_fill_1 FILLER_75_293 ();
 sg13g2_fill_1 FILLER_75_299 ();
 sg13g2_fill_1 FILLER_75_305 ();
 sg13g2_fill_1 FILLER_75_332 ();
 sg13g2_fill_1 FILLER_75_343 ();
 sg13g2_fill_1 FILLER_75_348 ();
 sg13g2_fill_2 FILLER_75_354 ();
 sg13g2_fill_2 FILLER_75_387 ();
 sg13g2_fill_2 FILLER_75_394 ();
 sg13g2_fill_1 FILLER_75_396 ();
 sg13g2_decap_4 FILLER_75_404 ();
 sg13g2_decap_8 FILLER_75_413 ();
 sg13g2_decap_8 FILLER_75_420 ();
 sg13g2_fill_2 FILLER_75_427 ();
 sg13g2_fill_1 FILLER_75_429 ();
 sg13g2_decap_8 FILLER_76_0 ();
 sg13g2_decap_8 FILLER_76_7 ();
 sg13g2_decap_8 FILLER_76_14 ();
 sg13g2_decap_8 FILLER_76_21 ();
 sg13g2_fill_2 FILLER_76_28 ();
 sg13g2_decap_8 FILLER_76_34 ();
 sg13g2_decap_8 FILLER_76_41 ();
 sg13g2_decap_4 FILLER_76_72 ();
 sg13g2_fill_2 FILLER_76_81 ();
 sg13g2_decap_8 FILLER_76_109 ();
 sg13g2_fill_2 FILLER_76_116 ();
 sg13g2_fill_1 FILLER_76_121 ();
 sg13g2_fill_2 FILLER_76_127 ();
 sg13g2_fill_1 FILLER_76_144 ();
 sg13g2_fill_1 FILLER_76_150 ();
 sg13g2_fill_2 FILLER_76_177 ();
 sg13g2_fill_1 FILLER_76_223 ();
 sg13g2_fill_1 FILLER_76_229 ();
 sg13g2_fill_2 FILLER_76_234 ();
 sg13g2_fill_2 FILLER_76_260 ();
 sg13g2_fill_2 FILLER_76_270 ();
 sg13g2_fill_1 FILLER_76_276 ();
 sg13g2_fill_2 FILLER_76_290 ();
 sg13g2_fill_2 FILLER_76_307 ();
 sg13g2_fill_1 FILLER_76_309 ();
 sg13g2_fill_1 FILLER_76_314 ();
 sg13g2_decap_8 FILLER_76_323 ();
 sg13g2_fill_1 FILLER_76_344 ();
 sg13g2_fill_1 FILLER_76_355 ();
 sg13g2_fill_2 FILLER_76_373 ();
 sg13g2_fill_1 FILLER_76_375 ();
 sg13g2_decap_8 FILLER_76_407 ();
 sg13g2_decap_8 FILLER_76_414 ();
 sg13g2_decap_8 FILLER_76_421 ();
 sg13g2_fill_2 FILLER_76_428 ();
 sg13g2_decap_8 FILLER_77_0 ();
 sg13g2_fill_1 FILLER_77_7 ();
 sg13g2_fill_2 FILLER_77_38 ();
 sg13g2_fill_2 FILLER_77_52 ();
 sg13g2_fill_1 FILLER_77_54 ();
 sg13g2_fill_2 FILLER_77_95 ();
 sg13g2_fill_1 FILLER_77_97 ();
 sg13g2_decap_8 FILLER_77_106 ();
 sg13g2_fill_1 FILLER_77_113 ();
 sg13g2_fill_1 FILLER_77_132 ();
 sg13g2_fill_2 FILLER_77_153 ();
 sg13g2_fill_1 FILLER_77_189 ();
 sg13g2_fill_1 FILLER_77_287 ();
 sg13g2_fill_2 FILLER_77_298 ();
 sg13g2_fill_2 FILLER_77_304 ();
 sg13g2_fill_2 FILLER_77_315 ();
 sg13g2_fill_1 FILLER_77_317 ();
 sg13g2_fill_2 FILLER_77_331 ();
 sg13g2_fill_1 FILLER_77_339 ();
 sg13g2_fill_1 FILLER_77_347 ();
 sg13g2_fill_1 FILLER_77_361 ();
 sg13g2_fill_1 FILLER_77_376 ();
 sg13g2_decap_8 FILLER_77_402 ();
 sg13g2_decap_8 FILLER_77_409 ();
 sg13g2_decap_8 FILLER_77_416 ();
 sg13g2_decap_8 FILLER_77_423 ();
 sg13g2_decap_8 FILLER_78_0 ();
 sg13g2_decap_8 FILLER_78_7 ();
 sg13g2_fill_2 FILLER_78_14 ();
 sg13g2_fill_1 FILLER_78_55 ();
 sg13g2_fill_1 FILLER_78_69 ();
 sg13g2_fill_1 FILLER_78_75 ();
 sg13g2_fill_1 FILLER_78_80 ();
 sg13g2_fill_1 FILLER_78_90 ();
 sg13g2_fill_2 FILLER_78_117 ();
 sg13g2_fill_1 FILLER_78_141 ();
 sg13g2_fill_2 FILLER_78_151 ();
 sg13g2_decap_8 FILLER_78_162 ();
 sg13g2_fill_2 FILLER_78_169 ();
 sg13g2_fill_1 FILLER_78_180 ();
 sg13g2_decap_4 FILLER_78_211 ();
 sg13g2_fill_1 FILLER_78_215 ();
 sg13g2_fill_2 FILLER_78_221 ();
 sg13g2_fill_1 FILLER_78_223 ();
 sg13g2_decap_4 FILLER_78_315 ();
 sg13g2_fill_2 FILLER_78_343 ();
 sg13g2_fill_1 FILLER_78_382 ();
 sg13g2_decap_8 FILLER_78_413 ();
 sg13g2_decap_8 FILLER_78_420 ();
 sg13g2_fill_2 FILLER_78_427 ();
 sg13g2_fill_1 FILLER_78_429 ();
 sg13g2_decap_8 FILLER_79_0 ();
 sg13g2_decap_8 FILLER_79_7 ();
 sg13g2_decap_4 FILLER_79_14 ();
 sg13g2_fill_1 FILLER_79_18 ();
 sg13g2_fill_1 FILLER_79_23 ();
 sg13g2_fill_2 FILLER_79_32 ();
 sg13g2_fill_2 FILLER_79_64 ();
 sg13g2_fill_2 FILLER_79_92 ();
 sg13g2_fill_1 FILLER_79_94 ();
 sg13g2_fill_2 FILLER_79_125 ();
 sg13g2_decap_4 FILLER_79_205 ();
 sg13g2_decap_8 FILLER_79_213 ();
 sg13g2_fill_1 FILLER_79_220 ();
 sg13g2_decap_4 FILLER_79_229 ();
 sg13g2_fill_1 FILLER_79_246 ();
 sg13g2_fill_1 FILLER_79_251 ();
 sg13g2_fill_2 FILLER_79_257 ();
 sg13g2_fill_2 FILLER_79_263 ();
 sg13g2_decap_4 FILLER_79_269 ();
 sg13g2_decap_8 FILLER_79_278 ();
 sg13g2_fill_2 FILLER_79_285 ();
 sg13g2_fill_1 FILLER_79_287 ();
 sg13g2_fill_1 FILLER_79_344 ();
 sg13g2_fill_1 FILLER_79_398 ();
 sg13g2_decap_8 FILLER_79_404 ();
 sg13g2_decap_8 FILLER_79_411 ();
 sg13g2_decap_8 FILLER_79_418 ();
 sg13g2_decap_4 FILLER_79_425 ();
 sg13g2_fill_1 FILLER_79_429 ();
 sg13g2_decap_8 FILLER_80_0 ();
 sg13g2_decap_8 FILLER_80_7 ();
 sg13g2_decap_8 FILLER_80_14 ();
 sg13g2_decap_8 FILLER_80_21 ();
 sg13g2_fill_2 FILLER_80_28 ();
 sg13g2_fill_1 FILLER_80_30 ();
 sg13g2_decap_4 FILLER_80_35 ();
 sg13g2_fill_2 FILLER_80_39 ();
 sg13g2_decap_8 FILLER_80_45 ();
 sg13g2_fill_1 FILLER_80_56 ();
 sg13g2_fill_2 FILLER_80_62 ();
 sg13g2_decap_4 FILLER_80_67 ();
 sg13g2_fill_1 FILLER_80_71 ();
 sg13g2_fill_1 FILLER_80_96 ();
 sg13g2_fill_2 FILLER_80_125 ();
 sg13g2_fill_2 FILLER_80_147 ();
 sg13g2_fill_1 FILLER_80_153 ();
 sg13g2_fill_1 FILLER_80_158 ();
 sg13g2_fill_1 FILLER_80_163 ();
 sg13g2_fill_1 FILLER_80_168 ();
 sg13g2_fill_1 FILLER_80_177 ();
 sg13g2_fill_2 FILLER_80_194 ();
 sg13g2_fill_1 FILLER_80_204 ();
 sg13g2_fill_2 FILLER_80_209 ();
 sg13g2_fill_2 FILLER_80_215 ();
 sg13g2_fill_1 FILLER_80_221 ();
 sg13g2_fill_1 FILLER_80_226 ();
 sg13g2_fill_1 FILLER_80_235 ();
 sg13g2_fill_1 FILLER_80_240 ();
 sg13g2_fill_1 FILLER_80_253 ();
 sg13g2_fill_2 FILLER_80_258 ();
 sg13g2_decap_8 FILLER_80_264 ();
 sg13g2_decap_8 FILLER_80_271 ();
 sg13g2_decap_4 FILLER_80_278 ();
 sg13g2_fill_2 FILLER_80_282 ();
 sg13g2_decap_8 FILLER_80_288 ();
 sg13g2_fill_2 FILLER_80_303 ();
 sg13g2_decap_8 FILLER_80_312 ();
 sg13g2_decap_4 FILLER_80_319 ();
 sg13g2_fill_1 FILLER_80_323 ();
 sg13g2_decap_8 FILLER_80_328 ();
 sg13g2_decap_8 FILLER_80_335 ();
 sg13g2_decap_8 FILLER_80_342 ();
 sg13g2_decap_8 FILLER_80_349 ();
 sg13g2_decap_8 FILLER_80_356 ();
 sg13g2_decap_8 FILLER_80_363 ();
 sg13g2_decap_8 FILLER_80_370 ();
 sg13g2_decap_8 FILLER_80_377 ();
 sg13g2_decap_8 FILLER_80_384 ();
 sg13g2_decap_8 FILLER_80_391 ();
 sg13g2_decap_8 FILLER_80_398 ();
 sg13g2_decap_8 FILLER_80_405 ();
 sg13g2_decap_8 FILLER_80_412 ();
 sg13g2_decap_8 FILLER_80_419 ();
 sg13g2_decap_4 FILLER_80_426 ();
endmodule
