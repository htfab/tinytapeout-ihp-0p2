module tt_um_tomkeddie_a (clk,
    ena,
    rst_n,
    ui_in,
    uio_in,
    uio_oe,
    uio_out,
    uo_out);
 input clk;
 input ena;
 input rst_n;
 input [7:0] ui_in;
 input [7:0] uio_in;
 output [7:0] uio_oe;
 output [7:0] uio_out;
 output [7:0] uo_out;

 wire _0000_;
 wire _0001_;
 wire _0002_;
 wire _0003_;
 wire _0004_;
 wire _0005_;
 wire _0006_;
 wire _0007_;
 wire _0008_;
 wire _0009_;
 wire _0010_;
 wire _0011_;
 wire _0012_;
 wire _0013_;
 wire _0014_;
 wire _0015_;
 wire _0016_;
 wire _0017_;
 wire _0018_;
 wire _0019_;
 wire _0020_;
 wire _0021_;
 wire _0022_;
 wire _0023_;
 wire _0024_;
 wire _0025_;
 wire _0026_;
 wire _0027_;
 wire _0028_;
 wire _0029_;
 wire _0030_;
 wire _0031_;
 wire _0032_;
 wire _0033_;
 wire _0034_;
 wire _0035_;
 wire _0036_;
 wire _0037_;
 wire _0038_;
 wire _0039_;
 wire _0040_;
 wire _0041_;
 wire _0042_;
 wire _0043_;
 wire _0044_;
 wire _0045_;
 wire _0046_;
 wire _0047_;
 wire _0048_;
 wire _0049_;
 wire _0050_;
 wire _0051_;
 wire _0052_;
 wire _0053_;
 wire _0054_;
 wire _0055_;
 wire _0056_;
 wire _0057_;
 wire _0058_;
 wire _0059_;
 wire _0060_;
 wire _0061_;
 wire _0062_;
 wire _0063_;
 wire _0064_;
 wire _0065_;
 wire _0066_;
 wire _0067_;
 wire _0068_;
 wire _0069_;
 wire _0070_;
 wire _0071_;
 wire _0072_;
 wire _0073_;
 wire _0074_;
 wire _0075_;
 wire _0076_;
 wire _0077_;
 wire _0078_;
 wire _0079_;
 wire _0080_;
 wire _0081_;
 wire _0082_;
 wire _0083_;
 wire _0084_;
 wire _0085_;
 wire _0086_;
 wire _0087_;
 wire _0088_;
 wire _0089_;
 wire _0090_;
 wire _0091_;
 wire _0092_;
 wire _0093_;
 wire _0094_;
 wire _0095_;
 wire _0096_;
 wire _0097_;
 wire _0098_;
 wire _0099_;
 wire _0100_;
 wire _0101_;
 wire _0102_;
 wire _0103_;
 wire _0104_;
 wire _0105_;
 wire _0106_;
 wire _0107_;
 wire _0108_;
 wire _0109_;
 wire _0110_;
 wire _0111_;
 wire _0112_;
 wire _0113_;
 wire _0114_;
 wire _0115_;
 wire _0116_;
 wire _0117_;
 wire _0118_;
 wire _0119_;
 wire _0120_;
 wire _0121_;
 wire _0122_;
 wire _0123_;
 wire _0124_;
 wire _0125_;
 wire _0126_;
 wire _0127_;
 wire _0128_;
 wire _0129_;
 wire _0130_;
 wire _0131_;
 wire _0132_;
 wire _0133_;
 wire _0134_;
 wire _0135_;
 wire _0136_;
 wire _0137_;
 wire _0138_;
 wire _0139_;
 wire _0140_;
 wire _0141_;
 wire _0142_;
 wire _0143_;
 wire _0144_;
 wire _0145_;
 wire _0146_;
 wire _0147_;
 wire _0148_;
 wire _0149_;
 wire _0150_;
 wire _0151_;
 wire _0152_;
 wire _0153_;
 wire _0154_;
 wire _0155_;
 wire _0156_;
 wire _0157_;
 wire _0158_;
 wire _0159_;
 wire _0160_;
 wire _0161_;
 wire _0162_;
 wire _0163_;
 wire _0164_;
 wire _0165_;
 wire _0166_;
 wire _0167_;
 wire _0168_;
 wire _0169_;
 wire _0170_;
 wire _0171_;
 wire _0172_;
 wire _0173_;
 wire _0174_;
 wire _0175_;
 wire _0176_;
 wire _0177_;
 wire _0178_;
 wire _0179_;
 wire _0180_;
 wire _0181_;
 wire _0182_;
 wire _0183_;
 wire _0184_;
 wire _0185_;
 wire _0186_;
 wire _0187_;
 wire _0188_;
 wire _0189_;
 wire _0190_;
 wire _0191_;
 wire _0192_;
 wire _0193_;
 wire _0194_;
 wire _0195_;
 wire _0196_;
 wire _0197_;
 wire _0198_;
 wire _0199_;
 wire _0200_;
 wire _0201_;
 wire _0202_;
 wire _0203_;
 wire _0204_;
 wire _0205_;
 wire _0206_;
 wire _0207_;
 wire _0208_;
 wire _0209_;
 wire _0210_;
 wire _0211_;
 wire _0212_;
 wire _0213_;
 wire _0214_;
 wire _0215_;
 wire _0216_;
 wire _0217_;
 wire _0218_;
 wire _0219_;
 wire _0220_;
 wire _0221_;
 wire _0222_;
 wire _0223_;
 wire _0224_;
 wire _0225_;
 wire _0226_;
 wire _0227_;
 wire _0228_;
 wire _0229_;
 wire _0230_;
 wire _0231_;
 wire _0232_;
 wire _0233_;
 wire _0234_;
 wire _0235_;
 wire _0236_;
 wire _0237_;
 wire _0238_;
 wire _0239_;
 wire _0240_;
 wire _0241_;
 wire _0242_;
 wire _0243_;
 wire _0244_;
 wire _0245_;
 wire _0246_;
 wire _0247_;
 wire _0248_;
 wire _0249_;
 wire _0250_;
 wire _0251_;
 wire _0252_;
 wire _0253_;
 wire _0254_;
 wire _0255_;
 wire _0256_;
 wire _0257_;
 wire _0258_;
 wire _0259_;
 wire _0260_;
 wire _0261_;
 wire _0262_;
 wire _0263_;
 wire _0264_;
 wire _0265_;
 wire _0266_;
 wire _0267_;
 wire _0268_;
 wire _0269_;
 wire _0270_;
 wire _0271_;
 wire _0272_;
 wire _0273_;
 wire _0274_;
 wire _0275_;
 wire _0276_;
 wire _0277_;
 wire _0278_;
 wire _0279_;
 wire _0280_;
 wire _0281_;
 wire _0282_;
 wire _0283_;
 wire _0284_;
 wire _0285_;
 wire _0286_;
 wire _0287_;
 wire _0288_;
 wire _0289_;
 wire _0290_;
 wire _0291_;
 wire _0292_;
 wire _0293_;
 wire _0294_;
 wire _0295_;
 wire _0296_;
 wire _0297_;
 wire _0298_;
 wire _0299_;
 wire _0300_;
 wire _0301_;
 wire _0302_;
 wire _0303_;
 wire _0304_;
 wire _0305_;
 wire _0306_;
 wire _0307_;
 wire _0308_;
 wire _0309_;
 wire _0310_;
 wire _0311_;
 wire _0312_;
 wire _0313_;
 wire _0314_;
 wire _0315_;
 wire _0316_;
 wire _0317_;
 wire _0318_;
 wire _0319_;
 wire _0320_;
 wire _0321_;
 wire _0322_;
 wire _0323_;
 wire _0324_;
 wire _0325_;
 wire _0326_;
 wire _0327_;
 wire _0328_;
 wire _0329_;
 wire _0330_;
 wire _0331_;
 wire _0332_;
 wire _0333_;
 wire _0334_;
 wire _0335_;
 wire _0336_;
 wire _0337_;
 wire _0338_;
 wire _0339_;
 wire _0340_;
 wire _0341_;
 wire _0342_;
 wire _0343_;
 wire _0344_;
 wire _0345_;
 wire _0346_;
 wire _0347_;
 wire _0348_;
 wire _0349_;
 wire _0350_;
 wire _0351_;
 wire _0352_;
 wire _0353_;
 wire _0354_;
 wire _0355_;
 wire _0356_;
 wire _0357_;
 wire _0358_;
 wire _0359_;
 wire _0360_;
 wire _0361_;
 wire _0362_;
 wire _0363_;
 wire _0364_;
 wire _0365_;
 wire _0366_;
 wire _0367_;
 wire _0368_;
 wire _0369_;
 wire _0370_;
 wire _0371_;
 wire _0372_;
 wire _0373_;
 wire _0374_;
 wire _0375_;
 wire _0376_;
 wire _0377_;
 wire _0378_;
 wire _0379_;
 wire _0380_;
 wire _0381_;
 wire _0382_;
 wire _0383_;
 wire _0384_;
 wire _0385_;
 wire _0386_;
 wire _0387_;
 wire _0388_;
 wire _0389_;
 wire _0390_;
 wire _0391_;
 wire _0392_;
 wire _0393_;
 wire _0394_;
 wire _0395_;
 wire _0396_;
 wire _0397_;
 wire _0398_;
 wire _0399_;
 wire _0400_;
 wire _0401_;
 wire _0402_;
 wire _0403_;
 wire _0404_;
 wire _0405_;
 wire _0406_;
 wire _0407_;
 wire _0408_;
 wire _0409_;
 wire _0410_;
 wire _0411_;
 wire _0412_;
 wire _0413_;
 wire _0414_;
 wire _0415_;
 wire _0416_;
 wire _0417_;
 wire _0418_;
 wire _0419_;
 wire _0420_;
 wire _0421_;
 wire _0422_;
 wire _0423_;
 wire _0424_;
 wire _0425_;
 wire _0426_;
 wire _0427_;
 wire _0428_;
 wire _0429_;
 wire _0430_;
 wire _0431_;
 wire _0432_;
 wire _0433_;
 wire _0434_;
 wire _0435_;
 wire _0436_;
 wire _0437_;
 wire _0438_;
 wire _0439_;
 wire _0440_;
 wire _0441_;
 wire _0442_;
 wire _0443_;
 wire _0444_;
 wire _0445_;
 wire _0446_;
 wire _0447_;
 wire _0448_;
 wire _0449_;
 wire _0450_;
 wire _0451_;
 wire _0452_;
 wire _0453_;
 wire _0454_;
 wire _0455_;
 wire _0456_;
 wire _0457_;
 wire _0458_;
 wire _0459_;
 wire _0460_;
 wire _0461_;
 wire _0462_;
 wire _0463_;
 wire _0464_;
 wire _0465_;
 wire _0466_;
 wire _0467_;
 wire _0468_;
 wire _0469_;
 wire _0470_;
 wire _0471_;
 wire _0472_;
 wire _0473_;
 wire _0474_;
 wire _0475_;
 wire _0476_;
 wire _0477_;
 wire _0478_;
 wire _0479_;
 wire _0480_;
 wire _0481_;
 wire _0482_;
 wire _0483_;
 wire _0484_;
 wire _0485_;
 wire _0486_;
 wire _0487_;
 wire _0488_;
 wire _0489_;
 wire _0490_;
 wire _0491_;
 wire _0492_;
 wire _0493_;
 wire _0494_;
 wire _0495_;
 wire _0496_;
 wire _0497_;
 wire _0498_;
 wire _0499_;
 wire _0500_;
 wire _0501_;
 wire _0502_;
 wire _0503_;
 wire _0504_;
 wire _0505_;
 wire _0506_;
 wire _0507_;
 wire _0508_;
 wire _0509_;
 wire _0510_;
 wire _0511_;
 wire _0512_;
 wire _0513_;
 wire _0514_;
 wire _0515_;
 wire _0516_;
 wire _0517_;
 wire _0518_;
 wire _0519_;
 wire _0520_;
 wire _0521_;
 wire _0522_;
 wire _0523_;
 wire _0524_;
 wire _0525_;
 wire _0526_;
 wire _0527_;
 wire _0528_;
 wire _0529_;
 wire _0530_;
 wire _0531_;
 wire _0532_;
 wire _0533_;
 wire _0534_;
 wire _0535_;
 wire _0536_;
 wire _0537_;
 wire _0538_;
 wire _0539_;
 wire _0540_;
 wire _0541_;
 wire _0542_;
 wire _0543_;
 wire _0544_;
 wire _0545_;
 wire _0546_;
 wire _0547_;
 wire _0548_;
 wire _0549_;
 wire _0550_;
 wire _0551_;
 wire _0552_;
 wire _0553_;
 wire _0554_;
 wire _0555_;
 wire _0556_;
 wire _0557_;
 wire _0558_;
 wire _0559_;
 wire _0560_;
 wire _0561_;
 wire _0562_;
 wire _0563_;
 wire _0564_;
 wire _0565_;
 wire _0566_;
 wire _0567_;
 wire _0568_;
 wire _0569_;
 wire _0570_;
 wire _0571_;
 wire _0572_;
 wire _0573_;
 wire _0574_;
 wire _0575_;
 wire _0576_;
 wire _0577_;
 wire _0578_;
 wire _0579_;
 wire _0580_;
 wire _0581_;
 wire _0582_;
 wire _0583_;
 wire _0584_;
 wire _0585_;
 wire _0586_;
 wire _0587_;
 wire _0588_;
 wire _0589_;
 wire _0590_;
 wire _0591_;
 wire _0592_;
 wire _0593_;
 wire _0594_;
 wire _0595_;
 wire _0596_;
 wire _0597_;
 wire _0598_;
 wire _0599_;
 wire _0600_;
 wire _0601_;
 wire _0602_;
 wire _0603_;
 wire _0604_;
 wire _0605_;
 wire _0606_;
 wire _0607_;
 wire _0608_;
 wire _0609_;
 wire _0610_;
 wire _0611_;
 wire _0612_;
 wire _0613_;
 wire _0614_;
 wire _0615_;
 wire _0616_;
 wire _0617_;
 wire _0618_;
 wire _0619_;
 wire _0620_;
 wire _0621_;
 wire _0622_;
 wire _0623_;
 wire _0624_;
 wire _0625_;
 wire _0626_;
 wire _0627_;
 wire _0628_;
 wire _0629_;
 wire _0630_;
 wire _0631_;
 wire _0632_;
 wire _0633_;
 wire _0634_;
 wire _0635_;
 wire _0636_;
 wire _0637_;
 wire _0638_;
 wire _0639_;
 wire _0640_;
 wire _0641_;
 wire _0642_;
 wire _0643_;
 wire _0644_;
 wire _0645_;
 wire _0646_;
 wire _0647_;
 wire _0648_;
 wire _0649_;
 wire _0650_;
 wire _0651_;
 wire _0652_;
 wire _0653_;
 wire _0654_;
 wire _0655_;
 wire _0656_;
 wire _0657_;
 wire _0658_;
 wire _0659_;
 wire _0660_;
 wire _0661_;
 wire _0662_;
 wire _0663_;
 wire _0664_;
 wire _0665_;
 wire _0666_;
 wire _0667_;
 wire _0668_;
 wire _0669_;
 wire _0670_;
 wire _0671_;
 wire _0672_;
 wire _0673_;
 wire _0674_;
 wire _0675_;
 wire _0676_;
 wire _0677_;
 wire _0678_;
 wire _0679_;
 wire _0680_;
 wire _0681_;
 wire _0682_;
 wire _0683_;
 wire _0684_;
 wire _0685_;
 wire _0686_;
 wire _0687_;
 wire _0688_;
 wire _0689_;
 wire _0690_;
 wire _0691_;
 wire _0692_;
 wire _0693_;
 wire _0694_;
 wire _0695_;
 wire _0696_;
 wire _0697_;
 wire _0698_;
 wire _0699_;
 wire _0700_;
 wire _0701_;
 wire _0702_;
 wire _0703_;
 wire _0704_;
 wire _0705_;
 wire _0706_;
 wire _0707_;
 wire _0708_;
 wire _0709_;
 wire _0710_;
 wire _0711_;
 wire _0712_;
 wire _0713_;
 wire _0714_;
 wire _0715_;
 wire _0716_;
 wire _0717_;
 wire _0718_;
 wire _0719_;
 wire _0720_;
 wire _0721_;
 wire _0722_;
 wire _0723_;
 wire _0724_;
 wire _0725_;
 wire _0726_;
 wire _0727_;
 wire _0728_;
 wire _0729_;
 wire _0730_;
 wire _0731_;
 wire _0732_;
 wire _0733_;
 wire _0734_;
 wire _0735_;
 wire _0736_;
 wire _0737_;
 wire _0738_;
 wire _0739_;
 wire _0740_;
 wire _0741_;
 wire _0742_;
 wire _0743_;
 wire _0744_;
 wire _0745_;
 wire _0746_;
 wire _0747_;
 wire _0748_;
 wire _0749_;
 wire _0750_;
 wire _0751_;
 wire _0752_;
 wire _0753_;
 wire _0754_;
 wire _0755_;
 wire _0756_;
 wire _0757_;
 wire _0758_;
 wire _0759_;
 wire _0760_;
 wire _0761_;
 wire _0762_;
 wire _0763_;
 wire _0764_;
 wire _0765_;
 wire _0766_;
 wire _0767_;
 wire _0768_;
 wire _0769_;
 wire _0770_;
 wire _0771_;
 wire _0772_;
 wire _0773_;
 wire _0774_;
 wire _0775_;
 wire _0776_;
 wire _0777_;
 wire _0778_;
 wire _0779_;
 wire _0780_;
 wire _0781_;
 wire _0782_;
 wire _0783_;
 wire _0784_;
 wire _0785_;
 wire _0786_;
 wire _0787_;
 wire _0788_;
 wire _0789_;
 wire _0790_;
 wire _0791_;
 wire _0792_;
 wire _0793_;
 wire _0794_;
 wire _0795_;
 wire _0796_;
 wire _0797_;
 wire _0798_;
 wire _0799_;
 wire _0800_;
 wire _0801_;
 wire _0802_;
 wire _0803_;
 wire _0804_;
 wire _0805_;
 wire _0806_;
 wire _0807_;
 wire _0808_;
 wire _0809_;
 wire _0810_;
 wire _0811_;
 wire _0812_;
 wire _0813_;
 wire _0814_;
 wire _0815_;
 wire _0816_;
 wire _0817_;
 wire _0818_;
 wire _0819_;
 wire _0820_;
 wire _0821_;
 wire _0822_;
 wire _0823_;
 wire _0824_;
 wire _0825_;
 wire _0826_;
 wire _0827_;
 wire _0828_;
 wire _0829_;
 wire _0830_;
 wire _0831_;
 wire _0832_;
 wire _0833_;
 wire _0834_;
 wire _0835_;
 wire _0836_;
 wire _0837_;
 wire _0838_;
 wire _0839_;
 wire _0840_;
 wire _0841_;
 wire _0842_;
 wire _0843_;
 wire _0844_;
 wire _0845_;
 wire _0846_;
 wire _0847_;
 wire _0848_;
 wire _0849_;
 wire _0850_;
 wire _0851_;
 wire _0852_;
 wire _0853_;
 wire _0854_;
 wire _0855_;
 wire _0856_;
 wire _0857_;
 wire _0858_;
 wire _0859_;
 wire _0860_;
 wire _0861_;
 wire _0862_;
 wire _0863_;
 wire _0864_;
 wire _0865_;
 wire _0866_;
 wire _0867_;
 wire _0868_;
 wire _0869_;
 wire _0870_;
 wire _0871_;
 wire _0872_;
 wire _0873_;
 wire _0874_;
 wire _0875_;
 wire _0876_;
 wire _0877_;
 wire _0878_;
 wire _0879_;
 wire _0880_;
 wire _0881_;
 wire _0882_;
 wire _0883_;
 wire _0884_;
 wire _0885_;
 wire _0886_;
 wire _0887_;
 wire _0888_;
 wire _0889_;
 wire _0890_;
 wire _0891_;
 wire _0892_;
 wire _0893_;
 wire _0894_;
 wire _0895_;
 wire _0896_;
 wire _0897_;
 wire _0898_;
 wire _0899_;
 wire _0900_;
 wire _0901_;
 wire _0902_;
 wire _0903_;
 wire _0904_;
 wire _0905_;
 wire _0906_;
 wire _0907_;
 wire _0908_;
 wire _0909_;
 wire _0910_;
 wire _0911_;
 wire _0912_;
 wire _0913_;
 wire _0914_;
 wire _0915_;
 wire _0916_;
 wire _0917_;
 wire _0918_;
 wire _0919_;
 wire _0920_;
 wire _0921_;
 wire _0922_;
 wire _0923_;
 wire _0924_;
 wire _0925_;
 wire _0926_;
 wire _0927_;
 wire _0928_;
 wire _0929_;
 wire _0930_;
 wire _0931_;
 wire _0932_;
 wire _0933_;
 wire _0934_;
 wire _0935_;
 wire _0936_;
 wire _0937_;
 wire _0938_;
 wire _0939_;
 wire _0940_;
 wire _0941_;
 wire _0942_;
 wire _0943_;
 wire _0944_;
 wire _0945_;
 wire _0946_;
 wire _0947_;
 wire _0948_;
 wire _0949_;
 wire _0950_;
 wire _0951_;
 wire _0952_;
 wire _0953_;
 wire _0954_;
 wire _0955_;
 wire _0956_;
 wire _0957_;
 wire _0958_;
 wire _0959_;
 wire _0960_;
 wire _0961_;
 wire _0962_;
 wire _0963_;
 wire _0964_;
 wire _0965_;
 wire _0966_;
 wire _0967_;
 wire _0968_;
 wire _0969_;
 wire _0970_;
 wire _0971_;
 wire _0972_;
 wire _0973_;
 wire _0974_;
 wire _0975_;
 wire _0976_;
 wire _0977_;
 wire _0978_;
 wire _0979_;
 wire _0980_;
 wire _0981_;
 wire _0982_;
 wire _0983_;
 wire _0984_;
 wire _0985_;
 wire _0986_;
 wire _0987_;
 wire _0988_;
 wire _0989_;
 wire _0990_;
 wire _0991_;
 wire _0992_;
 wire _0993_;
 wire _0994_;
 wire _0995_;
 wire _0996_;
 wire _0997_;
 wire _0998_;
 wire _0999_;
 wire _1000_;
 wire _1001_;
 wire _1002_;
 wire _1003_;
 wire _1004_;
 wire _1005_;
 wire _1006_;
 wire _1007_;
 wire _1008_;
 wire _1009_;
 wire _1010_;
 wire _1011_;
 wire _1012_;
 wire _1013_;
 wire _1014_;
 wire _1015_;
 wire _1016_;
 wire _1017_;
 wire _1018_;
 wire _1019_;
 wire _1020_;
 wire _1021_;
 wire _1022_;
 wire _1023_;
 wire _1024_;
 wire _1025_;
 wire _1026_;
 wire _1027_;
 wire _1028_;
 wire _1029_;
 wire _1030_;
 wire _1031_;
 wire _1032_;
 wire _1033_;
 wire _1034_;
 wire _1035_;
 wire _1036_;
 wire _1037_;
 wire _1038_;
 wire _1039_;
 wire _1040_;
 wire _1041_;
 wire _1042_;
 wire _1043_;
 wire _1044_;
 wire _1045_;
 wire _1046_;
 wire _1047_;
 wire _1048_;
 wire _1049_;
 wire _1050_;
 wire _1051_;
 wire _1052_;
 wire _1053_;
 wire _1054_;
 wire _1055_;
 wire _1056_;
 wire _1057_;
 wire _1058_;
 wire _1059_;
 wire _1060_;
 wire _1061_;
 wire _1062_;
 wire _1063_;
 wire _1064_;
 wire _1065_;
 wire _1066_;
 wire _1067_;
 wire _1068_;
 wire _1069_;
 wire _1070_;
 wire _1071_;
 wire _1072_;
 wire _1073_;
 wire _1074_;
 wire _1075_;
 wire _1076_;
 wire _1077_;
 wire _1078_;
 wire _1079_;
 wire _1080_;
 wire _1081_;
 wire _1082_;
 wire _1083_;
 wire _1084_;
 wire _1085_;
 wire _1086_;
 wire _1087_;
 wire _1088_;
 wire _1089_;
 wire _1090_;
 wire _1091_;
 wire _1092_;
 wire _1093_;
 wire _1094_;
 wire _1095_;
 wire _1096_;
 wire _1097_;
 wire _1098_;
 wire _1099_;
 wire _1100_;
 wire _1101_;
 wire _1102_;
 wire _1103_;
 wire _1104_;
 wire _1105_;
 wire _1106_;
 wire _1107_;
 wire _1108_;
 wire _1109_;
 wire _1110_;
 wire _1111_;
 wire _1112_;
 wire _1113_;
 wire _1114_;
 wire _1115_;
 wire _1116_;
 wire _1117_;
 wire _1118_;
 wire _1119_;
 wire _1120_;
 wire _1121_;
 wire _1122_;
 wire _1123_;
 wire _1124_;
 wire _1125_;
 wire _1126_;
 wire _1127_;
 wire _1128_;
 wire _1129_;
 wire _1130_;
 wire _1131_;
 wire _1132_;
 wire _1133_;
 wire _1134_;
 wire _1135_;
 wire _1136_;
 wire _1137_;
 wire _1138_;
 wire _1139_;
 wire _1140_;
 wire _1141_;
 wire _1142_;
 wire _1143_;
 wire _1144_;
 wire _1145_;
 wire _1146_;
 wire _1147_;
 wire _1148_;
 wire _1149_;
 wire _1150_;
 wire _1151_;
 wire _1152_;
 wire _1153_;
 wire _1154_;
 wire _1155_;
 wire _1156_;
 wire _1157_;
 wire _1158_;
 wire _1159_;
 wire _1160_;
 wire _1161_;
 wire _1162_;
 wire _1163_;
 wire _1164_;
 wire _1165_;
 wire _1166_;
 wire _1167_;
 wire _1168_;
 wire _1169_;
 wire _1170_;
 wire _1171_;
 wire _1172_;
 wire _1173_;
 wire _1174_;
 wire _1175_;
 wire _1176_;
 wire _1177_;
 wire _1178_;
 wire _1179_;
 wire _1180_;
 wire _1181_;
 wire _1182_;
 wire _1183_;
 wire _1184_;
 wire _1185_;
 wire _1186_;
 wire _1187_;
 wire _1188_;
 wire _1189_;
 wire _1190_;
 wire _1191_;
 wire _1192_;
 wire _1193_;
 wire _1194_;
 wire _1195_;
 wire _1196_;
 wire _1197_;
 wire _1198_;
 wire _1199_;
 wire _1200_;
 wire _1201_;
 wire _1202_;
 wire _1203_;
 wire _1204_;
 wire _1205_;
 wire _1206_;
 wire _1207_;
 wire _1208_;
 wire _1209_;
 wire _1210_;
 wire _1211_;
 wire _1212_;
 wire _1213_;
 wire _1214_;
 wire _1215_;
 wire _1216_;
 wire _1217_;
 wire _1218_;
 wire _1219_;
 wire _1220_;
 wire _1221_;
 wire _1222_;
 wire _1223_;
 wire _1224_;
 wire _1225_;
 wire _1226_;
 wire _1227_;
 wire _1228_;
 wire _1229_;
 wire _1230_;
 wire _1231_;
 wire _1232_;
 wire _1233_;
 wire _1234_;
 wire _1235_;
 wire _1236_;
 wire _1237_;
 wire _1238_;
 wire _1239_;
 wire _1240_;
 wire _1241_;
 wire _1242_;
 wire _1243_;
 wire _1244_;
 wire _1245_;
 wire _1246_;
 wire _1247_;
 wire _1248_;
 wire _1249_;
 wire _1250_;
 wire _1251_;
 wire _1252_;
 wire _1253_;
 wire _1254_;
 wire _1255_;
 wire _1256_;
 wire _1257_;
 wire _1258_;
 wire _1259_;
 wire _1260_;
 wire _1261_;
 wire _1262_;
 wire _1263_;
 wire _1264_;
 wire _1265_;
 wire _1266_;
 wire _1267_;
 wire _1268_;
 wire _1269_;
 wire _1270_;
 wire _1271_;
 wire _1272_;
 wire _1273_;
 wire _1274_;
 wire _1275_;
 wire _1276_;
 wire _1277_;
 wire _1278_;
 wire _1279_;
 wire _1280_;
 wire _1281_;
 wire _1282_;
 wire _1283_;
 wire _1284_;
 wire _1285_;
 wire _1286_;
 wire _1287_;
 wire _1288_;
 wire _1289_;
 wire _1290_;
 wire _1291_;
 wire _1292_;
 wire _1293_;
 wire _1294_;
 wire _1295_;
 wire _1296_;
 wire _1297_;
 wire _1298_;
 wire _1299_;
 wire _1300_;
 wire _1301_;
 wire _1302_;
 wire _1303_;
 wire _1304_;
 wire _1305_;
 wire _1306_;
 wire _1307_;
 wire _1308_;
 wire _1309_;
 wire _1310_;
 wire _1311_;
 wire _1312_;
 wire _1313_;
 wire _1314_;
 wire _1315_;
 wire _1316_;
 wire _1317_;
 wire _1318_;
 wire _1319_;
 wire _1320_;
 wire _1321_;
 wire _1322_;
 wire _1323_;
 wire _1324_;
 wire _1325_;
 wire _1326_;
 wire _1327_;
 wire _1328_;
 wire _1329_;
 wire _1330_;
 wire _1331_;
 wire _1332_;
 wire _1333_;
 wire _1334_;
 wire _1335_;
 wire _1336_;
 wire _1337_;
 wire _1338_;
 wire _1339_;
 wire _1340_;
 wire _1341_;
 wire _1342_;
 wire _1343_;
 wire _1344_;
 wire _1345_;
 wire _1346_;
 wire _1347_;
 wire _1348_;
 wire _1349_;
 wire _1350_;
 wire _1351_;
 wire _1352_;
 wire _1353_;
 wire _1354_;
 wire _1355_;
 wire _1356_;
 wire _1357_;
 wire _1358_;
 wire _1359_;
 wire _1360_;
 wire _1361_;
 wire _1362_;
 wire _1363_;
 wire _1364_;
 wire _1365_;
 wire _1366_;
 wire _1367_;
 wire _1368_;
 wire _1369_;
 wire _1370_;
 wire _1371_;
 wire _1372_;
 wire _1373_;
 wire _1374_;
 wire _1375_;
 wire _1376_;
 wire _1377_;
 wire _1378_;
 wire _1379_;
 wire _1380_;
 wire _1381_;
 wire _1382_;
 wire _1383_;
 wire _1384_;
 wire _1385_;
 wire _1386_;
 wire _1387_;
 wire _1388_;
 wire _1389_;
 wire _1390_;
 wire _1391_;
 wire _1392_;
 wire _1393_;
 wire _1394_;
 wire _1395_;
 wire _1396_;
 wire _1397_;
 wire _1398_;
 wire _1399_;
 wire _1400_;
 wire _1401_;
 wire _1402_;
 wire _1403_;
 wire _1404_;
 wire _1405_;
 wire _1406_;
 wire _1407_;
 wire _1408_;
 wire _1409_;
 wire _1410_;
 wire _1411_;
 wire _1412_;
 wire _1413_;
 wire _1414_;
 wire _1415_;
 wire _1416_;
 wire _1417_;
 wire _1418_;
 wire _1419_;
 wire _1420_;
 wire _1421_;
 wire _1422_;
 wire _1423_;
 wire _1424_;
 wire _1425_;
 wire _1426_;
 wire _1427_;
 wire _1428_;
 wire _1429_;
 wire _1430_;
 wire _1431_;
 wire _1432_;
 wire _1433_;
 wire _1434_;
 wire _1435_;
 wire _1436_;
 wire _1437_;
 wire _1438_;
 wire _1439_;
 wire _1440_;
 wire _1441_;
 wire _1442_;
 wire _1443_;
 wire _1444_;
 wire _1445_;
 wire _1446_;
 wire _1447_;
 wire _1448_;
 wire _1449_;
 wire _1450_;
 wire _1451_;
 wire _1452_;
 wire _1453_;
 wire _1454_;
 wire _1455_;
 wire _1456_;
 wire _1457_;
 wire _1458_;
 wire _1459_;
 wire _1460_;
 wire _1461_;
 wire _1462_;
 wire _1463_;
 wire _1464_;
 wire _1465_;
 wire _1466_;
 wire _1467_;
 wire _1468_;
 wire _1469_;
 wire _1470_;
 wire _1471_;
 wire _1472_;
 wire _1473_;
 wire _1474_;
 wire _1475_;
 wire _1476_;
 wire _1477_;
 wire _1478_;
 wire _1479_;
 wire _1480_;
 wire _1481_;
 wire _1482_;
 wire _1483_;
 wire _1484_;
 wire _1485_;
 wire _1486_;
 wire _1487_;
 wire _1488_;
 wire _1489_;
 wire _1490_;
 wire _1491_;
 wire _1492_;
 wire _1493_;
 wire _1494_;
 wire _1495_;
 wire _1496_;
 wire _1497_;
 wire _1498_;
 wire _1499_;
 wire _1500_;
 wire _1501_;
 wire _1502_;
 wire _1503_;
 wire _1504_;
 wire _1505_;
 wire _1506_;
 wire _1507_;
 wire _1508_;
 wire _1509_;
 wire _1510_;
 wire _1511_;
 wire _1512_;
 wire _1513_;
 wire _1514_;
 wire _1515_;
 wire _1516_;
 wire _1517_;
 wire _1518_;
 wire _1519_;
 wire _1520_;
 wire _1521_;
 wire _1522_;
 wire _1523_;
 wire _1524_;
 wire _1525_;
 wire _1526_;
 wire _1527_;
 wire _1528_;
 wire _1529_;
 wire _1530_;
 wire _1531_;
 wire _1532_;
 wire _1533_;
 wire _1534_;
 wire _1535_;
 wire _1536_;
 wire _1537_;
 wire _1538_;
 wire _1539_;
 wire _1540_;
 wire _1541_;
 wire _1542_;
 wire _1543_;
 wire _1544_;
 wire _1545_;
 wire _1546_;
 wire _1547_;
 wire _1548_;
 wire _1549_;
 wire _1550_;
 wire _1551_;
 wire _1552_;
 wire _1553_;
 wire _1554_;
 wire _1555_;
 wire _1556_;
 wire _1557_;
 wire _1558_;
 wire _1559_;
 wire _1560_;
 wire _1561_;
 wire _1562_;
 wire _1563_;
 wire _1564_;
 wire _1565_;
 wire _1566_;
 wire _1567_;
 wire _1568_;
 wire _1569_;
 wire _1570_;
 wire _1571_;
 wire _1572_;
 wire _1573_;
 wire _1574_;
 wire _1575_;
 wire _1576_;
 wire _1577_;
 wire _1578_;
 wire _1579_;
 wire _1580_;
 wire _1581_;
 wire _1582_;
 wire _1583_;
 wire _1584_;
 wire _1585_;
 wire _1586_;
 wire _1587_;
 wire _1588_;
 wire _1589_;
 wire _1590_;
 wire _1591_;
 wire _1592_;
 wire _1593_;
 wire _1594_;
 wire _1595_;
 wire _1596_;
 wire _1597_;
 wire _1598_;
 wire _1599_;
 wire _1600_;
 wire _1601_;
 wire _1602_;
 wire _1603_;
 wire _1604_;
 wire _1605_;
 wire _1606_;
 wire _1607_;
 wire _1608_;
 wire _1609_;
 wire _1610_;
 wire _1611_;
 wire _1612_;
 wire _1613_;
 wire _1614_;
 wire _1615_;
 wire _1616_;
 wire _1617_;
 wire _1618_;
 wire _1619_;
 wire _1620_;
 wire _1621_;
 wire _1622_;
 wire _1623_;
 wire _1624_;
 wire _1625_;
 wire _1626_;
 wire _1627_;
 wire _1628_;
 wire _1629_;
 wire _1630_;
 wire _1631_;
 wire _1632_;
 wire _1633_;
 wire _1634_;
 wire _1635_;
 wire _1636_;
 wire _1637_;
 wire _1638_;
 wire _1639_;
 wire _1640_;
 wire _1641_;
 wire _1642_;
 wire _1643_;
 wire _1644_;
 wire _1645_;
 wire _1646_;
 wire _1647_;
 wire _1648_;
 wire _1649_;
 wire _1650_;
 wire _1651_;
 wire _1652_;
 wire _1653_;
 wire _1654_;
 wire _1655_;
 wire _1656_;
 wire _1657_;
 wire _1658_;
 wire _1659_;
 wire _1660_;
 wire _1661_;
 wire _1662_;
 wire _1663_;
 wire _1664_;
 wire _1665_;
 wire _1666_;
 wire _1667_;
 wire _1668_;
 wire _1669_;
 wire _1670_;
 wire _1671_;
 wire _1672_;
 wire _1673_;
 wire _1674_;
 wire _1675_;
 wire _1676_;
 wire _1677_;
 wire _1678_;
 wire _1679_;
 wire _1680_;
 wire _1681_;
 wire _1682_;
 wire _1683_;
 wire _1684_;
 wire _1685_;
 wire _1686_;
 wire _1687_;
 wire _1688_;
 wire _1689_;
 wire _1690_;
 wire _1691_;
 wire _1692_;
 wire _1693_;
 wire _1694_;
 wire _1695_;
 wire _1696_;
 wire _1697_;
 wire _1698_;
 wire _1699_;
 wire _1700_;
 wire _1701_;
 wire _1702_;
 wire _1703_;
 wire _1704_;
 wire _1705_;
 wire _1706_;
 wire _1707_;
 wire _1708_;
 wire _1709_;
 wire _1710_;
 wire _1711_;
 wire _1712_;
 wire _1713_;
 wire _1714_;
 wire _1715_;
 wire _1716_;
 wire _1717_;
 wire _1718_;
 wire _1719_;
 wire _1720_;
 wire _1721_;
 wire _1722_;
 wire _1723_;
 wire _1724_;
 wire _1725_;
 wire _1726_;
 wire _1727_;
 wire _1728_;
 wire _1729_;
 wire _1730_;
 wire _1731_;
 wire _1732_;
 wire _1733_;
 wire _1734_;
 wire _1735_;
 wire _1736_;
 wire _1737_;
 wire _1738_;
 wire _1739_;
 wire _1740_;
 wire _1741_;
 wire _1742_;
 wire _1743_;
 wire _1744_;
 wire _1745_;
 wire _1746_;
 wire _1747_;
 wire _1748_;
 wire _1749_;
 wire _1750_;
 wire _1751_;
 wire _1752_;
 wire _1753_;
 wire _1754_;
 wire _1755_;
 wire _1756_;
 wire _1757_;
 wire _1758_;
 wire _1759_;
 wire _1760_;
 wire _1761_;
 wire _1762_;
 wire _1763_;
 wire _1764_;
 wire _1765_;
 wire _1766_;
 wire _1767_;
 wire _1768_;
 wire _1769_;
 wire _1770_;
 wire _1771_;
 wire _1772_;
 wire _1773_;
 wire _1774_;
 wire _1775_;
 wire _1776_;
 wire _1777_;
 wire _1778_;
 wire _1779_;
 wire _1780_;
 wire _1781_;
 wire _1782_;
 wire _1783_;
 wire _1784_;
 wire _1785_;
 wire _1786_;
 wire _1787_;
 wire _1788_;
 wire _1789_;
 wire _1790_;
 wire _1791_;
 wire _1792_;
 wire _1793_;
 wire _1794_;
 wire _1795_;
 wire _1796_;
 wire _1797_;
 wire _1798_;
 wire _1799_;
 wire _1800_;
 wire _1801_;
 wire _1802_;
 wire _1803_;
 wire _1804_;
 wire _1805_;
 wire _1806_;
 wire _1807_;
 wire _1808_;
 wire _1809_;
 wire _1810_;
 wire _1811_;
 wire _1812_;
 wire _1813_;
 wire _1814_;
 wire _1815_;
 wire _1816_;
 wire _1817_;
 wire _1818_;
 wire _1819_;
 wire _1820_;
 wire _1821_;
 wire _1822_;
 wire _1823_;
 wire _1824_;
 wire _1825_;
 wire _1826_;
 wire _1827_;
 wire _1828_;
 wire _1829_;
 wire _1830_;
 wire _1831_;
 wire _1832_;
 wire _1833_;
 wire _1834_;
 wire _1835_;
 wire _1836_;
 wire _1837_;
 wire _1838_;
 wire _1839_;
 wire _1840_;
 wire _1841_;
 wire _1842_;
 wire _1843_;
 wire _1844_;
 wire _1845_;
 wire _1846_;
 wire _1847_;
 wire _1848_;
 wire _1849_;
 wire _1850_;
 wire _1851_;
 wire _1852_;
 wire _1853_;
 wire _1854_;
 wire _1855_;
 wire _1856_;
 wire _1857_;
 wire _1858_;
 wire _1859_;
 wire _1860_;
 wire _1861_;
 wire _1862_;
 wire _1863_;
 wire _1864_;
 wire _1865_;
 wire _1866_;
 wire _1867_;
 wire _1868_;
 wire _1869_;
 wire _1870_;
 wire _1871_;
 wire _1872_;
 wire _1873_;
 wire _1874_;
 wire _1875_;
 wire _1876_;
 wire _1877_;
 wire _1878_;
 wire _1879_;
 wire _1880_;
 wire _1881_;
 wire _1882_;
 wire _1883_;
 wire _1884_;
 wire _1885_;
 wire _1886_;
 wire _1887_;
 wire _1888_;
 wire _1889_;
 wire _1890_;
 wire _1891_;
 wire _1892_;
 wire _1893_;
 wire _1894_;
 wire _1895_;
 wire _1896_;
 wire _1897_;
 wire _1898_;
 wire _1899_;
 wire _1900_;
 wire _1901_;
 wire _1902_;
 wire _1903_;
 wire _1904_;
 wire _1905_;
 wire _1906_;
 wire _1907_;
 wire _1908_;
 wire _1909_;
 wire _1910_;
 wire _1911_;
 wire _1912_;
 wire _1913_;
 wire _1914_;
 wire _1915_;
 wire _1916_;
 wire _1917_;
 wire _1918_;
 wire _1919_;
 wire _1920_;
 wire _1921_;
 wire _1922_;
 wire _1923_;
 wire _1924_;
 wire _1925_;
 wire _1926_;
 wire _1927_;
 wire _1928_;
 wire _1929_;
 wire _1930_;
 wire _1931_;
 wire _1932_;
 wire _1933_;
 wire _1934_;
 wire _1935_;
 wire _1936_;
 wire _1937_;
 wire _1938_;
 wire _1939_;
 wire _1940_;
 wire _1941_;
 wire _1942_;
 wire _1943_;
 wire _1944_;
 wire _1945_;
 wire _1946_;
 wire _1947_;
 wire _1948_;
 wire _1949_;
 wire _1950_;
 wire _1951_;
 wire _1952_;
 wire _1953_;
 wire _1954_;
 wire _1955_;
 wire _1956_;
 wire _1957_;
 wire _1958_;
 wire _1959_;
 wire _1960_;
 wire _1961_;
 wire _1962_;
 wire _1963_;
 wire _1964_;
 wire _1965_;
 wire _1966_;
 wire _1967_;
 wire _1968_;
 wire _1969_;
 wire _1970_;
 wire _1971_;
 wire _1972_;
 wire _1973_;
 wire _1974_;
 wire _1975_;
 wire _1976_;
 wire _1977_;
 wire _1978_;
 wire _1979_;
 wire _1980_;
 wire _1981_;
 wire _1982_;
 wire _1983_;
 wire _1984_;
 wire _1985_;
 wire _1986_;
 wire _1987_;
 wire _1988_;
 wire _1989_;
 wire _1990_;
 wire _1991_;
 wire _1992_;
 wire _1993_;
 wire _1994_;
 wire _1995_;
 wire _1996_;
 wire _1997_;
 wire _1998_;
 wire _1999_;
 wire _2000_;
 wire _2001_;
 wire _2002_;
 wire _2003_;
 wire _2004_;
 wire _2005_;
 wire _2006_;
 wire _2007_;
 wire _2008_;
 wire _2009_;
 wire _2010_;
 wire _2011_;
 wire _2012_;
 wire _2013_;
 wire _2014_;
 wire _2015_;
 wire _2016_;
 wire _2017_;
 wire _2018_;
 wire _2019_;
 wire _2020_;
 wire _2021_;
 wire _2022_;
 wire _2023_;
 wire _2024_;
 wire _2025_;
 wire _2026_;
 wire _2027_;
 wire _2028_;
 wire _2029_;
 wire _2030_;
 wire _2031_;
 wire _2032_;
 wire _2033_;
 wire _2034_;
 wire _2035_;
 wire _2036_;
 wire _2037_;
 wire _2038_;
 wire _2039_;
 wire _2040_;
 wire _2041_;
 wire _2042_;
 wire _2043_;
 wire _2044_;
 wire _2045_;
 wire _2046_;
 wire _2047_;
 wire _2048_;
 wire _2049_;
 wire _2050_;
 wire _2051_;
 wire _2052_;
 wire _2053_;
 wire _2054_;
 wire _2055_;
 wire _2056_;
 wire _2057_;
 wire _2058_;
 wire _2059_;
 wire _2060_;
 wire _2061_;
 wire _2062_;
 wire _2063_;
 wire _2064_;
 wire _2065_;
 wire _2066_;
 wire _2067_;
 wire _2068_;
 wire _2069_;
 wire _2070_;
 wire _2071_;
 wire _2072_;
 wire _2073_;
 wire _2074_;
 wire _2075_;
 wire _2076_;
 wire _2077_;
 wire _2078_;
 wire _2079_;
 wire _2080_;
 wire _2081_;
 wire _2082_;
 wire _2083_;
 wire _2084_;
 wire _2085_;
 wire _2086_;
 wire _2087_;
 wire _2088_;
 wire _2089_;
 wire _2090_;
 wire _2091_;
 wire _2092_;
 wire _2093_;
 wire _2094_;
 wire _2095_;
 wire _2096_;
 wire _2097_;
 wire _2098_;
 wire _2099_;
 wire _2100_;
 wire _2101_;
 wire _2102_;
 wire _2103_;
 wire _2104_;
 wire _2105_;
 wire _2106_;
 wire _2107_;
 wire _2108_;
 wire _2109_;
 wire _2110_;
 wire _2111_;
 wire _2112_;
 wire _2113_;
 wire _2114_;
 wire _2115_;
 wire _2116_;
 wire _2117_;
 wire _2118_;
 wire _2119_;
 wire _2120_;
 wire _2121_;
 wire _2122_;
 wire _2123_;
 wire _2124_;
 wire _2125_;
 wire _2126_;
 wire _2127_;
 wire _2128_;
 wire _2129_;
 wire _2130_;
 wire _2131_;
 wire _2132_;
 wire _2133_;
 wire _2134_;
 wire _2135_;
 wire _2136_;
 wire _2137_;
 wire _2138_;
 wire _2139_;
 wire _2140_;
 wire _2141_;
 wire _2142_;
 wire _2143_;
 wire _2144_;
 wire _2145_;
 wire _2146_;
 wire _2147_;
 wire _2148_;
 wire _2149_;
 wire _2150_;
 wire _2151_;
 wire _2152_;
 wire _2153_;
 wire _2154_;
 wire _2155_;
 wire _2156_;
 wire _2157_;
 wire _2158_;
 wire _2159_;
 wire _2160_;
 wire _2161_;
 wire _2162_;
 wire _2163_;
 wire _2164_;
 wire _2165_;
 wire _2166_;
 wire _2167_;
 wire _2168_;
 wire _2169_;
 wire _2170_;
 wire _2171_;
 wire _2172_;
 wire _2173_;
 wire _2174_;
 wire _2175_;
 wire _2176_;
 wire _2177_;
 wire _2178_;
 wire _2179_;
 wire _2180_;
 wire _2181_;
 wire _2182_;
 wire _2183_;
 wire _2184_;
 wire _2185_;
 wire _2186_;
 wire _2187_;
 wire _2188_;
 wire _2189_;
 wire _2190_;
 wire _2191_;
 wire _2192_;
 wire _2193_;
 wire _2194_;
 wire _2195_;
 wire _2196_;
 wire _2197_;
 wire _2198_;
 wire _2199_;
 wire _2200_;
 wire _2201_;
 wire _2202_;
 wire _2203_;
 wire _2204_;
 wire _2205_;
 wire _2206_;
 wire _2207_;
 wire _2208_;
 wire _2209_;
 wire _2210_;
 wire _2211_;
 wire _2212_;
 wire _2213_;
 wire _2214_;
 wire _2215_;
 wire _2216_;
 wire _2217_;
 wire _2218_;
 wire _2219_;
 wire _2220_;
 wire _2221_;
 wire _2222_;
 wire _2223_;
 wire _2224_;
 wire _2225_;
 wire _2226_;
 wire clknet_0_clk;
 wire net151;
 wire b0;
 wire g0;
 wire hs;
 wire \vga.ball_angle[0] ;
 wire \vga.ball_angle[1] ;
 wire \vga.ball_angle[2] ;
 wire \vga.ball_angle[3] ;
 wire \vga.ball_motion_l ;
 wire \vga.ball_pos_h[0] ;
 wire \vga.ball_pos_h[1] ;
 wire \vga.ball_pos_h[2] ;
 wire \vga.ball_pos_h[3] ;
 wire \vga.ball_pos_h[4] ;
 wire \vga.ball_pos_h[5] ;
 wire \vga.ball_pos_h[6] ;
 wire \vga.ball_pos_h[7] ;
 wire \vga.ball_pos_h[8] ;
 wire \vga.ball_pos_h[9] ;
 wire \vga.ball_pos_v[0] ;
 wire \vga.ball_pos_v[1] ;
 wire \vga.ball_pos_v[2] ;
 wire \vga.ball_pos_v[3] ;
 wire \vga.ball_pos_v[4] ;
 wire \vga.ball_pos_v[5] ;
 wire \vga.ball_pos_v[6] ;
 wire \vga.ball_pos_v[7] ;
 wire \vga.ball_pos_v[8] ;
 wire \vga.ball_ratio[0] ;
 wire \vga.ball_ratio[1] ;
 wire \vga.ball_ratio[2] ;
 wire \vga.blank_h ;
 wire \vga.blank_v ;
 wire \vga.count_h[0] ;
 wire \vga.count_h[1] ;
 wire \vga.count_h[2] ;
 wire \vga.count_h[3] ;
 wire \vga.count_h[4] ;
 wire \vga.count_h[5] ;
 wire \vga.count_h[6] ;
 wire \vga.count_h[7] ;
 wire \vga.count_h[8] ;
 wire \vga.count_h[9] ;
 wire \vga.count_v[0] ;
 wire \vga.count_v[1] ;
 wire \vga.count_v[2] ;
 wire \vga.count_v[3] ;
 wire \vga.count_v[4] ;
 wire \vga.count_v[5] ;
 wire \vga.count_v[6] ;
 wire \vga.count_v[7] ;
 wire \vga.count_v[8] ;
 wire \vga.count_v[9] ;
 wire \vga.hs_out ;
 wire \vga.interval_counter[0] ;
 wire \vga.interval_counter[10] ;
 wire \vga.interval_counter[11] ;
 wire \vga.interval_counter[12] ;
 wire \vga.interval_counter[13] ;
 wire \vga.interval_counter[14] ;
 wire \vga.interval_counter[15] ;
 wire \vga.interval_counter[16] ;
 wire \vga.interval_counter[17] ;
 wire \vga.interval_counter[18] ;
 wire \vga.interval_counter[19] ;
 wire \vga.interval_counter[1] ;
 wire \vga.interval_counter[20] ;
 wire \vga.interval_counter[21] ;
 wire \vga.interval_counter[22] ;
 wire \vga.interval_counter[23] ;
 wire \vga.interval_counter[24] ;
 wire \vga.interval_counter[2] ;
 wire \vga.interval_counter[3] ;
 wire \vga.interval_counter[4] ;
 wire \vga.interval_counter[5] ;
 wire \vga.interval_counter[6] ;
 wire \vga.interval_counter[7] ;
 wire \vga.interval_counter[8] ;
 wire \vga.interval_counter[9] ;
 wire \vga.left_down_1d ;
 wire \vga.left_down_pressed ;
 wire \vga.left_up_1d ;
 wire \vga.left_up_pressed ;
 wire \vga.paddle_l_pos_v[0] ;
 wire \vga.paddle_l_pos_v[1] ;
 wire \vga.paddle_l_pos_v[2] ;
 wire \vga.paddle_l_pos_v[3] ;
 wire \vga.paddle_l_pos_v[4] ;
 wire \vga.paddle_l_pos_v[5] ;
 wire \vga.paddle_l_pos_v[6] ;
 wire \vga.paddle_l_pos_v[7] ;
 wire \vga.paddle_l_pos_v[8] ;
 wire \vga.paddle_r_pos_v[0] ;
 wire \vga.paddle_r_pos_v[1] ;
 wire \vga.paddle_r_pos_v[2] ;
 wire \vga.paddle_r_pos_v[3] ;
 wire \vga.paddle_r_pos_v[4] ;
 wire \vga.paddle_r_pos_v[5] ;
 wire \vga.paddle_r_pos_v[6] ;
 wire \vga.paddle_r_pos_v[7] ;
 wire \vga.paddle_r_pos_v[8] ;
 wire \vga.right_down_1d ;
 wire \vga.right_down_pressed ;
 wire \vga.right_up_1d ;
 wire \vga.right_up_pressed ;
 wire \vga.score_l[0] ;
 wire \vga.score_l[1] ;
 wire \vga.score_l[2] ;
 wire \vga.score_l[3] ;
 wire \vga.score_l[4] ;
 wire \vga.score_l_ten_enable ;
 wire \vga.score_l_unit_pixels[0] ;
 wire \vga.score_l_unit_pixels[1] ;
 wire \vga.score_l_unit_pixels[2] ;
 wire \vga.score_r[0] ;
 wire \vga.score_r[1] ;
 wire \vga.score_r[2] ;
 wire \vga.score_r[3] ;
 wire \vga.score_r[4] ;
 wire \vga.score_r_ten_enable ;
 wire \vga.score_r_unit_pixels[0] ;
 wire \vga.score_r_unit_pixels[1] ;
 wire \vga.score_r_unit_pixels[2] ;
 wire \vga.speed_lsb_1d ;
 wire \vga.speed_msb_1d ;
 wire \vga.vs ;
 wire \vga.vs_out ;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net150;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net180;
 wire net181;
 wire net182;
 wire net183;
 wire net184;
 wire net185;
 wire net186;
 wire net187;
 wire net188;
 wire net189;
 wire net190;
 wire net191;
 wire net192;
 wire net193;
 wire net194;
 wire net195;
 wire net196;
 wire net197;
 wire net198;
 wire net199;
 wire net200;
 wire net201;
 wire net202;
 wire net203;
 wire net204;
 wire net205;
 wire net206;
 wire net207;
 wire net208;
 wire net209;
 wire net210;
 wire net211;
 wire net212;
 wire net213;
 wire net214;
 wire net215;
 wire net216;
 wire net217;
 wire net218;
 wire net219;
 wire net220;
 wire net221;
 wire net222;
 wire net223;
 wire net224;
 wire net225;
 wire net226;
 wire net227;
 wire net228;
 wire net229;
 wire net230;
 wire net231;
 wire net232;
 wire net233;
 wire net234;
 wire net235;
 wire net236;
 wire net237;
 wire net238;
 wire net239;
 wire net240;
 wire net241;
 wire net242;
 wire net243;
 wire net244;
 wire net245;
 wire net246;
 wire net247;
 wire net248;
 wire net249;
 wire net250;
 wire net251;
 wire net252;
 wire net253;
 wire net254;
 wire net255;
 wire net256;
 wire net257;
 wire net258;
 wire net259;
 wire net260;
 wire net261;
 wire net262;
 wire net263;
 wire net264;
 wire net265;
 wire net266;
 wire net267;
 wire net268;
 wire net269;
 wire net270;
 wire net271;
 wire net272;
 wire net273;
 wire net274;
 wire net275;
 wire net276;
 wire net277;
 wire net278;
 wire net279;
 wire net280;
 wire net281;
 wire net282;
 wire net283;
 wire net284;
 wire net285;
 wire net286;
 wire net287;
 wire net288;
 wire net289;
 wire net290;
 wire net291;
 wire net292;
 wire net293;
 wire net294;
 wire net295;
 wire net296;
 wire clknet_4_0_0_clk;
 wire clknet_4_1_0_clk;
 wire clknet_4_2_0_clk;
 wire clknet_4_3_0_clk;
 wire clknet_4_4_0_clk;
 wire clknet_4_5_0_clk;
 wire clknet_4_6_0_clk;
 wire clknet_4_7_0_clk;
 wire clknet_4_8_0_clk;
 wire clknet_4_9_0_clk;
 wire clknet_4_10_0_clk;
 wire clknet_4_11_0_clk;
 wire clknet_4_12_0_clk;
 wire clknet_4_13_0_clk;
 wire clknet_4_14_0_clk;
 wire clknet_4_15_0_clk;
 wire clknet_5_0__leaf_clk;
 wire clknet_5_1__leaf_clk;
 wire clknet_5_2__leaf_clk;
 wire clknet_5_3__leaf_clk;
 wire clknet_5_4__leaf_clk;
 wire clknet_5_5__leaf_clk;
 wire clknet_5_6__leaf_clk;
 wire clknet_5_7__leaf_clk;
 wire clknet_5_8__leaf_clk;
 wire clknet_5_9__leaf_clk;
 wire clknet_5_10__leaf_clk;
 wire clknet_5_11__leaf_clk;
 wire clknet_5_12__leaf_clk;
 wire clknet_5_13__leaf_clk;
 wire clknet_5_14__leaf_clk;
 wire clknet_5_15__leaf_clk;
 wire clknet_5_16__leaf_clk;
 wire clknet_5_17__leaf_clk;
 wire clknet_5_18__leaf_clk;
 wire clknet_5_19__leaf_clk;
 wire clknet_5_20__leaf_clk;
 wire clknet_5_21__leaf_clk;
 wire clknet_5_22__leaf_clk;
 wire clknet_5_23__leaf_clk;
 wire clknet_5_24__leaf_clk;
 wire clknet_5_25__leaf_clk;
 wire clknet_5_26__leaf_clk;
 wire clknet_5_27__leaf_clk;
 wire clknet_5_28__leaf_clk;
 wire clknet_5_29__leaf_clk;
 wire clknet_5_30__leaf_clk;
 wire clknet_5_31__leaf_clk;

 sg13g2_buf_1 _2229_ (.A(\vga.score_l[3] ),
    .X(_1505_));
 sg13g2_and2_1 _2230_ (.A(net148),
    .B(\vga.score_l[4] ),
    .X(_1506_));
 sg13g2_buf_1 _2231_ (.A(_0072_),
    .X(_1507_));
 sg13g2_buf_1 _2232_ (.A(\vga.paddle_r_pos_v[1] ),
    .X(_1508_));
 sg13g2_inv_1 _2233_ (.Y(_1509_),
    .A(_1508_));
 sg13g2_buf_1 _2234_ (.A(\vga.ball_pos_v[1] ),
    .X(_1510_));
 sg13g2_buf_1 _2235_ (.A(\vga.ball_pos_v[0] ),
    .X(_1511_));
 sg13g2_buf_1 _2236_ (.A(\vga.paddle_r_pos_v[0] ),
    .X(_1512_));
 sg13g2_nand2b_1 _2237_ (.Y(_1513_),
    .B(_1512_),
    .A_N(net146));
 sg13g2_a21o_1 _2238_ (.A2(_1510_),
    .A1(_1509_),
    .B1(_1513_),
    .X(_1514_));
 sg13g2_buf_8 _2239_ (.A(\vga.paddle_r_pos_v[2] ),
    .X(_1515_));
 sg13g2_buf_1 _2240_ (.A(_1515_),
    .X(_1516_));
 sg13g2_inv_2 _2241_ (.Y(_1517_),
    .A(net116));
 sg13g2_buf_1 _2242_ (.A(\vga.ball_pos_v[2] ),
    .X(_1518_));
 sg13g2_inv_1 _2243_ (.Y(_1519_),
    .A(net145));
 sg13g2_inv_1 _2244_ (.Y(_1520_),
    .A(_1510_));
 sg13g2_a22oi_1 _2245_ (.Y(_1521_),
    .B1(_1520_),
    .B2(_1508_),
    .A2(_1519_),
    .A1(_1517_));
 sg13g2_buf_8 _2246_ (.A(\vga.paddle_r_pos_v[3] ),
    .X(_1522_));
 sg13g2_buf_1 _2247_ (.A(net144),
    .X(_1523_));
 sg13g2_buf_2 _2248_ (.A(\vga.ball_pos_v[3] ),
    .X(_1524_));
 sg13g2_inv_2 _2249_ (.Y(_1525_),
    .A(_1524_));
 sg13g2_o21ai_1 _2250_ (.B1(_1519_),
    .Y(_1526_),
    .A1(net115),
    .A2(_1525_));
 sg13g2_buf_1 _2251_ (.A(net116),
    .X(_1527_));
 sg13g2_and3_1 _2252_ (.X(_1528_),
    .A(net115),
    .B(_1517_),
    .C(_1524_));
 sg13g2_a221oi_1 _2253_ (.B2(net66),
    .C1(_1528_),
    .B1(_1526_),
    .A1(_1514_),
    .Y(_1529_),
    .A2(_1521_));
 sg13g2_buf_1 _2254_ (.A(\vga.ball_pos_v[4] ),
    .X(_1530_));
 sg13g2_buf_8 _2255_ (.A(\vga.paddle_r_pos_v[4] ),
    .X(_1531_));
 sg13g2_buf_1 _2256_ (.A(_1531_),
    .X(_1532_));
 sg13g2_nor2b_1 _2257_ (.A(net143),
    .B_N(net114),
    .Y(_1533_));
 sg13g2_nor2b_1 _2258_ (.A(_1531_),
    .B_N(net143),
    .Y(_1534_));
 sg13g2_buf_2 _2259_ (.A(_0069_),
    .X(_1535_));
 sg13g2_buf_2 _2260_ (.A(\vga.ball_pos_v[5] ),
    .X(_1536_));
 sg13g2_xnor2_1 _2261_ (.Y(_1537_),
    .A(_1535_),
    .B(_1536_));
 sg13g2_mux2_1 _2262_ (.A0(_1533_),
    .A1(_1534_),
    .S(_1537_),
    .X(_1538_));
 sg13g2_and2_1 _2263_ (.A(net144),
    .B(net116),
    .X(_1539_));
 sg13g2_buf_1 _2264_ (.A(_1539_),
    .X(_1540_));
 sg13g2_nor2_2 _2265_ (.A(net144),
    .B(_1516_),
    .Y(_1541_));
 sg13g2_a21oi_1 _2266_ (.A1(_1525_),
    .A2(_1540_),
    .Y(_1542_),
    .B1(_1541_));
 sg13g2_xnor2_1 _2267_ (.Y(_1543_),
    .A(_1531_),
    .B(_1530_));
 sg13g2_and4_1 _2268_ (.A(_1524_),
    .B(_1541_),
    .C(_1537_),
    .D(_1543_),
    .X(_1544_));
 sg13g2_a21oi_1 _2269_ (.A1(_1538_),
    .A2(_1542_),
    .Y(_1545_),
    .B1(_1544_));
 sg13g2_nor3_1 _2270_ (.A(net147),
    .B(_1529_),
    .C(_1545_),
    .Y(_1546_));
 sg13g2_and2_1 _2271_ (.A(_1541_),
    .B(_1534_),
    .X(_1547_));
 sg13g2_buf_2 _2272_ (.A(\vga.paddle_r_pos_v[5] ),
    .X(_1548_));
 sg13g2_buf_1 _2273_ (.A(_1548_),
    .X(_1549_));
 sg13g2_o21ai_1 _2274_ (.B1(_1531_),
    .Y(_1550_),
    .A1(\vga.paddle_r_pos_v[3] ),
    .A2(_1515_));
 sg13g2_buf_1 _2275_ (.A(_1550_),
    .X(_1551_));
 sg13g2_xnor2_1 _2276_ (.Y(_1552_),
    .A(net113),
    .B(net65));
 sg13g2_buf_1 _2277_ (.A(_0074_),
    .X(_1553_));
 sg13g2_inv_2 _2278_ (.Y(_1554_),
    .A(_1553_));
 sg13g2_nand2_1 _2279_ (.Y(_1555_),
    .A(net114),
    .B(net143));
 sg13g2_nor3_1 _2280_ (.A(_1541_),
    .B(_1537_),
    .C(_1555_),
    .Y(_1556_));
 sg13g2_a221oi_1 _2281_ (.B2(_1554_),
    .C1(_1556_),
    .B1(_1552_),
    .A1(_1537_),
    .Y(_1557_),
    .A2(_1547_));
 sg13g2_buf_2 _2282_ (.A(\vga.paddle_r_pos_v[6] ),
    .X(_1558_));
 sg13g2_inv_1 _2283_ (.Y(_1559_),
    .A(_1558_));
 sg13g2_or2_1 _2284_ (.X(_1560_),
    .B(_1515_),
    .A(net144));
 sg13g2_buf_1 _2285_ (.A(_1560_),
    .X(_1561_));
 sg13g2_nor2b_1 _2286_ (.A(net113),
    .B_N(_1532_),
    .Y(_1562_));
 sg13g2_inv_1 _2287_ (.Y(_1563_),
    .A(_1535_));
 sg13g2_a21oi_1 _2288_ (.A1(_1561_),
    .A2(_1562_),
    .Y(_1564_),
    .B1(_1563_));
 sg13g2_nor2_1 _2289_ (.A(_1559_),
    .B(_1564_),
    .Y(_1565_));
 sg13g2_o21ai_1 _2290_ (.B1(_1565_),
    .Y(_1566_),
    .A1(net147),
    .A2(_1557_));
 sg13g2_buf_2 _2291_ (.A(_0071_),
    .X(_1567_));
 sg13g2_nor2_1 _2292_ (.A(_1548_),
    .B(_1558_),
    .Y(_1568_));
 sg13g2_inv_1 _2293_ (.Y(_1569_),
    .A(_0070_));
 sg13g2_a21o_1 _2294_ (.A2(_1568_),
    .A1(net65),
    .B1(_1569_),
    .X(_1570_));
 sg13g2_nand3_1 _2295_ (.B(net65),
    .C(_1568_),
    .A(_1569_),
    .Y(_1571_));
 sg13g2_buf_1 _2296_ (.A(\vga.ball_pos_v[7] ),
    .X(_1572_));
 sg13g2_inv_1 _2297_ (.Y(_1573_),
    .A(_1572_));
 sg13g2_a21oi_1 _2298_ (.A1(_1570_),
    .A2(_1571_),
    .Y(_1574_),
    .B1(_1573_));
 sg13g2_and3_1 _2299_ (.X(_1575_),
    .A(_1573_),
    .B(_1570_),
    .C(_1571_));
 sg13g2_buf_1 _2300_ (.A(_1558_),
    .X(_1576_));
 sg13g2_o21ai_1 _2301_ (.B1(_1535_),
    .Y(_1577_),
    .A1(_1549_),
    .A2(net65));
 sg13g2_buf_2 _2302_ (.A(_1577_),
    .X(_1578_));
 sg13g2_nor2_1 _2303_ (.A(net112),
    .B(_1578_),
    .Y(_1579_));
 sg13g2_nor4_1 _2304_ (.A(_1567_),
    .B(_1574_),
    .C(_1575_),
    .D(_1579_),
    .Y(_1580_));
 sg13g2_o21ai_1 _2305_ (.B1(_1580_),
    .Y(_1581_),
    .A1(_1546_),
    .A2(_1566_));
 sg13g2_buf_1 _2306_ (.A(\vga.ball_pos_v[8] ),
    .X(_1582_));
 sg13g2_buf_1 _2307_ (.A(\vga.paddle_r_pos_v[7] ),
    .X(_1583_));
 sg13g2_inv_1 _2308_ (.Y(_1584_),
    .A(net141));
 sg13g2_nand2_1 _2309_ (.Y(_1585_),
    .A(_1584_),
    .B(_1559_));
 sg13g2_o21ai_1 _2310_ (.B1(_0068_),
    .Y(_1586_),
    .A1(_1585_),
    .A2(_1578_));
 sg13g2_or3_1 _2311_ (.A(_0068_),
    .B(_1585_),
    .C(_1578_),
    .X(_1587_));
 sg13g2_nand2_1 _2312_ (.Y(_1588_),
    .A(_1586_),
    .B(_1587_));
 sg13g2_nand2_1 _2313_ (.Y(_1589_),
    .A(_1551_),
    .B(_1568_));
 sg13g2_xnor2_1 _2314_ (.Y(_1590_),
    .A(_1584_),
    .B(_1589_));
 sg13g2_inv_1 _2315_ (.Y(_1591_),
    .A(_0073_));
 sg13g2_a22oi_1 _2316_ (.Y(_1592_),
    .B1(_1590_),
    .B2(_1591_),
    .A2(_1588_),
    .A1(net142));
 sg13g2_o21ai_1 _2317_ (.B1(net147),
    .Y(_1593_),
    .A1(_1559_),
    .A2(_1567_));
 sg13g2_nand2_1 _2318_ (.Y(_1594_),
    .A(_1567_),
    .B(_1564_));
 sg13g2_mux2_1 _2319_ (.A0(net147),
    .A1(_1593_),
    .S(_1594_),
    .X(_1595_));
 sg13g2_nor2_1 _2320_ (.A(_1574_),
    .B(_1575_),
    .Y(_1596_));
 sg13g2_o21ai_1 _2321_ (.B1(_1557_),
    .Y(_1597_),
    .A1(_1529_),
    .A2(_1545_));
 sg13g2_nand3b_1 _2322_ (.B(_1596_),
    .C(_1597_),
    .Y(_1598_),
    .A_N(_1595_));
 sg13g2_and3_1 _2323_ (.X(_1599_),
    .A(_1581_),
    .B(_1592_),
    .C(_1598_));
 sg13g2_buf_1 _2324_ (.A(_1599_),
    .X(_1600_));
 sg13g2_buf_2 _2325_ (.A(_0067_),
    .X(_1601_));
 sg13g2_buf_8 _2326_ (.A(_1601_),
    .X(_1602_));
 sg13g2_inv_2 _2327_ (.Y(_1603_),
    .A(_1602_));
 sg13g2_buf_1 _2328_ (.A(\vga.paddle_r_pos_v[8] ),
    .X(_1604_));
 sg13g2_nor4_2 _2329_ (.A(net141),
    .B(_1604_),
    .C(_1549_),
    .Y(_1605_),
    .D(net112));
 sg13g2_nand2_2 _2330_ (.Y(_1606_),
    .A(net65),
    .B(_1605_));
 sg13g2_nor2b_1 _2331_ (.A(net142),
    .B_N(_0068_),
    .Y(_1607_));
 sg13g2_o21ai_1 _2332_ (.B1(_1607_),
    .Y(_1608_),
    .A1(_1585_),
    .A2(_1578_));
 sg13g2_or4_1 _2333_ (.A(_0068_),
    .B(_1582_),
    .C(_1585_),
    .D(_1578_),
    .X(_1609_));
 sg13g2_nand4_1 _2334_ (.B(_1606_),
    .C(_1608_),
    .A(_1603_),
    .Y(_1610_),
    .D(_1609_));
 sg13g2_nand2_1 _2335_ (.Y(_1611_),
    .A(net111),
    .B(_1606_));
 sg13g2_a21o_1 _2336_ (.A2(_1587_),
    .A1(_1586_),
    .B1(_1611_),
    .X(_1612_));
 sg13g2_nand2_1 _2337_ (.Y(_1613_),
    .A(_1610_),
    .B(_1612_));
 sg13g2_xor2_1 _2338_ (.B(_1567_),
    .A(_1558_),
    .X(_1614_));
 sg13g2_a21o_1 _2339_ (.A2(_1515_),
    .A1(net144),
    .B1(_1531_),
    .X(_1615_));
 sg13g2_buf_1 _2340_ (.A(_1615_),
    .X(_1616_));
 sg13g2_nand3_1 _2341_ (.B(_1614_),
    .C(_1616_),
    .A(net113),
    .Y(_1617_));
 sg13g2_a21o_1 _2342_ (.A2(_1616_),
    .A1(net113),
    .B1(_1614_),
    .X(_1618_));
 sg13g2_buf_1 _2343_ (.A(_0061_),
    .X(_1619_));
 sg13g2_nand3b_1 _2344_ (.B(net144),
    .C(_1515_),
    .Y(_1620_),
    .A_N(_1531_));
 sg13g2_buf_2 _2345_ (.A(_1620_),
    .X(_1621_));
 sg13g2_or2_1 _2346_ (.X(_1622_),
    .B(_1536_),
    .A(net113));
 sg13g2_a21o_1 _2347_ (.A2(_1621_),
    .A1(net140),
    .B1(_1622_),
    .X(_1623_));
 sg13g2_inv_2 _2348_ (.Y(_1624_),
    .A(_1536_));
 sg13g2_nand4_1 _2349_ (.B(net140),
    .C(_1624_),
    .A(net113),
    .Y(_1625_),
    .D(_1621_));
 sg13g2_nand4_1 _2350_ (.B(_1618_),
    .C(_1623_),
    .A(_1617_),
    .Y(_1626_),
    .D(_1625_));
 sg13g2_and3_1 _2351_ (.X(_1627_),
    .A(net141),
    .B(_1548_),
    .C(_1558_));
 sg13g2_buf_1 _2352_ (.A(_1627_),
    .X(_1628_));
 sg13g2_a21oi_1 _2353_ (.A1(_1522_),
    .A2(net116),
    .Y(_1629_),
    .B1(net114));
 sg13g2_or2_1 _2354_ (.X(_1630_),
    .B(_1601_),
    .A(_1604_));
 sg13g2_nand4_1 _2355_ (.B(net114),
    .C(_1619_),
    .A(_1604_),
    .Y(_1631_),
    .D(_1601_));
 sg13g2_o21ai_1 _2356_ (.B1(_1631_),
    .Y(_1632_),
    .A1(_1629_),
    .A2(_1630_));
 sg13g2_nor2b_1 _2357_ (.A(net140),
    .B_N(_1604_),
    .Y(_1633_));
 sg13g2_o21ai_1 _2358_ (.B1(_1628_),
    .Y(_1634_),
    .A1(_1616_),
    .A2(_1633_));
 sg13g2_buf_1 _2359_ (.A(_1604_),
    .X(_1635_));
 sg13g2_xor2_1 _2360_ (.B(_1602_),
    .A(net110),
    .X(_1636_));
 sg13g2_a22oi_1 _2361_ (.Y(_1637_),
    .B1(_1634_),
    .B2(_1636_),
    .A2(_1632_),
    .A1(_1628_));
 sg13g2_nand2_1 _2362_ (.Y(_1638_),
    .A(_1548_),
    .B(_1558_));
 sg13g2_and2_1 _2363_ (.A(\vga.paddle_r_pos_v[7] ),
    .B(_0061_),
    .X(_1639_));
 sg13g2_a22oi_1 _2364_ (.Y(_1640_),
    .B1(_1639_),
    .B2(_1621_),
    .A2(_1638_),
    .A1(net141));
 sg13g2_nand3b_1 _2365_ (.B(_1548_),
    .C(_1558_),
    .Y(_1641_),
    .A_N(net141));
 sg13g2_a21o_1 _2366_ (.A2(_1621_),
    .A1(net140),
    .B1(_1641_),
    .X(_1642_));
 sg13g2_a21oi_1 _2367_ (.A1(_1640_),
    .A2(_1642_),
    .Y(_1643_),
    .B1(_1572_));
 sg13g2_and3_1 _2368_ (.X(_1644_),
    .A(_1572_),
    .B(_1640_),
    .C(_1642_));
 sg13g2_or4_1 _2369_ (.A(_1626_),
    .B(_1637_),
    .C(_1643_),
    .D(_1644_),
    .X(_1645_));
 sg13g2_buf_1 _2370_ (.A(_1536_),
    .X(_1646_));
 sg13g2_buf_1 _2371_ (.A(net113),
    .X(_1647_));
 sg13g2_o21ai_1 _2372_ (.B1(net140),
    .Y(_1648_),
    .A1(net114),
    .A2(net143));
 sg13g2_xnor2_1 _2373_ (.Y(_1649_),
    .A(net64),
    .B(_1648_));
 sg13g2_nand2_2 _2374_ (.Y(_1650_),
    .A(net144),
    .B(_1516_));
 sg13g2_xnor2_1 _2375_ (.Y(_1651_),
    .A(_1650_),
    .B(_1543_));
 sg13g2_a21oi_1 _2376_ (.A1(net109),
    .A2(_1649_),
    .Y(_1652_),
    .B1(_1651_));
 sg13g2_buf_1 _2377_ (.A(_1512_),
    .X(_1653_));
 sg13g2_xnor2_1 _2378_ (.Y(_1654_),
    .A(net108),
    .B(_1511_));
 sg13g2_buf_1 _2379_ (.A(_1508_),
    .X(_1655_));
 sg13g2_buf_1 _2380_ (.A(_1510_),
    .X(_1656_));
 sg13g2_xnor2_1 _2381_ (.Y(_1657_),
    .A(_1655_),
    .B(net106));
 sg13g2_buf_1 _2382_ (.A(net145),
    .X(_1658_));
 sg13g2_buf_1 _2383_ (.A(_0075_),
    .X(_1659_));
 sg13g2_xnor2_1 _2384_ (.Y(_1660_),
    .A(net144),
    .B(_1659_));
 sg13g2_nand2_1 _2385_ (.Y(_1661_),
    .A(net116),
    .B(_1660_));
 sg13g2_or3_1 _2386_ (.A(net116),
    .B(_1519_),
    .C(_1660_),
    .X(_1662_));
 sg13g2_o21ai_1 _2387_ (.B1(_1662_),
    .Y(_1663_),
    .A1(_1658_),
    .A2(_1661_));
 sg13g2_nand4_1 _2388_ (.B(_1654_),
    .C(_1657_),
    .A(_1652_),
    .Y(_1664_),
    .D(_1663_));
 sg13g2_nor2_1 _2389_ (.A(_1645_),
    .B(_1664_),
    .Y(_1665_));
 sg13g2_buf_1 _2390_ (.A(net143),
    .X(_1666_));
 sg13g2_xnor2_1 _2391_ (.Y(_1667_),
    .A(net114),
    .B(_1650_));
 sg13g2_nand2_1 _2392_ (.Y(_1668_),
    .A(net140),
    .B(_1621_));
 sg13g2_xnor2_1 _2393_ (.Y(_1669_),
    .A(net64),
    .B(_1668_));
 sg13g2_a22oi_1 _2394_ (.Y(_1670_),
    .B1(_1669_),
    .B2(net109),
    .A2(_1667_),
    .A1(net104));
 sg13g2_nand3_1 _2395_ (.B(net145),
    .C(_1660_),
    .A(net66),
    .Y(_1671_));
 sg13g2_nor2_1 _2396_ (.A(_1656_),
    .B(_1513_),
    .Y(_1672_));
 sg13g2_a21oi_1 _2397_ (.A1(_1656_),
    .A2(_1513_),
    .Y(_1673_),
    .B1(_1509_));
 sg13g2_a221oi_1 _2398_ (.B2(_1672_),
    .C1(_1673_),
    .B1(_1671_),
    .A1(_1661_),
    .Y(_1674_),
    .A2(_1662_));
 sg13g2_a21oi_1 _2399_ (.A1(_1518_),
    .A2(_1659_),
    .Y(_1675_),
    .B1(_1524_));
 sg13g2_buf_1 _2400_ (.A(_1524_),
    .X(_1676_));
 sg13g2_nor2b_1 _2401_ (.A(net139),
    .B_N(net145),
    .Y(_1677_));
 sg13g2_nor2b_1 _2402_ (.A(net115),
    .B_N(net116),
    .Y(_1678_));
 sg13g2_a22oi_1 _2403_ (.Y(_1679_),
    .B1(_1677_),
    .B2(_1678_),
    .A2(_1541_),
    .A1(_1676_));
 sg13g2_o21ai_1 _2404_ (.B1(_1679_),
    .Y(_1680_),
    .A1(_1650_),
    .A2(_1675_));
 sg13g2_o21ai_1 _2405_ (.B1(_1652_),
    .Y(_1681_),
    .A1(_1674_),
    .A2(_1680_));
 sg13g2_a21o_1 _2406_ (.A2(_1681_),
    .A1(_1670_),
    .B1(_1645_),
    .X(_1682_));
 sg13g2_buf_1 _2407_ (.A(_1572_),
    .X(_1683_));
 sg13g2_and2_1 _2408_ (.A(_1640_),
    .B(_1642_),
    .X(_1684_));
 sg13g2_buf_1 _2409_ (.A(_1684_),
    .X(_1685_));
 sg13g2_nand3_1 _2410_ (.B(_1559_),
    .C(_1616_),
    .A(net64),
    .Y(_1686_));
 sg13g2_inv_2 _2411_ (.Y(_1687_),
    .A(net113));
 sg13g2_o21ai_1 _2412_ (.B1(net112),
    .Y(_1688_),
    .A1(_1687_),
    .A2(_1629_));
 sg13g2_and3_1 _2413_ (.X(_1689_),
    .A(\vga.ball_pos_v[6] ),
    .B(_1686_),
    .C(_1688_));
 sg13g2_a21o_1 _2414_ (.A2(_1685_),
    .A1(_1683_),
    .B1(_1689_),
    .X(_1690_));
 sg13g2_nor2_1 _2415_ (.A(_1637_),
    .B(_1643_),
    .Y(_1691_));
 sg13g2_and2_1 _2416_ (.A(_1616_),
    .B(_1628_),
    .X(_1692_));
 sg13g2_nand4_1 _2417_ (.B(_1532_),
    .C(_1619_),
    .A(net110),
    .Y(_1693_),
    .D(_1628_));
 sg13g2_o21ai_1 _2418_ (.B1(_1693_),
    .Y(_1694_),
    .A1(net110),
    .A2(_1692_));
 sg13g2_and2_1 _2419_ (.A(_1582_),
    .B(_1694_),
    .X(_1695_));
 sg13g2_a221oi_1 _2420_ (.B2(_1691_),
    .C1(_1695_),
    .B1(_1690_),
    .A1(_1610_),
    .Y(_1696_),
    .A2(_1612_));
 sg13g2_a22oi_1 _2421_ (.Y(_1697_),
    .B1(_1682_),
    .B2(_1696_),
    .A2(_1665_),
    .A1(_1613_));
 sg13g2_inv_1 _2422_ (.Y(_1698_),
    .A(\vga.interval_counter[4] ));
 sg13g2_buf_1 _2423_ (.A(\vga.interval_counter[13] ),
    .X(_1699_));
 sg13g2_inv_1 _2424_ (.Y(_1700_),
    .A(_1699_));
 sg13g2_buf_2 _2425_ (.A(\vga.interval_counter[1] ),
    .X(_1701_));
 sg13g2_buf_1 _2426_ (.A(\vga.interval_counter[5] ),
    .X(_1702_));
 sg13g2_nor2_1 _2427_ (.A(_1701_),
    .B(_1702_),
    .Y(_1703_));
 sg13g2_buf_2 _2428_ (.A(\vga.interval_counter[0] ),
    .X(_1704_));
 sg13g2_buf_1 _2429_ (.A(\vga.interval_counter[12] ),
    .X(_1705_));
 sg13g2_buf_1 _2430_ (.A(\vga.interval_counter[15] ),
    .X(_1706_));
 sg13g2_nor3_1 _2431_ (.A(_1704_),
    .B(_1705_),
    .C(_1706_),
    .Y(_1707_));
 sg13g2_nand4_1 _2432_ (.B(_1700_),
    .C(_1703_),
    .A(_1698_),
    .Y(_1708_),
    .D(_1707_));
 sg13g2_buf_2 _2433_ (.A(\vga.interval_counter[3] ),
    .X(_1709_));
 sg13g2_buf_2 _2434_ (.A(\vga.interval_counter[7] ),
    .X(_1710_));
 sg13g2_buf_1 _2435_ (.A(\vga.interval_counter[17] ),
    .X(_1711_));
 sg13g2_nor4_1 _2436_ (.A(_1709_),
    .B(_1710_),
    .C(\vga.interval_counter[10] ),
    .D(_1711_),
    .Y(_1712_));
 sg13g2_buf_1 _2437_ (.A(\vga.interval_counter[8] ),
    .X(_1713_));
 sg13g2_buf_2 _2438_ (.A(\vga.interval_counter[9] ),
    .X(_1714_));
 sg13g2_nor3_1 _2439_ (.A(_1713_),
    .B(_1714_),
    .C(\vga.interval_counter[11] ),
    .Y(_1715_));
 sg13g2_nand2_1 _2440_ (.Y(_1716_),
    .A(_1712_),
    .B(_1715_));
 sg13g2_buf_1 _2441_ (.A(\vga.interval_counter[20] ),
    .X(_1717_));
 sg13g2_nor4_1 _2442_ (.A(_1717_),
    .B(\vga.interval_counter[23] ),
    .C(\vga.interval_counter[22] ),
    .D(\vga.interval_counter[24] ),
    .Y(_1718_));
 sg13g2_nand2b_1 _2443_ (.Y(_1719_),
    .B(_1718_),
    .A_N(\vga.interval_counter[21] ));
 sg13g2_buf_2 _2444_ (.A(\vga.interval_counter[2] ),
    .X(_1720_));
 sg13g2_buf_1 _2445_ (.A(\vga.interval_counter[6] ),
    .X(_1721_));
 sg13g2_buf_2 _2446_ (.A(\vga.interval_counter[14] ),
    .X(_1722_));
 sg13g2_nor3_1 _2447_ (.A(_1720_),
    .B(_1721_),
    .C(_1722_),
    .Y(_1723_));
 sg13g2_buf_1 _2448_ (.A(\vga.interval_counter[16] ),
    .X(_1724_));
 sg13g2_buf_1 _2449_ (.A(\vga.interval_counter[19] ),
    .X(_1725_));
 sg13g2_buf_1 _2450_ (.A(\vga.interval_counter[18] ),
    .X(_1726_));
 sg13g2_nor3_1 _2451_ (.A(_1724_),
    .B(_1725_),
    .C(_1726_),
    .Y(_1727_));
 sg13g2_nand2_1 _2452_ (.Y(_1728_),
    .A(_1723_),
    .B(_1727_));
 sg13g2_nor4_2 _2453_ (.A(_1708_),
    .B(_1716_),
    .C(_1719_),
    .Y(_1729_),
    .D(_1728_));
 sg13g2_buf_1 _2454_ (.A(\vga.ball_motion_l ),
    .X(_1730_));
 sg13g2_buf_1 _2455_ (.A(\vga.ball_pos_h[0] ),
    .X(_1731_));
 sg13g2_nand2_1 _2456_ (.Y(_1732_),
    .A(net138),
    .B(\vga.ball_pos_h[1] ));
 sg13g2_buf_1 _2457_ (.A(\vga.ball_pos_h[3] ),
    .X(_1733_));
 sg13g2_buf_1 _2458_ (.A(\vga.ball_pos_h[2] ),
    .X(_1734_));
 sg13g2_nand2_2 _2459_ (.Y(_1735_),
    .A(_1733_),
    .B(_1734_));
 sg13g2_or2_1 _2460_ (.X(_1736_),
    .B(_1735_),
    .A(_1732_));
 sg13g2_buf_1 _2461_ (.A(_1736_),
    .X(_1737_));
 sg13g2_buf_1 _2462_ (.A(\vga.ball_pos_h[6] ),
    .X(_1738_));
 sg13g2_buf_2 _2463_ (.A(\vga.ball_pos_h[9] ),
    .X(_1739_));
 sg13g2_buf_2 _2464_ (.A(\vga.ball_pos_h[4] ),
    .X(_1740_));
 sg13g2_buf_1 _2465_ (.A(\vga.ball_pos_h[5] ),
    .X(_1741_));
 sg13g2_inv_1 _2466_ (.Y(_1742_),
    .A(net136));
 sg13g2_nor2_1 _2467_ (.A(_1740_),
    .B(_1742_),
    .Y(_1743_));
 sg13g2_buf_1 _2468_ (.A(\vga.ball_pos_h[7] ),
    .X(_1744_));
 sg13g2_buf_1 _2469_ (.A(\vga.ball_pos_h[8] ),
    .X(_1745_));
 sg13g2_nor2_1 _2470_ (.A(_1744_),
    .B(_1745_),
    .Y(_1746_));
 sg13g2_nand4_1 _2471_ (.B(_1739_),
    .C(_1743_),
    .A(_1738_),
    .Y(_1747_),
    .D(_1746_));
 sg13g2_nor3_1 _2472_ (.A(_1730_),
    .B(_1737_),
    .C(_1747_),
    .Y(_1748_));
 sg13g2_buf_2 _2473_ (.A(_1748_),
    .X(_1749_));
 sg13g2_nand2_1 _2474_ (.Y(_1750_),
    .A(_1729_),
    .B(_1749_));
 sg13g2_inv_1 _2475_ (.Y(_1751_),
    .A(_1750_));
 sg13g2_o21ai_1 _2476_ (.B1(_1751_),
    .Y(_1752_),
    .A1(_1600_),
    .A2(_1697_));
 sg13g2_buf_2 _2477_ (.A(_1752_),
    .X(_1753_));
 sg13g2_buf_1 _2478_ (.A(\vga.score_l[1] ),
    .X(_1754_));
 sg13g2_buf_2 _2479_ (.A(\vga.score_l[0] ),
    .X(_1755_));
 sg13g2_buf_1 _2480_ (.A(\vga.score_l[2] ),
    .X(_1756_));
 sg13g2_nand3_1 _2481_ (.B(_1755_),
    .C(_1756_),
    .A(_1754_),
    .Y(_1757_));
 sg13g2_buf_1 _2482_ (.A(_1757_),
    .X(_1758_));
 sg13g2_nor2_1 _2483_ (.A(_1753_),
    .B(_1758_),
    .Y(_1759_));
 sg13g2_nand2_1 _2484_ (.Y(_1760_),
    .A(_1754_),
    .B(_1755_));
 sg13g2_or2_1 _2485_ (.X(_1761_),
    .B(_1760_),
    .A(_1756_));
 sg13g2_buf_1 _2486_ (.A(_1761_),
    .X(_1762_));
 sg13g2_inv_1 _2487_ (.Y(_1763_),
    .A(\vga.score_l[4] ));
 sg13g2_nand2_1 _2488_ (.Y(_1764_),
    .A(_1763_),
    .B(_1758_));
 sg13g2_a22oi_1 _2489_ (.Y(_1765_),
    .B1(_1764_),
    .B2(net148),
    .A2(_1762_),
    .A1(\vga.score_l[4] ));
 sg13g2_or2_1 _2490_ (.X(_1766_),
    .B(_1765_),
    .A(_1753_));
 sg13g2_buf_2 _2491_ (.A(ui_in[4]),
    .X(_1767_));
 sg13g2_inv_1 _2492_ (.Y(_1768_),
    .A(_1767_));
 sg13g2_nand2_1 _2493_ (.Y(_1769_),
    .A(\vga.score_l[4] ),
    .B(net135));
 sg13g2_buf_2 _2494_ (.A(rst_n),
    .X(_1770_));
 sg13g2_inv_1 _2495_ (.Y(_1771_),
    .A(_1770_));
 sg13g2_buf_1 _2496_ (.A(_1771_),
    .X(_1772_));
 sg13g2_a221oi_1 _2497_ (.B2(_1769_),
    .C1(net101),
    .B1(_1766_),
    .A1(_1506_),
    .Y(_1773_),
    .A2(_1759_));
 sg13g2_buf_1 _2498_ (.A(_1773_),
    .X(_1774_));
 sg13g2_buf_1 _2499_ (.A(_1774_),
    .X(_0200_));
 sg13g2_nor3_1 _2500_ (.A(net148),
    .B(_1763_),
    .C(_1762_),
    .Y(_1775_));
 sg13g2_nand2_1 _2501_ (.Y(_1776_),
    .A(_1756_),
    .B(_1760_));
 sg13g2_o21ai_1 _2502_ (.B1(_1776_),
    .Y(_1777_),
    .A1(_1762_),
    .A2(_1775_));
 sg13g2_nand2_1 _2503_ (.Y(_1778_),
    .A(_1770_),
    .B(_1777_));
 sg13g2_nor2_1 _2504_ (.A(net101),
    .B(_1767_),
    .Y(_1779_));
 sg13g2_nand2_1 _2505_ (.Y(_1780_),
    .A(_1756_),
    .B(_1779_));
 sg13g2_mux2_1 _2506_ (.A0(_1778_),
    .A1(_1780_),
    .S(_1753_),
    .X(_1781_));
 sg13g2_buf_2 _2507_ (.A(_1781_),
    .X(_1782_));
 sg13g2_inv_4 _2508_ (.A(_1782_),
    .Y(_0198_));
 sg13g2_nand3_1 _2509_ (.B(_1505_),
    .C(_1758_),
    .A(_1770_),
    .Y(_1783_));
 sg13g2_or3_1 _2510_ (.A(_1771_),
    .B(net148),
    .C(_1758_),
    .X(_1784_));
 sg13g2_a21oi_1 _2511_ (.A1(_1783_),
    .A2(_1784_),
    .Y(_1785_),
    .B1(_1753_));
 sg13g2_nand4_1 _2512_ (.B(_1505_),
    .C(net135),
    .A(_1770_),
    .Y(_1786_),
    .D(_1753_));
 sg13g2_nand2b_1 _2513_ (.Y(_1787_),
    .B(_1786_),
    .A_N(_1785_));
 sg13g2_buf_1 _2514_ (.A(_1787_),
    .X(_0199_));
 sg13g2_nor2_1 _2515_ (.A(net34),
    .B(net33),
    .Y(_1788_));
 sg13g2_inv_1 _2516_ (.Y(_1789_),
    .A(_1788_));
 sg13g2_mux2_1 _2517_ (.A0(_1758_),
    .A1(net135),
    .S(_1753_),
    .X(_1790_));
 sg13g2_nor3_1 _2518_ (.A(net148),
    .B(_1753_),
    .C(_1758_),
    .Y(_1791_));
 sg13g2_a21o_1 _2519_ (.A2(_1790_),
    .A1(net148),
    .B1(_1791_),
    .X(_1792_));
 sg13g2_nor2_1 _2520_ (.A(_1750_),
    .B(_1775_),
    .Y(_1793_));
 sg13g2_o21ai_1 _2521_ (.B1(_1793_),
    .Y(_1794_),
    .A1(_1600_),
    .A2(_1697_));
 sg13g2_nand3_1 _2522_ (.B(net135),
    .C(_1794_),
    .A(_1754_),
    .Y(_1795_));
 sg13g2_nand2b_1 _2523_ (.Y(_1796_),
    .B(_1754_),
    .A_N(_1755_));
 sg13g2_nand2b_1 _2524_ (.Y(_1797_),
    .B(_1755_),
    .A_N(_1754_));
 sg13g2_a21o_1 _2525_ (.A2(_1797_),
    .A1(_1796_),
    .B1(_1753_),
    .X(_1798_));
 sg13g2_nand2_1 _2526_ (.Y(_1799_),
    .A(_1795_),
    .B(_1798_));
 sg13g2_buf_2 _2527_ (.A(_1799_),
    .X(_1800_));
 sg13g2_buf_1 _2528_ (.A(_1770_),
    .X(_1801_));
 sg13g2_o21ai_1 _2529_ (.B1(net134),
    .Y(_1802_),
    .A1(_1792_),
    .A2(_1800_));
 sg13g2_a21o_1 _2530_ (.A2(_1800_),
    .A1(_1792_),
    .B1(_1802_),
    .X(_1803_));
 sg13g2_nor2_1 _2531_ (.A(net101),
    .B(_1755_),
    .Y(_1804_));
 sg13g2_and3_1 _2532_ (.X(_1805_),
    .A(_1770_),
    .B(_1755_),
    .C(net135));
 sg13g2_mux2_1 _2533_ (.A0(_1804_),
    .A1(_1805_),
    .S(_1794_),
    .X(_1806_));
 sg13g2_buf_1 _2534_ (.A(_1806_),
    .X(_1807_));
 sg13g2_buf_1 _2535_ (.A(_1807_),
    .X(_0196_));
 sg13g2_a221oi_1 _2536_ (.B2(net34),
    .C1(net39),
    .B1(_1803_),
    .A1(net31),
    .Y(_0008_),
    .A2(_1789_));
 sg13g2_buf_1 _2537_ (.A(\vga.score_r[3] ),
    .X(_1808_));
 sg13g2_buf_1 _2538_ (.A(\vga.paddle_l_pos_v[5] ),
    .X(_1809_));
 sg13g2_buf_8 _2539_ (.A(_1809_),
    .X(_1810_));
 sg13g2_or2_1 _2540_ (.X(_1811_),
    .B(_1553_),
    .A(net100));
 sg13g2_buf_1 _2541_ (.A(net100),
    .X(_1812_));
 sg13g2_nand2b_1 _2542_ (.Y(_1813_),
    .B(net63),
    .A_N(_1553_));
 sg13g2_buf_8 _2543_ (.A(\vga.paddle_l_pos_v[2] ),
    .X(_1814_));
 sg13g2_buf_8 _2544_ (.A(\vga.paddle_l_pos_v[4] ),
    .X(_1815_));
 sg13g2_o21ai_1 _2545_ (.B1(_1815_),
    .Y(_1816_),
    .A1(\vga.paddle_l_pos_v[3] ),
    .A2(_1814_));
 sg13g2_buf_8 _2546_ (.A(_1816_),
    .X(_1817_));
 sg13g2_mux2_1 _2547_ (.A0(_1811_),
    .A1(_1813_),
    .S(net62),
    .X(_1818_));
 sg13g2_buf_2 _2548_ (.A(_0077_),
    .X(_1819_));
 sg13g2_xnor2_1 _2549_ (.Y(_1820_),
    .A(_1536_),
    .B(_1819_));
 sg13g2_buf_1 _2550_ (.A(_1815_),
    .X(_1821_));
 sg13g2_buf_8 _2551_ (.A(\vga.paddle_l_pos_v[3] ),
    .X(_1822_));
 sg13g2_buf_1 _2552_ (.A(_1814_),
    .X(_1823_));
 sg13g2_nor2_1 _2553_ (.A(net132),
    .B(_1823_),
    .Y(_1824_));
 sg13g2_buf_2 _2554_ (.A(_1824_),
    .X(_1825_));
 sg13g2_nor2_1 _2555_ (.A(net143),
    .B(_1825_),
    .Y(_1826_));
 sg13g2_nand2_1 _2556_ (.Y(_1827_),
    .A(net104),
    .B(_1825_));
 sg13g2_o21ai_1 _2557_ (.B1(_1827_),
    .Y(_1828_),
    .A1(net99),
    .A2(_1826_));
 sg13g2_nor2_1 _2558_ (.A(net62),
    .B(_1820_),
    .Y(_1829_));
 sg13g2_a21oi_1 _2559_ (.A1(_1820_),
    .A2(_1828_),
    .Y(_1830_),
    .B1(_1829_));
 sg13g2_inv_1 _2560_ (.Y(_1831_),
    .A(net98));
 sg13g2_nand2_1 _2561_ (.Y(_1832_),
    .A(_1831_),
    .B(net105));
 sg13g2_buf_1 _2562_ (.A(\vga.paddle_l_pos_v[0] ),
    .X(_1833_));
 sg13g2_nor2b_1 _2563_ (.A(net146),
    .B_N(net131),
    .Y(_1834_));
 sg13g2_nand2b_1 _2564_ (.Y(_1835_),
    .B(\vga.paddle_l_pos_v[0] ),
    .A_N(net146));
 sg13g2_buf_2 _2565_ (.A(_1835_),
    .X(_1836_));
 sg13g2_inv_1 _2566_ (.Y(_1837_),
    .A(\vga.paddle_l_pos_v[1] ));
 sg13g2_a21oi_1 _2567_ (.A1(net106),
    .A2(_1836_),
    .Y(_1838_),
    .B1(_1837_));
 sg13g2_a221oi_1 _2568_ (.B2(_1520_),
    .C1(_1838_),
    .B1(_1834_),
    .A1(_1525_),
    .Y(_1839_),
    .A2(_1832_));
 sg13g2_buf_1 _2569_ (.A(net98),
    .X(_1840_));
 sg13g2_a21oi_1 _2570_ (.A1(net61),
    .A2(_1519_),
    .Y(_1841_),
    .B1(_1525_));
 sg13g2_buf_1 _2571_ (.A(net132),
    .X(_1842_));
 sg13g2_o21ai_1 _2572_ (.B1(net97),
    .Y(_1843_),
    .A1(_1839_),
    .A2(_1841_));
 sg13g2_nand3b_1 _2573_ (.B(_1825_),
    .C(_1820_),
    .Y(_1844_),
    .A_N(net99));
 sg13g2_nand2b_1 _2574_ (.Y(_1845_),
    .B(_1844_),
    .A_N(_1829_));
 sg13g2_o21ai_1 _2575_ (.B1(net105),
    .Y(_1846_),
    .A1(net106),
    .A2(_1836_));
 sg13g2_nor2b_1 _2576_ (.A(net97),
    .B_N(net98),
    .Y(_1847_));
 sg13g2_inv_1 _2577_ (.Y(_1848_),
    .A(_1847_));
 sg13g2_o21ai_1 _2578_ (.B1(_1848_),
    .Y(_1849_),
    .A1(_1838_),
    .A2(_1846_));
 sg13g2_buf_1 _2579_ (.A(\vga.paddle_l_pos_v[1] ),
    .X(_1850_));
 sg13g2_nand2b_1 _2580_ (.Y(_1851_),
    .B(net130),
    .A_N(net145));
 sg13g2_a21oi_1 _2581_ (.A1(net106),
    .A2(_1836_),
    .Y(_1852_),
    .B1(_1851_));
 sg13g2_or2_1 _2582_ (.X(_1853_),
    .B(_1510_),
    .A(net145));
 sg13g2_buf_1 _2583_ (.A(_1853_),
    .X(_1854_));
 sg13g2_o21ai_1 _2584_ (.B1(_1847_),
    .Y(_1855_),
    .A1(_1836_),
    .A2(_1854_));
 sg13g2_o21ai_1 _2585_ (.B1(_1818_),
    .Y(_1856_),
    .A1(_1852_),
    .A2(_1855_));
 sg13g2_a221oi_1 _2586_ (.B2(net103),
    .C1(_1856_),
    .B1(_1849_),
    .A1(net104),
    .Y(_1857_),
    .A2(_1845_));
 sg13g2_inv_2 _2587_ (.Y(_1858_),
    .A(net63));
 sg13g2_nand2b_1 _2588_ (.Y(_1859_),
    .B(_1858_),
    .A_N(net62));
 sg13g2_buf_2 _2589_ (.A(\vga.paddle_l_pos_v[7] ),
    .X(_1860_));
 sg13g2_buf_1 _2590_ (.A(_1860_),
    .X(_1861_));
 sg13g2_buf_2 _2591_ (.A(\vga.paddle_l_pos_v[6] ),
    .X(_1862_));
 sg13g2_buf_8 _2592_ (.A(_1862_),
    .X(_1863_));
 sg13g2_inv_1 _2593_ (.Y(_1864_),
    .A(_1819_));
 sg13g2_buf_2 _2594_ (.A(_0076_),
    .X(_1865_));
 sg13g2_xor2_1 _2595_ (.B(_1865_),
    .A(net111),
    .X(_1866_));
 sg13g2_nor4_1 _2596_ (.A(net96),
    .B(net95),
    .C(_1864_),
    .D(_1866_),
    .Y(_1867_));
 sg13g2_buf_1 _2597_ (.A(\vga.paddle_l_pos_v[8] ),
    .X(_1868_));
 sg13g2_nor3_1 _2598_ (.A(_1868_),
    .B(_1860_),
    .C(net95),
    .Y(_1869_));
 sg13g2_mux2_1 _2599_ (.A0(_1866_),
    .A1(_1869_),
    .S(net62),
    .X(_1870_));
 sg13g2_nor2_1 _2600_ (.A(net96),
    .B(net95),
    .Y(_1871_));
 sg13g2_xnor2_1 _2601_ (.Y(_1872_),
    .A(net111),
    .B(_1865_));
 sg13g2_a21oi_1 _2602_ (.A1(_1819_),
    .A2(_1871_),
    .Y(_1873_),
    .B1(_1872_));
 sg13g2_a221oi_1 _2603_ (.B2(_1858_),
    .C1(_1873_),
    .B1(_1870_),
    .A1(_1859_),
    .Y(_1874_),
    .A2(_1867_));
 sg13g2_nor2_1 _2604_ (.A(_1862_),
    .B(_1809_),
    .Y(_1875_));
 sg13g2_inv_1 _2605_ (.Y(_1876_),
    .A(_0078_));
 sg13g2_a21oi_1 _2606_ (.A1(_1817_),
    .A2(_1875_),
    .Y(_1877_),
    .B1(_1876_));
 sg13g2_and3_1 _2607_ (.X(_1878_),
    .A(_1876_),
    .B(_1816_),
    .C(_1875_));
 sg13g2_buf_1 _2608_ (.A(_1878_),
    .X(_1879_));
 sg13g2_o21ai_1 _2609_ (.B1(net102),
    .Y(_1880_),
    .A1(_1877_),
    .A2(_1879_));
 sg13g2_or3_1 _2610_ (.A(_1683_),
    .B(_1877_),
    .C(_1879_),
    .X(_1881_));
 sg13g2_o21ai_1 _2611_ (.B1(_1819_),
    .Y(_1882_),
    .A1(net100),
    .A2(_1817_));
 sg13g2_buf_2 _2612_ (.A(_1882_),
    .X(_1883_));
 sg13g2_buf_1 _2613_ (.A(_0079_),
    .X(_1884_));
 sg13g2_xnor2_1 _2614_ (.Y(_1885_),
    .A(_1567_),
    .B(_1884_));
 sg13g2_xnor2_1 _2615_ (.Y(_1886_),
    .A(_1883_),
    .B(_1885_));
 sg13g2_nand4_1 _2616_ (.B(_1880_),
    .C(_1881_),
    .A(_1874_),
    .Y(_1887_),
    .D(_1886_));
 sg13g2_a221oi_1 _2617_ (.B2(_1857_),
    .C1(_1887_),
    .B1(_1843_),
    .A1(_1818_),
    .Y(_1888_),
    .A2(_1830_));
 sg13g2_buf_1 _2618_ (.A(net95),
    .X(_1889_));
 sg13g2_nor3_1 _2619_ (.A(_1861_),
    .B(net60),
    .C(_1883_),
    .Y(_1890_));
 sg13g2_xor2_1 _2620_ (.B(_1890_),
    .A(_1865_),
    .X(_1891_));
 sg13g2_and2_1 _2621_ (.A(_1858_),
    .B(_1869_),
    .X(_1892_));
 sg13g2_nand2_1 _2622_ (.Y(_1893_),
    .A(net62),
    .B(_1892_));
 sg13g2_and2_1 _2623_ (.A(net142),
    .B(_1893_),
    .X(_1894_));
 sg13g2_inv_1 _2624_ (.Y(_1895_),
    .A(_1567_));
 sg13g2_xor2_1 _2625_ (.B(_1883_),
    .A(_1889_),
    .X(_1896_));
 sg13g2_and4_1 _2626_ (.A(_1895_),
    .B(_1880_),
    .C(_1881_),
    .D(_1896_),
    .X(_1897_));
 sg13g2_nand2_1 _2627_ (.Y(_1898_),
    .A(net62),
    .B(_1875_));
 sg13g2_xor2_1 _2628_ (.B(_1898_),
    .A(net96),
    .X(_1899_));
 sg13g2_and3_1 _2629_ (.X(_1900_),
    .A(_1591_),
    .B(_1874_),
    .C(_1899_));
 sg13g2_a221oi_1 _2630_ (.B2(_1874_),
    .C1(_1900_),
    .B1(_1897_),
    .A1(_1891_),
    .Y(_1901_),
    .A2(_1894_));
 sg13g2_nand2b_1 _2631_ (.Y(_1902_),
    .B(_1901_),
    .A_N(_1888_));
 sg13g2_a21o_1 _2632_ (.A2(_1814_),
    .A1(net132),
    .B1(_1815_),
    .X(_1903_));
 sg13g2_buf_2 _2633_ (.A(_1903_),
    .X(_1904_));
 sg13g2_nand3_1 _2634_ (.B(net132),
    .C(net98),
    .A(net99),
    .Y(_1905_));
 sg13g2_and2_1 _2635_ (.A(_1904_),
    .B(_1905_),
    .X(_1906_));
 sg13g2_xor2_1 _2636_ (.B(net145),
    .A(_1823_),
    .X(_1907_));
 sg13g2_o21ai_1 _2637_ (.B1(_1907_),
    .Y(_1908_),
    .A1(net106),
    .A2(_1836_));
 sg13g2_a21o_1 _2638_ (.A2(_1524_),
    .A1(net132),
    .B1(net145),
    .X(_1909_));
 sg13g2_a22oi_1 _2639_ (.Y(_1910_),
    .B1(_1825_),
    .B2(net103),
    .A2(_1909_),
    .A1(net61));
 sg13g2_o21ai_1 _2640_ (.B1(_1910_),
    .Y(_1911_),
    .A1(_1838_),
    .A2(_1908_));
 sg13g2_nor2b_1 _2641_ (.A(_1815_),
    .B_N(net132),
    .Y(_1912_));
 sg13g2_and2_1 _2642_ (.A(_1809_),
    .B(_1814_),
    .X(_1913_));
 sg13g2_buf_1 _2643_ (.A(_0059_),
    .X(_1914_));
 sg13g2_nor2b_1 _2644_ (.A(net100),
    .B_N(net129),
    .Y(_1915_));
 sg13g2_nand3b_1 _2645_ (.B(net132),
    .C(_1814_),
    .Y(_1916_),
    .A_N(_1815_));
 sg13g2_buf_2 _2646_ (.A(_1916_),
    .X(_1917_));
 sg13g2_nor2b_1 _2647_ (.A(net129),
    .B_N(net100),
    .Y(_1918_));
 sg13g2_a221oi_1 _2648_ (.B2(_1917_),
    .C1(_1918_),
    .B1(_1915_),
    .A1(_1912_),
    .Y(_1919_),
    .A2(_1913_));
 sg13g2_nor2_1 _2649_ (.A(_1524_),
    .B(net139),
    .Y(_1920_));
 sg13g2_xnor2_1 _2650_ (.Y(_1921_),
    .A(net132),
    .B(net98));
 sg13g2_mux2_1 _2651_ (.A0(net139),
    .A1(_1920_),
    .S(_1921_),
    .X(_1922_));
 sg13g2_nor2_1 _2652_ (.A(_1919_),
    .B(_1922_),
    .Y(_1923_));
 sg13g2_nand3_1 _2653_ (.B(_1911_),
    .C(_1923_),
    .A(_1906_),
    .Y(_1924_));
 sg13g2_nand3_1 _2654_ (.B(_1911_),
    .C(_1923_),
    .A(net104),
    .Y(_1925_));
 sg13g2_nand3_1 _2655_ (.B(_1904_),
    .C(_1905_),
    .A(net109),
    .Y(_1926_));
 sg13g2_nor2_1 _2656_ (.A(_1922_),
    .B(_1926_),
    .Y(_1927_));
 sg13g2_inv_2 _2657_ (.Y(_1928_),
    .A(net143));
 sg13g2_nor2_1 _2658_ (.A(_1624_),
    .B(_1928_),
    .Y(_1929_));
 sg13g2_nor2b_1 _2659_ (.A(_1922_),
    .B_N(_1929_),
    .Y(_1930_));
 sg13g2_o21ai_1 _2660_ (.B1(_1911_),
    .Y(_1931_),
    .A1(_1927_),
    .A2(_1930_));
 sg13g2_nand3_1 _2661_ (.B(_1904_),
    .C(_1905_),
    .A(net104),
    .Y(_1932_));
 sg13g2_a21oi_1 _2662_ (.A1(_1624_),
    .A2(_1932_),
    .Y(_1933_),
    .B1(_1919_));
 sg13g2_a21oi_1 _2663_ (.A1(_1906_),
    .A2(_1929_),
    .Y(_1934_),
    .B1(_1933_));
 sg13g2_nand4_1 _2664_ (.B(_1925_),
    .C(_1931_),
    .A(_1924_),
    .Y(_1935_),
    .D(_1934_));
 sg13g2_xnor2_1 _2665_ (.Y(_1936_),
    .A(_1624_),
    .B(_1919_));
 sg13g2_xnor2_1 _2666_ (.Y(_1937_),
    .A(net130),
    .B(net106));
 sg13g2_nand2b_1 _2667_ (.Y(_1938_),
    .B(net146),
    .A_N(\vga.paddle_l_pos_v[0] ));
 sg13g2_nand4_1 _2668_ (.B(_1907_),
    .C(_1836_),
    .A(_1937_),
    .Y(_1939_),
    .D(_1938_));
 sg13g2_and3_1 _2669_ (.X(_1940_),
    .A(_1860_),
    .B(_1862_),
    .C(_1809_));
 sg13g2_buf_1 _2670_ (.A(_1940_),
    .X(_1941_));
 sg13g2_inv_2 _2671_ (.Y(_1942_),
    .A(_1868_));
 sg13g2_a21oi_1 _2672_ (.A1(_1904_),
    .A2(_1941_),
    .Y(_1943_),
    .B1(_1942_));
 sg13g2_a21oi_1 _2673_ (.A1(_1822_),
    .A2(_1814_),
    .Y(_1944_),
    .B1(net99));
 sg13g2_nand3_1 _2674_ (.B(net95),
    .C(net100),
    .A(_1860_),
    .Y(_1945_));
 sg13g2_buf_1 _2675_ (.A(_1945_),
    .X(_1946_));
 sg13g2_nor3_1 _2676_ (.A(_1868_),
    .B(_1944_),
    .C(_1946_),
    .Y(_1947_));
 sg13g2_nand2_1 _2677_ (.Y(_1948_),
    .A(_1603_),
    .B(net142));
 sg13g2_nor3_1 _2678_ (.A(_1943_),
    .B(_1947_),
    .C(_1948_),
    .Y(_1949_));
 sg13g2_and2_1 _2679_ (.A(net98),
    .B(net139),
    .X(_1950_));
 sg13g2_nor2_1 _2680_ (.A(net98),
    .B(net139),
    .Y(_1951_));
 sg13g2_xor2_1 _2681_ (.B(net143),
    .A(_1815_),
    .X(_1952_));
 sg13g2_mux2_1 _2682_ (.A0(_1950_),
    .A1(_1951_),
    .S(_1952_),
    .X(_1953_));
 sg13g2_xnor2_1 _2683_ (.Y(_1954_),
    .A(net98),
    .B(net139));
 sg13g2_nor2_1 _2684_ (.A(net97),
    .B(_1954_),
    .Y(_1955_));
 sg13g2_a22oi_1 _2685_ (.Y(_1956_),
    .B1(_1955_),
    .B2(_1952_),
    .A2(_1953_),
    .A1(net97));
 sg13g2_nor4_2 _2686_ (.A(_1936_),
    .B(_1939_),
    .C(_1949_),
    .Y(_1957_),
    .D(_1956_));
 sg13g2_or2_1 _2687_ (.X(_1958_),
    .B(net142),
    .A(net111));
 sg13g2_nand2_1 _2688_ (.Y(_1959_),
    .A(_1904_),
    .B(_1941_));
 sg13g2_mux2_1 _2689_ (.A0(_1603_),
    .A1(_1958_),
    .S(_1959_),
    .X(_1960_));
 sg13g2_o21ai_1 _2690_ (.B1(_1821_),
    .Y(_1961_),
    .A1(net111),
    .A2(\vga.ball_pos_v[8] ));
 sg13g2_inv_1 _2691_ (.Y(_1962_),
    .A(net129));
 sg13g2_a21o_1 _2692_ (.A2(_1961_),
    .A1(_1904_),
    .B1(_1962_),
    .X(_1963_));
 sg13g2_a221oi_1 _2693_ (.B2(_1941_),
    .C1(_1942_),
    .B1(_1963_),
    .A1(net111),
    .Y(_1964_),
    .A2(_1959_));
 sg13g2_a21oi_1 _2694_ (.A1(_1942_),
    .A2(_1960_),
    .Y(_1965_),
    .B1(_1964_));
 sg13g2_nand2_1 _2695_ (.Y(_1966_),
    .A(_1863_),
    .B(_1810_));
 sg13g2_and2_1 _2696_ (.A(_1860_),
    .B(net129),
    .X(_1967_));
 sg13g2_a22oi_1 _2697_ (.Y(_1968_),
    .B1(_1967_),
    .B2(_1917_),
    .A2(_1966_),
    .A1(_1860_));
 sg13g2_buf_1 _2698_ (.A(_1968_),
    .X(_1969_));
 sg13g2_nand3b_1 _2699_ (.B(_1863_),
    .C(_1810_),
    .Y(_1970_),
    .A_N(_1860_));
 sg13g2_a21o_1 _2700_ (.A2(_1917_),
    .A1(net129),
    .B1(_1970_),
    .X(_1971_));
 sg13g2_a21o_1 _2701_ (.A2(_1971_),
    .A1(_1969_),
    .B1(_1573_),
    .X(_1972_));
 sg13g2_nand3_1 _2702_ (.B(_1969_),
    .C(_1971_),
    .A(_1573_),
    .Y(_1973_));
 sg13g2_and2_1 _2703_ (.A(_1972_),
    .B(_1973_),
    .X(_1974_));
 sg13g2_nand2_1 _2704_ (.Y(_1975_),
    .A(_1822_),
    .B(_1814_));
 sg13g2_nor2b_1 _2705_ (.A(net99),
    .B_N(net95),
    .Y(_1976_));
 sg13g2_nor2b_1 _2706_ (.A(net95),
    .B_N(net100),
    .Y(_1977_));
 sg13g2_nor2b_1 _2707_ (.A(net100),
    .B_N(net95),
    .Y(_1978_));
 sg13g2_a221oi_1 _2708_ (.B2(_1904_),
    .C1(_1978_),
    .B1(_1977_),
    .A1(_1975_),
    .Y(_1979_),
    .A2(_1976_));
 sg13g2_buf_1 _2709_ (.A(_1979_),
    .X(_1980_));
 sg13g2_xnor2_1 _2710_ (.Y(_1981_),
    .A(_1895_),
    .B(_1980_));
 sg13g2_nor4_2 _2711_ (.A(_1957_),
    .B(_1965_),
    .C(_1974_),
    .Y(_1982_),
    .D(_1981_));
 sg13g2_a21oi_1 _2712_ (.A1(_1972_),
    .A2(_1973_),
    .Y(_1983_),
    .B1(_1981_));
 sg13g2_buf_1 _2713_ (.A(\vga.ball_pos_v[6] ),
    .X(_1984_));
 sg13g2_a21o_1 _2714_ (.A2(_1980_),
    .A1(net128),
    .B1(net102),
    .X(_1985_));
 sg13g2_nand3_1 _2715_ (.B(_1971_),
    .C(_1985_),
    .A(_1969_),
    .Y(_1986_));
 sg13g2_nand3_1 _2716_ (.B(_1914_),
    .C(_1941_),
    .A(_1821_),
    .Y(_1987_));
 sg13g2_o21ai_1 _2717_ (.B1(_1942_),
    .Y(_1988_),
    .A1(_1944_),
    .A2(_1946_));
 sg13g2_o21ai_1 _2718_ (.B1(_1988_),
    .Y(_1989_),
    .A1(_1942_),
    .A2(_1987_));
 sg13g2_and2_1 _2719_ (.A(_1572_),
    .B(net128),
    .X(_1990_));
 sg13g2_buf_1 _2720_ (.A(_1990_),
    .X(_1991_));
 sg13g2_a22oi_1 _2721_ (.Y(_1992_),
    .B1(_1991_),
    .B2(_1980_),
    .A2(_1989_),
    .A1(net142));
 sg13g2_a221oi_1 _2722_ (.B2(_1992_),
    .C1(_1965_),
    .B1(_1986_),
    .A1(_1957_),
    .Y(_1993_),
    .A2(_1983_));
 sg13g2_a21oi_2 _2723_ (.B1(_1993_),
    .Y(_1994_),
    .A2(_1982_),
    .A1(_1935_));
 sg13g2_nor3_1 _2724_ (.A(_1740_),
    .B(net136),
    .C(\vga.ball_pos_h[6] ),
    .Y(_1995_));
 sg13g2_nand3b_1 _2725_ (.B(_1746_),
    .C(_1995_),
    .Y(_1996_),
    .A_N(_1739_));
 sg13g2_buf_1 _2726_ (.A(_1996_),
    .X(_1997_));
 sg13g2_buf_1 _2727_ (.A(\vga.ball_pos_h[1] ),
    .X(_1998_));
 sg13g2_nand2b_1 _2728_ (.Y(_1999_),
    .B(net138),
    .A_N(_1998_));
 sg13g2_nor3_1 _2729_ (.A(_1735_),
    .B(_1997_),
    .C(_1999_),
    .Y(_2000_));
 sg13g2_buf_2 _2730_ (.A(_2000_),
    .X(_2001_));
 sg13g2_and2_1 _2731_ (.A(_1730_),
    .B(_2001_),
    .X(_2002_));
 sg13g2_buf_2 _2732_ (.A(_2002_),
    .X(_2003_));
 sg13g2_nand2_1 _2733_ (.Y(_2004_),
    .A(_1729_),
    .B(_2003_));
 sg13g2_a21oi_1 _2734_ (.A1(_1902_),
    .A2(_1994_),
    .Y(_2005_),
    .B1(_2004_));
 sg13g2_buf_2 _2735_ (.A(_2005_),
    .X(_2006_));
 sg13g2_nand2_1 _2736_ (.Y(_2007_),
    .A(\vga.score_r[4] ),
    .B(net135));
 sg13g2_a21oi_1 _2737_ (.A1(net133),
    .A2(_2006_),
    .Y(_2008_),
    .B1(_2007_));
 sg13g2_buf_2 _2738_ (.A(\vga.score_r[2] ),
    .X(_2009_));
 sg13g2_inv_1 _2739_ (.Y(_2010_),
    .A(\vga.score_r[4] ));
 sg13g2_nor2_1 _2740_ (.A(_2009_),
    .B(_2010_),
    .Y(_2011_));
 sg13g2_inv_1 _2741_ (.Y(_2012_),
    .A(_2009_));
 sg13g2_buf_1 _2742_ (.A(\vga.score_r[1] ),
    .X(_2013_));
 sg13g2_nand2_1 _2743_ (.Y(_2014_),
    .A(net126),
    .B(\vga.score_r[0] ));
 sg13g2_nor3_1 _2744_ (.A(_2012_),
    .B(\vga.score_r[4] ),
    .C(_2014_),
    .Y(_2015_));
 sg13g2_o21ai_1 _2745_ (.B1(net133),
    .Y(_2016_),
    .A1(_2011_),
    .A2(_2015_));
 sg13g2_nor2_1 _2746_ (.A(\vga.score_r[3] ),
    .B(_2012_),
    .Y(_2017_));
 sg13g2_o21ai_1 _2747_ (.B1(\vga.score_r[4] ),
    .Y(_2018_),
    .A1(_2014_),
    .A2(_2017_));
 sg13g2_a21o_1 _2748_ (.A2(_1994_),
    .A1(_1902_),
    .B1(_2004_),
    .X(_2019_));
 sg13g2_buf_1 _2749_ (.A(_2019_),
    .X(_2020_));
 sg13g2_a21oi_1 _2750_ (.A1(_2016_),
    .A2(_2018_),
    .Y(_2021_),
    .B1(_2020_));
 sg13g2_nor2_1 _2751_ (.A(_2008_),
    .B(_2021_),
    .Y(_2022_));
 sg13g2_buf_1 _2752_ (.A(_2022_),
    .X(_2023_));
 sg13g2_nor2b_1 _2753_ (.A(_1767_),
    .B_N(net133),
    .Y(_2024_));
 sg13g2_buf_1 _2754_ (.A(\vga.score_r[0] ),
    .X(_2025_));
 sg13g2_nand3_1 _2755_ (.B(net125),
    .C(_2009_),
    .A(_2013_),
    .Y(_2026_));
 sg13g2_nand2_1 _2756_ (.Y(_2027_),
    .A(_1808_),
    .B(_2026_));
 sg13g2_or2_1 _2757_ (.X(_2028_),
    .B(_2026_),
    .A(_1808_));
 sg13g2_a221oi_1 _2758_ (.B2(_2028_),
    .C1(_2004_),
    .B1(_2027_),
    .A1(_1902_),
    .Y(_2029_),
    .A2(_1994_));
 sg13g2_a21oi_1 _2759_ (.A1(_2020_),
    .A2(_2024_),
    .Y(_2030_),
    .B1(_2029_));
 sg13g2_inv_2 _2760_ (.Y(_2031_),
    .A(_2030_));
 sg13g2_nor2b_1 _2761_ (.A(_1888_),
    .B_N(_1901_),
    .Y(_2032_));
 sg13g2_a21o_1 _2762_ (.A2(_1982_),
    .A1(_1935_),
    .B1(_1993_),
    .X(_2033_));
 sg13g2_or4_1 _2763_ (.A(_1708_),
    .B(_1716_),
    .C(_1719_),
    .D(_1728_),
    .X(_2034_));
 sg13g2_buf_1 _2764_ (.A(_2034_),
    .X(_2035_));
 sg13g2_nand2_1 _2765_ (.Y(_2036_),
    .A(_1730_),
    .B(_2001_));
 sg13g2_nor4_2 _2766_ (.A(\vga.score_r[3] ),
    .B(_2009_),
    .C(_2010_),
    .Y(_2037_),
    .D(_2014_));
 sg13g2_nor3_1 _2767_ (.A(_2035_),
    .B(_2036_),
    .C(_2037_),
    .Y(_2038_));
 sg13g2_o21ai_1 _2768_ (.B1(_2038_),
    .Y(_2039_),
    .A1(_2032_),
    .A2(_2033_));
 sg13g2_and2_1 _2769_ (.A(net135),
    .B(_2039_),
    .X(_2040_));
 sg13g2_inv_1 _2770_ (.Y(_2041_),
    .A(net125));
 sg13g2_nand2_1 _2771_ (.Y(_2042_),
    .A(_2013_),
    .B(_2041_));
 sg13g2_inv_1 _2772_ (.Y(_2043_),
    .A(net126));
 sg13g2_nand2_1 _2773_ (.Y(_2044_),
    .A(_2043_),
    .B(net125));
 sg13g2_a21oi_1 _2774_ (.A1(_2042_),
    .A2(_2044_),
    .Y(_2045_),
    .B1(_2020_));
 sg13g2_a21oi_1 _2775_ (.A1(net126),
    .A2(_2040_),
    .Y(_2046_),
    .B1(_2045_));
 sg13g2_buf_8 _2776_ (.A(_2046_),
    .X(_2047_));
 sg13g2_xnor2_1 _2777_ (.Y(_2048_),
    .A(net41),
    .B(_2047_));
 sg13g2_nor3_1 _2778_ (.A(_1772_),
    .B(_2012_),
    .C(_1767_),
    .Y(_2049_));
 sg13g2_a221oi_1 _2779_ (.B2(_2035_),
    .C1(_2012_),
    .B1(_1767_),
    .A1(net126),
    .Y(_2050_),
    .A2(net125));
 sg13g2_nor3_1 _2780_ (.A(_2009_),
    .B(_2035_),
    .C(_2014_),
    .Y(_2051_));
 sg13g2_nor3_1 _2781_ (.A(_1771_),
    .B(_2036_),
    .C(_2037_),
    .Y(_2052_));
 sg13g2_o21ai_1 _2782_ (.B1(_2052_),
    .Y(_2053_),
    .A1(_2050_),
    .A2(_2051_));
 sg13g2_a21oi_1 _2783_ (.A1(_1902_),
    .A2(_1994_),
    .Y(_2054_),
    .B1(_2053_));
 sg13g2_a21oi_1 _2784_ (.A1(_2020_),
    .A2(_2049_),
    .Y(_2055_),
    .B1(_2054_));
 sg13g2_buf_2 _2785_ (.A(_2055_),
    .X(_2056_));
 sg13g2_buf_1 _2786_ (.A(_2056_),
    .X(_2057_));
 sg13g2_and3_1 _2787_ (.X(_2058_),
    .A(net125),
    .B(_1768_),
    .C(_2039_));
 sg13g2_buf_2 _2788_ (.A(_2058_),
    .X(_2059_));
 sg13g2_nor2_2 _2789_ (.A(_2032_),
    .B(_2033_),
    .Y(_2060_));
 sg13g2_buf_1 _2790_ (.A(_1730_),
    .X(_2061_));
 sg13g2_nor3_1 _2791_ (.A(_1735_),
    .B(_1997_),
    .C(_1999_),
    .Y(_2062_));
 sg13g2_nand3_1 _2792_ (.B(_1729_),
    .C(_2062_),
    .A(net94),
    .Y(_2063_));
 sg13g2_nor3_2 _2793_ (.A(net125),
    .B(_2060_),
    .C(_2063_),
    .Y(_2064_));
 sg13g2_nor2_2 _2794_ (.A(_2059_),
    .B(_2064_),
    .Y(_2065_));
 sg13g2_nand2_1 _2795_ (.Y(_2066_),
    .A(net37),
    .B(_2065_));
 sg13g2_inv_2 _2796_ (.Y(_0207_),
    .A(_2056_));
 sg13g2_or2_1 _2797_ (.X(_2067_),
    .B(_2064_),
    .A(_2059_));
 sg13g2_buf_2 _2798_ (.A(_2067_),
    .X(_2068_));
 sg13g2_buf_1 _2799_ (.A(_2030_),
    .X(_2069_));
 sg13g2_a21o_1 _2800_ (.A2(_2040_),
    .A1(net126),
    .B1(_2045_),
    .X(_2070_));
 sg13g2_buf_1 _2801_ (.A(_2070_),
    .X(_2071_));
 sg13g2_nand4_1 _2802_ (.B(_2068_),
    .C(net40),
    .A(net36),
    .Y(_2072_),
    .D(_2071_));
 sg13g2_o21ai_1 _2803_ (.B1(_2072_),
    .Y(_2073_),
    .A1(_2048_),
    .A2(_2066_));
 sg13g2_nand2_1 _2804_ (.Y(_2074_),
    .A(net40),
    .B(_2047_));
 sg13g2_nand3b_1 _2805_ (.B(_2056_),
    .C(_2068_),
    .Y(_2075_),
    .A_N(net38));
 sg13g2_buf_1 _2806_ (.A(_1801_),
    .X(_2076_));
 sg13g2_o21ai_1 _2807_ (.B1(net93),
    .Y(_2077_),
    .A1(_2074_),
    .A2(_2075_));
 sg13g2_a21oi_1 _2808_ (.A1(net38),
    .A2(_2073_),
    .Y(_0006_),
    .B1(_2077_));
 sg13g2_nand3_1 _2809_ (.B(net41),
    .C(net35),
    .A(_2022_),
    .Y(_2078_));
 sg13g2_a21oi_1 _2810_ (.A1(_2074_),
    .A2(_2078_),
    .Y(_2079_),
    .B1(net36));
 sg13g2_nand2_1 _2811_ (.Y(_2080_),
    .A(net38),
    .B(net35));
 sg13g2_nor3_1 _2812_ (.A(net37),
    .B(net41),
    .C(_2080_),
    .Y(_2081_));
 sg13g2_o21ai_1 _2813_ (.B1(_1770_),
    .Y(_2082_),
    .A1(_2059_),
    .A2(_2064_));
 sg13g2_inv_1 _2814_ (.Y(_0205_),
    .A(_2082_));
 sg13g2_o21ai_1 _2815_ (.B1(_0205_),
    .Y(_0007_),
    .A1(_2079_),
    .A2(_2081_));
 sg13g2_nor2_1 _2816_ (.A(_1807_),
    .B(net34),
    .Y(_2083_));
 sg13g2_nor2b_1 _2817_ (.A(net31),
    .B_N(_2083_),
    .Y(_2084_));
 sg13g2_nor2b_1 _2818_ (.A(net33),
    .B_N(net39),
    .Y(_2085_));
 sg13g2_nor2_1 _2819_ (.A(_0198_),
    .B(_1800_),
    .Y(_2086_));
 sg13g2_and2_1 _2820_ (.A(_1795_),
    .B(_1798_),
    .X(_2087_));
 sg13g2_buf_8 _2821_ (.A(_2087_),
    .X(_2088_));
 sg13g2_nor3_1 _2822_ (.A(net31),
    .B(_1782_),
    .C(_2088_),
    .Y(_2089_));
 sg13g2_a21o_1 _2823_ (.A2(_2086_),
    .A1(_0200_),
    .B1(_2089_),
    .X(_2090_));
 sg13g2_a22oi_1 _2824_ (.Y(_0004_),
    .B1(_2085_),
    .B2(_2090_),
    .A2(_2084_),
    .A1(_1803_));
 sg13g2_nor2_1 _2825_ (.A(net31),
    .B(_2088_),
    .Y(_2091_));
 sg13g2_xnor2_1 _2826_ (.Y(_2092_),
    .A(_1782_),
    .B(net33));
 sg13g2_a22oi_1 _2827_ (.Y(_2093_),
    .B1(_2091_),
    .B2(_2092_),
    .A2(_2088_),
    .A1(_1788_));
 sg13g2_nand2b_1 _2828_ (.Y(_0005_),
    .B(_0196_),
    .A_N(_2093_));
 sg13g2_o21ai_1 _2829_ (.B1(_1770_),
    .Y(_2094_),
    .A1(_2008_),
    .A2(_2021_));
 sg13g2_buf_1 _2830_ (.A(_2094_),
    .X(_2095_));
 sg13g2_inv_1 _2831_ (.Y(_0209_),
    .A(_2095_));
 sg13g2_nand2_1 _2832_ (.Y(_2096_),
    .A(_2065_),
    .B(net40));
 sg13g2_nor4_1 _2833_ (.A(net36),
    .B(net40),
    .C(_2071_),
    .D(_2082_),
    .Y(_2097_));
 sg13g2_a21o_1 _2834_ (.A2(_2096_),
    .A1(_0209_),
    .B1(_2097_),
    .X(_2098_));
 sg13g2_nand3_1 _2835_ (.B(_2069_),
    .C(net35),
    .A(_2068_),
    .Y(_2099_));
 sg13g2_nand4_1 _2836_ (.B(_2065_),
    .C(net41),
    .A(net36),
    .Y(_2100_),
    .D(net35));
 sg13g2_o21ai_1 _2837_ (.B1(_2100_),
    .Y(_2101_),
    .A1(net37),
    .A2(_2099_));
 sg13g2_nor4_1 _2838_ (.A(net37),
    .B(_2068_),
    .C(net41),
    .D(net35),
    .Y(_2102_));
 sg13g2_nor2_1 _2839_ (.A(net38),
    .B(net37),
    .Y(_2103_));
 sg13g2_nor4_1 _2840_ (.A(_2098_),
    .B(_2101_),
    .C(_2102_),
    .D(_2103_),
    .Y(_0012_));
 sg13g2_or2_1 _2841_ (.X(_2104_),
    .B(net133),
    .A(net125));
 sg13g2_nand2_1 _2842_ (.Y(_2105_),
    .A(net125),
    .B(_2009_));
 sg13g2_mux2_1 _2843_ (.A0(_2104_),
    .A1(_2105_),
    .S(_2006_),
    .X(_2106_));
 sg13g2_o21ai_1 _2844_ (.B1(net133),
    .Y(_2107_),
    .A1(_2025_),
    .A2(_2006_));
 sg13g2_and3_1 _2845_ (.X(_2108_),
    .A(net126),
    .B(_2106_),
    .C(_2107_));
 sg13g2_nand2_1 _2846_ (.Y(_2109_),
    .A(_2025_),
    .B(net133));
 sg13g2_mux2_1 _2847_ (.A0(_2104_),
    .A1(_2109_),
    .S(_2006_),
    .X(_2110_));
 sg13g2_o21ai_1 _2848_ (.B1(_2095_),
    .Y(_2111_),
    .A1(net126),
    .A2(_2110_));
 sg13g2_o21ai_1 _2849_ (.B1(_2006_),
    .Y(_2112_),
    .A1(_2012_),
    .A2(_2109_));
 sg13g2_o21ai_1 _2850_ (.B1(_2112_),
    .Y(_2113_),
    .A1(_1767_),
    .A2(_2006_));
 sg13g2_nand3_1 _2851_ (.B(_0207_),
    .C(_2113_),
    .A(net134),
    .Y(_2114_));
 sg13g2_or3_1 _2852_ (.A(_2108_),
    .B(_2111_),
    .C(_2114_),
    .X(_2115_));
 sg13g2_nor2_1 _2853_ (.A(_2031_),
    .B(_2047_),
    .Y(_2116_));
 sg13g2_o21ai_1 _2854_ (.B1(net37),
    .Y(_2117_),
    .A1(_2116_),
    .A2(_2082_));
 sg13g2_a22oi_1 _2855_ (.Y(_0013_),
    .B1(_2115_),
    .B2(_2117_),
    .A2(_2096_),
    .A1(_0209_));
 sg13g2_nand3b_1 _2856_ (.B(_2056_),
    .C(_2047_),
    .Y(_2118_),
    .A_N(_2022_));
 sg13g2_nand3_1 _2857_ (.B(net36),
    .C(net35),
    .A(net38),
    .Y(_2119_));
 sg13g2_a21oi_1 _2858_ (.A1(_2118_),
    .A2(_2119_),
    .Y(_2120_),
    .B1(_2096_));
 sg13g2_nand3_1 _2859_ (.B(_2069_),
    .C(_2047_),
    .A(net38),
    .Y(_2121_));
 sg13g2_a21oi_1 _2860_ (.A1(_2078_),
    .A2(_2121_),
    .Y(_2122_),
    .B1(_2065_));
 sg13g2_buf_1 _2861_ (.A(_1801_),
    .X(_2123_));
 sg13g2_o21ai_1 _2862_ (.B1(net92),
    .Y(_0002_),
    .A1(_2120_),
    .A2(_2122_));
 sg13g2_nand3_1 _2863_ (.B(_2068_),
    .C(net40),
    .A(_2056_),
    .Y(_2124_));
 sg13g2_nand3_1 _2864_ (.B(net36),
    .C(net41),
    .A(net38),
    .Y(_2125_));
 sg13g2_a21oi_1 _2865_ (.A1(_2124_),
    .A2(_2125_),
    .Y(_2126_),
    .B1(net35));
 sg13g2_nand2_1 _2866_ (.Y(_2127_),
    .A(net37),
    .B(_2068_));
 sg13g2_nor3_1 _2867_ (.A(_2056_),
    .B(_2059_),
    .C(_2064_),
    .Y(_2128_));
 sg13g2_nand2b_1 _2868_ (.Y(_2129_),
    .B(net40),
    .A_N(_2128_));
 sg13g2_a21oi_1 _2869_ (.A1(_2127_),
    .A2(_2129_),
    .Y(_2130_),
    .B1(_2080_));
 sg13g2_o21ai_1 _2870_ (.B1(net92),
    .Y(_0003_),
    .A1(_2126_),
    .A2(_2130_));
 sg13g2_a21o_1 _2871_ (.A2(_2086_),
    .A1(_0199_),
    .B1(net31),
    .X(_2131_));
 sg13g2_xnor2_1 _2872_ (.Y(_0217_),
    .A(net33),
    .B(_2088_));
 sg13g2_inv_1 _2873_ (.Y(_0218_),
    .A(_1774_));
 sg13g2_o21ai_1 _2874_ (.B1(_0218_),
    .Y(_0219_),
    .A1(net39),
    .A2(_0217_));
 sg13g2_nand2_1 _2875_ (.Y(_0220_),
    .A(_0200_),
    .B(net33));
 sg13g2_a21oi_2 _2876_ (.B1(_1791_),
    .Y(_0221_),
    .A2(_1790_),
    .A1(net148));
 sg13g2_nand2_1 _2877_ (.Y(_0222_),
    .A(_1755_),
    .B(net135));
 sg13g2_mux2_1 _2878_ (.A0(_1755_),
    .A1(_0222_),
    .S(_1794_),
    .X(_0223_));
 sg13g2_nor2_1 _2879_ (.A(_0223_),
    .B(_1782_),
    .Y(_0224_));
 sg13g2_nand3_1 _2880_ (.B(_1800_),
    .C(_0224_),
    .A(_0221_),
    .Y(_0225_));
 sg13g2_nand2_1 _2881_ (.Y(_0226_),
    .A(_0220_),
    .B(_0225_));
 sg13g2_a221oi_1 _2882_ (.B2(net34),
    .C1(_0226_),
    .B1(_0219_),
    .A1(net39),
    .Y(_0010_),
    .A2(_2131_));
 sg13g2_nor2_1 _2883_ (.A(net33),
    .B(_2088_),
    .Y(_0227_));
 sg13g2_nor3_1 _2884_ (.A(_1782_),
    .B(_0221_),
    .C(_1800_),
    .Y(_0228_));
 sg13g2_nor4_1 _2885_ (.A(_2083_),
    .B(_0224_),
    .C(_0227_),
    .D(_0228_),
    .Y(_0229_));
 sg13g2_nor2_1 _2886_ (.A(_0218_),
    .B(_2083_),
    .Y(_0230_));
 sg13g2_nor3_1 _2887_ (.A(_0226_),
    .B(_0229_),
    .C(_0230_),
    .Y(_0011_));
 sg13g2_and2_1 _2888_ (.A(_1774_),
    .B(_1782_),
    .X(_0231_));
 sg13g2_nor2_1 _2889_ (.A(net31),
    .B(_1782_),
    .Y(_0232_));
 sg13g2_a22oi_1 _2890_ (.Y(_0233_),
    .B1(_0232_),
    .B2(_0227_),
    .A2(_0231_),
    .A1(_1802_));
 sg13g2_or2_1 _2891_ (.X(_0234_),
    .B(_0217_),
    .A(_1774_));
 sg13g2_buf_1 _2892_ (.A(_0234_),
    .X(_0235_));
 sg13g2_mux2_1 _2893_ (.A0(_0233_),
    .A1(_0235_),
    .S(net39),
    .X(_0000_));
 sg13g2_nor2_1 _2894_ (.A(net101),
    .B(net31),
    .Y(_0236_));
 sg13g2_nor2_1 _2895_ (.A(net34),
    .B(_2088_),
    .Y(_0237_));
 sg13g2_a21o_1 _2896_ (.A2(_0237_),
    .A1(_0221_),
    .B1(_0228_),
    .X(_0238_));
 sg13g2_nand2_1 _2897_ (.Y(_0239_),
    .A(_0196_),
    .B(_1800_));
 sg13g2_a21oi_1 _2898_ (.A1(net34),
    .A2(net33),
    .Y(_0240_),
    .B1(_0239_));
 sg13g2_and3_1 _2899_ (.X(_0241_),
    .A(net39),
    .B(_1788_),
    .C(_2088_));
 sg13g2_a221oi_1 _2900_ (.B2(_0218_),
    .C1(_0241_),
    .B1(_0240_),
    .A1(_0236_),
    .Y(_0001_),
    .A2(_0238_));
 sg13g2_nand2b_1 _2901_ (.Y(_0242_),
    .B(net41),
    .A_N(_2023_));
 sg13g2_a22oi_1 _2902_ (.Y(_0243_),
    .B1(_0242_),
    .B2(net37),
    .A2(_2048_),
    .A1(_2023_));
 sg13g2_o21ai_1 _2903_ (.B1(_2123_),
    .Y(_0009_),
    .A1(_2068_),
    .A2(_0243_));
 sg13g2_inv_1 _2904_ (.Y(_0244_),
    .A(_0015_));
 sg13g2_buf_2 _2905_ (.A(\vga.count_v[1] ),
    .X(_0245_));
 sg13g2_buf_1 _2906_ (.A(_0245_),
    .X(_0246_));
 sg13g2_buf_1 _2907_ (.A(\vga.count_v[2] ),
    .X(_0247_));
 sg13g2_buf_1 _2908_ (.A(_0247_),
    .X(_0248_));
 sg13g2_buf_1 _2909_ (.A(\vga.count_v[3] ),
    .X(_0249_));
 sg13g2_buf_2 _2910_ (.A(\vga.count_v[5] ),
    .X(_0250_));
 sg13g2_nand2b_1 _2911_ (.Y(_0251_),
    .B(_0250_),
    .A_N(_0249_));
 sg13g2_buf_1 _2912_ (.A(\vga.count_v[4] ),
    .X(_0252_));
 sg13g2_buf_1 _2913_ (.A(\vga.count_v[0] ),
    .X(_0253_));
 sg13g2_buf_1 _2914_ (.A(_0253_),
    .X(_0254_));
 sg13g2_buf_2 _2915_ (.A(\vga.count_v[9] ),
    .X(_0255_));
 sg13g2_buf_1 _2916_ (.A(\vga.count_v[7] ),
    .X(_0256_));
 sg13g2_or2_1 _2917_ (.X(_0257_),
    .B(\vga.count_v[8] ),
    .A(_0256_));
 sg13g2_buf_1 _2918_ (.A(_0257_),
    .X(_0258_));
 sg13g2_nor4_2 _2919_ (.A(net89),
    .B(\vga.count_v[6] ),
    .C(_0255_),
    .Y(_0259_),
    .D(_0258_));
 sg13g2_nand2_1 _2920_ (.Y(_0260_),
    .A(_0252_),
    .B(_0259_));
 sg13g2_nor4_1 _2921_ (.A(net91),
    .B(net90),
    .C(_0251_),
    .D(_0260_),
    .Y(_0261_));
 sg13g2_buf_1 _2922_ (.A(_0261_),
    .X(_0262_));
 sg13g2_nand2_1 _2923_ (.Y(_0263_),
    .A(_0247_),
    .B(_0249_));
 sg13g2_or3_1 _2924_ (.A(net91),
    .B(_0250_),
    .C(_0263_),
    .X(_0264_));
 sg13g2_or2_1 _2925_ (.X(_0265_),
    .B(_0260_),
    .A(_0264_));
 sg13g2_buf_2 _2926_ (.A(_0265_),
    .X(_0266_));
 sg13g2_nor2b_1 _2927_ (.A(_0262_),
    .B_N(_0266_),
    .Y(_0267_));
 sg13g2_nand2b_1 _2928_ (.Y(_0268_),
    .B(_0262_),
    .A_N(_0028_));
 sg13g2_o21ai_1 _2929_ (.B1(_0268_),
    .Y(_0269_),
    .A1(_0018_),
    .A2(_0266_));
 sg13g2_a21oi_1 _2930_ (.A1(_0244_),
    .A2(_0267_),
    .Y(_0270_),
    .B1(_0269_));
 sg13g2_buf_1 _2931_ (.A(_0249_),
    .X(_0271_));
 sg13g2_buf_1 _2932_ (.A(net88),
    .X(_0272_));
 sg13g2_buf_1 _2933_ (.A(_0250_),
    .X(_0273_));
 sg13g2_xnor2_1 _2934_ (.Y(_0274_),
    .A(net59),
    .B(net87));
 sg13g2_nor2_1 _2935_ (.A(net91),
    .B(_0251_),
    .Y(_0275_));
 sg13g2_a21oi_1 _2936_ (.A1(net91),
    .A2(_0274_),
    .Y(_0276_),
    .B1(_0275_));
 sg13g2_o21ai_1 _2937_ (.B1(_0264_),
    .Y(_0277_),
    .A1(net90),
    .A2(_0276_));
 sg13g2_inv_1 _2938_ (.Y(_0278_),
    .A(_0247_));
 sg13g2_inv_1 _2939_ (.Y(_0279_),
    .A(_0250_));
 sg13g2_nand2b_1 _2940_ (.Y(_0280_),
    .B(_0245_),
    .A_N(_0249_));
 sg13g2_nor4_1 _2941_ (.A(net86),
    .B(_0279_),
    .C(_0252_),
    .D(_0280_),
    .Y(_0281_));
 sg13g2_a21oi_1 _2942_ (.A1(_0252_),
    .A2(_0277_),
    .Y(_0282_),
    .B1(_0281_));
 sg13g2_nor2b_1 _2943_ (.A(_0282_),
    .B_N(_0259_),
    .Y(_0283_));
 sg13g2_buf_2 _2944_ (.A(_0283_),
    .X(_0284_));
 sg13g2_mux2_1 _2945_ (.A0(\vga.score_l_unit_pixels[0] ),
    .A1(_0270_),
    .S(_0284_),
    .X(_0202_));
 sg13g2_and2_1 _2946_ (.A(_0259_),
    .B(_0281_),
    .X(_0285_));
 sg13g2_buf_1 _2947_ (.A(_0285_),
    .X(_0286_));
 sg13g2_or2_1 _2948_ (.X(_0287_),
    .B(_0286_),
    .A(_0262_));
 sg13g2_buf_1 _2949_ (.A(_0287_),
    .X(_0288_));
 sg13g2_nand2b_1 _2950_ (.Y(_0289_),
    .B(_0286_),
    .A_N(_0024_));
 sg13g2_o21ai_1 _2951_ (.B1(_0289_),
    .Y(_0290_),
    .A1(_0032_),
    .A2(_0288_));
 sg13g2_nor2_1 _2952_ (.A(_0019_),
    .B(_0267_),
    .Y(_0291_));
 sg13g2_a21oi_1 _2953_ (.A1(_0266_),
    .A2(_0290_),
    .Y(_0292_),
    .B1(_0291_));
 sg13g2_or4_1 _2954_ (.A(net90),
    .B(net87),
    .C(_0280_),
    .D(_0260_),
    .X(_0293_));
 sg13g2_buf_2 _2955_ (.A(_0293_),
    .X(_0294_));
 sg13g2_mux2_1 _2956_ (.A0(_0014_),
    .A1(_0292_),
    .S(_0294_),
    .X(_0295_));
 sg13g2_mux2_1 _2957_ (.A0(\vga.score_l_unit_pixels[1] ),
    .A1(_0295_),
    .S(_0284_),
    .X(_0203_));
 sg13g2_inv_1 _2958_ (.Y(_0296_),
    .A(_0033_));
 sg13g2_a22oi_1 _2959_ (.Y(_0297_),
    .B1(_0286_),
    .B2(_0025_),
    .A2(_0262_),
    .A1(_0029_));
 sg13g2_o21ai_1 _2960_ (.B1(_0297_),
    .Y(_0298_),
    .A1(_0296_),
    .A2(_0288_));
 sg13g2_mux2_1 _2961_ (.A0(_0020_),
    .A1(_0298_),
    .S(_0266_),
    .X(_0299_));
 sg13g2_nor2_1 _2962_ (.A(_0244_),
    .B(_0294_),
    .Y(_0300_));
 sg13g2_a21oi_1 _2963_ (.A1(_0294_),
    .A2(_0299_),
    .Y(_0301_),
    .B1(_0300_));
 sg13g2_nor2_1 _2964_ (.A(\vga.score_l_unit_pixels[2] ),
    .B(_0284_),
    .Y(_0302_));
 sg13g2_a21oi_1 _2965_ (.A1(_0284_),
    .A2(_0301_),
    .Y(_0204_),
    .B1(_0302_));
 sg13g2_inv_1 _2966_ (.Y(_0303_),
    .A(_0017_));
 sg13g2_nand2b_1 _2967_ (.Y(_0304_),
    .B(_0262_),
    .A_N(_0030_));
 sg13g2_o21ai_1 _2968_ (.B1(_0304_),
    .Y(_0305_),
    .A1(_0021_),
    .A2(_0266_));
 sg13g2_a21oi_1 _2969_ (.A1(_0303_),
    .A2(_0267_),
    .Y(_0306_),
    .B1(_0305_));
 sg13g2_mux2_1 _2970_ (.A0(\vga.score_r_unit_pixels[0] ),
    .A1(_0306_),
    .S(_0284_),
    .X(_0211_));
 sg13g2_nand2b_1 _2971_ (.Y(_0307_),
    .B(_0286_),
    .A_N(_0026_));
 sg13g2_o21ai_1 _2972_ (.B1(_0307_),
    .Y(_0308_),
    .A1(_0034_),
    .A2(_0288_));
 sg13g2_nor2_1 _2973_ (.A(_0022_),
    .B(_0267_),
    .Y(_0309_));
 sg13g2_a21oi_1 _2974_ (.A1(_0266_),
    .A2(_0308_),
    .Y(_0310_),
    .B1(_0309_));
 sg13g2_mux2_1 _2975_ (.A0(_0016_),
    .A1(_0310_),
    .S(_0294_),
    .X(_0311_));
 sg13g2_mux2_1 _2976_ (.A0(\vga.score_r_unit_pixels[1] ),
    .A1(_0311_),
    .S(_0284_),
    .X(_0212_));
 sg13g2_inv_1 _2977_ (.Y(_0312_),
    .A(_0035_));
 sg13g2_a22oi_1 _2978_ (.Y(_0313_),
    .B1(_0286_),
    .B2(_0027_),
    .A2(_0262_),
    .A1(_0031_));
 sg13g2_o21ai_1 _2979_ (.B1(_0313_),
    .Y(_0314_),
    .A1(_0312_),
    .A2(_0288_));
 sg13g2_mux2_1 _2980_ (.A0(_0023_),
    .A1(_0314_),
    .S(_0266_),
    .X(_0315_));
 sg13g2_nor2_1 _2981_ (.A(_0303_),
    .B(_0294_),
    .Y(_0316_));
 sg13g2_a21oi_1 _2982_ (.A1(_0294_),
    .A2(_0315_),
    .Y(_0317_),
    .B1(_0316_));
 sg13g2_nor2_1 _2983_ (.A(\vga.score_r_unit_pixels[2] ),
    .B(_0284_),
    .Y(_0318_));
 sg13g2_a21oi_1 _2984_ (.A1(_0284_),
    .A2(_0317_),
    .Y(_0213_),
    .B1(_0318_));
 sg13g2_buf_1 _2985_ (.A(_1729_),
    .X(_0319_));
 sg13g2_mux2_1 _2986_ (.A0(\vga.left_down_1d ),
    .A1(net2),
    .S(net50),
    .X(_0169_));
 sg13g2_mux2_1 _2987_ (.A0(\vga.left_up_1d ),
    .A1(net1),
    .S(net50),
    .X(_0171_));
 sg13g2_mux2_1 _2988_ (.A0(\vga.right_down_1d ),
    .A1(net4),
    .S(net50),
    .X(_0192_));
 sg13g2_mux2_1 _2989_ (.A0(\vga.right_up_1d ),
    .A1(net3),
    .S(net50),
    .X(_0194_));
 sg13g2_o21ai_1 _2990_ (.B1(_2020_),
    .Y(_0320_),
    .A1(_2041_),
    .A2(_1767_));
 sg13g2_nor3_1 _2991_ (.A(_1767_),
    .B(_2006_),
    .C(_2042_),
    .Y(_0321_));
 sg13g2_a21oi_1 _2992_ (.A1(_2043_),
    .A2(_0320_),
    .Y(_0322_),
    .B1(_0321_));
 sg13g2_nor3_1 _2993_ (.A(net133),
    .B(_0207_),
    .C(_0322_),
    .Y(_0323_));
 sg13g2_o21ai_1 _2994_ (.B1(_2128_),
    .Y(_0324_),
    .A1(_1772_),
    .A2(_2047_));
 sg13g2_nand3_1 _2995_ (.B(_2068_),
    .C(net35),
    .A(_2056_),
    .Y(_0325_));
 sg13g2_a21oi_1 _2996_ (.A1(_0324_),
    .A2(_0325_),
    .Y(_0326_),
    .B1(net40));
 sg13g2_buf_1 _2997_ (.A(net101),
    .X(_0327_));
 sg13g2_nor3_1 _2998_ (.A(net58),
    .B(_2008_),
    .C(_2021_),
    .Y(_0328_));
 sg13g2_o21ai_1 _2999_ (.B1(_0328_),
    .Y(_0085_),
    .A1(_0323_),
    .A2(_0326_));
 sg13g2_nor2_1 _3000_ (.A(net101),
    .B(_2047_),
    .Y(_0206_));
 sg13g2_xnor2_1 _3001_ (.Y(_0329_),
    .A(net41),
    .B(_0206_));
 sg13g2_and4_1 _3002_ (.A(_2057_),
    .B(_0205_),
    .C(_2095_),
    .D(_0329_),
    .X(_0086_));
 sg13g2_nand4_1 _3003_ (.B(_0205_),
    .C(_2095_),
    .A(_2057_),
    .Y(_0087_),
    .D(_0329_));
 sg13g2_nand2_1 _3004_ (.Y(_0330_),
    .A(_1807_),
    .B(_1782_));
 sg13g2_or2_1 _3005_ (.X(_0088_),
    .B(_0330_),
    .A(_0235_));
 sg13g2_xnor2_1 _3006_ (.Y(_0331_),
    .A(net39),
    .B(_1792_));
 sg13g2_and2_1 _3007_ (.A(_0237_),
    .B(_0331_),
    .X(_0332_));
 sg13g2_nand2b_1 _3008_ (.Y(_0333_),
    .B(net34),
    .A_N(_1807_));
 sg13g2_mux2_1 _3009_ (.A0(_0333_),
    .A1(_0330_),
    .S(_0221_),
    .X(_0334_));
 sg13g2_nor2_1 _3010_ (.A(_1800_),
    .B(_0334_),
    .Y(_0335_));
 sg13g2_o21ai_1 _3011_ (.B1(_0236_),
    .Y(_0089_),
    .A1(_0332_),
    .A2(_0335_));
 sg13g2_nor2_1 _3012_ (.A(_0235_),
    .B(_0330_),
    .Y(_0090_));
 sg13g2_or2_1 _3013_ (.X(_0091_),
    .B(_0235_),
    .A(_0333_));
 sg13g2_nand2_1 _3014_ (.Y(_0336_),
    .A(net38),
    .B(_2065_));
 sg13g2_o21ai_1 _3015_ (.B1(net93),
    .Y(_0337_),
    .A1(_2048_),
    .A2(_0336_));
 sg13g2_nand2_1 _3016_ (.Y(_0092_),
    .A(net36),
    .B(_0337_));
 sg13g2_buf_1 _3017_ (.A(net101),
    .X(_0338_));
 sg13g2_buf_1 _3018_ (.A(\vga.count_h[8] ),
    .X(_0339_));
 sg13g2_buf_1 _3019_ (.A(_0339_),
    .X(_0340_));
 sg13g2_buf_1 _3020_ (.A(\vga.count_h[7] ),
    .X(_0341_));
 sg13g2_inv_2 _3021_ (.Y(_0342_),
    .A(\vga.count_h[9] ));
 sg13g2_nor3_1 _3022_ (.A(net85),
    .B(_0341_),
    .C(_0342_),
    .Y(_0343_));
 sg13g2_buf_1 _3023_ (.A(\vga.count_h[5] ),
    .X(_0344_));
 sg13g2_buf_2 _3024_ (.A(\vga.count_h[6] ),
    .X(_0345_));
 sg13g2_nand2_1 _3025_ (.Y(_0346_),
    .A(_0344_),
    .B(_0345_));
 sg13g2_buf_1 _3026_ (.A(\vga.count_h[4] ),
    .X(_0347_));
 sg13g2_buf_1 _3027_ (.A(_0347_),
    .X(_0348_));
 sg13g2_buf_2 _3028_ (.A(\vga.count_h[0] ),
    .X(_0349_));
 sg13g2_inv_2 _3029_ (.Y(_0350_),
    .A(_0349_));
 sg13g2_buf_1 _3030_ (.A(\vga.count_h[3] ),
    .X(_0351_));
 sg13g2_inv_2 _3031_ (.Y(_0352_),
    .A(net124));
 sg13g2_buf_1 _3032_ (.A(\vga.count_h[2] ),
    .X(_0353_));
 sg13g2_buf_1 _3033_ (.A(\vga.count_h[1] ),
    .X(_0354_));
 sg13g2_nand2_2 _3034_ (.Y(_0355_),
    .A(net123),
    .B(net122));
 sg13g2_nor3_2 _3035_ (.A(_0350_),
    .B(_0352_),
    .C(_0355_),
    .Y(_0356_));
 sg13g2_nand2_1 _3036_ (.Y(_0357_),
    .A(net84),
    .B(_0356_));
 sg13g2_nor2_2 _3037_ (.A(_0346_),
    .B(_0357_),
    .Y(_0358_));
 sg13g2_buf_1 _3038_ (.A(_0066_),
    .X(_0359_));
 sg13g2_nor2_1 _3039_ (.A(_0359_),
    .B(_0343_),
    .Y(_0360_));
 sg13g2_a21oi_1 _3040_ (.A1(_0343_),
    .A2(_0358_),
    .Y(_0361_),
    .B1(_0360_));
 sg13g2_buf_1 _3041_ (.A(_0341_),
    .X(_0362_));
 sg13g2_buf_1 _3042_ (.A(_0344_),
    .X(_0363_));
 sg13g2_nor3_1 _3043_ (.A(_0363_),
    .B(_0345_),
    .C(net84),
    .Y(_0364_));
 sg13g2_nor2_1 _3044_ (.A(_0339_),
    .B(_0342_),
    .Y(_0365_));
 sg13g2_nand3_1 _3045_ (.B(_0356_),
    .C(_0364_),
    .A(_0365_),
    .Y(_0366_));
 sg13g2_o21ai_1 _3046_ (.B1(_0366_),
    .Y(_0367_),
    .A1(_0359_),
    .A2(_0364_));
 sg13g2_nor2_1 _3047_ (.A(_0359_),
    .B(_0365_),
    .Y(_0368_));
 sg13g2_a21oi_1 _3048_ (.A1(net83),
    .A2(_0367_),
    .Y(_0369_),
    .B1(_0368_));
 sg13g2_inv_2 _3049_ (.Y(_0370_),
    .A(_0347_));
 sg13g2_nand3_1 _3050_ (.B(_0365_),
    .C(_0356_),
    .A(_0370_),
    .Y(_0371_));
 sg13g2_o21ai_1 _3051_ (.B1(_0371_),
    .Y(_0372_),
    .A1(_0370_),
    .A2(_0359_));
 sg13g2_nand4_1 _3052_ (.B(net82),
    .C(_0345_),
    .A(_0362_),
    .Y(_0373_),
    .D(_0372_));
 sg13g2_nand2b_1 _3053_ (.Y(_0374_),
    .B(_0373_),
    .A_N(_0368_));
 sg13g2_nor4_1 _3054_ (.A(net57),
    .B(_0361_),
    .C(_0369_),
    .D(_0374_),
    .Y(_0143_));
 sg13g2_inv_1 _3055_ (.Y(_0375_),
    .A(_0083_));
 sg13g2_xnor2_1 _3056_ (.Y(_0376_),
    .A(net5),
    .B(\vga.speed_lsb_1d ));
 sg13g2_buf_1 _3057_ (.A(ui_in[6]),
    .X(_0377_));
 sg13g2_xnor2_1 _3058_ (.Y(_0378_),
    .A(_0377_),
    .B(\vga.speed_msb_1d ));
 sg13g2_nand2_1 _3059_ (.Y(_0379_),
    .A(_1702_),
    .B(_1721_));
 sg13g2_or4_1 _3060_ (.A(\vga.interval_counter[4] ),
    .B(_1699_),
    .C(_1725_),
    .D(_1726_),
    .X(_0380_));
 sg13g2_nand2b_1 _3061_ (.Y(_0381_),
    .B(\vga.interval_counter[10] ),
    .A_N(\vga.interval_counter[11] ));
 sg13g2_nor3_1 _3062_ (.A(_1709_),
    .B(_1710_),
    .C(_0381_),
    .Y(_0382_));
 sg13g2_nor2_1 _3063_ (.A(net5),
    .B(_1704_),
    .Y(_0383_));
 sg13g2_nand4_1 _3064_ (.B(_1705_),
    .C(_0382_),
    .A(_1713_),
    .Y(_0384_),
    .D(_0383_));
 sg13g2_and4_1 _3065_ (.A(_1706_),
    .B(_1722_),
    .C(_1724_),
    .D(_1711_),
    .X(_0385_));
 sg13g2_buf_1 _3066_ (.A(_0385_),
    .X(_0386_));
 sg13g2_nand4_1 _3067_ (.B(_1720_),
    .C(_1714_),
    .A(_1701_),
    .Y(_0387_),
    .D(_0386_));
 sg13g2_nor4_1 _3068_ (.A(_0379_),
    .B(_0380_),
    .C(_0384_),
    .D(_0387_),
    .Y(_0388_));
 sg13g2_nand4_1 _3069_ (.B(_1706_),
    .C(_1703_),
    .A(\vga.interval_counter[4] ),
    .Y(_0389_),
    .D(_1723_));
 sg13g2_nand4_1 _3070_ (.B(_1710_),
    .C(_1713_),
    .A(net5),
    .Y(_0390_),
    .D(_1714_));
 sg13g2_nor2b_1 _3071_ (.A(_1699_),
    .B_N(_1704_),
    .Y(_0391_));
 sg13g2_inv_1 _3072_ (.Y(_0392_),
    .A(_1709_));
 sg13g2_nand2_1 _3073_ (.Y(_0393_),
    .A(\vga.interval_counter[11] ),
    .B(\vga.interval_counter[10] ));
 sg13g2_nor3_1 _3074_ (.A(_0392_),
    .B(_1705_),
    .C(_0393_),
    .Y(_0394_));
 sg13g2_nand4_1 _3075_ (.B(_1727_),
    .C(_0391_),
    .A(_1711_),
    .Y(_0395_),
    .D(_0394_));
 sg13g2_nor3_1 _3076_ (.A(_0389_),
    .B(_0390_),
    .C(_0395_),
    .Y(_0396_));
 sg13g2_nor2_1 _3077_ (.A(_0388_),
    .B(_0396_),
    .Y(_0397_));
 sg13g2_nand4_1 _3078_ (.B(_1720_),
    .C(_1721_),
    .A(_1709_),
    .Y(_0398_),
    .D(_1722_));
 sg13g2_nor4_1 _3079_ (.A(_1708_),
    .B(_0381_),
    .C(_0390_),
    .D(_0398_),
    .Y(_0399_));
 sg13g2_nor4_1 _3080_ (.A(_1714_),
    .B(_1700_),
    .C(_0384_),
    .D(_0389_),
    .Y(_0400_));
 sg13g2_nand2_1 _3081_ (.Y(_0401_),
    .A(_0377_),
    .B(_1724_));
 sg13g2_nor4_1 _3082_ (.A(_1711_),
    .B(_1725_),
    .C(_1726_),
    .D(_0401_),
    .Y(_0402_));
 sg13g2_o21ai_1 _3083_ (.B1(_0402_),
    .Y(_0403_),
    .A1(_0399_),
    .A2(_0400_));
 sg13g2_o21ai_1 _3084_ (.B1(_0403_),
    .Y(_0404_),
    .A1(_0377_),
    .A2(_0397_));
 sg13g2_nand2b_1 _3085_ (.Y(_0405_),
    .B(_0404_),
    .A_N(_1719_));
 sg13g2_nand4_1 _3086_ (.B(_0376_),
    .C(_0378_),
    .A(net134),
    .Y(_0406_),
    .D(_0405_));
 sg13g2_buf_1 _3087_ (.A(_0406_),
    .X(_0407_));
 sg13g2_buf_1 _3088_ (.A(_0407_),
    .X(_0408_));
 sg13g2_nor2_1 _3089_ (.A(_0375_),
    .B(net44),
    .Y(_0144_));
 sg13g2_inv_1 _3090_ (.Y(_0409_),
    .A(\vga.interval_counter[10] ));
 sg13g2_nand4_1 _3091_ (.B(_1704_),
    .C(_1709_),
    .A(_1701_),
    .Y(_0410_),
    .D(_1720_));
 sg13g2_buf_1 _3092_ (.A(_0410_),
    .X(_0411_));
 sg13g2_nor3_2 _3093_ (.A(_1698_),
    .B(_0379_),
    .C(_0411_),
    .Y(_0412_));
 sg13g2_nand4_1 _3094_ (.B(_1713_),
    .C(_1714_),
    .A(_1710_),
    .Y(_0413_),
    .D(_0412_));
 sg13g2_xnor2_1 _3095_ (.Y(_0414_),
    .A(_0409_),
    .B(_0413_));
 sg13g2_nor2_1 _3096_ (.A(net44),
    .B(_0414_),
    .Y(_0145_));
 sg13g2_nor2_1 _3097_ (.A(_0409_),
    .B(_0413_),
    .Y(_0415_));
 sg13g2_xnor2_1 _3098_ (.Y(_0416_),
    .A(\vga.interval_counter[11] ),
    .B(_0415_));
 sg13g2_nor2_1 _3099_ (.A(net44),
    .B(_0416_),
    .Y(_0146_));
 sg13g2_nor2_1 _3100_ (.A(_0393_),
    .B(_0413_),
    .Y(_0417_));
 sg13g2_xnor2_1 _3101_ (.Y(_0418_),
    .A(_1705_),
    .B(_0417_));
 sg13g2_nor2_1 _3102_ (.A(net44),
    .B(_0418_),
    .Y(_0147_));
 sg13g2_and2_1 _3103_ (.A(_1705_),
    .B(_0417_),
    .X(_0419_));
 sg13g2_xnor2_1 _3104_ (.Y(_0420_),
    .A(_1699_),
    .B(_0419_));
 sg13g2_nor2_1 _3105_ (.A(net44),
    .B(_0420_),
    .Y(_0148_));
 sg13g2_and2_1 _3106_ (.A(_1699_),
    .B(_0419_),
    .X(_0421_));
 sg13g2_buf_2 _3107_ (.A(_0421_),
    .X(_0422_));
 sg13g2_xnor2_1 _3108_ (.Y(_0423_),
    .A(_1722_),
    .B(_0422_));
 sg13g2_nor2_1 _3109_ (.A(net44),
    .B(_0423_),
    .Y(_0149_));
 sg13g2_nand2_1 _3110_ (.Y(_0424_),
    .A(_1722_),
    .B(_0422_));
 sg13g2_xor2_1 _3111_ (.B(_0424_),
    .A(_1706_),
    .X(_0425_));
 sg13g2_nor2_1 _3112_ (.A(net44),
    .B(_0425_),
    .Y(_0150_));
 sg13g2_nand3_1 _3113_ (.B(_1722_),
    .C(_0422_),
    .A(_1706_),
    .Y(_0426_));
 sg13g2_xor2_1 _3114_ (.B(_0426_),
    .A(_1724_),
    .X(_0427_));
 sg13g2_nor2_1 _3115_ (.A(net44),
    .B(_0427_),
    .Y(_0151_));
 sg13g2_nand4_1 _3116_ (.B(_1722_),
    .C(_1724_),
    .A(_1706_),
    .Y(_0428_),
    .D(_0422_));
 sg13g2_xor2_1 _3117_ (.B(_0428_),
    .A(_1711_),
    .X(_0429_));
 sg13g2_nor2_1 _3118_ (.A(_0408_),
    .B(_0429_),
    .Y(_0152_));
 sg13g2_nand2_1 _3119_ (.Y(_0430_),
    .A(_0386_),
    .B(_0422_));
 sg13g2_xor2_1 _3120_ (.B(_0430_),
    .A(_1726_),
    .X(_0431_));
 sg13g2_nor2_1 _3121_ (.A(_0408_),
    .B(_0431_),
    .Y(_0153_));
 sg13g2_buf_1 _3122_ (.A(_0407_),
    .X(_0432_));
 sg13g2_nand3_1 _3123_ (.B(_0386_),
    .C(_0422_),
    .A(_1726_),
    .Y(_0433_));
 sg13g2_xor2_1 _3124_ (.B(_0433_),
    .A(_1725_),
    .X(_0434_));
 sg13g2_nor2_1 _3125_ (.A(net43),
    .B(_0434_),
    .Y(_0154_));
 sg13g2_xnor2_1 _3126_ (.Y(_0435_),
    .A(_1701_),
    .B(_1704_));
 sg13g2_nor2_1 _3127_ (.A(net43),
    .B(_0435_),
    .Y(_0155_));
 sg13g2_and4_1 _3128_ (.A(_1725_),
    .B(_1726_),
    .C(_0386_),
    .D(_0422_),
    .X(_0436_));
 sg13g2_buf_1 _3129_ (.A(_0436_),
    .X(_0437_));
 sg13g2_xnor2_1 _3130_ (.Y(_0438_),
    .A(_1717_),
    .B(_0437_));
 sg13g2_nor2_1 _3131_ (.A(net43),
    .B(_0438_),
    .Y(_0156_));
 sg13g2_nand2_1 _3132_ (.Y(_0439_),
    .A(_1717_),
    .B(_0437_));
 sg13g2_xor2_1 _3133_ (.B(_0439_),
    .A(\vga.interval_counter[21] ),
    .X(_0440_));
 sg13g2_nor2_1 _3134_ (.A(net43),
    .B(_0440_),
    .Y(_0157_));
 sg13g2_inv_1 _3135_ (.Y(_0441_),
    .A(\vga.interval_counter[22] ));
 sg13g2_nand3_1 _3136_ (.B(_1717_),
    .C(_0437_),
    .A(\vga.interval_counter[21] ),
    .Y(_0442_));
 sg13g2_xnor2_1 _3137_ (.Y(_0443_),
    .A(_0441_),
    .B(_0442_));
 sg13g2_nor2_1 _3138_ (.A(net43),
    .B(_0443_),
    .Y(_0158_));
 sg13g2_nor2_1 _3139_ (.A(_0441_),
    .B(_0442_),
    .Y(_0444_));
 sg13g2_xnor2_1 _3140_ (.Y(_0445_),
    .A(\vga.interval_counter[23] ),
    .B(_0444_));
 sg13g2_nor2_1 _3141_ (.A(_0432_),
    .B(_0445_),
    .Y(_0159_));
 sg13g2_nand2_1 _3142_ (.Y(_0446_),
    .A(\vga.interval_counter[23] ),
    .B(_0444_));
 sg13g2_xor2_1 _3143_ (.B(_0446_),
    .A(\vga.interval_counter[24] ),
    .X(_0447_));
 sg13g2_nor2_1 _3144_ (.A(_0432_),
    .B(_0447_),
    .Y(_0160_));
 sg13g2_nand2_1 _3145_ (.Y(_0448_),
    .A(_1701_),
    .B(_1704_));
 sg13g2_xor2_1 _3146_ (.B(_0448_),
    .A(_1720_),
    .X(_0449_));
 sg13g2_nor2_1 _3147_ (.A(net43),
    .B(_0449_),
    .Y(_0161_));
 sg13g2_nand3_1 _3148_ (.B(_1704_),
    .C(_1720_),
    .A(_1701_),
    .Y(_0450_));
 sg13g2_xnor2_1 _3149_ (.Y(_0451_),
    .A(_0392_),
    .B(_0450_));
 sg13g2_nor2_1 _3150_ (.A(net43),
    .B(_0451_),
    .Y(_0162_));
 sg13g2_xnor2_1 _3151_ (.Y(_0452_),
    .A(_1698_),
    .B(_0411_));
 sg13g2_nor2_1 _3152_ (.A(net43),
    .B(_0452_),
    .Y(_0163_));
 sg13g2_nor2_1 _3153_ (.A(_1698_),
    .B(_0411_),
    .Y(_0453_));
 sg13g2_xnor2_1 _3154_ (.Y(_0454_),
    .A(_1702_),
    .B(_0453_));
 sg13g2_nor2_1 _3155_ (.A(_0407_),
    .B(_0454_),
    .Y(_0164_));
 sg13g2_nand2_1 _3156_ (.Y(_0455_),
    .A(_1702_),
    .B(_0453_));
 sg13g2_xor2_1 _3157_ (.B(_0455_),
    .A(_1721_),
    .X(_0456_));
 sg13g2_nor2_1 _3158_ (.A(_0407_),
    .B(_0456_),
    .Y(_0165_));
 sg13g2_xnor2_1 _3159_ (.Y(_0457_),
    .A(_1710_),
    .B(_0412_));
 sg13g2_nor2_1 _3160_ (.A(_0407_),
    .B(_0457_),
    .Y(_0166_));
 sg13g2_nand2_1 _3161_ (.Y(_0458_),
    .A(_1710_),
    .B(_0412_));
 sg13g2_xor2_1 _3162_ (.B(_0458_),
    .A(_1713_),
    .X(_0459_));
 sg13g2_nor2_1 _3163_ (.A(_0407_),
    .B(_0459_),
    .Y(_0167_));
 sg13g2_nand3_1 _3164_ (.B(_1713_),
    .C(_0412_),
    .A(_1710_),
    .Y(_0460_));
 sg13g2_xor2_1 _3165_ (.B(_0460_),
    .A(_1714_),
    .X(_0461_));
 sg13g2_nor2_1 _3166_ (.A(_0407_),
    .B(_0461_),
    .Y(_0168_));
 sg13g2_and3_1 _3167_ (.X(_0170_),
    .A(\vga.left_down_1d ),
    .B(net2),
    .C(net50));
 sg13g2_and3_1 _3168_ (.X(_0172_),
    .A(\vga.left_up_1d ),
    .B(net1),
    .C(net50));
 sg13g2_buf_2 _3169_ (.A(_0052_),
    .X(_0462_));
 sg13g2_nand3_1 _3170_ (.B(_1733_),
    .C(_1734_),
    .A(net127),
    .Y(_0463_));
 sg13g2_buf_1 _3171_ (.A(_0463_),
    .X(_0464_));
 sg13g2_and2_1 _3172_ (.A(_0462_),
    .B(_0464_),
    .X(_0465_));
 sg13g2_buf_1 _3173_ (.A(_1733_),
    .X(_0466_));
 sg13g2_buf_1 _3174_ (.A(_1734_),
    .X(_0467_));
 sg13g2_nand4_1 _3175_ (.B(net81),
    .C(net80),
    .A(net127),
    .Y(_0468_),
    .D(_1740_));
 sg13g2_nor2_1 _3176_ (.A(_0462_),
    .B(_0468_),
    .Y(_0469_));
 sg13g2_nand2_1 _3177_ (.Y(_0470_),
    .A(_1731_),
    .B(net136));
 sg13g2_a22oi_1 _3178_ (.Y(_0471_),
    .B1(_0469_),
    .B2(_0470_),
    .A2(_0465_),
    .A1(_1743_));
 sg13g2_buf_1 _3179_ (.A(_0046_),
    .X(_0472_));
 sg13g2_buf_1 _3180_ (.A(_1740_),
    .X(_0473_));
 sg13g2_nand2_1 _3181_ (.Y(_0474_),
    .A(net79),
    .B(net136));
 sg13g2_or2_1 _3182_ (.X(_0475_),
    .B(_0464_),
    .A(_0474_));
 sg13g2_nor2_1 _3183_ (.A(_0472_),
    .B(_0475_),
    .Y(_0476_));
 sg13g2_nand2_1 _3184_ (.Y(_0477_),
    .A(_0472_),
    .B(_0475_));
 sg13g2_nor2_1 _3185_ (.A(net137),
    .B(_0477_),
    .Y(_0478_));
 sg13g2_a21oi_1 _3186_ (.A1(net137),
    .A2(_0476_),
    .Y(_0479_),
    .B1(_0478_));
 sg13g2_nand3_1 _3187_ (.B(net136),
    .C(_1738_),
    .A(_1740_),
    .Y(_0480_));
 sg13g2_buf_1 _3188_ (.A(_0480_),
    .X(_0481_));
 sg13g2_nand3_1 _3189_ (.B(_1745_),
    .C(_1739_),
    .A(_1744_),
    .Y(_0482_));
 sg13g2_nor4_2 _3190_ (.A(_0057_),
    .B(_1735_),
    .C(_0481_),
    .Y(_0483_),
    .D(_0482_));
 sg13g2_buf_1 _3191_ (.A(_0047_),
    .X(_0484_));
 sg13g2_o21ai_1 _3192_ (.B1(_0484_),
    .Y(_0485_),
    .A1(_0481_),
    .A2(_0464_));
 sg13g2_buf_1 _3193_ (.A(_1745_),
    .X(_0486_));
 sg13g2_nand2b_1 _3194_ (.Y(_0487_),
    .B(net78),
    .A_N(_1744_));
 sg13g2_buf_1 _3195_ (.A(_1744_),
    .X(_0488_));
 sg13g2_inv_1 _3196_ (.Y(_0489_),
    .A(_0484_));
 sg13g2_nor2_1 _3197_ (.A(_0481_),
    .B(_0464_),
    .Y(_0490_));
 sg13g2_buf_1 _3198_ (.A(_0490_),
    .X(_0491_));
 sg13g2_o21ai_1 _3199_ (.B1(_1745_),
    .Y(_0492_),
    .A1(_1731_),
    .A2(_1742_));
 sg13g2_nand4_1 _3200_ (.B(_0489_),
    .C(_0491_),
    .A(net77),
    .Y(_0493_),
    .D(_0492_));
 sg13g2_o21ai_1 _3201_ (.B1(_0493_),
    .Y(_0494_),
    .A1(_0485_),
    .A2(_0487_));
 sg13g2_nor2_1 _3202_ (.A(_0483_),
    .B(_0494_),
    .Y(_0495_));
 sg13g2_o21ai_1 _3203_ (.B1(_0495_),
    .Y(_0496_),
    .A1(_0471_),
    .A2(_0479_));
 sg13g2_nor2_1 _3204_ (.A(_0472_),
    .B(_0471_),
    .Y(_0497_));
 sg13g2_nand3_1 _3205_ (.B(_0491_),
    .C(_0497_),
    .A(_0483_),
    .Y(_0498_));
 sg13g2_a21oi_1 _3206_ (.A1(_0484_),
    .A2(_0491_),
    .Y(_0499_),
    .B1(net78));
 sg13g2_a21oi_1 _3207_ (.A1(net78),
    .A2(_0485_),
    .Y(_0500_),
    .B1(net77));
 sg13g2_nor2_1 _3208_ (.A(_0499_),
    .B(_0500_),
    .Y(_0501_));
 sg13g2_nor3_1 _3209_ (.A(_0481_),
    .B(_0482_),
    .C(_0464_),
    .Y(_0502_));
 sg13g2_nor2_1 _3210_ (.A(_0483_),
    .B(_0502_),
    .Y(_0503_));
 sg13g2_o21ai_1 _3211_ (.B1(_0503_),
    .Y(_0504_),
    .A1(_1739_),
    .A2(_0501_));
 sg13g2_nand3_1 _3212_ (.B(_0498_),
    .C(_0504_),
    .A(_0496_),
    .Y(_0505_));
 sg13g2_nand3_1 _3213_ (.B(net78),
    .C(_0491_),
    .A(net77),
    .Y(_0506_));
 sg13g2_xnor2_1 _3214_ (.Y(_0507_),
    .A(_1739_),
    .B(_0506_));
 sg13g2_xnor2_1 _3215_ (.Y(_0508_),
    .A(_0494_),
    .B(_0507_));
 sg13g2_xnor2_1 _3216_ (.Y(_0509_),
    .A(_0359_),
    .B(_0508_));
 sg13g2_xor2_1 _3217_ (.B(_0497_),
    .A(net77),
    .X(_0510_));
 sg13g2_nor3_1 _3218_ (.A(net137),
    .B(_0471_),
    .C(_0477_),
    .Y(_0511_));
 sg13g2_a21oi_1 _3219_ (.A1(_0491_),
    .A2(_0510_),
    .Y(_0512_),
    .B1(_0511_));
 sg13g2_xnor2_1 _3220_ (.Y(_0513_),
    .A(_0484_),
    .B(_0512_));
 sg13g2_nand2b_1 _3221_ (.Y(_0514_),
    .B(_0054_),
    .A_N(_0513_));
 sg13g2_buf_1 _3222_ (.A(net138),
    .X(_0515_));
 sg13g2_nand2_1 _3223_ (.Y(_0516_),
    .A(net76),
    .B(_0491_));
 sg13g2_xnor2_1 _3224_ (.Y(_0517_),
    .A(_0472_),
    .B(_0516_));
 sg13g2_nor2_1 _3225_ (.A(net83),
    .B(_0517_),
    .Y(_0518_));
 sg13g2_nor2_1 _3226_ (.A(net138),
    .B(_0462_),
    .Y(_0519_));
 sg13g2_nor2_1 _3227_ (.A(_0464_),
    .B(_0519_),
    .Y(_0520_));
 sg13g2_mux2_1 _3228_ (.A0(_0465_),
    .A1(_0520_),
    .S(_1740_),
    .X(_0521_));
 sg13g2_mux2_1 _3229_ (.A0(_0469_),
    .A1(_0521_),
    .S(net136),
    .X(_0522_));
 sg13g2_xnor2_1 _3230_ (.Y(_0523_),
    .A(net137),
    .B(_0522_));
 sg13g2_xor2_1 _3231_ (.B(_0053_),
    .A(_1734_),
    .X(_0524_));
 sg13g2_nand2b_1 _3232_ (.Y(_0525_),
    .B(_0349_),
    .A_N(net138));
 sg13g2_nor2b_1 _3233_ (.A(net122),
    .B_N(net127),
    .Y(_0526_));
 sg13g2_nand2b_1 _3234_ (.Y(_0527_),
    .B(net122),
    .A_N(net127));
 sg13g2_o21ai_1 _3235_ (.B1(_0527_),
    .Y(_0528_),
    .A1(_0525_),
    .A2(_0526_));
 sg13g2_a21oi_1 _3236_ (.A1(net138),
    .A2(_1998_),
    .Y(_0529_),
    .B1(net80));
 sg13g2_nor2_1 _3237_ (.A(_1732_),
    .B(_0524_),
    .Y(_0530_));
 sg13g2_a221oi_1 _3238_ (.B2(net123),
    .C1(_0530_),
    .B1(_0529_),
    .A1(_0524_),
    .Y(_0531_),
    .A2(_0528_));
 sg13g2_nand3_1 _3239_ (.B(net127),
    .C(net80),
    .A(net138),
    .Y(_0532_));
 sg13g2_and2_1 _3240_ (.A(net81),
    .B(_0532_),
    .X(_0533_));
 sg13g2_o21ai_1 _3241_ (.B1(_0533_),
    .Y(_0534_),
    .A1(_0352_),
    .A2(_0531_));
 sg13g2_a21o_1 _3242_ (.A2(_0528_),
    .A1(_0524_),
    .B1(_0530_),
    .X(_0535_));
 sg13g2_inv_1 _3243_ (.Y(_0536_),
    .A(net123));
 sg13g2_o21ai_1 _3244_ (.B1(net124),
    .Y(_0537_),
    .A1(net81),
    .A2(_0532_));
 sg13g2_nor3_1 _3245_ (.A(net124),
    .B(net81),
    .C(_0529_),
    .Y(_0538_));
 sg13g2_a21oi_1 _3246_ (.A1(_0536_),
    .A2(_0537_),
    .Y(_0539_),
    .B1(_0538_));
 sg13g2_or2_1 _3247_ (.X(_0540_),
    .B(_0539_),
    .A(_0535_));
 sg13g2_inv_1 _3248_ (.Y(_0541_),
    .A(net81));
 sg13g2_nand3b_1 _3249_ (.B(_0541_),
    .C(_0352_),
    .Y(_0542_),
    .A_N(_0532_));
 sg13g2_inv_1 _3250_ (.Y(_0543_),
    .A(_1740_));
 sg13g2_xnor2_1 _3251_ (.Y(_0544_),
    .A(_0543_),
    .B(_1737_));
 sg13g2_nand2b_1 _3252_ (.Y(_0545_),
    .B(_0056_),
    .A_N(_0544_));
 sg13g2_and4_1 _3253_ (.A(_0534_),
    .B(_0540_),
    .C(_0542_),
    .D(_0545_),
    .X(_0546_));
 sg13g2_nor2b_1 _3254_ (.A(_0056_),
    .B_N(_0544_),
    .Y(_0547_));
 sg13g2_nor2_1 _3255_ (.A(_0543_),
    .B(_1737_),
    .Y(_0548_));
 sg13g2_xor2_1 _3256_ (.B(_0548_),
    .A(_0462_),
    .X(_0549_));
 sg13g2_xnor2_1 _3257_ (.Y(_0550_),
    .A(_0058_),
    .B(_0549_));
 sg13g2_o21ai_1 _3258_ (.B1(_0550_),
    .Y(_0551_),
    .A1(_0546_),
    .A2(_0547_));
 sg13g2_nand2_1 _3259_ (.Y(_0552_),
    .A(net82),
    .B(_0549_));
 sg13g2_inv_1 _3260_ (.Y(_0553_),
    .A(_0055_));
 sg13g2_xnor2_1 _3261_ (.Y(_0554_),
    .A(_0553_),
    .B(_0523_));
 sg13g2_a21oi_1 _3262_ (.A1(_0551_),
    .A2(_0552_),
    .Y(_0555_),
    .B1(_0554_));
 sg13g2_a221oi_1 _3263_ (.B2(_0345_),
    .C1(_0555_),
    .B1(_0523_),
    .A1(net83),
    .Y(_0556_),
    .A2(_0517_));
 sg13g2_nand2b_1 _3264_ (.Y(_0557_),
    .B(_0513_),
    .A_N(_0054_));
 sg13g2_o21ai_1 _3265_ (.B1(_0557_),
    .Y(_0558_),
    .A1(_0518_),
    .A2(_0556_));
 sg13g2_nand4_1 _3266_ (.B(_0509_),
    .C(_0514_),
    .A(_0505_),
    .Y(_0559_),
    .D(_0558_));
 sg13g2_buf_2 _3267_ (.A(_0042_),
    .X(_0560_));
 sg13g2_inv_2 _3268_ (.Y(_0561_),
    .A(_0560_));
 sg13g2_buf_1 _3269_ (.A(net106),
    .X(_0562_));
 sg13g2_nand2_2 _3270_ (.Y(_0563_),
    .A(net105),
    .B(net56));
 sg13g2_nor3_1 _3271_ (.A(_1928_),
    .B(_1525_),
    .C(_0563_),
    .Y(_0564_));
 sg13g2_xnor2_1 _3272_ (.Y(_0565_),
    .A(_1554_),
    .B(_0564_));
 sg13g2_buf_2 _3273_ (.A(_0038_),
    .X(_0566_));
 sg13g2_inv_2 _3274_ (.Y(_0567_),
    .A(_0253_));
 sg13g2_nand2_1 _3275_ (.Y(_0568_),
    .A(_0567_),
    .B(net146));
 sg13g2_nand2_1 _3276_ (.Y(_0569_),
    .A(net56),
    .B(_0568_));
 sg13g2_o21ai_1 _3277_ (.B1(_0245_),
    .Y(_0570_),
    .A1(net56),
    .A2(_0568_));
 sg13g2_nand3_1 _3278_ (.B(_0569_),
    .C(_0570_),
    .A(_0566_),
    .Y(_0571_));
 sg13g2_xor2_1 _3279_ (.B(_0039_),
    .A(net139),
    .X(_0572_));
 sg13g2_and2_1 _3280_ (.A(net105),
    .B(net56),
    .X(_0573_));
 sg13g2_buf_1 _3281_ (.A(_0573_),
    .X(_0574_));
 sg13g2_nand2_1 _3282_ (.Y(_0575_),
    .A(_0574_),
    .B(_0572_));
 sg13g2_o21ai_1 _3283_ (.B1(_0575_),
    .Y(_0576_),
    .A1(_1854_),
    .A2(_0572_));
 sg13g2_nor3_1 _3284_ (.A(_0566_),
    .B(_0574_),
    .C(_0572_),
    .Y(_0577_));
 sg13g2_nand2_1 _3285_ (.Y(_0578_),
    .A(_0569_),
    .B(_0570_));
 sg13g2_xnor2_1 _3286_ (.Y(_0579_),
    .A(net139),
    .B(_0563_));
 sg13g2_and2_1 _3287_ (.A(net88),
    .B(_0579_),
    .X(_0580_));
 sg13g2_a221oi_1 _3288_ (.B2(_0578_),
    .C1(_0580_),
    .B1(_0577_),
    .A1(_0571_),
    .Y(_0581_),
    .A2(_0576_));
 sg13g2_nand3_1 _3289_ (.B(net103),
    .C(_0574_),
    .A(net104),
    .Y(_0582_));
 sg13g2_buf_1 _3290_ (.A(_0582_),
    .X(_0583_));
 sg13g2_buf_2 _3291_ (.A(_0041_),
    .X(_0584_));
 sg13g2_xnor2_1 _3292_ (.Y(_0585_),
    .A(_1553_),
    .B(_0584_));
 sg13g2_nand2_1 _3293_ (.Y(_0586_),
    .A(_0583_),
    .B(_0585_));
 sg13g2_nand3_1 _3294_ (.B(_1658_),
    .C(_0562_),
    .A(net103),
    .Y(_0587_));
 sg13g2_nor2_1 _3295_ (.A(_0587_),
    .B(_0585_),
    .Y(_0588_));
 sg13g2_and2_1 _3296_ (.A(_1928_),
    .B(_0585_),
    .X(_0589_));
 sg13g2_a22oi_1 _3297_ (.Y(_0590_),
    .B1(_0589_),
    .B2(_0587_),
    .A2(_0588_),
    .A1(net104));
 sg13g2_o21ai_1 _3298_ (.B1(_0590_),
    .Y(_0591_),
    .A1(_0581_),
    .A2(_0586_));
 sg13g2_buf_1 _3299_ (.A(_0040_),
    .X(_0592_));
 sg13g2_inv_2 _3300_ (.Y(_0593_),
    .A(net121));
 sg13g2_nor2_1 _3301_ (.A(_0590_),
    .B(_0581_),
    .Y(_0594_));
 sg13g2_a221oi_1 _3302_ (.B2(_0593_),
    .C1(_0594_),
    .B1(_0591_),
    .A1(net87),
    .Y(_0595_),
    .A2(_0565_));
 sg13g2_buf_1 _3303_ (.A(\vga.count_v[6] ),
    .X(_0596_));
 sg13g2_nor2_1 _3304_ (.A(_1624_),
    .B(_0583_),
    .Y(_0597_));
 sg13g2_buf_1 _3305_ (.A(_0597_),
    .X(_0598_));
 sg13g2_xnor2_1 _3306_ (.Y(_0599_),
    .A(_1567_),
    .B(net47));
 sg13g2_nor2_1 _3307_ (.A(net120),
    .B(_0599_),
    .Y(_0600_));
 sg13g2_o21ai_1 _3308_ (.B1(_0600_),
    .Y(_0601_),
    .A1(_0561_),
    .A2(_0595_));
 sg13g2_o21ai_1 _3309_ (.B1(_0599_),
    .Y(_0602_),
    .A1(_0560_),
    .A2(_0595_));
 sg13g2_nand2_1 _3310_ (.Y(_0603_),
    .A(_1984_),
    .B(net47));
 sg13g2_xnor2_1 _3311_ (.Y(_0604_),
    .A(_0073_),
    .B(_0603_));
 sg13g2_buf_1 _3312_ (.A(_0256_),
    .X(_0605_));
 sg13g2_a22oi_1 _3313_ (.Y(_0606_),
    .B1(_0604_),
    .B2(net75),
    .A2(_0602_),
    .A1(_0601_));
 sg13g2_nand2_1 _3314_ (.Y(_0607_),
    .A(_1991_),
    .B(net47));
 sg13g2_buf_1 _3315_ (.A(_0065_),
    .X(_0608_));
 sg13g2_inv_1 _3316_ (.Y(_0609_),
    .A(_0608_));
 sg13g2_buf_1 _3317_ (.A(net142),
    .X(_0610_));
 sg13g2_buf_1 _3318_ (.A(_0044_),
    .X(_0611_));
 sg13g2_xor2_1 _3319_ (.B(net119),
    .A(net111),
    .X(_0612_));
 sg13g2_nand3_1 _3320_ (.B(net74),
    .C(_0612_),
    .A(_0609_),
    .Y(_0613_));
 sg13g2_a21oi_1 _3321_ (.A1(_1991_),
    .A2(net47),
    .Y(_0614_),
    .B1(_0612_));
 sg13g2_nand2b_1 _3322_ (.Y(_0615_),
    .B(_0612_),
    .A_N(net74));
 sg13g2_nor2_1 _3323_ (.A(_0607_),
    .B(_0615_),
    .Y(_0616_));
 sg13g2_buf_1 _3324_ (.A(_0608_),
    .X(_0617_));
 sg13g2_o21ai_1 _3325_ (.B1(net73),
    .Y(_0618_),
    .A1(_0614_),
    .A2(_0616_));
 sg13g2_o21ai_1 _3326_ (.B1(_0618_),
    .Y(_0619_),
    .A1(_0607_),
    .A2(_0613_));
 sg13g2_o21ai_1 _3327_ (.B1(_0619_),
    .Y(_0620_),
    .A1(net75),
    .A2(_0604_));
 sg13g2_or2_1 _3328_ (.X(_0621_),
    .B(_0620_),
    .A(_0606_));
 sg13g2_inv_2 _3329_ (.Y(_0622_),
    .A(net119));
 sg13g2_buf_1 _3330_ (.A(_0255_),
    .X(_0623_));
 sg13g2_nor3_1 _3331_ (.A(net103),
    .B(net105),
    .C(net106),
    .Y(_0624_));
 sg13g2_buf_2 _3332_ (.A(_0624_),
    .X(_0625_));
 sg13g2_nand2_1 _3333_ (.Y(_0626_),
    .A(_1928_),
    .B(_0625_));
 sg13g2_buf_2 _3334_ (.A(_0626_),
    .X(_0627_));
 sg13g2_nor4_2 _3335_ (.A(net102),
    .B(net109),
    .C(net128),
    .Y(_0628_),
    .D(_0627_));
 sg13g2_mux2_1 _3336_ (.A0(_1603_),
    .A1(_1948_),
    .S(_0628_),
    .X(_0629_));
 sg13g2_nor2b_1 _3337_ (.A(net74),
    .B_N(_0628_),
    .Y(_0630_));
 sg13g2_nand3_1 _3338_ (.B(_1603_),
    .C(_0630_),
    .A(net72),
    .Y(_0631_));
 sg13g2_o21ai_1 _3339_ (.B1(_0631_),
    .Y(_0632_),
    .A1(net72),
    .A2(_0629_));
 sg13g2_nand2_1 _3340_ (.Y(_0633_),
    .A(_0622_),
    .B(_0632_));
 sg13g2_nor3_1 _3341_ (.A(_1646_),
    .B(_1984_),
    .C(_0627_),
    .Y(_0634_));
 sg13g2_xnor2_1 _3342_ (.Y(_0635_),
    .A(_0073_),
    .B(_0634_));
 sg13g2_nor2_1 _3343_ (.A(net109),
    .B(_0627_),
    .Y(_0636_));
 sg13g2_xnor2_1 _3344_ (.Y(_0637_),
    .A(_1895_),
    .B(_0636_));
 sg13g2_xnor2_1 _3345_ (.Y(_0638_),
    .A(_1554_),
    .B(_0627_));
 sg13g2_xnor2_1 _3346_ (.Y(_0639_),
    .A(_0561_),
    .B(_0637_));
 sg13g2_a21oi_1 _3347_ (.A1(_0279_),
    .A2(_0638_),
    .Y(_0640_),
    .B1(_0639_));
 sg13g2_nand2b_1 _3348_ (.Y(_0641_),
    .B(_1666_),
    .A_N(_0625_));
 sg13g2_a21oi_1 _3349_ (.A1(_0627_),
    .A2(_0641_),
    .Y(_0642_),
    .B1(_0593_));
 sg13g2_and2_1 _3350_ (.A(net86),
    .B(_1854_),
    .X(_0643_));
 sg13g2_nand2_1 _3351_ (.Y(_0644_),
    .A(net88),
    .B(_0563_));
 sg13g2_o21ai_1 _3352_ (.B1(net103),
    .Y(_0645_),
    .A1(_0643_),
    .A2(_0644_));
 sg13g2_a21oi_1 _3353_ (.A1(_0248_),
    .A2(_0563_),
    .Y(_0646_),
    .B1(net88));
 sg13g2_nor2_1 _3354_ (.A(_0625_),
    .B(_0646_),
    .Y(_0647_));
 sg13g2_xnor2_1 _3355_ (.Y(_0648_),
    .A(_0249_),
    .B(net103));
 sg13g2_inv_1 _3356_ (.Y(_0649_),
    .A(_0566_));
 sg13g2_a21oi_1 _3357_ (.A1(_1854_),
    .A2(_0563_),
    .Y(_0650_),
    .B1(_0649_));
 sg13g2_a21oi_1 _3358_ (.A1(_0649_),
    .A2(_0563_),
    .Y(_0651_),
    .B1(_0650_));
 sg13g2_nor3_1 _3359_ (.A(_0566_),
    .B(_1854_),
    .C(_0648_),
    .Y(_0652_));
 sg13g2_a21o_1 _3360_ (.A2(_0651_),
    .A1(_0648_),
    .B1(_0652_),
    .X(_0653_));
 sg13g2_a22oi_1 _3361_ (.Y(_0654_),
    .B1(_0653_),
    .B2(_0578_),
    .A2(_0647_),
    .A1(_0645_));
 sg13g2_nand3_1 _3362_ (.B(_1554_),
    .C(_0625_),
    .A(_1928_),
    .Y(_0655_));
 sg13g2_o21ai_1 _3363_ (.B1(_0655_),
    .Y(_0656_),
    .A1(_1554_),
    .A2(_0625_));
 sg13g2_a22oi_1 _3364_ (.Y(_0657_),
    .B1(_0593_),
    .B2(_0625_),
    .A2(_1553_),
    .A1(_0250_));
 sg13g2_or3_1 _3365_ (.A(_1666_),
    .B(net121),
    .C(_0625_),
    .X(_0658_));
 sg13g2_o21ai_1 _3366_ (.B1(_0658_),
    .Y(_0659_),
    .A1(_1928_),
    .A2(_0657_));
 sg13g2_a21oi_1 _3367_ (.A1(_0250_),
    .A2(_0656_),
    .Y(_0660_),
    .B1(_0659_));
 sg13g2_o21ai_1 _3368_ (.B1(_0660_),
    .Y(_0661_),
    .A1(_0642_),
    .A2(_0654_));
 sg13g2_a22oi_1 _3369_ (.Y(_0662_),
    .B1(_0640_),
    .B2(_0661_),
    .A2(_0637_),
    .A1(net120));
 sg13g2_inv_1 _3370_ (.Y(_0663_),
    .A(_0605_));
 sg13g2_a21oi_1 _3371_ (.A1(_0635_),
    .A2(_0662_),
    .Y(_0664_),
    .B1(_0663_));
 sg13g2_nor2_1 _3372_ (.A(_0635_),
    .B(_0662_),
    .Y(_0665_));
 sg13g2_nand2_1 _3373_ (.Y(_0666_),
    .A(net74),
    .B(_0612_));
 sg13g2_mux2_1 _3374_ (.A0(_0612_),
    .A1(_0666_),
    .S(_0628_),
    .X(_0667_));
 sg13g2_nand3_1 _3375_ (.B(_0612_),
    .C(_0630_),
    .A(_0255_),
    .Y(_0668_));
 sg13g2_o21ai_1 _3376_ (.B1(_0668_),
    .Y(_0669_),
    .A1(net72),
    .A2(_0667_));
 sg13g2_o21ai_1 _3377_ (.B1(_0669_),
    .Y(_0670_),
    .A1(_0664_),
    .A2(_0665_));
 sg13g2_nand3_1 _3378_ (.B(_0633_),
    .C(_0670_),
    .A(net73),
    .Y(_0671_));
 sg13g2_buf_1 _3379_ (.A(\vga.count_h[9] ),
    .X(_0672_));
 sg13g2_and2_1 _3380_ (.A(net118),
    .B(_0508_),
    .X(_0673_));
 sg13g2_buf_1 _3381_ (.A(net127),
    .X(_0674_));
 sg13g2_nand2_1 _3382_ (.Y(_0675_),
    .A(_0350_),
    .B(net138));
 sg13g2_nand2b_1 _3383_ (.Y(_0676_),
    .B(_0675_),
    .A_N(_0524_));
 sg13g2_nand2_1 _3384_ (.Y(_0677_),
    .A(net71),
    .B(_0524_));
 sg13g2_o21ai_1 _3385_ (.B1(_0677_),
    .Y(_0678_),
    .A1(net71),
    .A2(_0676_));
 sg13g2_xor2_1 _3386_ (.B(net80),
    .A(net71),
    .X(_0679_));
 sg13g2_and3_1 _3387_ (.X(_0680_),
    .A(_0674_),
    .B(_0524_),
    .C(_0675_));
 sg13g2_a221oi_1 _3388_ (.B2(net123),
    .C1(_0680_),
    .B1(_0679_),
    .A1(net122),
    .Y(_0681_),
    .A2(_0678_));
 sg13g2_nand2b_1 _3389_ (.Y(_0682_),
    .B(net124),
    .A_N(_0681_));
 sg13g2_nor3_2 _3390_ (.A(net127),
    .B(_1733_),
    .C(net80),
    .Y(_0683_));
 sg13g2_xor2_1 _3391_ (.B(net79),
    .A(net84),
    .X(_0684_));
 sg13g2_nand2_1 _3392_ (.Y(_0685_),
    .A(_0683_),
    .B(_0684_));
 sg13g2_or3_1 _3393_ (.A(net127),
    .B(_0466_),
    .C(_0467_),
    .X(_0686_));
 sg13g2_buf_1 _3394_ (.A(_0686_),
    .X(_0687_));
 sg13g2_nor2_1 _3395_ (.A(net79),
    .B(_0687_),
    .Y(_0688_));
 sg13g2_mux2_1 _3396_ (.A0(_0688_),
    .A1(_0687_),
    .S(_0462_),
    .X(_0689_));
 sg13g2_nand2_1 _3397_ (.Y(_0690_),
    .A(net82),
    .B(_0462_));
 sg13g2_o21ai_1 _3398_ (.B1(_0690_),
    .Y(_0691_),
    .A1(_0056_),
    .A2(_0687_));
 sg13g2_nor3_1 _3399_ (.A(_0473_),
    .B(_0056_),
    .C(_0683_),
    .Y(_0692_));
 sg13g2_a221oi_1 _3400_ (.B2(_0473_),
    .C1(_0692_),
    .B1(_0691_),
    .A1(net82),
    .Y(_0693_),
    .A2(_0689_));
 sg13g2_o21ai_1 _3401_ (.B1(_0693_),
    .Y(_0694_),
    .A1(_0682_),
    .A2(_0685_));
 sg13g2_nand2_1 _3402_ (.Y(_0695_),
    .A(_0352_),
    .B(_0681_));
 sg13g2_o21ai_1 _3403_ (.B1(_0466_),
    .Y(_0696_),
    .A1(_0674_),
    .A2(_0467_));
 sg13g2_nand3_1 _3404_ (.B(_0695_),
    .C(_0696_),
    .A(_0687_),
    .Y(_0697_));
 sg13g2_or2_1 _3405_ (.X(_0698_),
    .B(_0682_),
    .A(_0541_));
 sg13g2_a21oi_1 _3406_ (.A1(_0697_),
    .A2(_0698_),
    .Y(_0699_),
    .B1(_0684_));
 sg13g2_inv_2 _3407_ (.Y(_0700_),
    .A(_0344_));
 sg13g2_xnor2_1 _3408_ (.Y(_0701_),
    .A(_0462_),
    .B(_0688_));
 sg13g2_nor3_1 _3409_ (.A(net79),
    .B(net136),
    .C(_0687_),
    .Y(_0702_));
 sg13g2_xnor2_1 _3410_ (.Y(_0703_),
    .A(net137),
    .B(_0702_));
 sg13g2_xnor2_1 _3411_ (.Y(_0704_),
    .A(_0345_),
    .B(_0703_));
 sg13g2_a21oi_1 _3412_ (.A1(_0700_),
    .A2(_0701_),
    .Y(_0705_),
    .B1(_0704_));
 sg13g2_o21ai_1 _3413_ (.B1(_0705_),
    .Y(_0706_),
    .A1(_0694_),
    .A2(_0699_));
 sg13g2_buf_1 _3414_ (.A(_0048_),
    .X(_0707_));
 sg13g2_nand2_1 _3415_ (.Y(_0708_),
    .A(_1995_),
    .B(_0683_));
 sg13g2_nor2_1 _3416_ (.A(_1744_),
    .B(_0708_),
    .Y(_0709_));
 sg13g2_nand2b_1 _3417_ (.Y(_0710_),
    .B(_0709_),
    .A_N(_1745_));
 sg13g2_buf_1 _3418_ (.A(_0710_),
    .X(_0711_));
 sg13g2_or2_1 _3419_ (.X(_0712_),
    .B(_0708_),
    .A(_1744_));
 sg13g2_buf_1 _3420_ (.A(_0712_),
    .X(_0713_));
 sg13g2_nand2_1 _3421_ (.Y(_0714_),
    .A(_0707_),
    .B(_0713_));
 sg13g2_o21ai_1 _3422_ (.B1(_0714_),
    .Y(_0715_),
    .A1(_0707_),
    .A2(_0711_));
 sg13g2_nand2_1 _3423_ (.Y(_0716_),
    .A(net118),
    .B(_0707_));
 sg13g2_o21ai_1 _3424_ (.B1(_0716_),
    .Y(_0717_),
    .A1(_0054_),
    .A2(_0713_));
 sg13g2_nor3_1 _3425_ (.A(_0486_),
    .B(_0054_),
    .C(_0709_),
    .Y(_0718_));
 sg13g2_a221oi_1 _3426_ (.B2(net78),
    .C1(_0718_),
    .B1(_0717_),
    .A1(net118),
    .Y(_0719_),
    .A2(_0715_));
 sg13g2_buf_1 _3427_ (.A(_0050_),
    .X(_0720_));
 sg13g2_and2_1 _3428_ (.A(net77),
    .B(_0708_),
    .X(_0721_));
 sg13g2_nor3_1 _3429_ (.A(_0720_),
    .B(_0709_),
    .C(_0721_),
    .Y(_0722_));
 sg13g2_a21oi_1 _3430_ (.A1(_0553_),
    .A2(_0703_),
    .Y(_0723_),
    .B1(_0722_));
 sg13g2_and2_1 _3431_ (.A(_0719_),
    .B(_0723_),
    .X(_0724_));
 sg13g2_xnor2_1 _3432_ (.Y(_0725_),
    .A(net75),
    .B(_0635_));
 sg13g2_buf_1 _3433_ (.A(net146),
    .X(_0726_));
 sg13g2_xor2_1 _3434_ (.B(net70),
    .A(net89),
    .X(_0727_));
 sg13g2_xnor2_1 _3435_ (.Y(_0728_),
    .A(net91),
    .B(_0562_));
 sg13g2_nor3_1 _3436_ (.A(_0642_),
    .B(_0727_),
    .C(_0728_),
    .Y(_0729_));
 sg13g2_nand4_1 _3437_ (.B(_0653_),
    .C(_0725_),
    .A(_0660_),
    .Y(_0730_),
    .D(_0729_));
 sg13g2_nand3b_1 _3438_ (.B(_0669_),
    .C(_0640_),
    .Y(_0731_),
    .A_N(_0730_));
 sg13g2_xnor2_1 _3439_ (.Y(_0732_),
    .A(net85),
    .B(_0486_));
 sg13g2_nand3_1 _3440_ (.B(_0720_),
    .C(_0708_),
    .A(_0488_),
    .Y(_0733_));
 sg13g2_nand3_1 _3441_ (.B(_0732_),
    .C(_0733_),
    .A(_0713_),
    .Y(_0734_));
 sg13g2_or3_1 _3442_ (.A(_0720_),
    .B(_0713_),
    .C(_0732_),
    .X(_0735_));
 sg13g2_nand3_1 _3443_ (.B(_0734_),
    .C(_0735_),
    .A(_0719_),
    .Y(_0736_));
 sg13g2_xor2_1 _3444_ (.B(_0610_),
    .A(_0608_),
    .X(_0737_));
 sg13g2_nand2_1 _3445_ (.Y(_0738_),
    .A(_1603_),
    .B(_0737_));
 sg13g2_nand3_1 _3446_ (.B(net111),
    .C(_0607_),
    .A(net73),
    .Y(_0739_));
 sg13g2_o21ai_1 _3447_ (.B1(_0739_),
    .Y(_0740_),
    .A1(_0607_),
    .A2(_0738_));
 sg13g2_xor2_1 _3448_ (.B(_0711_),
    .A(_0707_),
    .X(_0741_));
 sg13g2_or3_1 _3449_ (.A(net101),
    .B(\vga.blank_h ),
    .C(\vga.blank_v ),
    .X(_0742_));
 sg13g2_inv_1 _3450_ (.Y(_0122_),
    .A(_0742_));
 sg13g2_o21ai_1 _3451_ (.B1(_0122_),
    .Y(_0743_),
    .A1(_1739_),
    .A2(_0711_));
 sg13g2_a221oi_1 _3452_ (.B2(_0342_),
    .C1(_0743_),
    .B1(_0741_),
    .A1(\vga.count_v[8] ),
    .Y(_0744_),
    .A2(_0740_));
 sg13g2_nand3_1 _3453_ (.B(_1991_),
    .C(net47),
    .A(net74),
    .Y(_0745_));
 sg13g2_a21oi_1 _3454_ (.A1(net72),
    .A2(_0745_),
    .Y(_0746_),
    .B1(_0630_));
 sg13g2_nand4_1 _3455_ (.B(_0736_),
    .C(_0744_),
    .A(_0731_),
    .Y(_0747_),
    .D(_0746_));
 sg13g2_a221oi_1 _3456_ (.B2(_0724_),
    .C1(_0747_),
    .B1(_0706_),
    .A1(_0505_),
    .Y(_0748_),
    .A2(_0673_));
 sg13g2_nand4_1 _3457_ (.B(_0621_),
    .C(_0671_),
    .A(_0559_),
    .Y(_0749_),
    .D(_0748_));
 sg13g2_inv_1 _3458_ (.Y(_0750_),
    .A(net85));
 sg13g2_inv_1 _3459_ (.Y(_0751_),
    .A(net122));
 sg13g2_nand2_1 _3460_ (.Y(_0752_),
    .A(net123),
    .B(net124));
 sg13g2_a21oi_1 _3461_ (.A1(_0350_),
    .A2(_0751_),
    .Y(_0753_),
    .B1(_0752_));
 sg13g2_nor2_1 _3462_ (.A(_0700_),
    .B(_0370_),
    .Y(_0754_));
 sg13g2_or2_1 _3463_ (.X(_0755_),
    .B(_0345_),
    .A(_0341_));
 sg13g2_buf_1 _3464_ (.A(_0755_),
    .X(_0756_));
 sg13g2_a21oi_1 _3465_ (.A1(_0753_),
    .A2(_0754_),
    .Y(_0757_),
    .B1(_0756_));
 sg13g2_o21ai_1 _3466_ (.B1(_0342_),
    .Y(_0758_),
    .A1(_0750_),
    .A2(_0757_));
 sg13g2_inv_1 _3467_ (.Y(_0759_),
    .A(_0345_));
 sg13g2_nand2_2 _3468_ (.Y(_0760_),
    .A(_0339_),
    .B(_0342_));
 sg13g2_nor3_2 _3469_ (.A(_0341_),
    .B(_0759_),
    .C(_0760_),
    .Y(_0761_));
 sg13g2_nand2_1 _3470_ (.Y(_0762_),
    .A(_0370_),
    .B(_0352_));
 sg13g2_nor4_1 _3471_ (.A(net82),
    .B(net123),
    .C(net122),
    .D(_0762_),
    .Y(_0763_));
 sg13g2_a21oi_2 _3472_ (.B1(net118),
    .Y(_0764_),
    .A2(_0756_),
    .A1(net85));
 sg13g2_a21oi_1 _3473_ (.A1(_0761_),
    .A2(_0763_),
    .Y(_0765_),
    .B1(_0764_));
 sg13g2_nor2_1 _3474_ (.A(_0593_),
    .B(_0765_),
    .Y(_0766_));
 sg13g2_nor4_1 _3475_ (.A(_0349_),
    .B(net122),
    .C(_0752_),
    .D(_0760_),
    .Y(_0767_));
 sg13g2_nor3_1 _3476_ (.A(net83),
    .B(net84),
    .C(_0346_),
    .Y(_0768_));
 sg13g2_o21ai_1 _3477_ (.B1(net82),
    .Y(_0769_),
    .A1(_0348_),
    .A2(_0753_));
 sg13g2_a21oi_1 _3478_ (.A1(_0761_),
    .A2(_0769_),
    .Y(_0770_),
    .B1(_0764_));
 sg13g2_a21oi_1 _3479_ (.A1(_0767_),
    .A2(_0768_),
    .Y(_0771_),
    .B1(_0770_));
 sg13g2_nand2_2 _3480_ (.Y(_0772_),
    .A(_0349_),
    .B(net122));
 sg13g2_nor2_1 _3481_ (.A(net123),
    .B(net124),
    .Y(_0773_));
 sg13g2_nand2_1 _3482_ (.Y(_0774_),
    .A(_0772_),
    .B(_0773_));
 sg13g2_o21ai_1 _3483_ (.B1(net82),
    .Y(_0775_),
    .A1(net84),
    .A2(_0774_));
 sg13g2_a21oi_1 _3484_ (.A1(_0761_),
    .A2(_0775_),
    .Y(_0776_),
    .B1(_0764_));
 sg13g2_nand2_1 _3485_ (.Y(_0777_),
    .A(_0354_),
    .B(_0773_));
 sg13g2_nor3_1 _3486_ (.A(_0349_),
    .B(_0760_),
    .C(_0777_),
    .Y(_0778_));
 sg13g2_and2_1 _3487_ (.A(_0778_),
    .B(_0768_),
    .X(_0779_));
 sg13g2_o21ai_1 _3488_ (.B1(\vga.score_r_unit_pixels[2] ),
    .Y(_0780_),
    .A1(_0776_),
    .A2(_0779_));
 sg13g2_and2_1 _3489_ (.A(_0771_),
    .B(_0780_),
    .X(_0781_));
 sg13g2_nor3_1 _3490_ (.A(_0349_),
    .B(_0355_),
    .C(_0760_),
    .Y(_0782_));
 sg13g2_nor4_1 _3491_ (.A(net83),
    .B(_0370_),
    .C(net124),
    .D(_0346_),
    .Y(_0783_));
 sg13g2_nor2_1 _3492_ (.A(_0350_),
    .B(_0355_),
    .Y(_0784_));
 sg13g2_o21ai_1 _3493_ (.B1(_0754_),
    .Y(_0785_),
    .A1(net124),
    .A2(_0784_));
 sg13g2_a21oi_1 _3494_ (.A1(_0761_),
    .A2(_0785_),
    .Y(_0786_),
    .B1(_0764_));
 sg13g2_a21oi_1 _3495_ (.A1(_0782_),
    .A2(_0783_),
    .Y(_0787_),
    .B1(_0786_));
 sg13g2_a21oi_1 _3496_ (.A1(\vga.score_r_unit_pixels[1] ),
    .A2(_0787_),
    .Y(_0788_),
    .B1(_0771_));
 sg13g2_inv_1 _3497_ (.Y(_0789_),
    .A(\vga.score_r_unit_pixels[0] ));
 sg13g2_nand4_1 _3498_ (.B(_0759_),
    .C(_0350_),
    .A(net83),
    .Y(_0790_),
    .D(_0763_));
 sg13g2_a21oi_1 _3499_ (.A1(_0720_),
    .A2(_0790_),
    .Y(_0791_),
    .B1(_0750_));
 sg13g2_nor4_1 _3500_ (.A(_0672_),
    .B(_0789_),
    .C(_0787_),
    .D(_0791_),
    .Y(_0792_));
 sg13g2_o21ai_1 _3501_ (.B1(_0340_),
    .Y(_0793_),
    .A1(_0756_),
    .A2(_0754_));
 sg13g2_nand3_1 _3502_ (.B(\vga.score_l_unit_pixels[0] ),
    .C(_0793_),
    .A(_0342_),
    .Y(_0794_));
 sg13g2_nor2_1 _3503_ (.A(_0341_),
    .B(_0345_),
    .Y(_0795_));
 sg13g2_nand2_1 _3504_ (.Y(_0796_),
    .A(_0700_),
    .B(_0795_));
 sg13g2_a21o_1 _3505_ (.A2(_0753_),
    .A1(_0348_),
    .B1(_0796_),
    .X(_0797_));
 sg13g2_nor2_1 _3506_ (.A(_0370_),
    .B(_0796_),
    .Y(_0798_));
 sg13g2_a221oi_1 _3507_ (.B2(_0798_),
    .C1(net118),
    .B1(_0767_),
    .A1(_0339_),
    .Y(_0799_),
    .A2(_0797_));
 sg13g2_nand2b_1 _3508_ (.Y(_0800_),
    .B(\vga.score_l_unit_pixels[1] ),
    .A_N(_0799_));
 sg13g2_nor3_1 _3509_ (.A(_0700_),
    .B(_0756_),
    .C(_0762_),
    .Y(_0801_));
 sg13g2_o21ai_1 _3510_ (.B1(_0363_),
    .Y(_0802_),
    .A1(_0784_),
    .A2(_0762_));
 sg13g2_nand2_1 _3511_ (.Y(_0803_),
    .A(_0795_),
    .B(_0802_));
 sg13g2_a221oi_1 _3512_ (.B2(net85),
    .C1(net118),
    .B1(_0803_),
    .A1(_0782_),
    .Y(_0804_),
    .A2(_0801_));
 sg13g2_mux2_1 _3513_ (.A0(_0794_),
    .A1(_0800_),
    .S(_0804_),
    .X(_0805_));
 sg13g2_a21oi_1 _3514_ (.A1(_0772_),
    .A2(_0773_),
    .Y(_0806_),
    .B1(_0370_));
 sg13g2_nor2b_1 _3515_ (.A(net82),
    .B_N(\vga.score_r_ten_enable ),
    .Y(_0807_));
 sg13g2_nand2_1 _3516_ (.Y(_0808_),
    .A(_0349_),
    .B(_0751_));
 sg13g2_a21oi_1 _3517_ (.A1(_0051_),
    .A2(_0808_),
    .Y(_0809_),
    .B1(_0352_));
 sg13g2_o21ai_1 _3518_ (.B1(net123),
    .Y(_0810_),
    .A1(_0764_),
    .A2(_0809_));
 sg13g2_nand4_1 _3519_ (.B(_0806_),
    .C(_0807_),
    .A(_0761_),
    .Y(_0811_),
    .D(_0810_));
 sg13g2_a22oi_1 _3520_ (.Y(_0812_),
    .B1(_0809_),
    .B2(_0353_),
    .A2(_0773_),
    .A1(_0772_));
 sg13g2_nor3_1 _3521_ (.A(_0672_),
    .B(net84),
    .C(_0796_),
    .Y(_0813_));
 sg13g2_nand4_1 _3522_ (.B(\vga.score_l_ten_enable ),
    .C(_0812_),
    .A(net85),
    .Y(_0814_),
    .D(_0813_));
 sg13g2_o21ai_1 _3523_ (.B1(_0340_),
    .Y(_0815_),
    .A1(_0796_),
    .A2(_0806_));
 sg13g2_a21oi_1 _3524_ (.A1(_0798_),
    .A2(_0778_),
    .Y(_0816_),
    .B1(net118));
 sg13g2_nand2_1 _3525_ (.Y(_0817_),
    .A(_0815_),
    .B(_0816_));
 sg13g2_nand3_1 _3526_ (.B(_0799_),
    .C(_0817_),
    .A(\vga.score_l_unit_pixels[2] ),
    .Y(_0818_));
 sg13g2_nand4_1 _3527_ (.B(_0811_),
    .C(_0814_),
    .A(_0805_),
    .Y(_0819_),
    .D(_0818_));
 sg13g2_nor2_1 _3528_ (.A(_0792_),
    .B(_0819_),
    .Y(_0820_));
 sg13g2_o21ai_1 _3529_ (.B1(_0820_),
    .Y(_0821_),
    .A1(_0781_),
    .A2(_0788_));
 sg13g2_nand2_1 _3530_ (.Y(_0822_),
    .A(_0245_),
    .B(net89));
 sg13g2_nor2_1 _3531_ (.A(net90),
    .B(net59),
    .Y(_0823_));
 sg13g2_inv_1 _3532_ (.Y(_0824_),
    .A(_0252_));
 sg13g2_a21oi_1 _3533_ (.A1(_0822_),
    .A2(_0823_),
    .Y(_0825_),
    .B1(_0824_));
 sg13g2_nor3_1 _3534_ (.A(net87),
    .B(net120),
    .C(_0825_),
    .Y(_0826_));
 sg13g2_nand2b_1 _3535_ (.Y(_0827_),
    .B(net89),
    .A_N(net91));
 sg13g2_a21oi_1 _3536_ (.A1(_0080_),
    .A2(_0827_),
    .Y(_0828_),
    .B1(_0278_));
 sg13g2_nor4_1 _3537_ (.A(net59),
    .B(net87),
    .C(_0252_),
    .D(_0828_),
    .Y(_0829_));
 sg13g2_nor2b_1 _3538_ (.A(_0829_),
    .B_N(net120),
    .Y(_0830_));
 sg13g2_nor4_1 _3539_ (.A(_0623_),
    .B(_0258_),
    .C(_0826_),
    .D(_0830_),
    .Y(_0831_));
 sg13g2_a22oi_1 _3540_ (.Y(_0832_),
    .B1(_0821_),
    .B2(_0831_),
    .A2(_0766_),
    .A1(_0758_));
 sg13g2_nor2_2 _3541_ (.A(net107),
    .B(net108),
    .Y(_0833_));
 sg13g2_nand2b_1 _3542_ (.Y(_0834_),
    .B(_0833_),
    .A_N(_1621_));
 sg13g2_nor4_1 _3543_ (.A(_1584_),
    .B(net110),
    .C(_1638_),
    .D(_0834_),
    .Y(_0835_));
 sg13g2_nor2_1 _3544_ (.A(_1638_),
    .B(_0834_),
    .Y(_0836_));
 sg13g2_and2_1 _3545_ (.A(_1685_),
    .B(_0836_),
    .X(_0837_));
 sg13g2_nor2_1 _3546_ (.A(_1685_),
    .B(_0836_),
    .Y(_0838_));
 sg13g2_buf_1 _3547_ (.A(net114),
    .X(_0839_));
 sg13g2_nor2_1 _3548_ (.A(_1650_),
    .B(_0833_),
    .Y(_0840_));
 sg13g2_o21ai_1 _3549_ (.B1(net64),
    .Y(_0841_),
    .A1(net55),
    .A2(_0840_));
 sg13g2_xnor2_1 _3550_ (.Y(_0842_),
    .A(_1559_),
    .B(_0841_));
 sg13g2_nand2_1 _3551_ (.Y(_0843_),
    .A(net120),
    .B(_0842_));
 sg13g2_o21ai_1 _3552_ (.B1(_0843_),
    .Y(_0844_),
    .A1(_0837_),
    .A2(_0838_));
 sg13g2_xnor2_1 _3553_ (.Y(_0845_),
    .A(_1635_),
    .B(_1692_));
 sg13g2_a21oi_1 _3554_ (.A1(_1685_),
    .A2(_0845_),
    .Y(_0846_),
    .B1(_0611_));
 sg13g2_nor2_1 _3555_ (.A(_0838_),
    .B(_0843_),
    .Y(_0847_));
 sg13g2_a22oi_1 _3556_ (.Y(_0848_),
    .B1(_0846_),
    .B2(_0847_),
    .A2(_0844_),
    .A1(net75));
 sg13g2_nand2b_1 _3557_ (.Y(_0849_),
    .B(_0848_),
    .A_N(_0835_));
 sg13g2_xnor2_1 _3558_ (.Y(_0850_),
    .A(net66),
    .B(_0566_));
 sg13g2_nor4_1 _3559_ (.A(_0567_),
    .B(net107),
    .C(net108),
    .D(_0850_),
    .Y(_0851_));
 sg13g2_a21o_1 _3560_ (.A2(_0850_),
    .A1(net107),
    .B1(_0851_),
    .X(_0852_));
 sg13g2_nor2_1 _3561_ (.A(_1517_),
    .B(_0833_),
    .Y(_0853_));
 sg13g2_xnor2_1 _3562_ (.Y(_0854_),
    .A(net115),
    .B(_0853_));
 sg13g2_nor2_1 _3563_ (.A(_0567_),
    .B(net108),
    .Y(_0855_));
 sg13g2_mux2_1 _3564_ (.A0(net108),
    .A1(_0855_),
    .S(net107),
    .X(_0856_));
 sg13g2_xnor2_1 _3565_ (.Y(_0857_),
    .A(net66),
    .B(_0833_));
 sg13g2_nor2_1 _3566_ (.A(net86),
    .B(_0857_),
    .Y(_0858_));
 sg13g2_a21o_1 _3567_ (.A2(_0856_),
    .A1(_0850_),
    .B1(_0858_),
    .X(_0859_));
 sg13g2_a221oi_1 _3568_ (.B2(_0271_),
    .C1(_0859_),
    .B1(_0854_),
    .A1(_0245_),
    .Y(_0860_),
    .A2(_0852_));
 sg13g2_nor2_1 _3569_ (.A(net59),
    .B(_0854_),
    .Y(_0861_));
 sg13g2_xnor2_1 _3570_ (.Y(_0862_),
    .A(net55),
    .B(_0840_));
 sg13g2_nor3_1 _3571_ (.A(_0860_),
    .B(_0861_),
    .C(_0862_),
    .Y(_0863_));
 sg13g2_o21ai_1 _3572_ (.B1(_0862_),
    .Y(_0864_),
    .A1(_0860_),
    .A2(_0861_));
 sg13g2_o21ai_1 _3573_ (.B1(_0864_),
    .Y(_0865_),
    .A1(_0252_),
    .A2(_0863_));
 sg13g2_nand2_1 _3574_ (.Y(_0866_),
    .A(_1668_),
    .B(_0834_));
 sg13g2_xnor2_1 _3575_ (.Y(_0867_),
    .A(net64),
    .B(_0866_));
 sg13g2_o21ai_1 _3576_ (.B1(_0279_),
    .Y(_0868_),
    .A1(_0865_),
    .A2(_0867_));
 sg13g2_nand2b_1 _3577_ (.Y(_0869_),
    .B(_0845_),
    .A_N(_0837_));
 sg13g2_nand2_1 _3578_ (.Y(_0870_),
    .A(_0663_),
    .B(_0845_));
 sg13g2_o21ai_1 _3579_ (.B1(_0870_),
    .Y(_0871_),
    .A1(_0622_),
    .A2(_0835_));
 sg13g2_nor2_1 _3580_ (.A(_0622_),
    .B(_0845_),
    .Y(_0872_));
 sg13g2_nor2_1 _3581_ (.A(_0838_),
    .B(_0872_),
    .Y(_0873_));
 sg13g2_xnor2_1 _3582_ (.Y(_0874_),
    .A(_0560_),
    .B(_0842_));
 sg13g2_o21ai_1 _3583_ (.B1(_0874_),
    .Y(_0875_),
    .A1(net75),
    .A2(_0873_));
 sg13g2_a221oi_1 _3584_ (.B2(_0867_),
    .C1(_0875_),
    .B1(_0865_),
    .A1(_0869_),
    .Y(_0876_),
    .A2(_0871_));
 sg13g2_nand2_1 _3585_ (.Y(_0877_),
    .A(_0838_),
    .B(_0843_));
 sg13g2_o21ai_1 _3586_ (.B1(_0877_),
    .Y(_0878_),
    .A1(_0605_),
    .A2(_0847_));
 sg13g2_a21oi_1 _3587_ (.A1(_0611_),
    .A2(_0878_),
    .Y(_0879_),
    .B1(_0869_));
 sg13g2_a221oi_1 _3588_ (.B2(_0876_),
    .C1(_0879_),
    .B1(_0868_),
    .A1(_0622_),
    .Y(_0880_),
    .A2(_0849_));
 sg13g2_xnor2_1 _3589_ (.Y(_0881_),
    .A(_0255_),
    .B(_1606_));
 sg13g2_nor2_1 _3590_ (.A(_0609_),
    .B(_0881_),
    .Y(_0882_));
 sg13g2_o21ai_1 _3591_ (.B1(_0882_),
    .Y(_0883_),
    .A1(_0622_),
    .A2(_1588_));
 sg13g2_inv_1 _3592_ (.Y(_0884_),
    .A(_0836_));
 sg13g2_nand4_1 _3593_ (.B(_1668_),
    .C(_1628_),
    .A(net110),
    .Y(_0885_),
    .D(_0884_));
 sg13g2_mux2_1 _3594_ (.A0(_0883_),
    .A1(_0617_),
    .S(_0885_),
    .X(_0886_));
 sg13g2_inv_1 _3595_ (.Y(_0887_),
    .A(_0886_));
 sg13g2_a21oi_1 _3596_ (.A1(_0567_),
    .A2(net108),
    .Y(_0888_),
    .B1(net107));
 sg13g2_nand3_1 _3597_ (.B(net107),
    .C(net108),
    .A(_0567_),
    .Y(_0889_));
 sg13g2_o21ai_1 _3598_ (.B1(_0889_),
    .Y(_0890_),
    .A1(_0245_),
    .A2(_0888_));
 sg13g2_buf_2 _3599_ (.A(_0890_),
    .X(_0891_));
 sg13g2_o21ai_1 _3600_ (.B1(net86),
    .Y(_0892_),
    .A1(_1517_),
    .A2(_0891_));
 sg13g2_nand2_1 _3601_ (.Y(_0893_),
    .A(_1517_),
    .B(_0891_));
 sg13g2_a21oi_1 _3602_ (.A1(_0892_),
    .A2(_0893_),
    .Y(_0894_),
    .B1(net59));
 sg13g2_nand2_1 _3603_ (.Y(_0895_),
    .A(net86),
    .B(_0891_));
 sg13g2_a21oi_1 _3604_ (.A1(net59),
    .A2(_0895_),
    .Y(_0896_),
    .B1(_1650_));
 sg13g2_o21ai_1 _3605_ (.B1(net121),
    .Y(_0897_),
    .A1(_0894_),
    .A2(_0896_));
 sg13g2_or2_1 _3606_ (.X(_0898_),
    .B(net65),
    .A(_1687_));
 sg13g2_a21oi_1 _3607_ (.A1(_1563_),
    .A2(_0897_),
    .Y(_0899_),
    .B1(_0898_));
 sg13g2_and2_1 _3608_ (.A(_1687_),
    .B(net65),
    .X(_0900_));
 sg13g2_and2_1 _3609_ (.A(_1570_),
    .B(_1571_),
    .X(_0901_));
 sg13g2_nand2_1 _3610_ (.Y(_0902_),
    .A(_0256_),
    .B(_0901_));
 sg13g2_or2_1 _3611_ (.X(_0903_),
    .B(_0901_),
    .A(_0256_));
 sg13g2_nand3_1 _3612_ (.B(net147),
    .C(_0561_),
    .A(_1576_),
    .Y(_0904_));
 sg13g2_o21ai_1 _3613_ (.B1(_0904_),
    .Y(_0905_),
    .A1(net147),
    .A2(_0561_));
 sg13g2_nor3_1 _3614_ (.A(net112),
    .B(net147),
    .C(_0560_),
    .Y(_0906_));
 sg13g2_a21oi_1 _3615_ (.A1(net147),
    .A2(_0560_),
    .Y(_0907_),
    .B1(_0906_));
 sg13g2_nor2_1 _3616_ (.A(_1578_),
    .B(_0907_),
    .Y(_0908_));
 sg13g2_a221oi_1 _3617_ (.B2(_1578_),
    .C1(_0908_),
    .B1(_0905_),
    .A1(_0902_),
    .Y(_0909_),
    .A2(_0903_));
 sg13g2_inv_1 _3618_ (.Y(_0910_),
    .A(_0909_));
 sg13g2_or4_1 _3619_ (.A(_0584_),
    .B(_0899_),
    .C(_0900_),
    .D(_0910_),
    .X(_0911_));
 sg13g2_o21ai_1 _3620_ (.B1(net115),
    .Y(_0912_),
    .A1(net66),
    .A2(_0891_));
 sg13g2_a21oi_1 _3621_ (.A1(net66),
    .A2(_0891_),
    .Y(_0913_),
    .B1(net115));
 sg13g2_a21o_1 _3622_ (.A2(_0912_),
    .A1(net90),
    .B1(_0913_),
    .X(_0914_));
 sg13g2_o21ai_1 _3623_ (.B1(_0592_),
    .Y(_0915_),
    .A1(_1561_),
    .A2(_0891_));
 sg13g2_a21oi_1 _3624_ (.A1(_1540_),
    .A2(_0891_),
    .Y(_0916_),
    .B1(net121));
 sg13g2_a21o_1 _3625_ (.A2(_0915_),
    .A1(net90),
    .B1(_0916_),
    .X(_0917_));
 sg13g2_a221oi_1 _3626_ (.B2(net59),
    .C1(net55),
    .B1(_0917_),
    .A1(_0593_),
    .Y(_0918_),
    .A2(_0914_));
 sg13g2_or3_1 _3627_ (.A(_0592_),
    .B(_0263_),
    .C(_0891_),
    .X(_0919_));
 sg13g2_nand3_1 _3628_ (.B(_1541_),
    .C(_0919_),
    .A(net55),
    .Y(_0920_));
 sg13g2_nor2b_1 _3629_ (.A(_0918_),
    .B_N(_0920_),
    .Y(_0921_));
 sg13g2_inv_1 _3630_ (.Y(_0922_),
    .A(_0584_));
 sg13g2_nand4_1 _3631_ (.B(net55),
    .C(_0922_),
    .A(net64),
    .Y(_0923_),
    .D(_1561_));
 sg13g2_nand2_1 _3632_ (.Y(_0924_),
    .A(_0584_),
    .B(net65));
 sg13g2_xnor2_1 _3633_ (.Y(_0925_),
    .A(_1535_),
    .B(_0924_));
 sg13g2_and4_1 _3634_ (.A(_0897_),
    .B(_0909_),
    .C(_0923_),
    .D(_0925_),
    .X(_0926_));
 sg13g2_nand2_1 _3635_ (.Y(_0927_),
    .A(_0622_),
    .B(_1588_));
 sg13g2_inv_1 _3636_ (.Y(_0928_),
    .A(_0043_));
 sg13g2_a21oi_1 _3637_ (.A1(_0928_),
    .A2(_1590_),
    .Y(_0929_),
    .B1(_0609_));
 sg13g2_nor3_1 _3638_ (.A(_0560_),
    .B(_1579_),
    .C(_1565_),
    .Y(_0930_));
 sg13g2_nand2_1 _3639_ (.Y(_0931_),
    .A(_0909_),
    .B(_0930_));
 sg13g2_nand3_1 _3640_ (.B(_0929_),
    .C(_0931_),
    .A(_0927_),
    .Y(_0932_));
 sg13g2_a21oi_1 _3641_ (.A1(_0921_),
    .A2(_0926_),
    .Y(_0933_),
    .B1(_0932_));
 sg13g2_and4_1 _3642_ (.A(_0720_),
    .B(_0365_),
    .C(_0355_),
    .D(_0783_),
    .X(_0934_));
 sg13g2_nand2_1 _3643_ (.Y(_0935_),
    .A(net72),
    .B(_0885_));
 sg13g2_nand3_1 _3644_ (.B(_0934_),
    .C(_0935_),
    .A(_1606_),
    .Y(_0936_));
 sg13g2_a221oi_1 _3645_ (.B2(_0933_),
    .C1(_0936_),
    .B1(_0911_),
    .A1(_0617_),
    .Y(_0937_),
    .A2(_0883_));
 sg13g2_o21ai_1 _3646_ (.B1(_0937_),
    .Y(_0938_),
    .A1(_0880_),
    .A2(_0887_));
 sg13g2_a21o_1 _3647_ (.A2(_0938_),
    .A1(_0832_),
    .B1(_0742_),
    .X(_0939_));
 sg13g2_nor2_1 _3648_ (.A(_1943_),
    .B(_1947_),
    .Y(_0940_));
 sg13g2_or2_1 _3649_ (.X(_0941_),
    .B(net131),
    .A(_1850_));
 sg13g2_buf_1 _3650_ (.A(_0941_),
    .X(_0942_));
 sg13g2_nor3_1 _3651_ (.A(_1917_),
    .B(_1946_),
    .C(_0942_),
    .Y(_0943_));
 sg13g2_nand2_1 _3652_ (.Y(_0944_),
    .A(_0622_),
    .B(_0943_));
 sg13g2_xnor2_1 _3653_ (.Y(_0945_),
    .A(_1865_),
    .B(_1890_));
 sg13g2_nand2_1 _3654_ (.Y(_0946_),
    .A(net119),
    .B(_0945_));
 sg13g2_o21ai_1 _3655_ (.B1(_0946_),
    .Y(_0947_),
    .A1(_0940_),
    .A2(_0944_));
 sg13g2_nand2_1 _3656_ (.Y(_0948_),
    .A(_1914_),
    .B(_1917_));
 sg13g2_o21ai_1 _3657_ (.B1(_0948_),
    .Y(_0949_),
    .A1(_1917_),
    .A2(_0942_));
 sg13g2_buf_1 _3658_ (.A(_0949_),
    .X(_0950_));
 sg13g2_or3_1 _3659_ (.A(_1942_),
    .B(_1946_),
    .C(_0950_),
    .X(_0951_));
 sg13g2_buf_1 _3660_ (.A(_0951_),
    .X(_0952_));
 sg13g2_xor2_1 _3661_ (.B(_0566_),
    .A(net61),
    .X(_0953_));
 sg13g2_nor2_2 _3662_ (.A(net130),
    .B(net131),
    .Y(_0954_));
 sg13g2_nand3_1 _3663_ (.B(_0954_),
    .C(_0953_),
    .A(net89),
    .Y(_0955_));
 sg13g2_o21ai_1 _3664_ (.B1(_0955_),
    .Y(_0956_),
    .A1(_1837_),
    .A2(_0953_));
 sg13g2_nor2_1 _3665_ (.A(_1975_),
    .B(_0954_),
    .Y(_0957_));
 sg13g2_a21oi_1 _3666_ (.A1(net61),
    .A2(_0942_),
    .Y(_0958_),
    .B1(net97));
 sg13g2_or2_1 _3667_ (.X(_0959_),
    .B(_0958_),
    .A(_0957_));
 sg13g2_xnor2_1 _3668_ (.Y(_0960_),
    .A(net61),
    .B(_0954_));
 sg13g2_nand3b_1 _3669_ (.B(net130),
    .C(net89),
    .Y(_0961_),
    .A_N(net131));
 sg13g2_nand2b_1 _3670_ (.Y(_0962_),
    .B(net131),
    .A_N(net130));
 sg13g2_a21o_1 _3671_ (.A2(_0962_),
    .A1(_0961_),
    .B1(_0953_),
    .X(_0963_));
 sg13g2_o21ai_1 _3672_ (.B1(_0963_),
    .Y(_0964_),
    .A1(net86),
    .A2(_0960_));
 sg13g2_a221oi_1 _3673_ (.B2(_0271_),
    .C1(_0964_),
    .B1(_0959_),
    .A1(net91),
    .Y(_0965_),
    .A2(_0956_));
 sg13g2_nor2_1 _3674_ (.A(_0272_),
    .B(_0959_),
    .Y(_0966_));
 sg13g2_nor2_1 _3675_ (.A(_0965_),
    .B(_0966_),
    .Y(_0967_));
 sg13g2_buf_1 _3676_ (.A(net99),
    .X(_0968_));
 sg13g2_xor2_1 _3677_ (.B(_0957_),
    .A(net54),
    .X(_0969_));
 sg13g2_a21oi_1 _3678_ (.A1(_0593_),
    .A2(_0967_),
    .Y(_0970_),
    .B1(_0969_));
 sg13g2_xnor2_1 _3679_ (.Y(_0971_),
    .A(_1858_),
    .B(_0950_));
 sg13g2_xnor2_1 _3680_ (.Y(_0972_),
    .A(_0584_),
    .B(_0971_));
 sg13g2_o21ai_1 _3681_ (.B1(_0972_),
    .Y(_0973_),
    .A1(_0593_),
    .A2(_0967_));
 sg13g2_nand2_1 _3682_ (.Y(_0974_),
    .A(net87),
    .B(_0971_));
 sg13g2_o21ai_1 _3683_ (.B1(_0974_),
    .Y(_0975_),
    .A1(_0970_),
    .A2(_0973_));
 sg13g2_o21ai_1 _3684_ (.B1(net63),
    .Y(_0976_),
    .A1(net99),
    .A2(_0957_));
 sg13g2_xor2_1 _3685_ (.B(_0976_),
    .A(net60),
    .X(_0977_));
 sg13g2_xnor2_1 _3686_ (.Y(_0978_),
    .A(_0560_),
    .B(_0977_));
 sg13g2_nand2_1 _3687_ (.Y(_0979_),
    .A(_0975_),
    .B(_0978_));
 sg13g2_nor2_1 _3688_ (.A(_1966_),
    .B(_0950_),
    .Y(_0980_));
 sg13g2_xnor2_1 _3689_ (.Y(_0981_),
    .A(net96),
    .B(_0980_));
 sg13g2_nand2b_1 _3690_ (.Y(_0982_),
    .B(_0940_),
    .A_N(_0943_));
 sg13g2_nor2_1 _3691_ (.A(net119),
    .B(_0982_),
    .Y(_0983_));
 sg13g2_a221oi_1 _3692_ (.B2(net120),
    .C1(_0983_),
    .B1(_0977_),
    .A1(net75),
    .Y(_0984_),
    .A2(_0981_));
 sg13g2_o21ai_1 _3693_ (.B1(_1969_),
    .Y(_0985_),
    .A1(_1970_),
    .A2(_0950_));
 sg13g2_nand2_1 _3694_ (.Y(_0986_),
    .A(net75),
    .B(_0943_));
 sg13g2_o21ai_1 _3695_ (.B1(_0986_),
    .Y(_0987_),
    .A1(net119),
    .A2(_0985_));
 sg13g2_nand2b_1 _3696_ (.Y(_0988_),
    .B(_0987_),
    .A_N(_0940_));
 sg13g2_a21oi_1 _3697_ (.A1(net119),
    .A2(_0985_),
    .Y(_0989_),
    .B1(_0982_));
 sg13g2_a21oi_1 _3698_ (.A1(net119),
    .A2(_0982_),
    .Y(_0990_),
    .B1(_0663_));
 sg13g2_nor2_1 _3699_ (.A(_0989_),
    .B(_0990_),
    .Y(_0991_));
 sg13g2_a22oi_1 _3700_ (.Y(_0992_),
    .B1(_0988_),
    .B2(_0991_),
    .A2(_0984_),
    .A1(_0979_));
 sg13g2_a221oi_1 _3701_ (.B2(_0992_),
    .C1(net72),
    .B1(_0952_),
    .A1(net73),
    .Y(_0993_),
    .A2(_0947_));
 sg13g2_nor2_1 _3702_ (.A(_1877_),
    .B(_1879_),
    .Y(_0994_));
 sg13g2_xnor2_1 _3703_ (.Y(_0995_),
    .A(_0663_),
    .B(_0994_));
 sg13g2_nor2_1 _3704_ (.A(_0560_),
    .B(_0995_),
    .Y(_0996_));
 sg13g2_a21oi_1 _3705_ (.A1(_0928_),
    .A2(_1899_),
    .Y(_0997_),
    .B1(_0609_));
 sg13g2_o21ai_1 _3706_ (.B1(_0997_),
    .Y(_0998_),
    .A1(net119),
    .A2(_0945_));
 sg13g2_a21oi_1 _3707_ (.A1(_1896_),
    .A2(_0996_),
    .Y(_0999_),
    .B1(_0998_));
 sg13g2_nor2_1 _3708_ (.A(net63),
    .B(net62),
    .Y(_1000_));
 sg13g2_a21oi_1 _3709_ (.A1(_0567_),
    .A2(net131),
    .Y(_1001_),
    .B1(net130));
 sg13g2_nand2_1 _3710_ (.Y(_1002_),
    .A(net130),
    .B(net131));
 sg13g2_o21ai_1 _3711_ (.B1(_0245_),
    .Y(_1003_),
    .A1(net89),
    .A2(_1002_));
 sg13g2_nand2b_1 _3712_ (.Y(_1004_),
    .B(_1003_),
    .A_N(_1001_));
 sg13g2_a21oi_1 _3713_ (.A1(_1831_),
    .A2(_1004_),
    .Y(_1005_),
    .B1(net88));
 sg13g2_o21ai_1 _3714_ (.B1(net88),
    .Y(_1006_),
    .A1(_1831_),
    .A2(_1004_));
 sg13g2_o21ai_1 _3715_ (.B1(_1006_),
    .Y(_1007_),
    .A1(net86),
    .A2(_1005_));
 sg13g2_a21oi_1 _3716_ (.A1(net88),
    .A2(_1004_),
    .Y(_1008_),
    .B1(_1847_));
 sg13g2_o21ai_1 _3717_ (.B1(_1847_),
    .Y(_1009_),
    .A1(net88),
    .A2(_1004_));
 sg13g2_o21ai_1 _3718_ (.B1(_1009_),
    .Y(_1010_),
    .A1(net86),
    .A2(_1008_));
 sg13g2_a21oi_2 _3719_ (.B1(_1010_),
    .Y(_1011_),
    .A2(_1007_),
    .A1(_1842_));
 sg13g2_nor4_1 _3720_ (.A(net63),
    .B(_1864_),
    .C(net121),
    .D(_1011_),
    .Y(_1012_));
 sg13g2_nand3b_1 _3721_ (.B(_1819_),
    .C(_1825_),
    .Y(_1013_),
    .A_N(net54));
 sg13g2_nand2_1 _3722_ (.Y(_1014_),
    .A(net63),
    .B(_1864_));
 sg13g2_a22oi_1 _3723_ (.Y(_1015_),
    .B1(_1011_),
    .B2(net121),
    .A2(_1014_),
    .A1(_1013_));
 sg13g2_inv_1 _3724_ (.Y(_1016_),
    .A(net62));
 sg13g2_o21ai_1 _3725_ (.B1(_0922_),
    .Y(_1017_),
    .A1(_1858_),
    .A2(_1016_));
 sg13g2_nor4_1 _3726_ (.A(_1000_),
    .B(_1012_),
    .C(_1015_),
    .D(_1017_),
    .Y(_1018_));
 sg13g2_nand3b_1 _3727_ (.B(_1819_),
    .C(net54),
    .Y(_1019_),
    .A_N(_1825_));
 sg13g2_nand3b_1 _3728_ (.B(_1864_),
    .C(_1825_),
    .Y(_1020_),
    .A_N(net54));
 sg13g2_a22oi_1 _3729_ (.Y(_1021_),
    .B1(_1019_),
    .B2(_1020_),
    .A2(_1011_),
    .A1(net121));
 sg13g2_nor4_1 _3730_ (.A(_1819_),
    .B(net121),
    .C(_1016_),
    .D(_1011_),
    .Y(_1022_));
 sg13g2_nor3_1 _3731_ (.A(_0922_),
    .B(_1021_),
    .C(_1022_),
    .Y(_1023_));
 sg13g2_nor2_1 _3732_ (.A(_0561_),
    .B(_1883_),
    .Y(_1024_));
 sg13g2_a21oi_1 _3733_ (.A1(net60),
    .A2(_0561_),
    .Y(_1025_),
    .B1(_1024_));
 sg13g2_xor2_1 _3734_ (.B(_1025_),
    .A(_1884_),
    .X(_1026_));
 sg13g2_or4_1 _3735_ (.A(_0995_),
    .B(_1018_),
    .C(_1023_),
    .D(_1026_),
    .X(_1027_));
 sg13g2_nor2_1 _3736_ (.A(net73),
    .B(_0952_),
    .Y(_1028_));
 sg13g2_and4_1 _3737_ (.A(_0750_),
    .B(_0351_),
    .C(_0355_),
    .D(_0122_),
    .X(_1029_));
 sg13g2_a21oi_1 _3738_ (.A1(net73),
    .A2(_0947_),
    .Y(_1030_),
    .B1(net72));
 sg13g2_nand2b_1 _3739_ (.Y(_1031_),
    .B(_0952_),
    .A_N(_1030_));
 sg13g2_nand4_1 _3740_ (.B(_0813_),
    .C(_1029_),
    .A(_1893_),
    .Y(_1032_),
    .D(_1031_));
 sg13g2_a221oi_1 _3741_ (.B2(_0992_),
    .C1(_1032_),
    .B1(_1028_),
    .A1(_0999_),
    .Y(_1033_),
    .A2(_1027_));
 sg13g2_o21ai_1 _3742_ (.B1(_1033_),
    .Y(_1034_),
    .A1(_0609_),
    .A2(_0993_));
 sg13g2_nand3_1 _3743_ (.B(_0939_),
    .C(_1034_),
    .A(_0749_),
    .Y(_0191_));
 sg13g2_and3_1 _3744_ (.X(_0193_),
    .A(\vga.right_down_1d ),
    .B(net4),
    .C(_0319_));
 sg13g2_and3_1 _3745_ (.X(_0195_),
    .A(\vga.right_up_1d ),
    .B(net3),
    .C(_0319_));
 sg13g2_buf_1 _3746_ (.A(\vga.ball_angle[0] ),
    .X(_1035_));
 sg13g2_nor2_1 _3747_ (.A(_1737_),
    .B(_1747_),
    .Y(_1036_));
 sg13g2_buf_1 _3748_ (.A(_1036_),
    .X(_1037_));
 sg13g2_nor2b_1 _3749_ (.A(_2061_),
    .B_N(_1775_),
    .Y(_1038_));
 sg13g2_or2_1 _3750_ (.X(_1039_),
    .B(_1697_),
    .A(_1600_));
 sg13g2_mux2_1 _3751_ (.A0(_0064_),
    .A1(_1038_),
    .S(_1039_),
    .X(_1040_));
 sg13g2_nor2b_1 _3752_ (.A(_0064_),
    .B_N(_2037_),
    .Y(_1041_));
 sg13g2_mux2_1 _3753_ (.A0(_1041_),
    .A1(_2061_),
    .S(_2060_),
    .X(_1042_));
 sg13g2_a221oi_1 _3754_ (.B2(_2062_),
    .C1(_2035_),
    .B1(_1042_),
    .A1(net49),
    .Y(_1043_),
    .A2(_1040_));
 sg13g2_buf_2 _3755_ (.A(_1043_),
    .X(_1044_));
 sg13g2_nor2_2 _3756_ (.A(net94),
    .B(net49),
    .Y(_1045_));
 sg13g2_or3_1 _3757_ (.A(_1735_),
    .B(_1997_),
    .C(_1999_),
    .X(_1046_));
 sg13g2_buf_1 _3758_ (.A(_1046_),
    .X(_1047_));
 sg13g2_and2_1 _3759_ (.A(net94),
    .B(_1047_),
    .X(_1048_));
 sg13g2_buf_1 _3760_ (.A(_1048_),
    .X(_1049_));
 sg13g2_nor2_2 _3761_ (.A(_1045_),
    .B(_1049_),
    .Y(_1050_));
 sg13g2_and2_1 _3762_ (.A(_1044_),
    .B(_1050_),
    .X(_1051_));
 sg13g2_mux2_1 _3763_ (.A0(_1035_),
    .A1(_0084_),
    .S(_1051_),
    .X(_1052_));
 sg13g2_buf_1 _3764_ (.A(net134),
    .X(_1053_));
 sg13g2_nand2b_1 _3765_ (.Y(_0093_),
    .B(net69),
    .A_N(_1052_));
 sg13g2_buf_1 _3766_ (.A(net58),
    .X(_1054_));
 sg13g2_buf_1 _3767_ (.A(\vga.ball_angle[1] ),
    .X(_1055_));
 sg13g2_buf_8 _3768_ (.A(_1044_),
    .X(_1056_));
 sg13g2_buf_1 _3769_ (.A(_1050_),
    .X(_1057_));
 sg13g2_nand3b_1 _3770_ (.B(net32),
    .C(_1057_),
    .Y(_1058_),
    .A_N(_1035_));
 sg13g2_xor2_1 _3771_ (.B(_1058_),
    .A(_1055_),
    .X(_1059_));
 sg13g2_nor2_1 _3772_ (.A(net52),
    .B(_1059_),
    .Y(_0094_));
 sg13g2_nor2_1 _3773_ (.A(_1055_),
    .B(_1035_),
    .Y(_1060_));
 sg13g2_xor2_1 _3774_ (.B(_1060_),
    .A(_0063_),
    .X(_1061_));
 sg13g2_mux2_1 _3775_ (.A0(\vga.ball_angle[2] ),
    .A1(_1061_),
    .S(_1051_),
    .X(_1062_));
 sg13g2_and2_1 _3776_ (.A(_2076_),
    .B(_1062_),
    .X(_0095_));
 sg13g2_buf_1 _3777_ (.A(\vga.ball_angle[3] ),
    .X(_1063_));
 sg13g2_buf_1 _3778_ (.A(\vga.ball_ratio[0] ),
    .X(_1064_));
 sg13g2_xor2_1 _3779_ (.B(_1064_),
    .A(_1035_),
    .X(_1065_));
 sg13g2_buf_1 _3780_ (.A(\vga.ball_ratio[2] ),
    .X(_1066_));
 sg13g2_xor2_1 _3781_ (.B(\vga.ball_angle[2] ),
    .A(_1066_),
    .X(_1067_));
 sg13g2_xor2_1 _3782_ (.B(\vga.ball_ratio[1] ),
    .A(_1055_),
    .X(_1068_));
 sg13g2_nor3_2 _3783_ (.A(_1065_),
    .B(_1067_),
    .C(_1068_),
    .Y(_1069_));
 sg13g2_nand2_1 _3784_ (.Y(_1070_),
    .A(_0063_),
    .B(_1060_));
 sg13g2_and2_1 _3785_ (.A(_1069_),
    .B(_1070_),
    .X(_1071_));
 sg13g2_buf_1 _3786_ (.A(_1071_),
    .X(_1072_));
 sg13g2_buf_8 _3787_ (.A(net32),
    .X(_1073_));
 sg13g2_o21ai_1 _3788_ (.B1(_1073_),
    .Y(_1074_),
    .A1(net46),
    .A2(_1072_));
 sg13g2_inv_2 _3789_ (.Y(_1075_),
    .A(_1044_));
 sg13g2_buf_1 _3790_ (.A(_1075_),
    .X(_1076_));
 sg13g2_o21ai_1 _3791_ (.B1(\vga.ball_angle[2] ),
    .Y(_1077_),
    .A1(_1055_),
    .A2(_1035_));
 sg13g2_xor2_1 _3792_ (.B(_1077_),
    .A(_0049_),
    .X(_1078_));
 sg13g2_nand2_1 _3793_ (.Y(_1079_),
    .A(_1069_),
    .B(_1070_));
 sg13g2_buf_2 _3794_ (.A(_1079_),
    .X(_1080_));
 sg13g2_nand2_1 _3795_ (.Y(_1081_),
    .A(net142),
    .B(_1991_));
 sg13g2_a21o_1 _3796_ (.A2(_0583_),
    .A1(_1624_),
    .B1(_1081_),
    .X(_1082_));
 sg13g2_or4_1 _3797_ (.A(_1603_),
    .B(net102),
    .C(_1646_),
    .D(net128),
    .X(_1083_));
 sg13g2_buf_1 _3798_ (.A(_1083_),
    .X(_1084_));
 sg13g2_inv_1 _3799_ (.Y(_1085_),
    .A(_1084_));
 sg13g2_nor2_1 _3800_ (.A(net146),
    .B(\vga.ball_angle[3] ),
    .Y(_1086_));
 sg13g2_nor2b_1 _3801_ (.A(_0627_),
    .B_N(_1086_),
    .Y(_1087_));
 sg13g2_a22oi_1 _3802_ (.Y(_1088_),
    .B1(_1085_),
    .B2(_1087_),
    .A2(_1082_),
    .A1(net117));
 sg13g2_nor3_1 _3803_ (.A(net46),
    .B(_1080_),
    .C(_1088_),
    .Y(_1089_));
 sg13g2_a21oi_1 _3804_ (.A1(net46),
    .A2(_1078_),
    .Y(_1090_),
    .B1(_1089_));
 sg13g2_o21ai_1 _3805_ (.B1(net93),
    .Y(_1091_),
    .A1(net29),
    .A2(_1090_));
 sg13g2_a21o_1 _3806_ (.A2(_1074_),
    .A1(net117),
    .B1(_1091_),
    .X(_0096_));
 sg13g2_buf_1 _3807_ (.A(net94),
    .X(_1092_));
 sg13g2_buf_1 _3808_ (.A(_1092_),
    .X(_1093_));
 sg13g2_nand3_1 _3809_ (.B(_2060_),
    .C(_2001_),
    .A(net50),
    .Y(_1094_));
 sg13g2_o21ai_1 _3810_ (.B1(net93),
    .Y(_1095_),
    .A1(_1039_),
    .A2(_1750_));
 sg13g2_a21o_1 _3811_ (.A2(_1094_),
    .A1(net51),
    .B1(_1095_),
    .X(_0097_));
 sg13g2_buf_1 _3812_ (.A(net32),
    .X(_1096_));
 sg13g2_nor2_1 _3813_ (.A(net76),
    .B(net28),
    .Y(_1097_));
 sg13g2_buf_1 _3814_ (.A(_0045_),
    .X(_1098_));
 sg13g2_nor3_1 _3815_ (.A(_1098_),
    .B(net29),
    .C(net46),
    .Y(_1099_));
 sg13g2_o21ai_1 _3816_ (.B1(net92),
    .Y(_0098_),
    .A1(_1097_),
    .A2(_1099_));
 sg13g2_nor2_1 _3817_ (.A(net76),
    .B(net53),
    .Y(_1100_));
 sg13g2_a21oi_1 _3818_ (.A1(net76),
    .A2(_1049_),
    .Y(_1101_),
    .B1(_1100_));
 sg13g2_a21oi_1 _3819_ (.A1(net30),
    .A2(_1101_),
    .Y(_1102_),
    .B1(net71));
 sg13g2_xor2_1 _3820_ (.B(net53),
    .A(net76),
    .X(_1103_));
 sg13g2_and3_1 _3821_ (.X(_1104_),
    .A(net71),
    .B(net32),
    .C(_1103_));
 sg13g2_o21ai_1 _3822_ (.B1(net92),
    .Y(_0099_),
    .A1(_1102_),
    .A2(_1104_));
 sg13g2_or2_1 _3823_ (.X(_1105_),
    .B(net49),
    .A(_1730_));
 sg13g2_buf_1 _3824_ (.A(_1105_),
    .X(_1106_));
 sg13g2_nand2_1 _3825_ (.Y(_1107_),
    .A(_1730_),
    .B(_1047_));
 sg13g2_nand2_2 _3826_ (.Y(_1108_),
    .A(_1106_),
    .B(_1107_));
 sg13g2_nor2_1 _3827_ (.A(net76),
    .B(net71),
    .Y(_1109_));
 sg13g2_nor2_1 _3828_ (.A(net94),
    .B(_1732_),
    .Y(_1110_));
 sg13g2_a21oi_1 _3829_ (.A1(net53),
    .A2(_1109_),
    .Y(_1111_),
    .B1(_1110_));
 sg13g2_nand2_1 _3830_ (.Y(_1112_),
    .A(_1108_),
    .B(_1111_));
 sg13g2_a21oi_1 _3831_ (.A1(net30),
    .A2(_1112_),
    .Y(_1113_),
    .B1(net80));
 sg13g2_inv_1 _3832_ (.Y(_1114_),
    .A(net80));
 sg13g2_nor4_1 _3833_ (.A(_1114_),
    .B(_1075_),
    .C(net46),
    .D(_1111_),
    .Y(_1115_));
 sg13g2_o21ai_1 _3834_ (.B1(net92),
    .Y(_0100_),
    .A1(_1113_),
    .A2(_1115_));
 sg13g2_nor3_1 _3835_ (.A(_1114_),
    .B(_1098_),
    .C(_1049_),
    .Y(_1116_));
 sg13g2_nor2b_1 _3836_ (.A(net80),
    .B_N(_1098_),
    .Y(_1117_));
 sg13g2_o21ai_1 _3837_ (.B1(_1106_),
    .Y(_1118_),
    .A1(_1107_),
    .A2(_1117_));
 sg13g2_nand2b_1 _3838_ (.Y(_1119_),
    .B(_1118_),
    .A_N(_1116_));
 sg13g2_a21oi_1 _3839_ (.A1(net30),
    .A2(_1119_),
    .Y(_1120_),
    .B1(net81));
 sg13g2_nand3_1 _3840_ (.B(net94),
    .C(_1117_),
    .A(net81),
    .Y(_1121_));
 sg13g2_o21ai_1 _3841_ (.B1(_1121_),
    .Y(_1122_),
    .A1(net81),
    .A2(net53));
 sg13g2_nor2_1 _3842_ (.A(_1098_),
    .B(_1735_),
    .Y(_1123_));
 sg13g2_a22oi_1 _3843_ (.Y(_1124_),
    .B1(_1045_),
    .B2(_1123_),
    .A2(net53),
    .A1(_0541_));
 sg13g2_nand2_1 _3844_ (.Y(_1125_),
    .A(net71),
    .B(_1124_));
 sg13g2_o21ai_1 _3845_ (.B1(_1125_),
    .Y(_1126_),
    .A1(net71),
    .A2(_1122_));
 sg13g2_nor2_1 _3846_ (.A(net29),
    .B(_1126_),
    .Y(_1127_));
 sg13g2_o21ai_1 _3847_ (.B1(net92),
    .Y(_0101_),
    .A1(_1120_),
    .A2(_1127_));
 sg13g2_nor2_1 _3848_ (.A(_0515_),
    .B(_0687_),
    .Y(_1128_));
 sg13g2_nor2_1 _3849_ (.A(net94),
    .B(_1737_),
    .Y(_1129_));
 sg13g2_a22oi_1 _3850_ (.Y(_1130_),
    .B1(_1129_),
    .B2(_1747_),
    .A2(_1128_),
    .A1(_1092_));
 sg13g2_inv_1 _3851_ (.Y(_1131_),
    .A(_1130_));
 sg13g2_a21oi_1 _3852_ (.A1(net30),
    .A2(_1131_),
    .Y(_1132_),
    .B1(net79));
 sg13g2_o21ai_1 _3853_ (.B1(net53),
    .Y(_1133_),
    .A1(_2001_),
    .A2(_1128_));
 sg13g2_nand2b_1 _3854_ (.Y(_1134_),
    .B(_1133_),
    .A_N(_1129_));
 sg13g2_and3_1 _3855_ (.X(_1135_),
    .A(net79),
    .B(net32),
    .C(_1134_));
 sg13g2_nor3_1 _3856_ (.A(net57),
    .B(_1132_),
    .C(_1135_),
    .Y(_0102_));
 sg13g2_inv_1 _3857_ (.Y(_1136_),
    .A(_1128_));
 sg13g2_o21ai_1 _3858_ (.B1(net51),
    .Y(_1137_),
    .A1(net79),
    .A2(_1136_));
 sg13g2_a21oi_1 _3859_ (.A1(net30),
    .A2(_1137_),
    .Y(_1138_),
    .B1(_1742_));
 sg13g2_nor2_1 _3860_ (.A(_1098_),
    .B(_0468_),
    .Y(_1139_));
 sg13g2_xnor2_1 _3861_ (.Y(_1140_),
    .A(net136),
    .B(_1139_));
 sg13g2_nor3_1 _3862_ (.A(net79),
    .B(_1741_),
    .C(_1136_),
    .Y(_1141_));
 sg13g2_a21oi_1 _3863_ (.A1(net53),
    .A2(_1141_),
    .Y(_1142_),
    .B1(_2003_));
 sg13g2_o21ai_1 _3864_ (.B1(_1142_),
    .Y(_1143_),
    .A1(_1106_),
    .A2(_1140_));
 sg13g2_a21oi_1 _3865_ (.A1(net28),
    .A2(_1143_),
    .Y(_1144_),
    .B1(_0327_));
 sg13g2_nand2b_1 _3866_ (.Y(_0103_),
    .B(_1144_),
    .A_N(_1138_));
 sg13g2_inv_1 _3867_ (.Y(_1145_),
    .A(_1141_));
 sg13g2_or2_1 _3868_ (.X(_1146_),
    .B(_0474_),
    .A(_1737_));
 sg13g2_a22oi_1 _3869_ (.Y(_1147_),
    .B1(_1146_),
    .B2(_1045_),
    .A2(_1145_),
    .A1(net51));
 sg13g2_and3_1 _3870_ (.X(_1148_),
    .A(net137),
    .B(net32),
    .C(_1147_));
 sg13g2_nor2b_1 _3871_ (.A(net137),
    .B_N(_1146_),
    .Y(_1149_));
 sg13g2_nor3_1 _3872_ (.A(net94),
    .B(net49),
    .C(_1149_),
    .Y(_1150_));
 sg13g2_a21oi_1 _3873_ (.A1(net53),
    .A2(_1141_),
    .Y(_1151_),
    .B1(_1150_));
 sg13g2_nand2_1 _3874_ (.Y(_1152_),
    .A(_2036_),
    .B(_1151_));
 sg13g2_a21oi_1 _3875_ (.A1(net30),
    .A2(_1152_),
    .Y(_1153_),
    .B1(net137));
 sg13g2_o21ai_1 _3876_ (.B1(net92),
    .Y(_0104_),
    .A1(_1148_),
    .A2(_1153_));
 sg13g2_nor3_1 _3877_ (.A(_1098_),
    .B(_0481_),
    .C(_0464_),
    .Y(_1154_));
 sg13g2_o21ai_1 _3878_ (.B1(_1056_),
    .Y(_1155_),
    .A1(_1106_),
    .A2(_1154_));
 sg13g2_nand3_1 _3879_ (.B(_1995_),
    .C(_0683_),
    .A(_1098_),
    .Y(_1156_));
 sg13g2_xnor2_1 _3880_ (.Y(_1157_),
    .A(_0472_),
    .B(_1156_));
 sg13g2_nand3b_1 _3881_ (.B(_1045_),
    .C(_1154_),
    .Y(_1158_),
    .A_N(net77));
 sg13g2_o21ai_1 _3882_ (.B1(_1158_),
    .Y(_1159_),
    .A1(_1107_),
    .A2(_1157_));
 sg13g2_a22oi_1 _3883_ (.Y(_1160_),
    .B1(_1159_),
    .B2(_1096_),
    .A2(_1155_),
    .A1(net77));
 sg13g2_nor2_1 _3884_ (.A(net52),
    .B(_1160_),
    .Y(_0105_));
 sg13g2_and3_1 _3885_ (.X(_1161_),
    .A(net76),
    .B(_0488_),
    .C(_0491_));
 sg13g2_nand2_1 _3886_ (.Y(_1162_),
    .A(_1045_),
    .B(_1161_));
 sg13g2_nor2_1 _3887_ (.A(_0515_),
    .B(_0713_),
    .Y(_1163_));
 sg13g2_xnor2_1 _3888_ (.Y(_1164_),
    .A(_0484_),
    .B(_1163_));
 sg13g2_nand2_1 _3889_ (.Y(_1165_),
    .A(_1049_),
    .B(_1164_));
 sg13g2_o21ai_1 _3890_ (.B1(_1165_),
    .Y(_1166_),
    .A1(net78),
    .A2(_1162_));
 sg13g2_o21ai_1 _3891_ (.B1(_1056_),
    .Y(_1167_),
    .A1(_1106_),
    .A2(_1161_));
 sg13g2_a22oi_1 _3892_ (.Y(_1168_),
    .B1(_1167_),
    .B2(net78),
    .A2(_1166_),
    .A1(_1096_));
 sg13g2_nor2_1 _3893_ (.A(net52),
    .B(_1168_),
    .Y(_0106_));
 sg13g2_nor2_1 _3894_ (.A(_1739_),
    .B(net28),
    .Y(_1169_));
 sg13g2_and3_1 _3895_ (.X(_1170_),
    .A(net77),
    .B(net78),
    .C(_1154_));
 sg13g2_xnor2_1 _3896_ (.Y(_1171_),
    .A(_0707_),
    .B(_1170_));
 sg13g2_nand2b_1 _3897_ (.Y(_1172_),
    .B(_1128_),
    .A_N(_1997_));
 sg13g2_o21ai_1 _3898_ (.B1(_1739_),
    .Y(_1173_),
    .A1(net76),
    .A2(_0711_));
 sg13g2_nand3_1 _3899_ (.B(_1172_),
    .C(_1173_),
    .A(_1047_),
    .Y(_1174_));
 sg13g2_a221oi_1 _3900_ (.B2(net51),
    .C1(net29),
    .B1(_1174_),
    .A1(_1045_),
    .Y(_1175_),
    .A2(_1171_));
 sg13g2_o21ai_1 _3901_ (.B1(net92),
    .Y(_0107_),
    .A1(_1169_),
    .A2(_1175_));
 sg13g2_a21oi_1 _3902_ (.A1(_1624_),
    .A2(_0583_),
    .Y(_1176_),
    .B1(_1081_));
 sg13g2_a21oi_2 _3903_ (.B1(_1080_),
    .Y(_1177_),
    .A2(_1176_),
    .A1(_1063_));
 sg13g2_o21ai_1 _3904_ (.B1(net30),
    .Y(_1178_),
    .A1(net46),
    .A2(_1177_));
 sg13g2_inv_1 _3905_ (.Y(_1179_),
    .A(_1087_));
 sg13g2_o21ai_1 _3906_ (.B1(_1177_),
    .Y(_1180_),
    .A1(_1084_),
    .A2(_1179_));
 sg13g2_nor3_1 _3907_ (.A(net70),
    .B(_1050_),
    .C(_1180_),
    .Y(_1181_));
 sg13g2_a221oi_1 _3908_ (.B2(_1653_),
    .C1(_1181_),
    .B1(_2003_),
    .A1(net131),
    .Y(_1182_),
    .A2(_1749_));
 sg13g2_o21ai_1 _3909_ (.B1(net93),
    .Y(_1183_),
    .A1(net29),
    .A2(_1182_));
 sg13g2_a21o_1 _3910_ (.A2(_1178_),
    .A1(net70),
    .B1(_1183_),
    .X(_0108_));
 sg13g2_buf_1 _3911_ (.A(net134),
    .X(_1184_));
 sg13g2_o21ai_1 _3912_ (.B1(_1086_),
    .Y(_1185_),
    .A1(_0627_),
    .A2(_1084_));
 sg13g2_nand3_1 _3913_ (.B(net117),
    .C(_1082_),
    .A(net70),
    .Y(_1186_));
 sg13g2_a21oi_1 _3914_ (.A1(_1185_),
    .A2(_1186_),
    .Y(_1187_),
    .B1(_1080_));
 sg13g2_xnor2_1 _3915_ (.Y(_1188_),
    .A(net56),
    .B(_1187_));
 sg13g2_nand2_1 _3916_ (.Y(_1189_),
    .A(_1047_),
    .B(_1188_));
 sg13g2_o21ai_1 _3917_ (.B1(_1189_),
    .Y(_1190_),
    .A1(_1655_),
    .A2(_1047_));
 sg13g2_nand2_1 _3918_ (.Y(_1191_),
    .A(_1837_),
    .B(net49));
 sg13g2_nand2b_1 _3919_ (.Y(_1192_),
    .B(_1188_),
    .A_N(net49));
 sg13g2_a21oi_1 _3920_ (.A1(_1191_),
    .A2(_1192_),
    .Y(_1193_),
    .B1(net51));
 sg13g2_a21oi_1 _3921_ (.A1(net51),
    .A2(_1190_),
    .Y(_1194_),
    .B1(_1193_));
 sg13g2_nand2_1 _3922_ (.Y(_1195_),
    .A(net28),
    .B(_1194_));
 sg13g2_nand2_1 _3923_ (.Y(_1196_),
    .A(net56),
    .B(net29));
 sg13g2_nand3_1 _3924_ (.B(_1195_),
    .C(_1196_),
    .A(net68),
    .Y(_0109_));
 sg13g2_nor2_1 _3925_ (.A(net56),
    .B(_1185_),
    .Y(_1197_));
 sg13g2_and3_1 _3926_ (.X(_1198_),
    .A(net56),
    .B(net70),
    .C(net117));
 sg13g2_buf_1 _3927_ (.A(_1198_),
    .X(_1199_));
 sg13g2_o21ai_1 _3928_ (.B1(_1177_),
    .Y(_1200_),
    .A1(_1197_),
    .A2(_1199_));
 sg13g2_nor3_1 _3929_ (.A(net105),
    .B(_1050_),
    .C(_1200_),
    .Y(_1201_));
 sg13g2_a221oi_1 _3930_ (.B2(_1527_),
    .C1(_1201_),
    .B1(_2003_),
    .A1(net61),
    .Y(_1202_),
    .A2(_1749_));
 sg13g2_o21ai_1 _3931_ (.B1(net134),
    .Y(_1203_),
    .A1(_1075_),
    .A2(_1202_));
 sg13g2_nand2_1 _3932_ (.Y(_1204_),
    .A(_1108_),
    .B(_1200_));
 sg13g2_a21oi_1 _3933_ (.A1(net30),
    .A2(_1204_),
    .Y(_1205_),
    .B1(_1519_));
 sg13g2_or2_1 _3934_ (.X(_0110_),
    .B(_1205_),
    .A(_1203_));
 sg13g2_mux2_1 _3935_ (.A0(_1197_),
    .A1(_1199_),
    .S(net105),
    .X(_1206_));
 sg13g2_nand2_1 _3936_ (.Y(_1207_),
    .A(_1177_),
    .B(_1206_));
 sg13g2_nor3_1 _3937_ (.A(net103),
    .B(_1050_),
    .C(_1207_),
    .Y(_1208_));
 sg13g2_a221oi_1 _3938_ (.B2(_1523_),
    .C1(_1208_),
    .B1(_2003_),
    .A1(_1842_),
    .Y(_1209_),
    .A2(_1749_));
 sg13g2_o21ai_1 _3939_ (.B1(net134),
    .Y(_1210_),
    .A1(_1075_),
    .A2(_1209_));
 sg13g2_nand2_1 _3940_ (.Y(_1211_),
    .A(_1108_),
    .B(_1207_));
 sg13g2_a21oi_1 _3941_ (.A1(net32),
    .A2(_1211_),
    .Y(_1212_),
    .B1(_1525_));
 sg13g2_or2_1 _3942_ (.X(_0111_),
    .B(_1212_),
    .A(_1210_));
 sg13g2_nand3_1 _3943_ (.B(net105),
    .C(_1199_),
    .A(_1676_),
    .Y(_1213_));
 sg13g2_nand2_1 _3944_ (.Y(_1214_),
    .A(_0625_),
    .B(_1086_));
 sg13g2_a21oi_1 _3945_ (.A1(_1213_),
    .A2(_1214_),
    .Y(_1215_),
    .B1(_1180_));
 sg13g2_nand3_1 _3946_ (.B(_1108_),
    .C(_1215_),
    .A(_1928_),
    .Y(_1216_));
 sg13g2_a22oi_1 _3947_ (.Y(_1217_),
    .B1(_2003_),
    .B2(_0839_),
    .A2(_1749_),
    .A1(net54));
 sg13g2_nand2_1 _3948_ (.Y(_1218_),
    .A(_1216_),
    .B(_1217_));
 sg13g2_o21ai_1 _3949_ (.B1(net32),
    .Y(_1219_),
    .A1(net46),
    .A2(_1215_));
 sg13g2_a22oi_1 _3950_ (.Y(_1220_),
    .B1(_1219_),
    .B2(net104),
    .A2(_1218_),
    .A1(net28));
 sg13g2_nor2_1 _3951_ (.A(net52),
    .B(_1220_),
    .Y(_0112_));
 sg13g2_and4_1 _3952_ (.A(net146),
    .B(\vga.ball_angle[3] ),
    .C(_0564_),
    .D(_1081_),
    .X(_1221_));
 sg13g2_o21ai_1 _3953_ (.B1(_1072_),
    .Y(_1222_),
    .A1(_1087_),
    .A2(_1221_));
 sg13g2_a21oi_1 _3954_ (.A1(_1084_),
    .A2(_1087_),
    .Y(_1223_),
    .B1(_1221_));
 sg13g2_nor3_1 _3955_ (.A(net109),
    .B(_1080_),
    .C(_1223_),
    .Y(_1224_));
 sg13g2_a21o_1 _3956_ (.A2(_1222_),
    .A1(net109),
    .B1(_1224_),
    .X(_1225_));
 sg13g2_nand2_1 _3957_ (.Y(_1226_),
    .A(_1858_),
    .B(net49));
 sg13g2_o21ai_1 _3958_ (.B1(_1226_),
    .Y(_1227_),
    .A1(net49),
    .A2(_1225_));
 sg13g2_nor2_1 _3959_ (.A(_2001_),
    .B(_1225_),
    .Y(_1228_));
 sg13g2_a21oi_1 _3960_ (.A1(_1687_),
    .A2(_2001_),
    .Y(_1229_),
    .B1(_1228_));
 sg13g2_nand2_1 _3961_ (.Y(_1230_),
    .A(net51),
    .B(_1229_));
 sg13g2_o21ai_1 _3962_ (.B1(_1230_),
    .Y(_1231_),
    .A1(net51),
    .A2(_1227_));
 sg13g2_nand2_1 _3963_ (.Y(_1232_),
    .A(net28),
    .B(_1231_));
 sg13g2_nand2_1 _3964_ (.Y(_1233_),
    .A(net109),
    .B(net29));
 sg13g2_nand3_1 _3965_ (.B(_1232_),
    .C(_1233_),
    .A(net68),
    .Y(_0113_));
 sg13g2_a21o_1 _3966_ (.A2(net47),
    .A1(net70),
    .B1(_1176_),
    .X(_1234_));
 sg13g2_nand3_1 _3967_ (.B(_1084_),
    .C(_1086_),
    .A(_0636_),
    .Y(_1235_));
 sg13g2_inv_1 _3968_ (.Y(_1236_),
    .A(_1235_));
 sg13g2_a21oi_1 _3969_ (.A1(net117),
    .A2(_1234_),
    .Y(_1237_),
    .B1(_1236_));
 sg13g2_a22oi_1 _3970_ (.Y(_1238_),
    .B1(_2003_),
    .B2(_1576_),
    .A2(_1749_),
    .A1(_1889_));
 sg13g2_o21ai_1 _3971_ (.B1(_1238_),
    .Y(_1239_),
    .A1(_1080_),
    .A2(_1237_));
 sg13g2_a21oi_1 _3972_ (.A1(_1073_),
    .A2(_1239_),
    .Y(_1240_),
    .B1(net128));
 sg13g2_nand4_1 _3973_ (.B(_1063_),
    .C(net47),
    .A(net70),
    .Y(_1241_),
    .D(_1082_));
 sg13g2_nand2_1 _3974_ (.Y(_1242_),
    .A(net128),
    .B(_1072_));
 sg13g2_a21oi_1 _3975_ (.A1(_1235_),
    .A2(_1241_),
    .Y(_1243_),
    .B1(_1242_));
 sg13g2_o21ai_1 _3976_ (.B1(_1238_),
    .Y(_1244_),
    .A1(net46),
    .A2(_1243_));
 sg13g2_nor2_1 _3977_ (.A(net29),
    .B(_1244_),
    .Y(_1245_));
 sg13g2_buf_1 _3978_ (.A(net134),
    .X(_1246_));
 sg13g2_o21ai_1 _3979_ (.B1(_1246_),
    .Y(_0114_),
    .A1(_1240_),
    .A2(_1245_));
 sg13g2_nand3_1 _3980_ (.B(net117),
    .C(net47),
    .A(net70),
    .Y(_1247_));
 sg13g2_mux2_1 _3981_ (.A0(_1235_),
    .A1(_1247_),
    .S(net128),
    .X(_1248_));
 sg13g2_a21oi_1 _3982_ (.A1(_1177_),
    .A2(_1248_),
    .Y(_1249_),
    .B1(_1080_));
 sg13g2_nand3b_1 _3983_ (.B(_1177_),
    .C(net102),
    .Y(_1250_),
    .A_N(_1248_));
 sg13g2_o21ai_1 _3984_ (.B1(_1250_),
    .Y(_1251_),
    .A1(net102),
    .A2(_1249_));
 sg13g2_a22oi_1 _3985_ (.Y(_1252_),
    .B1(_2003_),
    .B2(_1583_),
    .A2(_1749_),
    .A1(_1861_));
 sg13g2_o21ai_1 _3986_ (.B1(_1252_),
    .Y(_1253_),
    .A1(_1057_),
    .A2(_1251_));
 sg13g2_nand2_1 _3987_ (.Y(_1254_),
    .A(net28),
    .B(_1253_));
 sg13g2_nand2_1 _3988_ (.Y(_1255_),
    .A(net102),
    .B(_1076_));
 sg13g2_nand3_1 _3989_ (.B(_1254_),
    .C(_1255_),
    .A(net68),
    .Y(_0115_));
 sg13g2_nand2_1 _3990_ (.Y(_1256_),
    .A(net74),
    .B(_1072_));
 sg13g2_nor3_1 _3991_ (.A(net102),
    .B(_0726_),
    .C(net128),
    .Y(_1257_));
 sg13g2_nand3_1 _3992_ (.B(_1084_),
    .C(_1257_),
    .A(_0636_),
    .Y(_1258_));
 sg13g2_mux2_1 _3993_ (.A0(_1256_),
    .A1(net74),
    .S(_1258_),
    .X(_1259_));
 sg13g2_nand3_1 _3994_ (.B(_1991_),
    .C(_0598_),
    .A(_0726_),
    .Y(_1260_));
 sg13g2_a21oi_1 _3995_ (.A1(net117),
    .A2(_1260_),
    .Y(_1261_),
    .B1(_1080_));
 sg13g2_or2_1 _3996_ (.X(_1262_),
    .B(_1261_),
    .A(net74));
 sg13g2_o21ai_1 _3997_ (.B1(_1262_),
    .Y(_1263_),
    .A1(net117),
    .A2(_1259_));
 sg13g2_nor2_1 _3998_ (.A(_2001_),
    .B(_1263_),
    .Y(_1264_));
 sg13g2_a21oi_1 _3999_ (.A1(_1635_),
    .A2(_2001_),
    .Y(_1265_),
    .B1(_1264_));
 sg13g2_nand2_1 _4000_ (.Y(_1266_),
    .A(_1868_),
    .B(_1037_));
 sg13g2_o21ai_1 _4001_ (.B1(_1266_),
    .Y(_1267_),
    .A1(_1037_),
    .A2(_1263_));
 sg13g2_nor2_1 _4002_ (.A(_1093_),
    .B(_1267_),
    .Y(_1268_));
 sg13g2_a21oi_1 _4003_ (.A1(_1093_),
    .A2(_1265_),
    .Y(_1269_),
    .B1(_1268_));
 sg13g2_nand2_1 _4004_ (.Y(_1270_),
    .A(net28),
    .B(_1269_));
 sg13g2_nand2_1 _4005_ (.Y(_1271_),
    .A(_0610_),
    .B(_1076_));
 sg13g2_a21oi_1 _4006_ (.A1(_1270_),
    .A2(_1271_),
    .Y(_0116_),
    .B1(net57));
 sg13g2_nand3_1 _4007_ (.B(_1108_),
    .C(_1070_),
    .A(net50),
    .Y(_1272_));
 sg13g2_buf_1 _4008_ (.A(_1272_),
    .X(_1273_));
 sg13g2_nor3_1 _4009_ (.A(_1064_),
    .B(_1069_),
    .C(_1273_),
    .Y(_1274_));
 sg13g2_a21oi_1 _4010_ (.A1(_1064_),
    .A2(_1273_),
    .Y(_1275_),
    .B1(_1274_));
 sg13g2_nor2_1 _4011_ (.A(net52),
    .B(_1275_),
    .Y(_0117_));
 sg13g2_inv_1 _4012_ (.Y(_1276_),
    .A(_1064_));
 sg13g2_or4_1 _4013_ (.A(_1276_),
    .B(\vga.ball_ratio[1] ),
    .C(_1069_),
    .D(_1273_),
    .X(_1277_));
 sg13g2_nor2_1 _4014_ (.A(_1064_),
    .B(_1069_),
    .Y(_1278_));
 sg13g2_o21ai_1 _4015_ (.B1(\vga.ball_ratio[1] ),
    .Y(_1279_),
    .A1(_1278_),
    .A2(_1273_));
 sg13g2_a21oi_1 _4016_ (.A1(_1277_),
    .A2(_1279_),
    .Y(_0118_),
    .B1(net57));
 sg13g2_nand2_1 _4017_ (.Y(_1280_),
    .A(_1064_),
    .B(\vga.ball_ratio[1] ));
 sg13g2_nor3_1 _4018_ (.A(_1066_),
    .B(_1273_),
    .C(_1280_),
    .Y(_1281_));
 sg13g2_a21oi_1 _4019_ (.A1(_1066_),
    .A2(_1280_),
    .Y(_1282_),
    .B1(_1281_));
 sg13g2_nor2_1 _4020_ (.A(_1069_),
    .B(_1282_),
    .Y(_1283_));
 sg13g2_a21oi_1 _4021_ (.A1(_1066_),
    .A2(_1273_),
    .Y(_1284_),
    .B1(_1283_));
 sg13g2_nor2_1 _4022_ (.A(net52),
    .B(_1284_),
    .Y(_0119_));
 sg13g2_nand3_1 _4023_ (.B(net84),
    .C(_0356_),
    .A(_0700_),
    .Y(_1285_));
 sg13g2_nand3_1 _4024_ (.B(_0795_),
    .C(_1285_),
    .A(_0058_),
    .Y(_1286_));
 sg13g2_nand3_1 _4025_ (.B(net118),
    .C(_1286_),
    .A(net85),
    .Y(_1287_));
 sg13g2_buf_1 _4026_ (.A(_1287_),
    .X(_1288_));
 sg13g2_nor2b_1 _4027_ (.A(_0361_),
    .B_N(_0374_),
    .Y(_1289_));
 sg13g2_nor2b_1 _4028_ (.A(_1288_),
    .B_N(_1289_),
    .Y(_1290_));
 sg13g2_buf_1 _4029_ (.A(_1290_),
    .X(_1291_));
 sg13g2_nand2b_1 _4030_ (.Y(_1292_),
    .B(\vga.blank_h ),
    .A_N(_1291_));
 sg13g2_nand2b_1 _4031_ (.Y(_1293_),
    .B(_0369_),
    .A_N(_0361_));
 sg13g2_nand3_1 _4032_ (.B(_1292_),
    .C(_1293_),
    .A(net68),
    .Y(_0120_));
 sg13g2_or2_1 _4033_ (.X(_1294_),
    .B(_0822_),
    .A(_0263_));
 sg13g2_buf_1 _4034_ (.A(_1294_),
    .X(_1295_));
 sg13g2_nor3_1 _4035_ (.A(_0250_),
    .B(net120),
    .C(_0258_),
    .Y(_1296_));
 sg13g2_nand3_1 _4036_ (.B(_0255_),
    .C(_1296_),
    .A(_0824_),
    .Y(_1297_));
 sg13g2_mux2_1 _4037_ (.A0(_1295_),
    .A1(net73),
    .S(_1297_),
    .X(_1298_));
 sg13g2_nand3_1 _4038_ (.B(net120),
    .C(\vga.count_v[8] ),
    .A(_0256_),
    .Y(_1299_));
 sg13g2_nor2_2 _4039_ (.A(_0824_),
    .B(_1295_),
    .Y(_1300_));
 sg13g2_nor2_1 _4040_ (.A(_0250_),
    .B(_1300_),
    .Y(_1301_));
 sg13g2_inv_1 _4041_ (.Y(_1302_),
    .A(_0255_));
 sg13g2_o21ai_1 _4042_ (.B1(_1302_),
    .Y(_1303_),
    .A1(_1299_),
    .A2(_1301_));
 sg13g2_buf_1 _4043_ (.A(_1303_),
    .X(_1304_));
 sg13g2_nand3b_1 _4044_ (.B(_1298_),
    .C(_1304_),
    .Y(_1305_),
    .A_N(_1288_));
 sg13g2_inv_1 _4045_ (.Y(_1306_),
    .A(_1304_));
 sg13g2_o21ai_1 _4046_ (.B1(\vga.blank_v ),
    .Y(_1307_),
    .A1(_1288_),
    .A2(_1306_));
 sg13g2_nand3_1 _4047_ (.B(_1305_),
    .C(_1307_),
    .A(net68),
    .Y(_0121_));
 sg13g2_nand2b_1 _4048_ (.Y(_1308_),
    .B(_0036_),
    .A_N(_1289_));
 sg13g2_buf_1 _4049_ (.A(_1288_),
    .X(_1309_));
 sg13g2_nand3_1 _4050_ (.B(net48),
    .C(_1289_),
    .A(_0350_),
    .Y(_1310_));
 sg13g2_nand3_1 _4051_ (.B(_1308_),
    .C(_1310_),
    .A(net68),
    .Y(_0123_));
 sg13g2_xnor2_1 _4052_ (.Y(_1311_),
    .A(_0349_),
    .B(_0354_));
 sg13g2_o21ai_1 _4053_ (.B1(net67),
    .Y(_0124_),
    .A1(net45),
    .A2(_1311_));
 sg13g2_xnor2_1 _4054_ (.Y(_1312_),
    .A(_0536_),
    .B(_0772_));
 sg13g2_o21ai_1 _4055_ (.B1(net67),
    .Y(_0125_),
    .A1(net45),
    .A2(_1312_));
 sg13g2_xnor2_1 _4056_ (.Y(_1313_),
    .A(_0351_),
    .B(_0784_));
 sg13g2_o21ai_1 _4057_ (.B1(net67),
    .Y(_0126_),
    .A1(net45),
    .A2(_1313_));
 sg13g2_xnor2_1 _4058_ (.Y(_1314_),
    .A(net84),
    .B(_0356_));
 sg13g2_o21ai_1 _4059_ (.B1(net67),
    .Y(_0127_),
    .A1(net45),
    .A2(_1314_));
 sg13g2_xnor2_1 _4060_ (.Y(_1315_),
    .A(_0700_),
    .B(_0357_));
 sg13g2_o21ai_1 _4061_ (.B1(net67),
    .Y(_0128_),
    .A1(net45),
    .A2(_1315_));
 sg13g2_nand2_1 _4062_ (.Y(_1316_),
    .A(_0356_),
    .B(_0754_));
 sg13g2_xnor2_1 _4063_ (.Y(_1317_),
    .A(_0759_),
    .B(_1316_));
 sg13g2_o21ai_1 _4064_ (.B1(net67),
    .Y(_0129_),
    .A1(net45),
    .A2(_1317_));
 sg13g2_xnor2_1 _4065_ (.Y(_1318_),
    .A(net83),
    .B(_0358_));
 sg13g2_o21ai_1 _4066_ (.B1(net67),
    .Y(_0130_),
    .A1(net45),
    .A2(_1318_));
 sg13g2_nand2_1 _4067_ (.Y(_1319_),
    .A(_0362_),
    .B(_0358_));
 sg13g2_xnor2_1 _4068_ (.Y(_1320_),
    .A(_0750_),
    .B(_1319_));
 sg13g2_o21ai_1 _4069_ (.B1(_1246_),
    .Y(_0131_),
    .A1(_1291_),
    .A2(_1320_));
 sg13g2_nand3_1 _4070_ (.B(net83),
    .C(_0358_),
    .A(net85),
    .Y(_1321_));
 sg13g2_xnor2_1 _4071_ (.Y(_1322_),
    .A(_0342_),
    .B(_1321_));
 sg13g2_o21ai_1 _4072_ (.B1(net67),
    .Y(_0132_),
    .A1(net45),
    .A2(_1322_));
 sg13g2_nand2_1 _4073_ (.Y(_1323_),
    .A(_0037_),
    .B(_1306_));
 sg13g2_nand3_1 _4074_ (.B(_1298_),
    .C(_1304_),
    .A(_0567_),
    .Y(_1324_));
 sg13g2_a21o_1 _4075_ (.A2(_1324_),
    .A1(_1323_),
    .B1(_1288_),
    .X(_1325_));
 sg13g2_nand2_1 _4076_ (.Y(_1326_),
    .A(_0254_),
    .B(net48));
 sg13g2_nand3_1 _4077_ (.B(_1325_),
    .C(_1326_),
    .A(net68),
    .Y(_0133_));
 sg13g2_inv_1 _4078_ (.Y(_1327_),
    .A(_1298_));
 sg13g2_a21oi_1 _4079_ (.A1(_1327_),
    .A2(_1304_),
    .Y(_1328_),
    .B1(_1288_));
 sg13g2_buf_1 _4080_ (.A(_1328_),
    .X(_1329_));
 sg13g2_a21oi_1 _4081_ (.A1(_0567_),
    .A2(net42),
    .Y(_1330_),
    .B1(_1288_));
 sg13g2_a21oi_1 _4082_ (.A1(_0254_),
    .A2(net42),
    .Y(_1331_),
    .B1(_0246_));
 sg13g2_a21oi_1 _4083_ (.A1(_0246_),
    .A2(_1330_),
    .Y(_1332_),
    .B1(_1331_));
 sg13g2_nand2b_1 _4084_ (.Y(_0134_),
    .B(_1053_),
    .A_N(_1332_));
 sg13g2_xor2_1 _4085_ (.B(_0822_),
    .A(_0566_),
    .X(_1333_));
 sg13g2_nand2_1 _4086_ (.Y(_1334_),
    .A(net42),
    .B(_1333_));
 sg13g2_a21oi_1 _4087_ (.A1(net90),
    .A2(net48),
    .Y(_1335_),
    .B1(net57));
 sg13g2_nand2_1 _4088_ (.Y(_0135_),
    .A(_1334_),
    .B(_1335_));
 sg13g2_nand3_1 _4089_ (.B(net89),
    .C(net90),
    .A(net91),
    .Y(_1336_));
 sg13g2_xor2_1 _4090_ (.B(_1336_),
    .A(_0039_),
    .X(_1337_));
 sg13g2_nand2_1 _4091_ (.Y(_1338_),
    .A(net42),
    .B(_1337_));
 sg13g2_a21oi_1 _4092_ (.A1(net59),
    .A2(net48),
    .Y(_1339_),
    .B1(net58));
 sg13g2_nand2_1 _4093_ (.Y(_0136_),
    .A(_1338_),
    .B(_1339_));
 sg13g2_xnor2_1 _4094_ (.Y(_1340_),
    .A(_0593_),
    .B(_1295_));
 sg13g2_nand2_1 _4095_ (.Y(_1341_),
    .A(_1329_),
    .B(_1340_));
 sg13g2_a21oi_1 _4096_ (.A1(_0252_),
    .A2(_1309_),
    .Y(_1342_),
    .B1(net58));
 sg13g2_nand2_1 _4097_ (.Y(_0137_),
    .A(_1341_),
    .B(_1342_));
 sg13g2_xnor2_1 _4098_ (.Y(_1343_),
    .A(_0584_),
    .B(_1300_));
 sg13g2_nand2_1 _4099_ (.Y(_1344_),
    .A(net42),
    .B(_1343_));
 sg13g2_a21oi_1 _4100_ (.A1(net87),
    .A2(net48),
    .Y(_1345_),
    .B1(net58));
 sg13g2_nand2_1 _4101_ (.Y(_0138_),
    .A(_1344_),
    .B(_1345_));
 sg13g2_nand2_1 _4102_ (.Y(_1346_),
    .A(net87),
    .B(_1300_));
 sg13g2_xnor2_1 _4103_ (.Y(_1347_),
    .A(_0561_),
    .B(_1346_));
 sg13g2_nand2_1 _4104_ (.Y(_1348_),
    .A(net42),
    .B(_1347_));
 sg13g2_a21oi_1 _4105_ (.A1(_0596_),
    .A2(net48),
    .Y(_1349_),
    .B1(net58));
 sg13g2_nand2_1 _4106_ (.Y(_0139_),
    .A(_1348_),
    .B(_1349_));
 sg13g2_nand3_1 _4107_ (.B(_0596_),
    .C(_1300_),
    .A(_0273_),
    .Y(_1350_));
 sg13g2_xnor2_1 _4108_ (.Y(_1351_),
    .A(_0928_),
    .B(_1350_));
 sg13g2_nand2_1 _4109_ (.Y(_1352_),
    .A(net42),
    .B(_1351_));
 sg13g2_a21oi_1 _4110_ (.A1(net75),
    .A2(net48),
    .Y(_1353_),
    .B1(net58));
 sg13g2_nand2_1 _4111_ (.Y(_0140_),
    .A(_1352_),
    .B(_1353_));
 sg13g2_or2_1 _4112_ (.X(_1354_),
    .B(_1350_),
    .A(_0663_));
 sg13g2_xnor2_1 _4113_ (.Y(_1355_),
    .A(_0622_),
    .B(_1354_));
 sg13g2_nand2_1 _4114_ (.Y(_1356_),
    .A(_1329_),
    .B(_1355_));
 sg13g2_a21oi_1 _4115_ (.A1(\vga.count_v[8] ),
    .A2(_1309_),
    .Y(_1357_),
    .B1(_0327_));
 sg13g2_nand2_1 _4116_ (.Y(_0141_),
    .A(_1356_),
    .B(_1357_));
 sg13g2_nor2_1 _4117_ (.A(_1299_),
    .B(_1346_),
    .Y(_1358_));
 sg13g2_xnor2_1 _4118_ (.Y(_1359_),
    .A(net73),
    .B(_1358_));
 sg13g2_a22oi_1 _4119_ (.Y(_1360_),
    .B1(net42),
    .B2(_1359_),
    .A2(net48),
    .A1(_0623_));
 sg13g2_nor2_1 _4120_ (.A(_1054_),
    .B(_1360_),
    .Y(_0142_));
 sg13g2_nor2b_1 _4121_ (.A(net130),
    .B_N(_0082_),
    .Y(_1361_));
 sg13g2_a21oi_1 _4122_ (.A1(net61),
    .A2(_1361_),
    .Y(_1362_),
    .B1(_0060_));
 sg13g2_o21ai_1 _4123_ (.B1(net99),
    .Y(_1363_),
    .A1(net97),
    .A2(_1362_));
 sg13g2_nand2_1 _4124_ (.Y(_1364_),
    .A(_1892_),
    .B(_1363_));
 sg13g2_a21o_1 _4125_ (.A2(_1833_),
    .A1(_1850_),
    .B1(net61),
    .X(_1365_));
 sg13g2_nand2b_1 _4126_ (.Y(_1366_),
    .B(net129),
    .A_N(net63));
 sg13g2_a21oi_1 _4127_ (.A1(_1912_),
    .A2(_1365_),
    .Y(_1367_),
    .B1(_1366_));
 sg13g2_nand3_1 _4128_ (.B(net96),
    .C(net60),
    .A(_1868_),
    .Y(_1368_));
 sg13g2_buf_1 _4129_ (.A(\vga.left_down_pressed ),
    .X(_1369_));
 sg13g2_o21ai_1 _4130_ (.B1(_1369_),
    .Y(_1370_),
    .A1(_1367_),
    .A2(_1368_));
 sg13g2_buf_2 _4131_ (.A(_1370_),
    .X(_1371_));
 sg13g2_inv_1 _4132_ (.Y(_1372_),
    .A(_1371_));
 sg13g2_a21oi_1 _4133_ (.A1(\vga.left_up_pressed ),
    .A2(_1364_),
    .Y(_1373_),
    .B1(_1372_));
 sg13g2_nand2_1 _4134_ (.Y(_1374_),
    .A(_1833_),
    .B(_1373_));
 sg13g2_nand2b_1 _4135_ (.Y(_1375_),
    .B(_0082_),
    .A_N(_1373_));
 sg13g2_nand3_1 _4136_ (.B(_1374_),
    .C(_1375_),
    .A(net68),
    .Y(_0173_));
 sg13g2_nand2_1 _4137_ (.Y(_1376_),
    .A(\vga.left_up_pressed ),
    .B(_1364_));
 sg13g2_nor2_1 _4138_ (.A(_1376_),
    .B(_1372_),
    .Y(_1377_));
 sg13g2_buf_2 _4139_ (.A(_1377_),
    .X(_1378_));
 sg13g2_nor2_1 _4140_ (.A(_0082_),
    .B(_1371_),
    .Y(_1379_));
 sg13g2_a21oi_1 _4141_ (.A1(_0082_),
    .A2(_1378_),
    .Y(_1380_),
    .B1(_1379_));
 sg13g2_xnor2_1 _4142_ (.Y(_1381_),
    .A(_1837_),
    .B(_1380_));
 sg13g2_nand2_1 _4143_ (.Y(_0174_),
    .A(net69),
    .B(_1381_));
 sg13g2_nor2_1 _4144_ (.A(_1002_),
    .B(_1371_),
    .Y(_1382_));
 sg13g2_nor3_1 _4145_ (.A(_0942_),
    .B(_1376_),
    .C(_1372_),
    .Y(_1383_));
 sg13g2_nor2_1 _4146_ (.A(_1382_),
    .B(_1383_),
    .Y(_1384_));
 sg13g2_xnor2_1 _4147_ (.Y(_1385_),
    .A(_1831_),
    .B(_1384_));
 sg13g2_nand2_1 _4148_ (.Y(_0175_),
    .A(net69),
    .B(_1385_));
 sg13g2_a21o_1 _4149_ (.A2(_1378_),
    .A1(_0060_),
    .B1(_1382_),
    .X(_1386_));
 sg13g2_a22oi_1 _4150_ (.Y(_1387_),
    .B1(_1386_),
    .B2(_1840_),
    .A2(_1383_),
    .A1(_0060_));
 sg13g2_xor2_1 _4151_ (.B(_1387_),
    .A(net97),
    .X(_1388_));
 sg13g2_nand2_1 _4152_ (.Y(_0176_),
    .A(net69),
    .B(_1388_));
 sg13g2_nor2b_1 _4153_ (.A(net97),
    .B_N(_0060_),
    .Y(_1389_));
 sg13g2_o21ai_1 _4154_ (.B1(_1389_),
    .Y(_1390_),
    .A1(_1840_),
    .A2(_0954_));
 sg13g2_nand2_1 _4155_ (.Y(_1391_),
    .A(_1371_),
    .B(_1390_));
 sg13g2_nor3_2 _4156_ (.A(_1975_),
    .B(_1002_),
    .C(_1371_),
    .Y(_1392_));
 sg13g2_a21oi_1 _4157_ (.A1(_1378_),
    .A2(_1391_),
    .Y(_1393_),
    .B1(_1392_));
 sg13g2_xor2_1 _4158_ (.B(_1393_),
    .A(net54),
    .X(_1394_));
 sg13g2_nor2_1 _4159_ (.A(net52),
    .B(_1394_),
    .Y(_0177_));
 sg13g2_a21oi_1 _4160_ (.A1(net129),
    .A2(_1378_),
    .Y(_1395_),
    .B1(_1392_));
 sg13g2_inv_1 _4161_ (.Y(_1396_),
    .A(_1392_));
 sg13g2_a21oi_1 _4162_ (.A1(_1396_),
    .A2(_1391_),
    .Y(_1397_),
    .B1(net54));
 sg13g2_nor2_1 _4163_ (.A(_1395_),
    .B(_1397_),
    .Y(_1398_));
 sg13g2_xnor2_1 _4164_ (.Y(_1399_),
    .A(net63),
    .B(_1398_));
 sg13g2_nand2_1 _4165_ (.Y(_0178_),
    .A(net69),
    .B(_1399_));
 sg13g2_and3_1 _4166_ (.X(_1400_),
    .A(_1812_),
    .B(net54),
    .C(_1392_));
 sg13g2_o21ai_1 _4167_ (.B1(net129),
    .Y(_1401_),
    .A1(_0968_),
    .A2(_1391_));
 sg13g2_o21ai_1 _4168_ (.B1(_1858_),
    .Y(_1402_),
    .A1(_1392_),
    .A2(_1401_));
 sg13g2_nand2_1 _4169_ (.Y(_1403_),
    .A(_1819_),
    .B(_1402_));
 sg13g2_a21oi_1 _4170_ (.A1(_1371_),
    .A2(_1403_),
    .Y(_1404_),
    .B1(_1400_));
 sg13g2_nand2_1 _4171_ (.Y(_1405_),
    .A(_1378_),
    .B(_1404_));
 sg13g2_nand3b_1 _4172_ (.B(_1405_),
    .C(net60),
    .Y(_1406_),
    .A_N(_1400_));
 sg13g2_xnor2_1 _4173_ (.Y(_1407_),
    .A(_1369_),
    .B(_1404_));
 sg13g2_or3_1 _4174_ (.A(net60),
    .B(_1373_),
    .C(_1407_),
    .X(_1408_));
 sg13g2_nand3_1 _4175_ (.B(_1406_),
    .C(_1408_),
    .A(net93),
    .Y(_0179_));
 sg13g2_nand4_1 _4176_ (.B(_1812_),
    .C(_0968_),
    .A(net60),
    .Y(_1409_),
    .D(_1392_));
 sg13g2_nor2_1 _4177_ (.A(net60),
    .B(_1369_),
    .Y(_1410_));
 sg13g2_nand2_1 _4178_ (.Y(_1411_),
    .A(_1403_),
    .B(_1410_));
 sg13g2_nand3_1 _4179_ (.B(_1371_),
    .C(_1411_),
    .A(_1884_),
    .Y(_1412_));
 sg13g2_a21oi_1 _4180_ (.A1(_1409_),
    .A2(_1412_),
    .Y(_1413_),
    .B1(_1373_));
 sg13g2_nor2_1 _4181_ (.A(_1369_),
    .B(_1376_),
    .Y(_1414_));
 sg13g2_o21ai_1 _4182_ (.B1(_1409_),
    .Y(_1415_),
    .A1(_1884_),
    .A2(_1372_));
 sg13g2_mux2_1 _4183_ (.A0(_1414_),
    .A1(_1369_),
    .S(_1415_),
    .X(_1416_));
 sg13g2_a21oi_1 _4184_ (.A1(_1411_),
    .A2(_1416_),
    .Y(_1417_),
    .B1(net96));
 sg13g2_a21oi_1 _4185_ (.A1(net96),
    .A2(_1413_),
    .Y(_1418_),
    .B1(_1417_));
 sg13g2_nand2b_1 _4186_ (.Y(_0180_),
    .B(_1053_),
    .A_N(_1418_));
 sg13g2_nand2_1 _4187_ (.Y(_1419_),
    .A(_0078_),
    .B(_1378_));
 sg13g2_nand2_1 _4188_ (.Y(_1420_),
    .A(_1409_),
    .B(_1419_));
 sg13g2_and4_1 _4189_ (.A(_0078_),
    .B(_1884_),
    .C(_1378_),
    .D(_1411_),
    .X(_1421_));
 sg13g2_a21oi_1 _4190_ (.A1(net96),
    .A2(_1420_),
    .Y(_1422_),
    .B1(_1421_));
 sg13g2_xnor2_1 _4191_ (.Y(_1423_),
    .A(_1942_),
    .B(_1422_));
 sg13g2_nor2_1 _4192_ (.A(net52),
    .B(_1423_),
    .Y(_0181_));
 sg13g2_nor2b_1 _4193_ (.A(net107),
    .B_N(_0081_),
    .Y(_1424_));
 sg13g2_a21oi_1 _4194_ (.A1(net66),
    .A2(_1424_),
    .Y(_1425_),
    .B1(_0062_));
 sg13g2_o21ai_1 _4195_ (.B1(net55),
    .Y(_1426_),
    .A1(net115),
    .A2(_1425_));
 sg13g2_nand2_1 _4196_ (.Y(_1427_),
    .A(_1605_),
    .B(_1426_));
 sg13g2_nand2_1 _4197_ (.Y(_1428_),
    .A(\vga.right_up_pressed ),
    .B(_1427_));
 sg13g2_buf_2 _4198_ (.A(\vga.right_down_pressed ),
    .X(_1429_));
 sg13g2_nand2b_1 _4199_ (.Y(_1430_),
    .B(_1522_),
    .A_N(net114));
 sg13g2_a21oi_1 _4200_ (.A1(_1508_),
    .A2(_1512_),
    .Y(_1431_),
    .B1(net116));
 sg13g2_o21ai_1 _4201_ (.B1(net140),
    .Y(_1432_),
    .A1(_1430_),
    .A2(_1431_));
 sg13g2_nand3_1 _4202_ (.B(net110),
    .C(net112),
    .A(_1583_),
    .Y(_1433_));
 sg13g2_inv_1 _4203_ (.Y(_1434_),
    .A(_1433_));
 sg13g2_o21ai_1 _4204_ (.B1(_1434_),
    .Y(_1435_),
    .A1(net64),
    .A2(_1432_));
 sg13g2_nand2_2 _4205_ (.Y(_1436_),
    .A(_1429_),
    .B(_1435_));
 sg13g2_and2_1 _4206_ (.A(_1428_),
    .B(_1436_),
    .X(_1437_));
 sg13g2_buf_1 _4207_ (.A(_1437_),
    .X(_1438_));
 sg13g2_nor2b_1 _4208_ (.A(net108),
    .B_N(_1438_),
    .Y(_1439_));
 sg13g2_nor2_1 _4209_ (.A(_0081_),
    .B(_1438_),
    .Y(_1440_));
 sg13g2_o21ai_1 _4210_ (.B1(_1184_),
    .Y(_0182_),
    .A1(_1439_),
    .A2(_1440_));
 sg13g2_nor2b_1 _4211_ (.A(_1428_),
    .B_N(_1436_),
    .Y(_1441_));
 sg13g2_buf_1 _4212_ (.A(_1441_),
    .X(_1442_));
 sg13g2_nor2_1 _4213_ (.A(_0081_),
    .B(_1436_),
    .Y(_1443_));
 sg13g2_a21oi_1 _4214_ (.A1(_0081_),
    .A2(_1442_),
    .Y(_1444_),
    .B1(_1443_));
 sg13g2_xnor2_1 _4215_ (.Y(_1445_),
    .A(_1509_),
    .B(_1444_));
 sg13g2_nand2_1 _4216_ (.Y(_0183_),
    .A(net69),
    .B(_1445_));
 sg13g2_and4_1 _4217_ (.A(net107),
    .B(_1653_),
    .C(_1429_),
    .D(_1435_),
    .X(_1446_));
 sg13g2_buf_1 _4218_ (.A(_1446_),
    .X(_1447_));
 sg13g2_and2_1 _4219_ (.A(_0833_),
    .B(_1442_),
    .X(_1448_));
 sg13g2_nor2_1 _4220_ (.A(_1447_),
    .B(_1448_),
    .Y(_1449_));
 sg13g2_xnor2_1 _4221_ (.Y(_1450_),
    .A(_1517_),
    .B(_1449_));
 sg13g2_nand2_1 _4222_ (.Y(_0184_),
    .A(net69),
    .B(_1450_));
 sg13g2_a21o_1 _4223_ (.A2(_1442_),
    .A1(_0062_),
    .B1(_1447_),
    .X(_1451_));
 sg13g2_a22oi_1 _4224_ (.Y(_1452_),
    .B1(_1451_),
    .B2(net66),
    .A2(_1448_),
    .A1(_0062_));
 sg13g2_xor2_1 _4225_ (.B(_1452_),
    .A(_1523_),
    .X(_1453_));
 sg13g2_nand2_1 _4226_ (.Y(_0185_),
    .A(net69),
    .B(_1453_));
 sg13g2_inv_1 _4227_ (.Y(_1454_),
    .A(_0062_));
 sg13g2_nor2_1 _4228_ (.A(_1527_),
    .B(_0833_),
    .Y(_1455_));
 sg13g2_nor3_1 _4229_ (.A(net115),
    .B(_1454_),
    .C(_1455_),
    .Y(_1456_));
 sg13g2_a22oi_1 _4230_ (.Y(_1457_),
    .B1(_1456_),
    .B2(_1442_),
    .A2(_1447_),
    .A1(_1540_));
 sg13g2_xor2_1 _4231_ (.B(_1457_),
    .A(net55),
    .X(_1458_));
 sg13g2_nor2_1 _4232_ (.A(net57),
    .B(_1458_),
    .Y(_0186_));
 sg13g2_o21ai_1 _4233_ (.B1(net140),
    .Y(_1459_),
    .A1(_0839_),
    .A2(_1456_));
 sg13g2_and3_1 _4234_ (.X(_1460_),
    .A(net55),
    .B(_1540_),
    .C(_1447_));
 sg13g2_a21o_1 _4235_ (.A2(_1459_),
    .A1(_1436_),
    .B1(_1460_),
    .X(_1461_));
 sg13g2_buf_1 _4236_ (.A(_1461_),
    .X(_1462_));
 sg13g2_nor2_1 _4237_ (.A(net64),
    .B(_1433_),
    .Y(_1463_));
 sg13g2_inv_1 _4238_ (.Y(_1464_),
    .A(_1429_));
 sg13g2_a21oi_1 _4239_ (.A1(_1432_),
    .A2(_1463_),
    .Y(_1465_),
    .B1(_1464_));
 sg13g2_nor3_1 _4240_ (.A(_1428_),
    .B(_1462_),
    .C(_1465_),
    .Y(_1466_));
 sg13g2_a21oi_1 _4241_ (.A1(_1462_),
    .A2(_1465_),
    .Y(_1467_),
    .B1(_1466_));
 sg13g2_inv_1 _4242_ (.Y(_1468_),
    .A(_1442_));
 sg13g2_nor2_1 _4243_ (.A(_1687_),
    .B(_1460_),
    .Y(_1469_));
 sg13g2_o21ai_1 _4244_ (.B1(_1469_),
    .Y(_1470_),
    .A1(_1468_),
    .A2(_1462_));
 sg13g2_o21ai_1 _4245_ (.B1(_1470_),
    .Y(_1471_),
    .A1(_1647_),
    .A2(_1467_));
 sg13g2_nand2b_1 _4246_ (.Y(_0187_),
    .B(_2123_),
    .A_N(_1471_));
 sg13g2_a21oi_1 _4247_ (.A1(_1647_),
    .A2(_1462_),
    .Y(_1472_),
    .B1(_1464_));
 sg13g2_nor2_1 _4248_ (.A(_1438_),
    .B(_1472_),
    .Y(_1473_));
 sg13g2_nor2_1 _4249_ (.A(net112),
    .B(_1473_),
    .Y(_1474_));
 sg13g2_nor2_1 _4250_ (.A(net112),
    .B(_1429_),
    .Y(_1475_));
 sg13g2_a21o_1 _4251_ (.A2(_1462_),
    .A1(_1687_),
    .B1(_1563_),
    .X(_1476_));
 sg13g2_nor2b_1 _4252_ (.A(_1638_),
    .B_N(_1460_),
    .Y(_1477_));
 sg13g2_a21oi_1 _4253_ (.A1(_1475_),
    .A2(_1476_),
    .Y(_1478_),
    .B1(_1477_));
 sg13g2_and3_1 _4254_ (.X(_1479_),
    .A(net110),
    .B(_1628_),
    .C(_1465_));
 sg13g2_nand2b_1 _4255_ (.Y(_1480_),
    .B(net112),
    .A_N(_1465_));
 sg13g2_a21oi_1 _4256_ (.A1(_1687_),
    .A2(_1462_),
    .Y(_1481_),
    .B1(_1480_));
 sg13g2_o21ai_1 _4257_ (.B1(_1535_),
    .Y(_1482_),
    .A1(_1479_),
    .A2(_1481_));
 sg13g2_a21oi_1 _4258_ (.A1(_1478_),
    .A2(_1482_),
    .Y(_1483_),
    .B1(_1438_));
 sg13g2_o21ai_1 _4259_ (.B1(_1184_),
    .Y(_0188_),
    .A1(_1474_),
    .A2(_1483_));
 sg13g2_and2_1 _4260_ (.A(_1507_),
    .B(_1478_),
    .X(_1484_));
 sg13g2_buf_1 _4261_ (.A(_1484_),
    .X(_1485_));
 sg13g2_inv_1 _4262_ (.Y(_1486_),
    .A(_1507_));
 sg13g2_a21oi_1 _4263_ (.A1(_1486_),
    .A2(_1436_),
    .Y(_1487_),
    .B1(_1477_));
 sg13g2_a21oi_1 _4264_ (.A1(_1429_),
    .A2(_1487_),
    .Y(_1488_),
    .B1(_1438_));
 sg13g2_o21ai_1 _4265_ (.B1(_1488_),
    .Y(_1489_),
    .A1(_1429_),
    .A2(_1485_));
 sg13g2_nand2b_1 _4266_ (.Y(_1490_),
    .B(net141),
    .A_N(_1477_));
 sg13g2_a21oi_1 _4267_ (.A1(_1442_),
    .A2(_1485_),
    .Y(_1491_),
    .B1(_1490_));
 sg13g2_nor2_1 _4268_ (.A(net58),
    .B(_1491_),
    .Y(_1492_));
 sg13g2_o21ai_1 _4269_ (.B1(_1492_),
    .Y(_0189_),
    .A1(net141),
    .A2(_1489_));
 sg13g2_nor2_1 _4270_ (.A(_1569_),
    .B(_1468_),
    .Y(_1493_));
 sg13g2_or2_1 _4271_ (.X(_1494_),
    .B(_1493_),
    .A(_1477_));
 sg13g2_a22oi_1 _4272_ (.Y(_1495_),
    .B1(_1494_),
    .B2(net141),
    .A2(_1493_),
    .A1(_1485_));
 sg13g2_xor2_1 _4273_ (.B(_1495_),
    .A(net110),
    .X(_1496_));
 sg13g2_nor2_1 _4274_ (.A(net57),
    .B(_1496_),
    .Y(_0190_));
 sg13g2_nor2_1 _4275_ (.A(net57),
    .B(_2088_),
    .Y(_0197_));
 sg13g2_o21ai_1 _4276_ (.B1(net148),
    .Y(_1497_),
    .A1(_1754_),
    .A2(_1756_));
 sg13g2_a21oi_1 _4277_ (.A1(_1763_),
    .A2(_1497_),
    .Y(_0201_),
    .B1(_0338_));
 sg13g2_nor2_1 _4278_ (.A(_1054_),
    .B(net40),
    .Y(_0208_));
 sg13g2_o21ai_1 _4279_ (.B1(net133),
    .Y(_1498_),
    .A1(net126),
    .A2(_2009_));
 sg13g2_a21oi_1 _4280_ (.A1(_2010_),
    .A2(_1498_),
    .Y(_0210_),
    .B1(_0338_));
 sg13g2_and2_1 _4281_ (.A(net93),
    .B(net5),
    .X(_0214_));
 sg13g2_and2_1 _4282_ (.A(_2076_),
    .B(_0377_),
    .X(_0215_));
 sg13g2_nand4_1 _4283_ (.B(_0272_),
    .C(_0273_),
    .A(_0248_),
    .Y(_1499_),
    .D(_0824_));
 sg13g2_nor4_1 _4284_ (.A(net72),
    .B(_0080_),
    .C(_1299_),
    .D(_1499_),
    .Y(_1500_));
 sg13g2_mux2_1 _4285_ (.A0(_1500_),
    .A1(\vga.vs_out ),
    .S(_1305_),
    .X(_1501_));
 sg13g2_and2_1 _4286_ (.A(net93),
    .B(_1501_),
    .X(_0216_));
 sg13g2_buf_1 _4287_ (.A(ui_in[7]),
    .X(_1502_));
 sg13g2_inv_1 _4288_ (.Y(net13),
    .A(_1502_));
 sg13g2_nor2b_1 _4289_ (.A(_1502_),
    .B_N(g0),
    .Y(_1503_));
 sg13g2_a21o_1 _4290_ (.A2(b0),
    .A1(_1502_),
    .B1(_1503_),
    .X(net22));
 sg13g2_a21o_1 _4291_ (.A2(\vga.vs ),
    .A1(_1502_),
    .B1(_1503_),
    .X(net23));
 sg13g2_nor2b_1 _4292_ (.A(_1502_),
    .B_N(b0),
    .Y(_1504_));
 sg13g2_a21o_1 _4293_ (.A2(g0),
    .A1(_1502_),
    .B1(_1504_),
    .X(net25));
 sg13g2_a21o_1 _4294_ (.A2(hs),
    .A1(_1502_),
    .B1(_1504_),
    .X(net27));
 sg13g2_dfrbp_1 _4295_ (.CLK(clknet_5_17__leaf_clk),
    .RESET_B(net151),
    .D(_0006_),
    .Q_N(_2214_),
    .Q(_0026_));
 sg13g2_dfrbp_1 _4296_ (.CLK(clknet_5_20__leaf_clk),
    .RESET_B(net152),
    .D(_0007_),
    .Q_N(_2213_),
    .Q(_0027_));
 sg13g2_dfrbp_1 _4297_ (.CLK(clknet_5_7__leaf_clk),
    .RESET_B(net153),
    .D(_0085_),
    .Q_N(_2212_),
    .Q(_0030_));
 sg13g2_dfrbp_1 _4298_ (.CLK(clknet_5_6__leaf_clk),
    .RESET_B(net154),
    .D(_0086_),
    .Q_N(_2215_),
    .Q(_0022_));
 sg13g2_dfrbp_1 _4299_ (.CLK(clknet_5_7__leaf_clk),
    .RESET_B(net155),
    .D(_0002_),
    .Q_N(_2216_),
    .Q(_0021_));
 sg13g2_dfrbp_1 _4300_ (.CLK(clknet_5_6__leaf_clk),
    .RESET_B(net156),
    .D(_0003_),
    .Q_N(_2217_),
    .Q(_0023_));
 sg13g2_dfrbp_1 _4301_ (.CLK(clknet_5_16__leaf_clk),
    .RESET_B(net157),
    .D(_0010_),
    .Q_N(_2218_),
    .Q(_0032_));
 sg13g2_dfrbp_1 _4302_ (.CLK(clknet_5_17__leaf_clk),
    .RESET_B(net158),
    .D(_0011_),
    .Q_N(_2219_),
    .Q(_0033_));
 sg13g2_dfrbp_1 _4303_ (.CLK(clknet_5_16__leaf_clk),
    .RESET_B(net159),
    .D(_0000_),
    .Q_N(_2220_),
    .Q(_0018_));
 sg13g2_dfrbp_1 _4304_ (.CLK(clknet_5_16__leaf_clk),
    .RESET_B(net160),
    .D(_0001_),
    .Q_N(_2211_),
    .Q(_0020_));
 sg13g2_dfrbp_1 _4305_ (.CLK(clknet_5_6__leaf_clk),
    .RESET_B(net161),
    .D(_0087_),
    .Q_N(_2221_),
    .Q(_0017_));
 sg13g2_dfrbp_1 _4306_ (.CLK(clknet_5_21__leaf_clk),
    .RESET_B(net162),
    .D(_0009_),
    .Q_N(_2222_),
    .Q(_0031_));
 sg13g2_dfrbp_1 _4307_ (.CLK(clknet_5_19__leaf_clk),
    .RESET_B(net163),
    .D(_0012_),
    .Q_N(_2223_),
    .Q(_0034_));
 sg13g2_dfrbp_1 _4308_ (.CLK(clknet_5_20__leaf_clk),
    .RESET_B(net164),
    .D(_0013_),
    .Q_N(_2210_),
    .Q(_0035_));
 sg13g2_dfrbp_1 _4309_ (.CLK(clknet_5_5__leaf_clk),
    .RESET_B(net165),
    .D(_0088_),
    .Q_N(_2224_),
    .Q(_0015_));
 sg13g2_dfrbp_1 _4310_ (.CLK(clknet_5_17__leaf_clk),
    .RESET_B(net166),
    .D(_0008_),
    .Q_N(_2209_),
    .Q(_0029_));
 sg13g2_dfrbp_1 _4311_ (.CLK(clknet_5_16__leaf_clk),
    .RESET_B(net167),
    .D(_0089_),
    .Q_N(_2208_),
    .Q(_0028_));
 sg13g2_dfrbp_1 _4312_ (.CLK(clknet_5_5__leaf_clk),
    .RESET_B(net168),
    .D(_0090_),
    .Q_N(_2207_),
    .Q(_0019_));
 sg13g2_dfrbp_1 _4313_ (.CLK(clknet_5_5__leaf_clk),
    .RESET_B(net169),
    .D(_0091_),
    .Q_N(_2225_),
    .Q(_0014_));
 sg13g2_dfrbp_1 _4314_ (.CLK(clknet_5_17__leaf_clk),
    .RESET_B(net170),
    .D(_0004_),
    .Q_N(_2226_),
    .Q(_0024_));
 sg13g2_dfrbp_1 _4315_ (.CLK(clknet_5_17__leaf_clk),
    .RESET_B(net171),
    .D(_0005_),
    .Q_N(_2206_),
    .Q(_0025_));
 sg13g2_dfrbp_1 _4316_ (.CLK(clknet_5_7__leaf_clk),
    .RESET_B(net172),
    .D(_0092_),
    .Q_N(_2205_),
    .Q(_0016_));
 sg13g2_buf_1 clkbuf_0_clk (.A(clk),
    .X(clknet_0_clk));
 sg13g2_tiehi _4295__151 (.L_HI(net151));
 sg13g2_buf_1 _4319_ (.A(net13),
    .X(net6));
 sg13g2_buf_1 _4320_ (.A(net13),
    .X(net7));
 sg13g2_buf_1 _4321_ (.A(net13),
    .X(net8));
 sg13g2_buf_1 _4322_ (.A(net13),
    .X(net9));
 sg13g2_buf_1 _4323_ (.A(net13),
    .X(net10));
 sg13g2_buf_1 _4324_ (.A(net13),
    .X(net11));
 sg13g2_buf_1 _4325_ (.A(net13),
    .X(net12));
 sg13g2_buf_1 _4326_ (.A(g0),
    .X(net14));
 sg13g2_buf_1 _4327_ (.A(g0),
    .X(net15));
 sg13g2_buf_1 _4328_ (.A(g0),
    .X(net16));
 sg13g2_buf_1 _4329_ (.A(g0),
    .X(net17));
 sg13g2_buf_1 _4330_ (.A(hs),
    .X(net18));
 sg13g2_buf_1 _4331_ (.A(\vga.vs ),
    .X(net19));
 sg13g2_buf_1 _4332_ (.A(net149),
    .X(uio_out[6]));
 sg13g2_buf_1 _4333_ (.A(net150),
    .X(uio_out[7]));
 sg13g2_buf_1 _4334_ (.A(g0),
    .X(net20));
 sg13g2_buf_1 _4335_ (.A(g0),
    .X(net21));
 sg13g2_buf_1 _4336_ (.A(net25),
    .X(net24));
 sg13g2_buf_1 _4337_ (.A(b0),
    .X(net26));
 sg13g2_dfrbp_1 \vga.ball_angle[0]$_SDFFE_PN1P_  (.CLK(clknet_5_13__leaf_clk),
    .RESET_B(net173),
    .D(_0093_),
    .Q_N(_0084_),
    .Q(\vga.ball_angle[0] ));
 sg13g2_dfrbp_1 \vga.ball_angle[1]$_SDFFE_PN0P_  (.CLK(clknet_5_18__leaf_clk),
    .RESET_B(net174),
    .D(_0094_),
    .Q_N(_2204_),
    .Q(\vga.ball_angle[1] ));
 sg13g2_dfrbp_1 \vga.ball_angle[2]$_SDFFE_PN0P_  (.CLK(clknet_5_1__leaf_clk),
    .RESET_B(net175),
    .D(_0095_),
    .Q_N(_0063_),
    .Q(\vga.ball_angle[2] ));
 sg13g2_dfrbp_1 \vga.ball_angle[3]$_SDFFE_PN1P_  (.CLK(clknet_5_14__leaf_clk),
    .RESET_B(net176),
    .D(_0096_),
    .Q_N(_0049_),
    .Q(\vga.ball_angle[3] ));
 sg13g2_dfrbp_1 \vga.ball_motion_l$_SDFFE_PN1N_  (.CLK(clknet_5_1__leaf_clk),
    .RESET_B(net177),
    .D(_0097_),
    .Q_N(_0064_),
    .Q(\vga.ball_motion_l ));
 sg13g2_dfrbp_1 \vga.ball_pos_h[0]$_SDFFE_PN1P_  (.CLK(clknet_5_9__leaf_clk),
    .RESET_B(net178),
    .D(_0098_),
    .Q_N(_0045_),
    .Q(\vga.ball_pos_h[0] ));
 sg13g2_dfrbp_1 \vga.ball_pos_h[1]$_SDFFE_PN1P_  (.CLK(clknet_5_8__leaf_clk),
    .RESET_B(net179),
    .D(_0099_),
    .Q_N(_0057_),
    .Q(\vga.ball_pos_h[1] ));
 sg13g2_dfrbp_1 \vga.ball_pos_h[2]$_SDFFE_PN1P_  (.CLK(clknet_5_9__leaf_clk),
    .RESET_B(net180),
    .D(_0100_),
    .Q_N(_2203_),
    .Q(\vga.ball_pos_h[2] ));
 sg13g2_dfrbp_1 \vga.ball_pos_h[3]$_SDFFE_PN1P_  (.CLK(clknet_5_8__leaf_clk),
    .RESET_B(net181),
    .D(_0101_),
    .Q_N(_2202_),
    .Q(\vga.ball_pos_h[3] ));
 sg13g2_dfrbp_1 \vga.ball_pos_h[4]$_SDFFE_PN0P_  (.CLK(clknet_5_8__leaf_clk),
    .RESET_B(net182),
    .D(_0102_),
    .Q_N(_2201_),
    .Q(\vga.ball_pos_h[4] ));
 sg13g2_dfrbp_1 \vga.ball_pos_h[5]$_SDFFE_PN1P_  (.CLK(clknet_5_9__leaf_clk),
    .RESET_B(net183),
    .D(_0103_),
    .Q_N(_0052_),
    .Q(\vga.ball_pos_h[5] ));
 sg13g2_dfrbp_1 \vga.ball_pos_h[6]$_SDFFE_PN1P_  (.CLK(clknet_5_12__leaf_clk),
    .RESET_B(net184),
    .D(_0104_),
    .Q_N(_2200_),
    .Q(\vga.ball_pos_h[6] ));
 sg13g2_dfrbp_1 \vga.ball_pos_h[7]$_SDFFE_PN0P_  (.CLK(clknet_5_12__leaf_clk),
    .RESET_B(net185),
    .D(_0105_),
    .Q_N(_0046_),
    .Q(\vga.ball_pos_h[7] ));
 sg13g2_dfrbp_1 \vga.ball_pos_h[8]$_SDFFE_PN0P_  (.CLK(clknet_5_12__leaf_clk),
    .RESET_B(net186),
    .D(_0106_),
    .Q_N(_0047_),
    .Q(\vga.ball_pos_h[8] ));
 sg13g2_dfrbp_1 \vga.ball_pos_h[9]$_SDFFE_PN1P_  (.CLK(clknet_5_14__leaf_clk),
    .RESET_B(net187),
    .D(_0107_),
    .Q_N(_0048_),
    .Q(\vga.ball_pos_h[9] ));
 sg13g2_dfrbp_1 \vga.ball_pos_v[0]$_SDFFE_PN1P_  (.CLK(clknet_5_14__leaf_clk),
    .RESET_B(net188),
    .D(_0108_),
    .Q_N(_2199_),
    .Q(\vga.ball_pos_v[0] ));
 sg13g2_dfrbp_1 \vga.ball_pos_v[1]$_SDFFE_PN1P_  (.CLK(clknet_5_8__leaf_clk),
    .RESET_B(net189),
    .D(_0109_),
    .Q_N(_2198_),
    .Q(\vga.ball_pos_v[1] ));
 sg13g2_dfrbp_1 \vga.ball_pos_v[2]$_SDFFE_PN1P_  (.CLK(clknet_5_11__leaf_clk),
    .RESET_B(net190),
    .D(_0110_),
    .Q_N(_2197_),
    .Q(\vga.ball_pos_v[2] ));
 sg13g2_dfrbp_1 \vga.ball_pos_v[3]$_SDFFE_PN1P_  (.CLK(clknet_5_11__leaf_clk),
    .RESET_B(net191),
    .D(_0111_),
    .Q_N(_0075_),
    .Q(\vga.ball_pos_v[3] ));
 sg13g2_dfrbp_1 \vga.ball_pos_v[4]$_SDFFE_PN0P_  (.CLK(clknet_5_11__leaf_clk),
    .RESET_B(net192),
    .D(_0112_),
    .Q_N(_2196_),
    .Q(\vga.ball_pos_v[4] ));
 sg13g2_dfrbp_1 \vga.ball_pos_v[5]$_SDFFE_PN1P_  (.CLK(clknet_5_8__leaf_clk),
    .RESET_B(net193),
    .D(_0113_),
    .Q_N(_0074_),
    .Q(\vga.ball_pos_v[5] ));
 sg13g2_dfrbp_1 \vga.ball_pos_v[6]$_SDFFE_PN1P_  (.CLK(clknet_5_2__leaf_clk),
    .RESET_B(net194),
    .D(_0114_),
    .Q_N(_0071_),
    .Q(\vga.ball_pos_v[6] ));
 sg13g2_dfrbp_1 \vga.ball_pos_v[7]$_SDFFE_PN1P_  (.CLK(clknet_5_15__leaf_clk),
    .RESET_B(net195),
    .D(_0115_),
    .Q_N(_0073_),
    .Q(\vga.ball_pos_v[7] ));
 sg13g2_dfrbp_1 \vga.ball_pos_v[8]$_SDFFE_PN0P_  (.CLK(clknet_5_2__leaf_clk),
    .RESET_B(net196),
    .D(_0116_),
    .Q_N(_0067_),
    .Q(\vga.ball_pos_v[8] ));
 sg13g2_dfrbp_1 \vga.ball_ratio[0]$_SDFFE_PN0P_  (.CLK(clknet_5_22__leaf_clk),
    .RESET_B(net197),
    .D(_0117_),
    .Q_N(_2195_),
    .Q(\vga.ball_ratio[0] ));
 sg13g2_dfrbp_1 \vga.ball_ratio[1]$_SDFFE_PN0P_  (.CLK(clknet_5_24__leaf_clk),
    .RESET_B(net198),
    .D(_0118_),
    .Q_N(_2194_),
    .Q(\vga.ball_ratio[1] ));
 sg13g2_dfrbp_1 \vga.ball_ratio[2]$_SDFFE_PN0P_  (.CLK(clknet_5_18__leaf_clk),
    .RESET_B(net199),
    .D(_0119_),
    .Q_N(_2193_),
    .Q(\vga.ball_ratio[2] ));
 sg13g2_dfrbp_1 \vga.blank_h$_SDFFE_PN1P_  (.CLK(clknet_5_0__leaf_clk),
    .RESET_B(net200),
    .D(_0120_),
    .Q_N(_2192_),
    .Q(\vga.blank_h ));
 sg13g2_dfrbp_1 \vga.blank_v$_SDFFE_PN1P_  (.CLK(clknet_5_0__leaf_clk),
    .RESET_B(net201),
    .D(_0121_),
    .Q_N(_2191_),
    .Q(\vga.blank_v ));
 sg13g2_dfrbp_1 \vga.blu$_SDFF_PN0_  (.CLK(clknet_5_21__leaf_clk),
    .RESET_B(net202),
    .D(_0122_),
    .Q_N(_2190_),
    .Q(b0));
 sg13g2_dfrbp_1 \vga.count_h[0]$_SDFF_PN1_  (.CLK(clknet_5_0__leaf_clk),
    .RESET_B(net203),
    .D(_0123_),
    .Q_N(_0036_),
    .Q(\vga.count_h[0] ));
 sg13g2_dfrbp_1 \vga.count_h[1]$_SDFF_PN1_  (.CLK(clknet_5_4__leaf_clk),
    .RESET_B(net204),
    .D(_0124_),
    .Q_N(_0051_),
    .Q(\vga.count_h[1] ));
 sg13g2_dfrbp_1 \vga.count_h[2]$_SDFF_PN1_  (.CLK(clknet_5_9__leaf_clk),
    .RESET_B(net205),
    .D(_0125_),
    .Q_N(_0053_),
    .Q(\vga.count_h[2] ));
 sg13g2_dfrbp_1 \vga.count_h[3]$_SDFF_PN1_  (.CLK(clknet_5_4__leaf_clk),
    .RESET_B(net206),
    .D(_0126_),
    .Q_N(_2189_),
    .Q(\vga.count_h[3] ));
 sg13g2_dfrbp_1 \vga.count_h[4]$_SDFF_PN1_  (.CLK(clknet_5_12__leaf_clk),
    .RESET_B(net207),
    .D(_0127_),
    .Q_N(_0056_),
    .Q(\vga.count_h[4] ));
 sg13g2_dfrbp_1 \vga.count_h[5]$_SDFF_PN1_  (.CLK(clknet_5_4__leaf_clk),
    .RESET_B(net208),
    .D(_0128_),
    .Q_N(_0058_),
    .Q(\vga.count_h[5] ));
 sg13g2_dfrbp_1 \vga.count_h[6]$_SDFF_PN1_  (.CLK(clknet_5_12__leaf_clk),
    .RESET_B(net209),
    .D(_0129_),
    .Q_N(_0055_),
    .Q(\vga.count_h[6] ));
 sg13g2_dfrbp_1 \vga.count_h[7]$_SDFF_PN1_  (.CLK(clknet_5_13__leaf_clk),
    .RESET_B(net210),
    .D(_0130_),
    .Q_N(_0050_),
    .Q(\vga.count_h[7] ));
 sg13g2_dfrbp_1 \vga.count_h[8]$_SDFF_PN1_  (.CLK(clknet_5_13__leaf_clk),
    .RESET_B(net211),
    .D(_0131_),
    .Q_N(_0054_),
    .Q(\vga.count_h[8] ));
 sg13g2_dfrbp_1 \vga.count_h[9]$_SDFF_PN1_  (.CLK(clknet_5_13__leaf_clk),
    .RESET_B(net212),
    .D(_0132_),
    .Q_N(_0066_),
    .Q(\vga.count_h[9] ));
 sg13g2_dfrbp_1 \vga.count_v[0]$_SDFFE_PN1N_  (.CLK(clknet_5_3__leaf_clk),
    .RESET_B(net213),
    .D(_0133_),
    .Q_N(_0037_),
    .Q(\vga.count_v[0] ));
 sg13g2_dfrbp_1 \vga.count_v[1]$_SDFFE_PN1N_  (.CLK(clknet_5_15__leaf_clk),
    .RESET_B(net214),
    .D(_0134_),
    .Q_N(_0080_),
    .Q(\vga.count_v[1] ));
 sg13g2_dfrbp_1 \vga.count_v[2]$_SDFFE_PN1N_  (.CLK(clknet_5_3__leaf_clk),
    .RESET_B(net215),
    .D(_0135_),
    .Q_N(_0038_),
    .Q(\vga.count_v[2] ));
 sg13g2_dfrbp_1 \vga.count_v[3]$_SDFFE_PN1N_  (.CLK(clknet_5_3__leaf_clk),
    .RESET_B(net216),
    .D(_0136_),
    .Q_N(_0039_),
    .Q(\vga.count_v[3] ));
 sg13g2_dfrbp_1 \vga.count_v[4]$_SDFFE_PN1N_  (.CLK(clknet_5_3__leaf_clk),
    .RESET_B(net217),
    .D(_0137_),
    .Q_N(_0040_),
    .Q(\vga.count_v[4] ));
 sg13g2_dfrbp_1 \vga.count_v[5]$_SDFFE_PN1N_  (.CLK(clknet_5_24__leaf_clk),
    .RESET_B(net218),
    .D(_0138_),
    .Q_N(_0041_),
    .Q(\vga.count_v[5] ));
 sg13g2_dfrbp_1 \vga.count_v[6]$_SDFFE_PN1N_  (.CLK(clknet_5_18__leaf_clk),
    .RESET_B(net219),
    .D(_0139_),
    .Q_N(_0042_),
    .Q(\vga.count_v[6] ));
 sg13g2_dfrbp_1 \vga.count_v[7]$_SDFFE_PN1N_  (.CLK(clknet_5_24__leaf_clk),
    .RESET_B(net220),
    .D(_0140_),
    .Q_N(_0043_),
    .Q(\vga.count_v[7] ));
 sg13g2_dfrbp_1 \vga.count_v[8]$_SDFFE_PN1N_  (.CLK(clknet_5_1__leaf_clk),
    .RESET_B(net221),
    .D(_0141_),
    .Q_N(_0044_),
    .Q(\vga.count_v[8] ));
 sg13g2_dfrbp_1 \vga.count_v[9]$_SDFFE_PN0N_  (.CLK(clknet_5_15__leaf_clk),
    .RESET_B(net222),
    .D(_0142_),
    .Q_N(_0065_),
    .Q(\vga.count_v[9] ));
 sg13g2_dfrbp_1 \vga.hs_out$_SDFF_PP0_  (.CLK(clknet_5_21__leaf_clk),
    .RESET_B(net223),
    .D(_0143_),
    .Q_N(hs),
    .Q(\vga.hs_out ));
 sg13g2_dfrbp_1 \vga.interval_counter[0]$_SDFF_PP0_  (.CLK(clknet_5_29__leaf_clk),
    .RESET_B(net224),
    .D(_0144_),
    .Q_N(_0083_),
    .Q(\vga.interval_counter[0] ));
 sg13g2_dfrbp_1 \vga.interval_counter[10]$_SDFF_PP0_  (.CLK(clknet_5_29__leaf_clk),
    .RESET_B(net225),
    .D(_0145_),
    .Q_N(_2188_),
    .Q(\vga.interval_counter[10] ));
 sg13g2_dfrbp_1 \vga.interval_counter[11]$_SDFF_PP0_  (.CLK(clknet_5_23__leaf_clk),
    .RESET_B(net226),
    .D(_0146_),
    .Q_N(_2187_),
    .Q(\vga.interval_counter[11] ));
 sg13g2_dfrbp_1 \vga.interval_counter[12]$_SDFF_PP0_  (.CLK(clknet_5_29__leaf_clk),
    .RESET_B(net227),
    .D(_0147_),
    .Q_N(_2186_),
    .Q(\vga.interval_counter[12] ));
 sg13g2_dfrbp_1 \vga.interval_counter[13]$_SDFF_PP0_  (.CLK(clknet_5_29__leaf_clk),
    .RESET_B(net228),
    .D(_0148_),
    .Q_N(_2185_),
    .Q(\vga.interval_counter[13] ));
 sg13g2_dfrbp_1 \vga.interval_counter[14]$_SDFF_PP0_  (.CLK(clknet_5_31__leaf_clk),
    .RESET_B(net229),
    .D(_0149_),
    .Q_N(_2184_),
    .Q(\vga.interval_counter[14] ));
 sg13g2_dfrbp_1 \vga.interval_counter[15]$_SDFF_PP0_  (.CLK(clknet_5_31__leaf_clk),
    .RESET_B(net230),
    .D(_0150_),
    .Q_N(_2183_),
    .Q(\vga.interval_counter[15] ));
 sg13g2_dfrbp_1 \vga.interval_counter[16]$_SDFF_PP0_  (.CLK(clknet_5_28__leaf_clk),
    .RESET_B(net231),
    .D(_0151_),
    .Q_N(_2182_),
    .Q(\vga.interval_counter[16] ));
 sg13g2_dfrbp_1 \vga.interval_counter[17]$_SDFF_PP0_  (.CLK(clknet_5_28__leaf_clk),
    .RESET_B(net232),
    .D(_0152_),
    .Q_N(_2181_),
    .Q(\vga.interval_counter[17] ));
 sg13g2_dfrbp_1 \vga.interval_counter[18]$_SDFF_PP0_  (.CLK(clknet_5_28__leaf_clk),
    .RESET_B(net233),
    .D(_0153_),
    .Q_N(_2180_),
    .Q(\vga.interval_counter[18] ));
 sg13g2_dfrbp_1 \vga.interval_counter[19]$_SDFF_PP0_  (.CLK(clknet_5_28__leaf_clk),
    .RESET_B(net234),
    .D(_0154_),
    .Q_N(_2179_),
    .Q(\vga.interval_counter[19] ));
 sg13g2_dfrbp_1 \vga.interval_counter[1]$_SDFF_PP0_  (.CLK(clknet_5_24__leaf_clk),
    .RESET_B(net235),
    .D(_0155_),
    .Q_N(_2178_),
    .Q(\vga.interval_counter[1] ));
 sg13g2_dfrbp_1 \vga.interval_counter[20]$_SDFF_PP0_  (.CLK(clknet_5_30__leaf_clk),
    .RESET_B(net236),
    .D(_0156_),
    .Q_N(_2177_),
    .Q(\vga.interval_counter[20] ));
 sg13g2_dfrbp_1 \vga.interval_counter[21]$_SDFF_PP0_  (.CLK(clknet_5_30__leaf_clk),
    .RESET_B(net237),
    .D(_0157_),
    .Q_N(_2176_),
    .Q(\vga.interval_counter[21] ));
 sg13g2_dfrbp_1 \vga.interval_counter[22]$_SDFF_PP0_  (.CLK(clknet_5_31__leaf_clk),
    .RESET_B(net238),
    .D(_0158_),
    .Q_N(_2175_),
    .Q(\vga.interval_counter[22] ));
 sg13g2_dfrbp_1 \vga.interval_counter[23]$_SDFF_PP0_  (.CLK(clknet_5_31__leaf_clk),
    .RESET_B(net239),
    .D(_0159_),
    .Q_N(_2174_),
    .Q(\vga.interval_counter[23] ));
 sg13g2_dfrbp_1 \vga.interval_counter[24]$_SDFF_PP0_  (.CLK(clknet_5_30__leaf_clk),
    .RESET_B(net240),
    .D(_0160_),
    .Q_N(_2173_),
    .Q(\vga.interval_counter[24] ));
 sg13g2_dfrbp_1 \vga.interval_counter[2]$_SDFF_PP0_  (.CLK(clknet_5_25__leaf_clk),
    .RESET_B(net241),
    .D(_0161_),
    .Q_N(_2172_),
    .Q(\vga.interval_counter[2] ));
 sg13g2_dfrbp_1 \vga.interval_counter[3]$_SDFF_PP0_  (.CLK(clknet_5_24__leaf_clk),
    .RESET_B(net242),
    .D(_0162_),
    .Q_N(_2171_),
    .Q(\vga.interval_counter[3] ));
 sg13g2_dfrbp_1 \vga.interval_counter[4]$_SDFF_PP0_  (.CLK(clknet_5_28__leaf_clk),
    .RESET_B(net243),
    .D(_0163_),
    .Q_N(_2170_),
    .Q(\vga.interval_counter[4] ));
 sg13g2_dfrbp_1 \vga.interval_counter[5]$_SDFF_PP0_  (.CLK(clknet_5_18__leaf_clk),
    .RESET_B(net244),
    .D(_0164_),
    .Q_N(_2169_),
    .Q(\vga.interval_counter[5] ));
 sg13g2_dfrbp_1 \vga.interval_counter[6]$_SDFF_PP0_  (.CLK(clknet_5_22__leaf_clk),
    .RESET_B(net245),
    .D(_0165_),
    .Q_N(_2168_),
    .Q(\vga.interval_counter[6] ));
 sg13g2_dfrbp_1 \vga.interval_counter[7]$_SDFF_PP0_  (.CLK(clknet_5_22__leaf_clk),
    .RESET_B(net246),
    .D(_0166_),
    .Q_N(_2167_),
    .Q(\vga.interval_counter[7] ));
 sg13g2_dfrbp_1 \vga.interval_counter[8]$_SDFF_PP0_  (.CLK(clknet_5_22__leaf_clk),
    .RESET_B(net247),
    .D(_0167_),
    .Q_N(_2166_),
    .Q(\vga.interval_counter[8] ));
 sg13g2_dfrbp_1 \vga.interval_counter[9]$_SDFF_PP0_  (.CLK(clknet_5_22__leaf_clk),
    .RESET_B(net248),
    .D(_0168_),
    .Q_N(_2165_),
    .Q(\vga.interval_counter[9] ));
 sg13g2_dfrbp_1 \vga.left_down_1d$_DFFE_PN_  (.CLK(clknet_5_30__leaf_clk),
    .RESET_B(net249),
    .D(_0169_),
    .Q_N(_2164_),
    .Q(\vga.left_down_1d ));
 sg13g2_dfrbp_1 \vga.left_down_pressed$_SDFF_PP0_  (.CLK(clknet_5_27__leaf_clk),
    .RESET_B(net250),
    .D(_0170_),
    .Q_N(_2163_),
    .Q(\vga.left_down_pressed ));
 sg13g2_dfrbp_1 \vga.left_up_1d$_DFFE_PN_  (.CLK(clknet_5_30__leaf_clk),
    .RESET_B(net251),
    .D(_0171_),
    .Q_N(_2162_),
    .Q(\vga.left_up_1d ));
 sg13g2_dfrbp_1 \vga.left_up_pressed$_SDFF_PP0_  (.CLK(clknet_5_27__leaf_clk),
    .RESET_B(net252),
    .D(_0172_),
    .Q_N(_2161_),
    .Q(\vga.left_up_pressed ));
 sg13g2_dfrbp_1 \vga.paddle_l_pos_v[0]$_SDFFE_PN1P_  (.CLK(clknet_5_10__leaf_clk),
    .RESET_B(net253),
    .D(_0173_),
    .Q_N(_0082_),
    .Q(\vga.paddle_l_pos_v[0] ));
 sg13g2_dfrbp_1 \vga.paddle_l_pos_v[1]$_SDFFE_PN1P_  (.CLK(clknet_5_11__leaf_clk),
    .RESET_B(net254),
    .D(_0174_),
    .Q_N(_2160_),
    .Q(\vga.paddle_l_pos_v[1] ));
 sg13g2_dfrbp_1 \vga.paddle_l_pos_v[2]$_SDFFE_PN1P_  (.CLK(clknet_5_10__leaf_clk),
    .RESET_B(net255),
    .D(_0175_),
    .Q_N(_0060_),
    .Q(\vga.paddle_l_pos_v[2] ));
 sg13g2_dfrbp_1 \vga.paddle_l_pos_v[3]$_SDFFE_PN1P_  (.CLK(clknet_5_10__leaf_clk),
    .RESET_B(net256),
    .D(_0176_),
    .Q_N(_2159_),
    .Q(\vga.paddle_l_pos_v[3] ));
 sg13g2_dfrbp_1 \vga.paddle_l_pos_v[4]$_SDFFE_PN0P_  (.CLK(clknet_5_10__leaf_clk),
    .RESET_B(net257),
    .D(_0177_),
    .Q_N(_0059_),
    .Q(\vga.paddle_l_pos_v[4] ));
 sg13g2_dfrbp_1 \vga.paddle_l_pos_v[5]$_SDFFE_PN1P_  (.CLK(clknet_5_10__leaf_clk),
    .RESET_B(net258),
    .D(_0178_),
    .Q_N(_0077_),
    .Q(\vga.paddle_l_pos_v[5] ));
 sg13g2_dfrbp_1 \vga.paddle_l_pos_v[6]$_SDFFE_PN1P_  (.CLK(clknet_5_14__leaf_clk),
    .RESET_B(net259),
    .D(_0179_),
    .Q_N(_0079_),
    .Q(\vga.paddle_l_pos_v[6] ));
 sg13g2_dfrbp_1 \vga.paddle_l_pos_v[7]$_SDFFE_PN1P_  (.CLK(clknet_5_14__leaf_clk),
    .RESET_B(net260),
    .D(_0180_),
    .Q_N(_0078_),
    .Q(\vga.paddle_l_pos_v[7] ));
 sg13g2_dfrbp_1 \vga.paddle_l_pos_v[8]$_SDFFE_PN0P_  (.CLK(clknet_5_15__leaf_clk),
    .RESET_B(net261),
    .D(_0181_),
    .Q_N(_0076_),
    .Q(\vga.paddle_l_pos_v[8] ));
 sg13g2_dfrbp_1 \vga.paddle_r_pos_v[0]$_SDFFE_PN1P_  (.CLK(clknet_5_2__leaf_clk),
    .RESET_B(net262),
    .D(_0182_),
    .Q_N(_0081_),
    .Q(\vga.paddle_r_pos_v[0] ));
 sg13g2_dfrbp_1 \vga.paddle_r_pos_v[1]$_SDFFE_PN1P_  (.CLK(clknet_5_2__leaf_clk),
    .RESET_B(net263),
    .D(_0183_),
    .Q_N(_2158_),
    .Q(\vga.paddle_r_pos_v[1] ));
 sg13g2_dfrbp_1 \vga.paddle_r_pos_v[2]$_SDFFE_PN1P_  (.CLK(clknet_5_2__leaf_clk),
    .RESET_B(net264),
    .D(_0184_),
    .Q_N(_0062_),
    .Q(\vga.paddle_r_pos_v[2] ));
 sg13g2_dfrbp_1 \vga.paddle_r_pos_v[3]$_SDFFE_PN1P_  (.CLK(clknet_5_26__leaf_clk),
    .RESET_B(net265),
    .D(_0185_),
    .Q_N(_2157_),
    .Q(\vga.paddle_r_pos_v[3] ));
 sg13g2_dfrbp_1 \vga.paddle_r_pos_v[4]$_SDFFE_PN0P_  (.CLK(clknet_5_26__leaf_clk),
    .RESET_B(net266),
    .D(_0186_),
    .Q_N(_0061_),
    .Q(\vga.paddle_r_pos_v[4] ));
 sg13g2_dfrbp_1 \vga.paddle_r_pos_v[5]$_SDFFE_PN1P_  (.CLK(clknet_5_26__leaf_clk),
    .RESET_B(net267),
    .D(_0187_),
    .Q_N(_0069_),
    .Q(\vga.paddle_r_pos_v[5] ));
 sg13g2_dfrbp_1 \vga.paddle_r_pos_v[6]$_SDFFE_PN1P_  (.CLK(clknet_5_26__leaf_clk),
    .RESET_B(net268),
    .D(_0188_),
    .Q_N(_0072_),
    .Q(\vga.paddle_r_pos_v[6] ));
 sg13g2_dfrbp_1 \vga.paddle_r_pos_v[7]$_SDFFE_PN1P_  (.CLK(clknet_5_26__leaf_clk),
    .RESET_B(net269),
    .D(_0189_),
    .Q_N(_0070_),
    .Q(\vga.paddle_r_pos_v[7] ));
 sg13g2_dfrbp_1 \vga.paddle_r_pos_v[8]$_SDFFE_PN0P_  (.CLK(clknet_5_27__leaf_clk),
    .RESET_B(net270),
    .D(_0190_),
    .Q_N(_0068_),
    .Q(\vga.paddle_r_pos_v[8] ));
 sg13g2_dfrbp_1 \vga.red$_SDFF_PP0_  (.CLK(clknet_5_21__leaf_clk),
    .RESET_B(net271),
    .D(_0191_),
    .Q_N(_2156_),
    .Q(g0));
 sg13g2_dfrbp_1 \vga.right_down_1d$_DFFE_PN_  (.CLK(clknet_5_25__leaf_clk),
    .RESET_B(net272),
    .D(_0192_),
    .Q_N(_2155_),
    .Q(\vga.right_down_1d ));
 sg13g2_dfrbp_1 \vga.right_down_pressed$_SDFF_PP0_  (.CLK(clknet_5_27__leaf_clk),
    .RESET_B(net273),
    .D(_0193_),
    .Q_N(_2154_),
    .Q(\vga.right_down_pressed ));
 sg13g2_dfrbp_1 \vga.right_up_1d$_DFFE_PN_  (.CLK(clknet_5_25__leaf_clk),
    .RESET_B(net274),
    .D(_0194_),
    .Q_N(_2153_),
    .Q(\vga.right_up_1d ));
 sg13g2_dfrbp_1 \vga.right_up_pressed$_SDFF_PP0_  (.CLK(clknet_5_25__leaf_clk),
    .RESET_B(net275),
    .D(_0195_),
    .Q_N(_2152_),
    .Q(\vga.right_up_pressed ));
 sg13g2_dfrbp_1 \vga.score_l[0]$_SDFF_PN0_  (.CLK(clknet_5_19__leaf_clk),
    .RESET_B(net276),
    .D(net39),
    .Q_N(_2151_),
    .Q(\vga.score_l[0] ));
 sg13g2_dfrbp_1 \vga.score_l[1]$_SDFF_PN0_  (.CLK(clknet_5_18__leaf_clk),
    .RESET_B(net277),
    .D(_0197_),
    .Q_N(_2150_),
    .Q(\vga.score_l[1] ));
 sg13g2_dfrbp_1 \vga.score_l[2]$_SDFF_PN0_  (.CLK(clknet_5_19__leaf_clk),
    .RESET_B(net278),
    .D(net34),
    .Q_N(_2149_),
    .Q(\vga.score_l[2] ));
 sg13g2_dfrbp_1 \vga.score_l[3]$_SDFF_PN0_  (.CLK(clknet_5_19__leaf_clk),
    .RESET_B(net279),
    .D(net33),
    .Q_N(_2148_),
    .Q(\vga.score_l[3] ));
 sg13g2_dfrbp_1 \vga.score_l[4]$_SDFF_PN0_  (.CLK(clknet_5_16__leaf_clk),
    .RESET_B(net280),
    .D(net31),
    .Q_N(_2147_),
    .Q(\vga.score_l[4] ));
 sg13g2_dfrbp_1 \vga.score_l_ten_enable$_SDFF_PN0_  (.CLK(clknet_5_6__leaf_clk),
    .RESET_B(net281),
    .D(_0201_),
    .Q_N(_2146_),
    .Q(\vga.score_l_ten_enable ));
 sg13g2_dfrbp_1 \vga.score_l_unit_pixels[0]$_DFFE_PP_  (.CLK(clknet_5_4__leaf_clk),
    .RESET_B(net282),
    .D(_0202_),
    .Q_N(_2145_),
    .Q(\vga.score_l_unit_pixels[0] ));
 sg13g2_dfrbp_1 \vga.score_l_unit_pixels[1]$_DFFE_PP_  (.CLK(clknet_5_4__leaf_clk),
    .RESET_B(net283),
    .D(_0203_),
    .Q_N(_2144_),
    .Q(\vga.score_l_unit_pixels[1] ));
 sg13g2_dfrbp_1 \vga.score_l_unit_pixels[2]$_DFFE_PP_  (.CLK(clknet_5_5__leaf_clk),
    .RESET_B(net284),
    .D(_0204_),
    .Q_N(_2143_),
    .Q(\vga.score_l_unit_pixels[2] ));
 sg13g2_dfrbp_1 \vga.score_r[0]$_SDFF_PN0_  (.CLK(clknet_5_20__leaf_clk),
    .RESET_B(net285),
    .D(_0205_),
    .Q_N(_2142_),
    .Q(\vga.score_r[0] ));
 sg13g2_dfrbp_1 \vga.score_r[1]$_SDFF_PN0_  (.CLK(clknet_5_20__leaf_clk),
    .RESET_B(net286),
    .D(_0206_),
    .Q_N(_2141_),
    .Q(\vga.score_r[1] ));
 sg13g2_dfrbp_1 \vga.score_r[2]$_SDFF_PN0_  (.CLK(clknet_5_23__leaf_clk),
    .RESET_B(net287),
    .D(net36),
    .Q_N(_2140_),
    .Q(\vga.score_r[2] ));
 sg13g2_dfrbp_1 \vga.score_r[3]$_SDFF_PN0_  (.CLK(clknet_5_7__leaf_clk),
    .RESET_B(net288),
    .D(_0208_),
    .Q_N(_2139_),
    .Q(\vga.score_r[3] ));
 sg13g2_dfrbp_1 \vga.score_r[4]$_SDFF_PN0_  (.CLK(clknet_5_20__leaf_clk),
    .RESET_B(net289),
    .D(_0209_),
    .Q_N(_2138_),
    .Q(\vga.score_r[4] ));
 sg13g2_dfrbp_1 \vga.score_r_ten_enable$_SDFF_PN0_  (.CLK(clknet_5_1__leaf_clk),
    .RESET_B(net290),
    .D(_0210_),
    .Q_N(_2137_),
    .Q(\vga.score_r_ten_enable ));
 sg13g2_dfrbp_1 \vga.score_r_unit_pixels[0]$_DFFE_PP_  (.CLK(clknet_5_0__leaf_clk),
    .RESET_B(net291),
    .D(_0211_),
    .Q_N(_2136_),
    .Q(\vga.score_r_unit_pixels[0] ));
 sg13g2_dfrbp_1 \vga.score_r_unit_pixels[1]$_DFFE_PP_  (.CLK(clknet_5_0__leaf_clk),
    .RESET_B(net292),
    .D(_0212_),
    .Q_N(_2135_),
    .Q(\vga.score_r_unit_pixels[1] ));
 sg13g2_dfrbp_1 \vga.score_r_unit_pixels[2]$_DFFE_PP_  (.CLK(clknet_5_6__leaf_clk),
    .RESET_B(net293),
    .D(_0213_),
    .Q_N(_2134_),
    .Q(\vga.score_r_unit_pixels[2] ));
 sg13g2_dfrbp_1 \vga.speed_lsb_1d$_SDFF_PN0_  (.CLK(clknet_5_23__leaf_clk),
    .RESET_B(net294),
    .D(_0214_),
    .Q_N(_2133_),
    .Q(\vga.speed_lsb_1d ));
 sg13g2_dfrbp_1 \vga.speed_msb_1d$_SDFF_PN0_  (.CLK(clknet_5_23__leaf_clk),
    .RESET_B(net295),
    .D(_0215_),
    .Q_N(_2132_),
    .Q(\vga.speed_msb_1d ));
 sg13g2_dfrbp_1 \vga.vs_out$_SDFFE_PN0P_  (.CLK(clknet_5_1__leaf_clk),
    .RESET_B(net296),
    .D(_0216_),
    .Q_N(\vga.vs ),
    .Q(\vga.vs_out ));
 sg13g2_buf_1 input1 (.A(ui_in[0]),
    .X(net1));
 sg13g2_buf_1 input2 (.A(ui_in[1]),
    .X(net2));
 sg13g2_buf_1 input3 (.A(ui_in[2]),
    .X(net3));
 sg13g2_buf_1 input4 (.A(ui_in[3]),
    .X(net4));
 sg13g2_buf_1 input5 (.A(ui_in[5]),
    .X(net5));
 sg13g2_buf_1 output6 (.A(net6),
    .X(uio_oe[0]));
 sg13g2_buf_1 output7 (.A(net7),
    .X(uio_oe[1]));
 sg13g2_buf_1 output8 (.A(net8),
    .X(uio_oe[2]));
 sg13g2_buf_1 output9 (.A(net9),
    .X(uio_oe[3]));
 sg13g2_buf_1 output10 (.A(net10),
    .X(uio_oe[4]));
 sg13g2_buf_1 output11 (.A(net11),
    .X(uio_oe[5]));
 sg13g2_buf_1 output12 (.A(net12),
    .X(uio_oe[6]));
 sg13g2_buf_1 output13 (.A(net13),
    .X(uio_oe[7]));
 sg13g2_buf_1 output14 (.A(net14),
    .X(uio_out[0]));
 sg13g2_buf_1 output15 (.A(net15),
    .X(uio_out[1]));
 sg13g2_buf_1 output16 (.A(net16),
    .X(uio_out[2]));
 sg13g2_buf_1 output17 (.A(net17),
    .X(uio_out[3]));
 sg13g2_buf_1 output18 (.A(net18),
    .X(uio_out[4]));
 sg13g2_buf_1 output19 (.A(net19),
    .X(uio_out[5]));
 sg13g2_buf_1 output20 (.A(net20),
    .X(uo_out[0]));
 sg13g2_buf_1 output21 (.A(net21),
    .X(uo_out[1]));
 sg13g2_buf_1 output22 (.A(net22),
    .X(uo_out[2]));
 sg13g2_buf_1 output23 (.A(net23),
    .X(uo_out[3]));
 sg13g2_buf_1 output24 (.A(net24),
    .X(uo_out[4]));
 sg13g2_buf_1 output25 (.A(net25),
    .X(uo_out[5]));
 sg13g2_buf_1 output26 (.A(net26),
    .X(uo_out[6]));
 sg13g2_buf_1 output27 (.A(net27),
    .X(uo_out[7]));
 sg13g2_buf_2 fanout28 (.A(_1096_),
    .X(net28));
 sg13g2_buf_2 fanout29 (.A(_1076_),
    .X(net29));
 sg13g2_buf_2 fanout30 (.A(_1073_),
    .X(net30));
 sg13g2_buf_2 fanout31 (.A(_0200_),
    .X(net31));
 sg13g2_buf_2 fanout32 (.A(_1056_),
    .X(net32));
 sg13g2_buf_2 fanout33 (.A(_0199_),
    .X(net33));
 sg13g2_buf_2 fanout34 (.A(_0198_),
    .X(net34));
 sg13g2_buf_2 fanout35 (.A(_2071_),
    .X(net35));
 sg13g2_buf_2 fanout36 (.A(_0207_),
    .X(net36));
 sg13g2_buf_2 fanout37 (.A(_2057_),
    .X(net37));
 sg13g2_buf_2 fanout38 (.A(_2023_),
    .X(net38));
 sg13g2_buf_2 fanout39 (.A(_0196_),
    .X(net39));
 sg13g2_buf_2 fanout40 (.A(_2069_),
    .X(net40));
 sg13g2_buf_2 fanout41 (.A(_2031_),
    .X(net41));
 sg13g2_buf_2 fanout42 (.A(_1329_),
    .X(net42));
 sg13g2_buf_2 fanout43 (.A(_0432_),
    .X(net43));
 sg13g2_buf_2 fanout44 (.A(_0408_),
    .X(net44));
 sg13g2_buf_2 fanout45 (.A(_1291_),
    .X(net45));
 sg13g2_buf_2 fanout46 (.A(_1057_),
    .X(net46));
 sg13g2_buf_2 fanout47 (.A(_0598_),
    .X(net47));
 sg13g2_buf_2 fanout48 (.A(_1309_),
    .X(net48));
 sg13g2_buf_2 fanout49 (.A(_1037_),
    .X(net49));
 sg13g2_buf_2 fanout50 (.A(_0319_),
    .X(net50));
 sg13g2_buf_2 fanout51 (.A(_1093_),
    .X(net51));
 sg13g2_buf_2 fanout52 (.A(_1054_),
    .X(net52));
 sg13g2_buf_2 fanout53 (.A(_1092_),
    .X(net53));
 sg13g2_buf_2 fanout54 (.A(_0968_),
    .X(net54));
 sg13g2_buf_2 fanout55 (.A(_0839_),
    .X(net55));
 sg13g2_buf_2 fanout56 (.A(_0562_),
    .X(net56));
 sg13g2_buf_2 fanout57 (.A(_0338_),
    .X(net57));
 sg13g2_buf_2 fanout58 (.A(_0327_),
    .X(net58));
 sg13g2_buf_2 fanout59 (.A(_0272_),
    .X(net59));
 sg13g2_buf_2 fanout60 (.A(_1889_),
    .X(net60));
 sg13g2_buf_2 fanout61 (.A(_1840_),
    .X(net61));
 sg13g2_buf_2 fanout62 (.A(_1817_),
    .X(net62));
 sg13g2_buf_2 fanout63 (.A(_1812_),
    .X(net63));
 sg13g2_buf_2 fanout64 (.A(_1647_),
    .X(net64));
 sg13g2_buf_2 fanout65 (.A(_1551_),
    .X(net65));
 sg13g2_buf_2 fanout66 (.A(_1527_),
    .X(net66));
 sg13g2_buf_2 fanout67 (.A(_1246_),
    .X(net67));
 sg13g2_buf_2 fanout68 (.A(_1184_),
    .X(net68));
 sg13g2_buf_2 fanout69 (.A(_1053_),
    .X(net69));
 sg13g2_buf_2 fanout70 (.A(_0726_),
    .X(net70));
 sg13g2_buf_2 fanout71 (.A(_0674_),
    .X(net71));
 sg13g2_buf_2 fanout72 (.A(_0623_),
    .X(net72));
 sg13g2_buf_2 fanout73 (.A(_0617_),
    .X(net73));
 sg13g2_buf_2 fanout74 (.A(_0610_),
    .X(net74));
 sg13g2_buf_2 fanout75 (.A(_0605_),
    .X(net75));
 sg13g2_buf_2 fanout76 (.A(_0515_),
    .X(net76));
 sg13g2_buf_2 fanout77 (.A(_0488_),
    .X(net77));
 sg13g2_buf_2 fanout78 (.A(_0486_),
    .X(net78));
 sg13g2_buf_2 fanout79 (.A(_0473_),
    .X(net79));
 sg13g2_buf_2 fanout80 (.A(_0467_),
    .X(net80));
 sg13g2_buf_2 fanout81 (.A(_0466_),
    .X(net81));
 sg13g2_buf_2 fanout82 (.A(_0363_),
    .X(net82));
 sg13g2_buf_2 fanout83 (.A(_0362_),
    .X(net83));
 sg13g2_buf_2 fanout84 (.A(_0348_),
    .X(net84));
 sg13g2_buf_2 fanout85 (.A(_0340_),
    .X(net85));
 sg13g2_buf_2 fanout86 (.A(_0278_),
    .X(net86));
 sg13g2_buf_2 fanout87 (.A(_0273_),
    .X(net87));
 sg13g2_buf_2 fanout88 (.A(_0271_),
    .X(net88));
 sg13g2_buf_2 fanout89 (.A(_0254_),
    .X(net89));
 sg13g2_buf_2 fanout90 (.A(_0248_),
    .X(net90));
 sg13g2_buf_2 fanout91 (.A(_0246_),
    .X(net91));
 sg13g2_buf_2 fanout92 (.A(_2123_),
    .X(net92));
 sg13g2_buf_2 fanout93 (.A(_2076_),
    .X(net93));
 sg13g2_buf_2 fanout94 (.A(_2061_),
    .X(net94));
 sg13g2_buf_2 fanout95 (.A(_1863_),
    .X(net95));
 sg13g2_buf_2 fanout96 (.A(_1861_),
    .X(net96));
 sg13g2_buf_2 fanout97 (.A(_1842_),
    .X(net97));
 sg13g2_buf_2 fanout98 (.A(_1823_),
    .X(net98));
 sg13g2_buf_2 fanout99 (.A(_1821_),
    .X(net99));
 sg13g2_buf_2 fanout100 (.A(_1810_),
    .X(net100));
 sg13g2_buf_2 fanout101 (.A(_1772_),
    .X(net101));
 sg13g2_buf_2 fanout102 (.A(_1683_),
    .X(net102));
 sg13g2_buf_2 fanout103 (.A(_1676_),
    .X(net103));
 sg13g2_buf_2 fanout104 (.A(_1666_),
    .X(net104));
 sg13g2_buf_2 fanout105 (.A(_1658_),
    .X(net105));
 sg13g2_buf_2 fanout106 (.A(_1656_),
    .X(net106));
 sg13g2_buf_2 fanout107 (.A(_1655_),
    .X(net107));
 sg13g2_buf_2 fanout108 (.A(_1653_),
    .X(net108));
 sg13g2_buf_2 fanout109 (.A(_1646_),
    .X(net109));
 sg13g2_buf_2 fanout110 (.A(_1635_),
    .X(net110));
 sg13g2_buf_2 fanout111 (.A(_1602_),
    .X(net111));
 sg13g2_buf_2 fanout112 (.A(_1576_),
    .X(net112));
 sg13g2_buf_2 fanout113 (.A(_1549_),
    .X(net113));
 sg13g2_buf_2 fanout114 (.A(_1532_),
    .X(net114));
 sg13g2_buf_2 fanout115 (.A(_1523_),
    .X(net115));
 sg13g2_buf_2 fanout116 (.A(_1516_),
    .X(net116));
 sg13g2_buf_2 fanout117 (.A(_1063_),
    .X(net117));
 sg13g2_buf_2 fanout118 (.A(_0672_),
    .X(net118));
 sg13g2_buf_2 fanout119 (.A(_0611_),
    .X(net119));
 sg13g2_buf_2 fanout120 (.A(_0596_),
    .X(net120));
 sg13g2_buf_2 fanout121 (.A(_0592_),
    .X(net121));
 sg13g2_buf_2 fanout122 (.A(_0354_),
    .X(net122));
 sg13g2_buf_2 fanout123 (.A(_0353_),
    .X(net123));
 sg13g2_buf_2 fanout124 (.A(_0351_),
    .X(net124));
 sg13g2_buf_2 fanout125 (.A(_2025_),
    .X(net125));
 sg13g2_buf_2 fanout126 (.A(_2013_),
    .X(net126));
 sg13g2_buf_2 fanout127 (.A(_1998_),
    .X(net127));
 sg13g2_buf_2 fanout128 (.A(_1984_),
    .X(net128));
 sg13g2_buf_2 fanout129 (.A(_1914_),
    .X(net129));
 sg13g2_buf_2 fanout130 (.A(_1850_),
    .X(net130));
 sg13g2_buf_2 fanout131 (.A(_1833_),
    .X(net131));
 sg13g2_buf_2 fanout132 (.A(_1822_),
    .X(net132));
 sg13g2_buf_2 fanout133 (.A(_1808_),
    .X(net133));
 sg13g2_buf_2 fanout134 (.A(_1801_),
    .X(net134));
 sg13g2_buf_2 fanout135 (.A(_1768_),
    .X(net135));
 sg13g2_buf_2 fanout136 (.A(_1741_),
    .X(net136));
 sg13g2_buf_2 fanout137 (.A(_1738_),
    .X(net137));
 sg13g2_buf_2 fanout138 (.A(_1731_),
    .X(net138));
 sg13g2_buf_2 fanout139 (.A(_1659_),
    .X(net139));
 sg13g2_buf_2 fanout140 (.A(_1619_),
    .X(net140));
 sg13g2_buf_2 fanout141 (.A(_1583_),
    .X(net141));
 sg13g2_buf_2 fanout142 (.A(_1582_),
    .X(net142));
 sg13g2_buf_2 fanout143 (.A(_1530_),
    .X(net143));
 sg13g2_buf_2 fanout144 (.A(_1522_),
    .X(net144));
 sg13g2_buf_2 fanout145 (.A(_1518_),
    .X(net145));
 sg13g2_buf_2 fanout146 (.A(_1511_),
    .X(net146));
 sg13g2_buf_2 fanout147 (.A(_1507_),
    .X(net147));
 sg13g2_buf_2 fanout148 (.A(_1505_),
    .X(net148));
 sg13g2_tielo _4332__149 (.L_LO(net149));
 sg13g2_tielo _4333__150 (.L_LO(net150));
 sg13g2_tiehi _4296__152 (.L_HI(net152));
 sg13g2_tiehi _4297__153 (.L_HI(net153));
 sg13g2_tiehi _4298__154 (.L_HI(net154));
 sg13g2_tiehi _4299__155 (.L_HI(net155));
 sg13g2_tiehi _4300__156 (.L_HI(net156));
 sg13g2_tiehi _4301__157 (.L_HI(net157));
 sg13g2_tiehi _4302__158 (.L_HI(net158));
 sg13g2_tiehi _4303__159 (.L_HI(net159));
 sg13g2_tiehi _4304__160 (.L_HI(net160));
 sg13g2_tiehi _4305__161 (.L_HI(net161));
 sg13g2_tiehi _4306__162 (.L_HI(net162));
 sg13g2_tiehi _4307__163 (.L_HI(net163));
 sg13g2_tiehi _4308__164 (.L_HI(net164));
 sg13g2_tiehi _4309__165 (.L_HI(net165));
 sg13g2_tiehi _4310__166 (.L_HI(net166));
 sg13g2_tiehi _4311__167 (.L_HI(net167));
 sg13g2_tiehi _4312__168 (.L_HI(net168));
 sg13g2_tiehi _4313__169 (.L_HI(net169));
 sg13g2_tiehi _4314__170 (.L_HI(net170));
 sg13g2_tiehi _4315__171 (.L_HI(net171));
 sg13g2_tiehi _4316__172 (.L_HI(net172));
 sg13g2_tiehi \vga.ball_angle[0]$_SDFFE_PN1P__173  (.L_HI(net173));
 sg13g2_tiehi \vga.ball_angle[1]$_SDFFE_PN0P__174  (.L_HI(net174));
 sg13g2_tiehi \vga.ball_angle[2]$_SDFFE_PN0P__175  (.L_HI(net175));
 sg13g2_tiehi \vga.ball_angle[3]$_SDFFE_PN1P__176  (.L_HI(net176));
 sg13g2_tiehi \vga.ball_motion_l$_SDFFE_PN1N__177  (.L_HI(net177));
 sg13g2_tiehi \vga.ball_pos_h[0]$_SDFFE_PN1P__178  (.L_HI(net178));
 sg13g2_tiehi \vga.ball_pos_h[1]$_SDFFE_PN1P__179  (.L_HI(net179));
 sg13g2_tiehi \vga.ball_pos_h[2]$_SDFFE_PN1P__180  (.L_HI(net180));
 sg13g2_tiehi \vga.ball_pos_h[3]$_SDFFE_PN1P__181  (.L_HI(net181));
 sg13g2_tiehi \vga.ball_pos_h[4]$_SDFFE_PN0P__182  (.L_HI(net182));
 sg13g2_tiehi \vga.ball_pos_h[5]$_SDFFE_PN1P__183  (.L_HI(net183));
 sg13g2_tiehi \vga.ball_pos_h[6]$_SDFFE_PN1P__184  (.L_HI(net184));
 sg13g2_tiehi \vga.ball_pos_h[7]$_SDFFE_PN0P__185  (.L_HI(net185));
 sg13g2_tiehi \vga.ball_pos_h[8]$_SDFFE_PN0P__186  (.L_HI(net186));
 sg13g2_tiehi \vga.ball_pos_h[9]$_SDFFE_PN1P__187  (.L_HI(net187));
 sg13g2_tiehi \vga.ball_pos_v[0]$_SDFFE_PN1P__188  (.L_HI(net188));
 sg13g2_tiehi \vga.ball_pos_v[1]$_SDFFE_PN1P__189  (.L_HI(net189));
 sg13g2_tiehi \vga.ball_pos_v[2]$_SDFFE_PN1P__190  (.L_HI(net190));
 sg13g2_tiehi \vga.ball_pos_v[3]$_SDFFE_PN1P__191  (.L_HI(net191));
 sg13g2_tiehi \vga.ball_pos_v[4]$_SDFFE_PN0P__192  (.L_HI(net192));
 sg13g2_tiehi \vga.ball_pos_v[5]$_SDFFE_PN1P__193  (.L_HI(net193));
 sg13g2_tiehi \vga.ball_pos_v[6]$_SDFFE_PN1P__194  (.L_HI(net194));
 sg13g2_tiehi \vga.ball_pos_v[7]$_SDFFE_PN1P__195  (.L_HI(net195));
 sg13g2_tiehi \vga.ball_pos_v[8]$_SDFFE_PN0P__196  (.L_HI(net196));
 sg13g2_tiehi \vga.ball_ratio[0]$_SDFFE_PN0P__197  (.L_HI(net197));
 sg13g2_tiehi \vga.ball_ratio[1]$_SDFFE_PN0P__198  (.L_HI(net198));
 sg13g2_tiehi \vga.ball_ratio[2]$_SDFFE_PN0P__199  (.L_HI(net199));
 sg13g2_tiehi \vga.blank_h$_SDFFE_PN1P__200  (.L_HI(net200));
 sg13g2_tiehi \vga.blank_v$_SDFFE_PN1P__201  (.L_HI(net201));
 sg13g2_tiehi \vga.blu$_SDFF_PN0__202  (.L_HI(net202));
 sg13g2_tiehi \vga.count_h[0]$_SDFF_PN1__203  (.L_HI(net203));
 sg13g2_tiehi \vga.count_h[1]$_SDFF_PN1__204  (.L_HI(net204));
 sg13g2_tiehi \vga.count_h[2]$_SDFF_PN1__205  (.L_HI(net205));
 sg13g2_tiehi \vga.count_h[3]$_SDFF_PN1__206  (.L_HI(net206));
 sg13g2_tiehi \vga.count_h[4]$_SDFF_PN1__207  (.L_HI(net207));
 sg13g2_tiehi \vga.count_h[5]$_SDFF_PN1__208  (.L_HI(net208));
 sg13g2_tiehi \vga.count_h[6]$_SDFF_PN1__209  (.L_HI(net209));
 sg13g2_tiehi \vga.count_h[7]$_SDFF_PN1__210  (.L_HI(net210));
 sg13g2_tiehi \vga.count_h[8]$_SDFF_PN1__211  (.L_HI(net211));
 sg13g2_tiehi \vga.count_h[9]$_SDFF_PN1__212  (.L_HI(net212));
 sg13g2_tiehi \vga.count_v[0]$_SDFFE_PN1N__213  (.L_HI(net213));
 sg13g2_tiehi \vga.count_v[1]$_SDFFE_PN1N__214  (.L_HI(net214));
 sg13g2_tiehi \vga.count_v[2]$_SDFFE_PN1N__215  (.L_HI(net215));
 sg13g2_tiehi \vga.count_v[3]$_SDFFE_PN1N__216  (.L_HI(net216));
 sg13g2_tiehi \vga.count_v[4]$_SDFFE_PN1N__217  (.L_HI(net217));
 sg13g2_tiehi \vga.count_v[5]$_SDFFE_PN1N__218  (.L_HI(net218));
 sg13g2_tiehi \vga.count_v[6]$_SDFFE_PN1N__219  (.L_HI(net219));
 sg13g2_tiehi \vga.count_v[7]$_SDFFE_PN1N__220  (.L_HI(net220));
 sg13g2_tiehi \vga.count_v[8]$_SDFFE_PN1N__221  (.L_HI(net221));
 sg13g2_tiehi \vga.count_v[9]$_SDFFE_PN0N__222  (.L_HI(net222));
 sg13g2_tiehi \vga.hs_out$_SDFF_PP0__223  (.L_HI(net223));
 sg13g2_tiehi \vga.interval_counter[0]$_SDFF_PP0__224  (.L_HI(net224));
 sg13g2_tiehi \vga.interval_counter[10]$_SDFF_PP0__225  (.L_HI(net225));
 sg13g2_tiehi \vga.interval_counter[11]$_SDFF_PP0__226  (.L_HI(net226));
 sg13g2_tiehi \vga.interval_counter[12]$_SDFF_PP0__227  (.L_HI(net227));
 sg13g2_tiehi \vga.interval_counter[13]$_SDFF_PP0__228  (.L_HI(net228));
 sg13g2_tiehi \vga.interval_counter[14]$_SDFF_PP0__229  (.L_HI(net229));
 sg13g2_tiehi \vga.interval_counter[15]$_SDFF_PP0__230  (.L_HI(net230));
 sg13g2_tiehi \vga.interval_counter[16]$_SDFF_PP0__231  (.L_HI(net231));
 sg13g2_tiehi \vga.interval_counter[17]$_SDFF_PP0__232  (.L_HI(net232));
 sg13g2_tiehi \vga.interval_counter[18]$_SDFF_PP0__233  (.L_HI(net233));
 sg13g2_tiehi \vga.interval_counter[19]$_SDFF_PP0__234  (.L_HI(net234));
 sg13g2_tiehi \vga.interval_counter[1]$_SDFF_PP0__235  (.L_HI(net235));
 sg13g2_tiehi \vga.interval_counter[20]$_SDFF_PP0__236  (.L_HI(net236));
 sg13g2_tiehi \vga.interval_counter[21]$_SDFF_PP0__237  (.L_HI(net237));
 sg13g2_tiehi \vga.interval_counter[22]$_SDFF_PP0__238  (.L_HI(net238));
 sg13g2_tiehi \vga.interval_counter[23]$_SDFF_PP0__239  (.L_HI(net239));
 sg13g2_tiehi \vga.interval_counter[24]$_SDFF_PP0__240  (.L_HI(net240));
 sg13g2_tiehi \vga.interval_counter[2]$_SDFF_PP0__241  (.L_HI(net241));
 sg13g2_tiehi \vga.interval_counter[3]$_SDFF_PP0__242  (.L_HI(net242));
 sg13g2_tiehi \vga.interval_counter[4]$_SDFF_PP0__243  (.L_HI(net243));
 sg13g2_tiehi \vga.interval_counter[5]$_SDFF_PP0__244  (.L_HI(net244));
 sg13g2_tiehi \vga.interval_counter[6]$_SDFF_PP0__245  (.L_HI(net245));
 sg13g2_tiehi \vga.interval_counter[7]$_SDFF_PP0__246  (.L_HI(net246));
 sg13g2_tiehi \vga.interval_counter[8]$_SDFF_PP0__247  (.L_HI(net247));
 sg13g2_tiehi \vga.interval_counter[9]$_SDFF_PP0__248  (.L_HI(net248));
 sg13g2_tiehi \vga.left_down_1d$_DFFE_PN__249  (.L_HI(net249));
 sg13g2_tiehi \vga.left_down_pressed$_SDFF_PP0__250  (.L_HI(net250));
 sg13g2_tiehi \vga.left_up_1d$_DFFE_PN__251  (.L_HI(net251));
 sg13g2_tiehi \vga.left_up_pressed$_SDFF_PP0__252  (.L_HI(net252));
 sg13g2_tiehi \vga.paddle_l_pos_v[0]$_SDFFE_PN1P__253  (.L_HI(net253));
 sg13g2_tiehi \vga.paddle_l_pos_v[1]$_SDFFE_PN1P__254  (.L_HI(net254));
 sg13g2_tiehi \vga.paddle_l_pos_v[2]$_SDFFE_PN1P__255  (.L_HI(net255));
 sg13g2_tiehi \vga.paddle_l_pos_v[3]$_SDFFE_PN1P__256  (.L_HI(net256));
 sg13g2_tiehi \vga.paddle_l_pos_v[4]$_SDFFE_PN0P__257  (.L_HI(net257));
 sg13g2_tiehi \vga.paddle_l_pos_v[5]$_SDFFE_PN1P__258  (.L_HI(net258));
 sg13g2_tiehi \vga.paddle_l_pos_v[6]$_SDFFE_PN1P__259  (.L_HI(net259));
 sg13g2_tiehi \vga.paddle_l_pos_v[7]$_SDFFE_PN1P__260  (.L_HI(net260));
 sg13g2_tiehi \vga.paddle_l_pos_v[8]$_SDFFE_PN0P__261  (.L_HI(net261));
 sg13g2_tiehi \vga.paddle_r_pos_v[0]$_SDFFE_PN1P__262  (.L_HI(net262));
 sg13g2_tiehi \vga.paddle_r_pos_v[1]$_SDFFE_PN1P__263  (.L_HI(net263));
 sg13g2_tiehi \vga.paddle_r_pos_v[2]$_SDFFE_PN1P__264  (.L_HI(net264));
 sg13g2_tiehi \vga.paddle_r_pos_v[3]$_SDFFE_PN1P__265  (.L_HI(net265));
 sg13g2_tiehi \vga.paddle_r_pos_v[4]$_SDFFE_PN0P__266  (.L_HI(net266));
 sg13g2_tiehi \vga.paddle_r_pos_v[5]$_SDFFE_PN1P__267  (.L_HI(net267));
 sg13g2_tiehi \vga.paddle_r_pos_v[6]$_SDFFE_PN1P__268  (.L_HI(net268));
 sg13g2_tiehi \vga.paddle_r_pos_v[7]$_SDFFE_PN1P__269  (.L_HI(net269));
 sg13g2_tiehi \vga.paddle_r_pos_v[8]$_SDFFE_PN0P__270  (.L_HI(net270));
 sg13g2_tiehi \vga.red$_SDFF_PP0__271  (.L_HI(net271));
 sg13g2_tiehi \vga.right_down_1d$_DFFE_PN__272  (.L_HI(net272));
 sg13g2_tiehi \vga.right_down_pressed$_SDFF_PP0__273  (.L_HI(net273));
 sg13g2_tiehi \vga.right_up_1d$_DFFE_PN__274  (.L_HI(net274));
 sg13g2_tiehi \vga.right_up_pressed$_SDFF_PP0__275  (.L_HI(net275));
 sg13g2_tiehi \vga.score_l[0]$_SDFF_PN0__276  (.L_HI(net276));
 sg13g2_tiehi \vga.score_l[1]$_SDFF_PN0__277  (.L_HI(net277));
 sg13g2_tiehi \vga.score_l[2]$_SDFF_PN0__278  (.L_HI(net278));
 sg13g2_tiehi \vga.score_l[3]$_SDFF_PN0__279  (.L_HI(net279));
 sg13g2_tiehi \vga.score_l[4]$_SDFF_PN0__280  (.L_HI(net280));
 sg13g2_tiehi \vga.score_l_ten_enable$_SDFF_PN0__281  (.L_HI(net281));
 sg13g2_tiehi \vga.score_l_unit_pixels[0]$_DFFE_PP__282  (.L_HI(net282));
 sg13g2_tiehi \vga.score_l_unit_pixels[1]$_DFFE_PP__283  (.L_HI(net283));
 sg13g2_tiehi \vga.score_l_unit_pixels[2]$_DFFE_PP__284  (.L_HI(net284));
 sg13g2_tiehi \vga.score_r[0]$_SDFF_PN0__285  (.L_HI(net285));
 sg13g2_tiehi \vga.score_r[1]$_SDFF_PN0__286  (.L_HI(net286));
 sg13g2_tiehi \vga.score_r[2]$_SDFF_PN0__287  (.L_HI(net287));
 sg13g2_tiehi \vga.score_r[3]$_SDFF_PN0__288  (.L_HI(net288));
 sg13g2_tiehi \vga.score_r[4]$_SDFF_PN0__289  (.L_HI(net289));
 sg13g2_tiehi \vga.score_r_ten_enable$_SDFF_PN0__290  (.L_HI(net290));
 sg13g2_tiehi \vga.score_r_unit_pixels[0]$_DFFE_PP__291  (.L_HI(net291));
 sg13g2_tiehi \vga.score_r_unit_pixels[1]$_DFFE_PP__292  (.L_HI(net292));
 sg13g2_tiehi \vga.score_r_unit_pixels[2]$_DFFE_PP__293  (.L_HI(net293));
 sg13g2_tiehi \vga.speed_lsb_1d$_SDFF_PN0__294  (.L_HI(net294));
 sg13g2_tiehi \vga.speed_msb_1d$_SDFF_PN0__295  (.L_HI(net295));
 sg13g2_tiehi \vga.vs_out$_SDFFE_PN0P__296  (.L_HI(net296));
 sg13g2_buf_2 clkbuf_4_0_0_clk (.A(clknet_0_clk),
    .X(clknet_4_0_0_clk));
 sg13g2_buf_2 clkbuf_4_1_0_clk (.A(clknet_0_clk),
    .X(clknet_4_1_0_clk));
 sg13g2_buf_2 clkbuf_4_2_0_clk (.A(clknet_0_clk),
    .X(clknet_4_2_0_clk));
 sg13g2_buf_2 clkbuf_4_3_0_clk (.A(clknet_0_clk),
    .X(clknet_4_3_0_clk));
 sg13g2_buf_2 clkbuf_4_4_0_clk (.A(clknet_0_clk),
    .X(clknet_4_4_0_clk));
 sg13g2_buf_2 clkbuf_4_5_0_clk (.A(clknet_0_clk),
    .X(clknet_4_5_0_clk));
 sg13g2_buf_2 clkbuf_4_6_0_clk (.A(clknet_0_clk),
    .X(clknet_4_6_0_clk));
 sg13g2_buf_2 clkbuf_4_7_0_clk (.A(clknet_0_clk),
    .X(clknet_4_7_0_clk));
 sg13g2_buf_2 clkbuf_4_8_0_clk (.A(clknet_0_clk),
    .X(clknet_4_8_0_clk));
 sg13g2_buf_2 clkbuf_4_9_0_clk (.A(clknet_0_clk),
    .X(clknet_4_9_0_clk));
 sg13g2_buf_2 clkbuf_4_10_0_clk (.A(clknet_0_clk),
    .X(clknet_4_10_0_clk));
 sg13g2_buf_2 clkbuf_4_11_0_clk (.A(clknet_0_clk),
    .X(clknet_4_11_0_clk));
 sg13g2_buf_2 clkbuf_4_12_0_clk (.A(clknet_0_clk),
    .X(clknet_4_12_0_clk));
 sg13g2_buf_2 clkbuf_4_13_0_clk (.A(clknet_0_clk),
    .X(clknet_4_13_0_clk));
 sg13g2_buf_2 clkbuf_4_14_0_clk (.A(clknet_0_clk),
    .X(clknet_4_14_0_clk));
 sg13g2_buf_2 clkbuf_4_15_0_clk (.A(clknet_0_clk),
    .X(clknet_4_15_0_clk));
 sg13g2_buf_1 clkbuf_5_0__f_clk (.A(clknet_4_0_0_clk),
    .X(clknet_5_0__leaf_clk));
 sg13g2_buf_1 clkbuf_5_1__f_clk (.A(clknet_4_0_0_clk),
    .X(clknet_5_1__leaf_clk));
 sg13g2_buf_1 clkbuf_5_2__f_clk (.A(clknet_4_1_0_clk),
    .X(clknet_5_2__leaf_clk));
 sg13g2_buf_1 clkbuf_5_3__f_clk (.A(clknet_4_1_0_clk),
    .X(clknet_5_3__leaf_clk));
 sg13g2_buf_1 clkbuf_5_4__f_clk (.A(clknet_4_2_0_clk),
    .X(clknet_5_4__leaf_clk));
 sg13g2_buf_1 clkbuf_5_5__f_clk (.A(clknet_4_2_0_clk),
    .X(clknet_5_5__leaf_clk));
 sg13g2_buf_1 clkbuf_5_6__f_clk (.A(clknet_4_3_0_clk),
    .X(clknet_5_6__leaf_clk));
 sg13g2_buf_1 clkbuf_5_7__f_clk (.A(clknet_4_3_0_clk),
    .X(clknet_5_7__leaf_clk));
 sg13g2_buf_1 clkbuf_5_8__f_clk (.A(clknet_4_4_0_clk),
    .X(clknet_5_8__leaf_clk));
 sg13g2_buf_1 clkbuf_5_9__f_clk (.A(clknet_4_4_0_clk),
    .X(clknet_5_9__leaf_clk));
 sg13g2_buf_1 clkbuf_5_10__f_clk (.A(clknet_4_5_0_clk),
    .X(clknet_5_10__leaf_clk));
 sg13g2_buf_1 clkbuf_5_11__f_clk (.A(clknet_4_5_0_clk),
    .X(clknet_5_11__leaf_clk));
 sg13g2_buf_1 clkbuf_5_12__f_clk (.A(clknet_4_6_0_clk),
    .X(clknet_5_12__leaf_clk));
 sg13g2_buf_1 clkbuf_5_13__f_clk (.A(clknet_4_6_0_clk),
    .X(clknet_5_13__leaf_clk));
 sg13g2_buf_1 clkbuf_5_14__f_clk (.A(clknet_4_7_0_clk),
    .X(clknet_5_14__leaf_clk));
 sg13g2_buf_1 clkbuf_5_15__f_clk (.A(clknet_4_7_0_clk),
    .X(clknet_5_15__leaf_clk));
 sg13g2_buf_1 clkbuf_5_16__f_clk (.A(clknet_4_8_0_clk),
    .X(clknet_5_16__leaf_clk));
 sg13g2_buf_1 clkbuf_5_17__f_clk (.A(clknet_4_8_0_clk),
    .X(clknet_5_17__leaf_clk));
 sg13g2_buf_1 clkbuf_5_18__f_clk (.A(clknet_4_9_0_clk),
    .X(clknet_5_18__leaf_clk));
 sg13g2_buf_1 clkbuf_5_19__f_clk (.A(clknet_4_9_0_clk),
    .X(clknet_5_19__leaf_clk));
 sg13g2_buf_1 clkbuf_5_20__f_clk (.A(clknet_4_10_0_clk),
    .X(clknet_5_20__leaf_clk));
 sg13g2_buf_1 clkbuf_5_21__f_clk (.A(clknet_4_10_0_clk),
    .X(clknet_5_21__leaf_clk));
 sg13g2_buf_1 clkbuf_5_22__f_clk (.A(clknet_4_11_0_clk),
    .X(clknet_5_22__leaf_clk));
 sg13g2_buf_1 clkbuf_5_23__f_clk (.A(clknet_4_11_0_clk),
    .X(clknet_5_23__leaf_clk));
 sg13g2_buf_1 clkbuf_5_24__f_clk (.A(clknet_4_12_0_clk),
    .X(clknet_5_24__leaf_clk));
 sg13g2_buf_1 clkbuf_5_25__f_clk (.A(clknet_4_12_0_clk),
    .X(clknet_5_25__leaf_clk));
 sg13g2_buf_1 clkbuf_5_26__f_clk (.A(clknet_4_13_0_clk),
    .X(clknet_5_26__leaf_clk));
 sg13g2_buf_1 clkbuf_5_27__f_clk (.A(clknet_4_13_0_clk),
    .X(clknet_5_27__leaf_clk));
 sg13g2_buf_1 clkbuf_5_28__f_clk (.A(clknet_4_14_0_clk),
    .X(clknet_5_28__leaf_clk));
 sg13g2_buf_1 clkbuf_5_29__f_clk (.A(clknet_4_14_0_clk),
    .X(clknet_5_29__leaf_clk));
 sg13g2_buf_1 clkbuf_5_30__f_clk (.A(clknet_4_15_0_clk),
    .X(clknet_5_30__leaf_clk));
 sg13g2_buf_1 clkbuf_5_31__f_clk (.A(clknet_4_15_0_clk),
    .X(clknet_5_31__leaf_clk));
 sg13g2_inv_1 clkload0 (.A(clknet_5_3__leaf_clk));
 sg13g2_inv_1 clkload1 (.A(clknet_5_5__leaf_clk));
 sg13g2_inv_1 clkload2 (.A(clknet_5_7__leaf_clk));
 sg13g2_inv_1 clkload3 (.A(clknet_5_9__leaf_clk));
 sg13g2_inv_1 clkload4 (.A(clknet_5_11__leaf_clk));
 sg13g2_inv_1 clkload5 (.A(clknet_5_13__leaf_clk));
 sg13g2_inv_1 clkload6 (.A(clknet_5_15__leaf_clk));
 sg13g2_inv_1 clkload7 (.A(clknet_5_19__leaf_clk));
 sg13g2_inv_1 clkload8 (.A(clknet_5_21__leaf_clk));
 sg13g2_inv_1 clkload9 (.A(clknet_5_23__leaf_clk));
 sg13g2_inv_1 clkload10 (.A(clknet_5_25__leaf_clk));
 sg13g2_inv_1 clkload11 (.A(clknet_5_27__leaf_clk));
 sg13g2_inv_1 clkload12 (.A(clknet_5_29__leaf_clk));
 sg13g2_inv_1 clkload13 (.A(clknet_5_31__leaf_clk));
 sg13g2_antennanp ANTENNA_1 (.A(_0143_));
 sg13g2_antennanp ANTENNA_2 (.A(_0191_));
 sg13g2_antennanp ANTENNA_3 (.A(clk));
 sg13g2_antennanp ANTENNA_4 (.A(clk));
 sg13g2_antennanp ANTENNA_5 (.A(_0143_));
 sg13g2_antennanp ANTENNA_6 (.A(_0191_));
 sg13g2_antennanp ANTENNA_7 (.A(clk));
 sg13g2_antennanp ANTENNA_8 (.A(_0143_));
 sg13g2_antennanp ANTENNA_9 (.A(_0191_));
 sg13g2_antennanp ANTENNA_10 (.A(clk));
 sg13g2_antennanp ANTENNA_11 (.A(_0143_));
 sg13g2_antennanp ANTENNA_12 (.A(_0191_));
 sg13g2_antennanp ANTENNA_13 (.A(clk));
 sg13g2_antennanp ANTENNA_14 (.A(_0143_));
 sg13g2_antennanp ANTENNA_15 (.A(_0191_));
 sg13g2_antennanp ANTENNA_16 (.A(clk));
 sg13g2_antennanp ANTENNA_17 (.A(clk));
 sg13g2_antennanp ANTENNA_18 (.A(clk));
 sg13g2_decap_8 FILLER_0_0 ();
 sg13g2_decap_8 FILLER_0_7 ();
 sg13g2_decap_8 FILLER_0_14 ();
 sg13g2_decap_8 FILLER_0_21 ();
 sg13g2_decap_8 FILLER_0_28 ();
 sg13g2_decap_8 FILLER_0_35 ();
 sg13g2_decap_8 FILLER_0_42 ();
 sg13g2_decap_8 FILLER_0_49 ();
 sg13g2_decap_8 FILLER_0_56 ();
 sg13g2_decap_8 FILLER_0_63 ();
 sg13g2_decap_8 FILLER_0_70 ();
 sg13g2_decap_8 FILLER_0_77 ();
 sg13g2_decap_8 FILLER_0_84 ();
 sg13g2_decap_8 FILLER_0_91 ();
 sg13g2_decap_8 FILLER_0_98 ();
 sg13g2_decap_8 FILLER_0_105 ();
 sg13g2_decap_8 FILLER_0_112 ();
 sg13g2_decap_8 FILLER_0_119 ();
 sg13g2_decap_8 FILLER_0_126 ();
 sg13g2_decap_8 FILLER_0_133 ();
 sg13g2_decap_8 FILLER_0_140 ();
 sg13g2_decap_8 FILLER_0_147 ();
 sg13g2_decap_8 FILLER_0_154 ();
 sg13g2_decap_8 FILLER_0_161 ();
 sg13g2_decap_8 FILLER_0_168 ();
 sg13g2_decap_8 FILLER_0_175 ();
 sg13g2_decap_8 FILLER_0_182 ();
 sg13g2_decap_8 FILLER_0_189 ();
 sg13g2_decap_8 FILLER_0_196 ();
 sg13g2_decap_8 FILLER_0_203 ();
 sg13g2_decap_8 FILLER_0_210 ();
 sg13g2_decap_8 FILLER_0_217 ();
 sg13g2_decap_8 FILLER_0_224 ();
 sg13g2_decap_8 FILLER_0_231 ();
 sg13g2_decap_8 FILLER_0_238 ();
 sg13g2_decap_8 FILLER_0_245 ();
 sg13g2_decap_8 FILLER_0_252 ();
 sg13g2_decap_8 FILLER_0_259 ();
 sg13g2_decap_8 FILLER_0_266 ();
 sg13g2_decap_8 FILLER_0_273 ();
 sg13g2_decap_8 FILLER_0_280 ();
 sg13g2_decap_8 FILLER_0_287 ();
 sg13g2_decap_8 FILLER_0_294 ();
 sg13g2_decap_8 FILLER_0_301 ();
 sg13g2_decap_8 FILLER_0_308 ();
 sg13g2_decap_8 FILLER_0_315 ();
 sg13g2_decap_8 FILLER_0_322 ();
 sg13g2_fill_2 FILLER_0_329 ();
 sg13g2_decap_8 FILLER_0_335 ();
 sg13g2_decap_8 FILLER_0_342 ();
 sg13g2_decap_8 FILLER_0_349 ();
 sg13g2_decap_8 FILLER_0_356 ();
 sg13g2_decap_8 FILLER_0_363 ();
 sg13g2_decap_8 FILLER_0_370 ();
 sg13g2_decap_8 FILLER_0_377 ();
 sg13g2_decap_8 FILLER_0_384 ();
 sg13g2_decap_8 FILLER_0_391 ();
 sg13g2_decap_8 FILLER_0_398 ();
 sg13g2_decap_8 FILLER_0_405 ();
 sg13g2_decap_8 FILLER_0_412 ();
 sg13g2_decap_8 FILLER_0_419 ();
 sg13g2_decap_4 FILLER_0_426 ();
 sg13g2_decap_8 FILLER_1_0 ();
 sg13g2_decap_8 FILLER_1_7 ();
 sg13g2_decap_8 FILLER_1_14 ();
 sg13g2_decap_8 FILLER_1_21 ();
 sg13g2_decap_8 FILLER_1_28 ();
 sg13g2_decap_8 FILLER_1_35 ();
 sg13g2_decap_8 FILLER_1_42 ();
 sg13g2_decap_8 FILLER_1_49 ();
 sg13g2_decap_8 FILLER_1_56 ();
 sg13g2_decap_8 FILLER_1_63 ();
 sg13g2_decap_8 FILLER_1_70 ();
 sg13g2_decap_8 FILLER_1_77 ();
 sg13g2_decap_8 FILLER_1_84 ();
 sg13g2_decap_8 FILLER_1_91 ();
 sg13g2_decap_8 FILLER_1_98 ();
 sg13g2_decap_8 FILLER_1_105 ();
 sg13g2_decap_8 FILLER_1_112 ();
 sg13g2_decap_8 FILLER_1_119 ();
 sg13g2_decap_8 FILLER_1_126 ();
 sg13g2_decap_8 FILLER_1_133 ();
 sg13g2_decap_8 FILLER_1_140 ();
 sg13g2_decap_8 FILLER_1_147 ();
 sg13g2_decap_8 FILLER_1_154 ();
 sg13g2_decap_8 FILLER_1_161 ();
 sg13g2_decap_8 FILLER_1_168 ();
 sg13g2_decap_8 FILLER_1_175 ();
 sg13g2_decap_8 FILLER_1_182 ();
 sg13g2_decap_8 FILLER_1_189 ();
 sg13g2_decap_8 FILLER_1_196 ();
 sg13g2_decap_8 FILLER_1_203 ();
 sg13g2_decap_8 FILLER_1_210 ();
 sg13g2_decap_8 FILLER_1_217 ();
 sg13g2_decap_8 FILLER_1_224 ();
 sg13g2_decap_8 FILLER_1_231 ();
 sg13g2_decap_8 FILLER_1_238 ();
 sg13g2_decap_8 FILLER_1_245 ();
 sg13g2_decap_8 FILLER_1_252 ();
 sg13g2_decap_8 FILLER_1_259 ();
 sg13g2_decap_4 FILLER_1_266 ();
 sg13g2_decap_4 FILLER_1_305 ();
 sg13g2_fill_2 FILLER_1_361 ();
 sg13g2_decap_8 FILLER_1_371 ();
 sg13g2_decap_8 FILLER_1_378 ();
 sg13g2_decap_8 FILLER_1_385 ();
 sg13g2_decap_8 FILLER_1_392 ();
 sg13g2_decap_8 FILLER_1_399 ();
 sg13g2_decap_8 FILLER_1_406 ();
 sg13g2_decap_8 FILLER_1_413 ();
 sg13g2_decap_8 FILLER_1_420 ();
 sg13g2_fill_2 FILLER_1_427 ();
 sg13g2_fill_1 FILLER_1_429 ();
 sg13g2_decap_8 FILLER_2_0 ();
 sg13g2_decap_8 FILLER_2_7 ();
 sg13g2_decap_8 FILLER_2_14 ();
 sg13g2_decap_8 FILLER_2_21 ();
 sg13g2_decap_8 FILLER_2_28 ();
 sg13g2_decap_8 FILLER_2_35 ();
 sg13g2_decap_8 FILLER_2_42 ();
 sg13g2_decap_8 FILLER_2_49 ();
 sg13g2_decap_8 FILLER_2_56 ();
 sg13g2_decap_8 FILLER_2_63 ();
 sg13g2_decap_8 FILLER_2_70 ();
 sg13g2_decap_8 FILLER_2_77 ();
 sg13g2_decap_8 FILLER_2_84 ();
 sg13g2_decap_8 FILLER_2_91 ();
 sg13g2_decap_8 FILLER_2_98 ();
 sg13g2_decap_8 FILLER_2_105 ();
 sg13g2_decap_8 FILLER_2_112 ();
 sg13g2_decap_8 FILLER_2_119 ();
 sg13g2_decap_8 FILLER_2_126 ();
 sg13g2_decap_8 FILLER_2_133 ();
 sg13g2_decap_8 FILLER_2_140 ();
 sg13g2_decap_8 FILLER_2_147 ();
 sg13g2_decap_8 FILLER_2_154 ();
 sg13g2_decap_8 FILLER_2_161 ();
 sg13g2_decap_8 FILLER_2_168 ();
 sg13g2_decap_8 FILLER_2_175 ();
 sg13g2_decap_8 FILLER_2_182 ();
 sg13g2_decap_8 FILLER_2_189 ();
 sg13g2_decap_8 FILLER_2_196 ();
 sg13g2_decap_8 FILLER_2_203 ();
 sg13g2_decap_8 FILLER_2_210 ();
 sg13g2_decap_8 FILLER_2_217 ();
 sg13g2_decap_8 FILLER_2_224 ();
 sg13g2_decap_8 FILLER_2_231 ();
 sg13g2_decap_8 FILLER_2_238 ();
 sg13g2_decap_8 FILLER_2_245 ();
 sg13g2_decap_8 FILLER_2_252 ();
 sg13g2_fill_2 FILLER_2_259 ();
 sg13g2_fill_1 FILLER_2_261 ();
 sg13g2_decap_8 FILLER_2_266 ();
 sg13g2_decap_4 FILLER_2_273 ();
 sg13g2_fill_2 FILLER_2_277 ();
 sg13g2_fill_2 FILLER_2_283 ();
 sg13g2_fill_2 FILLER_2_329 ();
 sg13g2_fill_2 FILLER_2_341 ();
 sg13g2_fill_1 FILLER_2_343 ();
 sg13g2_fill_1 FILLER_2_350 ();
 sg13g2_decap_8 FILLER_2_390 ();
 sg13g2_decap_8 FILLER_2_397 ();
 sg13g2_decap_8 FILLER_2_404 ();
 sg13g2_decap_8 FILLER_2_411 ();
 sg13g2_decap_8 FILLER_2_418 ();
 sg13g2_decap_4 FILLER_2_425 ();
 sg13g2_fill_1 FILLER_2_429 ();
 sg13g2_decap_8 FILLER_3_0 ();
 sg13g2_decap_8 FILLER_3_7 ();
 sg13g2_decap_8 FILLER_3_14 ();
 sg13g2_decap_8 FILLER_3_21 ();
 sg13g2_decap_8 FILLER_3_28 ();
 sg13g2_decap_8 FILLER_3_35 ();
 sg13g2_decap_8 FILLER_3_42 ();
 sg13g2_decap_8 FILLER_3_49 ();
 sg13g2_decap_8 FILLER_3_56 ();
 sg13g2_decap_8 FILLER_3_63 ();
 sg13g2_decap_8 FILLER_3_70 ();
 sg13g2_decap_8 FILLER_3_77 ();
 sg13g2_decap_8 FILLER_3_84 ();
 sg13g2_decap_8 FILLER_3_91 ();
 sg13g2_decap_8 FILLER_3_98 ();
 sg13g2_decap_8 FILLER_3_105 ();
 sg13g2_decap_8 FILLER_3_112 ();
 sg13g2_decap_8 FILLER_3_119 ();
 sg13g2_decap_8 FILLER_3_126 ();
 sg13g2_decap_8 FILLER_3_133 ();
 sg13g2_decap_8 FILLER_3_140 ();
 sg13g2_decap_8 FILLER_3_147 ();
 sg13g2_decap_8 FILLER_3_154 ();
 sg13g2_decap_8 FILLER_3_187 ();
 sg13g2_decap_8 FILLER_3_194 ();
 sg13g2_decap_8 FILLER_3_205 ();
 sg13g2_decap_8 FILLER_3_212 ();
 sg13g2_decap_8 FILLER_3_219 ();
 sg13g2_decap_8 FILLER_3_226 ();
 sg13g2_decap_8 FILLER_3_233 ();
 sg13g2_decap_8 FILLER_3_240 ();
 sg13g2_decap_8 FILLER_3_247 ();
 sg13g2_fill_1 FILLER_3_254 ();
 sg13g2_decap_8 FILLER_3_281 ();
 sg13g2_fill_2 FILLER_3_288 ();
 sg13g2_fill_1 FILLER_3_290 ();
 sg13g2_decap_8 FILLER_3_295 ();
 sg13g2_decap_4 FILLER_3_302 ();
 sg13g2_fill_2 FILLER_3_306 ();
 sg13g2_fill_1 FILLER_3_327 ();
 sg13g2_decap_8 FILLER_3_333 ();
 sg13g2_decap_8 FILLER_3_340 ();
 sg13g2_decap_4 FILLER_3_347 ();
 sg13g2_fill_1 FILLER_3_351 ();
 sg13g2_decap_8 FILLER_3_356 ();
 sg13g2_fill_1 FILLER_3_363 ();
 sg13g2_decap_8 FILLER_3_403 ();
 sg13g2_decap_8 FILLER_3_410 ();
 sg13g2_decap_8 FILLER_3_417 ();
 sg13g2_decap_4 FILLER_3_424 ();
 sg13g2_fill_2 FILLER_3_428 ();
 sg13g2_decap_8 FILLER_4_0 ();
 sg13g2_decap_8 FILLER_4_7 ();
 sg13g2_decap_8 FILLER_4_14 ();
 sg13g2_decap_8 FILLER_4_21 ();
 sg13g2_decap_8 FILLER_4_28 ();
 sg13g2_decap_8 FILLER_4_35 ();
 sg13g2_decap_8 FILLER_4_42 ();
 sg13g2_decap_8 FILLER_4_49 ();
 sg13g2_decap_8 FILLER_4_56 ();
 sg13g2_decap_8 FILLER_4_63 ();
 sg13g2_decap_8 FILLER_4_70 ();
 sg13g2_decap_8 FILLER_4_77 ();
 sg13g2_decap_8 FILLER_4_84 ();
 sg13g2_decap_8 FILLER_4_91 ();
 sg13g2_decap_8 FILLER_4_98 ();
 sg13g2_decap_8 FILLER_4_105 ();
 sg13g2_decap_8 FILLER_4_112 ();
 sg13g2_decap_8 FILLER_4_119 ();
 sg13g2_decap_8 FILLER_4_126 ();
 sg13g2_decap_8 FILLER_4_133 ();
 sg13g2_decap_8 FILLER_4_140 ();
 sg13g2_decap_8 FILLER_4_147 ();
 sg13g2_decap_8 FILLER_4_154 ();
 sg13g2_decap_4 FILLER_4_161 ();
 sg13g2_fill_1 FILLER_4_165 ();
 sg13g2_decap_8 FILLER_4_170 ();
 sg13g2_fill_2 FILLER_4_177 ();
 sg13g2_fill_1 FILLER_4_179 ();
 sg13g2_decap_8 FILLER_4_188 ();
 sg13g2_decap_8 FILLER_4_221 ();
 sg13g2_decap_8 FILLER_4_228 ();
 sg13g2_decap_8 FILLER_4_235 ();
 sg13g2_decap_8 FILLER_4_242 ();
 sg13g2_decap_8 FILLER_4_253 ();
 sg13g2_decap_8 FILLER_4_260 ();
 sg13g2_decap_8 FILLER_4_267 ();
 sg13g2_decap_8 FILLER_4_278 ();
 sg13g2_decap_8 FILLER_4_285 ();
 sg13g2_decap_4 FILLER_4_292 ();
 sg13g2_fill_1 FILLER_4_296 ();
 sg13g2_decap_8 FILLER_4_310 ();
 sg13g2_fill_1 FILLER_4_317 ();
 sg13g2_decap_4 FILLER_4_334 ();
 sg13g2_decap_4 FILLER_4_351 ();
 sg13g2_fill_2 FILLER_4_355 ();
 sg13g2_decap_8 FILLER_4_381 ();
 sg13g2_decap_8 FILLER_4_388 ();
 sg13g2_decap_8 FILLER_4_395 ();
 sg13g2_decap_8 FILLER_4_402 ();
 sg13g2_decap_8 FILLER_4_409 ();
 sg13g2_decap_8 FILLER_4_416 ();
 sg13g2_decap_8 FILLER_4_423 ();
 sg13g2_decap_8 FILLER_5_0 ();
 sg13g2_decap_8 FILLER_5_7 ();
 sg13g2_decap_8 FILLER_5_14 ();
 sg13g2_decap_8 FILLER_5_21 ();
 sg13g2_decap_8 FILLER_5_28 ();
 sg13g2_decap_8 FILLER_5_35 ();
 sg13g2_decap_8 FILLER_5_42 ();
 sg13g2_decap_8 FILLER_5_49 ();
 sg13g2_decap_8 FILLER_5_56 ();
 sg13g2_decap_8 FILLER_5_63 ();
 sg13g2_decap_8 FILLER_5_70 ();
 sg13g2_decap_8 FILLER_5_77 ();
 sg13g2_decap_8 FILLER_5_84 ();
 sg13g2_decap_8 FILLER_5_91 ();
 sg13g2_decap_8 FILLER_5_98 ();
 sg13g2_decap_8 FILLER_5_105 ();
 sg13g2_decap_8 FILLER_5_112 ();
 sg13g2_decap_8 FILLER_5_119 ();
 sg13g2_decap_8 FILLER_5_126 ();
 sg13g2_fill_2 FILLER_5_133 ();
 sg13g2_decap_8 FILLER_5_161 ();
 sg13g2_decap_8 FILLER_5_168 ();
 sg13g2_decap_4 FILLER_5_175 ();
 sg13g2_fill_2 FILLER_5_179 ();
 sg13g2_decap_8 FILLER_5_186 ();
 sg13g2_decap_4 FILLER_5_193 ();
 sg13g2_fill_2 FILLER_5_197 ();
 sg13g2_decap_8 FILLER_5_207 ();
 sg13g2_decap_8 FILLER_5_223 ();
 sg13g2_decap_8 FILLER_5_230 ();
 sg13g2_decap_4 FILLER_5_237 ();
 sg13g2_fill_2 FILLER_5_293 ();
 sg13g2_decap_4 FILLER_5_300 ();
 sg13g2_fill_1 FILLER_5_304 ();
 sg13g2_decap_4 FILLER_5_314 ();
 sg13g2_fill_2 FILLER_5_318 ();
 sg13g2_decap_8 FILLER_5_340 ();
 sg13g2_decap_4 FILLER_5_347 ();
 sg13g2_fill_2 FILLER_5_351 ();
 sg13g2_fill_1 FILLER_5_369 ();
 sg13g2_decap_8 FILLER_5_375 ();
 sg13g2_fill_2 FILLER_5_382 ();
 sg13g2_decap_4 FILLER_5_389 ();
 sg13g2_decap_8 FILLER_5_406 ();
 sg13g2_decap_8 FILLER_5_413 ();
 sg13g2_decap_8 FILLER_5_420 ();
 sg13g2_fill_2 FILLER_5_427 ();
 sg13g2_fill_1 FILLER_5_429 ();
 sg13g2_decap_8 FILLER_6_0 ();
 sg13g2_decap_8 FILLER_6_7 ();
 sg13g2_decap_8 FILLER_6_14 ();
 sg13g2_decap_8 FILLER_6_21 ();
 sg13g2_decap_8 FILLER_6_28 ();
 sg13g2_decap_8 FILLER_6_35 ();
 sg13g2_decap_8 FILLER_6_42 ();
 sg13g2_decap_8 FILLER_6_49 ();
 sg13g2_decap_8 FILLER_6_56 ();
 sg13g2_decap_8 FILLER_6_63 ();
 sg13g2_decap_8 FILLER_6_70 ();
 sg13g2_decap_8 FILLER_6_77 ();
 sg13g2_decap_8 FILLER_6_84 ();
 sg13g2_decap_8 FILLER_6_91 ();
 sg13g2_decap_8 FILLER_6_98 ();
 sg13g2_decap_8 FILLER_6_105 ();
 sg13g2_decap_8 FILLER_6_112 ();
 sg13g2_decap_8 FILLER_6_119 ();
 sg13g2_decap_8 FILLER_6_126 ();
 sg13g2_decap_4 FILLER_6_133 ();
 sg13g2_fill_1 FILLER_6_137 ();
 sg13g2_fill_2 FILLER_6_173 ();
 sg13g2_fill_1 FILLER_6_175 ();
 sg13g2_fill_1 FILLER_6_189 ();
 sg13g2_decap_4 FILLER_6_195 ();
 sg13g2_fill_2 FILLER_6_210 ();
 sg13g2_decap_8 FILLER_6_238 ();
 sg13g2_fill_1 FILLER_6_278 ();
 sg13g2_fill_2 FILLER_6_283 ();
 sg13g2_fill_1 FILLER_6_285 ();
 sg13g2_decap_4 FILLER_6_294 ();
 sg13g2_fill_1 FILLER_6_298 ();
 sg13g2_fill_1 FILLER_6_303 ();
 sg13g2_fill_2 FILLER_6_311 ();
 sg13g2_decap_4 FILLER_6_317 ();
 sg13g2_fill_2 FILLER_6_321 ();
 sg13g2_decap_4 FILLER_6_331 ();
 sg13g2_fill_2 FILLER_6_343 ();
 sg13g2_fill_1 FILLER_6_345 ();
 sg13g2_decap_8 FILLER_6_354 ();
 sg13g2_fill_1 FILLER_6_361 ();
 sg13g2_fill_2 FILLER_6_367 ();
 sg13g2_fill_1 FILLER_6_374 ();
 sg13g2_decap_8 FILLER_6_405 ();
 sg13g2_decap_8 FILLER_6_412 ();
 sg13g2_decap_8 FILLER_6_419 ();
 sg13g2_decap_4 FILLER_6_426 ();
 sg13g2_decap_8 FILLER_7_0 ();
 sg13g2_decap_8 FILLER_7_7 ();
 sg13g2_decap_8 FILLER_7_14 ();
 sg13g2_decap_8 FILLER_7_21 ();
 sg13g2_decap_8 FILLER_7_28 ();
 sg13g2_decap_8 FILLER_7_35 ();
 sg13g2_decap_8 FILLER_7_42 ();
 sg13g2_decap_8 FILLER_7_49 ();
 sg13g2_decap_8 FILLER_7_56 ();
 sg13g2_decap_8 FILLER_7_63 ();
 sg13g2_decap_8 FILLER_7_70 ();
 sg13g2_decap_8 FILLER_7_77 ();
 sg13g2_decap_8 FILLER_7_84 ();
 sg13g2_decap_8 FILLER_7_91 ();
 sg13g2_decap_8 FILLER_7_98 ();
 sg13g2_decap_8 FILLER_7_105 ();
 sg13g2_decap_8 FILLER_7_112 ();
 sg13g2_decap_8 FILLER_7_119 ();
 sg13g2_fill_2 FILLER_7_126 ();
 sg13g2_fill_1 FILLER_7_128 ();
 sg13g2_decap_8 FILLER_7_133 ();
 sg13g2_fill_2 FILLER_7_140 ();
 sg13g2_fill_2 FILLER_7_150 ();
 sg13g2_fill_1 FILLER_7_156 ();
 sg13g2_decap_4 FILLER_7_161 ();
 sg13g2_fill_2 FILLER_7_179 ();
 sg13g2_fill_1 FILLER_7_210 ();
 sg13g2_fill_2 FILLER_7_220 ();
 sg13g2_fill_1 FILLER_7_222 ();
 sg13g2_fill_1 FILLER_7_227 ();
 sg13g2_fill_1 FILLER_7_245 ();
 sg13g2_decap_4 FILLER_7_250 ();
 sg13g2_decap_8 FILLER_7_258 ();
 sg13g2_fill_1 FILLER_7_265 ();
 sg13g2_decap_8 FILLER_7_296 ();
 sg13g2_fill_2 FILLER_7_303 ();
 sg13g2_fill_1 FILLER_7_305 ();
 sg13g2_decap_4 FILLER_7_311 ();
 sg13g2_fill_2 FILLER_7_320 ();
 sg13g2_fill_2 FILLER_7_347 ();
 sg13g2_fill_2 FILLER_7_354 ();
 sg13g2_fill_1 FILLER_7_374 ();
 sg13g2_decap_4 FILLER_7_379 ();
 sg13g2_decap_8 FILLER_7_387 ();
 sg13g2_decap_8 FILLER_7_394 ();
 sg13g2_decap_8 FILLER_7_401 ();
 sg13g2_decap_8 FILLER_7_408 ();
 sg13g2_decap_8 FILLER_7_415 ();
 sg13g2_decap_8 FILLER_7_422 ();
 sg13g2_fill_1 FILLER_7_429 ();
 sg13g2_decap_8 FILLER_8_0 ();
 sg13g2_decap_8 FILLER_8_7 ();
 sg13g2_decap_8 FILLER_8_14 ();
 sg13g2_decap_8 FILLER_8_21 ();
 sg13g2_decap_8 FILLER_8_28 ();
 sg13g2_decap_8 FILLER_8_35 ();
 sg13g2_decap_8 FILLER_8_42 ();
 sg13g2_decap_8 FILLER_8_49 ();
 sg13g2_decap_8 FILLER_8_56 ();
 sg13g2_decap_8 FILLER_8_63 ();
 sg13g2_decap_8 FILLER_8_70 ();
 sg13g2_decap_8 FILLER_8_77 ();
 sg13g2_decap_8 FILLER_8_84 ();
 sg13g2_decap_8 FILLER_8_91 ();
 sg13g2_decap_8 FILLER_8_98 ();
 sg13g2_decap_8 FILLER_8_105 ();
 sg13g2_decap_8 FILLER_8_112 ();
 sg13g2_fill_1 FILLER_8_119 ();
 sg13g2_fill_2 FILLER_8_150 ();
 sg13g2_fill_1 FILLER_8_152 ();
 sg13g2_fill_1 FILLER_8_157 ();
 sg13g2_decap_8 FILLER_8_162 ();
 sg13g2_decap_8 FILLER_8_202 ();
 sg13g2_fill_1 FILLER_8_216 ();
 sg13g2_decap_4 FILLER_8_232 ();
 sg13g2_fill_2 FILLER_8_236 ();
 sg13g2_decap_8 FILLER_8_247 ();
 sg13g2_fill_2 FILLER_8_254 ();
 sg13g2_fill_1 FILLER_8_256 ();
 sg13g2_decap_8 FILLER_8_263 ();
 sg13g2_fill_1 FILLER_8_270 ();
 sg13g2_fill_2 FILLER_8_275 ();
 sg13g2_decap_4 FILLER_8_281 ();
 sg13g2_fill_2 FILLER_8_298 ();
 sg13g2_fill_1 FILLER_8_314 ();
 sg13g2_fill_1 FILLER_8_319 ();
 sg13g2_fill_1 FILLER_8_387 ();
 sg13g2_decap_8 FILLER_8_392 ();
 sg13g2_decap_8 FILLER_8_399 ();
 sg13g2_decap_8 FILLER_8_406 ();
 sg13g2_decap_8 FILLER_8_413 ();
 sg13g2_decap_8 FILLER_8_420 ();
 sg13g2_fill_2 FILLER_8_427 ();
 sg13g2_fill_1 FILLER_8_429 ();
 sg13g2_decap_8 FILLER_9_0 ();
 sg13g2_decap_8 FILLER_9_7 ();
 sg13g2_decap_8 FILLER_9_14 ();
 sg13g2_decap_8 FILLER_9_21 ();
 sg13g2_decap_8 FILLER_9_28 ();
 sg13g2_decap_8 FILLER_9_35 ();
 sg13g2_decap_8 FILLER_9_42 ();
 sg13g2_decap_8 FILLER_9_49 ();
 sg13g2_decap_8 FILLER_9_56 ();
 sg13g2_decap_8 FILLER_9_63 ();
 sg13g2_decap_8 FILLER_9_70 ();
 sg13g2_decap_8 FILLER_9_77 ();
 sg13g2_decap_8 FILLER_9_84 ();
 sg13g2_decap_8 FILLER_9_91 ();
 sg13g2_decap_8 FILLER_9_98 ();
 sg13g2_decap_8 FILLER_9_105 ();
 sg13g2_decap_8 FILLER_9_112 ();
 sg13g2_decap_8 FILLER_9_119 ();
 sg13g2_decap_8 FILLER_9_126 ();
 sg13g2_decap_8 FILLER_9_133 ();
 sg13g2_decap_4 FILLER_9_140 ();
 sg13g2_fill_2 FILLER_9_149 ();
 sg13g2_fill_1 FILLER_9_151 ();
 sg13g2_decap_8 FILLER_9_158 ();
 sg13g2_fill_2 FILLER_9_165 ();
 sg13g2_fill_2 FILLER_9_177 ();
 sg13g2_fill_1 FILLER_9_179 ();
 sg13g2_fill_1 FILLER_9_188 ();
 sg13g2_decap_4 FILLER_9_199 ();
 sg13g2_fill_1 FILLER_9_203 ();
 sg13g2_fill_1 FILLER_9_209 ();
 sg13g2_fill_1 FILLER_9_213 ();
 sg13g2_decap_4 FILLER_9_227 ();
 sg13g2_fill_2 FILLER_9_253 ();
 sg13g2_fill_1 FILLER_9_260 ();
 sg13g2_decap_4 FILLER_9_279 ();
 sg13g2_fill_1 FILLER_9_287 ();
 sg13g2_fill_1 FILLER_9_294 ();
 sg13g2_fill_1 FILLER_9_300 ();
 sg13g2_fill_1 FILLER_9_306 ();
 sg13g2_fill_1 FILLER_9_311 ();
 sg13g2_decap_4 FILLER_9_317 ();
 sg13g2_fill_1 FILLER_9_321 ();
 sg13g2_fill_2 FILLER_9_341 ();
 sg13g2_decap_4 FILLER_9_346 ();
 sg13g2_decap_4 FILLER_9_367 ();
 sg13g2_fill_1 FILLER_9_371 ();
 sg13g2_decap_8 FILLER_9_407 ();
 sg13g2_decap_8 FILLER_9_414 ();
 sg13g2_decap_8 FILLER_9_421 ();
 sg13g2_fill_2 FILLER_9_428 ();
 sg13g2_decap_8 FILLER_10_0 ();
 sg13g2_decap_8 FILLER_10_7 ();
 sg13g2_decap_8 FILLER_10_14 ();
 sg13g2_decap_8 FILLER_10_21 ();
 sg13g2_decap_8 FILLER_10_28 ();
 sg13g2_decap_8 FILLER_10_35 ();
 sg13g2_decap_8 FILLER_10_42 ();
 sg13g2_decap_8 FILLER_10_49 ();
 sg13g2_decap_8 FILLER_10_56 ();
 sg13g2_decap_8 FILLER_10_63 ();
 sg13g2_decap_8 FILLER_10_70 ();
 sg13g2_decap_8 FILLER_10_77 ();
 sg13g2_decap_8 FILLER_10_84 ();
 sg13g2_decap_8 FILLER_10_91 ();
 sg13g2_decap_8 FILLER_10_98 ();
 sg13g2_decap_8 FILLER_10_105 ();
 sg13g2_decap_8 FILLER_10_112 ();
 sg13g2_decap_8 FILLER_10_119 ();
 sg13g2_fill_2 FILLER_10_152 ();
 sg13g2_decap_4 FILLER_10_163 ();
 sg13g2_fill_1 FILLER_10_167 ();
 sg13g2_fill_1 FILLER_10_172 ();
 sg13g2_fill_2 FILLER_10_179 ();
 sg13g2_decap_8 FILLER_10_194 ();
 sg13g2_fill_2 FILLER_10_201 ();
 sg13g2_fill_1 FILLER_10_225 ();
 sg13g2_fill_1 FILLER_10_234 ();
 sg13g2_fill_2 FILLER_10_250 ();
 sg13g2_fill_2 FILLER_10_257 ();
 sg13g2_fill_2 FILLER_10_264 ();
 sg13g2_fill_1 FILLER_10_279 ();
 sg13g2_fill_1 FILLER_10_302 ();
 sg13g2_fill_1 FILLER_10_308 ();
 sg13g2_fill_1 FILLER_10_314 ();
 sg13g2_fill_1 FILLER_10_320 ();
 sg13g2_fill_1 FILLER_10_329 ();
 sg13g2_decap_8 FILLER_10_335 ();
 sg13g2_decap_8 FILLER_10_346 ();
 sg13g2_fill_1 FILLER_10_359 ();
 sg13g2_fill_1 FILLER_10_367 ();
 sg13g2_fill_1 FILLER_10_373 ();
 sg13g2_fill_2 FILLER_10_383 ();
 sg13g2_fill_2 FILLER_10_390 ();
 sg13g2_decap_8 FILLER_10_396 ();
 sg13g2_decap_8 FILLER_10_403 ();
 sg13g2_decap_8 FILLER_10_410 ();
 sg13g2_decap_8 FILLER_10_417 ();
 sg13g2_decap_4 FILLER_10_424 ();
 sg13g2_fill_2 FILLER_10_428 ();
 sg13g2_decap_8 FILLER_11_0 ();
 sg13g2_decap_8 FILLER_11_7 ();
 sg13g2_decap_8 FILLER_11_14 ();
 sg13g2_decap_8 FILLER_11_21 ();
 sg13g2_decap_8 FILLER_11_28 ();
 sg13g2_decap_8 FILLER_11_35 ();
 sg13g2_decap_8 FILLER_11_42 ();
 sg13g2_decap_8 FILLER_11_49 ();
 sg13g2_decap_8 FILLER_11_56 ();
 sg13g2_decap_8 FILLER_11_63 ();
 sg13g2_decap_8 FILLER_11_70 ();
 sg13g2_decap_8 FILLER_11_77 ();
 sg13g2_decap_8 FILLER_11_84 ();
 sg13g2_decap_8 FILLER_11_91 ();
 sg13g2_decap_8 FILLER_11_98 ();
 sg13g2_decap_8 FILLER_11_105 ();
 sg13g2_decap_8 FILLER_11_112 ();
 sg13g2_decap_4 FILLER_11_119 ();
 sg13g2_fill_2 FILLER_11_140 ();
 sg13g2_fill_1 FILLER_11_142 ();
 sg13g2_fill_1 FILLER_11_147 ();
 sg13g2_decap_4 FILLER_11_152 ();
 sg13g2_fill_2 FILLER_11_156 ();
 sg13g2_decap_8 FILLER_11_167 ();
 sg13g2_decap_8 FILLER_11_174 ();
 sg13g2_decap_4 FILLER_11_184 ();
 sg13g2_decap_8 FILLER_11_198 ();
 sg13g2_fill_2 FILLER_11_205 ();
 sg13g2_fill_1 FILLER_11_207 ();
 sg13g2_fill_2 FILLER_11_218 ();
 sg13g2_decap_4 FILLER_11_226 ();
 sg13g2_fill_2 FILLER_11_239 ();
 sg13g2_decap_8 FILLER_11_250 ();
 sg13g2_decap_8 FILLER_11_257 ();
 sg13g2_decap_4 FILLER_11_264 ();
 sg13g2_decap_4 FILLER_11_272 ();
 sg13g2_fill_1 FILLER_11_294 ();
 sg13g2_fill_2 FILLER_11_315 ();
 sg13g2_fill_2 FILLER_11_322 ();
 sg13g2_fill_1 FILLER_11_324 ();
 sg13g2_fill_2 FILLER_11_333 ();
 sg13g2_fill_1 FILLER_11_335 ();
 sg13g2_fill_2 FILLER_11_340 ();
 sg13g2_fill_1 FILLER_11_346 ();
 sg13g2_decap_4 FILLER_11_352 ();
 sg13g2_fill_1 FILLER_11_356 ();
 sg13g2_decap_8 FILLER_11_372 ();
 sg13g2_decap_8 FILLER_11_379 ();
 sg13g2_fill_2 FILLER_11_386 ();
 sg13g2_fill_1 FILLER_11_388 ();
 sg13g2_decap_8 FILLER_11_402 ();
 sg13g2_decap_8 FILLER_11_409 ();
 sg13g2_decap_8 FILLER_11_416 ();
 sg13g2_decap_8 FILLER_11_423 ();
 sg13g2_decap_8 FILLER_12_0 ();
 sg13g2_decap_8 FILLER_12_7 ();
 sg13g2_decap_8 FILLER_12_14 ();
 sg13g2_decap_8 FILLER_12_21 ();
 sg13g2_decap_8 FILLER_12_28 ();
 sg13g2_decap_8 FILLER_12_35 ();
 sg13g2_decap_8 FILLER_12_42 ();
 sg13g2_decap_8 FILLER_12_49 ();
 sg13g2_decap_8 FILLER_12_56 ();
 sg13g2_decap_8 FILLER_12_63 ();
 sg13g2_decap_8 FILLER_12_70 ();
 sg13g2_decap_8 FILLER_12_77 ();
 sg13g2_decap_8 FILLER_12_84 ();
 sg13g2_decap_8 FILLER_12_91 ();
 sg13g2_decap_8 FILLER_12_98 ();
 sg13g2_decap_8 FILLER_12_105 ();
 sg13g2_decap_4 FILLER_12_112 ();
 sg13g2_fill_2 FILLER_12_116 ();
 sg13g2_decap_4 FILLER_12_164 ();
 sg13g2_fill_1 FILLER_12_168 ();
 sg13g2_decap_4 FILLER_12_173 ();
 sg13g2_fill_2 FILLER_12_200 ();
 sg13g2_fill_1 FILLER_12_210 ();
 sg13g2_fill_1 FILLER_12_216 ();
 sg13g2_decap_8 FILLER_12_221 ();
 sg13g2_decap_8 FILLER_12_228 ();
 sg13g2_decap_8 FILLER_12_235 ();
 sg13g2_fill_1 FILLER_12_242 ();
 sg13g2_decap_8 FILLER_12_251 ();
 sg13g2_decap_4 FILLER_12_258 ();
 sg13g2_fill_1 FILLER_12_262 ();
 sg13g2_decap_4 FILLER_12_280 ();
 sg13g2_fill_2 FILLER_12_284 ();
 sg13g2_fill_1 FILLER_12_289 ();
 sg13g2_fill_1 FILLER_12_295 ();
 sg13g2_fill_1 FILLER_12_316 ();
 sg13g2_decap_4 FILLER_12_322 ();
 sg13g2_fill_2 FILLER_12_326 ();
 sg13g2_fill_2 FILLER_12_353 ();
 sg13g2_fill_1 FILLER_12_389 ();
 sg13g2_decap_8 FILLER_12_394 ();
 sg13g2_decap_4 FILLER_12_401 ();
 sg13g2_fill_1 FILLER_12_405 ();
 sg13g2_decap_8 FILLER_12_411 ();
 sg13g2_decap_8 FILLER_12_418 ();
 sg13g2_decap_4 FILLER_12_425 ();
 sg13g2_fill_1 FILLER_12_429 ();
 sg13g2_decap_8 FILLER_13_0 ();
 sg13g2_decap_8 FILLER_13_7 ();
 sg13g2_decap_8 FILLER_13_14 ();
 sg13g2_decap_8 FILLER_13_21 ();
 sg13g2_decap_8 FILLER_13_28 ();
 sg13g2_decap_8 FILLER_13_35 ();
 sg13g2_decap_8 FILLER_13_42 ();
 sg13g2_decap_8 FILLER_13_49 ();
 sg13g2_decap_8 FILLER_13_56 ();
 sg13g2_decap_8 FILLER_13_63 ();
 sg13g2_decap_8 FILLER_13_70 ();
 sg13g2_decap_8 FILLER_13_77 ();
 sg13g2_decap_8 FILLER_13_84 ();
 sg13g2_decap_8 FILLER_13_91 ();
 sg13g2_decap_8 FILLER_13_98 ();
 sg13g2_fill_1 FILLER_13_105 ();
 sg13g2_decap_4 FILLER_13_136 ();
 sg13g2_fill_1 FILLER_13_140 ();
 sg13g2_fill_1 FILLER_13_146 ();
 sg13g2_fill_1 FILLER_13_157 ();
 sg13g2_fill_1 FILLER_13_168 ();
 sg13g2_fill_2 FILLER_13_181 ();
 sg13g2_fill_2 FILLER_13_187 ();
 sg13g2_fill_1 FILLER_13_189 ();
 sg13g2_fill_1 FILLER_13_214 ();
 sg13g2_fill_2 FILLER_13_220 ();
 sg13g2_decap_8 FILLER_13_227 ();
 sg13g2_fill_2 FILLER_13_234 ();
 sg13g2_decap_8 FILLER_13_246 ();
 sg13g2_decap_4 FILLER_13_253 ();
 sg13g2_decap_8 FILLER_13_281 ();
 sg13g2_decap_8 FILLER_13_288 ();
 sg13g2_decap_8 FILLER_13_295 ();
 sg13g2_fill_1 FILLER_13_319 ();
 sg13g2_fill_1 FILLER_13_341 ();
 sg13g2_decap_8 FILLER_13_350 ();
 sg13g2_fill_2 FILLER_13_357 ();
 sg13g2_fill_1 FILLER_13_359 ();
 sg13g2_decap_4 FILLER_13_382 ();
 sg13g2_fill_1 FILLER_13_386 ();
 sg13g2_decap_8 FILLER_13_417 ();
 sg13g2_decap_4 FILLER_13_424 ();
 sg13g2_fill_2 FILLER_13_428 ();
 sg13g2_decap_8 FILLER_14_0 ();
 sg13g2_decap_8 FILLER_14_7 ();
 sg13g2_decap_8 FILLER_14_14 ();
 sg13g2_decap_8 FILLER_14_21 ();
 sg13g2_decap_8 FILLER_14_28 ();
 sg13g2_decap_8 FILLER_14_35 ();
 sg13g2_decap_8 FILLER_14_42 ();
 sg13g2_decap_8 FILLER_14_49 ();
 sg13g2_decap_8 FILLER_14_56 ();
 sg13g2_decap_8 FILLER_14_63 ();
 sg13g2_decap_8 FILLER_14_70 ();
 sg13g2_decap_8 FILLER_14_77 ();
 sg13g2_decap_8 FILLER_14_84 ();
 sg13g2_decap_8 FILLER_14_91 ();
 sg13g2_decap_8 FILLER_14_98 ();
 sg13g2_decap_4 FILLER_14_105 ();
 sg13g2_fill_2 FILLER_14_109 ();
 sg13g2_decap_8 FILLER_14_115 ();
 sg13g2_decap_4 FILLER_14_122 ();
 sg13g2_fill_2 FILLER_14_126 ();
 sg13g2_decap_4 FILLER_14_132 ();
 sg13g2_fill_2 FILLER_14_136 ();
 sg13g2_fill_1 FILLER_14_145 ();
 sg13g2_fill_1 FILLER_14_151 ();
 sg13g2_fill_1 FILLER_14_160 ();
 sg13g2_fill_2 FILLER_14_166 ();
 sg13g2_fill_1 FILLER_14_190 ();
 sg13g2_fill_2 FILLER_14_195 ();
 sg13g2_fill_1 FILLER_14_207 ();
 sg13g2_fill_1 FILLER_14_215 ();
 sg13g2_fill_1 FILLER_14_221 ();
 sg13g2_fill_1 FILLER_14_234 ();
 sg13g2_fill_2 FILLER_14_239 ();
 sg13g2_fill_1 FILLER_14_241 ();
 sg13g2_fill_2 FILLER_14_250 ();
 sg13g2_decap_8 FILLER_14_271 ();
 sg13g2_decap_8 FILLER_14_278 ();
 sg13g2_fill_1 FILLER_14_285 ();
 sg13g2_fill_2 FILLER_14_318 ();
 sg13g2_fill_1 FILLER_14_320 ();
 sg13g2_fill_2 FILLER_14_326 ();
 sg13g2_fill_2 FILLER_14_333 ();
 sg13g2_fill_1 FILLER_14_335 ();
 sg13g2_decap_8 FILLER_14_351 ();
 sg13g2_decap_8 FILLER_14_358 ();
 sg13g2_fill_2 FILLER_14_365 ();
 sg13g2_fill_1 FILLER_14_381 ();
 sg13g2_fill_1 FILLER_14_387 ();
 sg13g2_decap_8 FILLER_14_392 ();
 sg13g2_fill_1 FILLER_14_403 ();
 sg13g2_decap_8 FILLER_14_408 ();
 sg13g2_decap_8 FILLER_14_415 ();
 sg13g2_decap_8 FILLER_14_422 ();
 sg13g2_fill_1 FILLER_14_429 ();
 sg13g2_decap_8 FILLER_15_0 ();
 sg13g2_decap_8 FILLER_15_7 ();
 sg13g2_decap_8 FILLER_15_14 ();
 sg13g2_decap_8 FILLER_15_21 ();
 sg13g2_decap_8 FILLER_15_28 ();
 sg13g2_decap_8 FILLER_15_35 ();
 sg13g2_decap_8 FILLER_15_42 ();
 sg13g2_decap_8 FILLER_15_49 ();
 sg13g2_decap_8 FILLER_15_56 ();
 sg13g2_decap_8 FILLER_15_63 ();
 sg13g2_decap_8 FILLER_15_70 ();
 sg13g2_decap_8 FILLER_15_77 ();
 sg13g2_decap_8 FILLER_15_84 ();
 sg13g2_decap_8 FILLER_15_91 ();
 sg13g2_decap_8 FILLER_15_98 ();
 sg13g2_decap_8 FILLER_15_105 ();
 sg13g2_decap_8 FILLER_15_112 ();
 sg13g2_decap_4 FILLER_15_119 ();
 sg13g2_fill_2 FILLER_15_123 ();
 sg13g2_decap_8 FILLER_15_129 ();
 sg13g2_fill_2 FILLER_15_136 ();
 sg13g2_fill_1 FILLER_15_138 ();
 sg13g2_decap_8 FILLER_15_156 ();
 sg13g2_decap_4 FILLER_15_167 ();
 sg13g2_decap_8 FILLER_15_181 ();
 sg13g2_fill_2 FILLER_15_193 ();
 sg13g2_fill_2 FILLER_15_201 ();
 sg13g2_fill_1 FILLER_15_203 ();
 sg13g2_fill_2 FILLER_15_207 ();
 sg13g2_fill_1 FILLER_15_209 ();
 sg13g2_fill_2 FILLER_15_214 ();
 sg13g2_fill_1 FILLER_15_216 ();
 sg13g2_decap_4 FILLER_15_227 ();
 sg13g2_fill_1 FILLER_15_231 ();
 sg13g2_fill_1 FILLER_15_241 ();
 sg13g2_fill_1 FILLER_15_247 ();
 sg13g2_fill_1 FILLER_15_258 ();
 sg13g2_fill_2 FILLER_15_263 ();
 sg13g2_fill_1 FILLER_15_265 ();
 sg13g2_decap_4 FILLER_15_271 ();
 sg13g2_decap_4 FILLER_15_290 ();
 sg13g2_decap_8 FILLER_15_318 ();
 sg13g2_decap_4 FILLER_15_325 ();
 sg13g2_fill_2 FILLER_15_335 ();
 sg13g2_decap_8 FILLER_15_342 ();
 sg13g2_fill_2 FILLER_15_349 ();
 sg13g2_fill_2 FILLER_15_383 ();
 sg13g2_fill_1 FILLER_15_385 ();
 sg13g2_decap_8 FILLER_15_391 ();
 sg13g2_decap_8 FILLER_15_398 ();
 sg13g2_decap_8 FILLER_15_405 ();
 sg13g2_decap_8 FILLER_15_412 ();
 sg13g2_decap_8 FILLER_15_419 ();
 sg13g2_decap_4 FILLER_15_426 ();
 sg13g2_decap_8 FILLER_16_0 ();
 sg13g2_decap_8 FILLER_16_7 ();
 sg13g2_decap_8 FILLER_16_14 ();
 sg13g2_decap_8 FILLER_16_21 ();
 sg13g2_decap_8 FILLER_16_28 ();
 sg13g2_decap_8 FILLER_16_35 ();
 sg13g2_decap_8 FILLER_16_42 ();
 sg13g2_decap_8 FILLER_16_49 ();
 sg13g2_decap_8 FILLER_16_56 ();
 sg13g2_decap_8 FILLER_16_63 ();
 sg13g2_decap_8 FILLER_16_70 ();
 sg13g2_decap_8 FILLER_16_77 ();
 sg13g2_decap_8 FILLER_16_84 ();
 sg13g2_decap_8 FILLER_16_91 ();
 sg13g2_decap_8 FILLER_16_98 ();
 sg13g2_decap_8 FILLER_16_105 ();
 sg13g2_decap_4 FILLER_16_112 ();
 sg13g2_fill_2 FILLER_16_116 ();
 sg13g2_fill_1 FILLER_16_125 ();
 sg13g2_fill_1 FILLER_16_131 ();
 sg13g2_fill_1 FILLER_16_139 ();
 sg13g2_fill_2 FILLER_16_148 ();
 sg13g2_decap_4 FILLER_16_158 ();
 sg13g2_decap_8 FILLER_16_178 ();
 sg13g2_fill_2 FILLER_16_192 ();
 sg13g2_fill_1 FILLER_16_194 ();
 sg13g2_decap_8 FILLER_16_199 ();
 sg13g2_decap_8 FILLER_16_206 ();
 sg13g2_fill_2 FILLER_16_213 ();
 sg13g2_fill_1 FILLER_16_215 ();
 sg13g2_fill_1 FILLER_16_220 ();
 sg13g2_decap_4 FILLER_16_232 ();
 sg13g2_fill_1 FILLER_16_236 ();
 sg13g2_fill_2 FILLER_16_244 ();
 sg13g2_decap_8 FILLER_16_265 ();
 sg13g2_decap_8 FILLER_16_272 ();
 sg13g2_fill_1 FILLER_16_279 ();
 sg13g2_decap_4 FILLER_16_286 ();
 sg13g2_fill_2 FILLER_16_290 ();
 sg13g2_decap_4 FILLER_16_300 ();
 sg13g2_fill_1 FILLER_16_304 ();
 sg13g2_decap_4 FILLER_16_310 ();
 sg13g2_decap_8 FILLER_16_322 ();
 sg13g2_fill_1 FILLER_16_329 ();
 sg13g2_decap_8 FILLER_16_339 ();
 sg13g2_fill_1 FILLER_16_346 ();
 sg13g2_decap_4 FILLER_16_351 ();
 sg13g2_fill_1 FILLER_16_355 ();
 sg13g2_fill_2 FILLER_16_360 ();
 sg13g2_fill_1 FILLER_16_362 ();
 sg13g2_decap_8 FILLER_16_368 ();
 sg13g2_decap_8 FILLER_16_375 ();
 sg13g2_decap_4 FILLER_16_382 ();
 sg13g2_fill_1 FILLER_16_386 ();
 sg13g2_decap_8 FILLER_16_395 ();
 sg13g2_decap_8 FILLER_16_402 ();
 sg13g2_decap_8 FILLER_16_409 ();
 sg13g2_decap_8 FILLER_16_416 ();
 sg13g2_decap_8 FILLER_16_423 ();
 sg13g2_decap_8 FILLER_17_0 ();
 sg13g2_decap_8 FILLER_17_7 ();
 sg13g2_decap_8 FILLER_17_14 ();
 sg13g2_decap_8 FILLER_17_21 ();
 sg13g2_decap_8 FILLER_17_28 ();
 sg13g2_decap_8 FILLER_17_35 ();
 sg13g2_decap_8 FILLER_17_42 ();
 sg13g2_decap_8 FILLER_17_49 ();
 sg13g2_decap_8 FILLER_17_56 ();
 sg13g2_decap_8 FILLER_17_63 ();
 sg13g2_decap_8 FILLER_17_70 ();
 sg13g2_decap_8 FILLER_17_77 ();
 sg13g2_decap_8 FILLER_17_84 ();
 sg13g2_decap_8 FILLER_17_91 ();
 sg13g2_decap_8 FILLER_17_98 ();
 sg13g2_decap_8 FILLER_17_105 ();
 sg13g2_fill_2 FILLER_17_112 ();
 sg13g2_fill_2 FILLER_17_140 ();
 sg13g2_fill_1 FILLER_17_142 ();
 sg13g2_decap_8 FILLER_17_148 ();
 sg13g2_fill_1 FILLER_17_159 ();
 sg13g2_fill_2 FILLER_17_169 ();
 sg13g2_fill_1 FILLER_17_171 ();
 sg13g2_fill_2 FILLER_17_177 ();
 sg13g2_fill_1 FILLER_17_179 ();
 sg13g2_fill_2 FILLER_17_185 ();
 sg13g2_decap_8 FILLER_17_218 ();
 sg13g2_fill_2 FILLER_17_234 ();
 sg13g2_fill_1 FILLER_17_236 ();
 sg13g2_fill_2 FILLER_17_249 ();
 sg13g2_decap_4 FILLER_17_255 ();
 sg13g2_decap_8 FILLER_17_269 ();
 sg13g2_decap_4 FILLER_17_276 ();
 sg13g2_decap_8 FILLER_17_288 ();
 sg13g2_fill_1 FILLER_17_295 ();
 sg13g2_decap_4 FILLER_17_304 ();
 sg13g2_fill_2 FILLER_17_314 ();
 sg13g2_decap_4 FILLER_17_321 ();
 sg13g2_fill_1 FILLER_17_348 ();
 sg13g2_fill_2 FILLER_17_364 ();
 sg13g2_fill_1 FILLER_17_366 ();
 sg13g2_fill_2 FILLER_17_371 ();
 sg13g2_fill_2 FILLER_17_401 ();
 sg13g2_decap_8 FILLER_17_407 ();
 sg13g2_decap_8 FILLER_17_414 ();
 sg13g2_decap_8 FILLER_17_421 ();
 sg13g2_fill_2 FILLER_17_428 ();
 sg13g2_decap_8 FILLER_18_0 ();
 sg13g2_decap_8 FILLER_18_7 ();
 sg13g2_decap_8 FILLER_18_14 ();
 sg13g2_decap_8 FILLER_18_21 ();
 sg13g2_decap_8 FILLER_18_28 ();
 sg13g2_decap_8 FILLER_18_35 ();
 sg13g2_decap_8 FILLER_18_42 ();
 sg13g2_decap_8 FILLER_18_49 ();
 sg13g2_decap_8 FILLER_18_56 ();
 sg13g2_decap_8 FILLER_18_63 ();
 sg13g2_decap_8 FILLER_18_70 ();
 sg13g2_decap_8 FILLER_18_77 ();
 sg13g2_decap_8 FILLER_18_84 ();
 sg13g2_decap_8 FILLER_18_91 ();
 sg13g2_decap_8 FILLER_18_98 ();
 sg13g2_decap_8 FILLER_18_105 ();
 sg13g2_fill_2 FILLER_18_112 ();
 sg13g2_fill_1 FILLER_18_114 ();
 sg13g2_fill_2 FILLER_18_120 ();
 sg13g2_decap_4 FILLER_18_131 ();
 sg13g2_fill_2 FILLER_18_135 ();
 sg13g2_decap_4 FILLER_18_141 ();
 sg13g2_decap_4 FILLER_18_149 ();
 sg13g2_fill_2 FILLER_18_153 ();
 sg13g2_fill_1 FILLER_18_178 ();
 sg13g2_fill_2 FILLER_18_184 ();
 sg13g2_fill_2 FILLER_18_192 ();
 sg13g2_decap_8 FILLER_18_197 ();
 sg13g2_decap_4 FILLER_18_204 ();
 sg13g2_fill_1 FILLER_18_208 ();
 sg13g2_decap_4 FILLER_18_214 ();
 sg13g2_fill_2 FILLER_18_218 ();
 sg13g2_decap_8 FILLER_18_225 ();
 sg13g2_decap_8 FILLER_18_232 ();
 sg13g2_decap_8 FILLER_18_239 ();
 sg13g2_fill_2 FILLER_18_246 ();
 sg13g2_fill_1 FILLER_18_248 ();
 sg13g2_fill_1 FILLER_18_254 ();
 sg13g2_fill_2 FILLER_18_259 ();
 sg13g2_fill_2 FILLER_18_265 ();
 sg13g2_fill_1 FILLER_18_267 ();
 sg13g2_fill_2 FILLER_18_281 ();
 sg13g2_fill_1 FILLER_18_287 ();
 sg13g2_decap_8 FILLER_18_298 ();
 sg13g2_decap_8 FILLER_18_305 ();
 sg13g2_fill_1 FILLER_18_312 ();
 sg13g2_fill_1 FILLER_18_321 ();
 sg13g2_fill_2 FILLER_18_347 ();
 sg13g2_fill_1 FILLER_18_349 ();
 sg13g2_fill_1 FILLER_18_354 ();
 sg13g2_decap_8 FILLER_18_366 ();
 sg13g2_fill_2 FILLER_18_373 ();
 sg13g2_fill_1 FILLER_18_375 ();
 sg13g2_fill_2 FILLER_18_381 ();
 sg13g2_fill_1 FILLER_18_402 ();
 sg13g2_decap_8 FILLER_18_411 ();
 sg13g2_decap_8 FILLER_18_418 ();
 sg13g2_decap_4 FILLER_18_425 ();
 sg13g2_fill_1 FILLER_18_429 ();
 sg13g2_decap_8 FILLER_19_0 ();
 sg13g2_decap_8 FILLER_19_7 ();
 sg13g2_decap_8 FILLER_19_14 ();
 sg13g2_decap_8 FILLER_19_21 ();
 sg13g2_decap_8 FILLER_19_28 ();
 sg13g2_decap_8 FILLER_19_35 ();
 sg13g2_decap_8 FILLER_19_42 ();
 sg13g2_decap_8 FILLER_19_49 ();
 sg13g2_decap_8 FILLER_19_56 ();
 sg13g2_decap_8 FILLER_19_63 ();
 sg13g2_decap_8 FILLER_19_70 ();
 sg13g2_decap_8 FILLER_19_77 ();
 sg13g2_decap_8 FILLER_19_84 ();
 sg13g2_decap_8 FILLER_19_91 ();
 sg13g2_decap_8 FILLER_19_98 ();
 sg13g2_decap_4 FILLER_19_105 ();
 sg13g2_decap_8 FILLER_19_129 ();
 sg13g2_fill_2 FILLER_19_136 ();
 sg13g2_fill_2 FILLER_19_143 ();
 sg13g2_decap_8 FILLER_19_153 ();
 sg13g2_fill_2 FILLER_19_160 ();
 sg13g2_fill_2 FILLER_19_175 ();
 sg13g2_fill_1 FILLER_19_187 ();
 sg13g2_decap_8 FILLER_19_193 ();
 sg13g2_fill_2 FILLER_19_200 ();
 sg13g2_fill_1 FILLER_19_202 ();
 sg13g2_decap_8 FILLER_19_218 ();
 sg13g2_decap_8 FILLER_19_225 ();
 sg13g2_decap_8 FILLER_19_232 ();
 sg13g2_decap_4 FILLER_19_239 ();
 sg13g2_fill_2 FILLER_19_243 ();
 sg13g2_fill_2 FILLER_19_265 ();
 sg13g2_fill_1 FILLER_19_287 ();
 sg13g2_decap_4 FILLER_19_297 ();
 sg13g2_fill_1 FILLER_19_301 ();
 sg13g2_fill_1 FILLER_19_307 ();
 sg13g2_decap_8 FILLER_19_316 ();
 sg13g2_decap_8 FILLER_19_323 ();
 sg13g2_fill_2 FILLER_19_330 ();
 sg13g2_fill_2 FILLER_19_344 ();
 sg13g2_fill_1 FILLER_19_346 ();
 sg13g2_decap_8 FILLER_19_351 ();
 sg13g2_decap_8 FILLER_19_358 ();
 sg13g2_decap_4 FILLER_19_365 ();
 sg13g2_fill_1 FILLER_19_369 ();
 sg13g2_decap_4 FILLER_19_373 ();
 sg13g2_fill_2 FILLER_19_382 ();
 sg13g2_fill_1 FILLER_19_384 ();
 sg13g2_fill_1 FILLER_19_396 ();
 sg13g2_decap_8 FILLER_19_407 ();
 sg13g2_decap_8 FILLER_19_414 ();
 sg13g2_decap_8 FILLER_19_421 ();
 sg13g2_fill_2 FILLER_19_428 ();
 sg13g2_decap_8 FILLER_20_0 ();
 sg13g2_decap_8 FILLER_20_7 ();
 sg13g2_decap_8 FILLER_20_14 ();
 sg13g2_decap_8 FILLER_20_21 ();
 sg13g2_decap_8 FILLER_20_28 ();
 sg13g2_decap_8 FILLER_20_35 ();
 sg13g2_decap_8 FILLER_20_42 ();
 sg13g2_decap_8 FILLER_20_49 ();
 sg13g2_decap_8 FILLER_20_56 ();
 sg13g2_decap_8 FILLER_20_63 ();
 sg13g2_decap_8 FILLER_20_70 ();
 sg13g2_decap_8 FILLER_20_77 ();
 sg13g2_decap_8 FILLER_20_84 ();
 sg13g2_decap_8 FILLER_20_91 ();
 sg13g2_decap_8 FILLER_20_98 ();
 sg13g2_decap_4 FILLER_20_105 ();
 sg13g2_fill_2 FILLER_20_109 ();
 sg13g2_fill_2 FILLER_20_135 ();
 sg13g2_fill_2 FILLER_20_157 ();
 sg13g2_fill_1 FILLER_20_159 ();
 sg13g2_decap_4 FILLER_20_164 ();
 sg13g2_fill_2 FILLER_20_177 ();
 sg13g2_decap_8 FILLER_20_184 ();
 sg13g2_decap_8 FILLER_20_191 ();
 sg13g2_decap_8 FILLER_20_198 ();
 sg13g2_decap_8 FILLER_20_205 ();
 sg13g2_decap_4 FILLER_20_212 ();
 sg13g2_fill_2 FILLER_20_216 ();
 sg13g2_decap_4 FILLER_20_222 ();
 sg13g2_fill_2 FILLER_20_226 ();
 sg13g2_fill_2 FILLER_20_262 ();
 sg13g2_fill_1 FILLER_20_264 ();
 sg13g2_decap_4 FILLER_20_269 ();
 sg13g2_fill_1 FILLER_20_273 ();
 sg13g2_decap_4 FILLER_20_282 ();
 sg13g2_fill_2 FILLER_20_286 ();
 sg13g2_decap_8 FILLER_20_293 ();
 sg13g2_decap_8 FILLER_20_300 ();
 sg13g2_fill_2 FILLER_20_307 ();
 sg13g2_fill_2 FILLER_20_317 ();
 sg13g2_fill_1 FILLER_20_319 ();
 sg13g2_fill_2 FILLER_20_328 ();
 sg13g2_fill_1 FILLER_20_330 ();
 sg13g2_decap_8 FILLER_20_344 ();
 sg13g2_decap_8 FILLER_20_351 ();
 sg13g2_decap_8 FILLER_20_358 ();
 sg13g2_decap_8 FILLER_20_365 ();
 sg13g2_decap_8 FILLER_20_372 ();
 sg13g2_decap_8 FILLER_20_379 ();
 sg13g2_fill_2 FILLER_20_386 ();
 sg13g2_decap_8 FILLER_20_408 ();
 sg13g2_decap_8 FILLER_20_415 ();
 sg13g2_decap_8 FILLER_20_422 ();
 sg13g2_fill_1 FILLER_20_429 ();
 sg13g2_decap_8 FILLER_21_0 ();
 sg13g2_decap_8 FILLER_21_7 ();
 sg13g2_decap_8 FILLER_21_14 ();
 sg13g2_decap_8 FILLER_21_21 ();
 sg13g2_decap_8 FILLER_21_28 ();
 sg13g2_decap_8 FILLER_21_35 ();
 sg13g2_decap_8 FILLER_21_42 ();
 sg13g2_decap_8 FILLER_21_49 ();
 sg13g2_decap_8 FILLER_21_56 ();
 sg13g2_decap_8 FILLER_21_63 ();
 sg13g2_decap_8 FILLER_21_70 ();
 sg13g2_decap_8 FILLER_21_77 ();
 sg13g2_decap_8 FILLER_21_84 ();
 sg13g2_decap_8 FILLER_21_91 ();
 sg13g2_decap_8 FILLER_21_98 ();
 sg13g2_decap_8 FILLER_21_105 ();
 sg13g2_fill_1 FILLER_21_112 ();
 sg13g2_decap_8 FILLER_21_162 ();
 sg13g2_decap_4 FILLER_21_169 ();
 sg13g2_fill_1 FILLER_21_185 ();
 sg13g2_fill_1 FILLER_21_193 ();
 sg13g2_fill_2 FILLER_21_199 ();
 sg13g2_fill_2 FILLER_21_205 ();
 sg13g2_fill_2 FILLER_21_211 ();
 sg13g2_decap_8 FILLER_21_218 ();
 sg13g2_fill_2 FILLER_21_270 ();
 sg13g2_decap_8 FILLER_21_323 ();
 sg13g2_decap_8 FILLER_21_330 ();
 sg13g2_decap_8 FILLER_21_337 ();
 sg13g2_fill_1 FILLER_21_344 ();
 sg13g2_decap_4 FILLER_21_354 ();
 sg13g2_fill_2 FILLER_21_367 ();
 sg13g2_decap_8 FILLER_21_385 ();
 sg13g2_fill_1 FILLER_21_392 ();
 sg13g2_decap_4 FILLER_21_403 ();
 sg13g2_decap_8 FILLER_21_411 ();
 sg13g2_decap_8 FILLER_21_418 ();
 sg13g2_decap_4 FILLER_21_425 ();
 sg13g2_fill_1 FILLER_21_429 ();
 sg13g2_decap_8 FILLER_22_0 ();
 sg13g2_decap_8 FILLER_22_7 ();
 sg13g2_decap_8 FILLER_22_14 ();
 sg13g2_decap_8 FILLER_22_21 ();
 sg13g2_decap_8 FILLER_22_28 ();
 sg13g2_decap_8 FILLER_22_35 ();
 sg13g2_decap_8 FILLER_22_42 ();
 sg13g2_decap_8 FILLER_22_49 ();
 sg13g2_decap_8 FILLER_22_56 ();
 sg13g2_decap_8 FILLER_22_63 ();
 sg13g2_decap_8 FILLER_22_70 ();
 sg13g2_decap_8 FILLER_22_77 ();
 sg13g2_decap_8 FILLER_22_84 ();
 sg13g2_decap_8 FILLER_22_91 ();
 sg13g2_decap_8 FILLER_22_98 ();
 sg13g2_decap_8 FILLER_22_105 ();
 sg13g2_fill_1 FILLER_22_117 ();
 sg13g2_fill_2 FILLER_22_123 ();
 sg13g2_fill_1 FILLER_22_148 ();
 sg13g2_decap_8 FILLER_22_157 ();
 sg13g2_decap_8 FILLER_22_164 ();
 sg13g2_fill_1 FILLER_22_171 ();
 sg13g2_fill_2 FILLER_22_176 ();
 sg13g2_fill_1 FILLER_22_178 ();
 sg13g2_fill_2 FILLER_22_184 ();
 sg13g2_fill_1 FILLER_22_192 ();
 sg13g2_fill_2 FILLER_22_251 ();
 sg13g2_decap_8 FILLER_22_265 ();
 sg13g2_decap_8 FILLER_22_272 ();
 sg13g2_decap_4 FILLER_22_279 ();
 sg13g2_fill_1 FILLER_22_294 ();
 sg13g2_decap_4 FILLER_22_302 ();
 sg13g2_fill_2 FILLER_22_306 ();
 sg13g2_fill_1 FILLER_22_312 ();
 sg13g2_fill_1 FILLER_22_326 ();
 sg13g2_decap_8 FILLER_22_331 ();
 sg13g2_fill_2 FILLER_22_338 ();
 sg13g2_fill_1 FILLER_22_340 ();
 sg13g2_decap_4 FILLER_22_345 ();
 sg13g2_fill_1 FILLER_22_361 ();
 sg13g2_fill_2 FILLER_22_367 ();
 sg13g2_fill_1 FILLER_22_386 ();
 sg13g2_fill_1 FILLER_22_391 ();
 sg13g2_fill_1 FILLER_22_396 ();
 sg13g2_fill_1 FILLER_22_405 ();
 sg13g2_decap_8 FILLER_22_411 ();
 sg13g2_decap_8 FILLER_22_418 ();
 sg13g2_decap_4 FILLER_22_425 ();
 sg13g2_fill_1 FILLER_22_429 ();
 sg13g2_decap_8 FILLER_23_0 ();
 sg13g2_decap_8 FILLER_23_7 ();
 sg13g2_decap_8 FILLER_23_14 ();
 sg13g2_decap_8 FILLER_23_21 ();
 sg13g2_decap_8 FILLER_23_28 ();
 sg13g2_decap_8 FILLER_23_35 ();
 sg13g2_decap_8 FILLER_23_42 ();
 sg13g2_decap_8 FILLER_23_49 ();
 sg13g2_decap_8 FILLER_23_56 ();
 sg13g2_decap_8 FILLER_23_63 ();
 sg13g2_decap_8 FILLER_23_70 ();
 sg13g2_decap_8 FILLER_23_77 ();
 sg13g2_decap_8 FILLER_23_84 ();
 sg13g2_decap_8 FILLER_23_91 ();
 sg13g2_decap_8 FILLER_23_98 ();
 sg13g2_decap_8 FILLER_23_105 ();
 sg13g2_decap_8 FILLER_23_112 ();
 sg13g2_decap_8 FILLER_23_119 ();
 sg13g2_decap_8 FILLER_23_130 ();
 sg13g2_fill_1 FILLER_23_137 ();
 sg13g2_decap_8 FILLER_23_143 ();
 sg13g2_decap_4 FILLER_23_150 ();
 sg13g2_decap_8 FILLER_23_159 ();
 sg13g2_decap_4 FILLER_23_174 ();
 sg13g2_fill_1 FILLER_23_199 ();
 sg13g2_fill_1 FILLER_23_204 ();
 sg13g2_fill_1 FILLER_23_210 ();
 sg13g2_fill_1 FILLER_23_216 ();
 sg13g2_decap_8 FILLER_23_225 ();
 sg13g2_decap_8 FILLER_23_232 ();
 sg13g2_decap_8 FILLER_23_239 ();
 sg13g2_decap_8 FILLER_23_246 ();
 sg13g2_fill_2 FILLER_23_253 ();
 sg13g2_fill_1 FILLER_23_255 ();
 sg13g2_fill_2 FILLER_23_263 ();
 sg13g2_decap_8 FILLER_23_273 ();
 sg13g2_fill_1 FILLER_23_280 ();
 sg13g2_decap_4 FILLER_23_301 ();
 sg13g2_decap_8 FILLER_23_309 ();
 sg13g2_decap_8 FILLER_23_316 ();
 sg13g2_fill_2 FILLER_23_323 ();
 sg13g2_fill_1 FILLER_23_325 ();
 sg13g2_decap_4 FILLER_23_330 ();
 sg13g2_fill_2 FILLER_23_343 ();
 sg13g2_fill_1 FILLER_23_345 ();
 sg13g2_decap_4 FILLER_23_361 ();
 sg13g2_fill_2 FILLER_23_375 ();
 sg13g2_fill_1 FILLER_23_382 ();
 sg13g2_fill_2 FILLER_23_388 ();
 sg13g2_decap_8 FILLER_23_421 ();
 sg13g2_fill_2 FILLER_23_428 ();
 sg13g2_decap_8 FILLER_24_0 ();
 sg13g2_decap_8 FILLER_24_7 ();
 sg13g2_decap_8 FILLER_24_14 ();
 sg13g2_decap_8 FILLER_24_21 ();
 sg13g2_decap_8 FILLER_24_28 ();
 sg13g2_decap_8 FILLER_24_35 ();
 sg13g2_decap_8 FILLER_24_42 ();
 sg13g2_decap_8 FILLER_24_49 ();
 sg13g2_decap_8 FILLER_24_56 ();
 sg13g2_decap_8 FILLER_24_63 ();
 sg13g2_decap_8 FILLER_24_70 ();
 sg13g2_decap_8 FILLER_24_77 ();
 sg13g2_decap_8 FILLER_24_84 ();
 sg13g2_decap_8 FILLER_24_91 ();
 sg13g2_decap_8 FILLER_24_98 ();
 sg13g2_decap_8 FILLER_24_105 ();
 sg13g2_fill_1 FILLER_24_112 ();
 sg13g2_decap_8 FILLER_24_116 ();
 sg13g2_fill_1 FILLER_24_123 ();
 sg13g2_decap_8 FILLER_24_128 ();
 sg13g2_decap_4 FILLER_24_135 ();
 sg13g2_fill_1 FILLER_24_139 ();
 sg13g2_fill_1 FILLER_24_145 ();
 sg13g2_decap_4 FILLER_24_189 ();
 sg13g2_fill_2 FILLER_24_193 ();
 sg13g2_decap_8 FILLER_24_221 ();
 sg13g2_decap_8 FILLER_24_228 ();
 sg13g2_decap_4 FILLER_24_235 ();
 sg13g2_fill_1 FILLER_24_239 ();
 sg13g2_decap_4 FILLER_24_254 ();
 sg13g2_decap_4 FILLER_24_267 ();
 sg13g2_fill_2 FILLER_24_271 ();
 sg13g2_decap_8 FILLER_24_288 ();
 sg13g2_decap_8 FILLER_24_295 ();
 sg13g2_decap_8 FILLER_24_302 ();
 sg13g2_fill_1 FILLER_24_309 ();
 sg13g2_decap_8 FILLER_24_314 ();
 sg13g2_fill_2 FILLER_24_358 ();
 sg13g2_fill_1 FILLER_24_360 ();
 sg13g2_fill_1 FILLER_24_387 ();
 sg13g2_decap_8 FILLER_24_392 ();
 sg13g2_decap_4 FILLER_24_399 ();
 sg13g2_fill_1 FILLER_24_403 ();
 sg13g2_decap_8 FILLER_24_408 ();
 sg13g2_decap_8 FILLER_24_415 ();
 sg13g2_decap_8 FILLER_24_422 ();
 sg13g2_fill_1 FILLER_24_429 ();
 sg13g2_decap_8 FILLER_25_0 ();
 sg13g2_decap_8 FILLER_25_7 ();
 sg13g2_decap_8 FILLER_25_14 ();
 sg13g2_decap_8 FILLER_25_21 ();
 sg13g2_decap_8 FILLER_25_28 ();
 sg13g2_decap_8 FILLER_25_35 ();
 sg13g2_decap_8 FILLER_25_42 ();
 sg13g2_decap_8 FILLER_25_49 ();
 sg13g2_decap_8 FILLER_25_56 ();
 sg13g2_decap_8 FILLER_25_63 ();
 sg13g2_decap_8 FILLER_25_70 ();
 sg13g2_decap_8 FILLER_25_77 ();
 sg13g2_decap_8 FILLER_25_84 ();
 sg13g2_decap_8 FILLER_25_91 ();
 sg13g2_decap_8 FILLER_25_98 ();
 sg13g2_decap_8 FILLER_25_105 ();
 sg13g2_decap_8 FILLER_25_112 ();
 sg13g2_decap_8 FILLER_25_119 ();
 sg13g2_decap_8 FILLER_25_126 ();
 sg13g2_decap_4 FILLER_25_133 ();
 sg13g2_fill_2 FILLER_25_137 ();
 sg13g2_fill_2 FILLER_25_151 ();
 sg13g2_fill_1 FILLER_25_153 ();
 sg13g2_decap_8 FILLER_25_163 ();
 sg13g2_fill_1 FILLER_25_170 ();
 sg13g2_decap_8 FILLER_25_175 ();
 sg13g2_decap_8 FILLER_25_182 ();
 sg13g2_fill_2 FILLER_25_189 ();
 sg13g2_fill_2 FILLER_25_198 ();
 sg13g2_fill_2 FILLER_25_204 ();
 sg13g2_decap_8 FILLER_25_218 ();
 sg13g2_decap_8 FILLER_25_225 ();
 sg13g2_decap_8 FILLER_25_232 ();
 sg13g2_decap_4 FILLER_25_259 ();
 sg13g2_decap_8 FILLER_25_267 ();
 sg13g2_decap_4 FILLER_25_274 ();
 sg13g2_decap_8 FILLER_25_284 ();
 sg13g2_decap_8 FILLER_25_291 ();
 sg13g2_decap_4 FILLER_25_298 ();
 sg13g2_decap_4 FILLER_25_323 ();
 sg13g2_fill_2 FILLER_25_327 ();
 sg13g2_decap_4 FILLER_25_338 ();
 sg13g2_decap_4 FILLER_25_357 ();
 sg13g2_fill_1 FILLER_25_361 ();
 sg13g2_fill_2 FILLER_25_366 ();
 sg13g2_fill_2 FILLER_25_376 ();
 sg13g2_fill_1 FILLER_25_378 ();
 sg13g2_decap_8 FILLER_25_386 ();
 sg13g2_decap_8 FILLER_25_393 ();
 sg13g2_decap_8 FILLER_25_400 ();
 sg13g2_decap_8 FILLER_25_407 ();
 sg13g2_decap_8 FILLER_25_414 ();
 sg13g2_decap_8 FILLER_25_421 ();
 sg13g2_fill_2 FILLER_25_428 ();
 sg13g2_decap_8 FILLER_26_0 ();
 sg13g2_decap_8 FILLER_26_7 ();
 sg13g2_decap_8 FILLER_26_14 ();
 sg13g2_decap_8 FILLER_26_21 ();
 sg13g2_decap_8 FILLER_26_28 ();
 sg13g2_decap_8 FILLER_26_35 ();
 sg13g2_decap_8 FILLER_26_42 ();
 sg13g2_decap_8 FILLER_26_49 ();
 sg13g2_decap_8 FILLER_26_56 ();
 sg13g2_decap_8 FILLER_26_63 ();
 sg13g2_decap_8 FILLER_26_70 ();
 sg13g2_decap_8 FILLER_26_77 ();
 sg13g2_decap_8 FILLER_26_84 ();
 sg13g2_decap_8 FILLER_26_91 ();
 sg13g2_decap_8 FILLER_26_98 ();
 sg13g2_fill_2 FILLER_26_105 ();
 sg13g2_decap_8 FILLER_26_133 ();
 sg13g2_fill_2 FILLER_26_140 ();
 sg13g2_fill_1 FILLER_26_142 ();
 sg13g2_decap_8 FILLER_26_159 ();
 sg13g2_decap_8 FILLER_26_166 ();
 sg13g2_fill_2 FILLER_26_173 ();
 sg13g2_decap_8 FILLER_26_197 ();
 sg13g2_fill_2 FILLER_26_204 ();
 sg13g2_decap_8 FILLER_26_214 ();
 sg13g2_decap_8 FILLER_26_221 ();
 sg13g2_fill_2 FILLER_26_247 ();
 sg13g2_fill_2 FILLER_26_254 ();
 sg13g2_fill_1 FILLER_26_256 ();
 sg13g2_fill_2 FILLER_26_267 ();
 sg13g2_fill_2 FILLER_26_277 ();
 sg13g2_decap_8 FILLER_26_287 ();
 sg13g2_decap_8 FILLER_26_294 ();
 sg13g2_fill_2 FILLER_26_301 ();
 sg13g2_fill_1 FILLER_26_317 ();
 sg13g2_decap_8 FILLER_26_328 ();
 sg13g2_decap_8 FILLER_26_335 ();
 sg13g2_decap_8 FILLER_26_342 ();
 sg13g2_decap_4 FILLER_26_349 ();
 sg13g2_fill_2 FILLER_26_353 ();
 sg13g2_fill_2 FILLER_26_383 ();
 sg13g2_fill_1 FILLER_26_398 ();
 sg13g2_decap_8 FILLER_26_404 ();
 sg13g2_decap_8 FILLER_26_411 ();
 sg13g2_decap_8 FILLER_26_418 ();
 sg13g2_decap_4 FILLER_26_425 ();
 sg13g2_fill_1 FILLER_26_429 ();
 sg13g2_decap_8 FILLER_27_0 ();
 sg13g2_decap_8 FILLER_27_7 ();
 sg13g2_decap_8 FILLER_27_14 ();
 sg13g2_decap_8 FILLER_27_21 ();
 sg13g2_decap_8 FILLER_27_28 ();
 sg13g2_decap_8 FILLER_27_35 ();
 sg13g2_decap_8 FILLER_27_42 ();
 sg13g2_decap_8 FILLER_27_49 ();
 sg13g2_decap_8 FILLER_27_56 ();
 sg13g2_decap_8 FILLER_27_63 ();
 sg13g2_decap_8 FILLER_27_70 ();
 sg13g2_decap_8 FILLER_27_77 ();
 sg13g2_decap_8 FILLER_27_84 ();
 sg13g2_decap_8 FILLER_27_91 ();
 sg13g2_decap_8 FILLER_27_98 ();
 sg13g2_decap_4 FILLER_27_105 ();
 sg13g2_fill_2 FILLER_27_109 ();
 sg13g2_fill_1 FILLER_27_119 ();
 sg13g2_fill_1 FILLER_27_124 ();
 sg13g2_fill_1 FILLER_27_151 ();
 sg13g2_fill_2 FILLER_27_155 ();
 sg13g2_fill_1 FILLER_27_169 ();
 sg13g2_fill_2 FILLER_27_175 ();
 sg13g2_decap_8 FILLER_27_205 ();
 sg13g2_decap_8 FILLER_27_212 ();
 sg13g2_decap_8 FILLER_27_219 ();
 sg13g2_fill_1 FILLER_27_226 ();
 sg13g2_fill_2 FILLER_27_236 ();
 sg13g2_decap_4 FILLER_27_243 ();
 sg13g2_fill_2 FILLER_27_254 ();
 sg13g2_fill_2 FILLER_27_260 ();
 sg13g2_fill_1 FILLER_27_262 ();
 sg13g2_fill_2 FILLER_27_267 ();
 sg13g2_fill_1 FILLER_27_269 ();
 sg13g2_fill_2 FILLER_27_278 ();
 sg13g2_decap_4 FILLER_27_293 ();
 sg13g2_decap_8 FILLER_27_301 ();
 sg13g2_decap_4 FILLER_27_308 ();
 sg13g2_fill_1 FILLER_27_312 ();
 sg13g2_decap_8 FILLER_27_322 ();
 sg13g2_fill_1 FILLER_27_341 ();
 sg13g2_fill_1 FILLER_27_353 ();
 sg13g2_fill_1 FILLER_27_378 ();
 sg13g2_fill_2 FILLER_27_387 ();
 sg13g2_decap_8 FILLER_27_415 ();
 sg13g2_decap_8 FILLER_27_422 ();
 sg13g2_fill_1 FILLER_27_429 ();
 sg13g2_decap_8 FILLER_28_0 ();
 sg13g2_decap_8 FILLER_28_7 ();
 sg13g2_decap_8 FILLER_28_14 ();
 sg13g2_decap_8 FILLER_28_21 ();
 sg13g2_decap_8 FILLER_28_28 ();
 sg13g2_decap_8 FILLER_28_35 ();
 sg13g2_decap_8 FILLER_28_42 ();
 sg13g2_decap_8 FILLER_28_49 ();
 sg13g2_decap_8 FILLER_28_56 ();
 sg13g2_decap_8 FILLER_28_63 ();
 sg13g2_decap_8 FILLER_28_70 ();
 sg13g2_decap_8 FILLER_28_77 ();
 sg13g2_decap_8 FILLER_28_84 ();
 sg13g2_decap_8 FILLER_28_91 ();
 sg13g2_decap_8 FILLER_28_98 ();
 sg13g2_decap_4 FILLER_28_115 ();
 sg13g2_fill_2 FILLER_28_125 ();
 sg13g2_fill_1 FILLER_28_127 ();
 sg13g2_decap_8 FILLER_28_136 ();
 sg13g2_fill_2 FILLER_28_143 ();
 sg13g2_decap_8 FILLER_28_150 ();
 sg13g2_decap_8 FILLER_28_157 ();
 sg13g2_decap_4 FILLER_28_164 ();
 sg13g2_fill_1 FILLER_28_168 ();
 sg13g2_fill_1 FILLER_28_174 ();
 sg13g2_fill_1 FILLER_28_180 ();
 sg13g2_fill_2 FILLER_28_191 ();
 sg13g2_decap_8 FILLER_28_197 ();
 sg13g2_fill_1 FILLER_28_213 ();
 sg13g2_decap_8 FILLER_28_219 ();
 sg13g2_fill_2 FILLER_28_226 ();
 sg13g2_fill_1 FILLER_28_228 ();
 sg13g2_decap_8 FILLER_28_234 ();
 sg13g2_fill_2 FILLER_28_241 ();
 sg13g2_fill_1 FILLER_28_243 ();
 sg13g2_decap_4 FILLER_28_249 ();
 sg13g2_decap_8 FILLER_28_262 ();
 sg13g2_decap_4 FILLER_28_269 ();
 sg13g2_fill_2 FILLER_28_273 ();
 sg13g2_fill_1 FILLER_28_279 ();
 sg13g2_fill_1 FILLER_28_285 ();
 sg13g2_decap_4 FILLER_28_300 ();
 sg13g2_fill_2 FILLER_28_304 ();
 sg13g2_fill_2 FILLER_28_312 ();
 sg13g2_fill_1 FILLER_28_314 ();
 sg13g2_decap_4 FILLER_28_320 ();
 sg13g2_fill_2 FILLER_28_324 ();
 sg13g2_fill_1 FILLER_28_358 ();
 sg13g2_fill_1 FILLER_28_363 ();
 sg13g2_fill_1 FILLER_28_369 ();
 sg13g2_decap_4 FILLER_28_403 ();
 sg13g2_fill_1 FILLER_28_407 ();
 sg13g2_decap_8 FILLER_28_412 ();
 sg13g2_decap_8 FILLER_28_419 ();
 sg13g2_decap_4 FILLER_28_426 ();
 sg13g2_decap_8 FILLER_29_0 ();
 sg13g2_decap_8 FILLER_29_7 ();
 sg13g2_decap_8 FILLER_29_14 ();
 sg13g2_decap_8 FILLER_29_21 ();
 sg13g2_decap_8 FILLER_29_28 ();
 sg13g2_decap_8 FILLER_29_35 ();
 sg13g2_decap_8 FILLER_29_42 ();
 sg13g2_decap_8 FILLER_29_49 ();
 sg13g2_decap_8 FILLER_29_56 ();
 sg13g2_decap_8 FILLER_29_63 ();
 sg13g2_decap_8 FILLER_29_70 ();
 sg13g2_decap_8 FILLER_29_77 ();
 sg13g2_decap_8 FILLER_29_84 ();
 sg13g2_decap_8 FILLER_29_91 ();
 sg13g2_decap_8 FILLER_29_98 ();
 sg13g2_decap_8 FILLER_29_105 ();
 sg13g2_decap_4 FILLER_29_112 ();
 sg13g2_fill_1 FILLER_29_116 ();
 sg13g2_fill_1 FILLER_29_125 ();
 sg13g2_fill_1 FILLER_29_135 ();
 sg13g2_fill_2 FILLER_29_150 ();
 sg13g2_fill_1 FILLER_29_152 ();
 sg13g2_decap_8 FILLER_29_157 ();
 sg13g2_decap_8 FILLER_29_164 ();
 sg13g2_decap_8 FILLER_29_171 ();
 sg13g2_fill_1 FILLER_29_178 ();
 sg13g2_fill_1 FILLER_29_190 ();
 sg13g2_fill_1 FILLER_29_196 ();
 sg13g2_fill_2 FILLER_29_227 ();
 sg13g2_fill_1 FILLER_29_229 ();
 sg13g2_decap_8 FILLER_29_235 ();
 sg13g2_decap_4 FILLER_29_242 ();
 sg13g2_fill_1 FILLER_29_256 ();
 sg13g2_fill_1 FILLER_29_279 ();
 sg13g2_fill_1 FILLER_29_285 ();
 sg13g2_decap_8 FILLER_29_294 ();
 sg13g2_decap_8 FILLER_29_301 ();
 sg13g2_decap_4 FILLER_29_308 ();
 sg13g2_decap_8 FILLER_29_327 ();
 sg13g2_fill_2 FILLER_29_334 ();
 sg13g2_fill_1 FILLER_29_336 ();
 sg13g2_decap_8 FILLER_29_345 ();
 sg13g2_fill_2 FILLER_29_352 ();
 sg13g2_fill_1 FILLER_29_354 ();
 sg13g2_fill_2 FILLER_29_384 ();
 sg13g2_decap_8 FILLER_29_390 ();
 sg13g2_decap_8 FILLER_29_397 ();
 sg13g2_decap_8 FILLER_29_404 ();
 sg13g2_decap_8 FILLER_29_411 ();
 sg13g2_decap_8 FILLER_29_418 ();
 sg13g2_decap_4 FILLER_29_425 ();
 sg13g2_fill_1 FILLER_29_429 ();
 sg13g2_decap_8 FILLER_30_0 ();
 sg13g2_decap_8 FILLER_30_7 ();
 sg13g2_decap_8 FILLER_30_14 ();
 sg13g2_decap_8 FILLER_30_21 ();
 sg13g2_decap_8 FILLER_30_28 ();
 sg13g2_decap_8 FILLER_30_35 ();
 sg13g2_decap_8 FILLER_30_42 ();
 sg13g2_decap_8 FILLER_30_49 ();
 sg13g2_decap_8 FILLER_30_56 ();
 sg13g2_decap_8 FILLER_30_63 ();
 sg13g2_decap_8 FILLER_30_70 ();
 sg13g2_decap_8 FILLER_30_77 ();
 sg13g2_decap_8 FILLER_30_84 ();
 sg13g2_decap_8 FILLER_30_91 ();
 sg13g2_decap_8 FILLER_30_98 ();
 sg13g2_decap_8 FILLER_30_105 ();
 sg13g2_decap_8 FILLER_30_112 ();
 sg13g2_fill_2 FILLER_30_119 ();
 sg13g2_fill_2 FILLER_30_129 ();
 sg13g2_fill_1 FILLER_30_131 ();
 sg13g2_fill_1 FILLER_30_140 ();
 sg13g2_fill_1 FILLER_30_146 ();
 sg13g2_fill_2 FILLER_30_173 ();
 sg13g2_fill_1 FILLER_30_183 ();
 sg13g2_fill_2 FILLER_30_192 ();
 sg13g2_fill_2 FILLER_30_207 ();
 sg13g2_fill_1 FILLER_30_209 ();
 sg13g2_decap_8 FILLER_30_219 ();
 sg13g2_decap_8 FILLER_30_226 ();
 sg13g2_decap_4 FILLER_30_237 ();
 sg13g2_fill_1 FILLER_30_241 ();
 sg13g2_fill_2 FILLER_30_247 ();
 sg13g2_fill_1 FILLER_30_259 ();
 sg13g2_fill_2 FILLER_30_287 ();
 sg13g2_fill_1 FILLER_30_289 ();
 sg13g2_fill_2 FILLER_30_303 ();
 sg13g2_fill_1 FILLER_30_305 ();
 sg13g2_fill_2 FILLER_30_323 ();
 sg13g2_fill_1 FILLER_30_325 ();
 sg13g2_fill_2 FILLER_30_329 ();
 sg13g2_decap_8 FILLER_30_344 ();
 sg13g2_decap_8 FILLER_30_404 ();
 sg13g2_decap_8 FILLER_30_411 ();
 sg13g2_decap_8 FILLER_30_418 ();
 sg13g2_decap_4 FILLER_30_425 ();
 sg13g2_fill_1 FILLER_30_429 ();
 sg13g2_decap_8 FILLER_31_0 ();
 sg13g2_decap_8 FILLER_31_7 ();
 sg13g2_decap_8 FILLER_31_14 ();
 sg13g2_decap_8 FILLER_31_21 ();
 sg13g2_decap_8 FILLER_31_28 ();
 sg13g2_decap_8 FILLER_31_35 ();
 sg13g2_decap_8 FILLER_31_42 ();
 sg13g2_decap_8 FILLER_31_49 ();
 sg13g2_decap_8 FILLER_31_56 ();
 sg13g2_decap_8 FILLER_31_63 ();
 sg13g2_decap_8 FILLER_31_70 ();
 sg13g2_decap_8 FILLER_31_77 ();
 sg13g2_decap_8 FILLER_31_84 ();
 sg13g2_decap_8 FILLER_31_91 ();
 sg13g2_decap_4 FILLER_31_98 ();
 sg13g2_fill_1 FILLER_31_102 ();
 sg13g2_fill_2 FILLER_31_138 ();
 sg13g2_decap_4 FILLER_31_178 ();
 sg13g2_fill_2 FILLER_31_187 ();
 sg13g2_fill_1 FILLER_31_194 ();
 sg13g2_fill_1 FILLER_31_200 ();
 sg13g2_fill_2 FILLER_31_209 ();
 sg13g2_fill_1 FILLER_31_211 ();
 sg13g2_fill_2 FILLER_31_218 ();
 sg13g2_decap_8 FILLER_31_226 ();
 sg13g2_fill_2 FILLER_31_268 ();
 sg13g2_decap_8 FILLER_31_289 ();
 sg13g2_fill_2 FILLER_31_296 ();
 sg13g2_fill_1 FILLER_31_298 ();
 sg13g2_fill_2 FILLER_31_312 ();
 sg13g2_decap_4 FILLER_31_318 ();
 sg13g2_fill_2 FILLER_31_326 ();
 sg13g2_fill_1 FILLER_31_348 ();
 sg13g2_decap_8 FILLER_31_373 ();
 sg13g2_fill_1 FILLER_31_397 ();
 sg13g2_decap_8 FILLER_31_402 ();
 sg13g2_decap_8 FILLER_31_409 ();
 sg13g2_decap_8 FILLER_31_416 ();
 sg13g2_decap_8 FILLER_31_423 ();
 sg13g2_decap_8 FILLER_32_0 ();
 sg13g2_decap_8 FILLER_32_7 ();
 sg13g2_decap_8 FILLER_32_14 ();
 sg13g2_decap_8 FILLER_32_21 ();
 sg13g2_decap_8 FILLER_32_28 ();
 sg13g2_decap_8 FILLER_32_35 ();
 sg13g2_decap_8 FILLER_32_42 ();
 sg13g2_decap_8 FILLER_32_49 ();
 sg13g2_decap_8 FILLER_32_56 ();
 sg13g2_decap_8 FILLER_32_63 ();
 sg13g2_decap_8 FILLER_32_70 ();
 sg13g2_decap_8 FILLER_32_77 ();
 sg13g2_decap_8 FILLER_32_84 ();
 sg13g2_decap_8 FILLER_32_91 ();
 sg13g2_decap_8 FILLER_32_98 ();
 sg13g2_decap_8 FILLER_32_105 ();
 sg13g2_decap_4 FILLER_32_112 ();
 sg13g2_fill_2 FILLER_32_116 ();
 sg13g2_decap_8 FILLER_32_122 ();
 sg13g2_fill_2 FILLER_32_133 ();
 sg13g2_fill_2 FILLER_32_141 ();
 sg13g2_fill_2 FILLER_32_147 ();
 sg13g2_fill_1 FILLER_32_149 ();
 sg13g2_fill_2 FILLER_32_154 ();
 sg13g2_fill_2 FILLER_32_161 ();
 sg13g2_fill_1 FILLER_32_168 ();
 sg13g2_fill_1 FILLER_32_177 ();
 sg13g2_decap_8 FILLER_32_214 ();
 sg13g2_decap_8 FILLER_32_221 ();
 sg13g2_decap_4 FILLER_32_228 ();
 sg13g2_fill_2 FILLER_32_232 ();
 sg13g2_fill_1 FILLER_32_243 ();
 sg13g2_decap_8 FILLER_32_249 ();
 sg13g2_fill_1 FILLER_32_256 ();
 sg13g2_decap_8 FILLER_32_262 ();
 sg13g2_decap_4 FILLER_32_269 ();
 sg13g2_decap_8 FILLER_32_277 ();
 sg13g2_decap_8 FILLER_32_284 ();
 sg13g2_decap_8 FILLER_32_291 ();
 sg13g2_decap_4 FILLER_32_298 ();
 sg13g2_fill_2 FILLER_32_307 ();
 sg13g2_decap_8 FILLER_32_330 ();
 sg13g2_decap_8 FILLER_32_337 ();
 sg13g2_decap_4 FILLER_32_344 ();
 sg13g2_fill_2 FILLER_32_348 ();
 sg13g2_decap_8 FILLER_32_378 ();
 sg13g2_decap_8 FILLER_32_385 ();
 sg13g2_decap_8 FILLER_32_392 ();
 sg13g2_decap_8 FILLER_32_399 ();
 sg13g2_decap_8 FILLER_32_406 ();
 sg13g2_decap_8 FILLER_32_413 ();
 sg13g2_decap_8 FILLER_32_420 ();
 sg13g2_fill_2 FILLER_32_427 ();
 sg13g2_fill_1 FILLER_32_429 ();
 sg13g2_decap_8 FILLER_33_0 ();
 sg13g2_decap_8 FILLER_33_7 ();
 sg13g2_decap_8 FILLER_33_14 ();
 sg13g2_decap_8 FILLER_33_21 ();
 sg13g2_decap_8 FILLER_33_28 ();
 sg13g2_decap_8 FILLER_33_35 ();
 sg13g2_decap_8 FILLER_33_42 ();
 sg13g2_decap_8 FILLER_33_49 ();
 sg13g2_decap_8 FILLER_33_56 ();
 sg13g2_decap_8 FILLER_33_63 ();
 sg13g2_decap_8 FILLER_33_70 ();
 sg13g2_decap_8 FILLER_33_77 ();
 sg13g2_decap_8 FILLER_33_84 ();
 sg13g2_decap_8 FILLER_33_91 ();
 sg13g2_decap_8 FILLER_33_98 ();
 sg13g2_decap_8 FILLER_33_105 ();
 sg13g2_decap_8 FILLER_33_112 ();
 sg13g2_decap_8 FILLER_33_119 ();
 sg13g2_decap_8 FILLER_33_126 ();
 sg13g2_fill_1 FILLER_33_133 ();
 sg13g2_decap_8 FILLER_33_151 ();
 sg13g2_fill_1 FILLER_33_158 ();
 sg13g2_decap_8 FILLER_33_172 ();
 sg13g2_decap_4 FILLER_33_179 ();
 sg13g2_fill_2 FILLER_33_183 ();
 sg13g2_decap_8 FILLER_33_189 ();
 sg13g2_decap_8 FILLER_33_196 ();
 sg13g2_decap_8 FILLER_33_203 ();
 sg13g2_fill_2 FILLER_33_210 ();
 sg13g2_decap_8 FILLER_33_225 ();
 sg13g2_fill_1 FILLER_33_232 ();
 sg13g2_decap_4 FILLER_33_237 ();
 sg13g2_fill_2 FILLER_33_245 ();
 sg13g2_fill_1 FILLER_33_247 ();
 sg13g2_fill_1 FILLER_33_286 ();
 sg13g2_fill_1 FILLER_33_292 ();
 sg13g2_fill_1 FILLER_33_312 ();
 sg13g2_decap_8 FILLER_33_318 ();
 sg13g2_fill_1 FILLER_33_325 ();
 sg13g2_decap_8 FILLER_33_333 ();
 sg13g2_decap_8 FILLER_33_340 ();
 sg13g2_decap_8 FILLER_33_347 ();
 sg13g2_decap_8 FILLER_33_354 ();
 sg13g2_decap_8 FILLER_33_361 ();
 sg13g2_decap_8 FILLER_33_368 ();
 sg13g2_decap_8 FILLER_33_401 ();
 sg13g2_decap_8 FILLER_33_408 ();
 sg13g2_decap_8 FILLER_33_415 ();
 sg13g2_decap_8 FILLER_33_422 ();
 sg13g2_fill_1 FILLER_33_429 ();
 sg13g2_decap_8 FILLER_34_0 ();
 sg13g2_decap_8 FILLER_34_7 ();
 sg13g2_decap_8 FILLER_34_14 ();
 sg13g2_decap_8 FILLER_34_21 ();
 sg13g2_decap_8 FILLER_34_28 ();
 sg13g2_decap_8 FILLER_34_35 ();
 sg13g2_decap_8 FILLER_34_42 ();
 sg13g2_decap_8 FILLER_34_49 ();
 sg13g2_decap_8 FILLER_34_56 ();
 sg13g2_decap_8 FILLER_34_63 ();
 sg13g2_decap_8 FILLER_34_70 ();
 sg13g2_decap_8 FILLER_34_77 ();
 sg13g2_decap_8 FILLER_34_84 ();
 sg13g2_fill_2 FILLER_34_91 ();
 sg13g2_fill_1 FILLER_34_93 ();
 sg13g2_fill_1 FILLER_34_124 ();
 sg13g2_fill_1 FILLER_34_143 ();
 sg13g2_decap_8 FILLER_34_148 ();
 sg13g2_decap_8 FILLER_34_155 ();
 sg13g2_fill_2 FILLER_34_162 ();
 sg13g2_decap_4 FILLER_34_178 ();
 sg13g2_fill_1 FILLER_34_182 ();
 sg13g2_decap_8 FILLER_34_191 ();
 sg13g2_decap_8 FILLER_34_198 ();
 sg13g2_decap_8 FILLER_34_205 ();
 sg13g2_decap_4 FILLER_34_212 ();
 sg13g2_fill_2 FILLER_34_216 ();
 sg13g2_fill_1 FILLER_34_231 ();
 sg13g2_fill_2 FILLER_34_259 ();
 sg13g2_fill_2 FILLER_34_266 ();
 sg13g2_fill_1 FILLER_34_281 ();
 sg13g2_fill_1 FILLER_34_313 ();
 sg13g2_fill_1 FILLER_34_318 ();
 sg13g2_fill_2 FILLER_34_324 ();
 sg13g2_fill_1 FILLER_34_336 ();
 sg13g2_fill_2 FILLER_34_341 ();
 sg13g2_fill_1 FILLER_34_343 ();
 sg13g2_decap_4 FILLER_34_351 ();
 sg13g2_fill_1 FILLER_34_355 ();
 sg13g2_decap_8 FILLER_34_361 ();
 sg13g2_decap_8 FILLER_34_372 ();
 sg13g2_decap_4 FILLER_34_379 ();
 sg13g2_decap_4 FILLER_34_387 ();
 sg13g2_decap_8 FILLER_34_395 ();
 sg13g2_decap_8 FILLER_34_402 ();
 sg13g2_decap_8 FILLER_34_409 ();
 sg13g2_decap_8 FILLER_34_416 ();
 sg13g2_decap_8 FILLER_34_423 ();
 sg13g2_decap_8 FILLER_35_0 ();
 sg13g2_decap_8 FILLER_35_7 ();
 sg13g2_decap_8 FILLER_35_14 ();
 sg13g2_decap_8 FILLER_35_21 ();
 sg13g2_decap_8 FILLER_35_28 ();
 sg13g2_decap_8 FILLER_35_35 ();
 sg13g2_decap_8 FILLER_35_42 ();
 sg13g2_decap_8 FILLER_35_49 ();
 sg13g2_decap_8 FILLER_35_56 ();
 sg13g2_decap_8 FILLER_35_63 ();
 sg13g2_decap_8 FILLER_35_70 ();
 sg13g2_decap_8 FILLER_35_77 ();
 sg13g2_decap_8 FILLER_35_84 ();
 sg13g2_decap_8 FILLER_35_91 ();
 sg13g2_fill_2 FILLER_35_98 ();
 sg13g2_fill_1 FILLER_35_100 ();
 sg13g2_fill_1 FILLER_35_110 ();
 sg13g2_fill_1 FILLER_35_119 ();
 sg13g2_fill_1 FILLER_35_126 ();
 sg13g2_decap_8 FILLER_35_149 ();
 sg13g2_fill_1 FILLER_35_156 ();
 sg13g2_decap_8 FILLER_35_205 ();
 sg13g2_decap_4 FILLER_35_212 ();
 sg13g2_fill_2 FILLER_35_216 ();
 sg13g2_decap_4 FILLER_35_223 ();
 sg13g2_fill_2 FILLER_35_227 ();
 sg13g2_fill_2 FILLER_35_236 ();
 sg13g2_fill_1 FILLER_35_238 ();
 sg13g2_fill_2 FILLER_35_244 ();
 sg13g2_fill_1 FILLER_35_255 ();
 sg13g2_fill_2 FILLER_35_277 ();
 sg13g2_fill_1 FILLER_35_279 ();
 sg13g2_fill_1 FILLER_35_345 ();
 sg13g2_fill_1 FILLER_35_351 ();
 sg13g2_decap_8 FILLER_35_397 ();
 sg13g2_decap_8 FILLER_35_404 ();
 sg13g2_decap_8 FILLER_35_411 ();
 sg13g2_decap_8 FILLER_35_418 ();
 sg13g2_decap_4 FILLER_35_425 ();
 sg13g2_fill_1 FILLER_35_429 ();
 sg13g2_decap_8 FILLER_36_0 ();
 sg13g2_decap_8 FILLER_36_7 ();
 sg13g2_decap_8 FILLER_36_14 ();
 sg13g2_decap_8 FILLER_36_21 ();
 sg13g2_decap_8 FILLER_36_28 ();
 sg13g2_decap_8 FILLER_36_35 ();
 sg13g2_decap_8 FILLER_36_42 ();
 sg13g2_decap_8 FILLER_36_49 ();
 sg13g2_decap_8 FILLER_36_56 ();
 sg13g2_decap_8 FILLER_36_63 ();
 sg13g2_decap_8 FILLER_36_70 ();
 sg13g2_decap_8 FILLER_36_77 ();
 sg13g2_decap_8 FILLER_36_84 ();
 sg13g2_decap_8 FILLER_36_91 ();
 sg13g2_decap_8 FILLER_36_98 ();
 sg13g2_decap_8 FILLER_36_105 ();
 sg13g2_decap_8 FILLER_36_112 ();
 sg13g2_fill_1 FILLER_36_128 ();
 sg13g2_fill_1 FILLER_36_133 ();
 sg13g2_fill_1 FILLER_36_151 ();
 sg13g2_fill_2 FILLER_36_167 ();
 sg13g2_fill_1 FILLER_36_169 ();
 sg13g2_decap_8 FILLER_36_176 ();
 sg13g2_fill_2 FILLER_36_183 ();
 sg13g2_decap_8 FILLER_36_189 ();
 sg13g2_fill_1 FILLER_36_204 ();
 sg13g2_decap_8 FILLER_36_235 ();
 sg13g2_decap_8 FILLER_36_242 ();
 sg13g2_fill_2 FILLER_36_249 ();
 sg13g2_fill_1 FILLER_36_251 ();
 sg13g2_decap_8 FILLER_36_260 ();
 sg13g2_fill_1 FILLER_36_267 ();
 sg13g2_decap_8 FILLER_36_271 ();
 sg13g2_decap_8 FILLER_36_278 ();
 sg13g2_fill_1 FILLER_36_285 ();
 sg13g2_decap_8 FILLER_36_290 ();
 sg13g2_fill_1 FILLER_36_297 ();
 sg13g2_decap_4 FILLER_36_303 ();
 sg13g2_decap_8 FILLER_36_314 ();
 sg13g2_fill_2 FILLER_36_321 ();
 sg13g2_fill_1 FILLER_36_323 ();
 sg13g2_decap_8 FILLER_36_339 ();
 sg13g2_fill_1 FILLER_36_351 ();
 sg13g2_fill_2 FILLER_36_369 ();
 sg13g2_fill_1 FILLER_36_371 ();
 sg13g2_decap_8 FILLER_36_377 ();
 sg13g2_decap_8 FILLER_36_384 ();
 sg13g2_decap_8 FILLER_36_391 ();
 sg13g2_decap_8 FILLER_36_398 ();
 sg13g2_decap_8 FILLER_36_405 ();
 sg13g2_decap_8 FILLER_36_412 ();
 sg13g2_decap_8 FILLER_36_419 ();
 sg13g2_decap_4 FILLER_36_426 ();
 sg13g2_decap_8 FILLER_37_0 ();
 sg13g2_decap_8 FILLER_37_7 ();
 sg13g2_decap_8 FILLER_37_14 ();
 sg13g2_decap_8 FILLER_37_21 ();
 sg13g2_decap_8 FILLER_37_28 ();
 sg13g2_decap_8 FILLER_37_35 ();
 sg13g2_decap_8 FILLER_37_42 ();
 sg13g2_decap_8 FILLER_37_49 ();
 sg13g2_decap_8 FILLER_37_56 ();
 sg13g2_decap_8 FILLER_37_63 ();
 sg13g2_decap_8 FILLER_37_70 ();
 sg13g2_decap_8 FILLER_37_77 ();
 sg13g2_decap_8 FILLER_37_84 ();
 sg13g2_decap_8 FILLER_37_91 ();
 sg13g2_decap_8 FILLER_37_98 ();
 sg13g2_decap_4 FILLER_37_105 ();
 sg13g2_fill_2 FILLER_37_109 ();
 sg13g2_fill_1 FILLER_37_124 ();
 sg13g2_fill_1 FILLER_37_162 ();
 sg13g2_fill_1 FILLER_37_168 ();
 sg13g2_fill_2 FILLER_37_173 ();
 sg13g2_decap_8 FILLER_37_184 ();
 sg13g2_decap_8 FILLER_37_191 ();
 sg13g2_decap_8 FILLER_37_198 ();
 sg13g2_decap_8 FILLER_37_205 ();
 sg13g2_decap_4 FILLER_37_216 ();
 sg13g2_fill_1 FILLER_37_220 ();
 sg13g2_decap_8 FILLER_37_236 ();
 sg13g2_decap_8 FILLER_37_243 ();
 sg13g2_fill_2 FILLER_37_250 ();
 sg13g2_decap_4 FILLER_37_256 ();
 sg13g2_decap_8 FILLER_37_264 ();
 sg13g2_decap_8 FILLER_37_271 ();
 sg13g2_decap_4 FILLER_37_278 ();
 sg13g2_fill_1 FILLER_37_282 ();
 sg13g2_fill_2 FILLER_37_287 ();
 sg13g2_decap_8 FILLER_37_293 ();
 sg13g2_decap_8 FILLER_37_300 ();
 sg13g2_decap_8 FILLER_37_307 ();
 sg13g2_decap_8 FILLER_37_314 ();
 sg13g2_decap_4 FILLER_37_321 ();
 sg13g2_decap_4 FILLER_37_363 ();
 sg13g2_fill_1 FILLER_37_367 ();
 sg13g2_decap_8 FILLER_37_372 ();
 sg13g2_fill_1 FILLER_37_379 ();
 sg13g2_fill_2 FILLER_37_390 ();
 sg13g2_fill_1 FILLER_37_392 ();
 sg13g2_fill_2 FILLER_37_397 ();
 sg13g2_fill_2 FILLER_37_404 ();
 sg13g2_fill_1 FILLER_37_410 ();
 sg13g2_decap_8 FILLER_37_415 ();
 sg13g2_decap_8 FILLER_37_422 ();
 sg13g2_fill_1 FILLER_37_429 ();
 sg13g2_decap_8 FILLER_38_0 ();
 sg13g2_decap_8 FILLER_38_7 ();
 sg13g2_decap_8 FILLER_38_14 ();
 sg13g2_decap_8 FILLER_38_21 ();
 sg13g2_decap_8 FILLER_38_28 ();
 sg13g2_decap_8 FILLER_38_35 ();
 sg13g2_decap_8 FILLER_38_42 ();
 sg13g2_decap_8 FILLER_38_49 ();
 sg13g2_decap_8 FILLER_38_56 ();
 sg13g2_decap_8 FILLER_38_63 ();
 sg13g2_decap_8 FILLER_38_70 ();
 sg13g2_decap_8 FILLER_38_77 ();
 sg13g2_decap_8 FILLER_38_84 ();
 sg13g2_decap_8 FILLER_38_91 ();
 sg13g2_decap_4 FILLER_38_98 ();
 sg13g2_fill_1 FILLER_38_102 ();
 sg13g2_decap_8 FILLER_38_116 ();
 sg13g2_fill_2 FILLER_38_123 ();
 sg13g2_fill_1 FILLER_38_158 ();
 sg13g2_fill_1 FILLER_38_163 ();
 sg13g2_fill_2 FILLER_38_169 ();
 sg13g2_fill_1 FILLER_38_193 ();
 sg13g2_decap_8 FILLER_38_199 ();
 sg13g2_decap_4 FILLER_38_206 ();
 sg13g2_decap_8 FILLER_38_220 ();
 sg13g2_fill_1 FILLER_38_231 ();
 sg13g2_fill_2 FILLER_38_258 ();
 sg13g2_fill_2 FILLER_38_265 ();
 sg13g2_fill_2 FILLER_38_271 ();
 sg13g2_fill_1 FILLER_38_273 ();
 sg13g2_decap_8 FILLER_38_308 ();
 sg13g2_decap_4 FILLER_38_320 ();
 sg13g2_fill_2 FILLER_38_330 ();
 sg13g2_decap_4 FILLER_38_337 ();
 sg13g2_fill_1 FILLER_38_341 ();
 sg13g2_decap_8 FILLER_38_346 ();
 sg13g2_fill_2 FILLER_38_353 ();
 sg13g2_fill_1 FILLER_38_355 ();
 sg13g2_fill_1 FILLER_38_362 ();
 sg13g2_fill_2 FILLER_38_368 ();
 sg13g2_fill_1 FILLER_38_370 ();
 sg13g2_fill_2 FILLER_38_384 ();
 sg13g2_fill_1 FILLER_38_386 ();
 sg13g2_fill_2 FILLER_38_397 ();
 sg13g2_decap_4 FILLER_38_425 ();
 sg13g2_fill_1 FILLER_38_429 ();
 sg13g2_decap_8 FILLER_39_0 ();
 sg13g2_decap_8 FILLER_39_7 ();
 sg13g2_decap_8 FILLER_39_14 ();
 sg13g2_decap_8 FILLER_39_21 ();
 sg13g2_decap_8 FILLER_39_28 ();
 sg13g2_decap_8 FILLER_39_35 ();
 sg13g2_decap_8 FILLER_39_42 ();
 sg13g2_decap_8 FILLER_39_49 ();
 sg13g2_decap_8 FILLER_39_56 ();
 sg13g2_decap_8 FILLER_39_63 ();
 sg13g2_decap_8 FILLER_39_70 ();
 sg13g2_decap_8 FILLER_39_77 ();
 sg13g2_decap_8 FILLER_39_84 ();
 sg13g2_decap_4 FILLER_39_91 ();
 sg13g2_decap_8 FILLER_39_129 ();
 sg13g2_decap_8 FILLER_39_136 ();
 sg13g2_decap_4 FILLER_39_143 ();
 sg13g2_fill_1 FILLER_39_147 ();
 sg13g2_decap_8 FILLER_39_154 ();
 sg13g2_decap_8 FILLER_39_161 ();
 sg13g2_fill_2 FILLER_39_168 ();
 sg13g2_fill_1 FILLER_39_170 ();
 sg13g2_fill_1 FILLER_39_176 ();
 sg13g2_fill_1 FILLER_39_183 ();
 sg13g2_fill_1 FILLER_39_189 ();
 sg13g2_decap_8 FILLER_39_195 ();
 sg13g2_decap_8 FILLER_39_206 ();
 sg13g2_decap_8 FILLER_39_213 ();
 sg13g2_decap_8 FILLER_39_220 ();
 sg13g2_decap_8 FILLER_39_227 ();
 sg13g2_fill_2 FILLER_39_234 ();
 sg13g2_decap_8 FILLER_39_241 ();
 sg13g2_decap_8 FILLER_39_248 ();
 sg13g2_fill_1 FILLER_39_295 ();
 sg13g2_fill_1 FILLER_39_304 ();
 sg13g2_fill_2 FILLER_39_313 ();
 sg13g2_fill_1 FILLER_39_315 ();
 sg13g2_fill_1 FILLER_39_331 ();
 sg13g2_fill_2 FILLER_39_340 ();
 sg13g2_decap_4 FILLER_39_346 ();
 sg13g2_fill_2 FILLER_39_350 ();
 sg13g2_fill_2 FILLER_39_357 ();
 sg13g2_fill_2 FILLER_39_363 ();
 sg13g2_fill_1 FILLER_39_365 ();
 sg13g2_fill_1 FILLER_39_386 ();
 sg13g2_fill_2 FILLER_39_405 ();
 sg13g2_decap_8 FILLER_39_411 ();
 sg13g2_decap_8 FILLER_39_418 ();
 sg13g2_decap_4 FILLER_39_425 ();
 sg13g2_fill_1 FILLER_39_429 ();
 sg13g2_decap_8 FILLER_40_0 ();
 sg13g2_decap_8 FILLER_40_7 ();
 sg13g2_decap_8 FILLER_40_14 ();
 sg13g2_decap_8 FILLER_40_21 ();
 sg13g2_decap_8 FILLER_40_28 ();
 sg13g2_decap_8 FILLER_40_35 ();
 sg13g2_decap_8 FILLER_40_42 ();
 sg13g2_decap_8 FILLER_40_49 ();
 sg13g2_decap_8 FILLER_40_56 ();
 sg13g2_decap_8 FILLER_40_63 ();
 sg13g2_decap_8 FILLER_40_70 ();
 sg13g2_decap_8 FILLER_40_77 ();
 sg13g2_decap_8 FILLER_40_84 ();
 sg13g2_decap_8 FILLER_40_91 ();
 sg13g2_fill_2 FILLER_40_98 ();
 sg13g2_fill_1 FILLER_40_100 ();
 sg13g2_fill_1 FILLER_40_144 ();
 sg13g2_decap_8 FILLER_40_150 ();
 sg13g2_decap_8 FILLER_40_157 ();
 sg13g2_decap_8 FILLER_40_164 ();
 sg13g2_decap_8 FILLER_40_171 ();
 sg13g2_decap_4 FILLER_40_178 ();
 sg13g2_fill_1 FILLER_40_182 ();
 sg13g2_decap_4 FILLER_40_188 ();
 sg13g2_fill_1 FILLER_40_192 ();
 sg13g2_fill_2 FILLER_40_219 ();
 sg13g2_fill_2 FILLER_40_225 ();
 sg13g2_fill_1 FILLER_40_237 ();
 sg13g2_decap_4 FILLER_40_243 ();
 sg13g2_fill_1 FILLER_40_251 ();
 sg13g2_fill_2 FILLER_40_268 ();
 sg13g2_fill_1 FILLER_40_279 ();
 sg13g2_fill_2 FILLER_40_303 ();
 sg13g2_fill_2 FILLER_40_317 ();
 sg13g2_decap_8 FILLER_40_337 ();
 sg13g2_decap_8 FILLER_40_344 ();
 sg13g2_decap_8 FILLER_40_351 ();
 sg13g2_decap_8 FILLER_40_363 ();
 sg13g2_fill_2 FILLER_40_370 ();
 sg13g2_fill_1 FILLER_40_384 ();
 sg13g2_decap_8 FILLER_40_406 ();
 sg13g2_fill_1 FILLER_40_413 ();
 sg13g2_fill_2 FILLER_40_427 ();
 sg13g2_fill_1 FILLER_40_429 ();
 sg13g2_decap_8 FILLER_41_0 ();
 sg13g2_decap_8 FILLER_41_7 ();
 sg13g2_decap_8 FILLER_41_14 ();
 sg13g2_decap_8 FILLER_41_21 ();
 sg13g2_decap_8 FILLER_41_28 ();
 sg13g2_decap_8 FILLER_41_35 ();
 sg13g2_decap_8 FILLER_41_42 ();
 sg13g2_decap_8 FILLER_41_49 ();
 sg13g2_decap_8 FILLER_41_56 ();
 sg13g2_decap_8 FILLER_41_63 ();
 sg13g2_decap_8 FILLER_41_70 ();
 sg13g2_decap_8 FILLER_41_77 ();
 sg13g2_decap_8 FILLER_41_84 ();
 sg13g2_decap_8 FILLER_41_91 ();
 sg13g2_decap_8 FILLER_41_98 ();
 sg13g2_decap_8 FILLER_41_105 ();
 sg13g2_fill_1 FILLER_41_112 ();
 sg13g2_fill_1 FILLER_41_133 ();
 sg13g2_fill_2 FILLER_41_144 ();
 sg13g2_decap_4 FILLER_41_153 ();
 sg13g2_decap_4 FILLER_41_162 ();
 sg13g2_fill_1 FILLER_41_166 ();
 sg13g2_decap_8 FILLER_41_172 ();
 sg13g2_fill_1 FILLER_41_179 ();
 sg13g2_fill_1 FILLER_41_183 ();
 sg13g2_decap_8 FILLER_41_194 ();
 sg13g2_decap_8 FILLER_41_201 ();
 sg13g2_decap_8 FILLER_41_208 ();
 sg13g2_fill_2 FILLER_41_215 ();
 sg13g2_fill_1 FILLER_41_217 ();
 sg13g2_fill_2 FILLER_41_228 ();
 sg13g2_fill_2 FILLER_41_256 ();
 sg13g2_fill_1 FILLER_41_258 ();
 sg13g2_fill_2 FILLER_41_274 ();
 sg13g2_decap_4 FILLER_41_290 ();
 sg13g2_fill_1 FILLER_41_294 ();
 sg13g2_decap_8 FILLER_41_329 ();
 sg13g2_fill_2 FILLER_41_336 ();
 sg13g2_fill_1 FILLER_41_338 ();
 sg13g2_fill_1 FILLER_41_351 ();
 sg13g2_fill_1 FILLER_41_363 ();
 sg13g2_decap_8 FILLER_41_368 ();
 sg13g2_decap_4 FILLER_41_375 ();
 sg13g2_fill_1 FILLER_41_379 ();
 sg13g2_fill_1 FILLER_41_389 ();
 sg13g2_fill_2 FILLER_41_394 ();
 sg13g2_decap_8 FILLER_41_422 ();
 sg13g2_fill_1 FILLER_41_429 ();
 sg13g2_decap_8 FILLER_42_0 ();
 sg13g2_decap_8 FILLER_42_7 ();
 sg13g2_decap_8 FILLER_42_14 ();
 sg13g2_decap_8 FILLER_42_21 ();
 sg13g2_decap_8 FILLER_42_28 ();
 sg13g2_decap_8 FILLER_42_35 ();
 sg13g2_decap_8 FILLER_42_42 ();
 sg13g2_decap_8 FILLER_42_49 ();
 sg13g2_decap_8 FILLER_42_56 ();
 sg13g2_decap_8 FILLER_42_63 ();
 sg13g2_decap_8 FILLER_42_70 ();
 sg13g2_decap_8 FILLER_42_77 ();
 sg13g2_decap_8 FILLER_42_84 ();
 sg13g2_decap_8 FILLER_42_91 ();
 sg13g2_decap_8 FILLER_42_98 ();
 sg13g2_decap_8 FILLER_42_105 ();
 sg13g2_decap_4 FILLER_42_112 ();
 sg13g2_fill_1 FILLER_42_116 ();
 sg13g2_fill_1 FILLER_42_126 ();
 sg13g2_fill_1 FILLER_42_155 ();
 sg13g2_fill_2 FILLER_42_164 ();
 sg13g2_fill_1 FILLER_42_172 ();
 sg13g2_fill_2 FILLER_42_199 ();
 sg13g2_fill_1 FILLER_42_201 ();
 sg13g2_fill_2 FILLER_42_244 ();
 sg13g2_fill_1 FILLER_42_246 ();
 sg13g2_fill_2 FILLER_42_257 ();
 sg13g2_fill_1 FILLER_42_264 ();
 sg13g2_fill_1 FILLER_42_269 ();
 sg13g2_decap_8 FILLER_42_290 ();
 sg13g2_decap_4 FILLER_42_297 ();
 sg13g2_fill_2 FILLER_42_301 ();
 sg13g2_decap_8 FILLER_42_308 ();
 sg13g2_decap_8 FILLER_42_315 ();
 sg13g2_decap_8 FILLER_42_322 ();
 sg13g2_decap_8 FILLER_42_329 ();
 sg13g2_decap_4 FILLER_42_336 ();
 sg13g2_fill_1 FILLER_42_354 ();
 sg13g2_fill_1 FILLER_42_360 ();
 sg13g2_decap_8 FILLER_42_370 ();
 sg13g2_decap_8 FILLER_42_377 ();
 sg13g2_decap_8 FILLER_42_384 ();
 sg13g2_decap_8 FILLER_42_391 ();
 sg13g2_fill_2 FILLER_42_398 ();
 sg13g2_decap_8 FILLER_42_408 ();
 sg13g2_decap_8 FILLER_42_415 ();
 sg13g2_decap_8 FILLER_42_422 ();
 sg13g2_fill_1 FILLER_42_429 ();
 sg13g2_decap_8 FILLER_43_0 ();
 sg13g2_decap_8 FILLER_43_7 ();
 sg13g2_decap_8 FILLER_43_14 ();
 sg13g2_decap_8 FILLER_43_21 ();
 sg13g2_decap_8 FILLER_43_28 ();
 sg13g2_decap_8 FILLER_43_35 ();
 sg13g2_decap_8 FILLER_43_42 ();
 sg13g2_decap_8 FILLER_43_49 ();
 sg13g2_decap_8 FILLER_43_56 ();
 sg13g2_decap_8 FILLER_43_63 ();
 sg13g2_decap_8 FILLER_43_70 ();
 sg13g2_decap_8 FILLER_43_77 ();
 sg13g2_decap_8 FILLER_43_84 ();
 sg13g2_decap_8 FILLER_43_91 ();
 sg13g2_decap_8 FILLER_43_98 ();
 sg13g2_decap_8 FILLER_43_105 ();
 sg13g2_decap_8 FILLER_43_112 ();
 sg13g2_fill_1 FILLER_43_119 ();
 sg13g2_fill_1 FILLER_43_151 ();
 sg13g2_fill_1 FILLER_43_157 ();
 sg13g2_decap_8 FILLER_43_173 ();
 sg13g2_fill_2 FILLER_43_185 ();
 sg13g2_decap_8 FILLER_43_195 ();
 sg13g2_decap_8 FILLER_43_202 ();
 sg13g2_decap_4 FILLER_43_213 ();
 sg13g2_decap_8 FILLER_43_237 ();
 sg13g2_decap_8 FILLER_43_244 ();
 sg13g2_fill_2 FILLER_43_251 ();
 sg13g2_decap_4 FILLER_43_292 ();
 sg13g2_fill_1 FILLER_43_296 ();
 sg13g2_fill_1 FILLER_43_307 ();
 sg13g2_decap_4 FILLER_43_313 ();
 sg13g2_fill_2 FILLER_43_317 ();
 sg13g2_decap_4 FILLER_43_323 ();
 sg13g2_fill_1 FILLER_43_327 ();
 sg13g2_decap_8 FILLER_43_357 ();
 sg13g2_fill_1 FILLER_43_364 ();
 sg13g2_decap_8 FILLER_43_374 ();
 sg13g2_decap_8 FILLER_43_400 ();
 sg13g2_decap_8 FILLER_43_407 ();
 sg13g2_decap_8 FILLER_43_414 ();
 sg13g2_decap_8 FILLER_43_421 ();
 sg13g2_fill_2 FILLER_43_428 ();
 sg13g2_decap_8 FILLER_44_0 ();
 sg13g2_decap_8 FILLER_44_7 ();
 sg13g2_decap_8 FILLER_44_14 ();
 sg13g2_decap_8 FILLER_44_21 ();
 sg13g2_decap_8 FILLER_44_28 ();
 sg13g2_decap_8 FILLER_44_35 ();
 sg13g2_decap_8 FILLER_44_42 ();
 sg13g2_decap_8 FILLER_44_49 ();
 sg13g2_decap_8 FILLER_44_56 ();
 sg13g2_decap_8 FILLER_44_63 ();
 sg13g2_decap_8 FILLER_44_70 ();
 sg13g2_decap_8 FILLER_44_77 ();
 sg13g2_decap_8 FILLER_44_84 ();
 sg13g2_decap_8 FILLER_44_91 ();
 sg13g2_decap_8 FILLER_44_98 ();
 sg13g2_decap_8 FILLER_44_105 ();
 sg13g2_decap_8 FILLER_44_112 ();
 sg13g2_decap_8 FILLER_44_119 ();
 sg13g2_decap_4 FILLER_44_126 ();
 sg13g2_fill_2 FILLER_44_130 ();
 sg13g2_fill_1 FILLER_44_141 ();
 sg13g2_fill_2 FILLER_44_147 ();
 sg13g2_fill_1 FILLER_44_155 ();
 sg13g2_fill_2 FILLER_44_162 ();
 sg13g2_fill_1 FILLER_44_169 ();
 sg13g2_fill_2 FILLER_44_174 ();
 sg13g2_fill_2 FILLER_44_181 ();
 sg13g2_fill_1 FILLER_44_183 ();
 sg13g2_fill_2 FILLER_44_190 ();
 sg13g2_decap_4 FILLER_44_196 ();
 sg13g2_fill_2 FILLER_44_200 ();
 sg13g2_fill_2 FILLER_44_212 ();
 sg13g2_fill_1 FILLER_44_224 ();
 sg13g2_decap_8 FILLER_44_230 ();
 sg13g2_decap_4 FILLER_44_237 ();
 sg13g2_fill_2 FILLER_44_241 ();
 sg13g2_fill_1 FILLER_44_267 ();
 sg13g2_fill_1 FILLER_44_272 ();
 sg13g2_fill_1 FILLER_44_277 ();
 sg13g2_fill_2 FILLER_44_282 ();
 sg13g2_fill_1 FILLER_44_292 ();
 sg13g2_decap_8 FILLER_44_303 ();
 sg13g2_decap_4 FILLER_44_310 ();
 sg13g2_fill_1 FILLER_44_314 ();
 sg13g2_fill_1 FILLER_44_328 ();
 sg13g2_fill_2 FILLER_44_334 ();
 sg13g2_fill_1 FILLER_44_341 ();
 sg13g2_fill_2 FILLER_44_357 ();
 sg13g2_decap_8 FILLER_44_372 ();
 sg13g2_fill_1 FILLER_44_379 ();
 sg13g2_decap_8 FILLER_44_386 ();
 sg13g2_fill_2 FILLER_44_399 ();
 sg13g2_fill_2 FILLER_44_427 ();
 sg13g2_fill_1 FILLER_44_429 ();
 sg13g2_decap_8 FILLER_45_0 ();
 sg13g2_decap_8 FILLER_45_7 ();
 sg13g2_decap_8 FILLER_45_14 ();
 sg13g2_decap_8 FILLER_45_21 ();
 sg13g2_decap_8 FILLER_45_28 ();
 sg13g2_decap_8 FILLER_45_35 ();
 sg13g2_decap_8 FILLER_45_42 ();
 sg13g2_decap_8 FILLER_45_49 ();
 sg13g2_decap_8 FILLER_45_56 ();
 sg13g2_decap_8 FILLER_45_63 ();
 sg13g2_decap_8 FILLER_45_70 ();
 sg13g2_decap_8 FILLER_45_77 ();
 sg13g2_decap_8 FILLER_45_84 ();
 sg13g2_decap_8 FILLER_45_91 ();
 sg13g2_fill_2 FILLER_45_98 ();
 sg13g2_decap_8 FILLER_45_126 ();
 sg13g2_decap_8 FILLER_45_148 ();
 sg13g2_fill_2 FILLER_45_155 ();
 sg13g2_fill_1 FILLER_45_157 ();
 sg13g2_decap_8 FILLER_45_163 ();
 sg13g2_fill_2 FILLER_45_170 ();
 sg13g2_decap_4 FILLER_45_175 ();
 sg13g2_fill_2 FILLER_45_179 ();
 sg13g2_fill_2 FILLER_45_216 ();
 sg13g2_fill_1 FILLER_45_218 ();
 sg13g2_decap_4 FILLER_45_226 ();
 sg13g2_decap_8 FILLER_45_238 ();
 sg13g2_fill_2 FILLER_45_245 ();
 sg13g2_decap_8 FILLER_45_276 ();
 sg13g2_decap_4 FILLER_45_292 ();
 sg13g2_fill_1 FILLER_45_301 ();
 sg13g2_fill_2 FILLER_45_306 ();
 sg13g2_fill_1 FILLER_45_308 ();
 sg13g2_fill_1 FILLER_45_329 ();
 sg13g2_fill_1 FILLER_45_344 ();
 sg13g2_decap_8 FILLER_45_349 ();
 sg13g2_fill_2 FILLER_45_356 ();
 sg13g2_fill_2 FILLER_45_372 ();
 sg13g2_fill_1 FILLER_45_379 ();
 sg13g2_fill_2 FILLER_45_385 ();
 sg13g2_fill_1 FILLER_45_392 ();
 sg13g2_decap_8 FILLER_45_398 ();
 sg13g2_decap_4 FILLER_45_405 ();
 sg13g2_fill_1 FILLER_45_409 ();
 sg13g2_fill_2 FILLER_45_427 ();
 sg13g2_fill_1 FILLER_45_429 ();
 sg13g2_decap_8 FILLER_46_0 ();
 sg13g2_decap_8 FILLER_46_7 ();
 sg13g2_decap_8 FILLER_46_14 ();
 sg13g2_decap_8 FILLER_46_21 ();
 sg13g2_decap_8 FILLER_46_28 ();
 sg13g2_decap_8 FILLER_46_35 ();
 sg13g2_decap_8 FILLER_46_42 ();
 sg13g2_decap_8 FILLER_46_49 ();
 sg13g2_decap_8 FILLER_46_56 ();
 sg13g2_decap_8 FILLER_46_63 ();
 sg13g2_decap_8 FILLER_46_70 ();
 sg13g2_decap_8 FILLER_46_77 ();
 sg13g2_decap_8 FILLER_46_84 ();
 sg13g2_decap_8 FILLER_46_91 ();
 sg13g2_fill_2 FILLER_46_98 ();
 sg13g2_decap_8 FILLER_46_140 ();
 sg13g2_decap_8 FILLER_46_147 ();
 sg13g2_decap_8 FILLER_46_154 ();
 sg13g2_decap_8 FILLER_46_161 ();
 sg13g2_fill_1 FILLER_46_168 ();
 sg13g2_decap_8 FILLER_46_188 ();
 sg13g2_decap_8 FILLER_46_195 ();
 sg13g2_decap_8 FILLER_46_202 ();
 sg13g2_decap_4 FILLER_46_209 ();
 sg13g2_decap_8 FILLER_46_218 ();
 sg13g2_decap_8 FILLER_46_225 ();
 sg13g2_fill_1 FILLER_46_232 ();
 sg13g2_fill_1 FILLER_46_269 ();
 sg13g2_fill_1 FILLER_46_274 ();
 sg13g2_decap_8 FILLER_46_281 ();
 sg13g2_decap_8 FILLER_46_288 ();
 sg13g2_decap_8 FILLER_46_295 ();
 sg13g2_fill_2 FILLER_46_323 ();
 sg13g2_fill_1 FILLER_46_325 ();
 sg13g2_decap_4 FILLER_46_332 ();
 sg13g2_fill_1 FILLER_46_346 ();
 sg13g2_decap_4 FILLER_46_358 ();
 sg13g2_fill_2 FILLER_46_389 ();
 sg13g2_fill_1 FILLER_46_391 ();
 sg13g2_fill_2 FILLER_46_395 ();
 sg13g2_decap_8 FILLER_46_404 ();
 sg13g2_decap_8 FILLER_46_416 ();
 sg13g2_decap_8 FILLER_46_423 ();
 sg13g2_decap_8 FILLER_47_0 ();
 sg13g2_decap_8 FILLER_47_7 ();
 sg13g2_decap_8 FILLER_47_14 ();
 sg13g2_decap_8 FILLER_47_21 ();
 sg13g2_decap_8 FILLER_47_28 ();
 sg13g2_decap_8 FILLER_47_35 ();
 sg13g2_decap_8 FILLER_47_42 ();
 sg13g2_decap_8 FILLER_47_49 ();
 sg13g2_decap_8 FILLER_47_56 ();
 sg13g2_decap_8 FILLER_47_63 ();
 sg13g2_decap_8 FILLER_47_70 ();
 sg13g2_decap_8 FILLER_47_77 ();
 sg13g2_decap_8 FILLER_47_84 ();
 sg13g2_decap_8 FILLER_47_91 ();
 sg13g2_decap_8 FILLER_47_98 ();
 sg13g2_decap_4 FILLER_47_105 ();
 sg13g2_fill_2 FILLER_47_109 ();
 sg13g2_fill_1 FILLER_47_115 ();
 sg13g2_decap_8 FILLER_47_130 ();
 sg13g2_decap_8 FILLER_47_137 ();
 sg13g2_decap_8 FILLER_47_144 ();
 sg13g2_decap_8 FILLER_47_151 ();
 sg13g2_fill_2 FILLER_47_158 ();
 sg13g2_fill_1 FILLER_47_174 ();
 sg13g2_decap_8 FILLER_47_201 ();
 sg13g2_decap_8 FILLER_47_208 ();
 sg13g2_decap_4 FILLER_47_215 ();
 sg13g2_fill_1 FILLER_47_219 ();
 sg13g2_decap_4 FILLER_47_230 ();
 sg13g2_fill_2 FILLER_47_234 ();
 sg13g2_fill_2 FILLER_47_245 ();
 sg13g2_fill_1 FILLER_47_258 ();
 sg13g2_decap_8 FILLER_47_273 ();
 sg13g2_decap_8 FILLER_47_280 ();
 sg13g2_decap_8 FILLER_47_287 ();
 sg13g2_decap_8 FILLER_47_294 ();
 sg13g2_decap_8 FILLER_47_301 ();
 sg13g2_fill_2 FILLER_47_308 ();
 sg13g2_fill_1 FILLER_47_310 ();
 sg13g2_decap_8 FILLER_47_316 ();
 sg13g2_decap_8 FILLER_47_323 ();
 sg13g2_fill_1 FILLER_47_330 ();
 sg13g2_decap_8 FILLER_47_359 ();
 sg13g2_decap_4 FILLER_47_370 ();
 sg13g2_fill_1 FILLER_47_374 ();
 sg13g2_decap_4 FILLER_47_380 ();
 sg13g2_fill_1 FILLER_47_384 ();
 sg13g2_fill_1 FILLER_47_389 ();
 sg13g2_decap_8 FILLER_47_406 ();
 sg13g2_decap_8 FILLER_47_413 ();
 sg13g2_decap_8 FILLER_47_420 ();
 sg13g2_fill_2 FILLER_47_427 ();
 sg13g2_fill_1 FILLER_47_429 ();
 sg13g2_decap_8 FILLER_48_0 ();
 sg13g2_decap_8 FILLER_48_7 ();
 sg13g2_decap_8 FILLER_48_14 ();
 sg13g2_decap_8 FILLER_48_21 ();
 sg13g2_decap_8 FILLER_48_28 ();
 sg13g2_decap_8 FILLER_48_35 ();
 sg13g2_decap_8 FILLER_48_42 ();
 sg13g2_decap_8 FILLER_48_49 ();
 sg13g2_decap_8 FILLER_48_56 ();
 sg13g2_decap_8 FILLER_48_63 ();
 sg13g2_decap_8 FILLER_48_70 ();
 sg13g2_decap_8 FILLER_48_77 ();
 sg13g2_decap_8 FILLER_48_84 ();
 sg13g2_decap_8 FILLER_48_91 ();
 sg13g2_decap_8 FILLER_48_98 ();
 sg13g2_decap_8 FILLER_48_105 ();
 sg13g2_decap_8 FILLER_48_112 ();
 sg13g2_decap_4 FILLER_48_122 ();
 sg13g2_fill_1 FILLER_48_126 ();
 sg13g2_fill_2 FILLER_48_153 ();
 sg13g2_decap_8 FILLER_48_185 ();
 sg13g2_fill_2 FILLER_48_192 ();
 sg13g2_fill_2 FILLER_48_198 ();
 sg13g2_fill_1 FILLER_48_200 ();
 sg13g2_decap_4 FILLER_48_251 ();
 sg13g2_fill_2 FILLER_48_262 ();
 sg13g2_fill_2 FILLER_48_268 ();
 sg13g2_fill_1 FILLER_48_270 ();
 sg13g2_decap_4 FILLER_48_301 ();
 sg13g2_decap_4 FILLER_48_310 ();
 sg13g2_fill_1 FILLER_48_314 ();
 sg13g2_decap_8 FILLER_48_328 ();
 sg13g2_fill_2 FILLER_48_335 ();
 sg13g2_decap_4 FILLER_48_345 ();
 sg13g2_fill_1 FILLER_48_349 ();
 sg13g2_fill_1 FILLER_48_356 ();
 sg13g2_decap_8 FILLER_48_364 ();
 sg13g2_fill_1 FILLER_48_371 ();
 sg13g2_fill_1 FILLER_48_385 ();
 sg13g2_decap_4 FILLER_48_396 ();
 sg13g2_fill_1 FILLER_48_400 ();
 sg13g2_decap_8 FILLER_48_405 ();
 sg13g2_decap_4 FILLER_48_412 ();
 sg13g2_fill_1 FILLER_48_416 ();
 sg13g2_decap_8 FILLER_49_0 ();
 sg13g2_decap_8 FILLER_49_7 ();
 sg13g2_decap_8 FILLER_49_14 ();
 sg13g2_decap_8 FILLER_49_21 ();
 sg13g2_decap_8 FILLER_49_28 ();
 sg13g2_decap_8 FILLER_49_35 ();
 sg13g2_decap_8 FILLER_49_42 ();
 sg13g2_decap_8 FILLER_49_49 ();
 sg13g2_decap_8 FILLER_49_56 ();
 sg13g2_decap_8 FILLER_49_63 ();
 sg13g2_decap_8 FILLER_49_70 ();
 sg13g2_decap_8 FILLER_49_77 ();
 sg13g2_decap_4 FILLER_49_84 ();
 sg13g2_fill_2 FILLER_49_88 ();
 sg13g2_decap_8 FILLER_49_120 ();
 sg13g2_fill_1 FILLER_49_127 ();
 sg13g2_fill_1 FILLER_49_133 ();
 sg13g2_fill_1 FILLER_49_142 ();
 sg13g2_decap_8 FILLER_49_174 ();
 sg13g2_decap_4 FILLER_49_181 ();
 sg13g2_decap_4 FILLER_49_190 ();
 sg13g2_fill_1 FILLER_49_194 ();
 sg13g2_decap_8 FILLER_49_199 ();
 sg13g2_fill_2 FILLER_49_206 ();
 sg13g2_fill_1 FILLER_49_208 ();
 sg13g2_decap_8 FILLER_49_213 ();
 sg13g2_decap_4 FILLER_49_220 ();
 sg13g2_fill_1 FILLER_49_224 ();
 sg13g2_decap_4 FILLER_49_230 ();
 sg13g2_fill_1 FILLER_49_243 ();
 sg13g2_fill_1 FILLER_49_272 ();
 sg13g2_fill_2 FILLER_49_282 ();
 sg13g2_fill_1 FILLER_49_284 ();
 sg13g2_fill_2 FILLER_49_293 ();
 sg13g2_fill_1 FILLER_49_313 ();
 sg13g2_fill_1 FILLER_49_319 ();
 sg13g2_decap_4 FILLER_49_338 ();
 sg13g2_decap_4 FILLER_49_347 ();
 sg13g2_fill_2 FILLER_49_351 ();
 sg13g2_decap_4 FILLER_49_367 ();
 sg13g2_fill_1 FILLER_49_371 ();
 sg13g2_fill_2 FILLER_49_388 ();
 sg13g2_fill_1 FILLER_49_390 ();
 sg13g2_decap_4 FILLER_49_399 ();
 sg13g2_fill_1 FILLER_49_403 ();
 sg13g2_decap_8 FILLER_50_0 ();
 sg13g2_decap_8 FILLER_50_7 ();
 sg13g2_decap_8 FILLER_50_14 ();
 sg13g2_decap_8 FILLER_50_21 ();
 sg13g2_decap_8 FILLER_50_28 ();
 sg13g2_decap_8 FILLER_50_35 ();
 sg13g2_decap_8 FILLER_50_42 ();
 sg13g2_decap_8 FILLER_50_49 ();
 sg13g2_decap_8 FILLER_50_56 ();
 sg13g2_decap_8 FILLER_50_63 ();
 sg13g2_decap_8 FILLER_50_70 ();
 sg13g2_decap_8 FILLER_50_77 ();
 sg13g2_fill_2 FILLER_50_84 ();
 sg13g2_fill_1 FILLER_50_86 ();
 sg13g2_fill_2 FILLER_50_117 ();
 sg13g2_decap_8 FILLER_50_137 ();
 sg13g2_decap_4 FILLER_50_144 ();
 sg13g2_decap_8 FILLER_50_152 ();
 sg13g2_decap_8 FILLER_50_159 ();
 sg13g2_decap_8 FILLER_50_166 ();
 sg13g2_decap_8 FILLER_50_173 ();
 sg13g2_decap_4 FILLER_50_180 ();
 sg13g2_fill_2 FILLER_50_184 ();
 sg13g2_fill_1 FILLER_50_225 ();
 sg13g2_fill_2 FILLER_50_241 ();
 sg13g2_fill_1 FILLER_50_248 ();
 sg13g2_fill_1 FILLER_50_267 ();
 sg13g2_decap_8 FILLER_50_273 ();
 sg13g2_decap_8 FILLER_50_280 ();
 sg13g2_fill_2 FILLER_50_287 ();
 sg13g2_fill_2 FILLER_50_302 ();
 sg13g2_fill_2 FILLER_50_312 ();
 sg13g2_fill_2 FILLER_50_322 ();
 sg13g2_fill_2 FILLER_50_328 ();
 sg13g2_fill_1 FILLER_50_330 ();
 sg13g2_fill_2 FILLER_50_351 ();
 sg13g2_fill_1 FILLER_50_366 ();
 sg13g2_decap_8 FILLER_50_380 ();
 sg13g2_fill_2 FILLER_50_390 ();
 sg13g2_fill_1 FILLER_50_392 ();
 sg13g2_fill_1 FILLER_50_398 ();
 sg13g2_decap_8 FILLER_50_404 ();
 sg13g2_decap_8 FILLER_50_415 ();
 sg13g2_decap_8 FILLER_50_422 ();
 sg13g2_fill_1 FILLER_50_429 ();
 sg13g2_decap_8 FILLER_51_0 ();
 sg13g2_decap_8 FILLER_51_7 ();
 sg13g2_decap_8 FILLER_51_14 ();
 sg13g2_decap_8 FILLER_51_21 ();
 sg13g2_decap_8 FILLER_51_28 ();
 sg13g2_decap_8 FILLER_51_35 ();
 sg13g2_decap_8 FILLER_51_42 ();
 sg13g2_decap_8 FILLER_51_49 ();
 sg13g2_decap_8 FILLER_51_56 ();
 sg13g2_decap_8 FILLER_51_63 ();
 sg13g2_decap_8 FILLER_51_70 ();
 sg13g2_decap_8 FILLER_51_77 ();
 sg13g2_decap_4 FILLER_51_84 ();
 sg13g2_decap_8 FILLER_51_93 ();
 sg13g2_decap_4 FILLER_51_100 ();
 sg13g2_decap_8 FILLER_51_108 ();
 sg13g2_decap_8 FILLER_51_115 ();
 sg13g2_fill_2 FILLER_51_122 ();
 sg13g2_fill_1 FILLER_51_124 ();
 sg13g2_decap_8 FILLER_51_134 ();
 sg13g2_decap_8 FILLER_51_141 ();
 sg13g2_decap_8 FILLER_51_148 ();
 sg13g2_fill_1 FILLER_51_155 ();
 sg13g2_fill_2 FILLER_51_161 ();
 sg13g2_decap_8 FILLER_51_190 ();
 sg13g2_fill_2 FILLER_51_197 ();
 sg13g2_fill_1 FILLER_51_199 ();
 sg13g2_fill_1 FILLER_51_211 ();
 sg13g2_decap_8 FILLER_51_220 ();
 sg13g2_decap_8 FILLER_51_227 ();
 sg13g2_decap_4 FILLER_51_234 ();
 sg13g2_fill_2 FILLER_51_238 ();
 sg13g2_decap_8 FILLER_51_245 ();
 sg13g2_decap_8 FILLER_51_252 ();
 sg13g2_fill_1 FILLER_51_259 ();
 sg13g2_decap_4 FILLER_51_269 ();
 sg13g2_decap_8 FILLER_51_277 ();
 sg13g2_fill_1 FILLER_51_284 ();
 sg13g2_decap_8 FILLER_51_288 ();
 sg13g2_decap_8 FILLER_51_295 ();
 sg13g2_decap_8 FILLER_51_302 ();
 sg13g2_decap_8 FILLER_51_309 ();
 sg13g2_decap_8 FILLER_51_316 ();
 sg13g2_decap_8 FILLER_51_323 ();
 sg13g2_decap_4 FILLER_51_330 ();
 sg13g2_fill_1 FILLER_51_334 ();
 sg13g2_decap_4 FILLER_51_346 ();
 sg13g2_fill_1 FILLER_51_350 ();
 sg13g2_fill_1 FILLER_51_372 ();
 sg13g2_decap_8 FILLER_51_379 ();
 sg13g2_decap_8 FILLER_51_418 ();
 sg13g2_decap_4 FILLER_51_425 ();
 sg13g2_fill_1 FILLER_51_429 ();
 sg13g2_decap_8 FILLER_52_0 ();
 sg13g2_decap_8 FILLER_52_7 ();
 sg13g2_decap_8 FILLER_52_14 ();
 sg13g2_decap_8 FILLER_52_21 ();
 sg13g2_decap_8 FILLER_52_28 ();
 sg13g2_decap_8 FILLER_52_35 ();
 sg13g2_decap_8 FILLER_52_42 ();
 sg13g2_decap_8 FILLER_52_49 ();
 sg13g2_decap_8 FILLER_52_56 ();
 sg13g2_decap_8 FILLER_52_63 ();
 sg13g2_decap_8 FILLER_52_70 ();
 sg13g2_decap_8 FILLER_52_77 ();
 sg13g2_decap_8 FILLER_52_84 ();
 sg13g2_fill_1 FILLER_52_91 ();
 sg13g2_fill_1 FILLER_52_131 ();
 sg13g2_fill_1 FILLER_52_158 ();
 sg13g2_fill_2 FILLER_52_185 ();
 sg13g2_fill_2 FILLER_52_190 ();
 sg13g2_decap_8 FILLER_52_226 ();
 sg13g2_decap_4 FILLER_52_233 ();
 sg13g2_decap_8 FILLER_52_245 ();
 sg13g2_fill_2 FILLER_52_252 ();
 sg13g2_fill_1 FILLER_52_254 ();
 sg13g2_decap_8 FILLER_52_260 ();
 sg13g2_fill_2 FILLER_52_267 ();
 sg13g2_fill_1 FILLER_52_269 ();
 sg13g2_decap_8 FILLER_52_280 ();
 sg13g2_fill_2 FILLER_52_287 ();
 sg13g2_fill_1 FILLER_52_289 ();
 sg13g2_fill_2 FILLER_52_294 ();
 sg13g2_fill_1 FILLER_52_304 ();
 sg13g2_fill_2 FILLER_52_313 ();
 sg13g2_fill_1 FILLER_52_315 ();
 sg13g2_decap_4 FILLER_52_321 ();
 sg13g2_fill_1 FILLER_52_325 ();
 sg13g2_fill_2 FILLER_52_337 ();
 sg13g2_fill_1 FILLER_52_343 ();
 sg13g2_fill_1 FILLER_52_379 ();
 sg13g2_decap_8 FILLER_52_385 ();
 sg13g2_fill_2 FILLER_52_392 ();
 sg13g2_decap_8 FILLER_52_408 ();
 sg13g2_decap_8 FILLER_52_415 ();
 sg13g2_decap_8 FILLER_52_422 ();
 sg13g2_fill_1 FILLER_52_429 ();
 sg13g2_decap_8 FILLER_53_0 ();
 sg13g2_decap_8 FILLER_53_7 ();
 sg13g2_decap_8 FILLER_53_14 ();
 sg13g2_decap_8 FILLER_53_21 ();
 sg13g2_decap_8 FILLER_53_28 ();
 sg13g2_decap_8 FILLER_53_35 ();
 sg13g2_decap_8 FILLER_53_42 ();
 sg13g2_decap_8 FILLER_53_49 ();
 sg13g2_decap_8 FILLER_53_56 ();
 sg13g2_decap_8 FILLER_53_63 ();
 sg13g2_decap_8 FILLER_53_70 ();
 sg13g2_decap_8 FILLER_53_77 ();
 sg13g2_decap_8 FILLER_53_84 ();
 sg13g2_fill_1 FILLER_53_122 ();
 sg13g2_fill_1 FILLER_53_128 ();
 sg13g2_fill_1 FILLER_53_139 ();
 sg13g2_fill_1 FILLER_53_144 ();
 sg13g2_decap_4 FILLER_53_197 ();
 sg13g2_fill_1 FILLER_53_201 ();
 sg13g2_fill_2 FILLER_53_227 ();
 sg13g2_fill_1 FILLER_53_229 ();
 sg13g2_fill_2 FILLER_53_235 ();
 sg13g2_fill_1 FILLER_53_237 ();
 sg13g2_fill_2 FILLER_53_319 ();
 sg13g2_fill_2 FILLER_53_326 ();
 sg13g2_fill_1 FILLER_53_345 ();
 sg13g2_fill_2 FILLER_53_351 ();
 sg13g2_fill_1 FILLER_53_353 ();
 sg13g2_decap_4 FILLER_53_361 ();
 sg13g2_decap_4 FILLER_53_369 ();
 sg13g2_decap_4 FILLER_53_379 ();
 sg13g2_fill_1 FILLER_53_383 ();
 sg13g2_fill_2 FILLER_53_409 ();
 sg13g2_fill_1 FILLER_53_411 ();
 sg13g2_decap_8 FILLER_53_417 ();
 sg13g2_decap_4 FILLER_53_424 ();
 sg13g2_fill_2 FILLER_53_428 ();
 sg13g2_decap_8 FILLER_54_0 ();
 sg13g2_decap_8 FILLER_54_7 ();
 sg13g2_decap_8 FILLER_54_14 ();
 sg13g2_decap_8 FILLER_54_21 ();
 sg13g2_decap_8 FILLER_54_28 ();
 sg13g2_decap_8 FILLER_54_35 ();
 sg13g2_decap_8 FILLER_54_42 ();
 sg13g2_decap_8 FILLER_54_49 ();
 sg13g2_decap_8 FILLER_54_56 ();
 sg13g2_decap_8 FILLER_54_63 ();
 sg13g2_decap_8 FILLER_54_70 ();
 sg13g2_decap_8 FILLER_54_77 ();
 sg13g2_decap_8 FILLER_54_84 ();
 sg13g2_decap_8 FILLER_54_91 ();
 sg13g2_fill_1 FILLER_54_98 ();
 sg13g2_decap_4 FILLER_54_103 ();
 sg13g2_fill_2 FILLER_54_107 ();
 sg13g2_decap_8 FILLER_54_140 ();
 sg13g2_decap_4 FILLER_54_147 ();
 sg13g2_fill_2 FILLER_54_151 ();
 sg13g2_decap_4 FILLER_54_157 ();
 sg13g2_fill_1 FILLER_54_161 ();
 sg13g2_fill_1 FILLER_54_166 ();
 sg13g2_fill_2 FILLER_54_180 ();
 sg13g2_decap_8 FILLER_54_186 ();
 sg13g2_decap_8 FILLER_54_193 ();
 sg13g2_decap_4 FILLER_54_200 ();
 sg13g2_fill_1 FILLER_54_204 ();
 sg13g2_fill_1 FILLER_54_220 ();
 sg13g2_decap_4 FILLER_54_230 ();
 sg13g2_fill_2 FILLER_54_234 ();
 sg13g2_fill_1 FILLER_54_245 ();
 sg13g2_fill_2 FILLER_54_263 ();
 sg13g2_fill_1 FILLER_54_265 ();
 sg13g2_fill_2 FILLER_54_307 ();
 sg13g2_fill_1 FILLER_54_314 ();
 sg13g2_fill_1 FILLER_54_320 ();
 sg13g2_decap_8 FILLER_54_333 ();
 sg13g2_fill_2 FILLER_54_346 ();
 sg13g2_fill_2 FILLER_54_356 ();
 sg13g2_fill_2 FILLER_54_363 ();
 sg13g2_fill_1 FILLER_54_365 ();
 sg13g2_fill_1 FILLER_54_373 ();
 sg13g2_fill_2 FILLER_54_392 ();
 sg13g2_fill_2 FILLER_54_412 ();
 sg13g2_fill_1 FILLER_54_414 ();
 sg13g2_decap_8 FILLER_54_419 ();
 sg13g2_decap_4 FILLER_54_426 ();
 sg13g2_decap_8 FILLER_55_0 ();
 sg13g2_decap_8 FILLER_55_7 ();
 sg13g2_decap_8 FILLER_55_14 ();
 sg13g2_decap_8 FILLER_55_21 ();
 sg13g2_decap_8 FILLER_55_28 ();
 sg13g2_decap_8 FILLER_55_35 ();
 sg13g2_decap_8 FILLER_55_42 ();
 sg13g2_decap_8 FILLER_55_49 ();
 sg13g2_decap_8 FILLER_55_56 ();
 sg13g2_decap_8 FILLER_55_63 ();
 sg13g2_decap_8 FILLER_55_70 ();
 sg13g2_decap_8 FILLER_55_77 ();
 sg13g2_decap_8 FILLER_55_84 ();
 sg13g2_fill_2 FILLER_55_91 ();
 sg13g2_decap_8 FILLER_55_123 ();
 sg13g2_decap_8 FILLER_55_130 ();
 sg13g2_fill_1 FILLER_55_137 ();
 sg13g2_decap_8 FILLER_55_142 ();
 sg13g2_decap_8 FILLER_55_149 ();
 sg13g2_decap_8 FILLER_55_156 ();
 sg13g2_decap_8 FILLER_55_163 ();
 sg13g2_decap_4 FILLER_55_170 ();
 sg13g2_fill_2 FILLER_55_174 ();
 sg13g2_decap_8 FILLER_55_180 ();
 sg13g2_decap_8 FILLER_55_187 ();
 sg13g2_decap_4 FILLER_55_194 ();
 sg13g2_fill_2 FILLER_55_198 ();
 sg13g2_decap_8 FILLER_55_212 ();
 sg13g2_decap_8 FILLER_55_219 ();
 sg13g2_fill_2 FILLER_55_226 ();
 sg13g2_decap_4 FILLER_55_250 ();
 sg13g2_fill_2 FILLER_55_254 ();
 sg13g2_decap_4 FILLER_55_261 ();
 sg13g2_fill_2 FILLER_55_269 ();
 sg13g2_fill_1 FILLER_55_271 ();
 sg13g2_fill_1 FILLER_55_281 ();
 sg13g2_fill_1 FILLER_55_287 ();
 sg13g2_decap_4 FILLER_55_293 ();
 sg13g2_fill_1 FILLER_55_297 ();
 sg13g2_fill_1 FILLER_55_319 ();
 sg13g2_decap_8 FILLER_55_328 ();
 sg13g2_decap_8 FILLER_55_335 ();
 sg13g2_decap_8 FILLER_55_342 ();
 sg13g2_fill_1 FILLER_55_349 ();
 sg13g2_fill_2 FILLER_55_356 ();
 sg13g2_decap_8 FILLER_55_375 ();
 sg13g2_fill_2 FILLER_55_382 ();
 sg13g2_fill_1 FILLER_55_384 ();
 sg13g2_fill_1 FILLER_55_399 ();
 sg13g2_fill_1 FILLER_55_418 ();
 sg13g2_decap_8 FILLER_55_422 ();
 sg13g2_fill_1 FILLER_55_429 ();
 sg13g2_decap_8 FILLER_56_0 ();
 sg13g2_decap_8 FILLER_56_7 ();
 sg13g2_decap_8 FILLER_56_14 ();
 sg13g2_decap_8 FILLER_56_21 ();
 sg13g2_decap_8 FILLER_56_28 ();
 sg13g2_decap_8 FILLER_56_35 ();
 sg13g2_decap_8 FILLER_56_42 ();
 sg13g2_decap_8 FILLER_56_49 ();
 sg13g2_decap_8 FILLER_56_56 ();
 sg13g2_decap_8 FILLER_56_63 ();
 sg13g2_decap_8 FILLER_56_70 ();
 sg13g2_decap_8 FILLER_56_77 ();
 sg13g2_fill_2 FILLER_56_84 ();
 sg13g2_decap_4 FILLER_56_96 ();
 sg13g2_fill_2 FILLER_56_100 ();
 sg13g2_decap_4 FILLER_56_106 ();
 sg13g2_fill_1 FILLER_56_110 ();
 sg13g2_decap_8 FILLER_56_115 ();
 sg13g2_decap_4 FILLER_56_122 ();
 sg13g2_fill_1 FILLER_56_126 ();
 sg13g2_fill_2 FILLER_56_142 ();
 sg13g2_decap_8 FILLER_56_149 ();
 sg13g2_decap_8 FILLER_56_161 ();
 sg13g2_decap_4 FILLER_56_168 ();
 sg13g2_fill_2 FILLER_56_172 ();
 sg13g2_decap_8 FILLER_56_210 ();
 sg13g2_decap_8 FILLER_56_247 ();
 sg13g2_fill_2 FILLER_56_254 ();
 sg13g2_fill_1 FILLER_56_256 ();
 sg13g2_decap_8 FILLER_56_261 ();
 sg13g2_fill_1 FILLER_56_268 ();
 sg13g2_decap_4 FILLER_56_273 ();
 sg13g2_decap_8 FILLER_56_286 ();
 sg13g2_decap_8 FILLER_56_293 ();
 sg13g2_fill_2 FILLER_56_300 ();
 sg13g2_fill_1 FILLER_56_302 ();
 sg13g2_decap_8 FILLER_56_316 ();
 sg13g2_decap_8 FILLER_56_323 ();
 sg13g2_decap_8 FILLER_56_330 ();
 sg13g2_decap_8 FILLER_56_337 ();
 sg13g2_decap_8 FILLER_56_344 ();
 sg13g2_decap_4 FILLER_56_351 ();
 sg13g2_fill_2 FILLER_56_355 ();
 sg13g2_fill_1 FILLER_56_364 ();
 sg13g2_decap_8 FILLER_56_371 ();
 sg13g2_fill_2 FILLER_56_394 ();
 sg13g2_fill_1 FILLER_56_396 ();
 sg13g2_fill_2 FILLER_56_402 ();
 sg13g2_decap_8 FILLER_57_0 ();
 sg13g2_decap_8 FILLER_57_7 ();
 sg13g2_decap_8 FILLER_57_14 ();
 sg13g2_decap_8 FILLER_57_21 ();
 sg13g2_decap_8 FILLER_57_28 ();
 sg13g2_decap_8 FILLER_57_35 ();
 sg13g2_decap_8 FILLER_57_42 ();
 sg13g2_decap_8 FILLER_57_49 ();
 sg13g2_decap_8 FILLER_57_56 ();
 sg13g2_decap_8 FILLER_57_63 ();
 sg13g2_decap_8 FILLER_57_70 ();
 sg13g2_decap_4 FILLER_57_77 ();
 sg13g2_fill_2 FILLER_57_81 ();
 sg13g2_fill_2 FILLER_57_96 ();
 sg13g2_fill_1 FILLER_57_102 ();
 sg13g2_fill_1 FILLER_57_137 ();
 sg13g2_fill_2 FILLER_57_167 ();
 sg13g2_fill_1 FILLER_57_169 ();
 sg13g2_decap_8 FILLER_57_206 ();
 sg13g2_fill_1 FILLER_57_213 ();
 sg13g2_decap_8 FILLER_57_223 ();
 sg13g2_fill_2 FILLER_57_240 ();
 sg13g2_fill_1 FILLER_57_242 ();
 sg13g2_decap_8 FILLER_57_247 ();
 sg13g2_decap_8 FILLER_57_254 ();
 sg13g2_fill_2 FILLER_57_261 ();
 sg13g2_decap_4 FILLER_57_289 ();
 sg13g2_fill_2 FILLER_57_293 ();
 sg13g2_decap_8 FILLER_57_298 ();
 sg13g2_fill_2 FILLER_57_305 ();
 sg13g2_fill_1 FILLER_57_307 ();
 sg13g2_fill_1 FILLER_57_312 ();
 sg13g2_fill_2 FILLER_57_336 ();
 sg13g2_decap_4 FILLER_57_343 ();
 sg13g2_fill_1 FILLER_57_372 ();
 sg13g2_decap_4 FILLER_57_377 ();
 sg13g2_decap_4 FILLER_57_401 ();
 sg13g2_decap_8 FILLER_57_422 ();
 sg13g2_fill_1 FILLER_57_429 ();
 sg13g2_decap_8 FILLER_58_0 ();
 sg13g2_decap_8 FILLER_58_7 ();
 sg13g2_decap_8 FILLER_58_14 ();
 sg13g2_decap_8 FILLER_58_21 ();
 sg13g2_decap_8 FILLER_58_28 ();
 sg13g2_decap_8 FILLER_58_35 ();
 sg13g2_decap_8 FILLER_58_42 ();
 sg13g2_decap_8 FILLER_58_49 ();
 sg13g2_decap_8 FILLER_58_56 ();
 sg13g2_decap_8 FILLER_58_63 ();
 sg13g2_decap_8 FILLER_58_70 ();
 sg13g2_fill_2 FILLER_58_77 ();
 sg13g2_fill_1 FILLER_58_79 ();
 sg13g2_fill_2 FILLER_58_85 ();
 sg13g2_fill_1 FILLER_58_87 ();
 sg13g2_fill_1 FILLER_58_101 ();
 sg13g2_fill_1 FILLER_58_106 ();
 sg13g2_fill_1 FILLER_58_124 ();
 sg13g2_fill_1 FILLER_58_129 ();
 sg13g2_fill_1 FILLER_58_135 ();
 sg13g2_fill_1 FILLER_58_141 ();
 sg13g2_fill_1 FILLER_58_146 ();
 sg13g2_fill_1 FILLER_58_152 ();
 sg13g2_fill_2 FILLER_58_157 ();
 sg13g2_decap_4 FILLER_58_193 ();
 sg13g2_fill_1 FILLER_58_202 ();
 sg13g2_decap_8 FILLER_58_208 ();
 sg13g2_fill_2 FILLER_58_215 ();
 sg13g2_fill_1 FILLER_58_222 ();
 sg13g2_decap_8 FILLER_58_237 ();
 sg13g2_decap_8 FILLER_58_244 ();
 sg13g2_decap_8 FILLER_58_251 ();
 sg13g2_decap_4 FILLER_58_284 ();
 sg13g2_fill_1 FILLER_58_288 ();
 sg13g2_decap_8 FILLER_58_299 ();
 sg13g2_fill_1 FILLER_58_311 ();
 sg13g2_decap_4 FILLER_58_317 ();
 sg13g2_fill_1 FILLER_58_325 ();
 sg13g2_fill_2 FILLER_58_330 ();
 sg13g2_fill_1 FILLER_58_332 ();
 sg13g2_decap_4 FILLER_58_343 ();
 sg13g2_fill_1 FILLER_58_347 ();
 sg13g2_fill_1 FILLER_58_351 ();
 sg13g2_fill_2 FILLER_58_369 ();
 sg13g2_fill_2 FILLER_58_380 ();
 sg13g2_fill_1 FILLER_58_382 ();
 sg13g2_fill_2 FILLER_58_395 ();
 sg13g2_fill_1 FILLER_58_401 ();
 sg13g2_fill_2 FILLER_58_428 ();
 sg13g2_decap_8 FILLER_59_0 ();
 sg13g2_decap_8 FILLER_59_7 ();
 sg13g2_decap_8 FILLER_59_14 ();
 sg13g2_decap_8 FILLER_59_21 ();
 sg13g2_decap_8 FILLER_59_28 ();
 sg13g2_decap_8 FILLER_59_35 ();
 sg13g2_decap_8 FILLER_59_42 ();
 sg13g2_decap_8 FILLER_59_49 ();
 sg13g2_decap_8 FILLER_59_56 ();
 sg13g2_decap_8 FILLER_59_63 ();
 sg13g2_decap_8 FILLER_59_70 ();
 sg13g2_decap_8 FILLER_59_77 ();
 sg13g2_fill_2 FILLER_59_84 ();
 sg13g2_fill_1 FILLER_59_100 ();
 sg13g2_fill_1 FILLER_59_109 ();
 sg13g2_fill_2 FILLER_59_137 ();
 sg13g2_fill_2 FILLER_59_144 ();
 sg13g2_fill_1 FILLER_59_146 ();
 sg13g2_decap_8 FILLER_59_152 ();
 sg13g2_fill_1 FILLER_59_159 ();
 sg13g2_fill_2 FILLER_59_164 ();
 sg13g2_decap_8 FILLER_59_170 ();
 sg13g2_decap_8 FILLER_59_177 ();
 sg13g2_decap_8 FILLER_59_184 ();
 sg13g2_decap_8 FILLER_59_191 ();
 sg13g2_decap_8 FILLER_59_198 ();
 sg13g2_decap_4 FILLER_59_205 ();
 sg13g2_fill_1 FILLER_59_209 ();
 sg13g2_fill_2 FILLER_59_219 ();
 sg13g2_fill_1 FILLER_59_221 ();
 sg13g2_decap_8 FILLER_59_256 ();
 sg13g2_decap_4 FILLER_59_263 ();
 sg13g2_fill_1 FILLER_59_306 ();
 sg13g2_decap_4 FILLER_59_312 ();
 sg13g2_fill_2 FILLER_59_316 ();
 sg13g2_decap_4 FILLER_59_351 ();
 sg13g2_fill_1 FILLER_59_355 ();
 sg13g2_fill_1 FILLER_59_363 ();
 sg13g2_decap_8 FILLER_59_378 ();
 sg13g2_decap_8 FILLER_59_385 ();
 sg13g2_decap_8 FILLER_59_392 ();
 sg13g2_decap_4 FILLER_59_404 ();
 sg13g2_fill_1 FILLER_59_408 ();
 sg13g2_decap_8 FILLER_59_413 ();
 sg13g2_decap_4 FILLER_59_424 ();
 sg13g2_fill_2 FILLER_59_428 ();
 sg13g2_decap_8 FILLER_60_0 ();
 sg13g2_decap_8 FILLER_60_7 ();
 sg13g2_decap_8 FILLER_60_14 ();
 sg13g2_decap_8 FILLER_60_21 ();
 sg13g2_decap_8 FILLER_60_28 ();
 sg13g2_decap_8 FILLER_60_35 ();
 sg13g2_decap_8 FILLER_60_42 ();
 sg13g2_decap_8 FILLER_60_49 ();
 sg13g2_decap_8 FILLER_60_56 ();
 sg13g2_decap_8 FILLER_60_63 ();
 sg13g2_decap_8 FILLER_60_70 ();
 sg13g2_decap_8 FILLER_60_77 ();
 sg13g2_fill_2 FILLER_60_84 ();
 sg13g2_fill_1 FILLER_60_86 ();
 sg13g2_fill_1 FILLER_60_92 ();
 sg13g2_fill_2 FILLER_60_98 ();
 sg13g2_fill_1 FILLER_60_100 ();
 sg13g2_fill_1 FILLER_60_105 ();
 sg13g2_fill_2 FILLER_60_111 ();
 sg13g2_decap_8 FILLER_60_117 ();
 sg13g2_decap_8 FILLER_60_124 ();
 sg13g2_decap_8 FILLER_60_131 ();
 sg13g2_fill_2 FILLER_60_138 ();
 sg13g2_fill_2 FILLER_60_144 ();
 sg13g2_fill_1 FILLER_60_146 ();
 sg13g2_decap_8 FILLER_60_156 ();
 sg13g2_decap_8 FILLER_60_163 ();
 sg13g2_decap_8 FILLER_60_170 ();
 sg13g2_decap_8 FILLER_60_177 ();
 sg13g2_decap_4 FILLER_60_184 ();
 sg13g2_fill_2 FILLER_60_200 ();
 sg13g2_decap_4 FILLER_60_207 ();
 sg13g2_decap_8 FILLER_60_214 ();
 sg13g2_decap_8 FILLER_60_221 ();
 sg13g2_fill_2 FILLER_60_228 ();
 sg13g2_decap_8 FILLER_60_234 ();
 sg13g2_decap_4 FILLER_60_269 ();
 sg13g2_fill_2 FILLER_60_273 ();
 sg13g2_decap_4 FILLER_60_279 ();
 sg13g2_decap_8 FILLER_60_287 ();
 sg13g2_decap_8 FILLER_60_294 ();
 sg13g2_decap_8 FILLER_60_301 ();
 sg13g2_fill_1 FILLER_60_308 ();
 sg13g2_fill_2 FILLER_60_326 ();
 sg13g2_fill_2 FILLER_60_337 ();
 sg13g2_fill_2 FILLER_60_346 ();
 sg13g2_fill_1 FILLER_60_348 ();
 sg13g2_fill_2 FILLER_60_353 ();
 sg13g2_fill_1 FILLER_60_355 ();
 sg13g2_fill_2 FILLER_60_361 ();
 sg13g2_fill_1 FILLER_60_363 ();
 sg13g2_decap_4 FILLER_60_390 ();
 sg13g2_decap_8 FILLER_60_399 ();
 sg13g2_decap_8 FILLER_60_406 ();
 sg13g2_decap_8 FILLER_60_413 ();
 sg13g2_decap_8 FILLER_60_420 ();
 sg13g2_fill_2 FILLER_60_427 ();
 sg13g2_fill_1 FILLER_60_429 ();
 sg13g2_decap_8 FILLER_61_0 ();
 sg13g2_decap_8 FILLER_61_7 ();
 sg13g2_decap_8 FILLER_61_14 ();
 sg13g2_decap_8 FILLER_61_21 ();
 sg13g2_decap_8 FILLER_61_28 ();
 sg13g2_decap_8 FILLER_61_35 ();
 sg13g2_decap_8 FILLER_61_42 ();
 sg13g2_decap_8 FILLER_61_49 ();
 sg13g2_decap_8 FILLER_61_56 ();
 sg13g2_decap_8 FILLER_61_63 ();
 sg13g2_decap_8 FILLER_61_70 ();
 sg13g2_decap_4 FILLER_61_77 ();
 sg13g2_fill_2 FILLER_61_85 ();
 sg13g2_fill_1 FILLER_61_87 ();
 sg13g2_decap_8 FILLER_61_115 ();
 sg13g2_decap_8 FILLER_61_122 ();
 sg13g2_decap_8 FILLER_61_129 ();
 sg13g2_fill_1 FILLER_61_136 ();
 sg13g2_decap_8 FILLER_61_154 ();
 sg13g2_decap_8 FILLER_61_161 ();
 sg13g2_decap_8 FILLER_61_168 ();
 sg13g2_decap_8 FILLER_61_223 ();
 sg13g2_decap_8 FILLER_61_230 ();
 sg13g2_decap_8 FILLER_61_237 ();
 sg13g2_fill_1 FILLER_61_244 ();
 sg13g2_decap_8 FILLER_61_275 ();
 sg13g2_decap_8 FILLER_61_282 ();
 sg13g2_decap_8 FILLER_61_289 ();
 sg13g2_decap_8 FILLER_61_296 ();
 sg13g2_decap_8 FILLER_61_303 ();
 sg13g2_fill_2 FILLER_61_310 ();
 sg13g2_fill_1 FILLER_61_312 ();
 sg13g2_decap_4 FILLER_61_322 ();
 sg13g2_fill_2 FILLER_61_340 ();
 sg13g2_fill_1 FILLER_61_373 ();
 sg13g2_fill_2 FILLER_61_378 ();
 sg13g2_fill_1 FILLER_61_380 ();
 sg13g2_decap_8 FILLER_61_412 ();
 sg13g2_decap_8 FILLER_61_419 ();
 sg13g2_decap_4 FILLER_61_426 ();
 sg13g2_decap_8 FILLER_62_0 ();
 sg13g2_decap_8 FILLER_62_7 ();
 sg13g2_decap_8 FILLER_62_14 ();
 sg13g2_decap_8 FILLER_62_21 ();
 sg13g2_decap_8 FILLER_62_28 ();
 sg13g2_decap_8 FILLER_62_35 ();
 sg13g2_decap_8 FILLER_62_42 ();
 sg13g2_decap_8 FILLER_62_49 ();
 sg13g2_decap_8 FILLER_62_56 ();
 sg13g2_decap_8 FILLER_62_63 ();
 sg13g2_decap_8 FILLER_62_70 ();
 sg13g2_decap_8 FILLER_62_77 ();
 sg13g2_decap_4 FILLER_62_84 ();
 sg13g2_fill_1 FILLER_62_88 ();
 sg13g2_decap_4 FILLER_62_93 ();
 sg13g2_fill_1 FILLER_62_106 ();
 sg13g2_fill_2 FILLER_62_115 ();
 sg13g2_fill_1 FILLER_62_117 ();
 sg13g2_decap_8 FILLER_62_154 ();
 sg13g2_fill_2 FILLER_62_161 ();
 sg13g2_fill_2 FILLER_62_166 ();
 sg13g2_fill_1 FILLER_62_168 ();
 sg13g2_fill_1 FILLER_62_179 ();
 sg13g2_decap_4 FILLER_62_194 ();
 sg13g2_fill_2 FILLER_62_208 ();
 sg13g2_fill_1 FILLER_62_218 ();
 sg13g2_decap_8 FILLER_62_231 ();
 sg13g2_decap_4 FILLER_62_238 ();
 sg13g2_decap_4 FILLER_62_247 ();
 sg13g2_fill_2 FILLER_62_251 ();
 sg13g2_decap_8 FILLER_62_288 ();
 sg13g2_decap_8 FILLER_62_295 ();
 sg13g2_decap_4 FILLER_62_302 ();
 sg13g2_fill_2 FILLER_62_306 ();
 sg13g2_decap_8 FILLER_62_312 ();
 sg13g2_decap_8 FILLER_62_319 ();
 sg13g2_decap_8 FILLER_62_326 ();
 sg13g2_decap_8 FILLER_62_333 ();
 sg13g2_fill_1 FILLER_62_340 ();
 sg13g2_decap_8 FILLER_62_345 ();
 sg13g2_decap_8 FILLER_62_352 ();
 sg13g2_decap_8 FILLER_62_359 ();
 sg13g2_decap_4 FILLER_62_366 ();
 sg13g2_fill_1 FILLER_62_370 ();
 sg13g2_decap_8 FILLER_62_375 ();
 sg13g2_decap_4 FILLER_62_382 ();
 sg13g2_fill_1 FILLER_62_386 ();
 sg13g2_fill_2 FILLER_62_392 ();
 sg13g2_decap_8 FILLER_62_408 ();
 sg13g2_decap_8 FILLER_62_415 ();
 sg13g2_decap_8 FILLER_62_422 ();
 sg13g2_fill_1 FILLER_62_429 ();
 sg13g2_decap_8 FILLER_63_0 ();
 sg13g2_decap_8 FILLER_63_7 ();
 sg13g2_decap_8 FILLER_63_14 ();
 sg13g2_decap_8 FILLER_63_21 ();
 sg13g2_decap_8 FILLER_63_28 ();
 sg13g2_decap_8 FILLER_63_35 ();
 sg13g2_decap_8 FILLER_63_42 ();
 sg13g2_decap_8 FILLER_63_49 ();
 sg13g2_decap_8 FILLER_63_56 ();
 sg13g2_decap_8 FILLER_63_63 ();
 sg13g2_decap_8 FILLER_63_70 ();
 sg13g2_decap_8 FILLER_63_77 ();
 sg13g2_fill_2 FILLER_63_108 ();
 sg13g2_fill_1 FILLER_63_110 ();
 sg13g2_decap_4 FILLER_63_141 ();
 sg13g2_fill_1 FILLER_63_145 ();
 sg13g2_decap_8 FILLER_63_179 ();
 sg13g2_fill_2 FILLER_63_186 ();
 sg13g2_fill_2 FILLER_63_206 ();
 sg13g2_fill_1 FILLER_63_258 ();
 sg13g2_decap_4 FILLER_63_263 ();
 sg13g2_fill_2 FILLER_63_267 ();
 sg13g2_decap_8 FILLER_63_273 ();
 sg13g2_decap_8 FILLER_63_284 ();
 sg13g2_decap_8 FILLER_63_291 ();
 sg13g2_decap_8 FILLER_63_298 ();
 sg13g2_fill_1 FILLER_63_305 ();
 sg13g2_decap_8 FILLER_63_336 ();
 sg13g2_decap_8 FILLER_63_343 ();
 sg13g2_decap_8 FILLER_63_350 ();
 sg13g2_decap_8 FILLER_63_357 ();
 sg13g2_decap_8 FILLER_63_364 ();
 sg13g2_decap_8 FILLER_63_371 ();
 sg13g2_decap_4 FILLER_63_378 ();
 sg13g2_fill_2 FILLER_63_382 ();
 sg13g2_fill_2 FILLER_63_391 ();
 sg13g2_decap_8 FILLER_63_419 ();
 sg13g2_decap_4 FILLER_63_426 ();
 sg13g2_decap_8 FILLER_64_0 ();
 sg13g2_decap_8 FILLER_64_7 ();
 sg13g2_decap_8 FILLER_64_14 ();
 sg13g2_decap_8 FILLER_64_21 ();
 sg13g2_decap_8 FILLER_64_28 ();
 sg13g2_decap_8 FILLER_64_35 ();
 sg13g2_decap_8 FILLER_64_42 ();
 sg13g2_decap_8 FILLER_64_49 ();
 sg13g2_decap_8 FILLER_64_56 ();
 sg13g2_decap_8 FILLER_64_63 ();
 sg13g2_decap_8 FILLER_64_70 ();
 sg13g2_decap_8 FILLER_64_77 ();
 sg13g2_fill_1 FILLER_64_84 ();
 sg13g2_fill_1 FILLER_64_98 ();
 sg13g2_fill_2 FILLER_64_112 ();
 sg13g2_decap_4 FILLER_64_128 ();
 sg13g2_decap_4 FILLER_64_148 ();
 sg13g2_fill_1 FILLER_64_152 ();
 sg13g2_decap_4 FILLER_64_163 ();
 sg13g2_fill_2 FILLER_64_172 ();
 sg13g2_decap_8 FILLER_64_184 ();
 sg13g2_fill_1 FILLER_64_191 ();
 sg13g2_fill_1 FILLER_64_208 ();
 sg13g2_fill_1 FILLER_64_234 ();
 sg13g2_fill_1 FILLER_64_248 ();
 sg13g2_decap_8 FILLER_64_258 ();
 sg13g2_decap_8 FILLER_64_269 ();
 sg13g2_fill_2 FILLER_64_306 ();
 sg13g2_fill_1 FILLER_64_308 ();
 sg13g2_decap_4 FILLER_64_317 ();
 sg13g2_fill_2 FILLER_64_347 ();
 sg13g2_fill_1 FILLER_64_375 ();
 sg13g2_fill_2 FILLER_64_402 ();
 sg13g2_decap_8 FILLER_64_408 ();
 sg13g2_decap_8 FILLER_64_415 ();
 sg13g2_decap_8 FILLER_64_422 ();
 sg13g2_fill_1 FILLER_64_429 ();
 sg13g2_decap_8 FILLER_65_0 ();
 sg13g2_decap_8 FILLER_65_7 ();
 sg13g2_decap_8 FILLER_65_14 ();
 sg13g2_decap_8 FILLER_65_21 ();
 sg13g2_decap_8 FILLER_65_28 ();
 sg13g2_decap_8 FILLER_65_35 ();
 sg13g2_decap_8 FILLER_65_42 ();
 sg13g2_decap_8 FILLER_65_49 ();
 sg13g2_decap_8 FILLER_65_56 ();
 sg13g2_decap_8 FILLER_65_63 ();
 sg13g2_decap_8 FILLER_65_70 ();
 sg13g2_decap_4 FILLER_65_77 ();
 sg13g2_decap_4 FILLER_65_86 ();
 sg13g2_decap_8 FILLER_65_105 ();
 sg13g2_decap_8 FILLER_65_112 ();
 sg13g2_fill_2 FILLER_65_119 ();
 sg13g2_fill_1 FILLER_65_121 ();
 sg13g2_decap_8 FILLER_65_148 ();
 sg13g2_decap_4 FILLER_65_155 ();
 sg13g2_fill_2 FILLER_65_174 ();
 sg13g2_fill_1 FILLER_65_180 ();
 sg13g2_fill_1 FILLER_65_186 ();
 sg13g2_decap_4 FILLER_65_192 ();
 sg13g2_fill_1 FILLER_65_196 ();
 sg13g2_decap_8 FILLER_65_211 ();
 sg13g2_decap_8 FILLER_65_223 ();
 sg13g2_fill_2 FILLER_65_230 ();
 sg13g2_fill_1 FILLER_65_232 ();
 sg13g2_decap_8 FILLER_65_237 ();
 sg13g2_fill_1 FILLER_65_244 ();
 sg13g2_decap_8 FILLER_65_271 ();
 sg13g2_decap_4 FILLER_65_278 ();
 sg13g2_fill_1 FILLER_65_282 ();
 sg13g2_decap_8 FILLER_65_287 ();
 sg13g2_fill_1 FILLER_65_294 ();
 sg13g2_fill_2 FILLER_65_303 ();
 sg13g2_fill_1 FILLER_65_305 ();
 sg13g2_fill_2 FILLER_65_310 ();
 sg13g2_fill_2 FILLER_65_333 ();
 sg13g2_decap_8 FILLER_65_340 ();
 sg13g2_decap_4 FILLER_65_347 ();
 sg13g2_decap_4 FILLER_65_377 ();
 sg13g2_fill_2 FILLER_65_381 ();
 sg13g2_decap_8 FILLER_65_387 ();
 sg13g2_decap_8 FILLER_65_394 ();
 sg13g2_decap_8 FILLER_65_401 ();
 sg13g2_decap_8 FILLER_65_408 ();
 sg13g2_decap_8 FILLER_65_415 ();
 sg13g2_decap_8 FILLER_65_422 ();
 sg13g2_fill_1 FILLER_65_429 ();
 sg13g2_decap_8 FILLER_66_0 ();
 sg13g2_decap_8 FILLER_66_7 ();
 sg13g2_decap_8 FILLER_66_14 ();
 sg13g2_decap_8 FILLER_66_21 ();
 sg13g2_decap_8 FILLER_66_28 ();
 sg13g2_decap_8 FILLER_66_35 ();
 sg13g2_decap_8 FILLER_66_42 ();
 sg13g2_decap_8 FILLER_66_49 ();
 sg13g2_decap_8 FILLER_66_56 ();
 sg13g2_decap_8 FILLER_66_63 ();
 sg13g2_decap_8 FILLER_66_70 ();
 sg13g2_decap_8 FILLER_66_77 ();
 sg13g2_fill_1 FILLER_66_84 ();
 sg13g2_fill_1 FILLER_66_101 ();
 sg13g2_decap_8 FILLER_66_106 ();
 sg13g2_decap_8 FILLER_66_113 ();
 sg13g2_decap_4 FILLER_66_120 ();
 sg13g2_fill_2 FILLER_66_124 ();
 sg13g2_decap_8 FILLER_66_145 ();
 sg13g2_fill_1 FILLER_66_152 ();
 sg13g2_fill_1 FILLER_66_162 ();
 sg13g2_decap_8 FILLER_66_187 ();
 sg13g2_decap_4 FILLER_66_194 ();
 sg13g2_fill_1 FILLER_66_198 ();
 sg13g2_fill_1 FILLER_66_203 ();
 sg13g2_fill_1 FILLER_66_214 ();
 sg13g2_decap_8 FILLER_66_219 ();
 sg13g2_decap_4 FILLER_66_226 ();
 sg13g2_fill_2 FILLER_66_230 ();
 sg13g2_decap_4 FILLER_66_319 ();
 sg13g2_fill_1 FILLER_66_323 ();
 sg13g2_fill_2 FILLER_66_346 ();
 sg13g2_decap_4 FILLER_66_352 ();
 sg13g2_fill_1 FILLER_66_356 ();
 sg13g2_decap_4 FILLER_66_364 ();
 sg13g2_decap_8 FILLER_66_405 ();
 sg13g2_decap_8 FILLER_66_412 ();
 sg13g2_decap_8 FILLER_66_419 ();
 sg13g2_decap_4 FILLER_66_426 ();
 sg13g2_decap_8 FILLER_67_0 ();
 sg13g2_decap_8 FILLER_67_7 ();
 sg13g2_decap_8 FILLER_67_14 ();
 sg13g2_decap_8 FILLER_67_21 ();
 sg13g2_decap_8 FILLER_67_28 ();
 sg13g2_decap_8 FILLER_67_35 ();
 sg13g2_decap_8 FILLER_67_42 ();
 sg13g2_decap_8 FILLER_67_49 ();
 sg13g2_decap_8 FILLER_67_56 ();
 sg13g2_decap_8 FILLER_67_63 ();
 sg13g2_decap_8 FILLER_67_70 ();
 sg13g2_decap_4 FILLER_67_77 ();
 sg13g2_fill_2 FILLER_67_81 ();
 sg13g2_fill_2 FILLER_67_90 ();
 sg13g2_fill_1 FILLER_67_132 ();
 sg13g2_fill_1 FILLER_67_146 ();
 sg13g2_fill_1 FILLER_67_164 ();
 sg13g2_fill_1 FILLER_67_175 ();
 sg13g2_fill_2 FILLER_67_195 ();
 sg13g2_decap_4 FILLER_67_201 ();
 sg13g2_fill_1 FILLER_67_205 ();
 sg13g2_fill_2 FILLER_67_209 ();
 sg13g2_fill_1 FILLER_67_223 ();
 sg13g2_fill_1 FILLER_67_229 ();
 sg13g2_decap_4 FILLER_67_239 ();
 sg13g2_decap_8 FILLER_67_255 ();
 sg13g2_decap_8 FILLER_67_262 ();
 sg13g2_decap_8 FILLER_67_269 ();
 sg13g2_decap_4 FILLER_67_276 ();
 sg13g2_fill_1 FILLER_67_280 ();
 sg13g2_fill_2 FILLER_67_301 ();
 sg13g2_fill_1 FILLER_67_333 ();
 sg13g2_decap_4 FILLER_67_338 ();
 sg13g2_decap_4 FILLER_67_378 ();
 sg13g2_decap_4 FILLER_67_386 ();
 sg13g2_fill_1 FILLER_67_390 ();
 sg13g2_decap_8 FILLER_67_417 ();
 sg13g2_decap_4 FILLER_67_424 ();
 sg13g2_fill_2 FILLER_67_428 ();
 sg13g2_decap_8 FILLER_68_0 ();
 sg13g2_decap_8 FILLER_68_7 ();
 sg13g2_decap_8 FILLER_68_14 ();
 sg13g2_decap_8 FILLER_68_21 ();
 sg13g2_decap_8 FILLER_68_28 ();
 sg13g2_decap_8 FILLER_68_35 ();
 sg13g2_decap_8 FILLER_68_42 ();
 sg13g2_decap_8 FILLER_68_49 ();
 sg13g2_decap_8 FILLER_68_56 ();
 sg13g2_decap_8 FILLER_68_63 ();
 sg13g2_decap_8 FILLER_68_70 ();
 sg13g2_decap_8 FILLER_68_77 ();
 sg13g2_fill_1 FILLER_68_89 ();
 sg13g2_fill_1 FILLER_68_98 ();
 sg13g2_fill_2 FILLER_68_139 ();
 sg13g2_fill_2 FILLER_68_145 ();
 sg13g2_fill_1 FILLER_68_147 ();
 sg13g2_fill_2 FILLER_68_157 ();
 sg13g2_fill_2 FILLER_68_193 ();
 sg13g2_fill_1 FILLER_68_205 ();
 sg13g2_fill_1 FILLER_68_220 ();
 sg13g2_decap_8 FILLER_68_231 ();
 sg13g2_decap_4 FILLER_68_238 ();
 sg13g2_decap_8 FILLER_68_251 ();
 sg13g2_decap_8 FILLER_68_258 ();
 sg13g2_decap_4 FILLER_68_265 ();
 sg13g2_decap_8 FILLER_68_273 ();
 sg13g2_decap_8 FILLER_68_280 ();
 sg13g2_decap_8 FILLER_68_287 ();
 sg13g2_fill_1 FILLER_68_298 ();
 sg13g2_fill_2 FILLER_68_307 ();
 sg13g2_fill_1 FILLER_68_309 ();
 sg13g2_fill_2 FILLER_68_316 ();
 sg13g2_decap_8 FILLER_68_322 ();
 sg13g2_decap_8 FILLER_68_329 ();
 sg13g2_fill_2 FILLER_68_336 ();
 sg13g2_decap_4 FILLER_68_397 ();
 sg13g2_fill_2 FILLER_68_401 ();
 sg13g2_fill_1 FILLER_68_429 ();
 sg13g2_decap_8 FILLER_69_0 ();
 sg13g2_decap_8 FILLER_69_7 ();
 sg13g2_decap_8 FILLER_69_14 ();
 sg13g2_decap_8 FILLER_69_21 ();
 sg13g2_decap_8 FILLER_69_28 ();
 sg13g2_decap_8 FILLER_69_35 ();
 sg13g2_decap_8 FILLER_69_42 ();
 sg13g2_decap_8 FILLER_69_49 ();
 sg13g2_decap_8 FILLER_69_56 ();
 sg13g2_decap_8 FILLER_69_63 ();
 sg13g2_decap_8 FILLER_69_70 ();
 sg13g2_decap_8 FILLER_69_77 ();
 sg13g2_fill_2 FILLER_69_84 ();
 sg13g2_fill_1 FILLER_69_86 ();
 sg13g2_decap_4 FILLER_69_107 ();
 sg13g2_fill_2 FILLER_69_111 ();
 sg13g2_decap_8 FILLER_69_143 ();
 sg13g2_decap_4 FILLER_69_150 ();
 sg13g2_fill_1 FILLER_69_154 ();
 sg13g2_fill_2 FILLER_69_159 ();
 sg13g2_fill_1 FILLER_69_166 ();
 sg13g2_fill_1 FILLER_69_172 ();
 sg13g2_fill_1 FILLER_69_181 ();
 sg13g2_fill_1 FILLER_69_185 ();
 sg13g2_fill_2 FILLER_69_212 ();
 sg13g2_fill_1 FILLER_69_214 ();
 sg13g2_fill_2 FILLER_69_223 ();
 sg13g2_decap_8 FILLER_69_235 ();
 sg13g2_decap_8 FILLER_69_242 ();
 sg13g2_decap_4 FILLER_69_249 ();
 sg13g2_fill_1 FILLER_69_253 ();
 sg13g2_decap_8 FILLER_69_293 ();
 sg13g2_decap_4 FILLER_69_300 ();
 sg13g2_fill_1 FILLER_69_304 ();
 sg13g2_decap_8 FILLER_69_320 ();
 sg13g2_decap_8 FILLER_69_327 ();
 sg13g2_decap_4 FILLER_69_334 ();
 sg13g2_fill_1 FILLER_69_342 ();
 sg13g2_decap_8 FILLER_69_347 ();
 sg13g2_fill_2 FILLER_69_354 ();
 sg13g2_decap_8 FILLER_69_360 ();
 sg13g2_decap_4 FILLER_69_367 ();
 sg13g2_decap_4 FILLER_69_375 ();
 sg13g2_decap_8 FILLER_69_419 ();
 sg13g2_decap_4 FILLER_69_426 ();
 sg13g2_decap_8 FILLER_70_0 ();
 sg13g2_decap_8 FILLER_70_7 ();
 sg13g2_decap_8 FILLER_70_14 ();
 sg13g2_decap_8 FILLER_70_21 ();
 sg13g2_decap_8 FILLER_70_28 ();
 sg13g2_decap_8 FILLER_70_35 ();
 sg13g2_decap_8 FILLER_70_42 ();
 sg13g2_decap_8 FILLER_70_49 ();
 sg13g2_decap_8 FILLER_70_56 ();
 sg13g2_decap_8 FILLER_70_63 ();
 sg13g2_decap_8 FILLER_70_70 ();
 sg13g2_decap_8 FILLER_70_77 ();
 sg13g2_decap_8 FILLER_70_84 ();
 sg13g2_decap_8 FILLER_70_91 ();
 sg13g2_decap_8 FILLER_70_98 ();
 sg13g2_decap_8 FILLER_70_105 ();
 sg13g2_decap_8 FILLER_70_112 ();
 sg13g2_fill_2 FILLER_70_119 ();
 sg13g2_fill_1 FILLER_70_121 ();
 sg13g2_decap_8 FILLER_70_130 ();
 sg13g2_decap_8 FILLER_70_137 ();
 sg13g2_decap_8 FILLER_70_144 ();
 sg13g2_decap_4 FILLER_70_155 ();
 sg13g2_fill_1 FILLER_70_159 ();
 sg13g2_decap_8 FILLER_70_168 ();
 sg13g2_decap_4 FILLER_70_175 ();
 sg13g2_fill_1 FILLER_70_179 ();
 sg13g2_decap_4 FILLER_70_189 ();
 sg13g2_fill_2 FILLER_70_193 ();
 sg13g2_decap_8 FILLER_70_199 ();
 sg13g2_decap_8 FILLER_70_206 ();
 sg13g2_decap_8 FILLER_70_213 ();
 sg13g2_decap_4 FILLER_70_225 ();
 sg13g2_decap_8 FILLER_70_233 ();
 sg13g2_decap_8 FILLER_70_240 ();
 sg13g2_decap_4 FILLER_70_247 ();
 sg13g2_decap_8 FILLER_70_255 ();
 sg13g2_decap_8 FILLER_70_262 ();
 sg13g2_decap_4 FILLER_70_269 ();
 sg13g2_fill_1 FILLER_70_273 ();
 sg13g2_fill_2 FILLER_70_282 ();
 sg13g2_decap_4 FILLER_70_292 ();
 sg13g2_fill_1 FILLER_70_311 ();
 sg13g2_decap_4 FILLER_70_317 ();
 sg13g2_fill_2 FILLER_70_321 ();
 sg13g2_decap_8 FILLER_70_329 ();
 sg13g2_fill_2 FILLER_70_349 ();
 sg13g2_decap_4 FILLER_70_355 ();
 sg13g2_decap_8 FILLER_70_364 ();
 sg13g2_decap_8 FILLER_70_371 ();
 sg13g2_decap_8 FILLER_70_378 ();
 sg13g2_fill_2 FILLER_70_385 ();
 sg13g2_decap_8 FILLER_70_408 ();
 sg13g2_decap_8 FILLER_70_415 ();
 sg13g2_decap_8 FILLER_70_422 ();
 sg13g2_fill_1 FILLER_70_429 ();
 sg13g2_decap_8 FILLER_71_0 ();
 sg13g2_decap_8 FILLER_71_7 ();
 sg13g2_decap_8 FILLER_71_14 ();
 sg13g2_decap_8 FILLER_71_21 ();
 sg13g2_decap_8 FILLER_71_28 ();
 sg13g2_decap_8 FILLER_71_35 ();
 sg13g2_decap_8 FILLER_71_42 ();
 sg13g2_decap_8 FILLER_71_49 ();
 sg13g2_decap_8 FILLER_71_56 ();
 sg13g2_decap_8 FILLER_71_63 ();
 sg13g2_decap_8 FILLER_71_70 ();
 sg13g2_decap_8 FILLER_71_77 ();
 sg13g2_decap_8 FILLER_71_84 ();
 sg13g2_decap_8 FILLER_71_91 ();
 sg13g2_decap_8 FILLER_71_98 ();
 sg13g2_decap_8 FILLER_71_105 ();
 sg13g2_decap_4 FILLER_71_112 ();
 sg13g2_fill_1 FILLER_71_116 ();
 sg13g2_decap_8 FILLER_71_121 ();
 sg13g2_decap_8 FILLER_71_128 ();
 sg13g2_decap_8 FILLER_71_135 ();
 sg13g2_fill_2 FILLER_71_142 ();
 sg13g2_fill_1 FILLER_71_144 ();
 sg13g2_fill_2 FILLER_71_176 ();
 sg13g2_decap_8 FILLER_71_186 ();
 sg13g2_decap_8 FILLER_71_193 ();
 sg13g2_decap_8 FILLER_71_200 ();
 sg13g2_fill_1 FILLER_71_207 ();
 sg13g2_fill_2 FILLER_71_215 ();
 sg13g2_fill_1 FILLER_71_222 ();
 sg13g2_fill_2 FILLER_71_227 ();
 sg13g2_decap_8 FILLER_71_234 ();
 sg13g2_fill_2 FILLER_71_241 ();
 sg13g2_fill_1 FILLER_71_243 ();
 sg13g2_decap_4 FILLER_71_283 ();
 sg13g2_fill_2 FILLER_71_287 ();
 sg13g2_decap_8 FILLER_71_301 ();
 sg13g2_fill_2 FILLER_71_308 ();
 sg13g2_fill_1 FILLER_71_318 ();
 sg13g2_fill_2 FILLER_71_325 ();
 sg13g2_fill_1 FILLER_71_370 ();
 sg13g2_decap_8 FILLER_71_375 ();
 sg13g2_decap_8 FILLER_71_382 ();
 sg13g2_decap_8 FILLER_71_389 ();
 sg13g2_decap_8 FILLER_71_396 ();
 sg13g2_decap_8 FILLER_71_403 ();
 sg13g2_decap_8 FILLER_71_410 ();
 sg13g2_decap_8 FILLER_71_417 ();
 sg13g2_decap_4 FILLER_71_424 ();
 sg13g2_fill_2 FILLER_71_428 ();
 sg13g2_decap_8 FILLER_72_0 ();
 sg13g2_decap_8 FILLER_72_7 ();
 sg13g2_decap_8 FILLER_72_14 ();
 sg13g2_decap_8 FILLER_72_21 ();
 sg13g2_decap_8 FILLER_72_28 ();
 sg13g2_decap_8 FILLER_72_35 ();
 sg13g2_decap_8 FILLER_72_42 ();
 sg13g2_decap_8 FILLER_72_49 ();
 sg13g2_decap_8 FILLER_72_56 ();
 sg13g2_decap_8 FILLER_72_63 ();
 sg13g2_decap_8 FILLER_72_70 ();
 sg13g2_decap_8 FILLER_72_77 ();
 sg13g2_decap_8 FILLER_72_84 ();
 sg13g2_decap_8 FILLER_72_121 ();
 sg13g2_decap_8 FILLER_72_128 ();
 sg13g2_decap_8 FILLER_72_135 ();
 sg13g2_decap_8 FILLER_72_142 ();
 sg13g2_fill_2 FILLER_72_149 ();
 sg13g2_fill_1 FILLER_72_151 ();
 sg13g2_fill_1 FILLER_72_169 ();
 sg13g2_fill_1 FILLER_72_187 ();
 sg13g2_decap_8 FILLER_72_196 ();
 sg13g2_fill_1 FILLER_72_203 ();
 sg13g2_decap_8 FILLER_72_245 ();
 sg13g2_decap_8 FILLER_72_256 ();
 sg13g2_decap_8 FILLER_72_263 ();
 sg13g2_decap_4 FILLER_72_270 ();
 sg13g2_fill_2 FILLER_72_282 ();
 sg13g2_fill_1 FILLER_72_284 ();
 sg13g2_fill_1 FILLER_72_298 ();
 sg13g2_decap_4 FILLER_72_328 ();
 sg13g2_fill_2 FILLER_72_338 ();
 sg13g2_fill_1 FILLER_72_348 ();
 sg13g2_fill_2 FILLER_72_357 ();
 sg13g2_fill_2 FILLER_72_389 ();
 sg13g2_fill_1 FILLER_72_391 ();
 sg13g2_decap_4 FILLER_72_408 ();
 sg13g2_decap_8 FILLER_72_416 ();
 sg13g2_decap_8 FILLER_72_423 ();
 sg13g2_decap_8 FILLER_73_0 ();
 sg13g2_decap_8 FILLER_73_7 ();
 sg13g2_decap_8 FILLER_73_14 ();
 sg13g2_decap_8 FILLER_73_21 ();
 sg13g2_decap_8 FILLER_73_28 ();
 sg13g2_decap_8 FILLER_73_35 ();
 sg13g2_decap_8 FILLER_73_42 ();
 sg13g2_decap_8 FILLER_73_49 ();
 sg13g2_decap_8 FILLER_73_56 ();
 sg13g2_decap_8 FILLER_73_63 ();
 sg13g2_decap_8 FILLER_73_70 ();
 sg13g2_decap_8 FILLER_73_77 ();
 sg13g2_decap_8 FILLER_73_84 ();
 sg13g2_fill_1 FILLER_73_91 ();
 sg13g2_fill_1 FILLER_73_127 ();
 sg13g2_decap_8 FILLER_73_141 ();
 sg13g2_fill_2 FILLER_73_148 ();
 sg13g2_decap_4 FILLER_73_156 ();
 sg13g2_decap_4 FILLER_73_165 ();
 sg13g2_decap_4 FILLER_73_239 ();
 sg13g2_fill_2 FILLER_73_285 ();
 sg13g2_fill_1 FILLER_73_296 ();
 sg13g2_fill_2 FILLER_73_318 ();
 sg13g2_fill_1 FILLER_73_334 ();
 sg13g2_fill_2 FILLER_73_373 ();
 sg13g2_fill_1 FILLER_73_375 ();
 sg13g2_fill_2 FILLER_73_428 ();
 sg13g2_decap_8 FILLER_74_0 ();
 sg13g2_decap_8 FILLER_74_7 ();
 sg13g2_decap_8 FILLER_74_14 ();
 sg13g2_decap_8 FILLER_74_21 ();
 sg13g2_decap_8 FILLER_74_28 ();
 sg13g2_decap_8 FILLER_74_35 ();
 sg13g2_decap_8 FILLER_74_42 ();
 sg13g2_decap_8 FILLER_74_49 ();
 sg13g2_decap_8 FILLER_74_56 ();
 sg13g2_decap_8 FILLER_74_63 ();
 sg13g2_decap_8 FILLER_74_70 ();
 sg13g2_fill_2 FILLER_74_77 ();
 sg13g2_fill_1 FILLER_74_79 ();
 sg13g2_fill_2 FILLER_74_138 ();
 sg13g2_decap_8 FILLER_74_149 ();
 sg13g2_decap_8 FILLER_74_156 ();
 sg13g2_decap_8 FILLER_74_163 ();
 sg13g2_decap_8 FILLER_74_170 ();
 sg13g2_decap_4 FILLER_74_177 ();
 sg13g2_fill_2 FILLER_74_181 ();
 sg13g2_decap_4 FILLER_74_250 ();
 sg13g2_fill_2 FILLER_74_254 ();
 sg13g2_decap_8 FILLER_74_270 ();
 sg13g2_decap_8 FILLER_74_277 ();
 sg13g2_decap_4 FILLER_74_284 ();
 sg13g2_fill_2 FILLER_74_288 ();
 sg13g2_decap_4 FILLER_74_327 ();
 sg13g2_fill_2 FILLER_74_331 ();
 sg13g2_decap_4 FILLER_74_337 ();
 sg13g2_fill_2 FILLER_74_345 ();
 sg13g2_fill_1 FILLER_74_347 ();
 sg13g2_decap_4 FILLER_74_353 ();
 sg13g2_fill_1 FILLER_74_357 ();
 sg13g2_decap_4 FILLER_74_362 ();
 sg13g2_fill_1 FILLER_74_366 ();
 sg13g2_decap_8 FILLER_74_371 ();
 sg13g2_fill_2 FILLER_74_382 ();
 sg13g2_decap_4 FILLER_74_400 ();
 sg13g2_fill_2 FILLER_74_409 ();
 sg13g2_decap_8 FILLER_74_415 ();
 sg13g2_decap_8 FILLER_74_422 ();
 sg13g2_fill_1 FILLER_74_429 ();
 sg13g2_decap_8 FILLER_75_0 ();
 sg13g2_decap_8 FILLER_75_7 ();
 sg13g2_decap_8 FILLER_75_14 ();
 sg13g2_decap_8 FILLER_75_21 ();
 sg13g2_decap_8 FILLER_75_28 ();
 sg13g2_decap_8 FILLER_75_35 ();
 sg13g2_decap_8 FILLER_75_42 ();
 sg13g2_decap_8 FILLER_75_49 ();
 sg13g2_decap_8 FILLER_75_56 ();
 sg13g2_decap_8 FILLER_75_63 ();
 sg13g2_decap_8 FILLER_75_70 ();
 sg13g2_decap_8 FILLER_75_77 ();
 sg13g2_decap_8 FILLER_75_88 ();
 sg13g2_decap_8 FILLER_75_95 ();
 sg13g2_decap_4 FILLER_75_102 ();
 sg13g2_fill_2 FILLER_75_106 ();
 sg13g2_fill_2 FILLER_75_138 ();
 sg13g2_decap_4 FILLER_75_186 ();
 sg13g2_fill_1 FILLER_75_190 ();
 sg13g2_decap_8 FILLER_75_195 ();
 sg13g2_decap_8 FILLER_75_207 ();
 sg13g2_decap_4 FILLER_75_219 ();
 sg13g2_fill_2 FILLER_75_232 ();
 sg13g2_decap_8 FILLER_75_265 ();
 sg13g2_decap_8 FILLER_75_272 ();
 sg13g2_decap_8 FILLER_75_279 ();
 sg13g2_decap_8 FILLER_75_286 ();
 sg13g2_fill_2 FILLER_75_293 ();
 sg13g2_fill_1 FILLER_75_295 ();
 sg13g2_decap_4 FILLER_75_300 ();
 sg13g2_fill_2 FILLER_75_309 ();
 sg13g2_fill_1 FILLER_75_311 ();
 sg13g2_decap_8 FILLER_75_317 ();
 sg13g2_decap_4 FILLER_75_324 ();
 sg13g2_fill_2 FILLER_75_328 ();
 sg13g2_decap_8 FILLER_75_335 ();
 sg13g2_fill_1 FILLER_75_342 ();
 sg13g2_decap_8 FILLER_75_381 ();
 sg13g2_fill_2 FILLER_75_388 ();
 sg13g2_decap_4 FILLER_75_395 ();
 sg13g2_decap_8 FILLER_75_405 ();
 sg13g2_decap_8 FILLER_75_412 ();
 sg13g2_decap_8 FILLER_75_419 ();
 sg13g2_decap_4 FILLER_75_426 ();
 sg13g2_decap_8 FILLER_76_0 ();
 sg13g2_decap_8 FILLER_76_7 ();
 sg13g2_decap_8 FILLER_76_14 ();
 sg13g2_decap_8 FILLER_76_21 ();
 sg13g2_decap_8 FILLER_76_28 ();
 sg13g2_decap_8 FILLER_76_35 ();
 sg13g2_decap_8 FILLER_76_42 ();
 sg13g2_decap_8 FILLER_76_49 ();
 sg13g2_decap_8 FILLER_76_56 ();
 sg13g2_decap_8 FILLER_76_63 ();
 sg13g2_decap_8 FILLER_76_70 ();
 sg13g2_decap_8 FILLER_76_77 ();
 sg13g2_decap_8 FILLER_76_84 ();
 sg13g2_decap_8 FILLER_76_91 ();
 sg13g2_decap_8 FILLER_76_98 ();
 sg13g2_decap_8 FILLER_76_105 ();
 sg13g2_decap_8 FILLER_76_112 ();
 sg13g2_decap_8 FILLER_76_123 ();
 sg13g2_decap_8 FILLER_76_130 ();
 sg13g2_decap_8 FILLER_76_137 ();
 sg13g2_fill_1 FILLER_76_170 ();
 sg13g2_decap_4 FILLER_76_176 ();
 sg13g2_decap_4 FILLER_76_232 ();
 sg13g2_fill_1 FILLER_76_236 ();
 sg13g2_decap_4 FILLER_76_243 ();
 sg13g2_decap_4 FILLER_76_251 ();
 sg13g2_fill_1 FILLER_76_255 ();
 sg13g2_fill_2 FILLER_76_261 ();
 sg13g2_fill_1 FILLER_76_263 ();
 sg13g2_decap_4 FILLER_76_276 ();
 sg13g2_decap_4 FILLER_76_295 ();
 sg13g2_fill_1 FILLER_76_299 ();
 sg13g2_decap_4 FILLER_76_304 ();
 sg13g2_fill_2 FILLER_76_308 ();
 sg13g2_decap_8 FILLER_76_336 ();
 sg13g2_decap_8 FILLER_76_343 ();
 sg13g2_decap_8 FILLER_76_354 ();
 sg13g2_decap_8 FILLER_76_361 ();
 sg13g2_fill_2 FILLER_76_368 ();
 sg13g2_decap_4 FILLER_76_377 ();
 sg13g2_fill_1 FILLER_76_393 ();
 sg13g2_fill_1 FILLER_76_397 ();
 sg13g2_fill_2 FILLER_76_402 ();
 sg13g2_decap_8 FILLER_77_0 ();
 sg13g2_decap_8 FILLER_77_7 ();
 sg13g2_decap_8 FILLER_77_14 ();
 sg13g2_decap_8 FILLER_77_21 ();
 sg13g2_decap_8 FILLER_77_28 ();
 sg13g2_decap_8 FILLER_77_35 ();
 sg13g2_decap_8 FILLER_77_42 ();
 sg13g2_decap_8 FILLER_77_49 ();
 sg13g2_decap_8 FILLER_77_56 ();
 sg13g2_decap_8 FILLER_77_63 ();
 sg13g2_decap_8 FILLER_77_70 ();
 sg13g2_decap_8 FILLER_77_77 ();
 sg13g2_decap_8 FILLER_77_84 ();
 sg13g2_decap_8 FILLER_77_91 ();
 sg13g2_decap_8 FILLER_77_98 ();
 sg13g2_decap_8 FILLER_77_105 ();
 sg13g2_decap_8 FILLER_77_112 ();
 sg13g2_decap_8 FILLER_77_119 ();
 sg13g2_decap_8 FILLER_77_126 ();
 sg13g2_decap_8 FILLER_77_133 ();
 sg13g2_decap_8 FILLER_77_140 ();
 sg13g2_decap_4 FILLER_77_147 ();
 sg13g2_fill_1 FILLER_77_151 ();
 sg13g2_fill_2 FILLER_77_156 ();
 sg13g2_fill_1 FILLER_77_158 ();
 sg13g2_fill_1 FILLER_77_188 ();
 sg13g2_decap_8 FILLER_77_193 ();
 sg13g2_decap_4 FILLER_77_200 ();
 sg13g2_fill_2 FILLER_77_204 ();
 sg13g2_decap_8 FILLER_77_209 ();
 sg13g2_decap_4 FILLER_77_216 ();
 sg13g2_fill_2 FILLER_77_220 ();
 sg13g2_fill_2 FILLER_77_231 ();
 sg13g2_fill_2 FILLER_77_270 ();
 sg13g2_fill_2 FILLER_77_298 ();
 sg13g2_decap_8 FILLER_77_331 ();
 sg13g2_decap_8 FILLER_77_338 ();
 sg13g2_fill_2 FILLER_77_345 ();
 sg13g2_fill_1 FILLER_77_351 ();
 sg13g2_decap_8 FILLER_77_378 ();
 sg13g2_decap_8 FILLER_77_385 ();
 sg13g2_decap_4 FILLER_77_392 ();
 sg13g2_decap_4 FILLER_77_408 ();
 sg13g2_decap_8 FILLER_77_416 ();
 sg13g2_decap_8 FILLER_77_423 ();
 sg13g2_decap_8 FILLER_78_0 ();
 sg13g2_decap_8 FILLER_78_7 ();
 sg13g2_decap_8 FILLER_78_14 ();
 sg13g2_decap_8 FILLER_78_21 ();
 sg13g2_decap_8 FILLER_78_28 ();
 sg13g2_decap_8 FILLER_78_35 ();
 sg13g2_decap_8 FILLER_78_42 ();
 sg13g2_decap_8 FILLER_78_49 ();
 sg13g2_decap_8 FILLER_78_56 ();
 sg13g2_decap_8 FILLER_78_63 ();
 sg13g2_decap_8 FILLER_78_70 ();
 sg13g2_decap_8 FILLER_78_77 ();
 sg13g2_decap_8 FILLER_78_84 ();
 sg13g2_decap_8 FILLER_78_91 ();
 sg13g2_decap_8 FILLER_78_98 ();
 sg13g2_decap_8 FILLER_78_105 ();
 sg13g2_decap_8 FILLER_78_112 ();
 sg13g2_decap_8 FILLER_78_119 ();
 sg13g2_decap_8 FILLER_78_126 ();
 sg13g2_decap_8 FILLER_78_133 ();
 sg13g2_decap_8 FILLER_78_140 ();
 sg13g2_decap_4 FILLER_78_147 ();
 sg13g2_fill_1 FILLER_78_151 ();
 sg13g2_fill_1 FILLER_78_188 ();
 sg13g2_fill_1 FILLER_78_196 ();
 sg13g2_fill_1 FILLER_78_204 ();
 sg13g2_fill_2 FILLER_78_210 ();
 sg13g2_fill_1 FILLER_78_212 ();
 sg13g2_decap_4 FILLER_78_248 ();
 sg13g2_decap_8 FILLER_78_256 ();
 sg13g2_decap_8 FILLER_78_263 ();
 sg13g2_fill_1 FILLER_78_270 ();
 sg13g2_fill_1 FILLER_78_292 ();
 sg13g2_decap_8 FILLER_78_297 ();
 sg13g2_fill_2 FILLER_78_304 ();
 sg13g2_fill_1 FILLER_78_306 ();
 sg13g2_fill_2 FILLER_78_311 ();
 sg13g2_fill_1 FILLER_78_317 ();
 sg13g2_fill_1 FILLER_78_331 ();
 sg13g2_fill_1 FILLER_78_341 ();
 sg13g2_fill_2 FILLER_78_428 ();
 sg13g2_decap_8 FILLER_79_0 ();
 sg13g2_decap_8 FILLER_79_7 ();
 sg13g2_decap_8 FILLER_79_14 ();
 sg13g2_decap_8 FILLER_79_21 ();
 sg13g2_decap_8 FILLER_79_28 ();
 sg13g2_decap_8 FILLER_79_35 ();
 sg13g2_decap_8 FILLER_79_42 ();
 sg13g2_decap_8 FILLER_79_49 ();
 sg13g2_decap_8 FILLER_79_56 ();
 sg13g2_decap_8 FILLER_79_63 ();
 sg13g2_decap_8 FILLER_79_70 ();
 sg13g2_decap_4 FILLER_79_77 ();
 sg13g2_decap_8 FILLER_79_85 ();
 sg13g2_decap_8 FILLER_79_92 ();
 sg13g2_decap_8 FILLER_79_99 ();
 sg13g2_decap_8 FILLER_79_106 ();
 sg13g2_decap_8 FILLER_79_113 ();
 sg13g2_decap_8 FILLER_79_120 ();
 sg13g2_decap_8 FILLER_79_127 ();
 sg13g2_decap_8 FILLER_79_134 ();
 sg13g2_decap_8 FILLER_79_141 ();
 sg13g2_decap_8 FILLER_79_148 ();
 sg13g2_decap_4 FILLER_79_155 ();
 sg13g2_fill_1 FILLER_79_159 ();
 sg13g2_decap_4 FILLER_79_163 ();
 sg13g2_fill_1 FILLER_79_167 ();
 sg13g2_fill_2 FILLER_79_172 ();
 sg13g2_fill_1 FILLER_79_181 ();
 sg13g2_fill_1 FILLER_79_208 ();
 sg13g2_fill_1 FILLER_79_216 ();
 sg13g2_fill_1 FILLER_79_221 ();
 sg13g2_fill_1 FILLER_79_229 ();
 sg13g2_fill_1 FILLER_79_235 ();
 sg13g2_fill_1 FILLER_79_243 ();
 sg13g2_fill_2 FILLER_79_249 ();
 sg13g2_decap_8 FILLER_79_255 ();
 sg13g2_fill_1 FILLER_79_262 ();
 sg13g2_fill_1 FILLER_79_289 ();
 sg13g2_fill_1 FILLER_79_342 ();
 sg13g2_fill_2 FILLER_79_359 ();
 sg13g2_decap_4 FILLER_79_374 ();
 sg13g2_fill_1 FILLER_79_378 ();
 sg13g2_fill_1 FILLER_79_383 ();
 sg13g2_decap_4 FILLER_79_388 ();
 sg13g2_decap_8 FILLER_79_404 ();
 sg13g2_decap_8 FILLER_79_415 ();
 sg13g2_decap_8 FILLER_79_422 ();
 sg13g2_fill_1 FILLER_79_429 ();
 sg13g2_decap_8 FILLER_80_0 ();
 sg13g2_decap_8 FILLER_80_7 ();
 sg13g2_decap_8 FILLER_80_14 ();
 sg13g2_decap_8 FILLER_80_21 ();
 sg13g2_decap_8 FILLER_80_28 ();
 sg13g2_decap_8 FILLER_80_35 ();
 sg13g2_decap_8 FILLER_80_42 ();
 sg13g2_decap_8 FILLER_80_49 ();
 sg13g2_decap_8 FILLER_80_56 ();
 sg13g2_decap_8 FILLER_80_63 ();
 sg13g2_decap_8 FILLER_80_70 ();
 sg13g2_fill_2 FILLER_80_77 ();
 sg13g2_fill_1 FILLER_80_79 ();
 sg13g2_fill_2 FILLER_80_144 ();
 sg13g2_decap_8 FILLER_80_154 ();
 sg13g2_decap_8 FILLER_80_161 ();
 sg13g2_fill_1 FILLER_80_212 ();
 sg13g2_fill_1 FILLER_80_221 ();
 sg13g2_fill_1 FILLER_80_226 ();
 sg13g2_fill_2 FILLER_80_258 ();
 sg13g2_decap_8 FILLER_80_264 ();
 sg13g2_decap_4 FILLER_80_275 ();
 sg13g2_decap_8 FILLER_80_283 ();
 sg13g2_decap_8 FILLER_80_290 ();
 sg13g2_fill_1 FILLER_80_297 ();
 sg13g2_decap_8 FILLER_80_302 ();
 sg13g2_decap_8 FILLER_80_309 ();
 sg13g2_decap_4 FILLER_80_316 ();
 sg13g2_fill_2 FILLER_80_320 ();
 sg13g2_fill_2 FILLER_80_326 ();
 sg13g2_fill_1 FILLER_80_328 ();
 sg13g2_decap_8 FILLER_80_333 ();
 sg13g2_fill_1 FILLER_80_340 ();
 sg13g2_decap_8 FILLER_80_345 ();
 sg13g2_decap_4 FILLER_80_352 ();
 sg13g2_fill_2 FILLER_80_356 ();
 sg13g2_decap_4 FILLER_80_362 ();
 sg13g2_fill_2 FILLER_80_366 ();
 sg13g2_decap_8 FILLER_80_376 ();
 sg13g2_fill_1 FILLER_80_383 ();
 sg13g2_decap_4 FILLER_80_388 ();
 sg13g2_decap_8 FILLER_80_396 ();
 sg13g2_decap_8 FILLER_80_403 ();
 sg13g2_decap_8 FILLER_80_410 ();
 sg13g2_decap_8 FILLER_80_417 ();
 sg13g2_decap_4 FILLER_80_424 ();
 sg13g2_fill_2 FILLER_80_428 ();
endmodule
